
module aes_comb ( clk, rst, g_input, e_input, o );
  input [1279:0] g_input;
  input [127:0] e_input;
  output [127:0] o;
  input clk, rst;
  wire   \w0[1][127] , \w0[1][126] , \w0[1][125] , \w0[1][124] , \w0[1][123] ,
         \w0[1][122] , \w0[1][121] , \w0[1][120] , \w0[1][119] , \w0[1][118] ,
         \w0[1][117] , \w0[1][116] , \w0[1][115] , \w0[1][114] , \w0[1][113] ,
         \w0[1][112] , \w0[1][111] , \w0[1][110] , \w0[1][109] , \w0[1][108] ,
         \w0[1][107] , \w0[1][106] , \w0[1][105] , \w0[1][104] , \w0[1][103] ,
         \w0[1][102] , \w0[1][101] , \w0[1][100] , \w0[1][99] , \w0[1][98] ,
         \w0[1][97] , \w0[1][96] , \w0[1][95] , \w0[1][94] , \w0[1][93] ,
         \w0[1][92] , \w0[1][91] , \w0[1][90] , \w0[1][89] , \w0[1][88] ,
         \w0[1][87] , \w0[1][86] , \w0[1][85] , \w0[1][84] , \w0[1][83] ,
         \w0[1][82] , \w0[1][81] , \w0[1][80] , \w0[1][79] , \w0[1][78] ,
         \w0[1][77] , \w0[1][76] , \w0[1][75] , \w0[1][74] , \w0[1][73] ,
         \w0[1][72] , \w0[1][71] , \w0[1][70] , \w0[1][69] , \w0[1][68] ,
         \w0[1][67] , \w0[1][66] , \w0[1][65] , \w0[1][64] , \w0[1][63] ,
         \w0[1][62] , \w0[1][61] , \w0[1][60] , \w0[1][59] , \w0[1][58] ,
         \w0[1][57] , \w0[1][56] , \w0[1][55] , \w0[1][54] , \w0[1][53] ,
         \w0[1][52] , \w0[1][51] , \w0[1][50] , \w0[1][49] , \w0[1][48] ,
         \w0[1][47] , \w0[1][46] , \w0[1][45] , \w0[1][44] , \w0[1][43] ,
         \w0[1][42] , \w0[1][41] , \w0[1][40] , \w0[1][39] , \w0[1][38] ,
         \w0[1][37] , \w0[1][36] , \w0[1][35] , \w0[1][34] , \w0[1][33] ,
         \w0[1][32] , \w0[1][31] , \w0[1][30] , \w0[1][29] , \w0[1][28] ,
         \w0[1][27] , \w0[1][26] , \w0[1][25] , \w0[1][24] , \w0[1][23] ,
         \w0[1][22] , \w0[1][21] , \w0[1][20] , \w0[1][19] , \w0[1][18] ,
         \w0[1][17] , \w0[1][16] , \w0[1][15] , \w0[1][14] , \w0[1][13] ,
         \w0[1][12] , \w0[1][11] , \w0[1][10] , \w0[1][9] , \w0[1][8] ,
         \w0[1][7] , \w0[1][6] , \w0[1][5] , \w0[1][4] , \w0[1][3] ,
         \w0[1][2] , \w0[1][1] , \w0[1][0] , \w0[9][127] , \w0[9][126] ,
         \w0[9][125] , \w0[9][124] , \w0[9][123] , \w0[9][122] , \w0[9][121] ,
         \w0[9][120] , \w0[9][119] , \w0[9][118] , \w0[9][117] , \w0[9][116] ,
         \w0[9][115] , \w0[9][114] , \w0[9][113] , \w0[9][112] , \w0[9][111] ,
         \w0[9][110] , \w0[9][109] , \w0[9][108] , \w0[9][107] , \w0[9][106] ,
         \w0[9][105] , \w0[9][104] , \w0[9][103] , \w0[9][102] , \w0[9][101] ,
         \w0[9][100] , \w0[9][99] , \w0[9][98] , \w0[9][97] , \w0[9][96] ,
         \w0[9][95] , \w0[9][94] , \w0[9][93] , \w0[9][92] , \w0[9][91] ,
         \w0[9][90] , \w0[9][89] , \w0[9][88] , \w0[9][87] , \w0[9][86] ,
         \w0[9][85] , \w0[9][84] , \w0[9][83] , \w0[9][82] , \w0[9][81] ,
         \w0[9][80] , \w0[9][79] , \w0[9][78] , \w0[9][77] , \w0[9][76] ,
         \w0[9][75] , \w0[9][74] , \w0[9][73] , \w0[9][72] , \w0[9][71] ,
         \w0[9][70] , \w0[9][69] , \w0[9][68] , \w0[9][67] , \w0[9][66] ,
         \w0[9][65] , \w0[9][64] , \w0[9][63] , \w0[9][62] , \w0[9][61] ,
         \w0[9][60] , \w0[9][59] , \w0[9][58] , \w0[9][57] , \w0[9][56] ,
         \w0[9][55] , \w0[9][54] , \w0[9][53] , \w0[9][52] , \w0[9][51] ,
         \w0[9][50] , \w0[9][49] , \w0[9][48] , \w0[9][47] , \w0[9][46] ,
         \w0[9][45] , \w0[9][44] , \w0[9][43] , \w0[9][42] , \w0[9][41] ,
         \w0[9][40] , \w0[9][39] , \w0[9][38] , \w0[9][37] , \w0[9][36] ,
         \w0[9][35] , \w0[9][34] , \w0[9][33] , \w0[9][32] , \w0[9][31] ,
         \w0[9][30] , \w0[9][29] , \w0[9][28] , \w0[9][27] , \w0[9][26] ,
         \w0[9][25] , \w0[9][24] , \w0[9][23] , \w0[9][22] , \w0[9][21] ,
         \w0[9][20] , \w0[9][19] , \w0[9][18] , \w0[9][17] , \w0[9][16] ,
         \w0[9][15] , \w0[9][14] , \w0[9][13] , \w0[9][12] , \w0[9][11] ,
         \w0[9][10] , \w0[9][9] , \w0[9][8] , \w0[9][7] , \w0[9][6] ,
         \w0[9][5] , \w0[9][4] , \w0[9][3] , \w0[9][2] , \w0[9][1] ,
         \w0[9][0] , \w0[8][127] , \w0[8][126] , \w0[8][125] , \w0[8][124] ,
         \w0[8][123] , \w0[8][122] , \w0[8][121] , \w0[8][120] , \w0[8][119] ,
         \w0[8][118] , \w0[8][117] , \w0[8][116] , \w0[8][115] , \w0[8][114] ,
         \w0[8][113] , \w0[8][112] , \w0[8][111] , \w0[8][110] , \w0[8][109] ,
         \w0[8][108] , \w0[8][107] , \w0[8][106] , \w0[8][105] , \w0[8][104] ,
         \w0[8][103] , \w0[8][102] , \w0[8][101] , \w0[8][100] , \w0[8][99] ,
         \w0[8][98] , \w0[8][97] , \w0[8][96] , \w0[8][95] , \w0[8][94] ,
         \w0[8][93] , \w0[8][92] , \w0[8][91] , \w0[8][90] , \w0[8][89] ,
         \w0[8][88] , \w0[8][87] , \w0[8][86] , \w0[8][85] , \w0[8][84] ,
         \w0[8][83] , \w0[8][82] , \w0[8][81] , \w0[8][80] , \w0[8][79] ,
         \w0[8][78] , \w0[8][77] , \w0[8][76] , \w0[8][75] , \w0[8][74] ,
         \w0[8][73] , \w0[8][72] , \w0[8][71] , \w0[8][70] , \w0[8][69] ,
         \w0[8][68] , \w0[8][67] , \w0[8][66] , \w0[8][65] , \w0[8][64] ,
         \w0[8][63] , \w0[8][62] , \w0[8][61] , \w0[8][60] , \w0[8][59] ,
         \w0[8][58] , \w0[8][57] , \w0[8][56] , \w0[8][55] , \w0[8][54] ,
         \w0[8][53] , \w0[8][52] , \w0[8][51] , \w0[8][50] , \w0[8][49] ,
         \w0[8][48] , \w0[8][47] , \w0[8][46] , \w0[8][45] , \w0[8][44] ,
         \w0[8][43] , \w0[8][42] , \w0[8][41] , \w0[8][40] , \w0[8][39] ,
         \w0[8][38] , \w0[8][37] , \w0[8][36] , \w0[8][35] , \w0[8][34] ,
         \w0[8][33] , \w0[8][32] , \w0[8][31] , \w0[8][30] , \w0[8][29] ,
         \w0[8][28] , \w0[8][27] , \w0[8][26] , \w0[8][25] , \w0[8][24] ,
         \w0[8][23] , \w0[8][22] , \w0[8][21] , \w0[8][20] , \w0[8][19] ,
         \w0[8][18] , \w0[8][17] , \w0[8][16] , \w0[8][15] , \w0[8][14] ,
         \w0[8][13] , \w0[8][12] , \w0[8][11] , \w0[8][10] , \w0[8][9] ,
         \w0[8][8] , \w0[8][7] , \w0[8][6] , \w0[8][5] , \w0[8][4] ,
         \w0[8][3] , \w0[8][2] , \w0[8][1] , \w0[8][0] , \w0[7][127] ,
         \w0[7][126] , \w0[7][125] , \w0[7][124] , \w0[7][123] , \w0[7][122] ,
         \w0[7][121] , \w0[7][120] , \w0[7][119] , \w0[7][118] , \w0[7][117] ,
         \w0[7][116] , \w0[7][115] , \w0[7][114] , \w0[7][113] , \w0[7][112] ,
         \w0[7][111] , \w0[7][110] , \w0[7][109] , \w0[7][108] , \w0[7][107] ,
         \w0[7][106] , \w0[7][105] , \w0[7][104] , \w0[7][103] , \w0[7][102] ,
         \w0[7][101] , \w0[7][100] , \w0[7][99] , \w0[7][98] , \w0[7][97] ,
         \w0[7][96] , \w0[7][95] , \w0[7][94] , \w0[7][93] , \w0[7][92] ,
         \w0[7][91] , \w0[7][90] , \w0[7][89] , \w0[7][88] , \w0[7][87] ,
         \w0[7][86] , \w0[7][85] , \w0[7][84] , \w0[7][83] , \w0[7][82] ,
         \w0[7][81] , \w0[7][80] , \w0[7][79] , \w0[7][78] , \w0[7][77] ,
         \w0[7][76] , \w0[7][75] , \w0[7][74] , \w0[7][73] , \w0[7][72] ,
         \w0[7][71] , \w0[7][70] , \w0[7][69] , \w0[7][68] , \w0[7][67] ,
         \w0[7][66] , \w0[7][65] , \w0[7][64] , \w0[7][63] , \w0[7][62] ,
         \w0[7][61] , \w0[7][60] , \w0[7][59] , \w0[7][58] , \w0[7][57] ,
         \w0[7][56] , \w0[7][55] , \w0[7][54] , \w0[7][53] , \w0[7][52] ,
         \w0[7][51] , \w0[7][50] , \w0[7][49] , \w0[7][48] , \w0[7][47] ,
         \w0[7][46] , \w0[7][45] , \w0[7][44] , \w0[7][43] , \w0[7][42] ,
         \w0[7][41] , \w0[7][40] , \w0[7][39] , \w0[7][38] , \w0[7][37] ,
         \w0[7][36] , \w0[7][35] , \w0[7][34] , \w0[7][33] , \w0[7][32] ,
         \w0[7][31] , \w0[7][30] , \w0[7][29] , \w0[7][28] , \w0[7][27] ,
         \w0[7][26] , \w0[7][25] , \w0[7][24] , \w0[7][23] , \w0[7][22] ,
         \w0[7][21] , \w0[7][20] , \w0[7][19] , \w0[7][18] , \w0[7][17] ,
         \w0[7][16] , \w0[7][15] , \w0[7][14] , \w0[7][13] , \w0[7][12] ,
         \w0[7][11] , \w0[7][10] , \w0[7][9] , \w0[7][8] , \w0[7][7] ,
         \w0[7][6] , \w0[7][5] , \w0[7][4] , \w0[7][3] , \w0[7][2] ,
         \w0[7][1] , \w0[7][0] , \w0[6][127] , \w0[6][126] , \w0[6][125] ,
         \w0[6][124] , \w0[6][123] , \w0[6][122] , \w0[6][121] , \w0[6][120] ,
         \w0[6][119] , \w0[6][118] , \w0[6][117] , \w0[6][116] , \w0[6][115] ,
         \w0[6][114] , \w0[6][113] , \w0[6][112] , \w0[6][111] , \w0[6][110] ,
         \w0[6][109] , \w0[6][108] , \w0[6][107] , \w0[6][106] , \w0[6][105] ,
         \w0[6][104] , \w0[6][103] , \w0[6][102] , \w0[6][101] , \w0[6][100] ,
         \w0[6][99] , \w0[6][98] , \w0[6][97] , \w0[6][96] , \w0[6][95] ,
         \w0[6][94] , \w0[6][93] , \w0[6][92] , \w0[6][91] , \w0[6][90] ,
         \w0[6][89] , \w0[6][88] , \w0[6][87] , \w0[6][86] , \w0[6][85] ,
         \w0[6][84] , \w0[6][83] , \w0[6][82] , \w0[6][81] , \w0[6][80] ,
         \w0[6][79] , \w0[6][78] , \w0[6][77] , \w0[6][76] , \w0[6][75] ,
         \w0[6][74] , \w0[6][73] , \w0[6][72] , \w0[6][71] , \w0[6][70] ,
         \w0[6][69] , \w0[6][68] , \w0[6][67] , \w0[6][66] , \w0[6][65] ,
         \w0[6][64] , \w0[6][63] , \w0[6][62] , \w0[6][61] , \w0[6][60] ,
         \w0[6][59] , \w0[6][58] , \w0[6][57] , \w0[6][56] , \w0[6][55] ,
         \w0[6][54] , \w0[6][53] , \w0[6][52] , \w0[6][51] , \w0[6][50] ,
         \w0[6][49] , \w0[6][48] , \w0[6][47] , \w0[6][46] , \w0[6][45] ,
         \w0[6][44] , \w0[6][43] , \w0[6][42] , \w0[6][41] , \w0[6][40] ,
         \w0[6][39] , \w0[6][38] , \w0[6][37] , \w0[6][36] , \w0[6][35] ,
         \w0[6][34] , \w0[6][33] , \w0[6][32] , \w0[6][31] , \w0[6][30] ,
         \w0[6][29] , \w0[6][28] , \w0[6][27] , \w0[6][26] , \w0[6][25] ,
         \w0[6][24] , \w0[6][23] , \w0[6][22] , \w0[6][21] , \w0[6][20] ,
         \w0[6][19] , \w0[6][18] , \w0[6][17] , \w0[6][16] , \w0[6][15] ,
         \w0[6][14] , \w0[6][13] , \w0[6][12] , \w0[6][11] , \w0[6][10] ,
         \w0[6][9] , \w0[6][8] , \w0[6][7] , \w0[6][6] , \w0[6][5] ,
         \w0[6][4] , \w0[6][3] , \w0[6][2] , \w0[6][1] , \w0[6][0] ,
         \w0[5][127] , \w0[5][126] , \w0[5][125] , \w0[5][124] , \w0[5][123] ,
         \w0[5][122] , \w0[5][121] , \w0[5][120] , \w0[5][119] , \w0[5][118] ,
         \w0[5][117] , \w0[5][116] , \w0[5][115] , \w0[5][114] , \w0[5][113] ,
         \w0[5][112] , \w0[5][111] , \w0[5][110] , \w0[5][109] , \w0[5][108] ,
         \w0[5][107] , \w0[5][106] , \w0[5][105] , \w0[5][104] , \w0[5][103] ,
         \w0[5][102] , \w0[5][101] , \w0[5][100] , \w0[5][99] , \w0[5][98] ,
         \w0[5][97] , \w0[5][96] , \w0[5][95] , \w0[5][94] , \w0[5][93] ,
         \w0[5][92] , \w0[5][91] , \w0[5][90] , \w0[5][89] , \w0[5][88] ,
         \w0[5][87] , \w0[5][86] , \w0[5][85] , \w0[5][84] , \w0[5][83] ,
         \w0[5][82] , \w0[5][81] , \w0[5][80] , \w0[5][79] , \w0[5][78] ,
         \w0[5][77] , \w0[5][76] , \w0[5][75] , \w0[5][74] , \w0[5][73] ,
         \w0[5][72] , \w0[5][71] , \w0[5][70] , \w0[5][69] , \w0[5][68] ,
         \w0[5][67] , \w0[5][66] , \w0[5][65] , \w0[5][64] , \w0[5][63] ,
         \w0[5][62] , \w0[5][61] , \w0[5][60] , \w0[5][59] , \w0[5][58] ,
         \w0[5][57] , \w0[5][56] , \w0[5][55] , \w0[5][54] , \w0[5][53] ,
         \w0[5][52] , \w0[5][51] , \w0[5][50] , \w0[5][49] , \w0[5][48] ,
         \w0[5][47] , \w0[5][46] , \w0[5][45] , \w0[5][44] , \w0[5][43] ,
         \w0[5][42] , \w0[5][41] , \w0[5][40] , \w0[5][39] , \w0[5][38] ,
         \w0[5][37] , \w0[5][36] , \w0[5][35] , \w0[5][34] , \w0[5][33] ,
         \w0[5][32] , \w0[5][31] , \w0[5][30] , \w0[5][29] , \w0[5][28] ,
         \w0[5][27] , \w0[5][26] , \w0[5][25] , \w0[5][24] , \w0[5][23] ,
         \w0[5][22] , \w0[5][21] , \w0[5][20] , \w0[5][19] , \w0[5][18] ,
         \w0[5][17] , \w0[5][16] , \w0[5][15] , \w0[5][14] , \w0[5][13] ,
         \w0[5][12] , \w0[5][11] , \w0[5][10] , \w0[5][9] , \w0[5][8] ,
         \w0[5][7] , \w0[5][6] , \w0[5][5] , \w0[5][4] , \w0[5][3] ,
         \w0[5][2] , \w0[5][1] , \w0[5][0] , \w0[4][127] , \w0[4][126] ,
         \w0[4][125] , \w0[4][124] , \w0[4][123] , \w0[4][122] , \w0[4][121] ,
         \w0[4][120] , \w0[4][119] , \w0[4][118] , \w0[4][117] , \w0[4][116] ,
         \w0[4][115] , \w0[4][114] , \w0[4][113] , \w0[4][112] , \w0[4][111] ,
         \w0[4][110] , \w0[4][109] , \w0[4][108] , \w0[4][107] , \w0[4][106] ,
         \w0[4][105] , \w0[4][104] , \w0[4][103] , \w0[4][102] , \w0[4][101] ,
         \w0[4][100] , \w0[4][99] , \w0[4][98] , \w0[4][97] , \w0[4][96] ,
         \w0[4][95] , \w0[4][94] , \w0[4][93] , \w0[4][92] , \w0[4][91] ,
         \w0[4][90] , \w0[4][89] , \w0[4][88] , \w0[4][87] , \w0[4][86] ,
         \w0[4][85] , \w0[4][84] , \w0[4][83] , \w0[4][82] , \w0[4][81] ,
         \w0[4][80] , \w0[4][79] , \w0[4][78] , \w0[4][77] , \w0[4][76] ,
         \w0[4][75] , \w0[4][74] , \w0[4][73] , \w0[4][72] , \w0[4][71] ,
         \w0[4][70] , \w0[4][69] , \w0[4][68] , \w0[4][67] , \w0[4][66] ,
         \w0[4][65] , \w0[4][64] , \w0[4][63] , \w0[4][62] , \w0[4][61] ,
         \w0[4][60] , \w0[4][59] , \w0[4][58] , \w0[4][57] , \w0[4][56] ,
         \w0[4][55] , \w0[4][54] , \w0[4][53] , \w0[4][52] , \w0[4][51] ,
         \w0[4][50] , \w0[4][49] , \w0[4][48] , \w0[4][47] , \w0[4][46] ,
         \w0[4][45] , \w0[4][44] , \w0[4][43] , \w0[4][42] , \w0[4][41] ,
         \w0[4][40] , \w0[4][39] , \w0[4][38] , \w0[4][37] , \w0[4][36] ,
         \w0[4][35] , \w0[4][34] , \w0[4][33] , \w0[4][32] , \w0[4][31] ,
         \w0[4][30] , \w0[4][29] , \w0[4][28] , \w0[4][27] , \w0[4][26] ,
         \w0[4][25] , \w0[4][24] , \w0[4][23] , \w0[4][22] , \w0[4][21] ,
         \w0[4][20] , \w0[4][19] , \w0[4][18] , \w0[4][17] , \w0[4][16] ,
         \w0[4][15] , \w0[4][14] , \w0[4][13] , \w0[4][12] , \w0[4][11] ,
         \w0[4][10] , \w0[4][9] , \w0[4][8] , \w0[4][7] , \w0[4][6] ,
         \w0[4][5] , \w0[4][4] , \w0[4][3] , \w0[4][2] , \w0[4][1] ,
         \w0[4][0] , \w0[3][127] , \w0[3][126] , \w0[3][125] , \w0[3][124] ,
         \w0[3][123] , \w0[3][122] , \w0[3][121] , \w0[3][120] , \w0[3][119] ,
         \w0[3][118] , \w0[3][117] , \w0[3][116] , \w0[3][115] , \w0[3][114] ,
         \w0[3][113] , \w0[3][112] , \w0[3][111] , \w0[3][110] , \w0[3][109] ,
         \w0[3][108] , \w0[3][107] , \w0[3][106] , \w0[3][105] , \w0[3][104] ,
         \w0[3][103] , \w0[3][102] , \w0[3][101] , \w0[3][100] , \w0[3][99] ,
         \w0[3][98] , \w0[3][97] , \w0[3][96] , \w0[3][95] , \w0[3][94] ,
         \w0[3][93] , \w0[3][92] , \w0[3][91] , \w0[3][90] , \w0[3][89] ,
         \w0[3][88] , \w0[3][87] , \w0[3][86] , \w0[3][85] , \w0[3][84] ,
         \w0[3][83] , \w0[3][82] , \w0[3][81] , \w0[3][80] , \w0[3][79] ,
         \w0[3][78] , \w0[3][77] , \w0[3][76] , \w0[3][75] , \w0[3][74] ,
         \w0[3][73] , \w0[3][72] , \w0[3][71] , \w0[3][70] , \w0[3][69] ,
         \w0[3][68] , \w0[3][67] , \w0[3][66] , \w0[3][65] , \w0[3][64] ,
         \w0[3][63] , \w0[3][62] , \w0[3][61] , \w0[3][60] , \w0[3][59] ,
         \w0[3][58] , \w0[3][57] , \w0[3][56] , \w0[3][55] , \w0[3][54] ,
         \w0[3][53] , \w0[3][52] , \w0[3][51] , \w0[3][50] , \w0[3][49] ,
         \w0[3][48] , \w0[3][47] , \w0[3][46] , \w0[3][45] , \w0[3][44] ,
         \w0[3][43] , \w0[3][42] , \w0[3][41] , \w0[3][40] , \w0[3][39] ,
         \w0[3][38] , \w0[3][37] , \w0[3][36] , \w0[3][35] , \w0[3][34] ,
         \w0[3][33] , \w0[3][32] , \w0[3][31] , \w0[3][30] , \w0[3][29] ,
         \w0[3][28] , \w0[3][27] , \w0[3][26] , \w0[3][25] , \w0[3][24] ,
         \w0[3][23] , \w0[3][22] , \w0[3][21] , \w0[3][20] , \w0[3][19] ,
         \w0[3][18] , \w0[3][17] , \w0[3][16] , \w0[3][15] , \w0[3][14] ,
         \w0[3][13] , \w0[3][12] , \w0[3][11] , \w0[3][10] , \w0[3][9] ,
         \w0[3][8] , \w0[3][7] , \w0[3][6] , \w0[3][5] , \w0[3][4] ,
         \w0[3][3] , \w0[3][2] , \w0[3][1] , \w0[3][0] , \w0[2][127] ,
         \w0[2][126] , \w0[2][125] , \w0[2][124] , \w0[2][123] , \w0[2][122] ,
         \w0[2][121] , \w0[2][120] , \w0[2][119] , \w0[2][118] , \w0[2][117] ,
         \w0[2][116] , \w0[2][115] , \w0[2][114] , \w0[2][113] , \w0[2][112] ,
         \w0[2][111] , \w0[2][110] , \w0[2][109] , \w0[2][108] , \w0[2][107] ,
         \w0[2][106] , \w0[2][105] , \w0[2][104] , \w0[2][103] , \w0[2][102] ,
         \w0[2][101] , \w0[2][100] , \w0[2][99] , \w0[2][98] , \w0[2][97] ,
         \w0[2][96] , \w0[2][95] , \w0[2][94] , \w0[2][93] , \w0[2][92] ,
         \w0[2][91] , \w0[2][90] , \w0[2][89] , \w0[2][88] , \w0[2][87] ,
         \w0[2][86] , \w0[2][85] , \w0[2][84] , \w0[2][83] , \w0[2][82] ,
         \w0[2][81] , \w0[2][80] , \w0[2][79] , \w0[2][78] , \w0[2][77] ,
         \w0[2][76] , \w0[2][75] , \w0[2][74] , \w0[2][73] , \w0[2][72] ,
         \w0[2][71] , \w0[2][70] , \w0[2][69] , \w0[2][68] , \w0[2][67] ,
         \w0[2][66] , \w0[2][65] , \w0[2][64] , \w0[2][63] , \w0[2][62] ,
         \w0[2][61] , \w0[2][60] , \w0[2][59] , \w0[2][58] , \w0[2][57] ,
         \w0[2][56] , \w0[2][55] , \w0[2][54] , \w0[2][53] , \w0[2][52] ,
         \w0[2][51] , \w0[2][50] , \w0[2][49] , \w0[2][48] , \w0[2][47] ,
         \w0[2][46] , \w0[2][45] , \w0[2][44] , \w0[2][43] , \w0[2][42] ,
         \w0[2][41] , \w0[2][40] , \w0[2][39] , \w0[2][38] , \w0[2][37] ,
         \w0[2][36] , \w0[2][35] , \w0[2][34] , \w0[2][33] , \w0[2][32] ,
         \w0[2][31] , \w0[2][30] , \w0[2][29] , \w0[2][28] , \w0[2][27] ,
         \w0[2][26] , \w0[2][25] , \w0[2][24] , \w0[2][23] , \w0[2][22] ,
         \w0[2][21] , \w0[2][20] , \w0[2][19] , \w0[2][18] , \w0[2][17] ,
         \w0[2][16] , \w0[2][15] , \w0[2][14] , \w0[2][13] , \w0[2][12] ,
         \w0[2][11] , \w0[2][10] , \w0[2][9] , \w0[2][8] , \w0[2][7] ,
         \w0[2][6] , \w0[2][5] , \w0[2][4] , \w0[2][3] , \w0[2][2] ,
         \w0[2][1] , \w0[2][0] , \w1[9][127] , \w1[9][126] , \w1[9][125] ,
         \w1[9][124] , \w1[9][123] , \w1[9][122] , \w1[9][121] , \w1[9][120] ,
         \w1[9][119] , \w1[9][118] , \w1[9][117] , \w1[9][116] , \w1[9][115] ,
         \w1[9][114] , \w1[9][113] , \w1[9][112] , \w1[9][111] , \w1[9][110] ,
         \w1[9][109] , \w1[9][108] , \w1[9][107] , \w1[9][106] , \w1[9][105] ,
         \w1[9][104] , \w1[9][103] , \w1[9][102] , \w1[9][101] , \w1[9][100] ,
         \w1[9][99] , \w1[9][98] , \w1[9][97] , \w1[9][96] , \w1[9][95] ,
         \w1[9][94] , \w1[9][93] , \w1[9][92] , \w1[9][91] , \w1[9][90] ,
         \w1[9][89] , \w1[9][88] , \w1[9][87] , \w1[9][86] , \w1[9][85] ,
         \w1[9][84] , \w1[9][83] , \w1[9][82] , \w1[9][81] , \w1[9][80] ,
         \w1[9][79] , \w1[9][78] , \w1[9][77] , \w1[9][76] , \w1[9][75] ,
         \w1[9][74] , \w1[9][73] , \w1[9][72] , \w1[9][71] , \w1[9][70] ,
         \w1[9][69] , \w1[9][68] , \w1[9][67] , \w1[9][66] , \w1[9][65] ,
         \w1[9][64] , \w1[9][63] , \w1[9][62] , \w1[9][61] , \w1[9][60] ,
         \w1[9][59] , \w1[9][58] , \w1[9][57] , \w1[9][56] , \w1[9][55] ,
         \w1[9][54] , \w1[9][53] , \w1[9][52] , \w1[9][51] , \w1[9][50] ,
         \w1[9][49] , \w1[9][48] , \w1[9][47] , \w1[9][46] , \w1[9][45] ,
         \w1[9][44] , \w1[9][43] , \w1[9][42] , \w1[9][41] , \w1[9][40] ,
         \w1[9][39] , \w1[9][38] , \w1[9][37] , \w1[9][36] , \w1[9][35] ,
         \w1[9][34] , \w1[9][33] , \w1[9][32] , \w1[9][31] , \w1[9][30] ,
         \w1[9][29] , \w1[9][28] , \w1[9][27] , \w1[9][26] , \w1[9][25] ,
         \w1[9][24] , \w1[9][23] , \w1[9][22] , \w1[9][21] , \w1[9][20] ,
         \w1[9][19] , \w1[9][18] , \w1[9][17] , \w1[9][16] , \w1[9][15] ,
         \w1[9][14] , \w1[9][13] , \w1[9][12] , \w1[9][11] , \w1[9][10] ,
         \w1[9][9] , \w1[9][8] , \w1[9][7] , \w1[9][6] , \w1[9][5] ,
         \w1[9][4] , \w1[9][3] , \w1[9][2] , \w1[9][1] , \w1[9][0] ,
         \w1[8][127] , \w1[8][126] , \w1[8][125] , \w1[8][124] , \w1[8][123] ,
         \w1[8][122] , \w1[8][121] , \w1[8][120] , \w1[8][119] , \w1[8][118] ,
         \w1[8][117] , \w1[8][116] , \w1[8][115] , \w1[8][114] , \w1[8][113] ,
         \w1[8][112] , \w1[8][111] , \w1[8][110] , \w1[8][109] , \w1[8][108] ,
         \w1[8][107] , \w1[8][106] , \w1[8][105] , \w1[8][104] , \w1[8][103] ,
         \w1[8][102] , \w1[8][101] , \w1[8][100] , \w1[8][99] , \w1[8][98] ,
         \w1[8][97] , \w1[8][96] , \w1[8][95] , \w1[8][94] , \w1[8][93] ,
         \w1[8][92] , \w1[8][91] , \w1[8][90] , \w1[8][89] , \w1[8][88] ,
         \w1[8][87] , \w1[8][86] , \w1[8][85] , \w1[8][84] , \w1[8][83] ,
         \w1[8][82] , \w1[8][81] , \w1[8][80] , \w1[8][79] , \w1[8][78] ,
         \w1[8][77] , \w1[8][76] , \w1[8][75] , \w1[8][74] , \w1[8][73] ,
         \w1[8][72] , \w1[8][71] , \w1[8][70] , \w1[8][69] , \w1[8][68] ,
         \w1[8][67] , \w1[8][66] , \w1[8][65] , \w1[8][64] , \w1[8][63] ,
         \w1[8][62] , \w1[8][61] , \w1[8][60] , \w1[8][59] , \w1[8][58] ,
         \w1[8][57] , \w1[8][56] , \w1[8][55] , \w1[8][54] , \w1[8][53] ,
         \w1[8][52] , \w1[8][51] , \w1[8][50] , \w1[8][49] , \w1[8][48] ,
         \w1[8][47] , \w1[8][46] , \w1[8][45] , \w1[8][44] , \w1[8][43] ,
         \w1[8][42] , \w1[8][41] , \w1[8][40] , \w1[8][39] , \w1[8][38] ,
         \w1[8][37] , \w1[8][36] , \w1[8][35] , \w1[8][34] , \w1[8][33] ,
         \w1[8][32] , \w1[8][31] , \w1[8][30] , \w1[8][29] , \w1[8][28] ,
         \w1[8][27] , \w1[8][26] , \w1[8][25] , \w1[8][24] , \w1[8][23] ,
         \w1[8][22] , \w1[8][21] , \w1[8][20] , \w1[8][19] , \w1[8][18] ,
         \w1[8][17] , \w1[8][16] , \w1[8][15] , \w1[8][14] , \w1[8][13] ,
         \w1[8][12] , \w1[8][11] , \w1[8][10] , \w1[8][9] , \w1[8][8] ,
         \w1[8][7] , \w1[8][6] , \w1[8][5] , \w1[8][4] , \w1[8][3] ,
         \w1[8][2] , \w1[8][1] , \w1[8][0] , \w1[7][127] , \w1[7][126] ,
         \w1[7][125] , \w1[7][124] , \w1[7][123] , \w1[7][122] , \w1[7][121] ,
         \w1[7][120] , \w1[7][119] , \w1[7][118] , \w1[7][117] , \w1[7][116] ,
         \w1[7][115] , \w1[7][114] , \w1[7][113] , \w1[7][112] , \w1[7][111] ,
         \w1[7][110] , \w1[7][109] , \w1[7][108] , \w1[7][107] , \w1[7][106] ,
         \w1[7][105] , \w1[7][104] , \w1[7][103] , \w1[7][102] , \w1[7][101] ,
         \w1[7][100] , \w1[7][99] , \w1[7][98] , \w1[7][97] , \w1[7][96] ,
         \w1[7][95] , \w1[7][94] , \w1[7][93] , \w1[7][92] , \w1[7][91] ,
         \w1[7][90] , \w1[7][89] , \w1[7][88] , \w1[7][87] , \w1[7][86] ,
         \w1[7][85] , \w1[7][84] , \w1[7][83] , \w1[7][82] , \w1[7][81] ,
         \w1[7][80] , \w1[7][79] , \w1[7][78] , \w1[7][77] , \w1[7][76] ,
         \w1[7][75] , \w1[7][74] , \w1[7][73] , \w1[7][72] , \w1[7][71] ,
         \w1[7][70] , \w1[7][69] , \w1[7][68] , \w1[7][67] , \w1[7][66] ,
         \w1[7][65] , \w1[7][64] , \w1[7][63] , \w1[7][62] , \w1[7][61] ,
         \w1[7][60] , \w1[7][59] , \w1[7][58] , \w1[7][57] , \w1[7][56] ,
         \w1[7][55] , \w1[7][54] , \w1[7][53] , \w1[7][52] , \w1[7][51] ,
         \w1[7][50] , \w1[7][49] , \w1[7][48] , \w1[7][47] , \w1[7][46] ,
         \w1[7][45] , \w1[7][44] , \w1[7][43] , \w1[7][42] , \w1[7][41] ,
         \w1[7][40] , \w1[7][39] , \w1[7][38] , \w1[7][37] , \w1[7][36] ,
         \w1[7][35] , \w1[7][34] , \w1[7][33] , \w1[7][32] , \w1[7][31] ,
         \w1[7][30] , \w1[7][29] , \w1[7][28] , \w1[7][27] , \w1[7][26] ,
         \w1[7][25] , \w1[7][24] , \w1[7][23] , \w1[7][22] , \w1[7][21] ,
         \w1[7][20] , \w1[7][19] , \w1[7][18] , \w1[7][17] , \w1[7][16] ,
         \w1[7][15] , \w1[7][14] , \w1[7][13] , \w1[7][12] , \w1[7][11] ,
         \w1[7][10] , \w1[7][9] , \w1[7][8] , \w1[7][7] , \w1[7][6] ,
         \w1[7][5] , \w1[7][4] , \w1[7][3] , \w1[7][2] , \w1[7][1] ,
         \w1[7][0] , \w1[6][127] , \w1[6][126] , \w1[6][125] , \w1[6][124] ,
         \w1[6][123] , \w1[6][122] , \w1[6][121] , \w1[6][120] , \w1[6][119] ,
         \w1[6][118] , \w1[6][117] , \w1[6][116] , \w1[6][115] , \w1[6][114] ,
         \w1[6][113] , \w1[6][112] , \w1[6][111] , \w1[6][110] , \w1[6][109] ,
         \w1[6][108] , \w1[6][107] , \w1[6][106] , \w1[6][105] , \w1[6][104] ,
         \w1[6][103] , \w1[6][102] , \w1[6][101] , \w1[6][100] , \w1[6][99] ,
         \w1[6][98] , \w1[6][97] , \w1[6][96] , \w1[6][95] , \w1[6][94] ,
         \w1[6][93] , \w1[6][92] , \w1[6][91] , \w1[6][90] , \w1[6][89] ,
         \w1[6][88] , \w1[6][87] , \w1[6][86] , \w1[6][85] , \w1[6][84] ,
         \w1[6][83] , \w1[6][82] , \w1[6][81] , \w1[6][80] , \w1[6][79] ,
         \w1[6][78] , \w1[6][77] , \w1[6][76] , \w1[6][75] , \w1[6][74] ,
         \w1[6][73] , \w1[6][72] , \w1[6][71] , \w1[6][70] , \w1[6][69] ,
         \w1[6][68] , \w1[6][67] , \w1[6][66] , \w1[6][65] , \w1[6][64] ,
         \w1[6][63] , \w1[6][62] , \w1[6][61] , \w1[6][60] , \w1[6][59] ,
         \w1[6][58] , \w1[6][57] , \w1[6][56] , \w1[6][55] , \w1[6][54] ,
         \w1[6][53] , \w1[6][52] , \w1[6][51] , \w1[6][50] , \w1[6][49] ,
         \w1[6][48] , \w1[6][47] , \w1[6][46] , \w1[6][45] , \w1[6][44] ,
         \w1[6][43] , \w1[6][42] , \w1[6][41] , \w1[6][40] , \w1[6][39] ,
         \w1[6][38] , \w1[6][37] , \w1[6][36] , \w1[6][35] , \w1[6][34] ,
         \w1[6][33] , \w1[6][32] , \w1[6][31] , \w1[6][30] , \w1[6][29] ,
         \w1[6][28] , \w1[6][27] , \w1[6][26] , \w1[6][25] , \w1[6][24] ,
         \w1[6][23] , \w1[6][22] , \w1[6][21] , \w1[6][20] , \w1[6][19] ,
         \w1[6][18] , \w1[6][17] , \w1[6][16] , \w1[6][15] , \w1[6][14] ,
         \w1[6][13] , \w1[6][12] , \w1[6][11] , \w1[6][10] , \w1[6][9] ,
         \w1[6][8] , \w1[6][7] , \w1[6][6] , \w1[6][5] , \w1[6][4] ,
         \w1[6][3] , \w1[6][2] , \w1[6][1] , \w1[6][0] , \w1[5][127] ,
         \w1[5][126] , \w1[5][125] , \w1[5][124] , \w1[5][123] , \w1[5][122] ,
         \w1[5][121] , \w1[5][120] , \w1[5][119] , \w1[5][118] , \w1[5][117] ,
         \w1[5][116] , \w1[5][115] , \w1[5][114] , \w1[5][113] , \w1[5][112] ,
         \w1[5][111] , \w1[5][110] , \w1[5][109] , \w1[5][108] , \w1[5][107] ,
         \w1[5][106] , \w1[5][105] , \w1[5][104] , \w1[5][103] , \w1[5][102] ,
         \w1[5][101] , \w1[5][100] , \w1[5][99] , \w1[5][98] , \w1[5][97] ,
         \w1[5][96] , \w1[5][95] , \w1[5][94] , \w1[5][93] , \w1[5][92] ,
         \w1[5][91] , \w1[5][90] , \w1[5][89] , \w1[5][88] , \w1[5][87] ,
         \w1[5][86] , \w1[5][85] , \w1[5][84] , \w1[5][83] , \w1[5][82] ,
         \w1[5][81] , \w1[5][80] , \w1[5][79] , \w1[5][78] , \w1[5][77] ,
         \w1[5][76] , \w1[5][75] , \w1[5][74] , \w1[5][73] , \w1[5][72] ,
         \w1[5][71] , \w1[5][70] , \w1[5][69] , \w1[5][68] , \w1[5][67] ,
         \w1[5][66] , \w1[5][65] , \w1[5][64] , \w1[5][63] , \w1[5][62] ,
         \w1[5][61] , \w1[5][60] , \w1[5][59] , \w1[5][58] , \w1[5][57] ,
         \w1[5][56] , \w1[5][55] , \w1[5][54] , \w1[5][53] , \w1[5][52] ,
         \w1[5][51] , \w1[5][50] , \w1[5][49] , \w1[5][48] , \w1[5][47] ,
         \w1[5][46] , \w1[5][45] , \w1[5][44] , \w1[5][43] , \w1[5][42] ,
         \w1[5][41] , \w1[5][40] , \w1[5][39] , \w1[5][38] , \w1[5][37] ,
         \w1[5][36] , \w1[5][35] , \w1[5][34] , \w1[5][33] , \w1[5][32] ,
         \w1[5][31] , \w1[5][30] , \w1[5][29] , \w1[5][28] , \w1[5][27] ,
         \w1[5][26] , \w1[5][25] , \w1[5][24] , \w1[5][23] , \w1[5][22] ,
         \w1[5][21] , \w1[5][20] , \w1[5][19] , \w1[5][18] , \w1[5][17] ,
         \w1[5][16] , \w1[5][15] , \w1[5][14] , \w1[5][13] , \w1[5][12] ,
         \w1[5][11] , \w1[5][10] , \w1[5][9] , \w1[5][8] , \w1[5][7] ,
         \w1[5][6] , \w1[5][5] , \w1[5][4] , \w1[5][3] , \w1[5][2] ,
         \w1[5][1] , \w1[5][0] , \w1[4][127] , \w1[4][126] , \w1[4][125] ,
         \w1[4][124] , \w1[4][123] , \w1[4][122] , \w1[4][121] , \w1[4][120] ,
         \w1[4][119] , \w1[4][118] , \w1[4][117] , \w1[4][116] , \w1[4][115] ,
         \w1[4][114] , \w1[4][113] , \w1[4][112] , \w1[4][111] , \w1[4][110] ,
         \w1[4][109] , \w1[4][108] , \w1[4][107] , \w1[4][106] , \w1[4][105] ,
         \w1[4][104] , \w1[4][103] , \w1[4][102] , \w1[4][101] , \w1[4][100] ,
         \w1[4][99] , \w1[4][98] , \w1[4][97] , \w1[4][96] , \w1[4][95] ,
         \w1[4][94] , \w1[4][93] , \w1[4][92] , \w1[4][91] , \w1[4][90] ,
         \w1[4][89] , \w1[4][88] , \w1[4][87] , \w1[4][86] , \w1[4][85] ,
         \w1[4][84] , \w1[4][83] , \w1[4][82] , \w1[4][81] , \w1[4][80] ,
         \w1[4][79] , \w1[4][78] , \w1[4][77] , \w1[4][76] , \w1[4][75] ,
         \w1[4][74] , \w1[4][73] , \w1[4][72] , \w1[4][71] , \w1[4][70] ,
         \w1[4][69] , \w1[4][68] , \w1[4][67] , \w1[4][66] , \w1[4][65] ,
         \w1[4][64] , \w1[4][63] , \w1[4][62] , \w1[4][61] , \w1[4][60] ,
         \w1[4][59] , \w1[4][58] , \w1[4][57] , \w1[4][56] , \w1[4][55] ,
         \w1[4][54] , \w1[4][53] , \w1[4][52] , \w1[4][51] , \w1[4][50] ,
         \w1[4][49] , \w1[4][48] , \w1[4][47] , \w1[4][46] , \w1[4][45] ,
         \w1[4][44] , \w1[4][43] , \w1[4][42] , \w1[4][41] , \w1[4][40] ,
         \w1[4][39] , \w1[4][38] , \w1[4][37] , \w1[4][36] , \w1[4][35] ,
         \w1[4][34] , \w1[4][33] , \w1[4][32] , \w1[4][31] , \w1[4][30] ,
         \w1[4][29] , \w1[4][28] , \w1[4][27] , \w1[4][26] , \w1[4][25] ,
         \w1[4][24] , \w1[4][23] , \w1[4][22] , \w1[4][21] , \w1[4][20] ,
         \w1[4][19] , \w1[4][18] , \w1[4][17] , \w1[4][16] , \w1[4][15] ,
         \w1[4][14] , \w1[4][13] , \w1[4][12] , \w1[4][11] , \w1[4][10] ,
         \w1[4][9] , \w1[4][8] , \w1[4][7] , \w1[4][6] , \w1[4][5] ,
         \w1[4][4] , \w1[4][3] , \w1[4][2] , \w1[4][1] , \w1[4][0] ,
         \w1[3][127] , \w1[3][126] , \w1[3][125] , \w1[3][124] , \w1[3][123] ,
         \w1[3][122] , \w1[3][121] , \w1[3][120] , \w1[3][119] , \w1[3][118] ,
         \w1[3][117] , \w1[3][116] , \w1[3][115] , \w1[3][114] , \w1[3][113] ,
         \w1[3][112] , \w1[3][111] , \w1[3][110] , \w1[3][109] , \w1[3][108] ,
         \w1[3][107] , \w1[3][106] , \w1[3][105] , \w1[3][104] , \w1[3][103] ,
         \w1[3][102] , \w1[3][101] , \w1[3][100] , \w1[3][99] , \w1[3][98] ,
         \w1[3][97] , \w1[3][96] , \w1[3][95] , \w1[3][94] , \w1[3][93] ,
         \w1[3][92] , \w1[3][91] , \w1[3][90] , \w1[3][89] , \w1[3][88] ,
         \w1[3][87] , \w1[3][86] , \w1[3][85] , \w1[3][84] , \w1[3][83] ,
         \w1[3][82] , \w1[3][81] , \w1[3][80] , \w1[3][79] , \w1[3][78] ,
         \w1[3][77] , \w1[3][76] , \w1[3][75] , \w1[3][74] , \w1[3][73] ,
         \w1[3][72] , \w1[3][71] , \w1[3][70] , \w1[3][69] , \w1[3][68] ,
         \w1[3][67] , \w1[3][66] , \w1[3][65] , \w1[3][64] , \w1[3][63] ,
         \w1[3][62] , \w1[3][61] , \w1[3][60] , \w1[3][59] , \w1[3][58] ,
         \w1[3][57] , \w1[3][56] , \w1[3][55] , \w1[3][54] , \w1[3][53] ,
         \w1[3][52] , \w1[3][51] , \w1[3][50] , \w1[3][49] , \w1[3][48] ,
         \w1[3][47] , \w1[3][46] , \w1[3][45] , \w1[3][44] , \w1[3][43] ,
         \w1[3][42] , \w1[3][41] , \w1[3][40] , \w1[3][39] , \w1[3][38] ,
         \w1[3][37] , \w1[3][36] , \w1[3][35] , \w1[3][34] , \w1[3][33] ,
         \w1[3][32] , \w1[3][31] , \w1[3][30] , \w1[3][29] , \w1[3][28] ,
         \w1[3][27] , \w1[3][26] , \w1[3][25] , \w1[3][24] , \w1[3][23] ,
         \w1[3][22] , \w1[3][21] , \w1[3][20] , \w1[3][19] , \w1[3][18] ,
         \w1[3][17] , \w1[3][16] , \w1[3][15] , \w1[3][14] , \w1[3][13] ,
         \w1[3][12] , \w1[3][11] , \w1[3][10] , \w1[3][9] , \w1[3][8] ,
         \w1[3][7] , \w1[3][6] , \w1[3][5] , \w1[3][4] , \w1[3][3] ,
         \w1[3][2] , \w1[3][1] , \w1[3][0] , \w1[2][127] , \w1[2][126] ,
         \w1[2][125] , \w1[2][124] , \w1[2][123] , \w1[2][122] , \w1[2][121] ,
         \w1[2][120] , \w1[2][119] , \w1[2][118] , \w1[2][117] , \w1[2][116] ,
         \w1[2][115] , \w1[2][114] , \w1[2][113] , \w1[2][112] , \w1[2][111] ,
         \w1[2][110] , \w1[2][109] , \w1[2][108] , \w1[2][107] , \w1[2][106] ,
         \w1[2][105] , \w1[2][104] , \w1[2][103] , \w1[2][102] , \w1[2][101] ,
         \w1[2][100] , \w1[2][99] , \w1[2][98] , \w1[2][97] , \w1[2][96] ,
         \w1[2][95] , \w1[2][94] , \w1[2][93] , \w1[2][92] , \w1[2][91] ,
         \w1[2][90] , \w1[2][89] , \w1[2][88] , \w1[2][87] , \w1[2][86] ,
         \w1[2][85] , \w1[2][84] , \w1[2][83] , \w1[2][82] , \w1[2][81] ,
         \w1[2][80] , \w1[2][79] , \w1[2][78] , \w1[2][77] , \w1[2][76] ,
         \w1[2][75] , \w1[2][74] , \w1[2][73] , \w1[2][72] , \w1[2][71] ,
         \w1[2][70] , \w1[2][69] , \w1[2][68] , \w1[2][67] , \w1[2][66] ,
         \w1[2][65] , \w1[2][64] , \w1[2][63] , \w1[2][62] , \w1[2][61] ,
         \w1[2][60] , \w1[2][59] , \w1[2][58] , \w1[2][57] , \w1[2][56] ,
         \w1[2][55] , \w1[2][54] , \w1[2][53] , \w1[2][52] , \w1[2][51] ,
         \w1[2][50] , \w1[2][49] , \w1[2][48] , \w1[2][47] , \w1[2][46] ,
         \w1[2][45] , \w1[2][44] , \w1[2][43] , \w1[2][42] , \w1[2][41] ,
         \w1[2][40] , \w1[2][39] , \w1[2][38] , \w1[2][37] , \w1[2][36] ,
         \w1[2][35] , \w1[2][34] , \w1[2][33] , \w1[2][32] , \w1[2][31] ,
         \w1[2][30] , \w1[2][29] , \w1[2][28] , \w1[2][27] , \w1[2][26] ,
         \w1[2][25] , \w1[2][24] , \w1[2][23] , \w1[2][22] , \w1[2][21] ,
         \w1[2][20] , \w1[2][19] , \w1[2][18] , \w1[2][17] , \w1[2][16] ,
         \w1[2][15] , \w1[2][14] , \w1[2][13] , \w1[2][12] , \w1[2][11] ,
         \w1[2][10] , \w1[2][9] , \w1[2][8] , \w1[2][7] , \w1[2][6] ,
         \w1[2][5] , \w1[2][4] , \w1[2][3] , \w1[2][2] , \w1[2][1] ,
         \w1[2][0] , \w1[1][127] , \w1[1][126] , \w1[1][125] , \w1[1][124] ,
         \w1[1][123] , \w1[1][122] , \w1[1][121] , \w1[1][120] , \w1[1][119] ,
         \w1[1][118] , \w1[1][117] , \w1[1][116] , \w1[1][115] , \w1[1][114] ,
         \w1[1][113] , \w1[1][112] , \w1[1][111] , \w1[1][110] , \w1[1][109] ,
         \w1[1][108] , \w1[1][107] , \w1[1][106] , \w1[1][105] , \w1[1][104] ,
         \w1[1][103] , \w1[1][102] , \w1[1][101] , \w1[1][100] , \w1[1][99] ,
         \w1[1][98] , \w1[1][97] , \w1[1][96] , \w1[1][95] , \w1[1][94] ,
         \w1[1][93] , \w1[1][92] , \w1[1][91] , \w1[1][90] , \w1[1][89] ,
         \w1[1][88] , \w1[1][87] , \w1[1][86] , \w1[1][85] , \w1[1][84] ,
         \w1[1][83] , \w1[1][82] , \w1[1][81] , \w1[1][80] , \w1[1][79] ,
         \w1[1][78] , \w1[1][77] , \w1[1][76] , \w1[1][75] , \w1[1][74] ,
         \w1[1][73] , \w1[1][72] , \w1[1][71] , \w1[1][70] , \w1[1][69] ,
         \w1[1][68] , \w1[1][67] , \w1[1][66] , \w1[1][65] , \w1[1][64] ,
         \w1[1][63] , \w1[1][62] , \w1[1][61] , \w1[1][60] , \w1[1][59] ,
         \w1[1][58] , \w1[1][57] , \w1[1][56] , \w1[1][55] , \w1[1][54] ,
         \w1[1][53] , \w1[1][52] , \w1[1][51] , \w1[1][50] , \w1[1][49] ,
         \w1[1][48] , \w1[1][47] , \w1[1][46] , \w1[1][45] , \w1[1][44] ,
         \w1[1][43] , \w1[1][42] , \w1[1][41] , \w1[1][40] , \w1[1][39] ,
         \w1[1][38] , \w1[1][37] , \w1[1][36] , \w1[1][35] , \w1[1][34] ,
         \w1[1][33] , \w1[1][32] , \w1[1][31] , \w1[1][30] , \w1[1][29] ,
         \w1[1][28] , \w1[1][27] , \w1[1][26] , \w1[1][25] , \w1[1][24] ,
         \w1[1][23] , \w1[1][22] , \w1[1][21] , \w1[1][20] , \w1[1][19] ,
         \w1[1][18] , \w1[1][17] , \w1[1][16] , \w1[1][15] , \w1[1][14] ,
         \w1[1][13] , \w1[1][12] , \w1[1][11] , \w1[1][10] , \w1[1][9] ,
         \w1[1][8] , \w1[1][7] , \w1[1][6] , \w1[1][5] , \w1[1][4] ,
         \w1[1][3] , \w1[1][2] , \w1[1][1] , \w1[1][0] , \w1[0][127] ,
         \w1[0][126] , \w1[0][125] , \w1[0][124] , \w1[0][123] , \w1[0][122] ,
         \w1[0][121] , \w1[0][120] , \w1[0][119] , \w1[0][118] , \w1[0][117] ,
         \w1[0][116] , \w1[0][115] , \w1[0][114] , \w1[0][113] , \w1[0][112] ,
         \w1[0][111] , \w1[0][110] , \w1[0][109] , \w1[0][108] , \w1[0][107] ,
         \w1[0][106] , \w1[0][105] , \w1[0][104] , \w1[0][103] , \w1[0][102] ,
         \w1[0][101] , \w1[0][100] , \w1[0][99] , \w1[0][98] , \w1[0][97] ,
         \w1[0][96] , \w1[0][95] , \w1[0][94] , \w1[0][93] , \w1[0][92] ,
         \w1[0][91] , \w1[0][90] , \w1[0][89] , \w1[0][88] , \w1[0][87] ,
         \w1[0][86] , \w1[0][85] , \w1[0][84] , \w1[0][83] , \w1[0][82] ,
         \w1[0][81] , \w1[0][80] , \w1[0][79] , \w1[0][78] , \w1[0][77] ,
         \w1[0][76] , \w1[0][75] , \w1[0][74] , \w1[0][73] , \w1[0][72] ,
         \w1[0][71] , \w1[0][70] , \w1[0][69] , \w1[0][68] , \w1[0][67] ,
         \w1[0][66] , \w1[0][65] , \w1[0][64] , \w1[0][63] , \w1[0][62] ,
         \w1[0][61] , \w1[0][60] , \w1[0][59] , \w1[0][58] , \w1[0][57] ,
         \w1[0][56] , \w1[0][55] , \w1[0][54] , \w1[0][53] , \w1[0][52] ,
         \w1[0][51] , \w1[0][50] , \w1[0][49] , \w1[0][48] , \w1[0][47] ,
         \w1[0][46] , \w1[0][45] , \w1[0][44] , \w1[0][43] , \w1[0][42] ,
         \w1[0][41] , \w1[0][40] , \w1[0][39] , \w1[0][38] , \w1[0][37] ,
         \w1[0][36] , \w1[0][35] , \w1[0][34] , \w1[0][33] , \w1[0][32] ,
         \w1[0][31] , \w1[0][30] , \w1[0][29] , \w1[0][28] , \w1[0][27] ,
         \w1[0][26] , \w1[0][25] , \w1[0][24] , \w1[0][23] , \w1[0][22] ,
         \w1[0][21] , \w1[0][20] , \w1[0][19] , \w1[0][18] , \w1[0][17] ,
         \w1[0][16] , \w1[0][15] , \w1[0][14] , \w1[0][13] , \w1[0][12] ,
         \w1[0][11] , \w1[0][10] , \w1[0][9] , \w1[0][8] , \w1[0][7] ,
         \w1[0][6] , \w1[0][5] , \w1[0][4] , \w1[0][3] , \w1[0][2] ,
         \w1[0][1] , \w1[0][0] , \w3[8][122] , \w3[8][114] , \w3[8][106] ,
         \w3[8][98] , \w3[8][90] , \w3[8][82] , \w3[8][74] , \w3[8][66] ,
         \w3[8][58] , \w3[8][50] , \w3[8][42] , \w3[8][34] , \w3[8][26] ,
         \w3[8][18] , \w3[8][10] , \w3[8][2] , \w3[7][122] , \w3[7][114] ,
         \w3[7][106] , \w3[7][98] , \w3[7][90] , \w3[7][82] , \w3[7][74] ,
         \w3[7][66] , \w3[7][58] , \w3[7][50] , \w3[7][42] , \w3[7][34] ,
         \w3[7][26] , \w3[7][18] , \w3[7][10] , \w3[7][2] , \w3[6][122] ,
         \w3[6][114] , \w3[6][106] , \w3[6][98] , \w3[6][90] , \w3[6][82] ,
         \w3[6][74] , \w3[6][66] , \w3[6][58] , \w3[6][50] , \w3[6][42] ,
         \w3[6][34] , \w3[6][26] , \w3[6][18] , \w3[6][10] , \w3[6][2] ,
         \w3[5][122] , \w3[5][114] , \w3[5][106] , \w3[5][98] , \w3[5][90] ,
         \w3[5][82] , \w3[5][74] , \w3[5][66] , \w3[5][58] , \w3[5][50] ,
         \w3[5][42] , \w3[5][34] , \w3[5][26] , \w3[5][18] , \w3[5][10] ,
         \w3[5][2] , \w3[4][122] , \w3[4][114] , \w3[4][106] , \w3[4][98] ,
         \w3[4][90] , \w3[4][82] , \w3[4][74] , \w3[4][66] , \w3[4][58] ,
         \w3[4][50] , \w3[4][42] , \w3[4][34] , \w3[4][26] , \w3[4][18] ,
         \w3[4][10] , \w3[4][2] , \w3[3][122] , \w3[3][114] , \w3[3][106] ,
         \w3[3][98] , \w3[3][90] , \w3[3][82] , \w3[3][74] , \w3[3][66] ,
         \w3[3][58] , \w3[3][50] , \w3[3][42] , \w3[3][34] , \w3[3][26] ,
         \w3[3][18] , \w3[3][10] , \w3[3][2] , \w3[2][122] , \w3[2][114] ,
         \w3[2][106] , \w3[2][98] , \w3[2][90] , \w3[2][82] , \w3[2][74] ,
         \w3[2][66] , \w3[2][58] , \w3[2][50] , \w3[2][42] , \w3[2][34] ,
         \w3[2][26] , \w3[2][18] , \w3[2][10] , \w3[2][2] , \w3[1][122] ,
         \w3[1][114] , \w3[1][106] , \w3[1][98] , \w3[1][90] , \w3[1][82] ,
         \w3[1][74] , \w3[1][66] , \w3[1][58] , \w3[1][50] , \w3[1][42] ,
         \w3[1][34] , \w3[1][26] , \w3[1][18] , \w3[1][10] , \w3[1][2] ,
         \w3[0][122] , \w3[0][114] , \w3[0][106] , \w3[0][98] , \w3[0][90] ,
         \w3[0][82] , \w3[0][74] , \w3[0][66] , \w3[0][58] , \w3[0][50] ,
         \w3[0][42] , \w3[0][34] , \w3[0][26] , \w3[0][18] , \w3[0][10] ,
         \w3[0][2] , \SUBBYTES[0].a/n1739 , \SUBBYTES[0].a/n1731 ,
         \SUBBYTES[0].a/n1723 , \SUBBYTES[0].a/n1715 , \SUBBYTES[0].a/n1707 ,
         \SUBBYTES[0].a/n1699 , \SUBBYTES[0].a/n1691 , \SUBBYTES[0].a/n1683 ,
         \SUBBYTES[0].a/n1675 , \SUBBYTES[0].a/n1667 , \SUBBYTES[0].a/n1659 ,
         \SUBBYTES[0].a/n1651 , \SUBBYTES[0].a/n1643 , \SUBBYTES[0].a/n1635 ,
         \SUBBYTES[0].a/n1627 , \SUBBYTES[0].a/n1619 , \SUBBYTES[0].a/n1616 ,
         \SUBBYTES[0].a/n1615 , \SUBBYTES[0].a/n1614 , \SUBBYTES[0].a/n1613 ,
         \SUBBYTES[0].a/n1612 , \SUBBYTES[0].a/n1611 , \SUBBYTES[0].a/n1610 ,
         \SUBBYTES[0].a/n1609 , \SUBBYTES[0].a/n1608 , \SUBBYTES[0].a/n1607 ,
         \SUBBYTES[0].a/n1606 , \SUBBYTES[0].a/n1605 , \SUBBYTES[0].a/n1604 ,
         \SUBBYTES[0].a/n1603 , \SUBBYTES[0].a/n1602 , \SUBBYTES[0].a/n1601 ,
         \SUBBYTES[0].a/n1600 , \SUBBYTES[0].a/n1599 , \SUBBYTES[0].a/n1598 ,
         \SUBBYTES[0].a/n1597 , \SUBBYTES[0].a/n1596 , \SUBBYTES[0].a/n1595 ,
         \SUBBYTES[0].a/n1594 , \SUBBYTES[0].a/n1593 , \SUBBYTES[0].a/n1592 ,
         \SUBBYTES[0].a/n1591 , \SUBBYTES[0].a/n1590 , \SUBBYTES[0].a/n1589 ,
         \SUBBYTES[0].a/n1588 , \SUBBYTES[0].a/n1587 , \SUBBYTES[0].a/n1586 ,
         \SUBBYTES[0].a/n1585 , \SUBBYTES[0].a/n1584 , \SUBBYTES[0].a/n1583 ,
         \SUBBYTES[0].a/n1582 , \SUBBYTES[0].a/n1581 , \SUBBYTES[0].a/n1580 ,
         \SUBBYTES[0].a/n1579 , \SUBBYTES[0].a/n1578 , \SUBBYTES[0].a/n1577 ,
         \SUBBYTES[0].a/n1576 , \SUBBYTES[0].a/n1575 , \SUBBYTES[0].a/n1574 ,
         \SUBBYTES[0].a/n1573 , \SUBBYTES[0].a/n1572 , \SUBBYTES[0].a/n1571 ,
         \SUBBYTES[0].a/n1570 , \SUBBYTES[0].a/n1569 , \SUBBYTES[0].a/n1568 ,
         \SUBBYTES[0].a/n1567 , \SUBBYTES[0].a/n1566 , \SUBBYTES[0].a/n1565 ,
         \SUBBYTES[0].a/n1564 , \SUBBYTES[0].a/n1563 , \SUBBYTES[0].a/n1562 ,
         \SUBBYTES[0].a/n1561 , \SUBBYTES[0].a/n1560 , \SUBBYTES[0].a/n1559 ,
         \SUBBYTES[0].a/n1558 , \SUBBYTES[0].a/n1557 , \SUBBYTES[0].a/n1556 ,
         \SUBBYTES[0].a/n1555 , \SUBBYTES[0].a/n1554 , \SUBBYTES[0].a/n1553 ,
         \SUBBYTES[0].a/n1552 , \SUBBYTES[0].a/n1551 , \SUBBYTES[0].a/n1550 ,
         \SUBBYTES[0].a/n1549 , \SUBBYTES[0].a/n1548 , \SUBBYTES[0].a/n1547 ,
         \SUBBYTES[0].a/n1546 , \SUBBYTES[0].a/n1545 , \SUBBYTES[0].a/n1544 ,
         \SUBBYTES[0].a/n1543 , \SUBBYTES[0].a/n1542 , \SUBBYTES[0].a/n1541 ,
         \SUBBYTES[0].a/n1540 , \SUBBYTES[0].a/n1539 , \SUBBYTES[0].a/n1538 ,
         \SUBBYTES[0].a/n1537 , \SUBBYTES[0].a/n1536 , \SUBBYTES[0].a/n1535 ,
         \SUBBYTES[0].a/n1534 , \SUBBYTES[0].a/n1533 , \SUBBYTES[0].a/n1532 ,
         \SUBBYTES[0].a/n1531 , \SUBBYTES[0].a/n1530 , \SUBBYTES[0].a/n1529 ,
         \SUBBYTES[0].a/n1528 , \SUBBYTES[0].a/n1527 , \SUBBYTES[0].a/n1526 ,
         \SUBBYTES[0].a/n1525 , \SUBBYTES[0].a/n1524 , \SUBBYTES[0].a/n1523 ,
         \SUBBYTES[0].a/n1522 , \SUBBYTES[0].a/n1521 , \SUBBYTES[0].a/n1520 ,
         \SUBBYTES[0].a/n1519 , \SUBBYTES[0].a/n1518 , \SUBBYTES[0].a/n1517 ,
         \SUBBYTES[0].a/n1516 , \SUBBYTES[0].a/n1515 , \SUBBYTES[0].a/n1514 ,
         \SUBBYTES[0].a/n1513 , \SUBBYTES[0].a/n1512 , \SUBBYTES[0].a/n1511 ,
         \SUBBYTES[0].a/n1510 , \SUBBYTES[0].a/n1509 , \SUBBYTES[0].a/n1508 ,
         \SUBBYTES[0].a/n1507 , \SUBBYTES[0].a/n1506 , \SUBBYTES[0].a/n1505 ,
         \SUBBYTES[0].a/n1504 , \SUBBYTES[0].a/n1503 , \SUBBYTES[0].a/n1502 ,
         \SUBBYTES[0].a/n1501 , \SUBBYTES[0].a/n1500 , \SUBBYTES[0].a/n1499 ,
         \SUBBYTES[0].a/n1498 , \SUBBYTES[0].a/n1497 , \SUBBYTES[0].a/n1496 ,
         \SUBBYTES[0].a/n1495 , \SUBBYTES[0].a/n1494 , \SUBBYTES[0].a/n1493 ,
         \SUBBYTES[0].a/n1492 , \SUBBYTES[0].a/n1491 , \SUBBYTES[0].a/n1490 ,
         \SUBBYTES[0].a/n1489 , \SUBBYTES[0].a/n1488 , \SUBBYTES[0].a/n1487 ,
         \SUBBYTES[0].a/n1486 , \SUBBYTES[0].a/n1485 , \SUBBYTES[0].a/n1484 ,
         \SUBBYTES[0].a/n1483 , \SUBBYTES[0].a/n1482 , \SUBBYTES[0].a/n1481 ,
         \SUBBYTES[0].a/n1480 , \SUBBYTES[0].a/n1479 , \SUBBYTES[0].a/n1478 ,
         \SUBBYTES[0].a/n1477 , \SUBBYTES[0].a/n1476 , \SUBBYTES[0].a/n1475 ,
         \SUBBYTES[0].a/n1474 , \SUBBYTES[0].a/n1473 , \SUBBYTES[0].a/n1472 ,
         \SUBBYTES[0].a/n1471 , \SUBBYTES[0].a/n1470 , \SUBBYTES[0].a/n1469 ,
         \SUBBYTES[0].a/n1468 , \SUBBYTES[0].a/n1467 , \SUBBYTES[0].a/n1466 ,
         \SUBBYTES[0].a/n1465 , \SUBBYTES[0].a/n1464 , \SUBBYTES[0].a/n1463 ,
         \SUBBYTES[0].a/n1462 , \SUBBYTES[0].a/n1461 , \SUBBYTES[0].a/n1460 ,
         \SUBBYTES[0].a/n1459 , \SUBBYTES[0].a/n1458 , \SUBBYTES[0].a/n1457 ,
         \SUBBYTES[0].a/n1456 , \SUBBYTES[0].a/n1455 , \SUBBYTES[0].a/n1454 ,
         \SUBBYTES[0].a/n1453 , \SUBBYTES[0].a/n1452 , \SUBBYTES[0].a/n1451 ,
         \SUBBYTES[0].a/n1450 , \SUBBYTES[0].a/n1449 , \SUBBYTES[0].a/n1448 ,
         \SUBBYTES[0].a/n1447 , \SUBBYTES[0].a/n1446 , \SUBBYTES[0].a/n1445 ,
         \SUBBYTES[0].a/n1444 , \SUBBYTES[0].a/n1443 , \SUBBYTES[0].a/n1442 ,
         \SUBBYTES[0].a/n1441 , \SUBBYTES[0].a/n1440 , \SUBBYTES[0].a/n1439 ,
         \SUBBYTES[0].a/n1438 , \SUBBYTES[0].a/n1437 , \SUBBYTES[0].a/n1436 ,
         \SUBBYTES[0].a/n1435 , \SUBBYTES[0].a/n1434 , \SUBBYTES[0].a/n1433 ,
         \SUBBYTES[0].a/n1432 , \SUBBYTES[0].a/n1431 , \SUBBYTES[0].a/n1430 ,
         \SUBBYTES[0].a/n1429 , \SUBBYTES[0].a/n1428 , \SUBBYTES[0].a/n1427 ,
         \SUBBYTES[0].a/n1426 , \SUBBYTES[0].a/n1425 , \SUBBYTES[0].a/n1424 ,
         \SUBBYTES[0].a/n1423 , \SUBBYTES[0].a/n1422 , \SUBBYTES[0].a/n1421 ,
         \SUBBYTES[0].a/n1420 , \SUBBYTES[0].a/n1419 , \SUBBYTES[0].a/n1418 ,
         \SUBBYTES[0].a/n1417 , \SUBBYTES[0].a/n1416 , \SUBBYTES[0].a/n1415 ,
         \SUBBYTES[0].a/n1414 , \SUBBYTES[0].a/n1413 , \SUBBYTES[0].a/n1412 ,
         \SUBBYTES[0].a/n1411 , \SUBBYTES[0].a/n1410 , \SUBBYTES[0].a/n1409 ,
         \SUBBYTES[0].a/n1408 , \SUBBYTES[0].a/n1407 , \SUBBYTES[0].a/n1406 ,
         \SUBBYTES[0].a/n1405 , \SUBBYTES[0].a/n1404 , \SUBBYTES[0].a/n1403 ,
         \SUBBYTES[0].a/n1402 , \SUBBYTES[0].a/n1401 , \SUBBYTES[0].a/n1400 ,
         \SUBBYTES[0].a/n1399 , \SUBBYTES[0].a/n1398 , \SUBBYTES[0].a/n1397 ,
         \SUBBYTES[0].a/n1396 , \SUBBYTES[0].a/n1395 , \SUBBYTES[0].a/n1394 ,
         \SUBBYTES[0].a/n1393 , \SUBBYTES[0].a/n1392 , \SUBBYTES[0].a/n1391 ,
         \SUBBYTES[0].a/n1390 , \SUBBYTES[0].a/n1389 , \SUBBYTES[0].a/n1388 ,
         \SUBBYTES[0].a/n1387 , \SUBBYTES[0].a/n1386 , \SUBBYTES[0].a/n1385 ,
         \SUBBYTES[0].a/n1384 , \SUBBYTES[0].a/n1383 , \SUBBYTES[0].a/n1382 ,
         \SUBBYTES[0].a/n1381 , \SUBBYTES[0].a/n1380 , \SUBBYTES[0].a/n1379 ,
         \SUBBYTES[0].a/n1378 , \SUBBYTES[0].a/n1377 , \SUBBYTES[0].a/n1376 ,
         \SUBBYTES[0].a/n1375 , \SUBBYTES[0].a/n1374 , \SUBBYTES[0].a/n1373 ,
         \SUBBYTES[0].a/n1372 , \SUBBYTES[0].a/n1371 , \SUBBYTES[0].a/n1370 ,
         \SUBBYTES[0].a/n1369 , \SUBBYTES[0].a/n1368 , \SUBBYTES[0].a/n1367 ,
         \SUBBYTES[0].a/n1366 , \SUBBYTES[0].a/n1365 , \SUBBYTES[0].a/n1364 ,
         \SUBBYTES[0].a/n1363 , \SUBBYTES[0].a/n1362 , \SUBBYTES[0].a/n1361 ,
         \SUBBYTES[0].a/n1360 , \SUBBYTES[0].a/n1359 , \SUBBYTES[0].a/n1358 ,
         \SUBBYTES[0].a/n1357 , \SUBBYTES[0].a/n1356 , \SUBBYTES[0].a/n1355 ,
         \SUBBYTES[0].a/n1354 , \SUBBYTES[0].a/n1353 , \SUBBYTES[0].a/n1352 ,
         \SUBBYTES[0].a/n1351 , \SUBBYTES[0].a/n1350 , \SUBBYTES[0].a/n1349 ,
         \SUBBYTES[0].a/n1348 , \SUBBYTES[0].a/n1347 , \SUBBYTES[0].a/n1346 ,
         \SUBBYTES[0].a/n1345 , \SUBBYTES[0].a/n1344 , \SUBBYTES[0].a/n1343 ,
         \SUBBYTES[0].a/n1342 , \SUBBYTES[0].a/n1341 , \SUBBYTES[0].a/n1340 ,
         \SUBBYTES[0].a/n1339 , \SUBBYTES[0].a/n1338 , \SUBBYTES[0].a/n1337 ,
         \SUBBYTES[0].a/n1336 , \SUBBYTES[0].a/n1335 , \SUBBYTES[0].a/n1334 ,
         \SUBBYTES[0].a/n1333 , \SUBBYTES[0].a/n1332 , \SUBBYTES[0].a/n1331 ,
         \SUBBYTES[0].a/n1330 , \SUBBYTES[0].a/n1329 , \SUBBYTES[0].a/n1328 ,
         \SUBBYTES[0].a/n1327 , \SUBBYTES[0].a/n1326 , \SUBBYTES[0].a/n1325 ,
         \SUBBYTES[0].a/n1324 , \SUBBYTES[0].a/n1323 , \SUBBYTES[0].a/n1322 ,
         \SUBBYTES[0].a/n1321 , \SUBBYTES[0].a/n1320 , \SUBBYTES[0].a/n1319 ,
         \SUBBYTES[0].a/n1318 , \SUBBYTES[0].a/n1317 , \SUBBYTES[0].a/n1316 ,
         \SUBBYTES[0].a/n1315 , \SUBBYTES[0].a/n1314 , \SUBBYTES[0].a/n1313 ,
         \SUBBYTES[0].a/n1312 , \SUBBYTES[0].a/n1311 , \SUBBYTES[0].a/n1310 ,
         \SUBBYTES[0].a/n1309 , \SUBBYTES[0].a/n1308 , \SUBBYTES[0].a/n1307 ,
         \SUBBYTES[0].a/n1306 , \SUBBYTES[0].a/n1305 , \SUBBYTES[0].a/n1304 ,
         \SUBBYTES[0].a/n1303 , \SUBBYTES[0].a/n1302 , \SUBBYTES[0].a/n1301 ,
         \SUBBYTES[0].a/n1300 , \SUBBYTES[0].a/n1299 , \SUBBYTES[0].a/n1298 ,
         \SUBBYTES[0].a/n1297 , \SUBBYTES[0].a/n1296 , \SUBBYTES[0].a/n1295 ,
         \SUBBYTES[0].a/n1294 , \SUBBYTES[0].a/n1293 , \SUBBYTES[0].a/n1292 ,
         \SUBBYTES[0].a/n1291 , \SUBBYTES[0].a/n1290 , \SUBBYTES[0].a/n1289 ,
         \SUBBYTES[0].a/n1288 , \SUBBYTES[0].a/n1287 , \SUBBYTES[0].a/n1286 ,
         \SUBBYTES[0].a/n1285 , \SUBBYTES[0].a/n1284 , \SUBBYTES[0].a/n1283 ,
         \SUBBYTES[0].a/n1282 , \SUBBYTES[0].a/n1281 , \SUBBYTES[0].a/n1280 ,
         \SUBBYTES[0].a/n1279 , \SUBBYTES[0].a/n1278 , \SUBBYTES[0].a/n1277 ,
         \SUBBYTES[0].a/n1276 , \SUBBYTES[0].a/n1275 , \SUBBYTES[0].a/n1274 ,
         \SUBBYTES[0].a/n1273 , \SUBBYTES[0].a/n1272 , \SUBBYTES[0].a/n1271 ,
         \SUBBYTES[0].a/n1270 , \SUBBYTES[0].a/n1269 , \SUBBYTES[0].a/n1268 ,
         \SUBBYTES[0].a/n1267 , \SUBBYTES[0].a/n1266 , \SUBBYTES[0].a/n1265 ,
         \SUBBYTES[0].a/n1264 , \SUBBYTES[0].a/n1263 , \SUBBYTES[0].a/n1262 ,
         \SUBBYTES[0].a/n1261 , \SUBBYTES[0].a/n1260 , \SUBBYTES[0].a/n1259 ,
         \SUBBYTES[0].a/n1258 , \SUBBYTES[0].a/n1257 , \SUBBYTES[0].a/n1256 ,
         \SUBBYTES[0].a/n1255 , \SUBBYTES[0].a/n1254 , \SUBBYTES[0].a/n1253 ,
         \SUBBYTES[0].a/n1252 , \SUBBYTES[0].a/n1251 , \SUBBYTES[0].a/n1250 ,
         \SUBBYTES[0].a/n1249 , \SUBBYTES[0].a/n1248 , \SUBBYTES[0].a/n1247 ,
         \SUBBYTES[0].a/n1246 , \SUBBYTES[0].a/n1245 , \SUBBYTES[0].a/n1244 ,
         \SUBBYTES[0].a/n1243 , \SUBBYTES[0].a/n1242 , \SUBBYTES[0].a/n1241 ,
         \SUBBYTES[0].a/n1240 , \SUBBYTES[0].a/n1239 , \SUBBYTES[0].a/n1238 ,
         \SUBBYTES[0].a/n1237 , \SUBBYTES[0].a/n1236 , \SUBBYTES[0].a/n1235 ,
         \SUBBYTES[0].a/n1234 , \SUBBYTES[0].a/n1233 , \SUBBYTES[0].a/n1232 ,
         \SUBBYTES[0].a/n1231 , \SUBBYTES[0].a/n1230 , \SUBBYTES[0].a/n1229 ,
         \SUBBYTES[0].a/n1228 , \SUBBYTES[0].a/n1227 , \SUBBYTES[0].a/n1226 ,
         \SUBBYTES[0].a/n1225 , \SUBBYTES[0].a/n1224 , \SUBBYTES[0].a/n1223 ,
         \SUBBYTES[0].a/n1222 , \SUBBYTES[0].a/n1221 , \SUBBYTES[0].a/n1220 ,
         \SUBBYTES[0].a/n1219 , \SUBBYTES[0].a/n1218 , \SUBBYTES[0].a/n1217 ,
         \SUBBYTES[0].a/n1216 , \SUBBYTES[0].a/n1215 , \SUBBYTES[0].a/n1214 ,
         \SUBBYTES[0].a/n1213 , \SUBBYTES[0].a/n1212 , \SUBBYTES[0].a/n1211 ,
         \SUBBYTES[0].a/n1210 , \SUBBYTES[0].a/n1209 , \SUBBYTES[0].a/n1208 ,
         \SUBBYTES[0].a/n1207 , \SUBBYTES[0].a/n1206 , \SUBBYTES[0].a/n1205 ,
         \SUBBYTES[0].a/n1204 , \SUBBYTES[0].a/n1203 , \SUBBYTES[0].a/n1202 ,
         \SUBBYTES[0].a/n1201 , \SUBBYTES[0].a/n1200 , \SUBBYTES[0].a/n1199 ,
         \SUBBYTES[0].a/n1198 , \SUBBYTES[0].a/n1197 , \SUBBYTES[0].a/n1196 ,
         \SUBBYTES[0].a/n1195 , \SUBBYTES[0].a/n1194 , \SUBBYTES[0].a/n1193 ,
         \SUBBYTES[0].a/n1192 , \SUBBYTES[0].a/n1191 , \SUBBYTES[0].a/n1190 ,
         \SUBBYTES[0].a/n1189 , \SUBBYTES[0].a/n1188 , \SUBBYTES[0].a/n1187 ,
         \SUBBYTES[0].a/n1186 , \SUBBYTES[0].a/n1185 , \SUBBYTES[0].a/n1184 ,
         \SUBBYTES[0].a/n1183 , \SUBBYTES[0].a/n1182 , \SUBBYTES[0].a/n1181 ,
         \SUBBYTES[0].a/n1180 , \SUBBYTES[0].a/n1179 , \SUBBYTES[0].a/n1178 ,
         \SUBBYTES[0].a/n1177 , \SUBBYTES[0].a/n1176 , \SUBBYTES[0].a/n1175 ,
         \SUBBYTES[0].a/n1174 , \SUBBYTES[0].a/n1173 , \SUBBYTES[0].a/n1172 ,
         \SUBBYTES[0].a/n1171 , \SUBBYTES[0].a/n1170 , \SUBBYTES[0].a/n1169 ,
         \SUBBYTES[0].a/n1168 , \SUBBYTES[0].a/n1167 , \SUBBYTES[0].a/n1166 ,
         \SUBBYTES[0].a/n1165 , \SUBBYTES[0].a/n1164 , \SUBBYTES[0].a/n1163 ,
         \SUBBYTES[0].a/n1162 , \SUBBYTES[0].a/n1161 , \SUBBYTES[0].a/n1160 ,
         \SUBBYTES[0].a/n1159 , \SUBBYTES[0].a/n1158 , \SUBBYTES[0].a/n1157 ,
         \SUBBYTES[0].a/n1156 , \SUBBYTES[0].a/n1155 , \SUBBYTES[0].a/n1154 ,
         \SUBBYTES[0].a/n1153 , \SUBBYTES[0].a/n1152 , \SUBBYTES[0].a/n1151 ,
         \SUBBYTES[0].a/n1150 , \SUBBYTES[0].a/n1149 , \SUBBYTES[0].a/n1148 ,
         \SUBBYTES[0].a/n1147 , \SUBBYTES[0].a/n1146 , \SUBBYTES[0].a/n1145 ,
         \SUBBYTES[0].a/n1144 , \SUBBYTES[0].a/n1143 , \SUBBYTES[0].a/n1142 ,
         \SUBBYTES[0].a/n1141 , \SUBBYTES[0].a/n1140 , \SUBBYTES[0].a/n1139 ,
         \SUBBYTES[0].a/n1138 , \SUBBYTES[0].a/n1137 , \SUBBYTES[0].a/n1136 ,
         \SUBBYTES[0].a/n1135 , \SUBBYTES[0].a/n1134 , \SUBBYTES[0].a/n1133 ,
         \SUBBYTES[0].a/n1132 , \SUBBYTES[0].a/n1131 , \SUBBYTES[0].a/n1130 ,
         \SUBBYTES[0].a/n1129 , \SUBBYTES[0].a/n1128 , \SUBBYTES[0].a/n1127 ,
         \SUBBYTES[0].a/n1126 , \SUBBYTES[0].a/n1125 , \SUBBYTES[0].a/n1124 ,
         \SUBBYTES[0].a/n1123 , \SUBBYTES[0].a/n1122 , \SUBBYTES[0].a/n1121 ,
         \SUBBYTES[0].a/n1120 , \SUBBYTES[0].a/n1119 , \SUBBYTES[0].a/n1118 ,
         \SUBBYTES[0].a/n1117 , \SUBBYTES[0].a/n1116 , \SUBBYTES[0].a/n1115 ,
         \SUBBYTES[0].a/n1114 , \SUBBYTES[0].a/n1113 , \SUBBYTES[0].a/n1112 ,
         \SUBBYTES[0].a/n1111 , \SUBBYTES[0].a/n1110 , \SUBBYTES[0].a/n1109 ,
         \SUBBYTES[0].a/n1108 , \SUBBYTES[0].a/n1107 , \SUBBYTES[0].a/n1106 ,
         \SUBBYTES[0].a/n1105 , \SUBBYTES[0].a/n1104 , \SUBBYTES[0].a/n1103 ,
         \SUBBYTES[0].a/n1102 , \SUBBYTES[0].a/n1101 , \SUBBYTES[0].a/n1100 ,
         \SUBBYTES[0].a/n1099 , \SUBBYTES[0].a/n1098 , \SUBBYTES[0].a/n1097 ,
         \SUBBYTES[0].a/n1096 , \SUBBYTES[0].a/n1095 , \SUBBYTES[0].a/n1094 ,
         \SUBBYTES[0].a/n1093 , \SUBBYTES[0].a/n1092 , \SUBBYTES[0].a/n1091 ,
         \SUBBYTES[0].a/n1090 , \SUBBYTES[0].a/n1089 , \SUBBYTES[0].a/n1088 ,
         \SUBBYTES[0].a/n1087 , \SUBBYTES[0].a/n1086 , \SUBBYTES[0].a/n1085 ,
         \SUBBYTES[0].a/n1084 , \SUBBYTES[0].a/n1083 , \SUBBYTES[0].a/n1082 ,
         \SUBBYTES[0].a/n1081 , \SUBBYTES[0].a/n1080 , \SUBBYTES[0].a/n1079 ,
         \SUBBYTES[0].a/n1078 , \SUBBYTES[0].a/n1077 , \SUBBYTES[0].a/n1076 ,
         \SUBBYTES[0].a/n1075 , \SUBBYTES[0].a/n1074 , \SUBBYTES[0].a/n1073 ,
         \SUBBYTES[0].a/n1072 , \SUBBYTES[0].a/n1071 , \SUBBYTES[0].a/n1070 ,
         \SUBBYTES[0].a/n1069 , \SUBBYTES[0].a/n1068 , \SUBBYTES[0].a/n1067 ,
         \SUBBYTES[0].a/n1066 , \SUBBYTES[0].a/n1065 , \SUBBYTES[0].a/n1064 ,
         \SUBBYTES[0].a/n1063 , \SUBBYTES[0].a/n1062 , \SUBBYTES[0].a/n1061 ,
         \SUBBYTES[0].a/n1060 , \SUBBYTES[0].a/n1059 , \SUBBYTES[0].a/n1058 ,
         \SUBBYTES[0].a/n1057 , \SUBBYTES[0].a/n1056 , \SUBBYTES[0].a/n1055 ,
         \SUBBYTES[0].a/n1054 , \SUBBYTES[0].a/n1053 , \SUBBYTES[0].a/n1052 ,
         \SUBBYTES[0].a/n1051 , \SUBBYTES[0].a/n1050 , \SUBBYTES[0].a/n1049 ,
         \SUBBYTES[0].a/n1048 , \SUBBYTES[0].a/n1047 , \SUBBYTES[0].a/n1046 ,
         \SUBBYTES[0].a/n1045 , \SUBBYTES[0].a/n1044 , \SUBBYTES[0].a/n1043 ,
         \SUBBYTES[0].a/n1042 , \SUBBYTES[0].a/n1041 , \SUBBYTES[0].a/n1040 ,
         \SUBBYTES[0].a/n1039 , \SUBBYTES[0].a/n1038 , \SUBBYTES[0].a/n1037 ,
         \SUBBYTES[0].a/n1036 , \SUBBYTES[0].a/n1035 , \SUBBYTES[0].a/n1034 ,
         \SUBBYTES[0].a/n1033 , \SUBBYTES[0].a/n1032 , \SUBBYTES[0].a/n1031 ,
         \SUBBYTES[0].a/n1030 , \SUBBYTES[0].a/n1029 , \SUBBYTES[0].a/n1028 ,
         \SUBBYTES[0].a/n1027 , \SUBBYTES[0].a/n1026 , \SUBBYTES[0].a/n1025 ,
         \SUBBYTES[0].a/n1024 , \SUBBYTES[0].a/n1023 , \SUBBYTES[0].a/n1022 ,
         \SUBBYTES[0].a/n1021 , \SUBBYTES[0].a/n1020 , \SUBBYTES[0].a/n1019 ,
         \SUBBYTES[0].a/n1018 , \SUBBYTES[0].a/n1017 , \SUBBYTES[0].a/n1016 ,
         \SUBBYTES[0].a/n1015 , \SUBBYTES[0].a/n1014 , \SUBBYTES[0].a/n1013 ,
         \SUBBYTES[0].a/n1012 , \SUBBYTES[0].a/n1011 , \SUBBYTES[0].a/n1010 ,
         \SUBBYTES[0].a/n1009 , \SUBBYTES[0].a/n1008 , \SUBBYTES[0].a/n1007 ,
         \SUBBYTES[0].a/n1006 , \SUBBYTES[0].a/n1005 , \SUBBYTES[0].a/n1004 ,
         \SUBBYTES[0].a/n1003 , \SUBBYTES[0].a/n1002 , \SUBBYTES[0].a/n1001 ,
         \SUBBYTES[0].a/n1000 , \SUBBYTES[0].a/n999 , \SUBBYTES[0].a/n998 ,
         \SUBBYTES[0].a/n997 , \SUBBYTES[0].a/n996 , \SUBBYTES[0].a/n995 ,
         \SUBBYTES[0].a/n994 , \SUBBYTES[0].a/n993 , \SUBBYTES[0].a/n992 ,
         \SUBBYTES[0].a/n991 , \SUBBYTES[0].a/n990 , \SUBBYTES[0].a/n989 ,
         \SUBBYTES[0].a/n988 , \SUBBYTES[0].a/n987 , \SUBBYTES[0].a/n986 ,
         \SUBBYTES[0].a/n985 , \SUBBYTES[0].a/n984 , \SUBBYTES[0].a/n983 ,
         \SUBBYTES[0].a/n982 , \SUBBYTES[0].a/n981 , \SUBBYTES[0].a/n980 ,
         \SUBBYTES[0].a/n979 , \SUBBYTES[0].a/n978 , \SUBBYTES[0].a/n977 ,
         \SUBBYTES[0].a/n976 , \SUBBYTES[0].a/n975 , \SUBBYTES[0].a/n974 ,
         \SUBBYTES[0].a/n973 , \SUBBYTES[0].a/n972 , \SUBBYTES[0].a/n971 ,
         \SUBBYTES[0].a/n970 , \SUBBYTES[0].a/n969 , \SUBBYTES[0].a/n968 ,
         \SUBBYTES[0].a/n967 , \SUBBYTES[0].a/n966 , \SUBBYTES[0].a/n965 ,
         \SUBBYTES[0].a/n964 , \SUBBYTES[0].a/n963 , \SUBBYTES[0].a/n962 ,
         \SUBBYTES[0].a/n961 , \SUBBYTES[0].a/n960 , \SUBBYTES[0].a/n959 ,
         \SUBBYTES[0].a/n958 , \SUBBYTES[0].a/n957 , \SUBBYTES[0].a/n956 ,
         \SUBBYTES[0].a/n955 , \SUBBYTES[0].a/n954 , \SUBBYTES[0].a/n953 ,
         \SUBBYTES[0].a/n952 , \SUBBYTES[0].a/n951 , \SUBBYTES[0].a/n950 ,
         \SUBBYTES[0].a/n949 , \SUBBYTES[0].a/n948 , \SUBBYTES[0].a/n947 ,
         \SUBBYTES[0].a/n946 , \SUBBYTES[0].a/n945 , \SUBBYTES[0].a/n944 ,
         \SUBBYTES[0].a/n943 , \SUBBYTES[0].a/n942 , \SUBBYTES[0].a/n941 ,
         \SUBBYTES[0].a/n940 , \SUBBYTES[0].a/n939 , \SUBBYTES[0].a/n938 ,
         \SUBBYTES[0].a/n937 , \SUBBYTES[0].a/n936 , \SUBBYTES[0].a/n935 ,
         \SUBBYTES[0].a/n934 , \SUBBYTES[0].a/n933 , \SUBBYTES[0].a/n932 ,
         \SUBBYTES[0].a/n931 , \SUBBYTES[0].a/n930 , \SUBBYTES[0].a/n929 ,
         \SUBBYTES[0].a/n928 , \SUBBYTES[0].a/n927 , \SUBBYTES[0].a/n926 ,
         \SUBBYTES[0].a/n925 , \SUBBYTES[0].a/n924 , \SUBBYTES[0].a/n923 ,
         \SUBBYTES[0].a/n922 , \SUBBYTES[0].a/n921 , \SUBBYTES[0].a/n920 ,
         \SUBBYTES[0].a/n919 , \SUBBYTES[0].a/n918 , \SUBBYTES[0].a/n917 ,
         \SUBBYTES[0].a/n916 , \SUBBYTES[0].a/n915 , \SUBBYTES[0].a/n914 ,
         \SUBBYTES[0].a/n913 , \SUBBYTES[0].a/n912 , \SUBBYTES[0].a/n911 ,
         \SUBBYTES[0].a/n910 , \SUBBYTES[0].a/n909 , \SUBBYTES[0].a/n908 ,
         \SUBBYTES[0].a/n907 , \SUBBYTES[0].a/n906 , \SUBBYTES[0].a/n905 ,
         \SUBBYTES[0].a/n904 , \SUBBYTES[0].a/n903 , \SUBBYTES[0].a/n902 ,
         \SUBBYTES[0].a/n901 , \SUBBYTES[0].a/n900 , \SUBBYTES[0].a/n899 ,
         \SUBBYTES[0].a/n898 , \SUBBYTES[0].a/n897 , \SUBBYTES[0].a/n896 ,
         \SUBBYTES[0].a/n895 , \SUBBYTES[0].a/n894 , \SUBBYTES[0].a/n893 ,
         \SUBBYTES[0].a/n892 , \SUBBYTES[0].a/n891 , \SUBBYTES[0].a/n890 ,
         \SUBBYTES[0].a/n889 , \SUBBYTES[0].a/n888 , \SUBBYTES[0].a/n887 ,
         \SUBBYTES[0].a/n886 , \SUBBYTES[0].a/n885 , \SUBBYTES[0].a/n884 ,
         \SUBBYTES[0].a/n883 , \SUBBYTES[0].a/n882 , \SUBBYTES[0].a/n881 ,
         \SUBBYTES[0].a/n880 , \SUBBYTES[0].a/n879 , \SUBBYTES[0].a/n878 ,
         \SUBBYTES[0].a/n877 , \SUBBYTES[0].a/n876 , \SUBBYTES[0].a/n875 ,
         \SUBBYTES[0].a/n874 , \SUBBYTES[0].a/n873 , \SUBBYTES[0].a/n872 ,
         \SUBBYTES[0].a/n871 , \SUBBYTES[0].a/n870 , \SUBBYTES[0].a/n869 ,
         \SUBBYTES[0].a/n868 , \SUBBYTES[0].a/n867 , \SUBBYTES[0].a/n866 ,
         \SUBBYTES[0].a/n865 , \SUBBYTES[0].a/n864 , \SUBBYTES[0].a/n863 ,
         \SUBBYTES[0].a/n862 , \SUBBYTES[0].a/n861 , \SUBBYTES[0].a/n860 ,
         \SUBBYTES[0].a/n859 , \SUBBYTES[0].a/n858 , \SUBBYTES[0].a/n857 ,
         \SUBBYTES[0].a/n856 , \SUBBYTES[0].a/n855 , \SUBBYTES[0].a/n854 ,
         \SUBBYTES[0].a/n853 , \SUBBYTES[0].a/n852 , \SUBBYTES[0].a/n851 ,
         \SUBBYTES[0].a/n850 , \SUBBYTES[0].a/n849 , \SUBBYTES[0].a/n848 ,
         \SUBBYTES[0].a/n847 , \SUBBYTES[0].a/n846 , \SUBBYTES[0].a/n845 ,
         \SUBBYTES[0].a/n844 , \SUBBYTES[0].a/n843 , \SUBBYTES[0].a/n842 ,
         \SUBBYTES[0].a/n841 , \SUBBYTES[0].a/n840 , \SUBBYTES[0].a/n839 ,
         \SUBBYTES[0].a/n838 , \SUBBYTES[0].a/n837 , \SUBBYTES[0].a/n836 ,
         \SUBBYTES[0].a/n835 , \SUBBYTES[0].a/n834 , \SUBBYTES[0].a/n833 ,
         \SUBBYTES[0].a/n832 , \SUBBYTES[0].a/n831 , \SUBBYTES[0].a/n830 ,
         \SUBBYTES[0].a/n829 , \SUBBYTES[0].a/n828 , \SUBBYTES[0].a/n827 ,
         \SUBBYTES[0].a/n826 , \SUBBYTES[0].a/n825 , \SUBBYTES[0].a/n824 ,
         \SUBBYTES[0].a/n823 , \SUBBYTES[0].a/n822 , \SUBBYTES[0].a/n821 ,
         \SUBBYTES[0].a/n820 , \SUBBYTES[0].a/n819 , \SUBBYTES[0].a/n818 ,
         \SUBBYTES[0].a/n817 , \SUBBYTES[0].a/n816 , \SUBBYTES[0].a/n815 ,
         \SUBBYTES[0].a/n814 , \SUBBYTES[0].a/n813 , \SUBBYTES[0].a/n812 ,
         \SUBBYTES[0].a/n811 , \SUBBYTES[0].a/n810 , \SUBBYTES[0].a/n809 ,
         \SUBBYTES[0].a/n808 , \SUBBYTES[0].a/n807 , \SUBBYTES[0].a/n806 ,
         \SUBBYTES[0].a/n805 , \SUBBYTES[0].a/n804 , \SUBBYTES[0].a/n803 ,
         \SUBBYTES[0].a/n802 , \SUBBYTES[0].a/n801 , \SUBBYTES[0].a/n800 ,
         \SUBBYTES[0].a/n799 , \SUBBYTES[0].a/n798 , \SUBBYTES[0].a/n797 ,
         \SUBBYTES[0].a/n796 , \SUBBYTES[0].a/n795 , \SUBBYTES[0].a/n794 ,
         \SUBBYTES[0].a/n793 , \SUBBYTES[0].a/n792 , \SUBBYTES[0].a/n791 ,
         \SUBBYTES[0].a/n790 , \SUBBYTES[0].a/n789 , \SUBBYTES[0].a/n788 ,
         \SUBBYTES[0].a/n787 , \SUBBYTES[0].a/n786 , \SUBBYTES[0].a/n785 ,
         \SUBBYTES[0].a/n784 , \SUBBYTES[0].a/n783 , \SUBBYTES[0].a/n782 ,
         \SUBBYTES[0].a/n781 , \SUBBYTES[0].a/n780 , \SUBBYTES[0].a/n779 ,
         \SUBBYTES[0].a/n778 , \SUBBYTES[0].a/n777 , \SUBBYTES[0].a/n776 ,
         \SUBBYTES[0].a/n775 , \SUBBYTES[0].a/n774 , \SUBBYTES[0].a/n773 ,
         \SUBBYTES[0].a/n772 , \SUBBYTES[0].a/n771 , \SUBBYTES[0].a/n770 ,
         \SUBBYTES[0].a/n769 , \SUBBYTES[0].a/n768 , \SUBBYTES[0].a/n767 ,
         \SUBBYTES[0].a/n766 , \SUBBYTES[0].a/n765 , \SUBBYTES[0].a/n764 ,
         \SUBBYTES[0].a/n763 , \SUBBYTES[0].a/n762 , \SUBBYTES[0].a/n761 ,
         \SUBBYTES[0].a/n760 , \SUBBYTES[0].a/n759 , \SUBBYTES[0].a/n758 ,
         \SUBBYTES[0].a/n757 , \SUBBYTES[0].a/n756 , \SUBBYTES[0].a/n755 ,
         \SUBBYTES[0].a/n754 , \SUBBYTES[0].a/n753 , \SUBBYTES[0].a/n752 ,
         \SUBBYTES[0].a/n751 , \SUBBYTES[0].a/n750 , \SUBBYTES[0].a/n749 ,
         \SUBBYTES[0].a/n748 , \SUBBYTES[0].a/n747 , \SUBBYTES[0].a/n746 ,
         \SUBBYTES[0].a/n745 , \SUBBYTES[0].a/n744 , \SUBBYTES[0].a/n743 ,
         \SUBBYTES[0].a/n742 , \SUBBYTES[0].a/n741 , \SUBBYTES[0].a/n740 ,
         \SUBBYTES[0].a/n739 , \SUBBYTES[0].a/n738 , \SUBBYTES[0].a/n737 ,
         \SUBBYTES[0].a/n736 , \SUBBYTES[0].a/n735 , \SUBBYTES[0].a/n734 ,
         \SUBBYTES[0].a/n733 , \SUBBYTES[0].a/n732 , \SUBBYTES[0].a/n731 ,
         \SUBBYTES[0].a/n730 , \SUBBYTES[0].a/n729 , \SUBBYTES[0].a/n728 ,
         \SUBBYTES[0].a/n727 , \SUBBYTES[0].a/n726 , \SUBBYTES[0].a/n725 ,
         \SUBBYTES[0].a/n724 , \SUBBYTES[0].a/n723 , \SUBBYTES[0].a/n722 ,
         \SUBBYTES[0].a/n721 , \SUBBYTES[0].a/n720 , \SUBBYTES[0].a/n719 ,
         \SUBBYTES[0].a/n718 , \SUBBYTES[0].a/n717 , \SUBBYTES[0].a/n716 ,
         \SUBBYTES[0].a/n715 , \SUBBYTES[0].a/n714 , \SUBBYTES[0].a/n713 ,
         \SUBBYTES[0].a/n712 , \SUBBYTES[0].a/n711 , \SUBBYTES[0].a/n710 ,
         \SUBBYTES[0].a/n709 , \SUBBYTES[0].a/n708 , \SUBBYTES[0].a/n707 ,
         \SUBBYTES[0].a/n706 , \SUBBYTES[0].a/n705 , \SUBBYTES[0].a/n704 ,
         \SUBBYTES[0].a/n703 , \SUBBYTES[0].a/n702 , \SUBBYTES[0].a/n701 ,
         \SUBBYTES[0].a/n700 , \SUBBYTES[0].a/n699 , \SUBBYTES[0].a/n698 ,
         \SUBBYTES[0].a/n697 , \SUBBYTES[0].a/n696 , \SUBBYTES[0].a/n695 ,
         \SUBBYTES[0].a/n694 , \SUBBYTES[0].a/n693 , \SUBBYTES[0].a/n692 ,
         \SUBBYTES[0].a/n691 , \SUBBYTES[0].a/n690 , \SUBBYTES[0].a/n689 ,
         \SUBBYTES[0].a/n688 , \SUBBYTES[0].a/n687 , \SUBBYTES[0].a/n686 ,
         \SUBBYTES[0].a/n685 , \SUBBYTES[0].a/n684 , \SUBBYTES[0].a/n683 ,
         \SUBBYTES[0].a/n682 , \SUBBYTES[0].a/n681 , \SUBBYTES[0].a/n680 ,
         \SUBBYTES[0].a/n679 , \SUBBYTES[0].a/n678 , \SUBBYTES[0].a/n677 ,
         \SUBBYTES[0].a/n676 , \SUBBYTES[0].a/n675 , \SUBBYTES[0].a/n674 ,
         \SUBBYTES[0].a/n673 , \SUBBYTES[0].a/n672 , \SUBBYTES[0].a/n671 ,
         \SUBBYTES[0].a/n670 , \SUBBYTES[0].a/n669 , \SUBBYTES[0].a/n668 ,
         \SUBBYTES[0].a/n667 , \SUBBYTES[0].a/n666 , \SUBBYTES[0].a/n665 ,
         \SUBBYTES[0].a/n664 , \SUBBYTES[0].a/n663 , \SUBBYTES[0].a/n662 ,
         \SUBBYTES[0].a/n661 , \SUBBYTES[0].a/n660 , \SUBBYTES[0].a/n659 ,
         \SUBBYTES[0].a/n658 , \SUBBYTES[0].a/n657 , \SUBBYTES[0].a/n656 ,
         \SUBBYTES[0].a/n655 , \SUBBYTES[0].a/n654 , \SUBBYTES[0].a/n653 ,
         \SUBBYTES[0].a/n652 , \SUBBYTES[0].a/n651 , \SUBBYTES[0].a/n650 ,
         \SUBBYTES[0].a/n649 , \SUBBYTES[0].a/n648 , \SUBBYTES[0].a/n647 ,
         \SUBBYTES[0].a/n646 , \SUBBYTES[0].a/n645 , \SUBBYTES[0].a/n644 ,
         \SUBBYTES[0].a/n643 , \SUBBYTES[0].a/n642 , \SUBBYTES[0].a/n641 ,
         \SUBBYTES[0].a/n640 , \SUBBYTES[0].a/n639 , \SUBBYTES[0].a/n638 ,
         \SUBBYTES[0].a/n637 , \SUBBYTES[0].a/n636 , \SUBBYTES[0].a/n635 ,
         \SUBBYTES[0].a/n634 , \SUBBYTES[0].a/n633 , \SUBBYTES[0].a/n632 ,
         \SUBBYTES[0].a/n631 , \SUBBYTES[0].a/n630 , \SUBBYTES[0].a/n629 ,
         \SUBBYTES[0].a/n628 , \SUBBYTES[0].a/n627 , \SUBBYTES[0].a/n626 ,
         \SUBBYTES[0].a/n625 , \SUBBYTES[0].a/n624 , \SUBBYTES[0].a/n623 ,
         \SUBBYTES[0].a/n622 , \SUBBYTES[0].a/n621 , \SUBBYTES[0].a/n620 ,
         \SUBBYTES[0].a/n619 , \SUBBYTES[0].a/n618 , \SUBBYTES[0].a/n617 ,
         \SUBBYTES[0].a/n616 , \SUBBYTES[0].a/n615 , \SUBBYTES[0].a/n614 ,
         \SUBBYTES[0].a/n613 , \SUBBYTES[0].a/n612 , \SUBBYTES[0].a/n611 ,
         \SUBBYTES[0].a/n610 , \SUBBYTES[0].a/n609 , \SUBBYTES[0].a/n608 ,
         \SUBBYTES[0].a/n607 , \SUBBYTES[0].a/n606 , \SUBBYTES[0].a/n605 ,
         \SUBBYTES[0].a/n604 , \SUBBYTES[0].a/n603 , \SUBBYTES[0].a/n602 ,
         \SUBBYTES[0].a/n601 , \SUBBYTES[0].a/n600 , \SUBBYTES[0].a/n599 ,
         \SUBBYTES[0].a/n598 , \SUBBYTES[0].a/n597 , \SUBBYTES[0].a/n596 ,
         \SUBBYTES[0].a/n595 , \SUBBYTES[0].a/n594 , \SUBBYTES[0].a/n593 ,
         \SUBBYTES[0].a/n592 , \SUBBYTES[0].a/n591 , \SUBBYTES[0].a/n590 ,
         \SUBBYTES[0].a/n589 , \SUBBYTES[0].a/n588 , \SUBBYTES[0].a/n587 ,
         \SUBBYTES[0].a/n586 , \SUBBYTES[0].a/n585 , \SUBBYTES[0].a/n584 ,
         \SUBBYTES[0].a/n583 , \SUBBYTES[0].a/n582 , \SUBBYTES[0].a/n581 ,
         \SUBBYTES[0].a/n580 , \SUBBYTES[0].a/n579 , \SUBBYTES[0].a/n578 ,
         \SUBBYTES[0].a/n577 , \SUBBYTES[0].a/n576 , \SUBBYTES[0].a/n575 ,
         \SUBBYTES[0].a/n574 , \SUBBYTES[0].a/n573 , \SUBBYTES[0].a/n572 ,
         \SUBBYTES[0].a/n571 , \SUBBYTES[0].a/n570 , \SUBBYTES[0].a/n569 ,
         \SUBBYTES[0].a/n568 , \SUBBYTES[0].a/n567 , \SUBBYTES[0].a/n566 ,
         \SUBBYTES[0].a/n565 , \SUBBYTES[0].a/n564 , \SUBBYTES[0].a/n563 ,
         \SUBBYTES[0].a/n562 , \SUBBYTES[0].a/n561 , \SUBBYTES[0].a/n560 ,
         \SUBBYTES[0].a/n559 , \SUBBYTES[0].a/n558 , \SUBBYTES[0].a/n557 ,
         \SUBBYTES[0].a/n556 , \SUBBYTES[0].a/n555 , \SUBBYTES[0].a/n554 ,
         \SUBBYTES[0].a/n553 , \SUBBYTES[0].a/n552 , \SUBBYTES[0].a/n551 ,
         \SUBBYTES[0].a/n550 , \SUBBYTES[0].a/n549 , \SUBBYTES[0].a/n548 ,
         \SUBBYTES[0].a/n547 , \SUBBYTES[0].a/n546 , \SUBBYTES[0].a/n545 ,
         \SUBBYTES[0].a/n544 , \SUBBYTES[0].a/n543 , \SUBBYTES[0].a/n542 ,
         \SUBBYTES[0].a/n541 , \SUBBYTES[0].a/n540 , \SUBBYTES[0].a/n539 ,
         \SUBBYTES[0].a/n538 , \SUBBYTES[0].a/n537 , \SUBBYTES[0].a/n536 ,
         \SUBBYTES[0].a/n535 , \SUBBYTES[0].a/n534 , \SUBBYTES[0].a/n533 ,
         \SUBBYTES[0].a/n532 , \SUBBYTES[0].a/n531 , \SUBBYTES[0].a/n530 ,
         \SUBBYTES[0].a/n529 , \SUBBYTES[0].a/n528 , \SUBBYTES[0].a/n527 ,
         \SUBBYTES[0].a/n526 , \SUBBYTES[0].a/n525 , \SUBBYTES[0].a/n524 ,
         \SUBBYTES[0].a/n523 , \SUBBYTES[0].a/n522 , \SUBBYTES[0].a/n521 ,
         \SUBBYTES[0].a/n520 , \SUBBYTES[0].a/n519 , \SUBBYTES[0].a/n518 ,
         \SUBBYTES[0].a/n517 , \SUBBYTES[0].a/n516 , \SUBBYTES[0].a/n515 ,
         \SUBBYTES[0].a/n514 , \SUBBYTES[0].a/n513 , \SUBBYTES[0].a/n512 ,
         \SUBBYTES[0].a/n511 , \SUBBYTES[0].a/n510 , \SUBBYTES[0].a/n509 ,
         \SUBBYTES[0].a/n508 , \SUBBYTES[0].a/n507 , \SUBBYTES[0].a/n506 ,
         \SUBBYTES[0].a/n505 , \SUBBYTES[0].a/n504 , \SUBBYTES[0].a/n503 ,
         \SUBBYTES[0].a/n502 , \SUBBYTES[0].a/n501 , \SUBBYTES[0].a/n500 ,
         \SUBBYTES[0].a/n499 , \SUBBYTES[0].a/n498 , \SUBBYTES[0].a/n497 ,
         \SUBBYTES[0].a/n496 , \SUBBYTES[0].a/n495 , \SUBBYTES[0].a/n494 ,
         \SUBBYTES[0].a/n493 , \SUBBYTES[0].a/n492 , \SUBBYTES[0].a/n491 ,
         \SUBBYTES[0].a/n490 , \SUBBYTES[0].a/n489 , \SUBBYTES[0].a/n488 ,
         \SUBBYTES[0].a/n487 , \SUBBYTES[0].a/n486 , \SUBBYTES[0].a/n485 ,
         \SUBBYTES[0].a/n484 , \SUBBYTES[0].a/n483 , \SUBBYTES[0].a/n482 ,
         \SUBBYTES[0].a/n481 , \SUBBYTES[0].a/n480 , \SUBBYTES[0].a/n479 ,
         \SUBBYTES[0].a/n478 , \SUBBYTES[0].a/n477 , \SUBBYTES[0].a/n476 ,
         \SUBBYTES[0].a/n475 , \SUBBYTES[0].a/n474 , \SUBBYTES[0].a/n473 ,
         \SUBBYTES[0].a/n472 , \SUBBYTES[0].a/n471 , \SUBBYTES[0].a/n470 ,
         \SUBBYTES[0].a/n469 , \SUBBYTES[0].a/n468 , \SUBBYTES[0].a/n467 ,
         \SUBBYTES[0].a/n466 , \SUBBYTES[0].a/n465 , \SUBBYTES[0].a/n464 ,
         \SUBBYTES[0].a/n463 , \SUBBYTES[0].a/n462 , \SUBBYTES[0].a/n461 ,
         \SUBBYTES[0].a/n460 , \SUBBYTES[0].a/n459 , \SUBBYTES[0].a/n458 ,
         \SUBBYTES[0].a/n457 , \SUBBYTES[0].a/n456 , \SUBBYTES[0].a/n455 ,
         \SUBBYTES[0].a/n454 , \SUBBYTES[0].a/n453 , \SUBBYTES[0].a/n452 ,
         \SUBBYTES[0].a/n451 , \SUBBYTES[0].a/n450 , \SUBBYTES[0].a/n449 ,
         \SUBBYTES[0].a/n448 , \SUBBYTES[0].a/n447 , \SUBBYTES[0].a/n446 ,
         \SUBBYTES[0].a/n445 , \SUBBYTES[0].a/n444 , \SUBBYTES[0].a/n443 ,
         \SUBBYTES[0].a/n442 , \SUBBYTES[0].a/n441 , \SUBBYTES[0].a/n440 ,
         \SUBBYTES[0].a/n439 , \SUBBYTES[0].a/n438 , \SUBBYTES[0].a/n437 ,
         \SUBBYTES[0].a/n436 , \SUBBYTES[0].a/n435 , \SUBBYTES[0].a/n434 ,
         \SUBBYTES[0].a/n433 , \SUBBYTES[0].a/n432 , \SUBBYTES[0].a/n431 ,
         \SUBBYTES[0].a/n430 , \SUBBYTES[0].a/n429 , \SUBBYTES[0].a/n428 ,
         \SUBBYTES[0].a/n427 , \SUBBYTES[0].a/n426 , \SUBBYTES[0].a/n425 ,
         \SUBBYTES[0].a/n424 , \SUBBYTES[0].a/n423 , \SUBBYTES[0].a/n422 ,
         \SUBBYTES[0].a/n421 , \SUBBYTES[0].a/n420 , \SUBBYTES[0].a/n419 ,
         \SUBBYTES[0].a/n418 , \SUBBYTES[0].a/n417 , \SUBBYTES[0].a/n416 ,
         \SUBBYTES[0].a/n415 , \SUBBYTES[0].a/n414 , \SUBBYTES[0].a/n413 ,
         \SUBBYTES[0].a/n412 , \SUBBYTES[0].a/n411 , \SUBBYTES[0].a/n410 ,
         \SUBBYTES[0].a/n409 , \SUBBYTES[0].a/n408 , \SUBBYTES[0].a/n407 ,
         \SUBBYTES[0].a/n406 , \SUBBYTES[0].a/n405 , \SUBBYTES[0].a/n404 ,
         \SUBBYTES[0].a/n403 , \SUBBYTES[0].a/n402 , \SUBBYTES[0].a/n401 ,
         \SUBBYTES[0].a/n400 , \SUBBYTES[0].a/n399 , \SUBBYTES[0].a/n398 ,
         \SUBBYTES[0].a/n397 , \SUBBYTES[0].a/n396 , \SUBBYTES[0].a/n395 ,
         \SUBBYTES[0].a/n394 , \SUBBYTES[0].a/n393 , \SUBBYTES[0].a/n392 ,
         \SUBBYTES[0].a/n391 , \SUBBYTES[0].a/n390 , \SUBBYTES[0].a/n389 ,
         \SUBBYTES[0].a/n388 , \SUBBYTES[0].a/n387 , \SUBBYTES[0].a/n386 ,
         \SUBBYTES[0].a/n385 , \SUBBYTES[0].a/n160 , \SUBBYTES[0].a/n159 ,
         \SUBBYTES[0].a/n150 , \SUBBYTES[0].a/n149 , \SUBBYTES[0].a/n140 ,
         \SUBBYTES[0].a/n139 , \SUBBYTES[0].a/n130 , \SUBBYTES[0].a/n129 ,
         \SUBBYTES[0].a/n120 , \SUBBYTES[0].a/n119 , \SUBBYTES[0].a/n110 ,
         \SUBBYTES[0].a/n109 , \SUBBYTES[0].a/n100 , \SUBBYTES[0].a/n99 ,
         \SUBBYTES[0].a/n90 , \SUBBYTES[0].a/n89 , \SUBBYTES[0].a/n80 ,
         \SUBBYTES[0].a/n79 , \SUBBYTES[0].a/n70 , \SUBBYTES[0].a/n69 ,
         \SUBBYTES[0].a/n60 , \SUBBYTES[0].a/n59 , \SUBBYTES[0].a/n50 ,
         \SUBBYTES[0].a/n49 , \SUBBYTES[0].a/n40 , \SUBBYTES[0].a/n39 ,
         \SUBBYTES[0].a/n30 , \SUBBYTES[0].a/n29 , \SUBBYTES[0].a/n20 ,
         \SUBBYTES[0].a/n19 , \SUBBYTES[0].a/n10 , \SUBBYTES[0].a/n9 ,
         \SUBBYTES[0].a/w3400 , \SUBBYTES[0].a/w3398 , \SUBBYTES[0].a/w3397 ,
         \SUBBYTES[0].a/w3396 , \SUBBYTES[0].a/w3393 , \SUBBYTES[0].a/w3391 ,
         \SUBBYTES[0].a/w3390 , \SUBBYTES[0].a/w3389 , \SUBBYTES[0].a/w3385 ,
         \SUBBYTES[0].a/w3383 , \SUBBYTES[0].a/w3382 , \SUBBYTES[0].a/w3381 ,
         \SUBBYTES[0].a/w3380 , \SUBBYTES[0].a/w3379 , \SUBBYTES[0].a/w3378 ,
         \SUBBYTES[0].a/w3377 , \SUBBYTES[0].a/w3376 , \SUBBYTES[0].a/w3368 ,
         \SUBBYTES[0].a/w3366 , \SUBBYTES[0].a/w3365 , \SUBBYTES[0].a/w3361 ,
         \SUBBYTES[0].a/w3359 , \SUBBYTES[0].a/w3358 , \SUBBYTES[0].a/w3357 ,
         \SUBBYTES[0].a/w3353 , \SUBBYTES[0].a/w3351 , \SUBBYTES[0].a/w3350 ,
         \SUBBYTES[0].a/w3337 , \SUBBYTES[0].a/w3336 , \SUBBYTES[0].a/w3335 ,
         \SUBBYTES[0].a/w3333 , \SUBBYTES[0].a/w3330 , \SUBBYTES[0].a/w3329 ,
         \SUBBYTES[0].a/w3327 , \SUBBYTES[0].a/w3326 , \SUBBYTES[0].a/w3324 ,
         \SUBBYTES[0].a/w3322 , \SUBBYTES[0].a/w3321 , \SUBBYTES[0].a/w3315 ,
         \SUBBYTES[0].a/w3314 , \SUBBYTES[0].a/w3313 , \SUBBYTES[0].a/w3312 ,
         \SUBBYTES[0].a/w3306 , \SUBBYTES[0].a/w3304 , \SUBBYTES[0].a/w3303 ,
         \SUBBYTES[0].a/w3299 , \SUBBYTES[0].a/w3297 , \SUBBYTES[0].a/w3296 ,
         \SUBBYTES[0].a/w3291 , \SUBBYTES[0].a/w3289 , \SUBBYTES[0].a/w3288 ,
         \SUBBYTES[0].a/w3272 , \SUBBYTES[0].a/w3271 , \SUBBYTES[0].a/w3270 ,
         \SUBBYTES[0].a/w3269 , \SUBBYTES[0].a/w3268 , \SUBBYTES[0].a/w3266 ,
         \SUBBYTES[0].a/w3265 , \SUBBYTES[0].a/w3193 , \SUBBYTES[0].a/w3191 ,
         \SUBBYTES[0].a/w3190 , \SUBBYTES[0].a/w3189 , \SUBBYTES[0].a/w3186 ,
         \SUBBYTES[0].a/w3184 , \SUBBYTES[0].a/w3183 , \SUBBYTES[0].a/w3182 ,
         \SUBBYTES[0].a/w3178 , \SUBBYTES[0].a/w3176 , \SUBBYTES[0].a/w3175 ,
         \SUBBYTES[0].a/w3174 , \SUBBYTES[0].a/w3173 , \SUBBYTES[0].a/w3172 ,
         \SUBBYTES[0].a/w3171 , \SUBBYTES[0].a/w3170 , \SUBBYTES[0].a/w3169 ,
         \SUBBYTES[0].a/w3161 , \SUBBYTES[0].a/w3159 , \SUBBYTES[0].a/w3158 ,
         \SUBBYTES[0].a/w3154 , \SUBBYTES[0].a/w3152 , \SUBBYTES[0].a/w3151 ,
         \SUBBYTES[0].a/w3150 , \SUBBYTES[0].a/w3146 , \SUBBYTES[0].a/w3144 ,
         \SUBBYTES[0].a/w3143 , \SUBBYTES[0].a/w3130 , \SUBBYTES[0].a/w3129 ,
         \SUBBYTES[0].a/w3128 , \SUBBYTES[0].a/w3126 , \SUBBYTES[0].a/w3123 ,
         \SUBBYTES[0].a/w3122 , \SUBBYTES[0].a/w3120 , \SUBBYTES[0].a/w3119 ,
         \SUBBYTES[0].a/w3117 , \SUBBYTES[0].a/w3115 , \SUBBYTES[0].a/w3114 ,
         \SUBBYTES[0].a/w3108 , \SUBBYTES[0].a/w3107 , \SUBBYTES[0].a/w3106 ,
         \SUBBYTES[0].a/w3105 , \SUBBYTES[0].a/w3099 , \SUBBYTES[0].a/w3097 ,
         \SUBBYTES[0].a/w3096 , \SUBBYTES[0].a/w3092 , \SUBBYTES[0].a/w3090 ,
         \SUBBYTES[0].a/w3089 , \SUBBYTES[0].a/w3084 , \SUBBYTES[0].a/w3082 ,
         \SUBBYTES[0].a/w3081 , \SUBBYTES[0].a/w3065 , \SUBBYTES[0].a/w3064 ,
         \SUBBYTES[0].a/w3063 , \SUBBYTES[0].a/w3062 , \SUBBYTES[0].a/w3061 ,
         \SUBBYTES[0].a/w3059 , \SUBBYTES[0].a/w3058 , \SUBBYTES[0].a/w2986 ,
         \SUBBYTES[0].a/w2984 , \SUBBYTES[0].a/w2983 , \SUBBYTES[0].a/w2982 ,
         \SUBBYTES[0].a/w2979 , \SUBBYTES[0].a/w2977 , \SUBBYTES[0].a/w2976 ,
         \SUBBYTES[0].a/w2975 , \SUBBYTES[0].a/w2971 , \SUBBYTES[0].a/w2969 ,
         \SUBBYTES[0].a/w2968 , \SUBBYTES[0].a/w2967 , \SUBBYTES[0].a/w2966 ,
         \SUBBYTES[0].a/w2965 , \SUBBYTES[0].a/w2964 , \SUBBYTES[0].a/w2963 ,
         \SUBBYTES[0].a/w2962 , \SUBBYTES[0].a/w2954 , \SUBBYTES[0].a/w2952 ,
         \SUBBYTES[0].a/w2951 , \SUBBYTES[0].a/w2947 , \SUBBYTES[0].a/w2945 ,
         \SUBBYTES[0].a/w2944 , \SUBBYTES[0].a/w2943 , \SUBBYTES[0].a/w2939 ,
         \SUBBYTES[0].a/w2937 , \SUBBYTES[0].a/w2936 , \SUBBYTES[0].a/w2923 ,
         \SUBBYTES[0].a/w2922 , \SUBBYTES[0].a/w2921 , \SUBBYTES[0].a/w2919 ,
         \SUBBYTES[0].a/w2916 , \SUBBYTES[0].a/w2915 , \SUBBYTES[0].a/w2913 ,
         \SUBBYTES[0].a/w2912 , \SUBBYTES[0].a/w2910 , \SUBBYTES[0].a/w2908 ,
         \SUBBYTES[0].a/w2907 , \SUBBYTES[0].a/w2901 , \SUBBYTES[0].a/w2900 ,
         \SUBBYTES[0].a/w2899 , \SUBBYTES[0].a/w2898 , \SUBBYTES[0].a/w2892 ,
         \SUBBYTES[0].a/w2890 , \SUBBYTES[0].a/w2889 , \SUBBYTES[0].a/w2885 ,
         \SUBBYTES[0].a/w2883 , \SUBBYTES[0].a/w2882 , \SUBBYTES[0].a/w2877 ,
         \SUBBYTES[0].a/w2875 , \SUBBYTES[0].a/w2874 , \SUBBYTES[0].a/w2858 ,
         \SUBBYTES[0].a/w2857 , \SUBBYTES[0].a/w2856 , \SUBBYTES[0].a/w2855 ,
         \SUBBYTES[0].a/w2854 , \SUBBYTES[0].a/w2852 , \SUBBYTES[0].a/w2851 ,
         \SUBBYTES[0].a/w2779 , \SUBBYTES[0].a/w2777 , \SUBBYTES[0].a/w2776 ,
         \SUBBYTES[0].a/w2775 , \SUBBYTES[0].a/w2772 , \SUBBYTES[0].a/w2770 ,
         \SUBBYTES[0].a/w2769 , \SUBBYTES[0].a/w2768 , \SUBBYTES[0].a/w2764 ,
         \SUBBYTES[0].a/w2762 , \SUBBYTES[0].a/w2761 , \SUBBYTES[0].a/w2760 ,
         \SUBBYTES[0].a/w2759 , \SUBBYTES[0].a/w2758 , \SUBBYTES[0].a/w2757 ,
         \SUBBYTES[0].a/w2756 , \SUBBYTES[0].a/w2755 , \SUBBYTES[0].a/w2747 ,
         \SUBBYTES[0].a/w2745 , \SUBBYTES[0].a/w2744 , \SUBBYTES[0].a/w2740 ,
         \SUBBYTES[0].a/w2738 , \SUBBYTES[0].a/w2737 , \SUBBYTES[0].a/w2736 ,
         \SUBBYTES[0].a/w2732 , \SUBBYTES[0].a/w2730 , \SUBBYTES[0].a/w2729 ,
         \SUBBYTES[0].a/w2716 , \SUBBYTES[0].a/w2715 , \SUBBYTES[0].a/w2714 ,
         \SUBBYTES[0].a/w2712 , \SUBBYTES[0].a/w2709 , \SUBBYTES[0].a/w2708 ,
         \SUBBYTES[0].a/w2706 , \SUBBYTES[0].a/w2705 , \SUBBYTES[0].a/w2703 ,
         \SUBBYTES[0].a/w2701 , \SUBBYTES[0].a/w2700 , \SUBBYTES[0].a/w2694 ,
         \SUBBYTES[0].a/w2693 , \SUBBYTES[0].a/w2692 , \SUBBYTES[0].a/w2691 ,
         \SUBBYTES[0].a/w2685 , \SUBBYTES[0].a/w2683 , \SUBBYTES[0].a/w2682 ,
         \SUBBYTES[0].a/w2678 , \SUBBYTES[0].a/w2676 , \SUBBYTES[0].a/w2675 ,
         \SUBBYTES[0].a/w2670 , \SUBBYTES[0].a/w2668 , \SUBBYTES[0].a/w2667 ,
         \SUBBYTES[0].a/w2651 , \SUBBYTES[0].a/w2650 , \SUBBYTES[0].a/w2649 ,
         \SUBBYTES[0].a/w2648 , \SUBBYTES[0].a/w2647 , \SUBBYTES[0].a/w2645 ,
         \SUBBYTES[0].a/w2644 , \SUBBYTES[0].a/w2572 , \SUBBYTES[0].a/w2570 ,
         \SUBBYTES[0].a/w2569 , \SUBBYTES[0].a/w2568 , \SUBBYTES[0].a/w2565 ,
         \SUBBYTES[0].a/w2563 , \SUBBYTES[0].a/w2562 , \SUBBYTES[0].a/w2561 ,
         \SUBBYTES[0].a/w2557 , \SUBBYTES[0].a/w2555 , \SUBBYTES[0].a/w2554 ,
         \SUBBYTES[0].a/w2553 , \SUBBYTES[0].a/w2552 , \SUBBYTES[0].a/w2551 ,
         \SUBBYTES[0].a/w2550 , \SUBBYTES[0].a/w2549 , \SUBBYTES[0].a/w2548 ,
         \SUBBYTES[0].a/w2540 , \SUBBYTES[0].a/w2538 , \SUBBYTES[0].a/w2537 ,
         \SUBBYTES[0].a/w2533 , \SUBBYTES[0].a/w2531 , \SUBBYTES[0].a/w2530 ,
         \SUBBYTES[0].a/w2529 , \SUBBYTES[0].a/w2525 , \SUBBYTES[0].a/w2523 ,
         \SUBBYTES[0].a/w2522 , \SUBBYTES[0].a/w2509 , \SUBBYTES[0].a/w2508 ,
         \SUBBYTES[0].a/w2507 , \SUBBYTES[0].a/w2505 , \SUBBYTES[0].a/w2502 ,
         \SUBBYTES[0].a/w2501 , \SUBBYTES[0].a/w2499 , \SUBBYTES[0].a/w2498 ,
         \SUBBYTES[0].a/w2496 , \SUBBYTES[0].a/w2494 , \SUBBYTES[0].a/w2493 ,
         \SUBBYTES[0].a/w2487 , \SUBBYTES[0].a/w2486 , \SUBBYTES[0].a/w2485 ,
         \SUBBYTES[0].a/w2484 , \SUBBYTES[0].a/w2478 , \SUBBYTES[0].a/w2476 ,
         \SUBBYTES[0].a/w2475 , \SUBBYTES[0].a/w2471 , \SUBBYTES[0].a/w2469 ,
         \SUBBYTES[0].a/w2468 , \SUBBYTES[0].a/w2463 , \SUBBYTES[0].a/w2461 ,
         \SUBBYTES[0].a/w2460 , \SUBBYTES[0].a/w2444 , \SUBBYTES[0].a/w2443 ,
         \SUBBYTES[0].a/w2442 , \SUBBYTES[0].a/w2441 , \SUBBYTES[0].a/w2440 ,
         \SUBBYTES[0].a/w2438 , \SUBBYTES[0].a/w2437 , \SUBBYTES[0].a/w2365 ,
         \SUBBYTES[0].a/w2363 , \SUBBYTES[0].a/w2362 , \SUBBYTES[0].a/w2361 ,
         \SUBBYTES[0].a/w2358 , \SUBBYTES[0].a/w2356 , \SUBBYTES[0].a/w2355 ,
         \SUBBYTES[0].a/w2354 , \SUBBYTES[0].a/w2350 , \SUBBYTES[0].a/w2348 ,
         \SUBBYTES[0].a/w2347 , \SUBBYTES[0].a/w2346 , \SUBBYTES[0].a/w2345 ,
         \SUBBYTES[0].a/w2344 , \SUBBYTES[0].a/w2343 , \SUBBYTES[0].a/w2342 ,
         \SUBBYTES[0].a/w2341 , \SUBBYTES[0].a/w2333 , \SUBBYTES[0].a/w2331 ,
         \SUBBYTES[0].a/w2330 , \SUBBYTES[0].a/w2326 , \SUBBYTES[0].a/w2324 ,
         \SUBBYTES[0].a/w2323 , \SUBBYTES[0].a/w2322 , \SUBBYTES[0].a/w2318 ,
         \SUBBYTES[0].a/w2316 , \SUBBYTES[0].a/w2315 , \SUBBYTES[0].a/w2302 ,
         \SUBBYTES[0].a/w2301 , \SUBBYTES[0].a/w2300 , \SUBBYTES[0].a/w2298 ,
         \SUBBYTES[0].a/w2295 , \SUBBYTES[0].a/w2294 , \SUBBYTES[0].a/w2292 ,
         \SUBBYTES[0].a/w2291 , \SUBBYTES[0].a/w2289 , \SUBBYTES[0].a/w2287 ,
         \SUBBYTES[0].a/w2286 , \SUBBYTES[0].a/w2280 , \SUBBYTES[0].a/w2279 ,
         \SUBBYTES[0].a/w2278 , \SUBBYTES[0].a/w2277 , \SUBBYTES[0].a/w2271 ,
         \SUBBYTES[0].a/w2269 , \SUBBYTES[0].a/w2268 , \SUBBYTES[0].a/w2264 ,
         \SUBBYTES[0].a/w2262 , \SUBBYTES[0].a/w2261 , \SUBBYTES[0].a/w2256 ,
         \SUBBYTES[0].a/w2254 , \SUBBYTES[0].a/w2253 , \SUBBYTES[0].a/w2237 ,
         \SUBBYTES[0].a/w2236 , \SUBBYTES[0].a/w2235 , \SUBBYTES[0].a/w2234 ,
         \SUBBYTES[0].a/w2233 , \SUBBYTES[0].a/w2231 , \SUBBYTES[0].a/w2230 ,
         \SUBBYTES[0].a/w2158 , \SUBBYTES[0].a/w2156 , \SUBBYTES[0].a/w2155 ,
         \SUBBYTES[0].a/w2154 , \SUBBYTES[0].a/w2151 , \SUBBYTES[0].a/w2149 ,
         \SUBBYTES[0].a/w2148 , \SUBBYTES[0].a/w2147 , \SUBBYTES[0].a/w2143 ,
         \SUBBYTES[0].a/w2141 , \SUBBYTES[0].a/w2140 , \SUBBYTES[0].a/w2139 ,
         \SUBBYTES[0].a/w2138 , \SUBBYTES[0].a/w2137 , \SUBBYTES[0].a/w2136 ,
         \SUBBYTES[0].a/w2135 , \SUBBYTES[0].a/w2134 , \SUBBYTES[0].a/w2126 ,
         \SUBBYTES[0].a/w2124 , \SUBBYTES[0].a/w2123 , \SUBBYTES[0].a/w2119 ,
         \SUBBYTES[0].a/w2117 , \SUBBYTES[0].a/w2116 , \SUBBYTES[0].a/w2115 ,
         \SUBBYTES[0].a/w2111 , \SUBBYTES[0].a/w2109 , \SUBBYTES[0].a/w2108 ,
         \SUBBYTES[0].a/w2095 , \SUBBYTES[0].a/w2094 , \SUBBYTES[0].a/w2093 ,
         \SUBBYTES[0].a/w2091 , \SUBBYTES[0].a/w2088 , \SUBBYTES[0].a/w2087 ,
         \SUBBYTES[0].a/w2085 , \SUBBYTES[0].a/w2084 , \SUBBYTES[0].a/w2082 ,
         \SUBBYTES[0].a/w2080 , \SUBBYTES[0].a/w2079 , \SUBBYTES[0].a/w2073 ,
         \SUBBYTES[0].a/w2072 , \SUBBYTES[0].a/w2071 , \SUBBYTES[0].a/w2070 ,
         \SUBBYTES[0].a/w2064 , \SUBBYTES[0].a/w2062 , \SUBBYTES[0].a/w2061 ,
         \SUBBYTES[0].a/w2057 , \SUBBYTES[0].a/w2055 , \SUBBYTES[0].a/w2054 ,
         \SUBBYTES[0].a/w2049 , \SUBBYTES[0].a/w2047 , \SUBBYTES[0].a/w2046 ,
         \SUBBYTES[0].a/w2030 , \SUBBYTES[0].a/w2029 , \SUBBYTES[0].a/w2028 ,
         \SUBBYTES[0].a/w2027 , \SUBBYTES[0].a/w2026 , \SUBBYTES[0].a/w2024 ,
         \SUBBYTES[0].a/w2023 , \SUBBYTES[0].a/w1951 , \SUBBYTES[0].a/w1949 ,
         \SUBBYTES[0].a/w1948 , \SUBBYTES[0].a/w1947 , \SUBBYTES[0].a/w1944 ,
         \SUBBYTES[0].a/w1942 , \SUBBYTES[0].a/w1941 , \SUBBYTES[0].a/w1940 ,
         \SUBBYTES[0].a/w1936 , \SUBBYTES[0].a/w1934 , \SUBBYTES[0].a/w1933 ,
         \SUBBYTES[0].a/w1932 , \SUBBYTES[0].a/w1931 , \SUBBYTES[0].a/w1930 ,
         \SUBBYTES[0].a/w1929 , \SUBBYTES[0].a/w1928 , \SUBBYTES[0].a/w1927 ,
         \SUBBYTES[0].a/w1919 , \SUBBYTES[0].a/w1917 , \SUBBYTES[0].a/w1916 ,
         \SUBBYTES[0].a/w1912 , \SUBBYTES[0].a/w1910 , \SUBBYTES[0].a/w1909 ,
         \SUBBYTES[0].a/w1908 , \SUBBYTES[0].a/w1904 , \SUBBYTES[0].a/w1902 ,
         \SUBBYTES[0].a/w1901 , \SUBBYTES[0].a/w1888 , \SUBBYTES[0].a/w1887 ,
         \SUBBYTES[0].a/w1886 , \SUBBYTES[0].a/w1884 , \SUBBYTES[0].a/w1881 ,
         \SUBBYTES[0].a/w1880 , \SUBBYTES[0].a/w1878 , \SUBBYTES[0].a/w1877 ,
         \SUBBYTES[0].a/w1875 , \SUBBYTES[0].a/w1873 , \SUBBYTES[0].a/w1872 ,
         \SUBBYTES[0].a/w1866 , \SUBBYTES[0].a/w1865 , \SUBBYTES[0].a/w1864 ,
         \SUBBYTES[0].a/w1863 , \SUBBYTES[0].a/w1857 , \SUBBYTES[0].a/w1855 ,
         \SUBBYTES[0].a/w1854 , \SUBBYTES[0].a/w1850 , \SUBBYTES[0].a/w1848 ,
         \SUBBYTES[0].a/w1847 , \SUBBYTES[0].a/w1842 , \SUBBYTES[0].a/w1840 ,
         \SUBBYTES[0].a/w1839 , \SUBBYTES[0].a/w1823 , \SUBBYTES[0].a/w1822 ,
         \SUBBYTES[0].a/w1821 , \SUBBYTES[0].a/w1820 , \SUBBYTES[0].a/w1819 ,
         \SUBBYTES[0].a/w1817 , \SUBBYTES[0].a/w1816 , \SUBBYTES[0].a/w1744 ,
         \SUBBYTES[0].a/w1742 , \SUBBYTES[0].a/w1741 , \SUBBYTES[0].a/w1740 ,
         \SUBBYTES[0].a/w1737 , \SUBBYTES[0].a/w1735 , \SUBBYTES[0].a/w1734 ,
         \SUBBYTES[0].a/w1733 , \SUBBYTES[0].a/w1729 , \SUBBYTES[0].a/w1727 ,
         \SUBBYTES[0].a/w1726 , \SUBBYTES[0].a/w1725 , \SUBBYTES[0].a/w1724 ,
         \SUBBYTES[0].a/w1723 , \SUBBYTES[0].a/w1722 , \SUBBYTES[0].a/w1721 ,
         \SUBBYTES[0].a/w1720 , \SUBBYTES[0].a/w1712 , \SUBBYTES[0].a/w1710 ,
         \SUBBYTES[0].a/w1709 , \SUBBYTES[0].a/w1705 , \SUBBYTES[0].a/w1703 ,
         \SUBBYTES[0].a/w1702 , \SUBBYTES[0].a/w1701 , \SUBBYTES[0].a/w1697 ,
         \SUBBYTES[0].a/w1695 , \SUBBYTES[0].a/w1694 , \SUBBYTES[0].a/w1681 ,
         \SUBBYTES[0].a/w1680 , \SUBBYTES[0].a/w1679 , \SUBBYTES[0].a/w1677 ,
         \SUBBYTES[0].a/w1674 , \SUBBYTES[0].a/w1673 , \SUBBYTES[0].a/w1671 ,
         \SUBBYTES[0].a/w1670 , \SUBBYTES[0].a/w1668 , \SUBBYTES[0].a/w1666 ,
         \SUBBYTES[0].a/w1665 , \SUBBYTES[0].a/w1659 , \SUBBYTES[0].a/w1658 ,
         \SUBBYTES[0].a/w1657 , \SUBBYTES[0].a/w1656 , \SUBBYTES[0].a/w1650 ,
         \SUBBYTES[0].a/w1648 , \SUBBYTES[0].a/w1647 , \SUBBYTES[0].a/w1643 ,
         \SUBBYTES[0].a/w1641 , \SUBBYTES[0].a/w1640 , \SUBBYTES[0].a/w1635 ,
         \SUBBYTES[0].a/w1633 , \SUBBYTES[0].a/w1632 , \SUBBYTES[0].a/w1616 ,
         \SUBBYTES[0].a/w1615 , \SUBBYTES[0].a/w1614 , \SUBBYTES[0].a/w1613 ,
         \SUBBYTES[0].a/w1612 , \SUBBYTES[0].a/w1610 , \SUBBYTES[0].a/w1609 ,
         \SUBBYTES[0].a/w1537 , \SUBBYTES[0].a/w1535 , \SUBBYTES[0].a/w1534 ,
         \SUBBYTES[0].a/w1533 , \SUBBYTES[0].a/w1530 , \SUBBYTES[0].a/w1528 ,
         \SUBBYTES[0].a/w1527 , \SUBBYTES[0].a/w1526 , \SUBBYTES[0].a/w1522 ,
         \SUBBYTES[0].a/w1520 , \SUBBYTES[0].a/w1519 , \SUBBYTES[0].a/w1518 ,
         \SUBBYTES[0].a/w1517 , \SUBBYTES[0].a/w1516 , \SUBBYTES[0].a/w1515 ,
         \SUBBYTES[0].a/w1514 , \SUBBYTES[0].a/w1513 , \SUBBYTES[0].a/w1505 ,
         \SUBBYTES[0].a/w1503 , \SUBBYTES[0].a/w1502 , \SUBBYTES[0].a/w1498 ,
         \SUBBYTES[0].a/w1496 , \SUBBYTES[0].a/w1495 , \SUBBYTES[0].a/w1494 ,
         \SUBBYTES[0].a/w1490 , \SUBBYTES[0].a/w1488 , \SUBBYTES[0].a/w1487 ,
         \SUBBYTES[0].a/w1474 , \SUBBYTES[0].a/w1473 , \SUBBYTES[0].a/w1472 ,
         \SUBBYTES[0].a/w1470 , \SUBBYTES[0].a/w1467 , \SUBBYTES[0].a/w1466 ,
         \SUBBYTES[0].a/w1464 , \SUBBYTES[0].a/w1463 , \SUBBYTES[0].a/w1461 ,
         \SUBBYTES[0].a/w1459 , \SUBBYTES[0].a/w1458 , \SUBBYTES[0].a/w1452 ,
         \SUBBYTES[0].a/w1451 , \SUBBYTES[0].a/w1450 , \SUBBYTES[0].a/w1449 ,
         \SUBBYTES[0].a/w1443 , \SUBBYTES[0].a/w1441 , \SUBBYTES[0].a/w1440 ,
         \SUBBYTES[0].a/w1436 , \SUBBYTES[0].a/w1434 , \SUBBYTES[0].a/w1433 ,
         \SUBBYTES[0].a/w1428 , \SUBBYTES[0].a/w1426 , \SUBBYTES[0].a/w1425 ,
         \SUBBYTES[0].a/w1409 , \SUBBYTES[0].a/w1408 , \SUBBYTES[0].a/w1407 ,
         \SUBBYTES[0].a/w1406 , \SUBBYTES[0].a/w1405 , \SUBBYTES[0].a/w1403 ,
         \SUBBYTES[0].a/w1402 , \SUBBYTES[0].a/w1330 , \SUBBYTES[0].a/w1328 ,
         \SUBBYTES[0].a/w1327 , \SUBBYTES[0].a/w1326 , \SUBBYTES[0].a/w1323 ,
         \SUBBYTES[0].a/w1321 , \SUBBYTES[0].a/w1320 , \SUBBYTES[0].a/w1319 ,
         \SUBBYTES[0].a/w1315 , \SUBBYTES[0].a/w1313 , \SUBBYTES[0].a/w1312 ,
         \SUBBYTES[0].a/w1311 , \SUBBYTES[0].a/w1310 , \SUBBYTES[0].a/w1309 ,
         \SUBBYTES[0].a/w1308 , \SUBBYTES[0].a/w1307 , \SUBBYTES[0].a/w1306 ,
         \SUBBYTES[0].a/w1298 , \SUBBYTES[0].a/w1296 , \SUBBYTES[0].a/w1295 ,
         \SUBBYTES[0].a/w1291 , \SUBBYTES[0].a/w1289 , \SUBBYTES[0].a/w1288 ,
         \SUBBYTES[0].a/w1287 , \SUBBYTES[0].a/w1283 , \SUBBYTES[0].a/w1281 ,
         \SUBBYTES[0].a/w1280 , \SUBBYTES[0].a/w1267 , \SUBBYTES[0].a/w1266 ,
         \SUBBYTES[0].a/w1265 , \SUBBYTES[0].a/w1263 , \SUBBYTES[0].a/w1260 ,
         \SUBBYTES[0].a/w1259 , \SUBBYTES[0].a/w1257 , \SUBBYTES[0].a/w1256 ,
         \SUBBYTES[0].a/w1254 , \SUBBYTES[0].a/w1252 , \SUBBYTES[0].a/w1251 ,
         \SUBBYTES[0].a/w1245 , \SUBBYTES[0].a/w1244 , \SUBBYTES[0].a/w1243 ,
         \SUBBYTES[0].a/w1242 , \SUBBYTES[0].a/w1236 , \SUBBYTES[0].a/w1234 ,
         \SUBBYTES[0].a/w1233 , \SUBBYTES[0].a/w1229 , \SUBBYTES[0].a/w1227 ,
         \SUBBYTES[0].a/w1226 , \SUBBYTES[0].a/w1221 , \SUBBYTES[0].a/w1219 ,
         \SUBBYTES[0].a/w1218 , \SUBBYTES[0].a/w1202 , \SUBBYTES[0].a/w1201 ,
         \SUBBYTES[0].a/w1200 , \SUBBYTES[0].a/w1199 , \SUBBYTES[0].a/w1198 ,
         \SUBBYTES[0].a/w1196 , \SUBBYTES[0].a/w1195 , \SUBBYTES[0].a/w1123 ,
         \SUBBYTES[0].a/w1121 , \SUBBYTES[0].a/w1120 , \SUBBYTES[0].a/w1119 ,
         \SUBBYTES[0].a/w1116 , \SUBBYTES[0].a/w1114 , \SUBBYTES[0].a/w1113 ,
         \SUBBYTES[0].a/w1112 , \SUBBYTES[0].a/w1108 , \SUBBYTES[0].a/w1106 ,
         \SUBBYTES[0].a/w1105 , \SUBBYTES[0].a/w1104 , \SUBBYTES[0].a/w1103 ,
         \SUBBYTES[0].a/w1102 , \SUBBYTES[0].a/w1101 , \SUBBYTES[0].a/w1100 ,
         \SUBBYTES[0].a/w1099 , \SUBBYTES[0].a/w1091 , \SUBBYTES[0].a/w1089 ,
         \SUBBYTES[0].a/w1088 , \SUBBYTES[0].a/w1084 , \SUBBYTES[0].a/w1082 ,
         \SUBBYTES[0].a/w1081 , \SUBBYTES[0].a/w1080 , \SUBBYTES[0].a/w1076 ,
         \SUBBYTES[0].a/w1074 , \SUBBYTES[0].a/w1073 , \SUBBYTES[0].a/w1060 ,
         \SUBBYTES[0].a/w1059 , \SUBBYTES[0].a/w1058 , \SUBBYTES[0].a/w1056 ,
         \SUBBYTES[0].a/w1053 , \SUBBYTES[0].a/w1052 , \SUBBYTES[0].a/w1050 ,
         \SUBBYTES[0].a/w1049 , \SUBBYTES[0].a/w1047 , \SUBBYTES[0].a/w1045 ,
         \SUBBYTES[0].a/w1044 , \SUBBYTES[0].a/w1038 , \SUBBYTES[0].a/w1037 ,
         \SUBBYTES[0].a/w1036 , \SUBBYTES[0].a/w1035 , \SUBBYTES[0].a/w1029 ,
         \SUBBYTES[0].a/w1027 , \SUBBYTES[0].a/w1026 , \SUBBYTES[0].a/w1022 ,
         \SUBBYTES[0].a/w1020 , \SUBBYTES[0].a/w1019 , \SUBBYTES[0].a/w1014 ,
         \SUBBYTES[0].a/w1012 , \SUBBYTES[0].a/w1011 , \SUBBYTES[0].a/w995 ,
         \SUBBYTES[0].a/w994 , \SUBBYTES[0].a/w993 , \SUBBYTES[0].a/w992 ,
         \SUBBYTES[0].a/w991 , \SUBBYTES[0].a/w989 , \SUBBYTES[0].a/w988 ,
         \SUBBYTES[0].a/w916 , \SUBBYTES[0].a/w914 , \SUBBYTES[0].a/w913 ,
         \SUBBYTES[0].a/w912 , \SUBBYTES[0].a/w909 , \SUBBYTES[0].a/w907 ,
         \SUBBYTES[0].a/w906 , \SUBBYTES[0].a/w905 , \SUBBYTES[0].a/w901 ,
         \SUBBYTES[0].a/w899 , \SUBBYTES[0].a/w898 , \SUBBYTES[0].a/w897 ,
         \SUBBYTES[0].a/w896 , \SUBBYTES[0].a/w895 , \SUBBYTES[0].a/w894 ,
         \SUBBYTES[0].a/w893 , \SUBBYTES[0].a/w892 , \SUBBYTES[0].a/w884 ,
         \SUBBYTES[0].a/w882 , \SUBBYTES[0].a/w881 , \SUBBYTES[0].a/w877 ,
         \SUBBYTES[0].a/w875 , \SUBBYTES[0].a/w874 , \SUBBYTES[0].a/w873 ,
         \SUBBYTES[0].a/w869 , \SUBBYTES[0].a/w867 , \SUBBYTES[0].a/w866 ,
         \SUBBYTES[0].a/w853 , \SUBBYTES[0].a/w852 , \SUBBYTES[0].a/w851 ,
         \SUBBYTES[0].a/w849 , \SUBBYTES[0].a/w846 , \SUBBYTES[0].a/w845 ,
         \SUBBYTES[0].a/w843 , \SUBBYTES[0].a/w842 , \SUBBYTES[0].a/w840 ,
         \SUBBYTES[0].a/w838 , \SUBBYTES[0].a/w837 , \SUBBYTES[0].a/w831 ,
         \SUBBYTES[0].a/w830 , \SUBBYTES[0].a/w829 , \SUBBYTES[0].a/w828 ,
         \SUBBYTES[0].a/w822 , \SUBBYTES[0].a/w820 , \SUBBYTES[0].a/w819 ,
         \SUBBYTES[0].a/w815 , \SUBBYTES[0].a/w813 , \SUBBYTES[0].a/w812 ,
         \SUBBYTES[0].a/w807 , \SUBBYTES[0].a/w805 , \SUBBYTES[0].a/w804 ,
         \SUBBYTES[0].a/w788 , \SUBBYTES[0].a/w787 , \SUBBYTES[0].a/w786 ,
         \SUBBYTES[0].a/w785 , \SUBBYTES[0].a/w784 , \SUBBYTES[0].a/w782 ,
         \SUBBYTES[0].a/w781 , \SUBBYTES[0].a/w709 , \SUBBYTES[0].a/w707 ,
         \SUBBYTES[0].a/w706 , \SUBBYTES[0].a/w705 , \SUBBYTES[0].a/w702 ,
         \SUBBYTES[0].a/w700 , \SUBBYTES[0].a/w699 , \SUBBYTES[0].a/w698 ,
         \SUBBYTES[0].a/w694 , \SUBBYTES[0].a/w692 , \SUBBYTES[0].a/w691 ,
         \SUBBYTES[0].a/w690 , \SUBBYTES[0].a/w689 , \SUBBYTES[0].a/w688 ,
         \SUBBYTES[0].a/w687 , \SUBBYTES[0].a/w686 , \SUBBYTES[0].a/w685 ,
         \SUBBYTES[0].a/w677 , \SUBBYTES[0].a/w675 , \SUBBYTES[0].a/w674 ,
         \SUBBYTES[0].a/w670 , \SUBBYTES[0].a/w668 , \SUBBYTES[0].a/w667 ,
         \SUBBYTES[0].a/w666 , \SUBBYTES[0].a/w662 , \SUBBYTES[0].a/w660 ,
         \SUBBYTES[0].a/w659 , \SUBBYTES[0].a/w646 , \SUBBYTES[0].a/w645 ,
         \SUBBYTES[0].a/w644 , \SUBBYTES[0].a/w642 , \SUBBYTES[0].a/w639 ,
         \SUBBYTES[0].a/w638 , \SUBBYTES[0].a/w636 , \SUBBYTES[0].a/w635 ,
         \SUBBYTES[0].a/w633 , \SUBBYTES[0].a/w631 , \SUBBYTES[0].a/w630 ,
         \SUBBYTES[0].a/w624 , \SUBBYTES[0].a/w623 , \SUBBYTES[0].a/w622 ,
         \SUBBYTES[0].a/w621 , \SUBBYTES[0].a/w615 , \SUBBYTES[0].a/w613 ,
         \SUBBYTES[0].a/w612 , \SUBBYTES[0].a/w608 , \SUBBYTES[0].a/w606 ,
         \SUBBYTES[0].a/w605 , \SUBBYTES[0].a/w600 , \SUBBYTES[0].a/w598 ,
         \SUBBYTES[0].a/w597 , \SUBBYTES[0].a/w581 , \SUBBYTES[0].a/w580 ,
         \SUBBYTES[0].a/w579 , \SUBBYTES[0].a/w578 , \SUBBYTES[0].a/w577 ,
         \SUBBYTES[0].a/w575 , \SUBBYTES[0].a/w574 , \SUBBYTES[0].a/w502 ,
         \SUBBYTES[0].a/w500 , \SUBBYTES[0].a/w499 , \SUBBYTES[0].a/w498 ,
         \SUBBYTES[0].a/w495 , \SUBBYTES[0].a/w493 , \SUBBYTES[0].a/w492 ,
         \SUBBYTES[0].a/w491 , \SUBBYTES[0].a/w487 , \SUBBYTES[0].a/w485 ,
         \SUBBYTES[0].a/w484 , \SUBBYTES[0].a/w483 , \SUBBYTES[0].a/w482 ,
         \SUBBYTES[0].a/w481 , \SUBBYTES[0].a/w480 , \SUBBYTES[0].a/w479 ,
         \SUBBYTES[0].a/w478 , \SUBBYTES[0].a/w470 , \SUBBYTES[0].a/w468 ,
         \SUBBYTES[0].a/w467 , \SUBBYTES[0].a/w463 , \SUBBYTES[0].a/w461 ,
         \SUBBYTES[0].a/w460 , \SUBBYTES[0].a/w459 , \SUBBYTES[0].a/w455 ,
         \SUBBYTES[0].a/w453 , \SUBBYTES[0].a/w452 , \SUBBYTES[0].a/w439 ,
         \SUBBYTES[0].a/w438 , \SUBBYTES[0].a/w437 , \SUBBYTES[0].a/w435 ,
         \SUBBYTES[0].a/w432 , \SUBBYTES[0].a/w431 , \SUBBYTES[0].a/w429 ,
         \SUBBYTES[0].a/w428 , \SUBBYTES[0].a/w426 , \SUBBYTES[0].a/w424 ,
         \SUBBYTES[0].a/w423 , \SUBBYTES[0].a/w417 , \SUBBYTES[0].a/w416 ,
         \SUBBYTES[0].a/w415 , \SUBBYTES[0].a/w414 , \SUBBYTES[0].a/w408 ,
         \SUBBYTES[0].a/w406 , \SUBBYTES[0].a/w405 , \SUBBYTES[0].a/w401 ,
         \SUBBYTES[0].a/w399 , \SUBBYTES[0].a/w398 , \SUBBYTES[0].a/w393 ,
         \SUBBYTES[0].a/w391 , \SUBBYTES[0].a/w390 , \SUBBYTES[0].a/w374 ,
         \SUBBYTES[0].a/w373 , \SUBBYTES[0].a/w372 , \SUBBYTES[0].a/w371 ,
         \SUBBYTES[0].a/w370 , \SUBBYTES[0].a/w368 , \SUBBYTES[0].a/w367 ,
         \SUBBYTES[0].a/w295 , \SUBBYTES[0].a/w293 , \SUBBYTES[0].a/w292 ,
         \SUBBYTES[0].a/w291 , \SUBBYTES[0].a/w288 , \SUBBYTES[0].a/w286 ,
         \SUBBYTES[0].a/w285 , \SUBBYTES[0].a/w284 , \SUBBYTES[0].a/w280 ,
         \SUBBYTES[0].a/w278 , \SUBBYTES[0].a/w277 , \SUBBYTES[0].a/w276 ,
         \SUBBYTES[0].a/w275 , \SUBBYTES[0].a/w274 , \SUBBYTES[0].a/w273 ,
         \SUBBYTES[0].a/w272 , \SUBBYTES[0].a/w271 , \SUBBYTES[0].a/w263 ,
         \SUBBYTES[0].a/w261 , \SUBBYTES[0].a/w260 , \SUBBYTES[0].a/w256 ,
         \SUBBYTES[0].a/w254 , \SUBBYTES[0].a/w253 , \SUBBYTES[0].a/w252 ,
         \SUBBYTES[0].a/w248 , \SUBBYTES[0].a/w246 , \SUBBYTES[0].a/w245 ,
         \SUBBYTES[0].a/w232 , \SUBBYTES[0].a/w231 , \SUBBYTES[0].a/w230 ,
         \SUBBYTES[0].a/w228 , \SUBBYTES[0].a/w225 , \SUBBYTES[0].a/w224 ,
         \SUBBYTES[0].a/w222 , \SUBBYTES[0].a/w221 , \SUBBYTES[0].a/w219 ,
         \SUBBYTES[0].a/w217 , \SUBBYTES[0].a/w216 , \SUBBYTES[0].a/w210 ,
         \SUBBYTES[0].a/w209 , \SUBBYTES[0].a/w208 , \SUBBYTES[0].a/w207 ,
         \SUBBYTES[0].a/w201 , \SUBBYTES[0].a/w199 , \SUBBYTES[0].a/w198 ,
         \SUBBYTES[0].a/w194 , \SUBBYTES[0].a/w192 , \SUBBYTES[0].a/w191 ,
         \SUBBYTES[0].a/w186 , \SUBBYTES[0].a/w184 , \SUBBYTES[0].a/w183 ,
         \SUBBYTES[0].a/w167 , \SUBBYTES[0].a/w166 , \SUBBYTES[0].a/w165 ,
         \SUBBYTES[0].a/w164 , \SUBBYTES[0].a/w163 , \SUBBYTES[0].a/w161 ,
         \SUBBYTES[0].a/w160 , \MIXCOLUMNS[0].d/n304 , \MIXCOLUMNS[0].d/n303 ,
         \MIXCOLUMNS[0].d/n302 , \MIXCOLUMNS[0].d/n301 ,
         \MIXCOLUMNS[0].d/n300 , \MIXCOLUMNS[0].d/n299 ,
         \MIXCOLUMNS[0].d/n298 , \MIXCOLUMNS[0].d/n297 ,
         \MIXCOLUMNS[0].d/n296 , \MIXCOLUMNS[0].d/n295 ,
         \MIXCOLUMNS[0].d/n294 , \MIXCOLUMNS[0].d/n293 ,
         \MIXCOLUMNS[0].d/n292 , \MIXCOLUMNS[0].d/n291 ,
         \MIXCOLUMNS[0].d/n290 , \MIXCOLUMNS[0].d/n289 ,
         \MIXCOLUMNS[0].d/n288 , \MIXCOLUMNS[0].d/n287 ,
         \MIXCOLUMNS[0].d/n286 , \MIXCOLUMNS[0].d/n285 ,
         \MIXCOLUMNS[0].d/n284 , \MIXCOLUMNS[0].d/n283 ,
         \MIXCOLUMNS[0].d/n282 , \MIXCOLUMNS[0].d/n281 ,
         \MIXCOLUMNS[0].d/n280 , \MIXCOLUMNS[0].d/n279 ,
         \MIXCOLUMNS[0].d/n278 , \MIXCOLUMNS[0].d/n277 ,
         \MIXCOLUMNS[0].d/n276 , \MIXCOLUMNS[0].d/n275 ,
         \MIXCOLUMNS[0].d/n274 , \MIXCOLUMNS[0].d/n273 ,
         \MIXCOLUMNS[0].d/n272 , \MIXCOLUMNS[0].d/n271 ,
         \MIXCOLUMNS[0].d/n270 , \MIXCOLUMNS[0].d/n269 ,
         \MIXCOLUMNS[0].d/n268 , \MIXCOLUMNS[0].d/n267 ,
         \MIXCOLUMNS[0].d/n266 , \MIXCOLUMNS[0].d/n265 ,
         \MIXCOLUMNS[0].d/n264 , \MIXCOLUMNS[0].d/n263 ,
         \MIXCOLUMNS[0].d/n262 , \MIXCOLUMNS[0].d/n261 ,
         \MIXCOLUMNS[0].d/n260 , \MIXCOLUMNS[0].d/n259 ,
         \MIXCOLUMNS[0].d/n258 , \MIXCOLUMNS[0].d/n257 ,
         \MIXCOLUMNS[0].d/n256 , \MIXCOLUMNS[0].d/n255 ,
         \MIXCOLUMNS[0].d/n254 , \MIXCOLUMNS[0].d/n253 ,
         \MIXCOLUMNS[0].d/n252 , \MIXCOLUMNS[0].d/n251 ,
         \MIXCOLUMNS[0].d/n250 , \MIXCOLUMNS[0].d/n249 ,
         \MIXCOLUMNS[0].d/n248 , \MIXCOLUMNS[0].d/n247 ,
         \MIXCOLUMNS[0].d/n246 , \MIXCOLUMNS[0].d/n245 ,
         \MIXCOLUMNS[0].d/n244 , \MIXCOLUMNS[0].d/n243 ,
         \MIXCOLUMNS[0].d/n242 , \MIXCOLUMNS[0].d/n241 ,
         \MIXCOLUMNS[0].d/n240 , \MIXCOLUMNS[0].d/n239 ,
         \MIXCOLUMNS[0].d/n238 , \MIXCOLUMNS[0].d/n237 ,
         \MIXCOLUMNS[0].d/n236 , \MIXCOLUMNS[0].d/n235 ,
         \MIXCOLUMNS[0].d/n234 , \MIXCOLUMNS[0].d/n233 ,
         \MIXCOLUMNS[0].d/n232 , \MIXCOLUMNS[0].d/n231 ,
         \MIXCOLUMNS[0].d/n230 , \MIXCOLUMNS[0].d/n229 ,
         \MIXCOLUMNS[0].d/n228 , \MIXCOLUMNS[0].d/n227 ,
         \MIXCOLUMNS[0].d/n226 , \MIXCOLUMNS[0].d/n225 ,
         \MIXCOLUMNS[0].d/n224 , \MIXCOLUMNS[0].d/n223 ,
         \MIXCOLUMNS[0].d/n222 , \MIXCOLUMNS[0].d/n221 ,
         \MIXCOLUMNS[0].d/n220 , \MIXCOLUMNS[0].d/n219 ,
         \MIXCOLUMNS[0].d/n218 , \MIXCOLUMNS[0].d/n217 ,
         \MIXCOLUMNS[0].d/n216 , \MIXCOLUMNS[0].d/n215 ,
         \MIXCOLUMNS[0].d/n214 , \MIXCOLUMNS[0].d/n213 ,
         \MIXCOLUMNS[0].d/n212 , \MIXCOLUMNS[0].d/n211 ,
         \MIXCOLUMNS[0].d/n210 , \MIXCOLUMNS[0].d/n209 ,
         \MIXCOLUMNS[0].d/n208 , \MIXCOLUMNS[0].d/n207 ,
         \MIXCOLUMNS[0].d/n206 , \MIXCOLUMNS[0].d/n205 ,
         \MIXCOLUMNS[0].d/n204 , \MIXCOLUMNS[0].d/n203 ,
         \MIXCOLUMNS[0].d/n202 , \MIXCOLUMNS[0].d/n201 ,
         \MIXCOLUMNS[0].d/n200 , \MIXCOLUMNS[0].d/n199 ,
         \MIXCOLUMNS[0].d/n198 , \MIXCOLUMNS[0].d/n197 ,
         \MIXCOLUMNS[0].d/n196 , \MIXCOLUMNS[0].d/n195 ,
         \MIXCOLUMNS[0].d/n194 , \MIXCOLUMNS[0].d/n193 ,
         \MIXCOLUMNS[0].d/n192 , \MIXCOLUMNS[0].d/n191 ,
         \MIXCOLUMNS[0].d/n190 , \MIXCOLUMNS[0].d/n189 ,
         \MIXCOLUMNS[0].d/n188 , \MIXCOLUMNS[0].d/n187 ,
         \MIXCOLUMNS[0].d/n186 , \MIXCOLUMNS[0].d/n185 ,
         \MIXCOLUMNS[0].d/n184 , \MIXCOLUMNS[0].d/n183 ,
         \MIXCOLUMNS[0].d/n182 , \MIXCOLUMNS[0].d/n181 ,
         \MIXCOLUMNS[0].d/n180 , \MIXCOLUMNS[0].d/n179 ,
         \MIXCOLUMNS[0].d/n178 , \MIXCOLUMNS[0].d/n177 ,
         \MIXCOLUMNS[0].d/n176 , \MIXCOLUMNS[0].d/n175 ,
         \MIXCOLUMNS[0].d/n174 , \MIXCOLUMNS[0].d/n173 ,
         \MIXCOLUMNS[0].d/n172 , \MIXCOLUMNS[0].d/n171 ,
         \MIXCOLUMNS[0].d/n170 , \MIXCOLUMNS[0].d/n169 ,
         \MIXCOLUMNS[0].d/n168 , \MIXCOLUMNS[0].d/n167 ,
         \MIXCOLUMNS[0].d/n166 , \MIXCOLUMNS[0].d/n165 ,
         \MIXCOLUMNS[0].d/n164 , \MIXCOLUMNS[0].d/n163 ,
         \MIXCOLUMNS[0].d/n162 , \MIXCOLUMNS[0].d/n161 ,
         \MIXCOLUMNS[0].d/n160 , \MIXCOLUMNS[0].d/n159 ,
         \MIXCOLUMNS[0].d/n158 , \MIXCOLUMNS[0].d/n157 ,
         \MIXCOLUMNS[0].d/n156 , \MIXCOLUMNS[0].d/n155 ,
         \MIXCOLUMNS[0].d/n154 , \MIXCOLUMNS[0].d/n153 ,
         \MIXCOLUMNS[0].d/n152 , \MIXCOLUMNS[0].d/n151 ,
         \MIXCOLUMNS[0].d/n150 , \MIXCOLUMNS[0].d/n149 ,
         \MIXCOLUMNS[0].d/n148 , \MIXCOLUMNS[0].d/n147 ,
         \MIXCOLUMNS[0].d/n146 , \MIXCOLUMNS[0].d/n145 ,
         \MIXCOLUMNS[0].d/n144 , \MIXCOLUMNS[0].d/n143 ,
         \MIXCOLUMNS[0].d/n142 , \MIXCOLUMNS[0].d/n141 ,
         \MIXCOLUMNS[0].d/n140 , \MIXCOLUMNS[0].d/n139 ,
         \MIXCOLUMNS[0].d/n138 , \MIXCOLUMNS[0].d/n137 ,
         \MIXCOLUMNS[0].d/n136 , \MIXCOLUMNS[0].d/n135 ,
         \MIXCOLUMNS[0].d/n134 , \MIXCOLUMNS[0].d/n133 ,
         \MIXCOLUMNS[0].d/n132 , \MIXCOLUMNS[0].d/n131 ,
         \MIXCOLUMNS[0].d/n130 , \MIXCOLUMNS[0].d/n129 ,
         \MIXCOLUMNS[0].d/n128 , \MIXCOLUMNS[0].d/n127 ,
         \MIXCOLUMNS[0].d/n126 , \MIXCOLUMNS[0].d/n125 ,
         \MIXCOLUMNS[0].d/n124 , \MIXCOLUMNS[0].d/n123 ,
         \MIXCOLUMNS[0].d/n122 , \MIXCOLUMNS[0].d/n121 ,
         \MIXCOLUMNS[0].d/n120 , \MIXCOLUMNS[0].d/n119 ,
         \MIXCOLUMNS[0].d/n118 , \MIXCOLUMNS[0].d/n117 ,
         \MIXCOLUMNS[0].d/n116 , \MIXCOLUMNS[0].d/n115 ,
         \MIXCOLUMNS[0].d/n114 , \MIXCOLUMNS[0].d/n113 ,
         \MIXCOLUMNS[0].d/n112 , \MIXCOLUMNS[0].d/n111 ,
         \MIXCOLUMNS[0].d/n110 , \MIXCOLUMNS[0].d/n109 ,
         \MIXCOLUMNS[0].d/n108 , \MIXCOLUMNS[0].d/n107 ,
         \MIXCOLUMNS[0].d/n106 , \MIXCOLUMNS[0].d/n105 ,
         \MIXCOLUMNS[0].d/n104 , \MIXCOLUMNS[0].d/n103 ,
         \MIXCOLUMNS[0].d/n102 , \MIXCOLUMNS[0].d/n101 ,
         \MIXCOLUMNS[0].d/n100 , \MIXCOLUMNS[0].d/n99 , \MIXCOLUMNS[0].d/n98 ,
         \MIXCOLUMNS[0].d/n97 , \MIXCOLUMNS[0].d/n96 , \MIXCOLUMNS[0].d/n95 ,
         \MIXCOLUMNS[0].d/n94 , \MIXCOLUMNS[0].d/n93 , \MIXCOLUMNS[0].d/n92 ,
         \MIXCOLUMNS[0].d/n91 , \MIXCOLUMNS[0].d/n90 , \MIXCOLUMNS[0].d/n89 ,
         \MIXCOLUMNS[0].d/n88 , \MIXCOLUMNS[0].d/n87 , \MIXCOLUMNS[0].d/n86 ,
         \MIXCOLUMNS[0].d/n85 , \MIXCOLUMNS[0].d/n84 , \MIXCOLUMNS[0].d/n83 ,
         \MIXCOLUMNS[0].d/n82 , \MIXCOLUMNS[0].d/n81 , \MIXCOLUMNS[0].d/n80 ,
         \MIXCOLUMNS[0].d/n79 , \MIXCOLUMNS[0].d/n78 , \MIXCOLUMNS[0].d/n77 ,
         \MIXCOLUMNS[0].d/n76 , \MIXCOLUMNS[0].d/n75 , \MIXCOLUMNS[0].d/n74 ,
         \MIXCOLUMNS[0].d/n73 , \MIXCOLUMNS[0].d/n72 , \MIXCOLUMNS[0].d/n71 ,
         \MIXCOLUMNS[0].d/n70 , \MIXCOLUMNS[0].d/n69 , \MIXCOLUMNS[0].d/n68 ,
         \MIXCOLUMNS[0].d/n67 , \MIXCOLUMNS[0].d/n66 , \MIXCOLUMNS[0].d/n65 ,
         \MIXCOLUMNS[0].d/n64 , \MIXCOLUMNS[0].d/n63 , \MIXCOLUMNS[0].d/n62 ,
         \MIXCOLUMNS[0].d/n61 , \MIXCOLUMNS[0].d/n60 , \MIXCOLUMNS[0].d/n59 ,
         \MIXCOLUMNS[0].d/n58 , \MIXCOLUMNS[0].d/n57 , \MIXCOLUMNS[0].d/n56 ,
         \MIXCOLUMNS[0].d/n55 , \MIXCOLUMNS[0].d/n54 , \MIXCOLUMNS[0].d/n53 ,
         \MIXCOLUMNS[0].d/n52 , \MIXCOLUMNS[0].d/n51 , \MIXCOLUMNS[0].d/n50 ,
         \MIXCOLUMNS[0].d/n49 , \MIXCOLUMNS[0].d/n48 , \MIXCOLUMNS[0].d/n47 ,
         \MIXCOLUMNS[0].d/n46 , \MIXCOLUMNS[0].d/n45 , \MIXCOLUMNS[0].d/n44 ,
         \MIXCOLUMNS[0].d/n43 , \MIXCOLUMNS[0].d/n42 , \MIXCOLUMNS[0].d/n41 ,
         \MIXCOLUMNS[0].d/n40 , \MIXCOLUMNS[0].d/n39 , \MIXCOLUMNS[0].d/n38 ,
         \MIXCOLUMNS[0].d/n37 , \MIXCOLUMNS[0].d/n36 , \MIXCOLUMNS[0].d/n35 ,
         \MIXCOLUMNS[0].d/n34 , \MIXCOLUMNS[0].d/n33 , \MIXCOLUMNS[0].d/n32 ,
         \MIXCOLUMNS[0].d/n31 , \MIXCOLUMNS[0].d/n30 , \MIXCOLUMNS[0].d/n29 ,
         \MIXCOLUMNS[0].d/n28 , \MIXCOLUMNS[0].d/n27 , \MIXCOLUMNS[0].d/n26 ,
         \MIXCOLUMNS[0].d/n25 , \MIXCOLUMNS[0].d/n24 , \MIXCOLUMNS[0].d/n23 ,
         \MIXCOLUMNS[0].d/n22 , \MIXCOLUMNS[0].d/n21 , \MIXCOLUMNS[0].d/n20 ,
         \MIXCOLUMNS[0].d/n19 , \MIXCOLUMNS[0].d/n18 , \MIXCOLUMNS[0].d/n17 ,
         \MIXCOLUMNS[0].d/n16 , \MIXCOLUMNS[0].d/n15 , \MIXCOLUMNS[0].d/n14 ,
         \MIXCOLUMNS[0].d/n13 , \MIXCOLUMNS[0].d/n12 , \MIXCOLUMNS[0].d/n11 ,
         \MIXCOLUMNS[0].d/n10 , \MIXCOLUMNS[0].d/n9 , \MIXCOLUMNS[0].d/n8 ,
         \MIXCOLUMNS[0].d/n7 , \MIXCOLUMNS[0].d/n6 , \MIXCOLUMNS[0].d/n5 ,
         \MIXCOLUMNS[0].d/n4 , \MIXCOLUMNS[0].d/n3 , \MIXCOLUMNS[0].d/n2 ,
         \MIXCOLUMNS[0].d/n1 , \SUBBYTES[9].a/w3400 , \SUBBYTES[9].a/w3398 ,
         \SUBBYTES[9].a/w3397 , \SUBBYTES[9].a/w3396 , \SUBBYTES[9].a/w3393 ,
         \SUBBYTES[9].a/w3391 , \SUBBYTES[9].a/w3390 , \SUBBYTES[9].a/w3389 ,
         \SUBBYTES[9].a/w3385 , \SUBBYTES[9].a/w3383 , \SUBBYTES[9].a/w3382 ,
         \SUBBYTES[9].a/w3381 , \SUBBYTES[9].a/w3380 , \SUBBYTES[9].a/w3379 ,
         \SUBBYTES[9].a/w3378 , \SUBBYTES[9].a/w3377 , \SUBBYTES[9].a/w3376 ,
         \SUBBYTES[9].a/w3368 , \SUBBYTES[9].a/w3366 , \SUBBYTES[9].a/w3365 ,
         \SUBBYTES[9].a/w3361 , \SUBBYTES[9].a/w3359 , \SUBBYTES[9].a/w3358 ,
         \SUBBYTES[9].a/w3357 , \SUBBYTES[9].a/w3353 , \SUBBYTES[9].a/w3351 ,
         \SUBBYTES[9].a/w3350 , \SUBBYTES[9].a/w3337 , \SUBBYTES[9].a/w3336 ,
         \SUBBYTES[9].a/w3335 , \SUBBYTES[9].a/w3333 , \SUBBYTES[9].a/w3330 ,
         \SUBBYTES[9].a/w3329 , \SUBBYTES[9].a/w3327 , \SUBBYTES[9].a/w3326 ,
         \SUBBYTES[9].a/w3324 , \SUBBYTES[9].a/w3322 , \SUBBYTES[9].a/w3321 ,
         \SUBBYTES[9].a/w3315 , \SUBBYTES[9].a/w3314 , \SUBBYTES[9].a/w3313 ,
         \SUBBYTES[9].a/w3312 , \SUBBYTES[9].a/w3306 , \SUBBYTES[9].a/w3304 ,
         \SUBBYTES[9].a/w3303 , \SUBBYTES[9].a/w3299 , \SUBBYTES[9].a/w3297 ,
         \SUBBYTES[9].a/w3296 , \SUBBYTES[9].a/w3291 , \SUBBYTES[9].a/w3289 ,
         \SUBBYTES[9].a/w3288 , \SUBBYTES[9].a/w3272 , \SUBBYTES[9].a/w3271 ,
         \SUBBYTES[9].a/w3270 , \SUBBYTES[9].a/w3269 , \SUBBYTES[9].a/w3268 ,
         \SUBBYTES[9].a/w3266 , \SUBBYTES[9].a/w3265 , \SUBBYTES[9].a/w3193 ,
         \SUBBYTES[9].a/w3191 , \SUBBYTES[9].a/w3190 , \SUBBYTES[9].a/w3189 ,
         \SUBBYTES[9].a/w3186 , \SUBBYTES[9].a/w3184 , \SUBBYTES[9].a/w3183 ,
         \SUBBYTES[9].a/w3182 , \SUBBYTES[9].a/w3178 , \SUBBYTES[9].a/w3176 ,
         \SUBBYTES[9].a/w3175 , \SUBBYTES[9].a/w3174 , \SUBBYTES[9].a/w3173 ,
         \SUBBYTES[9].a/w3172 , \SUBBYTES[9].a/w3171 , \SUBBYTES[9].a/w3170 ,
         \SUBBYTES[9].a/w3169 , \SUBBYTES[9].a/w3161 , \SUBBYTES[9].a/w3159 ,
         \SUBBYTES[9].a/w3158 , \SUBBYTES[9].a/w3154 , \SUBBYTES[9].a/w3152 ,
         \SUBBYTES[9].a/w3151 , \SUBBYTES[9].a/w3150 , \SUBBYTES[9].a/w3146 ,
         \SUBBYTES[9].a/w3144 , \SUBBYTES[9].a/w3143 , \SUBBYTES[9].a/w3130 ,
         \SUBBYTES[9].a/w3129 , \SUBBYTES[9].a/w3128 , \SUBBYTES[9].a/w3126 ,
         \SUBBYTES[9].a/w3123 , \SUBBYTES[9].a/w3122 , \SUBBYTES[9].a/w3120 ,
         \SUBBYTES[9].a/w3119 , \SUBBYTES[9].a/w3117 , \SUBBYTES[9].a/w3115 ,
         \SUBBYTES[9].a/w3114 , \SUBBYTES[9].a/w3108 , \SUBBYTES[9].a/w3107 ,
         \SUBBYTES[9].a/w3106 , \SUBBYTES[9].a/w3105 , \SUBBYTES[9].a/w3099 ,
         \SUBBYTES[9].a/w3097 , \SUBBYTES[9].a/w3096 , \SUBBYTES[9].a/w3092 ,
         \SUBBYTES[9].a/w3090 , \SUBBYTES[9].a/w3089 , \SUBBYTES[9].a/w3084 ,
         \SUBBYTES[9].a/w3082 , \SUBBYTES[9].a/w3081 , \SUBBYTES[9].a/w3065 ,
         \SUBBYTES[9].a/w3064 , \SUBBYTES[9].a/w3063 , \SUBBYTES[9].a/w3062 ,
         \SUBBYTES[9].a/w3061 , \SUBBYTES[9].a/w3059 , \SUBBYTES[9].a/w3058 ,
         \SUBBYTES[9].a/w2986 , \SUBBYTES[9].a/w2984 , \SUBBYTES[9].a/w2983 ,
         \SUBBYTES[9].a/w2982 , \SUBBYTES[9].a/w2979 , \SUBBYTES[9].a/w2977 ,
         \SUBBYTES[9].a/w2976 , \SUBBYTES[9].a/w2975 , \SUBBYTES[9].a/w2971 ,
         \SUBBYTES[9].a/w2969 , \SUBBYTES[9].a/w2968 , \SUBBYTES[9].a/w2967 ,
         \SUBBYTES[9].a/w2966 , \SUBBYTES[9].a/w2965 , \SUBBYTES[9].a/w2964 ,
         \SUBBYTES[9].a/w2963 , \SUBBYTES[9].a/w2962 , \SUBBYTES[9].a/w2954 ,
         \SUBBYTES[9].a/w2952 , \SUBBYTES[9].a/w2951 , \SUBBYTES[9].a/w2947 ,
         \SUBBYTES[9].a/w2945 , \SUBBYTES[9].a/w2944 , \SUBBYTES[9].a/w2943 ,
         \SUBBYTES[9].a/w2939 , \SUBBYTES[9].a/w2937 , \SUBBYTES[9].a/w2936 ,
         \SUBBYTES[9].a/w2923 , \SUBBYTES[9].a/w2922 , \SUBBYTES[9].a/w2921 ,
         \SUBBYTES[9].a/w2919 , \SUBBYTES[9].a/w2916 , \SUBBYTES[9].a/w2915 ,
         \SUBBYTES[9].a/w2913 , \SUBBYTES[9].a/w2912 , \SUBBYTES[9].a/w2910 ,
         \SUBBYTES[9].a/w2908 , \SUBBYTES[9].a/w2907 , \SUBBYTES[9].a/w2901 ,
         \SUBBYTES[9].a/w2900 , \SUBBYTES[9].a/w2899 , \SUBBYTES[9].a/w2898 ,
         \SUBBYTES[9].a/w2892 , \SUBBYTES[9].a/w2890 , \SUBBYTES[9].a/w2889 ,
         \SUBBYTES[9].a/w2885 , \SUBBYTES[9].a/w2883 , \SUBBYTES[9].a/w2882 ,
         \SUBBYTES[9].a/w2877 , \SUBBYTES[9].a/w2875 , \SUBBYTES[9].a/w2874 ,
         \SUBBYTES[9].a/w2858 , \SUBBYTES[9].a/w2857 , \SUBBYTES[9].a/w2856 ,
         \SUBBYTES[9].a/w2855 , \SUBBYTES[9].a/w2854 , \SUBBYTES[9].a/w2852 ,
         \SUBBYTES[9].a/w2851 , \SUBBYTES[9].a/w2779 , \SUBBYTES[9].a/w2777 ,
         \SUBBYTES[9].a/w2776 , \SUBBYTES[9].a/w2775 , \SUBBYTES[9].a/w2772 ,
         \SUBBYTES[9].a/w2770 , \SUBBYTES[9].a/w2769 , \SUBBYTES[9].a/w2768 ,
         \SUBBYTES[9].a/w2764 , \SUBBYTES[9].a/w2762 , \SUBBYTES[9].a/w2761 ,
         \SUBBYTES[9].a/w2760 , \SUBBYTES[9].a/w2759 , \SUBBYTES[9].a/w2758 ,
         \SUBBYTES[9].a/w2757 , \SUBBYTES[9].a/w2756 , \SUBBYTES[9].a/w2755 ,
         \SUBBYTES[9].a/w2747 , \SUBBYTES[9].a/w2745 , \SUBBYTES[9].a/w2744 ,
         \SUBBYTES[9].a/w2740 , \SUBBYTES[9].a/w2738 , \SUBBYTES[9].a/w2737 ,
         \SUBBYTES[9].a/w2736 , \SUBBYTES[9].a/w2732 , \SUBBYTES[9].a/w2730 ,
         \SUBBYTES[9].a/w2729 , \SUBBYTES[9].a/w2716 , \SUBBYTES[9].a/w2715 ,
         \SUBBYTES[9].a/w2714 , \SUBBYTES[9].a/w2712 , \SUBBYTES[9].a/w2709 ,
         \SUBBYTES[9].a/w2708 , \SUBBYTES[9].a/w2706 , \SUBBYTES[9].a/w2705 ,
         \SUBBYTES[9].a/w2703 , \SUBBYTES[9].a/w2701 , \SUBBYTES[9].a/w2700 ,
         \SUBBYTES[9].a/w2694 , \SUBBYTES[9].a/w2693 , \SUBBYTES[9].a/w2692 ,
         \SUBBYTES[9].a/w2691 , \SUBBYTES[9].a/w2685 , \SUBBYTES[9].a/w2683 ,
         \SUBBYTES[9].a/w2682 , \SUBBYTES[9].a/w2678 , \SUBBYTES[9].a/w2676 ,
         \SUBBYTES[9].a/w2675 , \SUBBYTES[9].a/w2670 , \SUBBYTES[9].a/w2668 ,
         \SUBBYTES[9].a/w2667 , \SUBBYTES[9].a/w2651 , \SUBBYTES[9].a/w2650 ,
         \SUBBYTES[9].a/w2649 , \SUBBYTES[9].a/w2648 , \SUBBYTES[9].a/w2647 ,
         \SUBBYTES[9].a/w2645 , \SUBBYTES[9].a/w2644 , \SUBBYTES[9].a/w2572 ,
         \SUBBYTES[9].a/w2570 , \SUBBYTES[9].a/w2569 , \SUBBYTES[9].a/w2568 ,
         \SUBBYTES[9].a/w2565 , \SUBBYTES[9].a/w2563 , \SUBBYTES[9].a/w2562 ,
         \SUBBYTES[9].a/w2561 , \SUBBYTES[9].a/w2557 , \SUBBYTES[9].a/w2555 ,
         \SUBBYTES[9].a/w2554 , \SUBBYTES[9].a/w2553 , \SUBBYTES[9].a/w2552 ,
         \SUBBYTES[9].a/w2551 , \SUBBYTES[9].a/w2550 , \SUBBYTES[9].a/w2549 ,
         \SUBBYTES[9].a/w2548 , \SUBBYTES[9].a/w2540 , \SUBBYTES[9].a/w2538 ,
         \SUBBYTES[9].a/w2537 , \SUBBYTES[9].a/w2533 , \SUBBYTES[9].a/w2531 ,
         \SUBBYTES[9].a/w2530 , \SUBBYTES[9].a/w2529 , \SUBBYTES[9].a/w2525 ,
         \SUBBYTES[9].a/w2523 , \SUBBYTES[9].a/w2522 , \SUBBYTES[9].a/w2509 ,
         \SUBBYTES[9].a/w2508 , \SUBBYTES[9].a/w2507 , \SUBBYTES[9].a/w2505 ,
         \SUBBYTES[9].a/w2502 , \SUBBYTES[9].a/w2501 , \SUBBYTES[9].a/w2499 ,
         \SUBBYTES[9].a/w2498 , \SUBBYTES[9].a/w2496 , \SUBBYTES[9].a/w2494 ,
         \SUBBYTES[9].a/w2493 , \SUBBYTES[9].a/w2487 , \SUBBYTES[9].a/w2486 ,
         \SUBBYTES[9].a/w2485 , \SUBBYTES[9].a/w2484 , \SUBBYTES[9].a/w2478 ,
         \SUBBYTES[9].a/w2476 , \SUBBYTES[9].a/w2475 , \SUBBYTES[9].a/w2471 ,
         \SUBBYTES[9].a/w2469 , \SUBBYTES[9].a/w2468 , \SUBBYTES[9].a/w2463 ,
         \SUBBYTES[9].a/w2461 , \SUBBYTES[9].a/w2460 , \SUBBYTES[9].a/w2444 ,
         \SUBBYTES[9].a/w2443 , \SUBBYTES[9].a/w2442 , \SUBBYTES[9].a/w2441 ,
         \SUBBYTES[9].a/w2440 , \SUBBYTES[9].a/w2438 , \SUBBYTES[9].a/w2437 ,
         \SUBBYTES[9].a/w2365 , \SUBBYTES[9].a/w2363 , \SUBBYTES[9].a/w2362 ,
         \SUBBYTES[9].a/w2361 , \SUBBYTES[9].a/w2358 , \SUBBYTES[9].a/w2356 ,
         \SUBBYTES[9].a/w2355 , \SUBBYTES[9].a/w2354 , \SUBBYTES[9].a/w2350 ,
         \SUBBYTES[9].a/w2348 , \SUBBYTES[9].a/w2347 , \SUBBYTES[9].a/w2346 ,
         \SUBBYTES[9].a/w2345 , \SUBBYTES[9].a/w2344 , \SUBBYTES[9].a/w2343 ,
         \SUBBYTES[9].a/w2342 , \SUBBYTES[9].a/w2341 , \SUBBYTES[9].a/w2333 ,
         \SUBBYTES[9].a/w2331 , \SUBBYTES[9].a/w2330 , \SUBBYTES[9].a/w2326 ,
         \SUBBYTES[9].a/w2324 , \SUBBYTES[9].a/w2323 , \SUBBYTES[9].a/w2322 ,
         \SUBBYTES[9].a/w2318 , \SUBBYTES[9].a/w2316 , \SUBBYTES[9].a/w2315 ,
         \SUBBYTES[9].a/w2302 , \SUBBYTES[9].a/w2301 , \SUBBYTES[9].a/w2300 ,
         \SUBBYTES[9].a/w2298 , \SUBBYTES[9].a/w2295 , \SUBBYTES[9].a/w2294 ,
         \SUBBYTES[9].a/w2292 , \SUBBYTES[9].a/w2291 , \SUBBYTES[9].a/w2289 ,
         \SUBBYTES[9].a/w2287 , \SUBBYTES[9].a/w2286 , \SUBBYTES[9].a/w2280 ,
         \SUBBYTES[9].a/w2279 , \SUBBYTES[9].a/w2278 , \SUBBYTES[9].a/w2277 ,
         \SUBBYTES[9].a/w2271 , \SUBBYTES[9].a/w2269 , \SUBBYTES[9].a/w2268 ,
         \SUBBYTES[9].a/w2264 , \SUBBYTES[9].a/w2262 , \SUBBYTES[9].a/w2261 ,
         \SUBBYTES[9].a/w2256 , \SUBBYTES[9].a/w2254 , \SUBBYTES[9].a/w2253 ,
         \SUBBYTES[9].a/w2237 , \SUBBYTES[9].a/w2236 , \SUBBYTES[9].a/w2235 ,
         \SUBBYTES[9].a/w2234 , \SUBBYTES[9].a/w2233 , \SUBBYTES[9].a/w2231 ,
         \SUBBYTES[9].a/w2230 , \SUBBYTES[9].a/w2158 , \SUBBYTES[9].a/w2156 ,
         \SUBBYTES[9].a/w2155 , \SUBBYTES[9].a/w2154 , \SUBBYTES[9].a/w2151 ,
         \SUBBYTES[9].a/w2149 , \SUBBYTES[9].a/w2148 , \SUBBYTES[9].a/w2147 ,
         \SUBBYTES[9].a/w2143 , \SUBBYTES[9].a/w2141 , \SUBBYTES[9].a/w2140 ,
         \SUBBYTES[9].a/w2139 , \SUBBYTES[9].a/w2138 , \SUBBYTES[9].a/w2137 ,
         \SUBBYTES[9].a/w2136 , \SUBBYTES[9].a/w2135 , \SUBBYTES[9].a/w2134 ,
         \SUBBYTES[9].a/w2126 , \SUBBYTES[9].a/w2124 , \SUBBYTES[9].a/w2123 ,
         \SUBBYTES[9].a/w2119 , \SUBBYTES[9].a/w2117 , \SUBBYTES[9].a/w2116 ,
         \SUBBYTES[9].a/w2115 , \SUBBYTES[9].a/w2111 , \SUBBYTES[9].a/w2109 ,
         \SUBBYTES[9].a/w2108 , \SUBBYTES[9].a/w2095 , \SUBBYTES[9].a/w2094 ,
         \SUBBYTES[9].a/w2093 , \SUBBYTES[9].a/w2091 , \SUBBYTES[9].a/w2088 ,
         \SUBBYTES[9].a/w2087 , \SUBBYTES[9].a/w2085 , \SUBBYTES[9].a/w2084 ,
         \SUBBYTES[9].a/w2082 , \SUBBYTES[9].a/w2080 , \SUBBYTES[9].a/w2079 ,
         \SUBBYTES[9].a/w2073 , \SUBBYTES[9].a/w2072 , \SUBBYTES[9].a/w2071 ,
         \SUBBYTES[9].a/w2070 , \SUBBYTES[9].a/w2064 , \SUBBYTES[9].a/w2062 ,
         \SUBBYTES[9].a/w2061 , \SUBBYTES[9].a/w2057 , \SUBBYTES[9].a/w2055 ,
         \SUBBYTES[9].a/w2054 , \SUBBYTES[9].a/w2049 , \SUBBYTES[9].a/w2047 ,
         \SUBBYTES[9].a/w2046 , \SUBBYTES[9].a/w2030 , \SUBBYTES[9].a/w2029 ,
         \SUBBYTES[9].a/w2028 , \SUBBYTES[9].a/w2027 , \SUBBYTES[9].a/w2026 ,
         \SUBBYTES[9].a/w2024 , \SUBBYTES[9].a/w2023 , \SUBBYTES[9].a/w1951 ,
         \SUBBYTES[9].a/w1949 , \SUBBYTES[9].a/w1948 , \SUBBYTES[9].a/w1947 ,
         \SUBBYTES[9].a/w1944 , \SUBBYTES[9].a/w1942 , \SUBBYTES[9].a/w1941 ,
         \SUBBYTES[9].a/w1940 , \SUBBYTES[9].a/w1936 , \SUBBYTES[9].a/w1934 ,
         \SUBBYTES[9].a/w1933 , \SUBBYTES[9].a/w1932 , \SUBBYTES[9].a/w1931 ,
         \SUBBYTES[9].a/w1930 , \SUBBYTES[9].a/w1929 , \SUBBYTES[9].a/w1928 ,
         \SUBBYTES[9].a/w1927 , \SUBBYTES[9].a/w1919 , \SUBBYTES[9].a/w1917 ,
         \SUBBYTES[9].a/w1916 , \SUBBYTES[9].a/w1912 , \SUBBYTES[9].a/w1910 ,
         \SUBBYTES[9].a/w1909 , \SUBBYTES[9].a/w1908 , \SUBBYTES[9].a/w1904 ,
         \SUBBYTES[9].a/w1902 , \SUBBYTES[9].a/w1901 , \SUBBYTES[9].a/w1888 ,
         \SUBBYTES[9].a/w1887 , \SUBBYTES[9].a/w1886 , \SUBBYTES[9].a/w1884 ,
         \SUBBYTES[9].a/w1881 , \SUBBYTES[9].a/w1880 , \SUBBYTES[9].a/w1878 ,
         \SUBBYTES[9].a/w1877 , \SUBBYTES[9].a/w1875 , \SUBBYTES[9].a/w1873 ,
         \SUBBYTES[9].a/w1872 , \SUBBYTES[9].a/w1866 , \SUBBYTES[9].a/w1865 ,
         \SUBBYTES[9].a/w1864 , \SUBBYTES[9].a/w1863 , \SUBBYTES[9].a/w1857 ,
         \SUBBYTES[9].a/w1855 , \SUBBYTES[9].a/w1854 , \SUBBYTES[9].a/w1850 ,
         \SUBBYTES[9].a/w1848 , \SUBBYTES[9].a/w1847 , \SUBBYTES[9].a/w1842 ,
         \SUBBYTES[9].a/w1840 , \SUBBYTES[9].a/w1839 , \SUBBYTES[9].a/w1823 ,
         \SUBBYTES[9].a/w1822 , \SUBBYTES[9].a/w1821 , \SUBBYTES[9].a/w1820 ,
         \SUBBYTES[9].a/w1819 , \SUBBYTES[9].a/w1817 , \SUBBYTES[9].a/w1816 ,
         \SUBBYTES[9].a/w1744 , \SUBBYTES[9].a/w1742 , \SUBBYTES[9].a/w1741 ,
         \SUBBYTES[9].a/w1740 , \SUBBYTES[9].a/w1737 , \SUBBYTES[9].a/w1735 ,
         \SUBBYTES[9].a/w1734 , \SUBBYTES[9].a/w1733 , \SUBBYTES[9].a/w1729 ,
         \SUBBYTES[9].a/w1727 , \SUBBYTES[9].a/w1726 , \SUBBYTES[9].a/w1725 ,
         \SUBBYTES[9].a/w1724 , \SUBBYTES[9].a/w1723 , \SUBBYTES[9].a/w1722 ,
         \SUBBYTES[9].a/w1721 , \SUBBYTES[9].a/w1720 , \SUBBYTES[9].a/w1712 ,
         \SUBBYTES[9].a/w1710 , \SUBBYTES[9].a/w1709 , \SUBBYTES[9].a/w1705 ,
         \SUBBYTES[9].a/w1703 , \SUBBYTES[9].a/w1702 , \SUBBYTES[9].a/w1701 ,
         \SUBBYTES[9].a/w1697 , \SUBBYTES[9].a/w1695 , \SUBBYTES[9].a/w1694 ,
         \SUBBYTES[9].a/w1681 , \SUBBYTES[9].a/w1680 , \SUBBYTES[9].a/w1679 ,
         \SUBBYTES[9].a/w1677 , \SUBBYTES[9].a/w1674 , \SUBBYTES[9].a/w1673 ,
         \SUBBYTES[9].a/w1671 , \SUBBYTES[9].a/w1670 , \SUBBYTES[9].a/w1668 ,
         \SUBBYTES[9].a/w1666 , \SUBBYTES[9].a/w1665 , \SUBBYTES[9].a/w1659 ,
         \SUBBYTES[9].a/w1658 , \SUBBYTES[9].a/w1657 , \SUBBYTES[9].a/w1656 ,
         \SUBBYTES[9].a/w1650 , \SUBBYTES[9].a/w1648 , \SUBBYTES[9].a/w1647 ,
         \SUBBYTES[9].a/w1643 , \SUBBYTES[9].a/w1641 , \SUBBYTES[9].a/w1640 ,
         \SUBBYTES[9].a/w1635 , \SUBBYTES[9].a/w1633 , \SUBBYTES[9].a/w1632 ,
         \SUBBYTES[9].a/w1616 , \SUBBYTES[9].a/w1615 , \SUBBYTES[9].a/w1614 ,
         \SUBBYTES[9].a/w1613 , \SUBBYTES[9].a/w1612 , \SUBBYTES[9].a/w1610 ,
         \SUBBYTES[9].a/w1609 , \SUBBYTES[9].a/w1537 , \SUBBYTES[9].a/w1535 ,
         \SUBBYTES[9].a/w1534 , \SUBBYTES[9].a/w1533 , \SUBBYTES[9].a/w1530 ,
         \SUBBYTES[9].a/w1528 , \SUBBYTES[9].a/w1527 , \SUBBYTES[9].a/w1526 ,
         \SUBBYTES[9].a/w1522 , \SUBBYTES[9].a/w1520 , \SUBBYTES[9].a/w1519 ,
         \SUBBYTES[9].a/w1518 , \SUBBYTES[9].a/w1517 , \SUBBYTES[9].a/w1516 ,
         \SUBBYTES[9].a/w1515 , \SUBBYTES[9].a/w1514 , \SUBBYTES[9].a/w1513 ,
         \SUBBYTES[9].a/w1505 , \SUBBYTES[9].a/w1503 , \SUBBYTES[9].a/w1502 ,
         \SUBBYTES[9].a/w1498 , \SUBBYTES[9].a/w1496 , \SUBBYTES[9].a/w1495 ,
         \SUBBYTES[9].a/w1494 , \SUBBYTES[9].a/w1490 , \SUBBYTES[9].a/w1488 ,
         \SUBBYTES[9].a/w1487 , \SUBBYTES[9].a/w1474 , \SUBBYTES[9].a/w1473 ,
         \SUBBYTES[9].a/w1472 , \SUBBYTES[9].a/w1470 , \SUBBYTES[9].a/w1467 ,
         \SUBBYTES[9].a/w1466 , \SUBBYTES[9].a/w1464 , \SUBBYTES[9].a/w1463 ,
         \SUBBYTES[9].a/w1461 , \SUBBYTES[9].a/w1459 , \SUBBYTES[9].a/w1458 ,
         \SUBBYTES[9].a/w1452 , \SUBBYTES[9].a/w1451 , \SUBBYTES[9].a/w1450 ,
         \SUBBYTES[9].a/w1449 , \SUBBYTES[9].a/w1443 , \SUBBYTES[9].a/w1441 ,
         \SUBBYTES[9].a/w1440 , \SUBBYTES[9].a/w1436 , \SUBBYTES[9].a/w1434 ,
         \SUBBYTES[9].a/w1433 , \SUBBYTES[9].a/w1428 , \SUBBYTES[9].a/w1426 ,
         \SUBBYTES[9].a/w1425 , \SUBBYTES[9].a/w1409 , \SUBBYTES[9].a/w1408 ,
         \SUBBYTES[9].a/w1407 , \SUBBYTES[9].a/w1406 , \SUBBYTES[9].a/w1405 ,
         \SUBBYTES[9].a/w1403 , \SUBBYTES[9].a/w1402 , \SUBBYTES[9].a/w1330 ,
         \SUBBYTES[9].a/w1328 , \SUBBYTES[9].a/w1327 , \SUBBYTES[9].a/w1326 ,
         \SUBBYTES[9].a/w1323 , \SUBBYTES[9].a/w1321 , \SUBBYTES[9].a/w1320 ,
         \SUBBYTES[9].a/w1319 , \SUBBYTES[9].a/w1315 , \SUBBYTES[9].a/w1313 ,
         \SUBBYTES[9].a/w1312 , \SUBBYTES[9].a/w1311 , \SUBBYTES[9].a/w1310 ,
         \SUBBYTES[9].a/w1309 , \SUBBYTES[9].a/w1308 , \SUBBYTES[9].a/w1307 ,
         \SUBBYTES[9].a/w1306 , \SUBBYTES[9].a/w1298 , \SUBBYTES[9].a/w1296 ,
         \SUBBYTES[9].a/w1295 , \SUBBYTES[9].a/w1291 , \SUBBYTES[9].a/w1289 ,
         \SUBBYTES[9].a/w1288 , \SUBBYTES[9].a/w1287 , \SUBBYTES[9].a/w1283 ,
         \SUBBYTES[9].a/w1281 , \SUBBYTES[9].a/w1280 , \SUBBYTES[9].a/w1267 ,
         \SUBBYTES[9].a/w1266 , \SUBBYTES[9].a/w1265 , \SUBBYTES[9].a/w1263 ,
         \SUBBYTES[9].a/w1260 , \SUBBYTES[9].a/w1259 , \SUBBYTES[9].a/w1257 ,
         \SUBBYTES[9].a/w1256 , \SUBBYTES[9].a/w1254 , \SUBBYTES[9].a/w1252 ,
         \SUBBYTES[9].a/w1251 , \SUBBYTES[9].a/w1245 , \SUBBYTES[9].a/w1244 ,
         \SUBBYTES[9].a/w1243 , \SUBBYTES[9].a/w1242 , \SUBBYTES[9].a/w1236 ,
         \SUBBYTES[9].a/w1234 , \SUBBYTES[9].a/w1233 , \SUBBYTES[9].a/w1229 ,
         \SUBBYTES[9].a/w1227 , \SUBBYTES[9].a/w1226 , \SUBBYTES[9].a/w1221 ,
         \SUBBYTES[9].a/w1219 , \SUBBYTES[9].a/w1218 , \SUBBYTES[9].a/w1202 ,
         \SUBBYTES[9].a/w1201 , \SUBBYTES[9].a/w1200 , \SUBBYTES[9].a/w1199 ,
         \SUBBYTES[9].a/w1198 , \SUBBYTES[9].a/w1196 , \SUBBYTES[9].a/w1195 ,
         \SUBBYTES[9].a/w1123 , \SUBBYTES[9].a/w1121 , \SUBBYTES[9].a/w1120 ,
         \SUBBYTES[9].a/w1119 , \SUBBYTES[9].a/w1116 , \SUBBYTES[9].a/w1114 ,
         \SUBBYTES[9].a/w1113 , \SUBBYTES[9].a/w1112 , \SUBBYTES[9].a/w1108 ,
         \SUBBYTES[9].a/w1106 , \SUBBYTES[9].a/w1105 , \SUBBYTES[9].a/w1104 ,
         \SUBBYTES[9].a/w1103 , \SUBBYTES[9].a/w1102 , \SUBBYTES[9].a/w1101 ,
         \SUBBYTES[9].a/w1100 , \SUBBYTES[9].a/w1099 , \SUBBYTES[9].a/w1091 ,
         \SUBBYTES[9].a/w1089 , \SUBBYTES[9].a/w1088 , \SUBBYTES[9].a/w1084 ,
         \SUBBYTES[9].a/w1082 , \SUBBYTES[9].a/w1081 , \SUBBYTES[9].a/w1080 ,
         \SUBBYTES[9].a/w1076 , \SUBBYTES[9].a/w1074 , \SUBBYTES[9].a/w1073 ,
         \SUBBYTES[9].a/w1060 , \SUBBYTES[9].a/w1059 , \SUBBYTES[9].a/w1058 ,
         \SUBBYTES[9].a/w1056 , \SUBBYTES[9].a/w1053 , \SUBBYTES[9].a/w1052 ,
         \SUBBYTES[9].a/w1050 , \SUBBYTES[9].a/w1049 , \SUBBYTES[9].a/w1047 ,
         \SUBBYTES[9].a/w1045 , \SUBBYTES[9].a/w1044 , \SUBBYTES[9].a/w1038 ,
         \SUBBYTES[9].a/w1037 , \SUBBYTES[9].a/w1036 , \SUBBYTES[9].a/w1035 ,
         \SUBBYTES[9].a/w1029 , \SUBBYTES[9].a/w1027 , \SUBBYTES[9].a/w1026 ,
         \SUBBYTES[9].a/w1022 , \SUBBYTES[9].a/w1020 , \SUBBYTES[9].a/w1019 ,
         \SUBBYTES[9].a/w1014 , \SUBBYTES[9].a/w1012 , \SUBBYTES[9].a/w1011 ,
         \SUBBYTES[9].a/w995 , \SUBBYTES[9].a/w994 , \SUBBYTES[9].a/w993 ,
         \SUBBYTES[9].a/w992 , \SUBBYTES[9].a/w991 , \SUBBYTES[9].a/w989 ,
         \SUBBYTES[9].a/w988 , \SUBBYTES[9].a/w916 , \SUBBYTES[9].a/w914 ,
         \SUBBYTES[9].a/w913 , \SUBBYTES[9].a/w912 , \SUBBYTES[9].a/w909 ,
         \SUBBYTES[9].a/w907 , \SUBBYTES[9].a/w906 , \SUBBYTES[9].a/w905 ,
         \SUBBYTES[9].a/w901 , \SUBBYTES[9].a/w899 , \SUBBYTES[9].a/w898 ,
         \SUBBYTES[9].a/w897 , \SUBBYTES[9].a/w896 , \SUBBYTES[9].a/w895 ,
         \SUBBYTES[9].a/w894 , \SUBBYTES[9].a/w893 , \SUBBYTES[9].a/w892 ,
         \SUBBYTES[9].a/w884 , \SUBBYTES[9].a/w882 , \SUBBYTES[9].a/w881 ,
         \SUBBYTES[9].a/w877 , \SUBBYTES[9].a/w875 , \SUBBYTES[9].a/w874 ,
         \SUBBYTES[9].a/w873 , \SUBBYTES[9].a/w869 , \SUBBYTES[9].a/w867 ,
         \SUBBYTES[9].a/w866 , \SUBBYTES[9].a/w853 , \SUBBYTES[9].a/w852 ,
         \SUBBYTES[9].a/w851 , \SUBBYTES[9].a/w849 , \SUBBYTES[9].a/w846 ,
         \SUBBYTES[9].a/w845 , \SUBBYTES[9].a/w843 , \SUBBYTES[9].a/w842 ,
         \SUBBYTES[9].a/w840 , \SUBBYTES[9].a/w838 , \SUBBYTES[9].a/w837 ,
         \SUBBYTES[9].a/w831 , \SUBBYTES[9].a/w830 , \SUBBYTES[9].a/w829 ,
         \SUBBYTES[9].a/w828 , \SUBBYTES[9].a/w822 , \SUBBYTES[9].a/w820 ,
         \SUBBYTES[9].a/w819 , \SUBBYTES[9].a/w815 , \SUBBYTES[9].a/w813 ,
         \SUBBYTES[9].a/w812 , \SUBBYTES[9].a/w807 , \SUBBYTES[9].a/w805 ,
         \SUBBYTES[9].a/w804 , \SUBBYTES[9].a/w788 , \SUBBYTES[9].a/w787 ,
         \SUBBYTES[9].a/w786 , \SUBBYTES[9].a/w785 , \SUBBYTES[9].a/w784 ,
         \SUBBYTES[9].a/w782 , \SUBBYTES[9].a/w781 , \SUBBYTES[9].a/w709 ,
         \SUBBYTES[9].a/w707 , \SUBBYTES[9].a/w706 , \SUBBYTES[9].a/w705 ,
         \SUBBYTES[9].a/w702 , \SUBBYTES[9].a/w700 , \SUBBYTES[9].a/w699 ,
         \SUBBYTES[9].a/w698 , \SUBBYTES[9].a/w694 , \SUBBYTES[9].a/w692 ,
         \SUBBYTES[9].a/w691 , \SUBBYTES[9].a/w690 , \SUBBYTES[9].a/w689 ,
         \SUBBYTES[9].a/w688 , \SUBBYTES[9].a/w687 , \SUBBYTES[9].a/w686 ,
         \SUBBYTES[9].a/w685 , \SUBBYTES[9].a/w677 , \SUBBYTES[9].a/w675 ,
         \SUBBYTES[9].a/w674 , \SUBBYTES[9].a/w670 , \SUBBYTES[9].a/w668 ,
         \SUBBYTES[9].a/w667 , \SUBBYTES[9].a/w666 , \SUBBYTES[9].a/w662 ,
         \SUBBYTES[9].a/w660 , \SUBBYTES[9].a/w659 , \SUBBYTES[9].a/w646 ,
         \SUBBYTES[9].a/w645 , \SUBBYTES[9].a/w644 , \SUBBYTES[9].a/w642 ,
         \SUBBYTES[9].a/w639 , \SUBBYTES[9].a/w638 , \SUBBYTES[9].a/w636 ,
         \SUBBYTES[9].a/w635 , \SUBBYTES[9].a/w633 , \SUBBYTES[9].a/w631 ,
         \SUBBYTES[9].a/w630 , \SUBBYTES[9].a/w624 , \SUBBYTES[9].a/w623 ,
         \SUBBYTES[9].a/w622 , \SUBBYTES[9].a/w621 , \SUBBYTES[9].a/w615 ,
         \SUBBYTES[9].a/w613 , \SUBBYTES[9].a/w612 , \SUBBYTES[9].a/w608 ,
         \SUBBYTES[9].a/w606 , \SUBBYTES[9].a/w605 , \SUBBYTES[9].a/w600 ,
         \SUBBYTES[9].a/w598 , \SUBBYTES[9].a/w597 , \SUBBYTES[9].a/w581 ,
         \SUBBYTES[9].a/w580 , \SUBBYTES[9].a/w579 , \SUBBYTES[9].a/w578 ,
         \SUBBYTES[9].a/w577 , \SUBBYTES[9].a/w575 , \SUBBYTES[9].a/w574 ,
         \SUBBYTES[9].a/w502 , \SUBBYTES[9].a/w500 , \SUBBYTES[9].a/w499 ,
         \SUBBYTES[9].a/w498 , \SUBBYTES[9].a/w495 , \SUBBYTES[9].a/w493 ,
         \SUBBYTES[9].a/w492 , \SUBBYTES[9].a/w491 , \SUBBYTES[9].a/w487 ,
         \SUBBYTES[9].a/w485 , \SUBBYTES[9].a/w484 , \SUBBYTES[9].a/w483 ,
         \SUBBYTES[9].a/w482 , \SUBBYTES[9].a/w481 , \SUBBYTES[9].a/w480 ,
         \SUBBYTES[9].a/w479 , \SUBBYTES[9].a/w478 , \SUBBYTES[9].a/w470 ,
         \SUBBYTES[9].a/w468 , \SUBBYTES[9].a/w467 , \SUBBYTES[9].a/w463 ,
         \SUBBYTES[9].a/w461 , \SUBBYTES[9].a/w460 , \SUBBYTES[9].a/w459 ,
         \SUBBYTES[9].a/w455 , \SUBBYTES[9].a/w453 , \SUBBYTES[9].a/w452 ,
         \SUBBYTES[9].a/w439 , \SUBBYTES[9].a/w438 , \SUBBYTES[9].a/w437 ,
         \SUBBYTES[9].a/w435 , \SUBBYTES[9].a/w432 , \SUBBYTES[9].a/w431 ,
         \SUBBYTES[9].a/w429 , \SUBBYTES[9].a/w428 , \SUBBYTES[9].a/w426 ,
         \SUBBYTES[9].a/w424 , \SUBBYTES[9].a/w423 , \SUBBYTES[9].a/w417 ,
         \SUBBYTES[9].a/w416 , \SUBBYTES[9].a/w415 , \SUBBYTES[9].a/w414 ,
         \SUBBYTES[9].a/w408 , \SUBBYTES[9].a/w406 , \SUBBYTES[9].a/w405 ,
         \SUBBYTES[9].a/w401 , \SUBBYTES[9].a/w399 , \SUBBYTES[9].a/w398 ,
         \SUBBYTES[9].a/w393 , \SUBBYTES[9].a/w391 , \SUBBYTES[9].a/w390 ,
         \SUBBYTES[9].a/w374 , \SUBBYTES[9].a/w373 , \SUBBYTES[9].a/w372 ,
         \SUBBYTES[9].a/w371 , \SUBBYTES[9].a/w370 , \SUBBYTES[9].a/w368 ,
         \SUBBYTES[9].a/w367 , \SUBBYTES[9].a/w295 , \SUBBYTES[9].a/w293 ,
         \SUBBYTES[9].a/w292 , \SUBBYTES[9].a/w291 , \SUBBYTES[9].a/w288 ,
         \SUBBYTES[9].a/w286 , \SUBBYTES[9].a/w285 , \SUBBYTES[9].a/w284 ,
         \SUBBYTES[9].a/w280 , \SUBBYTES[9].a/w278 , \SUBBYTES[9].a/w277 ,
         \SUBBYTES[9].a/w276 , \SUBBYTES[9].a/w275 , \SUBBYTES[9].a/w274 ,
         \SUBBYTES[9].a/w273 , \SUBBYTES[9].a/w272 , \SUBBYTES[9].a/w271 ,
         \SUBBYTES[9].a/w263 , \SUBBYTES[9].a/w261 , \SUBBYTES[9].a/w260 ,
         \SUBBYTES[9].a/w256 , \SUBBYTES[9].a/w254 , \SUBBYTES[9].a/w253 ,
         \SUBBYTES[9].a/w252 , \SUBBYTES[9].a/w248 , \SUBBYTES[9].a/w246 ,
         \SUBBYTES[9].a/w245 , \SUBBYTES[9].a/w232 , \SUBBYTES[9].a/w231 ,
         \SUBBYTES[9].a/w230 , \SUBBYTES[9].a/w228 , \SUBBYTES[9].a/w225 ,
         \SUBBYTES[9].a/w224 , \SUBBYTES[9].a/w222 , \SUBBYTES[9].a/w221 ,
         \SUBBYTES[9].a/w219 , \SUBBYTES[9].a/w217 , \SUBBYTES[9].a/w216 ,
         \SUBBYTES[9].a/w210 , \SUBBYTES[9].a/w209 , \SUBBYTES[9].a/w208 ,
         \SUBBYTES[9].a/w207 , \SUBBYTES[9].a/w201 , \SUBBYTES[9].a/w199 ,
         \SUBBYTES[9].a/w198 , \SUBBYTES[9].a/w194 , \SUBBYTES[9].a/w192 ,
         \SUBBYTES[9].a/w191 , \SUBBYTES[9].a/w186 , \SUBBYTES[9].a/w184 ,
         \SUBBYTES[9].a/w183 , \SUBBYTES[9].a/w167 , \SUBBYTES[9].a/w166 ,
         \SUBBYTES[9].a/w165 , \SUBBYTES[9].a/w164 , \SUBBYTES[9].a/w163 ,
         \SUBBYTES[9].a/w161 , \SUBBYTES[9].a/w160 , \SUBBYTES[8].a/w3400 ,
         \SUBBYTES[8].a/w3398 , \SUBBYTES[8].a/w3397 , \SUBBYTES[8].a/w3396 ,
         \SUBBYTES[8].a/w3393 , \SUBBYTES[8].a/w3391 , \SUBBYTES[8].a/w3390 ,
         \SUBBYTES[8].a/w3389 , \SUBBYTES[8].a/w3385 , \SUBBYTES[8].a/w3383 ,
         \SUBBYTES[8].a/w3382 , \SUBBYTES[8].a/w3381 , \SUBBYTES[8].a/w3380 ,
         \SUBBYTES[8].a/w3379 , \SUBBYTES[8].a/w3378 , \SUBBYTES[8].a/w3377 ,
         \SUBBYTES[8].a/w3376 , \SUBBYTES[8].a/w3368 , \SUBBYTES[8].a/w3366 ,
         \SUBBYTES[8].a/w3365 , \SUBBYTES[8].a/w3361 , \SUBBYTES[8].a/w3359 ,
         \SUBBYTES[8].a/w3358 , \SUBBYTES[8].a/w3357 , \SUBBYTES[8].a/w3353 ,
         \SUBBYTES[8].a/w3351 , \SUBBYTES[8].a/w3350 , \SUBBYTES[8].a/w3337 ,
         \SUBBYTES[8].a/w3336 , \SUBBYTES[8].a/w3335 , \SUBBYTES[8].a/w3333 ,
         \SUBBYTES[8].a/w3330 , \SUBBYTES[8].a/w3329 , \SUBBYTES[8].a/w3327 ,
         \SUBBYTES[8].a/w3326 , \SUBBYTES[8].a/w3324 , \SUBBYTES[8].a/w3322 ,
         \SUBBYTES[8].a/w3321 , \SUBBYTES[8].a/w3315 , \SUBBYTES[8].a/w3314 ,
         \SUBBYTES[8].a/w3313 , \SUBBYTES[8].a/w3312 , \SUBBYTES[8].a/w3306 ,
         \SUBBYTES[8].a/w3304 , \SUBBYTES[8].a/w3303 , \SUBBYTES[8].a/w3299 ,
         \SUBBYTES[8].a/w3297 , \SUBBYTES[8].a/w3296 , \SUBBYTES[8].a/w3291 ,
         \SUBBYTES[8].a/w3289 , \SUBBYTES[8].a/w3288 , \SUBBYTES[8].a/w3272 ,
         \SUBBYTES[8].a/w3271 , \SUBBYTES[8].a/w3270 , \SUBBYTES[8].a/w3269 ,
         \SUBBYTES[8].a/w3268 , \SUBBYTES[8].a/w3266 , \SUBBYTES[8].a/w3265 ,
         \SUBBYTES[8].a/w3193 , \SUBBYTES[8].a/w3191 , \SUBBYTES[8].a/w3190 ,
         \SUBBYTES[8].a/w3189 , \SUBBYTES[8].a/w3186 , \SUBBYTES[8].a/w3184 ,
         \SUBBYTES[8].a/w3183 , \SUBBYTES[8].a/w3182 , \SUBBYTES[8].a/w3178 ,
         \SUBBYTES[8].a/w3176 , \SUBBYTES[8].a/w3175 , \SUBBYTES[8].a/w3174 ,
         \SUBBYTES[8].a/w3173 , \SUBBYTES[8].a/w3172 , \SUBBYTES[8].a/w3171 ,
         \SUBBYTES[8].a/w3170 , \SUBBYTES[8].a/w3169 , \SUBBYTES[8].a/w3161 ,
         \SUBBYTES[8].a/w3159 , \SUBBYTES[8].a/w3158 , \SUBBYTES[8].a/w3154 ,
         \SUBBYTES[8].a/w3152 , \SUBBYTES[8].a/w3151 , \SUBBYTES[8].a/w3150 ,
         \SUBBYTES[8].a/w3146 , \SUBBYTES[8].a/w3144 , \SUBBYTES[8].a/w3143 ,
         \SUBBYTES[8].a/w3130 , \SUBBYTES[8].a/w3129 , \SUBBYTES[8].a/w3128 ,
         \SUBBYTES[8].a/w3126 , \SUBBYTES[8].a/w3123 , \SUBBYTES[8].a/w3122 ,
         \SUBBYTES[8].a/w3120 , \SUBBYTES[8].a/w3119 , \SUBBYTES[8].a/w3117 ,
         \SUBBYTES[8].a/w3115 , \SUBBYTES[8].a/w3114 , \SUBBYTES[8].a/w3108 ,
         \SUBBYTES[8].a/w3107 , \SUBBYTES[8].a/w3106 , \SUBBYTES[8].a/w3105 ,
         \SUBBYTES[8].a/w3099 , \SUBBYTES[8].a/w3097 , \SUBBYTES[8].a/w3096 ,
         \SUBBYTES[8].a/w3092 , \SUBBYTES[8].a/w3090 , \SUBBYTES[8].a/w3089 ,
         \SUBBYTES[8].a/w3084 , \SUBBYTES[8].a/w3082 , \SUBBYTES[8].a/w3081 ,
         \SUBBYTES[8].a/w3065 , \SUBBYTES[8].a/w3064 , \SUBBYTES[8].a/w3063 ,
         \SUBBYTES[8].a/w3062 , \SUBBYTES[8].a/w3061 , \SUBBYTES[8].a/w3059 ,
         \SUBBYTES[8].a/w3058 , \SUBBYTES[8].a/w2986 , \SUBBYTES[8].a/w2984 ,
         \SUBBYTES[8].a/w2983 , \SUBBYTES[8].a/w2982 , \SUBBYTES[8].a/w2979 ,
         \SUBBYTES[8].a/w2977 , \SUBBYTES[8].a/w2976 , \SUBBYTES[8].a/w2975 ,
         \SUBBYTES[8].a/w2971 , \SUBBYTES[8].a/w2969 , \SUBBYTES[8].a/w2968 ,
         \SUBBYTES[8].a/w2967 , \SUBBYTES[8].a/w2966 , \SUBBYTES[8].a/w2965 ,
         \SUBBYTES[8].a/w2964 , \SUBBYTES[8].a/w2963 , \SUBBYTES[8].a/w2962 ,
         \SUBBYTES[8].a/w2954 , \SUBBYTES[8].a/w2952 , \SUBBYTES[8].a/w2951 ,
         \SUBBYTES[8].a/w2947 , \SUBBYTES[8].a/w2945 , \SUBBYTES[8].a/w2944 ,
         \SUBBYTES[8].a/w2943 , \SUBBYTES[8].a/w2939 , \SUBBYTES[8].a/w2937 ,
         \SUBBYTES[8].a/w2936 , \SUBBYTES[8].a/w2923 , \SUBBYTES[8].a/w2922 ,
         \SUBBYTES[8].a/w2921 , \SUBBYTES[8].a/w2919 , \SUBBYTES[8].a/w2916 ,
         \SUBBYTES[8].a/w2915 , \SUBBYTES[8].a/w2913 , \SUBBYTES[8].a/w2912 ,
         \SUBBYTES[8].a/w2910 , \SUBBYTES[8].a/w2908 , \SUBBYTES[8].a/w2907 ,
         \SUBBYTES[8].a/w2901 , \SUBBYTES[8].a/w2900 , \SUBBYTES[8].a/w2899 ,
         \SUBBYTES[8].a/w2898 , \SUBBYTES[8].a/w2892 , \SUBBYTES[8].a/w2890 ,
         \SUBBYTES[8].a/w2889 , \SUBBYTES[8].a/w2885 , \SUBBYTES[8].a/w2883 ,
         \SUBBYTES[8].a/w2882 , \SUBBYTES[8].a/w2877 , \SUBBYTES[8].a/w2875 ,
         \SUBBYTES[8].a/w2874 , \SUBBYTES[8].a/w2858 , \SUBBYTES[8].a/w2857 ,
         \SUBBYTES[8].a/w2856 , \SUBBYTES[8].a/w2855 , \SUBBYTES[8].a/w2854 ,
         \SUBBYTES[8].a/w2852 , \SUBBYTES[8].a/w2851 , \SUBBYTES[8].a/w2779 ,
         \SUBBYTES[8].a/w2777 , \SUBBYTES[8].a/w2776 , \SUBBYTES[8].a/w2775 ,
         \SUBBYTES[8].a/w2772 , \SUBBYTES[8].a/w2770 , \SUBBYTES[8].a/w2769 ,
         \SUBBYTES[8].a/w2768 , \SUBBYTES[8].a/w2764 , \SUBBYTES[8].a/w2762 ,
         \SUBBYTES[8].a/w2761 , \SUBBYTES[8].a/w2760 , \SUBBYTES[8].a/w2759 ,
         \SUBBYTES[8].a/w2758 , \SUBBYTES[8].a/w2757 , \SUBBYTES[8].a/w2756 ,
         \SUBBYTES[8].a/w2755 , \SUBBYTES[8].a/w2747 , \SUBBYTES[8].a/w2745 ,
         \SUBBYTES[8].a/w2744 , \SUBBYTES[8].a/w2740 , \SUBBYTES[8].a/w2738 ,
         \SUBBYTES[8].a/w2737 , \SUBBYTES[8].a/w2736 , \SUBBYTES[8].a/w2732 ,
         \SUBBYTES[8].a/w2730 , \SUBBYTES[8].a/w2729 , \SUBBYTES[8].a/w2716 ,
         \SUBBYTES[8].a/w2715 , \SUBBYTES[8].a/w2714 , \SUBBYTES[8].a/w2712 ,
         \SUBBYTES[8].a/w2709 , \SUBBYTES[8].a/w2708 , \SUBBYTES[8].a/w2706 ,
         \SUBBYTES[8].a/w2705 , \SUBBYTES[8].a/w2703 , \SUBBYTES[8].a/w2701 ,
         \SUBBYTES[8].a/w2700 , \SUBBYTES[8].a/w2694 , \SUBBYTES[8].a/w2693 ,
         \SUBBYTES[8].a/w2692 , \SUBBYTES[8].a/w2691 , \SUBBYTES[8].a/w2685 ,
         \SUBBYTES[8].a/w2683 , \SUBBYTES[8].a/w2682 , \SUBBYTES[8].a/w2678 ,
         \SUBBYTES[8].a/w2676 , \SUBBYTES[8].a/w2675 , \SUBBYTES[8].a/w2670 ,
         \SUBBYTES[8].a/w2668 , \SUBBYTES[8].a/w2667 , \SUBBYTES[8].a/w2651 ,
         \SUBBYTES[8].a/w2650 , \SUBBYTES[8].a/w2649 , \SUBBYTES[8].a/w2648 ,
         \SUBBYTES[8].a/w2647 , \SUBBYTES[8].a/w2645 , \SUBBYTES[8].a/w2644 ,
         \SUBBYTES[8].a/w2572 , \SUBBYTES[8].a/w2570 , \SUBBYTES[8].a/w2569 ,
         \SUBBYTES[8].a/w2568 , \SUBBYTES[8].a/w2565 , \SUBBYTES[8].a/w2563 ,
         \SUBBYTES[8].a/w2562 , \SUBBYTES[8].a/w2561 , \SUBBYTES[8].a/w2557 ,
         \SUBBYTES[8].a/w2555 , \SUBBYTES[8].a/w2554 , \SUBBYTES[8].a/w2553 ,
         \SUBBYTES[8].a/w2552 , \SUBBYTES[8].a/w2551 , \SUBBYTES[8].a/w2550 ,
         \SUBBYTES[8].a/w2549 , \SUBBYTES[8].a/w2548 , \SUBBYTES[8].a/w2540 ,
         \SUBBYTES[8].a/w2538 , \SUBBYTES[8].a/w2537 , \SUBBYTES[8].a/w2533 ,
         \SUBBYTES[8].a/w2531 , \SUBBYTES[8].a/w2530 , \SUBBYTES[8].a/w2529 ,
         \SUBBYTES[8].a/w2525 , \SUBBYTES[8].a/w2523 , \SUBBYTES[8].a/w2522 ,
         \SUBBYTES[8].a/w2509 , \SUBBYTES[8].a/w2508 , \SUBBYTES[8].a/w2507 ,
         \SUBBYTES[8].a/w2505 , \SUBBYTES[8].a/w2502 , \SUBBYTES[8].a/w2501 ,
         \SUBBYTES[8].a/w2499 , \SUBBYTES[8].a/w2498 , \SUBBYTES[8].a/w2496 ,
         \SUBBYTES[8].a/w2494 , \SUBBYTES[8].a/w2493 , \SUBBYTES[8].a/w2487 ,
         \SUBBYTES[8].a/w2486 , \SUBBYTES[8].a/w2485 , \SUBBYTES[8].a/w2484 ,
         \SUBBYTES[8].a/w2478 , \SUBBYTES[8].a/w2476 , \SUBBYTES[8].a/w2475 ,
         \SUBBYTES[8].a/w2471 , \SUBBYTES[8].a/w2469 , \SUBBYTES[8].a/w2468 ,
         \SUBBYTES[8].a/w2463 , \SUBBYTES[8].a/w2461 , \SUBBYTES[8].a/w2460 ,
         \SUBBYTES[8].a/w2444 , \SUBBYTES[8].a/w2443 , \SUBBYTES[8].a/w2442 ,
         \SUBBYTES[8].a/w2441 , \SUBBYTES[8].a/w2440 , \SUBBYTES[8].a/w2438 ,
         \SUBBYTES[8].a/w2437 , \SUBBYTES[8].a/w2365 , \SUBBYTES[8].a/w2363 ,
         \SUBBYTES[8].a/w2362 , \SUBBYTES[8].a/w2361 , \SUBBYTES[8].a/w2358 ,
         \SUBBYTES[8].a/w2356 , \SUBBYTES[8].a/w2355 , \SUBBYTES[8].a/w2354 ,
         \SUBBYTES[8].a/w2350 , \SUBBYTES[8].a/w2348 , \SUBBYTES[8].a/w2347 ,
         \SUBBYTES[8].a/w2346 , \SUBBYTES[8].a/w2345 , \SUBBYTES[8].a/w2344 ,
         \SUBBYTES[8].a/w2343 , \SUBBYTES[8].a/w2342 , \SUBBYTES[8].a/w2341 ,
         \SUBBYTES[8].a/w2333 , \SUBBYTES[8].a/w2331 , \SUBBYTES[8].a/w2330 ,
         \SUBBYTES[8].a/w2326 , \SUBBYTES[8].a/w2324 , \SUBBYTES[8].a/w2323 ,
         \SUBBYTES[8].a/w2322 , \SUBBYTES[8].a/w2318 , \SUBBYTES[8].a/w2316 ,
         \SUBBYTES[8].a/w2315 , \SUBBYTES[8].a/w2302 , \SUBBYTES[8].a/w2301 ,
         \SUBBYTES[8].a/w2300 , \SUBBYTES[8].a/w2298 , \SUBBYTES[8].a/w2295 ,
         \SUBBYTES[8].a/w2294 , \SUBBYTES[8].a/w2292 , \SUBBYTES[8].a/w2291 ,
         \SUBBYTES[8].a/w2289 , \SUBBYTES[8].a/w2287 , \SUBBYTES[8].a/w2286 ,
         \SUBBYTES[8].a/w2280 , \SUBBYTES[8].a/w2279 , \SUBBYTES[8].a/w2278 ,
         \SUBBYTES[8].a/w2277 , \SUBBYTES[8].a/w2271 , \SUBBYTES[8].a/w2269 ,
         \SUBBYTES[8].a/w2268 , \SUBBYTES[8].a/w2264 , \SUBBYTES[8].a/w2262 ,
         \SUBBYTES[8].a/w2261 , \SUBBYTES[8].a/w2256 , \SUBBYTES[8].a/w2254 ,
         \SUBBYTES[8].a/w2253 , \SUBBYTES[8].a/w2237 , \SUBBYTES[8].a/w2236 ,
         \SUBBYTES[8].a/w2235 , \SUBBYTES[8].a/w2234 , \SUBBYTES[8].a/w2233 ,
         \SUBBYTES[8].a/w2231 , \SUBBYTES[8].a/w2230 , \SUBBYTES[8].a/w2158 ,
         \SUBBYTES[8].a/w2156 , \SUBBYTES[8].a/w2155 , \SUBBYTES[8].a/w2154 ,
         \SUBBYTES[8].a/w2151 , \SUBBYTES[8].a/w2149 , \SUBBYTES[8].a/w2148 ,
         \SUBBYTES[8].a/w2147 , \SUBBYTES[8].a/w2143 , \SUBBYTES[8].a/w2141 ,
         \SUBBYTES[8].a/w2140 , \SUBBYTES[8].a/w2139 , \SUBBYTES[8].a/w2138 ,
         \SUBBYTES[8].a/w2137 , \SUBBYTES[8].a/w2136 , \SUBBYTES[8].a/w2135 ,
         \SUBBYTES[8].a/w2134 , \SUBBYTES[8].a/w2126 , \SUBBYTES[8].a/w2124 ,
         \SUBBYTES[8].a/w2123 , \SUBBYTES[8].a/w2119 , \SUBBYTES[8].a/w2117 ,
         \SUBBYTES[8].a/w2116 , \SUBBYTES[8].a/w2115 , \SUBBYTES[8].a/w2111 ,
         \SUBBYTES[8].a/w2109 , \SUBBYTES[8].a/w2108 , \SUBBYTES[8].a/w2095 ,
         \SUBBYTES[8].a/w2094 , \SUBBYTES[8].a/w2093 , \SUBBYTES[8].a/w2091 ,
         \SUBBYTES[8].a/w2088 , \SUBBYTES[8].a/w2087 , \SUBBYTES[8].a/w2085 ,
         \SUBBYTES[8].a/w2084 , \SUBBYTES[8].a/w2082 , \SUBBYTES[8].a/w2080 ,
         \SUBBYTES[8].a/w2079 , \SUBBYTES[8].a/w2073 , \SUBBYTES[8].a/w2072 ,
         \SUBBYTES[8].a/w2071 , \SUBBYTES[8].a/w2070 , \SUBBYTES[8].a/w2064 ,
         \SUBBYTES[8].a/w2062 , \SUBBYTES[8].a/w2061 , \SUBBYTES[8].a/w2057 ,
         \SUBBYTES[8].a/w2055 , \SUBBYTES[8].a/w2054 , \SUBBYTES[8].a/w2049 ,
         \SUBBYTES[8].a/w2047 , \SUBBYTES[8].a/w2046 , \SUBBYTES[8].a/w2030 ,
         \SUBBYTES[8].a/w2029 , \SUBBYTES[8].a/w2028 , \SUBBYTES[8].a/w2027 ,
         \SUBBYTES[8].a/w2026 , \SUBBYTES[8].a/w2024 , \SUBBYTES[8].a/w2023 ,
         \SUBBYTES[8].a/w1951 , \SUBBYTES[8].a/w1949 , \SUBBYTES[8].a/w1948 ,
         \SUBBYTES[8].a/w1947 , \SUBBYTES[8].a/w1944 , \SUBBYTES[8].a/w1942 ,
         \SUBBYTES[8].a/w1941 , \SUBBYTES[8].a/w1940 , \SUBBYTES[8].a/w1936 ,
         \SUBBYTES[8].a/w1934 , \SUBBYTES[8].a/w1933 , \SUBBYTES[8].a/w1932 ,
         \SUBBYTES[8].a/w1931 , \SUBBYTES[8].a/w1930 , \SUBBYTES[8].a/w1929 ,
         \SUBBYTES[8].a/w1928 , \SUBBYTES[8].a/w1927 , \SUBBYTES[8].a/w1919 ,
         \SUBBYTES[8].a/w1917 , \SUBBYTES[8].a/w1916 , \SUBBYTES[8].a/w1912 ,
         \SUBBYTES[8].a/w1910 , \SUBBYTES[8].a/w1909 , \SUBBYTES[8].a/w1908 ,
         \SUBBYTES[8].a/w1904 , \SUBBYTES[8].a/w1902 , \SUBBYTES[8].a/w1901 ,
         \SUBBYTES[8].a/w1888 , \SUBBYTES[8].a/w1887 , \SUBBYTES[8].a/w1886 ,
         \SUBBYTES[8].a/w1884 , \SUBBYTES[8].a/w1881 , \SUBBYTES[8].a/w1880 ,
         \SUBBYTES[8].a/w1878 , \SUBBYTES[8].a/w1877 , \SUBBYTES[8].a/w1875 ,
         \SUBBYTES[8].a/w1873 , \SUBBYTES[8].a/w1872 , \SUBBYTES[8].a/w1866 ,
         \SUBBYTES[8].a/w1865 , \SUBBYTES[8].a/w1864 , \SUBBYTES[8].a/w1863 ,
         \SUBBYTES[8].a/w1857 , \SUBBYTES[8].a/w1855 , \SUBBYTES[8].a/w1854 ,
         \SUBBYTES[8].a/w1850 , \SUBBYTES[8].a/w1848 , \SUBBYTES[8].a/w1847 ,
         \SUBBYTES[8].a/w1842 , \SUBBYTES[8].a/w1840 , \SUBBYTES[8].a/w1839 ,
         \SUBBYTES[8].a/w1823 , \SUBBYTES[8].a/w1822 , \SUBBYTES[8].a/w1821 ,
         \SUBBYTES[8].a/w1820 , \SUBBYTES[8].a/w1819 , \SUBBYTES[8].a/w1817 ,
         \SUBBYTES[8].a/w1816 , \SUBBYTES[8].a/w1744 , \SUBBYTES[8].a/w1742 ,
         \SUBBYTES[8].a/w1741 , \SUBBYTES[8].a/w1740 , \SUBBYTES[8].a/w1737 ,
         \SUBBYTES[8].a/w1735 , \SUBBYTES[8].a/w1734 , \SUBBYTES[8].a/w1733 ,
         \SUBBYTES[8].a/w1729 , \SUBBYTES[8].a/w1727 , \SUBBYTES[8].a/w1726 ,
         \SUBBYTES[8].a/w1725 , \SUBBYTES[8].a/w1724 , \SUBBYTES[8].a/w1723 ,
         \SUBBYTES[8].a/w1722 , \SUBBYTES[8].a/w1721 , \SUBBYTES[8].a/w1720 ,
         \SUBBYTES[8].a/w1712 , \SUBBYTES[8].a/w1710 , \SUBBYTES[8].a/w1709 ,
         \SUBBYTES[8].a/w1705 , \SUBBYTES[8].a/w1703 , \SUBBYTES[8].a/w1702 ,
         \SUBBYTES[8].a/w1701 , \SUBBYTES[8].a/w1697 , \SUBBYTES[8].a/w1695 ,
         \SUBBYTES[8].a/w1694 , \SUBBYTES[8].a/w1681 , \SUBBYTES[8].a/w1680 ,
         \SUBBYTES[8].a/w1679 , \SUBBYTES[8].a/w1677 , \SUBBYTES[8].a/w1674 ,
         \SUBBYTES[8].a/w1673 , \SUBBYTES[8].a/w1671 , \SUBBYTES[8].a/w1670 ,
         \SUBBYTES[8].a/w1668 , \SUBBYTES[8].a/w1666 , \SUBBYTES[8].a/w1665 ,
         \SUBBYTES[8].a/w1659 , \SUBBYTES[8].a/w1658 , \SUBBYTES[8].a/w1657 ,
         \SUBBYTES[8].a/w1656 , \SUBBYTES[8].a/w1650 , \SUBBYTES[8].a/w1648 ,
         \SUBBYTES[8].a/w1647 , \SUBBYTES[8].a/w1643 , \SUBBYTES[8].a/w1641 ,
         \SUBBYTES[8].a/w1640 , \SUBBYTES[8].a/w1635 , \SUBBYTES[8].a/w1633 ,
         \SUBBYTES[8].a/w1632 , \SUBBYTES[8].a/w1616 , \SUBBYTES[8].a/w1615 ,
         \SUBBYTES[8].a/w1614 , \SUBBYTES[8].a/w1613 , \SUBBYTES[8].a/w1612 ,
         \SUBBYTES[8].a/w1610 , \SUBBYTES[8].a/w1609 , \SUBBYTES[8].a/w1537 ,
         \SUBBYTES[8].a/w1535 , \SUBBYTES[8].a/w1534 , \SUBBYTES[8].a/w1533 ,
         \SUBBYTES[8].a/w1530 , \SUBBYTES[8].a/w1528 , \SUBBYTES[8].a/w1527 ,
         \SUBBYTES[8].a/w1526 , \SUBBYTES[8].a/w1522 , \SUBBYTES[8].a/w1520 ,
         \SUBBYTES[8].a/w1519 , \SUBBYTES[8].a/w1518 , \SUBBYTES[8].a/w1517 ,
         \SUBBYTES[8].a/w1516 , \SUBBYTES[8].a/w1515 , \SUBBYTES[8].a/w1514 ,
         \SUBBYTES[8].a/w1513 , \SUBBYTES[8].a/w1505 , \SUBBYTES[8].a/w1503 ,
         \SUBBYTES[8].a/w1502 , \SUBBYTES[8].a/w1498 , \SUBBYTES[8].a/w1496 ,
         \SUBBYTES[8].a/w1495 , \SUBBYTES[8].a/w1494 , \SUBBYTES[8].a/w1490 ,
         \SUBBYTES[8].a/w1488 , \SUBBYTES[8].a/w1487 , \SUBBYTES[8].a/w1474 ,
         \SUBBYTES[8].a/w1473 , \SUBBYTES[8].a/w1472 , \SUBBYTES[8].a/w1470 ,
         \SUBBYTES[8].a/w1467 , \SUBBYTES[8].a/w1466 , \SUBBYTES[8].a/w1464 ,
         \SUBBYTES[8].a/w1463 , \SUBBYTES[8].a/w1461 , \SUBBYTES[8].a/w1459 ,
         \SUBBYTES[8].a/w1458 , \SUBBYTES[8].a/w1452 , \SUBBYTES[8].a/w1451 ,
         \SUBBYTES[8].a/w1450 , \SUBBYTES[8].a/w1449 , \SUBBYTES[8].a/w1443 ,
         \SUBBYTES[8].a/w1441 , \SUBBYTES[8].a/w1440 , \SUBBYTES[8].a/w1436 ,
         \SUBBYTES[8].a/w1434 , \SUBBYTES[8].a/w1433 , \SUBBYTES[8].a/w1428 ,
         \SUBBYTES[8].a/w1426 , \SUBBYTES[8].a/w1425 , \SUBBYTES[8].a/w1409 ,
         \SUBBYTES[8].a/w1408 , \SUBBYTES[8].a/w1407 , \SUBBYTES[8].a/w1406 ,
         \SUBBYTES[8].a/w1405 , \SUBBYTES[8].a/w1403 , \SUBBYTES[8].a/w1402 ,
         \SUBBYTES[8].a/w1330 , \SUBBYTES[8].a/w1328 , \SUBBYTES[8].a/w1327 ,
         \SUBBYTES[8].a/w1326 , \SUBBYTES[8].a/w1323 , \SUBBYTES[8].a/w1321 ,
         \SUBBYTES[8].a/w1320 , \SUBBYTES[8].a/w1319 , \SUBBYTES[8].a/w1315 ,
         \SUBBYTES[8].a/w1313 , \SUBBYTES[8].a/w1312 , \SUBBYTES[8].a/w1311 ,
         \SUBBYTES[8].a/w1310 , \SUBBYTES[8].a/w1309 , \SUBBYTES[8].a/w1308 ,
         \SUBBYTES[8].a/w1307 , \SUBBYTES[8].a/w1306 , \SUBBYTES[8].a/w1298 ,
         \SUBBYTES[8].a/w1296 , \SUBBYTES[8].a/w1295 , \SUBBYTES[8].a/w1291 ,
         \SUBBYTES[8].a/w1289 , \SUBBYTES[8].a/w1288 , \SUBBYTES[8].a/w1287 ,
         \SUBBYTES[8].a/w1283 , \SUBBYTES[8].a/w1281 , \SUBBYTES[8].a/w1280 ,
         \SUBBYTES[8].a/w1267 , \SUBBYTES[8].a/w1266 , \SUBBYTES[8].a/w1265 ,
         \SUBBYTES[8].a/w1263 , \SUBBYTES[8].a/w1260 , \SUBBYTES[8].a/w1259 ,
         \SUBBYTES[8].a/w1257 , \SUBBYTES[8].a/w1256 , \SUBBYTES[8].a/w1254 ,
         \SUBBYTES[8].a/w1252 , \SUBBYTES[8].a/w1251 , \SUBBYTES[8].a/w1245 ,
         \SUBBYTES[8].a/w1244 , \SUBBYTES[8].a/w1243 , \SUBBYTES[8].a/w1242 ,
         \SUBBYTES[8].a/w1236 , \SUBBYTES[8].a/w1234 , \SUBBYTES[8].a/w1233 ,
         \SUBBYTES[8].a/w1229 , \SUBBYTES[8].a/w1227 , \SUBBYTES[8].a/w1226 ,
         \SUBBYTES[8].a/w1221 , \SUBBYTES[8].a/w1219 , \SUBBYTES[8].a/w1218 ,
         \SUBBYTES[8].a/w1202 , \SUBBYTES[8].a/w1201 , \SUBBYTES[8].a/w1200 ,
         \SUBBYTES[8].a/w1199 , \SUBBYTES[8].a/w1198 , \SUBBYTES[8].a/w1196 ,
         \SUBBYTES[8].a/w1195 , \SUBBYTES[8].a/w1123 , \SUBBYTES[8].a/w1121 ,
         \SUBBYTES[8].a/w1120 , \SUBBYTES[8].a/w1119 , \SUBBYTES[8].a/w1116 ,
         \SUBBYTES[8].a/w1114 , \SUBBYTES[8].a/w1113 , \SUBBYTES[8].a/w1112 ,
         \SUBBYTES[8].a/w1108 , \SUBBYTES[8].a/w1106 , \SUBBYTES[8].a/w1105 ,
         \SUBBYTES[8].a/w1104 , \SUBBYTES[8].a/w1103 , \SUBBYTES[8].a/w1102 ,
         \SUBBYTES[8].a/w1101 , \SUBBYTES[8].a/w1100 , \SUBBYTES[8].a/w1099 ,
         \SUBBYTES[8].a/w1091 , \SUBBYTES[8].a/w1089 , \SUBBYTES[8].a/w1088 ,
         \SUBBYTES[8].a/w1084 , \SUBBYTES[8].a/w1082 , \SUBBYTES[8].a/w1081 ,
         \SUBBYTES[8].a/w1080 , \SUBBYTES[8].a/w1076 , \SUBBYTES[8].a/w1074 ,
         \SUBBYTES[8].a/w1073 , \SUBBYTES[8].a/w1060 , \SUBBYTES[8].a/w1059 ,
         \SUBBYTES[8].a/w1058 , \SUBBYTES[8].a/w1056 , \SUBBYTES[8].a/w1053 ,
         \SUBBYTES[8].a/w1052 , \SUBBYTES[8].a/w1050 , \SUBBYTES[8].a/w1049 ,
         \SUBBYTES[8].a/w1047 , \SUBBYTES[8].a/w1045 , \SUBBYTES[8].a/w1044 ,
         \SUBBYTES[8].a/w1038 , \SUBBYTES[8].a/w1037 , \SUBBYTES[8].a/w1036 ,
         \SUBBYTES[8].a/w1035 , \SUBBYTES[8].a/w1029 , \SUBBYTES[8].a/w1027 ,
         \SUBBYTES[8].a/w1026 , \SUBBYTES[8].a/w1022 , \SUBBYTES[8].a/w1020 ,
         \SUBBYTES[8].a/w1019 , \SUBBYTES[8].a/w1014 , \SUBBYTES[8].a/w1012 ,
         \SUBBYTES[8].a/w1011 , \SUBBYTES[8].a/w995 , \SUBBYTES[8].a/w994 ,
         \SUBBYTES[8].a/w993 , \SUBBYTES[8].a/w992 , \SUBBYTES[8].a/w991 ,
         \SUBBYTES[8].a/w989 , \SUBBYTES[8].a/w988 , \SUBBYTES[8].a/w916 ,
         \SUBBYTES[8].a/w914 , \SUBBYTES[8].a/w913 , \SUBBYTES[8].a/w912 ,
         \SUBBYTES[8].a/w909 , \SUBBYTES[8].a/w907 , \SUBBYTES[8].a/w906 ,
         \SUBBYTES[8].a/w905 , \SUBBYTES[8].a/w901 , \SUBBYTES[8].a/w899 ,
         \SUBBYTES[8].a/w898 , \SUBBYTES[8].a/w897 , \SUBBYTES[8].a/w896 ,
         \SUBBYTES[8].a/w895 , \SUBBYTES[8].a/w894 , \SUBBYTES[8].a/w893 ,
         \SUBBYTES[8].a/w892 , \SUBBYTES[8].a/w884 , \SUBBYTES[8].a/w882 ,
         \SUBBYTES[8].a/w881 , \SUBBYTES[8].a/w877 , \SUBBYTES[8].a/w875 ,
         \SUBBYTES[8].a/w874 , \SUBBYTES[8].a/w873 , \SUBBYTES[8].a/w869 ,
         \SUBBYTES[8].a/w867 , \SUBBYTES[8].a/w866 , \SUBBYTES[8].a/w853 ,
         \SUBBYTES[8].a/w852 , \SUBBYTES[8].a/w851 , \SUBBYTES[8].a/w849 ,
         \SUBBYTES[8].a/w846 , \SUBBYTES[8].a/w845 , \SUBBYTES[8].a/w843 ,
         \SUBBYTES[8].a/w842 , \SUBBYTES[8].a/w840 , \SUBBYTES[8].a/w838 ,
         \SUBBYTES[8].a/w837 , \SUBBYTES[8].a/w831 , \SUBBYTES[8].a/w830 ,
         \SUBBYTES[8].a/w829 , \SUBBYTES[8].a/w828 , \SUBBYTES[8].a/w822 ,
         \SUBBYTES[8].a/w820 , \SUBBYTES[8].a/w819 , \SUBBYTES[8].a/w815 ,
         \SUBBYTES[8].a/w813 , \SUBBYTES[8].a/w812 , \SUBBYTES[8].a/w807 ,
         \SUBBYTES[8].a/w805 , \SUBBYTES[8].a/w804 , \SUBBYTES[8].a/w788 ,
         \SUBBYTES[8].a/w787 , \SUBBYTES[8].a/w786 , \SUBBYTES[8].a/w785 ,
         \SUBBYTES[8].a/w784 , \SUBBYTES[8].a/w782 , \SUBBYTES[8].a/w781 ,
         \SUBBYTES[8].a/w709 , \SUBBYTES[8].a/w707 , \SUBBYTES[8].a/w706 ,
         \SUBBYTES[8].a/w705 , \SUBBYTES[8].a/w702 , \SUBBYTES[8].a/w700 ,
         \SUBBYTES[8].a/w699 , \SUBBYTES[8].a/w698 , \SUBBYTES[8].a/w694 ,
         \SUBBYTES[8].a/w692 , \SUBBYTES[8].a/w691 , \SUBBYTES[8].a/w690 ,
         \SUBBYTES[8].a/w689 , \SUBBYTES[8].a/w688 , \SUBBYTES[8].a/w687 ,
         \SUBBYTES[8].a/w686 , \SUBBYTES[8].a/w685 , \SUBBYTES[8].a/w677 ,
         \SUBBYTES[8].a/w675 , \SUBBYTES[8].a/w674 , \SUBBYTES[8].a/w670 ,
         \SUBBYTES[8].a/w668 , \SUBBYTES[8].a/w667 , \SUBBYTES[8].a/w666 ,
         \SUBBYTES[8].a/w662 , \SUBBYTES[8].a/w660 , \SUBBYTES[8].a/w659 ,
         \SUBBYTES[8].a/w646 , \SUBBYTES[8].a/w645 , \SUBBYTES[8].a/w644 ,
         \SUBBYTES[8].a/w642 , \SUBBYTES[8].a/w639 , \SUBBYTES[8].a/w638 ,
         \SUBBYTES[8].a/w636 , \SUBBYTES[8].a/w635 , \SUBBYTES[8].a/w633 ,
         \SUBBYTES[8].a/w631 , \SUBBYTES[8].a/w630 , \SUBBYTES[8].a/w624 ,
         \SUBBYTES[8].a/w623 , \SUBBYTES[8].a/w622 , \SUBBYTES[8].a/w621 ,
         \SUBBYTES[8].a/w615 , \SUBBYTES[8].a/w613 , \SUBBYTES[8].a/w612 ,
         \SUBBYTES[8].a/w608 , \SUBBYTES[8].a/w606 , \SUBBYTES[8].a/w605 ,
         \SUBBYTES[8].a/w600 , \SUBBYTES[8].a/w598 , \SUBBYTES[8].a/w597 ,
         \SUBBYTES[8].a/w581 , \SUBBYTES[8].a/w580 , \SUBBYTES[8].a/w579 ,
         \SUBBYTES[8].a/w578 , \SUBBYTES[8].a/w577 , \SUBBYTES[8].a/w575 ,
         \SUBBYTES[8].a/w574 , \SUBBYTES[8].a/w502 , \SUBBYTES[8].a/w500 ,
         \SUBBYTES[8].a/w499 , \SUBBYTES[8].a/w498 , \SUBBYTES[8].a/w495 ,
         \SUBBYTES[8].a/w493 , \SUBBYTES[8].a/w492 , \SUBBYTES[8].a/w491 ,
         \SUBBYTES[8].a/w487 , \SUBBYTES[8].a/w485 , \SUBBYTES[8].a/w484 ,
         \SUBBYTES[8].a/w483 , \SUBBYTES[8].a/w482 , \SUBBYTES[8].a/w481 ,
         \SUBBYTES[8].a/w480 , \SUBBYTES[8].a/w479 , \SUBBYTES[8].a/w478 ,
         \SUBBYTES[8].a/w470 , \SUBBYTES[8].a/w468 , \SUBBYTES[8].a/w467 ,
         \SUBBYTES[8].a/w463 , \SUBBYTES[8].a/w461 , \SUBBYTES[8].a/w460 ,
         \SUBBYTES[8].a/w459 , \SUBBYTES[8].a/w455 , \SUBBYTES[8].a/w453 ,
         \SUBBYTES[8].a/w452 , \SUBBYTES[8].a/w439 , \SUBBYTES[8].a/w438 ,
         \SUBBYTES[8].a/w437 , \SUBBYTES[8].a/w435 , \SUBBYTES[8].a/w432 ,
         \SUBBYTES[8].a/w431 , \SUBBYTES[8].a/w429 , \SUBBYTES[8].a/w428 ,
         \SUBBYTES[8].a/w426 , \SUBBYTES[8].a/w424 , \SUBBYTES[8].a/w423 ,
         \SUBBYTES[8].a/w417 , \SUBBYTES[8].a/w416 , \SUBBYTES[8].a/w415 ,
         \SUBBYTES[8].a/w414 , \SUBBYTES[8].a/w408 , \SUBBYTES[8].a/w406 ,
         \SUBBYTES[8].a/w405 , \SUBBYTES[8].a/w401 , \SUBBYTES[8].a/w399 ,
         \SUBBYTES[8].a/w398 , \SUBBYTES[8].a/w393 , \SUBBYTES[8].a/w391 ,
         \SUBBYTES[8].a/w390 , \SUBBYTES[8].a/w374 , \SUBBYTES[8].a/w373 ,
         \SUBBYTES[8].a/w372 , \SUBBYTES[8].a/w371 , \SUBBYTES[8].a/w370 ,
         \SUBBYTES[8].a/w368 , \SUBBYTES[8].a/w367 , \SUBBYTES[8].a/w295 ,
         \SUBBYTES[8].a/w293 , \SUBBYTES[8].a/w292 , \SUBBYTES[8].a/w291 ,
         \SUBBYTES[8].a/w288 , \SUBBYTES[8].a/w286 , \SUBBYTES[8].a/w285 ,
         \SUBBYTES[8].a/w284 , \SUBBYTES[8].a/w280 , \SUBBYTES[8].a/w278 ,
         \SUBBYTES[8].a/w277 , \SUBBYTES[8].a/w276 , \SUBBYTES[8].a/w275 ,
         \SUBBYTES[8].a/w274 , \SUBBYTES[8].a/w273 , \SUBBYTES[8].a/w272 ,
         \SUBBYTES[8].a/w271 , \SUBBYTES[8].a/w263 , \SUBBYTES[8].a/w261 ,
         \SUBBYTES[8].a/w260 , \SUBBYTES[8].a/w256 , \SUBBYTES[8].a/w254 ,
         \SUBBYTES[8].a/w253 , \SUBBYTES[8].a/w252 , \SUBBYTES[8].a/w248 ,
         \SUBBYTES[8].a/w246 , \SUBBYTES[8].a/w245 , \SUBBYTES[8].a/w232 ,
         \SUBBYTES[8].a/w231 , \SUBBYTES[8].a/w230 , \SUBBYTES[8].a/w228 ,
         \SUBBYTES[8].a/w225 , \SUBBYTES[8].a/w224 , \SUBBYTES[8].a/w222 ,
         \SUBBYTES[8].a/w221 , \SUBBYTES[8].a/w219 , \SUBBYTES[8].a/w217 ,
         \SUBBYTES[8].a/w216 , \SUBBYTES[8].a/w210 , \SUBBYTES[8].a/w209 ,
         \SUBBYTES[8].a/w208 , \SUBBYTES[8].a/w207 , \SUBBYTES[8].a/w201 ,
         \SUBBYTES[8].a/w199 , \SUBBYTES[8].a/w198 , \SUBBYTES[8].a/w194 ,
         \SUBBYTES[8].a/w192 , \SUBBYTES[8].a/w191 , \SUBBYTES[8].a/w186 ,
         \SUBBYTES[8].a/w184 , \SUBBYTES[8].a/w183 , \SUBBYTES[8].a/w167 ,
         \SUBBYTES[8].a/w166 , \SUBBYTES[8].a/w165 , \SUBBYTES[8].a/w164 ,
         \SUBBYTES[8].a/w163 , \SUBBYTES[8].a/w161 , \SUBBYTES[8].a/w160 ,
         \SUBBYTES[7].a/w3400 , \SUBBYTES[7].a/w3398 , \SUBBYTES[7].a/w3397 ,
         \SUBBYTES[7].a/w3396 , \SUBBYTES[7].a/w3393 , \SUBBYTES[7].a/w3391 ,
         \SUBBYTES[7].a/w3390 , \SUBBYTES[7].a/w3389 , \SUBBYTES[7].a/w3385 ,
         \SUBBYTES[7].a/w3383 , \SUBBYTES[7].a/w3382 , \SUBBYTES[7].a/w3381 ,
         \SUBBYTES[7].a/w3380 , \SUBBYTES[7].a/w3379 , \SUBBYTES[7].a/w3378 ,
         \SUBBYTES[7].a/w3377 , \SUBBYTES[7].a/w3376 , \SUBBYTES[7].a/w3368 ,
         \SUBBYTES[7].a/w3366 , \SUBBYTES[7].a/w3365 , \SUBBYTES[7].a/w3361 ,
         \SUBBYTES[7].a/w3359 , \SUBBYTES[7].a/w3358 , \SUBBYTES[7].a/w3357 ,
         \SUBBYTES[7].a/w3353 , \SUBBYTES[7].a/w3351 , \SUBBYTES[7].a/w3350 ,
         \SUBBYTES[7].a/w3337 , \SUBBYTES[7].a/w3336 , \SUBBYTES[7].a/w3335 ,
         \SUBBYTES[7].a/w3333 , \SUBBYTES[7].a/w3330 , \SUBBYTES[7].a/w3329 ,
         \SUBBYTES[7].a/w3327 , \SUBBYTES[7].a/w3326 , \SUBBYTES[7].a/w3324 ,
         \SUBBYTES[7].a/w3322 , \SUBBYTES[7].a/w3321 , \SUBBYTES[7].a/w3315 ,
         \SUBBYTES[7].a/w3314 , \SUBBYTES[7].a/w3313 , \SUBBYTES[7].a/w3312 ,
         \SUBBYTES[7].a/w3306 , \SUBBYTES[7].a/w3304 , \SUBBYTES[7].a/w3303 ,
         \SUBBYTES[7].a/w3299 , \SUBBYTES[7].a/w3297 , \SUBBYTES[7].a/w3296 ,
         \SUBBYTES[7].a/w3291 , \SUBBYTES[7].a/w3289 , \SUBBYTES[7].a/w3288 ,
         \SUBBYTES[7].a/w3272 , \SUBBYTES[7].a/w3271 , \SUBBYTES[7].a/w3270 ,
         \SUBBYTES[7].a/w3269 , \SUBBYTES[7].a/w3268 , \SUBBYTES[7].a/w3266 ,
         \SUBBYTES[7].a/w3265 , \SUBBYTES[7].a/w3193 , \SUBBYTES[7].a/w3191 ,
         \SUBBYTES[7].a/w3190 , \SUBBYTES[7].a/w3189 , \SUBBYTES[7].a/w3186 ,
         \SUBBYTES[7].a/w3184 , \SUBBYTES[7].a/w3183 , \SUBBYTES[7].a/w3182 ,
         \SUBBYTES[7].a/w3178 , \SUBBYTES[7].a/w3176 , \SUBBYTES[7].a/w3175 ,
         \SUBBYTES[7].a/w3174 , \SUBBYTES[7].a/w3173 , \SUBBYTES[7].a/w3172 ,
         \SUBBYTES[7].a/w3171 , \SUBBYTES[7].a/w3170 , \SUBBYTES[7].a/w3169 ,
         \SUBBYTES[7].a/w3161 , \SUBBYTES[7].a/w3159 , \SUBBYTES[7].a/w3158 ,
         \SUBBYTES[7].a/w3154 , \SUBBYTES[7].a/w3152 , \SUBBYTES[7].a/w3151 ,
         \SUBBYTES[7].a/w3150 , \SUBBYTES[7].a/w3146 , \SUBBYTES[7].a/w3144 ,
         \SUBBYTES[7].a/w3143 , \SUBBYTES[7].a/w3130 , \SUBBYTES[7].a/w3129 ,
         \SUBBYTES[7].a/w3128 , \SUBBYTES[7].a/w3126 , \SUBBYTES[7].a/w3123 ,
         \SUBBYTES[7].a/w3122 , \SUBBYTES[7].a/w3120 , \SUBBYTES[7].a/w3119 ,
         \SUBBYTES[7].a/w3117 , \SUBBYTES[7].a/w3115 , \SUBBYTES[7].a/w3114 ,
         \SUBBYTES[7].a/w3108 , \SUBBYTES[7].a/w3107 , \SUBBYTES[7].a/w3106 ,
         \SUBBYTES[7].a/w3105 , \SUBBYTES[7].a/w3099 , \SUBBYTES[7].a/w3097 ,
         \SUBBYTES[7].a/w3096 , \SUBBYTES[7].a/w3092 , \SUBBYTES[7].a/w3090 ,
         \SUBBYTES[7].a/w3089 , \SUBBYTES[7].a/w3084 , \SUBBYTES[7].a/w3082 ,
         \SUBBYTES[7].a/w3081 , \SUBBYTES[7].a/w3065 , \SUBBYTES[7].a/w3064 ,
         \SUBBYTES[7].a/w3063 , \SUBBYTES[7].a/w3062 , \SUBBYTES[7].a/w3061 ,
         \SUBBYTES[7].a/w3059 , \SUBBYTES[7].a/w3058 , \SUBBYTES[7].a/w2986 ,
         \SUBBYTES[7].a/w2984 , \SUBBYTES[7].a/w2983 , \SUBBYTES[7].a/w2982 ,
         \SUBBYTES[7].a/w2979 , \SUBBYTES[7].a/w2977 , \SUBBYTES[7].a/w2976 ,
         \SUBBYTES[7].a/w2975 , \SUBBYTES[7].a/w2971 , \SUBBYTES[7].a/w2969 ,
         \SUBBYTES[7].a/w2968 , \SUBBYTES[7].a/w2967 , \SUBBYTES[7].a/w2966 ,
         \SUBBYTES[7].a/w2965 , \SUBBYTES[7].a/w2964 , \SUBBYTES[7].a/w2963 ,
         \SUBBYTES[7].a/w2962 , \SUBBYTES[7].a/w2954 , \SUBBYTES[7].a/w2952 ,
         \SUBBYTES[7].a/w2951 , \SUBBYTES[7].a/w2947 , \SUBBYTES[7].a/w2945 ,
         \SUBBYTES[7].a/w2944 , \SUBBYTES[7].a/w2943 , \SUBBYTES[7].a/w2939 ,
         \SUBBYTES[7].a/w2937 , \SUBBYTES[7].a/w2936 , \SUBBYTES[7].a/w2923 ,
         \SUBBYTES[7].a/w2922 , \SUBBYTES[7].a/w2921 , \SUBBYTES[7].a/w2919 ,
         \SUBBYTES[7].a/w2916 , \SUBBYTES[7].a/w2915 , \SUBBYTES[7].a/w2913 ,
         \SUBBYTES[7].a/w2912 , \SUBBYTES[7].a/w2910 , \SUBBYTES[7].a/w2908 ,
         \SUBBYTES[7].a/w2907 , \SUBBYTES[7].a/w2901 , \SUBBYTES[7].a/w2900 ,
         \SUBBYTES[7].a/w2899 , \SUBBYTES[7].a/w2898 , \SUBBYTES[7].a/w2892 ,
         \SUBBYTES[7].a/w2890 , \SUBBYTES[7].a/w2889 , \SUBBYTES[7].a/w2885 ,
         \SUBBYTES[7].a/w2883 , \SUBBYTES[7].a/w2882 , \SUBBYTES[7].a/w2877 ,
         \SUBBYTES[7].a/w2875 , \SUBBYTES[7].a/w2874 , \SUBBYTES[7].a/w2858 ,
         \SUBBYTES[7].a/w2857 , \SUBBYTES[7].a/w2856 , \SUBBYTES[7].a/w2855 ,
         \SUBBYTES[7].a/w2854 , \SUBBYTES[7].a/w2852 , \SUBBYTES[7].a/w2851 ,
         \SUBBYTES[7].a/w2779 , \SUBBYTES[7].a/w2777 , \SUBBYTES[7].a/w2776 ,
         \SUBBYTES[7].a/w2775 , \SUBBYTES[7].a/w2772 , \SUBBYTES[7].a/w2770 ,
         \SUBBYTES[7].a/w2769 , \SUBBYTES[7].a/w2768 , \SUBBYTES[7].a/w2764 ,
         \SUBBYTES[7].a/w2762 , \SUBBYTES[7].a/w2761 , \SUBBYTES[7].a/w2760 ,
         \SUBBYTES[7].a/w2759 , \SUBBYTES[7].a/w2758 , \SUBBYTES[7].a/w2757 ,
         \SUBBYTES[7].a/w2756 , \SUBBYTES[7].a/w2755 , \SUBBYTES[7].a/w2747 ,
         \SUBBYTES[7].a/w2745 , \SUBBYTES[7].a/w2744 , \SUBBYTES[7].a/w2740 ,
         \SUBBYTES[7].a/w2738 , \SUBBYTES[7].a/w2737 , \SUBBYTES[7].a/w2736 ,
         \SUBBYTES[7].a/w2732 , \SUBBYTES[7].a/w2730 , \SUBBYTES[7].a/w2729 ,
         \SUBBYTES[7].a/w2716 , \SUBBYTES[7].a/w2715 , \SUBBYTES[7].a/w2714 ,
         \SUBBYTES[7].a/w2712 , \SUBBYTES[7].a/w2709 , \SUBBYTES[7].a/w2708 ,
         \SUBBYTES[7].a/w2706 , \SUBBYTES[7].a/w2705 , \SUBBYTES[7].a/w2703 ,
         \SUBBYTES[7].a/w2701 , \SUBBYTES[7].a/w2700 , \SUBBYTES[7].a/w2694 ,
         \SUBBYTES[7].a/w2693 , \SUBBYTES[7].a/w2692 , \SUBBYTES[7].a/w2691 ,
         \SUBBYTES[7].a/w2685 , \SUBBYTES[7].a/w2683 , \SUBBYTES[7].a/w2682 ,
         \SUBBYTES[7].a/w2678 , \SUBBYTES[7].a/w2676 , \SUBBYTES[7].a/w2675 ,
         \SUBBYTES[7].a/w2670 , \SUBBYTES[7].a/w2668 , \SUBBYTES[7].a/w2667 ,
         \SUBBYTES[7].a/w2651 , \SUBBYTES[7].a/w2650 , \SUBBYTES[7].a/w2649 ,
         \SUBBYTES[7].a/w2648 , \SUBBYTES[7].a/w2647 , \SUBBYTES[7].a/w2645 ,
         \SUBBYTES[7].a/w2644 , \SUBBYTES[7].a/w2572 , \SUBBYTES[7].a/w2570 ,
         \SUBBYTES[7].a/w2569 , \SUBBYTES[7].a/w2568 , \SUBBYTES[7].a/w2565 ,
         \SUBBYTES[7].a/w2563 , \SUBBYTES[7].a/w2562 , \SUBBYTES[7].a/w2561 ,
         \SUBBYTES[7].a/w2557 , \SUBBYTES[7].a/w2555 , \SUBBYTES[7].a/w2554 ,
         \SUBBYTES[7].a/w2553 , \SUBBYTES[7].a/w2552 , \SUBBYTES[7].a/w2551 ,
         \SUBBYTES[7].a/w2550 , \SUBBYTES[7].a/w2549 , \SUBBYTES[7].a/w2548 ,
         \SUBBYTES[7].a/w2540 , \SUBBYTES[7].a/w2538 , \SUBBYTES[7].a/w2537 ,
         \SUBBYTES[7].a/w2533 , \SUBBYTES[7].a/w2531 , \SUBBYTES[7].a/w2530 ,
         \SUBBYTES[7].a/w2529 , \SUBBYTES[7].a/w2525 , \SUBBYTES[7].a/w2523 ,
         \SUBBYTES[7].a/w2522 , \SUBBYTES[7].a/w2509 , \SUBBYTES[7].a/w2508 ,
         \SUBBYTES[7].a/w2507 , \SUBBYTES[7].a/w2505 , \SUBBYTES[7].a/w2502 ,
         \SUBBYTES[7].a/w2501 , \SUBBYTES[7].a/w2499 , \SUBBYTES[7].a/w2498 ,
         \SUBBYTES[7].a/w2496 , \SUBBYTES[7].a/w2494 , \SUBBYTES[7].a/w2493 ,
         \SUBBYTES[7].a/w2487 , \SUBBYTES[7].a/w2486 , \SUBBYTES[7].a/w2485 ,
         \SUBBYTES[7].a/w2484 , \SUBBYTES[7].a/w2478 , \SUBBYTES[7].a/w2476 ,
         \SUBBYTES[7].a/w2475 , \SUBBYTES[7].a/w2471 , \SUBBYTES[7].a/w2469 ,
         \SUBBYTES[7].a/w2468 , \SUBBYTES[7].a/w2463 , \SUBBYTES[7].a/w2461 ,
         \SUBBYTES[7].a/w2460 , \SUBBYTES[7].a/w2444 , \SUBBYTES[7].a/w2443 ,
         \SUBBYTES[7].a/w2442 , \SUBBYTES[7].a/w2441 , \SUBBYTES[7].a/w2440 ,
         \SUBBYTES[7].a/w2438 , \SUBBYTES[7].a/w2437 , \SUBBYTES[7].a/w2365 ,
         \SUBBYTES[7].a/w2363 , \SUBBYTES[7].a/w2362 , \SUBBYTES[7].a/w2361 ,
         \SUBBYTES[7].a/w2358 , \SUBBYTES[7].a/w2356 , \SUBBYTES[7].a/w2355 ,
         \SUBBYTES[7].a/w2354 , \SUBBYTES[7].a/w2350 , \SUBBYTES[7].a/w2348 ,
         \SUBBYTES[7].a/w2347 , \SUBBYTES[7].a/w2346 , \SUBBYTES[7].a/w2345 ,
         \SUBBYTES[7].a/w2344 , \SUBBYTES[7].a/w2343 , \SUBBYTES[7].a/w2342 ,
         \SUBBYTES[7].a/w2341 , \SUBBYTES[7].a/w2333 , \SUBBYTES[7].a/w2331 ,
         \SUBBYTES[7].a/w2330 , \SUBBYTES[7].a/w2326 , \SUBBYTES[7].a/w2324 ,
         \SUBBYTES[7].a/w2323 , \SUBBYTES[7].a/w2322 , \SUBBYTES[7].a/w2318 ,
         \SUBBYTES[7].a/w2316 , \SUBBYTES[7].a/w2315 , \SUBBYTES[7].a/w2302 ,
         \SUBBYTES[7].a/w2301 , \SUBBYTES[7].a/w2300 , \SUBBYTES[7].a/w2298 ,
         \SUBBYTES[7].a/w2295 , \SUBBYTES[7].a/w2294 , \SUBBYTES[7].a/w2292 ,
         \SUBBYTES[7].a/w2291 , \SUBBYTES[7].a/w2289 , \SUBBYTES[7].a/w2287 ,
         \SUBBYTES[7].a/w2286 , \SUBBYTES[7].a/w2280 , \SUBBYTES[7].a/w2279 ,
         \SUBBYTES[7].a/w2278 , \SUBBYTES[7].a/w2277 , \SUBBYTES[7].a/w2271 ,
         \SUBBYTES[7].a/w2269 , \SUBBYTES[7].a/w2268 , \SUBBYTES[7].a/w2264 ,
         \SUBBYTES[7].a/w2262 , \SUBBYTES[7].a/w2261 , \SUBBYTES[7].a/w2256 ,
         \SUBBYTES[7].a/w2254 , \SUBBYTES[7].a/w2253 , \SUBBYTES[7].a/w2237 ,
         \SUBBYTES[7].a/w2236 , \SUBBYTES[7].a/w2235 , \SUBBYTES[7].a/w2234 ,
         \SUBBYTES[7].a/w2233 , \SUBBYTES[7].a/w2231 , \SUBBYTES[7].a/w2230 ,
         \SUBBYTES[7].a/w2158 , \SUBBYTES[7].a/w2156 , \SUBBYTES[7].a/w2155 ,
         \SUBBYTES[7].a/w2154 , \SUBBYTES[7].a/w2151 , \SUBBYTES[7].a/w2149 ,
         \SUBBYTES[7].a/w2148 , \SUBBYTES[7].a/w2147 , \SUBBYTES[7].a/w2143 ,
         \SUBBYTES[7].a/w2141 , \SUBBYTES[7].a/w2140 , \SUBBYTES[7].a/w2139 ,
         \SUBBYTES[7].a/w2138 , \SUBBYTES[7].a/w2137 , \SUBBYTES[7].a/w2136 ,
         \SUBBYTES[7].a/w2135 , \SUBBYTES[7].a/w2134 , \SUBBYTES[7].a/w2126 ,
         \SUBBYTES[7].a/w2124 , \SUBBYTES[7].a/w2123 , \SUBBYTES[7].a/w2119 ,
         \SUBBYTES[7].a/w2117 , \SUBBYTES[7].a/w2116 , \SUBBYTES[7].a/w2115 ,
         \SUBBYTES[7].a/w2111 , \SUBBYTES[7].a/w2109 , \SUBBYTES[7].a/w2108 ,
         \SUBBYTES[7].a/w2095 , \SUBBYTES[7].a/w2094 , \SUBBYTES[7].a/w2093 ,
         \SUBBYTES[7].a/w2091 , \SUBBYTES[7].a/w2088 , \SUBBYTES[7].a/w2087 ,
         \SUBBYTES[7].a/w2085 , \SUBBYTES[7].a/w2084 , \SUBBYTES[7].a/w2082 ,
         \SUBBYTES[7].a/w2080 , \SUBBYTES[7].a/w2079 , \SUBBYTES[7].a/w2073 ,
         \SUBBYTES[7].a/w2072 , \SUBBYTES[7].a/w2071 , \SUBBYTES[7].a/w2070 ,
         \SUBBYTES[7].a/w2064 , \SUBBYTES[7].a/w2062 , \SUBBYTES[7].a/w2061 ,
         \SUBBYTES[7].a/w2057 , \SUBBYTES[7].a/w2055 , \SUBBYTES[7].a/w2054 ,
         \SUBBYTES[7].a/w2049 , \SUBBYTES[7].a/w2047 , \SUBBYTES[7].a/w2046 ,
         \SUBBYTES[7].a/w2030 , \SUBBYTES[7].a/w2029 , \SUBBYTES[7].a/w2028 ,
         \SUBBYTES[7].a/w2027 , \SUBBYTES[7].a/w2026 , \SUBBYTES[7].a/w2024 ,
         \SUBBYTES[7].a/w2023 , \SUBBYTES[7].a/w1951 , \SUBBYTES[7].a/w1949 ,
         \SUBBYTES[7].a/w1948 , \SUBBYTES[7].a/w1947 , \SUBBYTES[7].a/w1944 ,
         \SUBBYTES[7].a/w1942 , \SUBBYTES[7].a/w1941 , \SUBBYTES[7].a/w1940 ,
         \SUBBYTES[7].a/w1936 , \SUBBYTES[7].a/w1934 , \SUBBYTES[7].a/w1933 ,
         \SUBBYTES[7].a/w1932 , \SUBBYTES[7].a/w1931 , \SUBBYTES[7].a/w1930 ,
         \SUBBYTES[7].a/w1929 , \SUBBYTES[7].a/w1928 , \SUBBYTES[7].a/w1927 ,
         \SUBBYTES[7].a/w1919 , \SUBBYTES[7].a/w1917 , \SUBBYTES[7].a/w1916 ,
         \SUBBYTES[7].a/w1912 , \SUBBYTES[7].a/w1910 , \SUBBYTES[7].a/w1909 ,
         \SUBBYTES[7].a/w1908 , \SUBBYTES[7].a/w1904 , \SUBBYTES[7].a/w1902 ,
         \SUBBYTES[7].a/w1901 , \SUBBYTES[7].a/w1888 , \SUBBYTES[7].a/w1887 ,
         \SUBBYTES[7].a/w1886 , \SUBBYTES[7].a/w1884 , \SUBBYTES[7].a/w1881 ,
         \SUBBYTES[7].a/w1880 , \SUBBYTES[7].a/w1878 , \SUBBYTES[7].a/w1877 ,
         \SUBBYTES[7].a/w1875 , \SUBBYTES[7].a/w1873 , \SUBBYTES[7].a/w1872 ,
         \SUBBYTES[7].a/w1866 , \SUBBYTES[7].a/w1865 , \SUBBYTES[7].a/w1864 ,
         \SUBBYTES[7].a/w1863 , \SUBBYTES[7].a/w1857 , \SUBBYTES[7].a/w1855 ,
         \SUBBYTES[7].a/w1854 , \SUBBYTES[7].a/w1850 , \SUBBYTES[7].a/w1848 ,
         \SUBBYTES[7].a/w1847 , \SUBBYTES[7].a/w1842 , \SUBBYTES[7].a/w1840 ,
         \SUBBYTES[7].a/w1839 , \SUBBYTES[7].a/w1823 , \SUBBYTES[7].a/w1822 ,
         \SUBBYTES[7].a/w1821 , \SUBBYTES[7].a/w1820 , \SUBBYTES[7].a/w1819 ,
         \SUBBYTES[7].a/w1817 , \SUBBYTES[7].a/w1816 , \SUBBYTES[7].a/w1744 ,
         \SUBBYTES[7].a/w1742 , \SUBBYTES[7].a/w1741 , \SUBBYTES[7].a/w1740 ,
         \SUBBYTES[7].a/w1737 , \SUBBYTES[7].a/w1735 , \SUBBYTES[7].a/w1734 ,
         \SUBBYTES[7].a/w1733 , \SUBBYTES[7].a/w1729 , \SUBBYTES[7].a/w1727 ,
         \SUBBYTES[7].a/w1726 , \SUBBYTES[7].a/w1725 , \SUBBYTES[7].a/w1724 ,
         \SUBBYTES[7].a/w1723 , \SUBBYTES[7].a/w1722 , \SUBBYTES[7].a/w1721 ,
         \SUBBYTES[7].a/w1720 , \SUBBYTES[7].a/w1712 , \SUBBYTES[7].a/w1710 ,
         \SUBBYTES[7].a/w1709 , \SUBBYTES[7].a/w1705 , \SUBBYTES[7].a/w1703 ,
         \SUBBYTES[7].a/w1702 , \SUBBYTES[7].a/w1701 , \SUBBYTES[7].a/w1697 ,
         \SUBBYTES[7].a/w1695 , \SUBBYTES[7].a/w1694 , \SUBBYTES[7].a/w1681 ,
         \SUBBYTES[7].a/w1680 , \SUBBYTES[7].a/w1679 , \SUBBYTES[7].a/w1677 ,
         \SUBBYTES[7].a/w1674 , \SUBBYTES[7].a/w1673 , \SUBBYTES[7].a/w1671 ,
         \SUBBYTES[7].a/w1670 , \SUBBYTES[7].a/w1668 , \SUBBYTES[7].a/w1666 ,
         \SUBBYTES[7].a/w1665 , \SUBBYTES[7].a/w1659 , \SUBBYTES[7].a/w1658 ,
         \SUBBYTES[7].a/w1657 , \SUBBYTES[7].a/w1656 , \SUBBYTES[7].a/w1650 ,
         \SUBBYTES[7].a/w1648 , \SUBBYTES[7].a/w1647 , \SUBBYTES[7].a/w1643 ,
         \SUBBYTES[7].a/w1641 , \SUBBYTES[7].a/w1640 , \SUBBYTES[7].a/w1635 ,
         \SUBBYTES[7].a/w1633 , \SUBBYTES[7].a/w1632 , \SUBBYTES[7].a/w1616 ,
         \SUBBYTES[7].a/w1615 , \SUBBYTES[7].a/w1614 , \SUBBYTES[7].a/w1613 ,
         \SUBBYTES[7].a/w1612 , \SUBBYTES[7].a/w1610 , \SUBBYTES[7].a/w1609 ,
         \SUBBYTES[7].a/w1537 , \SUBBYTES[7].a/w1535 , \SUBBYTES[7].a/w1534 ,
         \SUBBYTES[7].a/w1533 , \SUBBYTES[7].a/w1530 , \SUBBYTES[7].a/w1528 ,
         \SUBBYTES[7].a/w1527 , \SUBBYTES[7].a/w1526 , \SUBBYTES[7].a/w1522 ,
         \SUBBYTES[7].a/w1520 , \SUBBYTES[7].a/w1519 , \SUBBYTES[7].a/w1518 ,
         \SUBBYTES[7].a/w1517 , \SUBBYTES[7].a/w1516 , \SUBBYTES[7].a/w1515 ,
         \SUBBYTES[7].a/w1514 , \SUBBYTES[7].a/w1513 , \SUBBYTES[7].a/w1505 ,
         \SUBBYTES[7].a/w1503 , \SUBBYTES[7].a/w1502 , \SUBBYTES[7].a/w1498 ,
         \SUBBYTES[7].a/w1496 , \SUBBYTES[7].a/w1495 , \SUBBYTES[7].a/w1494 ,
         \SUBBYTES[7].a/w1490 , \SUBBYTES[7].a/w1488 , \SUBBYTES[7].a/w1487 ,
         \SUBBYTES[7].a/w1474 , \SUBBYTES[7].a/w1473 , \SUBBYTES[7].a/w1472 ,
         \SUBBYTES[7].a/w1470 , \SUBBYTES[7].a/w1467 , \SUBBYTES[7].a/w1466 ,
         \SUBBYTES[7].a/w1464 , \SUBBYTES[7].a/w1463 , \SUBBYTES[7].a/w1461 ,
         \SUBBYTES[7].a/w1459 , \SUBBYTES[7].a/w1458 , \SUBBYTES[7].a/w1452 ,
         \SUBBYTES[7].a/w1451 , \SUBBYTES[7].a/w1450 , \SUBBYTES[7].a/w1449 ,
         \SUBBYTES[7].a/w1443 , \SUBBYTES[7].a/w1441 , \SUBBYTES[7].a/w1440 ,
         \SUBBYTES[7].a/w1436 , \SUBBYTES[7].a/w1434 , \SUBBYTES[7].a/w1433 ,
         \SUBBYTES[7].a/w1428 , \SUBBYTES[7].a/w1426 , \SUBBYTES[7].a/w1425 ,
         \SUBBYTES[7].a/w1409 , \SUBBYTES[7].a/w1408 , \SUBBYTES[7].a/w1407 ,
         \SUBBYTES[7].a/w1406 , \SUBBYTES[7].a/w1405 , \SUBBYTES[7].a/w1403 ,
         \SUBBYTES[7].a/w1402 , \SUBBYTES[7].a/w1330 , \SUBBYTES[7].a/w1328 ,
         \SUBBYTES[7].a/w1327 , \SUBBYTES[7].a/w1326 , \SUBBYTES[7].a/w1323 ,
         \SUBBYTES[7].a/w1321 , \SUBBYTES[7].a/w1320 , \SUBBYTES[7].a/w1319 ,
         \SUBBYTES[7].a/w1315 , \SUBBYTES[7].a/w1313 , \SUBBYTES[7].a/w1312 ,
         \SUBBYTES[7].a/w1311 , \SUBBYTES[7].a/w1310 , \SUBBYTES[7].a/w1309 ,
         \SUBBYTES[7].a/w1308 , \SUBBYTES[7].a/w1307 , \SUBBYTES[7].a/w1306 ,
         \SUBBYTES[7].a/w1298 , \SUBBYTES[7].a/w1296 , \SUBBYTES[7].a/w1295 ,
         \SUBBYTES[7].a/w1291 , \SUBBYTES[7].a/w1289 , \SUBBYTES[7].a/w1288 ,
         \SUBBYTES[7].a/w1287 , \SUBBYTES[7].a/w1283 , \SUBBYTES[7].a/w1281 ,
         \SUBBYTES[7].a/w1280 , \SUBBYTES[7].a/w1267 , \SUBBYTES[7].a/w1266 ,
         \SUBBYTES[7].a/w1265 , \SUBBYTES[7].a/w1263 , \SUBBYTES[7].a/w1260 ,
         \SUBBYTES[7].a/w1259 , \SUBBYTES[7].a/w1257 , \SUBBYTES[7].a/w1256 ,
         \SUBBYTES[7].a/w1254 , \SUBBYTES[7].a/w1252 , \SUBBYTES[7].a/w1251 ,
         \SUBBYTES[7].a/w1245 , \SUBBYTES[7].a/w1244 , \SUBBYTES[7].a/w1243 ,
         \SUBBYTES[7].a/w1242 , \SUBBYTES[7].a/w1236 , \SUBBYTES[7].a/w1234 ,
         \SUBBYTES[7].a/w1233 , \SUBBYTES[7].a/w1229 , \SUBBYTES[7].a/w1227 ,
         \SUBBYTES[7].a/w1226 , \SUBBYTES[7].a/w1221 , \SUBBYTES[7].a/w1219 ,
         \SUBBYTES[7].a/w1218 , \SUBBYTES[7].a/w1202 , \SUBBYTES[7].a/w1201 ,
         \SUBBYTES[7].a/w1200 , \SUBBYTES[7].a/w1199 , \SUBBYTES[7].a/w1198 ,
         \SUBBYTES[7].a/w1196 , \SUBBYTES[7].a/w1195 , \SUBBYTES[7].a/w1123 ,
         \SUBBYTES[7].a/w1121 , \SUBBYTES[7].a/w1120 , \SUBBYTES[7].a/w1119 ,
         \SUBBYTES[7].a/w1116 , \SUBBYTES[7].a/w1114 , \SUBBYTES[7].a/w1113 ,
         \SUBBYTES[7].a/w1112 , \SUBBYTES[7].a/w1108 , \SUBBYTES[7].a/w1106 ,
         \SUBBYTES[7].a/w1105 , \SUBBYTES[7].a/w1104 , \SUBBYTES[7].a/w1103 ,
         \SUBBYTES[7].a/w1102 , \SUBBYTES[7].a/w1101 , \SUBBYTES[7].a/w1100 ,
         \SUBBYTES[7].a/w1099 , \SUBBYTES[7].a/w1091 , \SUBBYTES[7].a/w1089 ,
         \SUBBYTES[7].a/w1088 , \SUBBYTES[7].a/w1084 , \SUBBYTES[7].a/w1082 ,
         \SUBBYTES[7].a/w1081 , \SUBBYTES[7].a/w1080 , \SUBBYTES[7].a/w1076 ,
         \SUBBYTES[7].a/w1074 , \SUBBYTES[7].a/w1073 , \SUBBYTES[7].a/w1060 ,
         \SUBBYTES[7].a/w1059 , \SUBBYTES[7].a/w1058 , \SUBBYTES[7].a/w1056 ,
         \SUBBYTES[7].a/w1053 , \SUBBYTES[7].a/w1052 , \SUBBYTES[7].a/w1050 ,
         \SUBBYTES[7].a/w1049 , \SUBBYTES[7].a/w1047 , \SUBBYTES[7].a/w1045 ,
         \SUBBYTES[7].a/w1044 , \SUBBYTES[7].a/w1038 , \SUBBYTES[7].a/w1037 ,
         \SUBBYTES[7].a/w1036 , \SUBBYTES[7].a/w1035 , \SUBBYTES[7].a/w1029 ,
         \SUBBYTES[7].a/w1027 , \SUBBYTES[7].a/w1026 , \SUBBYTES[7].a/w1022 ,
         \SUBBYTES[7].a/w1020 , \SUBBYTES[7].a/w1019 , \SUBBYTES[7].a/w1014 ,
         \SUBBYTES[7].a/w1012 , \SUBBYTES[7].a/w1011 , \SUBBYTES[7].a/w995 ,
         \SUBBYTES[7].a/w994 , \SUBBYTES[7].a/w993 , \SUBBYTES[7].a/w992 ,
         \SUBBYTES[7].a/w991 , \SUBBYTES[7].a/w989 , \SUBBYTES[7].a/w988 ,
         \SUBBYTES[7].a/w916 , \SUBBYTES[7].a/w914 , \SUBBYTES[7].a/w913 ,
         \SUBBYTES[7].a/w912 , \SUBBYTES[7].a/w909 , \SUBBYTES[7].a/w907 ,
         \SUBBYTES[7].a/w906 , \SUBBYTES[7].a/w905 , \SUBBYTES[7].a/w901 ,
         \SUBBYTES[7].a/w899 , \SUBBYTES[7].a/w898 , \SUBBYTES[7].a/w897 ,
         \SUBBYTES[7].a/w896 , \SUBBYTES[7].a/w895 , \SUBBYTES[7].a/w894 ,
         \SUBBYTES[7].a/w893 , \SUBBYTES[7].a/w892 , \SUBBYTES[7].a/w884 ,
         \SUBBYTES[7].a/w882 , \SUBBYTES[7].a/w881 , \SUBBYTES[7].a/w877 ,
         \SUBBYTES[7].a/w875 , \SUBBYTES[7].a/w874 , \SUBBYTES[7].a/w873 ,
         \SUBBYTES[7].a/w869 , \SUBBYTES[7].a/w867 , \SUBBYTES[7].a/w866 ,
         \SUBBYTES[7].a/w853 , \SUBBYTES[7].a/w852 , \SUBBYTES[7].a/w851 ,
         \SUBBYTES[7].a/w849 , \SUBBYTES[7].a/w846 , \SUBBYTES[7].a/w845 ,
         \SUBBYTES[7].a/w843 , \SUBBYTES[7].a/w842 , \SUBBYTES[7].a/w840 ,
         \SUBBYTES[7].a/w838 , \SUBBYTES[7].a/w837 , \SUBBYTES[7].a/w831 ,
         \SUBBYTES[7].a/w830 , \SUBBYTES[7].a/w829 , \SUBBYTES[7].a/w828 ,
         \SUBBYTES[7].a/w822 , \SUBBYTES[7].a/w820 , \SUBBYTES[7].a/w819 ,
         \SUBBYTES[7].a/w815 , \SUBBYTES[7].a/w813 , \SUBBYTES[7].a/w812 ,
         \SUBBYTES[7].a/w807 , \SUBBYTES[7].a/w805 , \SUBBYTES[7].a/w804 ,
         \SUBBYTES[7].a/w788 , \SUBBYTES[7].a/w787 , \SUBBYTES[7].a/w786 ,
         \SUBBYTES[7].a/w785 , \SUBBYTES[7].a/w784 , \SUBBYTES[7].a/w782 ,
         \SUBBYTES[7].a/w781 , \SUBBYTES[7].a/w709 , \SUBBYTES[7].a/w707 ,
         \SUBBYTES[7].a/w706 , \SUBBYTES[7].a/w705 , \SUBBYTES[7].a/w702 ,
         \SUBBYTES[7].a/w700 , \SUBBYTES[7].a/w699 , \SUBBYTES[7].a/w698 ,
         \SUBBYTES[7].a/w694 , \SUBBYTES[7].a/w692 , \SUBBYTES[7].a/w691 ,
         \SUBBYTES[7].a/w690 , \SUBBYTES[7].a/w689 , \SUBBYTES[7].a/w688 ,
         \SUBBYTES[7].a/w687 , \SUBBYTES[7].a/w686 , \SUBBYTES[7].a/w685 ,
         \SUBBYTES[7].a/w677 , \SUBBYTES[7].a/w675 , \SUBBYTES[7].a/w674 ,
         \SUBBYTES[7].a/w670 , \SUBBYTES[7].a/w668 , \SUBBYTES[7].a/w667 ,
         \SUBBYTES[7].a/w666 , \SUBBYTES[7].a/w662 , \SUBBYTES[7].a/w660 ,
         \SUBBYTES[7].a/w659 , \SUBBYTES[7].a/w646 , \SUBBYTES[7].a/w645 ,
         \SUBBYTES[7].a/w644 , \SUBBYTES[7].a/w642 , \SUBBYTES[7].a/w639 ,
         \SUBBYTES[7].a/w638 , \SUBBYTES[7].a/w636 , \SUBBYTES[7].a/w635 ,
         \SUBBYTES[7].a/w633 , \SUBBYTES[7].a/w631 , \SUBBYTES[7].a/w630 ,
         \SUBBYTES[7].a/w624 , \SUBBYTES[7].a/w623 , \SUBBYTES[7].a/w622 ,
         \SUBBYTES[7].a/w621 , \SUBBYTES[7].a/w615 , \SUBBYTES[7].a/w613 ,
         \SUBBYTES[7].a/w612 , \SUBBYTES[7].a/w608 , \SUBBYTES[7].a/w606 ,
         \SUBBYTES[7].a/w605 , \SUBBYTES[7].a/w600 , \SUBBYTES[7].a/w598 ,
         \SUBBYTES[7].a/w597 , \SUBBYTES[7].a/w581 , \SUBBYTES[7].a/w580 ,
         \SUBBYTES[7].a/w579 , \SUBBYTES[7].a/w578 , \SUBBYTES[7].a/w577 ,
         \SUBBYTES[7].a/w575 , \SUBBYTES[7].a/w574 , \SUBBYTES[7].a/w502 ,
         \SUBBYTES[7].a/w500 , \SUBBYTES[7].a/w499 , \SUBBYTES[7].a/w498 ,
         \SUBBYTES[7].a/w495 , \SUBBYTES[7].a/w493 , \SUBBYTES[7].a/w492 ,
         \SUBBYTES[7].a/w491 , \SUBBYTES[7].a/w487 , \SUBBYTES[7].a/w485 ,
         \SUBBYTES[7].a/w484 , \SUBBYTES[7].a/w483 , \SUBBYTES[7].a/w482 ,
         \SUBBYTES[7].a/w481 , \SUBBYTES[7].a/w480 , \SUBBYTES[7].a/w479 ,
         \SUBBYTES[7].a/w478 , \SUBBYTES[7].a/w470 , \SUBBYTES[7].a/w468 ,
         \SUBBYTES[7].a/w467 , \SUBBYTES[7].a/w463 , \SUBBYTES[7].a/w461 ,
         \SUBBYTES[7].a/w460 , \SUBBYTES[7].a/w459 , \SUBBYTES[7].a/w455 ,
         \SUBBYTES[7].a/w453 , \SUBBYTES[7].a/w452 , \SUBBYTES[7].a/w439 ,
         \SUBBYTES[7].a/w438 , \SUBBYTES[7].a/w437 , \SUBBYTES[7].a/w435 ,
         \SUBBYTES[7].a/w432 , \SUBBYTES[7].a/w431 , \SUBBYTES[7].a/w429 ,
         \SUBBYTES[7].a/w428 , \SUBBYTES[7].a/w426 , \SUBBYTES[7].a/w424 ,
         \SUBBYTES[7].a/w423 , \SUBBYTES[7].a/w417 , \SUBBYTES[7].a/w416 ,
         \SUBBYTES[7].a/w415 , \SUBBYTES[7].a/w414 , \SUBBYTES[7].a/w408 ,
         \SUBBYTES[7].a/w406 , \SUBBYTES[7].a/w405 , \SUBBYTES[7].a/w401 ,
         \SUBBYTES[7].a/w399 , \SUBBYTES[7].a/w398 , \SUBBYTES[7].a/w393 ,
         \SUBBYTES[7].a/w391 , \SUBBYTES[7].a/w390 , \SUBBYTES[7].a/w374 ,
         \SUBBYTES[7].a/w373 , \SUBBYTES[7].a/w372 , \SUBBYTES[7].a/w371 ,
         \SUBBYTES[7].a/w370 , \SUBBYTES[7].a/w368 , \SUBBYTES[7].a/w367 ,
         \SUBBYTES[7].a/w295 , \SUBBYTES[7].a/w293 , \SUBBYTES[7].a/w292 ,
         \SUBBYTES[7].a/w291 , \SUBBYTES[7].a/w288 , \SUBBYTES[7].a/w286 ,
         \SUBBYTES[7].a/w285 , \SUBBYTES[7].a/w284 , \SUBBYTES[7].a/w280 ,
         \SUBBYTES[7].a/w278 , \SUBBYTES[7].a/w277 , \SUBBYTES[7].a/w276 ,
         \SUBBYTES[7].a/w275 , \SUBBYTES[7].a/w274 , \SUBBYTES[7].a/w273 ,
         \SUBBYTES[7].a/w272 , \SUBBYTES[7].a/w271 , \SUBBYTES[7].a/w263 ,
         \SUBBYTES[7].a/w261 , \SUBBYTES[7].a/w260 , \SUBBYTES[7].a/w256 ,
         \SUBBYTES[7].a/w254 , \SUBBYTES[7].a/w253 , \SUBBYTES[7].a/w252 ,
         \SUBBYTES[7].a/w248 , \SUBBYTES[7].a/w246 , \SUBBYTES[7].a/w245 ,
         \SUBBYTES[7].a/w232 , \SUBBYTES[7].a/w231 , \SUBBYTES[7].a/w230 ,
         \SUBBYTES[7].a/w228 , \SUBBYTES[7].a/w225 , \SUBBYTES[7].a/w224 ,
         \SUBBYTES[7].a/w222 , \SUBBYTES[7].a/w221 , \SUBBYTES[7].a/w219 ,
         \SUBBYTES[7].a/w217 , \SUBBYTES[7].a/w216 , \SUBBYTES[7].a/w210 ,
         \SUBBYTES[7].a/w209 , \SUBBYTES[7].a/w208 , \SUBBYTES[7].a/w207 ,
         \SUBBYTES[7].a/w201 , \SUBBYTES[7].a/w199 , \SUBBYTES[7].a/w198 ,
         \SUBBYTES[7].a/w194 , \SUBBYTES[7].a/w192 , \SUBBYTES[7].a/w191 ,
         \SUBBYTES[7].a/w186 , \SUBBYTES[7].a/w184 , \SUBBYTES[7].a/w183 ,
         \SUBBYTES[7].a/w167 , \SUBBYTES[7].a/w166 , \SUBBYTES[7].a/w165 ,
         \SUBBYTES[7].a/w164 , \SUBBYTES[7].a/w163 , \SUBBYTES[7].a/w161 ,
         \SUBBYTES[7].a/w160 , \SUBBYTES[6].a/w3400 , \SUBBYTES[6].a/w3398 ,
         \SUBBYTES[6].a/w3397 , \SUBBYTES[6].a/w3396 , \SUBBYTES[6].a/w3393 ,
         \SUBBYTES[6].a/w3391 , \SUBBYTES[6].a/w3390 , \SUBBYTES[6].a/w3389 ,
         \SUBBYTES[6].a/w3385 , \SUBBYTES[6].a/w3383 , \SUBBYTES[6].a/w3382 ,
         \SUBBYTES[6].a/w3381 , \SUBBYTES[6].a/w3380 , \SUBBYTES[6].a/w3379 ,
         \SUBBYTES[6].a/w3378 , \SUBBYTES[6].a/w3377 , \SUBBYTES[6].a/w3376 ,
         \SUBBYTES[6].a/w3368 , \SUBBYTES[6].a/w3366 , \SUBBYTES[6].a/w3365 ,
         \SUBBYTES[6].a/w3361 , \SUBBYTES[6].a/w3359 , \SUBBYTES[6].a/w3358 ,
         \SUBBYTES[6].a/w3357 , \SUBBYTES[6].a/w3353 , \SUBBYTES[6].a/w3351 ,
         \SUBBYTES[6].a/w3350 , \SUBBYTES[6].a/w3337 , \SUBBYTES[6].a/w3336 ,
         \SUBBYTES[6].a/w3335 , \SUBBYTES[6].a/w3333 , \SUBBYTES[6].a/w3330 ,
         \SUBBYTES[6].a/w3329 , \SUBBYTES[6].a/w3327 , \SUBBYTES[6].a/w3326 ,
         \SUBBYTES[6].a/w3324 , \SUBBYTES[6].a/w3322 , \SUBBYTES[6].a/w3321 ,
         \SUBBYTES[6].a/w3315 , \SUBBYTES[6].a/w3314 , \SUBBYTES[6].a/w3313 ,
         \SUBBYTES[6].a/w3312 , \SUBBYTES[6].a/w3306 , \SUBBYTES[6].a/w3304 ,
         \SUBBYTES[6].a/w3303 , \SUBBYTES[6].a/w3299 , \SUBBYTES[6].a/w3297 ,
         \SUBBYTES[6].a/w3296 , \SUBBYTES[6].a/w3291 , \SUBBYTES[6].a/w3289 ,
         \SUBBYTES[6].a/w3288 , \SUBBYTES[6].a/w3272 , \SUBBYTES[6].a/w3271 ,
         \SUBBYTES[6].a/w3270 , \SUBBYTES[6].a/w3269 , \SUBBYTES[6].a/w3268 ,
         \SUBBYTES[6].a/w3266 , \SUBBYTES[6].a/w3265 , \SUBBYTES[6].a/w3193 ,
         \SUBBYTES[6].a/w3191 , \SUBBYTES[6].a/w3190 , \SUBBYTES[6].a/w3189 ,
         \SUBBYTES[6].a/w3186 , \SUBBYTES[6].a/w3184 , \SUBBYTES[6].a/w3183 ,
         \SUBBYTES[6].a/w3182 , \SUBBYTES[6].a/w3178 , \SUBBYTES[6].a/w3176 ,
         \SUBBYTES[6].a/w3175 , \SUBBYTES[6].a/w3174 , \SUBBYTES[6].a/w3173 ,
         \SUBBYTES[6].a/w3172 , \SUBBYTES[6].a/w3171 , \SUBBYTES[6].a/w3170 ,
         \SUBBYTES[6].a/w3169 , \SUBBYTES[6].a/w3161 , \SUBBYTES[6].a/w3159 ,
         \SUBBYTES[6].a/w3158 , \SUBBYTES[6].a/w3154 , \SUBBYTES[6].a/w3152 ,
         \SUBBYTES[6].a/w3151 , \SUBBYTES[6].a/w3150 , \SUBBYTES[6].a/w3146 ,
         \SUBBYTES[6].a/w3144 , \SUBBYTES[6].a/w3143 , \SUBBYTES[6].a/w3130 ,
         \SUBBYTES[6].a/w3129 , \SUBBYTES[6].a/w3128 , \SUBBYTES[6].a/w3126 ,
         \SUBBYTES[6].a/w3123 , \SUBBYTES[6].a/w3122 , \SUBBYTES[6].a/w3120 ,
         \SUBBYTES[6].a/w3119 , \SUBBYTES[6].a/w3117 , \SUBBYTES[6].a/w3115 ,
         \SUBBYTES[6].a/w3114 , \SUBBYTES[6].a/w3108 , \SUBBYTES[6].a/w3107 ,
         \SUBBYTES[6].a/w3106 , \SUBBYTES[6].a/w3105 , \SUBBYTES[6].a/w3099 ,
         \SUBBYTES[6].a/w3097 , \SUBBYTES[6].a/w3096 , \SUBBYTES[6].a/w3092 ,
         \SUBBYTES[6].a/w3090 , \SUBBYTES[6].a/w3089 , \SUBBYTES[6].a/w3084 ,
         \SUBBYTES[6].a/w3082 , \SUBBYTES[6].a/w3081 , \SUBBYTES[6].a/w3065 ,
         \SUBBYTES[6].a/w3064 , \SUBBYTES[6].a/w3063 , \SUBBYTES[6].a/w3062 ,
         \SUBBYTES[6].a/w3061 , \SUBBYTES[6].a/w3059 , \SUBBYTES[6].a/w3058 ,
         \SUBBYTES[6].a/w2986 , \SUBBYTES[6].a/w2984 , \SUBBYTES[6].a/w2983 ,
         \SUBBYTES[6].a/w2982 , \SUBBYTES[6].a/w2979 , \SUBBYTES[6].a/w2977 ,
         \SUBBYTES[6].a/w2976 , \SUBBYTES[6].a/w2975 , \SUBBYTES[6].a/w2971 ,
         \SUBBYTES[6].a/w2969 , \SUBBYTES[6].a/w2968 , \SUBBYTES[6].a/w2967 ,
         \SUBBYTES[6].a/w2966 , \SUBBYTES[6].a/w2965 , \SUBBYTES[6].a/w2964 ,
         \SUBBYTES[6].a/w2963 , \SUBBYTES[6].a/w2962 , \SUBBYTES[6].a/w2954 ,
         \SUBBYTES[6].a/w2952 , \SUBBYTES[6].a/w2951 , \SUBBYTES[6].a/w2947 ,
         \SUBBYTES[6].a/w2945 , \SUBBYTES[6].a/w2944 , \SUBBYTES[6].a/w2943 ,
         \SUBBYTES[6].a/w2939 , \SUBBYTES[6].a/w2937 , \SUBBYTES[6].a/w2936 ,
         \SUBBYTES[6].a/w2923 , \SUBBYTES[6].a/w2922 , \SUBBYTES[6].a/w2921 ,
         \SUBBYTES[6].a/w2919 , \SUBBYTES[6].a/w2916 , \SUBBYTES[6].a/w2915 ,
         \SUBBYTES[6].a/w2913 , \SUBBYTES[6].a/w2912 , \SUBBYTES[6].a/w2910 ,
         \SUBBYTES[6].a/w2908 , \SUBBYTES[6].a/w2907 , \SUBBYTES[6].a/w2901 ,
         \SUBBYTES[6].a/w2900 , \SUBBYTES[6].a/w2899 , \SUBBYTES[6].a/w2898 ,
         \SUBBYTES[6].a/w2892 , \SUBBYTES[6].a/w2890 , \SUBBYTES[6].a/w2889 ,
         \SUBBYTES[6].a/w2885 , \SUBBYTES[6].a/w2883 , \SUBBYTES[6].a/w2882 ,
         \SUBBYTES[6].a/w2877 , \SUBBYTES[6].a/w2875 , \SUBBYTES[6].a/w2874 ,
         \SUBBYTES[6].a/w2858 , \SUBBYTES[6].a/w2857 , \SUBBYTES[6].a/w2856 ,
         \SUBBYTES[6].a/w2855 , \SUBBYTES[6].a/w2854 , \SUBBYTES[6].a/w2852 ,
         \SUBBYTES[6].a/w2851 , \SUBBYTES[6].a/w2779 , \SUBBYTES[6].a/w2777 ,
         \SUBBYTES[6].a/w2776 , \SUBBYTES[6].a/w2775 , \SUBBYTES[6].a/w2772 ,
         \SUBBYTES[6].a/w2770 , \SUBBYTES[6].a/w2769 , \SUBBYTES[6].a/w2768 ,
         \SUBBYTES[6].a/w2764 , \SUBBYTES[6].a/w2762 , \SUBBYTES[6].a/w2761 ,
         \SUBBYTES[6].a/w2760 , \SUBBYTES[6].a/w2759 , \SUBBYTES[6].a/w2758 ,
         \SUBBYTES[6].a/w2757 , \SUBBYTES[6].a/w2756 , \SUBBYTES[6].a/w2755 ,
         \SUBBYTES[6].a/w2747 , \SUBBYTES[6].a/w2745 , \SUBBYTES[6].a/w2744 ,
         \SUBBYTES[6].a/w2740 , \SUBBYTES[6].a/w2738 , \SUBBYTES[6].a/w2737 ,
         \SUBBYTES[6].a/w2736 , \SUBBYTES[6].a/w2732 , \SUBBYTES[6].a/w2730 ,
         \SUBBYTES[6].a/w2729 , \SUBBYTES[6].a/w2716 , \SUBBYTES[6].a/w2715 ,
         \SUBBYTES[6].a/w2714 , \SUBBYTES[6].a/w2712 , \SUBBYTES[6].a/w2709 ,
         \SUBBYTES[6].a/w2708 , \SUBBYTES[6].a/w2706 , \SUBBYTES[6].a/w2705 ,
         \SUBBYTES[6].a/w2703 , \SUBBYTES[6].a/w2701 , \SUBBYTES[6].a/w2700 ,
         \SUBBYTES[6].a/w2694 , \SUBBYTES[6].a/w2693 , \SUBBYTES[6].a/w2692 ,
         \SUBBYTES[6].a/w2691 , \SUBBYTES[6].a/w2685 , \SUBBYTES[6].a/w2683 ,
         \SUBBYTES[6].a/w2682 , \SUBBYTES[6].a/w2678 , \SUBBYTES[6].a/w2676 ,
         \SUBBYTES[6].a/w2675 , \SUBBYTES[6].a/w2670 , \SUBBYTES[6].a/w2668 ,
         \SUBBYTES[6].a/w2667 , \SUBBYTES[6].a/w2651 , \SUBBYTES[6].a/w2650 ,
         \SUBBYTES[6].a/w2649 , \SUBBYTES[6].a/w2648 , \SUBBYTES[6].a/w2647 ,
         \SUBBYTES[6].a/w2645 , \SUBBYTES[6].a/w2644 , \SUBBYTES[6].a/w2572 ,
         \SUBBYTES[6].a/w2570 , \SUBBYTES[6].a/w2569 , \SUBBYTES[6].a/w2568 ,
         \SUBBYTES[6].a/w2565 , \SUBBYTES[6].a/w2563 , \SUBBYTES[6].a/w2562 ,
         \SUBBYTES[6].a/w2561 , \SUBBYTES[6].a/w2557 , \SUBBYTES[6].a/w2555 ,
         \SUBBYTES[6].a/w2554 , \SUBBYTES[6].a/w2553 , \SUBBYTES[6].a/w2552 ,
         \SUBBYTES[6].a/w2551 , \SUBBYTES[6].a/w2550 , \SUBBYTES[6].a/w2549 ,
         \SUBBYTES[6].a/w2548 , \SUBBYTES[6].a/w2540 , \SUBBYTES[6].a/w2538 ,
         \SUBBYTES[6].a/w2537 , \SUBBYTES[6].a/w2533 , \SUBBYTES[6].a/w2531 ,
         \SUBBYTES[6].a/w2530 , \SUBBYTES[6].a/w2529 , \SUBBYTES[6].a/w2525 ,
         \SUBBYTES[6].a/w2523 , \SUBBYTES[6].a/w2522 , \SUBBYTES[6].a/w2509 ,
         \SUBBYTES[6].a/w2508 , \SUBBYTES[6].a/w2507 , \SUBBYTES[6].a/w2505 ,
         \SUBBYTES[6].a/w2502 , \SUBBYTES[6].a/w2501 , \SUBBYTES[6].a/w2499 ,
         \SUBBYTES[6].a/w2498 , \SUBBYTES[6].a/w2496 , \SUBBYTES[6].a/w2494 ,
         \SUBBYTES[6].a/w2493 , \SUBBYTES[6].a/w2487 , \SUBBYTES[6].a/w2486 ,
         \SUBBYTES[6].a/w2485 , \SUBBYTES[6].a/w2484 , \SUBBYTES[6].a/w2478 ,
         \SUBBYTES[6].a/w2476 , \SUBBYTES[6].a/w2475 , \SUBBYTES[6].a/w2471 ,
         \SUBBYTES[6].a/w2469 , \SUBBYTES[6].a/w2468 , \SUBBYTES[6].a/w2463 ,
         \SUBBYTES[6].a/w2461 , \SUBBYTES[6].a/w2460 , \SUBBYTES[6].a/w2444 ,
         \SUBBYTES[6].a/w2443 , \SUBBYTES[6].a/w2442 , \SUBBYTES[6].a/w2441 ,
         \SUBBYTES[6].a/w2440 , \SUBBYTES[6].a/w2438 , \SUBBYTES[6].a/w2437 ,
         \SUBBYTES[6].a/w2365 , \SUBBYTES[6].a/w2363 , \SUBBYTES[6].a/w2362 ,
         \SUBBYTES[6].a/w2361 , \SUBBYTES[6].a/w2358 , \SUBBYTES[6].a/w2356 ,
         \SUBBYTES[6].a/w2355 , \SUBBYTES[6].a/w2354 , \SUBBYTES[6].a/w2350 ,
         \SUBBYTES[6].a/w2348 , \SUBBYTES[6].a/w2347 , \SUBBYTES[6].a/w2346 ,
         \SUBBYTES[6].a/w2345 , \SUBBYTES[6].a/w2344 , \SUBBYTES[6].a/w2343 ,
         \SUBBYTES[6].a/w2342 , \SUBBYTES[6].a/w2341 , \SUBBYTES[6].a/w2333 ,
         \SUBBYTES[6].a/w2331 , \SUBBYTES[6].a/w2330 , \SUBBYTES[6].a/w2326 ,
         \SUBBYTES[6].a/w2324 , \SUBBYTES[6].a/w2323 , \SUBBYTES[6].a/w2322 ,
         \SUBBYTES[6].a/w2318 , \SUBBYTES[6].a/w2316 , \SUBBYTES[6].a/w2315 ,
         \SUBBYTES[6].a/w2302 , \SUBBYTES[6].a/w2301 , \SUBBYTES[6].a/w2300 ,
         \SUBBYTES[6].a/w2298 , \SUBBYTES[6].a/w2295 , \SUBBYTES[6].a/w2294 ,
         \SUBBYTES[6].a/w2292 , \SUBBYTES[6].a/w2291 , \SUBBYTES[6].a/w2289 ,
         \SUBBYTES[6].a/w2287 , \SUBBYTES[6].a/w2286 , \SUBBYTES[6].a/w2280 ,
         \SUBBYTES[6].a/w2279 , \SUBBYTES[6].a/w2278 , \SUBBYTES[6].a/w2277 ,
         \SUBBYTES[6].a/w2271 , \SUBBYTES[6].a/w2269 , \SUBBYTES[6].a/w2268 ,
         \SUBBYTES[6].a/w2264 , \SUBBYTES[6].a/w2262 , \SUBBYTES[6].a/w2261 ,
         \SUBBYTES[6].a/w2256 , \SUBBYTES[6].a/w2254 , \SUBBYTES[6].a/w2253 ,
         \SUBBYTES[6].a/w2237 , \SUBBYTES[6].a/w2236 , \SUBBYTES[6].a/w2235 ,
         \SUBBYTES[6].a/w2234 , \SUBBYTES[6].a/w2233 , \SUBBYTES[6].a/w2231 ,
         \SUBBYTES[6].a/w2230 , \SUBBYTES[6].a/w2158 , \SUBBYTES[6].a/w2156 ,
         \SUBBYTES[6].a/w2155 , \SUBBYTES[6].a/w2154 , \SUBBYTES[6].a/w2151 ,
         \SUBBYTES[6].a/w2149 , \SUBBYTES[6].a/w2148 , \SUBBYTES[6].a/w2147 ,
         \SUBBYTES[6].a/w2143 , \SUBBYTES[6].a/w2141 , \SUBBYTES[6].a/w2140 ,
         \SUBBYTES[6].a/w2139 , \SUBBYTES[6].a/w2138 , \SUBBYTES[6].a/w2137 ,
         \SUBBYTES[6].a/w2136 , \SUBBYTES[6].a/w2135 , \SUBBYTES[6].a/w2134 ,
         \SUBBYTES[6].a/w2126 , \SUBBYTES[6].a/w2124 , \SUBBYTES[6].a/w2123 ,
         \SUBBYTES[6].a/w2119 , \SUBBYTES[6].a/w2117 , \SUBBYTES[6].a/w2116 ,
         \SUBBYTES[6].a/w2115 , \SUBBYTES[6].a/w2111 , \SUBBYTES[6].a/w2109 ,
         \SUBBYTES[6].a/w2108 , \SUBBYTES[6].a/w2095 , \SUBBYTES[6].a/w2094 ,
         \SUBBYTES[6].a/w2093 , \SUBBYTES[6].a/w2091 , \SUBBYTES[6].a/w2088 ,
         \SUBBYTES[6].a/w2087 , \SUBBYTES[6].a/w2085 , \SUBBYTES[6].a/w2084 ,
         \SUBBYTES[6].a/w2082 , \SUBBYTES[6].a/w2080 , \SUBBYTES[6].a/w2079 ,
         \SUBBYTES[6].a/w2073 , \SUBBYTES[6].a/w2072 , \SUBBYTES[6].a/w2071 ,
         \SUBBYTES[6].a/w2070 , \SUBBYTES[6].a/w2064 , \SUBBYTES[6].a/w2062 ,
         \SUBBYTES[6].a/w2061 , \SUBBYTES[6].a/w2057 , \SUBBYTES[6].a/w2055 ,
         \SUBBYTES[6].a/w2054 , \SUBBYTES[6].a/w2049 , \SUBBYTES[6].a/w2047 ,
         \SUBBYTES[6].a/w2046 , \SUBBYTES[6].a/w2030 , \SUBBYTES[6].a/w2029 ,
         \SUBBYTES[6].a/w2028 , \SUBBYTES[6].a/w2027 , \SUBBYTES[6].a/w2026 ,
         \SUBBYTES[6].a/w2024 , \SUBBYTES[6].a/w2023 , \SUBBYTES[6].a/w1951 ,
         \SUBBYTES[6].a/w1949 , \SUBBYTES[6].a/w1948 , \SUBBYTES[6].a/w1947 ,
         \SUBBYTES[6].a/w1944 , \SUBBYTES[6].a/w1942 , \SUBBYTES[6].a/w1941 ,
         \SUBBYTES[6].a/w1940 , \SUBBYTES[6].a/w1936 , \SUBBYTES[6].a/w1934 ,
         \SUBBYTES[6].a/w1933 , \SUBBYTES[6].a/w1932 , \SUBBYTES[6].a/w1931 ,
         \SUBBYTES[6].a/w1930 , \SUBBYTES[6].a/w1929 , \SUBBYTES[6].a/w1928 ,
         \SUBBYTES[6].a/w1927 , \SUBBYTES[6].a/w1919 , \SUBBYTES[6].a/w1917 ,
         \SUBBYTES[6].a/w1916 , \SUBBYTES[6].a/w1912 , \SUBBYTES[6].a/w1910 ,
         \SUBBYTES[6].a/w1909 , \SUBBYTES[6].a/w1908 , \SUBBYTES[6].a/w1904 ,
         \SUBBYTES[6].a/w1902 , \SUBBYTES[6].a/w1901 , \SUBBYTES[6].a/w1888 ,
         \SUBBYTES[6].a/w1887 , \SUBBYTES[6].a/w1886 , \SUBBYTES[6].a/w1884 ,
         \SUBBYTES[6].a/w1881 , \SUBBYTES[6].a/w1880 , \SUBBYTES[6].a/w1878 ,
         \SUBBYTES[6].a/w1877 , \SUBBYTES[6].a/w1875 , \SUBBYTES[6].a/w1873 ,
         \SUBBYTES[6].a/w1872 , \SUBBYTES[6].a/w1866 , \SUBBYTES[6].a/w1865 ,
         \SUBBYTES[6].a/w1864 , \SUBBYTES[6].a/w1863 , \SUBBYTES[6].a/w1857 ,
         \SUBBYTES[6].a/w1855 , \SUBBYTES[6].a/w1854 , \SUBBYTES[6].a/w1850 ,
         \SUBBYTES[6].a/w1848 , \SUBBYTES[6].a/w1847 , \SUBBYTES[6].a/w1842 ,
         \SUBBYTES[6].a/w1840 , \SUBBYTES[6].a/w1839 , \SUBBYTES[6].a/w1823 ,
         \SUBBYTES[6].a/w1822 , \SUBBYTES[6].a/w1821 , \SUBBYTES[6].a/w1820 ,
         \SUBBYTES[6].a/w1819 , \SUBBYTES[6].a/w1817 , \SUBBYTES[6].a/w1816 ,
         \SUBBYTES[6].a/w1744 , \SUBBYTES[6].a/w1742 , \SUBBYTES[6].a/w1741 ,
         \SUBBYTES[6].a/w1740 , \SUBBYTES[6].a/w1737 , \SUBBYTES[6].a/w1735 ,
         \SUBBYTES[6].a/w1734 , \SUBBYTES[6].a/w1733 , \SUBBYTES[6].a/w1729 ,
         \SUBBYTES[6].a/w1727 , \SUBBYTES[6].a/w1726 , \SUBBYTES[6].a/w1725 ,
         \SUBBYTES[6].a/w1724 , \SUBBYTES[6].a/w1723 , \SUBBYTES[6].a/w1722 ,
         \SUBBYTES[6].a/w1721 , \SUBBYTES[6].a/w1720 , \SUBBYTES[6].a/w1712 ,
         \SUBBYTES[6].a/w1710 , \SUBBYTES[6].a/w1709 , \SUBBYTES[6].a/w1705 ,
         \SUBBYTES[6].a/w1703 , \SUBBYTES[6].a/w1702 , \SUBBYTES[6].a/w1701 ,
         \SUBBYTES[6].a/w1697 , \SUBBYTES[6].a/w1695 , \SUBBYTES[6].a/w1694 ,
         \SUBBYTES[6].a/w1681 , \SUBBYTES[6].a/w1680 , \SUBBYTES[6].a/w1679 ,
         \SUBBYTES[6].a/w1677 , \SUBBYTES[6].a/w1674 , \SUBBYTES[6].a/w1673 ,
         \SUBBYTES[6].a/w1671 , \SUBBYTES[6].a/w1670 , \SUBBYTES[6].a/w1668 ,
         \SUBBYTES[6].a/w1666 , \SUBBYTES[6].a/w1665 , \SUBBYTES[6].a/w1659 ,
         \SUBBYTES[6].a/w1658 , \SUBBYTES[6].a/w1657 , \SUBBYTES[6].a/w1656 ,
         \SUBBYTES[6].a/w1650 , \SUBBYTES[6].a/w1648 , \SUBBYTES[6].a/w1647 ,
         \SUBBYTES[6].a/w1643 , \SUBBYTES[6].a/w1641 , \SUBBYTES[6].a/w1640 ,
         \SUBBYTES[6].a/w1635 , \SUBBYTES[6].a/w1633 , \SUBBYTES[6].a/w1632 ,
         \SUBBYTES[6].a/w1616 , \SUBBYTES[6].a/w1615 , \SUBBYTES[6].a/w1614 ,
         \SUBBYTES[6].a/w1613 , \SUBBYTES[6].a/w1612 , \SUBBYTES[6].a/w1610 ,
         \SUBBYTES[6].a/w1609 , \SUBBYTES[6].a/w1537 , \SUBBYTES[6].a/w1535 ,
         \SUBBYTES[6].a/w1534 , \SUBBYTES[6].a/w1533 , \SUBBYTES[6].a/w1530 ,
         \SUBBYTES[6].a/w1528 , \SUBBYTES[6].a/w1527 , \SUBBYTES[6].a/w1526 ,
         \SUBBYTES[6].a/w1522 , \SUBBYTES[6].a/w1520 , \SUBBYTES[6].a/w1519 ,
         \SUBBYTES[6].a/w1518 , \SUBBYTES[6].a/w1517 , \SUBBYTES[6].a/w1516 ,
         \SUBBYTES[6].a/w1515 , \SUBBYTES[6].a/w1514 , \SUBBYTES[6].a/w1513 ,
         \SUBBYTES[6].a/w1505 , \SUBBYTES[6].a/w1503 , \SUBBYTES[6].a/w1502 ,
         \SUBBYTES[6].a/w1498 , \SUBBYTES[6].a/w1496 , \SUBBYTES[6].a/w1495 ,
         \SUBBYTES[6].a/w1494 , \SUBBYTES[6].a/w1490 , \SUBBYTES[6].a/w1488 ,
         \SUBBYTES[6].a/w1487 , \SUBBYTES[6].a/w1474 , \SUBBYTES[6].a/w1473 ,
         \SUBBYTES[6].a/w1472 , \SUBBYTES[6].a/w1470 , \SUBBYTES[6].a/w1467 ,
         \SUBBYTES[6].a/w1466 , \SUBBYTES[6].a/w1464 , \SUBBYTES[6].a/w1463 ,
         \SUBBYTES[6].a/w1461 , \SUBBYTES[6].a/w1459 , \SUBBYTES[6].a/w1458 ,
         \SUBBYTES[6].a/w1452 , \SUBBYTES[6].a/w1451 , \SUBBYTES[6].a/w1450 ,
         \SUBBYTES[6].a/w1449 , \SUBBYTES[6].a/w1443 , \SUBBYTES[6].a/w1441 ,
         \SUBBYTES[6].a/w1440 , \SUBBYTES[6].a/w1436 , \SUBBYTES[6].a/w1434 ,
         \SUBBYTES[6].a/w1433 , \SUBBYTES[6].a/w1428 , \SUBBYTES[6].a/w1426 ,
         \SUBBYTES[6].a/w1425 , \SUBBYTES[6].a/w1409 , \SUBBYTES[6].a/w1408 ,
         \SUBBYTES[6].a/w1407 , \SUBBYTES[6].a/w1406 , \SUBBYTES[6].a/w1405 ,
         \SUBBYTES[6].a/w1403 , \SUBBYTES[6].a/w1402 , \SUBBYTES[6].a/w1330 ,
         \SUBBYTES[6].a/w1328 , \SUBBYTES[6].a/w1327 , \SUBBYTES[6].a/w1326 ,
         \SUBBYTES[6].a/w1323 , \SUBBYTES[6].a/w1321 , \SUBBYTES[6].a/w1320 ,
         \SUBBYTES[6].a/w1319 , \SUBBYTES[6].a/w1315 , \SUBBYTES[6].a/w1313 ,
         \SUBBYTES[6].a/w1312 , \SUBBYTES[6].a/w1311 , \SUBBYTES[6].a/w1310 ,
         \SUBBYTES[6].a/w1309 , \SUBBYTES[6].a/w1308 , \SUBBYTES[6].a/w1307 ,
         \SUBBYTES[6].a/w1306 , \SUBBYTES[6].a/w1298 , \SUBBYTES[6].a/w1296 ,
         \SUBBYTES[6].a/w1295 , \SUBBYTES[6].a/w1291 , \SUBBYTES[6].a/w1289 ,
         \SUBBYTES[6].a/w1288 , \SUBBYTES[6].a/w1287 , \SUBBYTES[6].a/w1283 ,
         \SUBBYTES[6].a/w1281 , \SUBBYTES[6].a/w1280 , \SUBBYTES[6].a/w1267 ,
         \SUBBYTES[6].a/w1266 , \SUBBYTES[6].a/w1265 , \SUBBYTES[6].a/w1263 ,
         \SUBBYTES[6].a/w1260 , \SUBBYTES[6].a/w1259 , \SUBBYTES[6].a/w1257 ,
         \SUBBYTES[6].a/w1256 , \SUBBYTES[6].a/w1254 , \SUBBYTES[6].a/w1252 ,
         \SUBBYTES[6].a/w1251 , \SUBBYTES[6].a/w1245 , \SUBBYTES[6].a/w1244 ,
         \SUBBYTES[6].a/w1243 , \SUBBYTES[6].a/w1242 , \SUBBYTES[6].a/w1236 ,
         \SUBBYTES[6].a/w1234 , \SUBBYTES[6].a/w1233 , \SUBBYTES[6].a/w1229 ,
         \SUBBYTES[6].a/w1227 , \SUBBYTES[6].a/w1226 , \SUBBYTES[6].a/w1221 ,
         \SUBBYTES[6].a/w1219 , \SUBBYTES[6].a/w1218 , \SUBBYTES[6].a/w1202 ,
         \SUBBYTES[6].a/w1201 , \SUBBYTES[6].a/w1200 , \SUBBYTES[6].a/w1199 ,
         \SUBBYTES[6].a/w1198 , \SUBBYTES[6].a/w1196 , \SUBBYTES[6].a/w1195 ,
         \SUBBYTES[6].a/w1123 , \SUBBYTES[6].a/w1121 , \SUBBYTES[6].a/w1120 ,
         \SUBBYTES[6].a/w1119 , \SUBBYTES[6].a/w1116 , \SUBBYTES[6].a/w1114 ,
         \SUBBYTES[6].a/w1113 , \SUBBYTES[6].a/w1112 , \SUBBYTES[6].a/w1108 ,
         \SUBBYTES[6].a/w1106 , \SUBBYTES[6].a/w1105 , \SUBBYTES[6].a/w1104 ,
         \SUBBYTES[6].a/w1103 , \SUBBYTES[6].a/w1102 , \SUBBYTES[6].a/w1101 ,
         \SUBBYTES[6].a/w1100 , \SUBBYTES[6].a/w1099 , \SUBBYTES[6].a/w1091 ,
         \SUBBYTES[6].a/w1089 , \SUBBYTES[6].a/w1088 , \SUBBYTES[6].a/w1084 ,
         \SUBBYTES[6].a/w1082 , \SUBBYTES[6].a/w1081 , \SUBBYTES[6].a/w1080 ,
         \SUBBYTES[6].a/w1076 , \SUBBYTES[6].a/w1074 , \SUBBYTES[6].a/w1073 ,
         \SUBBYTES[6].a/w1060 , \SUBBYTES[6].a/w1059 , \SUBBYTES[6].a/w1058 ,
         \SUBBYTES[6].a/w1056 , \SUBBYTES[6].a/w1053 , \SUBBYTES[6].a/w1052 ,
         \SUBBYTES[6].a/w1050 , \SUBBYTES[6].a/w1049 , \SUBBYTES[6].a/w1047 ,
         \SUBBYTES[6].a/w1045 , \SUBBYTES[6].a/w1044 , \SUBBYTES[6].a/w1038 ,
         \SUBBYTES[6].a/w1037 , \SUBBYTES[6].a/w1036 , \SUBBYTES[6].a/w1035 ,
         \SUBBYTES[6].a/w1029 , \SUBBYTES[6].a/w1027 , \SUBBYTES[6].a/w1026 ,
         \SUBBYTES[6].a/w1022 , \SUBBYTES[6].a/w1020 , \SUBBYTES[6].a/w1019 ,
         \SUBBYTES[6].a/w1014 , \SUBBYTES[6].a/w1012 , \SUBBYTES[6].a/w1011 ,
         \SUBBYTES[6].a/w995 , \SUBBYTES[6].a/w994 , \SUBBYTES[6].a/w993 ,
         \SUBBYTES[6].a/w992 , \SUBBYTES[6].a/w991 , \SUBBYTES[6].a/w989 ,
         \SUBBYTES[6].a/w988 , \SUBBYTES[6].a/w916 , \SUBBYTES[6].a/w914 ,
         \SUBBYTES[6].a/w913 , \SUBBYTES[6].a/w912 , \SUBBYTES[6].a/w909 ,
         \SUBBYTES[6].a/w907 , \SUBBYTES[6].a/w906 , \SUBBYTES[6].a/w905 ,
         \SUBBYTES[6].a/w901 , \SUBBYTES[6].a/w899 , \SUBBYTES[6].a/w898 ,
         \SUBBYTES[6].a/w897 , \SUBBYTES[6].a/w896 , \SUBBYTES[6].a/w895 ,
         \SUBBYTES[6].a/w894 , \SUBBYTES[6].a/w893 , \SUBBYTES[6].a/w892 ,
         \SUBBYTES[6].a/w884 , \SUBBYTES[6].a/w882 , \SUBBYTES[6].a/w881 ,
         \SUBBYTES[6].a/w877 , \SUBBYTES[6].a/w875 , \SUBBYTES[6].a/w874 ,
         \SUBBYTES[6].a/w873 , \SUBBYTES[6].a/w869 , \SUBBYTES[6].a/w867 ,
         \SUBBYTES[6].a/w866 , \SUBBYTES[6].a/w853 , \SUBBYTES[6].a/w852 ,
         \SUBBYTES[6].a/w851 , \SUBBYTES[6].a/w849 , \SUBBYTES[6].a/w846 ,
         \SUBBYTES[6].a/w845 , \SUBBYTES[6].a/w843 , \SUBBYTES[6].a/w842 ,
         \SUBBYTES[6].a/w840 , \SUBBYTES[6].a/w838 , \SUBBYTES[6].a/w837 ,
         \SUBBYTES[6].a/w831 , \SUBBYTES[6].a/w830 , \SUBBYTES[6].a/w829 ,
         \SUBBYTES[6].a/w828 , \SUBBYTES[6].a/w822 , \SUBBYTES[6].a/w820 ,
         \SUBBYTES[6].a/w819 , \SUBBYTES[6].a/w815 , \SUBBYTES[6].a/w813 ,
         \SUBBYTES[6].a/w812 , \SUBBYTES[6].a/w807 , \SUBBYTES[6].a/w805 ,
         \SUBBYTES[6].a/w804 , \SUBBYTES[6].a/w788 , \SUBBYTES[6].a/w787 ,
         \SUBBYTES[6].a/w786 , \SUBBYTES[6].a/w785 , \SUBBYTES[6].a/w784 ,
         \SUBBYTES[6].a/w782 , \SUBBYTES[6].a/w781 , \SUBBYTES[6].a/w709 ,
         \SUBBYTES[6].a/w707 , \SUBBYTES[6].a/w706 , \SUBBYTES[6].a/w705 ,
         \SUBBYTES[6].a/w702 , \SUBBYTES[6].a/w700 , \SUBBYTES[6].a/w699 ,
         \SUBBYTES[6].a/w698 , \SUBBYTES[6].a/w694 , \SUBBYTES[6].a/w692 ,
         \SUBBYTES[6].a/w691 , \SUBBYTES[6].a/w690 , \SUBBYTES[6].a/w689 ,
         \SUBBYTES[6].a/w688 , \SUBBYTES[6].a/w687 , \SUBBYTES[6].a/w686 ,
         \SUBBYTES[6].a/w685 , \SUBBYTES[6].a/w677 , \SUBBYTES[6].a/w675 ,
         \SUBBYTES[6].a/w674 , \SUBBYTES[6].a/w670 , \SUBBYTES[6].a/w668 ,
         \SUBBYTES[6].a/w667 , \SUBBYTES[6].a/w666 , \SUBBYTES[6].a/w662 ,
         \SUBBYTES[6].a/w660 , \SUBBYTES[6].a/w659 , \SUBBYTES[6].a/w646 ,
         \SUBBYTES[6].a/w645 , \SUBBYTES[6].a/w644 , \SUBBYTES[6].a/w642 ,
         \SUBBYTES[6].a/w639 , \SUBBYTES[6].a/w638 , \SUBBYTES[6].a/w636 ,
         \SUBBYTES[6].a/w635 , \SUBBYTES[6].a/w633 , \SUBBYTES[6].a/w631 ,
         \SUBBYTES[6].a/w630 , \SUBBYTES[6].a/w624 , \SUBBYTES[6].a/w623 ,
         \SUBBYTES[6].a/w622 , \SUBBYTES[6].a/w621 , \SUBBYTES[6].a/w615 ,
         \SUBBYTES[6].a/w613 , \SUBBYTES[6].a/w612 , \SUBBYTES[6].a/w608 ,
         \SUBBYTES[6].a/w606 , \SUBBYTES[6].a/w605 , \SUBBYTES[6].a/w600 ,
         \SUBBYTES[6].a/w598 , \SUBBYTES[6].a/w597 , \SUBBYTES[6].a/w581 ,
         \SUBBYTES[6].a/w580 , \SUBBYTES[6].a/w579 , \SUBBYTES[6].a/w578 ,
         \SUBBYTES[6].a/w577 , \SUBBYTES[6].a/w575 , \SUBBYTES[6].a/w574 ,
         \SUBBYTES[6].a/w502 , \SUBBYTES[6].a/w500 , \SUBBYTES[6].a/w499 ,
         \SUBBYTES[6].a/w498 , \SUBBYTES[6].a/w495 , \SUBBYTES[6].a/w493 ,
         \SUBBYTES[6].a/w492 , \SUBBYTES[6].a/w491 , \SUBBYTES[6].a/w487 ,
         \SUBBYTES[6].a/w485 , \SUBBYTES[6].a/w484 , \SUBBYTES[6].a/w483 ,
         \SUBBYTES[6].a/w482 , \SUBBYTES[6].a/w481 , \SUBBYTES[6].a/w480 ,
         \SUBBYTES[6].a/w479 , \SUBBYTES[6].a/w478 , \SUBBYTES[6].a/w470 ,
         \SUBBYTES[6].a/w468 , \SUBBYTES[6].a/w467 , \SUBBYTES[6].a/w463 ,
         \SUBBYTES[6].a/w461 , \SUBBYTES[6].a/w460 , \SUBBYTES[6].a/w459 ,
         \SUBBYTES[6].a/w455 , \SUBBYTES[6].a/w453 , \SUBBYTES[6].a/w452 ,
         \SUBBYTES[6].a/w439 , \SUBBYTES[6].a/w438 , \SUBBYTES[6].a/w437 ,
         \SUBBYTES[6].a/w435 , \SUBBYTES[6].a/w432 , \SUBBYTES[6].a/w431 ,
         \SUBBYTES[6].a/w429 , \SUBBYTES[6].a/w428 , \SUBBYTES[6].a/w426 ,
         \SUBBYTES[6].a/w424 , \SUBBYTES[6].a/w423 , \SUBBYTES[6].a/w417 ,
         \SUBBYTES[6].a/w416 , \SUBBYTES[6].a/w415 , \SUBBYTES[6].a/w414 ,
         \SUBBYTES[6].a/w408 , \SUBBYTES[6].a/w406 , \SUBBYTES[6].a/w405 ,
         \SUBBYTES[6].a/w401 , \SUBBYTES[6].a/w399 , \SUBBYTES[6].a/w398 ,
         \SUBBYTES[6].a/w393 , \SUBBYTES[6].a/w391 , \SUBBYTES[6].a/w390 ,
         \SUBBYTES[6].a/w374 , \SUBBYTES[6].a/w373 , \SUBBYTES[6].a/w372 ,
         \SUBBYTES[6].a/w371 , \SUBBYTES[6].a/w370 , \SUBBYTES[6].a/w368 ,
         \SUBBYTES[6].a/w367 , \SUBBYTES[6].a/w295 , \SUBBYTES[6].a/w293 ,
         \SUBBYTES[6].a/w292 , \SUBBYTES[6].a/w291 , \SUBBYTES[6].a/w288 ,
         \SUBBYTES[6].a/w286 , \SUBBYTES[6].a/w285 , \SUBBYTES[6].a/w284 ,
         \SUBBYTES[6].a/w280 , \SUBBYTES[6].a/w278 , \SUBBYTES[6].a/w277 ,
         \SUBBYTES[6].a/w276 , \SUBBYTES[6].a/w275 , \SUBBYTES[6].a/w274 ,
         \SUBBYTES[6].a/w273 , \SUBBYTES[6].a/w272 , \SUBBYTES[6].a/w271 ,
         \SUBBYTES[6].a/w263 , \SUBBYTES[6].a/w261 , \SUBBYTES[6].a/w260 ,
         \SUBBYTES[6].a/w256 , \SUBBYTES[6].a/w254 , \SUBBYTES[6].a/w253 ,
         \SUBBYTES[6].a/w252 , \SUBBYTES[6].a/w248 , \SUBBYTES[6].a/w246 ,
         \SUBBYTES[6].a/w245 , \SUBBYTES[6].a/w232 , \SUBBYTES[6].a/w231 ,
         \SUBBYTES[6].a/w230 , \SUBBYTES[6].a/w228 , \SUBBYTES[6].a/w225 ,
         \SUBBYTES[6].a/w224 , \SUBBYTES[6].a/w222 , \SUBBYTES[6].a/w221 ,
         \SUBBYTES[6].a/w219 , \SUBBYTES[6].a/w217 , \SUBBYTES[6].a/w216 ,
         \SUBBYTES[6].a/w210 , \SUBBYTES[6].a/w209 , \SUBBYTES[6].a/w208 ,
         \SUBBYTES[6].a/w207 , \SUBBYTES[6].a/w201 , \SUBBYTES[6].a/w199 ,
         \SUBBYTES[6].a/w198 , \SUBBYTES[6].a/w194 , \SUBBYTES[6].a/w192 ,
         \SUBBYTES[6].a/w191 , \SUBBYTES[6].a/w186 , \SUBBYTES[6].a/w184 ,
         \SUBBYTES[6].a/w183 , \SUBBYTES[6].a/w167 , \SUBBYTES[6].a/w166 ,
         \SUBBYTES[6].a/w165 , \SUBBYTES[6].a/w164 , \SUBBYTES[6].a/w163 ,
         \SUBBYTES[6].a/w161 , \SUBBYTES[6].a/w160 , \SUBBYTES[5].a/w3400 ,
         \SUBBYTES[5].a/w3398 , \SUBBYTES[5].a/w3397 , \SUBBYTES[5].a/w3396 ,
         \SUBBYTES[5].a/w3393 , \SUBBYTES[5].a/w3391 , \SUBBYTES[5].a/w3390 ,
         \SUBBYTES[5].a/w3389 , \SUBBYTES[5].a/w3385 , \SUBBYTES[5].a/w3383 ,
         \SUBBYTES[5].a/w3382 , \SUBBYTES[5].a/w3381 , \SUBBYTES[5].a/w3380 ,
         \SUBBYTES[5].a/w3379 , \SUBBYTES[5].a/w3378 , \SUBBYTES[5].a/w3377 ,
         \SUBBYTES[5].a/w3376 , \SUBBYTES[5].a/w3368 , \SUBBYTES[5].a/w3366 ,
         \SUBBYTES[5].a/w3365 , \SUBBYTES[5].a/w3361 , \SUBBYTES[5].a/w3359 ,
         \SUBBYTES[5].a/w3358 , \SUBBYTES[5].a/w3357 , \SUBBYTES[5].a/w3353 ,
         \SUBBYTES[5].a/w3351 , \SUBBYTES[5].a/w3350 , \SUBBYTES[5].a/w3337 ,
         \SUBBYTES[5].a/w3336 , \SUBBYTES[5].a/w3335 , \SUBBYTES[5].a/w3333 ,
         \SUBBYTES[5].a/w3330 , \SUBBYTES[5].a/w3329 , \SUBBYTES[5].a/w3327 ,
         \SUBBYTES[5].a/w3326 , \SUBBYTES[5].a/w3324 , \SUBBYTES[5].a/w3322 ,
         \SUBBYTES[5].a/w3321 , \SUBBYTES[5].a/w3315 , \SUBBYTES[5].a/w3314 ,
         \SUBBYTES[5].a/w3313 , \SUBBYTES[5].a/w3312 , \SUBBYTES[5].a/w3306 ,
         \SUBBYTES[5].a/w3304 , \SUBBYTES[5].a/w3303 , \SUBBYTES[5].a/w3299 ,
         \SUBBYTES[5].a/w3297 , \SUBBYTES[5].a/w3296 , \SUBBYTES[5].a/w3291 ,
         \SUBBYTES[5].a/w3289 , \SUBBYTES[5].a/w3288 , \SUBBYTES[5].a/w3272 ,
         \SUBBYTES[5].a/w3271 , \SUBBYTES[5].a/w3270 , \SUBBYTES[5].a/w3269 ,
         \SUBBYTES[5].a/w3268 , \SUBBYTES[5].a/w3266 , \SUBBYTES[5].a/w3265 ,
         \SUBBYTES[5].a/w3193 , \SUBBYTES[5].a/w3191 , \SUBBYTES[5].a/w3190 ,
         \SUBBYTES[5].a/w3189 , \SUBBYTES[5].a/w3186 , \SUBBYTES[5].a/w3184 ,
         \SUBBYTES[5].a/w3183 , \SUBBYTES[5].a/w3182 , \SUBBYTES[5].a/w3178 ,
         \SUBBYTES[5].a/w3176 , \SUBBYTES[5].a/w3175 , \SUBBYTES[5].a/w3174 ,
         \SUBBYTES[5].a/w3173 , \SUBBYTES[5].a/w3172 , \SUBBYTES[5].a/w3171 ,
         \SUBBYTES[5].a/w3170 , \SUBBYTES[5].a/w3169 , \SUBBYTES[5].a/w3161 ,
         \SUBBYTES[5].a/w3159 , \SUBBYTES[5].a/w3158 , \SUBBYTES[5].a/w3154 ,
         \SUBBYTES[5].a/w3152 , \SUBBYTES[5].a/w3151 , \SUBBYTES[5].a/w3150 ,
         \SUBBYTES[5].a/w3146 , \SUBBYTES[5].a/w3144 , \SUBBYTES[5].a/w3143 ,
         \SUBBYTES[5].a/w3130 , \SUBBYTES[5].a/w3129 , \SUBBYTES[5].a/w3128 ,
         \SUBBYTES[5].a/w3126 , \SUBBYTES[5].a/w3123 , \SUBBYTES[5].a/w3122 ,
         \SUBBYTES[5].a/w3120 , \SUBBYTES[5].a/w3119 , \SUBBYTES[5].a/w3117 ,
         \SUBBYTES[5].a/w3115 , \SUBBYTES[5].a/w3114 , \SUBBYTES[5].a/w3108 ,
         \SUBBYTES[5].a/w3107 , \SUBBYTES[5].a/w3106 , \SUBBYTES[5].a/w3105 ,
         \SUBBYTES[5].a/w3099 , \SUBBYTES[5].a/w3097 , \SUBBYTES[5].a/w3096 ,
         \SUBBYTES[5].a/w3092 , \SUBBYTES[5].a/w3090 , \SUBBYTES[5].a/w3089 ,
         \SUBBYTES[5].a/w3084 , \SUBBYTES[5].a/w3082 , \SUBBYTES[5].a/w3081 ,
         \SUBBYTES[5].a/w3065 , \SUBBYTES[5].a/w3064 , \SUBBYTES[5].a/w3063 ,
         \SUBBYTES[5].a/w3062 , \SUBBYTES[5].a/w3061 , \SUBBYTES[5].a/w3059 ,
         \SUBBYTES[5].a/w3058 , \SUBBYTES[5].a/w2986 , \SUBBYTES[5].a/w2984 ,
         \SUBBYTES[5].a/w2983 , \SUBBYTES[5].a/w2982 , \SUBBYTES[5].a/w2979 ,
         \SUBBYTES[5].a/w2977 , \SUBBYTES[5].a/w2976 , \SUBBYTES[5].a/w2975 ,
         \SUBBYTES[5].a/w2971 , \SUBBYTES[5].a/w2969 , \SUBBYTES[5].a/w2968 ,
         \SUBBYTES[5].a/w2967 , \SUBBYTES[5].a/w2966 , \SUBBYTES[5].a/w2965 ,
         \SUBBYTES[5].a/w2964 , \SUBBYTES[5].a/w2963 , \SUBBYTES[5].a/w2962 ,
         \SUBBYTES[5].a/w2954 , \SUBBYTES[5].a/w2952 , \SUBBYTES[5].a/w2951 ,
         \SUBBYTES[5].a/w2947 , \SUBBYTES[5].a/w2945 , \SUBBYTES[5].a/w2944 ,
         \SUBBYTES[5].a/w2943 , \SUBBYTES[5].a/w2939 , \SUBBYTES[5].a/w2937 ,
         \SUBBYTES[5].a/w2936 , \SUBBYTES[5].a/w2923 , \SUBBYTES[5].a/w2922 ,
         \SUBBYTES[5].a/w2921 , \SUBBYTES[5].a/w2919 , \SUBBYTES[5].a/w2916 ,
         \SUBBYTES[5].a/w2915 , \SUBBYTES[5].a/w2913 , \SUBBYTES[5].a/w2912 ,
         \SUBBYTES[5].a/w2910 , \SUBBYTES[5].a/w2908 , \SUBBYTES[5].a/w2907 ,
         \SUBBYTES[5].a/w2901 , \SUBBYTES[5].a/w2900 , \SUBBYTES[5].a/w2899 ,
         \SUBBYTES[5].a/w2898 , \SUBBYTES[5].a/w2892 , \SUBBYTES[5].a/w2890 ,
         \SUBBYTES[5].a/w2889 , \SUBBYTES[5].a/w2885 , \SUBBYTES[5].a/w2883 ,
         \SUBBYTES[5].a/w2882 , \SUBBYTES[5].a/w2877 , \SUBBYTES[5].a/w2875 ,
         \SUBBYTES[5].a/w2874 , \SUBBYTES[5].a/w2858 , \SUBBYTES[5].a/w2857 ,
         \SUBBYTES[5].a/w2856 , \SUBBYTES[5].a/w2855 , \SUBBYTES[5].a/w2854 ,
         \SUBBYTES[5].a/w2852 , \SUBBYTES[5].a/w2851 , \SUBBYTES[5].a/w2779 ,
         \SUBBYTES[5].a/w2777 , \SUBBYTES[5].a/w2776 , \SUBBYTES[5].a/w2775 ,
         \SUBBYTES[5].a/w2772 , \SUBBYTES[5].a/w2770 , \SUBBYTES[5].a/w2769 ,
         \SUBBYTES[5].a/w2768 , \SUBBYTES[5].a/w2764 , \SUBBYTES[5].a/w2762 ,
         \SUBBYTES[5].a/w2761 , \SUBBYTES[5].a/w2760 , \SUBBYTES[5].a/w2759 ,
         \SUBBYTES[5].a/w2758 , \SUBBYTES[5].a/w2757 , \SUBBYTES[5].a/w2756 ,
         \SUBBYTES[5].a/w2755 , \SUBBYTES[5].a/w2747 , \SUBBYTES[5].a/w2745 ,
         \SUBBYTES[5].a/w2744 , \SUBBYTES[5].a/w2740 , \SUBBYTES[5].a/w2738 ,
         \SUBBYTES[5].a/w2737 , \SUBBYTES[5].a/w2736 , \SUBBYTES[5].a/w2732 ,
         \SUBBYTES[5].a/w2730 , \SUBBYTES[5].a/w2729 , \SUBBYTES[5].a/w2716 ,
         \SUBBYTES[5].a/w2715 , \SUBBYTES[5].a/w2714 , \SUBBYTES[5].a/w2712 ,
         \SUBBYTES[5].a/w2709 , \SUBBYTES[5].a/w2708 , \SUBBYTES[5].a/w2706 ,
         \SUBBYTES[5].a/w2705 , \SUBBYTES[5].a/w2703 , \SUBBYTES[5].a/w2701 ,
         \SUBBYTES[5].a/w2700 , \SUBBYTES[5].a/w2694 , \SUBBYTES[5].a/w2693 ,
         \SUBBYTES[5].a/w2692 , \SUBBYTES[5].a/w2691 , \SUBBYTES[5].a/w2685 ,
         \SUBBYTES[5].a/w2683 , \SUBBYTES[5].a/w2682 , \SUBBYTES[5].a/w2678 ,
         \SUBBYTES[5].a/w2676 , \SUBBYTES[5].a/w2675 , \SUBBYTES[5].a/w2670 ,
         \SUBBYTES[5].a/w2668 , \SUBBYTES[5].a/w2667 , \SUBBYTES[5].a/w2651 ,
         \SUBBYTES[5].a/w2650 , \SUBBYTES[5].a/w2649 , \SUBBYTES[5].a/w2648 ,
         \SUBBYTES[5].a/w2647 , \SUBBYTES[5].a/w2645 , \SUBBYTES[5].a/w2644 ,
         \SUBBYTES[5].a/w2572 , \SUBBYTES[5].a/w2570 , \SUBBYTES[5].a/w2569 ,
         \SUBBYTES[5].a/w2568 , \SUBBYTES[5].a/w2565 , \SUBBYTES[5].a/w2563 ,
         \SUBBYTES[5].a/w2562 , \SUBBYTES[5].a/w2561 , \SUBBYTES[5].a/w2557 ,
         \SUBBYTES[5].a/w2555 , \SUBBYTES[5].a/w2554 , \SUBBYTES[5].a/w2553 ,
         \SUBBYTES[5].a/w2552 , \SUBBYTES[5].a/w2551 , \SUBBYTES[5].a/w2550 ,
         \SUBBYTES[5].a/w2549 , \SUBBYTES[5].a/w2548 , \SUBBYTES[5].a/w2540 ,
         \SUBBYTES[5].a/w2538 , \SUBBYTES[5].a/w2537 , \SUBBYTES[5].a/w2533 ,
         \SUBBYTES[5].a/w2531 , \SUBBYTES[5].a/w2530 , \SUBBYTES[5].a/w2529 ,
         \SUBBYTES[5].a/w2525 , \SUBBYTES[5].a/w2523 , \SUBBYTES[5].a/w2522 ,
         \SUBBYTES[5].a/w2509 , \SUBBYTES[5].a/w2508 , \SUBBYTES[5].a/w2507 ,
         \SUBBYTES[5].a/w2505 , \SUBBYTES[5].a/w2502 , \SUBBYTES[5].a/w2501 ,
         \SUBBYTES[5].a/w2499 , \SUBBYTES[5].a/w2498 , \SUBBYTES[5].a/w2496 ,
         \SUBBYTES[5].a/w2494 , \SUBBYTES[5].a/w2493 , \SUBBYTES[5].a/w2487 ,
         \SUBBYTES[5].a/w2486 , \SUBBYTES[5].a/w2485 , \SUBBYTES[5].a/w2484 ,
         \SUBBYTES[5].a/w2478 , \SUBBYTES[5].a/w2476 , \SUBBYTES[5].a/w2475 ,
         \SUBBYTES[5].a/w2471 , \SUBBYTES[5].a/w2469 , \SUBBYTES[5].a/w2468 ,
         \SUBBYTES[5].a/w2463 , \SUBBYTES[5].a/w2461 , \SUBBYTES[5].a/w2460 ,
         \SUBBYTES[5].a/w2444 , \SUBBYTES[5].a/w2443 , \SUBBYTES[5].a/w2442 ,
         \SUBBYTES[5].a/w2441 , \SUBBYTES[5].a/w2440 , \SUBBYTES[5].a/w2438 ,
         \SUBBYTES[5].a/w2437 , \SUBBYTES[5].a/w2365 , \SUBBYTES[5].a/w2363 ,
         \SUBBYTES[5].a/w2362 , \SUBBYTES[5].a/w2361 , \SUBBYTES[5].a/w2358 ,
         \SUBBYTES[5].a/w2356 , \SUBBYTES[5].a/w2355 , \SUBBYTES[5].a/w2354 ,
         \SUBBYTES[5].a/w2350 , \SUBBYTES[5].a/w2348 , \SUBBYTES[5].a/w2347 ,
         \SUBBYTES[5].a/w2346 , \SUBBYTES[5].a/w2345 , \SUBBYTES[5].a/w2344 ,
         \SUBBYTES[5].a/w2343 , \SUBBYTES[5].a/w2342 , \SUBBYTES[5].a/w2341 ,
         \SUBBYTES[5].a/w2333 , \SUBBYTES[5].a/w2331 , \SUBBYTES[5].a/w2330 ,
         \SUBBYTES[5].a/w2326 , \SUBBYTES[5].a/w2324 , \SUBBYTES[5].a/w2323 ,
         \SUBBYTES[5].a/w2322 , \SUBBYTES[5].a/w2318 , \SUBBYTES[5].a/w2316 ,
         \SUBBYTES[5].a/w2315 , \SUBBYTES[5].a/w2302 , \SUBBYTES[5].a/w2301 ,
         \SUBBYTES[5].a/w2300 , \SUBBYTES[5].a/w2298 , \SUBBYTES[5].a/w2295 ,
         \SUBBYTES[5].a/w2294 , \SUBBYTES[5].a/w2292 , \SUBBYTES[5].a/w2291 ,
         \SUBBYTES[5].a/w2289 , \SUBBYTES[5].a/w2287 , \SUBBYTES[5].a/w2286 ,
         \SUBBYTES[5].a/w2280 , \SUBBYTES[5].a/w2279 , \SUBBYTES[5].a/w2278 ,
         \SUBBYTES[5].a/w2277 , \SUBBYTES[5].a/w2271 , \SUBBYTES[5].a/w2269 ,
         \SUBBYTES[5].a/w2268 , \SUBBYTES[5].a/w2264 , \SUBBYTES[5].a/w2262 ,
         \SUBBYTES[5].a/w2261 , \SUBBYTES[5].a/w2256 , \SUBBYTES[5].a/w2254 ,
         \SUBBYTES[5].a/w2253 , \SUBBYTES[5].a/w2237 , \SUBBYTES[5].a/w2236 ,
         \SUBBYTES[5].a/w2235 , \SUBBYTES[5].a/w2234 , \SUBBYTES[5].a/w2233 ,
         \SUBBYTES[5].a/w2231 , \SUBBYTES[5].a/w2230 , \SUBBYTES[5].a/w2158 ,
         \SUBBYTES[5].a/w2156 , \SUBBYTES[5].a/w2155 , \SUBBYTES[5].a/w2154 ,
         \SUBBYTES[5].a/w2151 , \SUBBYTES[5].a/w2149 , \SUBBYTES[5].a/w2148 ,
         \SUBBYTES[5].a/w2147 , \SUBBYTES[5].a/w2143 , \SUBBYTES[5].a/w2141 ,
         \SUBBYTES[5].a/w2140 , \SUBBYTES[5].a/w2139 , \SUBBYTES[5].a/w2138 ,
         \SUBBYTES[5].a/w2137 , \SUBBYTES[5].a/w2136 , \SUBBYTES[5].a/w2135 ,
         \SUBBYTES[5].a/w2134 , \SUBBYTES[5].a/w2126 , \SUBBYTES[5].a/w2124 ,
         \SUBBYTES[5].a/w2123 , \SUBBYTES[5].a/w2119 , \SUBBYTES[5].a/w2117 ,
         \SUBBYTES[5].a/w2116 , \SUBBYTES[5].a/w2115 , \SUBBYTES[5].a/w2111 ,
         \SUBBYTES[5].a/w2109 , \SUBBYTES[5].a/w2108 , \SUBBYTES[5].a/w2095 ,
         \SUBBYTES[5].a/w2094 , \SUBBYTES[5].a/w2093 , \SUBBYTES[5].a/w2091 ,
         \SUBBYTES[5].a/w2088 , \SUBBYTES[5].a/w2087 , \SUBBYTES[5].a/w2085 ,
         \SUBBYTES[5].a/w2084 , \SUBBYTES[5].a/w2082 , \SUBBYTES[5].a/w2080 ,
         \SUBBYTES[5].a/w2079 , \SUBBYTES[5].a/w2073 , \SUBBYTES[5].a/w2072 ,
         \SUBBYTES[5].a/w2071 , \SUBBYTES[5].a/w2070 , \SUBBYTES[5].a/w2064 ,
         \SUBBYTES[5].a/w2062 , \SUBBYTES[5].a/w2061 , \SUBBYTES[5].a/w2057 ,
         \SUBBYTES[5].a/w2055 , \SUBBYTES[5].a/w2054 , \SUBBYTES[5].a/w2049 ,
         \SUBBYTES[5].a/w2047 , \SUBBYTES[5].a/w2046 , \SUBBYTES[5].a/w2030 ,
         \SUBBYTES[5].a/w2029 , \SUBBYTES[5].a/w2028 , \SUBBYTES[5].a/w2027 ,
         \SUBBYTES[5].a/w2026 , \SUBBYTES[5].a/w2024 , \SUBBYTES[5].a/w2023 ,
         \SUBBYTES[5].a/w1951 , \SUBBYTES[5].a/w1949 , \SUBBYTES[5].a/w1948 ,
         \SUBBYTES[5].a/w1947 , \SUBBYTES[5].a/w1944 , \SUBBYTES[5].a/w1942 ,
         \SUBBYTES[5].a/w1941 , \SUBBYTES[5].a/w1940 , \SUBBYTES[5].a/w1936 ,
         \SUBBYTES[5].a/w1934 , \SUBBYTES[5].a/w1933 , \SUBBYTES[5].a/w1932 ,
         \SUBBYTES[5].a/w1931 , \SUBBYTES[5].a/w1930 , \SUBBYTES[5].a/w1929 ,
         \SUBBYTES[5].a/w1928 , \SUBBYTES[5].a/w1927 , \SUBBYTES[5].a/w1919 ,
         \SUBBYTES[5].a/w1917 , \SUBBYTES[5].a/w1916 , \SUBBYTES[5].a/w1912 ,
         \SUBBYTES[5].a/w1910 , \SUBBYTES[5].a/w1909 , \SUBBYTES[5].a/w1908 ,
         \SUBBYTES[5].a/w1904 , \SUBBYTES[5].a/w1902 , \SUBBYTES[5].a/w1901 ,
         \SUBBYTES[5].a/w1888 , \SUBBYTES[5].a/w1887 , \SUBBYTES[5].a/w1886 ,
         \SUBBYTES[5].a/w1884 , \SUBBYTES[5].a/w1881 , \SUBBYTES[5].a/w1880 ,
         \SUBBYTES[5].a/w1878 , \SUBBYTES[5].a/w1877 , \SUBBYTES[5].a/w1875 ,
         \SUBBYTES[5].a/w1873 , \SUBBYTES[5].a/w1872 , \SUBBYTES[5].a/w1866 ,
         \SUBBYTES[5].a/w1865 , \SUBBYTES[5].a/w1864 , \SUBBYTES[5].a/w1863 ,
         \SUBBYTES[5].a/w1857 , \SUBBYTES[5].a/w1855 , \SUBBYTES[5].a/w1854 ,
         \SUBBYTES[5].a/w1850 , \SUBBYTES[5].a/w1848 , \SUBBYTES[5].a/w1847 ,
         \SUBBYTES[5].a/w1842 , \SUBBYTES[5].a/w1840 , \SUBBYTES[5].a/w1839 ,
         \SUBBYTES[5].a/w1823 , \SUBBYTES[5].a/w1822 , \SUBBYTES[5].a/w1821 ,
         \SUBBYTES[5].a/w1820 , \SUBBYTES[5].a/w1819 , \SUBBYTES[5].a/w1817 ,
         \SUBBYTES[5].a/w1816 , \SUBBYTES[5].a/w1744 , \SUBBYTES[5].a/w1742 ,
         \SUBBYTES[5].a/w1741 , \SUBBYTES[5].a/w1740 , \SUBBYTES[5].a/w1737 ,
         \SUBBYTES[5].a/w1735 , \SUBBYTES[5].a/w1734 , \SUBBYTES[5].a/w1733 ,
         \SUBBYTES[5].a/w1729 , \SUBBYTES[5].a/w1727 , \SUBBYTES[5].a/w1726 ,
         \SUBBYTES[5].a/w1725 , \SUBBYTES[5].a/w1724 , \SUBBYTES[5].a/w1723 ,
         \SUBBYTES[5].a/w1722 , \SUBBYTES[5].a/w1721 , \SUBBYTES[5].a/w1720 ,
         \SUBBYTES[5].a/w1712 , \SUBBYTES[5].a/w1710 , \SUBBYTES[5].a/w1709 ,
         \SUBBYTES[5].a/w1705 , \SUBBYTES[5].a/w1703 , \SUBBYTES[5].a/w1702 ,
         \SUBBYTES[5].a/w1701 , \SUBBYTES[5].a/w1697 , \SUBBYTES[5].a/w1695 ,
         \SUBBYTES[5].a/w1694 , \SUBBYTES[5].a/w1681 , \SUBBYTES[5].a/w1680 ,
         \SUBBYTES[5].a/w1679 , \SUBBYTES[5].a/w1677 , \SUBBYTES[5].a/w1674 ,
         \SUBBYTES[5].a/w1673 , \SUBBYTES[5].a/w1671 , \SUBBYTES[5].a/w1670 ,
         \SUBBYTES[5].a/w1668 , \SUBBYTES[5].a/w1666 , \SUBBYTES[5].a/w1665 ,
         \SUBBYTES[5].a/w1659 , \SUBBYTES[5].a/w1658 , \SUBBYTES[5].a/w1657 ,
         \SUBBYTES[5].a/w1656 , \SUBBYTES[5].a/w1650 , \SUBBYTES[5].a/w1648 ,
         \SUBBYTES[5].a/w1647 , \SUBBYTES[5].a/w1643 , \SUBBYTES[5].a/w1641 ,
         \SUBBYTES[5].a/w1640 , \SUBBYTES[5].a/w1635 , \SUBBYTES[5].a/w1633 ,
         \SUBBYTES[5].a/w1632 , \SUBBYTES[5].a/w1616 , \SUBBYTES[5].a/w1615 ,
         \SUBBYTES[5].a/w1614 , \SUBBYTES[5].a/w1613 , \SUBBYTES[5].a/w1612 ,
         \SUBBYTES[5].a/w1610 , \SUBBYTES[5].a/w1609 , \SUBBYTES[5].a/w1537 ,
         \SUBBYTES[5].a/w1535 , \SUBBYTES[5].a/w1534 , \SUBBYTES[5].a/w1533 ,
         \SUBBYTES[5].a/w1530 , \SUBBYTES[5].a/w1528 , \SUBBYTES[5].a/w1527 ,
         \SUBBYTES[5].a/w1526 , \SUBBYTES[5].a/w1522 , \SUBBYTES[5].a/w1520 ,
         \SUBBYTES[5].a/w1519 , \SUBBYTES[5].a/w1518 , \SUBBYTES[5].a/w1517 ,
         \SUBBYTES[5].a/w1516 , \SUBBYTES[5].a/w1515 , \SUBBYTES[5].a/w1514 ,
         \SUBBYTES[5].a/w1513 , \SUBBYTES[5].a/w1505 , \SUBBYTES[5].a/w1503 ,
         \SUBBYTES[5].a/w1502 , \SUBBYTES[5].a/w1498 , \SUBBYTES[5].a/w1496 ,
         \SUBBYTES[5].a/w1495 , \SUBBYTES[5].a/w1494 , \SUBBYTES[5].a/w1490 ,
         \SUBBYTES[5].a/w1488 , \SUBBYTES[5].a/w1487 , \SUBBYTES[5].a/w1474 ,
         \SUBBYTES[5].a/w1473 , \SUBBYTES[5].a/w1472 , \SUBBYTES[5].a/w1470 ,
         \SUBBYTES[5].a/w1467 , \SUBBYTES[5].a/w1466 , \SUBBYTES[5].a/w1464 ,
         \SUBBYTES[5].a/w1463 , \SUBBYTES[5].a/w1461 , \SUBBYTES[5].a/w1459 ,
         \SUBBYTES[5].a/w1458 , \SUBBYTES[5].a/w1452 , \SUBBYTES[5].a/w1451 ,
         \SUBBYTES[5].a/w1450 , \SUBBYTES[5].a/w1449 , \SUBBYTES[5].a/w1443 ,
         \SUBBYTES[5].a/w1441 , \SUBBYTES[5].a/w1440 , \SUBBYTES[5].a/w1436 ,
         \SUBBYTES[5].a/w1434 , \SUBBYTES[5].a/w1433 , \SUBBYTES[5].a/w1428 ,
         \SUBBYTES[5].a/w1426 , \SUBBYTES[5].a/w1425 , \SUBBYTES[5].a/w1409 ,
         \SUBBYTES[5].a/w1408 , \SUBBYTES[5].a/w1407 , \SUBBYTES[5].a/w1406 ,
         \SUBBYTES[5].a/w1405 , \SUBBYTES[5].a/w1403 , \SUBBYTES[5].a/w1402 ,
         \SUBBYTES[5].a/w1330 , \SUBBYTES[5].a/w1328 , \SUBBYTES[5].a/w1327 ,
         \SUBBYTES[5].a/w1326 , \SUBBYTES[5].a/w1323 , \SUBBYTES[5].a/w1321 ,
         \SUBBYTES[5].a/w1320 , \SUBBYTES[5].a/w1319 , \SUBBYTES[5].a/w1315 ,
         \SUBBYTES[5].a/w1313 , \SUBBYTES[5].a/w1312 , \SUBBYTES[5].a/w1311 ,
         \SUBBYTES[5].a/w1310 , \SUBBYTES[5].a/w1309 , \SUBBYTES[5].a/w1308 ,
         \SUBBYTES[5].a/w1307 , \SUBBYTES[5].a/w1306 , \SUBBYTES[5].a/w1298 ,
         \SUBBYTES[5].a/w1296 , \SUBBYTES[5].a/w1295 , \SUBBYTES[5].a/w1291 ,
         \SUBBYTES[5].a/w1289 , \SUBBYTES[5].a/w1288 , \SUBBYTES[5].a/w1287 ,
         \SUBBYTES[5].a/w1283 , \SUBBYTES[5].a/w1281 , \SUBBYTES[5].a/w1280 ,
         \SUBBYTES[5].a/w1267 , \SUBBYTES[5].a/w1266 , \SUBBYTES[5].a/w1265 ,
         \SUBBYTES[5].a/w1263 , \SUBBYTES[5].a/w1260 , \SUBBYTES[5].a/w1259 ,
         \SUBBYTES[5].a/w1257 , \SUBBYTES[5].a/w1256 , \SUBBYTES[5].a/w1254 ,
         \SUBBYTES[5].a/w1252 , \SUBBYTES[5].a/w1251 , \SUBBYTES[5].a/w1245 ,
         \SUBBYTES[5].a/w1244 , \SUBBYTES[5].a/w1243 , \SUBBYTES[5].a/w1242 ,
         \SUBBYTES[5].a/w1236 , \SUBBYTES[5].a/w1234 , \SUBBYTES[5].a/w1233 ,
         \SUBBYTES[5].a/w1229 , \SUBBYTES[5].a/w1227 , \SUBBYTES[5].a/w1226 ,
         \SUBBYTES[5].a/w1221 , \SUBBYTES[5].a/w1219 , \SUBBYTES[5].a/w1218 ,
         \SUBBYTES[5].a/w1202 , \SUBBYTES[5].a/w1201 , \SUBBYTES[5].a/w1200 ,
         \SUBBYTES[5].a/w1199 , \SUBBYTES[5].a/w1198 , \SUBBYTES[5].a/w1196 ,
         \SUBBYTES[5].a/w1195 , \SUBBYTES[5].a/w1123 , \SUBBYTES[5].a/w1121 ,
         \SUBBYTES[5].a/w1120 , \SUBBYTES[5].a/w1119 , \SUBBYTES[5].a/w1116 ,
         \SUBBYTES[5].a/w1114 , \SUBBYTES[5].a/w1113 , \SUBBYTES[5].a/w1112 ,
         \SUBBYTES[5].a/w1108 , \SUBBYTES[5].a/w1106 , \SUBBYTES[5].a/w1105 ,
         \SUBBYTES[5].a/w1104 , \SUBBYTES[5].a/w1103 , \SUBBYTES[5].a/w1102 ,
         \SUBBYTES[5].a/w1101 , \SUBBYTES[5].a/w1100 , \SUBBYTES[5].a/w1099 ,
         \SUBBYTES[5].a/w1091 , \SUBBYTES[5].a/w1089 , \SUBBYTES[5].a/w1088 ,
         \SUBBYTES[5].a/w1084 , \SUBBYTES[5].a/w1082 , \SUBBYTES[5].a/w1081 ,
         \SUBBYTES[5].a/w1080 , \SUBBYTES[5].a/w1076 , \SUBBYTES[5].a/w1074 ,
         \SUBBYTES[5].a/w1073 , \SUBBYTES[5].a/w1060 , \SUBBYTES[5].a/w1059 ,
         \SUBBYTES[5].a/w1058 , \SUBBYTES[5].a/w1056 , \SUBBYTES[5].a/w1053 ,
         \SUBBYTES[5].a/w1052 , \SUBBYTES[5].a/w1050 , \SUBBYTES[5].a/w1049 ,
         \SUBBYTES[5].a/w1047 , \SUBBYTES[5].a/w1045 , \SUBBYTES[5].a/w1044 ,
         \SUBBYTES[5].a/w1038 , \SUBBYTES[5].a/w1037 , \SUBBYTES[5].a/w1036 ,
         \SUBBYTES[5].a/w1035 , \SUBBYTES[5].a/w1029 , \SUBBYTES[5].a/w1027 ,
         \SUBBYTES[5].a/w1026 , \SUBBYTES[5].a/w1022 , \SUBBYTES[5].a/w1020 ,
         \SUBBYTES[5].a/w1019 , \SUBBYTES[5].a/w1014 , \SUBBYTES[5].a/w1012 ,
         \SUBBYTES[5].a/w1011 , \SUBBYTES[5].a/w995 , \SUBBYTES[5].a/w994 ,
         \SUBBYTES[5].a/w993 , \SUBBYTES[5].a/w992 , \SUBBYTES[5].a/w991 ,
         \SUBBYTES[5].a/w989 , \SUBBYTES[5].a/w988 , \SUBBYTES[5].a/w916 ,
         \SUBBYTES[5].a/w914 , \SUBBYTES[5].a/w913 , \SUBBYTES[5].a/w912 ,
         \SUBBYTES[5].a/w909 , \SUBBYTES[5].a/w907 , \SUBBYTES[5].a/w906 ,
         \SUBBYTES[5].a/w905 , \SUBBYTES[5].a/w901 , \SUBBYTES[5].a/w899 ,
         \SUBBYTES[5].a/w898 , \SUBBYTES[5].a/w897 , \SUBBYTES[5].a/w896 ,
         \SUBBYTES[5].a/w895 , \SUBBYTES[5].a/w894 , \SUBBYTES[5].a/w893 ,
         \SUBBYTES[5].a/w892 , \SUBBYTES[5].a/w884 , \SUBBYTES[5].a/w882 ,
         \SUBBYTES[5].a/w881 , \SUBBYTES[5].a/w877 , \SUBBYTES[5].a/w875 ,
         \SUBBYTES[5].a/w874 , \SUBBYTES[5].a/w873 , \SUBBYTES[5].a/w869 ,
         \SUBBYTES[5].a/w867 , \SUBBYTES[5].a/w866 , \SUBBYTES[5].a/w853 ,
         \SUBBYTES[5].a/w852 , \SUBBYTES[5].a/w851 , \SUBBYTES[5].a/w849 ,
         \SUBBYTES[5].a/w846 , \SUBBYTES[5].a/w845 , \SUBBYTES[5].a/w843 ,
         \SUBBYTES[5].a/w842 , \SUBBYTES[5].a/w840 , \SUBBYTES[5].a/w838 ,
         \SUBBYTES[5].a/w837 , \SUBBYTES[5].a/w831 , \SUBBYTES[5].a/w830 ,
         \SUBBYTES[5].a/w829 , \SUBBYTES[5].a/w828 , \SUBBYTES[5].a/w822 ,
         \SUBBYTES[5].a/w820 , \SUBBYTES[5].a/w819 , \SUBBYTES[5].a/w815 ,
         \SUBBYTES[5].a/w813 , \SUBBYTES[5].a/w812 , \SUBBYTES[5].a/w807 ,
         \SUBBYTES[5].a/w805 , \SUBBYTES[5].a/w804 , \SUBBYTES[5].a/w788 ,
         \SUBBYTES[5].a/w787 , \SUBBYTES[5].a/w786 , \SUBBYTES[5].a/w785 ,
         \SUBBYTES[5].a/w784 , \SUBBYTES[5].a/w782 , \SUBBYTES[5].a/w781 ,
         \SUBBYTES[5].a/w709 , \SUBBYTES[5].a/w707 , \SUBBYTES[5].a/w706 ,
         \SUBBYTES[5].a/w705 , \SUBBYTES[5].a/w702 , \SUBBYTES[5].a/w700 ,
         \SUBBYTES[5].a/w699 , \SUBBYTES[5].a/w698 , \SUBBYTES[5].a/w694 ,
         \SUBBYTES[5].a/w692 , \SUBBYTES[5].a/w691 , \SUBBYTES[5].a/w690 ,
         \SUBBYTES[5].a/w689 , \SUBBYTES[5].a/w688 , \SUBBYTES[5].a/w687 ,
         \SUBBYTES[5].a/w686 , \SUBBYTES[5].a/w685 , \SUBBYTES[5].a/w677 ,
         \SUBBYTES[5].a/w675 , \SUBBYTES[5].a/w674 , \SUBBYTES[5].a/w670 ,
         \SUBBYTES[5].a/w668 , \SUBBYTES[5].a/w667 , \SUBBYTES[5].a/w666 ,
         \SUBBYTES[5].a/w662 , \SUBBYTES[5].a/w660 , \SUBBYTES[5].a/w659 ,
         \SUBBYTES[5].a/w646 , \SUBBYTES[5].a/w645 , \SUBBYTES[5].a/w644 ,
         \SUBBYTES[5].a/w642 , \SUBBYTES[5].a/w639 , \SUBBYTES[5].a/w638 ,
         \SUBBYTES[5].a/w636 , \SUBBYTES[5].a/w635 , \SUBBYTES[5].a/w633 ,
         \SUBBYTES[5].a/w631 , \SUBBYTES[5].a/w630 , \SUBBYTES[5].a/w624 ,
         \SUBBYTES[5].a/w623 , \SUBBYTES[5].a/w622 , \SUBBYTES[5].a/w621 ,
         \SUBBYTES[5].a/w615 , \SUBBYTES[5].a/w613 , \SUBBYTES[5].a/w612 ,
         \SUBBYTES[5].a/w608 , \SUBBYTES[5].a/w606 , \SUBBYTES[5].a/w605 ,
         \SUBBYTES[5].a/w600 , \SUBBYTES[5].a/w598 , \SUBBYTES[5].a/w597 ,
         \SUBBYTES[5].a/w581 , \SUBBYTES[5].a/w580 , \SUBBYTES[5].a/w579 ,
         \SUBBYTES[5].a/w578 , \SUBBYTES[5].a/w577 , \SUBBYTES[5].a/w575 ,
         \SUBBYTES[5].a/w574 , \SUBBYTES[5].a/w502 , \SUBBYTES[5].a/w500 ,
         \SUBBYTES[5].a/w499 , \SUBBYTES[5].a/w498 , \SUBBYTES[5].a/w495 ,
         \SUBBYTES[5].a/w493 , \SUBBYTES[5].a/w492 , \SUBBYTES[5].a/w491 ,
         \SUBBYTES[5].a/w487 , \SUBBYTES[5].a/w485 , \SUBBYTES[5].a/w484 ,
         \SUBBYTES[5].a/w483 , \SUBBYTES[5].a/w482 , \SUBBYTES[5].a/w481 ,
         \SUBBYTES[5].a/w480 , \SUBBYTES[5].a/w479 , \SUBBYTES[5].a/w478 ,
         \SUBBYTES[5].a/w470 , \SUBBYTES[5].a/w468 , \SUBBYTES[5].a/w467 ,
         \SUBBYTES[5].a/w463 , \SUBBYTES[5].a/w461 , \SUBBYTES[5].a/w460 ,
         \SUBBYTES[5].a/w459 , \SUBBYTES[5].a/w455 , \SUBBYTES[5].a/w453 ,
         \SUBBYTES[5].a/w452 , \SUBBYTES[5].a/w439 , \SUBBYTES[5].a/w438 ,
         \SUBBYTES[5].a/w437 , \SUBBYTES[5].a/w435 , \SUBBYTES[5].a/w432 ,
         \SUBBYTES[5].a/w431 , \SUBBYTES[5].a/w429 , \SUBBYTES[5].a/w428 ,
         \SUBBYTES[5].a/w426 , \SUBBYTES[5].a/w424 , \SUBBYTES[5].a/w423 ,
         \SUBBYTES[5].a/w417 , \SUBBYTES[5].a/w416 , \SUBBYTES[5].a/w415 ,
         \SUBBYTES[5].a/w414 , \SUBBYTES[5].a/w408 , \SUBBYTES[5].a/w406 ,
         \SUBBYTES[5].a/w405 , \SUBBYTES[5].a/w401 , \SUBBYTES[5].a/w399 ,
         \SUBBYTES[5].a/w398 , \SUBBYTES[5].a/w393 , \SUBBYTES[5].a/w391 ,
         \SUBBYTES[5].a/w390 , \SUBBYTES[5].a/w374 , \SUBBYTES[5].a/w373 ,
         \SUBBYTES[5].a/w372 , \SUBBYTES[5].a/w371 , \SUBBYTES[5].a/w370 ,
         \SUBBYTES[5].a/w368 , \SUBBYTES[5].a/w367 , \SUBBYTES[5].a/w295 ,
         \SUBBYTES[5].a/w293 , \SUBBYTES[5].a/w292 , \SUBBYTES[5].a/w291 ,
         \SUBBYTES[5].a/w288 , \SUBBYTES[5].a/w286 , \SUBBYTES[5].a/w285 ,
         \SUBBYTES[5].a/w284 , \SUBBYTES[5].a/w280 , \SUBBYTES[5].a/w278 ,
         \SUBBYTES[5].a/w277 , \SUBBYTES[5].a/w276 , \SUBBYTES[5].a/w275 ,
         \SUBBYTES[5].a/w274 , \SUBBYTES[5].a/w273 , \SUBBYTES[5].a/w272 ,
         \SUBBYTES[5].a/w271 , \SUBBYTES[5].a/w263 , \SUBBYTES[5].a/w261 ,
         \SUBBYTES[5].a/w260 , \SUBBYTES[5].a/w256 , \SUBBYTES[5].a/w254 ,
         \SUBBYTES[5].a/w253 , \SUBBYTES[5].a/w252 , \SUBBYTES[5].a/w248 ,
         \SUBBYTES[5].a/w246 , \SUBBYTES[5].a/w245 , \SUBBYTES[5].a/w232 ,
         \SUBBYTES[5].a/w231 , \SUBBYTES[5].a/w230 , \SUBBYTES[5].a/w228 ,
         \SUBBYTES[5].a/w225 , \SUBBYTES[5].a/w224 , \SUBBYTES[5].a/w222 ,
         \SUBBYTES[5].a/w221 , \SUBBYTES[5].a/w219 , \SUBBYTES[5].a/w217 ,
         \SUBBYTES[5].a/w216 , \SUBBYTES[5].a/w210 , \SUBBYTES[5].a/w209 ,
         \SUBBYTES[5].a/w208 , \SUBBYTES[5].a/w207 , \SUBBYTES[5].a/w201 ,
         \SUBBYTES[5].a/w199 , \SUBBYTES[5].a/w198 , \SUBBYTES[5].a/w194 ,
         \SUBBYTES[5].a/w192 , \SUBBYTES[5].a/w191 , \SUBBYTES[5].a/w186 ,
         \SUBBYTES[5].a/w184 , \SUBBYTES[5].a/w183 , \SUBBYTES[5].a/w167 ,
         \SUBBYTES[5].a/w166 , \SUBBYTES[5].a/w165 , \SUBBYTES[5].a/w164 ,
         \SUBBYTES[5].a/w163 , \SUBBYTES[5].a/w161 , \SUBBYTES[5].a/w160 ,
         \SUBBYTES[4].a/w3400 , \SUBBYTES[4].a/w3398 , \SUBBYTES[4].a/w3397 ,
         \SUBBYTES[4].a/w3396 , \SUBBYTES[4].a/w3393 , \SUBBYTES[4].a/w3391 ,
         \SUBBYTES[4].a/w3390 , \SUBBYTES[4].a/w3389 , \SUBBYTES[4].a/w3385 ,
         \SUBBYTES[4].a/w3383 , \SUBBYTES[4].a/w3382 , \SUBBYTES[4].a/w3381 ,
         \SUBBYTES[4].a/w3380 , \SUBBYTES[4].a/w3379 , \SUBBYTES[4].a/w3378 ,
         \SUBBYTES[4].a/w3377 , \SUBBYTES[4].a/w3376 , \SUBBYTES[4].a/w3368 ,
         \SUBBYTES[4].a/w3366 , \SUBBYTES[4].a/w3365 , \SUBBYTES[4].a/w3361 ,
         \SUBBYTES[4].a/w3359 , \SUBBYTES[4].a/w3358 , \SUBBYTES[4].a/w3357 ,
         \SUBBYTES[4].a/w3353 , \SUBBYTES[4].a/w3351 , \SUBBYTES[4].a/w3350 ,
         \SUBBYTES[4].a/w3337 , \SUBBYTES[4].a/w3336 , \SUBBYTES[4].a/w3335 ,
         \SUBBYTES[4].a/w3333 , \SUBBYTES[4].a/w3330 , \SUBBYTES[4].a/w3329 ,
         \SUBBYTES[4].a/w3327 , \SUBBYTES[4].a/w3326 , \SUBBYTES[4].a/w3324 ,
         \SUBBYTES[4].a/w3322 , \SUBBYTES[4].a/w3321 , \SUBBYTES[4].a/w3315 ,
         \SUBBYTES[4].a/w3314 , \SUBBYTES[4].a/w3313 , \SUBBYTES[4].a/w3312 ,
         \SUBBYTES[4].a/w3306 , \SUBBYTES[4].a/w3304 , \SUBBYTES[4].a/w3303 ,
         \SUBBYTES[4].a/w3299 , \SUBBYTES[4].a/w3297 , \SUBBYTES[4].a/w3296 ,
         \SUBBYTES[4].a/w3291 , \SUBBYTES[4].a/w3289 , \SUBBYTES[4].a/w3288 ,
         \SUBBYTES[4].a/w3272 , \SUBBYTES[4].a/w3271 , \SUBBYTES[4].a/w3270 ,
         \SUBBYTES[4].a/w3269 , \SUBBYTES[4].a/w3268 , \SUBBYTES[4].a/w3266 ,
         \SUBBYTES[4].a/w3265 , \SUBBYTES[4].a/w3193 , \SUBBYTES[4].a/w3191 ,
         \SUBBYTES[4].a/w3190 , \SUBBYTES[4].a/w3189 , \SUBBYTES[4].a/w3186 ,
         \SUBBYTES[4].a/w3184 , \SUBBYTES[4].a/w3183 , \SUBBYTES[4].a/w3182 ,
         \SUBBYTES[4].a/w3178 , \SUBBYTES[4].a/w3176 , \SUBBYTES[4].a/w3175 ,
         \SUBBYTES[4].a/w3174 , \SUBBYTES[4].a/w3173 , \SUBBYTES[4].a/w3172 ,
         \SUBBYTES[4].a/w3171 , \SUBBYTES[4].a/w3170 , \SUBBYTES[4].a/w3169 ,
         \SUBBYTES[4].a/w3161 , \SUBBYTES[4].a/w3159 , \SUBBYTES[4].a/w3158 ,
         \SUBBYTES[4].a/w3154 , \SUBBYTES[4].a/w3152 , \SUBBYTES[4].a/w3151 ,
         \SUBBYTES[4].a/w3150 , \SUBBYTES[4].a/w3146 , \SUBBYTES[4].a/w3144 ,
         \SUBBYTES[4].a/w3143 , \SUBBYTES[4].a/w3130 , \SUBBYTES[4].a/w3129 ,
         \SUBBYTES[4].a/w3128 , \SUBBYTES[4].a/w3126 , \SUBBYTES[4].a/w3123 ,
         \SUBBYTES[4].a/w3122 , \SUBBYTES[4].a/w3120 , \SUBBYTES[4].a/w3119 ,
         \SUBBYTES[4].a/w3117 , \SUBBYTES[4].a/w3115 , \SUBBYTES[4].a/w3114 ,
         \SUBBYTES[4].a/w3108 , \SUBBYTES[4].a/w3107 , \SUBBYTES[4].a/w3106 ,
         \SUBBYTES[4].a/w3105 , \SUBBYTES[4].a/w3099 , \SUBBYTES[4].a/w3097 ,
         \SUBBYTES[4].a/w3096 , \SUBBYTES[4].a/w3092 , \SUBBYTES[4].a/w3090 ,
         \SUBBYTES[4].a/w3089 , \SUBBYTES[4].a/w3084 , \SUBBYTES[4].a/w3082 ,
         \SUBBYTES[4].a/w3081 , \SUBBYTES[4].a/w3065 , \SUBBYTES[4].a/w3064 ,
         \SUBBYTES[4].a/w3063 , \SUBBYTES[4].a/w3062 , \SUBBYTES[4].a/w3061 ,
         \SUBBYTES[4].a/w3059 , \SUBBYTES[4].a/w3058 , \SUBBYTES[4].a/w2986 ,
         \SUBBYTES[4].a/w2984 , \SUBBYTES[4].a/w2983 , \SUBBYTES[4].a/w2982 ,
         \SUBBYTES[4].a/w2979 , \SUBBYTES[4].a/w2977 , \SUBBYTES[4].a/w2976 ,
         \SUBBYTES[4].a/w2975 , \SUBBYTES[4].a/w2971 , \SUBBYTES[4].a/w2969 ,
         \SUBBYTES[4].a/w2968 , \SUBBYTES[4].a/w2967 , \SUBBYTES[4].a/w2966 ,
         \SUBBYTES[4].a/w2965 , \SUBBYTES[4].a/w2964 , \SUBBYTES[4].a/w2963 ,
         \SUBBYTES[4].a/w2962 , \SUBBYTES[4].a/w2954 , \SUBBYTES[4].a/w2952 ,
         \SUBBYTES[4].a/w2951 , \SUBBYTES[4].a/w2947 , \SUBBYTES[4].a/w2945 ,
         \SUBBYTES[4].a/w2944 , \SUBBYTES[4].a/w2943 , \SUBBYTES[4].a/w2939 ,
         \SUBBYTES[4].a/w2937 , \SUBBYTES[4].a/w2936 , \SUBBYTES[4].a/w2923 ,
         \SUBBYTES[4].a/w2922 , \SUBBYTES[4].a/w2921 , \SUBBYTES[4].a/w2919 ,
         \SUBBYTES[4].a/w2916 , \SUBBYTES[4].a/w2915 , \SUBBYTES[4].a/w2913 ,
         \SUBBYTES[4].a/w2912 , \SUBBYTES[4].a/w2910 , \SUBBYTES[4].a/w2908 ,
         \SUBBYTES[4].a/w2907 , \SUBBYTES[4].a/w2901 , \SUBBYTES[4].a/w2900 ,
         \SUBBYTES[4].a/w2899 , \SUBBYTES[4].a/w2898 , \SUBBYTES[4].a/w2892 ,
         \SUBBYTES[4].a/w2890 , \SUBBYTES[4].a/w2889 , \SUBBYTES[4].a/w2885 ,
         \SUBBYTES[4].a/w2883 , \SUBBYTES[4].a/w2882 , \SUBBYTES[4].a/w2877 ,
         \SUBBYTES[4].a/w2875 , \SUBBYTES[4].a/w2874 , \SUBBYTES[4].a/w2858 ,
         \SUBBYTES[4].a/w2857 , \SUBBYTES[4].a/w2856 , \SUBBYTES[4].a/w2855 ,
         \SUBBYTES[4].a/w2854 , \SUBBYTES[4].a/w2852 , \SUBBYTES[4].a/w2851 ,
         \SUBBYTES[4].a/w2779 , \SUBBYTES[4].a/w2777 , \SUBBYTES[4].a/w2776 ,
         \SUBBYTES[4].a/w2775 , \SUBBYTES[4].a/w2772 , \SUBBYTES[4].a/w2770 ,
         \SUBBYTES[4].a/w2769 , \SUBBYTES[4].a/w2768 , \SUBBYTES[4].a/w2764 ,
         \SUBBYTES[4].a/w2762 , \SUBBYTES[4].a/w2761 , \SUBBYTES[4].a/w2760 ,
         \SUBBYTES[4].a/w2759 , \SUBBYTES[4].a/w2758 , \SUBBYTES[4].a/w2757 ,
         \SUBBYTES[4].a/w2756 , \SUBBYTES[4].a/w2755 , \SUBBYTES[4].a/w2747 ,
         \SUBBYTES[4].a/w2745 , \SUBBYTES[4].a/w2744 , \SUBBYTES[4].a/w2740 ,
         \SUBBYTES[4].a/w2738 , \SUBBYTES[4].a/w2737 , \SUBBYTES[4].a/w2736 ,
         \SUBBYTES[4].a/w2732 , \SUBBYTES[4].a/w2730 , \SUBBYTES[4].a/w2729 ,
         \SUBBYTES[4].a/w2716 , \SUBBYTES[4].a/w2715 , \SUBBYTES[4].a/w2714 ,
         \SUBBYTES[4].a/w2712 , \SUBBYTES[4].a/w2709 , \SUBBYTES[4].a/w2708 ,
         \SUBBYTES[4].a/w2706 , \SUBBYTES[4].a/w2705 , \SUBBYTES[4].a/w2703 ,
         \SUBBYTES[4].a/w2701 , \SUBBYTES[4].a/w2700 , \SUBBYTES[4].a/w2694 ,
         \SUBBYTES[4].a/w2693 , \SUBBYTES[4].a/w2692 , \SUBBYTES[4].a/w2691 ,
         \SUBBYTES[4].a/w2685 , \SUBBYTES[4].a/w2683 , \SUBBYTES[4].a/w2682 ,
         \SUBBYTES[4].a/w2678 , \SUBBYTES[4].a/w2676 , \SUBBYTES[4].a/w2675 ,
         \SUBBYTES[4].a/w2670 , \SUBBYTES[4].a/w2668 , \SUBBYTES[4].a/w2667 ,
         \SUBBYTES[4].a/w2651 , \SUBBYTES[4].a/w2650 , \SUBBYTES[4].a/w2649 ,
         \SUBBYTES[4].a/w2648 , \SUBBYTES[4].a/w2647 , \SUBBYTES[4].a/w2645 ,
         \SUBBYTES[4].a/w2644 , \SUBBYTES[4].a/w2572 , \SUBBYTES[4].a/w2570 ,
         \SUBBYTES[4].a/w2569 , \SUBBYTES[4].a/w2568 , \SUBBYTES[4].a/w2565 ,
         \SUBBYTES[4].a/w2563 , \SUBBYTES[4].a/w2562 , \SUBBYTES[4].a/w2561 ,
         \SUBBYTES[4].a/w2557 , \SUBBYTES[4].a/w2555 , \SUBBYTES[4].a/w2554 ,
         \SUBBYTES[4].a/w2553 , \SUBBYTES[4].a/w2552 , \SUBBYTES[4].a/w2551 ,
         \SUBBYTES[4].a/w2550 , \SUBBYTES[4].a/w2549 , \SUBBYTES[4].a/w2548 ,
         \SUBBYTES[4].a/w2540 , \SUBBYTES[4].a/w2538 , \SUBBYTES[4].a/w2537 ,
         \SUBBYTES[4].a/w2533 , \SUBBYTES[4].a/w2531 , \SUBBYTES[4].a/w2530 ,
         \SUBBYTES[4].a/w2529 , \SUBBYTES[4].a/w2525 , \SUBBYTES[4].a/w2523 ,
         \SUBBYTES[4].a/w2522 , \SUBBYTES[4].a/w2509 , \SUBBYTES[4].a/w2508 ,
         \SUBBYTES[4].a/w2507 , \SUBBYTES[4].a/w2505 , \SUBBYTES[4].a/w2502 ,
         \SUBBYTES[4].a/w2501 , \SUBBYTES[4].a/w2499 , \SUBBYTES[4].a/w2498 ,
         \SUBBYTES[4].a/w2496 , \SUBBYTES[4].a/w2494 , \SUBBYTES[4].a/w2493 ,
         \SUBBYTES[4].a/w2487 , \SUBBYTES[4].a/w2486 , \SUBBYTES[4].a/w2485 ,
         \SUBBYTES[4].a/w2484 , \SUBBYTES[4].a/w2478 , \SUBBYTES[4].a/w2476 ,
         \SUBBYTES[4].a/w2475 , \SUBBYTES[4].a/w2471 , \SUBBYTES[4].a/w2469 ,
         \SUBBYTES[4].a/w2468 , \SUBBYTES[4].a/w2463 , \SUBBYTES[4].a/w2461 ,
         \SUBBYTES[4].a/w2460 , \SUBBYTES[4].a/w2444 , \SUBBYTES[4].a/w2443 ,
         \SUBBYTES[4].a/w2442 , \SUBBYTES[4].a/w2441 , \SUBBYTES[4].a/w2440 ,
         \SUBBYTES[4].a/w2438 , \SUBBYTES[4].a/w2437 , \SUBBYTES[4].a/w2365 ,
         \SUBBYTES[4].a/w2363 , \SUBBYTES[4].a/w2362 , \SUBBYTES[4].a/w2361 ,
         \SUBBYTES[4].a/w2358 , \SUBBYTES[4].a/w2356 , \SUBBYTES[4].a/w2355 ,
         \SUBBYTES[4].a/w2354 , \SUBBYTES[4].a/w2350 , \SUBBYTES[4].a/w2348 ,
         \SUBBYTES[4].a/w2347 , \SUBBYTES[4].a/w2346 , \SUBBYTES[4].a/w2345 ,
         \SUBBYTES[4].a/w2344 , \SUBBYTES[4].a/w2343 , \SUBBYTES[4].a/w2342 ,
         \SUBBYTES[4].a/w2341 , \SUBBYTES[4].a/w2333 , \SUBBYTES[4].a/w2331 ,
         \SUBBYTES[4].a/w2330 , \SUBBYTES[4].a/w2326 , \SUBBYTES[4].a/w2324 ,
         \SUBBYTES[4].a/w2323 , \SUBBYTES[4].a/w2322 , \SUBBYTES[4].a/w2318 ,
         \SUBBYTES[4].a/w2316 , \SUBBYTES[4].a/w2315 , \SUBBYTES[4].a/w2302 ,
         \SUBBYTES[4].a/w2301 , \SUBBYTES[4].a/w2300 , \SUBBYTES[4].a/w2298 ,
         \SUBBYTES[4].a/w2295 , \SUBBYTES[4].a/w2294 , \SUBBYTES[4].a/w2292 ,
         \SUBBYTES[4].a/w2291 , \SUBBYTES[4].a/w2289 , \SUBBYTES[4].a/w2287 ,
         \SUBBYTES[4].a/w2286 , \SUBBYTES[4].a/w2280 , \SUBBYTES[4].a/w2279 ,
         \SUBBYTES[4].a/w2278 , \SUBBYTES[4].a/w2277 , \SUBBYTES[4].a/w2271 ,
         \SUBBYTES[4].a/w2269 , \SUBBYTES[4].a/w2268 , \SUBBYTES[4].a/w2264 ,
         \SUBBYTES[4].a/w2262 , \SUBBYTES[4].a/w2261 , \SUBBYTES[4].a/w2256 ,
         \SUBBYTES[4].a/w2254 , \SUBBYTES[4].a/w2253 , \SUBBYTES[4].a/w2237 ,
         \SUBBYTES[4].a/w2236 , \SUBBYTES[4].a/w2235 , \SUBBYTES[4].a/w2234 ,
         \SUBBYTES[4].a/w2233 , \SUBBYTES[4].a/w2231 , \SUBBYTES[4].a/w2230 ,
         \SUBBYTES[4].a/w2158 , \SUBBYTES[4].a/w2156 , \SUBBYTES[4].a/w2155 ,
         \SUBBYTES[4].a/w2154 , \SUBBYTES[4].a/w2151 , \SUBBYTES[4].a/w2149 ,
         \SUBBYTES[4].a/w2148 , \SUBBYTES[4].a/w2147 , \SUBBYTES[4].a/w2143 ,
         \SUBBYTES[4].a/w2141 , \SUBBYTES[4].a/w2140 , \SUBBYTES[4].a/w2139 ,
         \SUBBYTES[4].a/w2138 , \SUBBYTES[4].a/w2137 , \SUBBYTES[4].a/w2136 ,
         \SUBBYTES[4].a/w2135 , \SUBBYTES[4].a/w2134 , \SUBBYTES[4].a/w2126 ,
         \SUBBYTES[4].a/w2124 , \SUBBYTES[4].a/w2123 , \SUBBYTES[4].a/w2119 ,
         \SUBBYTES[4].a/w2117 , \SUBBYTES[4].a/w2116 , \SUBBYTES[4].a/w2115 ,
         \SUBBYTES[4].a/w2111 , \SUBBYTES[4].a/w2109 , \SUBBYTES[4].a/w2108 ,
         \SUBBYTES[4].a/w2095 , \SUBBYTES[4].a/w2094 , \SUBBYTES[4].a/w2093 ,
         \SUBBYTES[4].a/w2091 , \SUBBYTES[4].a/w2088 , \SUBBYTES[4].a/w2087 ,
         \SUBBYTES[4].a/w2085 , \SUBBYTES[4].a/w2084 , \SUBBYTES[4].a/w2082 ,
         \SUBBYTES[4].a/w2080 , \SUBBYTES[4].a/w2079 , \SUBBYTES[4].a/w2073 ,
         \SUBBYTES[4].a/w2072 , \SUBBYTES[4].a/w2071 , \SUBBYTES[4].a/w2070 ,
         \SUBBYTES[4].a/w2064 , \SUBBYTES[4].a/w2062 , \SUBBYTES[4].a/w2061 ,
         \SUBBYTES[4].a/w2057 , \SUBBYTES[4].a/w2055 , \SUBBYTES[4].a/w2054 ,
         \SUBBYTES[4].a/w2049 , \SUBBYTES[4].a/w2047 , \SUBBYTES[4].a/w2046 ,
         \SUBBYTES[4].a/w2030 , \SUBBYTES[4].a/w2029 , \SUBBYTES[4].a/w2028 ,
         \SUBBYTES[4].a/w2027 , \SUBBYTES[4].a/w2026 , \SUBBYTES[4].a/w2024 ,
         \SUBBYTES[4].a/w2023 , \SUBBYTES[4].a/w1951 , \SUBBYTES[4].a/w1949 ,
         \SUBBYTES[4].a/w1948 , \SUBBYTES[4].a/w1947 , \SUBBYTES[4].a/w1944 ,
         \SUBBYTES[4].a/w1942 , \SUBBYTES[4].a/w1941 , \SUBBYTES[4].a/w1940 ,
         \SUBBYTES[4].a/w1936 , \SUBBYTES[4].a/w1934 , \SUBBYTES[4].a/w1933 ,
         \SUBBYTES[4].a/w1932 , \SUBBYTES[4].a/w1931 , \SUBBYTES[4].a/w1930 ,
         \SUBBYTES[4].a/w1929 , \SUBBYTES[4].a/w1928 , \SUBBYTES[4].a/w1927 ,
         \SUBBYTES[4].a/w1919 , \SUBBYTES[4].a/w1917 , \SUBBYTES[4].a/w1916 ,
         \SUBBYTES[4].a/w1912 , \SUBBYTES[4].a/w1910 , \SUBBYTES[4].a/w1909 ,
         \SUBBYTES[4].a/w1908 , \SUBBYTES[4].a/w1904 , \SUBBYTES[4].a/w1902 ,
         \SUBBYTES[4].a/w1901 , \SUBBYTES[4].a/w1888 , \SUBBYTES[4].a/w1887 ,
         \SUBBYTES[4].a/w1886 , \SUBBYTES[4].a/w1884 , \SUBBYTES[4].a/w1881 ,
         \SUBBYTES[4].a/w1880 , \SUBBYTES[4].a/w1878 , \SUBBYTES[4].a/w1877 ,
         \SUBBYTES[4].a/w1875 , \SUBBYTES[4].a/w1873 , \SUBBYTES[4].a/w1872 ,
         \SUBBYTES[4].a/w1866 , \SUBBYTES[4].a/w1865 , \SUBBYTES[4].a/w1864 ,
         \SUBBYTES[4].a/w1863 , \SUBBYTES[4].a/w1857 , \SUBBYTES[4].a/w1855 ,
         \SUBBYTES[4].a/w1854 , \SUBBYTES[4].a/w1850 , \SUBBYTES[4].a/w1848 ,
         \SUBBYTES[4].a/w1847 , \SUBBYTES[4].a/w1842 , \SUBBYTES[4].a/w1840 ,
         \SUBBYTES[4].a/w1839 , \SUBBYTES[4].a/w1823 , \SUBBYTES[4].a/w1822 ,
         \SUBBYTES[4].a/w1821 , \SUBBYTES[4].a/w1820 , \SUBBYTES[4].a/w1819 ,
         \SUBBYTES[4].a/w1817 , \SUBBYTES[4].a/w1816 , \SUBBYTES[4].a/w1744 ,
         \SUBBYTES[4].a/w1742 , \SUBBYTES[4].a/w1741 , \SUBBYTES[4].a/w1740 ,
         \SUBBYTES[4].a/w1737 , \SUBBYTES[4].a/w1735 , \SUBBYTES[4].a/w1734 ,
         \SUBBYTES[4].a/w1733 , \SUBBYTES[4].a/w1729 , \SUBBYTES[4].a/w1727 ,
         \SUBBYTES[4].a/w1726 , \SUBBYTES[4].a/w1725 , \SUBBYTES[4].a/w1724 ,
         \SUBBYTES[4].a/w1723 , \SUBBYTES[4].a/w1722 , \SUBBYTES[4].a/w1721 ,
         \SUBBYTES[4].a/w1720 , \SUBBYTES[4].a/w1712 , \SUBBYTES[4].a/w1710 ,
         \SUBBYTES[4].a/w1709 , \SUBBYTES[4].a/w1705 , \SUBBYTES[4].a/w1703 ,
         \SUBBYTES[4].a/w1702 , \SUBBYTES[4].a/w1701 , \SUBBYTES[4].a/w1697 ,
         \SUBBYTES[4].a/w1695 , \SUBBYTES[4].a/w1694 , \SUBBYTES[4].a/w1681 ,
         \SUBBYTES[4].a/w1680 , \SUBBYTES[4].a/w1679 , \SUBBYTES[4].a/w1677 ,
         \SUBBYTES[4].a/w1674 , \SUBBYTES[4].a/w1673 , \SUBBYTES[4].a/w1671 ,
         \SUBBYTES[4].a/w1670 , \SUBBYTES[4].a/w1668 , \SUBBYTES[4].a/w1666 ,
         \SUBBYTES[4].a/w1665 , \SUBBYTES[4].a/w1659 , \SUBBYTES[4].a/w1658 ,
         \SUBBYTES[4].a/w1657 , \SUBBYTES[4].a/w1656 , \SUBBYTES[4].a/w1650 ,
         \SUBBYTES[4].a/w1648 , \SUBBYTES[4].a/w1647 , \SUBBYTES[4].a/w1643 ,
         \SUBBYTES[4].a/w1641 , \SUBBYTES[4].a/w1640 , \SUBBYTES[4].a/w1635 ,
         \SUBBYTES[4].a/w1633 , \SUBBYTES[4].a/w1632 , \SUBBYTES[4].a/w1616 ,
         \SUBBYTES[4].a/w1615 , \SUBBYTES[4].a/w1614 , \SUBBYTES[4].a/w1613 ,
         \SUBBYTES[4].a/w1612 , \SUBBYTES[4].a/w1610 , \SUBBYTES[4].a/w1609 ,
         \SUBBYTES[4].a/w1537 , \SUBBYTES[4].a/w1535 , \SUBBYTES[4].a/w1534 ,
         \SUBBYTES[4].a/w1533 , \SUBBYTES[4].a/w1530 , \SUBBYTES[4].a/w1528 ,
         \SUBBYTES[4].a/w1527 , \SUBBYTES[4].a/w1526 , \SUBBYTES[4].a/w1522 ,
         \SUBBYTES[4].a/w1520 , \SUBBYTES[4].a/w1519 , \SUBBYTES[4].a/w1518 ,
         \SUBBYTES[4].a/w1517 , \SUBBYTES[4].a/w1516 , \SUBBYTES[4].a/w1515 ,
         \SUBBYTES[4].a/w1514 , \SUBBYTES[4].a/w1513 , \SUBBYTES[4].a/w1505 ,
         \SUBBYTES[4].a/w1503 , \SUBBYTES[4].a/w1502 , \SUBBYTES[4].a/w1498 ,
         \SUBBYTES[4].a/w1496 , \SUBBYTES[4].a/w1495 , \SUBBYTES[4].a/w1494 ,
         \SUBBYTES[4].a/w1490 , \SUBBYTES[4].a/w1488 , \SUBBYTES[4].a/w1487 ,
         \SUBBYTES[4].a/w1474 , \SUBBYTES[4].a/w1473 , \SUBBYTES[4].a/w1472 ,
         \SUBBYTES[4].a/w1470 , \SUBBYTES[4].a/w1467 , \SUBBYTES[4].a/w1466 ,
         \SUBBYTES[4].a/w1464 , \SUBBYTES[4].a/w1463 , \SUBBYTES[4].a/w1461 ,
         \SUBBYTES[4].a/w1459 , \SUBBYTES[4].a/w1458 , \SUBBYTES[4].a/w1452 ,
         \SUBBYTES[4].a/w1451 , \SUBBYTES[4].a/w1450 , \SUBBYTES[4].a/w1449 ,
         \SUBBYTES[4].a/w1443 , \SUBBYTES[4].a/w1441 , \SUBBYTES[4].a/w1440 ,
         \SUBBYTES[4].a/w1436 , \SUBBYTES[4].a/w1434 , \SUBBYTES[4].a/w1433 ,
         \SUBBYTES[4].a/w1428 , \SUBBYTES[4].a/w1426 , \SUBBYTES[4].a/w1425 ,
         \SUBBYTES[4].a/w1409 , \SUBBYTES[4].a/w1408 , \SUBBYTES[4].a/w1407 ,
         \SUBBYTES[4].a/w1406 , \SUBBYTES[4].a/w1405 , \SUBBYTES[4].a/w1403 ,
         \SUBBYTES[4].a/w1402 , \SUBBYTES[4].a/w1330 , \SUBBYTES[4].a/w1328 ,
         \SUBBYTES[4].a/w1327 , \SUBBYTES[4].a/w1326 , \SUBBYTES[4].a/w1323 ,
         \SUBBYTES[4].a/w1321 , \SUBBYTES[4].a/w1320 , \SUBBYTES[4].a/w1319 ,
         \SUBBYTES[4].a/w1315 , \SUBBYTES[4].a/w1313 , \SUBBYTES[4].a/w1312 ,
         \SUBBYTES[4].a/w1311 , \SUBBYTES[4].a/w1310 , \SUBBYTES[4].a/w1309 ,
         \SUBBYTES[4].a/w1308 , \SUBBYTES[4].a/w1307 , \SUBBYTES[4].a/w1306 ,
         \SUBBYTES[4].a/w1298 , \SUBBYTES[4].a/w1296 , \SUBBYTES[4].a/w1295 ,
         \SUBBYTES[4].a/w1291 , \SUBBYTES[4].a/w1289 , \SUBBYTES[4].a/w1288 ,
         \SUBBYTES[4].a/w1287 , \SUBBYTES[4].a/w1283 , \SUBBYTES[4].a/w1281 ,
         \SUBBYTES[4].a/w1280 , \SUBBYTES[4].a/w1267 , \SUBBYTES[4].a/w1266 ,
         \SUBBYTES[4].a/w1265 , \SUBBYTES[4].a/w1263 , \SUBBYTES[4].a/w1260 ,
         \SUBBYTES[4].a/w1259 , \SUBBYTES[4].a/w1257 , \SUBBYTES[4].a/w1256 ,
         \SUBBYTES[4].a/w1254 , \SUBBYTES[4].a/w1252 , \SUBBYTES[4].a/w1251 ,
         \SUBBYTES[4].a/w1245 , \SUBBYTES[4].a/w1244 , \SUBBYTES[4].a/w1243 ,
         \SUBBYTES[4].a/w1242 , \SUBBYTES[4].a/w1236 , \SUBBYTES[4].a/w1234 ,
         \SUBBYTES[4].a/w1233 , \SUBBYTES[4].a/w1229 , \SUBBYTES[4].a/w1227 ,
         \SUBBYTES[4].a/w1226 , \SUBBYTES[4].a/w1221 , \SUBBYTES[4].a/w1219 ,
         \SUBBYTES[4].a/w1218 , \SUBBYTES[4].a/w1202 , \SUBBYTES[4].a/w1201 ,
         \SUBBYTES[4].a/w1200 , \SUBBYTES[4].a/w1199 , \SUBBYTES[4].a/w1198 ,
         \SUBBYTES[4].a/w1196 , \SUBBYTES[4].a/w1195 , \SUBBYTES[4].a/w1123 ,
         \SUBBYTES[4].a/w1121 , \SUBBYTES[4].a/w1120 , \SUBBYTES[4].a/w1119 ,
         \SUBBYTES[4].a/w1116 , \SUBBYTES[4].a/w1114 , \SUBBYTES[4].a/w1113 ,
         \SUBBYTES[4].a/w1112 , \SUBBYTES[4].a/w1108 , \SUBBYTES[4].a/w1106 ,
         \SUBBYTES[4].a/w1105 , \SUBBYTES[4].a/w1104 , \SUBBYTES[4].a/w1103 ,
         \SUBBYTES[4].a/w1102 , \SUBBYTES[4].a/w1101 , \SUBBYTES[4].a/w1100 ,
         \SUBBYTES[4].a/w1099 , \SUBBYTES[4].a/w1091 , \SUBBYTES[4].a/w1089 ,
         \SUBBYTES[4].a/w1088 , \SUBBYTES[4].a/w1084 , \SUBBYTES[4].a/w1082 ,
         \SUBBYTES[4].a/w1081 , \SUBBYTES[4].a/w1080 , \SUBBYTES[4].a/w1076 ,
         \SUBBYTES[4].a/w1074 , \SUBBYTES[4].a/w1073 , \SUBBYTES[4].a/w1060 ,
         \SUBBYTES[4].a/w1059 , \SUBBYTES[4].a/w1058 , \SUBBYTES[4].a/w1056 ,
         \SUBBYTES[4].a/w1053 , \SUBBYTES[4].a/w1052 , \SUBBYTES[4].a/w1050 ,
         \SUBBYTES[4].a/w1049 , \SUBBYTES[4].a/w1047 , \SUBBYTES[4].a/w1045 ,
         \SUBBYTES[4].a/w1044 , \SUBBYTES[4].a/w1038 , \SUBBYTES[4].a/w1037 ,
         \SUBBYTES[4].a/w1036 , \SUBBYTES[4].a/w1035 , \SUBBYTES[4].a/w1029 ,
         \SUBBYTES[4].a/w1027 , \SUBBYTES[4].a/w1026 , \SUBBYTES[4].a/w1022 ,
         \SUBBYTES[4].a/w1020 , \SUBBYTES[4].a/w1019 , \SUBBYTES[4].a/w1014 ,
         \SUBBYTES[4].a/w1012 , \SUBBYTES[4].a/w1011 , \SUBBYTES[4].a/w995 ,
         \SUBBYTES[4].a/w994 , \SUBBYTES[4].a/w993 , \SUBBYTES[4].a/w992 ,
         \SUBBYTES[4].a/w991 , \SUBBYTES[4].a/w989 , \SUBBYTES[4].a/w988 ,
         \SUBBYTES[4].a/w916 , \SUBBYTES[4].a/w914 , \SUBBYTES[4].a/w913 ,
         \SUBBYTES[4].a/w912 , \SUBBYTES[4].a/w909 , \SUBBYTES[4].a/w907 ,
         \SUBBYTES[4].a/w906 , \SUBBYTES[4].a/w905 , \SUBBYTES[4].a/w901 ,
         \SUBBYTES[4].a/w899 , \SUBBYTES[4].a/w898 , \SUBBYTES[4].a/w897 ,
         \SUBBYTES[4].a/w896 , \SUBBYTES[4].a/w895 , \SUBBYTES[4].a/w894 ,
         \SUBBYTES[4].a/w893 , \SUBBYTES[4].a/w892 , \SUBBYTES[4].a/w884 ,
         \SUBBYTES[4].a/w882 , \SUBBYTES[4].a/w881 , \SUBBYTES[4].a/w877 ,
         \SUBBYTES[4].a/w875 , \SUBBYTES[4].a/w874 , \SUBBYTES[4].a/w873 ,
         \SUBBYTES[4].a/w869 , \SUBBYTES[4].a/w867 , \SUBBYTES[4].a/w866 ,
         \SUBBYTES[4].a/w853 , \SUBBYTES[4].a/w852 , \SUBBYTES[4].a/w851 ,
         \SUBBYTES[4].a/w849 , \SUBBYTES[4].a/w846 , \SUBBYTES[4].a/w845 ,
         \SUBBYTES[4].a/w843 , \SUBBYTES[4].a/w842 , \SUBBYTES[4].a/w840 ,
         \SUBBYTES[4].a/w838 , \SUBBYTES[4].a/w837 , \SUBBYTES[4].a/w831 ,
         \SUBBYTES[4].a/w830 , \SUBBYTES[4].a/w829 , \SUBBYTES[4].a/w828 ,
         \SUBBYTES[4].a/w822 , \SUBBYTES[4].a/w820 , \SUBBYTES[4].a/w819 ,
         \SUBBYTES[4].a/w815 , \SUBBYTES[4].a/w813 , \SUBBYTES[4].a/w812 ,
         \SUBBYTES[4].a/w807 , \SUBBYTES[4].a/w805 , \SUBBYTES[4].a/w804 ,
         \SUBBYTES[4].a/w788 , \SUBBYTES[4].a/w787 , \SUBBYTES[4].a/w786 ,
         \SUBBYTES[4].a/w785 , \SUBBYTES[4].a/w784 , \SUBBYTES[4].a/w782 ,
         \SUBBYTES[4].a/w781 , \SUBBYTES[4].a/w709 , \SUBBYTES[4].a/w707 ,
         \SUBBYTES[4].a/w706 , \SUBBYTES[4].a/w705 , \SUBBYTES[4].a/w702 ,
         \SUBBYTES[4].a/w700 , \SUBBYTES[4].a/w699 , \SUBBYTES[4].a/w698 ,
         \SUBBYTES[4].a/w694 , \SUBBYTES[4].a/w692 , \SUBBYTES[4].a/w691 ,
         \SUBBYTES[4].a/w690 , \SUBBYTES[4].a/w689 , \SUBBYTES[4].a/w688 ,
         \SUBBYTES[4].a/w687 , \SUBBYTES[4].a/w686 , \SUBBYTES[4].a/w685 ,
         \SUBBYTES[4].a/w677 , \SUBBYTES[4].a/w675 , \SUBBYTES[4].a/w674 ,
         \SUBBYTES[4].a/w670 , \SUBBYTES[4].a/w668 , \SUBBYTES[4].a/w667 ,
         \SUBBYTES[4].a/w666 , \SUBBYTES[4].a/w662 , \SUBBYTES[4].a/w660 ,
         \SUBBYTES[4].a/w659 , \SUBBYTES[4].a/w646 , \SUBBYTES[4].a/w645 ,
         \SUBBYTES[4].a/w644 , \SUBBYTES[4].a/w642 , \SUBBYTES[4].a/w639 ,
         \SUBBYTES[4].a/w638 , \SUBBYTES[4].a/w636 , \SUBBYTES[4].a/w635 ,
         \SUBBYTES[4].a/w633 , \SUBBYTES[4].a/w631 , \SUBBYTES[4].a/w630 ,
         \SUBBYTES[4].a/w624 , \SUBBYTES[4].a/w623 , \SUBBYTES[4].a/w622 ,
         \SUBBYTES[4].a/w621 , \SUBBYTES[4].a/w615 , \SUBBYTES[4].a/w613 ,
         \SUBBYTES[4].a/w612 , \SUBBYTES[4].a/w608 , \SUBBYTES[4].a/w606 ,
         \SUBBYTES[4].a/w605 , \SUBBYTES[4].a/w600 , \SUBBYTES[4].a/w598 ,
         \SUBBYTES[4].a/w597 , \SUBBYTES[4].a/w581 , \SUBBYTES[4].a/w580 ,
         \SUBBYTES[4].a/w579 , \SUBBYTES[4].a/w578 , \SUBBYTES[4].a/w577 ,
         \SUBBYTES[4].a/w575 , \SUBBYTES[4].a/w574 , \SUBBYTES[4].a/w502 ,
         \SUBBYTES[4].a/w500 , \SUBBYTES[4].a/w499 , \SUBBYTES[4].a/w498 ,
         \SUBBYTES[4].a/w495 , \SUBBYTES[4].a/w493 , \SUBBYTES[4].a/w492 ,
         \SUBBYTES[4].a/w491 , \SUBBYTES[4].a/w487 , \SUBBYTES[4].a/w485 ,
         \SUBBYTES[4].a/w484 , \SUBBYTES[4].a/w483 , \SUBBYTES[4].a/w482 ,
         \SUBBYTES[4].a/w481 , \SUBBYTES[4].a/w480 , \SUBBYTES[4].a/w479 ,
         \SUBBYTES[4].a/w478 , \SUBBYTES[4].a/w470 , \SUBBYTES[4].a/w468 ,
         \SUBBYTES[4].a/w467 , \SUBBYTES[4].a/w463 , \SUBBYTES[4].a/w461 ,
         \SUBBYTES[4].a/w460 , \SUBBYTES[4].a/w459 , \SUBBYTES[4].a/w455 ,
         \SUBBYTES[4].a/w453 , \SUBBYTES[4].a/w452 , \SUBBYTES[4].a/w439 ,
         \SUBBYTES[4].a/w438 , \SUBBYTES[4].a/w437 , \SUBBYTES[4].a/w435 ,
         \SUBBYTES[4].a/w432 , \SUBBYTES[4].a/w431 , \SUBBYTES[4].a/w429 ,
         \SUBBYTES[4].a/w428 , \SUBBYTES[4].a/w426 , \SUBBYTES[4].a/w424 ,
         \SUBBYTES[4].a/w423 , \SUBBYTES[4].a/w417 , \SUBBYTES[4].a/w416 ,
         \SUBBYTES[4].a/w415 , \SUBBYTES[4].a/w414 , \SUBBYTES[4].a/w408 ,
         \SUBBYTES[4].a/w406 , \SUBBYTES[4].a/w405 , \SUBBYTES[4].a/w401 ,
         \SUBBYTES[4].a/w399 , \SUBBYTES[4].a/w398 , \SUBBYTES[4].a/w393 ,
         \SUBBYTES[4].a/w391 , \SUBBYTES[4].a/w390 , \SUBBYTES[4].a/w374 ,
         \SUBBYTES[4].a/w373 , \SUBBYTES[4].a/w372 , \SUBBYTES[4].a/w371 ,
         \SUBBYTES[4].a/w370 , \SUBBYTES[4].a/w368 , \SUBBYTES[4].a/w367 ,
         \SUBBYTES[4].a/w295 , \SUBBYTES[4].a/w293 , \SUBBYTES[4].a/w292 ,
         \SUBBYTES[4].a/w291 , \SUBBYTES[4].a/w288 , \SUBBYTES[4].a/w286 ,
         \SUBBYTES[4].a/w285 , \SUBBYTES[4].a/w284 , \SUBBYTES[4].a/w280 ,
         \SUBBYTES[4].a/w278 , \SUBBYTES[4].a/w277 , \SUBBYTES[4].a/w276 ,
         \SUBBYTES[4].a/w275 , \SUBBYTES[4].a/w274 , \SUBBYTES[4].a/w273 ,
         \SUBBYTES[4].a/w272 , \SUBBYTES[4].a/w271 , \SUBBYTES[4].a/w263 ,
         \SUBBYTES[4].a/w261 , \SUBBYTES[4].a/w260 , \SUBBYTES[4].a/w256 ,
         \SUBBYTES[4].a/w254 , \SUBBYTES[4].a/w253 , \SUBBYTES[4].a/w252 ,
         \SUBBYTES[4].a/w248 , \SUBBYTES[4].a/w246 , \SUBBYTES[4].a/w245 ,
         \SUBBYTES[4].a/w232 , \SUBBYTES[4].a/w231 , \SUBBYTES[4].a/w230 ,
         \SUBBYTES[4].a/w228 , \SUBBYTES[4].a/w225 , \SUBBYTES[4].a/w224 ,
         \SUBBYTES[4].a/w222 , \SUBBYTES[4].a/w221 , \SUBBYTES[4].a/w219 ,
         \SUBBYTES[4].a/w217 , \SUBBYTES[4].a/w216 , \SUBBYTES[4].a/w210 ,
         \SUBBYTES[4].a/w209 , \SUBBYTES[4].a/w208 , \SUBBYTES[4].a/w207 ,
         \SUBBYTES[4].a/w201 , \SUBBYTES[4].a/w199 , \SUBBYTES[4].a/w198 ,
         \SUBBYTES[4].a/w194 , \SUBBYTES[4].a/w192 , \SUBBYTES[4].a/w191 ,
         \SUBBYTES[4].a/w186 , \SUBBYTES[4].a/w184 , \SUBBYTES[4].a/w183 ,
         \SUBBYTES[4].a/w167 , \SUBBYTES[4].a/w166 , \SUBBYTES[4].a/w165 ,
         \SUBBYTES[4].a/w164 , \SUBBYTES[4].a/w163 , \SUBBYTES[4].a/w161 ,
         \SUBBYTES[4].a/w160 , \SUBBYTES[3].a/w3400 , \SUBBYTES[3].a/w3398 ,
         \SUBBYTES[3].a/w3397 , \SUBBYTES[3].a/w3396 , \SUBBYTES[3].a/w3393 ,
         \SUBBYTES[3].a/w3391 , \SUBBYTES[3].a/w3390 , \SUBBYTES[3].a/w3389 ,
         \SUBBYTES[3].a/w3385 , \SUBBYTES[3].a/w3383 , \SUBBYTES[3].a/w3382 ,
         \SUBBYTES[3].a/w3381 , \SUBBYTES[3].a/w3380 , \SUBBYTES[3].a/w3379 ,
         \SUBBYTES[3].a/w3378 , \SUBBYTES[3].a/w3377 , \SUBBYTES[3].a/w3376 ,
         \SUBBYTES[3].a/w3368 , \SUBBYTES[3].a/w3366 , \SUBBYTES[3].a/w3365 ,
         \SUBBYTES[3].a/w3361 , \SUBBYTES[3].a/w3359 , \SUBBYTES[3].a/w3358 ,
         \SUBBYTES[3].a/w3357 , \SUBBYTES[3].a/w3353 , \SUBBYTES[3].a/w3351 ,
         \SUBBYTES[3].a/w3350 , \SUBBYTES[3].a/w3337 , \SUBBYTES[3].a/w3336 ,
         \SUBBYTES[3].a/w3335 , \SUBBYTES[3].a/w3333 , \SUBBYTES[3].a/w3330 ,
         \SUBBYTES[3].a/w3329 , \SUBBYTES[3].a/w3327 , \SUBBYTES[3].a/w3326 ,
         \SUBBYTES[3].a/w3324 , \SUBBYTES[3].a/w3322 , \SUBBYTES[3].a/w3321 ,
         \SUBBYTES[3].a/w3315 , \SUBBYTES[3].a/w3314 , \SUBBYTES[3].a/w3313 ,
         \SUBBYTES[3].a/w3312 , \SUBBYTES[3].a/w3306 , \SUBBYTES[3].a/w3304 ,
         \SUBBYTES[3].a/w3303 , \SUBBYTES[3].a/w3299 , \SUBBYTES[3].a/w3297 ,
         \SUBBYTES[3].a/w3296 , \SUBBYTES[3].a/w3291 , \SUBBYTES[3].a/w3289 ,
         \SUBBYTES[3].a/w3288 , \SUBBYTES[3].a/w3272 , \SUBBYTES[3].a/w3271 ,
         \SUBBYTES[3].a/w3270 , \SUBBYTES[3].a/w3269 , \SUBBYTES[3].a/w3268 ,
         \SUBBYTES[3].a/w3266 , \SUBBYTES[3].a/w3265 , \SUBBYTES[3].a/w3193 ,
         \SUBBYTES[3].a/w3191 , \SUBBYTES[3].a/w3190 , \SUBBYTES[3].a/w3189 ,
         \SUBBYTES[3].a/w3186 , \SUBBYTES[3].a/w3184 , \SUBBYTES[3].a/w3183 ,
         \SUBBYTES[3].a/w3182 , \SUBBYTES[3].a/w3178 , \SUBBYTES[3].a/w3176 ,
         \SUBBYTES[3].a/w3175 , \SUBBYTES[3].a/w3174 , \SUBBYTES[3].a/w3173 ,
         \SUBBYTES[3].a/w3172 , \SUBBYTES[3].a/w3171 , \SUBBYTES[3].a/w3170 ,
         \SUBBYTES[3].a/w3169 , \SUBBYTES[3].a/w3161 , \SUBBYTES[3].a/w3159 ,
         \SUBBYTES[3].a/w3158 , \SUBBYTES[3].a/w3154 , \SUBBYTES[3].a/w3152 ,
         \SUBBYTES[3].a/w3151 , \SUBBYTES[3].a/w3150 , \SUBBYTES[3].a/w3146 ,
         \SUBBYTES[3].a/w3144 , \SUBBYTES[3].a/w3143 , \SUBBYTES[3].a/w3130 ,
         \SUBBYTES[3].a/w3129 , \SUBBYTES[3].a/w3128 , \SUBBYTES[3].a/w3126 ,
         \SUBBYTES[3].a/w3123 , \SUBBYTES[3].a/w3122 , \SUBBYTES[3].a/w3120 ,
         \SUBBYTES[3].a/w3119 , \SUBBYTES[3].a/w3117 , \SUBBYTES[3].a/w3115 ,
         \SUBBYTES[3].a/w3114 , \SUBBYTES[3].a/w3108 , \SUBBYTES[3].a/w3107 ,
         \SUBBYTES[3].a/w3106 , \SUBBYTES[3].a/w3105 , \SUBBYTES[3].a/w3099 ,
         \SUBBYTES[3].a/w3097 , \SUBBYTES[3].a/w3096 , \SUBBYTES[3].a/w3092 ,
         \SUBBYTES[3].a/w3090 , \SUBBYTES[3].a/w3089 , \SUBBYTES[3].a/w3084 ,
         \SUBBYTES[3].a/w3082 , \SUBBYTES[3].a/w3081 , \SUBBYTES[3].a/w3065 ,
         \SUBBYTES[3].a/w3064 , \SUBBYTES[3].a/w3063 , \SUBBYTES[3].a/w3062 ,
         \SUBBYTES[3].a/w3061 , \SUBBYTES[3].a/w3059 , \SUBBYTES[3].a/w3058 ,
         \SUBBYTES[3].a/w2986 , \SUBBYTES[3].a/w2984 , \SUBBYTES[3].a/w2983 ,
         \SUBBYTES[3].a/w2982 , \SUBBYTES[3].a/w2979 , \SUBBYTES[3].a/w2977 ,
         \SUBBYTES[3].a/w2976 , \SUBBYTES[3].a/w2975 , \SUBBYTES[3].a/w2971 ,
         \SUBBYTES[3].a/w2969 , \SUBBYTES[3].a/w2968 , \SUBBYTES[3].a/w2967 ,
         \SUBBYTES[3].a/w2966 , \SUBBYTES[3].a/w2965 , \SUBBYTES[3].a/w2964 ,
         \SUBBYTES[3].a/w2963 , \SUBBYTES[3].a/w2962 , \SUBBYTES[3].a/w2954 ,
         \SUBBYTES[3].a/w2952 , \SUBBYTES[3].a/w2951 , \SUBBYTES[3].a/w2947 ,
         \SUBBYTES[3].a/w2945 , \SUBBYTES[3].a/w2944 , \SUBBYTES[3].a/w2943 ,
         \SUBBYTES[3].a/w2939 , \SUBBYTES[3].a/w2937 , \SUBBYTES[3].a/w2936 ,
         \SUBBYTES[3].a/w2923 , \SUBBYTES[3].a/w2922 , \SUBBYTES[3].a/w2921 ,
         \SUBBYTES[3].a/w2919 , \SUBBYTES[3].a/w2916 , \SUBBYTES[3].a/w2915 ,
         \SUBBYTES[3].a/w2913 , \SUBBYTES[3].a/w2912 , \SUBBYTES[3].a/w2910 ,
         \SUBBYTES[3].a/w2908 , \SUBBYTES[3].a/w2907 , \SUBBYTES[3].a/w2901 ,
         \SUBBYTES[3].a/w2900 , \SUBBYTES[3].a/w2899 , \SUBBYTES[3].a/w2898 ,
         \SUBBYTES[3].a/w2892 , \SUBBYTES[3].a/w2890 , \SUBBYTES[3].a/w2889 ,
         \SUBBYTES[3].a/w2885 , \SUBBYTES[3].a/w2883 , \SUBBYTES[3].a/w2882 ,
         \SUBBYTES[3].a/w2877 , \SUBBYTES[3].a/w2875 , \SUBBYTES[3].a/w2874 ,
         \SUBBYTES[3].a/w2858 , \SUBBYTES[3].a/w2857 , \SUBBYTES[3].a/w2856 ,
         \SUBBYTES[3].a/w2855 , \SUBBYTES[3].a/w2854 , \SUBBYTES[3].a/w2852 ,
         \SUBBYTES[3].a/w2851 , \SUBBYTES[3].a/w2779 , \SUBBYTES[3].a/w2777 ,
         \SUBBYTES[3].a/w2776 , \SUBBYTES[3].a/w2775 , \SUBBYTES[3].a/w2772 ,
         \SUBBYTES[3].a/w2770 , \SUBBYTES[3].a/w2769 , \SUBBYTES[3].a/w2768 ,
         \SUBBYTES[3].a/w2764 , \SUBBYTES[3].a/w2762 , \SUBBYTES[3].a/w2761 ,
         \SUBBYTES[3].a/w2760 , \SUBBYTES[3].a/w2759 , \SUBBYTES[3].a/w2758 ,
         \SUBBYTES[3].a/w2757 , \SUBBYTES[3].a/w2756 , \SUBBYTES[3].a/w2755 ,
         \SUBBYTES[3].a/w2747 , \SUBBYTES[3].a/w2745 , \SUBBYTES[3].a/w2744 ,
         \SUBBYTES[3].a/w2740 , \SUBBYTES[3].a/w2738 , \SUBBYTES[3].a/w2737 ,
         \SUBBYTES[3].a/w2736 , \SUBBYTES[3].a/w2732 , \SUBBYTES[3].a/w2730 ,
         \SUBBYTES[3].a/w2729 , \SUBBYTES[3].a/w2716 , \SUBBYTES[3].a/w2715 ,
         \SUBBYTES[3].a/w2714 , \SUBBYTES[3].a/w2712 , \SUBBYTES[3].a/w2709 ,
         \SUBBYTES[3].a/w2708 , \SUBBYTES[3].a/w2706 , \SUBBYTES[3].a/w2705 ,
         \SUBBYTES[3].a/w2703 , \SUBBYTES[3].a/w2701 , \SUBBYTES[3].a/w2700 ,
         \SUBBYTES[3].a/w2694 , \SUBBYTES[3].a/w2693 , \SUBBYTES[3].a/w2692 ,
         \SUBBYTES[3].a/w2691 , \SUBBYTES[3].a/w2685 , \SUBBYTES[3].a/w2683 ,
         \SUBBYTES[3].a/w2682 , \SUBBYTES[3].a/w2678 , \SUBBYTES[3].a/w2676 ,
         \SUBBYTES[3].a/w2675 , \SUBBYTES[3].a/w2670 , \SUBBYTES[3].a/w2668 ,
         \SUBBYTES[3].a/w2667 , \SUBBYTES[3].a/w2651 , \SUBBYTES[3].a/w2650 ,
         \SUBBYTES[3].a/w2649 , \SUBBYTES[3].a/w2648 , \SUBBYTES[3].a/w2647 ,
         \SUBBYTES[3].a/w2645 , \SUBBYTES[3].a/w2644 , \SUBBYTES[3].a/w2572 ,
         \SUBBYTES[3].a/w2570 , \SUBBYTES[3].a/w2569 , \SUBBYTES[3].a/w2568 ,
         \SUBBYTES[3].a/w2565 , \SUBBYTES[3].a/w2563 , \SUBBYTES[3].a/w2562 ,
         \SUBBYTES[3].a/w2561 , \SUBBYTES[3].a/w2557 , \SUBBYTES[3].a/w2555 ,
         \SUBBYTES[3].a/w2554 , \SUBBYTES[3].a/w2553 , \SUBBYTES[3].a/w2552 ,
         \SUBBYTES[3].a/w2551 , \SUBBYTES[3].a/w2550 , \SUBBYTES[3].a/w2549 ,
         \SUBBYTES[3].a/w2548 , \SUBBYTES[3].a/w2540 , \SUBBYTES[3].a/w2538 ,
         \SUBBYTES[3].a/w2537 , \SUBBYTES[3].a/w2533 , \SUBBYTES[3].a/w2531 ,
         \SUBBYTES[3].a/w2530 , \SUBBYTES[3].a/w2529 , \SUBBYTES[3].a/w2525 ,
         \SUBBYTES[3].a/w2523 , \SUBBYTES[3].a/w2522 , \SUBBYTES[3].a/w2509 ,
         \SUBBYTES[3].a/w2508 , \SUBBYTES[3].a/w2507 , \SUBBYTES[3].a/w2505 ,
         \SUBBYTES[3].a/w2502 , \SUBBYTES[3].a/w2501 , \SUBBYTES[3].a/w2499 ,
         \SUBBYTES[3].a/w2498 , \SUBBYTES[3].a/w2496 , \SUBBYTES[3].a/w2494 ,
         \SUBBYTES[3].a/w2493 , \SUBBYTES[3].a/w2487 , \SUBBYTES[3].a/w2486 ,
         \SUBBYTES[3].a/w2485 , \SUBBYTES[3].a/w2484 , \SUBBYTES[3].a/w2478 ,
         \SUBBYTES[3].a/w2476 , \SUBBYTES[3].a/w2475 , \SUBBYTES[3].a/w2471 ,
         \SUBBYTES[3].a/w2469 , \SUBBYTES[3].a/w2468 , \SUBBYTES[3].a/w2463 ,
         \SUBBYTES[3].a/w2461 , \SUBBYTES[3].a/w2460 , \SUBBYTES[3].a/w2444 ,
         \SUBBYTES[3].a/w2443 , \SUBBYTES[3].a/w2442 , \SUBBYTES[3].a/w2441 ,
         \SUBBYTES[3].a/w2440 , \SUBBYTES[3].a/w2438 , \SUBBYTES[3].a/w2437 ,
         \SUBBYTES[3].a/w2365 , \SUBBYTES[3].a/w2363 , \SUBBYTES[3].a/w2362 ,
         \SUBBYTES[3].a/w2361 , \SUBBYTES[3].a/w2358 , \SUBBYTES[3].a/w2356 ,
         \SUBBYTES[3].a/w2355 , \SUBBYTES[3].a/w2354 , \SUBBYTES[3].a/w2350 ,
         \SUBBYTES[3].a/w2348 , \SUBBYTES[3].a/w2347 , \SUBBYTES[3].a/w2346 ,
         \SUBBYTES[3].a/w2345 , \SUBBYTES[3].a/w2344 , \SUBBYTES[3].a/w2343 ,
         \SUBBYTES[3].a/w2342 , \SUBBYTES[3].a/w2341 , \SUBBYTES[3].a/w2333 ,
         \SUBBYTES[3].a/w2331 , \SUBBYTES[3].a/w2330 , \SUBBYTES[3].a/w2326 ,
         \SUBBYTES[3].a/w2324 , \SUBBYTES[3].a/w2323 , \SUBBYTES[3].a/w2322 ,
         \SUBBYTES[3].a/w2318 , \SUBBYTES[3].a/w2316 , \SUBBYTES[3].a/w2315 ,
         \SUBBYTES[3].a/w2302 , \SUBBYTES[3].a/w2301 , \SUBBYTES[3].a/w2300 ,
         \SUBBYTES[3].a/w2298 , \SUBBYTES[3].a/w2295 , \SUBBYTES[3].a/w2294 ,
         \SUBBYTES[3].a/w2292 , \SUBBYTES[3].a/w2291 , \SUBBYTES[3].a/w2289 ,
         \SUBBYTES[3].a/w2287 , \SUBBYTES[3].a/w2286 , \SUBBYTES[3].a/w2280 ,
         \SUBBYTES[3].a/w2279 , \SUBBYTES[3].a/w2278 , \SUBBYTES[3].a/w2277 ,
         \SUBBYTES[3].a/w2271 , \SUBBYTES[3].a/w2269 , \SUBBYTES[3].a/w2268 ,
         \SUBBYTES[3].a/w2264 , \SUBBYTES[3].a/w2262 , \SUBBYTES[3].a/w2261 ,
         \SUBBYTES[3].a/w2256 , \SUBBYTES[3].a/w2254 , \SUBBYTES[3].a/w2253 ,
         \SUBBYTES[3].a/w2237 , \SUBBYTES[3].a/w2236 , \SUBBYTES[3].a/w2235 ,
         \SUBBYTES[3].a/w2234 , \SUBBYTES[3].a/w2233 , \SUBBYTES[3].a/w2231 ,
         \SUBBYTES[3].a/w2230 , \SUBBYTES[3].a/w2158 , \SUBBYTES[3].a/w2156 ,
         \SUBBYTES[3].a/w2155 , \SUBBYTES[3].a/w2154 , \SUBBYTES[3].a/w2151 ,
         \SUBBYTES[3].a/w2149 , \SUBBYTES[3].a/w2148 , \SUBBYTES[3].a/w2147 ,
         \SUBBYTES[3].a/w2143 , \SUBBYTES[3].a/w2141 , \SUBBYTES[3].a/w2140 ,
         \SUBBYTES[3].a/w2139 , \SUBBYTES[3].a/w2138 , \SUBBYTES[3].a/w2137 ,
         \SUBBYTES[3].a/w2136 , \SUBBYTES[3].a/w2135 , \SUBBYTES[3].a/w2134 ,
         \SUBBYTES[3].a/w2126 , \SUBBYTES[3].a/w2124 , \SUBBYTES[3].a/w2123 ,
         \SUBBYTES[3].a/w2119 , \SUBBYTES[3].a/w2117 , \SUBBYTES[3].a/w2116 ,
         \SUBBYTES[3].a/w2115 , \SUBBYTES[3].a/w2111 , \SUBBYTES[3].a/w2109 ,
         \SUBBYTES[3].a/w2108 , \SUBBYTES[3].a/w2095 , \SUBBYTES[3].a/w2094 ,
         \SUBBYTES[3].a/w2093 , \SUBBYTES[3].a/w2091 , \SUBBYTES[3].a/w2088 ,
         \SUBBYTES[3].a/w2087 , \SUBBYTES[3].a/w2085 , \SUBBYTES[3].a/w2084 ,
         \SUBBYTES[3].a/w2082 , \SUBBYTES[3].a/w2080 , \SUBBYTES[3].a/w2079 ,
         \SUBBYTES[3].a/w2073 , \SUBBYTES[3].a/w2072 , \SUBBYTES[3].a/w2071 ,
         \SUBBYTES[3].a/w2070 , \SUBBYTES[3].a/w2064 , \SUBBYTES[3].a/w2062 ,
         \SUBBYTES[3].a/w2061 , \SUBBYTES[3].a/w2057 , \SUBBYTES[3].a/w2055 ,
         \SUBBYTES[3].a/w2054 , \SUBBYTES[3].a/w2049 , \SUBBYTES[3].a/w2047 ,
         \SUBBYTES[3].a/w2046 , \SUBBYTES[3].a/w2030 , \SUBBYTES[3].a/w2029 ,
         \SUBBYTES[3].a/w2028 , \SUBBYTES[3].a/w2027 , \SUBBYTES[3].a/w2026 ,
         \SUBBYTES[3].a/w2024 , \SUBBYTES[3].a/w2023 , \SUBBYTES[3].a/w1951 ,
         \SUBBYTES[3].a/w1949 , \SUBBYTES[3].a/w1948 , \SUBBYTES[3].a/w1947 ,
         \SUBBYTES[3].a/w1944 , \SUBBYTES[3].a/w1942 , \SUBBYTES[3].a/w1941 ,
         \SUBBYTES[3].a/w1940 , \SUBBYTES[3].a/w1936 , \SUBBYTES[3].a/w1934 ,
         \SUBBYTES[3].a/w1933 , \SUBBYTES[3].a/w1932 , \SUBBYTES[3].a/w1931 ,
         \SUBBYTES[3].a/w1930 , \SUBBYTES[3].a/w1929 , \SUBBYTES[3].a/w1928 ,
         \SUBBYTES[3].a/w1927 , \SUBBYTES[3].a/w1919 , \SUBBYTES[3].a/w1917 ,
         \SUBBYTES[3].a/w1916 , \SUBBYTES[3].a/w1912 , \SUBBYTES[3].a/w1910 ,
         \SUBBYTES[3].a/w1909 , \SUBBYTES[3].a/w1908 , \SUBBYTES[3].a/w1904 ,
         \SUBBYTES[3].a/w1902 , \SUBBYTES[3].a/w1901 , \SUBBYTES[3].a/w1888 ,
         \SUBBYTES[3].a/w1887 , \SUBBYTES[3].a/w1886 , \SUBBYTES[3].a/w1884 ,
         \SUBBYTES[3].a/w1881 , \SUBBYTES[3].a/w1880 , \SUBBYTES[3].a/w1878 ,
         \SUBBYTES[3].a/w1877 , \SUBBYTES[3].a/w1875 , \SUBBYTES[3].a/w1873 ,
         \SUBBYTES[3].a/w1872 , \SUBBYTES[3].a/w1866 , \SUBBYTES[3].a/w1865 ,
         \SUBBYTES[3].a/w1864 , \SUBBYTES[3].a/w1863 , \SUBBYTES[3].a/w1857 ,
         \SUBBYTES[3].a/w1855 , \SUBBYTES[3].a/w1854 , \SUBBYTES[3].a/w1850 ,
         \SUBBYTES[3].a/w1848 , \SUBBYTES[3].a/w1847 , \SUBBYTES[3].a/w1842 ,
         \SUBBYTES[3].a/w1840 , \SUBBYTES[3].a/w1839 , \SUBBYTES[3].a/w1823 ,
         \SUBBYTES[3].a/w1822 , \SUBBYTES[3].a/w1821 , \SUBBYTES[3].a/w1820 ,
         \SUBBYTES[3].a/w1819 , \SUBBYTES[3].a/w1817 , \SUBBYTES[3].a/w1816 ,
         \SUBBYTES[3].a/w1744 , \SUBBYTES[3].a/w1742 , \SUBBYTES[3].a/w1741 ,
         \SUBBYTES[3].a/w1740 , \SUBBYTES[3].a/w1737 , \SUBBYTES[3].a/w1735 ,
         \SUBBYTES[3].a/w1734 , \SUBBYTES[3].a/w1733 , \SUBBYTES[3].a/w1729 ,
         \SUBBYTES[3].a/w1727 , \SUBBYTES[3].a/w1726 , \SUBBYTES[3].a/w1725 ,
         \SUBBYTES[3].a/w1724 , \SUBBYTES[3].a/w1723 , \SUBBYTES[3].a/w1722 ,
         \SUBBYTES[3].a/w1721 , \SUBBYTES[3].a/w1720 , \SUBBYTES[3].a/w1712 ,
         \SUBBYTES[3].a/w1710 , \SUBBYTES[3].a/w1709 , \SUBBYTES[3].a/w1705 ,
         \SUBBYTES[3].a/w1703 , \SUBBYTES[3].a/w1702 , \SUBBYTES[3].a/w1701 ,
         \SUBBYTES[3].a/w1697 , \SUBBYTES[3].a/w1695 , \SUBBYTES[3].a/w1694 ,
         \SUBBYTES[3].a/w1681 , \SUBBYTES[3].a/w1680 , \SUBBYTES[3].a/w1679 ,
         \SUBBYTES[3].a/w1677 , \SUBBYTES[3].a/w1674 , \SUBBYTES[3].a/w1673 ,
         \SUBBYTES[3].a/w1671 , \SUBBYTES[3].a/w1670 , \SUBBYTES[3].a/w1668 ,
         \SUBBYTES[3].a/w1666 , \SUBBYTES[3].a/w1665 , \SUBBYTES[3].a/w1659 ,
         \SUBBYTES[3].a/w1658 , \SUBBYTES[3].a/w1657 , \SUBBYTES[3].a/w1656 ,
         \SUBBYTES[3].a/w1650 , \SUBBYTES[3].a/w1648 , \SUBBYTES[3].a/w1647 ,
         \SUBBYTES[3].a/w1643 , \SUBBYTES[3].a/w1641 , \SUBBYTES[3].a/w1640 ,
         \SUBBYTES[3].a/w1635 , \SUBBYTES[3].a/w1633 , \SUBBYTES[3].a/w1632 ,
         \SUBBYTES[3].a/w1616 , \SUBBYTES[3].a/w1615 , \SUBBYTES[3].a/w1614 ,
         \SUBBYTES[3].a/w1613 , \SUBBYTES[3].a/w1612 , \SUBBYTES[3].a/w1610 ,
         \SUBBYTES[3].a/w1609 , \SUBBYTES[3].a/w1537 , \SUBBYTES[3].a/w1535 ,
         \SUBBYTES[3].a/w1534 , \SUBBYTES[3].a/w1533 , \SUBBYTES[3].a/w1530 ,
         \SUBBYTES[3].a/w1528 , \SUBBYTES[3].a/w1527 , \SUBBYTES[3].a/w1526 ,
         \SUBBYTES[3].a/w1522 , \SUBBYTES[3].a/w1520 , \SUBBYTES[3].a/w1519 ,
         \SUBBYTES[3].a/w1518 , \SUBBYTES[3].a/w1517 , \SUBBYTES[3].a/w1516 ,
         \SUBBYTES[3].a/w1515 , \SUBBYTES[3].a/w1514 , \SUBBYTES[3].a/w1513 ,
         \SUBBYTES[3].a/w1505 , \SUBBYTES[3].a/w1503 , \SUBBYTES[3].a/w1502 ,
         \SUBBYTES[3].a/w1498 , \SUBBYTES[3].a/w1496 , \SUBBYTES[3].a/w1495 ,
         \SUBBYTES[3].a/w1494 , \SUBBYTES[3].a/w1490 , \SUBBYTES[3].a/w1488 ,
         \SUBBYTES[3].a/w1487 , \SUBBYTES[3].a/w1474 , \SUBBYTES[3].a/w1473 ,
         \SUBBYTES[3].a/w1472 , \SUBBYTES[3].a/w1470 , \SUBBYTES[3].a/w1467 ,
         \SUBBYTES[3].a/w1466 , \SUBBYTES[3].a/w1464 , \SUBBYTES[3].a/w1463 ,
         \SUBBYTES[3].a/w1461 , \SUBBYTES[3].a/w1459 , \SUBBYTES[3].a/w1458 ,
         \SUBBYTES[3].a/w1452 , \SUBBYTES[3].a/w1451 , \SUBBYTES[3].a/w1450 ,
         \SUBBYTES[3].a/w1449 , \SUBBYTES[3].a/w1443 , \SUBBYTES[3].a/w1441 ,
         \SUBBYTES[3].a/w1440 , \SUBBYTES[3].a/w1436 , \SUBBYTES[3].a/w1434 ,
         \SUBBYTES[3].a/w1433 , \SUBBYTES[3].a/w1428 , \SUBBYTES[3].a/w1426 ,
         \SUBBYTES[3].a/w1425 , \SUBBYTES[3].a/w1409 , \SUBBYTES[3].a/w1408 ,
         \SUBBYTES[3].a/w1407 , \SUBBYTES[3].a/w1406 , \SUBBYTES[3].a/w1405 ,
         \SUBBYTES[3].a/w1403 , \SUBBYTES[3].a/w1402 , \SUBBYTES[3].a/w1330 ,
         \SUBBYTES[3].a/w1328 , \SUBBYTES[3].a/w1327 , \SUBBYTES[3].a/w1326 ,
         \SUBBYTES[3].a/w1323 , \SUBBYTES[3].a/w1321 , \SUBBYTES[3].a/w1320 ,
         \SUBBYTES[3].a/w1319 , \SUBBYTES[3].a/w1315 , \SUBBYTES[3].a/w1313 ,
         \SUBBYTES[3].a/w1312 , \SUBBYTES[3].a/w1311 , \SUBBYTES[3].a/w1310 ,
         \SUBBYTES[3].a/w1309 , \SUBBYTES[3].a/w1308 , \SUBBYTES[3].a/w1307 ,
         \SUBBYTES[3].a/w1306 , \SUBBYTES[3].a/w1298 , \SUBBYTES[3].a/w1296 ,
         \SUBBYTES[3].a/w1295 , \SUBBYTES[3].a/w1291 , \SUBBYTES[3].a/w1289 ,
         \SUBBYTES[3].a/w1288 , \SUBBYTES[3].a/w1287 , \SUBBYTES[3].a/w1283 ,
         \SUBBYTES[3].a/w1281 , \SUBBYTES[3].a/w1280 , \SUBBYTES[3].a/w1267 ,
         \SUBBYTES[3].a/w1266 , \SUBBYTES[3].a/w1265 , \SUBBYTES[3].a/w1263 ,
         \SUBBYTES[3].a/w1260 , \SUBBYTES[3].a/w1259 , \SUBBYTES[3].a/w1257 ,
         \SUBBYTES[3].a/w1256 , \SUBBYTES[3].a/w1254 , \SUBBYTES[3].a/w1252 ,
         \SUBBYTES[3].a/w1251 , \SUBBYTES[3].a/w1245 , \SUBBYTES[3].a/w1244 ,
         \SUBBYTES[3].a/w1243 , \SUBBYTES[3].a/w1242 , \SUBBYTES[3].a/w1236 ,
         \SUBBYTES[3].a/w1234 , \SUBBYTES[3].a/w1233 , \SUBBYTES[3].a/w1229 ,
         \SUBBYTES[3].a/w1227 , \SUBBYTES[3].a/w1226 , \SUBBYTES[3].a/w1221 ,
         \SUBBYTES[3].a/w1219 , \SUBBYTES[3].a/w1218 , \SUBBYTES[3].a/w1202 ,
         \SUBBYTES[3].a/w1201 , \SUBBYTES[3].a/w1200 , \SUBBYTES[3].a/w1199 ,
         \SUBBYTES[3].a/w1198 , \SUBBYTES[3].a/w1196 , \SUBBYTES[3].a/w1195 ,
         \SUBBYTES[3].a/w1123 , \SUBBYTES[3].a/w1121 , \SUBBYTES[3].a/w1120 ,
         \SUBBYTES[3].a/w1119 , \SUBBYTES[3].a/w1116 , \SUBBYTES[3].a/w1114 ,
         \SUBBYTES[3].a/w1113 , \SUBBYTES[3].a/w1112 , \SUBBYTES[3].a/w1108 ,
         \SUBBYTES[3].a/w1106 , \SUBBYTES[3].a/w1105 , \SUBBYTES[3].a/w1104 ,
         \SUBBYTES[3].a/w1103 , \SUBBYTES[3].a/w1102 , \SUBBYTES[3].a/w1101 ,
         \SUBBYTES[3].a/w1100 , \SUBBYTES[3].a/w1099 , \SUBBYTES[3].a/w1091 ,
         \SUBBYTES[3].a/w1089 , \SUBBYTES[3].a/w1088 , \SUBBYTES[3].a/w1084 ,
         \SUBBYTES[3].a/w1082 , \SUBBYTES[3].a/w1081 , \SUBBYTES[3].a/w1080 ,
         \SUBBYTES[3].a/w1076 , \SUBBYTES[3].a/w1074 , \SUBBYTES[3].a/w1073 ,
         \SUBBYTES[3].a/w1060 , \SUBBYTES[3].a/w1059 , \SUBBYTES[3].a/w1058 ,
         \SUBBYTES[3].a/w1056 , \SUBBYTES[3].a/w1053 , \SUBBYTES[3].a/w1052 ,
         \SUBBYTES[3].a/w1050 , \SUBBYTES[3].a/w1049 , \SUBBYTES[3].a/w1047 ,
         \SUBBYTES[3].a/w1045 , \SUBBYTES[3].a/w1044 , \SUBBYTES[3].a/w1038 ,
         \SUBBYTES[3].a/w1037 , \SUBBYTES[3].a/w1036 , \SUBBYTES[3].a/w1035 ,
         \SUBBYTES[3].a/w1029 , \SUBBYTES[3].a/w1027 , \SUBBYTES[3].a/w1026 ,
         \SUBBYTES[3].a/w1022 , \SUBBYTES[3].a/w1020 , \SUBBYTES[3].a/w1019 ,
         \SUBBYTES[3].a/w1014 , \SUBBYTES[3].a/w1012 , \SUBBYTES[3].a/w1011 ,
         \SUBBYTES[3].a/w995 , \SUBBYTES[3].a/w994 , \SUBBYTES[3].a/w993 ,
         \SUBBYTES[3].a/w992 , \SUBBYTES[3].a/w991 , \SUBBYTES[3].a/w989 ,
         \SUBBYTES[3].a/w988 , \SUBBYTES[3].a/w916 , \SUBBYTES[3].a/w914 ,
         \SUBBYTES[3].a/w913 , \SUBBYTES[3].a/w912 , \SUBBYTES[3].a/w909 ,
         \SUBBYTES[3].a/w907 , \SUBBYTES[3].a/w906 , \SUBBYTES[3].a/w905 ,
         \SUBBYTES[3].a/w901 , \SUBBYTES[3].a/w899 , \SUBBYTES[3].a/w898 ,
         \SUBBYTES[3].a/w897 , \SUBBYTES[3].a/w896 , \SUBBYTES[3].a/w895 ,
         \SUBBYTES[3].a/w894 , \SUBBYTES[3].a/w893 , \SUBBYTES[3].a/w892 ,
         \SUBBYTES[3].a/w884 , \SUBBYTES[3].a/w882 , \SUBBYTES[3].a/w881 ,
         \SUBBYTES[3].a/w877 , \SUBBYTES[3].a/w875 , \SUBBYTES[3].a/w874 ,
         \SUBBYTES[3].a/w873 , \SUBBYTES[3].a/w869 , \SUBBYTES[3].a/w867 ,
         \SUBBYTES[3].a/w866 , \SUBBYTES[3].a/w853 , \SUBBYTES[3].a/w852 ,
         \SUBBYTES[3].a/w851 , \SUBBYTES[3].a/w849 , \SUBBYTES[3].a/w846 ,
         \SUBBYTES[3].a/w845 , \SUBBYTES[3].a/w843 , \SUBBYTES[3].a/w842 ,
         \SUBBYTES[3].a/w840 , \SUBBYTES[3].a/w838 , \SUBBYTES[3].a/w837 ,
         \SUBBYTES[3].a/w831 , \SUBBYTES[3].a/w830 , \SUBBYTES[3].a/w829 ,
         \SUBBYTES[3].a/w828 , \SUBBYTES[3].a/w822 , \SUBBYTES[3].a/w820 ,
         \SUBBYTES[3].a/w819 , \SUBBYTES[3].a/w815 , \SUBBYTES[3].a/w813 ,
         \SUBBYTES[3].a/w812 , \SUBBYTES[3].a/w807 , \SUBBYTES[3].a/w805 ,
         \SUBBYTES[3].a/w804 , \SUBBYTES[3].a/w788 , \SUBBYTES[3].a/w787 ,
         \SUBBYTES[3].a/w786 , \SUBBYTES[3].a/w785 , \SUBBYTES[3].a/w784 ,
         \SUBBYTES[3].a/w782 , \SUBBYTES[3].a/w781 , \SUBBYTES[3].a/w709 ,
         \SUBBYTES[3].a/w707 , \SUBBYTES[3].a/w706 , \SUBBYTES[3].a/w705 ,
         \SUBBYTES[3].a/w702 , \SUBBYTES[3].a/w700 , \SUBBYTES[3].a/w699 ,
         \SUBBYTES[3].a/w698 , \SUBBYTES[3].a/w694 , \SUBBYTES[3].a/w692 ,
         \SUBBYTES[3].a/w691 , \SUBBYTES[3].a/w690 , \SUBBYTES[3].a/w689 ,
         \SUBBYTES[3].a/w688 , \SUBBYTES[3].a/w687 , \SUBBYTES[3].a/w686 ,
         \SUBBYTES[3].a/w685 , \SUBBYTES[3].a/w677 , \SUBBYTES[3].a/w675 ,
         \SUBBYTES[3].a/w674 , \SUBBYTES[3].a/w670 , \SUBBYTES[3].a/w668 ,
         \SUBBYTES[3].a/w667 , \SUBBYTES[3].a/w666 , \SUBBYTES[3].a/w662 ,
         \SUBBYTES[3].a/w660 , \SUBBYTES[3].a/w659 , \SUBBYTES[3].a/w646 ,
         \SUBBYTES[3].a/w645 , \SUBBYTES[3].a/w644 , \SUBBYTES[3].a/w642 ,
         \SUBBYTES[3].a/w639 , \SUBBYTES[3].a/w638 , \SUBBYTES[3].a/w636 ,
         \SUBBYTES[3].a/w635 , \SUBBYTES[3].a/w633 , \SUBBYTES[3].a/w631 ,
         \SUBBYTES[3].a/w630 , \SUBBYTES[3].a/w624 , \SUBBYTES[3].a/w623 ,
         \SUBBYTES[3].a/w622 , \SUBBYTES[3].a/w621 , \SUBBYTES[3].a/w615 ,
         \SUBBYTES[3].a/w613 , \SUBBYTES[3].a/w612 , \SUBBYTES[3].a/w608 ,
         \SUBBYTES[3].a/w606 , \SUBBYTES[3].a/w605 , \SUBBYTES[3].a/w600 ,
         \SUBBYTES[3].a/w598 , \SUBBYTES[3].a/w597 , \SUBBYTES[3].a/w581 ,
         \SUBBYTES[3].a/w580 , \SUBBYTES[3].a/w579 , \SUBBYTES[3].a/w578 ,
         \SUBBYTES[3].a/w577 , \SUBBYTES[3].a/w575 , \SUBBYTES[3].a/w574 ,
         \SUBBYTES[3].a/w502 , \SUBBYTES[3].a/w500 , \SUBBYTES[3].a/w499 ,
         \SUBBYTES[3].a/w498 , \SUBBYTES[3].a/w495 , \SUBBYTES[3].a/w493 ,
         \SUBBYTES[3].a/w492 , \SUBBYTES[3].a/w491 , \SUBBYTES[3].a/w487 ,
         \SUBBYTES[3].a/w485 , \SUBBYTES[3].a/w484 , \SUBBYTES[3].a/w483 ,
         \SUBBYTES[3].a/w482 , \SUBBYTES[3].a/w481 , \SUBBYTES[3].a/w480 ,
         \SUBBYTES[3].a/w479 , \SUBBYTES[3].a/w478 , \SUBBYTES[3].a/w470 ,
         \SUBBYTES[3].a/w468 , \SUBBYTES[3].a/w467 , \SUBBYTES[3].a/w463 ,
         \SUBBYTES[3].a/w461 , \SUBBYTES[3].a/w460 , \SUBBYTES[3].a/w459 ,
         \SUBBYTES[3].a/w455 , \SUBBYTES[3].a/w453 , \SUBBYTES[3].a/w452 ,
         \SUBBYTES[3].a/w439 , \SUBBYTES[3].a/w438 , \SUBBYTES[3].a/w437 ,
         \SUBBYTES[3].a/w435 , \SUBBYTES[3].a/w432 , \SUBBYTES[3].a/w431 ,
         \SUBBYTES[3].a/w429 , \SUBBYTES[3].a/w428 , \SUBBYTES[3].a/w426 ,
         \SUBBYTES[3].a/w424 , \SUBBYTES[3].a/w423 , \SUBBYTES[3].a/w417 ,
         \SUBBYTES[3].a/w416 , \SUBBYTES[3].a/w415 , \SUBBYTES[3].a/w414 ,
         \SUBBYTES[3].a/w408 , \SUBBYTES[3].a/w406 , \SUBBYTES[3].a/w405 ,
         \SUBBYTES[3].a/w401 , \SUBBYTES[3].a/w399 , \SUBBYTES[3].a/w398 ,
         \SUBBYTES[3].a/w393 , \SUBBYTES[3].a/w391 , \SUBBYTES[3].a/w390 ,
         \SUBBYTES[3].a/w374 , \SUBBYTES[3].a/w373 , \SUBBYTES[3].a/w372 ,
         \SUBBYTES[3].a/w371 , \SUBBYTES[3].a/w370 , \SUBBYTES[3].a/w368 ,
         \SUBBYTES[3].a/w367 , \SUBBYTES[3].a/w295 , \SUBBYTES[3].a/w293 ,
         \SUBBYTES[3].a/w292 , \SUBBYTES[3].a/w291 , \SUBBYTES[3].a/w288 ,
         \SUBBYTES[3].a/w286 , \SUBBYTES[3].a/w285 , \SUBBYTES[3].a/w284 ,
         \SUBBYTES[3].a/w280 , \SUBBYTES[3].a/w278 , \SUBBYTES[3].a/w277 ,
         \SUBBYTES[3].a/w276 , \SUBBYTES[3].a/w275 , \SUBBYTES[3].a/w274 ,
         \SUBBYTES[3].a/w273 , \SUBBYTES[3].a/w272 , \SUBBYTES[3].a/w271 ,
         \SUBBYTES[3].a/w263 , \SUBBYTES[3].a/w261 , \SUBBYTES[3].a/w260 ,
         \SUBBYTES[3].a/w256 , \SUBBYTES[3].a/w254 , \SUBBYTES[3].a/w253 ,
         \SUBBYTES[3].a/w252 , \SUBBYTES[3].a/w248 , \SUBBYTES[3].a/w246 ,
         \SUBBYTES[3].a/w245 , \SUBBYTES[3].a/w232 , \SUBBYTES[3].a/w231 ,
         \SUBBYTES[3].a/w230 , \SUBBYTES[3].a/w228 , \SUBBYTES[3].a/w225 ,
         \SUBBYTES[3].a/w224 , \SUBBYTES[3].a/w222 , \SUBBYTES[3].a/w221 ,
         \SUBBYTES[3].a/w219 , \SUBBYTES[3].a/w217 , \SUBBYTES[3].a/w216 ,
         \SUBBYTES[3].a/w210 , \SUBBYTES[3].a/w209 , \SUBBYTES[3].a/w208 ,
         \SUBBYTES[3].a/w207 , \SUBBYTES[3].a/w201 , \SUBBYTES[3].a/w199 ,
         \SUBBYTES[3].a/w198 , \SUBBYTES[3].a/w194 , \SUBBYTES[3].a/w192 ,
         \SUBBYTES[3].a/w191 , \SUBBYTES[3].a/w186 , \SUBBYTES[3].a/w184 ,
         \SUBBYTES[3].a/w183 , \SUBBYTES[3].a/w167 , \SUBBYTES[3].a/w166 ,
         \SUBBYTES[3].a/w165 , \SUBBYTES[3].a/w164 , \SUBBYTES[3].a/w163 ,
         \SUBBYTES[3].a/w161 , \SUBBYTES[3].a/w160 , \SUBBYTES[2].a/w3400 ,
         \SUBBYTES[2].a/w3398 , \SUBBYTES[2].a/w3397 , \SUBBYTES[2].a/w3396 ,
         \SUBBYTES[2].a/w3393 , \SUBBYTES[2].a/w3391 , \SUBBYTES[2].a/w3390 ,
         \SUBBYTES[2].a/w3389 , \SUBBYTES[2].a/w3385 , \SUBBYTES[2].a/w3383 ,
         \SUBBYTES[2].a/w3382 , \SUBBYTES[2].a/w3381 , \SUBBYTES[2].a/w3380 ,
         \SUBBYTES[2].a/w3379 , \SUBBYTES[2].a/w3378 , \SUBBYTES[2].a/w3377 ,
         \SUBBYTES[2].a/w3376 , \SUBBYTES[2].a/w3368 , \SUBBYTES[2].a/w3366 ,
         \SUBBYTES[2].a/w3365 , \SUBBYTES[2].a/w3361 , \SUBBYTES[2].a/w3359 ,
         \SUBBYTES[2].a/w3358 , \SUBBYTES[2].a/w3357 , \SUBBYTES[2].a/w3353 ,
         \SUBBYTES[2].a/w3351 , \SUBBYTES[2].a/w3350 , \SUBBYTES[2].a/w3337 ,
         \SUBBYTES[2].a/w3336 , \SUBBYTES[2].a/w3335 , \SUBBYTES[2].a/w3333 ,
         \SUBBYTES[2].a/w3330 , \SUBBYTES[2].a/w3329 , \SUBBYTES[2].a/w3327 ,
         \SUBBYTES[2].a/w3326 , \SUBBYTES[2].a/w3324 , \SUBBYTES[2].a/w3322 ,
         \SUBBYTES[2].a/w3321 , \SUBBYTES[2].a/w3315 , \SUBBYTES[2].a/w3314 ,
         \SUBBYTES[2].a/w3313 , \SUBBYTES[2].a/w3312 , \SUBBYTES[2].a/w3306 ,
         \SUBBYTES[2].a/w3304 , \SUBBYTES[2].a/w3303 , \SUBBYTES[2].a/w3299 ,
         \SUBBYTES[2].a/w3297 , \SUBBYTES[2].a/w3296 , \SUBBYTES[2].a/w3291 ,
         \SUBBYTES[2].a/w3289 , \SUBBYTES[2].a/w3288 , \SUBBYTES[2].a/w3272 ,
         \SUBBYTES[2].a/w3271 , \SUBBYTES[2].a/w3270 , \SUBBYTES[2].a/w3269 ,
         \SUBBYTES[2].a/w3268 , \SUBBYTES[2].a/w3266 , \SUBBYTES[2].a/w3265 ,
         \SUBBYTES[2].a/w3193 , \SUBBYTES[2].a/w3191 , \SUBBYTES[2].a/w3190 ,
         \SUBBYTES[2].a/w3189 , \SUBBYTES[2].a/w3186 , \SUBBYTES[2].a/w3184 ,
         \SUBBYTES[2].a/w3183 , \SUBBYTES[2].a/w3182 , \SUBBYTES[2].a/w3178 ,
         \SUBBYTES[2].a/w3176 , \SUBBYTES[2].a/w3175 , \SUBBYTES[2].a/w3174 ,
         \SUBBYTES[2].a/w3173 , \SUBBYTES[2].a/w3172 , \SUBBYTES[2].a/w3171 ,
         \SUBBYTES[2].a/w3170 , \SUBBYTES[2].a/w3169 , \SUBBYTES[2].a/w3161 ,
         \SUBBYTES[2].a/w3159 , \SUBBYTES[2].a/w3158 , \SUBBYTES[2].a/w3154 ,
         \SUBBYTES[2].a/w3152 , \SUBBYTES[2].a/w3151 , \SUBBYTES[2].a/w3150 ,
         \SUBBYTES[2].a/w3146 , \SUBBYTES[2].a/w3144 , \SUBBYTES[2].a/w3143 ,
         \SUBBYTES[2].a/w3130 , \SUBBYTES[2].a/w3129 , \SUBBYTES[2].a/w3128 ,
         \SUBBYTES[2].a/w3126 , \SUBBYTES[2].a/w3123 , \SUBBYTES[2].a/w3122 ,
         \SUBBYTES[2].a/w3120 , \SUBBYTES[2].a/w3119 , \SUBBYTES[2].a/w3117 ,
         \SUBBYTES[2].a/w3115 , \SUBBYTES[2].a/w3114 , \SUBBYTES[2].a/w3108 ,
         \SUBBYTES[2].a/w3107 , \SUBBYTES[2].a/w3106 , \SUBBYTES[2].a/w3105 ,
         \SUBBYTES[2].a/w3099 , \SUBBYTES[2].a/w3097 , \SUBBYTES[2].a/w3096 ,
         \SUBBYTES[2].a/w3092 , \SUBBYTES[2].a/w3090 , \SUBBYTES[2].a/w3089 ,
         \SUBBYTES[2].a/w3084 , \SUBBYTES[2].a/w3082 , \SUBBYTES[2].a/w3081 ,
         \SUBBYTES[2].a/w3065 , \SUBBYTES[2].a/w3064 , \SUBBYTES[2].a/w3063 ,
         \SUBBYTES[2].a/w3062 , \SUBBYTES[2].a/w3061 , \SUBBYTES[2].a/w3059 ,
         \SUBBYTES[2].a/w3058 , \SUBBYTES[2].a/w2986 , \SUBBYTES[2].a/w2984 ,
         \SUBBYTES[2].a/w2983 , \SUBBYTES[2].a/w2982 , \SUBBYTES[2].a/w2979 ,
         \SUBBYTES[2].a/w2977 , \SUBBYTES[2].a/w2976 , \SUBBYTES[2].a/w2975 ,
         \SUBBYTES[2].a/w2971 , \SUBBYTES[2].a/w2969 , \SUBBYTES[2].a/w2968 ,
         \SUBBYTES[2].a/w2967 , \SUBBYTES[2].a/w2966 , \SUBBYTES[2].a/w2965 ,
         \SUBBYTES[2].a/w2964 , \SUBBYTES[2].a/w2963 , \SUBBYTES[2].a/w2962 ,
         \SUBBYTES[2].a/w2954 , \SUBBYTES[2].a/w2952 , \SUBBYTES[2].a/w2951 ,
         \SUBBYTES[2].a/w2947 , \SUBBYTES[2].a/w2945 , \SUBBYTES[2].a/w2944 ,
         \SUBBYTES[2].a/w2943 , \SUBBYTES[2].a/w2939 , \SUBBYTES[2].a/w2937 ,
         \SUBBYTES[2].a/w2936 , \SUBBYTES[2].a/w2923 , \SUBBYTES[2].a/w2922 ,
         \SUBBYTES[2].a/w2921 , \SUBBYTES[2].a/w2919 , \SUBBYTES[2].a/w2916 ,
         \SUBBYTES[2].a/w2915 , \SUBBYTES[2].a/w2913 , \SUBBYTES[2].a/w2912 ,
         \SUBBYTES[2].a/w2910 , \SUBBYTES[2].a/w2908 , \SUBBYTES[2].a/w2907 ,
         \SUBBYTES[2].a/w2901 , \SUBBYTES[2].a/w2900 , \SUBBYTES[2].a/w2899 ,
         \SUBBYTES[2].a/w2898 , \SUBBYTES[2].a/w2892 , \SUBBYTES[2].a/w2890 ,
         \SUBBYTES[2].a/w2889 , \SUBBYTES[2].a/w2885 , \SUBBYTES[2].a/w2883 ,
         \SUBBYTES[2].a/w2882 , \SUBBYTES[2].a/w2877 , \SUBBYTES[2].a/w2875 ,
         \SUBBYTES[2].a/w2874 , \SUBBYTES[2].a/w2858 , \SUBBYTES[2].a/w2857 ,
         \SUBBYTES[2].a/w2856 , \SUBBYTES[2].a/w2855 , \SUBBYTES[2].a/w2854 ,
         \SUBBYTES[2].a/w2852 , \SUBBYTES[2].a/w2851 , \SUBBYTES[2].a/w2779 ,
         \SUBBYTES[2].a/w2777 , \SUBBYTES[2].a/w2776 , \SUBBYTES[2].a/w2775 ,
         \SUBBYTES[2].a/w2772 , \SUBBYTES[2].a/w2770 , \SUBBYTES[2].a/w2769 ,
         \SUBBYTES[2].a/w2768 , \SUBBYTES[2].a/w2764 , \SUBBYTES[2].a/w2762 ,
         \SUBBYTES[2].a/w2761 , \SUBBYTES[2].a/w2760 , \SUBBYTES[2].a/w2759 ,
         \SUBBYTES[2].a/w2758 , \SUBBYTES[2].a/w2757 , \SUBBYTES[2].a/w2756 ,
         \SUBBYTES[2].a/w2755 , \SUBBYTES[2].a/w2747 , \SUBBYTES[2].a/w2745 ,
         \SUBBYTES[2].a/w2744 , \SUBBYTES[2].a/w2740 , \SUBBYTES[2].a/w2738 ,
         \SUBBYTES[2].a/w2737 , \SUBBYTES[2].a/w2736 , \SUBBYTES[2].a/w2732 ,
         \SUBBYTES[2].a/w2730 , \SUBBYTES[2].a/w2729 , \SUBBYTES[2].a/w2716 ,
         \SUBBYTES[2].a/w2715 , \SUBBYTES[2].a/w2714 , \SUBBYTES[2].a/w2712 ,
         \SUBBYTES[2].a/w2709 , \SUBBYTES[2].a/w2708 , \SUBBYTES[2].a/w2706 ,
         \SUBBYTES[2].a/w2705 , \SUBBYTES[2].a/w2703 , \SUBBYTES[2].a/w2701 ,
         \SUBBYTES[2].a/w2700 , \SUBBYTES[2].a/w2694 , \SUBBYTES[2].a/w2693 ,
         \SUBBYTES[2].a/w2692 , \SUBBYTES[2].a/w2691 , \SUBBYTES[2].a/w2685 ,
         \SUBBYTES[2].a/w2683 , \SUBBYTES[2].a/w2682 , \SUBBYTES[2].a/w2678 ,
         \SUBBYTES[2].a/w2676 , \SUBBYTES[2].a/w2675 , \SUBBYTES[2].a/w2670 ,
         \SUBBYTES[2].a/w2668 , \SUBBYTES[2].a/w2667 , \SUBBYTES[2].a/w2651 ,
         \SUBBYTES[2].a/w2650 , \SUBBYTES[2].a/w2649 , \SUBBYTES[2].a/w2648 ,
         \SUBBYTES[2].a/w2647 , \SUBBYTES[2].a/w2645 , \SUBBYTES[2].a/w2644 ,
         \SUBBYTES[2].a/w2572 , \SUBBYTES[2].a/w2570 , \SUBBYTES[2].a/w2569 ,
         \SUBBYTES[2].a/w2568 , \SUBBYTES[2].a/w2565 , \SUBBYTES[2].a/w2563 ,
         \SUBBYTES[2].a/w2562 , \SUBBYTES[2].a/w2561 , \SUBBYTES[2].a/w2557 ,
         \SUBBYTES[2].a/w2555 , \SUBBYTES[2].a/w2554 , \SUBBYTES[2].a/w2553 ,
         \SUBBYTES[2].a/w2552 , \SUBBYTES[2].a/w2551 , \SUBBYTES[2].a/w2550 ,
         \SUBBYTES[2].a/w2549 , \SUBBYTES[2].a/w2548 , \SUBBYTES[2].a/w2540 ,
         \SUBBYTES[2].a/w2538 , \SUBBYTES[2].a/w2537 , \SUBBYTES[2].a/w2533 ,
         \SUBBYTES[2].a/w2531 , \SUBBYTES[2].a/w2530 , \SUBBYTES[2].a/w2529 ,
         \SUBBYTES[2].a/w2525 , \SUBBYTES[2].a/w2523 , \SUBBYTES[2].a/w2522 ,
         \SUBBYTES[2].a/w2509 , \SUBBYTES[2].a/w2508 , \SUBBYTES[2].a/w2507 ,
         \SUBBYTES[2].a/w2505 , \SUBBYTES[2].a/w2502 , \SUBBYTES[2].a/w2501 ,
         \SUBBYTES[2].a/w2499 , \SUBBYTES[2].a/w2498 , \SUBBYTES[2].a/w2496 ,
         \SUBBYTES[2].a/w2494 , \SUBBYTES[2].a/w2493 , \SUBBYTES[2].a/w2487 ,
         \SUBBYTES[2].a/w2486 , \SUBBYTES[2].a/w2485 , \SUBBYTES[2].a/w2484 ,
         \SUBBYTES[2].a/w2478 , \SUBBYTES[2].a/w2476 , \SUBBYTES[2].a/w2475 ,
         \SUBBYTES[2].a/w2471 , \SUBBYTES[2].a/w2469 , \SUBBYTES[2].a/w2468 ,
         \SUBBYTES[2].a/w2463 , \SUBBYTES[2].a/w2461 , \SUBBYTES[2].a/w2460 ,
         \SUBBYTES[2].a/w2444 , \SUBBYTES[2].a/w2443 , \SUBBYTES[2].a/w2442 ,
         \SUBBYTES[2].a/w2441 , \SUBBYTES[2].a/w2440 , \SUBBYTES[2].a/w2438 ,
         \SUBBYTES[2].a/w2437 , \SUBBYTES[2].a/w2365 , \SUBBYTES[2].a/w2363 ,
         \SUBBYTES[2].a/w2362 , \SUBBYTES[2].a/w2361 , \SUBBYTES[2].a/w2358 ,
         \SUBBYTES[2].a/w2356 , \SUBBYTES[2].a/w2355 , \SUBBYTES[2].a/w2354 ,
         \SUBBYTES[2].a/w2350 , \SUBBYTES[2].a/w2348 , \SUBBYTES[2].a/w2347 ,
         \SUBBYTES[2].a/w2346 , \SUBBYTES[2].a/w2345 , \SUBBYTES[2].a/w2344 ,
         \SUBBYTES[2].a/w2343 , \SUBBYTES[2].a/w2342 , \SUBBYTES[2].a/w2341 ,
         \SUBBYTES[2].a/w2333 , \SUBBYTES[2].a/w2331 , \SUBBYTES[2].a/w2330 ,
         \SUBBYTES[2].a/w2326 , \SUBBYTES[2].a/w2324 , \SUBBYTES[2].a/w2323 ,
         \SUBBYTES[2].a/w2322 , \SUBBYTES[2].a/w2318 , \SUBBYTES[2].a/w2316 ,
         \SUBBYTES[2].a/w2315 , \SUBBYTES[2].a/w2302 , \SUBBYTES[2].a/w2301 ,
         \SUBBYTES[2].a/w2300 , \SUBBYTES[2].a/w2298 , \SUBBYTES[2].a/w2295 ,
         \SUBBYTES[2].a/w2294 , \SUBBYTES[2].a/w2292 , \SUBBYTES[2].a/w2291 ,
         \SUBBYTES[2].a/w2289 , \SUBBYTES[2].a/w2287 , \SUBBYTES[2].a/w2286 ,
         \SUBBYTES[2].a/w2280 , \SUBBYTES[2].a/w2279 , \SUBBYTES[2].a/w2278 ,
         \SUBBYTES[2].a/w2277 , \SUBBYTES[2].a/w2271 , \SUBBYTES[2].a/w2269 ,
         \SUBBYTES[2].a/w2268 , \SUBBYTES[2].a/w2264 , \SUBBYTES[2].a/w2262 ,
         \SUBBYTES[2].a/w2261 , \SUBBYTES[2].a/w2256 , \SUBBYTES[2].a/w2254 ,
         \SUBBYTES[2].a/w2253 , \SUBBYTES[2].a/w2237 , \SUBBYTES[2].a/w2236 ,
         \SUBBYTES[2].a/w2235 , \SUBBYTES[2].a/w2234 , \SUBBYTES[2].a/w2233 ,
         \SUBBYTES[2].a/w2231 , \SUBBYTES[2].a/w2230 , \SUBBYTES[2].a/w2158 ,
         \SUBBYTES[2].a/w2156 , \SUBBYTES[2].a/w2155 , \SUBBYTES[2].a/w2154 ,
         \SUBBYTES[2].a/w2151 , \SUBBYTES[2].a/w2149 , \SUBBYTES[2].a/w2148 ,
         \SUBBYTES[2].a/w2147 , \SUBBYTES[2].a/w2143 , \SUBBYTES[2].a/w2141 ,
         \SUBBYTES[2].a/w2140 , \SUBBYTES[2].a/w2139 , \SUBBYTES[2].a/w2138 ,
         \SUBBYTES[2].a/w2137 , \SUBBYTES[2].a/w2136 , \SUBBYTES[2].a/w2135 ,
         \SUBBYTES[2].a/w2134 , \SUBBYTES[2].a/w2126 , \SUBBYTES[2].a/w2124 ,
         \SUBBYTES[2].a/w2123 , \SUBBYTES[2].a/w2119 , \SUBBYTES[2].a/w2117 ,
         \SUBBYTES[2].a/w2116 , \SUBBYTES[2].a/w2115 , \SUBBYTES[2].a/w2111 ,
         \SUBBYTES[2].a/w2109 , \SUBBYTES[2].a/w2108 , \SUBBYTES[2].a/w2095 ,
         \SUBBYTES[2].a/w2094 , \SUBBYTES[2].a/w2093 , \SUBBYTES[2].a/w2091 ,
         \SUBBYTES[2].a/w2088 , \SUBBYTES[2].a/w2087 , \SUBBYTES[2].a/w2085 ,
         \SUBBYTES[2].a/w2084 , \SUBBYTES[2].a/w2082 , \SUBBYTES[2].a/w2080 ,
         \SUBBYTES[2].a/w2079 , \SUBBYTES[2].a/w2073 , \SUBBYTES[2].a/w2072 ,
         \SUBBYTES[2].a/w2071 , \SUBBYTES[2].a/w2070 , \SUBBYTES[2].a/w2064 ,
         \SUBBYTES[2].a/w2062 , \SUBBYTES[2].a/w2061 , \SUBBYTES[2].a/w2057 ,
         \SUBBYTES[2].a/w2055 , \SUBBYTES[2].a/w2054 , \SUBBYTES[2].a/w2049 ,
         \SUBBYTES[2].a/w2047 , \SUBBYTES[2].a/w2046 , \SUBBYTES[2].a/w2030 ,
         \SUBBYTES[2].a/w2029 , \SUBBYTES[2].a/w2028 , \SUBBYTES[2].a/w2027 ,
         \SUBBYTES[2].a/w2026 , \SUBBYTES[2].a/w2024 , \SUBBYTES[2].a/w2023 ,
         \SUBBYTES[2].a/w1951 , \SUBBYTES[2].a/w1949 , \SUBBYTES[2].a/w1948 ,
         \SUBBYTES[2].a/w1947 , \SUBBYTES[2].a/w1944 , \SUBBYTES[2].a/w1942 ,
         \SUBBYTES[2].a/w1941 , \SUBBYTES[2].a/w1940 , \SUBBYTES[2].a/w1936 ,
         \SUBBYTES[2].a/w1934 , \SUBBYTES[2].a/w1933 , \SUBBYTES[2].a/w1932 ,
         \SUBBYTES[2].a/w1931 , \SUBBYTES[2].a/w1930 , \SUBBYTES[2].a/w1929 ,
         \SUBBYTES[2].a/w1928 , \SUBBYTES[2].a/w1927 , \SUBBYTES[2].a/w1919 ,
         \SUBBYTES[2].a/w1917 , \SUBBYTES[2].a/w1916 , \SUBBYTES[2].a/w1912 ,
         \SUBBYTES[2].a/w1910 , \SUBBYTES[2].a/w1909 , \SUBBYTES[2].a/w1908 ,
         \SUBBYTES[2].a/w1904 , \SUBBYTES[2].a/w1902 , \SUBBYTES[2].a/w1901 ,
         \SUBBYTES[2].a/w1888 , \SUBBYTES[2].a/w1887 , \SUBBYTES[2].a/w1886 ,
         \SUBBYTES[2].a/w1884 , \SUBBYTES[2].a/w1881 , \SUBBYTES[2].a/w1880 ,
         \SUBBYTES[2].a/w1878 , \SUBBYTES[2].a/w1877 , \SUBBYTES[2].a/w1875 ,
         \SUBBYTES[2].a/w1873 , \SUBBYTES[2].a/w1872 , \SUBBYTES[2].a/w1866 ,
         \SUBBYTES[2].a/w1865 , \SUBBYTES[2].a/w1864 , \SUBBYTES[2].a/w1863 ,
         \SUBBYTES[2].a/w1857 , \SUBBYTES[2].a/w1855 , \SUBBYTES[2].a/w1854 ,
         \SUBBYTES[2].a/w1850 , \SUBBYTES[2].a/w1848 , \SUBBYTES[2].a/w1847 ,
         \SUBBYTES[2].a/w1842 , \SUBBYTES[2].a/w1840 , \SUBBYTES[2].a/w1839 ,
         \SUBBYTES[2].a/w1823 , \SUBBYTES[2].a/w1822 , \SUBBYTES[2].a/w1821 ,
         \SUBBYTES[2].a/w1820 , \SUBBYTES[2].a/w1819 , \SUBBYTES[2].a/w1817 ,
         \SUBBYTES[2].a/w1816 , \SUBBYTES[2].a/w1744 , \SUBBYTES[2].a/w1742 ,
         \SUBBYTES[2].a/w1741 , \SUBBYTES[2].a/w1740 , \SUBBYTES[2].a/w1737 ,
         \SUBBYTES[2].a/w1735 , \SUBBYTES[2].a/w1734 , \SUBBYTES[2].a/w1733 ,
         \SUBBYTES[2].a/w1729 , \SUBBYTES[2].a/w1727 , \SUBBYTES[2].a/w1726 ,
         \SUBBYTES[2].a/w1725 , \SUBBYTES[2].a/w1724 , \SUBBYTES[2].a/w1723 ,
         \SUBBYTES[2].a/w1722 , \SUBBYTES[2].a/w1721 , \SUBBYTES[2].a/w1720 ,
         \SUBBYTES[2].a/w1712 , \SUBBYTES[2].a/w1710 , \SUBBYTES[2].a/w1709 ,
         \SUBBYTES[2].a/w1705 , \SUBBYTES[2].a/w1703 , \SUBBYTES[2].a/w1702 ,
         \SUBBYTES[2].a/w1701 , \SUBBYTES[2].a/w1697 , \SUBBYTES[2].a/w1695 ,
         \SUBBYTES[2].a/w1694 , \SUBBYTES[2].a/w1681 , \SUBBYTES[2].a/w1680 ,
         \SUBBYTES[2].a/w1679 , \SUBBYTES[2].a/w1677 , \SUBBYTES[2].a/w1674 ,
         \SUBBYTES[2].a/w1673 , \SUBBYTES[2].a/w1671 , \SUBBYTES[2].a/w1670 ,
         \SUBBYTES[2].a/w1668 , \SUBBYTES[2].a/w1666 , \SUBBYTES[2].a/w1665 ,
         \SUBBYTES[2].a/w1659 , \SUBBYTES[2].a/w1658 , \SUBBYTES[2].a/w1657 ,
         \SUBBYTES[2].a/w1656 , \SUBBYTES[2].a/w1650 , \SUBBYTES[2].a/w1648 ,
         \SUBBYTES[2].a/w1647 , \SUBBYTES[2].a/w1643 , \SUBBYTES[2].a/w1641 ,
         \SUBBYTES[2].a/w1640 , \SUBBYTES[2].a/w1635 , \SUBBYTES[2].a/w1633 ,
         \SUBBYTES[2].a/w1632 , \SUBBYTES[2].a/w1616 , \SUBBYTES[2].a/w1615 ,
         \SUBBYTES[2].a/w1614 , \SUBBYTES[2].a/w1613 , \SUBBYTES[2].a/w1612 ,
         \SUBBYTES[2].a/w1610 , \SUBBYTES[2].a/w1609 , \SUBBYTES[2].a/w1537 ,
         \SUBBYTES[2].a/w1535 , \SUBBYTES[2].a/w1534 , \SUBBYTES[2].a/w1533 ,
         \SUBBYTES[2].a/w1530 , \SUBBYTES[2].a/w1528 , \SUBBYTES[2].a/w1527 ,
         \SUBBYTES[2].a/w1526 , \SUBBYTES[2].a/w1522 , \SUBBYTES[2].a/w1520 ,
         \SUBBYTES[2].a/w1519 , \SUBBYTES[2].a/w1518 , \SUBBYTES[2].a/w1517 ,
         \SUBBYTES[2].a/w1516 , \SUBBYTES[2].a/w1515 , \SUBBYTES[2].a/w1514 ,
         \SUBBYTES[2].a/w1513 , \SUBBYTES[2].a/w1505 , \SUBBYTES[2].a/w1503 ,
         \SUBBYTES[2].a/w1502 , \SUBBYTES[2].a/w1498 , \SUBBYTES[2].a/w1496 ,
         \SUBBYTES[2].a/w1495 , \SUBBYTES[2].a/w1494 , \SUBBYTES[2].a/w1490 ,
         \SUBBYTES[2].a/w1488 , \SUBBYTES[2].a/w1487 , \SUBBYTES[2].a/w1474 ,
         \SUBBYTES[2].a/w1473 , \SUBBYTES[2].a/w1472 , \SUBBYTES[2].a/w1470 ,
         \SUBBYTES[2].a/w1467 , \SUBBYTES[2].a/w1466 , \SUBBYTES[2].a/w1464 ,
         \SUBBYTES[2].a/w1463 , \SUBBYTES[2].a/w1461 , \SUBBYTES[2].a/w1459 ,
         \SUBBYTES[2].a/w1458 , \SUBBYTES[2].a/w1452 , \SUBBYTES[2].a/w1451 ,
         \SUBBYTES[2].a/w1450 , \SUBBYTES[2].a/w1449 , \SUBBYTES[2].a/w1443 ,
         \SUBBYTES[2].a/w1441 , \SUBBYTES[2].a/w1440 , \SUBBYTES[2].a/w1436 ,
         \SUBBYTES[2].a/w1434 , \SUBBYTES[2].a/w1433 , \SUBBYTES[2].a/w1428 ,
         \SUBBYTES[2].a/w1426 , \SUBBYTES[2].a/w1425 , \SUBBYTES[2].a/w1409 ,
         \SUBBYTES[2].a/w1408 , \SUBBYTES[2].a/w1407 , \SUBBYTES[2].a/w1406 ,
         \SUBBYTES[2].a/w1405 , \SUBBYTES[2].a/w1403 , \SUBBYTES[2].a/w1402 ,
         \SUBBYTES[2].a/w1330 , \SUBBYTES[2].a/w1328 , \SUBBYTES[2].a/w1327 ,
         \SUBBYTES[2].a/w1326 , \SUBBYTES[2].a/w1323 , \SUBBYTES[2].a/w1321 ,
         \SUBBYTES[2].a/w1320 , \SUBBYTES[2].a/w1319 , \SUBBYTES[2].a/w1315 ,
         \SUBBYTES[2].a/w1313 , \SUBBYTES[2].a/w1312 , \SUBBYTES[2].a/w1311 ,
         \SUBBYTES[2].a/w1310 , \SUBBYTES[2].a/w1309 , \SUBBYTES[2].a/w1308 ,
         \SUBBYTES[2].a/w1307 , \SUBBYTES[2].a/w1306 , \SUBBYTES[2].a/w1298 ,
         \SUBBYTES[2].a/w1296 , \SUBBYTES[2].a/w1295 , \SUBBYTES[2].a/w1291 ,
         \SUBBYTES[2].a/w1289 , \SUBBYTES[2].a/w1288 , \SUBBYTES[2].a/w1287 ,
         \SUBBYTES[2].a/w1283 , \SUBBYTES[2].a/w1281 , \SUBBYTES[2].a/w1280 ,
         \SUBBYTES[2].a/w1267 , \SUBBYTES[2].a/w1266 , \SUBBYTES[2].a/w1265 ,
         \SUBBYTES[2].a/w1263 , \SUBBYTES[2].a/w1260 , \SUBBYTES[2].a/w1259 ,
         \SUBBYTES[2].a/w1257 , \SUBBYTES[2].a/w1256 , \SUBBYTES[2].a/w1254 ,
         \SUBBYTES[2].a/w1252 , \SUBBYTES[2].a/w1251 , \SUBBYTES[2].a/w1245 ,
         \SUBBYTES[2].a/w1244 , \SUBBYTES[2].a/w1243 , \SUBBYTES[2].a/w1242 ,
         \SUBBYTES[2].a/w1236 , \SUBBYTES[2].a/w1234 , \SUBBYTES[2].a/w1233 ,
         \SUBBYTES[2].a/w1229 , \SUBBYTES[2].a/w1227 , \SUBBYTES[2].a/w1226 ,
         \SUBBYTES[2].a/w1221 , \SUBBYTES[2].a/w1219 , \SUBBYTES[2].a/w1218 ,
         \SUBBYTES[2].a/w1202 , \SUBBYTES[2].a/w1201 , \SUBBYTES[2].a/w1200 ,
         \SUBBYTES[2].a/w1199 , \SUBBYTES[2].a/w1198 , \SUBBYTES[2].a/w1196 ,
         \SUBBYTES[2].a/w1195 , \SUBBYTES[2].a/w1123 , \SUBBYTES[2].a/w1121 ,
         \SUBBYTES[2].a/w1120 , \SUBBYTES[2].a/w1119 , \SUBBYTES[2].a/w1116 ,
         \SUBBYTES[2].a/w1114 , \SUBBYTES[2].a/w1113 , \SUBBYTES[2].a/w1112 ,
         \SUBBYTES[2].a/w1108 , \SUBBYTES[2].a/w1106 , \SUBBYTES[2].a/w1105 ,
         \SUBBYTES[2].a/w1104 , \SUBBYTES[2].a/w1103 , \SUBBYTES[2].a/w1102 ,
         \SUBBYTES[2].a/w1101 , \SUBBYTES[2].a/w1100 , \SUBBYTES[2].a/w1099 ,
         \SUBBYTES[2].a/w1091 , \SUBBYTES[2].a/w1089 , \SUBBYTES[2].a/w1088 ,
         \SUBBYTES[2].a/w1084 , \SUBBYTES[2].a/w1082 , \SUBBYTES[2].a/w1081 ,
         \SUBBYTES[2].a/w1080 , \SUBBYTES[2].a/w1076 , \SUBBYTES[2].a/w1074 ,
         \SUBBYTES[2].a/w1073 , \SUBBYTES[2].a/w1060 , \SUBBYTES[2].a/w1059 ,
         \SUBBYTES[2].a/w1058 , \SUBBYTES[2].a/w1056 , \SUBBYTES[2].a/w1053 ,
         \SUBBYTES[2].a/w1052 , \SUBBYTES[2].a/w1050 , \SUBBYTES[2].a/w1049 ,
         \SUBBYTES[2].a/w1047 , \SUBBYTES[2].a/w1045 , \SUBBYTES[2].a/w1044 ,
         \SUBBYTES[2].a/w1038 , \SUBBYTES[2].a/w1037 , \SUBBYTES[2].a/w1036 ,
         \SUBBYTES[2].a/w1035 , \SUBBYTES[2].a/w1029 , \SUBBYTES[2].a/w1027 ,
         \SUBBYTES[2].a/w1026 , \SUBBYTES[2].a/w1022 , \SUBBYTES[2].a/w1020 ,
         \SUBBYTES[2].a/w1019 , \SUBBYTES[2].a/w1014 , \SUBBYTES[2].a/w1012 ,
         \SUBBYTES[2].a/w1011 , \SUBBYTES[2].a/w995 , \SUBBYTES[2].a/w994 ,
         \SUBBYTES[2].a/w993 , \SUBBYTES[2].a/w992 , \SUBBYTES[2].a/w991 ,
         \SUBBYTES[2].a/w989 , \SUBBYTES[2].a/w988 , \SUBBYTES[2].a/w916 ,
         \SUBBYTES[2].a/w914 , \SUBBYTES[2].a/w913 , \SUBBYTES[2].a/w912 ,
         \SUBBYTES[2].a/w909 , \SUBBYTES[2].a/w907 , \SUBBYTES[2].a/w906 ,
         \SUBBYTES[2].a/w905 , \SUBBYTES[2].a/w901 , \SUBBYTES[2].a/w899 ,
         \SUBBYTES[2].a/w898 , \SUBBYTES[2].a/w897 , \SUBBYTES[2].a/w896 ,
         \SUBBYTES[2].a/w895 , \SUBBYTES[2].a/w894 , \SUBBYTES[2].a/w893 ,
         \SUBBYTES[2].a/w892 , \SUBBYTES[2].a/w884 , \SUBBYTES[2].a/w882 ,
         \SUBBYTES[2].a/w881 , \SUBBYTES[2].a/w877 , \SUBBYTES[2].a/w875 ,
         \SUBBYTES[2].a/w874 , \SUBBYTES[2].a/w873 , \SUBBYTES[2].a/w869 ,
         \SUBBYTES[2].a/w867 , \SUBBYTES[2].a/w866 , \SUBBYTES[2].a/w853 ,
         \SUBBYTES[2].a/w852 , \SUBBYTES[2].a/w851 , \SUBBYTES[2].a/w849 ,
         \SUBBYTES[2].a/w846 , \SUBBYTES[2].a/w845 , \SUBBYTES[2].a/w843 ,
         \SUBBYTES[2].a/w842 , \SUBBYTES[2].a/w840 , \SUBBYTES[2].a/w838 ,
         \SUBBYTES[2].a/w837 , \SUBBYTES[2].a/w831 , \SUBBYTES[2].a/w830 ,
         \SUBBYTES[2].a/w829 , \SUBBYTES[2].a/w828 , \SUBBYTES[2].a/w822 ,
         \SUBBYTES[2].a/w820 , \SUBBYTES[2].a/w819 , \SUBBYTES[2].a/w815 ,
         \SUBBYTES[2].a/w813 , \SUBBYTES[2].a/w812 , \SUBBYTES[2].a/w807 ,
         \SUBBYTES[2].a/w805 , \SUBBYTES[2].a/w804 , \SUBBYTES[2].a/w788 ,
         \SUBBYTES[2].a/w787 , \SUBBYTES[2].a/w786 , \SUBBYTES[2].a/w785 ,
         \SUBBYTES[2].a/w784 , \SUBBYTES[2].a/w782 , \SUBBYTES[2].a/w781 ,
         \SUBBYTES[2].a/w709 , \SUBBYTES[2].a/w707 , \SUBBYTES[2].a/w706 ,
         \SUBBYTES[2].a/w705 , \SUBBYTES[2].a/w702 , \SUBBYTES[2].a/w700 ,
         \SUBBYTES[2].a/w699 , \SUBBYTES[2].a/w698 , \SUBBYTES[2].a/w694 ,
         \SUBBYTES[2].a/w692 , \SUBBYTES[2].a/w691 , \SUBBYTES[2].a/w690 ,
         \SUBBYTES[2].a/w689 , \SUBBYTES[2].a/w688 , \SUBBYTES[2].a/w687 ,
         \SUBBYTES[2].a/w686 , \SUBBYTES[2].a/w685 , \SUBBYTES[2].a/w677 ,
         \SUBBYTES[2].a/w675 , \SUBBYTES[2].a/w674 , \SUBBYTES[2].a/w670 ,
         \SUBBYTES[2].a/w668 , \SUBBYTES[2].a/w667 , \SUBBYTES[2].a/w666 ,
         \SUBBYTES[2].a/w662 , \SUBBYTES[2].a/w660 , \SUBBYTES[2].a/w659 ,
         \SUBBYTES[2].a/w646 , \SUBBYTES[2].a/w645 , \SUBBYTES[2].a/w644 ,
         \SUBBYTES[2].a/w642 , \SUBBYTES[2].a/w639 , \SUBBYTES[2].a/w638 ,
         \SUBBYTES[2].a/w636 , \SUBBYTES[2].a/w635 , \SUBBYTES[2].a/w633 ,
         \SUBBYTES[2].a/w631 , \SUBBYTES[2].a/w630 , \SUBBYTES[2].a/w624 ,
         \SUBBYTES[2].a/w623 , \SUBBYTES[2].a/w622 , \SUBBYTES[2].a/w621 ,
         \SUBBYTES[2].a/w615 , \SUBBYTES[2].a/w613 , \SUBBYTES[2].a/w612 ,
         \SUBBYTES[2].a/w608 , \SUBBYTES[2].a/w606 , \SUBBYTES[2].a/w605 ,
         \SUBBYTES[2].a/w600 , \SUBBYTES[2].a/w598 , \SUBBYTES[2].a/w597 ,
         \SUBBYTES[2].a/w581 , \SUBBYTES[2].a/w580 , \SUBBYTES[2].a/w579 ,
         \SUBBYTES[2].a/w578 , \SUBBYTES[2].a/w577 , \SUBBYTES[2].a/w575 ,
         \SUBBYTES[2].a/w574 , \SUBBYTES[2].a/w502 , \SUBBYTES[2].a/w500 ,
         \SUBBYTES[2].a/w499 , \SUBBYTES[2].a/w498 , \SUBBYTES[2].a/w495 ,
         \SUBBYTES[2].a/w493 , \SUBBYTES[2].a/w492 , \SUBBYTES[2].a/w491 ,
         \SUBBYTES[2].a/w487 , \SUBBYTES[2].a/w485 , \SUBBYTES[2].a/w484 ,
         \SUBBYTES[2].a/w483 , \SUBBYTES[2].a/w482 , \SUBBYTES[2].a/w481 ,
         \SUBBYTES[2].a/w480 , \SUBBYTES[2].a/w479 , \SUBBYTES[2].a/w478 ,
         \SUBBYTES[2].a/w470 , \SUBBYTES[2].a/w468 , \SUBBYTES[2].a/w467 ,
         \SUBBYTES[2].a/w463 , \SUBBYTES[2].a/w461 , \SUBBYTES[2].a/w460 ,
         \SUBBYTES[2].a/w459 , \SUBBYTES[2].a/w455 , \SUBBYTES[2].a/w453 ,
         \SUBBYTES[2].a/w452 , \SUBBYTES[2].a/w439 , \SUBBYTES[2].a/w438 ,
         \SUBBYTES[2].a/w437 , \SUBBYTES[2].a/w435 , \SUBBYTES[2].a/w432 ,
         \SUBBYTES[2].a/w431 , \SUBBYTES[2].a/w429 , \SUBBYTES[2].a/w428 ,
         \SUBBYTES[2].a/w426 , \SUBBYTES[2].a/w424 , \SUBBYTES[2].a/w423 ,
         \SUBBYTES[2].a/w417 , \SUBBYTES[2].a/w416 , \SUBBYTES[2].a/w415 ,
         \SUBBYTES[2].a/w414 , \SUBBYTES[2].a/w408 , \SUBBYTES[2].a/w406 ,
         \SUBBYTES[2].a/w405 , \SUBBYTES[2].a/w401 , \SUBBYTES[2].a/w399 ,
         \SUBBYTES[2].a/w398 , \SUBBYTES[2].a/w393 , \SUBBYTES[2].a/w391 ,
         \SUBBYTES[2].a/w390 , \SUBBYTES[2].a/w374 , \SUBBYTES[2].a/w373 ,
         \SUBBYTES[2].a/w372 , \SUBBYTES[2].a/w371 , \SUBBYTES[2].a/w370 ,
         \SUBBYTES[2].a/w368 , \SUBBYTES[2].a/w367 , \SUBBYTES[2].a/w295 ,
         \SUBBYTES[2].a/w293 , \SUBBYTES[2].a/w292 , \SUBBYTES[2].a/w291 ,
         \SUBBYTES[2].a/w288 , \SUBBYTES[2].a/w286 , \SUBBYTES[2].a/w285 ,
         \SUBBYTES[2].a/w284 , \SUBBYTES[2].a/w280 , \SUBBYTES[2].a/w278 ,
         \SUBBYTES[2].a/w277 , \SUBBYTES[2].a/w276 , \SUBBYTES[2].a/w275 ,
         \SUBBYTES[2].a/w274 , \SUBBYTES[2].a/w273 , \SUBBYTES[2].a/w272 ,
         \SUBBYTES[2].a/w271 , \SUBBYTES[2].a/w263 , \SUBBYTES[2].a/w261 ,
         \SUBBYTES[2].a/w260 , \SUBBYTES[2].a/w256 , \SUBBYTES[2].a/w254 ,
         \SUBBYTES[2].a/w253 , \SUBBYTES[2].a/w252 , \SUBBYTES[2].a/w248 ,
         \SUBBYTES[2].a/w246 , \SUBBYTES[2].a/w245 , \SUBBYTES[2].a/w232 ,
         \SUBBYTES[2].a/w231 , \SUBBYTES[2].a/w230 , \SUBBYTES[2].a/w228 ,
         \SUBBYTES[2].a/w225 , \SUBBYTES[2].a/w224 , \SUBBYTES[2].a/w222 ,
         \SUBBYTES[2].a/w221 , \SUBBYTES[2].a/w219 , \SUBBYTES[2].a/w217 ,
         \SUBBYTES[2].a/w216 , \SUBBYTES[2].a/w210 , \SUBBYTES[2].a/w209 ,
         \SUBBYTES[2].a/w208 , \SUBBYTES[2].a/w207 , \SUBBYTES[2].a/w201 ,
         \SUBBYTES[2].a/w199 , \SUBBYTES[2].a/w198 , \SUBBYTES[2].a/w194 ,
         \SUBBYTES[2].a/w192 , \SUBBYTES[2].a/w191 , \SUBBYTES[2].a/w186 ,
         \SUBBYTES[2].a/w184 , \SUBBYTES[2].a/w183 , \SUBBYTES[2].a/w167 ,
         \SUBBYTES[2].a/w166 , \SUBBYTES[2].a/w165 , \SUBBYTES[2].a/w164 ,
         \SUBBYTES[2].a/w163 , \SUBBYTES[2].a/w161 , \SUBBYTES[2].a/w160 ,
         \SUBBYTES[1].a/w3400 , \SUBBYTES[1].a/w3398 , \SUBBYTES[1].a/w3397 ,
         \SUBBYTES[1].a/w3396 , \SUBBYTES[1].a/w3393 , \SUBBYTES[1].a/w3391 ,
         \SUBBYTES[1].a/w3390 , \SUBBYTES[1].a/w3389 , \SUBBYTES[1].a/w3385 ,
         \SUBBYTES[1].a/w3383 , \SUBBYTES[1].a/w3382 , \SUBBYTES[1].a/w3381 ,
         \SUBBYTES[1].a/w3380 , \SUBBYTES[1].a/w3379 , \SUBBYTES[1].a/w3378 ,
         \SUBBYTES[1].a/w3377 , \SUBBYTES[1].a/w3376 , \SUBBYTES[1].a/w3368 ,
         \SUBBYTES[1].a/w3366 , \SUBBYTES[1].a/w3365 , \SUBBYTES[1].a/w3361 ,
         \SUBBYTES[1].a/w3359 , \SUBBYTES[1].a/w3358 , \SUBBYTES[1].a/w3357 ,
         \SUBBYTES[1].a/w3353 , \SUBBYTES[1].a/w3351 , \SUBBYTES[1].a/w3350 ,
         \SUBBYTES[1].a/w3337 , \SUBBYTES[1].a/w3336 , \SUBBYTES[1].a/w3335 ,
         \SUBBYTES[1].a/w3333 , \SUBBYTES[1].a/w3330 , \SUBBYTES[1].a/w3329 ,
         \SUBBYTES[1].a/w3327 , \SUBBYTES[1].a/w3326 , \SUBBYTES[1].a/w3324 ,
         \SUBBYTES[1].a/w3322 , \SUBBYTES[1].a/w3321 , \SUBBYTES[1].a/w3315 ,
         \SUBBYTES[1].a/w3314 , \SUBBYTES[1].a/w3313 , \SUBBYTES[1].a/w3312 ,
         \SUBBYTES[1].a/w3306 , \SUBBYTES[1].a/w3304 , \SUBBYTES[1].a/w3303 ,
         \SUBBYTES[1].a/w3299 , \SUBBYTES[1].a/w3297 , \SUBBYTES[1].a/w3296 ,
         \SUBBYTES[1].a/w3291 , \SUBBYTES[1].a/w3289 , \SUBBYTES[1].a/w3288 ,
         \SUBBYTES[1].a/w3272 , \SUBBYTES[1].a/w3271 , \SUBBYTES[1].a/w3270 ,
         \SUBBYTES[1].a/w3269 , \SUBBYTES[1].a/w3268 , \SUBBYTES[1].a/w3266 ,
         \SUBBYTES[1].a/w3265 , \SUBBYTES[1].a/w3193 , \SUBBYTES[1].a/w3191 ,
         \SUBBYTES[1].a/w3190 , \SUBBYTES[1].a/w3189 , \SUBBYTES[1].a/w3186 ,
         \SUBBYTES[1].a/w3184 , \SUBBYTES[1].a/w3183 , \SUBBYTES[1].a/w3182 ,
         \SUBBYTES[1].a/w3178 , \SUBBYTES[1].a/w3176 , \SUBBYTES[1].a/w3175 ,
         \SUBBYTES[1].a/w3174 , \SUBBYTES[1].a/w3173 , \SUBBYTES[1].a/w3172 ,
         \SUBBYTES[1].a/w3171 , \SUBBYTES[1].a/w3170 , \SUBBYTES[1].a/w3169 ,
         \SUBBYTES[1].a/w3161 , \SUBBYTES[1].a/w3159 , \SUBBYTES[1].a/w3158 ,
         \SUBBYTES[1].a/w3154 , \SUBBYTES[1].a/w3152 , \SUBBYTES[1].a/w3151 ,
         \SUBBYTES[1].a/w3150 , \SUBBYTES[1].a/w3146 , \SUBBYTES[1].a/w3144 ,
         \SUBBYTES[1].a/w3143 , \SUBBYTES[1].a/w3130 , \SUBBYTES[1].a/w3129 ,
         \SUBBYTES[1].a/w3128 , \SUBBYTES[1].a/w3126 , \SUBBYTES[1].a/w3123 ,
         \SUBBYTES[1].a/w3122 , \SUBBYTES[1].a/w3120 , \SUBBYTES[1].a/w3119 ,
         \SUBBYTES[1].a/w3117 , \SUBBYTES[1].a/w3115 , \SUBBYTES[1].a/w3114 ,
         \SUBBYTES[1].a/w3108 , \SUBBYTES[1].a/w3107 , \SUBBYTES[1].a/w3106 ,
         \SUBBYTES[1].a/w3105 , \SUBBYTES[1].a/w3099 , \SUBBYTES[1].a/w3097 ,
         \SUBBYTES[1].a/w3096 , \SUBBYTES[1].a/w3092 , \SUBBYTES[1].a/w3090 ,
         \SUBBYTES[1].a/w3089 , \SUBBYTES[1].a/w3084 , \SUBBYTES[1].a/w3082 ,
         \SUBBYTES[1].a/w3081 , \SUBBYTES[1].a/w3065 , \SUBBYTES[1].a/w3064 ,
         \SUBBYTES[1].a/w3063 , \SUBBYTES[1].a/w3062 , \SUBBYTES[1].a/w3061 ,
         \SUBBYTES[1].a/w3059 , \SUBBYTES[1].a/w3058 , \SUBBYTES[1].a/w2986 ,
         \SUBBYTES[1].a/w2984 , \SUBBYTES[1].a/w2983 , \SUBBYTES[1].a/w2982 ,
         \SUBBYTES[1].a/w2979 , \SUBBYTES[1].a/w2977 , \SUBBYTES[1].a/w2976 ,
         \SUBBYTES[1].a/w2975 , \SUBBYTES[1].a/w2971 , \SUBBYTES[1].a/w2969 ,
         \SUBBYTES[1].a/w2968 , \SUBBYTES[1].a/w2967 , \SUBBYTES[1].a/w2966 ,
         \SUBBYTES[1].a/w2965 , \SUBBYTES[1].a/w2964 , \SUBBYTES[1].a/w2963 ,
         \SUBBYTES[1].a/w2962 , \SUBBYTES[1].a/w2954 , \SUBBYTES[1].a/w2952 ,
         \SUBBYTES[1].a/w2951 , \SUBBYTES[1].a/w2947 , \SUBBYTES[1].a/w2945 ,
         \SUBBYTES[1].a/w2944 , \SUBBYTES[1].a/w2943 , \SUBBYTES[1].a/w2939 ,
         \SUBBYTES[1].a/w2937 , \SUBBYTES[1].a/w2936 , \SUBBYTES[1].a/w2923 ,
         \SUBBYTES[1].a/w2922 , \SUBBYTES[1].a/w2921 , \SUBBYTES[1].a/w2919 ,
         \SUBBYTES[1].a/w2916 , \SUBBYTES[1].a/w2915 , \SUBBYTES[1].a/w2913 ,
         \SUBBYTES[1].a/w2912 , \SUBBYTES[1].a/w2910 , \SUBBYTES[1].a/w2908 ,
         \SUBBYTES[1].a/w2907 , \SUBBYTES[1].a/w2901 , \SUBBYTES[1].a/w2900 ,
         \SUBBYTES[1].a/w2899 , \SUBBYTES[1].a/w2898 , \SUBBYTES[1].a/w2892 ,
         \SUBBYTES[1].a/w2890 , \SUBBYTES[1].a/w2889 , \SUBBYTES[1].a/w2885 ,
         \SUBBYTES[1].a/w2883 , \SUBBYTES[1].a/w2882 , \SUBBYTES[1].a/w2877 ,
         \SUBBYTES[1].a/w2875 , \SUBBYTES[1].a/w2874 , \SUBBYTES[1].a/w2858 ,
         \SUBBYTES[1].a/w2857 , \SUBBYTES[1].a/w2856 , \SUBBYTES[1].a/w2855 ,
         \SUBBYTES[1].a/w2854 , \SUBBYTES[1].a/w2852 , \SUBBYTES[1].a/w2851 ,
         \SUBBYTES[1].a/w2779 , \SUBBYTES[1].a/w2777 , \SUBBYTES[1].a/w2776 ,
         \SUBBYTES[1].a/w2775 , \SUBBYTES[1].a/w2772 , \SUBBYTES[1].a/w2770 ,
         \SUBBYTES[1].a/w2769 , \SUBBYTES[1].a/w2768 , \SUBBYTES[1].a/w2764 ,
         \SUBBYTES[1].a/w2762 , \SUBBYTES[1].a/w2761 , \SUBBYTES[1].a/w2760 ,
         \SUBBYTES[1].a/w2759 , \SUBBYTES[1].a/w2758 , \SUBBYTES[1].a/w2757 ,
         \SUBBYTES[1].a/w2756 , \SUBBYTES[1].a/w2755 , \SUBBYTES[1].a/w2747 ,
         \SUBBYTES[1].a/w2745 , \SUBBYTES[1].a/w2744 , \SUBBYTES[1].a/w2740 ,
         \SUBBYTES[1].a/w2738 , \SUBBYTES[1].a/w2737 , \SUBBYTES[1].a/w2736 ,
         \SUBBYTES[1].a/w2732 , \SUBBYTES[1].a/w2730 , \SUBBYTES[1].a/w2729 ,
         \SUBBYTES[1].a/w2716 , \SUBBYTES[1].a/w2715 , \SUBBYTES[1].a/w2714 ,
         \SUBBYTES[1].a/w2712 , \SUBBYTES[1].a/w2709 , \SUBBYTES[1].a/w2708 ,
         \SUBBYTES[1].a/w2706 , \SUBBYTES[1].a/w2705 , \SUBBYTES[1].a/w2703 ,
         \SUBBYTES[1].a/w2701 , \SUBBYTES[1].a/w2700 , \SUBBYTES[1].a/w2694 ,
         \SUBBYTES[1].a/w2693 , \SUBBYTES[1].a/w2692 , \SUBBYTES[1].a/w2691 ,
         \SUBBYTES[1].a/w2685 , \SUBBYTES[1].a/w2683 , \SUBBYTES[1].a/w2682 ,
         \SUBBYTES[1].a/w2678 , \SUBBYTES[1].a/w2676 , \SUBBYTES[1].a/w2675 ,
         \SUBBYTES[1].a/w2670 , \SUBBYTES[1].a/w2668 , \SUBBYTES[1].a/w2667 ,
         \SUBBYTES[1].a/w2651 , \SUBBYTES[1].a/w2650 , \SUBBYTES[1].a/w2649 ,
         \SUBBYTES[1].a/w2648 , \SUBBYTES[1].a/w2647 , \SUBBYTES[1].a/w2645 ,
         \SUBBYTES[1].a/w2644 , \SUBBYTES[1].a/w2572 , \SUBBYTES[1].a/w2570 ,
         \SUBBYTES[1].a/w2569 , \SUBBYTES[1].a/w2568 , \SUBBYTES[1].a/w2565 ,
         \SUBBYTES[1].a/w2563 , \SUBBYTES[1].a/w2562 , \SUBBYTES[1].a/w2561 ,
         \SUBBYTES[1].a/w2557 , \SUBBYTES[1].a/w2555 , \SUBBYTES[1].a/w2554 ,
         \SUBBYTES[1].a/w2553 , \SUBBYTES[1].a/w2552 , \SUBBYTES[1].a/w2551 ,
         \SUBBYTES[1].a/w2550 , \SUBBYTES[1].a/w2549 , \SUBBYTES[1].a/w2548 ,
         \SUBBYTES[1].a/w2540 , \SUBBYTES[1].a/w2538 , \SUBBYTES[1].a/w2537 ,
         \SUBBYTES[1].a/w2533 , \SUBBYTES[1].a/w2531 , \SUBBYTES[1].a/w2530 ,
         \SUBBYTES[1].a/w2529 , \SUBBYTES[1].a/w2525 , \SUBBYTES[1].a/w2523 ,
         \SUBBYTES[1].a/w2522 , \SUBBYTES[1].a/w2509 , \SUBBYTES[1].a/w2508 ,
         \SUBBYTES[1].a/w2507 , \SUBBYTES[1].a/w2505 , \SUBBYTES[1].a/w2502 ,
         \SUBBYTES[1].a/w2501 , \SUBBYTES[1].a/w2499 , \SUBBYTES[1].a/w2498 ,
         \SUBBYTES[1].a/w2496 , \SUBBYTES[1].a/w2494 , \SUBBYTES[1].a/w2493 ,
         \SUBBYTES[1].a/w2487 , \SUBBYTES[1].a/w2486 , \SUBBYTES[1].a/w2485 ,
         \SUBBYTES[1].a/w2484 , \SUBBYTES[1].a/w2478 , \SUBBYTES[1].a/w2476 ,
         \SUBBYTES[1].a/w2475 , \SUBBYTES[1].a/w2471 , \SUBBYTES[1].a/w2469 ,
         \SUBBYTES[1].a/w2468 , \SUBBYTES[1].a/w2463 , \SUBBYTES[1].a/w2461 ,
         \SUBBYTES[1].a/w2460 , \SUBBYTES[1].a/w2444 , \SUBBYTES[1].a/w2443 ,
         \SUBBYTES[1].a/w2442 , \SUBBYTES[1].a/w2441 , \SUBBYTES[1].a/w2440 ,
         \SUBBYTES[1].a/w2438 , \SUBBYTES[1].a/w2437 , \SUBBYTES[1].a/w2365 ,
         \SUBBYTES[1].a/w2363 , \SUBBYTES[1].a/w2362 , \SUBBYTES[1].a/w2361 ,
         \SUBBYTES[1].a/w2358 , \SUBBYTES[1].a/w2356 , \SUBBYTES[1].a/w2355 ,
         \SUBBYTES[1].a/w2354 , \SUBBYTES[1].a/w2350 , \SUBBYTES[1].a/w2348 ,
         \SUBBYTES[1].a/w2347 , \SUBBYTES[1].a/w2346 , \SUBBYTES[1].a/w2345 ,
         \SUBBYTES[1].a/w2344 , \SUBBYTES[1].a/w2343 , \SUBBYTES[1].a/w2342 ,
         \SUBBYTES[1].a/w2341 , \SUBBYTES[1].a/w2333 , \SUBBYTES[1].a/w2331 ,
         \SUBBYTES[1].a/w2330 , \SUBBYTES[1].a/w2326 , \SUBBYTES[1].a/w2324 ,
         \SUBBYTES[1].a/w2323 , \SUBBYTES[1].a/w2322 , \SUBBYTES[1].a/w2318 ,
         \SUBBYTES[1].a/w2316 , \SUBBYTES[1].a/w2315 , \SUBBYTES[1].a/w2302 ,
         \SUBBYTES[1].a/w2301 , \SUBBYTES[1].a/w2300 , \SUBBYTES[1].a/w2298 ,
         \SUBBYTES[1].a/w2295 , \SUBBYTES[1].a/w2294 , \SUBBYTES[1].a/w2292 ,
         \SUBBYTES[1].a/w2291 , \SUBBYTES[1].a/w2289 , \SUBBYTES[1].a/w2287 ,
         \SUBBYTES[1].a/w2286 , \SUBBYTES[1].a/w2280 , \SUBBYTES[1].a/w2279 ,
         \SUBBYTES[1].a/w2278 , \SUBBYTES[1].a/w2277 , \SUBBYTES[1].a/w2271 ,
         \SUBBYTES[1].a/w2269 , \SUBBYTES[1].a/w2268 , \SUBBYTES[1].a/w2264 ,
         \SUBBYTES[1].a/w2262 , \SUBBYTES[1].a/w2261 , \SUBBYTES[1].a/w2256 ,
         \SUBBYTES[1].a/w2254 , \SUBBYTES[1].a/w2253 , \SUBBYTES[1].a/w2237 ,
         \SUBBYTES[1].a/w2236 , \SUBBYTES[1].a/w2235 , \SUBBYTES[1].a/w2234 ,
         \SUBBYTES[1].a/w2233 , \SUBBYTES[1].a/w2231 , \SUBBYTES[1].a/w2230 ,
         \SUBBYTES[1].a/w2158 , \SUBBYTES[1].a/w2156 , \SUBBYTES[1].a/w2155 ,
         \SUBBYTES[1].a/w2154 , \SUBBYTES[1].a/w2151 , \SUBBYTES[1].a/w2149 ,
         \SUBBYTES[1].a/w2148 , \SUBBYTES[1].a/w2147 , \SUBBYTES[1].a/w2143 ,
         \SUBBYTES[1].a/w2141 , \SUBBYTES[1].a/w2140 , \SUBBYTES[1].a/w2139 ,
         \SUBBYTES[1].a/w2138 , \SUBBYTES[1].a/w2137 , \SUBBYTES[1].a/w2136 ,
         \SUBBYTES[1].a/w2135 , \SUBBYTES[1].a/w2134 , \SUBBYTES[1].a/w2126 ,
         \SUBBYTES[1].a/w2124 , \SUBBYTES[1].a/w2123 , \SUBBYTES[1].a/w2119 ,
         \SUBBYTES[1].a/w2117 , \SUBBYTES[1].a/w2116 , \SUBBYTES[1].a/w2115 ,
         \SUBBYTES[1].a/w2111 , \SUBBYTES[1].a/w2109 , \SUBBYTES[1].a/w2108 ,
         \SUBBYTES[1].a/w2095 , \SUBBYTES[1].a/w2094 , \SUBBYTES[1].a/w2093 ,
         \SUBBYTES[1].a/w2091 , \SUBBYTES[1].a/w2088 , \SUBBYTES[1].a/w2087 ,
         \SUBBYTES[1].a/w2085 , \SUBBYTES[1].a/w2084 , \SUBBYTES[1].a/w2082 ,
         \SUBBYTES[1].a/w2080 , \SUBBYTES[1].a/w2079 , \SUBBYTES[1].a/w2073 ,
         \SUBBYTES[1].a/w2072 , \SUBBYTES[1].a/w2071 , \SUBBYTES[1].a/w2070 ,
         \SUBBYTES[1].a/w2064 , \SUBBYTES[1].a/w2062 , \SUBBYTES[1].a/w2061 ,
         \SUBBYTES[1].a/w2057 , \SUBBYTES[1].a/w2055 , \SUBBYTES[1].a/w2054 ,
         \SUBBYTES[1].a/w2049 , \SUBBYTES[1].a/w2047 , \SUBBYTES[1].a/w2046 ,
         \SUBBYTES[1].a/w2030 , \SUBBYTES[1].a/w2029 , \SUBBYTES[1].a/w2028 ,
         \SUBBYTES[1].a/w2027 , \SUBBYTES[1].a/w2026 , \SUBBYTES[1].a/w2024 ,
         \SUBBYTES[1].a/w2023 , \SUBBYTES[1].a/w1951 , \SUBBYTES[1].a/w1949 ,
         \SUBBYTES[1].a/w1948 , \SUBBYTES[1].a/w1947 , \SUBBYTES[1].a/w1944 ,
         \SUBBYTES[1].a/w1942 , \SUBBYTES[1].a/w1941 , \SUBBYTES[1].a/w1940 ,
         \SUBBYTES[1].a/w1936 , \SUBBYTES[1].a/w1934 , \SUBBYTES[1].a/w1933 ,
         \SUBBYTES[1].a/w1932 , \SUBBYTES[1].a/w1931 , \SUBBYTES[1].a/w1930 ,
         \SUBBYTES[1].a/w1929 , \SUBBYTES[1].a/w1928 , \SUBBYTES[1].a/w1927 ,
         \SUBBYTES[1].a/w1919 , \SUBBYTES[1].a/w1917 , \SUBBYTES[1].a/w1916 ,
         \SUBBYTES[1].a/w1912 , \SUBBYTES[1].a/w1910 , \SUBBYTES[1].a/w1909 ,
         \SUBBYTES[1].a/w1908 , \SUBBYTES[1].a/w1904 , \SUBBYTES[1].a/w1902 ,
         \SUBBYTES[1].a/w1901 , \SUBBYTES[1].a/w1888 , \SUBBYTES[1].a/w1887 ,
         \SUBBYTES[1].a/w1886 , \SUBBYTES[1].a/w1884 , \SUBBYTES[1].a/w1881 ,
         \SUBBYTES[1].a/w1880 , \SUBBYTES[1].a/w1878 , \SUBBYTES[1].a/w1877 ,
         \SUBBYTES[1].a/w1875 , \SUBBYTES[1].a/w1873 , \SUBBYTES[1].a/w1872 ,
         \SUBBYTES[1].a/w1866 , \SUBBYTES[1].a/w1865 , \SUBBYTES[1].a/w1864 ,
         \SUBBYTES[1].a/w1863 , \SUBBYTES[1].a/w1857 , \SUBBYTES[1].a/w1855 ,
         \SUBBYTES[1].a/w1854 , \SUBBYTES[1].a/w1850 , \SUBBYTES[1].a/w1848 ,
         \SUBBYTES[1].a/w1847 , \SUBBYTES[1].a/w1842 , \SUBBYTES[1].a/w1840 ,
         \SUBBYTES[1].a/w1839 , \SUBBYTES[1].a/w1823 , \SUBBYTES[1].a/w1822 ,
         \SUBBYTES[1].a/w1821 , \SUBBYTES[1].a/w1820 , \SUBBYTES[1].a/w1819 ,
         \SUBBYTES[1].a/w1817 , \SUBBYTES[1].a/w1816 , \SUBBYTES[1].a/w1744 ,
         \SUBBYTES[1].a/w1742 , \SUBBYTES[1].a/w1741 , \SUBBYTES[1].a/w1740 ,
         \SUBBYTES[1].a/w1737 , \SUBBYTES[1].a/w1735 , \SUBBYTES[1].a/w1734 ,
         \SUBBYTES[1].a/w1733 , \SUBBYTES[1].a/w1729 , \SUBBYTES[1].a/w1727 ,
         \SUBBYTES[1].a/w1726 , \SUBBYTES[1].a/w1725 , \SUBBYTES[1].a/w1724 ,
         \SUBBYTES[1].a/w1723 , \SUBBYTES[1].a/w1722 , \SUBBYTES[1].a/w1721 ,
         \SUBBYTES[1].a/w1720 , \SUBBYTES[1].a/w1712 , \SUBBYTES[1].a/w1710 ,
         \SUBBYTES[1].a/w1709 , \SUBBYTES[1].a/w1705 , \SUBBYTES[1].a/w1703 ,
         \SUBBYTES[1].a/w1702 , \SUBBYTES[1].a/w1701 , \SUBBYTES[1].a/w1697 ,
         \SUBBYTES[1].a/w1695 , \SUBBYTES[1].a/w1694 , \SUBBYTES[1].a/w1681 ,
         \SUBBYTES[1].a/w1680 , \SUBBYTES[1].a/w1679 , \SUBBYTES[1].a/w1677 ,
         \SUBBYTES[1].a/w1674 , \SUBBYTES[1].a/w1673 , \SUBBYTES[1].a/w1671 ,
         \SUBBYTES[1].a/w1670 , \SUBBYTES[1].a/w1668 , \SUBBYTES[1].a/w1666 ,
         \SUBBYTES[1].a/w1665 , \SUBBYTES[1].a/w1659 , \SUBBYTES[1].a/w1658 ,
         \SUBBYTES[1].a/w1657 , \SUBBYTES[1].a/w1656 , \SUBBYTES[1].a/w1650 ,
         \SUBBYTES[1].a/w1648 , \SUBBYTES[1].a/w1647 , \SUBBYTES[1].a/w1643 ,
         \SUBBYTES[1].a/w1641 , \SUBBYTES[1].a/w1640 , \SUBBYTES[1].a/w1635 ,
         \SUBBYTES[1].a/w1633 , \SUBBYTES[1].a/w1632 , \SUBBYTES[1].a/w1616 ,
         \SUBBYTES[1].a/w1615 , \SUBBYTES[1].a/w1614 , \SUBBYTES[1].a/w1613 ,
         \SUBBYTES[1].a/w1612 , \SUBBYTES[1].a/w1610 , \SUBBYTES[1].a/w1609 ,
         \SUBBYTES[1].a/w1537 , \SUBBYTES[1].a/w1535 , \SUBBYTES[1].a/w1534 ,
         \SUBBYTES[1].a/w1533 , \SUBBYTES[1].a/w1530 , \SUBBYTES[1].a/w1528 ,
         \SUBBYTES[1].a/w1527 , \SUBBYTES[1].a/w1526 , \SUBBYTES[1].a/w1522 ,
         \SUBBYTES[1].a/w1520 , \SUBBYTES[1].a/w1519 , \SUBBYTES[1].a/w1518 ,
         \SUBBYTES[1].a/w1517 , \SUBBYTES[1].a/w1516 , \SUBBYTES[1].a/w1515 ,
         \SUBBYTES[1].a/w1514 , \SUBBYTES[1].a/w1513 , \SUBBYTES[1].a/w1505 ,
         \SUBBYTES[1].a/w1503 , \SUBBYTES[1].a/w1502 , \SUBBYTES[1].a/w1498 ,
         \SUBBYTES[1].a/w1496 , \SUBBYTES[1].a/w1495 , \SUBBYTES[1].a/w1494 ,
         \SUBBYTES[1].a/w1490 , \SUBBYTES[1].a/w1488 , \SUBBYTES[1].a/w1487 ,
         \SUBBYTES[1].a/w1474 , \SUBBYTES[1].a/w1473 , \SUBBYTES[1].a/w1472 ,
         \SUBBYTES[1].a/w1470 , \SUBBYTES[1].a/w1467 , \SUBBYTES[1].a/w1466 ,
         \SUBBYTES[1].a/w1464 , \SUBBYTES[1].a/w1463 , \SUBBYTES[1].a/w1461 ,
         \SUBBYTES[1].a/w1459 , \SUBBYTES[1].a/w1458 , \SUBBYTES[1].a/w1452 ,
         \SUBBYTES[1].a/w1451 , \SUBBYTES[1].a/w1450 , \SUBBYTES[1].a/w1449 ,
         \SUBBYTES[1].a/w1443 , \SUBBYTES[1].a/w1441 , \SUBBYTES[1].a/w1440 ,
         \SUBBYTES[1].a/w1436 , \SUBBYTES[1].a/w1434 , \SUBBYTES[1].a/w1433 ,
         \SUBBYTES[1].a/w1428 , \SUBBYTES[1].a/w1426 , \SUBBYTES[1].a/w1425 ,
         \SUBBYTES[1].a/w1409 , \SUBBYTES[1].a/w1408 , \SUBBYTES[1].a/w1407 ,
         \SUBBYTES[1].a/w1406 , \SUBBYTES[1].a/w1405 , \SUBBYTES[1].a/w1403 ,
         \SUBBYTES[1].a/w1402 , \SUBBYTES[1].a/w1330 , \SUBBYTES[1].a/w1328 ,
         \SUBBYTES[1].a/w1327 , \SUBBYTES[1].a/w1326 , \SUBBYTES[1].a/w1323 ,
         \SUBBYTES[1].a/w1321 , \SUBBYTES[1].a/w1320 , \SUBBYTES[1].a/w1319 ,
         \SUBBYTES[1].a/w1315 , \SUBBYTES[1].a/w1313 , \SUBBYTES[1].a/w1312 ,
         \SUBBYTES[1].a/w1311 , \SUBBYTES[1].a/w1310 , \SUBBYTES[1].a/w1309 ,
         \SUBBYTES[1].a/w1308 , \SUBBYTES[1].a/w1307 , \SUBBYTES[1].a/w1306 ,
         \SUBBYTES[1].a/w1298 , \SUBBYTES[1].a/w1296 , \SUBBYTES[1].a/w1295 ,
         \SUBBYTES[1].a/w1291 , \SUBBYTES[1].a/w1289 , \SUBBYTES[1].a/w1288 ,
         \SUBBYTES[1].a/w1287 , \SUBBYTES[1].a/w1283 , \SUBBYTES[1].a/w1281 ,
         \SUBBYTES[1].a/w1280 , \SUBBYTES[1].a/w1267 , \SUBBYTES[1].a/w1266 ,
         \SUBBYTES[1].a/w1265 , \SUBBYTES[1].a/w1263 , \SUBBYTES[1].a/w1260 ,
         \SUBBYTES[1].a/w1259 , \SUBBYTES[1].a/w1257 , \SUBBYTES[1].a/w1256 ,
         \SUBBYTES[1].a/w1254 , \SUBBYTES[1].a/w1252 , \SUBBYTES[1].a/w1251 ,
         \SUBBYTES[1].a/w1245 , \SUBBYTES[1].a/w1244 , \SUBBYTES[1].a/w1243 ,
         \SUBBYTES[1].a/w1242 , \SUBBYTES[1].a/w1236 , \SUBBYTES[1].a/w1234 ,
         \SUBBYTES[1].a/w1233 , \SUBBYTES[1].a/w1229 , \SUBBYTES[1].a/w1227 ,
         \SUBBYTES[1].a/w1226 , \SUBBYTES[1].a/w1221 , \SUBBYTES[1].a/w1219 ,
         \SUBBYTES[1].a/w1218 , \SUBBYTES[1].a/w1202 , \SUBBYTES[1].a/w1201 ,
         \SUBBYTES[1].a/w1200 , \SUBBYTES[1].a/w1199 , \SUBBYTES[1].a/w1198 ,
         \SUBBYTES[1].a/w1196 , \SUBBYTES[1].a/w1195 , \SUBBYTES[1].a/w1123 ,
         \SUBBYTES[1].a/w1121 , \SUBBYTES[1].a/w1120 , \SUBBYTES[1].a/w1119 ,
         \SUBBYTES[1].a/w1116 , \SUBBYTES[1].a/w1114 , \SUBBYTES[1].a/w1113 ,
         \SUBBYTES[1].a/w1112 , \SUBBYTES[1].a/w1108 , \SUBBYTES[1].a/w1106 ,
         \SUBBYTES[1].a/w1105 , \SUBBYTES[1].a/w1104 , \SUBBYTES[1].a/w1103 ,
         \SUBBYTES[1].a/w1102 , \SUBBYTES[1].a/w1101 , \SUBBYTES[1].a/w1100 ,
         \SUBBYTES[1].a/w1099 , \SUBBYTES[1].a/w1091 , \SUBBYTES[1].a/w1089 ,
         \SUBBYTES[1].a/w1088 , \SUBBYTES[1].a/w1084 , \SUBBYTES[1].a/w1082 ,
         \SUBBYTES[1].a/w1081 , \SUBBYTES[1].a/w1080 , \SUBBYTES[1].a/w1076 ,
         \SUBBYTES[1].a/w1074 , \SUBBYTES[1].a/w1073 , \SUBBYTES[1].a/w1060 ,
         \SUBBYTES[1].a/w1059 , \SUBBYTES[1].a/w1058 , \SUBBYTES[1].a/w1056 ,
         \SUBBYTES[1].a/w1053 , \SUBBYTES[1].a/w1052 , \SUBBYTES[1].a/w1050 ,
         \SUBBYTES[1].a/w1049 , \SUBBYTES[1].a/w1047 , \SUBBYTES[1].a/w1045 ,
         \SUBBYTES[1].a/w1044 , \SUBBYTES[1].a/w1038 , \SUBBYTES[1].a/w1037 ,
         \SUBBYTES[1].a/w1036 , \SUBBYTES[1].a/w1035 , \SUBBYTES[1].a/w1029 ,
         \SUBBYTES[1].a/w1027 , \SUBBYTES[1].a/w1026 , \SUBBYTES[1].a/w1022 ,
         \SUBBYTES[1].a/w1020 , \SUBBYTES[1].a/w1019 , \SUBBYTES[1].a/w1014 ,
         \SUBBYTES[1].a/w1012 , \SUBBYTES[1].a/w1011 , \SUBBYTES[1].a/w995 ,
         \SUBBYTES[1].a/w994 , \SUBBYTES[1].a/w993 , \SUBBYTES[1].a/w992 ,
         \SUBBYTES[1].a/w991 , \SUBBYTES[1].a/w989 , \SUBBYTES[1].a/w988 ,
         \SUBBYTES[1].a/w916 , \SUBBYTES[1].a/w914 , \SUBBYTES[1].a/w913 ,
         \SUBBYTES[1].a/w912 , \SUBBYTES[1].a/w909 , \SUBBYTES[1].a/w907 ,
         \SUBBYTES[1].a/w906 , \SUBBYTES[1].a/w905 , \SUBBYTES[1].a/w901 ,
         \SUBBYTES[1].a/w899 , \SUBBYTES[1].a/w898 , \SUBBYTES[1].a/w897 ,
         \SUBBYTES[1].a/w896 , \SUBBYTES[1].a/w895 , \SUBBYTES[1].a/w894 ,
         \SUBBYTES[1].a/w893 , \SUBBYTES[1].a/w892 , \SUBBYTES[1].a/w884 ,
         \SUBBYTES[1].a/w882 , \SUBBYTES[1].a/w881 , \SUBBYTES[1].a/w877 ,
         \SUBBYTES[1].a/w875 , \SUBBYTES[1].a/w874 , \SUBBYTES[1].a/w873 ,
         \SUBBYTES[1].a/w869 , \SUBBYTES[1].a/w867 , \SUBBYTES[1].a/w866 ,
         \SUBBYTES[1].a/w853 , \SUBBYTES[1].a/w852 , \SUBBYTES[1].a/w851 ,
         \SUBBYTES[1].a/w849 , \SUBBYTES[1].a/w846 , \SUBBYTES[1].a/w845 ,
         \SUBBYTES[1].a/w843 , \SUBBYTES[1].a/w842 , \SUBBYTES[1].a/w840 ,
         \SUBBYTES[1].a/w838 , \SUBBYTES[1].a/w837 , \SUBBYTES[1].a/w831 ,
         \SUBBYTES[1].a/w830 , \SUBBYTES[1].a/w829 , \SUBBYTES[1].a/w828 ,
         \SUBBYTES[1].a/w822 , \SUBBYTES[1].a/w820 , \SUBBYTES[1].a/w819 ,
         \SUBBYTES[1].a/w815 , \SUBBYTES[1].a/w813 , \SUBBYTES[1].a/w812 ,
         \SUBBYTES[1].a/w807 , \SUBBYTES[1].a/w805 , \SUBBYTES[1].a/w804 ,
         \SUBBYTES[1].a/w788 , \SUBBYTES[1].a/w787 , \SUBBYTES[1].a/w786 ,
         \SUBBYTES[1].a/w785 , \SUBBYTES[1].a/w784 , \SUBBYTES[1].a/w782 ,
         \SUBBYTES[1].a/w781 , \SUBBYTES[1].a/w709 , \SUBBYTES[1].a/w707 ,
         \SUBBYTES[1].a/w706 , \SUBBYTES[1].a/w705 , \SUBBYTES[1].a/w702 ,
         \SUBBYTES[1].a/w700 , \SUBBYTES[1].a/w699 , \SUBBYTES[1].a/w698 ,
         \SUBBYTES[1].a/w694 , \SUBBYTES[1].a/w692 , \SUBBYTES[1].a/w691 ,
         \SUBBYTES[1].a/w690 , \SUBBYTES[1].a/w689 , \SUBBYTES[1].a/w688 ,
         \SUBBYTES[1].a/w687 , \SUBBYTES[1].a/w686 , \SUBBYTES[1].a/w685 ,
         \SUBBYTES[1].a/w677 , \SUBBYTES[1].a/w675 , \SUBBYTES[1].a/w674 ,
         \SUBBYTES[1].a/w670 , \SUBBYTES[1].a/w668 , \SUBBYTES[1].a/w667 ,
         \SUBBYTES[1].a/w666 , \SUBBYTES[1].a/w662 , \SUBBYTES[1].a/w660 ,
         \SUBBYTES[1].a/w659 , \SUBBYTES[1].a/w646 , \SUBBYTES[1].a/w645 ,
         \SUBBYTES[1].a/w644 , \SUBBYTES[1].a/w642 , \SUBBYTES[1].a/w639 ,
         \SUBBYTES[1].a/w638 , \SUBBYTES[1].a/w636 , \SUBBYTES[1].a/w635 ,
         \SUBBYTES[1].a/w633 , \SUBBYTES[1].a/w631 , \SUBBYTES[1].a/w630 ,
         \SUBBYTES[1].a/w624 , \SUBBYTES[1].a/w623 , \SUBBYTES[1].a/w622 ,
         \SUBBYTES[1].a/w621 , \SUBBYTES[1].a/w615 , \SUBBYTES[1].a/w613 ,
         \SUBBYTES[1].a/w612 , \SUBBYTES[1].a/w608 , \SUBBYTES[1].a/w606 ,
         \SUBBYTES[1].a/w605 , \SUBBYTES[1].a/w600 , \SUBBYTES[1].a/w598 ,
         \SUBBYTES[1].a/w597 , \SUBBYTES[1].a/w581 , \SUBBYTES[1].a/w580 ,
         \SUBBYTES[1].a/w579 , \SUBBYTES[1].a/w578 , \SUBBYTES[1].a/w577 ,
         \SUBBYTES[1].a/w575 , \SUBBYTES[1].a/w574 , \SUBBYTES[1].a/w502 ,
         \SUBBYTES[1].a/w500 , \SUBBYTES[1].a/w499 , \SUBBYTES[1].a/w498 ,
         \SUBBYTES[1].a/w495 , \SUBBYTES[1].a/w493 , \SUBBYTES[1].a/w492 ,
         \SUBBYTES[1].a/w491 , \SUBBYTES[1].a/w487 , \SUBBYTES[1].a/w485 ,
         \SUBBYTES[1].a/w484 , \SUBBYTES[1].a/w483 , \SUBBYTES[1].a/w482 ,
         \SUBBYTES[1].a/w481 , \SUBBYTES[1].a/w480 , \SUBBYTES[1].a/w479 ,
         \SUBBYTES[1].a/w478 , \SUBBYTES[1].a/w470 , \SUBBYTES[1].a/w468 ,
         \SUBBYTES[1].a/w467 , \SUBBYTES[1].a/w463 , \SUBBYTES[1].a/w461 ,
         \SUBBYTES[1].a/w460 , \SUBBYTES[1].a/w459 , \SUBBYTES[1].a/w455 ,
         \SUBBYTES[1].a/w453 , \SUBBYTES[1].a/w452 , \SUBBYTES[1].a/w439 ,
         \SUBBYTES[1].a/w438 , \SUBBYTES[1].a/w437 , \SUBBYTES[1].a/w435 ,
         \SUBBYTES[1].a/w432 , \SUBBYTES[1].a/w431 , \SUBBYTES[1].a/w429 ,
         \SUBBYTES[1].a/w428 , \SUBBYTES[1].a/w426 , \SUBBYTES[1].a/w424 ,
         \SUBBYTES[1].a/w423 , \SUBBYTES[1].a/w417 , \SUBBYTES[1].a/w416 ,
         \SUBBYTES[1].a/w415 , \SUBBYTES[1].a/w414 , \SUBBYTES[1].a/w408 ,
         \SUBBYTES[1].a/w406 , \SUBBYTES[1].a/w405 , \SUBBYTES[1].a/w401 ,
         \SUBBYTES[1].a/w399 , \SUBBYTES[1].a/w398 , \SUBBYTES[1].a/w393 ,
         \SUBBYTES[1].a/w391 , \SUBBYTES[1].a/w390 , \SUBBYTES[1].a/w374 ,
         \SUBBYTES[1].a/w373 , \SUBBYTES[1].a/w372 , \SUBBYTES[1].a/w371 ,
         \SUBBYTES[1].a/w370 , \SUBBYTES[1].a/w368 , \SUBBYTES[1].a/w367 ,
         \SUBBYTES[1].a/w295 , \SUBBYTES[1].a/w293 , \SUBBYTES[1].a/w292 ,
         \SUBBYTES[1].a/w291 , \SUBBYTES[1].a/w288 , \SUBBYTES[1].a/w286 ,
         \SUBBYTES[1].a/w285 , \SUBBYTES[1].a/w284 , \SUBBYTES[1].a/w280 ,
         \SUBBYTES[1].a/w278 , \SUBBYTES[1].a/w277 , \SUBBYTES[1].a/w276 ,
         \SUBBYTES[1].a/w275 , \SUBBYTES[1].a/w274 , \SUBBYTES[1].a/w273 ,
         \SUBBYTES[1].a/w272 , \SUBBYTES[1].a/w271 , \SUBBYTES[1].a/w263 ,
         \SUBBYTES[1].a/w261 , \SUBBYTES[1].a/w260 , \SUBBYTES[1].a/w256 ,
         \SUBBYTES[1].a/w254 , \SUBBYTES[1].a/w253 , \SUBBYTES[1].a/w252 ,
         \SUBBYTES[1].a/w248 , \SUBBYTES[1].a/w246 , \SUBBYTES[1].a/w245 ,
         \SUBBYTES[1].a/w232 , \SUBBYTES[1].a/w231 , \SUBBYTES[1].a/w230 ,
         \SUBBYTES[1].a/w228 , \SUBBYTES[1].a/w225 , \SUBBYTES[1].a/w224 ,
         \SUBBYTES[1].a/w222 , \SUBBYTES[1].a/w221 , \SUBBYTES[1].a/w219 ,
         \SUBBYTES[1].a/w217 , \SUBBYTES[1].a/w216 , \SUBBYTES[1].a/w210 ,
         \SUBBYTES[1].a/w209 , \SUBBYTES[1].a/w208 , \SUBBYTES[1].a/w207 ,
         \SUBBYTES[1].a/w201 , \SUBBYTES[1].a/w199 , \SUBBYTES[1].a/w198 ,
         \SUBBYTES[1].a/w194 , \SUBBYTES[1].a/w192 , \SUBBYTES[1].a/w191 ,
         \SUBBYTES[1].a/w186 , \SUBBYTES[1].a/w184 , \SUBBYTES[1].a/w183 ,
         \SUBBYTES[1].a/w167 , \SUBBYTES[1].a/w166 , \SUBBYTES[1].a/w165 ,
         \SUBBYTES[1].a/w164 , \SUBBYTES[1].a/w163 , \SUBBYTES[1].a/w161 ,
         \SUBBYTES[1].a/w160 , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107,
         n108, n109, n110, n111, n112, n113, n114, n115, n116, n117, n118,
         n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210, n211, n212, n213, n214, n215, n216, n217,
         n218, n219, n220, n221, n222, n223, n224, n225, n226, n227, n228,
         n229, n230, n231, n232, n233, n234, n235, n236, n237, n238, n239,
         n240, n241, n242, n243, n244, n245, n246, n247, n248, n249, n250,
         n251, n252, n253, n254, n255, n256, n257, n258, n259, n260, n261,
         n262, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n282, n283,
         n284, n285, n286, n287, n288, n289, n290, n291, n292, n293, n294,
         n295, n296, n297, n298, n299, n300, n301, n302, n303, n304, n305,
         n306, n307, n308, n309, n310, n311, n312, n313, n314, n315, n316,
         n317, n318, n319, n320, n321, n322, n323, n324, n325, n326, n327,
         n328, n329, n330, n331, n332, n333, n334, n335, n336, n337, n338,
         n339, n340, n341, n342, n343, n344, n345, n346, n347, n348, n349,
         n350, n351, n352, n353, n354, n355, n356, n357, n358, n359, n360,
         n361, n362, n363, n364, n365, n366, n367, n368, n369, n370, n371,
         n372, n373, n374, n375, n376, n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635,
         n636, n637, n638, n639, n640, n641, n642, n643, n644, n645, n646,
         n647, n648, n649, n650, n651, n652, n653, n654, n655, n656, n657,
         n658, n659, n660, n661, n662, n663, n664, n665, n666, n667, n668,
         n669, n670, n671, n672, n673, n674, n675, n676, n677, n678, n679,
         n680, n681, n682, n683, n684, n685, n686, n687, n688, n689, n690,
         n691, n692, n693, n694, n695, n696, n697, n698, n699, n700, n701,
         n702, n703, n704, n705, n706, n707, n708, n709, n710, n711, n712,
         n713, n714, n715, n716, n717, n718, n719, n720, n721, n722, n723,
         n724, n725, n726, n727, n728, n729, n730, n731, n732, n733, n734,
         n735, n736, n737, n738, n739, n740, n741, n742, n743, n744, n745,
         n746, n747, n748, n749, n750, n751, n752, n753, n754, n755, n756,
         n757, n758, n759, n760, n761, n762, n763, n764, n765, n766, n767,
         n768, n769, n770, n771, n772, n773, n774, n775, n776, n777, n778,
         n779, n780, n781, n782, n783, n784, n785, n786, n787, n788, n789,
         n790, n791, n792, n793, n794, n795, n796, n797, n798, n799, n800,
         n801, n802, n803, n804, n805, n806, n807, n808, n809, n810, n811,
         n812, n813, n814, n815, n816, n817, n818, n819, n820, n821, n822,
         n823, n824, n825, n826, n827, n828, n829, n830, n831, n832, n833,
         n834, n835, n836, n837, n838, n839, n840, n841, n842, n843, n844,
         n845, n846, n847, n848, n849, n850, n851, n852, n853, n854, n855,
         n856, n857, n858, n859, n860, n861, n862, n863, n864, n865, n866,
         n867, n868, n869, n870, n871, n872, n873, n874, n875, n876, n877,
         n878, n879, n880, n881, n882, n883, n884, n885, n886, n887, n888,
         n889, n890, n891, n892, n893, n894, n895, n896, n897, n898, n899,
         n900, n901, n902, n903, n904, n905, n906, n907, n908, n909, n910,
         n911, n912, n913, n914, n915, n916, n917, n918, n919, n920, n921,
         n922, n923, n924, n925, n926, n927, n928, n929, n930, n931, n932,
         n933, n934, n935, n936, n937, n938, n939, n940, n941, n942, n943,
         n944, n945, n946, n947, n948, n949, n950, n951, n952, n953, n954,
         n955, n956, n957, n958, n959, n960, n961, n962, n963, n964, n965,
         n966, n967, n968, n969, n970, n971, n972, n973, n974, n975, n976,
         n977, n978, n979, n980, n981, n982, n983, n984, n985, n986, n987,
         n988, n989, n990, n991, n992, n993, n994, n995, n996, n997, n998,
         n999, n1000, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1031, n1032, n1033, n1034, n1035, n1036, n1037, n1038,
         n1039, n1040, n1041, n1042, n1043, n1044, n1045, n1046, n1047, n1048,
         n1049, n1050, n1051, n1052, n1053, n1054, n1055, n1056, n1057, n1058,
         n1059, n1060, n1061, n1062, n1063, n1064, n1065, n1066, n1067, n1068,
         n1069, n1070, n1071, n1072, n1073, n1074, n1075, n1076, n1077, n1078,
         n1079, n1080, n1081, n1082, n1083, n1084, n1085, n1086, n1087, n1088,
         n1089, n1090, n1091, n1092, n1093, n1094, n1095, n1096, n1097, n1098,
         n1099, n1100, n1101, n1102, n1103, n1104, n1105, n1106, n1107, n1108,
         n1109, n1110, n1111, n1112, n1113, n1114, n1115, n1116, n1117, n1118,
         n1119, n1120, n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1327, n1328,
         n1329, n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338,
         n1339, n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348,
         n1349, n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358,
         n1359, n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368,
         n1369, n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378,
         n1379, n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388,
         n1389, n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398,
         n1399, n1400, n1401, n1402, n1403, n1404, n1405, n1406, n1407, n1408,
         n1409, n1410, n1411, n1412, n1413, n1414, n1415, n1416, n1417, n1418,
         n1419, n1420, n1421, n1422, n1423, n1424, n1425, n1426, n1427, n1428,
         n1429, n1430, n1431, n1432, n1433, n1434, n1435, n1436, n1437, n1438,
         n1439, n1440, n1441, n1442, n1443, n1444, n1445, n1446, n1447, n1448,
         n1449, n1450, n1451, n1452, n1453, n1454, n1455, n1456, n1457, n1458,
         n1459, n1460, n1461, n1462, n1463, n1464, n1465, n1466, n1467, n1468,
         n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476, n1477, n1478,
         n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486, n1487, n1488,
         n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496, n1497, n1498,
         n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506, n1507, n1508,
         n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516, n1517, n1518,
         n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526, n1527, n1528,
         n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536, n1537, n1538,
         n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546, n1547, n1548,
         n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556, n1557, n1558,
         n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566, n1567, n1568,
         n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576, n1577, n1578,
         n1579, n1580, n1581, n1582, n1583, n1584, n1585, n1586, n1587, n1588,
         n1589, n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598,
         n1599, n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608,
         n1609, n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618,
         n1619, n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628,
         n1629, n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638,
         n1639, n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648,
         n1649, n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658,
         n1659, n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668,
         n1669, n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678,
         n1679, n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688,
         n1689, n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698,
         n1699, n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708,
         n1709, n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718,
         n1719, n1720, n1721, n1722, n1723, n1724, n1725, n1726, n1727, n1728,
         n1729, n1730, n1731, n1732, n1733, n1734, n1735, n1736, n1737, n1738,
         n1739, n1740, n1741, n1742, n1743, n1744, n1745, n1746, n1747, n1748,
         n1749, n1750, n1751, n1752, n1753, n1754, n1755, n1756, n1757, n1758,
         n1759, n1760, n1761, n1762, n1763, n1764, n1765, n1766, n1767, n1768,
         n1769, n1770, n1771, n1772, n1773, n1774, n1775, n1776, n1777, n1778,
         n1779, n1780, n1781, n1782, n1783, n1784, n1785, n1786, n1787, n1788,
         n1789, n1790, n1791, n1792, n1793, n1794, n1795, n1796, n1797, n1798,
         n1799, n1800, n1801, n1802, n1803, n1804, n1805, n1806, n1807, n1808,
         n1809, n1810, n1811, n1812, n1813, n1814, n1815, n1816, n1817, n1818,
         n1819, n1820, n1821, n1822, n1823, n1824, n1825, n1826, n1827, n1828,
         n1829, n1830, n1831, n1832, n1833, n1834, n1835, n1836, n1837, n1838,
         n1839, n1840, n1841, n1842, n1843, n1844, n1845, n1846, n1847, n1848,
         n1849, n1850, n1851, n1852, n1853, n1854, n1855, n1856, n1857, n1858,
         n1859, n1860, n1861, n1862, n1863, n1864, n1865, n1866, n1867, n1868,
         n1869, n1870, n1871, n1872, n1873, n1874, n1875, n1876, n1877, n1878,
         n1879, n1880, n1881, n1882, n1883, n1884, n1885, n1886, n1887, n1888,
         n1889, n1890, n1891, n1892, n1893, n1894, n1895, n1896, n1897, n1898,
         n1899, n1900, n1901, n1902, n1903, n1904, n1905, n1906, n1907, n1908,
         n1909, n1910, n1911, n1912, n1913, n1914, n1915, n1916, n1917, n1918,
         n1919, n1920, n1921, n1922, n1923, n1924, n1925, n1926, n1927, n1928,
         n1929, n1930, n1931, n1932, n1933, n1934, n1935, n1936, n1937, n1938,
         n1939, n1940, n1941, n1942, n1943, n1944, n1945, n1946, n1947, n1948,
         n1949, n1950, n1951, n1952, n1953, n1954, n1955, n1956, n1957, n1958,
         n1959, n1960, n1961, n1962, n1963, n1964, n1965, n1966, n1967, n1968,
         n1969, n1970, n1971, n1972, n1973, n1974, n1975, n1976, n1977, n1978,
         n1979, n1980, n1981, n1982, n1983, n1984, n1985, n1986, n1987, n1988,
         n1989, n1990, n1991, n1992, n1993, n1994, n1995, n1996, n1997, n1998,
         n1999, n2000, n2001, n2002, n2003, n2004, n2005, n2006, n2007, n2008,
         n2009, n2010, n2011, n2012, n2013, n2014, n2015, n2016, n2017, n2018,
         n2019, n2020, n2021, n2022, n2023, n2024, n2025, n2026, n2027, n2028,
         n2029, n2030, n2031, n2032, n2033, n2034, n2035, n2036, n2037, n2038,
         n2039, n2040, n2041, n2042, n2043, n2044, n2045, n2046, n2047, n2048,
         n2049, n2050, n2051, n2052, n2053, n2054, n2055, n2056, n2057, n2058,
         n2059, n2060, n2061, n2062, n2063, n2064, n2065, n2066, n2067, n2068,
         n2069, n2070, n2071, n2072, n2073, n2074, n2075, n2076, n2077, n2078,
         n2079, n2080, n2081, n2082, n2083, n2084, n2085, n2086, n2087, n2088,
         n2089, n2090, n2091, n2092, n2093, n2094, n2095, n2096, n2097, n2098,
         n2099, n2100, n2101, n2102, n2103, n2104, n2105, n2106, n2107, n2108,
         n2109, n2110, n2111, n2112, n2113, n2114, n2115, n2116, n2117, n2118,
         n2119, n2120, n2121, n2122, n2123, n2124, n2125, n2126, n2127, n2128,
         n2129, n2130, n2131, n2132, n2133, n2134, n2135, n2136, n2137, n2138,
         n2139, n2140, n2141, n2142, n2143, n2144, n2145, n2146, n2147, n2148,
         n2149, n2150, n2151, n2152, n2153, n2154, n2155, n2156, n2157, n2158,
         n2159, n2160, n2161, n2162, n2163, n2164, n2165, n2166, n2167, n2168,
         n2169, n2170, n2171, n2172, n2173, n2174, n2175, n2176, n2177, n2178,
         n2179, n2180, n2181, n2182, n2183, n2184, n2185, n2186, n2187, n2188,
         n2189, n2190, n2191, n2192, n2193, n2194, n2195, n2196, n2197, n2198,
         n2199, n2200, n2201, n2202, n2203, n2204, n2205, n2206, n2207, n2208,
         n2209, n2210, n2211, n2212, n2213, n2214, n2215, n2216, n2217, n2218,
         n2219, n2220, n2221, n2222, n2223, n2224, n2225, n2226, n2227, n2228,
         n2229, n2230, n2231, n2232, n2233, n2234, n2235, n2236, n2237, n2238,
         n2239, n2240, n2241, n2242, n2243, n2244, n2245, n2246, n2247, n2248,
         n2249, n2250, n2251, n2252, n2253, n2254, n2255, n2256, n2257, n2258,
         n2259, n2260, n2261, n2262, n2263, n2264, n2265, n2266, n2267, n2268,
         n2269, n2270, n2271, n2272, n2273, n2274, n2275, n2276, n2277, n2278,
         n2279, n2280, n2281, n2282, n2283, n2284, n2285, n2286, n2287, n2288,
         n2289, n2290, n2291, n2292, n2293, n2294, n2295, n2296, n2297, n2298,
         n2299, n2300, n2301, n2302, n2303, n2304, n2305, n2306, n2307, n2308,
         n2309, n2310, n2311, n2312, n2313, n2314, n2315, n2316, n2317, n2318,
         n2319, n2320, n2321, n2322, n2323, n2324, n2325, n2326, n2327, n2328,
         n2329, n2330, n2331, n2332, n2333, n2334, n2335, n2336, n2337, n2338,
         n2339, n2340, n2341, n2342, n2343, n2344, n2345, n2346, n2347, n2348,
         n2349, n2350, n2351, n2352, n2353, n2354, n2355, n2356, n2357, n2358,
         n2359, n2360, n2361, n2362, n2363, n2364, n2365, n2366, n2367, n2368,
         n2369, n2370, n2371, n2372, n2373, n2374, n2375, n2376, n2377, n2378,
         n2379, n2380, n2381, n2382, n2383, n2384, n2385, n2386, n2387, n2388,
         n2389, n2390, n2391, n2392, n2393, n2394, n2395, n2396, n2397, n2398,
         n2399, n2400, n2401, n2402, n2403, n2404, n2405, n2406, n2407, n2408,
         n2409, n2410, n2411, n2412, n2413, n2414, n2415, n2416, n2417, n2418,
         n2419, n2420, n2421, n2422, n2423, n2424, n2425, n2426, n2427, n2428,
         n2429, n2430, n2431, n2432, n2433, n2434, n2435, n2436, n2437, n2438,
         n2439, n2440, n2441, n2442, n2443, n2444, n2445, n2446, n2447, n2448,
         n2449, n2450, n2451, n2452, n2453, n2454, n2455, n2456, n2457, n2458,
         n2459, n2460, n2461, n2462, n2463, n2464, n2465, n2466, n2467, n2468,
         n2469, n2470, n2471, n2472, n2473, n2474, n2475, n2476, n2477, n2478,
         n2479, n2480, n2481, n2482, n2483, n2484, n2485, n2486, n2487, n2488,
         n2489, n2490, n2491, n2492, n2493, n2494, n2495, n2496, n2497, n2498,
         n2499, n2500, n2501, n2502, n2503, n2504, n2505, n2506, n2507, n2508,
         n2509, n2510, n2511, n2512, n2513, n2514, n2515, n2516, n2517, n2518,
         n2519, n2520, n2521, n2522, n2523, n2524, n2525, n2526, n2527, n2528,
         n2529, n2530, n2531, n2532, n2533, n2534, n2535, n2536, n2537, n2538,
         n2539, n2540, n2541, n2542, n2543, n2544, n2545, n2546, n2547, n2548,
         n2549, n2550, n2551, n2552, n2553, n2554, n2555, n2556, n2557, n2558,
         n2559, n2560, n2561, n2562, n2563, n2564, n2565, n2566, n2567, n2568,
         n2569, n2570, n2571, n2572, n2573, n2574, n2575, n2576, n2577, n2578,
         n2579, n2580, n2581, n2582, n2583, n2584, n2585, n2586, n2587, n2588,
         n2589, n2590, n2591, n2592, n2593, n2594, n2595, n2596, n2597, n2598,
         n2599, n2600, n2601, n2602, n2603, n2604, n2605, n2606, n2607, n2608,
         n2609, n2610, n2611, n2612, n2613, n2614, n2615, n2616, n2617, n2618,
         n2619, n2620, n2621, n2622, n2623, n2624, n2625, n2626, n2627, n2628,
         n2629, n2630, n2631, n2632, n2633, n2634, n2635, n2636, n2637, n2638,
         n2639, n2640, n2641, n2642, n2643, n2644, n2645, n2646, n2647, n2648,
         n2649, n2650, n2651, n2652, n2653, n2654, n2655, n2656, n2657, n2658,
         n2659, n2660, n2661, n2662, n2663, n2664, n2665, n2666, n2667, n2668,
         n2669, n2670, n2671, n2672, n2673, n2674, n2675, n2676, n2677, n2678,
         n2679, n2680, n2681, n2682, n2683, n2684, n2685, n2686, n2687, n2688,
         n2689, n2690, n2691, n2692, n2693, n2694, n2695, n2696, n2697, n2698,
         n2699, n2700, n2701, n2702, n2703, n2704, n2705, n2706, n2707, n2708,
         n2709, n2710, n2711, n2712, n2713, n2714, n2715, n2716, n2717, n2718,
         n2719, n2720, n2721, n2722, n2723, n2724, n2725, n2726, n2727, n2728,
         n2729, n2730, n2731, n2732, n2733, n2734, n2735, n2736, n2737, n2738,
         n2739, n2740, n2741, n2742, n2743, n2744, n2745, n2746, n2747, n2748,
         n2749, n2750, n2751, n2752, n2753, n2754, n2755, n2756, n2757, n2758,
         n2759, n2760, n2761, n2762, n2763, n2764, n2765, n2766, n2767, n2768,
         n2769, n2770, n2771, n2772, n2773, n2774, n2775, n2776, n2777, n2778,
         n2779, n2780, n2781, n2782, n2783, n2784, n2785, n2786, n2787, n2788,
         n2789, n2790, n2791, n2792, n2793, n2794, n2795, n2796, n2797, n2798,
         n2799, n2800, n2801, n2802, n2803, n2804, n2805, n2806, n2807, n2808,
         n2809, n2810, n2811, n2812, n2813, n2814, n2815, n2816, n2817, n2818,
         n2819, n2820, n2821, n2822, n2823, n2824, n2825, n2826, n2827, n2828,
         n2829, n2830, n2831, n2832, n2833, n2834, n2835, n2836, n2837, n2838,
         n2839, n2840, n2841, n2842, n2843, n2844, n2845, n2846, n2847, n2848,
         n2849, n2850, n2851, n2852, n2853, n2854, n2855, n2856, n2857, n2858,
         n2859, n2860, n2861, n2862, n2863, n2864, n2865, n2866, n2867, n2868,
         n2869, n2870, n2871, n2872, n2873, n2874, n2875, n2876, n2877, n2878,
         n2879, n2880, n2881, n2882, n2883, n2884, n2885, n2886, n2887, n2888,
         n2889, n2890, n2891, n2892, n2893, n2894, n2895, n2896, n2897, n2898,
         n2899, n2900, n2901, n2902, n2903, n2904, n2905, n2906, n2907, n2908,
         n2909, n2910, n2911, n2912, n2913, n2914, n2915, n2916, n2917, n2918,
         n2919, n2920, n2921, n2922, n2923, n2924, n2925, n2926, n2927, n2928,
         n2929, n2930, n2931, n2932, n2933, n2934, n2935, n2936, n2937, n2938,
         n2939, n2940, n2941, n2942, n2943, n2944, n2945, n2946, n2947, n2948,
         n2949, n2950, n2951, n2952, n2953, n2954, n2955, n2956, n2957, n2958,
         n2959, n2960, n2961, n2962, n2963, n2964, n2965, n2966, n2967, n2968,
         n2969, n2970, n2971, n2972, n2973, n2974, n2975, n2976, n2977, n2978,
         n2979, n2980, n2981, n2982, n2983, n2984, n2985, n2986, n2987, n2988,
         n2989, n2990, n2991, n2992, n2993, n2994, n2995, n2996, n2997, n2998,
         n2999, n3000, n3001, n3002, n3003, n3004, n3005, n3006, n3007, n3008,
         n3009, n3010, n3011, n3012, n3013, n3014, n3015, n3016, n3017, n3018,
         n3019, n3020, n3021, n3022, n3023, n3024, n3025, n3026, n3027, n3028,
         n3029, n3030, n3031, n3032, n3033, n3034, n3035, n3036, n3037, n3038,
         n3039, n3040, n3041, n3042, n3043, n3044, n3045, n3046, n3047, n3048,
         n3049, n3050, n3051, n3052, n3053, n3054, n3055, n3056, n3057, n3058,
         n3059, n3060, n3061, n3062, n3063, n3064, n3065, n3066, n3067, n3068,
         n3069, n3070, n3071, n3072, n3073, n3074, n3075, n3076, n3077, n3078,
         n3079, n3080, n3081, n3082, n3083, n3084, n3085, n3086, n3087, n3088,
         n3089, n3090, n3091, n3092, n3093, n3094, n3095, n3096, n3097, n3098,
         n3099, n3100, n3101, n3102, n3103, n3104, n3105, n3106, n3107, n3108,
         n3109, n3110, n3111, n3112, n3113, n3114, n3115, n3116, n3117, n3118,
         n3119, n3120, n3121, n3122, n3123, n3124, n3125, n3126, n3127, n3128,
         n3129, n3130, n3131, n3132, n3133, n3134, n3135, n3136, n3137, n3138,
         n3139, n3140, n3141, n3142, n3143, n3144, n3145, n3146, n3147, n3148,
         n3149, n3150, n3151, n3152, n3153, n3154, n3155, n3156, n3157, n3158,
         n3159, n3160, n3161, n3162, n3163, n3164, n3165, n3166, n3167, n3168,
         n3169, n3170, n3171, n3172, n3173, n3174, n3175, n3176, n3177, n3178,
         n3179, n3180, n3181, n3182, n3183, n3184, n3185, n3186, n3187, n3188,
         n3189, n3190, n3191, n3192, n3193, n3194, n3195, n3196, n3197, n3198,
         n3199, n3200, n3201, n3202, n3203, n3204, n3205, n3206, n3207, n3208,
         n3209, n3210, n3211, n3212, n3213, n3214, n3215, n3216, n3217, n3218,
         n3219, n3220, n3221, n3222, n3223, n3224, n3225, n3226, n3227, n3228,
         n3229, n3230, n3231, n3232, n3233, n3234, n3235, n3236, n3237, n3238,
         n3239, n3240, n3241, n3242, n3243, n3244, n3245, n3246, n3247, n3248,
         n3249, n3250, n3251, n3252, n3253, n3254, n3255, n3256, n3257, n3258,
         n3259, n3260, n3261, n3262, n3263, n3264, n3265, n3266, n3267, n3268,
         n3269, n3270, n3271, n3272, n3273, n3274, n3275, n3276, n3277, n3278,
         n3279, n3280, n3281, n3282, n3283, n3284, n3285, n3286, n3287, n3288,
         n3289, n3290, n3291, n3292, n3293, n3294, n3295, n3296, n3297, n3298,
         n3299, n3300, n3301, n3302, n3303, n3304, n3305, n3306, n3307, n3308,
         n3309, n3310, n3311, n3312, n3313, n3314, n3315, n3316, n3317, n3318,
         n3319, n3320, n3321, n3322, n3323, n3324, n3325, n3326, n3327, n3328,
         n3329, n3330, n3331, n3332, n3333, n3334, n3335, n3336, n3337, n3338,
         n3339, n3340, n3341, n3342, n3343, n3344, n3345, n3346, n3347, n3348,
         n3349, n3350, n3351, n3352, n3353, n3354, n3355, n3356, n3357, n3358,
         n3359, n3360, n3361, n3362, n3363, n3364, n3365, n3366, n3367, n3368,
         n3369, n3370, n3371, n3372, n3373, n3374, n3375, n3376, n3377, n3378,
         n3379, n3380, n3381, n3382, n3383, n3384, n3385, n3386, n3387, n3388,
         n3389, n3390, n3391, n3392, n3393, n3394, n3395, n3396, n3397, n3398,
         n3399, n3400, n3401, n3402, n3403, n3404, n3405, n3406, n3407, n3408,
         n3409, n3410, n3411, n3412, n3413, n3414, n3415, n3416, n3417, n3418,
         n3419, n3420, n3421, n3422, n3423, n3424, n3425, n3426, n3427, n3428,
         n3429, n3430, n3431, n3432, n3433, n3434, n3435, n3436, n3437, n3438,
         n3439, n3440, n3441, n3442, n3443, n3444, n3445, n3446, n3447, n3448,
         n3449, n3450, n3451, n3452, n3453, n3454, n3455, n3456, n3457, n3458,
         n3459, n3460, n3461, n3462, n3463, n3464, n3465, n3466, n3467, n3468,
         n3469, n3470, n3471, n3472, n3473, n3474, n3475, n3476, n3477, n3478,
         n3479, n3480, n3481, n3482, n3483, n3484, n3485, n3486, n3487, n3488,
         n3489, n3490, n3491, n3492, n3493, n3494, n3495, n3496, n3497, n3498,
         n3499, n3500, n3501, n3502, n3503, n3504, n3505, n3506, n3507, n3508,
         n3509, n3510, n3511, n3512, n3513, n3514, n3515, n3516, n3517, n3518,
         n3519, n3520, n3521, n3522, n3523, n3524, n3525, n3526, n3527, n3528,
         n3529, n3530, n3531, n3532, n3533, n3534, n3535, n3536, n3537, n3538,
         n3539, n3540, n3541, n3542, n3543, n3544, n3545, n3546, n3547, n3548,
         n3549, n3550, n3551, n3552, n3553, n3554, n3555, n3556, n3557, n3558,
         n3559, n3560, n3561, n3562, n3563, n3564, n3565, n3566, n3567, n3568,
         n3569, n3570, n3571, n3572, n3573, n3574, n3575, n3576, n3577, n3578,
         n3579, n3580, n3581, n3582, n3583, n3584, n3585, n3586, n3587, n3588,
         n3589, n3590, n3591, n3592, n3593, n3594, n3595, n3596, n3597, n3598,
         n3599, n3600, n3601, n3602, n3603, n3604, n3605, n3606, n3607, n3608,
         n3609, n3610, n3611, n3612, n3613, n3614, n3615, n3616, n3617, n3618,
         n3619, n3620, n3621, n3622, n3623, n3624, n3625, n3626, n3627, n3628,
         n3629, n3630, n3631, n3632, n3633, n3634, n3635, n3636, n3637, n3638,
         n3639, n3640, n3641, n3642, n3643, n3644, n3645, n3646, n3647, n3648,
         n3649, n3650, n3651, n3652, n3653, n3654, n3655, n3656, n3657, n3658,
         n3659, n3660, n3661, n3662, n3663, n3664, n3665, n3666, n3667, n3668,
         n3669, n3670, n3671, n3672, n3673, n3674, n3675, n3676, n3677, n3678,
         n3679, n3680, n3681, n3682, n3683, n3684, n3685, n3686, n3687, n3688,
         n3689, n3690, n3691, n3692, n3693, n3694, n3695, n3696, n3697, n3698,
         n3699, n3700, n3701, n3702, n3703, n3704, n3705, n3706, n3707, n3708,
         n3709, n3710, n3711, n3712, n3713, n3714, n3715, n3716, n3717, n3718,
         n3719, n3720, n3721, n3722, n3723, n3724, n3725, n3726, n3727, n3728,
         n3729, n3730, n3731, n3732, n3733, n3734, n3735, n3736, n3737, n3738,
         n3739, n3740, n3741, n3742, n3743, n3744, n3745, n3746, n3747, n3748,
         n3749, n3750, n3751, n3752, n3753, n3754, n3755, n3756, n3757, n3758,
         n3759, n3760, n3761, n3762, n3763, n3764, n3765, n3766, n3767, n3768,
         n3769, n3770, n3771, n3772, n3773, n3774, n3775, n3776, n3777, n3778,
         n3779, n3780, n3781, n3782, n3783, n3784, n3785, n3786, n3787, n3788,
         n3789, n3790, n3791, n3792, n3793, n3794, n3795, n3796, n3797, n3798,
         n3799, n3800, n3801, n3802, n3803, n3804, n3805, n3806, n3807, n3808,
         n3809, n3810, n3811, n3812, n3813, n3814, n3815, n3816, n3817, n3818,
         n3819, n3820, n3821, n3822, n3823, n3824, n3825, n3826, n3827, n3828,
         n3829, n3830, n3831, n3832, n3833, n3834, n3835, n3836, n3837, n3838,
         n3839, n3840, n3841, n3842, n3843, n3844, n3845, n3846, n3847, n3848,
         n3849, n3850, n3851, n3852, n3853, n3854, n3855, n3856, n3857, n3858,
         n3859, n3860, n3861, n3862, n3863, n3864, n3865, n3866, n3867, n3868,
         n3869, n3870, n3871, n3872, n3873, n3874, n3875, n3876, n3877, n3878,
         n3879, n3880, n3881, n3882, n3883, n3884, n3885, n3886, n3887, n3888,
         n3889, n3890, n3891, n3892, n3893, n3894, n3895, n3896, n3897, n3898,
         n3899, n3900, n3901, n3902, n3903, n3904, n3905, n3906, n3907, n3908,
         n3909, n3910, n3911, n3912, n3913, n3914, n3915, n3916, n3917, n3918,
         n3919, n3920, n3921, n3922, n3923, n3924, n3925, n3926, n3927, n3928,
         n3929, n3930, n3931, n3932, n3933, n3934, n3935, n3936, n3937, n3938,
         n3939, n3940, n3941, n3942, n3943, n3944, n3945, n3946, n3947, n3948,
         n3949, n3950, n3951, n3952, n3953, n3954, n3955, n3956, n3957, n3958,
         n3959, n3960, n3961, n3962, n3963, n3964, n3965, n3966, n3967, n3968,
         n3969, n3970, n3971, n3972, n3973, n3974, n3975, n3976, n3977, n3978,
         n3979, n3980, n3981, n3982, n3983, n3984, n3985, n3986, n3987, n3988,
         n3989, n3990, n3991, n3992, n3993, n3994, n3995, n3996, n3997, n3998,
         n3999, n4000, n4001, n4002, n4003, n4004, n4005, n4006, n4007, n4008,
         n4009, n4010, n4011, n4012, n4013, n4014, n4015, n4016, n4017, n4018,
         n4019, n4020, n4021, n4022, n4023, n4024, n4025, n4026, n4027, n4028,
         n4029, n4030, n4031, n4032, n4033, n4034, n4035, n4036, n4037, n4038,
         n4039, n4040, n4041, n4042, n4043, n4044, n4045, n4046, n4047, n4048,
         n4049, n4050, n4051, n4052, n4053, n4054, n4055, n4056, n4057, n4058,
         n4059, n4060, n4061, n4062, n4063, n4064, n4065, n4066, n4067, n4068,
         n4069, n4070, n4071, n4072, n4073, n4074, n4075, n4076, n4077, n4078,
         n4079, n4080, n4081, n4082, n4083, n4084, n4085, n4086, n4087, n4088,
         n4089, n4090, n4091, n4092, n4093, n4094, n4095, n4096, n4097, n4098,
         n4099, n4100, n4101, n4102, n4103, n4104, n4105, n4106, n4107, n4108,
         n4109, n4110, n4111, n4112, n4113, n4114, n4115, n4116, n4117, n4118,
         n4119, n4120, n4121, n4122, n4123, n4124, n4125, n4126, n4127, n4128,
         n4129, n4130, n4131, n4132, n4133, n4134, n4135, n4136, n4137, n4138,
         n4139, n4140, n4141, n4142, n4143, n4144, n4145, n4146, n4147, n4148,
         n4149, n4150, n4151, n4152, n4153, n4154, n4155, n4156, n4157, n4158,
         n4159, n4160, n4161, n4162, n4163, n4164, n4165, n4166, n4167, n4168,
         n4169, n4170, n4171, n4172, n4173, n4174, n4175, n4176, n4177, n4178,
         n4179, n4180, n4181, n4182, n4183, n4184, n4185, n4186, n4187, n4188,
         n4189, n4190, n4191, n4192, n4193, n4194, n4195, n4196, n4197, n4198,
         n4199, n4200, n4201, n4202, n4203, n4204, n4205, n4206, n4207, n4208,
         n4209, n4210, n4211, n4212, n4213, n4214, n4215, n4216, n4217, n4218,
         n4219, n4220, n4221, n4222, n4223, n4224, n4225, n4226, n4227, n4228,
         n4229, n4230, n4231, n4232, n4233, n4234, n4235, n4236, n4237, n4238,
         n4239, n4240, n4241, n4242, n4243, n4244, n4245, n4246, n4247, n4248,
         n4249, n4250, n4251, n4252, n4253, n4254, n4255, n4256, n4257, n4258,
         n4259, n4260, n4261, n4262, n4263, n4264, n4265, n4266, n4267, n4268,
         n4269, n4270, n4271, n4272, n4273, n4274, n4275, n4276, n4277, n4278,
         n4279, n4280, n4281, n4282, n4283, n4284, n4285, n4286, n4287, n4288,
         n4289, n4290, n4291, n4292, n4293, n4294, n4295, n4296, n4297, n4298,
         n4299, n4300, n4301, n4302, n4303, n4304, n4305, n4306, n4307, n4308,
         n4309, n4310, n4311, n4312, n4313, n4314, n4315, n4316, n4317, n4318,
         n4319, n4320, n4321, n4322, n4323, n4324, n4325, n4326, n4327, n4328,
         n4329, n4330, n4331, n4332, n4333, n4334, n4335, n4336, n4337, n4338,
         n4339, n4340, n4341, n4342, n4343, n4344, n4345, n4346, n4347, n4348,
         n4349, n4350, n4351, n4352, n4353, n4354, n4355, n4356, n4357, n4358,
         n4359, n4360, n4361, n4362, n4363, n4364, n4365, n4366, n4367, n4368,
         n4369, n4370, n4371, n4372, n4373, n4374, n4375, n4376, n4377, n4378,
         n4379, n4380, n4381, n4382, n4383, n4384, n4385, n4386, n4387, n4388,
         n4389, n4390, n4391, n4392, n4393, n4394, n4395, n4396, n4397, n4398,
         n4399, n4400, n4401, n4402, n4403, n4404, n4405, n4406, n4407, n4408,
         n4409, n4410, n4411, n4412, n4413, n4414, n4415, n4416, n4417, n4418,
         n4419, n4420, n4421, n4422, n4423, n4424, n4425, n4426, n4427, n4428,
         n4429, n4430, n4431, n4432, n4433, n4434, n4435, n4436, n4437, n4438,
         n4439, n4440, n4441, n4442, n4443, n4444, n4445, n4446, n4447, n4448,
         n4449, n4450, n4451, n4452, n4453, n4454, n4455, n4456, n4457, n4458,
         n4459, n4460, n4461, n4462, n4463, n4464, n4465, n4466, n4467, n4468,
         n4469, n4470, n4471, n4472, n4473, n4474, n4475, n4476, n4477, n4478,
         n4479, n4480, n4481, n4482, n4483, n4484, n4485, n4486, n4487, n4488,
         n4489, n4490, n4491, n4492, n4493, n4494, n4495, n4496, n4497, n4498,
         n4499, n4500, n4501, n4502, n4503, n4504, n4505, n4506, n4507, n4508,
         n4509, n4510, n4511, n4512, n4513, n4514, n4515, n4516, n4517, n4518,
         n4519, n4520, n4521, n4522, n4523, n4524, n4525, n4526, n4527, n4528,
         n4529, n4530, n4531, n4532, n4533, n4534, n4535, n4536, n4537, n4538,
         n4539, n4540, n4541, n4542, n4543, n4544, n4545, n4546, n4547, n4548,
         n4549, n4550, n4551, n4552, n4553, n4554, n4555, n4556, n4557, n4558,
         n4559, n4560, n4561, n4562, n4563, n4564, n4565, n4566, n4567, n4568,
         n4569, n4570, n4571, n4572, n4573, n4574, n4575, n4576, n4577, n4578,
         n4579, n4580, n4581, n4582, n4583, n4584, n4585, n4586, n4587, n4588,
         n4589, n4590, n4591, n4592, n4593, n4594, n4595, n4596, n4597, n4598,
         n4599, n4600, n4601, n4602, n4603, n4604, n4605, n4606, n4607, n4608,
         n4609, n4610, n4611, n4612, n4613, n4614, n4615, n4616, n4617, n4618,
         n4619, n4620, n4621, n4622, n4623, n4624, n4625, n4626, n4627, n4628,
         n4629, n4630, n4631, n4632, n4633, n4634, n4635, n4636, n4637, n4638,
         n4639, n4640, n4641, n4642, n4643, n4644, n4645, n4646, n4647, n4648,
         n4649, n4650, n4651, n4652, n4653, n4654, n4655, n4656, n4657, n4658,
         n4659, n4660, n4661, n4662, n4663, n4664, n4665, n4666, n4667, n4668,
         n4669, n4670, n4671, n4672, n4673, n4674, n4675, n4676, n4677, n4678,
         n4679, n4680, n4681, n4682, n4683, n4684, n4685, n4686, n4687, n4688,
         n4689, n4690, n4691, n4692, n4693, n4694, n4695, n4696, n4697, n4698,
         n4699, n4700, n4701, n4702, n4703, n4704, n4705, n4706, n4707, n4708,
         n4709, n4710, n4711, n4712, n4713, n4714, n4715, n4716, n4717, n4718,
         n4719, n4720, n4721, n4722, n4723, n4724, n4725, n4726, n4727, n4728,
         n4729, n4730, n4731, n4732, n4733, n4734, n4735, n4736, n4737, n4738,
         n4739, n4740, n4741, n4742, n4743, n4744, n4745, n4746, n4747, n4748,
         n4749, n4750, n4751, n4752, n4753, n4754, n4755, n4756, n4757, n4758,
         n4759, n4760, n4761, n4762, n4763, n4764, n4765, n4766, n4767, n4768,
         n4769, n4770, n4771, n4772, n4773, n4774, n4775, n4776, n4777, n4778,
         n4779, n4780, n4781, n4782, n4783, n4784, n4785, n4786, n4787, n4788,
         n4789, n4790, n4791, n4792, n4793, n4794, n4795, n4796, n4797, n4798,
         n4799, n4800, n4801, n4802, n4803, n4804, n4805, n4806, n4807, n4808,
         n4809, n4810, n4811, n4812, n4813, n4814, n4815, n4816, n4817, n4818,
         n4819, n4820, n4821, n4822, n4823, n4824, n4825, n4826, n4827, n4828,
         n4829, n4830, n4831, n4832, n4833, n4834, n4835, n4836, n4837, n4838,
         n4839, n4840, n4841, n4842, n4843, n4844, n4845, n4846, n4847, n4848,
         n4849, n4850, n4851, n4852, n4853, n4854, n4855, n4856, n4857, n4858,
         n4859, n4860, n4861, n4862, n4863, n4864, n4865, n4866, n4867, n4868,
         n4869, n4870, n4871, n4872, n4873, n4874, n4875, n4876, n4877, n4878,
         n4879, n4880, n4881, n4882, n4883, n4884, n4885, n4886, n4887, n4888,
         n4889, n4890, n4891, n4892, n4893, n4894, n4895, n4896, n4897, n4898,
         n4899, n4900, n4901, n4902, n4903, n4904, n4905, n4906, n4907, n4908,
         n4909, n4910, n4911, n4912, n4913, n4914, n4915, n4916, n4917, n4918,
         n4919, n4920, n4921, n4922, n4923, n4924, n4925, n4926, n4927, n4928,
         n4929, n4930, n4931, n4932, n4933, n4934, n4935, n4936, n4937, n4938,
         n4939, n4940, n4941, n4942, n4943, n4944, n4945, n4946, n4947, n4948,
         n4949, n4950, n4951, n4952, n4953, n4954, n4955, n4956, n4957, n4958,
         n4959, n4960, n4961, n4962, n4963, n4964, n4965, n4966, n4967, n4968,
         n4969, n4970, n4971, n4972, n4973, n4974, n4975, n4976, n4977, n4978,
         n4979, n4980, n4981, n4982, n4983, n4984, n4985, n4986, n4987, n4988,
         n4989, n4990, n4991, n4992, n4993, n4994, n4995, n4996, n4997, n4998,
         n4999, n5000, n5001, n5002, n5003, n5004, n5005, n5006, n5007, n5008,
         n5009, n5010, n5011, n5012, n5013, n5014, n5015, n5016, n5017, n5018,
         n5019, n5020, n5021, n5022, n5023, n5024, n5025, n5026, n5027, n5028,
         n5029, n5030, n5031, n5032, n5033, n5034, n5035, n5036, n5037, n5038,
         n5039, n5040, n5041, n5042, n5043, n5044, n5045, n5046, n5047, n5048,
         n5049, n5050, n5051, n5052, n5053, n5054, n5055, n5056, n5057, n5058,
         n5059, n5060, n5061, n5062, n5063, n5064, n5065, n5066, n5067, n5068,
         n5069, n5070, n5071, n5072, n5073, n5074, n5075, n5076, n5077, n5078,
         n5079, n5080, n5081, n5082, n5083, n5084, n5085, n5086, n5087, n5088,
         n5089, n5090, n5091, n5092, n5093, n5094, n5095, n5096, n5097, n5098,
         n5099, n5100, n5101, n5102, n5103, n5104, n5105, n5106, n5107, n5108,
         n5109, n5110, n5111, n5112, n5113, n5114, n5115, n5116, n5117, n5118,
         n5119, n5120, n5121, n5122, n5123, n5124, n5125, n5126, n5127, n5128,
         n5129, n5130, n5131, n5132, n5133, n5134, n5135, n5136, n5137, n5138,
         n5139, n5140, n5141, n5142, n5143, n5144, n5145, n5146, n5147, n5148,
         n5149, n5150, n5151, n5152, n5153, n5154, n5155, n5156, n5157, n5158,
         n5159, n5160, n5161, n5162, n5163, n5164, n5165, n5166, n5167, n5168,
         n5169, n5170, n5171, n5172, n5173, n5174, n5175, n5176, n5177, n5178,
         n5179, n5180, n5181, n5182, n5183, n5184, n5185, n5186, n5187, n5188,
         n5189, n5190, n5191, n5192, n5193, n5194, n5195, n5196, n5197, n5198,
         n5199, n5200, n5201, n5202, n5203, n5204, n5205, n5206, n5207, n5208,
         n5209, n5210, n5211, n5212, n5213, n5214, n5215, n5216, n5217, n5218,
         n5219, n5220, n5221, n5222, n5223, n5224, n5225, n5226, n5227, n5228,
         n5229, n5230, n5231, n5232, n5233, n5234, n5235, n5236, n5237, n5238,
         n5239, n5240, n5241, n5242, n5243, n5244, n5245, n5246, n5247, n5248,
         n5249, n5250, n5251, n5252, n5253, n5254, n5255, n5256, n5257, n5258,
         n5259, n5260, n5261, n5262, n5263, n5264, n5265, n5266, n5267, n5268,
         n5269, n5270, n5271, n5272, n5273, n5274, n5275, n5276, n5277, n5278,
         n5279, n5280, n5281, n5282, n5283, n5284, n5285, n5286, n5287, n5288,
         n5289, n5290, n5291, n5292, n5293, n5294, n5295, n5296, n5297, n5298,
         n5299, n5300, n5301, n5302, n5303, n5304, n5305, n5306, n5307, n5308,
         n5309, n5310, n5311, n5312, n5313, n5314, n5315, n5316, n5317, n5318,
         n5319, n5320, n5321, n5322, n5323, n5324, n5325, n5326, n5327, n5328,
         n5329, n5330, n5331, n5332, n5333, n5334, n5335, n5336, n5337, n5338,
         n5339, n5340, n5341, n5342, n5343, n5344, n5345, n5346, n5347, n5348,
         n5349, n5350, n5351, n5352, n5353, n5354, n5355, n5356, n5357, n5358,
         n5359, n5360, n5361, n5362, n5363, n5364, n5365, n5366, n5367, n5368,
         n5369, n5370, n5371, n5372, n5373, n5374, n5375, n5376, n5377, n5378,
         n5379, n5380, n5381, n5382, n5383, n5384, n5385, n5386, n5387, n5388,
         n5389, n5390, n5391, n5392, n5393, n5394, n5395, n5396, n5397, n5398,
         n5399, n5400, n5401, n5402, n5403, n5404, n5405, n5406, n5407, n5408,
         n5409, n5410, n5411, n5412, n5413, n5414, n5415, n5416, n5417, n5418,
         n5419, n5420, n5421, n5422, n5423, n5424, n5425, n5426, n5427, n5428,
         n5429, n5430, n5431, n5432, n5433, n5434, n5435, n5436, n5437, n5438,
         n5439, n5440, n5441, n5442, n5443, n5444, n5445, n5446, n5447, n5448,
         n5449, n5450, n5451, n5452, n5453, n5454, n5455, n5456, n5457, n5458,
         n5459, n5460, n5461, n5462, n5463, n5464, n5465, n5466, n5467, n5468,
         n5469, n5470, n5471, n5472, n5473, n5474, n5475, n5476, n5477, n5478,
         n5479, n5480, n5481, n5482, n5483, n5484, n5485, n5486, n5487, n5488,
         n5489, n5490, n5491, n5492, n5493, n5494, n5495, n5496, n5497, n5498,
         n5499, n5500, n5501, n5502, n5503, n5504, n5505, n5506, n5507, n5508,
         n5509, n5510, n5511, n5512, n5513, n5514, n5515, n5516, n5517, n5518,
         n5519, n5520, n5521, n5522, n5523, n5524, n5525, n5526, n5527, n5528,
         n5529, n5530, n5531, n5532, n5533, n5534, n5535, n5536, n5537, n5538,
         n5539, n5540, n5541, n5542, n5543, n5544, n5545, n5546, n5547, n5548,
         n5549, n5550, n5551, n5552, n5553, n5554, n5555, n5556, n5557, n5558,
         n5559, n5560, n5561, n5562, n5563, n5564, n5565, n5566, n5567, n5568,
         n5569, n5570, n5571, n5572, n5573, n5574, n5575, n5576, n5577, n5578,
         n5579, n5580, n5581, n5582, n5583, n5584, n5585, n5586, n5587, n5588,
         n5589, n5590, n5591, n5592, n5593, n5594, n5595, n5596, n5597, n5598,
         n5599, n5600, n5601, n5602, n5603, n5604, n5605, n5606, n5607, n5608,
         n5609, n5610, n5611, n5612, n5613, n5614, n5615, n5616, n5617, n5618,
         n5619, n5620, n5621, n5622, n5623, n5624, n5625, n5626, n5627, n5628,
         n5629, n5630, n5631, n5632, n5633, n5634, n5635, n5636, n5637, n5638,
         n5639, n5640, n5641, n5642, n5643, n5644, n5645, n5646, n5647, n5648,
         n5649, n5650, n5651, n5652, n5653, n5654, n5655, n5656, n5657, n5658,
         n5659, n5660, n5661, n5662, n5663, n5664, n5665, n5666, n5667, n5668,
         n5669, n5670, n5671, n5672, n5673, n5674, n5675, n5676, n5677, n5678,
         n5679, n5680, n5681, n5682, n5683, n5684, n5685, n5686, n5687, n5688,
         n5689, n5690, n5691, n5692, n5693, n5694, n5695, n5696, n5697, n5698,
         n5699, n5700, n5701, n5702, n5703, n5704, n5705, n5706, n5707, n5708,
         n5709, n5710, n5711, n5712, n5713, n5714, n5715, n5716, n5717, n5718,
         n5719, n5720, n5721, n5722, n5723, n5724, n5725, n5726, n5727, n5728,
         n5729, n5730, n5731, n5732, n5733, n5734, n5735, n5736, n5737, n5738,
         n5739, n5740, n5741, n5742, n5743, n5744, n5745, n5746, n5747, n5748,
         n5749, n5750, n5751, n5752, n5753, n5754, n5755, n5756, n5757, n5758,
         n5759, n5760, n5761, n5762, n5763, n5764, n5765, n5766, n5767, n5768,
         n5769, n5770, n5771, n5772, n5773, n5774, n5775, n5776, n5777, n5778,
         n5779, n5780, n5781, n5782, n5783, n5784, n5785, n5786, n5787, n5788,
         n5789, n5790, n5791, n5792, n5793, n5794, n5795, n5796, n5797, n5798,
         n5799, n5800, n5801, n5802, n5803, n5804, n5805, n5806, n5807, n5808,
         n5809, n5810, n5811, n5812, n5813, n5814, n5815, n5816, n5817, n5818,
         n5819, n5820, n5821, n5822, n5823, n5824, n5825, n5826, n5827, n5828,
         n5829, n5830, n5831, n5832, n5833, n5834, n5835, n5836, n5837, n5838,
         n5839, n5840, n5841, n5842, n5843, n5844, n5845, n5846, n5847, n5848,
         n5849, n5850, n5851, n5852, n5853, n5854, n5855, n5856, n5857, n5858,
         n5859, n5860, n5861, n5862, n5863, n5864, n5865, n5866, n5867, n5868,
         n5869, n5870, n5871, n5872, n5873, n5874, n5875, n5876, n5877, n5878,
         n5879, n5880, n5881, n5882, n5883, n5884, n5885, n5886, n5887, n5888,
         n5889, n5890, n5891, n5892, n5893, n5894, n5895, n5896, n5897, n5898,
         n5899, n5900, n5901, n5902, n5903, n5904, n5905, n5906, n5907, n5908,
         n5909, n5910, n5911, n5912, n5913, n5914, n5915, n5916, n5917, n5918,
         n5919, n5920, n5921, n5922, n5923, n5924, n5925, n5926, n5927, n5928,
         n5929, n5930, n5931, n5932, n5933, n5934, n5935, n5936, n5937, n5938,
         n5939, n5940, n5941, n5942, n5943, n5944, n5945, n5946, n5947, n5948,
         n5949, n5950, n5951, n5952, n5953, n5954, n5955, n5956, n5957, n5958,
         n5959, n5960, n5961, n5962, n5963, n5964, n5965, n5966, n5967, n5968,
         n5969, n5970, n5971, n5972, n5973, n5974, n5975, n5976, n5977, n5978,
         n5979, n5980, n5981, n5982, n5983, n5984, n5985, n5986, n5987, n5988,
         n5989, n5990, n5991, n5992, n5993, n5994, n5995, n5996, n5997, n5998,
         n5999, n6000, n6001, n6002, n6003, n6004, n6005, n6006, n6007, n6008,
         n6009, n6010, n6011, n6012, n6013, n6014, n6015, n6016, n6017, n6018,
         n6019, n6020, n6021, n6022, n6023, n6024, n6025, n6026, n6027, n6028,
         n6029, n6030, n6031, n6032, n6033, n6034, n6035, n6036, n6037, n6038,
         n6039, n6040, n6041, n6042, n6043, n6044, n6045, n6046, n6047, n6048,
         n6049, n6050, n6051, n6052, n6053, n6054, n6055, n6056, n6057, n6058,
         n6059, n6060, n6061, n6062, n6063, n6064, n6065, n6066, n6067, n6068,
         n6069, n6070, n6071, n6072, n6073, n6074, n6075, n6076, n6077, n6078,
         n6079, n6080, n6081, n6082, n6083, n6084, n6085, n6086, n6087, n6088,
         n6089, n6090, n6091, n6092, n6093, n6094, n6095, n6096, n6097, n6098,
         n6099, n6100, n6101, n6102, n6103, n6104, n6105, n6106, n6107, n6108,
         n6109, n6110, n6111, n6112, n6113, n6114, n6115, n6116, n6117, n6118,
         n6119, n6120, n6121, n6122, n6123, n6124, n6125, n6126, n6127, n6128,
         n6129, n6130, n6131, n6132, n6133, n6134, n6135, n6136, n6137, n6138,
         n6139, n6140, n6141, n6142, n6143, n6144, n6145, n6146, n6147, n6148,
         n6149, n6150, n6151, n6152, n6153, n6154, n6155, n6156, n6157, n6158,
         n6159, n6160, n6161, n6162, n6163, n6164, n6165, n6166, n6167, n6168,
         n6169, n6170, n6171, n6172, n6173, n6174, n6175, n6176, n6177, n6178,
         n6179, n6180, n6181, n6182, n6183, n6184, n6185, n6186, n6187, n6188,
         n6189, n6190, n6191, n6192, n6193, n6194, n6195, n6196, n6197, n6198,
         n6199, n6200, n6201, n6202, n6203, n6204, n6205, n6206, n6207, n6208,
         n6209, n6210, n6211, n6212, n6213, n6214, n6215, n6216, n6217, n6218,
         n6219, n6220, n6221, n6222, n6223, n6224, n6225, n6226, n6227, n6228,
         n6229, n6230, n6231, n6232, n6233, n6234, n6235, n6236, n6237, n6238,
         n6239, n6240, n6241, n6242, n6243, n6244, n6245, n6246, n6247, n6248,
         n6249, n6250, n6251, n6252, n6253, n6254, n6255, n6256, n6257, n6258,
         n6259, n6260, n6261, n6262, n6263, n6264, n6265, n6266, n6267, n6268,
         n6269, n6270, n6271, n6272, n6273, n6274, n6275, n6276, n6277, n6278,
         n6279, n6280, n6281, n6282, n6283, n6284, n6285, n6286, n6287, n6288,
         n6289, n6290, n6291, n6292, n6293, n6294, n6295, n6296, n6297, n6298,
         n6299, n6300, n6301, n6302, n6303, n6304, n6305, n6306, n6307, n6308,
         n6309, n6310, n6311, n6312, n6313, n6314, n6315, n6316, n6317, n6318,
         n6319, n6320, n6321, n6322, n6323, n6324, n6325, n6326, n6327, n6328,
         n6329, n6330, n6331, n6332, n6333, n6334, n6335, n6336, n6337, n6338,
         n6339, n6340, n6341, n6342, n6343, n6344, n6345, n6346, n6347, n6348,
         n6349, n6350, n6351, n6352, n6353, n6354, n6355, n6356, n6357, n6358,
         n6359, n6360, n6361, n6362, n6363, n6364, n6365, n6366, n6367, n6368,
         n6369, n6370, n6371, n6372, n6373, n6374, n6375, n6376, n6377, n6378,
         n6379, n6380, n6381, n6382, n6383, n6384, n6385, n6386, n6387, n6388,
         n6389, n6390, n6391, n6392, n6393, n6394, n6395, n6396, n6397, n6398,
         n6399, n6400, n6401, n6402, n6403, n6404, n6405, n6406, n6407, n6408,
         n6409, n6410, n6411, n6412, n6413, n6414, n6415, n6416, n6417, n6418,
         n6419, n6420, n6421, n6422, n6423, n6424, n6425, n6426, n6427, n6428,
         n6429, n6430, n6431, n6432, n6433, n6434, n6435, n6436, n6437, n6438,
         n6439, n6440, n6441, n6442, n6443, n6444, n6445, n6446, n6447, n6448,
         n6449, n6450, n6451, n6452, n6453, n6454, n6455, n6456, n6457, n6458,
         n6459, n6460, n6461, n6462, n6463, n6464, n6465, n6466, n6467, n6468,
         n6469, n6470, n6471, n6472, n6473, n6474, n6475, n6476, n6477, n6478,
         n6479, n6480, n6481, n6482, n6483, n6484, n6485, n6486, n6487, n6488,
         n6489, n6490, n6491, n6492, n6493, n6494, n6495, n6496, n6497, n6498,
         n6499, n6500, n6501, n6502, n6503, n6504, n6505, n6506, n6507, n6508,
         n6509, n6510, n6511, n6512, n6513, n6514, n6515, n6516, n6517, n6518,
         n6519, n6520, n6521, n6522, n6523, n6524, n6525, n6526, n6527, n6528,
         n6529, n6530, n6531, n6532, n6533, n6534, n6535, n6536, n6537, n6538,
         n6539, n6540, n6541, n6542, n6543, n6544, n6545, n6546, n6547, n6548,
         n6549, n6550, n6551, n6552, n6553, n6554, n6555, n6556, n6557, n6558,
         n6559, n6560, n6561, n6562, n6563, n6564, n6565, n6566, n6567, n6568,
         n6569, n6570, n6571, n6572, n6573, n6574, n6575, n6576, n6577, n6578,
         n6579, n6580, n6581, n6582, n6583, n6584, n6585, n6586, n6587, n6588,
         n6589, n6590, n6591, n6592, n6593, n6594, n6595, n6596, n6597, n6598,
         n6599, n6600, n6601, n6602, n6603, n6604, n6605, n6606, n6607, n6608,
         n6609, n6610, n6611, n6612, n6613, n6614, n6615, n6616, n6617, n6618,
         n6619, n6620, n6621, n6622, n6623, n6624, n6625, n6626, n6627, n6628,
         n6629, n6630, n6631, n6632, n6633, n6634, n6635, n6636, n6637, n6638,
         n6639, n6640, n6641, n6642, n6643, n6644, n6645, n6646, n6647, n6648,
         n6649, n6650, n6651, n6652, n6653, n6654, n6655, n6656, n6657, n6658,
         n6659, n6660, n6661, n6662, n6663, n6664, n6665, n6666, n6667, n6668,
         n6669, n6670, n6671, n6672, n6673, n6674, n6675, n6676, n6677, n6678,
         n6679, n6680, n6681, n6682, n6683, n6684, n6685, n6686, n6687, n6688,
         n6689, n6690, n6691, n6692, n6693, n6694, n6695, n6696, n6697, n6698,
         n6699, n6700, n6701, n6702, n6703, n6704, n6705, n6706, n6707, n6708,
         n6709, n6710, n6711, n6712, n6713, n6714, n6715, n6716, n6717, n6718,
         n6719, n6720, n6721, n6722, n6723, n6724, n6725, n6726, n6727, n6728,
         n6729, n6730, n6731, n6732, n6733, n6734, n6735, n6736, n6737, n6738,
         n6739, n6740, n6741, n6742, n6743, n6744, n6745, n6746, n6747, n6748,
         n6749, n6750, n6751, n6752, n6753, n6754, n6755, n6756, n6757, n6758,
         n6759, n6760, n6761, n6762, n6763, n6764, n6765, n6766, n6767, n6768,
         n6769, n6770, n6771, n6772, n6773, n6774, n6775, n6776, n6777, n6778,
         n6779, n6780, n6781, n6782, n6783, n6784, n6785, n6786, n6787, n6788,
         n6789, n6790, n6791, n6792, n6793, n6794, n6795, n6796, n6797, n6798,
         n6799, n6800, n6801, n6802, n6803, n6804, n6805, n6806, n6807, n6808,
         n6809, n6810, n6811, n6812, n6813, n6814, n6815, n6816, n6817, n6818,
         n6819, n6820, n6821, n6822, n6823, n6824, n6825, n6826, n6827, n6828,
         n6829, n6830, n6831, n6832, n6833, n6834, n6835, n6836, n6837, n6838,
         n6839, n6840, n6841, n6842, n6843, n6844, n6845, n6846, n6847, n6848,
         n6849, n6850, n6851, n6852, n6853, n6854, n6855, n6856, n6857, n6858,
         n6859, n6860, n6861, n6862, n6863, n6864, n6865, n6866, n6867, n6868,
         n6869, n6870, n6871, n6872, n6873, n6874, n6875, n6876, n6877, n6878,
         n6879, n6880, n6881, n6882, n6883, n6884, n6885, n6886, n6887, n6888,
         n6889, n6890, n6891, n6892, n6893, n6894, n6895, n6896, n6897, n6898,
         n6899, n6900, n6901, n6902, n6903, n6904, n6905, n6906, n6907, n6908,
         n6909, n6910, n6911, n6912, n6913, n6914, n6915, n6916, n6917, n6918,
         n6919, n6920, n6921, n6922, n6923, n6924, n6925, n6926, n6927, n6928,
         n6929, n6930, n6931, n6932, n6933, n6934, n6935, n6936, n6937, n6938,
         n6939, n6940, n6941, n6942, n6943, n6944, n6945, n6946, n6947, n6948,
         n6949, n6950, n6951, n6952, n6953, n6954, n6955, n6956, n6957, n6958,
         n6959, n6960, n6961, n6962, n6963, n6964, n6965, n6966, n6967, n6968,
         n6969, n6970, n6971, n6972, n6973, n6974, n6975, n6976, n6977, n6978,
         n6979, n6980, n6981, n6982, n6983, n6984, n6985, n6986, n6987, n6988,
         n6989, n6990, n6991, n6992, n6993, n6994, n6995, n6996, n6997, n6998,
         n6999, n7000, n7001, n7002, n7003, n7004, n7005, n7006, n7007, n7008,
         n7009, n7010, n7011, n7012, n7013, n7014, n7015, n7016, n7017, n7018,
         n7019, n7020, n7021, n7022, n7023, n7024, n7025, n7026, n7027, n7028,
         n7029, n7030, n7031, n7032, n7033, n7034, n7035, n7036, n7037, n7038,
         n7039, n7040, n7041, n7042, n7043, n7044, n7045, n7046, n7047, n7048,
         n7049, n7050, n7051, n7052, n7053, n7054, n7055, n7056, n7057, n7058,
         n7059, n7060, n7061, n7062, n7063, n7064, n7065, n7066, n7067, n7068,
         n7069, n7070, n7071, n7072, n7073, n7074, n7075, n7076, n7077, n7078,
         n7079, n7080, n7081, n7082, n7083, n7084, n7085, n7086, n7087, n7088,
         n7089, n7090, n7091, n7092, n7093, n7094, n7095, n7096, n7097, n7098,
         n7099, n7100, n7101, n7102, n7103, n7104, n7105, n7106, n7107, n7108,
         n7109, n7110, n7111, n7112, n7113, n7114, n7115, n7116, n7117, n7118,
         n7119, n7120, n7121, n7122, n7123, n7124, n7125, n7126, n7127, n7128,
         n7129, n7130, n7131, n7132, n7133, n7134, n7135, n7136, n7137, n7138,
         n7139, n7140, n7141, n7142, n7143, n7144, n7145, n7146, n7147, n7148,
         n7149, n7150, n7151, n7152, n7153, n7154, n7155, n7156, n7157, n7158,
         n7159, n7160, n7161, n7162, n7163, n7164, n7165, n7166, n7167, n7168,
         n7169, n7170, n7171, n7172, n7173, n7174, n7175, n7176, n7177, n7178,
         n7179, n7180, n7181, n7182, n7183, n7184, n7185, n7186, n7187, n7188,
         n7189, n7190, n7191, n7192, n7193, n7194, n7195, n7196, n7197, n7198,
         n7199, n7200, n7201, n7202, n7203, n7204, n7205, n7206, n7207, n7208,
         n7209, n7210, n7211, n7212, n7213, n7214, n7215, n7216, n7217, n7218,
         n7219, n7220, n7221, n7222, n7223, n7224, n7225, n7226, n7227, n7228,
         n7229, n7230, n7231, n7232, n7233, n7234, n7235, n7236, n7237, n7238,
         n7239, n7240, n7241, n7242, n7243, n7244, n7245, n7246, n7247, n7248,
         n7249, n7250, n7251, n7252, n7253, n7254, n7255, n7256, n7257, n7258,
         n7259, n7260, n7261, n7262, n7263, n7264, n7265, n7266, n7267, n7268,
         n7269, n7270, n7271, n7272, n7273, n7274, n7275, n7276, n7277, n7278,
         n7279, n7280, n7281, n7282, n7283, n7284, n7285, n7286, n7287, n7288,
         n7289, n7290, n7291, n7292, n7293, n7294, n7295, n7296, n7297, n7298,
         n7299, n7300, n7301, n7302, n7303, n7304, n7305, n7306, n7307, n7308,
         n7309, n7310, n7311, n7312, n7313, n7314, n7315, n7316, n7317, n7318,
         n7319, n7320, n7321, n7322, n7323, n7324, n7325, n7326, n7327, n7328,
         n7329, n7330, n7331, n7332, n7333, n7334, n7335, n7336, n7337, n7338,
         n7339, n7340, n7341, n7342, n7343, n7344, n7345, n7346, n7347, n7348,
         n7349, n7350, n7351, n7352, n7353, n7354, n7355, n7356, n7357, n7358,
         n7359, n7360, n7361, n7362, n7363, n7364, n7365, n7366, n7367, n7368,
         n7369, n7370, n7371, n7372, n7373, n7374, n7375, n7376, n7377, n7378,
         n7379, n7380, n7381, n7382, n7383, n7384, n7385, n7386, n7387, n7388,
         n7389, n7390, n7391, n7392, n7393, n7394, n7395, n7396, n7397, n7398,
         n7399, n7400, n7401, n7402, n7403, n7404, n7405, n7406, n7407, n7408,
         n7409, n7410, n7411, n7412, n7413, n7414, n7415, n7416, n7417, n7418,
         n7419, n7420, n7421, n7422, n7423, n7424, n7425, n7426, n7427, n7428,
         n7429, n7430, n7431, n7432, n7433, n7434, n7435, n7436, n7437, n7438,
         n7439, n7440, n7441, n7442, n7443, n7444, n7445, n7446, n7447, n7448,
         n7449, n7450, n7451, n7452, n7453, n7454, n7455, n7456, n7457, n7458,
         n7459, n7460, n7461, n7462, n7463, n7464, n7465, n7466, n7467, n7468,
         n7469, n7470, n7471, n7472, n7473, n7474, n7475, n7476, n7477, n7478,
         n7479, n7480, n7481, n7482, n7483, n7484, n7485, n7486, n7487, n7488,
         n7489, n7490, n7491, n7492, n7493, n7494, n7495, n7496, n7497, n7498,
         n7499, n7500, n7501, n7502, n7503, n7504, n7505, n7506, n7507, n7508,
         n7509, n7510, n7511, n7512, n7513, n7514, n7515, n7516, n7517, n7518,
         n7519, n7520, n7521, n7522, n7523, n7524, n7525, n7526, n7527, n7528,
         n7529, n7530, n7531, n7532, n7533, n7534, n7535, n7536, n7537, n7538,
         n7539, n7540, n7541, n7542, n7543, n7544, n7545, n7546, n7547, n7548,
         n7549, n7550, n7551, n7552, n7553, n7554, n7555, n7556, n7557, n7558,
         n7559, n7560, n7561, n7562, n7563, n7564, n7565, n7566, n7567, n7568,
         n7569, n7570, n7571, n7572, n7573, n7574, n7575, n7576, n7577, n7578,
         n7579, n7580, n7581, n7582, n7583, n7584, n7585, n7586, n7587, n7588,
         n7589, n7590, n7591, n7592, n7593, n7594, n7595, n7596, n7597, n7598,
         n7599, n7600, n7601, n7602, n7603, n7604, n7605, n7606, n7607, n7608,
         n7609, n7610, n7611, n7612, n7613, n7614, n7615, n7616, n7617, n7618,
         n7619, n7620, n7621, n7622, n7623, n7624, n7625, n7626, n7627, n7628,
         n7629, n7630, n7631, n7632, n7633, n7634, n7635, n7636, n7637, n7638,
         n7639, n7640, n7641, n7642, n7643, n7644, n7645, n7646, n7647, n7648,
         n7649, n7650, n7651, n7652, n7653, n7654, n7655, n7656, n7657, n7658,
         n7659, n7660, n7661, n7662, n7663, n7664, n7665, n7666, n7667, n7668,
         n7669, n7670, n7671, n7672, n7673, n7674, n7675, n7676, n7677, n7678,
         n7679, n7680, n7681, n7682, n7683, n7684, n7685, n7686, n7687, n7688,
         n7689, n7690, n7691, n7692, n7693, n7694, n7695, n7696, n7697, n7698,
         n7699, n7700, n7701, n7702, n7703, n7704, n7705, n7706, n7707, n7708,
         n7709, n7710, n7711, n7712, n7713, n7714, n7715, n7716, n7717, n7718,
         n7719, n7720, n7721, n7722, n7723, n7724, n7725, n7726, n7727, n7728,
         n7729, n7730, n7731, n7732, n7733, n7734, n7735, n7736, n7737, n7738,
         n7739, n7740, n7741, n7742, n7743, n7744, n7745, n7746, n7747, n7748,
         n7749, n7750, n7751, n7752, n7753, n7754, n7755, n7756, n7757, n7758,
         n7759, n7760, n7761, n7762, n7763, n7764, n7765, n7766, n7767, n7768,
         n7769, n7770, n7771, n7772, n7773, n7774, n7775, n7776, n7777, n7778,
         n7779, n7780, n7781, n7782, n7783, n7784, n7785, n7786, n7787, n7788,
         n7789, n7790, n7791, n7792, n7793, n7794, n7795, n7796, n7797, n7798,
         n7799, n7800, n7801, n7802, n7803, n7804, n7805, n7806, n7807, n7808,
         n7809, n7810, n7811, n7812, n7813, n7814, n7815, n7816, n7817, n7818,
         n7819, n7820, n7821, n7822, n7823, n7824, n7825, n7826, n7827, n7828,
         n7829, n7830, n7831, n7832, n7833, n7834, n7835, n7836, n7837, n7838,
         n7839, n7840, n7841, n7842, n7843, n7844, n7845, n7846, n7847, n7848,
         n7849, n7850, n7851, n7852, n7853, n7854, n7855, n7856, n7857, n7858,
         n7859, n7860, n7861, n7862, n7863, n7864, n7865, n7866, n7867, n7868,
         n7869, n7870, n7871, n7872, n7873, n7874, n7875, n7876, n7877, n7878,
         n7879, n7880, n7881, n7882, n7883, n7884, n7885, n7886, n7887, n7888,
         n7889, n7890, n7891, n7892, n7893, n7894, n7895, n7896, n7897, n7898,
         n7899, n7900, n7901, n7902, n7903, n7904, n7905, n7906, n7907, n7908,
         n7909, n7910, n7911, n7912, n7913, n7914, n7915, n7916, n7917, n7918,
         n7919, n7920, n7921, n7922, n7923, n7924, n7925, n7926, n7927, n7928,
         n7929, n7930, n7931, n7932, n7933, n7934, n7935, n7936, n7937, n7938,
         n7939, n7940, n7941, n7942, n7943, n7944, n7945, n7946, n7947, n7948,
         n7949, n7950, n7951, n7952, n7953, n7954, n7955, n7956, n7957, n7958,
         n7959, n7960, n7961, n7962, n7963, n7964, n7965, n7966, n7967, n7968,
         n7969, n7970, n7971, n7972, n7973, n7974, n7975, n7976, n7977, n7978,
         n7979, n7980, n7981, n7982, n7983, n7984, n7985, n7986, n7987, n7988,
         n7989, n7990, n7991, n7992, n7993, n7994, n7995, n7996, n7997, n7998,
         n7999, n8000, n8001, n8002, n8003, n8004, n8005, n8006, n8007, n8008,
         n8009, n8010, n8011, n8012, n8013, n8014, n8015, n8016, n8017, n8018,
         n8019, n8020, n8021, n8022, n8023, n8024, n8025, n8026, n8027, n8028,
         n8029, n8030, n8031, n8032, n8033, n8034, n8035, n8036, n8037, n8038,
         n8039, n8040, n8041, n8042, n8043, n8044, n8045, n8046, n8047, n8048,
         n8049, n8050, n8051, n8052, n8053, n8054, n8055, n8056, n8057, n8058,
         n8059, n8060, n8061, n8062, n8063, n8064, n8065, n8066, n8067, n8068,
         n8069, n8070, n8071, n8072, n8073, n8074, n8075, n8076, n8077, n8078,
         n8079, n8080, n8081, n8082, n8083, n8084, n8085, n8086, n8087, n8088,
         n8089, n8090, n8091, n8092, n8093, n8094, n8095, n8096, n8097, n8098,
         n8099, n8100, n8101, n8102, n8103, n8104, n8105, n8106, n8107, n8108,
         n8109, n8110, n8111, n8112, n8113, n8114, n8115, n8116, n8117, n8118,
         n8119, n8120, n8121, n8122, n8123, n8124, n8125, n8126, n8127, n8128,
         n8129, n8130, n8131, n8132, n8133, n8134, n8135, n8136, n8137, n8138,
         n8139, n8140, n8141, n8142, n8143, n8144, n8145, n8146, n8147, n8148,
         n8149, n8150, n8151, n8152, n8153, n8154, n8155, n8156, n8157, n8158,
         n8159, n8160, n8161, n8162, n8163, n8164, n8165, n8166, n8167, n8168,
         n8169, n8170, n8171, n8172, n8173, n8174, n8175, n8176, n8177, n8178,
         n8179, n8180, n8181, n8182, n8183, n8184, n8185, n8186, n8187, n8188,
         n8189, n8190, n8191, n8192, n8193, n8194, n8195, n8196, n8197, n8198,
         n8199, n8200, n8201, n8202, n8203, n8204, n8205, n8206, n8207, n8208,
         n8209, n8210, n8211, n8212, n8213, n8214, n8215, n8216, n8217, n8218,
         n8219, n8220, n8221, n8222, n8223, n8224, n8225, n8226, n8227, n8228,
         n8229, n8230, n8231, n8232, n8233, n8234, n8235, n8236, n8237, n8238,
         n8239, n8240, n8241, n8242, n8243, n8244, n8245, n8246, n8247, n8248,
         n8249, n8250, n8251, n8252, n8253, n8254, n8255, n8256, n8257, n8258,
         n8259, n8260, n8261, n8262, n8263, n8264, n8265, n8266, n8267, n8268,
         n8269, n8270, n8271, n8272, n8273, n8274, n8275, n8276, n8277, n8278,
         n8279, n8280, n8281, n8282, n8283, n8284, n8285, n8286, n8287, n8288,
         n8289, n8290, n8291, n8292, n8293, n8294, n8295, n8296, n8297, n8298,
         n8299, n8300, n8301, n8302, n8303, n8304, n8305, n8306, n8307, n8308,
         n8309, n8310, n8311, n8312, n8313, n8314, n8315, n8316, n8317, n8318,
         n8319, n8320, n8321, n8322, n8323, n8324, n8325, n8326, n8327, n8328,
         n8329, n8330, n8331, n8332, n8333, n8334, n8335, n8336, n8337, n8338,
         n8339, n8340, n8341, n8342, n8343, n8344, n8345, n8346, n8347, n8348,
         n8349, n8350, n8351, n8352, n8353, n8354, n8355, n8356, n8357, n8358,
         n8359, n8360, n8361, n8362, n8363, n8364, n8365, n8366, n8367, n8368,
         n8369, n8370, n8371, n8372, n8373, n8374, n8375, n8376, n8377, n8378,
         n8379, n8380, n8381, n8382, n8383, n8384, n8385, n8386, n8387, n8388,
         n8389, n8390, n8391, n8392, n8393, n8394, n8395, n8396, n8397, n8398,
         n8399, n8400, n8401, n8402, n8403, n8404, n8405, n8406, n8407, n8408,
         n8409, n8410, n8411, n8412, n8413, n8414, n8415, n8416, n8417, n8418,
         n8419, n8420, n8421, n8422, n8423, n8424, n8425, n8426, n8427, n8428,
         n8429, n8430, n8431, n8432, n8433, n8434, n8435, n8436, n8437, n8438,
         n8439, n8440, n8441, n8442, n8443, n8444, n8445, n8446, n8447, n8448,
         n8449, n8450, n8451, n8452, n8453, n8454, n8455, n8456, n8457, n8458,
         n8459, n8460, n8461, n8462, n8463, n8464, n8465, n8466, n8467, n8468,
         n8469, n8470, n8471, n8472, n8473, n8474, n8475, n8476, n8477, n8478,
         n8479, n8480, n8481, n8482, n8483, n8484, n8485, n8486, n8487, n8488,
         n8489, n8490, n8491, n8492, n8493, n8494, n8495, n8496, n8497, n8498,
         n8499, n8500, n8501, n8502, n8503, n8504, n8505, n8506, n8507, n8508,
         n8509, n8510, n8511, n8512, n8513, n8514, n8515, n8516, n8517, n8518,
         n8519, n8520, n8521, n8522, n8523, n8524, n8525, n8526, n8527, n8528,
         n8529, n8530, n8531, n8532, n8533, n8534, n8535, n8536, n8537, n8538,
         n8539, n8540, n8541, n8542, n8543, n8544, n8545, n8546, n8547, n8548,
         n8549, n8550, n8551, n8552, n8553, n8554, n8555, n8556, n8557, n8558,
         n8559, n8560, n8561, n8562, n8563, n8564, n8565, n8566, n8567, n8568,
         n8569, n8570, n8571, n8572, n8573, n8574, n8575, n8576, n8577, n8578,
         n8579, n8580, n8581, n8582, n8583, n8584, n8585, n8586, n8587, n8588,
         n8589, n8590, n8591, n8592, n8593, n8594, n8595, n8596, n8597, n8598,
         n8599, n8600, n8601, n8602, n8603, n8604, n8605, n8606, n8607, n8608,
         n8609, n8610, n8611, n8612, n8613, n8614, n8615, n8616, n8617, n8618,
         n8619, n8620, n8621, n8622, n8623, n8624, n8625, n8626, n8627, n8628,
         n8629, n8630, n8631, n8632, n8633, n8634, n8635, n8636, n8637, n8638,
         n8639, n8640, n8641, n8642, n8643, n8644, n8645, n8646, n8647, n8648,
         n8649, n8650, n8651, n8652, n8653, n8654, n8655, n8656, n8657, n8658,
         n8659, n8660, n8661, n8662, n8663, n8664, n8665, n8666, n8667, n8668,
         n8669, n8670, n8671, n8672, n8673, n8674, n8675, n8676, n8677, n8678,
         n8679, n8680, n8681, n8682, n8683, n8684, n8685, n8686, n8687, n8688,
         n8689, n8690, n8691, n8692, n8693, n8694, n8695, n8696, n8697, n8698,
         n8699, n8700, n8701, n8702, n8703, n8704, n8705, n8706, n8707, n8708,
         n8709, n8710, n8711, n8712, n8713, n8714, n8715, n8716, n8717, n8718,
         n8719, n8720, n8721, n8722, n8723, n8724, n8725, n8726, n8727, n8728,
         n8729, n8730, n8731, n8732, n8733, n8734, n8735, n8736, n8737, n8738,
         n8739, n8740, n8741, n8742, n8743, n8744, n8745, n8746, n8747, n8748,
         n8749, n8750, n8751, n8752, n8753, n8754, n8755, n8756, n8757, n8758,
         n8759, n8760, n8761, n8762, n8763, n8764, n8765, n8766, n8767, n8768,
         n8769, n8770, n8771, n8772, n8773, n8774, n8775, n8776, n8777, n8778,
         n8779, n8780, n8781, n8782, n8783, n8784, n8785, n8786, n8787, n8788,
         n8789, n8790, n8791, n8792, n8793, n8794, n8795, n8796, n8797, n8798,
         n8799, n8800, n8801, n8802, n8803, n8804, n8805, n8806, n8807, n8808,
         n8809, n8810, n8811, n8812, n8813, n8814, n8815, n8816, n8817, n8818,
         n8819, n8820, n8821, n8822, n8823, n8824, n8825, n8826, n8827, n8828,
         n8829, n8830, n8831, n8832, n8833, n8834, n8835, n8836, n8837, n8838,
         n8839, n8840, n8841, n8842, n8843, n8844, n8845, n8846, n8847, n8848,
         n8849, n8850, n8851, n8852, n8853, n8854, n8855, n8856, n8857, n8858,
         n8859, n8860, n8861, n8862, n8863, n8864, n8865, n8866, n8867, n8868,
         n8869, n8870, n8871, n8872, n8873, n8874, n8875, n8876, n8877, n8878,
         n8879, n8880, n8881, n8882, n8883, n8884, n8885, n8886, n8887, n8888,
         n8889, n8890, n8891, n8892, n8893, n8894, n8895, n8896, n8897, n8898,
         n8899, n8900, n8901, n8902, n8903, n8904, n8905, n8906, n8907, n8908,
         n8909, n8910, n8911, n8912, n8913, n8914, n8915, n8916, n8917, n8918,
         n8919, n8920, n8921, n8922, n8923, n8924, n8925, n8926, n8927, n8928,
         n8929, n8930, n8931, n8932, n8933, n8934, n8935, n8936, n8937, n8938,
         n8939, n8940, n8941, n8942, n8943, n8944, n8945, n8946, n8947, n8948,
         n8949, n8950, n8951, n8952, n8953, n8954, n8955, n8956, n8957, n8958,
         n8959, n8960, n8961, n8962, n8963, n8964, n8965, n8966, n8967, n8968,
         n8969, n8970, n8971, n8972, n8973, n8974, n8975, n8976, n8977, n8978,
         n8979, n8980, n8981, n8982, n8983, n8984, n8985, n8986, n8987, n8988,
         n8989, n8990, n8991, n8992, n8993, n8994, n8995, n8996, n8997, n8998,
         n8999, n9000, n9001, n9002, n9003, n9004, n9005, n9006, n9007, n9008,
         n9009, n9010, n9011, n9012, n9013, n9014, n9015, n9016, n9017, n9018,
         n9019, n9020, n9021, n9022, n9023, n9024, n9025, n9026, n9027, n9028,
         n9029, n9030, n9031, n9032, n9033, n9034, n9035, n9036, n9037, n9038,
         n9039, n9040, n9041, n9042, n9043, n9044, n9045, n9046, n9047, n9048,
         n9049, n9050, n9051, n9052, n9053, n9054, n9055, n9056, n9057, n9058,
         n9059, n9060, n9061, n9062, n9063, n9064, n9065, n9066, n9067, n9068,
         n9069, n9070, n9071, n9072, n9073, n9074, n9075, n9076, n9077, n9078,
         n9079, n9080, n9081, n9082, n9083, n9084, n9085, n9086, n9087, n9088,
         n9089, n9090, n9091, n9092, n9093, n9094, n9095, n9096, n9097, n9098,
         n9099, n9100, n9101, n9102, n9103, n9104, n9105, n9106, n9107, n9108,
         n9109, n9110, n9111, n9112, n9113, n9114, n9115, n9116, n9117, n9118,
         n9119, n9120, n9121, n9122, n9123, n9124, n9125, n9126, n9127, n9128,
         n9129, n9130, n9131, n9132, n9133, n9134, n9135, n9136, n9137, n9138,
         n9139, n9140, n9141, n9142, n9143, n9144, n9145, n9146, n9147, n9148,
         n9149, n9150, n9151, n9152, n9153, n9154, n9155, n9156, n9157, n9158,
         n9159, n9160, n9161, n9162, n9163, n9164, n9165, n9166, n9167, n9168,
         n9169, n9170, n9171, n9172, n9173, n9174, n9175, n9176, n9177, n9178,
         n9179, n9180, n9181, n9182, n9183, n9184, n9185, n9186, n9187, n9188,
         n9189, n9190, n9191, n9192, n9193, n9194, n9195, n9196, n9197, n9198,
         n9199, n9200, n9201, n9202, n9203, n9204, n9205, n9206, n9207, n9208,
         n9209, n9210, n9211, n9212, n9213, n9214, n9215, n9216, n9217, n9218,
         n9219, n9220, n9221, n9222, n9223, n9224, n9225, n9226, n9227, n9228,
         n9229, n9230, n9231, n9232, n9233, n9234, n9235, n9236, n9237, n9238,
         n9239, n9240, n9241, n9242, n9243, n9244, n9245, n9246, n9247, n9248,
         n9249, n9250, n9251, n9252, n9253, n9254, n9255, n9256, n9257, n9258,
         n9259, n9260, n9261, n9262, n9263, n9264, n9265, n9266, n9267, n9268,
         n9269, n9270, n9271, n9272, n9273, n9274, n9275, n9276, n9277, n9278,
         n9279, n9280, n9281, n9282, n9283, n9284, n9285, n9286, n9287, n9288,
         n9289, n9290, n9291, n9292, n9293, n9294, n9295, n9296, n9297, n9298,
         n9299, n9300, n9301, n9302, n9303, n9304, n9305, n9306, n9307, n9308,
         n9309, n9310, n9311, n9312, n9313, n9314, n9315, n9316, n9317, n9318,
         n9319, n9320, n9321, n9322, n9323, n9324, n9325, n9326, n9327, n9328,
         n9329, n9330, n9331, n9332, n9333, n9334, n9335, n9336, n9337, n9338,
         n9339, n9340, n9341, n9342, n9343, n9344, n9345, n9346, n9347, n9348,
         n9349, n9350, n9351, n9352, n9353, n9354, n9355, n9356, n9357, n9358,
         n9359, n9360, n9361, n9362, n9363, n9364, n9365, n9366, n9367, n9368,
         n9369, n9370, n9371, n9372, n9373, n9374, n9375, n9376, n9377, n9378,
         n9379, n9380, n9381, n9382, n9383, n9384, n9385, n9386, n9387, n9388,
         n9389, n9390, n9391, n9392, n9393, n9394, n9395, n9396, n9397, n9398,
         n9399, n9400, n9401, n9402, n9403, n9404, n9405, n9406, n9407, n9408,
         n9409, n9410, n9411, n9412, n9413, n9414, n9415, n9416, n9417, n9418,
         n9419, n9420, n9421, n9422, n9423, n9424, n9425, n9426, n9427, n9428,
         n9429, n9430, n9431, n9432, n9433, n9434, n9435, n9436, n9437, n9438,
         n9439, n9440, n9441, n9442, n9443, n9444, n9445, n9446, n9447, n9448,
         n9449, n9450, n9451, n9452, n9453, n9454, n9455, n9456, n9457, n9458,
         n9459, n9460, n9461, n9462, n9463, n9464, n9465, n9466, n9467, n9468,
         n9469, n9470, n9471, n9472, n9473, n9474, n9475, n9476, n9477, n9478,
         n9479, n9480, n9481, n9482, n9483, n9484, n9485, n9486, n9487, n9488,
         n9489, n9490, n9491, n9492, n9493, n9494, n9495, n9496, n9497, n9498,
         n9499, n9500, n9501, n9502, n9503, n9504, n9505, n9506, n9507, n9508,
         n9509, n9510, n9511, n9512, n9513, n9514, n9515, n9516, n9517, n9518,
         n9519, n9520, n9521, n9522, n9523, n9524, n9525, n9526, n9527, n9528,
         n9529, n9530, n9531, n9532, n9533, n9534, n9535, n9536, n9537, n9538,
         n9539, n9540, n9541, n9542, n9543, n9544, n9545, n9546, n9547, n9548,
         n9549, n9550, n9551, n9552, n9553, n9554, n9555, n9556, n9557, n9558,
         n9559, n9560, n9561, n9562, n9563, n9564, n9565, n9566, n9567, n9568,
         n9569, n9570, n9571, n9572, n9573, n9574, n9575, n9576, n9577, n9578,
         n9579, n9580, n9581, n9582, n9583, n9584, n9585, n9586, n9587, n9588,
         n9589, n9590, n9591, n9592, n9593, n9594, n9595, n9596, n9597, n9598,
         n9599, n9600, n9601, n9602, n9603, n9604, n9605, n9606, n9607, n9608,
         n9609, n9610, n9611, n9612, n9613, n9614, n9615, n9616, n9617, n9618,
         n9619, n9620, n9621, n9622, n9623, n9624, n9625, n9626, n9627, n9628,
         n9629, n9630, n9631, n9632, n9633, n9634, n9635, n9636, n9637, n9638,
         n9639, n9640, n9641, n9642, n9643, n9644, n9645, n9646, n9647, n9648,
         n9649, n9650, n9651, n9652, n9653, n9654, n9655, n9656, n9657, n9658,
         n9659, n9660, n9661, n9662, n9663, n9664, n9665, n9666, n9667, n9668,
         n9669, n9670, n9671, n9672, n9673, n9674, n9675, n9676, n9677, n9678,
         n9679, n9680, n9681, n9682, n9683, n9684, n9685, n9686, n9687, n9688,
         n9689, n9690, n9691, n9692, n9693, n9694, n9695, n9696, n9697, n9698,
         n9699, n9700, n9701, n9702, n9703, n9704, n9705, n9706, n9707, n9708,
         n9709, n9710, n9711, n9712, n9713, n9714, n9715, n9716, n9717, n9718,
         n9719, n9720, n9721, n9722, n9723, n9724, n9725, n9726, n9727, n9728,
         n9729, n9730, n9731, n9732, n9733, n9734, n9735, n9736, n9737, n9738,
         n9739, n9740, n9741, n9742, n9743, n9744, n9745, n9746, n9747, n9748,
         n9749, n9750, n9751, n9752, n9753, n9754, n9755, n9756, n9757, n9758,
         n9759, n9760, n9761, n9762, n9763, n9764, n9765, n9766, n9767, n9768,
         n9769, n9770, n9771, n9772, n9773, n9774, n9775, n9776, n9777, n9778,
         n9779, n9780, n9781, n9782, n9783, n9784, n9785, n9786, n9787, n9788,
         n9789, n9790, n9791, n9792, n9793, n9794, n9795, n9796, n9797, n9798,
         n9799, n9800, n9801, n9802, n9803, n9804, n9805, n9806, n9807, n9808,
         n9809, n9810, n9811, n9812, n9813, n9814, n9815, n9816, n9817, n9818,
         n9819, n9820, n9821, n9822, n9823, n9824, n9825, n9826, n9827, n9828,
         n9829, n9830, n9831, n9832, n9833, n9834, n9835, n9836, n9837, n9838,
         n9839, n9840, n9841, n9842, n9843, n9844, n9845, n9846, n9847, n9848,
         n9849, n9850, n9851, n9852, n9853, n9854, n9855, n9856, n9857, n9858,
         n9859, n9860, n9861, n9862, n9863, n9864, n9865, n9866, n9867, n9868,
         n9869, n9870, n9871, n9872, n9873, n9874, n9875, n9876, n9877, n9878,
         n9879, n9880, n9881, n9882, n9883, n9884, n9885, n9886, n9887, n9888,
         n9889, n9890, n9891, n9892, n9893, n9894, n9895, n9896, n9897, n9898,
         n9899, n9900, n9901, n9902, n9903, n9904, n9905, n9906, n9907, n9908,
         n9909, n9910, n9911, n9912, n9913, n9914, n9915, n9916, n9917, n9918,
         n9919, n9920, n9921, n9922, n9923, n9924, n9925, n9926, n9927, n9928,
         n9929, n9930, n9931, n9932, n9933, n9934, n9935, n9936, n9937, n9938,
         n9939, n9940, n9941, n9942, n9943, n9944, n9945, n9946, n9947, n9948,
         n9949, n9950, n9951, n9952, n9953, n9954, n9955, n9956, n9957, n9958,
         n9959, n9960, n9961, n9962, n9963, n9964, n9965, n9966, n9967, n9968,
         n9969, n9970, n9971, n9972, n9973, n9974, n9975, n9976, n9977, n9978,
         n9979, n9980, n9981, n9982, n9983, n9984, n9985, n9986, n9987, n9988,
         n9989, n9990, n9991, n9992, n9993, n9994, n9995, n9996, n9997, n9998,
         n9999, n10000, n10001, n10002, n10003, n10004, n10005, n10006, n10007,
         n10008, n10009, n10010, n10011, n10012, n10013, n10014, n10015,
         n10016, n10017, n10018, n10019, n10020, n10021, n10022, n10023,
         n10024, n10025, n10026, n10027, n10028, n10029, n10030, n10031,
         n10032, n10033, n10034, n10035, n10036, n10037, n10038, n10039,
         n10040, n10041, n10042, n10043, n10044, n10045, n10046, n10047,
         n10048, n10049, n10050, n10051, n10052, n10053, n10054, n10055,
         n10056, n10057, n10058, n10059, n10060, n10061, n10062, n10063,
         n10064, n10065, n10066, n10067, n10068, n10069, n10070, n10071,
         n10072, n10073, n10074, n10075, n10076, n10077, n10078, n10079,
         n10080, n10081, n10082, n10083, n10084, n10085, n10086, n10087,
         n10088, n10089, n10090, n10091, n10092, n10093, n10094, n10095,
         n10096, n10097, n10098, n10099, n10100, n10101, n10102, n10103,
         n10104, n10105, n10106, n10107, n10108, n10109, n10110, n10111,
         n10112, n10113, n10114, n10115, n10116, n10117, n10118, n10119,
         n10120, n10121, n10122, n10123, n10124, n10125, n10126, n10127,
         n10128, n10129, n10130, n10131, n10132, n10133, n10134, n10135,
         n10136, n10137, n10138, n10139, n10140, n10141, n10142, n10143,
         n10144, n10145, n10146, n10147, n10148, n10149, n10150, n10151,
         n10152, n10153, n10154, n10155, n10156, n10157, n10158, n10159,
         n10160, n10161, n10162, n10163, n10164, n10165, n10166, n10167,
         n10168, n10169, n10170, n10171, n10172, n10173, n10174, n10175,
         n10176, n10177, n10178, n10179, n10180, n10181, n10182, n10183,
         n10184, n10185, n10186, n10187, n10188, n10189, n10190, n10191,
         n10192, n10193, n10194, n10195, n10196, n10197, n10198, n10199,
         n10200, n10201, n10202, n10203, n10204, n10205, n10206, n10207,
         n10208, n10209, n10210, n10211, n10212, n10213, n10214, n10215,
         n10216, n10217, n10218, n10219, n10220, n10221, n10222, n10223,
         n10224, n10225, n10226, n10227, n10228, n10229, n10230, n10231,
         n10232, n10233, n10234, n10235, n10236, n10237, n10238, n10239,
         n10240, n10241, n10242, n10243, n10244, n10245, n10246, n10247,
         n10248, n10249, n10250, n10251, n10252, n10253, n10254, n10255,
         n10256, n10257, n10258, n10259, n10260, n10261, n10262, n10263,
         n10264, n10265, n10266, n10267, n10268, n10269, n10270, n10271,
         n10272, n10273, n10274, n10275, n10276, n10277, n10278, n10279,
         n10280, n10281, n10282, n10283, n10284, n10285, n10286, n10287,
         n10288, n10289, n10290, n10291, n10292, n10293, n10294, n10295,
         n10296, n10297, n10298, n10299, n10300, n10301, n10302, n10303,
         n10304, n10305, n10306, n10307, n10308, n10309, n10310, n10311,
         n10312, n10313, n10314, n10315, n10316, n10317, n10318, n10319,
         n10320, n10321, n10322, n10323, n10324, n10325, n10326, n10327,
         n10328, n10329, n10330, n10331, n10332, n10333, n10334, n10335,
         n10336, n10337, n10338, n10339, n10340, n10341, n10342, n10343,
         n10344, n10345, n10346, n10347, n10348, n10349, n10350, n10351,
         n10352, n10353, n10354, n10355, n10356, n10357, n10358, n10359,
         n10360, n10361, n10362, n10363, n10364, n10365, n10366, n10367,
         n10368, n10369, n10370, n10371, n10372, n10373, n10374, n10375,
         n10376, n10377, n10378, n10379, n10380, n10381, n10382, n10383,
         n10384, n10385, n10386, n10387, n10388, n10389, n10390, n10391,
         n10392, n10393, n10394, n10395, n10396, n10397, n10398, n10399,
         n10400, n10401, n10402, n10403, n10404, n10405, n10406, n10407,
         n10408, n10409, n10410, n10411, n10412, n10413, n10414, n10415,
         n10416, n10417, n10418, n10419, n10420, n10421, n10422, n10423,
         n10424, n10425, n10426, n10427, n10428, n10429, n10430, n10431,
         n10432, n10433, n10434, n10435, n10436, n10437, n10438, n10439,
         n10440, n10441, n10442, n10443, n10444, n10445, n10446, n10447,
         n10448, n10449, n10450, n10451, n10452, n10453, n10454, n10455,
         n10456, n10457, n10458, n10459, n10460, n10461, n10462, n10463,
         n10464, n10465, n10466, n10467, n10468, n10469, n10470, n10471,
         n10472, n10473, n10474, n10475, n10476, n10477, n10478, n10479,
         n10480, n10481, n10482, n10483, n10484, n10485, n10486, n10487,
         n10488, n10489, n10490, n10491, n10492, n10493, n10494, n10495,
         n10496, n10497, n10498, n10499, n10500, n10501, n10502, n10503,
         n10504, n10505, n10506, n10507, n10508, n10509, n10510, n10511,
         n10512, n10513, n10514, n10515, n10516, n10517, n10518, n10519,
         n10520, n10521, n10522, n10523, n10524, n10525, n10526, n10527,
         n10528, n10529, n10530, n10531, n10532, n10533, n10534, n10535,
         n10536, n10537, n10538, n10539, n10540, n10541, n10542, n10543,
         n10544, n10545, n10546, n10547, n10548, n10549, n10550, n10551,
         n10552, n10553, n10554, n10555, n10556, n10557, n10558, n10559,
         n10560, n10561, n10562, n10563, n10564, n10565, n10566, n10567,
         n10568, n10569, n10570, n10571, n10572, n10573, n10574, n10575,
         n10576, n10577, n10578, n10579, n10580, n10581, n10582, n10583,
         n10584, n10585, n10586, n10587, n10588, n10589, n10590, n10591,
         n10592, n10593, n10594, n10595, n10596, n10597, n10598, n10599,
         n10600, n10601, n10602, n10603, n10604, n10605, n10606, n10607,
         n10608, n10609, n10610, n10611, n10612, n10613, n10614, n10615,
         n10616, n10617, n10618, n10619, n10620, n10621, n10622, n10623,
         n10624, n10625, n10626, n10627, n10628, n10629, n10630, n10631,
         n10632, n10633, n10634, n10635, n10636, n10637, n10638, n10639,
         n10640, n10641, n10642, n10643, n10644, n10645, n10646, n10647,
         n10648, n10649, n10650, n10651, n10652, n10653, n10654, n10655,
         n10656, n10657, n10658, n10659, n10660, n10661, n10662, n10663,
         n10664, n10665, n10666, n10667, n10668, n10669, n10670, n10671,
         n10672, n10673, n10674, n10675, n10676, n10677, n10678, n10679,
         n10680, n10681, n10682, n10683, n10684, n10685, n10686, n10687,
         n10688, n10689, n10690, n10691, n10692, n10693, n10694, n10695,
         n10696, n10697, n10698, n10699, n10700, n10701, n10702, n10703,
         n10704, n10705, n10706, n10707, n10708, n10709, n10710, n10711,
         n10712, n10713, n10714, n10715, n10716, n10717, n10718, n10719,
         n10720, n10721, n10722, n10723, n10724, n10725, n10726, n10727,
         n10728, n10729, n10730, n10731, n10732, n10733, n10734, n10735,
         n10736, n10737, n10738, n10739, n10740, n10741, n10742, n10743,
         n10744, n10745, n10746, n10747, n10748, n10749, n10750, n10751,
         n10752, n10753, n10754, n10755, n10756, n10757, n10758, n10759,
         n10760, n10761, n10762, n10763, n10764, n10765, n10766, n10767,
         n10768, n10769, n10770, n10771, n10772, n10773, n10774, n10775,
         n10776, n10777, n10778, n10779, n10780, n10781, n10782, n10783,
         n10784, n10785, n10786, n10787, n10788, n10789, n10790, n10791,
         n10792, n10793, n10794, n10795, n10796, n10797, n10798, n10799,
         n10800, n10801, n10802, n10803, n10804, n10805, n10806, n10807,
         n10808, n10809, n10810, n10811, n10812, n10813, n10814, n10815,
         n10816, n10817, n10818, n10819, n10820, n10821, n10822, n10823,
         n10824, n10825, n10826, n10827, n10828, n10829, n10830, n10831,
         n10832, n10833, n10834, n10835, n10836, n10837, n10838, n10839,
         n10840, n10841, n10842, n10843, n10844, n10845, n10846, n10847,
         n10848, n10849, n10850, n10851, n10852, n10853, n10854, n10855,
         n10856, n10857, n10858, n10859, n10860, n10861, n10862, n10863,
         n10864, n10865, n10866, n10867, n10868, n10869, n10870, n10871,
         n10872, n10873, n10874, n10875, n10876, n10877, n10878, n10879,
         n10880, n10881, n10882, n10883, n10884, n10885, n10886, n10887,
         n10888, n10889, n10890, n10891, n10892, n10893, n10894, n10895,
         n10896, n10897, n10898, n10899, n10900, n10901, n10902, n10903,
         n10904, n10905, n10906, n10907, n10908, n10909, n10910, n10911,
         n10912, n10913, n10914, n10915, n10916, n10917, n10918, n10919,
         n10920, n10921, n10922, n10923, n10924, n10925, n10926, n10927,
         n10928, n10929, n10930, n10931, n10932, n10933, n10934, n10935,
         n10936, n10937, n10938, n10939, n10940, n10941, n10942, n10943,
         n10944, n10945, n10946, n10947, n10948, n10949, n10950, n10951,
         n10952, n10953, n10954, n10955, n10956, n10957, n10958, n10959,
         n10960, n10961, n10962, n10963, n10964, n10965, n10966, n10967,
         n10968, n10969, n10970, n10971, n10972, n10973, n10974, n10975,
         n10976, n10977, n10978, n10979, n10980, n10981, n10982, n10983,
         n10984, n10985, n10986, n10987, n10988, n10989, n10990, n10991,
         n10992, n10993, n10994, n10995, n10996, n10997, n10998, n10999,
         n11000, n11001, n11002, n11003, n11004, n11005, n11006, n11007,
         n11008, n11009, n11010, n11011, n11012, n11013, n11014, n11015,
         n11016, n11017, n11018, n11019, n11020, n11021, n11022, n11023,
         n11024, n11025, n11026, n11027, n11028, n11029, n11030, n11031,
         n11032, n11033, n11034, n11035, n11036, n11037, n11038, n11039,
         n11040, n11041, n11042, n11043, n11044, n11045, n11046, n11047,
         n11048, n11049, n11050, n11051, n11052, n11053, n11054, n11055,
         n11056, n11057, n11058, n11059, n11060, n11061, n11062, n11063,
         n11064, n11065, n11066, n11067, n11068, n11069, n11070, n11071,
         n11072, n11073, n11074, n11075, n11076, n11077, n11078, n11079,
         n11080, n11081, n11082, n11083, n11084, n11085, n11086, n11087,
         n11088, n11089, n11090, n11091, n11092, n11093, n11094, n11095,
         n11096, n11097, n11098, n11099, n11100, n11101, n11102, n11103,
         n11104, n11105, n11106, n11107, n11108, n11109, n11110, n11111,
         n11112, n11113, n11114, n11115, n11116, n11117, n11118, n11119,
         n11120, n11121, n11122, n11123, n11124, n11125, n11126, n11127,
         n11128, n11129, n11130, n11131, n11132, n11133, n11134, n11135,
         n11136, n11137, n11138, n11139, n11140, n11141, n11142, n11143,
         n11144, n11145, n11146, n11147, n11148, n11149, n11150, n11151,
         n11152, n11153, n11154, n11155, n11156, n11157, n11158, n11159,
         n11160, n11161, n11162, n11163, n11164, n11165, n11166, n11167,
         n11168, n11169, n11170, n11171, n11172, n11173, n11174, n11175,
         n11176, n11177, n11178, n11179, n11180, n11181, n11182, n11183,
         n11184, n11185, n11186, n11187, n11188, n11189, n11190, n11191,
         n11192, n11193, n11194, n11195, n11196, n11197, n11198, n11199,
         n11200, n11201, n11202, n11203, n11204, n11205, n11206, n11207,
         n11208, n11209, n11210, n11211, n11212, n11213, n11214, n11215,
         n11216, n11217, n11218, n11219, n11220, n11221, n11222, n11223,
         n11224, n11225, n11226, n11227, n11228, n11229, n11230, n11231,
         n11232, n11233, n11234, n11235, n11236, n11237, n11238, n11239,
         n11240, n11241, n11242, n11243, n11244, n11245, n11246, n11247,
         n11248, n11249, n11250, n11251, n11252, n11253, n11254, n11255,
         n11256, n11257, n11258, n11259, n11260, n11261, n11262, n11263,
         n11264, n11265, n11266, n11267, n11268, n11269, n11270, n11271,
         n11272, n11273, n11274, n11275, n11276, n11277, n11278, n11279,
         n11280, n11281, n11282, n11283, n11284, n11285, n11286, n11287,
         n11288, n11289, n11290, n11291, n11292, n11293, n11294, n11295,
         n11296, n11297, n11298, n11299, n11300, n11301, n11302, n11303,
         n11304, n11305, n11306, n11307, n11308, n11309, n11310, n11311,
         n11312, n11313, n11314, n11315, n11316, n11317, n11318, n11319,
         n11320, n11321, n11322, n11323, n11324, n11325, n11326, n11327,
         n11328, n11329, n11330, n11331, n11332, n11333, n11334, n11335,
         n11336, n11337, n11338, n11339, n11340, n11341, n11342, n11343,
         n11344, n11345, n11346, n11347, n11348, n11349, n11350, n11351,
         n11352, n11353, n11354, n11355, n11356, n11357, n11358, n11359,
         n11360, n11361, n11362, n11363, n11364, n11365, n11366, n11367,
         n11368, n11369, n11370, n11371, n11372, n11373, n11374, n11375,
         n11376, n11377, n11378, n11379, n11380, n11381, n11382, n11383,
         n11384, n11385, n11386, n11387, n11388, n11389, n11390, n11391,
         n11392, n11393, n11394, n11395, n11396, n11397, n11398, n11399,
         n11400, n11401, n11402, n11403, n11404, n11405, n11406, n11407,
         n11408, n11409, n11410, n11411, n11412, n11413, n11414, n11415,
         n11416, n11417, n11418, n11419, n11420, n11421, n11422, n11423,
         n11424, n11425, n11426, n11427, n11428, n11429, n11430, n11431,
         n11432, n11433, n11434, n11435, n11436, n11437, n11438, n11439,
         n11440, n11441, n11442, n11443, n11444, n11445, n11446, n11447,
         n11448, n11449, n11450, n11451, n11452, n11453, n11454, n11455,
         n11456, n11457, n11458, n11459, n11460, n11461, n11462, n11463,
         n11464, n11465, n11466, n11467, n11468, n11469, n11470, n11471,
         n11472, n11473, n11474, n11475, n11476, n11477, n11478, n11479,
         n11480, n11481, n11482, n11483, n11484, n11485, n11486, n11487,
         n11488, n11489, n11490, n11491, n11492, n11493, n11494, n11495,
         n11496, n11497, n11498, n11499, n11500, n11501, n11502, n11503,
         n11504, n11505, n11506, n11507, n11508, n11509, n11510, n11511,
         n11512, n11513, n11514, n11515, n11516, n11517, n11518, n11519,
         n11520, n11521, n11522, n11523, n11524, n11525, n11526, n11527,
         n11528, n11529, n11530, n11531, n11532, n11533, n11534, n11535,
         n11536, n11537, n11538, n11539, n11540, n11541, n11542, n11543,
         n11544, n11545, n11546, n11547, n11548, n11549, n11550, n11551,
         n11552, n11553, n11554, n11555, n11556, n11557, n11558, n11559,
         n11560, n11561, n11562, n11563, n11564, n11565, n11566, n11567,
         n11568, n11569, n11570, n11571, n11572, n11573, n11574, n11575,
         n11576, n11577, n11578, n11579, n11580, n11581, n11582, n11583,
         n11584, n11585, n11586, n11587, n11588, n11589, n11590, n11591,
         n11592, n11593, n11594, n11595, n11596, n11597, n11598, n11599,
         n11600, n11601, n11602, n11603, n11604, n11605, n11606, n11607,
         n11608, n11609, n11610, n11611, n11612, n11613, n11614, n11615,
         n11616, n11617, n11618, n11619, n11620, n11621, n11622, n11623,
         n11624, n11625, n11626, n11627, n11628, n11629, n11630, n11631,
         n11632, n11633, n11634, n11635, n11636, n11637, n11638, n11639,
         n11640, n11641, n11642, n11643, n11644, n11645, n11646, n11647,
         n11648, n11649, n11650, n11651, n11652, n11653, n11654, n11655,
         n11656, n11657, n11658, n11659, n11660, n11661, n11662, n11663,
         n11664, n11665, n11666, n11667, n11668, n11669, n11670, n11671,
         n11672, n11673, n11674, n11675, n11676, n11677, n11678, n11679,
         n11680, n11681, n11682, n11683, n11684, n11685, n11686, n11687,
         n11688, n11689, n11690, n11691, n11692, n11693, n11694, n11695,
         n11696, n11697, n11698, n11699, n11700, n11701, n11702, n11703,
         n11704, n11705, n11706, n11707, n11708, n11709, n11710, n11711,
         n11712, n11713, n11714, n11715, n11716, n11717, n11718, n11719,
         n11720, n11721, n11722, n11723, n11724, n11725, n11726, n11727,
         n11728, n11729, n11730, n11731, n11732, n11733, n11734, n11735,
         n11736, n11737, n11738, n11739, n11740, n11741, n11742, n11743,
         n11744, n11745, n11746, n11747, n11748, n11749, n11750, n11751,
         n11752, n11753, n11754, n11755, n11756, n11757, n11758, n11759,
         n11760, n11761, n11762, n11763, n11764, n11765, n11766, n11767,
         n11768, n11769, n11770, n11771, n11772, n11773, n11774, n11775,
         n11776, n11777, n11778, n11779, n11780, n11781, n11782, n11783,
         n11784, n11785, n11786, n11787, n11788, n11789, n11790, n11791,
         n11792, n11793, n11794, n11795, n11796, n11797, n11798, n11799,
         n11800, n11801, n11802, n11803, n11804, n11805, n11806, n11807,
         n11808, n11809, n11810, n11811, n11812, n11813, n11814, n11815,
         n11816, n11817, n11818, n11819, n11820, n11821, n11822, n11823,
         n11824, n11825, n11826, n11827, n11828, n11829, n11830, n11831,
         n11832, n11833, n11834, n11835, n11836, n11837, n11838, n11839,
         n11840, n11841, n11842, n11843, n11844, n11845, n11846, n11847,
         n11848, n11849, n11850, n11851, n11852, n11853, n11854, n11855,
         n11856, n11857, n11858, n11859, n11860, n11861, n11862, n11863,
         n11864, n11865, n11866, n11867, n11868, n11869, n11870, n11871,
         n11872, n11873, n11874, n11875, n11876, n11877, n11878, n11879,
         n11880, n11881, n11882, n11883, n11884, n11885, n11886, n11887,
         n11888, n11889, n11890, n11891, n11892, n11893, n11894, n11895,
         n11896, n11897, n11898, n11899, n11900, n11901, n11902, n11903,
         n11904, n11905, n11906, n11907, n11908, n11909, n11910, n11911,
         n11912, n11913, n11914, n11915, n11916, n11917, n11918, n11919,
         n11920, n11921, n11922, n11923, n11924, n11925, n11926, n11927,
         n11928, n11929, n11930, n11931, n11932, n11933, n11934, n11935,
         n11936, n11937, n11938, n11939, n11940, n11941, n11942, n11943,
         n11944, n11945, n11946, n11947, n11948, n11949, n11950, n11951,
         n11952, n11953, n11954, n11955, n11956, n11957, n11958, n11959,
         n11960, n11961, n11962, n11963, n11964, n11965, n11966, n11967,
         n11968, n11969, n11970, n11971, n11972, n11973, n11974, n11975,
         n11976, n11977, n11978, n11979, n11980, n11981, n11982, n11983,
         n11984, n11985, n11986, n11987, n11988, n11989, n11990, n11991,
         n11992, n11993, n11994, n11995, n11996, n11997, n11998, n11999,
         n12000, n12001, n12002, n12003, n12004, n12005, n12006, n12007,
         n12008, n12009, n12010, n12011, n12012, n12013, n12014, n12015,
         n12016, n12017, n12018, n12019, n12020, n12021, n12022, n12023,
         n12024, n12025, n12026, n12027, n12028, n12029, n12030, n12031,
         n12032, n12033, n12034, n12035, n12036, n12037, n12038, n12039,
         n12040, n12041, n12042, n12043, n12044, n12045, n12046, n12047,
         n12048, n12049, n12050, n12051, n12052, n12053, n12054, n12055,
         n12056, n12057, n12058, n12059, n12060, n12061, n12062, n12063,
         n12064, n12065, n12066, n12067, n12068, n12069, n12070, n12071,
         n12072, n12073, n12074, n12075, n12076, n12077, n12078, n12079,
         n12080, n12081, n12082, n12083, n12084, n12085, n12086, n12087,
         n12088, n12089, n12090, n12091, n12092, n12093, n12094, n12095,
         n12096, n12097, n12098, n12099, n12100, n12101, n12102, n12103,
         n12104, n12105, n12106, n12107, n12108, n12109, n12110, n12111,
         n12112, n12113, n12114, n12115, n12116, n12117, n12118, n12119,
         n12120, n12121, n12122, n12123, n12124, n12125, n12126, n12127,
         n12128, n12129, n12130, n12131, n12132, n12133, n12134, n12135,
         n12136, n12137, n12138, n12139, n12140, n12141, n12142, n12143,
         n12144, n12145, n12146, n12147, n12148, n12149, n12150, n12151,
         n12152, n12153, n12154, n12155, n12156, n12157, n12158, n12159,
         n12160, n12161, n12162, n12163, n12164, n12165, n12166, n12167,
         n12168, n12169, n12170, n12171, n12172, n12173, n12174, n12175,
         n12176, n12177, n12178, n12179, n12180, n12181, n12182, n12183,
         n12184, n12185, n12186, n12187, n12188, n12189, n12190, n12191,
         n12192, n12193, n12194, n12195, n12196, n12197, n12198, n12199,
         n12200, n12201, n12202, n12203, n12204, n12205, n12206, n12207,
         n12208, n12209, n12210, n12211, n12212, n12213, n12214, n12215,
         n12216, n12217, n12218, n12219, n12220, n12221, n12222, n12223,
         n12224, n12225, n12226, n12227, n12228, n12229, n12230, n12231,
         n12232, n12233, n12234, n12235, n12236, n12237, n12238, n12239,
         n12240, n12241, n12242, n12243, n12244, n12245, n12246, n12247,
         n12248, n12249, n12250, n12251, n12252, n12253, n12254, n12255,
         n12256, n12257, n12258, n12259, n12260, n12261, n12262, n12263,
         n12264, n12265, n12266, n12267, n12268, n12269, n12270, n12271,
         n12272, n12273, n12274, n12275, n12276, n12277, n12278, n12279,
         n12280, n12281, n12282, n12283, n12284, n12285, n12286, n12287,
         n12288, n12289, n12290, n12291, n12292, n12293, n12294, n12295,
         n12296, n12297, n12298, n12299, n12300, n12301, n12302, n12303,
         n12304, n12305, n12306, n12307, n12308, n12309, n12310, n12311,
         n12312, n12313, n12314, n12315, n12316, n12317, n12318, n12319,
         n12320, n12321, n12322, n12323, n12324, n12325, n12326, n12327,
         n12328, n12329, n12330, n12331, n12332, n12333, n12334, n12335,
         n12336, n12337, n12338, n12339, n12340, n12341, n12342, n12343,
         n12344, n12345, n12346, n12347, n12348, n12349, n12350, n12351,
         n12352, n12353, n12354, n12355, n12356, n12357, n12358, n12359,
         n12360, n12361, n12362, n12363, n12364, n12365, n12366, n12367,
         n12368, n12369, n12370, n12371, n12372, n12373, n12374, n12375,
         n12376, n12377, n12378, n12379, n12380, n12381, n12382, n12383,
         n12384, n12385, n12386, n12387, n12388, n12389, n12390, n12391,
         n12392, n12393, n12394, n12395, n12396, n12397, n12398, n12399,
         n12400, n12401, n12402, n12403, n12404, n12405, n12406, n12407,
         n12408, n12409, n12410, n12411, n12412, n12413, n12414, n12415,
         n12416, n12417, n12418, n12419, n12420, n12421, n12422, n12423,
         n12424, n12425, n12426, n12427, n12428, n12429, n12430, n12431,
         n12432, n12433, n12434, n12435, n12436, n12437, n12438, n12439,
         n12440, n12441, n12442, n12443, n12444, n12445, n12446, n12447,
         n12448, n12449, n12450, n12451, n12452, n12453, n12454, n12455,
         n12456, n12457, n12458, n12459, n12460, n12461, n12462, n12463,
         n12464, n12465, n12466, n12467, n12468, n12469, n12470, n12471,
         n12472, n12473, n12474, n12475, n12476, n12477, n12478, n12479,
         n12480, n12481, n12482, n12483, n12484, n12485, n12486, n12487,
         n12488, n12489, n12490, n12491, n12492, n12493, n12494, n12495,
         n12496, n12497, n12498, n12499, n12500, n12501, n12502, n12503,
         n12504, n12505, n12506, n12507, n12508, n12509, n12510, n12511,
         n12512, n12513, n12514, n12515, n12516, n12517, n12518, n12519,
         n12520, n12521, n12522, n12523, n12524, n12525, n12526, n12527,
         n12528, n12529, n12530, n12531, n12532, n12533, n12534, n12535,
         n12536, n12537, n12538, n12539, n12540, n12541, n12542, n12543,
         n12544, n12545, n12546, n12547, n12548, n12549, n12550, n12551,
         n12552, n12553, n12554, n12555, n12556, n12557, n12558, n12559,
         n12560, n12561, n12562, n12563, n12564, n12565, n12566, n12567,
         n12568, n12569, n12570, n12571, n12572, n12573, n12574, n12575,
         n12576, n12577, n12578, n12579, n12580, n12581, n12582, n12583,
         n12584, n12585, n12586, n12587, n12588, n12589, n12590, n12591,
         n12592, n12593, n12594, n12595, n12596, n12597, n12598, n12599,
         n12600, n12601, n12602, n12603, n12604, n12605, n12606, n12607,
         n12608, n12609, n12610, n12611, n12612, n12613, n12614, n12615,
         n12616, n12617, n12618, n12619, n12620, n12621, n12622, n12623,
         n12624, n12625, n12626, n12627, n12628, n12629, n12630, n12631,
         n12632, n12633, n12634, n12635, n12636, n12637, n12638, n12639,
         n12640, n12641, n12642, n12643, n12644, n12645, n12646, n12647,
         n12648, n12649, n12650, n12651, n12652, n12653, n12654, n12655,
         n12656, n12657, n12658, n12659, n12660, n12661, n12662, n12663,
         n12664, n12665, n12666, n12667, n12668, n12669, n12670, n12671,
         n12672, n12673, n12674, n12675, n12676, n12677, n12678, n12679,
         n12680, n12681, n12682, n12683, n12684, n12685, n12686, n12687,
         n12688, n12689, n12690, n12691, n12692, n12693, n12694, n12695,
         n12696, n12697, n12698, n12699, n12700, n12701, n12702, n12703,
         n12704, n12705, n12706, n12707, n12708, n12709, n12710, n12711,
         n12712, n12713, n12714, n12715, n12716, n12717, n12718, n12719,
         n12720, n12721, n12722, n12723, n12724, n12725, n12726, n12727,
         n12728, n12729, n12730, n12731, n12732, n12733, n12734, n12735,
         n12736, n12737, n12738, n12739, n12740, n12741, n12742, n12743,
         n12744, n12745, n12746, n12747, n12748, n12749, n12750, n12751,
         n12752, n12753, n12754, n12755, n12756, n12757, n12758, n12759,
         n12760, n12761, n12762, n12763, n12764, n12765, n12766, n12767,
         n12768, n12769, n12770, n12771, n12772, n12773, n12774, n12775,
         n12776, n12777, n12778, n12779, n12780, n12781, n12782, n12783,
         n12784, n12785, n12786, n12787, n12788, n12789, n12790, n12791,
         n12792, n12793, n12794, n12795, n12796, n12797, n12798, n12799,
         n12800, n12801, n12802, n12803, n12804, n12805, n12806, n12807,
         n12808, n12809, n12810, n12811, n12812, n12813, n12814, n12815,
         n12816, n12817, n12818, n12819, n12820, n12821, n12822, n12823,
         n12824, n12825, n12826, n12827, n12828, n12829, n12830, n12831,
         n12832, n12833, n12834, n12835, n12836, n12837, n12838, n12839,
         n12840, n12841, n12842, n12843, n12844, n12845, n12846, n12847,
         n12848, n12849, n12850, n12851, n12852, n12853, n12854, n12855,
         n12856, n12857, n12858, n12859, n12860, n12861, n12862, n12863,
         n12864, n12865, n12866, n12867, n12868, n12869, n12870, n12871,
         n12872, n12873, n12874, n12875, n12876, n12877, n12878, n12879,
         n12880, n12881, n12882, n12883, n12884, n12885, n12886, n12887,
         n12888, n12889, n12890, n12891, n12892, n12893, n12894, n12895,
         n12896, n12897, n12898, n12899, n12900, n12901, n12902, n12903,
         n12904, n12905, n12906, n12907, n12908, n12909, n12910, n12911,
         n12912, n12913, n12914, n12915, n12916, n12917, n12918, n12919,
         n12920, n12921, n12922, n12923, n12924, n12925, n12926, n12927,
         n12928, n12929, n12930, n12931, n12932, n12933, n12934, n12935,
         n12936, n12937, n12938, n12939, n12940, n12941, n12942, n12943,
         n12944, n12945, n12946, n12947, n12948, n12949, n12950, n12951,
         n12952, n12953, n12954, n12955, n12956, n12957, n12958, n12959,
         n12960, n12961, n12962, n12963, n12964, n12965, n12966, n12967,
         n12968, n12969, n12970, n12971, n12972, n12973, n12974, n12975,
         n12976, n12977, n12978, n12979, n12980, n12981, n12982, n12983,
         n12984, n12985, n12986, n12987, n12988, n12989, n12990, n12991,
         n12992, n12993, n12994, n12995, n12996, n12997, n12998, n12999,
         n13000, n13001, n13002, n13003, n13004, n13005, n13006, n13007,
         n13008, n13009, n13010, n13011, n13012, n13013, n13014, n13015,
         n13016, n13017, n13018, n13019, n13020, n13021, n13022, n13023,
         n13024, n13025, n13026, n13027, n13028, n13029, n13030, n13031,
         n13032, n13033, n13034, n13035, n13036, n13037, n13038, n13039,
         n13040, n13041, n13042, n13043, n13044, n13045, n13046, n13047,
         n13048, n13049, n13050, n13051, n13052, n13053, n13054, n13055,
         n13056, n13057, n13058, n13059, n13060, n13061, n13062, n13063,
         n13064, n13065, n13066, n13067, n13068, n13069, n13070, n13071,
         n13072, n13073, n13074, n13075, n13076, n13077, n13078, n13079,
         n13080, n13081, n13082, n13083, n13084, n13085, n13086, n13087,
         n13088, n13089, n13090, n13091, n13092, n13093, n13094, n13095,
         n13096, n13097, n13098, n13099, n13100, n13101, n13102, n13103,
         n13104, n13105, n13106, n13107, n13108, n13109, n13110, n13111,
         n13112, n13113, n13114, n13115, n13116, n13117, n13118, n13119,
         n13120, n13121, n13122, n13123, n13124, n13125, n13126, n13127,
         n13128, n13129, n13130, n13131, n13132, n13133, n13134, n13135,
         n13136, n13137, n13138, n13139, n13140, n13141, n13142, n13143,
         n13144, n13145, n13146, n13147, n13148, n13149, n13150, n13151,
         n13152, n13153, n13154, n13155, n13156, n13157, n13158, n13159,
         n13160, n13161, n13162, n13163, n13164, n13165, n13166, n13167,
         n13168, n13169, n13170, n13171, n13172, n13173, n13174, n13175,
         n13176, n13177, n13178, n13179, n13180, n13181, n13182, n13183,
         n13184, n13185, n13186, n13187, n13188, n13189, n13190, n13191,
         n13192, n13193, n13194, n13195, n13196, n13197, n13198, n13199,
         n13200, n13201, n13202, n13203, n13204, n13205, n13206, n13207,
         n13208, n13209, n13210, n13211, n13212, n13213, n13214, n13215,
         n13216, n13217, n13218, n13219, n13220, n13221, n13222, n13223,
         n13224, n13225, n13226, n13227, n13228, n13229, n13230, n13231,
         n13232, n13233, n13234, n13235, n13236, n13237, n13238, n13239,
         n13240, n13241, n13242, n13243, n13244, n13245, n13246, n13247,
         n13248, n13249, n13250, n13251, n13252, n13253, n13254, n13255,
         n13256, n13257, n13258, n13259, n13260, n13261, n13262, n13263,
         n13264, n13265, n13266, n13267, n13268, n13269, n13270, n13271,
         n13272, n13273, n13274, n13275, n13276, n13277, n13278, n13279,
         n13280, n13281, n13282, n13283, n13284, n13285, n13286, n13287,
         n13288, n13289, n13290, n13291, n13292, n13293, n13294, n13295,
         n13296, n13297, n13298, n13299, n13300, n13301, n13302, n13303,
         n13304, n13305, n13306, n13307, n13308, n13309, n13310, n13311,
         n13312, n13313, n13314, n13315, n13316, n13317, n13318, n13319,
         n13320, n13321, n13322, n13323, n13324, n13325, n13326, n13327,
         n13328, n13329, n13330, n13331, n13332, n13333, n13334, n13335,
         n13336, n13337, n13338, n13339, n13340, n13341, n13342, n13343,
         n13344, n13345, n13346, n13347, n13348, n13349, n13350, n13351,
         n13352, n13353, n13354, n13355, n13356, n13357, n13358, n13359,
         n13360, n13361, n13362, n13363, n13364, n13365, n13366, n13367,
         n13368, n13369, n13370, n13371, n13372, n13373, n13374, n13375,
         n13376, n13377, n13378, n13379, n13380, n13381, n13382, n13383,
         n13384, n13385, n13386, n13387, n13388, n13389, n13390, n13391,
         n13392, n13393, n13394, n13395, n13396, n13397, n13398, n13399,
         n13400, n13401, n13402, n13403, n13404, n13405, n13406, n13407,
         n13408, n13409, n13410, n13411, n13412, n13413, n13414, n13415,
         n13416, n13417, n13418, n13419, n13420, n13421, n13422, n13423,
         n13424, n13425, n13426, n13427, n13428, n13429, n13430, n13431,
         n13432, n13433, n13434, n13435, n13436, n13437, n13438, n13439,
         n13440, n13441, n13442, n13443, n13444, n13445, n13446, n13447,
         n13448, n13449, n13450, n13451, n13452, n13453, n13454, n13455,
         n13456, n13457, n13458, n13459, n13460, n13461, n13462, n13463,
         n13464, n13465, n13466, n13467, n13468, n13469, n13470, n13471,
         n13472, n13473, n13474, n13475, n13476, n13477, n13478, n13479,
         n13480, n13481, n13482, n13483, n13484, n13485, n13486, n13487,
         n13488, n13489, n13490, n13491, n13492, n13493, n13494, n13495,
         n13496, n13497, n13498, n13499, n13500, n13501, n13502, n13503,
         n13504, n13505, n13506, n13507, n13508, n13509, n13510, n13511,
         n13512, n13513, n13514, n13515, n13516, n13517, n13518, n13519,
         n13520, n13521, n13522, n13523, n13524, n13525, n13526, n13527,
         n13528, n13529, n13530, n13531, n13532, n13533, n13534, n13535,
         n13536, n13537, n13538, n13539, n13540, n13541, n13542, n13543,
         n13544, n13545, n13546, n13547, n13548, n13549, n13550, n13551,
         n13552, n13553, n13554, n13555, n13556, n13557, n13558, n13559,
         n13560, n13561, n13562, n13563, n13564, n13565, n13566, n13567,
         n13568, n13569, n13570, n13571, n13572, n13573, n13574, n13575,
         n13576, n13577, n13578, n13579, n13580, n13581, n13582, n13583,
         n13584, n13585, n13586, n13587, n13588, n13589, n13590, n13591,
         n13592, n13593, n13594, n13595, n13596, n13597, n13598, n13599,
         n13600, n13601, n13602, n13603, n13604, n13605, n13606, n13607,
         n13608, n13609, n13610, n13611, n13612, n13613, n13614, n13615,
         n13616, n13617, n13618, n13619, n13620, n13621, n13622, n13623,
         n13624, n13625, n13626, n13627, n13628, n13629, n13630, n13631,
         n13632, n13633, n13634, n13635, n13636, n13637, n13638, n13639,
         n13640, n13641, n13642, n13643, n13644, n13645, n13646, n13647,
         n13648, n13649, n13650, n13651, n13652, n13653, n13654, n13655,
         n13656, n13657, n13658, n13659, n13660, n13661, n13662, n13663,
         n13664, n13665, n13666, n13667, n13668, n13669, n13670, n13671,
         n13672, n13673, n13674, n13675, n13676, n13677, n13678, n13679,
         n13680, n13681, n13682, n13683, n13684, n13685, n13686, n13687,
         n13688, n13689, n13690, n13691, n13692, n13693, n13694, n13695,
         n13696, n13697, n13698, n13699, n13700, n13701, n13702, n13703,
         n13704, n13705, n13706, n13707, n13708, n13709, n13710, n13711,
         n13712, n13713, n13714, n13715, n13716, n13717, n13718, n13719,
         n13720, n13721, n13722, n13723, n13724, n13725, n13726, n13727,
         n13728, n13729, n13730, n13731, n13732, n13733, n13734, n13735,
         n13736, n13737, n13738, n13739, n13740, n13741, n13742, n13743,
         n13744, n13745, n13746, n13747, n13748, n13749, n13750, n13751,
         n13752, n13753, n13754, n13755, n13756, n13757, n13758, n13759,
         n13760, n13761, n13762, n13763, n13764, n13765, n13766, n13767,
         n13768, n13769, n13770, n13771, n13772, n13773, n13774, n13775,
         n13776, n13777, n13778, n13779, n13780, n13781, n13782, n13783,
         n13784, n13785, n13786, n13787, n13788, n13789, n13790, n13791,
         n13792, n13793, n13794, n13795, n13796, n13797, n13798, n13799,
         n13800, n13801, n13802, n13803, n13804, n13805, n13806, n13807,
         n13808, n13809, n13810, n13811, n13812, n13813, n13814, n13815,
         n13816, n13817, n13818, n13819, n13820, n13821, n13822, n13823,
         n13824, n13825, n13826, n13827, n13828, n13829, n13830, n13831,
         n13832, n13833, n13834, n13835, n13836, n13837, n13838, n13839,
         n13840, n13841, n13842, n13843, n13844, n13845, n13846, n13847,
         n13848, n13849, n13850, n13851, n13852, n13853, n13854, n13855,
         n13856, n13857, n13858, n13859, n13860, n13861, n13862, n13863,
         n13864, n13865, n13866, n13867, n13868, n13869, n13870, n13871,
         n13872, n13873, n13874, n13875, n13876, n13877, n13878, n13879,
         n13880, n13881, n13882, n13883, n13884, n13885, n13886, n13887,
         n13888, n13889, n13890, n13891, n13892, n13893, n13894, n13895,
         n13896, n13897, n13898, n13899, n13900, n13901, n13902, n13903,
         n13904, n13905, n13906, n13907, n13908, n13909, n13910, n13911,
         n13912, n13913, n13914, n13915, n13916, n13917, n13918, n13919,
         n13920, n13921, n13922, n13923, n13924, n13925, n13926, n13927,
         n13928, n13929, n13930, n13931, n13932, n13933, n13934, n13935,
         n13936, n13937, n13938, n13939, n13940, n13941, n13942, n13943,
         n13944, n13945, n13946, n13947, n13948, n13949, n13950, n13951,
         n13952, n13953, n13954, n13955, n13956, n13957, n13958, n13959,
         n13960, n13961, n13962, n13963, n13964, n13965, n13966, n13967,
         n13968, n13969, n13970, n13971, n13972, n13973, n13974, n13975,
         n13976, n13977, n13978, n13979, n13980, n13981, n13982, n13983,
         n13984, n13985, n13986, n13987, n13988, n13989, n13990, n13991,
         n13992, n13993, n13994, n13995, n13996, n13997, n13998, n13999,
         n14000, n14001, n14002, n14003, n14004, n14005, n14006, n14007,
         n14008, n14009, n14010, n14011, n14012, n14013, n14014, n14015,
         n14016, n14017, n14018, n14019, n14020, n14021, n14022, n14023,
         n14024, n14025, n14026, n14027, n14028, n14029, n14030, n14031,
         n14032, n14033, n14034, n14035, n14036, n14037, n14038, n14039,
         n14040, n14041, n14042, n14043, n14044, n14045, n14046, n14047,
         n14048, n14049, n14050, n14051, n14052, n14053, n14054, n14055,
         n14056, n14057, n14058, n14059, n14060, n14061, n14062, n14063,
         n14064, n14065, n14066, n14067, n14068, n14069, n14070, n14071,
         n14072, n14073, n14074, n14075, n14076, n14077, n14078, n14079,
         n14080, n14081, n14082, n14083, n14084, n14085, n14086, n14087,
         n14088, n14089, n14090, n14091, n14092, n14093, n14094, n14095,
         n14096, n14097, n14098, n14099, n14100, n14101, n14102, n14103,
         n14104, n14105, n14106, n14107, n14108, n14109, n14110, n14111,
         n14112, n14113, n14114, n14115, n14116, n14117, n14118, n14119,
         n14120, n14121, n14122, n14123, n14124, n14125, n14126, n14127,
         n14128, n14129, n14130, n14131, n14132, n14133, n14134, n14135,
         n14136, n14137, n14138, n14139, n14140, n14141, n14142, n14143,
         n14144, n14145, n14146, n14147, n14148, n14149, n14150, n14151,
         n14152, n14153, n14154, n14155, n14156, n14157, n14158, n14159,
         n14160, n14161, n14162, n14163, n14164, n14165, n14166, n14167,
         n14168, n14169, n14170, n14171, n14172, n14173, n14174, n14175,
         n14176, n14177, n14178, n14179, n14180, n14181, n14182, n14183,
         n14184, n14185, n14186, n14187, n14188, n14189, n14190, n14191,
         n14192, n14193, n14194, n14195, n14196, n14197, n14198, n14199,
         n14200, n14201, n14202, n14203, n14204, n14205, n14206, n14207,
         n14208, n14209, n14210, n14211, n14212, n14213, n14214, n14215,
         n14216, n14217, n14218, n14219, n14220, n14221, n14222, n14223,
         n14224, n14225, n14226, n14227, n14228, n14229, n14230, n14231,
         n14232, n14233, n14234, n14235, n14236, n14237, n14238, n14239,
         n14240, n14241, n14242, n14243, n14244, n14245, n14246, n14247,
         n14248, n14249, n14250, n14251, n14252, n14253, n14254, n14255,
         n14256, n14257, n14258, n14259, n14260, n14261, n14262, n14263,
         n14264, n14265, n14266, n14267, n14268, n14269, n14270, n14271,
         n14272, n14273, n14274, n14275, n14276, n14277, n14278, n14279,
         n14280, n14281, n14282, n14283, n14284, n14285, n14286, n14287,
         n14288, n14289, n14290, n14291, n14292, n14293, n14294, n14295,
         n14296, n14297, n14298, n14299, n14300, n14301, n14302, n14303,
         n14304, n14305, n14306, n14307, n14308, n14309, n14310, n14311,
         n14312, n14313, n14314, n14315, n14316, n14317, n14318, n14319,
         n14320, n14321, n14322, n14323, n14324, n14325, n14326, n14327,
         n14328, n14329, n14330, n14331, n14332, n14333, n14334, n14335,
         n14336, n14337, n14338, n14339, n14340, n14341, n14342, n14343,
         n14344, n14345, n14346, n14347, n14348, n14349, n14350, n14351,
         n14352, n14353, n14354, n14355, n14356, n14357, n14358, n14359,
         n14360, n14361, n14362, n14363, n14364, n14365, n14366, n14367,
         n14368, n14369, n14370, n14371, n14372, n14373, n14374, n14375,
         n14376, n14377, n14378, n14379, n14380, n14381, n14382, n14383,
         n14384, n14385, n14386, n14387, n14388, n14389, n14390, n14391,
         n14392, n14393, n14394, n14395, n14396, n14397, n14398, n14399,
         n14400, n14401, n14402, n14403, n14404, n14405, n14406, n14407,
         n14408, n14409, n14410, n14411, n14412, n14413, n14414, n14415,
         n14416, n14417, n14418, n14419, n14420, n14421, n14422, n14423,
         n14424, n14425, n14426, n14427, n14428, n14429, n14430, n14431,
         n14432, n14433, n14434, n14435, n14436, n14437, n14438, n14439,
         n14440, n14441, n14442, n14443, n14444, n14445, n14446, n14447,
         n14448, n14449, n14450, n14451, n14452, n14453, n14454, n14455,
         n14456, n14457, n14458, n14459, n14460, n14461, n14462, n14463,
         n14464, n14465, n14466, n14467, n14468, n14469, n14470, n14471,
         n14472, n14473, n14474, n14475, n14476, n14477, n14478, n14479,
         n14480, n14481, n14482, n14483, n14484, n14485, n14486, n14487,
         n14488, n14489, n14490, n14491, n14492, n14493, n14494, n14495,
         n14496, n14497, n14498, n14499, n14500, n14501, n14502, n14503,
         n14504, n14505, n14506, n14507, n14508, n14509, n14510, n14511,
         n14512, n14513, n14514, n14515, n14516, n14517, n14518, n14519,
         n14520, n14521, n14522, n14523, n14524, n14525, n14526, n14527,
         n14528, n14529, n14530, n14531, n14532, n14533, n14534, n14535,
         n14536, n14537, n14538, n14539, n14540, n14541, n14542, n14543,
         n14544, n14545, n14546, n14547, n14548, n14549, n14550, n14551,
         n14552, n14553, n14554, n14555, n14556, n14557, n14558, n14559,
         n14560, n14561, n14562, n14563, n14564, n14565, n14566, n14567,
         n14568, n14569, n14570, n14571, n14572, n14573, n14574, n14575,
         n14576, n14577, n14578, n14579, n14580, n14581, n14582, n14583,
         n14584, n14585, n14586, n14587, n14588, n14589, n14590, n14591,
         n14592, n14593, n14594, n14595, n14596, n14597, n14598, n14599,
         n14600, n14601, n14602, n14603, n14604, n14605, n14606, n14607,
         n14608, n14609, n14610, n14611, n14612, n14613, n14614, n14615,
         n14616, n14617, n14618, n14619, n14620, n14621, n14622, n14623,
         n14624, n14625, n14626, n14627, n14628, n14629, n14630, n14631,
         n14632, n14633, n14634, n14635, n14636, n14637, n14638, n14639,
         n14640, n14641, n14642, n14643, n14644, n14645, n14646, n14647,
         n14648, n14649, n14650, n14651, n14652, n14653, n14654, n14655,
         n14656, n14657, n14658, n14659, n14660, n14661, n14662, n14663,
         n14664, n14665, n14666, n14667, n14668, n14669, n14670, n14671,
         n14672, n14673, n14674, n14675, n14676, n14677, n14678, n14679,
         n14680, n14681, n14682, n14683, n14684, n14685, n14686, n14687,
         n14688, n14689, n14690, n14691, n14692, n14693, n14694, n14695,
         n14696, n14697, n14698, n14699, n14700, n14701, n14702, n14703,
         n14704, n14705, n14706, n14707, n14708, n14709, n14710, n14711,
         n14712, n14713, n14714, n14715, n14716, n14717, n14718, n14719,
         n14720, n14721, n14722, n14723, n14724, n14725, n14726, n14727,
         n14728, n14729, n14730, n14731, n14732, n14733, n14734, n14735,
         n14736, n14737, n14738, n14739, n14740, n14741, n14742, n14743,
         n14744, n14745, n14746, n14747, n14748, n14749, n14750, n14751,
         n14752, n14753, n14754, n14755, n14756, n14757, n14758, n14759,
         n14760, n14761, n14762, n14763, n14764, n14765, n14766, n14767,
         n14768, n14769, n14770, n14771, n14772, n14773, n14774, n14775,
         n14776, n14777, n14778, n14779, n14780, n14781, n14782, n14783,
         n14784, n14785, n14786, n14787, n14788, n14789, n14790, n14791,
         n14792, n14793, n14794, n14795, n14796, n14797, n14798, n14799,
         n14800, n14801, n14802, n14803, n14804, n14805, n14806, n14807,
         n14808, n14809, n14810, n14811, n14812, n14813, n14814, n14815,
         n14816, n14817, n14818, n14819, n14820, n14821, n14822, n14823,
         n14824, n14825, n14826, n14827, n14828, n14829, n14830, n14831,
         n14832, n14833, n14834, n14835, n14836, n14837, n14838, n14839,
         n14840, n14841, n14842, n14843, n14844, n14845, n14846, n14847,
         n14848, n14849, n14850, n14851, n14852, n14853, n14854, n14855,
         n14856, n14857, n14858, n14859, n14860, n14861, n14862, n14863,
         n14864, n14865, n14866, n14867, n14868, n14869, n14870, n14871,
         n14872, n14873, n14874, n14875, n14876, n14877, n14878, n14879,
         n14880, n14881, n14882, n14883, n14884, n14885, n14886, n14887,
         n14888, n14889, n14890, n14891, n14892, n14893, n14894, n14895,
         n14896, n14897, n14898, n14899, n14900, n14901, n14902, n14903,
         n14904, n14905, n14906, n14907, n14908, n14909, n14910, n14911,
         n14912, n14913, n14914, n14915, n14916, n14917, n14918, n14919,
         n14920, n14921, n14922, n14923, n14924, n14925, n14926, n14927,
         n14928, n14929, n14930, n14931, n14932, n14933, n14934, n14935,
         n14936, n14937, n14938, n14939, n14940, n14941, n14942, n14943,
         n14944, n14945, n14946, n14947, n14948, n14949, n14950, n14951,
         n14952, n14953, n14954, n14955, n14956, n14957, n14958, n14959,
         n14960, n14961, n14962, n14963, n14964, n14965, n14966, n14967,
         n14968, n14969, n14970, n14971, n14972, n14973, n14974, n14975,
         n14976, n14977, n14978, n14979, n14980, n14981, n14982, n14983,
         n14984, n14985, n14986, n14987, n14988, n14989, n14990, n14991,
         n14992, n14993, n14994, n14995, n14996, n14997, n14998, n14999,
         n15000, n15001, n15002, n15003, n15004, n15005, n15006, n15007,
         n15008, n15009, n15010, n15011, n15012, n15013, n15014, n15015,
         n15016, n15017, n15018, n15019, n15020, n15021, n15022, n15023,
         n15024, n15025, n15026, n15027, n15028, n15029, n15030, n15031,
         n15032, n15033, n15034, n15035, n15036, n15037, n15038, n15039,
         n15040, n15041, n15042, n15043, n15044, n15045, n15046, n15047,
         n15048, n15049, n15050, n15051, n15052, n15053, n15054, n15055,
         n15056, n15057, n15058, n15059, n15060, n15061, n15062, n15063,
         n15064, n15065, n15066, n15067, n15068, n15069, n15070, n15071,
         n15072, n15073, n15074, n15075, n15076, n15077, n15078, n15079,
         n15080, n15081, n15082, n15083, n15084, n15085, n15086, n15087,
         n15088, n15089, n15090, n15091, n15092, n15093, n15094, n15095,
         n15096, n15097, n15098, n15099, n15100, n15101, n15102, n15103,
         n15104, n15105, n15106, n15107, n15108, n15109, n15110, n15111,
         n15112, n15113, n15114, n15115, n15116, n15117, n15118, n15119,
         n15120, n15121, n15122, n15123, n15124, n15125, n15126, n15127,
         n15128, n15129, n15130, n15131, n15132, n15133, n15134, n15135,
         n15136, n15137, n15138, n15139, n15140, n15141, n15142, n15143,
         n15144, n15145, n15146, n15147, n15148, n15149, n15150, n15151,
         n15152, n15153, n15154, n15155, n15156, n15157, n15158, n15159,
         n15160, n15161, n15162, n15163, n15164, n15165, n15166, n15167,
         n15168, n15169, n15170, n15171, n15172, n15173, n15174, n15175,
         n15176, n15177, n15178, n15179, n15180, n15181, n15182, n15183,
         n15184, n15185, n15186, n15187, n15188, n15189, n15190, n15191,
         n15192, n15193, n15194, n15195, n15196, n15197, n15198, n15199,
         n15200, n15201, n15202, n15203, n15204, n15205, n15206, n15207,
         n15208, n15209, n15210, n15211, n15212, n15213, n15214, n15215,
         n15216, n15217, n15218, n15219, n15220, n15221, n15222, n15223,
         n15224, n15225, n15226, n15227, n15228, n15229, n15230, n15231,
         n15232, n15233, n15234, n15235, n15236, n15237, n15238, n15239,
         n15240, n15241, n15242, n15243, n15244, n15245, n15246, n15247,
         n15248, n15249, n15250, n15251, n15252, n15253, n15254, n15255,
         n15256, n15257, n15258, n15259, n15260, n15261, n15262, n15263,
         n15264, n15265, n15266, n15267, n15268, n15269, n15270, n15271,
         n15272, n15273, n15274, n15275, n15276, n15277, n15278, n15279,
         n15280, n15281, n15282, n15283, n15284, n15285, n15286, n15287,
         n15288, n15289, n15290, n15291, n15292, n15293, n15294, n15295,
         n15296, n15297, n15298, n15299, n15300, n15301, n15302, n15303,
         n15304, n15305, n15306, n15307, n15308, n15309, n15310, n15311,
         n15312, n15313, n15314, n15315, n15316, n15317, n15318, n15319,
         n15320, n15321, n15322, n15323, n15324, n15325, n15326, n15327,
         n15328, n15329, n15330, n15331, n15332, n15333, n15334, n15335,
         n15336, n15337, n15338, n15339, n15340, n15341, n15342, n15343,
         n15344, n15345, n15346, n15347, n15348, n15349, n15350, n15351,
         n15352, n15353, n15354, n15355, n15356, n15357, n15358, n15359,
         n15360, n15361, n15362, n15363, n15364, n15365, n15366, n15367,
         n15368, n15369, n15370, n15371, n15372, n15373, n15374, n15375,
         n15376, n15377, n15378, n15379, n15380, n15381, n15382, n15383,
         n15384, n15385, n15386, n15387, n15388, n15389, n15390, n15391,
         n15392, n15393, n15394, n15395, n15396, n15397, n15398, n15399,
         n15400, n15401, n15402, n15403, n15404, n15405, n15406, n15407,
         n15408, n15409, n15410, n15411, n15412, n15413, n15414, n15415,
         n15416, n15417, n15418, n15419, n15420, n15421, n15422, n15423,
         n15424, n15425, n15426, n15427, n15428, n15429, n15430, n15431,
         n15432, n15433, n15434, n15435, n15436, n15437, n15438, n15439,
         n15440, n15441, n15442, n15443, n15444, n15445, n15446, n15447,
         n15448, n15449, n15450, n15451, n15452, n15453, n15454, n15455,
         n15456, n15457, n15458, n15459, n15460, n15461, n15462, n15463,
         n15464, n15465, n15466, n15467, n15468, n15469, n15470, n15471,
         n15472, n15473, n15474, n15475, n15476, n15477, n15478, n15479,
         n15480, n15481, n15482, n15483, n15484, n15485, n15486, n15487,
         n15488, n15489, n15490, n15491, n15492, n15493, n15494, n15495,
         n15496, n15497, n15498, n15499, n15500, n15501, n15502, n15503,
         n15504, n15505, n15506, n15507, n15508, n15509, n15510, n15511,
         n15512, n15513, n15514, n15515, n15516, n15517, n15518, n15519,
         n15520, n15521, n15522, n15523, n15524, n15525, n15526, n15527,
         n15528, n15529, n15530, n15531, n15532, n15533, n15534, n15535,
         n15536, n15537, n15538, n15539, n15540, n15541, n15542, n15543,
         n15544, n15545, n15546, n15547, n15548, n15549, n15550, n15551,
         n15552, n15553, n15554, n15555, n15556, n15557, n15558, n15559,
         n15560, n15561, n15562, n15563, n15564, n15565, n15566, n15567,
         n15568, n15569, n15570, n15571, n15572, n15573, n15574, n15575,
         n15576, n15577, n15578, n15579, n15580, n15581, n15582, n15583,
         n15584, n15585, n15586, n15587, n15588, n15589, n15590, n15591,
         n15592, n15593, n15594, n15595, n15596, n15597, n15598, n15599,
         n15600, n15601, n15602, n15603, n15604, n15605, n15606, n15607,
         n15608, n15609, n15610, n15611, n15612, n15613, n15614, n15615,
         n15616, n15617, n15618, n15619, n15620, n15621, n15622, n15623,
         n15624, n15625, n15626, n15627, n15628, n15629, n15630, n15631,
         n15632, n15633, n15634, n15635, n15636, n15637, n15638, n15639,
         n15640, n15641, n15642, n15643, n15644, n15645, n15646, n15647,
         n15648, n15649, n15650, n15651, n15652, n15653, n15654, n15655,
         n15656, n15657, n15658, n15659, n15660, n15661, n15662, n15663,
         n15664, n15665, n15666, n15667, n15668, n15669, n15670, n15671,
         n15672, n15673, n15674, n15675, n15676, n15677, n15678, n15679,
         n15680, n15681, n15682, n15683, n15684, n15685, n15686, n15687,
         n15688, n15689, n15690, n15691, n15692, n15693, n15694, n15695,
         n15696, n15697, n15698, n15699, n15700, n15701, n15702, n15703,
         n15704, n15705, n15706, n15707, n15708, n15709, n15710, n15711,
         n15712, n15713, n15714, n15715, n15716, n15717, n15718, n15719,
         n15720, n15721, n15722, n15723, n15724, n15725, n15726, n15727,
         n15728, n15729, n15730, n15731, n15732, n15733, n15734, n15735,
         n15736, n15737, n15738, n15739, n15740, n15741, n15742, n15743,
         n15744, n15745, n15746, n15747, n15748, n15749, n15750, n15751,
         n15752, n15753, n15754, n15755, n15756, n15757, n15758, n15759,
         n15760, n15761, n15762, n15763, n15764, n15765, n15766, n15767,
         n15768, n15769, n15770, n15771, n15772, n15773, n15774, n15775,
         n15776, n15777, n15778, n15779, n15780, n15781, n15782, n15783,
         n15784, n15785, n15786, n15787, n15788, n15789, n15790, n15791,
         n15792, n15793, n15794, n15795, n15796, n15797, n15798, n15799,
         n15800, n15801, n15802, n15803, n15804, n15805, n15806, n15807,
         n15808, n15809, n15810, n15811, n15812, n15813, n15814, n15815,
         n15816, n15817, n15818, n15819, n15820, n15821, n15822, n15823,
         n15824, n15825, n15826, n15827, n15828, n15829, n15830, n15831,
         n15832, n15833, n15834, n15835, n15836, n15837, n15838, n15839,
         n15840, n15841, n15842, n15843, n15844, n15845, n15846, n15847,
         n15848, n15849, n15850, n15851, n15852, n15853, n15854, n15855,
         n15856, n15857, n15858, n15859, n15860, n15861, n15862, n15863,
         n15864, n15865, n15866, n15867, n15868, n15869, n15870, n15871,
         n15872, n15873, n15874, n15875, n15876, n15877, n15878, n15879,
         n15880, n15881, n15882, n15883, n15884, n15885, n15886, n15887,
         n15888, n15889, n15890, n15891, n15892, n15893, n15894, n15895,
         n15896, n15897, n15898, n15899, n15900, n15901, n15902, n15903,
         n15904, n15905, n15906, n15907, n15908, n15909, n15910, n15911,
         n15912, n15913, n15914, n15915, n15916, n15917, n15918, n15919,
         n15920, n15921, n15922, n15923, n15924, n15925, n15926, n15927,
         n15928, n15929, n15930, n15931, n15932, n15933, n15934, n15935,
         n15936, n15937, n15938, n15939, n15940, n15941, n15942, n15943,
         n15944, n15945, n15946, n15947, n15948, n15949, n15950, n15951,
         n15952, n15953, n15954, n15955, n15956, n15957, n15958, n15959,
         n15960, n15961, n15962, n15963, n15964, n15965, n15966, n15967,
         n15968, n15969, n15970, n15971, n15972, n15973, n15974, n15975,
         n15976, n15977, n15978, n15979, n15980, n15981, n15982, n15983,
         n15984, n15985, n15986, n15987, n15988, n15989, n15990, n15991,
         n15992, n15993, n15994, n15995, n15996, n15997, n15998, n15999,
         n16000, n16001, n16002, n16003, n16004, n16005, n16006, n16007,
         n16008, n16009, n16010, n16011, n16012, n16013, n16014, n16015,
         n16016, n16017, n16018, n16019, n16020, n16021, n16022, n16023,
         n16024, n16025, n16026, n16027, n16028, n16029, n16030, n16031,
         n16032, n16033, n16034, n16035, n16036, n16037, n16038, n16039,
         n16040, n16041, n16042, n16043, n16044, n16045, n16046, n16047,
         n16048, n16049, n16050, n16051, n16052, n16053, n16054, n16055,
         n16056, n16057, n16058, n16059, n16060, n16061, n16062, n16063,
         n16064, n16065, n16066, n16067, n16068, n16069, n16070, n16071,
         n16072, n16073, n16074, n16075, n16076, n16077, n16078, n16079,
         n16080, n16081, n16082, n16083, n16084, n16085, n16086, n16087,
         n16088, n16089, n16090, n16091, n16092, n16093, n16094, n16095,
         n16096, n16097, n16098, n16099, n16100, n16101, n16102, n16103,
         n16104, n16105, n16106, n16107, n16108, n16109, n16110, n16111,
         n16112, n16113, n16114, n16115, n16116, n16117, n16118, n16119,
         n16120, n16121, n16122, n16123, n16124, n16125, n16126, n16127,
         n16128, n16129, n16130, n16131, n16132, n16133, n16134, n16135,
         n16136, n16137, n16138, n16139, n16140, n16141, n16142, n16143,
         n16144, n16145, n16146, n16147, n16148, n16149, n16150, n16151,
         n16152, n16153, n16154, n16155, n16156, n16157, n16158, n16159,
         n16160, n16161, n16162, n16163, n16164, n16165, n16166, n16167,
         n16168, n16169, n16170, n16171, n16172, n16173, n16174, n16175,
         n16176, n16177, n16178, n16179, n16180, n16181, n16182, n16183,
         n16184, n16185, n16186, n16187, n16188, n16189, n16190, n16191,
         n16192, n16193, n16194, n16195, n16196, n16197, n16198, n16199,
         n16200, n16201, n16202, n16203, n16204, n16205, n16206, n16207,
         n16208, n16209, n16210, n16211, n16212, n16213, n16214, n16215,
         n16216, n16217, n16218, n16219, n16220, n16221, n16222, n16223,
         n16224, n16225, n16226, n16227, n16228, n16229, n16230, n16231,
         n16232, n16233, n16234, n16235, n16236, n16237, n16238, n16239,
         n16240, n16241, n16242, n16243, n16244, n16245, n16246, n16247,
         n16248, n16249, n16250, n16251, n16252, n16253, n16254, n16255,
         n16256, n16257, n16258, n16259, n16260, n16261, n16262, n16263,
         n16264, n16265, n16266, n16267, n16268, n16269, n16270, n16271,
         n16272, n16273, n16274, n16275, n16276, n16277, n16278, n16279,
         n16280, n16281, n16282, n16283, n16284, n16285, n16286, n16287,
         n16288, n16289, n16290, n16291, n16292, n16293, n16294, n16295,
         n16296, n16297, n16298, n16299, n16300, n16301, n16302, n16303,
         n16304, n16305, n16306, n16307, n16308, n16309, n16310, n16311,
         n16312, n16313, n16314, n16315, n16316, n16317, n16318, n16319,
         n16320, n16321, n16322, n16323, n16324, n16325, n16326, n16327,
         n16328, n16329, n16330, n16331, n16332, n16333, n16334, n16335,
         n16336, n16337, n16338, n16339, n16340, n16341, n16342, n16343,
         n16344, n16345, n16346, n16347, n16348, n16349, n16350, n16351,
         n16352, n16353, n16354, n16355, n16356, n16357, n16358, n16359,
         n16360, n16361, n16362, n16363, n16364, n16365, n16366, n16367,
         n16368, n16369, n16370, n16371, n16372, n16373, n16374, n16375,
         n16376, n16377, n16378, n16379, n16380, n16381, n16382, n16383,
         n16384, n16385, n16386, n16387, n16388, n16389, n16390, n16391,
         n16392, n16393, n16394, n16395, n16396, n16397, n16398, n16399,
         n16400, n16401, n16402, n16403, n16404, n16405, n16406, n16407,
         n16408, n16409, n16410, n16411, n16412, n16413, n16414, n16415,
         n16416, n16417, n16418, n16419, n16420, n16421, n16422, n16423,
         n16424, n16425, n16426, n16427, n16428, n16429, n16430, n16431,
         n16432, n16433, n16434, n16435, n16436, n16437, n16438, n16439,
         n16440, n16441, n16442, n16443, n16444, n16445, n16446, n16447,
         n16448, n16449, n16450, n16451, n16452, n16453, n16454, n16455,
         n16456, n16457, n16458, n16459, n16460, n16461, n16462, n16463,
         n16464, n16465, n16466, n16467, n16468, n16469, n16470, n16471,
         n16472, n16473, n16474, n16475, n16476, n16477, n16478, n16479,
         n16480, n16481, n16482, n16483, n16484, n16485, n16486, n16487,
         n16488, n16489, n16490, n16491, n16492, n16493, n16494, n16495,
         n16496, n16497, n16498, n16499, n16500, n16501, n16502, n16503,
         n16504, n16505, n16506, n16507, n16508, n16509, n16510, n16511,
         n16512, n16513, n16514, n16515, n16516, n16517, n16518, n16519,
         n16520, n16521, n16522, n16523, n16524, n16525, n16526, n16527,
         n16528, n16529, n16530, n16531, n16532, n16533, n16534, n16535,
         n16536, n16537, n16538, n16539, n16540, n16541, n16542, n16543,
         n16544, n16545, n16546, n16547, n16548, n16549, n16550, n16551,
         n16552, n16553, n16554, n16555, n16556, n16557, n16558, n16559,
         n16560, n16561, n16562, n16563, n16564, n16565, n16566, n16567,
         n16568, n16569, n16570, n16571, n16572, n16573, n16574, n16575,
         n16576, n16577, n16578, n16579, n16580, n16581, n16582, n16583,
         n16584, n16585, n16586, n16587, n16588, n16589, n16590, n16591,
         n16592, n16593, n16594, n16595, n16596, n16597, n16598, n16599,
         n16600, n16601, n16602, n16603, n16604, n16605, n16606, n16607,
         n16608, n16609, n16610, n16611, n16612, n16613, n16614, n16615,
         n16616, n16617, n16618, n16619, n16620, n16621, n16622, n16623,
         n16624, n16625, n16626, n16627, n16628, n16629, n16630, n16631,
         n16632, n16633, n16634, n16635, n16636, n16637, n16638, n16639,
         n16640, n16641, n16642, n16643, n16644, n16645, n16646, n16647,
         n16648, n16649, n16650, n16651, n16652, n16653, n16654, n16655,
         n16656, n16657, n16658, n16659, n16660, n16661, n16662, n16663,
         n16664, n16665, n16666, n16667, n16668, n16669, n16670, n16671,
         n16672, n16673, n16674, n16675, n16676, n16677, n16678, n16679,
         n16680, n16681, n16682, n16683, n16684, n16685, n16686, n16687,
         n16688, n16689, n16690, n16691, n16692, n16693, n16694, n16695,
         n16696, n16697, n16698, n16699, n16700, n16701, n16702, n16703,
         n16704, n16705, n16706, n16707, n16708, n16709, n16710, n16711,
         n16712, n16713, n16714, n16715, n16716, n16717, n16718, n16719,
         n16720, n16721, n16722, n16723, n16724, n16725, n16726, n16727,
         n16728, n16729, n16730, n16731, n16732, n16733, n16734, n16735,
         n16736, n16737, n16738, n16739, n16740, n16741, n16742, n16743,
         n16744, n16745, n16746, n16747, n16748, n16749, n16750, n16751,
         n16752, n16753, n16754, n16755, n16756, n16757, n16758, n16759,
         n16760, n16761, n16762, n16763, n16764, n16765, n16766, n16767,
         n16768, n16769, n16770, n16771, n16772, n16773, n16774, n16775,
         n16776, n16777, n16778, n16779, n16780, n16781, n16782, n16783,
         n16784, n16785, n16786, n16787, n16788, n16789, n16790, n16791,
         n16792, n16793, n16794, n16795, n16796, n16797, n16798, n16799,
         n16800, n16801, n16802, n16803, n16804, n16805, n16806, n16807,
         n16808, n16809, n16810, n16811, n16812, n16813, n16814, n16815,
         n16816, n16817, n16818, n16819, n16820, n16821, n16822, n16823,
         n16824, n16825, n16826, n16827, n16828, n16829, n16830, n16831,
         n16832, n16833, n16834, n16835, n16836, n16837, n16838, n16839,
         n16840, n16841, n16842, n16843, n16844, n16845, n16846, n16847,
         n16848, n16849, n16850, n16851, n16852, n16853, n16854, n16855,
         n16856, n16857, n16858, n16859, n16860, n16861, n16862, n16863,
         n16864, n16865, n16866, n16867, n16868, n16869, n16870, n16871,
         n16872, n16873, n16874, n16875, n16876, n16877, n16878, n16879,
         n16880, n16881, n16882, n16883, n16884, n16885, n16886, n16887,
         n16888, n16889, n16890, n16891, n16892, n16893, n16894, n16895,
         n16896, n16897, n16898, n16899, n16900, n16901, n16902, n16903,
         n16904, n16905, n16906, n16907, n16908, n16909, n16910, n16911,
         n16912, n16913, n16914, n16915, n16916, n16917, n16918, n16919,
         n16920, n16921, n16922, n16923, n16924, n16925, n16926, n16927,
         n16928, n16929, n16930, n16931, n16932, n16933, n16934, n16935,
         n16936, n16937, n16938, n16939, n16940, n16941, n16942, n16943,
         n16944, n16945, n16946, n16947, n16948, n16949, n16950, n16951,
         n16952, n16953, n16954, n16955, n16956, n16957, n16958, n16959,
         n16960, n16961, n16962, n16963, n16964, n16965, n16966, n16967,
         n16968, n16969, n16970, n16971, n16972, n16973, n16974, n16975,
         n16976, n16977, n16978, n16979, n16980, n16981, n16982, n16983,
         n16984, n16985, n16986, n16987, n16988, n16989, n16990, n16991,
         n16992, n16993, n16994, n16995, n16996, n16997, n16998, n16999,
         n17000, n17001, n17002, n17003, n17004, n17005, n17006, n17007,
         n17008, n17009, n17010, n17011, n17012, n17013, n17014, n17015,
         n17016, n17017, n17018, n17019, n17020, n17021, n17022, n17023,
         n17024, n17025, n17026, n17027, n17028, n17029, n17030, n17031,
         n17032, n17033, n17034, n17035, n17036, n17037, n17038, n17039,
         n17040, n17041, n17042, n17043, n17044, n17045, n17046, n17047,
         n17048, n17049, n17050, n17051, n17052, n17053, n17054, n17055,
         n17056, n17057, n17058, n17059, n17060, n17061, n17062, n17063,
         n17064, n17065, n17066, n17067, n17068, n17069, n17070, n17071,
         n17072, n17073, n17074, n17075, n17076, n17077, n17078, n17079,
         n17080, n17081, n17082, n17083, n17084, n17085, n17086, n17087,
         n17088, n17089, n17090, n17091, n17092, n17093, n17094, n17095,
         n17096, n17097, n17098, n17099, n17100, n17101, n17102, n17103,
         n17104, n17105, n17106, n17107, n17108, n17109, n17110, n17111,
         n17112, n17113, n17114, n17115, n17116, n17117, n17118, n17119,
         n17120, n17121, n17122, n17123, n17124, n17125, n17126, n17127,
         n17128, n17129, n17130, n17131, n17132, n17133, n17134, n17135,
         n17136, n17137, n17138, n17139, n17140, n17141, n17142, n17143,
         n17144, n17145, n17146, n17147, n17148, n17149, n17150, n17151,
         n17152, n17153, n17154, n17155, n17156, n17157, n17158, n17159,
         n17160, n17161, n17162, n17163, n17164, n17165, n17166, n17167,
         n17168, n17169, n17170, n17171, n17172, n17173, n17174, n17175,
         n17176, n17177, n17178, n17179, n17180, n17181, n17182, n17183,
         n17184, n17185, n17186, n17187, n17188, n17189, n17190, n17191,
         n17192, n17193, n17194, n17195, n17196, n17197, n17198, n17199,
         n17200, n17201, n17202, n17203, n17204, n17205, n17206, n17207,
         n17208, n17209, n17210, n17211, n17212, n17213, n17214, n17215,
         n17216, n17217, n17218, n17219, n17220, n17221, n17222, n17223,
         n17224, n17225, n17226, n17227, n17228, n17229, n17230, n17231,
         n17232, n17233, n17234, n17235, n17236, n17237, n17238, n17239,
         n17240, n17241, n17242, n17243, n17244, n17245, n17246, n17247,
         n17248, n17249, n17250, n17251, n17252, n17253, n17254, n17255,
         n17256, n17257, n17258, n17259, n17260, n17261, n17262, n17263,
         n17264, n17265, n17266, n17267, n17268, n17269, n17270, n17271,
         n17272, n17273, n17274, n17275, n17276, n17277, n17278, n17279,
         n17280, n17281, n17282, n17283, n17284, n17285, n17286, n17287,
         n17288, n17289, n17290, n17291, n17292, n17293, n17294, n17295,
         n17296, n17297, n17298, n17299, n17300, n17301, n17302, n17303,
         n17304, n17305, n17306, n17307, n17308, n17309, n17310, n17311,
         n17312, n17313, n17314, n17315, n17316, n17317, n17318, n17319,
         n17320, n17321, n17322, n17323, n17324, n17325, n17326, n17327,
         n17328, n17329, n17330, n17331, n17332, n17333, n17334, n17335,
         n17336, n17337, n17338, n17339, n17340, n17341, n17342, n17343,
         n17344, n17345, n17346, n17347, n17348, n17349, n17350, n17351,
         n17352, n17353, n17354, n17355, n17356, n17357, n17358, n17359,
         n17360, n17361, n17362, n17363, n17364, n17365, n17366, n17367,
         n17368, n17369, n17370, n17371, n17372, n17373, n17374, n17375,
         n17376, n17377, n17378, n17379, n17380, n17381, n17382, n17383,
         n17384, n17385, n17386, n17387, n17388, n17389, n17390, n17391,
         n17392, n17393, n17394, n17395, n17396, n17397, n17398, n17399,
         n17400, n17401, n17402, n17403, n17404, n17405, n17406, n17407,
         n17408, n17409, n17410, n17411, n17412, n17413, n17414, n17415,
         n17416, n17417, n17418, n17419, n17420, n17421, n17422, n17423,
         n17424, n17425, n17426, n17427, n17428, n17429, n17430, n17431,
         n17432, n17433, n17434, n17435, n17436, n17437, n17438, n17439,
         n17440, n17441, n17442, n17443, n17444, n17445, n17446, n17447,
         n17448, n17449, n17450, n17451, n17452, n17453, n17454, n17455,
         n17456, n17457, n17458, n17459, n17460, n17461, n17462, n17463;

  XOR \SUBBYTES[0].a/U5649  ( .A(\SUBBYTES[0].a/w3390 ), .B(
        \SUBBYTES[0].a/w3391 ), .Z(\SUBBYTES[0].a/n1426 ) );
  XOR \SUBBYTES[0].a/U5648  ( .A(\SUBBYTES[0].a/n1426 ), .B(
        \SUBBYTES[0].a/n385 ), .Z(\SUBBYTES[0].a/n1425 ) );
  XOR \SUBBYTES[0].a/U5647  ( .A(\SUBBYTES[0].a/w3383 ), .B(
        \SUBBYTES[0].a/w3400 ), .Z(\SUBBYTES[0].a/n385 ) );
  XOR \SUBBYTES[0].a/U5645  ( .A(\SUBBYTES[0].a/w3382 ), .B(
        \SUBBYTES[0].a/w3397 ), .Z(\SUBBYTES[0].a/n386 ) );
  XOR \SUBBYTES[0].a/U5644  ( .A(\SUBBYTES[0].a/n1426 ), .B(
        \SUBBYTES[0].a/n387 ), .Z(\SUBBYTES[0].a/n1619 ) );
  XOR \SUBBYTES[0].a/U5643  ( .A(\SUBBYTES[0].a/w3397 ), .B(
        \SUBBYTES[0].a/w3398 ), .Z(\SUBBYTES[0].a/n387 ) );
  XOR \SUBBYTES[0].a/U5642  ( .A(\SUBBYTES[0].a/w3359 ), .B(
        \SUBBYTES[0].a/n388 ), .Z(\SUBBYTES[0].a/n1428 ) );
  XOR \SUBBYTES[0].a/U5641  ( .A(\SUBBYTES[0].a/w3350 ), .B(
        \SUBBYTES[0].a/w3351 ), .Z(\SUBBYTES[0].a/n388 ) );
  XOR \SUBBYTES[0].a/U5639  ( .A(\SUBBYTES[0].a/w3361 ), .B(
        \SUBBYTES[0].a/n1619 ), .Z(\SUBBYTES[0].a/n389 ) );
  XOR \SUBBYTES[0].a/U5638  ( .A(\SUBBYTES[0].a/n391 ), .B(
        \SUBBYTES[0].a/n390 ), .Z(\SUBBYTES[0].a/n1429 ) );
  XOR \SUBBYTES[0].a/U5637  ( .A(\SUBBYTES[0].a/n393 ), .B(
        \SUBBYTES[0].a/n392 ), .Z(\SUBBYTES[0].a/n390 ) );
  XOR \SUBBYTES[0].a/U5636  ( .A(\SUBBYTES[0].a/w3397 ), .B(
        \SUBBYTES[0].a/w3398 ), .Z(\SUBBYTES[0].a/n391 ) );
  XOR \SUBBYTES[0].a/U5635  ( .A(\SUBBYTES[0].a/w3361 ), .B(
        \SUBBYTES[0].a/w3385 ), .Z(\SUBBYTES[0].a/n392 ) );
  XOR \SUBBYTES[0].a/U5634  ( .A(\SUBBYTES[0].a/w3350 ), .B(
        \SUBBYTES[0].a/w3359 ), .Z(\SUBBYTES[0].a/n393 ) );
  XOR \SUBBYTES[0].a/U5633  ( .A(\SUBBYTES[0].a/w3382 ), .B(
        \SUBBYTES[0].a/n394 ), .Z(\SUBBYTES[0].a/n1427 ) );
  XOR \SUBBYTES[0].a/U5632  ( .A(\SUBBYTES[0].a/w3365 ), .B(
        \SUBBYTES[0].a/w3368 ), .Z(\SUBBYTES[0].a/n394 ) );
  XOR \SUBBYTES[0].a/U5630  ( .A(\SUBBYTES[0].a/w3353 ), .B(
        \SUBBYTES[0].a/n1429 ), .Z(\SUBBYTES[0].a/n395 ) );
  XOR \SUBBYTES[0].a/U5628  ( .A(\SUBBYTES[0].a/w3385 ), .B(
        \SUBBYTES[0].a/w3398 ), .Z(\SUBBYTES[0].a/n396 ) );
  XOR \SUBBYTES[0].a/U5626  ( .A(\SUBBYTES[0].a/n400 ), .B(
        \SUBBYTES[0].a/n399 ), .Z(\SUBBYTES[0].a/n397 ) );
  XOR \SUBBYTES[0].a/U5625  ( .A(\SUBBYTES[0].a/n402 ), .B(
        \SUBBYTES[0].a/n401 ), .Z(\SUBBYTES[0].a/n398 ) );
  XOR \SUBBYTES[0].a/U5624  ( .A(\SUBBYTES[0].a/w3397 ), .B(
        \SUBBYTES[0].a/w3400 ), .Z(\SUBBYTES[0].a/n399 ) );
  XOR \SUBBYTES[0].a/U5623  ( .A(\SUBBYTES[0].a/w3390 ), .B(
        \SUBBYTES[0].a/w3393 ), .Z(\SUBBYTES[0].a/n400 ) );
  XOR \SUBBYTES[0].a/U5622  ( .A(\SUBBYTES[0].a/w3365 ), .B(
        \SUBBYTES[0].a/w3366 ), .Z(\SUBBYTES[0].a/n401 ) );
  XOR \SUBBYTES[0].a/U5621  ( .A(\SUBBYTES[0].a/w3350 ), .B(
        \SUBBYTES[0].a/w3353 ), .Z(\SUBBYTES[0].a/n402 ) );
  XOR \SUBBYTES[0].a/U5619  ( .A(\SUBBYTES[0].a/n1426 ), .B(
        \SUBBYTES[0].a/n405 ), .Z(\SUBBYTES[0].a/n403 ) );
  XOR \SUBBYTES[0].a/U5618  ( .A(\SUBBYTES[0].a/n1428 ), .B(
        \SUBBYTES[0].a/n1427 ), .Z(\SUBBYTES[0].a/n404 ) );
  XOR \SUBBYTES[0].a/U5617  ( .A(\SUBBYTES[0].a/w3358 ), .B(
        \SUBBYTES[0].a/w3385 ), .Z(\SUBBYTES[0].a/n405 ) );
  XOR \SUBBYTES[0].a/U5615  ( .A(\SUBBYTES[0].a/n1429 ), .B(
        \SUBBYTES[0].a/n408 ), .Z(\SUBBYTES[0].a/n406 ) );
  XOR \SUBBYTES[0].a/U5614  ( .A(\SUBBYTES[0].a/w3391 ), .B(
        \SUBBYTES[0].a/w3393 ), .Z(\SUBBYTES[0].a/n407 ) );
  XOR \SUBBYTES[0].a/U5613  ( .A(\SUBBYTES[0].a/w3351 ), .B(
        \SUBBYTES[0].a/w3383 ), .Z(\SUBBYTES[0].a/n408 ) );
  XOR \SUBBYTES[0].a/U5612  ( .A(\SUBBYTES[0].a/w3183 ), .B(
        \SUBBYTES[0].a/w3184 ), .Z(\SUBBYTES[0].a/n1431 ) );
  XOR \SUBBYTES[0].a/U5611  ( .A(\SUBBYTES[0].a/n1431 ), .B(
        \SUBBYTES[0].a/n409 ), .Z(\SUBBYTES[0].a/n1430 ) );
  XOR \SUBBYTES[0].a/U5610  ( .A(\SUBBYTES[0].a/w3176 ), .B(
        \SUBBYTES[0].a/w3193 ), .Z(\SUBBYTES[0].a/n409 ) );
  XOR \SUBBYTES[0].a/U5608  ( .A(\SUBBYTES[0].a/w3175 ), .B(
        \SUBBYTES[0].a/w3190 ), .Z(\SUBBYTES[0].a/n410 ) );
  XOR \SUBBYTES[0].a/U5607  ( .A(\SUBBYTES[0].a/n1431 ), .B(
        \SUBBYTES[0].a/n411 ), .Z(\SUBBYTES[0].a/n1627 ) );
  XOR \SUBBYTES[0].a/U5606  ( .A(\SUBBYTES[0].a/w3190 ), .B(
        \SUBBYTES[0].a/w3191 ), .Z(\SUBBYTES[0].a/n411 ) );
  XOR \SUBBYTES[0].a/U5605  ( .A(\SUBBYTES[0].a/w3152 ), .B(
        \SUBBYTES[0].a/n412 ), .Z(\SUBBYTES[0].a/n1433 ) );
  XOR \SUBBYTES[0].a/U5604  ( .A(\SUBBYTES[0].a/w3143 ), .B(
        \SUBBYTES[0].a/w3144 ), .Z(\SUBBYTES[0].a/n412 ) );
  XOR \SUBBYTES[0].a/U5602  ( .A(\SUBBYTES[0].a/w3154 ), .B(
        \SUBBYTES[0].a/n1627 ), .Z(\SUBBYTES[0].a/n413 ) );
  XOR \SUBBYTES[0].a/U5601  ( .A(\SUBBYTES[0].a/n415 ), .B(
        \SUBBYTES[0].a/n414 ), .Z(\SUBBYTES[0].a/n1434 ) );
  XOR \SUBBYTES[0].a/U5600  ( .A(\SUBBYTES[0].a/n417 ), .B(
        \SUBBYTES[0].a/n416 ), .Z(\SUBBYTES[0].a/n414 ) );
  XOR \SUBBYTES[0].a/U5599  ( .A(\SUBBYTES[0].a/w3190 ), .B(
        \SUBBYTES[0].a/w3191 ), .Z(\SUBBYTES[0].a/n415 ) );
  XOR \SUBBYTES[0].a/U5598  ( .A(\SUBBYTES[0].a/w3154 ), .B(
        \SUBBYTES[0].a/w3178 ), .Z(\SUBBYTES[0].a/n416 ) );
  XOR \SUBBYTES[0].a/U5597  ( .A(\SUBBYTES[0].a/w3143 ), .B(
        \SUBBYTES[0].a/w3152 ), .Z(\SUBBYTES[0].a/n417 ) );
  XOR \SUBBYTES[0].a/U5596  ( .A(\SUBBYTES[0].a/w3175 ), .B(
        \SUBBYTES[0].a/n418 ), .Z(\SUBBYTES[0].a/n1432 ) );
  XOR \SUBBYTES[0].a/U5595  ( .A(\SUBBYTES[0].a/w3158 ), .B(
        \SUBBYTES[0].a/w3161 ), .Z(\SUBBYTES[0].a/n418 ) );
  XOR \SUBBYTES[0].a/U5593  ( .A(\SUBBYTES[0].a/w3146 ), .B(
        \SUBBYTES[0].a/n1434 ), .Z(\SUBBYTES[0].a/n419 ) );
  XOR \SUBBYTES[0].a/U5591  ( .A(\SUBBYTES[0].a/w3178 ), .B(
        \SUBBYTES[0].a/w3191 ), .Z(\SUBBYTES[0].a/n420 ) );
  XOR \SUBBYTES[0].a/U5589  ( .A(\SUBBYTES[0].a/n424 ), .B(
        \SUBBYTES[0].a/n423 ), .Z(\SUBBYTES[0].a/n421 ) );
  XOR \SUBBYTES[0].a/U5588  ( .A(\SUBBYTES[0].a/n426 ), .B(
        \SUBBYTES[0].a/n425 ), .Z(\SUBBYTES[0].a/n422 ) );
  XOR \SUBBYTES[0].a/U5587  ( .A(\SUBBYTES[0].a/w3190 ), .B(
        \SUBBYTES[0].a/w3193 ), .Z(\SUBBYTES[0].a/n423 ) );
  XOR \SUBBYTES[0].a/U5586  ( .A(\SUBBYTES[0].a/w3183 ), .B(
        \SUBBYTES[0].a/w3186 ), .Z(\SUBBYTES[0].a/n424 ) );
  XOR \SUBBYTES[0].a/U5585  ( .A(\SUBBYTES[0].a/w3158 ), .B(
        \SUBBYTES[0].a/w3159 ), .Z(\SUBBYTES[0].a/n425 ) );
  XOR \SUBBYTES[0].a/U5584  ( .A(\SUBBYTES[0].a/w3143 ), .B(
        \SUBBYTES[0].a/w3146 ), .Z(\SUBBYTES[0].a/n426 ) );
  XOR \SUBBYTES[0].a/U5582  ( .A(\SUBBYTES[0].a/n1431 ), .B(
        \SUBBYTES[0].a/n429 ), .Z(\SUBBYTES[0].a/n427 ) );
  XOR \SUBBYTES[0].a/U5581  ( .A(\SUBBYTES[0].a/n1433 ), .B(
        \SUBBYTES[0].a/n1432 ), .Z(\SUBBYTES[0].a/n428 ) );
  XOR \SUBBYTES[0].a/U5580  ( .A(\SUBBYTES[0].a/w3151 ), .B(
        \SUBBYTES[0].a/w3178 ), .Z(\SUBBYTES[0].a/n429 ) );
  XOR \SUBBYTES[0].a/U5578  ( .A(\SUBBYTES[0].a/n1434 ), .B(
        \SUBBYTES[0].a/n432 ), .Z(\SUBBYTES[0].a/n430 ) );
  XOR \SUBBYTES[0].a/U5577  ( .A(\SUBBYTES[0].a/w3184 ), .B(
        \SUBBYTES[0].a/w3186 ), .Z(\SUBBYTES[0].a/n431 ) );
  XOR \SUBBYTES[0].a/U5576  ( .A(\SUBBYTES[0].a/w3144 ), .B(
        \SUBBYTES[0].a/w3176 ), .Z(\SUBBYTES[0].a/n432 ) );
  XOR \SUBBYTES[0].a/U5575  ( .A(\SUBBYTES[0].a/w2976 ), .B(
        \SUBBYTES[0].a/w2977 ), .Z(\SUBBYTES[0].a/n1436 ) );
  XOR \SUBBYTES[0].a/U5574  ( .A(\SUBBYTES[0].a/n1436 ), .B(
        \SUBBYTES[0].a/n433 ), .Z(\SUBBYTES[0].a/n1435 ) );
  XOR \SUBBYTES[0].a/U5573  ( .A(\SUBBYTES[0].a/w2969 ), .B(
        \SUBBYTES[0].a/w2986 ), .Z(\SUBBYTES[0].a/n433 ) );
  XOR \SUBBYTES[0].a/U5571  ( .A(\SUBBYTES[0].a/w2968 ), .B(
        \SUBBYTES[0].a/w2983 ), .Z(\SUBBYTES[0].a/n434 ) );
  XOR \SUBBYTES[0].a/U5570  ( .A(\SUBBYTES[0].a/n1436 ), .B(
        \SUBBYTES[0].a/n435 ), .Z(\SUBBYTES[0].a/n1635 ) );
  XOR \SUBBYTES[0].a/U5569  ( .A(\SUBBYTES[0].a/w2983 ), .B(
        \SUBBYTES[0].a/w2984 ), .Z(\SUBBYTES[0].a/n435 ) );
  XOR \SUBBYTES[0].a/U5568  ( .A(\SUBBYTES[0].a/w2945 ), .B(
        \SUBBYTES[0].a/n436 ), .Z(\SUBBYTES[0].a/n1438 ) );
  XOR \SUBBYTES[0].a/U5567  ( .A(\SUBBYTES[0].a/w2936 ), .B(
        \SUBBYTES[0].a/w2937 ), .Z(\SUBBYTES[0].a/n436 ) );
  XOR \SUBBYTES[0].a/U5565  ( .A(\SUBBYTES[0].a/w2947 ), .B(
        \SUBBYTES[0].a/n1635 ), .Z(\SUBBYTES[0].a/n437 ) );
  XOR \SUBBYTES[0].a/U5564  ( .A(\SUBBYTES[0].a/n439 ), .B(
        \SUBBYTES[0].a/n438 ), .Z(\SUBBYTES[0].a/n1439 ) );
  XOR \SUBBYTES[0].a/U5563  ( .A(\SUBBYTES[0].a/n441 ), .B(
        \SUBBYTES[0].a/n440 ), .Z(\SUBBYTES[0].a/n438 ) );
  XOR \SUBBYTES[0].a/U5562  ( .A(\SUBBYTES[0].a/w2983 ), .B(
        \SUBBYTES[0].a/w2984 ), .Z(\SUBBYTES[0].a/n439 ) );
  XOR \SUBBYTES[0].a/U5561  ( .A(\SUBBYTES[0].a/w2947 ), .B(
        \SUBBYTES[0].a/w2971 ), .Z(\SUBBYTES[0].a/n440 ) );
  XOR \SUBBYTES[0].a/U5560  ( .A(\SUBBYTES[0].a/w2936 ), .B(
        \SUBBYTES[0].a/w2945 ), .Z(\SUBBYTES[0].a/n441 ) );
  XOR \SUBBYTES[0].a/U5559  ( .A(\SUBBYTES[0].a/w2968 ), .B(
        \SUBBYTES[0].a/n442 ), .Z(\SUBBYTES[0].a/n1437 ) );
  XOR \SUBBYTES[0].a/U5558  ( .A(\SUBBYTES[0].a/w2951 ), .B(
        \SUBBYTES[0].a/w2954 ), .Z(\SUBBYTES[0].a/n442 ) );
  XOR \SUBBYTES[0].a/U5556  ( .A(\SUBBYTES[0].a/w2939 ), .B(
        \SUBBYTES[0].a/n1439 ), .Z(\SUBBYTES[0].a/n443 ) );
  XOR \SUBBYTES[0].a/U5554  ( .A(\SUBBYTES[0].a/w2971 ), .B(
        \SUBBYTES[0].a/w2984 ), .Z(\SUBBYTES[0].a/n444 ) );
  XOR \SUBBYTES[0].a/U5552  ( .A(\SUBBYTES[0].a/n448 ), .B(
        \SUBBYTES[0].a/n447 ), .Z(\SUBBYTES[0].a/n445 ) );
  XOR \SUBBYTES[0].a/U5551  ( .A(\SUBBYTES[0].a/n450 ), .B(
        \SUBBYTES[0].a/n449 ), .Z(\SUBBYTES[0].a/n446 ) );
  XOR \SUBBYTES[0].a/U5550  ( .A(\SUBBYTES[0].a/w2983 ), .B(
        \SUBBYTES[0].a/w2986 ), .Z(\SUBBYTES[0].a/n447 ) );
  XOR \SUBBYTES[0].a/U5549  ( .A(\SUBBYTES[0].a/w2976 ), .B(
        \SUBBYTES[0].a/w2979 ), .Z(\SUBBYTES[0].a/n448 ) );
  XOR \SUBBYTES[0].a/U5548  ( .A(\SUBBYTES[0].a/w2951 ), .B(
        \SUBBYTES[0].a/w2952 ), .Z(\SUBBYTES[0].a/n449 ) );
  XOR \SUBBYTES[0].a/U5547  ( .A(\SUBBYTES[0].a/w2936 ), .B(
        \SUBBYTES[0].a/w2939 ), .Z(\SUBBYTES[0].a/n450 ) );
  XOR \SUBBYTES[0].a/U5545  ( .A(\SUBBYTES[0].a/n1436 ), .B(
        \SUBBYTES[0].a/n453 ), .Z(\SUBBYTES[0].a/n451 ) );
  XOR \SUBBYTES[0].a/U5544  ( .A(\SUBBYTES[0].a/n1438 ), .B(
        \SUBBYTES[0].a/n1437 ), .Z(\SUBBYTES[0].a/n452 ) );
  XOR \SUBBYTES[0].a/U5543  ( .A(\SUBBYTES[0].a/w2944 ), .B(
        \SUBBYTES[0].a/w2971 ), .Z(\SUBBYTES[0].a/n453 ) );
  XOR \SUBBYTES[0].a/U5541  ( .A(\SUBBYTES[0].a/n1439 ), .B(
        \SUBBYTES[0].a/n456 ), .Z(\SUBBYTES[0].a/n454 ) );
  XOR \SUBBYTES[0].a/U5540  ( .A(\SUBBYTES[0].a/w2977 ), .B(
        \SUBBYTES[0].a/w2979 ), .Z(\SUBBYTES[0].a/n455 ) );
  XOR \SUBBYTES[0].a/U5539  ( .A(\SUBBYTES[0].a/w2937 ), .B(
        \SUBBYTES[0].a/w2969 ), .Z(\SUBBYTES[0].a/n456 ) );
  XOR \SUBBYTES[0].a/U5538  ( .A(\SUBBYTES[0].a/w2769 ), .B(
        \SUBBYTES[0].a/w2770 ), .Z(\SUBBYTES[0].a/n1441 ) );
  XOR \SUBBYTES[0].a/U5537  ( .A(\SUBBYTES[0].a/n1441 ), .B(
        \SUBBYTES[0].a/n457 ), .Z(\SUBBYTES[0].a/n1440 ) );
  XOR \SUBBYTES[0].a/U5536  ( .A(\SUBBYTES[0].a/w2762 ), .B(
        \SUBBYTES[0].a/w2779 ), .Z(\SUBBYTES[0].a/n457 ) );
  XOR \SUBBYTES[0].a/U5534  ( .A(\SUBBYTES[0].a/w2761 ), .B(
        \SUBBYTES[0].a/w2776 ), .Z(\SUBBYTES[0].a/n458 ) );
  XOR \SUBBYTES[0].a/U5533  ( .A(\SUBBYTES[0].a/n1441 ), .B(
        \SUBBYTES[0].a/n459 ), .Z(\SUBBYTES[0].a/n1643 ) );
  XOR \SUBBYTES[0].a/U5532  ( .A(\SUBBYTES[0].a/w2776 ), .B(
        \SUBBYTES[0].a/w2777 ), .Z(\SUBBYTES[0].a/n459 ) );
  XOR \SUBBYTES[0].a/U5531  ( .A(\SUBBYTES[0].a/w2738 ), .B(
        \SUBBYTES[0].a/n460 ), .Z(\SUBBYTES[0].a/n1443 ) );
  XOR \SUBBYTES[0].a/U5530  ( .A(\SUBBYTES[0].a/w2729 ), .B(
        \SUBBYTES[0].a/w2730 ), .Z(\SUBBYTES[0].a/n460 ) );
  XOR \SUBBYTES[0].a/U5528  ( .A(\SUBBYTES[0].a/w2740 ), .B(
        \SUBBYTES[0].a/n1643 ), .Z(\SUBBYTES[0].a/n461 ) );
  XOR \SUBBYTES[0].a/U5527  ( .A(\SUBBYTES[0].a/n463 ), .B(
        \SUBBYTES[0].a/n462 ), .Z(\SUBBYTES[0].a/n1444 ) );
  XOR \SUBBYTES[0].a/U5526  ( .A(\SUBBYTES[0].a/n465 ), .B(
        \SUBBYTES[0].a/n464 ), .Z(\SUBBYTES[0].a/n462 ) );
  XOR \SUBBYTES[0].a/U5525  ( .A(\SUBBYTES[0].a/w2776 ), .B(
        \SUBBYTES[0].a/w2777 ), .Z(\SUBBYTES[0].a/n463 ) );
  XOR \SUBBYTES[0].a/U5524  ( .A(\SUBBYTES[0].a/w2740 ), .B(
        \SUBBYTES[0].a/w2764 ), .Z(\SUBBYTES[0].a/n464 ) );
  XOR \SUBBYTES[0].a/U5523  ( .A(\SUBBYTES[0].a/w2729 ), .B(
        \SUBBYTES[0].a/w2738 ), .Z(\SUBBYTES[0].a/n465 ) );
  XOR \SUBBYTES[0].a/U5522  ( .A(\SUBBYTES[0].a/w2761 ), .B(
        \SUBBYTES[0].a/n466 ), .Z(\SUBBYTES[0].a/n1442 ) );
  XOR \SUBBYTES[0].a/U5521  ( .A(\SUBBYTES[0].a/w2744 ), .B(
        \SUBBYTES[0].a/w2747 ), .Z(\SUBBYTES[0].a/n466 ) );
  XOR \SUBBYTES[0].a/U5519  ( .A(\SUBBYTES[0].a/w2732 ), .B(
        \SUBBYTES[0].a/n1444 ), .Z(\SUBBYTES[0].a/n467 ) );
  XOR \SUBBYTES[0].a/U5517  ( .A(\SUBBYTES[0].a/w2764 ), .B(
        \SUBBYTES[0].a/w2777 ), .Z(\SUBBYTES[0].a/n468 ) );
  XOR \SUBBYTES[0].a/U5515  ( .A(\SUBBYTES[0].a/n472 ), .B(
        \SUBBYTES[0].a/n471 ), .Z(\SUBBYTES[0].a/n469 ) );
  XOR \SUBBYTES[0].a/U5514  ( .A(\SUBBYTES[0].a/n474 ), .B(
        \SUBBYTES[0].a/n473 ), .Z(\SUBBYTES[0].a/n470 ) );
  XOR \SUBBYTES[0].a/U5513  ( .A(\SUBBYTES[0].a/w2776 ), .B(
        \SUBBYTES[0].a/w2779 ), .Z(\SUBBYTES[0].a/n471 ) );
  XOR \SUBBYTES[0].a/U5512  ( .A(\SUBBYTES[0].a/w2769 ), .B(
        \SUBBYTES[0].a/w2772 ), .Z(\SUBBYTES[0].a/n472 ) );
  XOR \SUBBYTES[0].a/U5511  ( .A(\SUBBYTES[0].a/w2744 ), .B(
        \SUBBYTES[0].a/w2745 ), .Z(\SUBBYTES[0].a/n473 ) );
  XOR \SUBBYTES[0].a/U5510  ( .A(\SUBBYTES[0].a/w2729 ), .B(
        \SUBBYTES[0].a/w2732 ), .Z(\SUBBYTES[0].a/n474 ) );
  XOR \SUBBYTES[0].a/U5508  ( .A(\SUBBYTES[0].a/n1441 ), .B(
        \SUBBYTES[0].a/n477 ), .Z(\SUBBYTES[0].a/n475 ) );
  XOR \SUBBYTES[0].a/U5507  ( .A(\SUBBYTES[0].a/n1443 ), .B(
        \SUBBYTES[0].a/n1442 ), .Z(\SUBBYTES[0].a/n476 ) );
  XOR \SUBBYTES[0].a/U5506  ( .A(\SUBBYTES[0].a/w2737 ), .B(
        \SUBBYTES[0].a/w2764 ), .Z(\SUBBYTES[0].a/n477 ) );
  XOR \SUBBYTES[0].a/U5504  ( .A(\SUBBYTES[0].a/n1444 ), .B(
        \SUBBYTES[0].a/n480 ), .Z(\SUBBYTES[0].a/n478 ) );
  XOR \SUBBYTES[0].a/U5503  ( .A(\SUBBYTES[0].a/w2770 ), .B(
        \SUBBYTES[0].a/w2772 ), .Z(\SUBBYTES[0].a/n479 ) );
  XOR \SUBBYTES[0].a/U5502  ( .A(\SUBBYTES[0].a/w2730 ), .B(
        \SUBBYTES[0].a/w2762 ), .Z(\SUBBYTES[0].a/n480 ) );
  XOR \SUBBYTES[0].a/U5501  ( .A(\SUBBYTES[0].a/w2562 ), .B(
        \SUBBYTES[0].a/w2563 ), .Z(\SUBBYTES[0].a/n1446 ) );
  XOR \SUBBYTES[0].a/U5500  ( .A(\SUBBYTES[0].a/n1446 ), .B(
        \SUBBYTES[0].a/n481 ), .Z(\SUBBYTES[0].a/n1445 ) );
  XOR \SUBBYTES[0].a/U5499  ( .A(\SUBBYTES[0].a/w2555 ), .B(
        \SUBBYTES[0].a/w2572 ), .Z(\SUBBYTES[0].a/n481 ) );
  XOR \SUBBYTES[0].a/U5497  ( .A(\SUBBYTES[0].a/w2554 ), .B(
        \SUBBYTES[0].a/w2569 ), .Z(\SUBBYTES[0].a/n482 ) );
  XOR \SUBBYTES[0].a/U5496  ( .A(\SUBBYTES[0].a/n1446 ), .B(
        \SUBBYTES[0].a/n483 ), .Z(\SUBBYTES[0].a/n1651 ) );
  XOR \SUBBYTES[0].a/U5495  ( .A(\SUBBYTES[0].a/w2569 ), .B(
        \SUBBYTES[0].a/w2570 ), .Z(\SUBBYTES[0].a/n483 ) );
  XOR \SUBBYTES[0].a/U5494  ( .A(\SUBBYTES[0].a/w2531 ), .B(
        \SUBBYTES[0].a/n484 ), .Z(\SUBBYTES[0].a/n1448 ) );
  XOR \SUBBYTES[0].a/U5493  ( .A(\SUBBYTES[0].a/w2522 ), .B(
        \SUBBYTES[0].a/w2523 ), .Z(\SUBBYTES[0].a/n484 ) );
  XOR \SUBBYTES[0].a/U5491  ( .A(\SUBBYTES[0].a/w2533 ), .B(
        \SUBBYTES[0].a/n1651 ), .Z(\SUBBYTES[0].a/n485 ) );
  XOR \SUBBYTES[0].a/U5490  ( .A(\SUBBYTES[0].a/n487 ), .B(
        \SUBBYTES[0].a/n486 ), .Z(\SUBBYTES[0].a/n1449 ) );
  XOR \SUBBYTES[0].a/U5489  ( .A(\SUBBYTES[0].a/n489 ), .B(
        \SUBBYTES[0].a/n488 ), .Z(\SUBBYTES[0].a/n486 ) );
  XOR \SUBBYTES[0].a/U5488  ( .A(\SUBBYTES[0].a/w2569 ), .B(
        \SUBBYTES[0].a/w2570 ), .Z(\SUBBYTES[0].a/n487 ) );
  XOR \SUBBYTES[0].a/U5487  ( .A(\SUBBYTES[0].a/w2533 ), .B(
        \SUBBYTES[0].a/w2557 ), .Z(\SUBBYTES[0].a/n488 ) );
  XOR \SUBBYTES[0].a/U5486  ( .A(\SUBBYTES[0].a/w2522 ), .B(
        \SUBBYTES[0].a/w2531 ), .Z(\SUBBYTES[0].a/n489 ) );
  XOR \SUBBYTES[0].a/U5485  ( .A(\SUBBYTES[0].a/w2554 ), .B(
        \SUBBYTES[0].a/n490 ), .Z(\SUBBYTES[0].a/n1447 ) );
  XOR \SUBBYTES[0].a/U5484  ( .A(\SUBBYTES[0].a/w2537 ), .B(
        \SUBBYTES[0].a/w2540 ), .Z(\SUBBYTES[0].a/n490 ) );
  XOR \SUBBYTES[0].a/U5482  ( .A(\SUBBYTES[0].a/w2525 ), .B(
        \SUBBYTES[0].a/n1449 ), .Z(\SUBBYTES[0].a/n491 ) );
  XOR \SUBBYTES[0].a/U5480  ( .A(\SUBBYTES[0].a/w2557 ), .B(
        \SUBBYTES[0].a/w2570 ), .Z(\SUBBYTES[0].a/n492 ) );
  XOR \SUBBYTES[0].a/U5478  ( .A(\SUBBYTES[0].a/n496 ), .B(
        \SUBBYTES[0].a/n495 ), .Z(\SUBBYTES[0].a/n493 ) );
  XOR \SUBBYTES[0].a/U5477  ( .A(\SUBBYTES[0].a/n498 ), .B(
        \SUBBYTES[0].a/n497 ), .Z(\SUBBYTES[0].a/n494 ) );
  XOR \SUBBYTES[0].a/U5476  ( .A(\SUBBYTES[0].a/w2569 ), .B(
        \SUBBYTES[0].a/w2572 ), .Z(\SUBBYTES[0].a/n495 ) );
  XOR \SUBBYTES[0].a/U5475  ( .A(\SUBBYTES[0].a/w2562 ), .B(
        \SUBBYTES[0].a/w2565 ), .Z(\SUBBYTES[0].a/n496 ) );
  XOR \SUBBYTES[0].a/U5474  ( .A(\SUBBYTES[0].a/w2537 ), .B(
        \SUBBYTES[0].a/w2538 ), .Z(\SUBBYTES[0].a/n497 ) );
  XOR \SUBBYTES[0].a/U5473  ( .A(\SUBBYTES[0].a/w2522 ), .B(
        \SUBBYTES[0].a/w2525 ), .Z(\SUBBYTES[0].a/n498 ) );
  XOR \SUBBYTES[0].a/U5471  ( .A(\SUBBYTES[0].a/n1446 ), .B(
        \SUBBYTES[0].a/n501 ), .Z(\SUBBYTES[0].a/n499 ) );
  XOR \SUBBYTES[0].a/U5470  ( .A(\SUBBYTES[0].a/n1448 ), .B(
        \SUBBYTES[0].a/n1447 ), .Z(\SUBBYTES[0].a/n500 ) );
  XOR \SUBBYTES[0].a/U5469  ( .A(\SUBBYTES[0].a/w2530 ), .B(
        \SUBBYTES[0].a/w2557 ), .Z(\SUBBYTES[0].a/n501 ) );
  XOR \SUBBYTES[0].a/U5467  ( .A(\SUBBYTES[0].a/n1449 ), .B(
        \SUBBYTES[0].a/n504 ), .Z(\SUBBYTES[0].a/n502 ) );
  XOR \SUBBYTES[0].a/U5466  ( .A(\SUBBYTES[0].a/w2563 ), .B(
        \SUBBYTES[0].a/w2565 ), .Z(\SUBBYTES[0].a/n503 ) );
  XOR \SUBBYTES[0].a/U5465  ( .A(\SUBBYTES[0].a/w2523 ), .B(
        \SUBBYTES[0].a/w2555 ), .Z(\SUBBYTES[0].a/n504 ) );
  XOR \SUBBYTES[0].a/U5464  ( .A(\SUBBYTES[0].a/w2355 ), .B(
        \SUBBYTES[0].a/w2356 ), .Z(\SUBBYTES[0].a/n1451 ) );
  XOR \SUBBYTES[0].a/U5463  ( .A(\SUBBYTES[0].a/n1451 ), .B(
        \SUBBYTES[0].a/n505 ), .Z(\SUBBYTES[0].a/n1450 ) );
  XOR \SUBBYTES[0].a/U5462  ( .A(\SUBBYTES[0].a/w2348 ), .B(
        \SUBBYTES[0].a/w2365 ), .Z(\SUBBYTES[0].a/n505 ) );
  XOR \SUBBYTES[0].a/U5460  ( .A(\SUBBYTES[0].a/w2347 ), .B(
        \SUBBYTES[0].a/w2362 ), .Z(\SUBBYTES[0].a/n506 ) );
  XOR \SUBBYTES[0].a/U5459  ( .A(\SUBBYTES[0].a/n1451 ), .B(
        \SUBBYTES[0].a/n507 ), .Z(\SUBBYTES[0].a/n1659 ) );
  XOR \SUBBYTES[0].a/U5458  ( .A(\SUBBYTES[0].a/w2362 ), .B(
        \SUBBYTES[0].a/w2363 ), .Z(\SUBBYTES[0].a/n507 ) );
  XOR \SUBBYTES[0].a/U5457  ( .A(\SUBBYTES[0].a/w2324 ), .B(
        \SUBBYTES[0].a/n508 ), .Z(\SUBBYTES[0].a/n1453 ) );
  XOR \SUBBYTES[0].a/U5456  ( .A(\SUBBYTES[0].a/w2315 ), .B(
        \SUBBYTES[0].a/w2316 ), .Z(\SUBBYTES[0].a/n508 ) );
  XOR \SUBBYTES[0].a/U5454  ( .A(\SUBBYTES[0].a/w2326 ), .B(
        \SUBBYTES[0].a/n1659 ), .Z(\SUBBYTES[0].a/n509 ) );
  XOR \SUBBYTES[0].a/U5453  ( .A(\SUBBYTES[0].a/n511 ), .B(
        \SUBBYTES[0].a/n510 ), .Z(\SUBBYTES[0].a/n1454 ) );
  XOR \SUBBYTES[0].a/U5452  ( .A(\SUBBYTES[0].a/n513 ), .B(
        \SUBBYTES[0].a/n512 ), .Z(\SUBBYTES[0].a/n510 ) );
  XOR \SUBBYTES[0].a/U5451  ( .A(\SUBBYTES[0].a/w2362 ), .B(
        \SUBBYTES[0].a/w2363 ), .Z(\SUBBYTES[0].a/n511 ) );
  XOR \SUBBYTES[0].a/U5450  ( .A(\SUBBYTES[0].a/w2326 ), .B(
        \SUBBYTES[0].a/w2350 ), .Z(\SUBBYTES[0].a/n512 ) );
  XOR \SUBBYTES[0].a/U5449  ( .A(\SUBBYTES[0].a/w2315 ), .B(
        \SUBBYTES[0].a/w2324 ), .Z(\SUBBYTES[0].a/n513 ) );
  XOR \SUBBYTES[0].a/U5448  ( .A(\SUBBYTES[0].a/w2347 ), .B(
        \SUBBYTES[0].a/n514 ), .Z(\SUBBYTES[0].a/n1452 ) );
  XOR \SUBBYTES[0].a/U5447  ( .A(\SUBBYTES[0].a/w2330 ), .B(
        \SUBBYTES[0].a/w2333 ), .Z(\SUBBYTES[0].a/n514 ) );
  XOR \SUBBYTES[0].a/U5445  ( .A(\SUBBYTES[0].a/w2318 ), .B(
        \SUBBYTES[0].a/n1454 ), .Z(\SUBBYTES[0].a/n515 ) );
  XOR \SUBBYTES[0].a/U5443  ( .A(\SUBBYTES[0].a/w2350 ), .B(
        \SUBBYTES[0].a/w2363 ), .Z(\SUBBYTES[0].a/n516 ) );
  XOR \SUBBYTES[0].a/U5441  ( .A(\SUBBYTES[0].a/n520 ), .B(
        \SUBBYTES[0].a/n519 ), .Z(\SUBBYTES[0].a/n517 ) );
  XOR \SUBBYTES[0].a/U5440  ( .A(\SUBBYTES[0].a/n522 ), .B(
        \SUBBYTES[0].a/n521 ), .Z(\SUBBYTES[0].a/n518 ) );
  XOR \SUBBYTES[0].a/U5439  ( .A(\SUBBYTES[0].a/w2362 ), .B(
        \SUBBYTES[0].a/w2365 ), .Z(\SUBBYTES[0].a/n519 ) );
  XOR \SUBBYTES[0].a/U5438  ( .A(\SUBBYTES[0].a/w2355 ), .B(
        \SUBBYTES[0].a/w2358 ), .Z(\SUBBYTES[0].a/n520 ) );
  XOR \SUBBYTES[0].a/U5437  ( .A(\SUBBYTES[0].a/w2330 ), .B(
        \SUBBYTES[0].a/w2331 ), .Z(\SUBBYTES[0].a/n521 ) );
  XOR \SUBBYTES[0].a/U5436  ( .A(\SUBBYTES[0].a/w2315 ), .B(
        \SUBBYTES[0].a/w2318 ), .Z(\SUBBYTES[0].a/n522 ) );
  XOR \SUBBYTES[0].a/U5434  ( .A(\SUBBYTES[0].a/n1451 ), .B(
        \SUBBYTES[0].a/n525 ), .Z(\SUBBYTES[0].a/n523 ) );
  XOR \SUBBYTES[0].a/U5433  ( .A(\SUBBYTES[0].a/n1453 ), .B(
        \SUBBYTES[0].a/n1452 ), .Z(\SUBBYTES[0].a/n524 ) );
  XOR \SUBBYTES[0].a/U5432  ( .A(\SUBBYTES[0].a/w2323 ), .B(
        \SUBBYTES[0].a/w2350 ), .Z(\SUBBYTES[0].a/n525 ) );
  XOR \SUBBYTES[0].a/U5430  ( .A(\SUBBYTES[0].a/n1454 ), .B(
        \SUBBYTES[0].a/n528 ), .Z(\SUBBYTES[0].a/n526 ) );
  XOR \SUBBYTES[0].a/U5429  ( .A(\SUBBYTES[0].a/w2356 ), .B(
        \SUBBYTES[0].a/w2358 ), .Z(\SUBBYTES[0].a/n527 ) );
  XOR \SUBBYTES[0].a/U5428  ( .A(\SUBBYTES[0].a/w2316 ), .B(
        \SUBBYTES[0].a/w2348 ), .Z(\SUBBYTES[0].a/n528 ) );
  XOR \SUBBYTES[0].a/U5427  ( .A(\SUBBYTES[0].a/w2148 ), .B(
        \SUBBYTES[0].a/w2149 ), .Z(\SUBBYTES[0].a/n1456 ) );
  XOR \SUBBYTES[0].a/U5426  ( .A(\SUBBYTES[0].a/n1456 ), .B(
        \SUBBYTES[0].a/n529 ), .Z(\SUBBYTES[0].a/n1455 ) );
  XOR \SUBBYTES[0].a/U5425  ( .A(\SUBBYTES[0].a/w2141 ), .B(
        \SUBBYTES[0].a/w2158 ), .Z(\SUBBYTES[0].a/n529 ) );
  XOR \SUBBYTES[0].a/U5423  ( .A(\SUBBYTES[0].a/w2140 ), .B(
        \SUBBYTES[0].a/w2155 ), .Z(\SUBBYTES[0].a/n530 ) );
  XOR \SUBBYTES[0].a/U5422  ( .A(\SUBBYTES[0].a/n1456 ), .B(
        \SUBBYTES[0].a/n531 ), .Z(\SUBBYTES[0].a/n1667 ) );
  XOR \SUBBYTES[0].a/U5421  ( .A(\SUBBYTES[0].a/w2155 ), .B(
        \SUBBYTES[0].a/w2156 ), .Z(\SUBBYTES[0].a/n531 ) );
  XOR \SUBBYTES[0].a/U5420  ( .A(\SUBBYTES[0].a/w2117 ), .B(
        \SUBBYTES[0].a/n532 ), .Z(\SUBBYTES[0].a/n1458 ) );
  XOR \SUBBYTES[0].a/U5419  ( .A(\SUBBYTES[0].a/w2108 ), .B(
        \SUBBYTES[0].a/w2109 ), .Z(\SUBBYTES[0].a/n532 ) );
  XOR \SUBBYTES[0].a/U5417  ( .A(\SUBBYTES[0].a/w2119 ), .B(
        \SUBBYTES[0].a/n1667 ), .Z(\SUBBYTES[0].a/n533 ) );
  XOR \SUBBYTES[0].a/U5416  ( .A(\SUBBYTES[0].a/n535 ), .B(
        \SUBBYTES[0].a/n534 ), .Z(\SUBBYTES[0].a/n1459 ) );
  XOR \SUBBYTES[0].a/U5415  ( .A(\SUBBYTES[0].a/n537 ), .B(
        \SUBBYTES[0].a/n536 ), .Z(\SUBBYTES[0].a/n534 ) );
  XOR \SUBBYTES[0].a/U5414  ( .A(\SUBBYTES[0].a/w2155 ), .B(
        \SUBBYTES[0].a/w2156 ), .Z(\SUBBYTES[0].a/n535 ) );
  XOR \SUBBYTES[0].a/U5413  ( .A(\SUBBYTES[0].a/w2119 ), .B(
        \SUBBYTES[0].a/w2143 ), .Z(\SUBBYTES[0].a/n536 ) );
  XOR \SUBBYTES[0].a/U5412  ( .A(\SUBBYTES[0].a/w2108 ), .B(
        \SUBBYTES[0].a/w2117 ), .Z(\SUBBYTES[0].a/n537 ) );
  XOR \SUBBYTES[0].a/U5411  ( .A(\SUBBYTES[0].a/w2140 ), .B(
        \SUBBYTES[0].a/n538 ), .Z(\SUBBYTES[0].a/n1457 ) );
  XOR \SUBBYTES[0].a/U5410  ( .A(\SUBBYTES[0].a/w2123 ), .B(
        \SUBBYTES[0].a/w2126 ), .Z(\SUBBYTES[0].a/n538 ) );
  XOR \SUBBYTES[0].a/U5408  ( .A(\SUBBYTES[0].a/w2111 ), .B(
        \SUBBYTES[0].a/n1459 ), .Z(\SUBBYTES[0].a/n539 ) );
  XOR \SUBBYTES[0].a/U5406  ( .A(\SUBBYTES[0].a/w2143 ), .B(
        \SUBBYTES[0].a/w2156 ), .Z(\SUBBYTES[0].a/n540 ) );
  XOR \SUBBYTES[0].a/U5404  ( .A(\SUBBYTES[0].a/n544 ), .B(
        \SUBBYTES[0].a/n543 ), .Z(\SUBBYTES[0].a/n541 ) );
  XOR \SUBBYTES[0].a/U5403  ( .A(\SUBBYTES[0].a/n546 ), .B(
        \SUBBYTES[0].a/n545 ), .Z(\SUBBYTES[0].a/n542 ) );
  XOR \SUBBYTES[0].a/U5402  ( .A(\SUBBYTES[0].a/w2155 ), .B(
        \SUBBYTES[0].a/w2158 ), .Z(\SUBBYTES[0].a/n543 ) );
  XOR \SUBBYTES[0].a/U5401  ( .A(\SUBBYTES[0].a/w2148 ), .B(
        \SUBBYTES[0].a/w2151 ), .Z(\SUBBYTES[0].a/n544 ) );
  XOR \SUBBYTES[0].a/U5400  ( .A(\SUBBYTES[0].a/w2123 ), .B(
        \SUBBYTES[0].a/w2124 ), .Z(\SUBBYTES[0].a/n545 ) );
  XOR \SUBBYTES[0].a/U5399  ( .A(\SUBBYTES[0].a/w2108 ), .B(
        \SUBBYTES[0].a/w2111 ), .Z(\SUBBYTES[0].a/n546 ) );
  XOR \SUBBYTES[0].a/U5397  ( .A(\SUBBYTES[0].a/n1456 ), .B(
        \SUBBYTES[0].a/n549 ), .Z(\SUBBYTES[0].a/n547 ) );
  XOR \SUBBYTES[0].a/U5396  ( .A(\SUBBYTES[0].a/n1458 ), .B(
        \SUBBYTES[0].a/n1457 ), .Z(\SUBBYTES[0].a/n548 ) );
  XOR \SUBBYTES[0].a/U5395  ( .A(\SUBBYTES[0].a/w2116 ), .B(
        \SUBBYTES[0].a/w2143 ), .Z(\SUBBYTES[0].a/n549 ) );
  XOR \SUBBYTES[0].a/U5393  ( .A(\SUBBYTES[0].a/n1459 ), .B(
        \SUBBYTES[0].a/n552 ), .Z(\SUBBYTES[0].a/n550 ) );
  XOR \SUBBYTES[0].a/U5392  ( .A(\SUBBYTES[0].a/w2149 ), .B(
        \SUBBYTES[0].a/w2151 ), .Z(\SUBBYTES[0].a/n551 ) );
  XOR \SUBBYTES[0].a/U5391  ( .A(\SUBBYTES[0].a/w2109 ), .B(
        \SUBBYTES[0].a/w2141 ), .Z(\SUBBYTES[0].a/n552 ) );
  XOR \SUBBYTES[0].a/U5390  ( .A(\SUBBYTES[0].a/w1941 ), .B(
        \SUBBYTES[0].a/w1942 ), .Z(\SUBBYTES[0].a/n1461 ) );
  XOR \SUBBYTES[0].a/U5389  ( .A(\SUBBYTES[0].a/n1461 ), .B(
        \SUBBYTES[0].a/n553 ), .Z(\SUBBYTES[0].a/n1460 ) );
  XOR \SUBBYTES[0].a/U5388  ( .A(\SUBBYTES[0].a/w1934 ), .B(
        \SUBBYTES[0].a/w1951 ), .Z(\SUBBYTES[0].a/n553 ) );
  XOR \SUBBYTES[0].a/U5386  ( .A(\SUBBYTES[0].a/w1933 ), .B(
        \SUBBYTES[0].a/w1948 ), .Z(\SUBBYTES[0].a/n554 ) );
  XOR \SUBBYTES[0].a/U5385  ( .A(\SUBBYTES[0].a/n1461 ), .B(
        \SUBBYTES[0].a/n555 ), .Z(\SUBBYTES[0].a/n1675 ) );
  XOR \SUBBYTES[0].a/U5384  ( .A(\SUBBYTES[0].a/w1948 ), .B(
        \SUBBYTES[0].a/w1949 ), .Z(\SUBBYTES[0].a/n555 ) );
  XOR \SUBBYTES[0].a/U5383  ( .A(\SUBBYTES[0].a/w1910 ), .B(
        \SUBBYTES[0].a/n556 ), .Z(\SUBBYTES[0].a/n1463 ) );
  XOR \SUBBYTES[0].a/U5382  ( .A(\SUBBYTES[0].a/w1901 ), .B(
        \SUBBYTES[0].a/w1902 ), .Z(\SUBBYTES[0].a/n556 ) );
  XOR \SUBBYTES[0].a/U5380  ( .A(\SUBBYTES[0].a/w1912 ), .B(
        \SUBBYTES[0].a/n1675 ), .Z(\SUBBYTES[0].a/n557 ) );
  XOR \SUBBYTES[0].a/U5379  ( .A(\SUBBYTES[0].a/n559 ), .B(
        \SUBBYTES[0].a/n558 ), .Z(\SUBBYTES[0].a/n1464 ) );
  XOR \SUBBYTES[0].a/U5378  ( .A(\SUBBYTES[0].a/n561 ), .B(
        \SUBBYTES[0].a/n560 ), .Z(\SUBBYTES[0].a/n558 ) );
  XOR \SUBBYTES[0].a/U5377  ( .A(\SUBBYTES[0].a/w1948 ), .B(
        \SUBBYTES[0].a/w1949 ), .Z(\SUBBYTES[0].a/n559 ) );
  XOR \SUBBYTES[0].a/U5376  ( .A(\SUBBYTES[0].a/w1912 ), .B(
        \SUBBYTES[0].a/w1936 ), .Z(\SUBBYTES[0].a/n560 ) );
  XOR \SUBBYTES[0].a/U5375  ( .A(\SUBBYTES[0].a/w1901 ), .B(
        \SUBBYTES[0].a/w1910 ), .Z(\SUBBYTES[0].a/n561 ) );
  XOR \SUBBYTES[0].a/U5374  ( .A(\SUBBYTES[0].a/w1933 ), .B(
        \SUBBYTES[0].a/n562 ), .Z(\SUBBYTES[0].a/n1462 ) );
  XOR \SUBBYTES[0].a/U5373  ( .A(\SUBBYTES[0].a/w1916 ), .B(
        \SUBBYTES[0].a/w1919 ), .Z(\SUBBYTES[0].a/n562 ) );
  XOR \SUBBYTES[0].a/U5371  ( .A(\SUBBYTES[0].a/w1904 ), .B(
        \SUBBYTES[0].a/n1464 ), .Z(\SUBBYTES[0].a/n563 ) );
  XOR \SUBBYTES[0].a/U5369  ( .A(\SUBBYTES[0].a/w1936 ), .B(
        \SUBBYTES[0].a/w1949 ), .Z(\SUBBYTES[0].a/n564 ) );
  XOR \SUBBYTES[0].a/U5367  ( .A(\SUBBYTES[0].a/n568 ), .B(
        \SUBBYTES[0].a/n567 ), .Z(\SUBBYTES[0].a/n565 ) );
  XOR \SUBBYTES[0].a/U5366  ( .A(\SUBBYTES[0].a/n570 ), .B(
        \SUBBYTES[0].a/n569 ), .Z(\SUBBYTES[0].a/n566 ) );
  XOR \SUBBYTES[0].a/U5365  ( .A(\SUBBYTES[0].a/w1948 ), .B(
        \SUBBYTES[0].a/w1951 ), .Z(\SUBBYTES[0].a/n567 ) );
  XOR \SUBBYTES[0].a/U5364  ( .A(\SUBBYTES[0].a/w1941 ), .B(
        \SUBBYTES[0].a/w1944 ), .Z(\SUBBYTES[0].a/n568 ) );
  XOR \SUBBYTES[0].a/U5363  ( .A(\SUBBYTES[0].a/w1916 ), .B(
        \SUBBYTES[0].a/w1917 ), .Z(\SUBBYTES[0].a/n569 ) );
  XOR \SUBBYTES[0].a/U5362  ( .A(\SUBBYTES[0].a/w1901 ), .B(
        \SUBBYTES[0].a/w1904 ), .Z(\SUBBYTES[0].a/n570 ) );
  XOR \SUBBYTES[0].a/U5360  ( .A(\SUBBYTES[0].a/n1461 ), .B(
        \SUBBYTES[0].a/n573 ), .Z(\SUBBYTES[0].a/n571 ) );
  XOR \SUBBYTES[0].a/U5359  ( .A(\SUBBYTES[0].a/n1463 ), .B(
        \SUBBYTES[0].a/n1462 ), .Z(\SUBBYTES[0].a/n572 ) );
  XOR \SUBBYTES[0].a/U5358  ( .A(\SUBBYTES[0].a/w1909 ), .B(
        \SUBBYTES[0].a/w1936 ), .Z(\SUBBYTES[0].a/n573 ) );
  XOR \SUBBYTES[0].a/U5356  ( .A(\SUBBYTES[0].a/n1464 ), .B(
        \SUBBYTES[0].a/n576 ), .Z(\SUBBYTES[0].a/n574 ) );
  XOR \SUBBYTES[0].a/U5355  ( .A(\SUBBYTES[0].a/w1942 ), .B(
        \SUBBYTES[0].a/w1944 ), .Z(\SUBBYTES[0].a/n575 ) );
  XOR \SUBBYTES[0].a/U5354  ( .A(\SUBBYTES[0].a/w1902 ), .B(
        \SUBBYTES[0].a/w1934 ), .Z(\SUBBYTES[0].a/n576 ) );
  XOR \SUBBYTES[0].a/U5353  ( .A(\SUBBYTES[0].a/w1734 ), .B(
        \SUBBYTES[0].a/w1735 ), .Z(\SUBBYTES[0].a/n1466 ) );
  XOR \SUBBYTES[0].a/U5352  ( .A(\SUBBYTES[0].a/n1466 ), .B(
        \SUBBYTES[0].a/n577 ), .Z(\SUBBYTES[0].a/n1465 ) );
  XOR \SUBBYTES[0].a/U5351  ( .A(\SUBBYTES[0].a/w1727 ), .B(
        \SUBBYTES[0].a/w1744 ), .Z(\SUBBYTES[0].a/n577 ) );
  XOR \SUBBYTES[0].a/U5349  ( .A(\SUBBYTES[0].a/w1726 ), .B(
        \SUBBYTES[0].a/w1741 ), .Z(\SUBBYTES[0].a/n578 ) );
  XOR \SUBBYTES[0].a/U5348  ( .A(\SUBBYTES[0].a/n1466 ), .B(
        \SUBBYTES[0].a/n579 ), .Z(\SUBBYTES[0].a/n1683 ) );
  XOR \SUBBYTES[0].a/U5347  ( .A(\SUBBYTES[0].a/w1741 ), .B(
        \SUBBYTES[0].a/w1742 ), .Z(\SUBBYTES[0].a/n579 ) );
  XOR \SUBBYTES[0].a/U5346  ( .A(\SUBBYTES[0].a/w1703 ), .B(
        \SUBBYTES[0].a/n580 ), .Z(\SUBBYTES[0].a/n1468 ) );
  XOR \SUBBYTES[0].a/U5345  ( .A(\SUBBYTES[0].a/w1694 ), .B(
        \SUBBYTES[0].a/w1695 ), .Z(\SUBBYTES[0].a/n580 ) );
  XOR \SUBBYTES[0].a/U5343  ( .A(\SUBBYTES[0].a/w1705 ), .B(
        \SUBBYTES[0].a/n1683 ), .Z(\SUBBYTES[0].a/n581 ) );
  XOR \SUBBYTES[0].a/U5342  ( .A(\SUBBYTES[0].a/n583 ), .B(
        \SUBBYTES[0].a/n582 ), .Z(\SUBBYTES[0].a/n1469 ) );
  XOR \SUBBYTES[0].a/U5341  ( .A(\SUBBYTES[0].a/n585 ), .B(
        \SUBBYTES[0].a/n584 ), .Z(\SUBBYTES[0].a/n582 ) );
  XOR \SUBBYTES[0].a/U5340  ( .A(\SUBBYTES[0].a/w1741 ), .B(
        \SUBBYTES[0].a/w1742 ), .Z(\SUBBYTES[0].a/n583 ) );
  XOR \SUBBYTES[0].a/U5339  ( .A(\SUBBYTES[0].a/w1705 ), .B(
        \SUBBYTES[0].a/w1729 ), .Z(\SUBBYTES[0].a/n584 ) );
  XOR \SUBBYTES[0].a/U5338  ( .A(\SUBBYTES[0].a/w1694 ), .B(
        \SUBBYTES[0].a/w1703 ), .Z(\SUBBYTES[0].a/n585 ) );
  XOR \SUBBYTES[0].a/U5337  ( .A(\SUBBYTES[0].a/w1726 ), .B(
        \SUBBYTES[0].a/n586 ), .Z(\SUBBYTES[0].a/n1467 ) );
  XOR \SUBBYTES[0].a/U5336  ( .A(\SUBBYTES[0].a/w1709 ), .B(
        \SUBBYTES[0].a/w1712 ), .Z(\SUBBYTES[0].a/n586 ) );
  XOR \SUBBYTES[0].a/U5334  ( .A(\SUBBYTES[0].a/w1697 ), .B(
        \SUBBYTES[0].a/n1469 ), .Z(\SUBBYTES[0].a/n587 ) );
  XOR \SUBBYTES[0].a/U5332  ( .A(\SUBBYTES[0].a/w1729 ), .B(
        \SUBBYTES[0].a/w1742 ), .Z(\SUBBYTES[0].a/n588 ) );
  XOR \SUBBYTES[0].a/U5330  ( .A(\SUBBYTES[0].a/n592 ), .B(
        \SUBBYTES[0].a/n591 ), .Z(\SUBBYTES[0].a/n589 ) );
  XOR \SUBBYTES[0].a/U5329  ( .A(\SUBBYTES[0].a/n594 ), .B(
        \SUBBYTES[0].a/n593 ), .Z(\SUBBYTES[0].a/n590 ) );
  XOR \SUBBYTES[0].a/U5328  ( .A(\SUBBYTES[0].a/w1741 ), .B(
        \SUBBYTES[0].a/w1744 ), .Z(\SUBBYTES[0].a/n591 ) );
  XOR \SUBBYTES[0].a/U5327  ( .A(\SUBBYTES[0].a/w1734 ), .B(
        \SUBBYTES[0].a/w1737 ), .Z(\SUBBYTES[0].a/n592 ) );
  XOR \SUBBYTES[0].a/U5326  ( .A(\SUBBYTES[0].a/w1709 ), .B(
        \SUBBYTES[0].a/w1710 ), .Z(\SUBBYTES[0].a/n593 ) );
  XOR \SUBBYTES[0].a/U5325  ( .A(\SUBBYTES[0].a/w1694 ), .B(
        \SUBBYTES[0].a/w1697 ), .Z(\SUBBYTES[0].a/n594 ) );
  XOR \SUBBYTES[0].a/U5323  ( .A(\SUBBYTES[0].a/n1466 ), .B(
        \SUBBYTES[0].a/n597 ), .Z(\SUBBYTES[0].a/n595 ) );
  XOR \SUBBYTES[0].a/U5322  ( .A(\SUBBYTES[0].a/n1468 ), .B(
        \SUBBYTES[0].a/n1467 ), .Z(\SUBBYTES[0].a/n596 ) );
  XOR \SUBBYTES[0].a/U5321  ( .A(\SUBBYTES[0].a/w1702 ), .B(
        \SUBBYTES[0].a/w1729 ), .Z(\SUBBYTES[0].a/n597 ) );
  XOR \SUBBYTES[0].a/U5319  ( .A(\SUBBYTES[0].a/n1469 ), .B(
        \SUBBYTES[0].a/n600 ), .Z(\SUBBYTES[0].a/n598 ) );
  XOR \SUBBYTES[0].a/U5318  ( .A(\SUBBYTES[0].a/w1735 ), .B(
        \SUBBYTES[0].a/w1737 ), .Z(\SUBBYTES[0].a/n599 ) );
  XOR \SUBBYTES[0].a/U5317  ( .A(\SUBBYTES[0].a/w1695 ), .B(
        \SUBBYTES[0].a/w1727 ), .Z(\SUBBYTES[0].a/n600 ) );
  XOR \SUBBYTES[0].a/U5316  ( .A(\SUBBYTES[0].a/w1527 ), .B(
        \SUBBYTES[0].a/w1528 ), .Z(\SUBBYTES[0].a/n1471 ) );
  XOR \SUBBYTES[0].a/U5315  ( .A(\SUBBYTES[0].a/n1471 ), .B(
        \SUBBYTES[0].a/n601 ), .Z(\SUBBYTES[0].a/n1470 ) );
  XOR \SUBBYTES[0].a/U5314  ( .A(\SUBBYTES[0].a/w1520 ), .B(
        \SUBBYTES[0].a/w1537 ), .Z(\SUBBYTES[0].a/n601 ) );
  XOR \SUBBYTES[0].a/U5312  ( .A(\SUBBYTES[0].a/w1519 ), .B(
        \SUBBYTES[0].a/w1534 ), .Z(\SUBBYTES[0].a/n602 ) );
  XOR \SUBBYTES[0].a/U5311  ( .A(\SUBBYTES[0].a/n1471 ), .B(
        \SUBBYTES[0].a/n603 ), .Z(\SUBBYTES[0].a/n1691 ) );
  XOR \SUBBYTES[0].a/U5310  ( .A(\SUBBYTES[0].a/w1534 ), .B(
        \SUBBYTES[0].a/w1535 ), .Z(\SUBBYTES[0].a/n603 ) );
  XOR \SUBBYTES[0].a/U5309  ( .A(\SUBBYTES[0].a/w1496 ), .B(
        \SUBBYTES[0].a/n604 ), .Z(\SUBBYTES[0].a/n1473 ) );
  XOR \SUBBYTES[0].a/U5308  ( .A(\SUBBYTES[0].a/w1487 ), .B(
        \SUBBYTES[0].a/w1488 ), .Z(\SUBBYTES[0].a/n604 ) );
  XOR \SUBBYTES[0].a/U5306  ( .A(\SUBBYTES[0].a/w1498 ), .B(
        \SUBBYTES[0].a/n1691 ), .Z(\SUBBYTES[0].a/n605 ) );
  XOR \SUBBYTES[0].a/U5305  ( .A(\SUBBYTES[0].a/n607 ), .B(
        \SUBBYTES[0].a/n606 ), .Z(\SUBBYTES[0].a/n1474 ) );
  XOR \SUBBYTES[0].a/U5304  ( .A(\SUBBYTES[0].a/n609 ), .B(
        \SUBBYTES[0].a/n608 ), .Z(\SUBBYTES[0].a/n606 ) );
  XOR \SUBBYTES[0].a/U5303  ( .A(\SUBBYTES[0].a/w1534 ), .B(
        \SUBBYTES[0].a/w1535 ), .Z(\SUBBYTES[0].a/n607 ) );
  XOR \SUBBYTES[0].a/U5302  ( .A(\SUBBYTES[0].a/w1498 ), .B(
        \SUBBYTES[0].a/w1522 ), .Z(\SUBBYTES[0].a/n608 ) );
  XOR \SUBBYTES[0].a/U5301  ( .A(\SUBBYTES[0].a/w1487 ), .B(
        \SUBBYTES[0].a/w1496 ), .Z(\SUBBYTES[0].a/n609 ) );
  XOR \SUBBYTES[0].a/U5300  ( .A(\SUBBYTES[0].a/w1519 ), .B(
        \SUBBYTES[0].a/n610 ), .Z(\SUBBYTES[0].a/n1472 ) );
  XOR \SUBBYTES[0].a/U5299  ( .A(\SUBBYTES[0].a/w1502 ), .B(
        \SUBBYTES[0].a/w1505 ), .Z(\SUBBYTES[0].a/n610 ) );
  XOR \SUBBYTES[0].a/U5297  ( .A(\SUBBYTES[0].a/w1490 ), .B(
        \SUBBYTES[0].a/n1474 ), .Z(\SUBBYTES[0].a/n611 ) );
  XOR \SUBBYTES[0].a/U5295  ( .A(\SUBBYTES[0].a/w1522 ), .B(
        \SUBBYTES[0].a/w1535 ), .Z(\SUBBYTES[0].a/n612 ) );
  XOR \SUBBYTES[0].a/U5293  ( .A(\SUBBYTES[0].a/n616 ), .B(
        \SUBBYTES[0].a/n615 ), .Z(\SUBBYTES[0].a/n613 ) );
  XOR \SUBBYTES[0].a/U5292  ( .A(\SUBBYTES[0].a/n618 ), .B(
        \SUBBYTES[0].a/n617 ), .Z(\SUBBYTES[0].a/n614 ) );
  XOR \SUBBYTES[0].a/U5291  ( .A(\SUBBYTES[0].a/w1534 ), .B(
        \SUBBYTES[0].a/w1537 ), .Z(\SUBBYTES[0].a/n615 ) );
  XOR \SUBBYTES[0].a/U5290  ( .A(\SUBBYTES[0].a/w1527 ), .B(
        \SUBBYTES[0].a/w1530 ), .Z(\SUBBYTES[0].a/n616 ) );
  XOR \SUBBYTES[0].a/U5289  ( .A(\SUBBYTES[0].a/w1502 ), .B(
        \SUBBYTES[0].a/w1503 ), .Z(\SUBBYTES[0].a/n617 ) );
  XOR \SUBBYTES[0].a/U5288  ( .A(\SUBBYTES[0].a/w1487 ), .B(
        \SUBBYTES[0].a/w1490 ), .Z(\SUBBYTES[0].a/n618 ) );
  XOR \SUBBYTES[0].a/U5286  ( .A(\SUBBYTES[0].a/n1471 ), .B(
        \SUBBYTES[0].a/n621 ), .Z(\SUBBYTES[0].a/n619 ) );
  XOR \SUBBYTES[0].a/U5285  ( .A(\SUBBYTES[0].a/n1473 ), .B(
        \SUBBYTES[0].a/n1472 ), .Z(\SUBBYTES[0].a/n620 ) );
  XOR \SUBBYTES[0].a/U5284  ( .A(\SUBBYTES[0].a/w1495 ), .B(
        \SUBBYTES[0].a/w1522 ), .Z(\SUBBYTES[0].a/n621 ) );
  XOR \SUBBYTES[0].a/U5282  ( .A(\SUBBYTES[0].a/n1474 ), .B(
        \SUBBYTES[0].a/n624 ), .Z(\SUBBYTES[0].a/n622 ) );
  XOR \SUBBYTES[0].a/U5281  ( .A(\SUBBYTES[0].a/w1528 ), .B(
        \SUBBYTES[0].a/w1530 ), .Z(\SUBBYTES[0].a/n623 ) );
  XOR \SUBBYTES[0].a/U5280  ( .A(\SUBBYTES[0].a/w1488 ), .B(
        \SUBBYTES[0].a/w1520 ), .Z(\SUBBYTES[0].a/n624 ) );
  XOR \SUBBYTES[0].a/U5279  ( .A(\SUBBYTES[0].a/w1320 ), .B(
        \SUBBYTES[0].a/w1321 ), .Z(\SUBBYTES[0].a/n1476 ) );
  XOR \SUBBYTES[0].a/U5278  ( .A(\SUBBYTES[0].a/n1476 ), .B(
        \SUBBYTES[0].a/n625 ), .Z(\SUBBYTES[0].a/n1475 ) );
  XOR \SUBBYTES[0].a/U5277  ( .A(\SUBBYTES[0].a/w1313 ), .B(
        \SUBBYTES[0].a/w1330 ), .Z(\SUBBYTES[0].a/n625 ) );
  XOR \SUBBYTES[0].a/U5275  ( .A(\SUBBYTES[0].a/w1312 ), .B(
        \SUBBYTES[0].a/w1327 ), .Z(\SUBBYTES[0].a/n626 ) );
  XOR \SUBBYTES[0].a/U5274  ( .A(\SUBBYTES[0].a/n1476 ), .B(
        \SUBBYTES[0].a/n627 ), .Z(\SUBBYTES[0].a/n1699 ) );
  XOR \SUBBYTES[0].a/U5273  ( .A(\SUBBYTES[0].a/w1327 ), .B(
        \SUBBYTES[0].a/w1328 ), .Z(\SUBBYTES[0].a/n627 ) );
  XOR \SUBBYTES[0].a/U5272  ( .A(\SUBBYTES[0].a/w1289 ), .B(
        \SUBBYTES[0].a/n628 ), .Z(\SUBBYTES[0].a/n1478 ) );
  XOR \SUBBYTES[0].a/U5271  ( .A(\SUBBYTES[0].a/w1280 ), .B(
        \SUBBYTES[0].a/w1281 ), .Z(\SUBBYTES[0].a/n628 ) );
  XOR \SUBBYTES[0].a/U5269  ( .A(\SUBBYTES[0].a/w1291 ), .B(
        \SUBBYTES[0].a/n1699 ), .Z(\SUBBYTES[0].a/n629 ) );
  XOR \SUBBYTES[0].a/U5268  ( .A(\SUBBYTES[0].a/n631 ), .B(
        \SUBBYTES[0].a/n630 ), .Z(\SUBBYTES[0].a/n1479 ) );
  XOR \SUBBYTES[0].a/U5267  ( .A(\SUBBYTES[0].a/n633 ), .B(
        \SUBBYTES[0].a/n632 ), .Z(\SUBBYTES[0].a/n630 ) );
  XOR \SUBBYTES[0].a/U5266  ( .A(\SUBBYTES[0].a/w1327 ), .B(
        \SUBBYTES[0].a/w1328 ), .Z(\SUBBYTES[0].a/n631 ) );
  XOR \SUBBYTES[0].a/U5265  ( .A(\SUBBYTES[0].a/w1291 ), .B(
        \SUBBYTES[0].a/w1315 ), .Z(\SUBBYTES[0].a/n632 ) );
  XOR \SUBBYTES[0].a/U5264  ( .A(\SUBBYTES[0].a/w1280 ), .B(
        \SUBBYTES[0].a/w1289 ), .Z(\SUBBYTES[0].a/n633 ) );
  XOR \SUBBYTES[0].a/U5263  ( .A(\SUBBYTES[0].a/w1312 ), .B(
        \SUBBYTES[0].a/n634 ), .Z(\SUBBYTES[0].a/n1477 ) );
  XOR \SUBBYTES[0].a/U5262  ( .A(\SUBBYTES[0].a/w1295 ), .B(
        \SUBBYTES[0].a/w1298 ), .Z(\SUBBYTES[0].a/n634 ) );
  XOR \SUBBYTES[0].a/U5260  ( .A(\SUBBYTES[0].a/w1283 ), .B(
        \SUBBYTES[0].a/n1479 ), .Z(\SUBBYTES[0].a/n635 ) );
  XOR \SUBBYTES[0].a/U5258  ( .A(\SUBBYTES[0].a/w1315 ), .B(
        \SUBBYTES[0].a/w1328 ), .Z(\SUBBYTES[0].a/n636 ) );
  XOR \SUBBYTES[0].a/U5256  ( .A(\SUBBYTES[0].a/n640 ), .B(
        \SUBBYTES[0].a/n639 ), .Z(\SUBBYTES[0].a/n637 ) );
  XOR \SUBBYTES[0].a/U5255  ( .A(\SUBBYTES[0].a/n642 ), .B(
        \SUBBYTES[0].a/n641 ), .Z(\SUBBYTES[0].a/n638 ) );
  XOR \SUBBYTES[0].a/U5254  ( .A(\SUBBYTES[0].a/w1327 ), .B(
        \SUBBYTES[0].a/w1330 ), .Z(\SUBBYTES[0].a/n639 ) );
  XOR \SUBBYTES[0].a/U5253  ( .A(\SUBBYTES[0].a/w1320 ), .B(
        \SUBBYTES[0].a/w1323 ), .Z(\SUBBYTES[0].a/n640 ) );
  XOR \SUBBYTES[0].a/U5252  ( .A(\SUBBYTES[0].a/w1295 ), .B(
        \SUBBYTES[0].a/w1296 ), .Z(\SUBBYTES[0].a/n641 ) );
  XOR \SUBBYTES[0].a/U5251  ( .A(\SUBBYTES[0].a/w1280 ), .B(
        \SUBBYTES[0].a/w1283 ), .Z(\SUBBYTES[0].a/n642 ) );
  XOR \SUBBYTES[0].a/U5249  ( .A(\SUBBYTES[0].a/n1476 ), .B(
        \SUBBYTES[0].a/n645 ), .Z(\SUBBYTES[0].a/n643 ) );
  XOR \SUBBYTES[0].a/U5248  ( .A(\SUBBYTES[0].a/n1478 ), .B(
        \SUBBYTES[0].a/n1477 ), .Z(\SUBBYTES[0].a/n644 ) );
  XOR \SUBBYTES[0].a/U5247  ( .A(\SUBBYTES[0].a/w1288 ), .B(
        \SUBBYTES[0].a/w1315 ), .Z(\SUBBYTES[0].a/n645 ) );
  XOR \SUBBYTES[0].a/U5245  ( .A(\SUBBYTES[0].a/n1479 ), .B(
        \SUBBYTES[0].a/n648 ), .Z(\SUBBYTES[0].a/n646 ) );
  XOR \SUBBYTES[0].a/U5244  ( .A(\SUBBYTES[0].a/w1321 ), .B(
        \SUBBYTES[0].a/w1323 ), .Z(\SUBBYTES[0].a/n647 ) );
  XOR \SUBBYTES[0].a/U5243  ( .A(\SUBBYTES[0].a/w1281 ), .B(
        \SUBBYTES[0].a/w1313 ), .Z(\SUBBYTES[0].a/n648 ) );
  XOR \SUBBYTES[0].a/U5242  ( .A(\SUBBYTES[0].a/w1113 ), .B(
        \SUBBYTES[0].a/w1114 ), .Z(\SUBBYTES[0].a/n1481 ) );
  XOR \SUBBYTES[0].a/U5241  ( .A(\SUBBYTES[0].a/n1481 ), .B(
        \SUBBYTES[0].a/n649 ), .Z(\SUBBYTES[0].a/n1480 ) );
  XOR \SUBBYTES[0].a/U5240  ( .A(\SUBBYTES[0].a/w1106 ), .B(
        \SUBBYTES[0].a/w1123 ), .Z(\SUBBYTES[0].a/n649 ) );
  XOR \SUBBYTES[0].a/U5238  ( .A(\SUBBYTES[0].a/w1105 ), .B(
        \SUBBYTES[0].a/w1120 ), .Z(\SUBBYTES[0].a/n650 ) );
  XOR \SUBBYTES[0].a/U5237  ( .A(\SUBBYTES[0].a/n1481 ), .B(
        \SUBBYTES[0].a/n651 ), .Z(\SUBBYTES[0].a/n1707 ) );
  XOR \SUBBYTES[0].a/U5236  ( .A(\SUBBYTES[0].a/w1120 ), .B(
        \SUBBYTES[0].a/w1121 ), .Z(\SUBBYTES[0].a/n651 ) );
  XOR \SUBBYTES[0].a/U5235  ( .A(\SUBBYTES[0].a/w1082 ), .B(
        \SUBBYTES[0].a/n652 ), .Z(\SUBBYTES[0].a/n1483 ) );
  XOR \SUBBYTES[0].a/U5234  ( .A(\SUBBYTES[0].a/w1073 ), .B(
        \SUBBYTES[0].a/w1074 ), .Z(\SUBBYTES[0].a/n652 ) );
  XOR \SUBBYTES[0].a/U5232  ( .A(\SUBBYTES[0].a/w1084 ), .B(
        \SUBBYTES[0].a/n1707 ), .Z(\SUBBYTES[0].a/n653 ) );
  XOR \SUBBYTES[0].a/U5231  ( .A(\SUBBYTES[0].a/n655 ), .B(
        \SUBBYTES[0].a/n654 ), .Z(\SUBBYTES[0].a/n1484 ) );
  XOR \SUBBYTES[0].a/U5230  ( .A(\SUBBYTES[0].a/n657 ), .B(
        \SUBBYTES[0].a/n656 ), .Z(\SUBBYTES[0].a/n654 ) );
  XOR \SUBBYTES[0].a/U5229  ( .A(\SUBBYTES[0].a/w1120 ), .B(
        \SUBBYTES[0].a/w1121 ), .Z(\SUBBYTES[0].a/n655 ) );
  XOR \SUBBYTES[0].a/U5228  ( .A(\SUBBYTES[0].a/w1084 ), .B(
        \SUBBYTES[0].a/w1108 ), .Z(\SUBBYTES[0].a/n656 ) );
  XOR \SUBBYTES[0].a/U5227  ( .A(\SUBBYTES[0].a/w1073 ), .B(
        \SUBBYTES[0].a/w1082 ), .Z(\SUBBYTES[0].a/n657 ) );
  XOR \SUBBYTES[0].a/U5226  ( .A(\SUBBYTES[0].a/w1105 ), .B(
        \SUBBYTES[0].a/n658 ), .Z(\SUBBYTES[0].a/n1482 ) );
  XOR \SUBBYTES[0].a/U5225  ( .A(\SUBBYTES[0].a/w1088 ), .B(
        \SUBBYTES[0].a/w1091 ), .Z(\SUBBYTES[0].a/n658 ) );
  XOR \SUBBYTES[0].a/U5223  ( .A(\SUBBYTES[0].a/w1076 ), .B(
        \SUBBYTES[0].a/n1484 ), .Z(\SUBBYTES[0].a/n659 ) );
  XOR \SUBBYTES[0].a/U5221  ( .A(\SUBBYTES[0].a/w1108 ), .B(
        \SUBBYTES[0].a/w1121 ), .Z(\SUBBYTES[0].a/n660 ) );
  XOR \SUBBYTES[0].a/U5219  ( .A(\SUBBYTES[0].a/n664 ), .B(
        \SUBBYTES[0].a/n663 ), .Z(\SUBBYTES[0].a/n661 ) );
  XOR \SUBBYTES[0].a/U5218  ( .A(\SUBBYTES[0].a/n666 ), .B(
        \SUBBYTES[0].a/n665 ), .Z(\SUBBYTES[0].a/n662 ) );
  XOR \SUBBYTES[0].a/U5217  ( .A(\SUBBYTES[0].a/w1120 ), .B(
        \SUBBYTES[0].a/w1123 ), .Z(\SUBBYTES[0].a/n663 ) );
  XOR \SUBBYTES[0].a/U5216  ( .A(\SUBBYTES[0].a/w1113 ), .B(
        \SUBBYTES[0].a/w1116 ), .Z(\SUBBYTES[0].a/n664 ) );
  XOR \SUBBYTES[0].a/U5215  ( .A(\SUBBYTES[0].a/w1088 ), .B(
        \SUBBYTES[0].a/w1089 ), .Z(\SUBBYTES[0].a/n665 ) );
  XOR \SUBBYTES[0].a/U5214  ( .A(\SUBBYTES[0].a/w1073 ), .B(
        \SUBBYTES[0].a/w1076 ), .Z(\SUBBYTES[0].a/n666 ) );
  XOR \SUBBYTES[0].a/U5212  ( .A(\SUBBYTES[0].a/n1481 ), .B(
        \SUBBYTES[0].a/n669 ), .Z(\SUBBYTES[0].a/n667 ) );
  XOR \SUBBYTES[0].a/U5211  ( .A(\SUBBYTES[0].a/n1483 ), .B(
        \SUBBYTES[0].a/n1482 ), .Z(\SUBBYTES[0].a/n668 ) );
  XOR \SUBBYTES[0].a/U5210  ( .A(\SUBBYTES[0].a/w1081 ), .B(
        \SUBBYTES[0].a/w1108 ), .Z(\SUBBYTES[0].a/n669 ) );
  XOR \SUBBYTES[0].a/U5208  ( .A(\SUBBYTES[0].a/n1484 ), .B(
        \SUBBYTES[0].a/n672 ), .Z(\SUBBYTES[0].a/n670 ) );
  XOR \SUBBYTES[0].a/U5207  ( .A(\SUBBYTES[0].a/w1114 ), .B(
        \SUBBYTES[0].a/w1116 ), .Z(\SUBBYTES[0].a/n671 ) );
  XOR \SUBBYTES[0].a/U5206  ( .A(\SUBBYTES[0].a/w1074 ), .B(
        \SUBBYTES[0].a/w1106 ), .Z(\SUBBYTES[0].a/n672 ) );
  XOR \SUBBYTES[0].a/U5205  ( .A(\SUBBYTES[0].a/w906 ), .B(
        \SUBBYTES[0].a/w907 ), .Z(\SUBBYTES[0].a/n1486 ) );
  XOR \SUBBYTES[0].a/U5204  ( .A(\SUBBYTES[0].a/n1486 ), .B(
        \SUBBYTES[0].a/n673 ), .Z(\SUBBYTES[0].a/n1485 ) );
  XOR \SUBBYTES[0].a/U5203  ( .A(\SUBBYTES[0].a/w899 ), .B(
        \SUBBYTES[0].a/w916 ), .Z(\SUBBYTES[0].a/n673 ) );
  XOR \SUBBYTES[0].a/U5201  ( .A(\SUBBYTES[0].a/w898 ), .B(
        \SUBBYTES[0].a/w913 ), .Z(\SUBBYTES[0].a/n674 ) );
  XOR \SUBBYTES[0].a/U5200  ( .A(\SUBBYTES[0].a/n1486 ), .B(
        \SUBBYTES[0].a/n675 ), .Z(\SUBBYTES[0].a/n1715 ) );
  XOR \SUBBYTES[0].a/U5199  ( .A(\SUBBYTES[0].a/w913 ), .B(
        \SUBBYTES[0].a/w914 ), .Z(\SUBBYTES[0].a/n675 ) );
  XOR \SUBBYTES[0].a/U5198  ( .A(\SUBBYTES[0].a/w875 ), .B(
        \SUBBYTES[0].a/n676 ), .Z(\SUBBYTES[0].a/n1488 ) );
  XOR \SUBBYTES[0].a/U5197  ( .A(\SUBBYTES[0].a/w866 ), .B(
        \SUBBYTES[0].a/w867 ), .Z(\SUBBYTES[0].a/n676 ) );
  XOR \SUBBYTES[0].a/U5195  ( .A(\SUBBYTES[0].a/w877 ), .B(
        \SUBBYTES[0].a/n1715 ), .Z(\SUBBYTES[0].a/n677 ) );
  XOR \SUBBYTES[0].a/U5194  ( .A(\SUBBYTES[0].a/n679 ), .B(
        \SUBBYTES[0].a/n678 ), .Z(\SUBBYTES[0].a/n1489 ) );
  XOR \SUBBYTES[0].a/U5193  ( .A(\SUBBYTES[0].a/n681 ), .B(
        \SUBBYTES[0].a/n680 ), .Z(\SUBBYTES[0].a/n678 ) );
  XOR \SUBBYTES[0].a/U5192  ( .A(\SUBBYTES[0].a/w913 ), .B(
        \SUBBYTES[0].a/w914 ), .Z(\SUBBYTES[0].a/n679 ) );
  XOR \SUBBYTES[0].a/U5191  ( .A(\SUBBYTES[0].a/w877 ), .B(
        \SUBBYTES[0].a/w901 ), .Z(\SUBBYTES[0].a/n680 ) );
  XOR \SUBBYTES[0].a/U5190  ( .A(\SUBBYTES[0].a/w866 ), .B(
        \SUBBYTES[0].a/w875 ), .Z(\SUBBYTES[0].a/n681 ) );
  XOR \SUBBYTES[0].a/U5189  ( .A(\SUBBYTES[0].a/w898 ), .B(
        \SUBBYTES[0].a/n682 ), .Z(\SUBBYTES[0].a/n1487 ) );
  XOR \SUBBYTES[0].a/U5188  ( .A(\SUBBYTES[0].a/w881 ), .B(
        \SUBBYTES[0].a/w884 ), .Z(\SUBBYTES[0].a/n682 ) );
  XOR \SUBBYTES[0].a/U5186  ( .A(\SUBBYTES[0].a/w869 ), .B(
        \SUBBYTES[0].a/n1489 ), .Z(\SUBBYTES[0].a/n683 ) );
  XOR \SUBBYTES[0].a/U5184  ( .A(\SUBBYTES[0].a/w901 ), .B(
        \SUBBYTES[0].a/w914 ), .Z(\SUBBYTES[0].a/n684 ) );
  XOR \SUBBYTES[0].a/U5182  ( .A(\SUBBYTES[0].a/n688 ), .B(
        \SUBBYTES[0].a/n687 ), .Z(\SUBBYTES[0].a/n685 ) );
  XOR \SUBBYTES[0].a/U5181  ( .A(\SUBBYTES[0].a/n690 ), .B(
        \SUBBYTES[0].a/n689 ), .Z(\SUBBYTES[0].a/n686 ) );
  XOR \SUBBYTES[0].a/U5180  ( .A(\SUBBYTES[0].a/w913 ), .B(
        \SUBBYTES[0].a/w916 ), .Z(\SUBBYTES[0].a/n687 ) );
  XOR \SUBBYTES[0].a/U5179  ( .A(\SUBBYTES[0].a/w906 ), .B(
        \SUBBYTES[0].a/w909 ), .Z(\SUBBYTES[0].a/n688 ) );
  XOR \SUBBYTES[0].a/U5178  ( .A(\SUBBYTES[0].a/w881 ), .B(
        \SUBBYTES[0].a/w882 ), .Z(\SUBBYTES[0].a/n689 ) );
  XOR \SUBBYTES[0].a/U5177  ( .A(\SUBBYTES[0].a/w866 ), .B(
        \SUBBYTES[0].a/w869 ), .Z(\SUBBYTES[0].a/n690 ) );
  XOR \SUBBYTES[0].a/U5175  ( .A(\SUBBYTES[0].a/n1486 ), .B(
        \SUBBYTES[0].a/n693 ), .Z(\SUBBYTES[0].a/n691 ) );
  XOR \SUBBYTES[0].a/U5174  ( .A(\SUBBYTES[0].a/n1488 ), .B(
        \SUBBYTES[0].a/n1487 ), .Z(\SUBBYTES[0].a/n692 ) );
  XOR \SUBBYTES[0].a/U5173  ( .A(\SUBBYTES[0].a/w874 ), .B(
        \SUBBYTES[0].a/w901 ), .Z(\SUBBYTES[0].a/n693 ) );
  XOR \SUBBYTES[0].a/U5171  ( .A(\SUBBYTES[0].a/n1489 ), .B(
        \SUBBYTES[0].a/n696 ), .Z(\SUBBYTES[0].a/n694 ) );
  XOR \SUBBYTES[0].a/U5170  ( .A(\SUBBYTES[0].a/w907 ), .B(
        \SUBBYTES[0].a/w909 ), .Z(\SUBBYTES[0].a/n695 ) );
  XOR \SUBBYTES[0].a/U5169  ( .A(\SUBBYTES[0].a/w867 ), .B(
        \SUBBYTES[0].a/w899 ), .Z(\SUBBYTES[0].a/n696 ) );
  XOR \SUBBYTES[0].a/U5168  ( .A(\SUBBYTES[0].a/w699 ), .B(
        \SUBBYTES[0].a/w700 ), .Z(\SUBBYTES[0].a/n1491 ) );
  XOR \SUBBYTES[0].a/U5167  ( .A(\SUBBYTES[0].a/n1491 ), .B(
        \SUBBYTES[0].a/n697 ), .Z(\SUBBYTES[0].a/n1490 ) );
  XOR \SUBBYTES[0].a/U5166  ( .A(\SUBBYTES[0].a/w692 ), .B(
        \SUBBYTES[0].a/w709 ), .Z(\SUBBYTES[0].a/n697 ) );
  XOR \SUBBYTES[0].a/U5164  ( .A(\SUBBYTES[0].a/w691 ), .B(
        \SUBBYTES[0].a/w706 ), .Z(\SUBBYTES[0].a/n698 ) );
  XOR \SUBBYTES[0].a/U5163  ( .A(\SUBBYTES[0].a/n1491 ), .B(
        \SUBBYTES[0].a/n699 ), .Z(\SUBBYTES[0].a/n1723 ) );
  XOR \SUBBYTES[0].a/U5162  ( .A(\SUBBYTES[0].a/w706 ), .B(
        \SUBBYTES[0].a/w707 ), .Z(\SUBBYTES[0].a/n699 ) );
  XOR \SUBBYTES[0].a/U5161  ( .A(\SUBBYTES[0].a/w668 ), .B(
        \SUBBYTES[0].a/n700 ), .Z(\SUBBYTES[0].a/n1493 ) );
  XOR \SUBBYTES[0].a/U5160  ( .A(\SUBBYTES[0].a/w659 ), .B(
        \SUBBYTES[0].a/w660 ), .Z(\SUBBYTES[0].a/n700 ) );
  XOR \SUBBYTES[0].a/U5158  ( .A(\SUBBYTES[0].a/w670 ), .B(
        \SUBBYTES[0].a/n1723 ), .Z(\SUBBYTES[0].a/n701 ) );
  XOR \SUBBYTES[0].a/U5157  ( .A(\SUBBYTES[0].a/n703 ), .B(
        \SUBBYTES[0].a/n702 ), .Z(\SUBBYTES[0].a/n1494 ) );
  XOR \SUBBYTES[0].a/U5156  ( .A(\SUBBYTES[0].a/n705 ), .B(
        \SUBBYTES[0].a/n704 ), .Z(\SUBBYTES[0].a/n702 ) );
  XOR \SUBBYTES[0].a/U5155  ( .A(\SUBBYTES[0].a/w706 ), .B(
        \SUBBYTES[0].a/w707 ), .Z(\SUBBYTES[0].a/n703 ) );
  XOR \SUBBYTES[0].a/U5154  ( .A(\SUBBYTES[0].a/w670 ), .B(
        \SUBBYTES[0].a/w694 ), .Z(\SUBBYTES[0].a/n704 ) );
  XOR \SUBBYTES[0].a/U5153  ( .A(\SUBBYTES[0].a/w659 ), .B(
        \SUBBYTES[0].a/w668 ), .Z(\SUBBYTES[0].a/n705 ) );
  XOR \SUBBYTES[0].a/U5152  ( .A(\SUBBYTES[0].a/w691 ), .B(
        \SUBBYTES[0].a/n706 ), .Z(\SUBBYTES[0].a/n1492 ) );
  XOR \SUBBYTES[0].a/U5151  ( .A(\SUBBYTES[0].a/w674 ), .B(
        \SUBBYTES[0].a/w677 ), .Z(\SUBBYTES[0].a/n706 ) );
  XOR \SUBBYTES[0].a/U5149  ( .A(\SUBBYTES[0].a/w662 ), .B(
        \SUBBYTES[0].a/n1494 ), .Z(\SUBBYTES[0].a/n707 ) );
  XOR \SUBBYTES[0].a/U5147  ( .A(\SUBBYTES[0].a/w694 ), .B(
        \SUBBYTES[0].a/w707 ), .Z(\SUBBYTES[0].a/n708 ) );
  XOR \SUBBYTES[0].a/U5145  ( .A(\SUBBYTES[0].a/n712 ), .B(
        \SUBBYTES[0].a/n711 ), .Z(\SUBBYTES[0].a/n709 ) );
  XOR \SUBBYTES[0].a/U5144  ( .A(\SUBBYTES[0].a/n714 ), .B(
        \SUBBYTES[0].a/n713 ), .Z(\SUBBYTES[0].a/n710 ) );
  XOR \SUBBYTES[0].a/U5143  ( .A(\SUBBYTES[0].a/w706 ), .B(
        \SUBBYTES[0].a/w709 ), .Z(\SUBBYTES[0].a/n711 ) );
  XOR \SUBBYTES[0].a/U5142  ( .A(\SUBBYTES[0].a/w699 ), .B(
        \SUBBYTES[0].a/w702 ), .Z(\SUBBYTES[0].a/n712 ) );
  XOR \SUBBYTES[0].a/U5141  ( .A(\SUBBYTES[0].a/w674 ), .B(
        \SUBBYTES[0].a/w675 ), .Z(\SUBBYTES[0].a/n713 ) );
  XOR \SUBBYTES[0].a/U5140  ( .A(\SUBBYTES[0].a/w659 ), .B(
        \SUBBYTES[0].a/w662 ), .Z(\SUBBYTES[0].a/n714 ) );
  XOR \SUBBYTES[0].a/U5138  ( .A(\SUBBYTES[0].a/n1491 ), .B(
        \SUBBYTES[0].a/n717 ), .Z(\SUBBYTES[0].a/n715 ) );
  XOR \SUBBYTES[0].a/U5137  ( .A(\SUBBYTES[0].a/n1493 ), .B(
        \SUBBYTES[0].a/n1492 ), .Z(\SUBBYTES[0].a/n716 ) );
  XOR \SUBBYTES[0].a/U5136  ( .A(\SUBBYTES[0].a/w667 ), .B(
        \SUBBYTES[0].a/w694 ), .Z(\SUBBYTES[0].a/n717 ) );
  XOR \SUBBYTES[0].a/U5134  ( .A(\SUBBYTES[0].a/n1494 ), .B(
        \SUBBYTES[0].a/n720 ), .Z(\SUBBYTES[0].a/n718 ) );
  XOR \SUBBYTES[0].a/U5133  ( .A(\SUBBYTES[0].a/w700 ), .B(
        \SUBBYTES[0].a/w702 ), .Z(\SUBBYTES[0].a/n719 ) );
  XOR \SUBBYTES[0].a/U5132  ( .A(\SUBBYTES[0].a/w660 ), .B(
        \SUBBYTES[0].a/w692 ), .Z(\SUBBYTES[0].a/n720 ) );
  XOR \SUBBYTES[0].a/U5131  ( .A(\SUBBYTES[0].a/w492 ), .B(
        \SUBBYTES[0].a/w493 ), .Z(\SUBBYTES[0].a/n1496 ) );
  XOR \SUBBYTES[0].a/U5130  ( .A(\SUBBYTES[0].a/n1496 ), .B(
        \SUBBYTES[0].a/n721 ), .Z(\SUBBYTES[0].a/n1495 ) );
  XOR \SUBBYTES[0].a/U5129  ( .A(\SUBBYTES[0].a/w485 ), .B(
        \SUBBYTES[0].a/w502 ), .Z(\SUBBYTES[0].a/n721 ) );
  XOR \SUBBYTES[0].a/U5127  ( .A(\SUBBYTES[0].a/w484 ), .B(
        \SUBBYTES[0].a/w499 ), .Z(\SUBBYTES[0].a/n722 ) );
  XOR \SUBBYTES[0].a/U5126  ( .A(\SUBBYTES[0].a/n1496 ), .B(
        \SUBBYTES[0].a/n723 ), .Z(\SUBBYTES[0].a/n1731 ) );
  XOR \SUBBYTES[0].a/U5125  ( .A(\SUBBYTES[0].a/w499 ), .B(
        \SUBBYTES[0].a/w500 ), .Z(\SUBBYTES[0].a/n723 ) );
  XOR \SUBBYTES[0].a/U5124  ( .A(\SUBBYTES[0].a/w461 ), .B(
        \SUBBYTES[0].a/n724 ), .Z(\SUBBYTES[0].a/n1498 ) );
  XOR \SUBBYTES[0].a/U5123  ( .A(\SUBBYTES[0].a/w452 ), .B(
        \SUBBYTES[0].a/w453 ), .Z(\SUBBYTES[0].a/n724 ) );
  XOR \SUBBYTES[0].a/U5121  ( .A(\SUBBYTES[0].a/w463 ), .B(
        \SUBBYTES[0].a/n1731 ), .Z(\SUBBYTES[0].a/n725 ) );
  XOR \SUBBYTES[0].a/U5120  ( .A(\SUBBYTES[0].a/n727 ), .B(
        \SUBBYTES[0].a/n726 ), .Z(\SUBBYTES[0].a/n1499 ) );
  XOR \SUBBYTES[0].a/U5119  ( .A(\SUBBYTES[0].a/n729 ), .B(
        \SUBBYTES[0].a/n728 ), .Z(\SUBBYTES[0].a/n726 ) );
  XOR \SUBBYTES[0].a/U5118  ( .A(\SUBBYTES[0].a/w499 ), .B(
        \SUBBYTES[0].a/w500 ), .Z(\SUBBYTES[0].a/n727 ) );
  XOR \SUBBYTES[0].a/U5117  ( .A(\SUBBYTES[0].a/w463 ), .B(
        \SUBBYTES[0].a/w487 ), .Z(\SUBBYTES[0].a/n728 ) );
  XOR \SUBBYTES[0].a/U5116  ( .A(\SUBBYTES[0].a/w452 ), .B(
        \SUBBYTES[0].a/w461 ), .Z(\SUBBYTES[0].a/n729 ) );
  XOR \SUBBYTES[0].a/U5115  ( .A(\SUBBYTES[0].a/w484 ), .B(
        \SUBBYTES[0].a/n730 ), .Z(\SUBBYTES[0].a/n1497 ) );
  XOR \SUBBYTES[0].a/U5114  ( .A(\SUBBYTES[0].a/w467 ), .B(
        \SUBBYTES[0].a/w470 ), .Z(\SUBBYTES[0].a/n730 ) );
  XOR \SUBBYTES[0].a/U5112  ( .A(\SUBBYTES[0].a/w455 ), .B(
        \SUBBYTES[0].a/n1499 ), .Z(\SUBBYTES[0].a/n731 ) );
  XOR \SUBBYTES[0].a/U5110  ( .A(\SUBBYTES[0].a/w487 ), .B(
        \SUBBYTES[0].a/w500 ), .Z(\SUBBYTES[0].a/n732 ) );
  XOR \SUBBYTES[0].a/U5108  ( .A(\SUBBYTES[0].a/n736 ), .B(
        \SUBBYTES[0].a/n735 ), .Z(\SUBBYTES[0].a/n733 ) );
  XOR \SUBBYTES[0].a/U5107  ( .A(\SUBBYTES[0].a/n738 ), .B(
        \SUBBYTES[0].a/n737 ), .Z(\SUBBYTES[0].a/n734 ) );
  XOR \SUBBYTES[0].a/U5106  ( .A(\SUBBYTES[0].a/w499 ), .B(
        \SUBBYTES[0].a/w502 ), .Z(\SUBBYTES[0].a/n735 ) );
  XOR \SUBBYTES[0].a/U5105  ( .A(\SUBBYTES[0].a/w492 ), .B(
        \SUBBYTES[0].a/w495 ), .Z(\SUBBYTES[0].a/n736 ) );
  XOR \SUBBYTES[0].a/U5104  ( .A(\SUBBYTES[0].a/w467 ), .B(
        \SUBBYTES[0].a/w468 ), .Z(\SUBBYTES[0].a/n737 ) );
  XOR \SUBBYTES[0].a/U5103  ( .A(\SUBBYTES[0].a/w452 ), .B(
        \SUBBYTES[0].a/w455 ), .Z(\SUBBYTES[0].a/n738 ) );
  XOR \SUBBYTES[0].a/U5101  ( .A(\SUBBYTES[0].a/n1496 ), .B(
        \SUBBYTES[0].a/n741 ), .Z(\SUBBYTES[0].a/n739 ) );
  XOR \SUBBYTES[0].a/U5100  ( .A(\SUBBYTES[0].a/n1498 ), .B(
        \SUBBYTES[0].a/n1497 ), .Z(\SUBBYTES[0].a/n740 ) );
  XOR \SUBBYTES[0].a/U5099  ( .A(\SUBBYTES[0].a/w460 ), .B(
        \SUBBYTES[0].a/w487 ), .Z(\SUBBYTES[0].a/n741 ) );
  XOR \SUBBYTES[0].a/U5097  ( .A(\SUBBYTES[0].a/n1499 ), .B(
        \SUBBYTES[0].a/n744 ), .Z(\SUBBYTES[0].a/n742 ) );
  XOR \SUBBYTES[0].a/U5096  ( .A(\SUBBYTES[0].a/w493 ), .B(
        \SUBBYTES[0].a/w495 ), .Z(\SUBBYTES[0].a/n743 ) );
  XOR \SUBBYTES[0].a/U5095  ( .A(\SUBBYTES[0].a/w453 ), .B(
        \SUBBYTES[0].a/w485 ), .Z(\SUBBYTES[0].a/n744 ) );
  XOR \SUBBYTES[0].a/U5094  ( .A(\SUBBYTES[0].a/w285 ), .B(
        \SUBBYTES[0].a/w286 ), .Z(\SUBBYTES[0].a/n1501 ) );
  XOR \SUBBYTES[0].a/U5093  ( .A(\SUBBYTES[0].a/n1501 ), .B(
        \SUBBYTES[0].a/n745 ), .Z(\SUBBYTES[0].a/n1500 ) );
  XOR \SUBBYTES[0].a/U5092  ( .A(\SUBBYTES[0].a/w278 ), .B(
        \SUBBYTES[0].a/w295 ), .Z(\SUBBYTES[0].a/n745 ) );
  XOR \SUBBYTES[0].a/U5090  ( .A(\SUBBYTES[0].a/w277 ), .B(
        \SUBBYTES[0].a/w292 ), .Z(\SUBBYTES[0].a/n746 ) );
  XOR \SUBBYTES[0].a/U5089  ( .A(\SUBBYTES[0].a/n1501 ), .B(
        \SUBBYTES[0].a/n747 ), .Z(\SUBBYTES[0].a/n1739 ) );
  XOR \SUBBYTES[0].a/U5088  ( .A(\SUBBYTES[0].a/w292 ), .B(
        \SUBBYTES[0].a/w293 ), .Z(\SUBBYTES[0].a/n747 ) );
  XOR \SUBBYTES[0].a/U5087  ( .A(\SUBBYTES[0].a/w254 ), .B(
        \SUBBYTES[0].a/n748 ), .Z(\SUBBYTES[0].a/n1503 ) );
  XOR \SUBBYTES[0].a/U5086  ( .A(\SUBBYTES[0].a/w245 ), .B(
        \SUBBYTES[0].a/w246 ), .Z(\SUBBYTES[0].a/n748 ) );
  XOR \SUBBYTES[0].a/U5084  ( .A(\SUBBYTES[0].a/w256 ), .B(
        \SUBBYTES[0].a/n1739 ), .Z(\SUBBYTES[0].a/n749 ) );
  XOR \SUBBYTES[0].a/U5083  ( .A(\SUBBYTES[0].a/n751 ), .B(
        \SUBBYTES[0].a/n750 ), .Z(\SUBBYTES[0].a/n1504 ) );
  XOR \SUBBYTES[0].a/U5082  ( .A(\SUBBYTES[0].a/n753 ), .B(
        \SUBBYTES[0].a/n752 ), .Z(\SUBBYTES[0].a/n750 ) );
  XOR \SUBBYTES[0].a/U5081  ( .A(\SUBBYTES[0].a/w292 ), .B(
        \SUBBYTES[0].a/w293 ), .Z(\SUBBYTES[0].a/n751 ) );
  XOR \SUBBYTES[0].a/U5080  ( .A(\SUBBYTES[0].a/w256 ), .B(
        \SUBBYTES[0].a/w280 ), .Z(\SUBBYTES[0].a/n752 ) );
  XOR \SUBBYTES[0].a/U5079  ( .A(\SUBBYTES[0].a/w245 ), .B(
        \SUBBYTES[0].a/w254 ), .Z(\SUBBYTES[0].a/n753 ) );
  XOR \SUBBYTES[0].a/U5078  ( .A(\SUBBYTES[0].a/w277 ), .B(
        \SUBBYTES[0].a/n754 ), .Z(\SUBBYTES[0].a/n1502 ) );
  XOR \SUBBYTES[0].a/U5077  ( .A(\SUBBYTES[0].a/w260 ), .B(
        \SUBBYTES[0].a/w263 ), .Z(\SUBBYTES[0].a/n754 ) );
  XOR \SUBBYTES[0].a/U5075  ( .A(\SUBBYTES[0].a/w248 ), .B(
        \SUBBYTES[0].a/n1504 ), .Z(\SUBBYTES[0].a/n755 ) );
  XOR \SUBBYTES[0].a/U5073  ( .A(\SUBBYTES[0].a/w280 ), .B(
        \SUBBYTES[0].a/w293 ), .Z(\SUBBYTES[0].a/n756 ) );
  XOR \SUBBYTES[0].a/U5071  ( .A(\SUBBYTES[0].a/n760 ), .B(
        \SUBBYTES[0].a/n759 ), .Z(\SUBBYTES[0].a/n757 ) );
  XOR \SUBBYTES[0].a/U5070  ( .A(\SUBBYTES[0].a/n762 ), .B(
        \SUBBYTES[0].a/n761 ), .Z(\SUBBYTES[0].a/n758 ) );
  XOR \SUBBYTES[0].a/U5069  ( .A(\SUBBYTES[0].a/w292 ), .B(
        \SUBBYTES[0].a/w295 ), .Z(\SUBBYTES[0].a/n759 ) );
  XOR \SUBBYTES[0].a/U5068  ( .A(\SUBBYTES[0].a/w285 ), .B(
        \SUBBYTES[0].a/w288 ), .Z(\SUBBYTES[0].a/n760 ) );
  XOR \SUBBYTES[0].a/U5067  ( .A(\SUBBYTES[0].a/w260 ), .B(
        \SUBBYTES[0].a/w261 ), .Z(\SUBBYTES[0].a/n761 ) );
  XOR \SUBBYTES[0].a/U5066  ( .A(\SUBBYTES[0].a/w245 ), .B(
        \SUBBYTES[0].a/w248 ), .Z(\SUBBYTES[0].a/n762 ) );
  XOR \SUBBYTES[0].a/U5064  ( .A(\SUBBYTES[0].a/n1501 ), .B(
        \SUBBYTES[0].a/n765 ), .Z(\SUBBYTES[0].a/n763 ) );
  XOR \SUBBYTES[0].a/U5063  ( .A(\SUBBYTES[0].a/n1503 ), .B(
        \SUBBYTES[0].a/n1502 ), .Z(\SUBBYTES[0].a/n764 ) );
  XOR \SUBBYTES[0].a/U5062  ( .A(\SUBBYTES[0].a/w253 ), .B(
        \SUBBYTES[0].a/w280 ), .Z(\SUBBYTES[0].a/n765 ) );
  XOR \SUBBYTES[0].a/U5060  ( .A(\SUBBYTES[0].a/n1504 ), .B(
        \SUBBYTES[0].a/n768 ), .Z(\SUBBYTES[0].a/n766 ) );
  XOR \SUBBYTES[0].a/U5059  ( .A(\SUBBYTES[0].a/w286 ), .B(
        \SUBBYTES[0].a/w288 ), .Z(\SUBBYTES[0].a/n767 ) );
  XOR \SUBBYTES[0].a/U5058  ( .A(\SUBBYTES[0].a/w246 ), .B(
        \SUBBYTES[0].a/w278 ), .Z(\SUBBYTES[0].a/n768 ) );
  XOR \SUBBYTES[0].a/U5057  ( .A(\w1[0][1] ), .B(\SUBBYTES[0].a/n769 ), .Z(
        \SUBBYTES[0].a/n1505 ) );
  XOR \SUBBYTES[0].a/U5056  ( .A(\w1[0][3] ), .B(\w1[0][2] ), .Z(
        \SUBBYTES[0].a/n769 ) );
  XOR \SUBBYTES[0].a/U5055  ( .A(\w1[0][6] ), .B(\SUBBYTES[0].a/n1505 ), .Z(
        \SUBBYTES[0].a/w3378 ) );
  XOR \SUBBYTES[0].a/U5054  ( .A(\w1[0][0] ), .B(\SUBBYTES[0].a/w3378 ), .Z(
        \SUBBYTES[0].a/w3265 ) );
  XOR \SUBBYTES[0].a/U5053  ( .A(\w1[0][0] ), .B(\SUBBYTES[0].a/n770 ), .Z(
        \SUBBYTES[0].a/w3266 ) );
  XOR \SUBBYTES[0].a/U5052  ( .A(\w1[0][6] ), .B(\w1[0][5] ), .Z(
        \SUBBYTES[0].a/n770 ) );
  XOR \SUBBYTES[0].a/U5051  ( .A(\w1[0][5] ), .B(\SUBBYTES[0].a/n1505 ), .Z(
        \SUBBYTES[0].a/w3396 ) );
  XOR \SUBBYTES[0].a/U5050  ( .A(\SUBBYTES[0].a/n772 ), .B(
        \SUBBYTES[0].a/n771 ), .Z(\SUBBYTES[0].a/w3389 ) );
  XOR \SUBBYTES[0].a/U5049  ( .A(\w1[0][3] ), .B(\w1[0][1] ), .Z(
        \SUBBYTES[0].a/n771 ) );
  XOR \SUBBYTES[0].a/U5048  ( .A(\w1[0][7] ), .B(\w1[0][4] ), .Z(
        \SUBBYTES[0].a/n772 ) );
  XOR \SUBBYTES[0].a/U5047  ( .A(\w1[0][0] ), .B(\SUBBYTES[0].a/w3389 ), .Z(
        \SUBBYTES[0].a/w3268 ) );
  XOR \SUBBYTES[0].a/U5046  ( .A(\SUBBYTES[0].a/n774 ), .B(
        \SUBBYTES[0].a/n773 ), .Z(\SUBBYTES[0].a/w3376 ) );
  XOR \SUBBYTES[0].a/U5045  ( .A(\SUBBYTES[0].a/w3337 ), .B(n1168), .Z(
        \SUBBYTES[0].a/n773 ) );
  XOR \SUBBYTES[0].a/U5044  ( .A(\SUBBYTES[0].a/w3330 ), .B(
        \SUBBYTES[0].a/w3333 ), .Z(\SUBBYTES[0].a/n774 ) );
  XOR \SUBBYTES[0].a/U5043  ( .A(\SUBBYTES[0].a/n776 ), .B(
        \SUBBYTES[0].a/n775 ), .Z(\SUBBYTES[0].a/w3377 ) );
  XOR \SUBBYTES[0].a/U5042  ( .A(\SUBBYTES[0].a/w3337 ), .B(
        \SUBBYTES[0].a/n160 ), .Z(\SUBBYTES[0].a/n775 ) );
  XOR \SUBBYTES[0].a/U5041  ( .A(\SUBBYTES[0].a/w3330 ), .B(
        \SUBBYTES[0].a/n159 ), .Z(\SUBBYTES[0].a/n776 ) );
  XOR \SUBBYTES[0].a/U5040  ( .A(\SUBBYTES[0].a/w3389 ), .B(
        \SUBBYTES[0].a/n777 ), .Z(\SUBBYTES[0].a/w3379 ) );
  XOR \SUBBYTES[0].a/U5039  ( .A(\w1[0][6] ), .B(\w1[0][5] ), .Z(
        \SUBBYTES[0].a/n777 ) );
  XOR \SUBBYTES[0].a/U5038  ( .A(\SUBBYTES[0].a/n779 ), .B(
        \SUBBYTES[0].a/n778 ), .Z(\SUBBYTES[0].a/w3380 ) );
  XOR \SUBBYTES[0].a/U5037  ( .A(\SUBBYTES[0].a/n160 ), .B(n1168), .Z(
        \SUBBYTES[0].a/n778 ) );
  XOR \SUBBYTES[0].a/U5036  ( .A(\SUBBYTES[0].a/n159 ), .B(
        \SUBBYTES[0].a/w3333 ), .Z(\SUBBYTES[0].a/n779 ) );
  XOR \SUBBYTES[0].a/U5035  ( .A(\w1[0][7] ), .B(\w1[0][2] ), .Z(
        \SUBBYTES[0].a/n1511 ) );
  XOR \SUBBYTES[0].a/U5034  ( .A(\SUBBYTES[0].a/n1511 ), .B(
        \SUBBYTES[0].a/n780 ), .Z(\SUBBYTES[0].a/w3381 ) );
  XOR \SUBBYTES[0].a/U5033  ( .A(\w1[0][5] ), .B(\w1[0][4] ), .Z(
        \SUBBYTES[0].a/n780 ) );
  XOR \SUBBYTES[0].a/U5032  ( .A(\w1[0][7] ), .B(\SUBBYTES[0].a/w3266 ), .Z(
        \SUBBYTES[0].a/w3269 ) );
  XOR \SUBBYTES[0].a/U5031  ( .A(\w1[0][1] ), .B(\SUBBYTES[0].a/w3266 ), .Z(
        \SUBBYTES[0].a/w3270 ) );
  XOR \SUBBYTES[0].a/U5030  ( .A(\w1[0][4] ), .B(\SUBBYTES[0].a/w3266 ), .Z(
        \SUBBYTES[0].a/w3271 ) );
  XOR \SUBBYTES[0].a/U5029  ( .A(\SUBBYTES[0].a/w3270 ), .B(
        \SUBBYTES[0].a/n1511 ), .Z(\SUBBYTES[0].a/w3272 ) );
  XOR \SUBBYTES[0].a/U5028  ( .A(\SUBBYTES[0].a/n1511 ), .B(
        \SUBBYTES[0].a/n781 ), .Z(\SUBBYTES[0].a/w3357 ) );
  XOR \SUBBYTES[0].a/U5027  ( .A(\w1[0][4] ), .B(\w1[0][1] ), .Z(
        \SUBBYTES[0].a/n781 ) );
  XOR \SUBBYTES[0].a/U5026  ( .A(\SUBBYTES[0].a/n783 ), .B(
        \SUBBYTES[0].a/n782 ), .Z(\SUBBYTES[0].a/n1508 ) );
  XOR \SUBBYTES[0].a/U5025  ( .A(\w1[0][4] ), .B(\SUBBYTES[0].a/n784 ), .Z(
        \SUBBYTES[0].a/n782 ) );
  XOR \SUBBYTES[0].a/U5024  ( .A(\SUBBYTES[0].a/w3322 ), .B(\w1[0][6] ), .Z(
        \SUBBYTES[0].a/n783 ) );
  XOR \SUBBYTES[0].a/U5023  ( .A(\SUBBYTES[0].a/w3296 ), .B(
        \SUBBYTES[0].a/w3303 ), .Z(\SUBBYTES[0].a/n784 ) );
  XOR \SUBBYTES[0].a/U5022  ( .A(\SUBBYTES[0].a/n786 ), .B(
        \SUBBYTES[0].a/n785 ), .Z(\SUBBYTES[0].a/n1506 ) );
  XOR \SUBBYTES[0].a/U5021  ( .A(\w1[0][1] ), .B(\SUBBYTES[0].a/n787 ), .Z(
        \SUBBYTES[0].a/n785 ) );
  XOR \SUBBYTES[0].a/U5020  ( .A(\SUBBYTES[0].a/w3321 ), .B(\w1[0][5] ), .Z(
        \SUBBYTES[0].a/n786 ) );
  XOR \SUBBYTES[0].a/U5019  ( .A(\SUBBYTES[0].a/w3297 ), .B(
        \SUBBYTES[0].a/w3304 ), .Z(\SUBBYTES[0].a/n787 ) );
  XOR \SUBBYTES[0].a/U5018  ( .A(\SUBBYTES[0].a/n1508 ), .B(
        \SUBBYTES[0].a/n1506 ), .Z(\SUBBYTES[0].a/w3327 ) );
  XOR \SUBBYTES[0].a/U5017  ( .A(\w1[0][5] ), .B(\SUBBYTES[0].a/n788 ), .Z(
        \SUBBYTES[0].a/n1509 ) );
  XOR \SUBBYTES[0].a/U5016  ( .A(\SUBBYTES[0].a/w3289 ), .B(
        \SUBBYTES[0].a/w3299 ), .Z(\SUBBYTES[0].a/n788 ) );
  XOR \SUBBYTES[0].a/U5015  ( .A(\SUBBYTES[0].a/n790 ), .B(
        \SUBBYTES[0].a/n789 ), .Z(\SUBBYTES[0].a/w3314 ) );
  XOR \SUBBYTES[0].a/U5014  ( .A(\SUBBYTES[0].a/n1509 ), .B(
        \SUBBYTES[0].a/n791 ), .Z(\SUBBYTES[0].a/n789 ) );
  XOR \SUBBYTES[0].a/U5013  ( .A(\w1[0][4] ), .B(\SUBBYTES[0].a/w3378 ), .Z(
        \SUBBYTES[0].a/n790 ) );
  XOR \SUBBYTES[0].a/U5012  ( .A(\SUBBYTES[0].a/w3291 ), .B(
        \SUBBYTES[0].a/w3296 ), .Z(\SUBBYTES[0].a/n791 ) );
  XOR \SUBBYTES[0].a/U5011  ( .A(\SUBBYTES[0].a/n793 ), .B(
        \SUBBYTES[0].a/n792 ), .Z(\SUBBYTES[0].a/n1507 ) );
  XOR \SUBBYTES[0].a/U5010  ( .A(\SUBBYTES[0].a/w3324 ), .B(\w1[0][7] ), .Z(
        \SUBBYTES[0].a/n792 ) );
  XOR \SUBBYTES[0].a/U5009  ( .A(\SUBBYTES[0].a/w3299 ), .B(
        \SUBBYTES[0].a/w3306 ), .Z(\SUBBYTES[0].a/n793 ) );
  XOR \SUBBYTES[0].a/U5008  ( .A(\SUBBYTES[0].a/n1506 ), .B(
        \SUBBYTES[0].a/n1507 ), .Z(\SUBBYTES[0].a/w3326 ) );
  XOR \SUBBYTES[0].a/U5007  ( .A(\w1[0][3] ), .B(\SUBBYTES[0].a/n794 ), .Z(
        \SUBBYTES[0].a/n1510 ) );
  XOR \SUBBYTES[0].a/U5006  ( .A(\SUBBYTES[0].a/w3288 ), .B(
        \SUBBYTES[0].a/w3291 ), .Z(\SUBBYTES[0].a/n794 ) );
  XOR \SUBBYTES[0].a/U5005  ( .A(\SUBBYTES[0].a/n796 ), .B(
        \SUBBYTES[0].a/n795 ), .Z(\SUBBYTES[0].a/w3315 ) );
  XOR \SUBBYTES[0].a/U5004  ( .A(\SUBBYTES[0].a/n1510 ), .B(
        \SUBBYTES[0].a/n797 ), .Z(\SUBBYTES[0].a/n795 ) );
  XOR \SUBBYTES[0].a/U5003  ( .A(\w1[0][6] ), .B(\SUBBYTES[0].a/w3357 ), .Z(
        \SUBBYTES[0].a/n796 ) );
  XOR \SUBBYTES[0].a/U5002  ( .A(\SUBBYTES[0].a/w3296 ), .B(
        \SUBBYTES[0].a/w3297 ), .Z(\SUBBYTES[0].a/n797 ) );
  XOR \SUBBYTES[0].a/U5001  ( .A(\SUBBYTES[0].a/n1508 ), .B(
        \SUBBYTES[0].a/n1507 ), .Z(\SUBBYTES[0].a/w3335 ) );
  XOR \SUBBYTES[0].a/U5000  ( .A(\SUBBYTES[0].a/n799 ), .B(
        \SUBBYTES[0].a/n798 ), .Z(\SUBBYTES[0].a/w3336 ) );
  XOR \SUBBYTES[0].a/U4999  ( .A(\w1[0][7] ), .B(\SUBBYTES[0].a/n1509 ), .Z(
        \SUBBYTES[0].a/n798 ) );
  XOR \SUBBYTES[0].a/U4998  ( .A(\SUBBYTES[0].a/w3288 ), .B(
        \SUBBYTES[0].a/w3297 ), .Z(\SUBBYTES[0].a/n799 ) );
  XOR \SUBBYTES[0].a/U4997  ( .A(\SUBBYTES[0].a/n801 ), .B(
        \SUBBYTES[0].a/n800 ), .Z(\SUBBYTES[0].a/w3312 ) );
  XOR \SUBBYTES[0].a/U4996  ( .A(\SUBBYTES[0].a/n803 ), .B(
        \SUBBYTES[0].a/n802 ), .Z(\SUBBYTES[0].a/n800 ) );
  XOR \SUBBYTES[0].a/U4995  ( .A(\w1[0][7] ), .B(\SUBBYTES[0].a/w3396 ), .Z(
        \SUBBYTES[0].a/n801 ) );
  XOR \SUBBYTES[0].a/U4994  ( .A(\SUBBYTES[0].a/w3303 ), .B(
        \SUBBYTES[0].a/w3306 ), .Z(\SUBBYTES[0].a/n802 ) );
  XOR \SUBBYTES[0].a/U4993  ( .A(\SUBBYTES[0].a/w3289 ), .B(
        \SUBBYTES[0].a/w3291 ), .Z(\SUBBYTES[0].a/n803 ) );
  XOR \SUBBYTES[0].a/U4992  ( .A(\SUBBYTES[0].a/n805 ), .B(
        \SUBBYTES[0].a/n804 ), .Z(\SUBBYTES[0].a/w3313 ) );
  XOR \SUBBYTES[0].a/U4991  ( .A(\SUBBYTES[0].a/n1510 ), .B(
        \SUBBYTES[0].a/n806 ), .Z(\SUBBYTES[0].a/n804 ) );
  XOR \SUBBYTES[0].a/U4990  ( .A(\w1[0][5] ), .B(\SUBBYTES[0].a/n1511 ), .Z(
        \SUBBYTES[0].a/n805 ) );
  XOR \SUBBYTES[0].a/U4989  ( .A(\SUBBYTES[0].a/w3303 ), .B(
        \SUBBYTES[0].a/w3304 ), .Z(\SUBBYTES[0].a/n806 ) );
  XOR \SUBBYTES[0].a/U4988  ( .A(\SUBBYTES[0].a/n808 ), .B(
        \SUBBYTES[0].a/n807 ), .Z(\SUBBYTES[0].a/w3329 ) );
  XOR \SUBBYTES[0].a/U4987  ( .A(\w1[0][1] ), .B(\SUBBYTES[0].a/n809 ), .Z(
        \SUBBYTES[0].a/n807 ) );
  XOR \SUBBYTES[0].a/U4986  ( .A(\SUBBYTES[0].a/w3304 ), .B(
        \SUBBYTES[0].a/w3306 ), .Z(\SUBBYTES[0].a/n808 ) );
  XOR \SUBBYTES[0].a/U4985  ( .A(\SUBBYTES[0].a/w3288 ), .B(
        \SUBBYTES[0].a/w3289 ), .Z(\SUBBYTES[0].a/n809 ) );
  XOR \SUBBYTES[0].a/U4984  ( .A(\w1[0][9] ), .B(\SUBBYTES[0].a/n810 ), .Z(
        \SUBBYTES[0].a/n1512 ) );
  XOR \SUBBYTES[0].a/U4983  ( .A(\w1[0][11] ), .B(\w1[0][10] ), .Z(
        \SUBBYTES[0].a/n810 ) );
  XOR \SUBBYTES[0].a/U4982  ( .A(\w1[0][14] ), .B(\SUBBYTES[0].a/n1512 ), .Z(
        \SUBBYTES[0].a/w3171 ) );
  XOR \SUBBYTES[0].a/U4981  ( .A(\w1[0][8] ), .B(\SUBBYTES[0].a/w3171 ), .Z(
        \SUBBYTES[0].a/w3058 ) );
  XOR \SUBBYTES[0].a/U4980  ( .A(\w1[0][8] ), .B(\SUBBYTES[0].a/n811 ), .Z(
        \SUBBYTES[0].a/w3059 ) );
  XOR \SUBBYTES[0].a/U4979  ( .A(\w1[0][14] ), .B(\w1[0][13] ), .Z(
        \SUBBYTES[0].a/n811 ) );
  XOR \SUBBYTES[0].a/U4978  ( .A(\w1[0][13] ), .B(\SUBBYTES[0].a/n1512 ), .Z(
        \SUBBYTES[0].a/w3189 ) );
  XOR \SUBBYTES[0].a/U4977  ( .A(\SUBBYTES[0].a/n813 ), .B(
        \SUBBYTES[0].a/n812 ), .Z(\SUBBYTES[0].a/w3182 ) );
  XOR \SUBBYTES[0].a/U4976  ( .A(\w1[0][11] ), .B(\w1[0][9] ), .Z(
        \SUBBYTES[0].a/n812 ) );
  XOR \SUBBYTES[0].a/U4975  ( .A(\w1[0][15] ), .B(\w1[0][12] ), .Z(
        \SUBBYTES[0].a/n813 ) );
  XOR \SUBBYTES[0].a/U4974  ( .A(\w1[0][8] ), .B(\SUBBYTES[0].a/w3182 ), .Z(
        \SUBBYTES[0].a/w3061 ) );
  XOR \SUBBYTES[0].a/U4973  ( .A(\SUBBYTES[0].a/n815 ), .B(
        \SUBBYTES[0].a/n814 ), .Z(\SUBBYTES[0].a/w3169 ) );
  XOR \SUBBYTES[0].a/U4972  ( .A(\SUBBYTES[0].a/w3130 ), .B(n1167), .Z(
        \SUBBYTES[0].a/n814 ) );
  XOR \SUBBYTES[0].a/U4971  ( .A(\SUBBYTES[0].a/w3123 ), .B(
        \SUBBYTES[0].a/w3126 ), .Z(\SUBBYTES[0].a/n815 ) );
  XOR \SUBBYTES[0].a/U4970  ( .A(\SUBBYTES[0].a/n817 ), .B(
        \SUBBYTES[0].a/n816 ), .Z(\SUBBYTES[0].a/w3170 ) );
  XOR \SUBBYTES[0].a/U4969  ( .A(\SUBBYTES[0].a/w3130 ), .B(
        \SUBBYTES[0].a/n150 ), .Z(\SUBBYTES[0].a/n816 ) );
  XOR \SUBBYTES[0].a/U4968  ( .A(\SUBBYTES[0].a/w3123 ), .B(
        \SUBBYTES[0].a/n149 ), .Z(\SUBBYTES[0].a/n817 ) );
  XOR \SUBBYTES[0].a/U4967  ( .A(\SUBBYTES[0].a/w3182 ), .B(
        \SUBBYTES[0].a/n818 ), .Z(\SUBBYTES[0].a/w3172 ) );
  XOR \SUBBYTES[0].a/U4966  ( .A(\w1[0][14] ), .B(\w1[0][13] ), .Z(
        \SUBBYTES[0].a/n818 ) );
  XOR \SUBBYTES[0].a/U4965  ( .A(\SUBBYTES[0].a/n820 ), .B(
        \SUBBYTES[0].a/n819 ), .Z(\SUBBYTES[0].a/w3173 ) );
  XOR \SUBBYTES[0].a/U4964  ( .A(\SUBBYTES[0].a/n150 ), .B(n1167), .Z(
        \SUBBYTES[0].a/n819 ) );
  XOR \SUBBYTES[0].a/U4963  ( .A(\SUBBYTES[0].a/n149 ), .B(
        \SUBBYTES[0].a/w3126 ), .Z(\SUBBYTES[0].a/n820 ) );
  XOR \SUBBYTES[0].a/U4962  ( .A(\w1[0][15] ), .B(\w1[0][10] ), .Z(
        \SUBBYTES[0].a/n1518 ) );
  XOR \SUBBYTES[0].a/U4961  ( .A(\SUBBYTES[0].a/n1518 ), .B(
        \SUBBYTES[0].a/n821 ), .Z(\SUBBYTES[0].a/w3174 ) );
  XOR \SUBBYTES[0].a/U4960  ( .A(\w1[0][13] ), .B(\w1[0][12] ), .Z(
        \SUBBYTES[0].a/n821 ) );
  XOR \SUBBYTES[0].a/U4959  ( .A(\w1[0][15] ), .B(\SUBBYTES[0].a/w3059 ), .Z(
        \SUBBYTES[0].a/w3062 ) );
  XOR \SUBBYTES[0].a/U4958  ( .A(\w1[0][9] ), .B(\SUBBYTES[0].a/w3059 ), .Z(
        \SUBBYTES[0].a/w3063 ) );
  XOR \SUBBYTES[0].a/U4957  ( .A(\w1[0][12] ), .B(\SUBBYTES[0].a/w3059 ), .Z(
        \SUBBYTES[0].a/w3064 ) );
  XOR \SUBBYTES[0].a/U4956  ( .A(\SUBBYTES[0].a/w3063 ), .B(
        \SUBBYTES[0].a/n1518 ), .Z(\SUBBYTES[0].a/w3065 ) );
  XOR \SUBBYTES[0].a/U4955  ( .A(\SUBBYTES[0].a/n1518 ), .B(
        \SUBBYTES[0].a/n822 ), .Z(\SUBBYTES[0].a/w3150 ) );
  XOR \SUBBYTES[0].a/U4954  ( .A(\w1[0][12] ), .B(\w1[0][9] ), .Z(
        \SUBBYTES[0].a/n822 ) );
  XOR \SUBBYTES[0].a/U4953  ( .A(\SUBBYTES[0].a/n824 ), .B(
        \SUBBYTES[0].a/n823 ), .Z(\SUBBYTES[0].a/n1515 ) );
  XOR \SUBBYTES[0].a/U4952  ( .A(\w1[0][12] ), .B(\SUBBYTES[0].a/n825 ), .Z(
        \SUBBYTES[0].a/n823 ) );
  XOR \SUBBYTES[0].a/U4951  ( .A(\SUBBYTES[0].a/w3115 ), .B(\w1[0][14] ), .Z(
        \SUBBYTES[0].a/n824 ) );
  XOR \SUBBYTES[0].a/U4950  ( .A(\SUBBYTES[0].a/w3089 ), .B(
        \SUBBYTES[0].a/w3096 ), .Z(\SUBBYTES[0].a/n825 ) );
  XOR \SUBBYTES[0].a/U4949  ( .A(\SUBBYTES[0].a/n827 ), .B(
        \SUBBYTES[0].a/n826 ), .Z(\SUBBYTES[0].a/n1513 ) );
  XOR \SUBBYTES[0].a/U4948  ( .A(\w1[0][9] ), .B(\SUBBYTES[0].a/n828 ), .Z(
        \SUBBYTES[0].a/n826 ) );
  XOR \SUBBYTES[0].a/U4947  ( .A(\SUBBYTES[0].a/w3114 ), .B(\w1[0][13] ), .Z(
        \SUBBYTES[0].a/n827 ) );
  XOR \SUBBYTES[0].a/U4946  ( .A(\SUBBYTES[0].a/w3090 ), .B(
        \SUBBYTES[0].a/w3097 ), .Z(\SUBBYTES[0].a/n828 ) );
  XOR \SUBBYTES[0].a/U4945  ( .A(\SUBBYTES[0].a/n1515 ), .B(
        \SUBBYTES[0].a/n1513 ), .Z(\SUBBYTES[0].a/w3120 ) );
  XOR \SUBBYTES[0].a/U4944  ( .A(\w1[0][13] ), .B(\SUBBYTES[0].a/n829 ), .Z(
        \SUBBYTES[0].a/n1516 ) );
  XOR \SUBBYTES[0].a/U4943  ( .A(\SUBBYTES[0].a/w3082 ), .B(
        \SUBBYTES[0].a/w3092 ), .Z(\SUBBYTES[0].a/n829 ) );
  XOR \SUBBYTES[0].a/U4942  ( .A(\SUBBYTES[0].a/n831 ), .B(
        \SUBBYTES[0].a/n830 ), .Z(\SUBBYTES[0].a/w3107 ) );
  XOR \SUBBYTES[0].a/U4941  ( .A(\SUBBYTES[0].a/n1516 ), .B(
        \SUBBYTES[0].a/n832 ), .Z(\SUBBYTES[0].a/n830 ) );
  XOR \SUBBYTES[0].a/U4940  ( .A(\w1[0][12] ), .B(\SUBBYTES[0].a/w3171 ), .Z(
        \SUBBYTES[0].a/n831 ) );
  XOR \SUBBYTES[0].a/U4939  ( .A(\SUBBYTES[0].a/w3084 ), .B(
        \SUBBYTES[0].a/w3089 ), .Z(\SUBBYTES[0].a/n832 ) );
  XOR \SUBBYTES[0].a/U4938  ( .A(\SUBBYTES[0].a/n834 ), .B(
        \SUBBYTES[0].a/n833 ), .Z(\SUBBYTES[0].a/n1514 ) );
  XOR \SUBBYTES[0].a/U4937  ( .A(\SUBBYTES[0].a/w3117 ), .B(\w1[0][15] ), .Z(
        \SUBBYTES[0].a/n833 ) );
  XOR \SUBBYTES[0].a/U4936  ( .A(\SUBBYTES[0].a/w3092 ), .B(
        \SUBBYTES[0].a/w3099 ), .Z(\SUBBYTES[0].a/n834 ) );
  XOR \SUBBYTES[0].a/U4935  ( .A(\SUBBYTES[0].a/n1513 ), .B(
        \SUBBYTES[0].a/n1514 ), .Z(\SUBBYTES[0].a/w3119 ) );
  XOR \SUBBYTES[0].a/U4934  ( .A(\w1[0][11] ), .B(\SUBBYTES[0].a/n835 ), .Z(
        \SUBBYTES[0].a/n1517 ) );
  XOR \SUBBYTES[0].a/U4933  ( .A(\SUBBYTES[0].a/w3081 ), .B(
        \SUBBYTES[0].a/w3084 ), .Z(\SUBBYTES[0].a/n835 ) );
  XOR \SUBBYTES[0].a/U4932  ( .A(\SUBBYTES[0].a/n837 ), .B(
        \SUBBYTES[0].a/n836 ), .Z(\SUBBYTES[0].a/w3108 ) );
  XOR \SUBBYTES[0].a/U4931  ( .A(\SUBBYTES[0].a/n1517 ), .B(
        \SUBBYTES[0].a/n838 ), .Z(\SUBBYTES[0].a/n836 ) );
  XOR \SUBBYTES[0].a/U4930  ( .A(\w1[0][14] ), .B(\SUBBYTES[0].a/w3150 ), .Z(
        \SUBBYTES[0].a/n837 ) );
  XOR \SUBBYTES[0].a/U4929  ( .A(\SUBBYTES[0].a/w3089 ), .B(
        \SUBBYTES[0].a/w3090 ), .Z(\SUBBYTES[0].a/n838 ) );
  XOR \SUBBYTES[0].a/U4928  ( .A(\SUBBYTES[0].a/n1515 ), .B(
        \SUBBYTES[0].a/n1514 ), .Z(\SUBBYTES[0].a/w3128 ) );
  XOR \SUBBYTES[0].a/U4927  ( .A(\SUBBYTES[0].a/n840 ), .B(
        \SUBBYTES[0].a/n839 ), .Z(\SUBBYTES[0].a/w3129 ) );
  XOR \SUBBYTES[0].a/U4926  ( .A(\w1[0][15] ), .B(\SUBBYTES[0].a/n1516 ), .Z(
        \SUBBYTES[0].a/n839 ) );
  XOR \SUBBYTES[0].a/U4925  ( .A(\SUBBYTES[0].a/w3081 ), .B(
        \SUBBYTES[0].a/w3090 ), .Z(\SUBBYTES[0].a/n840 ) );
  XOR \SUBBYTES[0].a/U4924  ( .A(\SUBBYTES[0].a/n842 ), .B(
        \SUBBYTES[0].a/n841 ), .Z(\SUBBYTES[0].a/w3105 ) );
  XOR \SUBBYTES[0].a/U4923  ( .A(\SUBBYTES[0].a/n844 ), .B(
        \SUBBYTES[0].a/n843 ), .Z(\SUBBYTES[0].a/n841 ) );
  XOR \SUBBYTES[0].a/U4922  ( .A(\w1[0][15] ), .B(\SUBBYTES[0].a/w3189 ), .Z(
        \SUBBYTES[0].a/n842 ) );
  XOR \SUBBYTES[0].a/U4921  ( .A(\SUBBYTES[0].a/w3096 ), .B(
        \SUBBYTES[0].a/w3099 ), .Z(\SUBBYTES[0].a/n843 ) );
  XOR \SUBBYTES[0].a/U4920  ( .A(\SUBBYTES[0].a/w3082 ), .B(
        \SUBBYTES[0].a/w3084 ), .Z(\SUBBYTES[0].a/n844 ) );
  XOR \SUBBYTES[0].a/U4919  ( .A(\SUBBYTES[0].a/n846 ), .B(
        \SUBBYTES[0].a/n845 ), .Z(\SUBBYTES[0].a/w3106 ) );
  XOR \SUBBYTES[0].a/U4918  ( .A(\SUBBYTES[0].a/n1517 ), .B(
        \SUBBYTES[0].a/n847 ), .Z(\SUBBYTES[0].a/n845 ) );
  XOR \SUBBYTES[0].a/U4917  ( .A(\w1[0][13] ), .B(\SUBBYTES[0].a/n1518 ), .Z(
        \SUBBYTES[0].a/n846 ) );
  XOR \SUBBYTES[0].a/U4916  ( .A(\SUBBYTES[0].a/w3096 ), .B(
        \SUBBYTES[0].a/w3097 ), .Z(\SUBBYTES[0].a/n847 ) );
  XOR \SUBBYTES[0].a/U4915  ( .A(\SUBBYTES[0].a/n849 ), .B(
        \SUBBYTES[0].a/n848 ), .Z(\SUBBYTES[0].a/w3122 ) );
  XOR \SUBBYTES[0].a/U4914  ( .A(\w1[0][9] ), .B(\SUBBYTES[0].a/n850 ), .Z(
        \SUBBYTES[0].a/n848 ) );
  XOR \SUBBYTES[0].a/U4913  ( .A(\SUBBYTES[0].a/w3097 ), .B(
        \SUBBYTES[0].a/w3099 ), .Z(\SUBBYTES[0].a/n849 ) );
  XOR \SUBBYTES[0].a/U4912  ( .A(\SUBBYTES[0].a/w3081 ), .B(
        \SUBBYTES[0].a/w3082 ), .Z(\SUBBYTES[0].a/n850 ) );
  XOR \SUBBYTES[0].a/U4911  ( .A(\w1[0][17] ), .B(\SUBBYTES[0].a/n851 ), .Z(
        \SUBBYTES[0].a/n1519 ) );
  XOR \SUBBYTES[0].a/U4910  ( .A(\w1[0][19] ), .B(\w1[0][18] ), .Z(
        \SUBBYTES[0].a/n851 ) );
  XOR \SUBBYTES[0].a/U4909  ( .A(\w1[0][22] ), .B(\SUBBYTES[0].a/n1519 ), .Z(
        \SUBBYTES[0].a/w2964 ) );
  XOR \SUBBYTES[0].a/U4908  ( .A(\w1[0][16] ), .B(\SUBBYTES[0].a/w2964 ), .Z(
        \SUBBYTES[0].a/w2851 ) );
  XOR \SUBBYTES[0].a/U4907  ( .A(\w1[0][16] ), .B(\SUBBYTES[0].a/n852 ), .Z(
        \SUBBYTES[0].a/w2852 ) );
  XOR \SUBBYTES[0].a/U4906  ( .A(\w1[0][22] ), .B(\w1[0][21] ), .Z(
        \SUBBYTES[0].a/n852 ) );
  XOR \SUBBYTES[0].a/U4905  ( .A(\w1[0][21] ), .B(\SUBBYTES[0].a/n1519 ), .Z(
        \SUBBYTES[0].a/w2982 ) );
  XOR \SUBBYTES[0].a/U4904  ( .A(\SUBBYTES[0].a/n854 ), .B(
        \SUBBYTES[0].a/n853 ), .Z(\SUBBYTES[0].a/w2975 ) );
  XOR \SUBBYTES[0].a/U4903  ( .A(\w1[0][19] ), .B(\w1[0][17] ), .Z(
        \SUBBYTES[0].a/n853 ) );
  XOR \SUBBYTES[0].a/U4902  ( .A(\w1[0][23] ), .B(\w1[0][20] ), .Z(
        \SUBBYTES[0].a/n854 ) );
  XOR \SUBBYTES[0].a/U4901  ( .A(\w1[0][16] ), .B(\SUBBYTES[0].a/w2975 ), .Z(
        \SUBBYTES[0].a/w2854 ) );
  XOR \SUBBYTES[0].a/U4900  ( .A(\SUBBYTES[0].a/n856 ), .B(
        \SUBBYTES[0].a/n855 ), .Z(\SUBBYTES[0].a/w2962 ) );
  XOR \SUBBYTES[0].a/U4899  ( .A(\SUBBYTES[0].a/w2923 ), .B(n1166), .Z(
        \SUBBYTES[0].a/n855 ) );
  XOR \SUBBYTES[0].a/U4898  ( .A(\SUBBYTES[0].a/w2916 ), .B(
        \SUBBYTES[0].a/w2919 ), .Z(\SUBBYTES[0].a/n856 ) );
  XOR \SUBBYTES[0].a/U4897  ( .A(\SUBBYTES[0].a/n858 ), .B(
        \SUBBYTES[0].a/n857 ), .Z(\SUBBYTES[0].a/w2963 ) );
  XOR \SUBBYTES[0].a/U4896  ( .A(\SUBBYTES[0].a/w2923 ), .B(
        \SUBBYTES[0].a/n140 ), .Z(\SUBBYTES[0].a/n857 ) );
  XOR \SUBBYTES[0].a/U4895  ( .A(\SUBBYTES[0].a/w2916 ), .B(
        \SUBBYTES[0].a/n139 ), .Z(\SUBBYTES[0].a/n858 ) );
  XOR \SUBBYTES[0].a/U4894  ( .A(\SUBBYTES[0].a/w2975 ), .B(
        \SUBBYTES[0].a/n859 ), .Z(\SUBBYTES[0].a/w2965 ) );
  XOR \SUBBYTES[0].a/U4893  ( .A(\w1[0][22] ), .B(\w1[0][21] ), .Z(
        \SUBBYTES[0].a/n859 ) );
  XOR \SUBBYTES[0].a/U4892  ( .A(\SUBBYTES[0].a/n861 ), .B(
        \SUBBYTES[0].a/n860 ), .Z(\SUBBYTES[0].a/w2966 ) );
  XOR \SUBBYTES[0].a/U4891  ( .A(\SUBBYTES[0].a/n140 ), .B(n1166), .Z(
        \SUBBYTES[0].a/n860 ) );
  XOR \SUBBYTES[0].a/U4890  ( .A(\SUBBYTES[0].a/n139 ), .B(
        \SUBBYTES[0].a/w2919 ), .Z(\SUBBYTES[0].a/n861 ) );
  XOR \SUBBYTES[0].a/U4889  ( .A(\w1[0][23] ), .B(\w1[0][18] ), .Z(
        \SUBBYTES[0].a/n1525 ) );
  XOR \SUBBYTES[0].a/U4888  ( .A(\SUBBYTES[0].a/n1525 ), .B(
        \SUBBYTES[0].a/n862 ), .Z(\SUBBYTES[0].a/w2967 ) );
  XOR \SUBBYTES[0].a/U4887  ( .A(\w1[0][21] ), .B(\w1[0][20] ), .Z(
        \SUBBYTES[0].a/n862 ) );
  XOR \SUBBYTES[0].a/U4886  ( .A(\w1[0][23] ), .B(\SUBBYTES[0].a/w2852 ), .Z(
        \SUBBYTES[0].a/w2855 ) );
  XOR \SUBBYTES[0].a/U4885  ( .A(\w1[0][17] ), .B(\SUBBYTES[0].a/w2852 ), .Z(
        \SUBBYTES[0].a/w2856 ) );
  XOR \SUBBYTES[0].a/U4884  ( .A(\w1[0][20] ), .B(\SUBBYTES[0].a/w2852 ), .Z(
        \SUBBYTES[0].a/w2857 ) );
  XOR \SUBBYTES[0].a/U4883  ( .A(\SUBBYTES[0].a/w2856 ), .B(
        \SUBBYTES[0].a/n1525 ), .Z(\SUBBYTES[0].a/w2858 ) );
  XOR \SUBBYTES[0].a/U4882  ( .A(\SUBBYTES[0].a/n1525 ), .B(
        \SUBBYTES[0].a/n863 ), .Z(\SUBBYTES[0].a/w2943 ) );
  XOR \SUBBYTES[0].a/U4881  ( .A(\w1[0][20] ), .B(\w1[0][17] ), .Z(
        \SUBBYTES[0].a/n863 ) );
  XOR \SUBBYTES[0].a/U4880  ( .A(\SUBBYTES[0].a/n865 ), .B(
        \SUBBYTES[0].a/n864 ), .Z(\SUBBYTES[0].a/n1522 ) );
  XOR \SUBBYTES[0].a/U4879  ( .A(\w1[0][20] ), .B(\SUBBYTES[0].a/n866 ), .Z(
        \SUBBYTES[0].a/n864 ) );
  XOR \SUBBYTES[0].a/U4878  ( .A(\SUBBYTES[0].a/w2908 ), .B(\w1[0][22] ), .Z(
        \SUBBYTES[0].a/n865 ) );
  XOR \SUBBYTES[0].a/U4877  ( .A(\SUBBYTES[0].a/w2882 ), .B(
        \SUBBYTES[0].a/w2889 ), .Z(\SUBBYTES[0].a/n866 ) );
  XOR \SUBBYTES[0].a/U4876  ( .A(\SUBBYTES[0].a/n868 ), .B(
        \SUBBYTES[0].a/n867 ), .Z(\SUBBYTES[0].a/n1520 ) );
  XOR \SUBBYTES[0].a/U4875  ( .A(\w1[0][17] ), .B(\SUBBYTES[0].a/n869 ), .Z(
        \SUBBYTES[0].a/n867 ) );
  XOR \SUBBYTES[0].a/U4874  ( .A(\SUBBYTES[0].a/w2907 ), .B(\w1[0][21] ), .Z(
        \SUBBYTES[0].a/n868 ) );
  XOR \SUBBYTES[0].a/U4873  ( .A(\SUBBYTES[0].a/w2883 ), .B(
        \SUBBYTES[0].a/w2890 ), .Z(\SUBBYTES[0].a/n869 ) );
  XOR \SUBBYTES[0].a/U4872  ( .A(\SUBBYTES[0].a/n1522 ), .B(
        \SUBBYTES[0].a/n1520 ), .Z(\SUBBYTES[0].a/w2913 ) );
  XOR \SUBBYTES[0].a/U4871  ( .A(\w1[0][21] ), .B(\SUBBYTES[0].a/n870 ), .Z(
        \SUBBYTES[0].a/n1523 ) );
  XOR \SUBBYTES[0].a/U4870  ( .A(\SUBBYTES[0].a/w2875 ), .B(
        \SUBBYTES[0].a/w2885 ), .Z(\SUBBYTES[0].a/n870 ) );
  XOR \SUBBYTES[0].a/U4869  ( .A(\SUBBYTES[0].a/n872 ), .B(
        \SUBBYTES[0].a/n871 ), .Z(\SUBBYTES[0].a/w2900 ) );
  XOR \SUBBYTES[0].a/U4868  ( .A(\SUBBYTES[0].a/n1523 ), .B(
        \SUBBYTES[0].a/n873 ), .Z(\SUBBYTES[0].a/n871 ) );
  XOR \SUBBYTES[0].a/U4867  ( .A(\w1[0][20] ), .B(\SUBBYTES[0].a/w2964 ), .Z(
        \SUBBYTES[0].a/n872 ) );
  XOR \SUBBYTES[0].a/U4866  ( .A(\SUBBYTES[0].a/w2877 ), .B(
        \SUBBYTES[0].a/w2882 ), .Z(\SUBBYTES[0].a/n873 ) );
  XOR \SUBBYTES[0].a/U4865  ( .A(\SUBBYTES[0].a/n875 ), .B(
        \SUBBYTES[0].a/n874 ), .Z(\SUBBYTES[0].a/n1521 ) );
  XOR \SUBBYTES[0].a/U4864  ( .A(\SUBBYTES[0].a/w2910 ), .B(\w1[0][23] ), .Z(
        \SUBBYTES[0].a/n874 ) );
  XOR \SUBBYTES[0].a/U4863  ( .A(\SUBBYTES[0].a/w2885 ), .B(
        \SUBBYTES[0].a/w2892 ), .Z(\SUBBYTES[0].a/n875 ) );
  XOR \SUBBYTES[0].a/U4862  ( .A(\SUBBYTES[0].a/n1520 ), .B(
        \SUBBYTES[0].a/n1521 ), .Z(\SUBBYTES[0].a/w2912 ) );
  XOR \SUBBYTES[0].a/U4861  ( .A(\w1[0][19] ), .B(\SUBBYTES[0].a/n876 ), .Z(
        \SUBBYTES[0].a/n1524 ) );
  XOR \SUBBYTES[0].a/U4860  ( .A(\SUBBYTES[0].a/w2874 ), .B(
        \SUBBYTES[0].a/w2877 ), .Z(\SUBBYTES[0].a/n876 ) );
  XOR \SUBBYTES[0].a/U4859  ( .A(\SUBBYTES[0].a/n878 ), .B(
        \SUBBYTES[0].a/n877 ), .Z(\SUBBYTES[0].a/w2901 ) );
  XOR \SUBBYTES[0].a/U4858  ( .A(\SUBBYTES[0].a/n1524 ), .B(
        \SUBBYTES[0].a/n879 ), .Z(\SUBBYTES[0].a/n877 ) );
  XOR \SUBBYTES[0].a/U4857  ( .A(\w1[0][22] ), .B(\SUBBYTES[0].a/w2943 ), .Z(
        \SUBBYTES[0].a/n878 ) );
  XOR \SUBBYTES[0].a/U4856  ( .A(\SUBBYTES[0].a/w2882 ), .B(
        \SUBBYTES[0].a/w2883 ), .Z(\SUBBYTES[0].a/n879 ) );
  XOR \SUBBYTES[0].a/U4855  ( .A(\SUBBYTES[0].a/n1522 ), .B(
        \SUBBYTES[0].a/n1521 ), .Z(\SUBBYTES[0].a/w2921 ) );
  XOR \SUBBYTES[0].a/U4854  ( .A(\SUBBYTES[0].a/n881 ), .B(
        \SUBBYTES[0].a/n880 ), .Z(\SUBBYTES[0].a/w2922 ) );
  XOR \SUBBYTES[0].a/U4853  ( .A(\w1[0][23] ), .B(\SUBBYTES[0].a/n1523 ), .Z(
        \SUBBYTES[0].a/n880 ) );
  XOR \SUBBYTES[0].a/U4852  ( .A(\SUBBYTES[0].a/w2874 ), .B(
        \SUBBYTES[0].a/w2883 ), .Z(\SUBBYTES[0].a/n881 ) );
  XOR \SUBBYTES[0].a/U4851  ( .A(\SUBBYTES[0].a/n883 ), .B(
        \SUBBYTES[0].a/n882 ), .Z(\SUBBYTES[0].a/w2898 ) );
  XOR \SUBBYTES[0].a/U4850  ( .A(\SUBBYTES[0].a/n885 ), .B(
        \SUBBYTES[0].a/n884 ), .Z(\SUBBYTES[0].a/n882 ) );
  XOR \SUBBYTES[0].a/U4849  ( .A(\w1[0][23] ), .B(\SUBBYTES[0].a/w2982 ), .Z(
        \SUBBYTES[0].a/n883 ) );
  XOR \SUBBYTES[0].a/U4848  ( .A(\SUBBYTES[0].a/w2889 ), .B(
        \SUBBYTES[0].a/w2892 ), .Z(\SUBBYTES[0].a/n884 ) );
  XOR \SUBBYTES[0].a/U4847  ( .A(\SUBBYTES[0].a/w2875 ), .B(
        \SUBBYTES[0].a/w2877 ), .Z(\SUBBYTES[0].a/n885 ) );
  XOR \SUBBYTES[0].a/U4846  ( .A(\SUBBYTES[0].a/n887 ), .B(
        \SUBBYTES[0].a/n886 ), .Z(\SUBBYTES[0].a/w2899 ) );
  XOR \SUBBYTES[0].a/U4845  ( .A(\SUBBYTES[0].a/n1524 ), .B(
        \SUBBYTES[0].a/n888 ), .Z(\SUBBYTES[0].a/n886 ) );
  XOR \SUBBYTES[0].a/U4844  ( .A(\w1[0][21] ), .B(\SUBBYTES[0].a/n1525 ), .Z(
        \SUBBYTES[0].a/n887 ) );
  XOR \SUBBYTES[0].a/U4843  ( .A(\SUBBYTES[0].a/w2889 ), .B(
        \SUBBYTES[0].a/w2890 ), .Z(\SUBBYTES[0].a/n888 ) );
  XOR \SUBBYTES[0].a/U4842  ( .A(\SUBBYTES[0].a/n890 ), .B(
        \SUBBYTES[0].a/n889 ), .Z(\SUBBYTES[0].a/w2915 ) );
  XOR \SUBBYTES[0].a/U4841  ( .A(\w1[0][17] ), .B(\SUBBYTES[0].a/n891 ), .Z(
        \SUBBYTES[0].a/n889 ) );
  XOR \SUBBYTES[0].a/U4840  ( .A(\SUBBYTES[0].a/w2890 ), .B(
        \SUBBYTES[0].a/w2892 ), .Z(\SUBBYTES[0].a/n890 ) );
  XOR \SUBBYTES[0].a/U4839  ( .A(\SUBBYTES[0].a/w2874 ), .B(
        \SUBBYTES[0].a/w2875 ), .Z(\SUBBYTES[0].a/n891 ) );
  XOR \SUBBYTES[0].a/U4838  ( .A(\w1[0][25] ), .B(\SUBBYTES[0].a/n892 ), .Z(
        \SUBBYTES[0].a/n1526 ) );
  XOR \SUBBYTES[0].a/U4837  ( .A(\w1[0][27] ), .B(\w1[0][26] ), .Z(
        \SUBBYTES[0].a/n892 ) );
  XOR \SUBBYTES[0].a/U4836  ( .A(\w1[0][30] ), .B(\SUBBYTES[0].a/n1526 ), .Z(
        \SUBBYTES[0].a/w2757 ) );
  XOR \SUBBYTES[0].a/U4835  ( .A(\w1[0][24] ), .B(\SUBBYTES[0].a/w2757 ), .Z(
        \SUBBYTES[0].a/w2644 ) );
  XOR \SUBBYTES[0].a/U4834  ( .A(\w1[0][24] ), .B(\SUBBYTES[0].a/n893 ), .Z(
        \SUBBYTES[0].a/w2645 ) );
  XOR \SUBBYTES[0].a/U4833  ( .A(\w1[0][30] ), .B(\w1[0][29] ), .Z(
        \SUBBYTES[0].a/n893 ) );
  XOR \SUBBYTES[0].a/U4832  ( .A(\w1[0][29] ), .B(\SUBBYTES[0].a/n1526 ), .Z(
        \SUBBYTES[0].a/w2775 ) );
  XOR \SUBBYTES[0].a/U4831  ( .A(\SUBBYTES[0].a/n895 ), .B(
        \SUBBYTES[0].a/n894 ), .Z(\SUBBYTES[0].a/w2768 ) );
  XOR \SUBBYTES[0].a/U4830  ( .A(\w1[0][27] ), .B(\w1[0][25] ), .Z(
        \SUBBYTES[0].a/n894 ) );
  XOR \SUBBYTES[0].a/U4829  ( .A(\w1[0][31] ), .B(\w1[0][28] ), .Z(
        \SUBBYTES[0].a/n895 ) );
  XOR \SUBBYTES[0].a/U4828  ( .A(\w1[0][24] ), .B(\SUBBYTES[0].a/w2768 ), .Z(
        \SUBBYTES[0].a/w2647 ) );
  XOR \SUBBYTES[0].a/U4827  ( .A(\SUBBYTES[0].a/n897 ), .B(
        \SUBBYTES[0].a/n896 ), .Z(\SUBBYTES[0].a/w2755 ) );
  XOR \SUBBYTES[0].a/U4826  ( .A(\SUBBYTES[0].a/w2716 ), .B(n1165), .Z(
        \SUBBYTES[0].a/n896 ) );
  XOR \SUBBYTES[0].a/U4825  ( .A(\SUBBYTES[0].a/w2709 ), .B(
        \SUBBYTES[0].a/w2712 ), .Z(\SUBBYTES[0].a/n897 ) );
  XOR \SUBBYTES[0].a/U4824  ( .A(\SUBBYTES[0].a/n899 ), .B(
        \SUBBYTES[0].a/n898 ), .Z(\SUBBYTES[0].a/w2756 ) );
  XOR \SUBBYTES[0].a/U4823  ( .A(\SUBBYTES[0].a/w2716 ), .B(
        \SUBBYTES[0].a/n130 ), .Z(\SUBBYTES[0].a/n898 ) );
  XOR \SUBBYTES[0].a/U4822  ( .A(\SUBBYTES[0].a/w2709 ), .B(
        \SUBBYTES[0].a/n129 ), .Z(\SUBBYTES[0].a/n899 ) );
  XOR \SUBBYTES[0].a/U4821  ( .A(\SUBBYTES[0].a/w2768 ), .B(
        \SUBBYTES[0].a/n900 ), .Z(\SUBBYTES[0].a/w2758 ) );
  XOR \SUBBYTES[0].a/U4820  ( .A(\w1[0][30] ), .B(\w1[0][29] ), .Z(
        \SUBBYTES[0].a/n900 ) );
  XOR \SUBBYTES[0].a/U4819  ( .A(\SUBBYTES[0].a/n902 ), .B(
        \SUBBYTES[0].a/n901 ), .Z(\SUBBYTES[0].a/w2759 ) );
  XOR \SUBBYTES[0].a/U4818  ( .A(\SUBBYTES[0].a/n130 ), .B(n1165), .Z(
        \SUBBYTES[0].a/n901 ) );
  XOR \SUBBYTES[0].a/U4817  ( .A(\SUBBYTES[0].a/n129 ), .B(
        \SUBBYTES[0].a/w2712 ), .Z(\SUBBYTES[0].a/n902 ) );
  XOR \SUBBYTES[0].a/U4816  ( .A(\w1[0][31] ), .B(\w1[0][26] ), .Z(
        \SUBBYTES[0].a/n1532 ) );
  XOR \SUBBYTES[0].a/U4815  ( .A(\SUBBYTES[0].a/n1532 ), .B(
        \SUBBYTES[0].a/n903 ), .Z(\SUBBYTES[0].a/w2760 ) );
  XOR \SUBBYTES[0].a/U4814  ( .A(\w1[0][29] ), .B(\w1[0][28] ), .Z(
        \SUBBYTES[0].a/n903 ) );
  XOR \SUBBYTES[0].a/U4813  ( .A(\w1[0][31] ), .B(\SUBBYTES[0].a/w2645 ), .Z(
        \SUBBYTES[0].a/w2648 ) );
  XOR \SUBBYTES[0].a/U4812  ( .A(\w1[0][25] ), .B(\SUBBYTES[0].a/w2645 ), .Z(
        \SUBBYTES[0].a/w2649 ) );
  XOR \SUBBYTES[0].a/U4811  ( .A(\w1[0][28] ), .B(\SUBBYTES[0].a/w2645 ), .Z(
        \SUBBYTES[0].a/w2650 ) );
  XOR \SUBBYTES[0].a/U4810  ( .A(\SUBBYTES[0].a/w2649 ), .B(
        \SUBBYTES[0].a/n1532 ), .Z(\SUBBYTES[0].a/w2651 ) );
  XOR \SUBBYTES[0].a/U4809  ( .A(\SUBBYTES[0].a/n1532 ), .B(
        \SUBBYTES[0].a/n904 ), .Z(\SUBBYTES[0].a/w2736 ) );
  XOR \SUBBYTES[0].a/U4808  ( .A(\w1[0][28] ), .B(\w1[0][25] ), .Z(
        \SUBBYTES[0].a/n904 ) );
  XOR \SUBBYTES[0].a/U4807  ( .A(\SUBBYTES[0].a/n906 ), .B(
        \SUBBYTES[0].a/n905 ), .Z(\SUBBYTES[0].a/n1529 ) );
  XOR \SUBBYTES[0].a/U4806  ( .A(\w1[0][28] ), .B(\SUBBYTES[0].a/n907 ), .Z(
        \SUBBYTES[0].a/n905 ) );
  XOR \SUBBYTES[0].a/U4805  ( .A(\SUBBYTES[0].a/w2701 ), .B(\w1[0][30] ), .Z(
        \SUBBYTES[0].a/n906 ) );
  XOR \SUBBYTES[0].a/U4804  ( .A(\SUBBYTES[0].a/w2675 ), .B(
        \SUBBYTES[0].a/w2682 ), .Z(\SUBBYTES[0].a/n907 ) );
  XOR \SUBBYTES[0].a/U4803  ( .A(\SUBBYTES[0].a/n909 ), .B(
        \SUBBYTES[0].a/n908 ), .Z(\SUBBYTES[0].a/n1527 ) );
  XOR \SUBBYTES[0].a/U4802  ( .A(\w1[0][25] ), .B(\SUBBYTES[0].a/n910 ), .Z(
        \SUBBYTES[0].a/n908 ) );
  XOR \SUBBYTES[0].a/U4801  ( .A(\SUBBYTES[0].a/w2700 ), .B(\w1[0][29] ), .Z(
        \SUBBYTES[0].a/n909 ) );
  XOR \SUBBYTES[0].a/U4800  ( .A(\SUBBYTES[0].a/w2676 ), .B(
        \SUBBYTES[0].a/w2683 ), .Z(\SUBBYTES[0].a/n910 ) );
  XOR \SUBBYTES[0].a/U4799  ( .A(\SUBBYTES[0].a/n1529 ), .B(
        \SUBBYTES[0].a/n1527 ), .Z(\SUBBYTES[0].a/w2706 ) );
  XOR \SUBBYTES[0].a/U4798  ( .A(\w1[0][29] ), .B(\SUBBYTES[0].a/n911 ), .Z(
        \SUBBYTES[0].a/n1530 ) );
  XOR \SUBBYTES[0].a/U4797  ( .A(\SUBBYTES[0].a/w2668 ), .B(
        \SUBBYTES[0].a/w2678 ), .Z(\SUBBYTES[0].a/n911 ) );
  XOR \SUBBYTES[0].a/U4796  ( .A(\SUBBYTES[0].a/n913 ), .B(
        \SUBBYTES[0].a/n912 ), .Z(\SUBBYTES[0].a/w2693 ) );
  XOR \SUBBYTES[0].a/U4795  ( .A(\SUBBYTES[0].a/n1530 ), .B(
        \SUBBYTES[0].a/n914 ), .Z(\SUBBYTES[0].a/n912 ) );
  XOR \SUBBYTES[0].a/U4794  ( .A(\w1[0][28] ), .B(\SUBBYTES[0].a/w2757 ), .Z(
        \SUBBYTES[0].a/n913 ) );
  XOR \SUBBYTES[0].a/U4793  ( .A(\SUBBYTES[0].a/w2670 ), .B(
        \SUBBYTES[0].a/w2675 ), .Z(\SUBBYTES[0].a/n914 ) );
  XOR \SUBBYTES[0].a/U4792  ( .A(\SUBBYTES[0].a/n916 ), .B(
        \SUBBYTES[0].a/n915 ), .Z(\SUBBYTES[0].a/n1528 ) );
  XOR \SUBBYTES[0].a/U4791  ( .A(\SUBBYTES[0].a/w2703 ), .B(\w1[0][31] ), .Z(
        \SUBBYTES[0].a/n915 ) );
  XOR \SUBBYTES[0].a/U4790  ( .A(\SUBBYTES[0].a/w2678 ), .B(
        \SUBBYTES[0].a/w2685 ), .Z(\SUBBYTES[0].a/n916 ) );
  XOR \SUBBYTES[0].a/U4789  ( .A(\SUBBYTES[0].a/n1527 ), .B(
        \SUBBYTES[0].a/n1528 ), .Z(\SUBBYTES[0].a/w2705 ) );
  XOR \SUBBYTES[0].a/U4788  ( .A(\w1[0][27] ), .B(\SUBBYTES[0].a/n917 ), .Z(
        \SUBBYTES[0].a/n1531 ) );
  XOR \SUBBYTES[0].a/U4787  ( .A(\SUBBYTES[0].a/w2667 ), .B(
        \SUBBYTES[0].a/w2670 ), .Z(\SUBBYTES[0].a/n917 ) );
  XOR \SUBBYTES[0].a/U4786  ( .A(\SUBBYTES[0].a/n919 ), .B(
        \SUBBYTES[0].a/n918 ), .Z(\SUBBYTES[0].a/w2694 ) );
  XOR \SUBBYTES[0].a/U4785  ( .A(\SUBBYTES[0].a/n1531 ), .B(
        \SUBBYTES[0].a/n920 ), .Z(\SUBBYTES[0].a/n918 ) );
  XOR \SUBBYTES[0].a/U4784  ( .A(\w1[0][30] ), .B(\SUBBYTES[0].a/w2736 ), .Z(
        \SUBBYTES[0].a/n919 ) );
  XOR \SUBBYTES[0].a/U4783  ( .A(\SUBBYTES[0].a/w2675 ), .B(
        \SUBBYTES[0].a/w2676 ), .Z(\SUBBYTES[0].a/n920 ) );
  XOR \SUBBYTES[0].a/U4782  ( .A(\SUBBYTES[0].a/n1529 ), .B(
        \SUBBYTES[0].a/n1528 ), .Z(\SUBBYTES[0].a/w2714 ) );
  XOR \SUBBYTES[0].a/U4781  ( .A(\SUBBYTES[0].a/n922 ), .B(
        \SUBBYTES[0].a/n921 ), .Z(\SUBBYTES[0].a/w2715 ) );
  XOR \SUBBYTES[0].a/U4780  ( .A(\w1[0][31] ), .B(\SUBBYTES[0].a/n1530 ), .Z(
        \SUBBYTES[0].a/n921 ) );
  XOR \SUBBYTES[0].a/U4779  ( .A(\SUBBYTES[0].a/w2667 ), .B(
        \SUBBYTES[0].a/w2676 ), .Z(\SUBBYTES[0].a/n922 ) );
  XOR \SUBBYTES[0].a/U4778  ( .A(\SUBBYTES[0].a/n924 ), .B(
        \SUBBYTES[0].a/n923 ), .Z(\SUBBYTES[0].a/w2691 ) );
  XOR \SUBBYTES[0].a/U4777  ( .A(\SUBBYTES[0].a/n926 ), .B(
        \SUBBYTES[0].a/n925 ), .Z(\SUBBYTES[0].a/n923 ) );
  XOR \SUBBYTES[0].a/U4776  ( .A(\w1[0][31] ), .B(\SUBBYTES[0].a/w2775 ), .Z(
        \SUBBYTES[0].a/n924 ) );
  XOR \SUBBYTES[0].a/U4775  ( .A(\SUBBYTES[0].a/w2682 ), .B(
        \SUBBYTES[0].a/w2685 ), .Z(\SUBBYTES[0].a/n925 ) );
  XOR \SUBBYTES[0].a/U4774  ( .A(\SUBBYTES[0].a/w2668 ), .B(
        \SUBBYTES[0].a/w2670 ), .Z(\SUBBYTES[0].a/n926 ) );
  XOR \SUBBYTES[0].a/U4773  ( .A(\SUBBYTES[0].a/n928 ), .B(
        \SUBBYTES[0].a/n927 ), .Z(\SUBBYTES[0].a/w2692 ) );
  XOR \SUBBYTES[0].a/U4772  ( .A(\SUBBYTES[0].a/n1531 ), .B(
        \SUBBYTES[0].a/n929 ), .Z(\SUBBYTES[0].a/n927 ) );
  XOR \SUBBYTES[0].a/U4771  ( .A(\w1[0][29] ), .B(\SUBBYTES[0].a/n1532 ), .Z(
        \SUBBYTES[0].a/n928 ) );
  XOR \SUBBYTES[0].a/U4770  ( .A(\SUBBYTES[0].a/w2682 ), .B(
        \SUBBYTES[0].a/w2683 ), .Z(\SUBBYTES[0].a/n929 ) );
  XOR \SUBBYTES[0].a/U4769  ( .A(\SUBBYTES[0].a/n931 ), .B(
        \SUBBYTES[0].a/n930 ), .Z(\SUBBYTES[0].a/w2708 ) );
  XOR \SUBBYTES[0].a/U4768  ( .A(\w1[0][25] ), .B(\SUBBYTES[0].a/n932 ), .Z(
        \SUBBYTES[0].a/n930 ) );
  XOR \SUBBYTES[0].a/U4767  ( .A(\SUBBYTES[0].a/w2683 ), .B(
        \SUBBYTES[0].a/w2685 ), .Z(\SUBBYTES[0].a/n931 ) );
  XOR \SUBBYTES[0].a/U4766  ( .A(\SUBBYTES[0].a/w2667 ), .B(
        \SUBBYTES[0].a/w2668 ), .Z(\SUBBYTES[0].a/n932 ) );
  XOR \SUBBYTES[0].a/U4765  ( .A(\w1[0][33] ), .B(\SUBBYTES[0].a/n933 ), .Z(
        \SUBBYTES[0].a/n1533 ) );
  XOR \SUBBYTES[0].a/U4764  ( .A(\w1[0][35] ), .B(\w1[0][34] ), .Z(
        \SUBBYTES[0].a/n933 ) );
  XOR \SUBBYTES[0].a/U4763  ( .A(\w1[0][38] ), .B(\SUBBYTES[0].a/n1533 ), .Z(
        \SUBBYTES[0].a/w2550 ) );
  XOR \SUBBYTES[0].a/U4762  ( .A(\w1[0][32] ), .B(\SUBBYTES[0].a/w2550 ), .Z(
        \SUBBYTES[0].a/w2437 ) );
  XOR \SUBBYTES[0].a/U4761  ( .A(\w1[0][32] ), .B(\SUBBYTES[0].a/n934 ), .Z(
        \SUBBYTES[0].a/w2438 ) );
  XOR \SUBBYTES[0].a/U4760  ( .A(\w1[0][38] ), .B(\w1[0][37] ), .Z(
        \SUBBYTES[0].a/n934 ) );
  XOR \SUBBYTES[0].a/U4759  ( .A(\w1[0][37] ), .B(\SUBBYTES[0].a/n1533 ), .Z(
        \SUBBYTES[0].a/w2568 ) );
  XOR \SUBBYTES[0].a/U4758  ( .A(\SUBBYTES[0].a/n936 ), .B(
        \SUBBYTES[0].a/n935 ), .Z(\SUBBYTES[0].a/w2561 ) );
  XOR \SUBBYTES[0].a/U4757  ( .A(\w1[0][35] ), .B(\w1[0][33] ), .Z(
        \SUBBYTES[0].a/n935 ) );
  XOR \SUBBYTES[0].a/U4756  ( .A(\w1[0][39] ), .B(\w1[0][36] ), .Z(
        \SUBBYTES[0].a/n936 ) );
  XOR \SUBBYTES[0].a/U4755  ( .A(\w1[0][32] ), .B(\SUBBYTES[0].a/w2561 ), .Z(
        \SUBBYTES[0].a/w2440 ) );
  XOR \SUBBYTES[0].a/U4754  ( .A(\SUBBYTES[0].a/n938 ), .B(
        \SUBBYTES[0].a/n937 ), .Z(\SUBBYTES[0].a/w2548 ) );
  XOR \SUBBYTES[0].a/U4753  ( .A(\SUBBYTES[0].a/w2509 ), .B(n1164), .Z(
        \SUBBYTES[0].a/n937 ) );
  XOR \SUBBYTES[0].a/U4752  ( .A(\SUBBYTES[0].a/w2502 ), .B(
        \SUBBYTES[0].a/w2505 ), .Z(\SUBBYTES[0].a/n938 ) );
  XOR \SUBBYTES[0].a/U4751  ( .A(\SUBBYTES[0].a/n940 ), .B(
        \SUBBYTES[0].a/n939 ), .Z(\SUBBYTES[0].a/w2549 ) );
  XOR \SUBBYTES[0].a/U4750  ( .A(\SUBBYTES[0].a/w2509 ), .B(
        \SUBBYTES[0].a/n120 ), .Z(\SUBBYTES[0].a/n939 ) );
  XOR \SUBBYTES[0].a/U4749  ( .A(\SUBBYTES[0].a/w2502 ), .B(
        \SUBBYTES[0].a/n119 ), .Z(\SUBBYTES[0].a/n940 ) );
  XOR \SUBBYTES[0].a/U4748  ( .A(\SUBBYTES[0].a/w2561 ), .B(
        \SUBBYTES[0].a/n941 ), .Z(\SUBBYTES[0].a/w2551 ) );
  XOR \SUBBYTES[0].a/U4747  ( .A(\w1[0][38] ), .B(\w1[0][37] ), .Z(
        \SUBBYTES[0].a/n941 ) );
  XOR \SUBBYTES[0].a/U4746  ( .A(\SUBBYTES[0].a/n943 ), .B(
        \SUBBYTES[0].a/n942 ), .Z(\SUBBYTES[0].a/w2552 ) );
  XOR \SUBBYTES[0].a/U4745  ( .A(\SUBBYTES[0].a/n120 ), .B(n1164), .Z(
        \SUBBYTES[0].a/n942 ) );
  XOR \SUBBYTES[0].a/U4744  ( .A(\SUBBYTES[0].a/n119 ), .B(
        \SUBBYTES[0].a/w2505 ), .Z(\SUBBYTES[0].a/n943 ) );
  XOR \SUBBYTES[0].a/U4743  ( .A(\w1[0][39] ), .B(\w1[0][34] ), .Z(
        \SUBBYTES[0].a/n1539 ) );
  XOR \SUBBYTES[0].a/U4742  ( .A(\SUBBYTES[0].a/n1539 ), .B(
        \SUBBYTES[0].a/n944 ), .Z(\SUBBYTES[0].a/w2553 ) );
  XOR \SUBBYTES[0].a/U4741  ( .A(\w1[0][37] ), .B(\w1[0][36] ), .Z(
        \SUBBYTES[0].a/n944 ) );
  XOR \SUBBYTES[0].a/U4740  ( .A(\w1[0][39] ), .B(\SUBBYTES[0].a/w2438 ), .Z(
        \SUBBYTES[0].a/w2441 ) );
  XOR \SUBBYTES[0].a/U4739  ( .A(\w1[0][33] ), .B(\SUBBYTES[0].a/w2438 ), .Z(
        \SUBBYTES[0].a/w2442 ) );
  XOR \SUBBYTES[0].a/U4738  ( .A(\w1[0][36] ), .B(\SUBBYTES[0].a/w2438 ), .Z(
        \SUBBYTES[0].a/w2443 ) );
  XOR \SUBBYTES[0].a/U4737  ( .A(\SUBBYTES[0].a/w2442 ), .B(
        \SUBBYTES[0].a/n1539 ), .Z(\SUBBYTES[0].a/w2444 ) );
  XOR \SUBBYTES[0].a/U4736  ( .A(\SUBBYTES[0].a/n1539 ), .B(
        \SUBBYTES[0].a/n945 ), .Z(\SUBBYTES[0].a/w2529 ) );
  XOR \SUBBYTES[0].a/U4735  ( .A(\w1[0][36] ), .B(\w1[0][33] ), .Z(
        \SUBBYTES[0].a/n945 ) );
  XOR \SUBBYTES[0].a/U4734  ( .A(\SUBBYTES[0].a/n947 ), .B(
        \SUBBYTES[0].a/n946 ), .Z(\SUBBYTES[0].a/n1536 ) );
  XOR \SUBBYTES[0].a/U4733  ( .A(\w1[0][36] ), .B(\SUBBYTES[0].a/n948 ), .Z(
        \SUBBYTES[0].a/n946 ) );
  XOR \SUBBYTES[0].a/U4732  ( .A(\SUBBYTES[0].a/w2494 ), .B(\w1[0][38] ), .Z(
        \SUBBYTES[0].a/n947 ) );
  XOR \SUBBYTES[0].a/U4731  ( .A(\SUBBYTES[0].a/w2468 ), .B(
        \SUBBYTES[0].a/w2475 ), .Z(\SUBBYTES[0].a/n948 ) );
  XOR \SUBBYTES[0].a/U4730  ( .A(\SUBBYTES[0].a/n950 ), .B(
        \SUBBYTES[0].a/n949 ), .Z(\SUBBYTES[0].a/n1534 ) );
  XOR \SUBBYTES[0].a/U4729  ( .A(\w1[0][33] ), .B(\SUBBYTES[0].a/n951 ), .Z(
        \SUBBYTES[0].a/n949 ) );
  XOR \SUBBYTES[0].a/U4728  ( .A(\SUBBYTES[0].a/w2493 ), .B(\w1[0][37] ), .Z(
        \SUBBYTES[0].a/n950 ) );
  XOR \SUBBYTES[0].a/U4727  ( .A(\SUBBYTES[0].a/w2469 ), .B(
        \SUBBYTES[0].a/w2476 ), .Z(\SUBBYTES[0].a/n951 ) );
  XOR \SUBBYTES[0].a/U4726  ( .A(\SUBBYTES[0].a/n1536 ), .B(
        \SUBBYTES[0].a/n1534 ), .Z(\SUBBYTES[0].a/w2499 ) );
  XOR \SUBBYTES[0].a/U4725  ( .A(\w1[0][37] ), .B(\SUBBYTES[0].a/n952 ), .Z(
        \SUBBYTES[0].a/n1537 ) );
  XOR \SUBBYTES[0].a/U4724  ( .A(\SUBBYTES[0].a/w2461 ), .B(
        \SUBBYTES[0].a/w2471 ), .Z(\SUBBYTES[0].a/n952 ) );
  XOR \SUBBYTES[0].a/U4723  ( .A(\SUBBYTES[0].a/n954 ), .B(
        \SUBBYTES[0].a/n953 ), .Z(\SUBBYTES[0].a/w2486 ) );
  XOR \SUBBYTES[0].a/U4722  ( .A(\SUBBYTES[0].a/n1537 ), .B(
        \SUBBYTES[0].a/n955 ), .Z(\SUBBYTES[0].a/n953 ) );
  XOR \SUBBYTES[0].a/U4721  ( .A(\w1[0][36] ), .B(\SUBBYTES[0].a/w2550 ), .Z(
        \SUBBYTES[0].a/n954 ) );
  XOR \SUBBYTES[0].a/U4720  ( .A(\SUBBYTES[0].a/w2463 ), .B(
        \SUBBYTES[0].a/w2468 ), .Z(\SUBBYTES[0].a/n955 ) );
  XOR \SUBBYTES[0].a/U4719  ( .A(\SUBBYTES[0].a/n957 ), .B(
        \SUBBYTES[0].a/n956 ), .Z(\SUBBYTES[0].a/n1535 ) );
  XOR \SUBBYTES[0].a/U4718  ( .A(\SUBBYTES[0].a/w2496 ), .B(\w1[0][39] ), .Z(
        \SUBBYTES[0].a/n956 ) );
  XOR \SUBBYTES[0].a/U4717  ( .A(\SUBBYTES[0].a/w2471 ), .B(
        \SUBBYTES[0].a/w2478 ), .Z(\SUBBYTES[0].a/n957 ) );
  XOR \SUBBYTES[0].a/U4716  ( .A(\SUBBYTES[0].a/n1534 ), .B(
        \SUBBYTES[0].a/n1535 ), .Z(\SUBBYTES[0].a/w2498 ) );
  XOR \SUBBYTES[0].a/U4715  ( .A(\w1[0][35] ), .B(\SUBBYTES[0].a/n958 ), .Z(
        \SUBBYTES[0].a/n1538 ) );
  XOR \SUBBYTES[0].a/U4714  ( .A(\SUBBYTES[0].a/w2460 ), .B(
        \SUBBYTES[0].a/w2463 ), .Z(\SUBBYTES[0].a/n958 ) );
  XOR \SUBBYTES[0].a/U4713  ( .A(\SUBBYTES[0].a/n960 ), .B(
        \SUBBYTES[0].a/n959 ), .Z(\SUBBYTES[0].a/w2487 ) );
  XOR \SUBBYTES[0].a/U4712  ( .A(\SUBBYTES[0].a/n1538 ), .B(
        \SUBBYTES[0].a/n961 ), .Z(\SUBBYTES[0].a/n959 ) );
  XOR \SUBBYTES[0].a/U4711  ( .A(\w1[0][38] ), .B(\SUBBYTES[0].a/w2529 ), .Z(
        \SUBBYTES[0].a/n960 ) );
  XOR \SUBBYTES[0].a/U4710  ( .A(\SUBBYTES[0].a/w2468 ), .B(
        \SUBBYTES[0].a/w2469 ), .Z(\SUBBYTES[0].a/n961 ) );
  XOR \SUBBYTES[0].a/U4709  ( .A(\SUBBYTES[0].a/n1536 ), .B(
        \SUBBYTES[0].a/n1535 ), .Z(\SUBBYTES[0].a/w2507 ) );
  XOR \SUBBYTES[0].a/U4708  ( .A(\SUBBYTES[0].a/n963 ), .B(
        \SUBBYTES[0].a/n962 ), .Z(\SUBBYTES[0].a/w2508 ) );
  XOR \SUBBYTES[0].a/U4707  ( .A(\w1[0][39] ), .B(\SUBBYTES[0].a/n1537 ), .Z(
        \SUBBYTES[0].a/n962 ) );
  XOR \SUBBYTES[0].a/U4706  ( .A(\SUBBYTES[0].a/w2460 ), .B(
        \SUBBYTES[0].a/w2469 ), .Z(\SUBBYTES[0].a/n963 ) );
  XOR \SUBBYTES[0].a/U4705  ( .A(\SUBBYTES[0].a/n965 ), .B(
        \SUBBYTES[0].a/n964 ), .Z(\SUBBYTES[0].a/w2484 ) );
  XOR \SUBBYTES[0].a/U4704  ( .A(\SUBBYTES[0].a/n967 ), .B(
        \SUBBYTES[0].a/n966 ), .Z(\SUBBYTES[0].a/n964 ) );
  XOR \SUBBYTES[0].a/U4703  ( .A(\w1[0][39] ), .B(\SUBBYTES[0].a/w2568 ), .Z(
        \SUBBYTES[0].a/n965 ) );
  XOR \SUBBYTES[0].a/U4702  ( .A(\SUBBYTES[0].a/w2475 ), .B(
        \SUBBYTES[0].a/w2478 ), .Z(\SUBBYTES[0].a/n966 ) );
  XOR \SUBBYTES[0].a/U4701  ( .A(\SUBBYTES[0].a/w2461 ), .B(
        \SUBBYTES[0].a/w2463 ), .Z(\SUBBYTES[0].a/n967 ) );
  XOR \SUBBYTES[0].a/U4700  ( .A(\SUBBYTES[0].a/n969 ), .B(
        \SUBBYTES[0].a/n968 ), .Z(\SUBBYTES[0].a/w2485 ) );
  XOR \SUBBYTES[0].a/U4699  ( .A(\SUBBYTES[0].a/n1538 ), .B(
        \SUBBYTES[0].a/n970 ), .Z(\SUBBYTES[0].a/n968 ) );
  XOR \SUBBYTES[0].a/U4698  ( .A(\w1[0][37] ), .B(\SUBBYTES[0].a/n1539 ), .Z(
        \SUBBYTES[0].a/n969 ) );
  XOR \SUBBYTES[0].a/U4697  ( .A(\SUBBYTES[0].a/w2475 ), .B(
        \SUBBYTES[0].a/w2476 ), .Z(\SUBBYTES[0].a/n970 ) );
  XOR \SUBBYTES[0].a/U4696  ( .A(\SUBBYTES[0].a/n972 ), .B(
        \SUBBYTES[0].a/n971 ), .Z(\SUBBYTES[0].a/w2501 ) );
  XOR \SUBBYTES[0].a/U4695  ( .A(\w1[0][33] ), .B(\SUBBYTES[0].a/n973 ), .Z(
        \SUBBYTES[0].a/n971 ) );
  XOR \SUBBYTES[0].a/U4694  ( .A(\SUBBYTES[0].a/w2476 ), .B(
        \SUBBYTES[0].a/w2478 ), .Z(\SUBBYTES[0].a/n972 ) );
  XOR \SUBBYTES[0].a/U4693  ( .A(\SUBBYTES[0].a/w2460 ), .B(
        \SUBBYTES[0].a/w2461 ), .Z(\SUBBYTES[0].a/n973 ) );
  XOR \SUBBYTES[0].a/U4692  ( .A(\w1[0][41] ), .B(\SUBBYTES[0].a/n974 ), .Z(
        \SUBBYTES[0].a/n1540 ) );
  XOR \SUBBYTES[0].a/U4691  ( .A(\w1[0][43] ), .B(\w1[0][42] ), .Z(
        \SUBBYTES[0].a/n974 ) );
  XOR \SUBBYTES[0].a/U4690  ( .A(\w1[0][46] ), .B(\SUBBYTES[0].a/n1540 ), .Z(
        \SUBBYTES[0].a/w2343 ) );
  XOR \SUBBYTES[0].a/U4689  ( .A(\w1[0][40] ), .B(\SUBBYTES[0].a/w2343 ), .Z(
        \SUBBYTES[0].a/w2230 ) );
  XOR \SUBBYTES[0].a/U4688  ( .A(\w1[0][40] ), .B(\SUBBYTES[0].a/n975 ), .Z(
        \SUBBYTES[0].a/w2231 ) );
  XOR \SUBBYTES[0].a/U4687  ( .A(\w1[0][46] ), .B(\w1[0][45] ), .Z(
        \SUBBYTES[0].a/n975 ) );
  XOR \SUBBYTES[0].a/U4686  ( .A(\w1[0][45] ), .B(\SUBBYTES[0].a/n1540 ), .Z(
        \SUBBYTES[0].a/w2361 ) );
  XOR \SUBBYTES[0].a/U4685  ( .A(\SUBBYTES[0].a/n977 ), .B(
        \SUBBYTES[0].a/n976 ), .Z(\SUBBYTES[0].a/w2354 ) );
  XOR \SUBBYTES[0].a/U4684  ( .A(\w1[0][43] ), .B(\w1[0][41] ), .Z(
        \SUBBYTES[0].a/n976 ) );
  XOR \SUBBYTES[0].a/U4683  ( .A(\w1[0][47] ), .B(\w1[0][44] ), .Z(
        \SUBBYTES[0].a/n977 ) );
  XOR \SUBBYTES[0].a/U4682  ( .A(\w1[0][40] ), .B(\SUBBYTES[0].a/w2354 ), .Z(
        \SUBBYTES[0].a/w2233 ) );
  XOR \SUBBYTES[0].a/U4681  ( .A(\SUBBYTES[0].a/n979 ), .B(
        \SUBBYTES[0].a/n978 ), .Z(\SUBBYTES[0].a/w2341 ) );
  XOR \SUBBYTES[0].a/U4680  ( .A(\SUBBYTES[0].a/w2302 ), .B(n1163), .Z(
        \SUBBYTES[0].a/n978 ) );
  XOR \SUBBYTES[0].a/U4679  ( .A(\SUBBYTES[0].a/w2295 ), .B(
        \SUBBYTES[0].a/w2298 ), .Z(\SUBBYTES[0].a/n979 ) );
  XOR \SUBBYTES[0].a/U4678  ( .A(\SUBBYTES[0].a/n981 ), .B(
        \SUBBYTES[0].a/n980 ), .Z(\SUBBYTES[0].a/w2342 ) );
  XOR \SUBBYTES[0].a/U4677  ( .A(\SUBBYTES[0].a/w2302 ), .B(
        \SUBBYTES[0].a/n110 ), .Z(\SUBBYTES[0].a/n980 ) );
  XOR \SUBBYTES[0].a/U4676  ( .A(\SUBBYTES[0].a/w2295 ), .B(
        \SUBBYTES[0].a/n109 ), .Z(\SUBBYTES[0].a/n981 ) );
  XOR \SUBBYTES[0].a/U4675  ( .A(\SUBBYTES[0].a/w2354 ), .B(
        \SUBBYTES[0].a/n982 ), .Z(\SUBBYTES[0].a/w2344 ) );
  XOR \SUBBYTES[0].a/U4674  ( .A(\w1[0][46] ), .B(\w1[0][45] ), .Z(
        \SUBBYTES[0].a/n982 ) );
  XOR \SUBBYTES[0].a/U4673  ( .A(\SUBBYTES[0].a/n984 ), .B(
        \SUBBYTES[0].a/n983 ), .Z(\SUBBYTES[0].a/w2345 ) );
  XOR \SUBBYTES[0].a/U4672  ( .A(\SUBBYTES[0].a/n110 ), .B(n1163), .Z(
        \SUBBYTES[0].a/n983 ) );
  XOR \SUBBYTES[0].a/U4671  ( .A(\SUBBYTES[0].a/n109 ), .B(
        \SUBBYTES[0].a/w2298 ), .Z(\SUBBYTES[0].a/n984 ) );
  XOR \SUBBYTES[0].a/U4670  ( .A(\w1[0][47] ), .B(\w1[0][42] ), .Z(
        \SUBBYTES[0].a/n1546 ) );
  XOR \SUBBYTES[0].a/U4669  ( .A(\SUBBYTES[0].a/n1546 ), .B(
        \SUBBYTES[0].a/n985 ), .Z(\SUBBYTES[0].a/w2346 ) );
  XOR \SUBBYTES[0].a/U4668  ( .A(\w1[0][45] ), .B(\w1[0][44] ), .Z(
        \SUBBYTES[0].a/n985 ) );
  XOR \SUBBYTES[0].a/U4667  ( .A(\w1[0][47] ), .B(\SUBBYTES[0].a/w2231 ), .Z(
        \SUBBYTES[0].a/w2234 ) );
  XOR \SUBBYTES[0].a/U4666  ( .A(\w1[0][41] ), .B(\SUBBYTES[0].a/w2231 ), .Z(
        \SUBBYTES[0].a/w2235 ) );
  XOR \SUBBYTES[0].a/U4665  ( .A(\w1[0][44] ), .B(\SUBBYTES[0].a/w2231 ), .Z(
        \SUBBYTES[0].a/w2236 ) );
  XOR \SUBBYTES[0].a/U4664  ( .A(\SUBBYTES[0].a/w2235 ), .B(
        \SUBBYTES[0].a/n1546 ), .Z(\SUBBYTES[0].a/w2237 ) );
  XOR \SUBBYTES[0].a/U4663  ( .A(\SUBBYTES[0].a/n1546 ), .B(
        \SUBBYTES[0].a/n986 ), .Z(\SUBBYTES[0].a/w2322 ) );
  XOR \SUBBYTES[0].a/U4662  ( .A(\w1[0][44] ), .B(\w1[0][41] ), .Z(
        \SUBBYTES[0].a/n986 ) );
  XOR \SUBBYTES[0].a/U4661  ( .A(\SUBBYTES[0].a/n988 ), .B(
        \SUBBYTES[0].a/n987 ), .Z(\SUBBYTES[0].a/n1543 ) );
  XOR \SUBBYTES[0].a/U4660  ( .A(\w1[0][44] ), .B(\SUBBYTES[0].a/n989 ), .Z(
        \SUBBYTES[0].a/n987 ) );
  XOR \SUBBYTES[0].a/U4659  ( .A(\SUBBYTES[0].a/w2287 ), .B(\w1[0][46] ), .Z(
        \SUBBYTES[0].a/n988 ) );
  XOR \SUBBYTES[0].a/U4658  ( .A(\SUBBYTES[0].a/w2261 ), .B(
        \SUBBYTES[0].a/w2268 ), .Z(\SUBBYTES[0].a/n989 ) );
  XOR \SUBBYTES[0].a/U4657  ( .A(\SUBBYTES[0].a/n991 ), .B(
        \SUBBYTES[0].a/n990 ), .Z(\SUBBYTES[0].a/n1541 ) );
  XOR \SUBBYTES[0].a/U4656  ( .A(\w1[0][41] ), .B(\SUBBYTES[0].a/n992 ), .Z(
        \SUBBYTES[0].a/n990 ) );
  XOR \SUBBYTES[0].a/U4655  ( .A(\SUBBYTES[0].a/w2286 ), .B(\w1[0][45] ), .Z(
        \SUBBYTES[0].a/n991 ) );
  XOR \SUBBYTES[0].a/U4654  ( .A(\SUBBYTES[0].a/w2262 ), .B(
        \SUBBYTES[0].a/w2269 ), .Z(\SUBBYTES[0].a/n992 ) );
  XOR \SUBBYTES[0].a/U4653  ( .A(\SUBBYTES[0].a/n1543 ), .B(
        \SUBBYTES[0].a/n1541 ), .Z(\SUBBYTES[0].a/w2292 ) );
  XOR \SUBBYTES[0].a/U4652  ( .A(\w1[0][45] ), .B(\SUBBYTES[0].a/n993 ), .Z(
        \SUBBYTES[0].a/n1544 ) );
  XOR \SUBBYTES[0].a/U4651  ( .A(\SUBBYTES[0].a/w2254 ), .B(
        \SUBBYTES[0].a/w2264 ), .Z(\SUBBYTES[0].a/n993 ) );
  XOR \SUBBYTES[0].a/U4650  ( .A(\SUBBYTES[0].a/n995 ), .B(
        \SUBBYTES[0].a/n994 ), .Z(\SUBBYTES[0].a/w2279 ) );
  XOR \SUBBYTES[0].a/U4649  ( .A(\SUBBYTES[0].a/n1544 ), .B(
        \SUBBYTES[0].a/n996 ), .Z(\SUBBYTES[0].a/n994 ) );
  XOR \SUBBYTES[0].a/U4648  ( .A(\w1[0][44] ), .B(\SUBBYTES[0].a/w2343 ), .Z(
        \SUBBYTES[0].a/n995 ) );
  XOR \SUBBYTES[0].a/U4647  ( .A(\SUBBYTES[0].a/w2256 ), .B(
        \SUBBYTES[0].a/w2261 ), .Z(\SUBBYTES[0].a/n996 ) );
  XOR \SUBBYTES[0].a/U4646  ( .A(\SUBBYTES[0].a/n998 ), .B(
        \SUBBYTES[0].a/n997 ), .Z(\SUBBYTES[0].a/n1542 ) );
  XOR \SUBBYTES[0].a/U4645  ( .A(\SUBBYTES[0].a/w2289 ), .B(\w1[0][47] ), .Z(
        \SUBBYTES[0].a/n997 ) );
  XOR \SUBBYTES[0].a/U4644  ( .A(\SUBBYTES[0].a/w2264 ), .B(
        \SUBBYTES[0].a/w2271 ), .Z(\SUBBYTES[0].a/n998 ) );
  XOR \SUBBYTES[0].a/U4643  ( .A(\SUBBYTES[0].a/n1541 ), .B(
        \SUBBYTES[0].a/n1542 ), .Z(\SUBBYTES[0].a/w2291 ) );
  XOR \SUBBYTES[0].a/U4642  ( .A(\w1[0][43] ), .B(\SUBBYTES[0].a/n999 ), .Z(
        \SUBBYTES[0].a/n1545 ) );
  XOR \SUBBYTES[0].a/U4641  ( .A(\SUBBYTES[0].a/w2253 ), .B(
        \SUBBYTES[0].a/w2256 ), .Z(\SUBBYTES[0].a/n999 ) );
  XOR \SUBBYTES[0].a/U4640  ( .A(\SUBBYTES[0].a/n1001 ), .B(
        \SUBBYTES[0].a/n1000 ), .Z(\SUBBYTES[0].a/w2280 ) );
  XOR \SUBBYTES[0].a/U4639  ( .A(\SUBBYTES[0].a/n1545 ), .B(
        \SUBBYTES[0].a/n1002 ), .Z(\SUBBYTES[0].a/n1000 ) );
  XOR \SUBBYTES[0].a/U4638  ( .A(\w1[0][46] ), .B(\SUBBYTES[0].a/w2322 ), .Z(
        \SUBBYTES[0].a/n1001 ) );
  XOR \SUBBYTES[0].a/U4637  ( .A(\SUBBYTES[0].a/w2261 ), .B(
        \SUBBYTES[0].a/w2262 ), .Z(\SUBBYTES[0].a/n1002 ) );
  XOR \SUBBYTES[0].a/U4636  ( .A(\SUBBYTES[0].a/n1543 ), .B(
        \SUBBYTES[0].a/n1542 ), .Z(\SUBBYTES[0].a/w2300 ) );
  XOR \SUBBYTES[0].a/U4635  ( .A(\SUBBYTES[0].a/n1004 ), .B(
        \SUBBYTES[0].a/n1003 ), .Z(\SUBBYTES[0].a/w2301 ) );
  XOR \SUBBYTES[0].a/U4634  ( .A(\w1[0][47] ), .B(\SUBBYTES[0].a/n1544 ), .Z(
        \SUBBYTES[0].a/n1003 ) );
  XOR \SUBBYTES[0].a/U4633  ( .A(\SUBBYTES[0].a/w2253 ), .B(
        \SUBBYTES[0].a/w2262 ), .Z(\SUBBYTES[0].a/n1004 ) );
  XOR \SUBBYTES[0].a/U4632  ( .A(\SUBBYTES[0].a/n1006 ), .B(
        \SUBBYTES[0].a/n1005 ), .Z(\SUBBYTES[0].a/w2277 ) );
  XOR \SUBBYTES[0].a/U4631  ( .A(\SUBBYTES[0].a/n1008 ), .B(
        \SUBBYTES[0].a/n1007 ), .Z(\SUBBYTES[0].a/n1005 ) );
  XOR \SUBBYTES[0].a/U4630  ( .A(\w1[0][47] ), .B(\SUBBYTES[0].a/w2361 ), .Z(
        \SUBBYTES[0].a/n1006 ) );
  XOR \SUBBYTES[0].a/U4629  ( .A(\SUBBYTES[0].a/w2268 ), .B(
        \SUBBYTES[0].a/w2271 ), .Z(\SUBBYTES[0].a/n1007 ) );
  XOR \SUBBYTES[0].a/U4628  ( .A(\SUBBYTES[0].a/w2254 ), .B(
        \SUBBYTES[0].a/w2256 ), .Z(\SUBBYTES[0].a/n1008 ) );
  XOR \SUBBYTES[0].a/U4627  ( .A(\SUBBYTES[0].a/n1010 ), .B(
        \SUBBYTES[0].a/n1009 ), .Z(\SUBBYTES[0].a/w2278 ) );
  XOR \SUBBYTES[0].a/U4626  ( .A(\SUBBYTES[0].a/n1545 ), .B(
        \SUBBYTES[0].a/n1011 ), .Z(\SUBBYTES[0].a/n1009 ) );
  XOR \SUBBYTES[0].a/U4625  ( .A(\w1[0][45] ), .B(\SUBBYTES[0].a/n1546 ), .Z(
        \SUBBYTES[0].a/n1010 ) );
  XOR \SUBBYTES[0].a/U4624  ( .A(\SUBBYTES[0].a/w2268 ), .B(
        \SUBBYTES[0].a/w2269 ), .Z(\SUBBYTES[0].a/n1011 ) );
  XOR \SUBBYTES[0].a/U4623  ( .A(\SUBBYTES[0].a/n1013 ), .B(
        \SUBBYTES[0].a/n1012 ), .Z(\SUBBYTES[0].a/w2294 ) );
  XOR \SUBBYTES[0].a/U4622  ( .A(\w1[0][41] ), .B(\SUBBYTES[0].a/n1014 ), .Z(
        \SUBBYTES[0].a/n1012 ) );
  XOR \SUBBYTES[0].a/U4621  ( .A(\SUBBYTES[0].a/w2269 ), .B(
        \SUBBYTES[0].a/w2271 ), .Z(\SUBBYTES[0].a/n1013 ) );
  XOR \SUBBYTES[0].a/U4620  ( .A(\SUBBYTES[0].a/w2253 ), .B(
        \SUBBYTES[0].a/w2254 ), .Z(\SUBBYTES[0].a/n1014 ) );
  XOR \SUBBYTES[0].a/U4619  ( .A(\w1[0][49] ), .B(\SUBBYTES[0].a/n1015 ), .Z(
        \SUBBYTES[0].a/n1547 ) );
  XOR \SUBBYTES[0].a/U4618  ( .A(\w1[0][51] ), .B(\w1[0][50] ), .Z(
        \SUBBYTES[0].a/n1015 ) );
  XOR \SUBBYTES[0].a/U4617  ( .A(\w1[0][54] ), .B(\SUBBYTES[0].a/n1547 ), .Z(
        \SUBBYTES[0].a/w2136 ) );
  XOR \SUBBYTES[0].a/U4616  ( .A(\w1[0][48] ), .B(\SUBBYTES[0].a/w2136 ), .Z(
        \SUBBYTES[0].a/w2023 ) );
  XOR \SUBBYTES[0].a/U4615  ( .A(\w1[0][48] ), .B(\SUBBYTES[0].a/n1016 ), .Z(
        \SUBBYTES[0].a/w2024 ) );
  XOR \SUBBYTES[0].a/U4614  ( .A(\w1[0][54] ), .B(\w1[0][53] ), .Z(
        \SUBBYTES[0].a/n1016 ) );
  XOR \SUBBYTES[0].a/U4613  ( .A(\w1[0][53] ), .B(\SUBBYTES[0].a/n1547 ), .Z(
        \SUBBYTES[0].a/w2154 ) );
  XOR \SUBBYTES[0].a/U4612  ( .A(\SUBBYTES[0].a/n1018 ), .B(
        \SUBBYTES[0].a/n1017 ), .Z(\SUBBYTES[0].a/w2147 ) );
  XOR \SUBBYTES[0].a/U4611  ( .A(\w1[0][51] ), .B(\w1[0][49] ), .Z(
        \SUBBYTES[0].a/n1017 ) );
  XOR \SUBBYTES[0].a/U4610  ( .A(\w1[0][55] ), .B(\w1[0][52] ), .Z(
        \SUBBYTES[0].a/n1018 ) );
  XOR \SUBBYTES[0].a/U4609  ( .A(\w1[0][48] ), .B(\SUBBYTES[0].a/w2147 ), .Z(
        \SUBBYTES[0].a/w2026 ) );
  XOR \SUBBYTES[0].a/U4608  ( .A(\SUBBYTES[0].a/n1020 ), .B(
        \SUBBYTES[0].a/n1019 ), .Z(\SUBBYTES[0].a/w2134 ) );
  XOR \SUBBYTES[0].a/U4607  ( .A(\SUBBYTES[0].a/w2095 ), .B(n1162), .Z(
        \SUBBYTES[0].a/n1019 ) );
  XOR \SUBBYTES[0].a/U4606  ( .A(\SUBBYTES[0].a/w2088 ), .B(
        \SUBBYTES[0].a/w2091 ), .Z(\SUBBYTES[0].a/n1020 ) );
  XOR \SUBBYTES[0].a/U4605  ( .A(\SUBBYTES[0].a/n1022 ), .B(
        \SUBBYTES[0].a/n1021 ), .Z(\SUBBYTES[0].a/w2135 ) );
  XOR \SUBBYTES[0].a/U4604  ( .A(\SUBBYTES[0].a/w2095 ), .B(
        \SUBBYTES[0].a/n100 ), .Z(\SUBBYTES[0].a/n1021 ) );
  XOR \SUBBYTES[0].a/U4603  ( .A(\SUBBYTES[0].a/w2088 ), .B(
        \SUBBYTES[0].a/n99 ), .Z(\SUBBYTES[0].a/n1022 ) );
  XOR \SUBBYTES[0].a/U4602  ( .A(\SUBBYTES[0].a/w2147 ), .B(
        \SUBBYTES[0].a/n1023 ), .Z(\SUBBYTES[0].a/w2137 ) );
  XOR \SUBBYTES[0].a/U4601  ( .A(\w1[0][54] ), .B(\w1[0][53] ), .Z(
        \SUBBYTES[0].a/n1023 ) );
  XOR \SUBBYTES[0].a/U4600  ( .A(\SUBBYTES[0].a/n1025 ), .B(
        \SUBBYTES[0].a/n1024 ), .Z(\SUBBYTES[0].a/w2138 ) );
  XOR \SUBBYTES[0].a/U4599  ( .A(\SUBBYTES[0].a/n100 ), .B(n1162), .Z(
        \SUBBYTES[0].a/n1024 ) );
  XOR \SUBBYTES[0].a/U4598  ( .A(\SUBBYTES[0].a/n99 ), .B(
        \SUBBYTES[0].a/w2091 ), .Z(\SUBBYTES[0].a/n1025 ) );
  XOR \SUBBYTES[0].a/U4597  ( .A(\w1[0][55] ), .B(\w1[0][50] ), .Z(
        \SUBBYTES[0].a/n1553 ) );
  XOR \SUBBYTES[0].a/U4596  ( .A(\SUBBYTES[0].a/n1553 ), .B(
        \SUBBYTES[0].a/n1026 ), .Z(\SUBBYTES[0].a/w2139 ) );
  XOR \SUBBYTES[0].a/U4595  ( .A(\w1[0][53] ), .B(\w1[0][52] ), .Z(
        \SUBBYTES[0].a/n1026 ) );
  XOR \SUBBYTES[0].a/U4594  ( .A(\w1[0][55] ), .B(\SUBBYTES[0].a/w2024 ), .Z(
        \SUBBYTES[0].a/w2027 ) );
  XOR \SUBBYTES[0].a/U4593  ( .A(\w1[0][49] ), .B(\SUBBYTES[0].a/w2024 ), .Z(
        \SUBBYTES[0].a/w2028 ) );
  XOR \SUBBYTES[0].a/U4592  ( .A(\w1[0][52] ), .B(\SUBBYTES[0].a/w2024 ), .Z(
        \SUBBYTES[0].a/w2029 ) );
  XOR \SUBBYTES[0].a/U4591  ( .A(\SUBBYTES[0].a/w2028 ), .B(
        \SUBBYTES[0].a/n1553 ), .Z(\SUBBYTES[0].a/w2030 ) );
  XOR \SUBBYTES[0].a/U4590  ( .A(\SUBBYTES[0].a/n1553 ), .B(
        \SUBBYTES[0].a/n1027 ), .Z(\SUBBYTES[0].a/w2115 ) );
  XOR \SUBBYTES[0].a/U4589  ( .A(\w1[0][52] ), .B(\w1[0][49] ), .Z(
        \SUBBYTES[0].a/n1027 ) );
  XOR \SUBBYTES[0].a/U4588  ( .A(\SUBBYTES[0].a/n1029 ), .B(
        \SUBBYTES[0].a/n1028 ), .Z(\SUBBYTES[0].a/n1550 ) );
  XOR \SUBBYTES[0].a/U4587  ( .A(\w1[0][52] ), .B(\SUBBYTES[0].a/n1030 ), .Z(
        \SUBBYTES[0].a/n1028 ) );
  XOR \SUBBYTES[0].a/U4586  ( .A(\SUBBYTES[0].a/w2080 ), .B(\w1[0][54] ), .Z(
        \SUBBYTES[0].a/n1029 ) );
  XOR \SUBBYTES[0].a/U4585  ( .A(\SUBBYTES[0].a/w2054 ), .B(
        \SUBBYTES[0].a/w2061 ), .Z(\SUBBYTES[0].a/n1030 ) );
  XOR \SUBBYTES[0].a/U4584  ( .A(\SUBBYTES[0].a/n1032 ), .B(
        \SUBBYTES[0].a/n1031 ), .Z(\SUBBYTES[0].a/n1548 ) );
  XOR \SUBBYTES[0].a/U4583  ( .A(\w1[0][49] ), .B(\SUBBYTES[0].a/n1033 ), .Z(
        \SUBBYTES[0].a/n1031 ) );
  XOR \SUBBYTES[0].a/U4582  ( .A(\SUBBYTES[0].a/w2079 ), .B(\w1[0][53] ), .Z(
        \SUBBYTES[0].a/n1032 ) );
  XOR \SUBBYTES[0].a/U4581  ( .A(\SUBBYTES[0].a/w2055 ), .B(
        \SUBBYTES[0].a/w2062 ), .Z(\SUBBYTES[0].a/n1033 ) );
  XOR \SUBBYTES[0].a/U4580  ( .A(\SUBBYTES[0].a/n1550 ), .B(
        \SUBBYTES[0].a/n1548 ), .Z(\SUBBYTES[0].a/w2085 ) );
  XOR \SUBBYTES[0].a/U4579  ( .A(\w1[0][53] ), .B(\SUBBYTES[0].a/n1034 ), .Z(
        \SUBBYTES[0].a/n1551 ) );
  XOR \SUBBYTES[0].a/U4578  ( .A(\SUBBYTES[0].a/w2047 ), .B(
        \SUBBYTES[0].a/w2057 ), .Z(\SUBBYTES[0].a/n1034 ) );
  XOR \SUBBYTES[0].a/U4577  ( .A(\SUBBYTES[0].a/n1036 ), .B(
        \SUBBYTES[0].a/n1035 ), .Z(\SUBBYTES[0].a/w2072 ) );
  XOR \SUBBYTES[0].a/U4576  ( .A(\SUBBYTES[0].a/n1551 ), .B(
        \SUBBYTES[0].a/n1037 ), .Z(\SUBBYTES[0].a/n1035 ) );
  XOR \SUBBYTES[0].a/U4575  ( .A(\w1[0][52] ), .B(\SUBBYTES[0].a/w2136 ), .Z(
        \SUBBYTES[0].a/n1036 ) );
  XOR \SUBBYTES[0].a/U4574  ( .A(\SUBBYTES[0].a/w2049 ), .B(
        \SUBBYTES[0].a/w2054 ), .Z(\SUBBYTES[0].a/n1037 ) );
  XOR \SUBBYTES[0].a/U4573  ( .A(\SUBBYTES[0].a/n1039 ), .B(
        \SUBBYTES[0].a/n1038 ), .Z(\SUBBYTES[0].a/n1549 ) );
  XOR \SUBBYTES[0].a/U4572  ( .A(\SUBBYTES[0].a/w2082 ), .B(\w1[0][55] ), .Z(
        \SUBBYTES[0].a/n1038 ) );
  XOR \SUBBYTES[0].a/U4571  ( .A(\SUBBYTES[0].a/w2057 ), .B(
        \SUBBYTES[0].a/w2064 ), .Z(\SUBBYTES[0].a/n1039 ) );
  XOR \SUBBYTES[0].a/U4570  ( .A(\SUBBYTES[0].a/n1548 ), .B(
        \SUBBYTES[0].a/n1549 ), .Z(\SUBBYTES[0].a/w2084 ) );
  XOR \SUBBYTES[0].a/U4569  ( .A(\w1[0][51] ), .B(\SUBBYTES[0].a/n1040 ), .Z(
        \SUBBYTES[0].a/n1552 ) );
  XOR \SUBBYTES[0].a/U4568  ( .A(\SUBBYTES[0].a/w2046 ), .B(
        \SUBBYTES[0].a/w2049 ), .Z(\SUBBYTES[0].a/n1040 ) );
  XOR \SUBBYTES[0].a/U4567  ( .A(\SUBBYTES[0].a/n1042 ), .B(
        \SUBBYTES[0].a/n1041 ), .Z(\SUBBYTES[0].a/w2073 ) );
  XOR \SUBBYTES[0].a/U4566  ( .A(\SUBBYTES[0].a/n1552 ), .B(
        \SUBBYTES[0].a/n1043 ), .Z(\SUBBYTES[0].a/n1041 ) );
  XOR \SUBBYTES[0].a/U4565  ( .A(\w1[0][54] ), .B(\SUBBYTES[0].a/w2115 ), .Z(
        \SUBBYTES[0].a/n1042 ) );
  XOR \SUBBYTES[0].a/U4564  ( .A(\SUBBYTES[0].a/w2054 ), .B(
        \SUBBYTES[0].a/w2055 ), .Z(\SUBBYTES[0].a/n1043 ) );
  XOR \SUBBYTES[0].a/U4563  ( .A(\SUBBYTES[0].a/n1550 ), .B(
        \SUBBYTES[0].a/n1549 ), .Z(\SUBBYTES[0].a/w2093 ) );
  XOR \SUBBYTES[0].a/U4562  ( .A(\SUBBYTES[0].a/n1045 ), .B(
        \SUBBYTES[0].a/n1044 ), .Z(\SUBBYTES[0].a/w2094 ) );
  XOR \SUBBYTES[0].a/U4561  ( .A(\w1[0][55] ), .B(\SUBBYTES[0].a/n1551 ), .Z(
        \SUBBYTES[0].a/n1044 ) );
  XOR \SUBBYTES[0].a/U4560  ( .A(\SUBBYTES[0].a/w2046 ), .B(
        \SUBBYTES[0].a/w2055 ), .Z(\SUBBYTES[0].a/n1045 ) );
  XOR \SUBBYTES[0].a/U4559  ( .A(\SUBBYTES[0].a/n1047 ), .B(
        \SUBBYTES[0].a/n1046 ), .Z(\SUBBYTES[0].a/w2070 ) );
  XOR \SUBBYTES[0].a/U4558  ( .A(\SUBBYTES[0].a/n1049 ), .B(
        \SUBBYTES[0].a/n1048 ), .Z(\SUBBYTES[0].a/n1046 ) );
  XOR \SUBBYTES[0].a/U4557  ( .A(\w1[0][55] ), .B(\SUBBYTES[0].a/w2154 ), .Z(
        \SUBBYTES[0].a/n1047 ) );
  XOR \SUBBYTES[0].a/U4556  ( .A(\SUBBYTES[0].a/w2061 ), .B(
        \SUBBYTES[0].a/w2064 ), .Z(\SUBBYTES[0].a/n1048 ) );
  XOR \SUBBYTES[0].a/U4555  ( .A(\SUBBYTES[0].a/w2047 ), .B(
        \SUBBYTES[0].a/w2049 ), .Z(\SUBBYTES[0].a/n1049 ) );
  XOR \SUBBYTES[0].a/U4554  ( .A(\SUBBYTES[0].a/n1051 ), .B(
        \SUBBYTES[0].a/n1050 ), .Z(\SUBBYTES[0].a/w2071 ) );
  XOR \SUBBYTES[0].a/U4553  ( .A(\SUBBYTES[0].a/n1552 ), .B(
        \SUBBYTES[0].a/n1052 ), .Z(\SUBBYTES[0].a/n1050 ) );
  XOR \SUBBYTES[0].a/U4552  ( .A(\w1[0][53] ), .B(\SUBBYTES[0].a/n1553 ), .Z(
        \SUBBYTES[0].a/n1051 ) );
  XOR \SUBBYTES[0].a/U4551  ( .A(\SUBBYTES[0].a/w2061 ), .B(
        \SUBBYTES[0].a/w2062 ), .Z(\SUBBYTES[0].a/n1052 ) );
  XOR \SUBBYTES[0].a/U4550  ( .A(\SUBBYTES[0].a/n1054 ), .B(
        \SUBBYTES[0].a/n1053 ), .Z(\SUBBYTES[0].a/w2087 ) );
  XOR \SUBBYTES[0].a/U4549  ( .A(\w1[0][49] ), .B(\SUBBYTES[0].a/n1055 ), .Z(
        \SUBBYTES[0].a/n1053 ) );
  XOR \SUBBYTES[0].a/U4548  ( .A(\SUBBYTES[0].a/w2062 ), .B(
        \SUBBYTES[0].a/w2064 ), .Z(\SUBBYTES[0].a/n1054 ) );
  XOR \SUBBYTES[0].a/U4547  ( .A(\SUBBYTES[0].a/w2046 ), .B(
        \SUBBYTES[0].a/w2047 ), .Z(\SUBBYTES[0].a/n1055 ) );
  XOR \SUBBYTES[0].a/U4546  ( .A(\w1[0][57] ), .B(\SUBBYTES[0].a/n1056 ), .Z(
        \SUBBYTES[0].a/n1554 ) );
  XOR \SUBBYTES[0].a/U4545  ( .A(\w1[0][59] ), .B(\w1[0][58] ), .Z(
        \SUBBYTES[0].a/n1056 ) );
  XOR \SUBBYTES[0].a/U4544  ( .A(\w1[0][62] ), .B(\SUBBYTES[0].a/n1554 ), .Z(
        \SUBBYTES[0].a/w1929 ) );
  XOR \SUBBYTES[0].a/U4543  ( .A(\w1[0][56] ), .B(\SUBBYTES[0].a/w1929 ), .Z(
        \SUBBYTES[0].a/w1816 ) );
  XOR \SUBBYTES[0].a/U4542  ( .A(\w1[0][56] ), .B(\SUBBYTES[0].a/n1057 ), .Z(
        \SUBBYTES[0].a/w1817 ) );
  XOR \SUBBYTES[0].a/U4541  ( .A(\w1[0][62] ), .B(\w1[0][61] ), .Z(
        \SUBBYTES[0].a/n1057 ) );
  XOR \SUBBYTES[0].a/U4540  ( .A(\w1[0][61] ), .B(\SUBBYTES[0].a/n1554 ), .Z(
        \SUBBYTES[0].a/w1947 ) );
  XOR \SUBBYTES[0].a/U4539  ( .A(\SUBBYTES[0].a/n1059 ), .B(
        \SUBBYTES[0].a/n1058 ), .Z(\SUBBYTES[0].a/w1940 ) );
  XOR \SUBBYTES[0].a/U4538  ( .A(\w1[0][59] ), .B(\w1[0][57] ), .Z(
        \SUBBYTES[0].a/n1058 ) );
  XOR \SUBBYTES[0].a/U4537  ( .A(\w1[0][63] ), .B(\w1[0][60] ), .Z(
        \SUBBYTES[0].a/n1059 ) );
  XOR \SUBBYTES[0].a/U4536  ( .A(\w1[0][56] ), .B(\SUBBYTES[0].a/w1940 ), .Z(
        \SUBBYTES[0].a/w1819 ) );
  XOR \SUBBYTES[0].a/U4535  ( .A(\SUBBYTES[0].a/n1061 ), .B(
        \SUBBYTES[0].a/n1060 ), .Z(\SUBBYTES[0].a/w1927 ) );
  XOR \SUBBYTES[0].a/U4534  ( .A(\SUBBYTES[0].a/w1888 ), .B(n1161), .Z(
        \SUBBYTES[0].a/n1060 ) );
  XOR \SUBBYTES[0].a/U4533  ( .A(\SUBBYTES[0].a/w1881 ), .B(
        \SUBBYTES[0].a/w1884 ), .Z(\SUBBYTES[0].a/n1061 ) );
  XOR \SUBBYTES[0].a/U4532  ( .A(\SUBBYTES[0].a/n1063 ), .B(
        \SUBBYTES[0].a/n1062 ), .Z(\SUBBYTES[0].a/w1928 ) );
  XOR \SUBBYTES[0].a/U4531  ( .A(\SUBBYTES[0].a/w1888 ), .B(
        \SUBBYTES[0].a/n90 ), .Z(\SUBBYTES[0].a/n1062 ) );
  XOR \SUBBYTES[0].a/U4530  ( .A(\SUBBYTES[0].a/w1881 ), .B(
        \SUBBYTES[0].a/n89 ), .Z(\SUBBYTES[0].a/n1063 ) );
  XOR \SUBBYTES[0].a/U4529  ( .A(\SUBBYTES[0].a/w1940 ), .B(
        \SUBBYTES[0].a/n1064 ), .Z(\SUBBYTES[0].a/w1930 ) );
  XOR \SUBBYTES[0].a/U4528  ( .A(\w1[0][62] ), .B(\w1[0][61] ), .Z(
        \SUBBYTES[0].a/n1064 ) );
  XOR \SUBBYTES[0].a/U4527  ( .A(\SUBBYTES[0].a/n1066 ), .B(
        \SUBBYTES[0].a/n1065 ), .Z(\SUBBYTES[0].a/w1931 ) );
  XOR \SUBBYTES[0].a/U4526  ( .A(\SUBBYTES[0].a/n90 ), .B(n1161), .Z(
        \SUBBYTES[0].a/n1065 ) );
  XOR \SUBBYTES[0].a/U4525  ( .A(\SUBBYTES[0].a/n89 ), .B(
        \SUBBYTES[0].a/w1884 ), .Z(\SUBBYTES[0].a/n1066 ) );
  XOR \SUBBYTES[0].a/U4524  ( .A(\w1[0][63] ), .B(\w1[0][58] ), .Z(
        \SUBBYTES[0].a/n1560 ) );
  XOR \SUBBYTES[0].a/U4523  ( .A(\SUBBYTES[0].a/n1560 ), .B(
        \SUBBYTES[0].a/n1067 ), .Z(\SUBBYTES[0].a/w1932 ) );
  XOR \SUBBYTES[0].a/U4522  ( .A(\w1[0][61] ), .B(\w1[0][60] ), .Z(
        \SUBBYTES[0].a/n1067 ) );
  XOR \SUBBYTES[0].a/U4521  ( .A(\w1[0][63] ), .B(\SUBBYTES[0].a/w1817 ), .Z(
        \SUBBYTES[0].a/w1820 ) );
  XOR \SUBBYTES[0].a/U4520  ( .A(\w1[0][57] ), .B(\SUBBYTES[0].a/w1817 ), .Z(
        \SUBBYTES[0].a/w1821 ) );
  XOR \SUBBYTES[0].a/U4519  ( .A(\w1[0][60] ), .B(\SUBBYTES[0].a/w1817 ), .Z(
        \SUBBYTES[0].a/w1822 ) );
  XOR \SUBBYTES[0].a/U4518  ( .A(\SUBBYTES[0].a/w1821 ), .B(
        \SUBBYTES[0].a/n1560 ), .Z(\SUBBYTES[0].a/w1823 ) );
  XOR \SUBBYTES[0].a/U4517  ( .A(\SUBBYTES[0].a/n1560 ), .B(
        \SUBBYTES[0].a/n1068 ), .Z(\SUBBYTES[0].a/w1908 ) );
  XOR \SUBBYTES[0].a/U4516  ( .A(\w1[0][60] ), .B(\w1[0][57] ), .Z(
        \SUBBYTES[0].a/n1068 ) );
  XOR \SUBBYTES[0].a/U4515  ( .A(\SUBBYTES[0].a/n1070 ), .B(
        \SUBBYTES[0].a/n1069 ), .Z(\SUBBYTES[0].a/n1557 ) );
  XOR \SUBBYTES[0].a/U4514  ( .A(\w1[0][60] ), .B(\SUBBYTES[0].a/n1071 ), .Z(
        \SUBBYTES[0].a/n1069 ) );
  XOR \SUBBYTES[0].a/U4513  ( .A(\SUBBYTES[0].a/w1873 ), .B(\w1[0][62] ), .Z(
        \SUBBYTES[0].a/n1070 ) );
  XOR \SUBBYTES[0].a/U4512  ( .A(\SUBBYTES[0].a/w1847 ), .B(
        \SUBBYTES[0].a/w1854 ), .Z(\SUBBYTES[0].a/n1071 ) );
  XOR \SUBBYTES[0].a/U4511  ( .A(\SUBBYTES[0].a/n1073 ), .B(
        \SUBBYTES[0].a/n1072 ), .Z(\SUBBYTES[0].a/n1555 ) );
  XOR \SUBBYTES[0].a/U4510  ( .A(\w1[0][57] ), .B(\SUBBYTES[0].a/n1074 ), .Z(
        \SUBBYTES[0].a/n1072 ) );
  XOR \SUBBYTES[0].a/U4509  ( .A(\SUBBYTES[0].a/w1872 ), .B(\w1[0][61] ), .Z(
        \SUBBYTES[0].a/n1073 ) );
  XOR \SUBBYTES[0].a/U4508  ( .A(\SUBBYTES[0].a/w1848 ), .B(
        \SUBBYTES[0].a/w1855 ), .Z(\SUBBYTES[0].a/n1074 ) );
  XOR \SUBBYTES[0].a/U4507  ( .A(\SUBBYTES[0].a/n1557 ), .B(
        \SUBBYTES[0].a/n1555 ), .Z(\SUBBYTES[0].a/w1878 ) );
  XOR \SUBBYTES[0].a/U4506  ( .A(\w1[0][61] ), .B(\SUBBYTES[0].a/n1075 ), .Z(
        \SUBBYTES[0].a/n1558 ) );
  XOR \SUBBYTES[0].a/U4505  ( .A(\SUBBYTES[0].a/w1840 ), .B(
        \SUBBYTES[0].a/w1850 ), .Z(\SUBBYTES[0].a/n1075 ) );
  XOR \SUBBYTES[0].a/U4504  ( .A(\SUBBYTES[0].a/n1077 ), .B(
        \SUBBYTES[0].a/n1076 ), .Z(\SUBBYTES[0].a/w1865 ) );
  XOR \SUBBYTES[0].a/U4503  ( .A(\SUBBYTES[0].a/n1558 ), .B(
        \SUBBYTES[0].a/n1078 ), .Z(\SUBBYTES[0].a/n1076 ) );
  XOR \SUBBYTES[0].a/U4502  ( .A(\w1[0][60] ), .B(\SUBBYTES[0].a/w1929 ), .Z(
        \SUBBYTES[0].a/n1077 ) );
  XOR \SUBBYTES[0].a/U4501  ( .A(\SUBBYTES[0].a/w1842 ), .B(
        \SUBBYTES[0].a/w1847 ), .Z(\SUBBYTES[0].a/n1078 ) );
  XOR \SUBBYTES[0].a/U4500  ( .A(\SUBBYTES[0].a/n1080 ), .B(
        \SUBBYTES[0].a/n1079 ), .Z(\SUBBYTES[0].a/n1556 ) );
  XOR \SUBBYTES[0].a/U4499  ( .A(\SUBBYTES[0].a/w1875 ), .B(\w1[0][63] ), .Z(
        \SUBBYTES[0].a/n1079 ) );
  XOR \SUBBYTES[0].a/U4498  ( .A(\SUBBYTES[0].a/w1850 ), .B(
        \SUBBYTES[0].a/w1857 ), .Z(\SUBBYTES[0].a/n1080 ) );
  XOR \SUBBYTES[0].a/U4497  ( .A(\SUBBYTES[0].a/n1555 ), .B(
        \SUBBYTES[0].a/n1556 ), .Z(\SUBBYTES[0].a/w1877 ) );
  XOR \SUBBYTES[0].a/U4496  ( .A(\w1[0][59] ), .B(\SUBBYTES[0].a/n1081 ), .Z(
        \SUBBYTES[0].a/n1559 ) );
  XOR \SUBBYTES[0].a/U4495  ( .A(\SUBBYTES[0].a/w1839 ), .B(
        \SUBBYTES[0].a/w1842 ), .Z(\SUBBYTES[0].a/n1081 ) );
  XOR \SUBBYTES[0].a/U4494  ( .A(\SUBBYTES[0].a/n1083 ), .B(
        \SUBBYTES[0].a/n1082 ), .Z(\SUBBYTES[0].a/w1866 ) );
  XOR \SUBBYTES[0].a/U4493  ( .A(\SUBBYTES[0].a/n1559 ), .B(
        \SUBBYTES[0].a/n1084 ), .Z(\SUBBYTES[0].a/n1082 ) );
  XOR \SUBBYTES[0].a/U4492  ( .A(\w1[0][62] ), .B(\SUBBYTES[0].a/w1908 ), .Z(
        \SUBBYTES[0].a/n1083 ) );
  XOR \SUBBYTES[0].a/U4491  ( .A(\SUBBYTES[0].a/w1847 ), .B(
        \SUBBYTES[0].a/w1848 ), .Z(\SUBBYTES[0].a/n1084 ) );
  XOR \SUBBYTES[0].a/U4490  ( .A(\SUBBYTES[0].a/n1557 ), .B(
        \SUBBYTES[0].a/n1556 ), .Z(\SUBBYTES[0].a/w1886 ) );
  XOR \SUBBYTES[0].a/U4489  ( .A(\SUBBYTES[0].a/n1086 ), .B(
        \SUBBYTES[0].a/n1085 ), .Z(\SUBBYTES[0].a/w1887 ) );
  XOR \SUBBYTES[0].a/U4488  ( .A(\w1[0][63] ), .B(\SUBBYTES[0].a/n1558 ), .Z(
        \SUBBYTES[0].a/n1085 ) );
  XOR \SUBBYTES[0].a/U4487  ( .A(\SUBBYTES[0].a/w1839 ), .B(
        \SUBBYTES[0].a/w1848 ), .Z(\SUBBYTES[0].a/n1086 ) );
  XOR \SUBBYTES[0].a/U4486  ( .A(\SUBBYTES[0].a/n1088 ), .B(
        \SUBBYTES[0].a/n1087 ), .Z(\SUBBYTES[0].a/w1863 ) );
  XOR \SUBBYTES[0].a/U4485  ( .A(\SUBBYTES[0].a/n1090 ), .B(
        \SUBBYTES[0].a/n1089 ), .Z(\SUBBYTES[0].a/n1087 ) );
  XOR \SUBBYTES[0].a/U4484  ( .A(\w1[0][63] ), .B(\SUBBYTES[0].a/w1947 ), .Z(
        \SUBBYTES[0].a/n1088 ) );
  XOR \SUBBYTES[0].a/U4483  ( .A(\SUBBYTES[0].a/w1854 ), .B(
        \SUBBYTES[0].a/w1857 ), .Z(\SUBBYTES[0].a/n1089 ) );
  XOR \SUBBYTES[0].a/U4482  ( .A(\SUBBYTES[0].a/w1840 ), .B(
        \SUBBYTES[0].a/w1842 ), .Z(\SUBBYTES[0].a/n1090 ) );
  XOR \SUBBYTES[0].a/U4481  ( .A(\SUBBYTES[0].a/n1092 ), .B(
        \SUBBYTES[0].a/n1091 ), .Z(\SUBBYTES[0].a/w1864 ) );
  XOR \SUBBYTES[0].a/U4480  ( .A(\SUBBYTES[0].a/n1559 ), .B(
        \SUBBYTES[0].a/n1093 ), .Z(\SUBBYTES[0].a/n1091 ) );
  XOR \SUBBYTES[0].a/U4479  ( .A(\w1[0][61] ), .B(\SUBBYTES[0].a/n1560 ), .Z(
        \SUBBYTES[0].a/n1092 ) );
  XOR \SUBBYTES[0].a/U4478  ( .A(\SUBBYTES[0].a/w1854 ), .B(
        \SUBBYTES[0].a/w1855 ), .Z(\SUBBYTES[0].a/n1093 ) );
  XOR \SUBBYTES[0].a/U4477  ( .A(\SUBBYTES[0].a/n1095 ), .B(
        \SUBBYTES[0].a/n1094 ), .Z(\SUBBYTES[0].a/w1880 ) );
  XOR \SUBBYTES[0].a/U4476  ( .A(\w1[0][57] ), .B(\SUBBYTES[0].a/n1096 ), .Z(
        \SUBBYTES[0].a/n1094 ) );
  XOR \SUBBYTES[0].a/U4475  ( .A(\SUBBYTES[0].a/w1855 ), .B(
        \SUBBYTES[0].a/w1857 ), .Z(\SUBBYTES[0].a/n1095 ) );
  XOR \SUBBYTES[0].a/U4474  ( .A(\SUBBYTES[0].a/w1839 ), .B(
        \SUBBYTES[0].a/w1840 ), .Z(\SUBBYTES[0].a/n1096 ) );
  XOR \SUBBYTES[0].a/U4473  ( .A(\w1[0][65] ), .B(\SUBBYTES[0].a/n1097 ), .Z(
        \SUBBYTES[0].a/n1561 ) );
  XOR \SUBBYTES[0].a/U4472  ( .A(\w1[0][67] ), .B(\w1[0][66] ), .Z(
        \SUBBYTES[0].a/n1097 ) );
  XOR \SUBBYTES[0].a/U4471  ( .A(\w1[0][70] ), .B(\SUBBYTES[0].a/n1561 ), .Z(
        \SUBBYTES[0].a/w1722 ) );
  XOR \SUBBYTES[0].a/U4470  ( .A(\w1[0][64] ), .B(\SUBBYTES[0].a/w1722 ), .Z(
        \SUBBYTES[0].a/w1609 ) );
  XOR \SUBBYTES[0].a/U4469  ( .A(\w1[0][64] ), .B(\SUBBYTES[0].a/n1098 ), .Z(
        \SUBBYTES[0].a/w1610 ) );
  XOR \SUBBYTES[0].a/U4468  ( .A(\w1[0][70] ), .B(\w1[0][69] ), .Z(
        \SUBBYTES[0].a/n1098 ) );
  XOR \SUBBYTES[0].a/U4467  ( .A(\w1[0][69] ), .B(\SUBBYTES[0].a/n1561 ), .Z(
        \SUBBYTES[0].a/w1740 ) );
  XOR \SUBBYTES[0].a/U4466  ( .A(\SUBBYTES[0].a/n1100 ), .B(
        \SUBBYTES[0].a/n1099 ), .Z(\SUBBYTES[0].a/w1733 ) );
  XOR \SUBBYTES[0].a/U4465  ( .A(\w1[0][67] ), .B(\w1[0][65] ), .Z(
        \SUBBYTES[0].a/n1099 ) );
  XOR \SUBBYTES[0].a/U4464  ( .A(\w1[0][71] ), .B(\w1[0][68] ), .Z(
        \SUBBYTES[0].a/n1100 ) );
  XOR \SUBBYTES[0].a/U4463  ( .A(\w1[0][64] ), .B(\SUBBYTES[0].a/w1733 ), .Z(
        \SUBBYTES[0].a/w1612 ) );
  XOR \SUBBYTES[0].a/U4462  ( .A(\SUBBYTES[0].a/n1102 ), .B(
        \SUBBYTES[0].a/n1101 ), .Z(\SUBBYTES[0].a/w1720 ) );
  XOR \SUBBYTES[0].a/U4461  ( .A(\SUBBYTES[0].a/w1681 ), .B(n1160), .Z(
        \SUBBYTES[0].a/n1101 ) );
  XOR \SUBBYTES[0].a/U4460  ( .A(\SUBBYTES[0].a/w1674 ), .B(
        \SUBBYTES[0].a/w1677 ), .Z(\SUBBYTES[0].a/n1102 ) );
  XOR \SUBBYTES[0].a/U4459  ( .A(\SUBBYTES[0].a/n1104 ), .B(
        \SUBBYTES[0].a/n1103 ), .Z(\SUBBYTES[0].a/w1721 ) );
  XOR \SUBBYTES[0].a/U4458  ( .A(\SUBBYTES[0].a/w1681 ), .B(
        \SUBBYTES[0].a/n80 ), .Z(\SUBBYTES[0].a/n1103 ) );
  XOR \SUBBYTES[0].a/U4457  ( .A(\SUBBYTES[0].a/w1674 ), .B(
        \SUBBYTES[0].a/n79 ), .Z(\SUBBYTES[0].a/n1104 ) );
  XOR \SUBBYTES[0].a/U4456  ( .A(\SUBBYTES[0].a/w1733 ), .B(
        \SUBBYTES[0].a/n1105 ), .Z(\SUBBYTES[0].a/w1723 ) );
  XOR \SUBBYTES[0].a/U4455  ( .A(\w1[0][70] ), .B(\w1[0][69] ), .Z(
        \SUBBYTES[0].a/n1105 ) );
  XOR \SUBBYTES[0].a/U4454  ( .A(\SUBBYTES[0].a/n1107 ), .B(
        \SUBBYTES[0].a/n1106 ), .Z(\SUBBYTES[0].a/w1724 ) );
  XOR \SUBBYTES[0].a/U4453  ( .A(\SUBBYTES[0].a/n80 ), .B(n1160), .Z(
        \SUBBYTES[0].a/n1106 ) );
  XOR \SUBBYTES[0].a/U4452  ( .A(\SUBBYTES[0].a/n79 ), .B(
        \SUBBYTES[0].a/w1677 ), .Z(\SUBBYTES[0].a/n1107 ) );
  XOR \SUBBYTES[0].a/U4451  ( .A(\w1[0][71] ), .B(\w1[0][66] ), .Z(
        \SUBBYTES[0].a/n1567 ) );
  XOR \SUBBYTES[0].a/U4450  ( .A(\SUBBYTES[0].a/n1567 ), .B(
        \SUBBYTES[0].a/n1108 ), .Z(\SUBBYTES[0].a/w1725 ) );
  XOR \SUBBYTES[0].a/U4449  ( .A(\w1[0][69] ), .B(\w1[0][68] ), .Z(
        \SUBBYTES[0].a/n1108 ) );
  XOR \SUBBYTES[0].a/U4448  ( .A(\w1[0][71] ), .B(\SUBBYTES[0].a/w1610 ), .Z(
        \SUBBYTES[0].a/w1613 ) );
  XOR \SUBBYTES[0].a/U4447  ( .A(\w1[0][65] ), .B(\SUBBYTES[0].a/w1610 ), .Z(
        \SUBBYTES[0].a/w1614 ) );
  XOR \SUBBYTES[0].a/U4446  ( .A(\w1[0][68] ), .B(\SUBBYTES[0].a/w1610 ), .Z(
        \SUBBYTES[0].a/w1615 ) );
  XOR \SUBBYTES[0].a/U4445  ( .A(\SUBBYTES[0].a/w1614 ), .B(
        \SUBBYTES[0].a/n1567 ), .Z(\SUBBYTES[0].a/w1616 ) );
  XOR \SUBBYTES[0].a/U4444  ( .A(\SUBBYTES[0].a/n1567 ), .B(
        \SUBBYTES[0].a/n1109 ), .Z(\SUBBYTES[0].a/w1701 ) );
  XOR \SUBBYTES[0].a/U4443  ( .A(\w1[0][68] ), .B(\w1[0][65] ), .Z(
        \SUBBYTES[0].a/n1109 ) );
  XOR \SUBBYTES[0].a/U4442  ( .A(\SUBBYTES[0].a/n1111 ), .B(
        \SUBBYTES[0].a/n1110 ), .Z(\SUBBYTES[0].a/n1564 ) );
  XOR \SUBBYTES[0].a/U4441  ( .A(\w1[0][68] ), .B(\SUBBYTES[0].a/n1112 ), .Z(
        \SUBBYTES[0].a/n1110 ) );
  XOR \SUBBYTES[0].a/U4440  ( .A(\SUBBYTES[0].a/w1666 ), .B(\w1[0][70] ), .Z(
        \SUBBYTES[0].a/n1111 ) );
  XOR \SUBBYTES[0].a/U4439  ( .A(\SUBBYTES[0].a/w1640 ), .B(
        \SUBBYTES[0].a/w1647 ), .Z(\SUBBYTES[0].a/n1112 ) );
  XOR \SUBBYTES[0].a/U4438  ( .A(\SUBBYTES[0].a/n1114 ), .B(
        \SUBBYTES[0].a/n1113 ), .Z(\SUBBYTES[0].a/n1562 ) );
  XOR \SUBBYTES[0].a/U4437  ( .A(\w1[0][65] ), .B(\SUBBYTES[0].a/n1115 ), .Z(
        \SUBBYTES[0].a/n1113 ) );
  XOR \SUBBYTES[0].a/U4436  ( .A(\SUBBYTES[0].a/w1665 ), .B(\w1[0][69] ), .Z(
        \SUBBYTES[0].a/n1114 ) );
  XOR \SUBBYTES[0].a/U4435  ( .A(\SUBBYTES[0].a/w1641 ), .B(
        \SUBBYTES[0].a/w1648 ), .Z(\SUBBYTES[0].a/n1115 ) );
  XOR \SUBBYTES[0].a/U4434  ( .A(\SUBBYTES[0].a/n1564 ), .B(
        \SUBBYTES[0].a/n1562 ), .Z(\SUBBYTES[0].a/w1671 ) );
  XOR \SUBBYTES[0].a/U4433  ( .A(\w1[0][69] ), .B(\SUBBYTES[0].a/n1116 ), .Z(
        \SUBBYTES[0].a/n1565 ) );
  XOR \SUBBYTES[0].a/U4432  ( .A(\SUBBYTES[0].a/w1633 ), .B(
        \SUBBYTES[0].a/w1643 ), .Z(\SUBBYTES[0].a/n1116 ) );
  XOR \SUBBYTES[0].a/U4431  ( .A(\SUBBYTES[0].a/n1118 ), .B(
        \SUBBYTES[0].a/n1117 ), .Z(\SUBBYTES[0].a/w1658 ) );
  XOR \SUBBYTES[0].a/U4430  ( .A(\SUBBYTES[0].a/n1565 ), .B(
        \SUBBYTES[0].a/n1119 ), .Z(\SUBBYTES[0].a/n1117 ) );
  XOR \SUBBYTES[0].a/U4429  ( .A(\w1[0][68] ), .B(\SUBBYTES[0].a/w1722 ), .Z(
        \SUBBYTES[0].a/n1118 ) );
  XOR \SUBBYTES[0].a/U4428  ( .A(\SUBBYTES[0].a/w1635 ), .B(
        \SUBBYTES[0].a/w1640 ), .Z(\SUBBYTES[0].a/n1119 ) );
  XOR \SUBBYTES[0].a/U4427  ( .A(\SUBBYTES[0].a/n1121 ), .B(
        \SUBBYTES[0].a/n1120 ), .Z(\SUBBYTES[0].a/n1563 ) );
  XOR \SUBBYTES[0].a/U4426  ( .A(\SUBBYTES[0].a/w1668 ), .B(\w1[0][71] ), .Z(
        \SUBBYTES[0].a/n1120 ) );
  XOR \SUBBYTES[0].a/U4425  ( .A(\SUBBYTES[0].a/w1643 ), .B(
        \SUBBYTES[0].a/w1650 ), .Z(\SUBBYTES[0].a/n1121 ) );
  XOR \SUBBYTES[0].a/U4424  ( .A(\SUBBYTES[0].a/n1562 ), .B(
        \SUBBYTES[0].a/n1563 ), .Z(\SUBBYTES[0].a/w1670 ) );
  XOR \SUBBYTES[0].a/U4423  ( .A(\w1[0][67] ), .B(\SUBBYTES[0].a/n1122 ), .Z(
        \SUBBYTES[0].a/n1566 ) );
  XOR \SUBBYTES[0].a/U4422  ( .A(\SUBBYTES[0].a/w1632 ), .B(
        \SUBBYTES[0].a/w1635 ), .Z(\SUBBYTES[0].a/n1122 ) );
  XOR \SUBBYTES[0].a/U4421  ( .A(\SUBBYTES[0].a/n1124 ), .B(
        \SUBBYTES[0].a/n1123 ), .Z(\SUBBYTES[0].a/w1659 ) );
  XOR \SUBBYTES[0].a/U4420  ( .A(\SUBBYTES[0].a/n1566 ), .B(
        \SUBBYTES[0].a/n1125 ), .Z(\SUBBYTES[0].a/n1123 ) );
  XOR \SUBBYTES[0].a/U4419  ( .A(\w1[0][70] ), .B(\SUBBYTES[0].a/w1701 ), .Z(
        \SUBBYTES[0].a/n1124 ) );
  XOR \SUBBYTES[0].a/U4418  ( .A(\SUBBYTES[0].a/w1640 ), .B(
        \SUBBYTES[0].a/w1641 ), .Z(\SUBBYTES[0].a/n1125 ) );
  XOR \SUBBYTES[0].a/U4417  ( .A(\SUBBYTES[0].a/n1564 ), .B(
        \SUBBYTES[0].a/n1563 ), .Z(\SUBBYTES[0].a/w1679 ) );
  XOR \SUBBYTES[0].a/U4416  ( .A(\SUBBYTES[0].a/n1127 ), .B(
        \SUBBYTES[0].a/n1126 ), .Z(\SUBBYTES[0].a/w1680 ) );
  XOR \SUBBYTES[0].a/U4415  ( .A(\w1[0][71] ), .B(\SUBBYTES[0].a/n1565 ), .Z(
        \SUBBYTES[0].a/n1126 ) );
  XOR \SUBBYTES[0].a/U4414  ( .A(\SUBBYTES[0].a/w1632 ), .B(
        \SUBBYTES[0].a/w1641 ), .Z(\SUBBYTES[0].a/n1127 ) );
  XOR \SUBBYTES[0].a/U4413  ( .A(\SUBBYTES[0].a/n1129 ), .B(
        \SUBBYTES[0].a/n1128 ), .Z(\SUBBYTES[0].a/w1656 ) );
  XOR \SUBBYTES[0].a/U4412  ( .A(\SUBBYTES[0].a/n1131 ), .B(
        \SUBBYTES[0].a/n1130 ), .Z(\SUBBYTES[0].a/n1128 ) );
  XOR \SUBBYTES[0].a/U4411  ( .A(\w1[0][71] ), .B(\SUBBYTES[0].a/w1740 ), .Z(
        \SUBBYTES[0].a/n1129 ) );
  XOR \SUBBYTES[0].a/U4410  ( .A(\SUBBYTES[0].a/w1647 ), .B(
        \SUBBYTES[0].a/w1650 ), .Z(\SUBBYTES[0].a/n1130 ) );
  XOR \SUBBYTES[0].a/U4409  ( .A(\SUBBYTES[0].a/w1633 ), .B(
        \SUBBYTES[0].a/w1635 ), .Z(\SUBBYTES[0].a/n1131 ) );
  XOR \SUBBYTES[0].a/U4408  ( .A(\SUBBYTES[0].a/n1133 ), .B(
        \SUBBYTES[0].a/n1132 ), .Z(\SUBBYTES[0].a/w1657 ) );
  XOR \SUBBYTES[0].a/U4407  ( .A(\SUBBYTES[0].a/n1566 ), .B(
        \SUBBYTES[0].a/n1134 ), .Z(\SUBBYTES[0].a/n1132 ) );
  XOR \SUBBYTES[0].a/U4406  ( .A(\w1[0][69] ), .B(\SUBBYTES[0].a/n1567 ), .Z(
        \SUBBYTES[0].a/n1133 ) );
  XOR \SUBBYTES[0].a/U4405  ( .A(\SUBBYTES[0].a/w1647 ), .B(
        \SUBBYTES[0].a/w1648 ), .Z(\SUBBYTES[0].a/n1134 ) );
  XOR \SUBBYTES[0].a/U4404  ( .A(\SUBBYTES[0].a/n1136 ), .B(
        \SUBBYTES[0].a/n1135 ), .Z(\SUBBYTES[0].a/w1673 ) );
  XOR \SUBBYTES[0].a/U4403  ( .A(\w1[0][65] ), .B(\SUBBYTES[0].a/n1137 ), .Z(
        \SUBBYTES[0].a/n1135 ) );
  XOR \SUBBYTES[0].a/U4402  ( .A(\SUBBYTES[0].a/w1648 ), .B(
        \SUBBYTES[0].a/w1650 ), .Z(\SUBBYTES[0].a/n1136 ) );
  XOR \SUBBYTES[0].a/U4401  ( .A(\SUBBYTES[0].a/w1632 ), .B(
        \SUBBYTES[0].a/w1633 ), .Z(\SUBBYTES[0].a/n1137 ) );
  XOR \SUBBYTES[0].a/U4400  ( .A(\w1[0][73] ), .B(\SUBBYTES[0].a/n1138 ), .Z(
        \SUBBYTES[0].a/n1568 ) );
  XOR \SUBBYTES[0].a/U4399  ( .A(\w1[0][75] ), .B(\w1[0][74] ), .Z(
        \SUBBYTES[0].a/n1138 ) );
  XOR \SUBBYTES[0].a/U4398  ( .A(\w1[0][78] ), .B(\SUBBYTES[0].a/n1568 ), .Z(
        \SUBBYTES[0].a/w1515 ) );
  XOR \SUBBYTES[0].a/U4397  ( .A(\w1[0][72] ), .B(\SUBBYTES[0].a/w1515 ), .Z(
        \SUBBYTES[0].a/w1402 ) );
  XOR \SUBBYTES[0].a/U4396  ( .A(\w1[0][72] ), .B(\SUBBYTES[0].a/n1139 ), .Z(
        \SUBBYTES[0].a/w1403 ) );
  XOR \SUBBYTES[0].a/U4395  ( .A(\w1[0][78] ), .B(\w1[0][77] ), .Z(
        \SUBBYTES[0].a/n1139 ) );
  XOR \SUBBYTES[0].a/U4394  ( .A(\w1[0][77] ), .B(\SUBBYTES[0].a/n1568 ), .Z(
        \SUBBYTES[0].a/w1533 ) );
  XOR \SUBBYTES[0].a/U4393  ( .A(\SUBBYTES[0].a/n1141 ), .B(
        \SUBBYTES[0].a/n1140 ), .Z(\SUBBYTES[0].a/w1526 ) );
  XOR \SUBBYTES[0].a/U4392  ( .A(\w1[0][75] ), .B(\w1[0][73] ), .Z(
        \SUBBYTES[0].a/n1140 ) );
  XOR \SUBBYTES[0].a/U4391  ( .A(\w1[0][79] ), .B(\w1[0][76] ), .Z(
        \SUBBYTES[0].a/n1141 ) );
  XOR \SUBBYTES[0].a/U4390  ( .A(\w1[0][72] ), .B(\SUBBYTES[0].a/w1526 ), .Z(
        \SUBBYTES[0].a/w1405 ) );
  XOR \SUBBYTES[0].a/U4389  ( .A(\SUBBYTES[0].a/n1143 ), .B(
        \SUBBYTES[0].a/n1142 ), .Z(\SUBBYTES[0].a/w1513 ) );
  XOR \SUBBYTES[0].a/U4388  ( .A(\SUBBYTES[0].a/w1474 ), .B(n1159), .Z(
        \SUBBYTES[0].a/n1142 ) );
  XOR \SUBBYTES[0].a/U4387  ( .A(\SUBBYTES[0].a/w1467 ), .B(
        \SUBBYTES[0].a/w1470 ), .Z(\SUBBYTES[0].a/n1143 ) );
  XOR \SUBBYTES[0].a/U4386  ( .A(\SUBBYTES[0].a/n1145 ), .B(
        \SUBBYTES[0].a/n1144 ), .Z(\SUBBYTES[0].a/w1514 ) );
  XOR \SUBBYTES[0].a/U4385  ( .A(\SUBBYTES[0].a/w1474 ), .B(
        \SUBBYTES[0].a/n70 ), .Z(\SUBBYTES[0].a/n1144 ) );
  XOR \SUBBYTES[0].a/U4384  ( .A(\SUBBYTES[0].a/w1467 ), .B(
        \SUBBYTES[0].a/n69 ), .Z(\SUBBYTES[0].a/n1145 ) );
  XOR \SUBBYTES[0].a/U4383  ( .A(\SUBBYTES[0].a/w1526 ), .B(
        \SUBBYTES[0].a/n1146 ), .Z(\SUBBYTES[0].a/w1516 ) );
  XOR \SUBBYTES[0].a/U4382  ( .A(\w1[0][78] ), .B(\w1[0][77] ), .Z(
        \SUBBYTES[0].a/n1146 ) );
  XOR \SUBBYTES[0].a/U4381  ( .A(\SUBBYTES[0].a/n1148 ), .B(
        \SUBBYTES[0].a/n1147 ), .Z(\SUBBYTES[0].a/w1517 ) );
  XOR \SUBBYTES[0].a/U4380  ( .A(\SUBBYTES[0].a/n70 ), .B(n1159), .Z(
        \SUBBYTES[0].a/n1147 ) );
  XOR \SUBBYTES[0].a/U4379  ( .A(\SUBBYTES[0].a/n69 ), .B(
        \SUBBYTES[0].a/w1470 ), .Z(\SUBBYTES[0].a/n1148 ) );
  XOR \SUBBYTES[0].a/U4378  ( .A(\w1[0][79] ), .B(\w1[0][74] ), .Z(
        \SUBBYTES[0].a/n1574 ) );
  XOR \SUBBYTES[0].a/U4377  ( .A(\SUBBYTES[0].a/n1574 ), .B(
        \SUBBYTES[0].a/n1149 ), .Z(\SUBBYTES[0].a/w1518 ) );
  XOR \SUBBYTES[0].a/U4376  ( .A(\w1[0][77] ), .B(\w1[0][76] ), .Z(
        \SUBBYTES[0].a/n1149 ) );
  XOR \SUBBYTES[0].a/U4375  ( .A(\w1[0][79] ), .B(\SUBBYTES[0].a/w1403 ), .Z(
        \SUBBYTES[0].a/w1406 ) );
  XOR \SUBBYTES[0].a/U4374  ( .A(\w1[0][73] ), .B(\SUBBYTES[0].a/w1403 ), .Z(
        \SUBBYTES[0].a/w1407 ) );
  XOR \SUBBYTES[0].a/U4373  ( .A(\w1[0][76] ), .B(\SUBBYTES[0].a/w1403 ), .Z(
        \SUBBYTES[0].a/w1408 ) );
  XOR \SUBBYTES[0].a/U4372  ( .A(\SUBBYTES[0].a/w1407 ), .B(
        \SUBBYTES[0].a/n1574 ), .Z(\SUBBYTES[0].a/w1409 ) );
  XOR \SUBBYTES[0].a/U4371  ( .A(\SUBBYTES[0].a/n1574 ), .B(
        \SUBBYTES[0].a/n1150 ), .Z(\SUBBYTES[0].a/w1494 ) );
  XOR \SUBBYTES[0].a/U4370  ( .A(\w1[0][76] ), .B(\w1[0][73] ), .Z(
        \SUBBYTES[0].a/n1150 ) );
  XOR \SUBBYTES[0].a/U4369  ( .A(\SUBBYTES[0].a/n1152 ), .B(
        \SUBBYTES[0].a/n1151 ), .Z(\SUBBYTES[0].a/n1571 ) );
  XOR \SUBBYTES[0].a/U4368  ( .A(\w1[0][76] ), .B(\SUBBYTES[0].a/n1153 ), .Z(
        \SUBBYTES[0].a/n1151 ) );
  XOR \SUBBYTES[0].a/U4367  ( .A(\SUBBYTES[0].a/w1459 ), .B(\w1[0][78] ), .Z(
        \SUBBYTES[0].a/n1152 ) );
  XOR \SUBBYTES[0].a/U4366  ( .A(\SUBBYTES[0].a/w1433 ), .B(
        \SUBBYTES[0].a/w1440 ), .Z(\SUBBYTES[0].a/n1153 ) );
  XOR \SUBBYTES[0].a/U4365  ( .A(\SUBBYTES[0].a/n1155 ), .B(
        \SUBBYTES[0].a/n1154 ), .Z(\SUBBYTES[0].a/n1569 ) );
  XOR \SUBBYTES[0].a/U4364  ( .A(\w1[0][73] ), .B(\SUBBYTES[0].a/n1156 ), .Z(
        \SUBBYTES[0].a/n1154 ) );
  XOR \SUBBYTES[0].a/U4363  ( .A(\SUBBYTES[0].a/w1458 ), .B(\w1[0][77] ), .Z(
        \SUBBYTES[0].a/n1155 ) );
  XOR \SUBBYTES[0].a/U4362  ( .A(\SUBBYTES[0].a/w1434 ), .B(
        \SUBBYTES[0].a/w1441 ), .Z(\SUBBYTES[0].a/n1156 ) );
  XOR \SUBBYTES[0].a/U4361  ( .A(\SUBBYTES[0].a/n1571 ), .B(
        \SUBBYTES[0].a/n1569 ), .Z(\SUBBYTES[0].a/w1464 ) );
  XOR \SUBBYTES[0].a/U4360  ( .A(\w1[0][77] ), .B(\SUBBYTES[0].a/n1157 ), .Z(
        \SUBBYTES[0].a/n1572 ) );
  XOR \SUBBYTES[0].a/U4359  ( .A(\SUBBYTES[0].a/w1426 ), .B(
        \SUBBYTES[0].a/w1436 ), .Z(\SUBBYTES[0].a/n1157 ) );
  XOR \SUBBYTES[0].a/U4358  ( .A(\SUBBYTES[0].a/n1159 ), .B(
        \SUBBYTES[0].a/n1158 ), .Z(\SUBBYTES[0].a/w1451 ) );
  XOR \SUBBYTES[0].a/U4357  ( .A(\SUBBYTES[0].a/n1572 ), .B(
        \SUBBYTES[0].a/n1160 ), .Z(\SUBBYTES[0].a/n1158 ) );
  XOR \SUBBYTES[0].a/U4356  ( .A(\w1[0][76] ), .B(\SUBBYTES[0].a/w1515 ), .Z(
        \SUBBYTES[0].a/n1159 ) );
  XOR \SUBBYTES[0].a/U4355  ( .A(\SUBBYTES[0].a/w1428 ), .B(
        \SUBBYTES[0].a/w1433 ), .Z(\SUBBYTES[0].a/n1160 ) );
  XOR \SUBBYTES[0].a/U4354  ( .A(\SUBBYTES[0].a/n1162 ), .B(
        \SUBBYTES[0].a/n1161 ), .Z(\SUBBYTES[0].a/n1570 ) );
  XOR \SUBBYTES[0].a/U4353  ( .A(\SUBBYTES[0].a/w1461 ), .B(\w1[0][79] ), .Z(
        \SUBBYTES[0].a/n1161 ) );
  XOR \SUBBYTES[0].a/U4352  ( .A(\SUBBYTES[0].a/w1436 ), .B(
        \SUBBYTES[0].a/w1443 ), .Z(\SUBBYTES[0].a/n1162 ) );
  XOR \SUBBYTES[0].a/U4351  ( .A(\SUBBYTES[0].a/n1569 ), .B(
        \SUBBYTES[0].a/n1570 ), .Z(\SUBBYTES[0].a/w1463 ) );
  XOR \SUBBYTES[0].a/U4350  ( .A(\w1[0][75] ), .B(\SUBBYTES[0].a/n1163 ), .Z(
        \SUBBYTES[0].a/n1573 ) );
  XOR \SUBBYTES[0].a/U4349  ( .A(\SUBBYTES[0].a/w1425 ), .B(
        \SUBBYTES[0].a/w1428 ), .Z(\SUBBYTES[0].a/n1163 ) );
  XOR \SUBBYTES[0].a/U4348  ( .A(\SUBBYTES[0].a/n1165 ), .B(
        \SUBBYTES[0].a/n1164 ), .Z(\SUBBYTES[0].a/w1452 ) );
  XOR \SUBBYTES[0].a/U4347  ( .A(\SUBBYTES[0].a/n1573 ), .B(
        \SUBBYTES[0].a/n1166 ), .Z(\SUBBYTES[0].a/n1164 ) );
  XOR \SUBBYTES[0].a/U4346  ( .A(\w1[0][78] ), .B(\SUBBYTES[0].a/w1494 ), .Z(
        \SUBBYTES[0].a/n1165 ) );
  XOR \SUBBYTES[0].a/U4345  ( .A(\SUBBYTES[0].a/w1433 ), .B(
        \SUBBYTES[0].a/w1434 ), .Z(\SUBBYTES[0].a/n1166 ) );
  XOR \SUBBYTES[0].a/U4344  ( .A(\SUBBYTES[0].a/n1571 ), .B(
        \SUBBYTES[0].a/n1570 ), .Z(\SUBBYTES[0].a/w1472 ) );
  XOR \SUBBYTES[0].a/U4343  ( .A(\SUBBYTES[0].a/n1168 ), .B(
        \SUBBYTES[0].a/n1167 ), .Z(\SUBBYTES[0].a/w1473 ) );
  XOR \SUBBYTES[0].a/U4342  ( .A(\w1[0][79] ), .B(\SUBBYTES[0].a/n1572 ), .Z(
        \SUBBYTES[0].a/n1167 ) );
  XOR \SUBBYTES[0].a/U4341  ( .A(\SUBBYTES[0].a/w1425 ), .B(
        \SUBBYTES[0].a/w1434 ), .Z(\SUBBYTES[0].a/n1168 ) );
  XOR \SUBBYTES[0].a/U4340  ( .A(\SUBBYTES[0].a/n1170 ), .B(
        \SUBBYTES[0].a/n1169 ), .Z(\SUBBYTES[0].a/w1449 ) );
  XOR \SUBBYTES[0].a/U4339  ( .A(\SUBBYTES[0].a/n1172 ), .B(
        \SUBBYTES[0].a/n1171 ), .Z(\SUBBYTES[0].a/n1169 ) );
  XOR \SUBBYTES[0].a/U4338  ( .A(\w1[0][79] ), .B(\SUBBYTES[0].a/w1533 ), .Z(
        \SUBBYTES[0].a/n1170 ) );
  XOR \SUBBYTES[0].a/U4337  ( .A(\SUBBYTES[0].a/w1440 ), .B(
        \SUBBYTES[0].a/w1443 ), .Z(\SUBBYTES[0].a/n1171 ) );
  XOR \SUBBYTES[0].a/U4336  ( .A(\SUBBYTES[0].a/w1426 ), .B(
        \SUBBYTES[0].a/w1428 ), .Z(\SUBBYTES[0].a/n1172 ) );
  XOR \SUBBYTES[0].a/U4335  ( .A(\SUBBYTES[0].a/n1174 ), .B(
        \SUBBYTES[0].a/n1173 ), .Z(\SUBBYTES[0].a/w1450 ) );
  XOR \SUBBYTES[0].a/U4334  ( .A(\SUBBYTES[0].a/n1573 ), .B(
        \SUBBYTES[0].a/n1175 ), .Z(\SUBBYTES[0].a/n1173 ) );
  XOR \SUBBYTES[0].a/U4333  ( .A(\w1[0][77] ), .B(\SUBBYTES[0].a/n1574 ), .Z(
        \SUBBYTES[0].a/n1174 ) );
  XOR \SUBBYTES[0].a/U4332  ( .A(\SUBBYTES[0].a/w1440 ), .B(
        \SUBBYTES[0].a/w1441 ), .Z(\SUBBYTES[0].a/n1175 ) );
  XOR \SUBBYTES[0].a/U4331  ( .A(\SUBBYTES[0].a/n1177 ), .B(
        \SUBBYTES[0].a/n1176 ), .Z(\SUBBYTES[0].a/w1466 ) );
  XOR \SUBBYTES[0].a/U4330  ( .A(\w1[0][73] ), .B(\SUBBYTES[0].a/n1178 ), .Z(
        \SUBBYTES[0].a/n1176 ) );
  XOR \SUBBYTES[0].a/U4329  ( .A(\SUBBYTES[0].a/w1441 ), .B(
        \SUBBYTES[0].a/w1443 ), .Z(\SUBBYTES[0].a/n1177 ) );
  XOR \SUBBYTES[0].a/U4328  ( .A(\SUBBYTES[0].a/w1425 ), .B(
        \SUBBYTES[0].a/w1426 ), .Z(\SUBBYTES[0].a/n1178 ) );
  XOR \SUBBYTES[0].a/U4327  ( .A(\w1[0][81] ), .B(\SUBBYTES[0].a/n1179 ), .Z(
        \SUBBYTES[0].a/n1575 ) );
  XOR \SUBBYTES[0].a/U4326  ( .A(\w1[0][83] ), .B(\w1[0][82] ), .Z(
        \SUBBYTES[0].a/n1179 ) );
  XOR \SUBBYTES[0].a/U4325  ( .A(\w1[0][86] ), .B(\SUBBYTES[0].a/n1575 ), .Z(
        \SUBBYTES[0].a/w1308 ) );
  XOR \SUBBYTES[0].a/U4324  ( .A(\w1[0][80] ), .B(\SUBBYTES[0].a/w1308 ), .Z(
        \SUBBYTES[0].a/w1195 ) );
  XOR \SUBBYTES[0].a/U4323  ( .A(\w1[0][80] ), .B(\SUBBYTES[0].a/n1180 ), .Z(
        \SUBBYTES[0].a/w1196 ) );
  XOR \SUBBYTES[0].a/U4322  ( .A(\w1[0][86] ), .B(\w1[0][85] ), .Z(
        \SUBBYTES[0].a/n1180 ) );
  XOR \SUBBYTES[0].a/U4321  ( .A(\w1[0][85] ), .B(\SUBBYTES[0].a/n1575 ), .Z(
        \SUBBYTES[0].a/w1326 ) );
  XOR \SUBBYTES[0].a/U4320  ( .A(\SUBBYTES[0].a/n1182 ), .B(
        \SUBBYTES[0].a/n1181 ), .Z(\SUBBYTES[0].a/w1319 ) );
  XOR \SUBBYTES[0].a/U4319  ( .A(\w1[0][83] ), .B(\w1[0][81] ), .Z(
        \SUBBYTES[0].a/n1181 ) );
  XOR \SUBBYTES[0].a/U4318  ( .A(\w1[0][87] ), .B(\w1[0][84] ), .Z(
        \SUBBYTES[0].a/n1182 ) );
  XOR \SUBBYTES[0].a/U4317  ( .A(\w1[0][80] ), .B(\SUBBYTES[0].a/w1319 ), .Z(
        \SUBBYTES[0].a/w1198 ) );
  XOR \SUBBYTES[0].a/U4316  ( .A(\SUBBYTES[0].a/n1184 ), .B(
        \SUBBYTES[0].a/n1183 ), .Z(\SUBBYTES[0].a/w1306 ) );
  XOR \SUBBYTES[0].a/U4315  ( .A(\SUBBYTES[0].a/w1267 ), .B(n1158), .Z(
        \SUBBYTES[0].a/n1183 ) );
  XOR \SUBBYTES[0].a/U4314  ( .A(\SUBBYTES[0].a/w1260 ), .B(
        \SUBBYTES[0].a/w1263 ), .Z(\SUBBYTES[0].a/n1184 ) );
  XOR \SUBBYTES[0].a/U4313  ( .A(\SUBBYTES[0].a/n1186 ), .B(
        \SUBBYTES[0].a/n1185 ), .Z(\SUBBYTES[0].a/w1307 ) );
  XOR \SUBBYTES[0].a/U4312  ( .A(\SUBBYTES[0].a/w1267 ), .B(
        \SUBBYTES[0].a/n60 ), .Z(\SUBBYTES[0].a/n1185 ) );
  XOR \SUBBYTES[0].a/U4311  ( .A(\SUBBYTES[0].a/w1260 ), .B(
        \SUBBYTES[0].a/n59 ), .Z(\SUBBYTES[0].a/n1186 ) );
  XOR \SUBBYTES[0].a/U4310  ( .A(\SUBBYTES[0].a/w1319 ), .B(
        \SUBBYTES[0].a/n1187 ), .Z(\SUBBYTES[0].a/w1309 ) );
  XOR \SUBBYTES[0].a/U4309  ( .A(\w1[0][86] ), .B(\w1[0][85] ), .Z(
        \SUBBYTES[0].a/n1187 ) );
  XOR \SUBBYTES[0].a/U4308  ( .A(\SUBBYTES[0].a/n1189 ), .B(
        \SUBBYTES[0].a/n1188 ), .Z(\SUBBYTES[0].a/w1310 ) );
  XOR \SUBBYTES[0].a/U4307  ( .A(\SUBBYTES[0].a/n60 ), .B(n1158), .Z(
        \SUBBYTES[0].a/n1188 ) );
  XOR \SUBBYTES[0].a/U4306  ( .A(\SUBBYTES[0].a/n59 ), .B(
        \SUBBYTES[0].a/w1263 ), .Z(\SUBBYTES[0].a/n1189 ) );
  XOR \SUBBYTES[0].a/U4305  ( .A(\w1[0][87] ), .B(\w1[0][82] ), .Z(
        \SUBBYTES[0].a/n1581 ) );
  XOR \SUBBYTES[0].a/U4304  ( .A(\SUBBYTES[0].a/n1581 ), .B(
        \SUBBYTES[0].a/n1190 ), .Z(\SUBBYTES[0].a/w1311 ) );
  XOR \SUBBYTES[0].a/U4303  ( .A(\w1[0][85] ), .B(\w1[0][84] ), .Z(
        \SUBBYTES[0].a/n1190 ) );
  XOR \SUBBYTES[0].a/U4302  ( .A(\w1[0][87] ), .B(\SUBBYTES[0].a/w1196 ), .Z(
        \SUBBYTES[0].a/w1199 ) );
  XOR \SUBBYTES[0].a/U4301  ( .A(\w1[0][81] ), .B(\SUBBYTES[0].a/w1196 ), .Z(
        \SUBBYTES[0].a/w1200 ) );
  XOR \SUBBYTES[0].a/U4300  ( .A(\w1[0][84] ), .B(\SUBBYTES[0].a/w1196 ), .Z(
        \SUBBYTES[0].a/w1201 ) );
  XOR \SUBBYTES[0].a/U4299  ( .A(\SUBBYTES[0].a/w1200 ), .B(
        \SUBBYTES[0].a/n1581 ), .Z(\SUBBYTES[0].a/w1202 ) );
  XOR \SUBBYTES[0].a/U4298  ( .A(\SUBBYTES[0].a/n1581 ), .B(
        \SUBBYTES[0].a/n1191 ), .Z(\SUBBYTES[0].a/w1287 ) );
  XOR \SUBBYTES[0].a/U4297  ( .A(\w1[0][84] ), .B(\w1[0][81] ), .Z(
        \SUBBYTES[0].a/n1191 ) );
  XOR \SUBBYTES[0].a/U4296  ( .A(\SUBBYTES[0].a/n1193 ), .B(
        \SUBBYTES[0].a/n1192 ), .Z(\SUBBYTES[0].a/n1578 ) );
  XOR \SUBBYTES[0].a/U4295  ( .A(\w1[0][84] ), .B(\SUBBYTES[0].a/n1194 ), .Z(
        \SUBBYTES[0].a/n1192 ) );
  XOR \SUBBYTES[0].a/U4294  ( .A(\SUBBYTES[0].a/w1252 ), .B(\w1[0][86] ), .Z(
        \SUBBYTES[0].a/n1193 ) );
  XOR \SUBBYTES[0].a/U4293  ( .A(\SUBBYTES[0].a/w1226 ), .B(
        \SUBBYTES[0].a/w1233 ), .Z(\SUBBYTES[0].a/n1194 ) );
  XOR \SUBBYTES[0].a/U4292  ( .A(\SUBBYTES[0].a/n1196 ), .B(
        \SUBBYTES[0].a/n1195 ), .Z(\SUBBYTES[0].a/n1576 ) );
  XOR \SUBBYTES[0].a/U4291  ( .A(\w1[0][81] ), .B(\SUBBYTES[0].a/n1197 ), .Z(
        \SUBBYTES[0].a/n1195 ) );
  XOR \SUBBYTES[0].a/U4290  ( .A(\SUBBYTES[0].a/w1251 ), .B(\w1[0][85] ), .Z(
        \SUBBYTES[0].a/n1196 ) );
  XOR \SUBBYTES[0].a/U4289  ( .A(\SUBBYTES[0].a/w1227 ), .B(
        \SUBBYTES[0].a/w1234 ), .Z(\SUBBYTES[0].a/n1197 ) );
  XOR \SUBBYTES[0].a/U4288  ( .A(\SUBBYTES[0].a/n1578 ), .B(
        \SUBBYTES[0].a/n1576 ), .Z(\SUBBYTES[0].a/w1257 ) );
  XOR \SUBBYTES[0].a/U4287  ( .A(\w1[0][85] ), .B(\SUBBYTES[0].a/n1198 ), .Z(
        \SUBBYTES[0].a/n1579 ) );
  XOR \SUBBYTES[0].a/U4286  ( .A(\SUBBYTES[0].a/w1219 ), .B(
        \SUBBYTES[0].a/w1229 ), .Z(\SUBBYTES[0].a/n1198 ) );
  XOR \SUBBYTES[0].a/U4285  ( .A(\SUBBYTES[0].a/n1200 ), .B(
        \SUBBYTES[0].a/n1199 ), .Z(\SUBBYTES[0].a/w1244 ) );
  XOR \SUBBYTES[0].a/U4284  ( .A(\SUBBYTES[0].a/n1579 ), .B(
        \SUBBYTES[0].a/n1201 ), .Z(\SUBBYTES[0].a/n1199 ) );
  XOR \SUBBYTES[0].a/U4283  ( .A(\w1[0][84] ), .B(\SUBBYTES[0].a/w1308 ), .Z(
        \SUBBYTES[0].a/n1200 ) );
  XOR \SUBBYTES[0].a/U4282  ( .A(\SUBBYTES[0].a/w1221 ), .B(
        \SUBBYTES[0].a/w1226 ), .Z(\SUBBYTES[0].a/n1201 ) );
  XOR \SUBBYTES[0].a/U4281  ( .A(\SUBBYTES[0].a/n1203 ), .B(
        \SUBBYTES[0].a/n1202 ), .Z(\SUBBYTES[0].a/n1577 ) );
  XOR \SUBBYTES[0].a/U4280  ( .A(\SUBBYTES[0].a/w1254 ), .B(\w1[0][87] ), .Z(
        \SUBBYTES[0].a/n1202 ) );
  XOR \SUBBYTES[0].a/U4279  ( .A(\SUBBYTES[0].a/w1229 ), .B(
        \SUBBYTES[0].a/w1236 ), .Z(\SUBBYTES[0].a/n1203 ) );
  XOR \SUBBYTES[0].a/U4278  ( .A(\SUBBYTES[0].a/n1576 ), .B(
        \SUBBYTES[0].a/n1577 ), .Z(\SUBBYTES[0].a/w1256 ) );
  XOR \SUBBYTES[0].a/U4277  ( .A(\w1[0][83] ), .B(\SUBBYTES[0].a/n1204 ), .Z(
        \SUBBYTES[0].a/n1580 ) );
  XOR \SUBBYTES[0].a/U4276  ( .A(\SUBBYTES[0].a/w1218 ), .B(
        \SUBBYTES[0].a/w1221 ), .Z(\SUBBYTES[0].a/n1204 ) );
  XOR \SUBBYTES[0].a/U4275  ( .A(\SUBBYTES[0].a/n1206 ), .B(
        \SUBBYTES[0].a/n1205 ), .Z(\SUBBYTES[0].a/w1245 ) );
  XOR \SUBBYTES[0].a/U4274  ( .A(\SUBBYTES[0].a/n1580 ), .B(
        \SUBBYTES[0].a/n1207 ), .Z(\SUBBYTES[0].a/n1205 ) );
  XOR \SUBBYTES[0].a/U4273  ( .A(\w1[0][86] ), .B(\SUBBYTES[0].a/w1287 ), .Z(
        \SUBBYTES[0].a/n1206 ) );
  XOR \SUBBYTES[0].a/U4272  ( .A(\SUBBYTES[0].a/w1226 ), .B(
        \SUBBYTES[0].a/w1227 ), .Z(\SUBBYTES[0].a/n1207 ) );
  XOR \SUBBYTES[0].a/U4271  ( .A(\SUBBYTES[0].a/n1578 ), .B(
        \SUBBYTES[0].a/n1577 ), .Z(\SUBBYTES[0].a/w1265 ) );
  XOR \SUBBYTES[0].a/U4270  ( .A(\SUBBYTES[0].a/n1209 ), .B(
        \SUBBYTES[0].a/n1208 ), .Z(\SUBBYTES[0].a/w1266 ) );
  XOR \SUBBYTES[0].a/U4269  ( .A(\w1[0][87] ), .B(\SUBBYTES[0].a/n1579 ), .Z(
        \SUBBYTES[0].a/n1208 ) );
  XOR \SUBBYTES[0].a/U4268  ( .A(\SUBBYTES[0].a/w1218 ), .B(
        \SUBBYTES[0].a/w1227 ), .Z(\SUBBYTES[0].a/n1209 ) );
  XOR \SUBBYTES[0].a/U4267  ( .A(\SUBBYTES[0].a/n1211 ), .B(
        \SUBBYTES[0].a/n1210 ), .Z(\SUBBYTES[0].a/w1242 ) );
  XOR \SUBBYTES[0].a/U4266  ( .A(\SUBBYTES[0].a/n1213 ), .B(
        \SUBBYTES[0].a/n1212 ), .Z(\SUBBYTES[0].a/n1210 ) );
  XOR \SUBBYTES[0].a/U4265  ( .A(\w1[0][87] ), .B(\SUBBYTES[0].a/w1326 ), .Z(
        \SUBBYTES[0].a/n1211 ) );
  XOR \SUBBYTES[0].a/U4264  ( .A(\SUBBYTES[0].a/w1233 ), .B(
        \SUBBYTES[0].a/w1236 ), .Z(\SUBBYTES[0].a/n1212 ) );
  XOR \SUBBYTES[0].a/U4263  ( .A(\SUBBYTES[0].a/w1219 ), .B(
        \SUBBYTES[0].a/w1221 ), .Z(\SUBBYTES[0].a/n1213 ) );
  XOR \SUBBYTES[0].a/U4262  ( .A(\SUBBYTES[0].a/n1215 ), .B(
        \SUBBYTES[0].a/n1214 ), .Z(\SUBBYTES[0].a/w1243 ) );
  XOR \SUBBYTES[0].a/U4261  ( .A(\SUBBYTES[0].a/n1580 ), .B(
        \SUBBYTES[0].a/n1216 ), .Z(\SUBBYTES[0].a/n1214 ) );
  XOR \SUBBYTES[0].a/U4260  ( .A(\w1[0][85] ), .B(\SUBBYTES[0].a/n1581 ), .Z(
        \SUBBYTES[0].a/n1215 ) );
  XOR \SUBBYTES[0].a/U4259  ( .A(\SUBBYTES[0].a/w1233 ), .B(
        \SUBBYTES[0].a/w1234 ), .Z(\SUBBYTES[0].a/n1216 ) );
  XOR \SUBBYTES[0].a/U4258  ( .A(\SUBBYTES[0].a/n1218 ), .B(
        \SUBBYTES[0].a/n1217 ), .Z(\SUBBYTES[0].a/w1259 ) );
  XOR \SUBBYTES[0].a/U4257  ( .A(\w1[0][81] ), .B(\SUBBYTES[0].a/n1219 ), .Z(
        \SUBBYTES[0].a/n1217 ) );
  XOR \SUBBYTES[0].a/U4256  ( .A(\SUBBYTES[0].a/w1234 ), .B(
        \SUBBYTES[0].a/w1236 ), .Z(\SUBBYTES[0].a/n1218 ) );
  XOR \SUBBYTES[0].a/U4255  ( .A(\SUBBYTES[0].a/w1218 ), .B(
        \SUBBYTES[0].a/w1219 ), .Z(\SUBBYTES[0].a/n1219 ) );
  XOR \SUBBYTES[0].a/U4254  ( .A(\w1[0][89] ), .B(\SUBBYTES[0].a/n1220 ), .Z(
        \SUBBYTES[0].a/n1582 ) );
  XOR \SUBBYTES[0].a/U4253  ( .A(\w1[0][91] ), .B(\w1[0][90] ), .Z(
        \SUBBYTES[0].a/n1220 ) );
  XOR \SUBBYTES[0].a/U4252  ( .A(\w1[0][94] ), .B(\SUBBYTES[0].a/n1582 ), .Z(
        \SUBBYTES[0].a/w1101 ) );
  XOR \SUBBYTES[0].a/U4251  ( .A(\w1[0][88] ), .B(\SUBBYTES[0].a/w1101 ), .Z(
        \SUBBYTES[0].a/w988 ) );
  XOR \SUBBYTES[0].a/U4250  ( .A(\w1[0][88] ), .B(\SUBBYTES[0].a/n1221 ), .Z(
        \SUBBYTES[0].a/w989 ) );
  XOR \SUBBYTES[0].a/U4249  ( .A(\w1[0][94] ), .B(\w1[0][93] ), .Z(
        \SUBBYTES[0].a/n1221 ) );
  XOR \SUBBYTES[0].a/U4248  ( .A(\w1[0][93] ), .B(\SUBBYTES[0].a/n1582 ), .Z(
        \SUBBYTES[0].a/w1119 ) );
  XOR \SUBBYTES[0].a/U4247  ( .A(\SUBBYTES[0].a/n1223 ), .B(
        \SUBBYTES[0].a/n1222 ), .Z(\SUBBYTES[0].a/w1112 ) );
  XOR \SUBBYTES[0].a/U4246  ( .A(\w1[0][91] ), .B(\w1[0][89] ), .Z(
        \SUBBYTES[0].a/n1222 ) );
  XOR \SUBBYTES[0].a/U4245  ( .A(\w1[0][95] ), .B(\w1[0][92] ), .Z(
        \SUBBYTES[0].a/n1223 ) );
  XOR \SUBBYTES[0].a/U4244  ( .A(\w1[0][88] ), .B(\SUBBYTES[0].a/w1112 ), .Z(
        \SUBBYTES[0].a/w991 ) );
  XOR \SUBBYTES[0].a/U4243  ( .A(\SUBBYTES[0].a/n1225 ), .B(
        \SUBBYTES[0].a/n1224 ), .Z(\SUBBYTES[0].a/w1099 ) );
  XOR \SUBBYTES[0].a/U4242  ( .A(\SUBBYTES[0].a/w1060 ), .B(n1157), .Z(
        \SUBBYTES[0].a/n1224 ) );
  XOR \SUBBYTES[0].a/U4241  ( .A(\SUBBYTES[0].a/w1053 ), .B(
        \SUBBYTES[0].a/w1056 ), .Z(\SUBBYTES[0].a/n1225 ) );
  XOR \SUBBYTES[0].a/U4240  ( .A(\SUBBYTES[0].a/n1227 ), .B(
        \SUBBYTES[0].a/n1226 ), .Z(\SUBBYTES[0].a/w1100 ) );
  XOR \SUBBYTES[0].a/U4239  ( .A(\SUBBYTES[0].a/w1060 ), .B(
        \SUBBYTES[0].a/n50 ), .Z(\SUBBYTES[0].a/n1226 ) );
  XOR \SUBBYTES[0].a/U4238  ( .A(\SUBBYTES[0].a/w1053 ), .B(
        \SUBBYTES[0].a/n49 ), .Z(\SUBBYTES[0].a/n1227 ) );
  XOR \SUBBYTES[0].a/U4237  ( .A(\SUBBYTES[0].a/w1112 ), .B(
        \SUBBYTES[0].a/n1228 ), .Z(\SUBBYTES[0].a/w1102 ) );
  XOR \SUBBYTES[0].a/U4236  ( .A(\w1[0][94] ), .B(\w1[0][93] ), .Z(
        \SUBBYTES[0].a/n1228 ) );
  XOR \SUBBYTES[0].a/U4235  ( .A(\SUBBYTES[0].a/n1230 ), .B(
        \SUBBYTES[0].a/n1229 ), .Z(\SUBBYTES[0].a/w1103 ) );
  XOR \SUBBYTES[0].a/U4234  ( .A(\SUBBYTES[0].a/n50 ), .B(n1157), .Z(
        \SUBBYTES[0].a/n1229 ) );
  XOR \SUBBYTES[0].a/U4233  ( .A(\SUBBYTES[0].a/n49 ), .B(
        \SUBBYTES[0].a/w1056 ), .Z(\SUBBYTES[0].a/n1230 ) );
  XOR \SUBBYTES[0].a/U4232  ( .A(\w1[0][95] ), .B(\w1[0][90] ), .Z(
        \SUBBYTES[0].a/n1588 ) );
  XOR \SUBBYTES[0].a/U4231  ( .A(\SUBBYTES[0].a/n1588 ), .B(
        \SUBBYTES[0].a/n1231 ), .Z(\SUBBYTES[0].a/w1104 ) );
  XOR \SUBBYTES[0].a/U4230  ( .A(\w1[0][93] ), .B(\w1[0][92] ), .Z(
        \SUBBYTES[0].a/n1231 ) );
  XOR \SUBBYTES[0].a/U4229  ( .A(\w1[0][95] ), .B(\SUBBYTES[0].a/w989 ), .Z(
        \SUBBYTES[0].a/w992 ) );
  XOR \SUBBYTES[0].a/U4228  ( .A(\w1[0][89] ), .B(\SUBBYTES[0].a/w989 ), .Z(
        \SUBBYTES[0].a/w993 ) );
  XOR \SUBBYTES[0].a/U4227  ( .A(\w1[0][92] ), .B(\SUBBYTES[0].a/w989 ), .Z(
        \SUBBYTES[0].a/w994 ) );
  XOR \SUBBYTES[0].a/U4226  ( .A(\SUBBYTES[0].a/w993 ), .B(
        \SUBBYTES[0].a/n1588 ), .Z(\SUBBYTES[0].a/w995 ) );
  XOR \SUBBYTES[0].a/U4225  ( .A(\SUBBYTES[0].a/n1588 ), .B(
        \SUBBYTES[0].a/n1232 ), .Z(\SUBBYTES[0].a/w1080 ) );
  XOR \SUBBYTES[0].a/U4224  ( .A(\w1[0][92] ), .B(\w1[0][89] ), .Z(
        \SUBBYTES[0].a/n1232 ) );
  XOR \SUBBYTES[0].a/U4223  ( .A(\SUBBYTES[0].a/n1234 ), .B(
        \SUBBYTES[0].a/n1233 ), .Z(\SUBBYTES[0].a/n1585 ) );
  XOR \SUBBYTES[0].a/U4222  ( .A(\w1[0][92] ), .B(\SUBBYTES[0].a/n1235 ), .Z(
        \SUBBYTES[0].a/n1233 ) );
  XOR \SUBBYTES[0].a/U4221  ( .A(\SUBBYTES[0].a/w1045 ), .B(\w1[0][94] ), .Z(
        \SUBBYTES[0].a/n1234 ) );
  XOR \SUBBYTES[0].a/U4220  ( .A(\SUBBYTES[0].a/w1019 ), .B(
        \SUBBYTES[0].a/w1026 ), .Z(\SUBBYTES[0].a/n1235 ) );
  XOR \SUBBYTES[0].a/U4219  ( .A(\SUBBYTES[0].a/n1237 ), .B(
        \SUBBYTES[0].a/n1236 ), .Z(\SUBBYTES[0].a/n1583 ) );
  XOR \SUBBYTES[0].a/U4218  ( .A(\w1[0][89] ), .B(\SUBBYTES[0].a/n1238 ), .Z(
        \SUBBYTES[0].a/n1236 ) );
  XOR \SUBBYTES[0].a/U4217  ( .A(\SUBBYTES[0].a/w1044 ), .B(\w1[0][93] ), .Z(
        \SUBBYTES[0].a/n1237 ) );
  XOR \SUBBYTES[0].a/U4216  ( .A(\SUBBYTES[0].a/w1020 ), .B(
        \SUBBYTES[0].a/w1027 ), .Z(\SUBBYTES[0].a/n1238 ) );
  XOR \SUBBYTES[0].a/U4215  ( .A(\SUBBYTES[0].a/n1585 ), .B(
        \SUBBYTES[0].a/n1583 ), .Z(\SUBBYTES[0].a/w1050 ) );
  XOR \SUBBYTES[0].a/U4214  ( .A(\w1[0][93] ), .B(\SUBBYTES[0].a/n1239 ), .Z(
        \SUBBYTES[0].a/n1586 ) );
  XOR \SUBBYTES[0].a/U4213  ( .A(\SUBBYTES[0].a/w1012 ), .B(
        \SUBBYTES[0].a/w1022 ), .Z(\SUBBYTES[0].a/n1239 ) );
  XOR \SUBBYTES[0].a/U4212  ( .A(\SUBBYTES[0].a/n1241 ), .B(
        \SUBBYTES[0].a/n1240 ), .Z(\SUBBYTES[0].a/w1037 ) );
  XOR \SUBBYTES[0].a/U4211  ( .A(\SUBBYTES[0].a/n1586 ), .B(
        \SUBBYTES[0].a/n1242 ), .Z(\SUBBYTES[0].a/n1240 ) );
  XOR \SUBBYTES[0].a/U4210  ( .A(\w1[0][92] ), .B(\SUBBYTES[0].a/w1101 ), .Z(
        \SUBBYTES[0].a/n1241 ) );
  XOR \SUBBYTES[0].a/U4209  ( .A(\SUBBYTES[0].a/w1014 ), .B(
        \SUBBYTES[0].a/w1019 ), .Z(\SUBBYTES[0].a/n1242 ) );
  XOR \SUBBYTES[0].a/U4208  ( .A(\SUBBYTES[0].a/n1244 ), .B(
        \SUBBYTES[0].a/n1243 ), .Z(\SUBBYTES[0].a/n1584 ) );
  XOR \SUBBYTES[0].a/U4207  ( .A(\SUBBYTES[0].a/w1047 ), .B(\w1[0][95] ), .Z(
        \SUBBYTES[0].a/n1243 ) );
  XOR \SUBBYTES[0].a/U4206  ( .A(\SUBBYTES[0].a/w1022 ), .B(
        \SUBBYTES[0].a/w1029 ), .Z(\SUBBYTES[0].a/n1244 ) );
  XOR \SUBBYTES[0].a/U4205  ( .A(\SUBBYTES[0].a/n1583 ), .B(
        \SUBBYTES[0].a/n1584 ), .Z(\SUBBYTES[0].a/w1049 ) );
  XOR \SUBBYTES[0].a/U4204  ( .A(\w1[0][91] ), .B(\SUBBYTES[0].a/n1245 ), .Z(
        \SUBBYTES[0].a/n1587 ) );
  XOR \SUBBYTES[0].a/U4203  ( .A(\SUBBYTES[0].a/w1011 ), .B(
        \SUBBYTES[0].a/w1014 ), .Z(\SUBBYTES[0].a/n1245 ) );
  XOR \SUBBYTES[0].a/U4202  ( .A(\SUBBYTES[0].a/n1247 ), .B(
        \SUBBYTES[0].a/n1246 ), .Z(\SUBBYTES[0].a/w1038 ) );
  XOR \SUBBYTES[0].a/U4201  ( .A(\SUBBYTES[0].a/n1587 ), .B(
        \SUBBYTES[0].a/n1248 ), .Z(\SUBBYTES[0].a/n1246 ) );
  XOR \SUBBYTES[0].a/U4200  ( .A(\w1[0][94] ), .B(\SUBBYTES[0].a/w1080 ), .Z(
        \SUBBYTES[0].a/n1247 ) );
  XOR \SUBBYTES[0].a/U4199  ( .A(\SUBBYTES[0].a/w1019 ), .B(
        \SUBBYTES[0].a/w1020 ), .Z(\SUBBYTES[0].a/n1248 ) );
  XOR \SUBBYTES[0].a/U4198  ( .A(\SUBBYTES[0].a/n1585 ), .B(
        \SUBBYTES[0].a/n1584 ), .Z(\SUBBYTES[0].a/w1058 ) );
  XOR \SUBBYTES[0].a/U4197  ( .A(\SUBBYTES[0].a/n1250 ), .B(
        \SUBBYTES[0].a/n1249 ), .Z(\SUBBYTES[0].a/w1059 ) );
  XOR \SUBBYTES[0].a/U4196  ( .A(\w1[0][95] ), .B(\SUBBYTES[0].a/n1586 ), .Z(
        \SUBBYTES[0].a/n1249 ) );
  XOR \SUBBYTES[0].a/U4195  ( .A(\SUBBYTES[0].a/w1011 ), .B(
        \SUBBYTES[0].a/w1020 ), .Z(\SUBBYTES[0].a/n1250 ) );
  XOR \SUBBYTES[0].a/U4194  ( .A(\SUBBYTES[0].a/n1252 ), .B(
        \SUBBYTES[0].a/n1251 ), .Z(\SUBBYTES[0].a/w1035 ) );
  XOR \SUBBYTES[0].a/U4193  ( .A(\SUBBYTES[0].a/n1254 ), .B(
        \SUBBYTES[0].a/n1253 ), .Z(\SUBBYTES[0].a/n1251 ) );
  XOR \SUBBYTES[0].a/U4192  ( .A(\w1[0][95] ), .B(\SUBBYTES[0].a/w1119 ), .Z(
        \SUBBYTES[0].a/n1252 ) );
  XOR \SUBBYTES[0].a/U4191  ( .A(\SUBBYTES[0].a/w1026 ), .B(
        \SUBBYTES[0].a/w1029 ), .Z(\SUBBYTES[0].a/n1253 ) );
  XOR \SUBBYTES[0].a/U4190  ( .A(\SUBBYTES[0].a/w1012 ), .B(
        \SUBBYTES[0].a/w1014 ), .Z(\SUBBYTES[0].a/n1254 ) );
  XOR \SUBBYTES[0].a/U4189  ( .A(\SUBBYTES[0].a/n1256 ), .B(
        \SUBBYTES[0].a/n1255 ), .Z(\SUBBYTES[0].a/w1036 ) );
  XOR \SUBBYTES[0].a/U4188  ( .A(\SUBBYTES[0].a/n1587 ), .B(
        \SUBBYTES[0].a/n1257 ), .Z(\SUBBYTES[0].a/n1255 ) );
  XOR \SUBBYTES[0].a/U4187  ( .A(\w1[0][93] ), .B(\SUBBYTES[0].a/n1588 ), .Z(
        \SUBBYTES[0].a/n1256 ) );
  XOR \SUBBYTES[0].a/U4186  ( .A(\SUBBYTES[0].a/w1026 ), .B(
        \SUBBYTES[0].a/w1027 ), .Z(\SUBBYTES[0].a/n1257 ) );
  XOR \SUBBYTES[0].a/U4185  ( .A(\SUBBYTES[0].a/n1259 ), .B(
        \SUBBYTES[0].a/n1258 ), .Z(\SUBBYTES[0].a/w1052 ) );
  XOR \SUBBYTES[0].a/U4184  ( .A(\w1[0][89] ), .B(\SUBBYTES[0].a/n1260 ), .Z(
        \SUBBYTES[0].a/n1258 ) );
  XOR \SUBBYTES[0].a/U4183  ( .A(\SUBBYTES[0].a/w1027 ), .B(
        \SUBBYTES[0].a/w1029 ), .Z(\SUBBYTES[0].a/n1259 ) );
  XOR \SUBBYTES[0].a/U4182  ( .A(\SUBBYTES[0].a/w1011 ), .B(
        \SUBBYTES[0].a/w1012 ), .Z(\SUBBYTES[0].a/n1260 ) );
  XOR \SUBBYTES[0].a/U4181  ( .A(\w1[0][97] ), .B(\SUBBYTES[0].a/n1261 ), .Z(
        \SUBBYTES[0].a/n1589 ) );
  XOR \SUBBYTES[0].a/U4180  ( .A(\w1[0][99] ), .B(\w1[0][98] ), .Z(
        \SUBBYTES[0].a/n1261 ) );
  XOR \SUBBYTES[0].a/U4179  ( .A(\w1[0][102] ), .B(\SUBBYTES[0].a/n1589 ), .Z(
        \SUBBYTES[0].a/w894 ) );
  XOR \SUBBYTES[0].a/U4178  ( .A(\w1[0][96] ), .B(\SUBBYTES[0].a/w894 ), .Z(
        \SUBBYTES[0].a/w781 ) );
  XOR \SUBBYTES[0].a/U4177  ( .A(\w1[0][96] ), .B(\SUBBYTES[0].a/n1262 ), .Z(
        \SUBBYTES[0].a/w782 ) );
  XOR \SUBBYTES[0].a/U4176  ( .A(\w1[0][102] ), .B(\w1[0][101] ), .Z(
        \SUBBYTES[0].a/n1262 ) );
  XOR \SUBBYTES[0].a/U4175  ( .A(\w1[0][101] ), .B(\SUBBYTES[0].a/n1589 ), .Z(
        \SUBBYTES[0].a/w912 ) );
  XOR \SUBBYTES[0].a/U4174  ( .A(\SUBBYTES[0].a/n1264 ), .B(
        \SUBBYTES[0].a/n1263 ), .Z(\SUBBYTES[0].a/w905 ) );
  XOR \SUBBYTES[0].a/U4173  ( .A(\w1[0][99] ), .B(\w1[0][97] ), .Z(
        \SUBBYTES[0].a/n1263 ) );
  XOR \SUBBYTES[0].a/U4172  ( .A(\w1[0][103] ), .B(\w1[0][100] ), .Z(
        \SUBBYTES[0].a/n1264 ) );
  XOR \SUBBYTES[0].a/U4171  ( .A(\w1[0][96] ), .B(\SUBBYTES[0].a/w905 ), .Z(
        \SUBBYTES[0].a/w784 ) );
  XOR \SUBBYTES[0].a/U4170  ( .A(\SUBBYTES[0].a/n1266 ), .B(
        \SUBBYTES[0].a/n1265 ), .Z(\SUBBYTES[0].a/w892 ) );
  XOR \SUBBYTES[0].a/U4169  ( .A(\SUBBYTES[0].a/w853 ), .B(n1156), .Z(
        \SUBBYTES[0].a/n1265 ) );
  XOR \SUBBYTES[0].a/U4168  ( .A(\SUBBYTES[0].a/w846 ), .B(
        \SUBBYTES[0].a/w849 ), .Z(\SUBBYTES[0].a/n1266 ) );
  XOR \SUBBYTES[0].a/U4167  ( .A(\SUBBYTES[0].a/n1268 ), .B(
        \SUBBYTES[0].a/n1267 ), .Z(\SUBBYTES[0].a/w893 ) );
  XOR \SUBBYTES[0].a/U4166  ( .A(\SUBBYTES[0].a/w853 ), .B(\SUBBYTES[0].a/n40 ), .Z(\SUBBYTES[0].a/n1267 ) );
  XOR \SUBBYTES[0].a/U4165  ( .A(\SUBBYTES[0].a/w846 ), .B(\SUBBYTES[0].a/n39 ), .Z(\SUBBYTES[0].a/n1268 ) );
  XOR \SUBBYTES[0].a/U4164  ( .A(\SUBBYTES[0].a/w905 ), .B(
        \SUBBYTES[0].a/n1269 ), .Z(\SUBBYTES[0].a/w895 ) );
  XOR \SUBBYTES[0].a/U4163  ( .A(\w1[0][102] ), .B(\w1[0][101] ), .Z(
        \SUBBYTES[0].a/n1269 ) );
  XOR \SUBBYTES[0].a/U4162  ( .A(\SUBBYTES[0].a/n1271 ), .B(
        \SUBBYTES[0].a/n1270 ), .Z(\SUBBYTES[0].a/w896 ) );
  XOR \SUBBYTES[0].a/U4161  ( .A(\SUBBYTES[0].a/n40 ), .B(n1156), .Z(
        \SUBBYTES[0].a/n1270 ) );
  XOR \SUBBYTES[0].a/U4160  ( .A(\SUBBYTES[0].a/n39 ), .B(\SUBBYTES[0].a/w849 ), .Z(\SUBBYTES[0].a/n1271 ) );
  XOR \SUBBYTES[0].a/U4159  ( .A(\w1[0][103] ), .B(\w1[0][98] ), .Z(
        \SUBBYTES[0].a/n1595 ) );
  XOR \SUBBYTES[0].a/U4158  ( .A(\SUBBYTES[0].a/n1595 ), .B(
        \SUBBYTES[0].a/n1272 ), .Z(\SUBBYTES[0].a/w897 ) );
  XOR \SUBBYTES[0].a/U4157  ( .A(\w1[0][101] ), .B(\w1[0][100] ), .Z(
        \SUBBYTES[0].a/n1272 ) );
  XOR \SUBBYTES[0].a/U4156  ( .A(\w1[0][103] ), .B(\SUBBYTES[0].a/w782 ), .Z(
        \SUBBYTES[0].a/w785 ) );
  XOR \SUBBYTES[0].a/U4155  ( .A(\w1[0][97] ), .B(\SUBBYTES[0].a/w782 ), .Z(
        \SUBBYTES[0].a/w786 ) );
  XOR \SUBBYTES[0].a/U4154  ( .A(\w1[0][100] ), .B(\SUBBYTES[0].a/w782 ), .Z(
        \SUBBYTES[0].a/w787 ) );
  XOR \SUBBYTES[0].a/U4153  ( .A(\SUBBYTES[0].a/w786 ), .B(
        \SUBBYTES[0].a/n1595 ), .Z(\SUBBYTES[0].a/w788 ) );
  XOR \SUBBYTES[0].a/U4152  ( .A(\SUBBYTES[0].a/n1595 ), .B(
        \SUBBYTES[0].a/n1273 ), .Z(\SUBBYTES[0].a/w873 ) );
  XOR \SUBBYTES[0].a/U4151  ( .A(\w1[0][100] ), .B(\w1[0][97] ), .Z(
        \SUBBYTES[0].a/n1273 ) );
  XOR \SUBBYTES[0].a/U4150  ( .A(\SUBBYTES[0].a/n1275 ), .B(
        \SUBBYTES[0].a/n1274 ), .Z(\SUBBYTES[0].a/n1592 ) );
  XOR \SUBBYTES[0].a/U4149  ( .A(\w1[0][100] ), .B(\SUBBYTES[0].a/n1276 ), .Z(
        \SUBBYTES[0].a/n1274 ) );
  XOR \SUBBYTES[0].a/U4148  ( .A(\SUBBYTES[0].a/w838 ), .B(\w1[0][102] ), .Z(
        \SUBBYTES[0].a/n1275 ) );
  XOR \SUBBYTES[0].a/U4147  ( .A(\SUBBYTES[0].a/w812 ), .B(
        \SUBBYTES[0].a/w819 ), .Z(\SUBBYTES[0].a/n1276 ) );
  XOR \SUBBYTES[0].a/U4146  ( .A(\SUBBYTES[0].a/n1278 ), .B(
        \SUBBYTES[0].a/n1277 ), .Z(\SUBBYTES[0].a/n1590 ) );
  XOR \SUBBYTES[0].a/U4145  ( .A(\w1[0][97] ), .B(\SUBBYTES[0].a/n1279 ), .Z(
        \SUBBYTES[0].a/n1277 ) );
  XOR \SUBBYTES[0].a/U4144  ( .A(\SUBBYTES[0].a/w837 ), .B(\w1[0][101] ), .Z(
        \SUBBYTES[0].a/n1278 ) );
  XOR \SUBBYTES[0].a/U4143  ( .A(\SUBBYTES[0].a/w813 ), .B(
        \SUBBYTES[0].a/w820 ), .Z(\SUBBYTES[0].a/n1279 ) );
  XOR \SUBBYTES[0].a/U4142  ( .A(\SUBBYTES[0].a/n1592 ), .B(
        \SUBBYTES[0].a/n1590 ), .Z(\SUBBYTES[0].a/w843 ) );
  XOR \SUBBYTES[0].a/U4141  ( .A(\w1[0][101] ), .B(\SUBBYTES[0].a/n1280 ), .Z(
        \SUBBYTES[0].a/n1593 ) );
  XOR \SUBBYTES[0].a/U4140  ( .A(\SUBBYTES[0].a/w805 ), .B(
        \SUBBYTES[0].a/w815 ), .Z(\SUBBYTES[0].a/n1280 ) );
  XOR \SUBBYTES[0].a/U4139  ( .A(\SUBBYTES[0].a/n1282 ), .B(
        \SUBBYTES[0].a/n1281 ), .Z(\SUBBYTES[0].a/w830 ) );
  XOR \SUBBYTES[0].a/U4138  ( .A(\SUBBYTES[0].a/n1593 ), .B(
        \SUBBYTES[0].a/n1283 ), .Z(\SUBBYTES[0].a/n1281 ) );
  XOR \SUBBYTES[0].a/U4137  ( .A(\w1[0][100] ), .B(\SUBBYTES[0].a/w894 ), .Z(
        \SUBBYTES[0].a/n1282 ) );
  XOR \SUBBYTES[0].a/U4136  ( .A(\SUBBYTES[0].a/w807 ), .B(
        \SUBBYTES[0].a/w812 ), .Z(\SUBBYTES[0].a/n1283 ) );
  XOR \SUBBYTES[0].a/U4135  ( .A(\SUBBYTES[0].a/n1285 ), .B(
        \SUBBYTES[0].a/n1284 ), .Z(\SUBBYTES[0].a/n1591 ) );
  XOR \SUBBYTES[0].a/U4134  ( .A(\SUBBYTES[0].a/w840 ), .B(\w1[0][103] ), .Z(
        \SUBBYTES[0].a/n1284 ) );
  XOR \SUBBYTES[0].a/U4133  ( .A(\SUBBYTES[0].a/w815 ), .B(
        \SUBBYTES[0].a/w822 ), .Z(\SUBBYTES[0].a/n1285 ) );
  XOR \SUBBYTES[0].a/U4132  ( .A(\SUBBYTES[0].a/n1590 ), .B(
        \SUBBYTES[0].a/n1591 ), .Z(\SUBBYTES[0].a/w842 ) );
  XOR \SUBBYTES[0].a/U4131  ( .A(\w1[0][99] ), .B(\SUBBYTES[0].a/n1286 ), .Z(
        \SUBBYTES[0].a/n1594 ) );
  XOR \SUBBYTES[0].a/U4130  ( .A(\SUBBYTES[0].a/w804 ), .B(
        \SUBBYTES[0].a/w807 ), .Z(\SUBBYTES[0].a/n1286 ) );
  XOR \SUBBYTES[0].a/U4129  ( .A(\SUBBYTES[0].a/n1288 ), .B(
        \SUBBYTES[0].a/n1287 ), .Z(\SUBBYTES[0].a/w831 ) );
  XOR \SUBBYTES[0].a/U4128  ( .A(\SUBBYTES[0].a/n1594 ), .B(
        \SUBBYTES[0].a/n1289 ), .Z(\SUBBYTES[0].a/n1287 ) );
  XOR \SUBBYTES[0].a/U4127  ( .A(\w1[0][102] ), .B(\SUBBYTES[0].a/w873 ), .Z(
        \SUBBYTES[0].a/n1288 ) );
  XOR \SUBBYTES[0].a/U4126  ( .A(\SUBBYTES[0].a/w812 ), .B(
        \SUBBYTES[0].a/w813 ), .Z(\SUBBYTES[0].a/n1289 ) );
  XOR \SUBBYTES[0].a/U4125  ( .A(\SUBBYTES[0].a/n1592 ), .B(
        \SUBBYTES[0].a/n1591 ), .Z(\SUBBYTES[0].a/w851 ) );
  XOR \SUBBYTES[0].a/U4124  ( .A(\SUBBYTES[0].a/n1291 ), .B(
        \SUBBYTES[0].a/n1290 ), .Z(\SUBBYTES[0].a/w852 ) );
  XOR \SUBBYTES[0].a/U4123  ( .A(\w1[0][103] ), .B(\SUBBYTES[0].a/n1593 ), .Z(
        \SUBBYTES[0].a/n1290 ) );
  XOR \SUBBYTES[0].a/U4122  ( .A(\SUBBYTES[0].a/w804 ), .B(
        \SUBBYTES[0].a/w813 ), .Z(\SUBBYTES[0].a/n1291 ) );
  XOR \SUBBYTES[0].a/U4121  ( .A(\SUBBYTES[0].a/n1293 ), .B(
        \SUBBYTES[0].a/n1292 ), .Z(\SUBBYTES[0].a/w828 ) );
  XOR \SUBBYTES[0].a/U4120  ( .A(\SUBBYTES[0].a/n1295 ), .B(
        \SUBBYTES[0].a/n1294 ), .Z(\SUBBYTES[0].a/n1292 ) );
  XOR \SUBBYTES[0].a/U4119  ( .A(\w1[0][103] ), .B(\SUBBYTES[0].a/w912 ), .Z(
        \SUBBYTES[0].a/n1293 ) );
  XOR \SUBBYTES[0].a/U4118  ( .A(\SUBBYTES[0].a/w819 ), .B(
        \SUBBYTES[0].a/w822 ), .Z(\SUBBYTES[0].a/n1294 ) );
  XOR \SUBBYTES[0].a/U4117  ( .A(\SUBBYTES[0].a/w805 ), .B(
        \SUBBYTES[0].a/w807 ), .Z(\SUBBYTES[0].a/n1295 ) );
  XOR \SUBBYTES[0].a/U4116  ( .A(\SUBBYTES[0].a/n1297 ), .B(
        \SUBBYTES[0].a/n1296 ), .Z(\SUBBYTES[0].a/w829 ) );
  XOR \SUBBYTES[0].a/U4115  ( .A(\SUBBYTES[0].a/n1594 ), .B(
        \SUBBYTES[0].a/n1298 ), .Z(\SUBBYTES[0].a/n1296 ) );
  XOR \SUBBYTES[0].a/U4114  ( .A(\w1[0][101] ), .B(\SUBBYTES[0].a/n1595 ), .Z(
        \SUBBYTES[0].a/n1297 ) );
  XOR \SUBBYTES[0].a/U4113  ( .A(\SUBBYTES[0].a/w819 ), .B(
        \SUBBYTES[0].a/w820 ), .Z(\SUBBYTES[0].a/n1298 ) );
  XOR \SUBBYTES[0].a/U4112  ( .A(\SUBBYTES[0].a/n1300 ), .B(
        \SUBBYTES[0].a/n1299 ), .Z(\SUBBYTES[0].a/w845 ) );
  XOR \SUBBYTES[0].a/U4111  ( .A(\w1[0][97] ), .B(\SUBBYTES[0].a/n1301 ), .Z(
        \SUBBYTES[0].a/n1299 ) );
  XOR \SUBBYTES[0].a/U4110  ( .A(\SUBBYTES[0].a/w820 ), .B(
        \SUBBYTES[0].a/w822 ), .Z(\SUBBYTES[0].a/n1300 ) );
  XOR \SUBBYTES[0].a/U4109  ( .A(\SUBBYTES[0].a/w804 ), .B(
        \SUBBYTES[0].a/w805 ), .Z(\SUBBYTES[0].a/n1301 ) );
  XOR \SUBBYTES[0].a/U4108  ( .A(\w1[0][105] ), .B(\SUBBYTES[0].a/n1302 ), .Z(
        \SUBBYTES[0].a/n1596 ) );
  XOR \SUBBYTES[0].a/U4107  ( .A(\w1[0][107] ), .B(\w1[0][106] ), .Z(
        \SUBBYTES[0].a/n1302 ) );
  XOR \SUBBYTES[0].a/U4106  ( .A(\w1[0][110] ), .B(\SUBBYTES[0].a/n1596 ), .Z(
        \SUBBYTES[0].a/w687 ) );
  XOR \SUBBYTES[0].a/U4105  ( .A(\w1[0][104] ), .B(\SUBBYTES[0].a/w687 ), .Z(
        \SUBBYTES[0].a/w574 ) );
  XOR \SUBBYTES[0].a/U4104  ( .A(\w1[0][104] ), .B(\SUBBYTES[0].a/n1303 ), .Z(
        \SUBBYTES[0].a/w575 ) );
  XOR \SUBBYTES[0].a/U4103  ( .A(\w1[0][110] ), .B(\w1[0][109] ), .Z(
        \SUBBYTES[0].a/n1303 ) );
  XOR \SUBBYTES[0].a/U4102  ( .A(\w1[0][109] ), .B(\SUBBYTES[0].a/n1596 ), .Z(
        \SUBBYTES[0].a/w705 ) );
  XOR \SUBBYTES[0].a/U4101  ( .A(\SUBBYTES[0].a/n1305 ), .B(
        \SUBBYTES[0].a/n1304 ), .Z(\SUBBYTES[0].a/w698 ) );
  XOR \SUBBYTES[0].a/U4100  ( .A(\w1[0][107] ), .B(\w1[0][105] ), .Z(
        \SUBBYTES[0].a/n1304 ) );
  XOR \SUBBYTES[0].a/U4099  ( .A(\w1[0][111] ), .B(\w1[0][108] ), .Z(
        \SUBBYTES[0].a/n1305 ) );
  XOR \SUBBYTES[0].a/U4098  ( .A(\w1[0][104] ), .B(\SUBBYTES[0].a/w698 ), .Z(
        \SUBBYTES[0].a/w577 ) );
  XOR \SUBBYTES[0].a/U4097  ( .A(\SUBBYTES[0].a/n1307 ), .B(
        \SUBBYTES[0].a/n1306 ), .Z(\SUBBYTES[0].a/w685 ) );
  XOR \SUBBYTES[0].a/U4096  ( .A(\SUBBYTES[0].a/w646 ), .B(n1155), .Z(
        \SUBBYTES[0].a/n1306 ) );
  XOR \SUBBYTES[0].a/U4095  ( .A(\SUBBYTES[0].a/w639 ), .B(
        \SUBBYTES[0].a/w642 ), .Z(\SUBBYTES[0].a/n1307 ) );
  XOR \SUBBYTES[0].a/U4094  ( .A(\SUBBYTES[0].a/n1309 ), .B(
        \SUBBYTES[0].a/n1308 ), .Z(\SUBBYTES[0].a/w686 ) );
  XOR \SUBBYTES[0].a/U4093  ( .A(\SUBBYTES[0].a/w646 ), .B(\SUBBYTES[0].a/n30 ), .Z(\SUBBYTES[0].a/n1308 ) );
  XOR \SUBBYTES[0].a/U4092  ( .A(\SUBBYTES[0].a/w639 ), .B(\SUBBYTES[0].a/n29 ), .Z(\SUBBYTES[0].a/n1309 ) );
  XOR \SUBBYTES[0].a/U4091  ( .A(\SUBBYTES[0].a/w698 ), .B(
        \SUBBYTES[0].a/n1310 ), .Z(\SUBBYTES[0].a/w688 ) );
  XOR \SUBBYTES[0].a/U4090  ( .A(\w1[0][110] ), .B(\w1[0][109] ), .Z(
        \SUBBYTES[0].a/n1310 ) );
  XOR \SUBBYTES[0].a/U4089  ( .A(\SUBBYTES[0].a/n1312 ), .B(
        \SUBBYTES[0].a/n1311 ), .Z(\SUBBYTES[0].a/w689 ) );
  XOR \SUBBYTES[0].a/U4088  ( .A(\SUBBYTES[0].a/n30 ), .B(n1155), .Z(
        \SUBBYTES[0].a/n1311 ) );
  XOR \SUBBYTES[0].a/U4087  ( .A(\SUBBYTES[0].a/n29 ), .B(\SUBBYTES[0].a/w642 ), .Z(\SUBBYTES[0].a/n1312 ) );
  XOR \SUBBYTES[0].a/U4086  ( .A(\w1[0][111] ), .B(\w1[0][106] ), .Z(
        \SUBBYTES[0].a/n1602 ) );
  XOR \SUBBYTES[0].a/U4085  ( .A(\SUBBYTES[0].a/n1602 ), .B(
        \SUBBYTES[0].a/n1313 ), .Z(\SUBBYTES[0].a/w690 ) );
  XOR \SUBBYTES[0].a/U4084  ( .A(\w1[0][109] ), .B(\w1[0][108] ), .Z(
        \SUBBYTES[0].a/n1313 ) );
  XOR \SUBBYTES[0].a/U4083  ( .A(\w1[0][111] ), .B(\SUBBYTES[0].a/w575 ), .Z(
        \SUBBYTES[0].a/w578 ) );
  XOR \SUBBYTES[0].a/U4082  ( .A(\w1[0][105] ), .B(\SUBBYTES[0].a/w575 ), .Z(
        \SUBBYTES[0].a/w579 ) );
  XOR \SUBBYTES[0].a/U4081  ( .A(\w1[0][108] ), .B(\SUBBYTES[0].a/w575 ), .Z(
        \SUBBYTES[0].a/w580 ) );
  XOR \SUBBYTES[0].a/U4080  ( .A(\SUBBYTES[0].a/w579 ), .B(
        \SUBBYTES[0].a/n1602 ), .Z(\SUBBYTES[0].a/w581 ) );
  XOR \SUBBYTES[0].a/U4079  ( .A(\SUBBYTES[0].a/n1602 ), .B(
        \SUBBYTES[0].a/n1314 ), .Z(\SUBBYTES[0].a/w666 ) );
  XOR \SUBBYTES[0].a/U4078  ( .A(\w1[0][108] ), .B(\w1[0][105] ), .Z(
        \SUBBYTES[0].a/n1314 ) );
  XOR \SUBBYTES[0].a/U4077  ( .A(\SUBBYTES[0].a/n1316 ), .B(
        \SUBBYTES[0].a/n1315 ), .Z(\SUBBYTES[0].a/n1599 ) );
  XOR \SUBBYTES[0].a/U4076  ( .A(\w1[0][108] ), .B(\SUBBYTES[0].a/n1317 ), .Z(
        \SUBBYTES[0].a/n1315 ) );
  XOR \SUBBYTES[0].a/U4075  ( .A(\SUBBYTES[0].a/w631 ), .B(\w1[0][110] ), .Z(
        \SUBBYTES[0].a/n1316 ) );
  XOR \SUBBYTES[0].a/U4074  ( .A(\SUBBYTES[0].a/w605 ), .B(
        \SUBBYTES[0].a/w612 ), .Z(\SUBBYTES[0].a/n1317 ) );
  XOR \SUBBYTES[0].a/U4073  ( .A(\SUBBYTES[0].a/n1319 ), .B(
        \SUBBYTES[0].a/n1318 ), .Z(\SUBBYTES[0].a/n1597 ) );
  XOR \SUBBYTES[0].a/U4072  ( .A(\w1[0][105] ), .B(\SUBBYTES[0].a/n1320 ), .Z(
        \SUBBYTES[0].a/n1318 ) );
  XOR \SUBBYTES[0].a/U4071  ( .A(\SUBBYTES[0].a/w630 ), .B(\w1[0][109] ), .Z(
        \SUBBYTES[0].a/n1319 ) );
  XOR \SUBBYTES[0].a/U4070  ( .A(\SUBBYTES[0].a/w606 ), .B(
        \SUBBYTES[0].a/w613 ), .Z(\SUBBYTES[0].a/n1320 ) );
  XOR \SUBBYTES[0].a/U4069  ( .A(\SUBBYTES[0].a/n1599 ), .B(
        \SUBBYTES[0].a/n1597 ), .Z(\SUBBYTES[0].a/w636 ) );
  XOR \SUBBYTES[0].a/U4068  ( .A(\w1[0][109] ), .B(\SUBBYTES[0].a/n1321 ), .Z(
        \SUBBYTES[0].a/n1600 ) );
  XOR \SUBBYTES[0].a/U4067  ( .A(\SUBBYTES[0].a/w598 ), .B(
        \SUBBYTES[0].a/w608 ), .Z(\SUBBYTES[0].a/n1321 ) );
  XOR \SUBBYTES[0].a/U4066  ( .A(\SUBBYTES[0].a/n1323 ), .B(
        \SUBBYTES[0].a/n1322 ), .Z(\SUBBYTES[0].a/w623 ) );
  XOR \SUBBYTES[0].a/U4065  ( .A(\SUBBYTES[0].a/n1600 ), .B(
        \SUBBYTES[0].a/n1324 ), .Z(\SUBBYTES[0].a/n1322 ) );
  XOR \SUBBYTES[0].a/U4064  ( .A(\w1[0][108] ), .B(\SUBBYTES[0].a/w687 ), .Z(
        \SUBBYTES[0].a/n1323 ) );
  XOR \SUBBYTES[0].a/U4063  ( .A(\SUBBYTES[0].a/w600 ), .B(
        \SUBBYTES[0].a/w605 ), .Z(\SUBBYTES[0].a/n1324 ) );
  XOR \SUBBYTES[0].a/U4062  ( .A(\SUBBYTES[0].a/n1326 ), .B(
        \SUBBYTES[0].a/n1325 ), .Z(\SUBBYTES[0].a/n1598 ) );
  XOR \SUBBYTES[0].a/U4061  ( .A(\SUBBYTES[0].a/w633 ), .B(\w1[0][111] ), .Z(
        \SUBBYTES[0].a/n1325 ) );
  XOR \SUBBYTES[0].a/U4060  ( .A(\SUBBYTES[0].a/w608 ), .B(
        \SUBBYTES[0].a/w615 ), .Z(\SUBBYTES[0].a/n1326 ) );
  XOR \SUBBYTES[0].a/U4059  ( .A(\SUBBYTES[0].a/n1597 ), .B(
        \SUBBYTES[0].a/n1598 ), .Z(\SUBBYTES[0].a/w635 ) );
  XOR \SUBBYTES[0].a/U4058  ( .A(\w1[0][107] ), .B(\SUBBYTES[0].a/n1327 ), .Z(
        \SUBBYTES[0].a/n1601 ) );
  XOR \SUBBYTES[0].a/U4057  ( .A(\SUBBYTES[0].a/w597 ), .B(
        \SUBBYTES[0].a/w600 ), .Z(\SUBBYTES[0].a/n1327 ) );
  XOR \SUBBYTES[0].a/U4056  ( .A(\SUBBYTES[0].a/n1329 ), .B(
        \SUBBYTES[0].a/n1328 ), .Z(\SUBBYTES[0].a/w624 ) );
  XOR \SUBBYTES[0].a/U4055  ( .A(\SUBBYTES[0].a/n1601 ), .B(
        \SUBBYTES[0].a/n1330 ), .Z(\SUBBYTES[0].a/n1328 ) );
  XOR \SUBBYTES[0].a/U4054  ( .A(\w1[0][110] ), .B(\SUBBYTES[0].a/w666 ), .Z(
        \SUBBYTES[0].a/n1329 ) );
  XOR \SUBBYTES[0].a/U4053  ( .A(\SUBBYTES[0].a/w605 ), .B(
        \SUBBYTES[0].a/w606 ), .Z(\SUBBYTES[0].a/n1330 ) );
  XOR \SUBBYTES[0].a/U4052  ( .A(\SUBBYTES[0].a/n1599 ), .B(
        \SUBBYTES[0].a/n1598 ), .Z(\SUBBYTES[0].a/w644 ) );
  XOR \SUBBYTES[0].a/U4051  ( .A(\SUBBYTES[0].a/n1332 ), .B(
        \SUBBYTES[0].a/n1331 ), .Z(\SUBBYTES[0].a/w645 ) );
  XOR \SUBBYTES[0].a/U4050  ( .A(\w1[0][111] ), .B(\SUBBYTES[0].a/n1600 ), .Z(
        \SUBBYTES[0].a/n1331 ) );
  XOR \SUBBYTES[0].a/U4049  ( .A(\SUBBYTES[0].a/w597 ), .B(
        \SUBBYTES[0].a/w606 ), .Z(\SUBBYTES[0].a/n1332 ) );
  XOR \SUBBYTES[0].a/U4048  ( .A(\SUBBYTES[0].a/n1334 ), .B(
        \SUBBYTES[0].a/n1333 ), .Z(\SUBBYTES[0].a/w621 ) );
  XOR \SUBBYTES[0].a/U4047  ( .A(\SUBBYTES[0].a/n1336 ), .B(
        \SUBBYTES[0].a/n1335 ), .Z(\SUBBYTES[0].a/n1333 ) );
  XOR \SUBBYTES[0].a/U4046  ( .A(\w1[0][111] ), .B(\SUBBYTES[0].a/w705 ), .Z(
        \SUBBYTES[0].a/n1334 ) );
  XOR \SUBBYTES[0].a/U4045  ( .A(\SUBBYTES[0].a/w612 ), .B(
        \SUBBYTES[0].a/w615 ), .Z(\SUBBYTES[0].a/n1335 ) );
  XOR \SUBBYTES[0].a/U4044  ( .A(\SUBBYTES[0].a/w598 ), .B(
        \SUBBYTES[0].a/w600 ), .Z(\SUBBYTES[0].a/n1336 ) );
  XOR \SUBBYTES[0].a/U4043  ( .A(\SUBBYTES[0].a/n1338 ), .B(
        \SUBBYTES[0].a/n1337 ), .Z(\SUBBYTES[0].a/w622 ) );
  XOR \SUBBYTES[0].a/U4042  ( .A(\SUBBYTES[0].a/n1601 ), .B(
        \SUBBYTES[0].a/n1339 ), .Z(\SUBBYTES[0].a/n1337 ) );
  XOR \SUBBYTES[0].a/U4041  ( .A(\w1[0][109] ), .B(\SUBBYTES[0].a/n1602 ), .Z(
        \SUBBYTES[0].a/n1338 ) );
  XOR \SUBBYTES[0].a/U4040  ( .A(\SUBBYTES[0].a/w612 ), .B(
        \SUBBYTES[0].a/w613 ), .Z(\SUBBYTES[0].a/n1339 ) );
  XOR \SUBBYTES[0].a/U4039  ( .A(\SUBBYTES[0].a/n1341 ), .B(
        \SUBBYTES[0].a/n1340 ), .Z(\SUBBYTES[0].a/w638 ) );
  XOR \SUBBYTES[0].a/U4038  ( .A(\w1[0][105] ), .B(\SUBBYTES[0].a/n1342 ), .Z(
        \SUBBYTES[0].a/n1340 ) );
  XOR \SUBBYTES[0].a/U4037  ( .A(\SUBBYTES[0].a/w613 ), .B(
        \SUBBYTES[0].a/w615 ), .Z(\SUBBYTES[0].a/n1341 ) );
  XOR \SUBBYTES[0].a/U4036  ( .A(\SUBBYTES[0].a/w597 ), .B(
        \SUBBYTES[0].a/w598 ), .Z(\SUBBYTES[0].a/n1342 ) );
  XOR \SUBBYTES[0].a/U4035  ( .A(\w1[0][113] ), .B(\SUBBYTES[0].a/n1343 ), .Z(
        \SUBBYTES[0].a/n1603 ) );
  XOR \SUBBYTES[0].a/U4034  ( .A(\w1[0][115] ), .B(\w1[0][114] ), .Z(
        \SUBBYTES[0].a/n1343 ) );
  XOR \SUBBYTES[0].a/U4033  ( .A(\w1[0][118] ), .B(\SUBBYTES[0].a/n1603 ), .Z(
        \SUBBYTES[0].a/w480 ) );
  XOR \SUBBYTES[0].a/U4032  ( .A(\w1[0][112] ), .B(\SUBBYTES[0].a/w480 ), .Z(
        \SUBBYTES[0].a/w367 ) );
  XOR \SUBBYTES[0].a/U4031  ( .A(\w1[0][112] ), .B(\SUBBYTES[0].a/n1344 ), .Z(
        \SUBBYTES[0].a/w368 ) );
  XOR \SUBBYTES[0].a/U4030  ( .A(\w1[0][118] ), .B(\w1[0][117] ), .Z(
        \SUBBYTES[0].a/n1344 ) );
  XOR \SUBBYTES[0].a/U4029  ( .A(\w1[0][117] ), .B(\SUBBYTES[0].a/n1603 ), .Z(
        \SUBBYTES[0].a/w498 ) );
  XOR \SUBBYTES[0].a/U4028  ( .A(\SUBBYTES[0].a/n1346 ), .B(
        \SUBBYTES[0].a/n1345 ), .Z(\SUBBYTES[0].a/w491 ) );
  XOR \SUBBYTES[0].a/U4027  ( .A(\w1[0][115] ), .B(\w1[0][113] ), .Z(
        \SUBBYTES[0].a/n1345 ) );
  XOR \SUBBYTES[0].a/U4026  ( .A(\w1[0][119] ), .B(\w1[0][116] ), .Z(
        \SUBBYTES[0].a/n1346 ) );
  XOR \SUBBYTES[0].a/U4025  ( .A(\w1[0][112] ), .B(\SUBBYTES[0].a/w491 ), .Z(
        \SUBBYTES[0].a/w370 ) );
  XOR \SUBBYTES[0].a/U4024  ( .A(\SUBBYTES[0].a/n1348 ), .B(
        \SUBBYTES[0].a/n1347 ), .Z(\SUBBYTES[0].a/w478 ) );
  XOR \SUBBYTES[0].a/U4023  ( .A(\SUBBYTES[0].a/w439 ), .B(n1154), .Z(
        \SUBBYTES[0].a/n1347 ) );
  XOR \SUBBYTES[0].a/U4022  ( .A(\SUBBYTES[0].a/w432 ), .B(
        \SUBBYTES[0].a/w435 ), .Z(\SUBBYTES[0].a/n1348 ) );
  XOR \SUBBYTES[0].a/U4021  ( .A(\SUBBYTES[0].a/n1350 ), .B(
        \SUBBYTES[0].a/n1349 ), .Z(\SUBBYTES[0].a/w479 ) );
  XOR \SUBBYTES[0].a/U4020  ( .A(\SUBBYTES[0].a/w439 ), .B(\SUBBYTES[0].a/n20 ), .Z(\SUBBYTES[0].a/n1349 ) );
  XOR \SUBBYTES[0].a/U4019  ( .A(\SUBBYTES[0].a/w432 ), .B(\SUBBYTES[0].a/n19 ), .Z(\SUBBYTES[0].a/n1350 ) );
  XOR \SUBBYTES[0].a/U4018  ( .A(\SUBBYTES[0].a/w491 ), .B(
        \SUBBYTES[0].a/n1351 ), .Z(\SUBBYTES[0].a/w481 ) );
  XOR \SUBBYTES[0].a/U4017  ( .A(\w1[0][118] ), .B(\w1[0][117] ), .Z(
        \SUBBYTES[0].a/n1351 ) );
  XOR \SUBBYTES[0].a/U4016  ( .A(\SUBBYTES[0].a/n1353 ), .B(
        \SUBBYTES[0].a/n1352 ), .Z(\SUBBYTES[0].a/w482 ) );
  XOR \SUBBYTES[0].a/U4015  ( .A(\SUBBYTES[0].a/n20 ), .B(n1154), .Z(
        \SUBBYTES[0].a/n1352 ) );
  XOR \SUBBYTES[0].a/U4014  ( .A(\SUBBYTES[0].a/n19 ), .B(\SUBBYTES[0].a/w435 ), .Z(\SUBBYTES[0].a/n1353 ) );
  XOR \SUBBYTES[0].a/U4013  ( .A(\w1[0][119] ), .B(\w1[0][114] ), .Z(
        \SUBBYTES[0].a/n1609 ) );
  XOR \SUBBYTES[0].a/U4012  ( .A(\SUBBYTES[0].a/n1609 ), .B(
        \SUBBYTES[0].a/n1354 ), .Z(\SUBBYTES[0].a/w483 ) );
  XOR \SUBBYTES[0].a/U4011  ( .A(\w1[0][117] ), .B(\w1[0][116] ), .Z(
        \SUBBYTES[0].a/n1354 ) );
  XOR \SUBBYTES[0].a/U4010  ( .A(\w1[0][119] ), .B(\SUBBYTES[0].a/w368 ), .Z(
        \SUBBYTES[0].a/w371 ) );
  XOR \SUBBYTES[0].a/U4009  ( .A(\w1[0][113] ), .B(\SUBBYTES[0].a/w368 ), .Z(
        \SUBBYTES[0].a/w372 ) );
  XOR \SUBBYTES[0].a/U4008  ( .A(\w1[0][116] ), .B(\SUBBYTES[0].a/w368 ), .Z(
        \SUBBYTES[0].a/w373 ) );
  XOR \SUBBYTES[0].a/U4007  ( .A(\SUBBYTES[0].a/w372 ), .B(
        \SUBBYTES[0].a/n1609 ), .Z(\SUBBYTES[0].a/w374 ) );
  XOR \SUBBYTES[0].a/U4006  ( .A(\SUBBYTES[0].a/n1609 ), .B(
        \SUBBYTES[0].a/n1355 ), .Z(\SUBBYTES[0].a/w459 ) );
  XOR \SUBBYTES[0].a/U4005  ( .A(\w1[0][116] ), .B(\w1[0][113] ), .Z(
        \SUBBYTES[0].a/n1355 ) );
  XOR \SUBBYTES[0].a/U4004  ( .A(\SUBBYTES[0].a/n1357 ), .B(
        \SUBBYTES[0].a/n1356 ), .Z(\SUBBYTES[0].a/n1606 ) );
  XOR \SUBBYTES[0].a/U4003  ( .A(\w1[0][116] ), .B(\SUBBYTES[0].a/n1358 ), .Z(
        \SUBBYTES[0].a/n1356 ) );
  XOR \SUBBYTES[0].a/U4002  ( .A(\SUBBYTES[0].a/w424 ), .B(\w1[0][118] ), .Z(
        \SUBBYTES[0].a/n1357 ) );
  XOR \SUBBYTES[0].a/U4001  ( .A(\SUBBYTES[0].a/w398 ), .B(
        \SUBBYTES[0].a/w405 ), .Z(\SUBBYTES[0].a/n1358 ) );
  XOR \SUBBYTES[0].a/U4000  ( .A(\SUBBYTES[0].a/n1360 ), .B(
        \SUBBYTES[0].a/n1359 ), .Z(\SUBBYTES[0].a/n1604 ) );
  XOR \SUBBYTES[0].a/U3999  ( .A(\w1[0][113] ), .B(\SUBBYTES[0].a/n1361 ), .Z(
        \SUBBYTES[0].a/n1359 ) );
  XOR \SUBBYTES[0].a/U3998  ( .A(\SUBBYTES[0].a/w423 ), .B(\w1[0][117] ), .Z(
        \SUBBYTES[0].a/n1360 ) );
  XOR \SUBBYTES[0].a/U3997  ( .A(\SUBBYTES[0].a/w399 ), .B(
        \SUBBYTES[0].a/w406 ), .Z(\SUBBYTES[0].a/n1361 ) );
  XOR \SUBBYTES[0].a/U3996  ( .A(\SUBBYTES[0].a/n1606 ), .B(
        \SUBBYTES[0].a/n1604 ), .Z(\SUBBYTES[0].a/w429 ) );
  XOR \SUBBYTES[0].a/U3995  ( .A(\w1[0][117] ), .B(\SUBBYTES[0].a/n1362 ), .Z(
        \SUBBYTES[0].a/n1607 ) );
  XOR \SUBBYTES[0].a/U3994  ( .A(\SUBBYTES[0].a/w391 ), .B(
        \SUBBYTES[0].a/w401 ), .Z(\SUBBYTES[0].a/n1362 ) );
  XOR \SUBBYTES[0].a/U3993  ( .A(\SUBBYTES[0].a/n1364 ), .B(
        \SUBBYTES[0].a/n1363 ), .Z(\SUBBYTES[0].a/w416 ) );
  XOR \SUBBYTES[0].a/U3992  ( .A(\SUBBYTES[0].a/n1607 ), .B(
        \SUBBYTES[0].a/n1365 ), .Z(\SUBBYTES[0].a/n1363 ) );
  XOR \SUBBYTES[0].a/U3991  ( .A(\w1[0][116] ), .B(\SUBBYTES[0].a/w480 ), .Z(
        \SUBBYTES[0].a/n1364 ) );
  XOR \SUBBYTES[0].a/U3990  ( .A(\SUBBYTES[0].a/w393 ), .B(
        \SUBBYTES[0].a/w398 ), .Z(\SUBBYTES[0].a/n1365 ) );
  XOR \SUBBYTES[0].a/U3989  ( .A(\SUBBYTES[0].a/n1367 ), .B(
        \SUBBYTES[0].a/n1366 ), .Z(\SUBBYTES[0].a/n1605 ) );
  XOR \SUBBYTES[0].a/U3988  ( .A(\SUBBYTES[0].a/w426 ), .B(\w1[0][119] ), .Z(
        \SUBBYTES[0].a/n1366 ) );
  XOR \SUBBYTES[0].a/U3987  ( .A(\SUBBYTES[0].a/w401 ), .B(
        \SUBBYTES[0].a/w408 ), .Z(\SUBBYTES[0].a/n1367 ) );
  XOR \SUBBYTES[0].a/U3986  ( .A(\SUBBYTES[0].a/n1604 ), .B(
        \SUBBYTES[0].a/n1605 ), .Z(\SUBBYTES[0].a/w428 ) );
  XOR \SUBBYTES[0].a/U3985  ( .A(\w1[0][115] ), .B(\SUBBYTES[0].a/n1368 ), .Z(
        \SUBBYTES[0].a/n1608 ) );
  XOR \SUBBYTES[0].a/U3984  ( .A(\SUBBYTES[0].a/w390 ), .B(
        \SUBBYTES[0].a/w393 ), .Z(\SUBBYTES[0].a/n1368 ) );
  XOR \SUBBYTES[0].a/U3983  ( .A(\SUBBYTES[0].a/n1370 ), .B(
        \SUBBYTES[0].a/n1369 ), .Z(\SUBBYTES[0].a/w417 ) );
  XOR \SUBBYTES[0].a/U3982  ( .A(\SUBBYTES[0].a/n1608 ), .B(
        \SUBBYTES[0].a/n1371 ), .Z(\SUBBYTES[0].a/n1369 ) );
  XOR \SUBBYTES[0].a/U3981  ( .A(\w1[0][118] ), .B(\SUBBYTES[0].a/w459 ), .Z(
        \SUBBYTES[0].a/n1370 ) );
  XOR \SUBBYTES[0].a/U3980  ( .A(\SUBBYTES[0].a/w398 ), .B(
        \SUBBYTES[0].a/w399 ), .Z(\SUBBYTES[0].a/n1371 ) );
  XOR \SUBBYTES[0].a/U3979  ( .A(\SUBBYTES[0].a/n1606 ), .B(
        \SUBBYTES[0].a/n1605 ), .Z(\SUBBYTES[0].a/w437 ) );
  XOR \SUBBYTES[0].a/U3978  ( .A(\SUBBYTES[0].a/n1373 ), .B(
        \SUBBYTES[0].a/n1372 ), .Z(\SUBBYTES[0].a/w438 ) );
  XOR \SUBBYTES[0].a/U3977  ( .A(\w1[0][119] ), .B(\SUBBYTES[0].a/n1607 ), .Z(
        \SUBBYTES[0].a/n1372 ) );
  XOR \SUBBYTES[0].a/U3976  ( .A(\SUBBYTES[0].a/w390 ), .B(
        \SUBBYTES[0].a/w399 ), .Z(\SUBBYTES[0].a/n1373 ) );
  XOR \SUBBYTES[0].a/U3975  ( .A(\SUBBYTES[0].a/n1375 ), .B(
        \SUBBYTES[0].a/n1374 ), .Z(\SUBBYTES[0].a/w414 ) );
  XOR \SUBBYTES[0].a/U3974  ( .A(\SUBBYTES[0].a/n1377 ), .B(
        \SUBBYTES[0].a/n1376 ), .Z(\SUBBYTES[0].a/n1374 ) );
  XOR \SUBBYTES[0].a/U3973  ( .A(\w1[0][119] ), .B(\SUBBYTES[0].a/w498 ), .Z(
        \SUBBYTES[0].a/n1375 ) );
  XOR \SUBBYTES[0].a/U3972  ( .A(\SUBBYTES[0].a/w405 ), .B(
        \SUBBYTES[0].a/w408 ), .Z(\SUBBYTES[0].a/n1376 ) );
  XOR \SUBBYTES[0].a/U3971  ( .A(\SUBBYTES[0].a/w391 ), .B(
        \SUBBYTES[0].a/w393 ), .Z(\SUBBYTES[0].a/n1377 ) );
  XOR \SUBBYTES[0].a/U3970  ( .A(\SUBBYTES[0].a/n1379 ), .B(
        \SUBBYTES[0].a/n1378 ), .Z(\SUBBYTES[0].a/w415 ) );
  XOR \SUBBYTES[0].a/U3969  ( .A(\SUBBYTES[0].a/n1608 ), .B(
        \SUBBYTES[0].a/n1380 ), .Z(\SUBBYTES[0].a/n1378 ) );
  XOR \SUBBYTES[0].a/U3968  ( .A(\w1[0][117] ), .B(\SUBBYTES[0].a/n1609 ), .Z(
        \SUBBYTES[0].a/n1379 ) );
  XOR \SUBBYTES[0].a/U3967  ( .A(\SUBBYTES[0].a/w405 ), .B(
        \SUBBYTES[0].a/w406 ), .Z(\SUBBYTES[0].a/n1380 ) );
  XOR \SUBBYTES[0].a/U3966  ( .A(\SUBBYTES[0].a/n1382 ), .B(
        \SUBBYTES[0].a/n1381 ), .Z(\SUBBYTES[0].a/w431 ) );
  XOR \SUBBYTES[0].a/U3965  ( .A(\w1[0][113] ), .B(\SUBBYTES[0].a/n1383 ), .Z(
        \SUBBYTES[0].a/n1381 ) );
  XOR \SUBBYTES[0].a/U3964  ( .A(\SUBBYTES[0].a/w406 ), .B(
        \SUBBYTES[0].a/w408 ), .Z(\SUBBYTES[0].a/n1382 ) );
  XOR \SUBBYTES[0].a/U3963  ( .A(\SUBBYTES[0].a/w390 ), .B(
        \SUBBYTES[0].a/w391 ), .Z(\SUBBYTES[0].a/n1383 ) );
  XOR \SUBBYTES[0].a/U3962  ( .A(\w1[0][121] ), .B(\SUBBYTES[0].a/n1384 ), .Z(
        \SUBBYTES[0].a/n1610 ) );
  XOR \SUBBYTES[0].a/U3961  ( .A(\w1[0][123] ), .B(\w1[0][122] ), .Z(
        \SUBBYTES[0].a/n1384 ) );
  XOR \SUBBYTES[0].a/U3960  ( .A(\w1[0][126] ), .B(\SUBBYTES[0].a/n1610 ), .Z(
        \SUBBYTES[0].a/w273 ) );
  XOR \SUBBYTES[0].a/U3959  ( .A(\w1[0][120] ), .B(\SUBBYTES[0].a/w273 ), .Z(
        \SUBBYTES[0].a/w160 ) );
  XOR \SUBBYTES[0].a/U3958  ( .A(\w1[0][120] ), .B(\SUBBYTES[0].a/n1385 ), .Z(
        \SUBBYTES[0].a/w161 ) );
  XOR \SUBBYTES[0].a/U3957  ( .A(\w1[0][126] ), .B(\w1[0][125] ), .Z(
        \SUBBYTES[0].a/n1385 ) );
  XOR \SUBBYTES[0].a/U3956  ( .A(\w1[0][125] ), .B(\SUBBYTES[0].a/n1610 ), .Z(
        \SUBBYTES[0].a/w291 ) );
  XOR \SUBBYTES[0].a/U3955  ( .A(\SUBBYTES[0].a/n1387 ), .B(
        \SUBBYTES[0].a/n1386 ), .Z(\SUBBYTES[0].a/w284 ) );
  XOR \SUBBYTES[0].a/U3954  ( .A(\w1[0][123] ), .B(\w1[0][121] ), .Z(
        \SUBBYTES[0].a/n1386 ) );
  XOR \SUBBYTES[0].a/U3953  ( .A(\w1[0][127] ), .B(\w1[0][124] ), .Z(
        \SUBBYTES[0].a/n1387 ) );
  XOR \SUBBYTES[0].a/U3952  ( .A(\w1[0][120] ), .B(\SUBBYTES[0].a/w284 ), .Z(
        \SUBBYTES[0].a/w163 ) );
  XOR \SUBBYTES[0].a/U3951  ( .A(\SUBBYTES[0].a/n1389 ), .B(
        \SUBBYTES[0].a/n1388 ), .Z(\SUBBYTES[0].a/w271 ) );
  XOR \SUBBYTES[0].a/U3950  ( .A(\SUBBYTES[0].a/w232 ), .B(n1153), .Z(
        \SUBBYTES[0].a/n1388 ) );
  XOR \SUBBYTES[0].a/U3949  ( .A(\SUBBYTES[0].a/w225 ), .B(
        \SUBBYTES[0].a/w228 ), .Z(\SUBBYTES[0].a/n1389 ) );
  XOR \SUBBYTES[0].a/U3948  ( .A(\SUBBYTES[0].a/n1391 ), .B(
        \SUBBYTES[0].a/n1390 ), .Z(\SUBBYTES[0].a/w272 ) );
  XOR \SUBBYTES[0].a/U3947  ( .A(\SUBBYTES[0].a/w232 ), .B(\SUBBYTES[0].a/n10 ), .Z(\SUBBYTES[0].a/n1390 ) );
  XOR \SUBBYTES[0].a/U3946  ( .A(\SUBBYTES[0].a/w225 ), .B(\SUBBYTES[0].a/n9 ), 
        .Z(\SUBBYTES[0].a/n1391 ) );
  XOR \SUBBYTES[0].a/U3945  ( .A(\SUBBYTES[0].a/w284 ), .B(
        \SUBBYTES[0].a/n1392 ), .Z(\SUBBYTES[0].a/w274 ) );
  XOR \SUBBYTES[0].a/U3944  ( .A(\w1[0][126] ), .B(\w1[0][125] ), .Z(
        \SUBBYTES[0].a/n1392 ) );
  XOR \SUBBYTES[0].a/U3943  ( .A(\SUBBYTES[0].a/n1394 ), .B(
        \SUBBYTES[0].a/n1393 ), .Z(\SUBBYTES[0].a/w275 ) );
  XOR \SUBBYTES[0].a/U3942  ( .A(\SUBBYTES[0].a/n10 ), .B(n1153), .Z(
        \SUBBYTES[0].a/n1393 ) );
  XOR \SUBBYTES[0].a/U3941  ( .A(\SUBBYTES[0].a/n9 ), .B(\SUBBYTES[0].a/w228 ), 
        .Z(\SUBBYTES[0].a/n1394 ) );
  XOR \SUBBYTES[0].a/U3940  ( .A(\w1[0][127] ), .B(\w1[0][122] ), .Z(
        \SUBBYTES[0].a/n1616 ) );
  XOR \SUBBYTES[0].a/U3939  ( .A(\SUBBYTES[0].a/n1616 ), .B(
        \SUBBYTES[0].a/n1395 ), .Z(\SUBBYTES[0].a/w276 ) );
  XOR \SUBBYTES[0].a/U3938  ( .A(\w1[0][125] ), .B(\w1[0][124] ), .Z(
        \SUBBYTES[0].a/n1395 ) );
  XOR \SUBBYTES[0].a/U3937  ( .A(\w1[0][127] ), .B(\SUBBYTES[0].a/w161 ), .Z(
        \SUBBYTES[0].a/w164 ) );
  XOR \SUBBYTES[0].a/U3936  ( .A(\w1[0][121] ), .B(\SUBBYTES[0].a/w161 ), .Z(
        \SUBBYTES[0].a/w165 ) );
  XOR \SUBBYTES[0].a/U3935  ( .A(\w1[0][124] ), .B(\SUBBYTES[0].a/w161 ), .Z(
        \SUBBYTES[0].a/w166 ) );
  XOR \SUBBYTES[0].a/U3934  ( .A(\SUBBYTES[0].a/w165 ), .B(
        \SUBBYTES[0].a/n1616 ), .Z(\SUBBYTES[0].a/w167 ) );
  XOR \SUBBYTES[0].a/U3933  ( .A(\SUBBYTES[0].a/n1616 ), .B(
        \SUBBYTES[0].a/n1396 ), .Z(\SUBBYTES[0].a/w252 ) );
  XOR \SUBBYTES[0].a/U3932  ( .A(\w1[0][124] ), .B(\w1[0][121] ), .Z(
        \SUBBYTES[0].a/n1396 ) );
  XOR \SUBBYTES[0].a/U3931  ( .A(\SUBBYTES[0].a/n1398 ), .B(
        \SUBBYTES[0].a/n1397 ), .Z(\SUBBYTES[0].a/n1613 ) );
  XOR \SUBBYTES[0].a/U3930  ( .A(\w1[0][124] ), .B(\SUBBYTES[0].a/n1399 ), .Z(
        \SUBBYTES[0].a/n1397 ) );
  XOR \SUBBYTES[0].a/U3929  ( .A(\SUBBYTES[0].a/w217 ), .B(\w1[0][126] ), .Z(
        \SUBBYTES[0].a/n1398 ) );
  XOR \SUBBYTES[0].a/U3928  ( .A(\SUBBYTES[0].a/w191 ), .B(
        \SUBBYTES[0].a/w198 ), .Z(\SUBBYTES[0].a/n1399 ) );
  XOR \SUBBYTES[0].a/U3927  ( .A(\SUBBYTES[0].a/n1401 ), .B(
        \SUBBYTES[0].a/n1400 ), .Z(\SUBBYTES[0].a/n1611 ) );
  XOR \SUBBYTES[0].a/U3926  ( .A(\w1[0][121] ), .B(\SUBBYTES[0].a/n1402 ), .Z(
        \SUBBYTES[0].a/n1400 ) );
  XOR \SUBBYTES[0].a/U3925  ( .A(\SUBBYTES[0].a/w216 ), .B(\w1[0][125] ), .Z(
        \SUBBYTES[0].a/n1401 ) );
  XOR \SUBBYTES[0].a/U3924  ( .A(\SUBBYTES[0].a/w192 ), .B(
        \SUBBYTES[0].a/w199 ), .Z(\SUBBYTES[0].a/n1402 ) );
  XOR \SUBBYTES[0].a/U3923  ( .A(\SUBBYTES[0].a/n1613 ), .B(
        \SUBBYTES[0].a/n1611 ), .Z(\SUBBYTES[0].a/w222 ) );
  XOR \SUBBYTES[0].a/U3922  ( .A(\w1[0][125] ), .B(\SUBBYTES[0].a/n1403 ), .Z(
        \SUBBYTES[0].a/n1614 ) );
  XOR \SUBBYTES[0].a/U3921  ( .A(\SUBBYTES[0].a/w184 ), .B(
        \SUBBYTES[0].a/w194 ), .Z(\SUBBYTES[0].a/n1403 ) );
  XOR \SUBBYTES[0].a/U3920  ( .A(\SUBBYTES[0].a/n1405 ), .B(
        \SUBBYTES[0].a/n1404 ), .Z(\SUBBYTES[0].a/w209 ) );
  XOR \SUBBYTES[0].a/U3919  ( .A(\SUBBYTES[0].a/n1614 ), .B(
        \SUBBYTES[0].a/n1406 ), .Z(\SUBBYTES[0].a/n1404 ) );
  XOR \SUBBYTES[0].a/U3918  ( .A(\w1[0][124] ), .B(\SUBBYTES[0].a/w273 ), .Z(
        \SUBBYTES[0].a/n1405 ) );
  XOR \SUBBYTES[0].a/U3917  ( .A(\SUBBYTES[0].a/w186 ), .B(
        \SUBBYTES[0].a/w191 ), .Z(\SUBBYTES[0].a/n1406 ) );
  XOR \SUBBYTES[0].a/U3916  ( .A(\SUBBYTES[0].a/n1408 ), .B(
        \SUBBYTES[0].a/n1407 ), .Z(\SUBBYTES[0].a/n1612 ) );
  XOR \SUBBYTES[0].a/U3915  ( .A(\SUBBYTES[0].a/w219 ), .B(\w1[0][127] ), .Z(
        \SUBBYTES[0].a/n1407 ) );
  XOR \SUBBYTES[0].a/U3914  ( .A(\SUBBYTES[0].a/w194 ), .B(
        \SUBBYTES[0].a/w201 ), .Z(\SUBBYTES[0].a/n1408 ) );
  XOR \SUBBYTES[0].a/U3913  ( .A(\SUBBYTES[0].a/n1611 ), .B(
        \SUBBYTES[0].a/n1612 ), .Z(\SUBBYTES[0].a/w221 ) );
  XOR \SUBBYTES[0].a/U3912  ( .A(\w1[0][123] ), .B(\SUBBYTES[0].a/n1409 ), .Z(
        \SUBBYTES[0].a/n1615 ) );
  XOR \SUBBYTES[0].a/U3911  ( .A(\SUBBYTES[0].a/w183 ), .B(
        \SUBBYTES[0].a/w186 ), .Z(\SUBBYTES[0].a/n1409 ) );
  XOR \SUBBYTES[0].a/U3910  ( .A(\SUBBYTES[0].a/n1411 ), .B(
        \SUBBYTES[0].a/n1410 ), .Z(\SUBBYTES[0].a/w210 ) );
  XOR \SUBBYTES[0].a/U3909  ( .A(\SUBBYTES[0].a/n1615 ), .B(
        \SUBBYTES[0].a/n1412 ), .Z(\SUBBYTES[0].a/n1410 ) );
  XOR \SUBBYTES[0].a/U3908  ( .A(\w1[0][126] ), .B(\SUBBYTES[0].a/w252 ), .Z(
        \SUBBYTES[0].a/n1411 ) );
  XOR \SUBBYTES[0].a/U3907  ( .A(\SUBBYTES[0].a/w191 ), .B(
        \SUBBYTES[0].a/w192 ), .Z(\SUBBYTES[0].a/n1412 ) );
  XOR \SUBBYTES[0].a/U3906  ( .A(\SUBBYTES[0].a/n1613 ), .B(
        \SUBBYTES[0].a/n1612 ), .Z(\SUBBYTES[0].a/w230 ) );
  XOR \SUBBYTES[0].a/U3905  ( .A(\SUBBYTES[0].a/n1414 ), .B(
        \SUBBYTES[0].a/n1413 ), .Z(\SUBBYTES[0].a/w231 ) );
  XOR \SUBBYTES[0].a/U3904  ( .A(\w1[0][127] ), .B(\SUBBYTES[0].a/n1614 ), .Z(
        \SUBBYTES[0].a/n1413 ) );
  XOR \SUBBYTES[0].a/U3903  ( .A(\SUBBYTES[0].a/w183 ), .B(
        \SUBBYTES[0].a/w192 ), .Z(\SUBBYTES[0].a/n1414 ) );
  XOR \SUBBYTES[0].a/U3902  ( .A(\SUBBYTES[0].a/n1416 ), .B(
        \SUBBYTES[0].a/n1415 ), .Z(\SUBBYTES[0].a/w207 ) );
  XOR \SUBBYTES[0].a/U3901  ( .A(\SUBBYTES[0].a/n1418 ), .B(
        \SUBBYTES[0].a/n1417 ), .Z(\SUBBYTES[0].a/n1415 ) );
  XOR \SUBBYTES[0].a/U3900  ( .A(\w1[0][127] ), .B(\SUBBYTES[0].a/w291 ), .Z(
        \SUBBYTES[0].a/n1416 ) );
  XOR \SUBBYTES[0].a/U3899  ( .A(\SUBBYTES[0].a/w198 ), .B(
        \SUBBYTES[0].a/w201 ), .Z(\SUBBYTES[0].a/n1417 ) );
  XOR \SUBBYTES[0].a/U3898  ( .A(\SUBBYTES[0].a/w184 ), .B(
        \SUBBYTES[0].a/w186 ), .Z(\SUBBYTES[0].a/n1418 ) );
  XOR \SUBBYTES[0].a/U3897  ( .A(\SUBBYTES[0].a/n1420 ), .B(
        \SUBBYTES[0].a/n1419 ), .Z(\SUBBYTES[0].a/w208 ) );
  XOR \SUBBYTES[0].a/U3896  ( .A(\SUBBYTES[0].a/n1615 ), .B(
        \SUBBYTES[0].a/n1421 ), .Z(\SUBBYTES[0].a/n1419 ) );
  XOR \SUBBYTES[0].a/U3895  ( .A(\w1[0][125] ), .B(\SUBBYTES[0].a/n1616 ), .Z(
        \SUBBYTES[0].a/n1420 ) );
  XOR \SUBBYTES[0].a/U3894  ( .A(\SUBBYTES[0].a/w198 ), .B(
        \SUBBYTES[0].a/w199 ), .Z(\SUBBYTES[0].a/n1421 ) );
  XOR \SUBBYTES[0].a/U3893  ( .A(\SUBBYTES[0].a/n1423 ), .B(
        \SUBBYTES[0].a/n1422 ), .Z(\SUBBYTES[0].a/w224 ) );
  XOR \SUBBYTES[0].a/U3892  ( .A(\w1[0][121] ), .B(\SUBBYTES[0].a/n1424 ), .Z(
        \SUBBYTES[0].a/n1422 ) );
  XOR \SUBBYTES[0].a/U3891  ( .A(\SUBBYTES[0].a/w199 ), .B(
        \SUBBYTES[0].a/w201 ), .Z(\SUBBYTES[0].a/n1423 ) );
  XOR \SUBBYTES[0].a/U3890  ( .A(\SUBBYTES[0].a/w183 ), .B(
        \SUBBYTES[0].a/w184 ), .Z(\SUBBYTES[0].a/n1424 ) );
  XOR \MIXCOLUMNS[0].d/U432  ( .A(n1152), .B(n540), .Z(\MIXCOLUMNS[0].d/n250 )
         );
  XOR \MIXCOLUMNS[0].d/U431  ( .A(\MIXCOLUMNS[0].d/n2 ), .B(
        \MIXCOLUMNS[0].d/n1 ), .Z(\w0[1][0] ) );
  XOR \MIXCOLUMNS[0].d/U430  ( .A(n1151), .B(\MIXCOLUMNS[0].d/n250 ), .Z(
        \MIXCOLUMNS[0].d/n1 ) );
  XOR \MIXCOLUMNS[0].d/U429  ( .A(n1150), .B(n36), .Z(\MIXCOLUMNS[0].d/n2 ) );
  XOR \MIXCOLUMNS[0].d/U428  ( .A(n1150), .B(n539), .Z(\MIXCOLUMNS[0].d/n235 )
         );
  XOR \MIXCOLUMNS[0].d/U427  ( .A(\MIXCOLUMNS[0].d/n4 ), .B(
        \MIXCOLUMNS[0].d/n3 ), .Z(\w0[1][1] ) );
  XOR \MIXCOLUMNS[0].d/U426  ( .A(\w3[0][2] ), .B(\MIXCOLUMNS[0].d/n235 ), .Z(
        \MIXCOLUMNS[0].d/n3 ) );
  XOR \MIXCOLUMNS[0].d/U425  ( .A(\w3[0][26] ), .B(n538), .Z(
        \MIXCOLUMNS[0].d/n4 ) );
  XOR \MIXCOLUMNS[0].d/U424  ( .A(\w3[0][26] ), .B(\w3[0][18] ), .Z(
        \MIXCOLUMNS[0].d/n238 ) );
  XOR \MIXCOLUMNS[0].d/U423  ( .A(\MIXCOLUMNS[0].d/n6 ), .B(
        \MIXCOLUMNS[0].d/n5 ), .Z(\w0[1][2] ) );
  XOR \MIXCOLUMNS[0].d/U422  ( .A(n1149), .B(\MIXCOLUMNS[0].d/n238 ), .Z(
        \MIXCOLUMNS[0].d/n5 ) );
  XOR \MIXCOLUMNS[0].d/U421  ( .A(n1148), .B(\w3[0][10] ), .Z(
        \MIXCOLUMNS[0].d/n6 ) );
  XOR \MIXCOLUMNS[0].d/U420  ( .A(n1152), .B(n537), .Z(\MIXCOLUMNS[0].d/n233 )
         );
  XOR \MIXCOLUMNS[0].d/U419  ( .A(n1148), .B(n536), .Z(\MIXCOLUMNS[0].d/n240 )
         );
  XOR \MIXCOLUMNS[0].d/U418  ( .A(\MIXCOLUMNS[0].d/n8 ), .B(
        \MIXCOLUMNS[0].d/n7 ), .Z(\w0[1][3] ) );
  XOR \MIXCOLUMNS[0].d/U417  ( .A(\MIXCOLUMNS[0].d/n240 ), .B(
        \MIXCOLUMNS[0].d/n9 ), .Z(\MIXCOLUMNS[0].d/n7 ) );
  XOR \MIXCOLUMNS[0].d/U416  ( .A(n1147), .B(\MIXCOLUMNS[0].d/n233 ), .Z(
        \MIXCOLUMNS[0].d/n8 ) );
  XOR \MIXCOLUMNS[0].d/U415  ( .A(n1146), .B(n535), .Z(\MIXCOLUMNS[0].d/n9 )
         );
  XOR \MIXCOLUMNS[0].d/U414  ( .A(n1146), .B(n534), .Z(\MIXCOLUMNS[0].d/n242 )
         );
  XOR \MIXCOLUMNS[0].d/U413  ( .A(\MIXCOLUMNS[0].d/n11 ), .B(
        \MIXCOLUMNS[0].d/n10 ), .Z(\w0[1][4] ) );
  XOR \MIXCOLUMNS[0].d/U412  ( .A(\MIXCOLUMNS[0].d/n242 ), .B(
        \MIXCOLUMNS[0].d/n12 ), .Z(\MIXCOLUMNS[0].d/n10 ) );
  XOR \MIXCOLUMNS[0].d/U411  ( .A(n1145), .B(\MIXCOLUMNS[0].d/n233 ), .Z(
        \MIXCOLUMNS[0].d/n11 ) );
  XOR \MIXCOLUMNS[0].d/U410  ( .A(n1144), .B(n533), .Z(\MIXCOLUMNS[0].d/n12 )
         );
  XOR \MIXCOLUMNS[0].d/U409  ( .A(n1144), .B(n532), .Z(\MIXCOLUMNS[0].d/n244 )
         );
  XOR \MIXCOLUMNS[0].d/U408  ( .A(\MIXCOLUMNS[0].d/n14 ), .B(
        \MIXCOLUMNS[0].d/n13 ), .Z(\w0[1][5] ) );
  XOR \MIXCOLUMNS[0].d/U407  ( .A(n1143), .B(\MIXCOLUMNS[0].d/n244 ), .Z(
        \MIXCOLUMNS[0].d/n13 ) );
  XOR \MIXCOLUMNS[0].d/U406  ( .A(n1142), .B(n531), .Z(\MIXCOLUMNS[0].d/n14 )
         );
  XOR \MIXCOLUMNS[0].d/U405  ( .A(n1142), .B(n530), .Z(\MIXCOLUMNS[0].d/n246 )
         );
  XOR \MIXCOLUMNS[0].d/U404  ( .A(\MIXCOLUMNS[0].d/n16 ), .B(
        \MIXCOLUMNS[0].d/n15 ), .Z(\w0[1][6] ) );
  XOR \MIXCOLUMNS[0].d/U403  ( .A(\MIXCOLUMNS[0].d/n246 ), .B(
        \MIXCOLUMNS[0].d/n17 ), .Z(\MIXCOLUMNS[0].d/n15 ) );
  XOR \MIXCOLUMNS[0].d/U402  ( .A(n1141), .B(\MIXCOLUMNS[0].d/n233 ), .Z(
        \MIXCOLUMNS[0].d/n16 ) );
  XOR \MIXCOLUMNS[0].d/U401  ( .A(n1140), .B(n529), .Z(\MIXCOLUMNS[0].d/n17 )
         );
  XOR \MIXCOLUMNS[0].d/U400  ( .A(n1140), .B(n528), .Z(\MIXCOLUMNS[0].d/n248 )
         );
  XOR \MIXCOLUMNS[0].d/U399  ( .A(\MIXCOLUMNS[0].d/n248 ), .B(
        \MIXCOLUMNS[0].d/n18 ), .Z(\w0[1][7] ) );
  XOR \MIXCOLUMNS[0].d/U398  ( .A(n527), .B(\MIXCOLUMNS[0].d/n233 ), .Z(
        \MIXCOLUMNS[0].d/n18 ) );
  XOR \MIXCOLUMNS[0].d/U397  ( .A(n538), .B(n1151), .Z(\MIXCOLUMNS[0].d/n237 )
         );
  XOR \MIXCOLUMNS[0].d/U396  ( .A(\MIXCOLUMNS[0].d/n237 ), .B(
        \MIXCOLUMNS[0].d/n19 ), .Z(\w0[1][8] ) );
  XOR \MIXCOLUMNS[0].d/U395  ( .A(n537), .B(\MIXCOLUMNS[0].d/n250 ), .Z(
        \MIXCOLUMNS[0].d/n19 ) );
  XOR \MIXCOLUMNS[0].d/U394  ( .A(\w3[0][10] ), .B(\w3[0][2] ), .Z(
        \MIXCOLUMNS[0].d/n239 ) );
  XOR \MIXCOLUMNS[0].d/U393  ( .A(\MIXCOLUMNS[0].d/n239 ), .B(
        \MIXCOLUMNS[0].d/n20 ), .Z(\w0[1][9] ) );
  XOR \MIXCOLUMNS[0].d/U392  ( .A(n1151), .B(\MIXCOLUMNS[0].d/n235 ), .Z(
        \MIXCOLUMNS[0].d/n20 ) );
  XOR \MIXCOLUMNS[0].d/U391  ( .A(n535), .B(n1149), .Z(\MIXCOLUMNS[0].d/n241 )
         );
  XOR \MIXCOLUMNS[0].d/U390  ( .A(\MIXCOLUMNS[0].d/n241 ), .B(
        \MIXCOLUMNS[0].d/n21 ), .Z(\w0[1][10] ) );
  XOR \MIXCOLUMNS[0].d/U389  ( .A(\w3[0][2] ), .B(\MIXCOLUMNS[0].d/n238 ), .Z(
        \MIXCOLUMNS[0].d/n21 ) );
  XOR \MIXCOLUMNS[0].d/U388  ( .A(n36), .B(n537), .Z(\MIXCOLUMNS[0].d/n236 )
         );
  XOR \MIXCOLUMNS[0].d/U387  ( .A(n533), .B(n1147), .Z(\MIXCOLUMNS[0].d/n243 )
         );
  XOR \MIXCOLUMNS[0].d/U386  ( .A(\MIXCOLUMNS[0].d/n23 ), .B(
        \MIXCOLUMNS[0].d/n22 ), .Z(\w0[1][11] ) );
  XOR \MIXCOLUMNS[0].d/U385  ( .A(\MIXCOLUMNS[0].d/n240 ), .B(
        \MIXCOLUMNS[0].d/n243 ), .Z(\MIXCOLUMNS[0].d/n22 ) );
  XOR \MIXCOLUMNS[0].d/U384  ( .A(n1149), .B(\MIXCOLUMNS[0].d/n236 ), .Z(
        \MIXCOLUMNS[0].d/n23 ) );
  XOR \MIXCOLUMNS[0].d/U383  ( .A(n531), .B(n1145), .Z(\MIXCOLUMNS[0].d/n245 )
         );
  XOR \MIXCOLUMNS[0].d/U382  ( .A(\MIXCOLUMNS[0].d/n25 ), .B(
        \MIXCOLUMNS[0].d/n24 ), .Z(\w0[1][12] ) );
  XOR \MIXCOLUMNS[0].d/U381  ( .A(\MIXCOLUMNS[0].d/n242 ), .B(
        \MIXCOLUMNS[0].d/n245 ), .Z(\MIXCOLUMNS[0].d/n24 ) );
  XOR \MIXCOLUMNS[0].d/U380  ( .A(n1147), .B(\MIXCOLUMNS[0].d/n236 ), .Z(
        \MIXCOLUMNS[0].d/n25 ) );
  XOR \MIXCOLUMNS[0].d/U379  ( .A(n529), .B(n1143), .Z(\MIXCOLUMNS[0].d/n247 )
         );
  XOR \MIXCOLUMNS[0].d/U378  ( .A(\MIXCOLUMNS[0].d/n247 ), .B(
        \MIXCOLUMNS[0].d/n26 ), .Z(\w0[1][13] ) );
  XOR \MIXCOLUMNS[0].d/U377  ( .A(n1145), .B(\MIXCOLUMNS[0].d/n244 ), .Z(
        \MIXCOLUMNS[0].d/n26 ) );
  XOR \MIXCOLUMNS[0].d/U376  ( .A(n527), .B(n1141), .Z(\MIXCOLUMNS[0].d/n249 )
         );
  XOR \MIXCOLUMNS[0].d/U375  ( .A(\MIXCOLUMNS[0].d/n28 ), .B(
        \MIXCOLUMNS[0].d/n27 ), .Z(\w0[1][14] ) );
  XOR \MIXCOLUMNS[0].d/U374  ( .A(\MIXCOLUMNS[0].d/n246 ), .B(
        \MIXCOLUMNS[0].d/n249 ), .Z(\MIXCOLUMNS[0].d/n27 ) );
  XOR \MIXCOLUMNS[0].d/U373  ( .A(n1143), .B(\MIXCOLUMNS[0].d/n236 ), .Z(
        \MIXCOLUMNS[0].d/n28 ) );
  XOR \MIXCOLUMNS[0].d/U372  ( .A(\MIXCOLUMNS[0].d/n248 ), .B(
        \MIXCOLUMNS[0].d/n29 ), .Z(\w0[1][15] ) );
  XOR \MIXCOLUMNS[0].d/U371  ( .A(n1141), .B(\MIXCOLUMNS[0].d/n236 ), .Z(
        \MIXCOLUMNS[0].d/n29 ) );
  XOR \MIXCOLUMNS[0].d/U370  ( .A(\MIXCOLUMNS[0].d/n31 ), .B(
        \MIXCOLUMNS[0].d/n30 ), .Z(\w0[1][16] ) );
  XOR \MIXCOLUMNS[0].d/U369  ( .A(n538), .B(\MIXCOLUMNS[0].d/n236 ), .Z(
        \MIXCOLUMNS[0].d/n30 ) );
  XOR \MIXCOLUMNS[0].d/U368  ( .A(n1152), .B(n539), .Z(\MIXCOLUMNS[0].d/n31 )
         );
  XOR \MIXCOLUMNS[0].d/U367  ( .A(\MIXCOLUMNS[0].d/n33 ), .B(
        \MIXCOLUMNS[0].d/n32 ), .Z(\w0[1][17] ) );
  XOR \MIXCOLUMNS[0].d/U366  ( .A(\w3[0][10] ), .B(\MIXCOLUMNS[0].d/n237 ), 
        .Z(\MIXCOLUMNS[0].d/n32 ) );
  XOR \MIXCOLUMNS[0].d/U365  ( .A(n1150), .B(\w3[0][18] ), .Z(
        \MIXCOLUMNS[0].d/n33 ) );
  XOR \MIXCOLUMNS[0].d/U364  ( .A(\MIXCOLUMNS[0].d/n35 ), .B(
        \MIXCOLUMNS[0].d/n34 ), .Z(\w0[1][18] ) );
  XOR \MIXCOLUMNS[0].d/U363  ( .A(n535), .B(\MIXCOLUMNS[0].d/n239 ), .Z(
        \MIXCOLUMNS[0].d/n34 ) );
  XOR \MIXCOLUMNS[0].d/U362  ( .A(\w3[0][26] ), .B(n536), .Z(
        \MIXCOLUMNS[0].d/n35 ) );
  XOR \MIXCOLUMNS[0].d/U361  ( .A(n540), .B(n36), .Z(\MIXCOLUMNS[0].d/n234 )
         );
  XOR \MIXCOLUMNS[0].d/U360  ( .A(\MIXCOLUMNS[0].d/n37 ), .B(
        \MIXCOLUMNS[0].d/n36 ), .Z(\w0[1][19] ) );
  XOR \MIXCOLUMNS[0].d/U359  ( .A(\MIXCOLUMNS[0].d/n241 ), .B(
        \MIXCOLUMNS[0].d/n38 ), .Z(\MIXCOLUMNS[0].d/n36 ) );
  XOR \MIXCOLUMNS[0].d/U358  ( .A(n533), .B(\MIXCOLUMNS[0].d/n234 ), .Z(
        \MIXCOLUMNS[0].d/n37 ) );
  XOR \MIXCOLUMNS[0].d/U357  ( .A(n1148), .B(n534), .Z(\MIXCOLUMNS[0].d/n38 )
         );
  XOR \MIXCOLUMNS[0].d/U356  ( .A(\MIXCOLUMNS[0].d/n40 ), .B(
        \MIXCOLUMNS[0].d/n39 ), .Z(\w0[1][20] ) );
  XOR \MIXCOLUMNS[0].d/U355  ( .A(\MIXCOLUMNS[0].d/n243 ), .B(
        \MIXCOLUMNS[0].d/n41 ), .Z(\MIXCOLUMNS[0].d/n39 ) );
  XOR \MIXCOLUMNS[0].d/U354  ( .A(n531), .B(\MIXCOLUMNS[0].d/n234 ), .Z(
        \MIXCOLUMNS[0].d/n40 ) );
  XOR \MIXCOLUMNS[0].d/U353  ( .A(n1146), .B(n532), .Z(\MIXCOLUMNS[0].d/n41 )
         );
  XOR \MIXCOLUMNS[0].d/U352  ( .A(\MIXCOLUMNS[0].d/n43 ), .B(
        \MIXCOLUMNS[0].d/n42 ), .Z(\w0[1][21] ) );
  XOR \MIXCOLUMNS[0].d/U351  ( .A(n529), .B(\MIXCOLUMNS[0].d/n245 ), .Z(
        \MIXCOLUMNS[0].d/n42 ) );
  XOR \MIXCOLUMNS[0].d/U350  ( .A(n1144), .B(n530), .Z(\MIXCOLUMNS[0].d/n43 )
         );
  XOR \MIXCOLUMNS[0].d/U349  ( .A(\MIXCOLUMNS[0].d/n45 ), .B(
        \MIXCOLUMNS[0].d/n44 ), .Z(\w0[1][22] ) );
  XOR \MIXCOLUMNS[0].d/U348  ( .A(\MIXCOLUMNS[0].d/n247 ), .B(
        \MIXCOLUMNS[0].d/n46 ), .Z(\MIXCOLUMNS[0].d/n44 ) );
  XOR \MIXCOLUMNS[0].d/U347  ( .A(n527), .B(\MIXCOLUMNS[0].d/n234 ), .Z(
        \MIXCOLUMNS[0].d/n45 ) );
  XOR \MIXCOLUMNS[0].d/U346  ( .A(n1142), .B(n528), .Z(\MIXCOLUMNS[0].d/n46 )
         );
  XOR \MIXCOLUMNS[0].d/U345  ( .A(\MIXCOLUMNS[0].d/n249 ), .B(
        \MIXCOLUMNS[0].d/n47 ), .Z(\w0[1][23] ) );
  XOR \MIXCOLUMNS[0].d/U344  ( .A(n1140), .B(\MIXCOLUMNS[0].d/n234 ), .Z(
        \MIXCOLUMNS[0].d/n47 ) );
  XOR \MIXCOLUMNS[0].d/U343  ( .A(\MIXCOLUMNS[0].d/n235 ), .B(
        \MIXCOLUMNS[0].d/n48 ), .Z(\w0[1][24] ) );
  XOR \MIXCOLUMNS[0].d/U342  ( .A(n540), .B(\MIXCOLUMNS[0].d/n236 ), .Z(
        \MIXCOLUMNS[0].d/n48 ) );
  XOR \MIXCOLUMNS[0].d/U341  ( .A(\MIXCOLUMNS[0].d/n237 ), .B(
        \MIXCOLUMNS[0].d/n49 ), .Z(\w0[1][25] ) );
  XOR \MIXCOLUMNS[0].d/U340  ( .A(n539), .B(\MIXCOLUMNS[0].d/n238 ), .Z(
        \MIXCOLUMNS[0].d/n49 ) );
  XOR \MIXCOLUMNS[0].d/U339  ( .A(\MIXCOLUMNS[0].d/n239 ), .B(
        \MIXCOLUMNS[0].d/n50 ), .Z(\w0[1][26] ) );
  XOR \MIXCOLUMNS[0].d/U338  ( .A(\w3[0][18] ), .B(\MIXCOLUMNS[0].d/n240 ), 
        .Z(\MIXCOLUMNS[0].d/n50 ) );
  XOR \MIXCOLUMNS[0].d/U337  ( .A(\MIXCOLUMNS[0].d/n52 ), .B(
        \MIXCOLUMNS[0].d/n51 ), .Z(\w0[1][27] ) );
  XOR \MIXCOLUMNS[0].d/U336  ( .A(\MIXCOLUMNS[0].d/n242 ), .B(
        \MIXCOLUMNS[0].d/n241 ), .Z(\MIXCOLUMNS[0].d/n51 ) );
  XOR \MIXCOLUMNS[0].d/U335  ( .A(n536), .B(\MIXCOLUMNS[0].d/n250 ), .Z(
        \MIXCOLUMNS[0].d/n52 ) );
  XOR \MIXCOLUMNS[0].d/U334  ( .A(\MIXCOLUMNS[0].d/n54 ), .B(
        \MIXCOLUMNS[0].d/n53 ), .Z(\w0[1][28] ) );
  XOR \MIXCOLUMNS[0].d/U333  ( .A(\MIXCOLUMNS[0].d/n244 ), .B(
        \MIXCOLUMNS[0].d/n243 ), .Z(\MIXCOLUMNS[0].d/n53 ) );
  XOR \MIXCOLUMNS[0].d/U332  ( .A(n534), .B(\MIXCOLUMNS[0].d/n250 ), .Z(
        \MIXCOLUMNS[0].d/n54 ) );
  XOR \MIXCOLUMNS[0].d/U331  ( .A(\MIXCOLUMNS[0].d/n245 ), .B(
        \MIXCOLUMNS[0].d/n55 ), .Z(\w0[1][29] ) );
  XOR \MIXCOLUMNS[0].d/U330  ( .A(n532), .B(\MIXCOLUMNS[0].d/n246 ), .Z(
        \MIXCOLUMNS[0].d/n55 ) );
  XOR \MIXCOLUMNS[0].d/U329  ( .A(\MIXCOLUMNS[0].d/n57 ), .B(
        \MIXCOLUMNS[0].d/n56 ), .Z(\w0[1][30] ) );
  XOR \MIXCOLUMNS[0].d/U328  ( .A(\MIXCOLUMNS[0].d/n248 ), .B(
        \MIXCOLUMNS[0].d/n247 ), .Z(\MIXCOLUMNS[0].d/n56 ) );
  XOR \MIXCOLUMNS[0].d/U327  ( .A(n530), .B(\MIXCOLUMNS[0].d/n250 ), .Z(
        \MIXCOLUMNS[0].d/n57 ) );
  XOR \MIXCOLUMNS[0].d/U326  ( .A(\MIXCOLUMNS[0].d/n249 ), .B(
        \MIXCOLUMNS[0].d/n58 ), .Z(\w0[1][31] ) );
  XOR \MIXCOLUMNS[0].d/U325  ( .A(n528), .B(\MIXCOLUMNS[0].d/n250 ), .Z(
        \MIXCOLUMNS[0].d/n58 ) );
  XOR \MIXCOLUMNS[0].d/U324  ( .A(n1139), .B(n526), .Z(\MIXCOLUMNS[0].d/n268 )
         );
  XOR \MIXCOLUMNS[0].d/U323  ( .A(\MIXCOLUMNS[0].d/n60 ), .B(
        \MIXCOLUMNS[0].d/n59 ), .Z(\w0[1][32] ) );
  XOR \MIXCOLUMNS[0].d/U322  ( .A(n1138), .B(\MIXCOLUMNS[0].d/n268 ), .Z(
        \MIXCOLUMNS[0].d/n59 ) );
  XOR \MIXCOLUMNS[0].d/U321  ( .A(n1137), .B(n35), .Z(\MIXCOLUMNS[0].d/n60 )
         );
  XOR \MIXCOLUMNS[0].d/U320  ( .A(n1137), .B(n525), .Z(\MIXCOLUMNS[0].d/n253 )
         );
  XOR \MIXCOLUMNS[0].d/U319  ( .A(\MIXCOLUMNS[0].d/n62 ), .B(
        \MIXCOLUMNS[0].d/n61 ), .Z(\w0[1][33] ) );
  XOR \MIXCOLUMNS[0].d/U318  ( .A(\w3[0][34] ), .B(\MIXCOLUMNS[0].d/n253 ), 
        .Z(\MIXCOLUMNS[0].d/n61 ) );
  XOR \MIXCOLUMNS[0].d/U317  ( .A(\w3[0][58] ), .B(n524), .Z(
        \MIXCOLUMNS[0].d/n62 ) );
  XOR \MIXCOLUMNS[0].d/U316  ( .A(\w3[0][58] ), .B(\w3[0][50] ), .Z(
        \MIXCOLUMNS[0].d/n256 ) );
  XOR \MIXCOLUMNS[0].d/U315  ( .A(\MIXCOLUMNS[0].d/n64 ), .B(
        \MIXCOLUMNS[0].d/n63 ), .Z(\w0[1][34] ) );
  XOR \MIXCOLUMNS[0].d/U314  ( .A(n1136), .B(\MIXCOLUMNS[0].d/n256 ), .Z(
        \MIXCOLUMNS[0].d/n63 ) );
  XOR \MIXCOLUMNS[0].d/U313  ( .A(n1135), .B(\w3[0][42] ), .Z(
        \MIXCOLUMNS[0].d/n64 ) );
  XOR \MIXCOLUMNS[0].d/U312  ( .A(n1139), .B(n523), .Z(\MIXCOLUMNS[0].d/n251 )
         );
  XOR \MIXCOLUMNS[0].d/U311  ( .A(n1135), .B(n522), .Z(\MIXCOLUMNS[0].d/n258 )
         );
  XOR \MIXCOLUMNS[0].d/U310  ( .A(\MIXCOLUMNS[0].d/n66 ), .B(
        \MIXCOLUMNS[0].d/n65 ), .Z(\w0[1][35] ) );
  XOR \MIXCOLUMNS[0].d/U309  ( .A(\MIXCOLUMNS[0].d/n258 ), .B(
        \MIXCOLUMNS[0].d/n67 ), .Z(\MIXCOLUMNS[0].d/n65 ) );
  XOR \MIXCOLUMNS[0].d/U308  ( .A(n1134), .B(\MIXCOLUMNS[0].d/n251 ), .Z(
        \MIXCOLUMNS[0].d/n66 ) );
  XOR \MIXCOLUMNS[0].d/U307  ( .A(n1133), .B(n521), .Z(\MIXCOLUMNS[0].d/n67 )
         );
  XOR \MIXCOLUMNS[0].d/U306  ( .A(n1133), .B(n520), .Z(\MIXCOLUMNS[0].d/n260 )
         );
  XOR \MIXCOLUMNS[0].d/U305  ( .A(\MIXCOLUMNS[0].d/n69 ), .B(
        \MIXCOLUMNS[0].d/n68 ), .Z(\w0[1][36] ) );
  XOR \MIXCOLUMNS[0].d/U304  ( .A(\MIXCOLUMNS[0].d/n260 ), .B(
        \MIXCOLUMNS[0].d/n70 ), .Z(\MIXCOLUMNS[0].d/n68 ) );
  XOR \MIXCOLUMNS[0].d/U303  ( .A(n1132), .B(\MIXCOLUMNS[0].d/n251 ), .Z(
        \MIXCOLUMNS[0].d/n69 ) );
  XOR \MIXCOLUMNS[0].d/U302  ( .A(n1131), .B(n519), .Z(\MIXCOLUMNS[0].d/n70 )
         );
  XOR \MIXCOLUMNS[0].d/U301  ( .A(n1131), .B(n518), .Z(\MIXCOLUMNS[0].d/n262 )
         );
  XOR \MIXCOLUMNS[0].d/U300  ( .A(\MIXCOLUMNS[0].d/n72 ), .B(
        \MIXCOLUMNS[0].d/n71 ), .Z(\w0[1][37] ) );
  XOR \MIXCOLUMNS[0].d/U299  ( .A(n1130), .B(\MIXCOLUMNS[0].d/n262 ), .Z(
        \MIXCOLUMNS[0].d/n71 ) );
  XOR \MIXCOLUMNS[0].d/U298  ( .A(n1129), .B(n517), .Z(\MIXCOLUMNS[0].d/n72 )
         );
  XOR \MIXCOLUMNS[0].d/U297  ( .A(n1129), .B(n516), .Z(\MIXCOLUMNS[0].d/n264 )
         );
  XOR \MIXCOLUMNS[0].d/U296  ( .A(\MIXCOLUMNS[0].d/n74 ), .B(
        \MIXCOLUMNS[0].d/n73 ), .Z(\w0[1][38] ) );
  XOR \MIXCOLUMNS[0].d/U295  ( .A(\MIXCOLUMNS[0].d/n264 ), .B(
        \MIXCOLUMNS[0].d/n75 ), .Z(\MIXCOLUMNS[0].d/n73 ) );
  XOR \MIXCOLUMNS[0].d/U294  ( .A(n1128), .B(\MIXCOLUMNS[0].d/n251 ), .Z(
        \MIXCOLUMNS[0].d/n74 ) );
  XOR \MIXCOLUMNS[0].d/U293  ( .A(n1127), .B(n515), .Z(\MIXCOLUMNS[0].d/n75 )
         );
  XOR \MIXCOLUMNS[0].d/U292  ( .A(n1127), .B(n514), .Z(\MIXCOLUMNS[0].d/n266 )
         );
  XOR \MIXCOLUMNS[0].d/U291  ( .A(\MIXCOLUMNS[0].d/n266 ), .B(
        \MIXCOLUMNS[0].d/n76 ), .Z(\w0[1][39] ) );
  XOR \MIXCOLUMNS[0].d/U290  ( .A(n513), .B(\MIXCOLUMNS[0].d/n251 ), .Z(
        \MIXCOLUMNS[0].d/n76 ) );
  XOR \MIXCOLUMNS[0].d/U289  ( .A(n524), .B(n1138), .Z(\MIXCOLUMNS[0].d/n255 )
         );
  XOR \MIXCOLUMNS[0].d/U288  ( .A(\MIXCOLUMNS[0].d/n255 ), .B(
        \MIXCOLUMNS[0].d/n77 ), .Z(\w0[1][40] ) );
  XOR \MIXCOLUMNS[0].d/U287  ( .A(n523), .B(\MIXCOLUMNS[0].d/n268 ), .Z(
        \MIXCOLUMNS[0].d/n77 ) );
  XOR \MIXCOLUMNS[0].d/U286  ( .A(\w3[0][42] ), .B(\w3[0][34] ), .Z(
        \MIXCOLUMNS[0].d/n257 ) );
  XOR \MIXCOLUMNS[0].d/U285  ( .A(\MIXCOLUMNS[0].d/n257 ), .B(
        \MIXCOLUMNS[0].d/n78 ), .Z(\w0[1][41] ) );
  XOR \MIXCOLUMNS[0].d/U284  ( .A(n1138), .B(\MIXCOLUMNS[0].d/n253 ), .Z(
        \MIXCOLUMNS[0].d/n78 ) );
  XOR \MIXCOLUMNS[0].d/U283  ( .A(n521), .B(n1136), .Z(\MIXCOLUMNS[0].d/n259 )
         );
  XOR \MIXCOLUMNS[0].d/U282  ( .A(\MIXCOLUMNS[0].d/n259 ), .B(
        \MIXCOLUMNS[0].d/n79 ), .Z(\w0[1][42] ) );
  XOR \MIXCOLUMNS[0].d/U281  ( .A(\w3[0][34] ), .B(\MIXCOLUMNS[0].d/n256 ), 
        .Z(\MIXCOLUMNS[0].d/n79 ) );
  XOR \MIXCOLUMNS[0].d/U280  ( .A(n35), .B(n523), .Z(\MIXCOLUMNS[0].d/n254 )
         );
  XOR \MIXCOLUMNS[0].d/U279  ( .A(n519), .B(n1134), .Z(\MIXCOLUMNS[0].d/n261 )
         );
  XOR \MIXCOLUMNS[0].d/U278  ( .A(\MIXCOLUMNS[0].d/n81 ), .B(
        \MIXCOLUMNS[0].d/n80 ), .Z(\w0[1][43] ) );
  XOR \MIXCOLUMNS[0].d/U277  ( .A(\MIXCOLUMNS[0].d/n258 ), .B(
        \MIXCOLUMNS[0].d/n261 ), .Z(\MIXCOLUMNS[0].d/n80 ) );
  XOR \MIXCOLUMNS[0].d/U276  ( .A(n1136), .B(\MIXCOLUMNS[0].d/n254 ), .Z(
        \MIXCOLUMNS[0].d/n81 ) );
  XOR \MIXCOLUMNS[0].d/U275  ( .A(n517), .B(n1132), .Z(\MIXCOLUMNS[0].d/n263 )
         );
  XOR \MIXCOLUMNS[0].d/U274  ( .A(\MIXCOLUMNS[0].d/n83 ), .B(
        \MIXCOLUMNS[0].d/n82 ), .Z(\w0[1][44] ) );
  XOR \MIXCOLUMNS[0].d/U273  ( .A(\MIXCOLUMNS[0].d/n260 ), .B(
        \MIXCOLUMNS[0].d/n263 ), .Z(\MIXCOLUMNS[0].d/n82 ) );
  XOR \MIXCOLUMNS[0].d/U272  ( .A(n1134), .B(\MIXCOLUMNS[0].d/n254 ), .Z(
        \MIXCOLUMNS[0].d/n83 ) );
  XOR \MIXCOLUMNS[0].d/U271  ( .A(n515), .B(n1130), .Z(\MIXCOLUMNS[0].d/n265 )
         );
  XOR \MIXCOLUMNS[0].d/U270  ( .A(\MIXCOLUMNS[0].d/n265 ), .B(
        \MIXCOLUMNS[0].d/n84 ), .Z(\w0[1][45] ) );
  XOR \MIXCOLUMNS[0].d/U269  ( .A(n1132), .B(\MIXCOLUMNS[0].d/n262 ), .Z(
        \MIXCOLUMNS[0].d/n84 ) );
  XOR \MIXCOLUMNS[0].d/U268  ( .A(n513), .B(n1128), .Z(\MIXCOLUMNS[0].d/n267 )
         );
  XOR \MIXCOLUMNS[0].d/U267  ( .A(\MIXCOLUMNS[0].d/n86 ), .B(
        \MIXCOLUMNS[0].d/n85 ), .Z(\w0[1][46] ) );
  XOR \MIXCOLUMNS[0].d/U266  ( .A(\MIXCOLUMNS[0].d/n264 ), .B(
        \MIXCOLUMNS[0].d/n267 ), .Z(\MIXCOLUMNS[0].d/n85 ) );
  XOR \MIXCOLUMNS[0].d/U265  ( .A(n1130), .B(\MIXCOLUMNS[0].d/n254 ), .Z(
        \MIXCOLUMNS[0].d/n86 ) );
  XOR \MIXCOLUMNS[0].d/U264  ( .A(\MIXCOLUMNS[0].d/n266 ), .B(
        \MIXCOLUMNS[0].d/n87 ), .Z(\w0[1][47] ) );
  XOR \MIXCOLUMNS[0].d/U263  ( .A(n1128), .B(\MIXCOLUMNS[0].d/n254 ), .Z(
        \MIXCOLUMNS[0].d/n87 ) );
  XOR \MIXCOLUMNS[0].d/U262  ( .A(\MIXCOLUMNS[0].d/n89 ), .B(
        \MIXCOLUMNS[0].d/n88 ), .Z(\w0[1][48] ) );
  XOR \MIXCOLUMNS[0].d/U261  ( .A(n524), .B(\MIXCOLUMNS[0].d/n254 ), .Z(
        \MIXCOLUMNS[0].d/n88 ) );
  XOR \MIXCOLUMNS[0].d/U260  ( .A(n1139), .B(n525), .Z(\MIXCOLUMNS[0].d/n89 )
         );
  XOR \MIXCOLUMNS[0].d/U259  ( .A(\MIXCOLUMNS[0].d/n91 ), .B(
        \MIXCOLUMNS[0].d/n90 ), .Z(\w0[1][49] ) );
  XOR \MIXCOLUMNS[0].d/U258  ( .A(\w3[0][42] ), .B(\MIXCOLUMNS[0].d/n255 ), 
        .Z(\MIXCOLUMNS[0].d/n90 ) );
  XOR \MIXCOLUMNS[0].d/U257  ( .A(n1137), .B(\w3[0][50] ), .Z(
        \MIXCOLUMNS[0].d/n91 ) );
  XOR \MIXCOLUMNS[0].d/U256  ( .A(\MIXCOLUMNS[0].d/n93 ), .B(
        \MIXCOLUMNS[0].d/n92 ), .Z(\w0[1][50] ) );
  XOR \MIXCOLUMNS[0].d/U255  ( .A(n521), .B(\MIXCOLUMNS[0].d/n257 ), .Z(
        \MIXCOLUMNS[0].d/n92 ) );
  XOR \MIXCOLUMNS[0].d/U254  ( .A(\w3[0][58] ), .B(n522), .Z(
        \MIXCOLUMNS[0].d/n93 ) );
  XOR \MIXCOLUMNS[0].d/U253  ( .A(n526), .B(n35), .Z(\MIXCOLUMNS[0].d/n252 )
         );
  XOR \MIXCOLUMNS[0].d/U252  ( .A(\MIXCOLUMNS[0].d/n95 ), .B(
        \MIXCOLUMNS[0].d/n94 ), .Z(\w0[1][51] ) );
  XOR \MIXCOLUMNS[0].d/U251  ( .A(\MIXCOLUMNS[0].d/n259 ), .B(
        \MIXCOLUMNS[0].d/n96 ), .Z(\MIXCOLUMNS[0].d/n94 ) );
  XOR \MIXCOLUMNS[0].d/U250  ( .A(n519), .B(\MIXCOLUMNS[0].d/n252 ), .Z(
        \MIXCOLUMNS[0].d/n95 ) );
  XOR \MIXCOLUMNS[0].d/U249  ( .A(n1135), .B(n520), .Z(\MIXCOLUMNS[0].d/n96 )
         );
  XOR \MIXCOLUMNS[0].d/U248  ( .A(\MIXCOLUMNS[0].d/n98 ), .B(
        \MIXCOLUMNS[0].d/n97 ), .Z(\w0[1][52] ) );
  XOR \MIXCOLUMNS[0].d/U247  ( .A(\MIXCOLUMNS[0].d/n261 ), .B(
        \MIXCOLUMNS[0].d/n99 ), .Z(\MIXCOLUMNS[0].d/n97 ) );
  XOR \MIXCOLUMNS[0].d/U246  ( .A(n517), .B(\MIXCOLUMNS[0].d/n252 ), .Z(
        \MIXCOLUMNS[0].d/n98 ) );
  XOR \MIXCOLUMNS[0].d/U245  ( .A(n1133), .B(n518), .Z(\MIXCOLUMNS[0].d/n99 )
         );
  XOR \MIXCOLUMNS[0].d/U244  ( .A(\MIXCOLUMNS[0].d/n101 ), .B(
        \MIXCOLUMNS[0].d/n100 ), .Z(\w0[1][53] ) );
  XOR \MIXCOLUMNS[0].d/U243  ( .A(n515), .B(\MIXCOLUMNS[0].d/n263 ), .Z(
        \MIXCOLUMNS[0].d/n100 ) );
  XOR \MIXCOLUMNS[0].d/U242  ( .A(n1131), .B(n516), .Z(\MIXCOLUMNS[0].d/n101 )
         );
  XOR \MIXCOLUMNS[0].d/U241  ( .A(\MIXCOLUMNS[0].d/n103 ), .B(
        \MIXCOLUMNS[0].d/n102 ), .Z(\w0[1][54] ) );
  XOR \MIXCOLUMNS[0].d/U240  ( .A(\MIXCOLUMNS[0].d/n265 ), .B(
        \MIXCOLUMNS[0].d/n104 ), .Z(\MIXCOLUMNS[0].d/n102 ) );
  XOR \MIXCOLUMNS[0].d/U239  ( .A(n513), .B(\MIXCOLUMNS[0].d/n252 ), .Z(
        \MIXCOLUMNS[0].d/n103 ) );
  XOR \MIXCOLUMNS[0].d/U238  ( .A(n1129), .B(n514), .Z(\MIXCOLUMNS[0].d/n104 )
         );
  XOR \MIXCOLUMNS[0].d/U237  ( .A(\MIXCOLUMNS[0].d/n267 ), .B(
        \MIXCOLUMNS[0].d/n105 ), .Z(\w0[1][55] ) );
  XOR \MIXCOLUMNS[0].d/U236  ( .A(n1127), .B(\MIXCOLUMNS[0].d/n252 ), .Z(
        \MIXCOLUMNS[0].d/n105 ) );
  XOR \MIXCOLUMNS[0].d/U235  ( .A(\MIXCOLUMNS[0].d/n253 ), .B(
        \MIXCOLUMNS[0].d/n106 ), .Z(\w0[1][56] ) );
  XOR \MIXCOLUMNS[0].d/U234  ( .A(n526), .B(\MIXCOLUMNS[0].d/n254 ), .Z(
        \MIXCOLUMNS[0].d/n106 ) );
  XOR \MIXCOLUMNS[0].d/U233  ( .A(\MIXCOLUMNS[0].d/n255 ), .B(
        \MIXCOLUMNS[0].d/n107 ), .Z(\w0[1][57] ) );
  XOR \MIXCOLUMNS[0].d/U232  ( .A(n525), .B(\MIXCOLUMNS[0].d/n256 ), .Z(
        \MIXCOLUMNS[0].d/n107 ) );
  XOR \MIXCOLUMNS[0].d/U231  ( .A(\MIXCOLUMNS[0].d/n257 ), .B(
        \MIXCOLUMNS[0].d/n108 ), .Z(\w0[1][58] ) );
  XOR \MIXCOLUMNS[0].d/U230  ( .A(\w3[0][50] ), .B(\MIXCOLUMNS[0].d/n258 ), 
        .Z(\MIXCOLUMNS[0].d/n108 ) );
  XOR \MIXCOLUMNS[0].d/U229  ( .A(\MIXCOLUMNS[0].d/n110 ), .B(
        \MIXCOLUMNS[0].d/n109 ), .Z(\w0[1][59] ) );
  XOR \MIXCOLUMNS[0].d/U228  ( .A(\MIXCOLUMNS[0].d/n260 ), .B(
        \MIXCOLUMNS[0].d/n259 ), .Z(\MIXCOLUMNS[0].d/n109 ) );
  XOR \MIXCOLUMNS[0].d/U227  ( .A(n522), .B(\MIXCOLUMNS[0].d/n268 ), .Z(
        \MIXCOLUMNS[0].d/n110 ) );
  XOR \MIXCOLUMNS[0].d/U226  ( .A(\MIXCOLUMNS[0].d/n112 ), .B(
        \MIXCOLUMNS[0].d/n111 ), .Z(\w0[1][60] ) );
  XOR \MIXCOLUMNS[0].d/U225  ( .A(\MIXCOLUMNS[0].d/n262 ), .B(
        \MIXCOLUMNS[0].d/n261 ), .Z(\MIXCOLUMNS[0].d/n111 ) );
  XOR \MIXCOLUMNS[0].d/U224  ( .A(n520), .B(\MIXCOLUMNS[0].d/n268 ), .Z(
        \MIXCOLUMNS[0].d/n112 ) );
  XOR \MIXCOLUMNS[0].d/U223  ( .A(\MIXCOLUMNS[0].d/n263 ), .B(
        \MIXCOLUMNS[0].d/n113 ), .Z(\w0[1][61] ) );
  XOR \MIXCOLUMNS[0].d/U222  ( .A(n518), .B(\MIXCOLUMNS[0].d/n264 ), .Z(
        \MIXCOLUMNS[0].d/n113 ) );
  XOR \MIXCOLUMNS[0].d/U221  ( .A(\MIXCOLUMNS[0].d/n115 ), .B(
        \MIXCOLUMNS[0].d/n114 ), .Z(\w0[1][62] ) );
  XOR \MIXCOLUMNS[0].d/U220  ( .A(\MIXCOLUMNS[0].d/n266 ), .B(
        \MIXCOLUMNS[0].d/n265 ), .Z(\MIXCOLUMNS[0].d/n114 ) );
  XOR \MIXCOLUMNS[0].d/U219  ( .A(n516), .B(\MIXCOLUMNS[0].d/n268 ), .Z(
        \MIXCOLUMNS[0].d/n115 ) );
  XOR \MIXCOLUMNS[0].d/U218  ( .A(\MIXCOLUMNS[0].d/n267 ), .B(
        \MIXCOLUMNS[0].d/n116 ), .Z(\w0[1][63] ) );
  XOR \MIXCOLUMNS[0].d/U217  ( .A(n514), .B(\MIXCOLUMNS[0].d/n268 ), .Z(
        \MIXCOLUMNS[0].d/n116 ) );
  XOR \MIXCOLUMNS[0].d/U216  ( .A(n1126), .B(n512), .Z(\MIXCOLUMNS[0].d/n286 )
         );
  XOR \MIXCOLUMNS[0].d/U215  ( .A(\MIXCOLUMNS[0].d/n118 ), .B(
        \MIXCOLUMNS[0].d/n117 ), .Z(\w0[1][64] ) );
  XOR \MIXCOLUMNS[0].d/U214  ( .A(n1125), .B(\MIXCOLUMNS[0].d/n286 ), .Z(
        \MIXCOLUMNS[0].d/n117 ) );
  XOR \MIXCOLUMNS[0].d/U213  ( .A(n1124), .B(n34), .Z(\MIXCOLUMNS[0].d/n118 )
         );
  XOR \MIXCOLUMNS[0].d/U212  ( .A(n1124), .B(n511), .Z(\MIXCOLUMNS[0].d/n271 )
         );
  XOR \MIXCOLUMNS[0].d/U211  ( .A(\MIXCOLUMNS[0].d/n120 ), .B(
        \MIXCOLUMNS[0].d/n119 ), .Z(\w0[1][65] ) );
  XOR \MIXCOLUMNS[0].d/U210  ( .A(\w3[0][66] ), .B(\MIXCOLUMNS[0].d/n271 ), 
        .Z(\MIXCOLUMNS[0].d/n119 ) );
  XOR \MIXCOLUMNS[0].d/U209  ( .A(\w3[0][90] ), .B(n510), .Z(
        \MIXCOLUMNS[0].d/n120 ) );
  XOR \MIXCOLUMNS[0].d/U208  ( .A(\w3[0][90] ), .B(\w3[0][82] ), .Z(
        \MIXCOLUMNS[0].d/n274 ) );
  XOR \MIXCOLUMNS[0].d/U207  ( .A(\MIXCOLUMNS[0].d/n122 ), .B(
        \MIXCOLUMNS[0].d/n121 ), .Z(\w0[1][66] ) );
  XOR \MIXCOLUMNS[0].d/U206  ( .A(n1123), .B(\MIXCOLUMNS[0].d/n274 ), .Z(
        \MIXCOLUMNS[0].d/n121 ) );
  XOR \MIXCOLUMNS[0].d/U205  ( .A(n1122), .B(\w3[0][74] ), .Z(
        \MIXCOLUMNS[0].d/n122 ) );
  XOR \MIXCOLUMNS[0].d/U204  ( .A(n1126), .B(n509), .Z(\MIXCOLUMNS[0].d/n269 )
         );
  XOR \MIXCOLUMNS[0].d/U203  ( .A(n1122), .B(n508), .Z(\MIXCOLUMNS[0].d/n276 )
         );
  XOR \MIXCOLUMNS[0].d/U202  ( .A(\MIXCOLUMNS[0].d/n124 ), .B(
        \MIXCOLUMNS[0].d/n123 ), .Z(\w0[1][67] ) );
  XOR \MIXCOLUMNS[0].d/U201  ( .A(\MIXCOLUMNS[0].d/n276 ), .B(
        \MIXCOLUMNS[0].d/n125 ), .Z(\MIXCOLUMNS[0].d/n123 ) );
  XOR \MIXCOLUMNS[0].d/U200  ( .A(n1121), .B(\MIXCOLUMNS[0].d/n269 ), .Z(
        \MIXCOLUMNS[0].d/n124 ) );
  XOR \MIXCOLUMNS[0].d/U199  ( .A(n1120), .B(n507), .Z(\MIXCOLUMNS[0].d/n125 )
         );
  XOR \MIXCOLUMNS[0].d/U198  ( .A(n1120), .B(n506), .Z(\MIXCOLUMNS[0].d/n278 )
         );
  XOR \MIXCOLUMNS[0].d/U197  ( .A(\MIXCOLUMNS[0].d/n127 ), .B(
        \MIXCOLUMNS[0].d/n126 ), .Z(\w0[1][68] ) );
  XOR \MIXCOLUMNS[0].d/U196  ( .A(\MIXCOLUMNS[0].d/n278 ), .B(
        \MIXCOLUMNS[0].d/n128 ), .Z(\MIXCOLUMNS[0].d/n126 ) );
  XOR \MIXCOLUMNS[0].d/U195  ( .A(n1119), .B(\MIXCOLUMNS[0].d/n269 ), .Z(
        \MIXCOLUMNS[0].d/n127 ) );
  XOR \MIXCOLUMNS[0].d/U194  ( .A(n1118), .B(n505), .Z(\MIXCOLUMNS[0].d/n128 )
         );
  XOR \MIXCOLUMNS[0].d/U193  ( .A(n1118), .B(n504), .Z(\MIXCOLUMNS[0].d/n280 )
         );
  XOR \MIXCOLUMNS[0].d/U192  ( .A(\MIXCOLUMNS[0].d/n130 ), .B(
        \MIXCOLUMNS[0].d/n129 ), .Z(\w0[1][69] ) );
  XOR \MIXCOLUMNS[0].d/U191  ( .A(n1117), .B(\MIXCOLUMNS[0].d/n280 ), .Z(
        \MIXCOLUMNS[0].d/n129 ) );
  XOR \MIXCOLUMNS[0].d/U190  ( .A(n1116), .B(n503), .Z(\MIXCOLUMNS[0].d/n130 )
         );
  XOR \MIXCOLUMNS[0].d/U189  ( .A(n1116), .B(n502), .Z(\MIXCOLUMNS[0].d/n282 )
         );
  XOR \MIXCOLUMNS[0].d/U188  ( .A(\MIXCOLUMNS[0].d/n132 ), .B(
        \MIXCOLUMNS[0].d/n131 ), .Z(\w0[1][70] ) );
  XOR \MIXCOLUMNS[0].d/U187  ( .A(\MIXCOLUMNS[0].d/n282 ), .B(
        \MIXCOLUMNS[0].d/n133 ), .Z(\MIXCOLUMNS[0].d/n131 ) );
  XOR \MIXCOLUMNS[0].d/U186  ( .A(n1115), .B(\MIXCOLUMNS[0].d/n269 ), .Z(
        \MIXCOLUMNS[0].d/n132 ) );
  XOR \MIXCOLUMNS[0].d/U185  ( .A(n1114), .B(n501), .Z(\MIXCOLUMNS[0].d/n133 )
         );
  XOR \MIXCOLUMNS[0].d/U184  ( .A(n1114), .B(n500), .Z(\MIXCOLUMNS[0].d/n284 )
         );
  XOR \MIXCOLUMNS[0].d/U183  ( .A(\MIXCOLUMNS[0].d/n284 ), .B(
        \MIXCOLUMNS[0].d/n134 ), .Z(\w0[1][71] ) );
  XOR \MIXCOLUMNS[0].d/U182  ( .A(n499), .B(\MIXCOLUMNS[0].d/n269 ), .Z(
        \MIXCOLUMNS[0].d/n134 ) );
  XOR \MIXCOLUMNS[0].d/U181  ( .A(n510), .B(n1125), .Z(\MIXCOLUMNS[0].d/n273 )
         );
  XOR \MIXCOLUMNS[0].d/U180  ( .A(\MIXCOLUMNS[0].d/n273 ), .B(
        \MIXCOLUMNS[0].d/n135 ), .Z(\w0[1][72] ) );
  XOR \MIXCOLUMNS[0].d/U179  ( .A(n509), .B(\MIXCOLUMNS[0].d/n286 ), .Z(
        \MIXCOLUMNS[0].d/n135 ) );
  XOR \MIXCOLUMNS[0].d/U178  ( .A(\w3[0][74] ), .B(\w3[0][66] ), .Z(
        \MIXCOLUMNS[0].d/n275 ) );
  XOR \MIXCOLUMNS[0].d/U177  ( .A(\MIXCOLUMNS[0].d/n275 ), .B(
        \MIXCOLUMNS[0].d/n136 ), .Z(\w0[1][73] ) );
  XOR \MIXCOLUMNS[0].d/U176  ( .A(n1125), .B(\MIXCOLUMNS[0].d/n271 ), .Z(
        \MIXCOLUMNS[0].d/n136 ) );
  XOR \MIXCOLUMNS[0].d/U175  ( .A(n507), .B(n1123), .Z(\MIXCOLUMNS[0].d/n277 )
         );
  XOR \MIXCOLUMNS[0].d/U174  ( .A(\MIXCOLUMNS[0].d/n277 ), .B(
        \MIXCOLUMNS[0].d/n137 ), .Z(\w0[1][74] ) );
  XOR \MIXCOLUMNS[0].d/U173  ( .A(\w3[0][66] ), .B(\MIXCOLUMNS[0].d/n274 ), 
        .Z(\MIXCOLUMNS[0].d/n137 ) );
  XOR \MIXCOLUMNS[0].d/U172  ( .A(n34), .B(n509), .Z(\MIXCOLUMNS[0].d/n272 )
         );
  XOR \MIXCOLUMNS[0].d/U171  ( .A(n505), .B(n1121), .Z(\MIXCOLUMNS[0].d/n279 )
         );
  XOR \MIXCOLUMNS[0].d/U170  ( .A(\MIXCOLUMNS[0].d/n139 ), .B(
        \MIXCOLUMNS[0].d/n138 ), .Z(\w0[1][75] ) );
  XOR \MIXCOLUMNS[0].d/U169  ( .A(\MIXCOLUMNS[0].d/n276 ), .B(
        \MIXCOLUMNS[0].d/n279 ), .Z(\MIXCOLUMNS[0].d/n138 ) );
  XOR \MIXCOLUMNS[0].d/U168  ( .A(n1123), .B(\MIXCOLUMNS[0].d/n272 ), .Z(
        \MIXCOLUMNS[0].d/n139 ) );
  XOR \MIXCOLUMNS[0].d/U167  ( .A(n503), .B(n1119), .Z(\MIXCOLUMNS[0].d/n281 )
         );
  XOR \MIXCOLUMNS[0].d/U166  ( .A(\MIXCOLUMNS[0].d/n141 ), .B(
        \MIXCOLUMNS[0].d/n140 ), .Z(\w0[1][76] ) );
  XOR \MIXCOLUMNS[0].d/U165  ( .A(\MIXCOLUMNS[0].d/n278 ), .B(
        \MIXCOLUMNS[0].d/n281 ), .Z(\MIXCOLUMNS[0].d/n140 ) );
  XOR \MIXCOLUMNS[0].d/U164  ( .A(n1121), .B(\MIXCOLUMNS[0].d/n272 ), .Z(
        \MIXCOLUMNS[0].d/n141 ) );
  XOR \MIXCOLUMNS[0].d/U163  ( .A(n501), .B(n1117), .Z(\MIXCOLUMNS[0].d/n283 )
         );
  XOR \MIXCOLUMNS[0].d/U162  ( .A(\MIXCOLUMNS[0].d/n283 ), .B(
        \MIXCOLUMNS[0].d/n142 ), .Z(\w0[1][77] ) );
  XOR \MIXCOLUMNS[0].d/U161  ( .A(n1119), .B(\MIXCOLUMNS[0].d/n280 ), .Z(
        \MIXCOLUMNS[0].d/n142 ) );
  XOR \MIXCOLUMNS[0].d/U160  ( .A(n499), .B(n1115), .Z(\MIXCOLUMNS[0].d/n285 )
         );
  XOR \MIXCOLUMNS[0].d/U159  ( .A(\MIXCOLUMNS[0].d/n144 ), .B(
        \MIXCOLUMNS[0].d/n143 ), .Z(\w0[1][78] ) );
  XOR \MIXCOLUMNS[0].d/U158  ( .A(\MIXCOLUMNS[0].d/n282 ), .B(
        \MIXCOLUMNS[0].d/n285 ), .Z(\MIXCOLUMNS[0].d/n143 ) );
  XOR \MIXCOLUMNS[0].d/U157  ( .A(n1117), .B(\MIXCOLUMNS[0].d/n272 ), .Z(
        \MIXCOLUMNS[0].d/n144 ) );
  XOR \MIXCOLUMNS[0].d/U156  ( .A(\MIXCOLUMNS[0].d/n284 ), .B(
        \MIXCOLUMNS[0].d/n145 ), .Z(\w0[1][79] ) );
  XOR \MIXCOLUMNS[0].d/U155  ( .A(n1115), .B(\MIXCOLUMNS[0].d/n272 ), .Z(
        \MIXCOLUMNS[0].d/n145 ) );
  XOR \MIXCOLUMNS[0].d/U154  ( .A(\MIXCOLUMNS[0].d/n147 ), .B(
        \MIXCOLUMNS[0].d/n146 ), .Z(\w0[1][80] ) );
  XOR \MIXCOLUMNS[0].d/U153  ( .A(n510), .B(\MIXCOLUMNS[0].d/n272 ), .Z(
        \MIXCOLUMNS[0].d/n146 ) );
  XOR \MIXCOLUMNS[0].d/U152  ( .A(n1126), .B(n511), .Z(\MIXCOLUMNS[0].d/n147 )
         );
  XOR \MIXCOLUMNS[0].d/U151  ( .A(\MIXCOLUMNS[0].d/n149 ), .B(
        \MIXCOLUMNS[0].d/n148 ), .Z(\w0[1][81] ) );
  XOR \MIXCOLUMNS[0].d/U150  ( .A(\w3[0][74] ), .B(\MIXCOLUMNS[0].d/n273 ), 
        .Z(\MIXCOLUMNS[0].d/n148 ) );
  XOR \MIXCOLUMNS[0].d/U149  ( .A(n1124), .B(\w3[0][82] ), .Z(
        \MIXCOLUMNS[0].d/n149 ) );
  XOR \MIXCOLUMNS[0].d/U148  ( .A(\MIXCOLUMNS[0].d/n151 ), .B(
        \MIXCOLUMNS[0].d/n150 ), .Z(\w0[1][82] ) );
  XOR \MIXCOLUMNS[0].d/U147  ( .A(n507), .B(\MIXCOLUMNS[0].d/n275 ), .Z(
        \MIXCOLUMNS[0].d/n150 ) );
  XOR \MIXCOLUMNS[0].d/U146  ( .A(\w3[0][90] ), .B(n508), .Z(
        \MIXCOLUMNS[0].d/n151 ) );
  XOR \MIXCOLUMNS[0].d/U145  ( .A(n512), .B(n34), .Z(\MIXCOLUMNS[0].d/n270 )
         );
  XOR \MIXCOLUMNS[0].d/U144  ( .A(\MIXCOLUMNS[0].d/n153 ), .B(
        \MIXCOLUMNS[0].d/n152 ), .Z(\w0[1][83] ) );
  XOR \MIXCOLUMNS[0].d/U143  ( .A(\MIXCOLUMNS[0].d/n277 ), .B(
        \MIXCOLUMNS[0].d/n154 ), .Z(\MIXCOLUMNS[0].d/n152 ) );
  XOR \MIXCOLUMNS[0].d/U142  ( .A(n505), .B(\MIXCOLUMNS[0].d/n270 ), .Z(
        \MIXCOLUMNS[0].d/n153 ) );
  XOR \MIXCOLUMNS[0].d/U141  ( .A(n1122), .B(n506), .Z(\MIXCOLUMNS[0].d/n154 )
         );
  XOR \MIXCOLUMNS[0].d/U140  ( .A(\MIXCOLUMNS[0].d/n156 ), .B(
        \MIXCOLUMNS[0].d/n155 ), .Z(\w0[1][84] ) );
  XOR \MIXCOLUMNS[0].d/U139  ( .A(\MIXCOLUMNS[0].d/n279 ), .B(
        \MIXCOLUMNS[0].d/n157 ), .Z(\MIXCOLUMNS[0].d/n155 ) );
  XOR \MIXCOLUMNS[0].d/U138  ( .A(n503), .B(\MIXCOLUMNS[0].d/n270 ), .Z(
        \MIXCOLUMNS[0].d/n156 ) );
  XOR \MIXCOLUMNS[0].d/U137  ( .A(n1120), .B(n504), .Z(\MIXCOLUMNS[0].d/n157 )
         );
  XOR \MIXCOLUMNS[0].d/U136  ( .A(\MIXCOLUMNS[0].d/n159 ), .B(
        \MIXCOLUMNS[0].d/n158 ), .Z(\w0[1][85] ) );
  XOR \MIXCOLUMNS[0].d/U135  ( .A(n501), .B(\MIXCOLUMNS[0].d/n281 ), .Z(
        \MIXCOLUMNS[0].d/n158 ) );
  XOR \MIXCOLUMNS[0].d/U134  ( .A(n1118), .B(n502), .Z(\MIXCOLUMNS[0].d/n159 )
         );
  XOR \MIXCOLUMNS[0].d/U133  ( .A(\MIXCOLUMNS[0].d/n161 ), .B(
        \MIXCOLUMNS[0].d/n160 ), .Z(\w0[1][86] ) );
  XOR \MIXCOLUMNS[0].d/U132  ( .A(\MIXCOLUMNS[0].d/n283 ), .B(
        \MIXCOLUMNS[0].d/n162 ), .Z(\MIXCOLUMNS[0].d/n160 ) );
  XOR \MIXCOLUMNS[0].d/U131  ( .A(n499), .B(\MIXCOLUMNS[0].d/n270 ), .Z(
        \MIXCOLUMNS[0].d/n161 ) );
  XOR \MIXCOLUMNS[0].d/U130  ( .A(n1116), .B(n500), .Z(\MIXCOLUMNS[0].d/n162 )
         );
  XOR \MIXCOLUMNS[0].d/U129  ( .A(\MIXCOLUMNS[0].d/n285 ), .B(
        \MIXCOLUMNS[0].d/n163 ), .Z(\w0[1][87] ) );
  XOR \MIXCOLUMNS[0].d/U128  ( .A(n1114), .B(\MIXCOLUMNS[0].d/n270 ), .Z(
        \MIXCOLUMNS[0].d/n163 ) );
  XOR \MIXCOLUMNS[0].d/U127  ( .A(\MIXCOLUMNS[0].d/n271 ), .B(
        \MIXCOLUMNS[0].d/n164 ), .Z(\w0[1][88] ) );
  XOR \MIXCOLUMNS[0].d/U126  ( .A(n512), .B(\MIXCOLUMNS[0].d/n272 ), .Z(
        \MIXCOLUMNS[0].d/n164 ) );
  XOR \MIXCOLUMNS[0].d/U125  ( .A(\MIXCOLUMNS[0].d/n273 ), .B(
        \MIXCOLUMNS[0].d/n165 ), .Z(\w0[1][89] ) );
  XOR \MIXCOLUMNS[0].d/U124  ( .A(n511), .B(\MIXCOLUMNS[0].d/n274 ), .Z(
        \MIXCOLUMNS[0].d/n165 ) );
  XOR \MIXCOLUMNS[0].d/U123  ( .A(\MIXCOLUMNS[0].d/n275 ), .B(
        \MIXCOLUMNS[0].d/n166 ), .Z(\w0[1][90] ) );
  XOR \MIXCOLUMNS[0].d/U122  ( .A(\w3[0][82] ), .B(\MIXCOLUMNS[0].d/n276 ), 
        .Z(\MIXCOLUMNS[0].d/n166 ) );
  XOR \MIXCOLUMNS[0].d/U121  ( .A(\MIXCOLUMNS[0].d/n168 ), .B(
        \MIXCOLUMNS[0].d/n167 ), .Z(\w0[1][91] ) );
  XOR \MIXCOLUMNS[0].d/U120  ( .A(\MIXCOLUMNS[0].d/n278 ), .B(
        \MIXCOLUMNS[0].d/n277 ), .Z(\MIXCOLUMNS[0].d/n167 ) );
  XOR \MIXCOLUMNS[0].d/U119  ( .A(n508), .B(\MIXCOLUMNS[0].d/n286 ), .Z(
        \MIXCOLUMNS[0].d/n168 ) );
  XOR \MIXCOLUMNS[0].d/U118  ( .A(\MIXCOLUMNS[0].d/n170 ), .B(
        \MIXCOLUMNS[0].d/n169 ), .Z(\w0[1][92] ) );
  XOR \MIXCOLUMNS[0].d/U117  ( .A(\MIXCOLUMNS[0].d/n280 ), .B(
        \MIXCOLUMNS[0].d/n279 ), .Z(\MIXCOLUMNS[0].d/n169 ) );
  XOR \MIXCOLUMNS[0].d/U116  ( .A(n506), .B(\MIXCOLUMNS[0].d/n286 ), .Z(
        \MIXCOLUMNS[0].d/n170 ) );
  XOR \MIXCOLUMNS[0].d/U115  ( .A(\MIXCOLUMNS[0].d/n281 ), .B(
        \MIXCOLUMNS[0].d/n171 ), .Z(\w0[1][93] ) );
  XOR \MIXCOLUMNS[0].d/U114  ( .A(n504), .B(\MIXCOLUMNS[0].d/n282 ), .Z(
        \MIXCOLUMNS[0].d/n171 ) );
  XOR \MIXCOLUMNS[0].d/U113  ( .A(\MIXCOLUMNS[0].d/n173 ), .B(
        \MIXCOLUMNS[0].d/n172 ), .Z(\w0[1][94] ) );
  XOR \MIXCOLUMNS[0].d/U112  ( .A(\MIXCOLUMNS[0].d/n284 ), .B(
        \MIXCOLUMNS[0].d/n283 ), .Z(\MIXCOLUMNS[0].d/n172 ) );
  XOR \MIXCOLUMNS[0].d/U111  ( .A(n502), .B(\MIXCOLUMNS[0].d/n286 ), .Z(
        \MIXCOLUMNS[0].d/n173 ) );
  XOR \MIXCOLUMNS[0].d/U110  ( .A(\MIXCOLUMNS[0].d/n285 ), .B(
        \MIXCOLUMNS[0].d/n174 ), .Z(\w0[1][95] ) );
  XOR \MIXCOLUMNS[0].d/U109  ( .A(n500), .B(\MIXCOLUMNS[0].d/n286 ), .Z(
        \MIXCOLUMNS[0].d/n174 ) );
  XOR \MIXCOLUMNS[0].d/U108  ( .A(n1113), .B(n498), .Z(\MIXCOLUMNS[0].d/n304 )
         );
  XOR \MIXCOLUMNS[0].d/U107  ( .A(\MIXCOLUMNS[0].d/n176 ), .B(
        \MIXCOLUMNS[0].d/n175 ), .Z(\w0[1][96] ) );
  XOR \MIXCOLUMNS[0].d/U106  ( .A(n1112), .B(\MIXCOLUMNS[0].d/n304 ), .Z(
        \MIXCOLUMNS[0].d/n175 ) );
  XOR \MIXCOLUMNS[0].d/U105  ( .A(n1111), .B(n33), .Z(\MIXCOLUMNS[0].d/n176 )
         );
  XOR \MIXCOLUMNS[0].d/U104  ( .A(n1111), .B(n497), .Z(\MIXCOLUMNS[0].d/n289 )
         );
  XOR \MIXCOLUMNS[0].d/U103  ( .A(\MIXCOLUMNS[0].d/n178 ), .B(
        \MIXCOLUMNS[0].d/n177 ), .Z(\w0[1][97] ) );
  XOR \MIXCOLUMNS[0].d/U102  ( .A(\w3[0][98] ), .B(\MIXCOLUMNS[0].d/n289 ), 
        .Z(\MIXCOLUMNS[0].d/n177 ) );
  XOR \MIXCOLUMNS[0].d/U101  ( .A(\w3[0][122] ), .B(n496), .Z(
        \MIXCOLUMNS[0].d/n178 ) );
  XOR \MIXCOLUMNS[0].d/U100  ( .A(\w3[0][122] ), .B(\w3[0][114] ), .Z(
        \MIXCOLUMNS[0].d/n292 ) );
  XOR \MIXCOLUMNS[0].d/U99  ( .A(\MIXCOLUMNS[0].d/n180 ), .B(
        \MIXCOLUMNS[0].d/n179 ), .Z(\w0[1][98] ) );
  XOR \MIXCOLUMNS[0].d/U98  ( .A(n1110), .B(\MIXCOLUMNS[0].d/n292 ), .Z(
        \MIXCOLUMNS[0].d/n179 ) );
  XOR \MIXCOLUMNS[0].d/U97  ( .A(n1109), .B(\w3[0][106] ), .Z(
        \MIXCOLUMNS[0].d/n180 ) );
  XOR \MIXCOLUMNS[0].d/U96  ( .A(n1113), .B(n495), .Z(\MIXCOLUMNS[0].d/n287 )
         );
  XOR \MIXCOLUMNS[0].d/U95  ( .A(n1109), .B(n494), .Z(\MIXCOLUMNS[0].d/n294 )
         );
  XOR \MIXCOLUMNS[0].d/U94  ( .A(\MIXCOLUMNS[0].d/n182 ), .B(
        \MIXCOLUMNS[0].d/n181 ), .Z(\w0[1][99] ) );
  XOR \MIXCOLUMNS[0].d/U93  ( .A(\MIXCOLUMNS[0].d/n294 ), .B(
        \MIXCOLUMNS[0].d/n183 ), .Z(\MIXCOLUMNS[0].d/n181 ) );
  XOR \MIXCOLUMNS[0].d/U92  ( .A(n1108), .B(\MIXCOLUMNS[0].d/n287 ), .Z(
        \MIXCOLUMNS[0].d/n182 ) );
  XOR \MIXCOLUMNS[0].d/U91  ( .A(n1107), .B(n493), .Z(\MIXCOLUMNS[0].d/n183 )
         );
  XOR \MIXCOLUMNS[0].d/U90  ( .A(n1107), .B(n492), .Z(\MIXCOLUMNS[0].d/n296 )
         );
  XOR \MIXCOLUMNS[0].d/U89  ( .A(\MIXCOLUMNS[0].d/n185 ), .B(
        \MIXCOLUMNS[0].d/n184 ), .Z(\w0[1][100] ) );
  XOR \MIXCOLUMNS[0].d/U88  ( .A(\MIXCOLUMNS[0].d/n296 ), .B(
        \MIXCOLUMNS[0].d/n186 ), .Z(\MIXCOLUMNS[0].d/n184 ) );
  XOR \MIXCOLUMNS[0].d/U87  ( .A(n1106), .B(\MIXCOLUMNS[0].d/n287 ), .Z(
        \MIXCOLUMNS[0].d/n185 ) );
  XOR \MIXCOLUMNS[0].d/U86  ( .A(n1105), .B(n491), .Z(\MIXCOLUMNS[0].d/n186 )
         );
  XOR \MIXCOLUMNS[0].d/U85  ( .A(n1105), .B(n490), .Z(\MIXCOLUMNS[0].d/n298 )
         );
  XOR \MIXCOLUMNS[0].d/U84  ( .A(\MIXCOLUMNS[0].d/n188 ), .B(
        \MIXCOLUMNS[0].d/n187 ), .Z(\w0[1][101] ) );
  XOR \MIXCOLUMNS[0].d/U83  ( .A(n1104), .B(\MIXCOLUMNS[0].d/n298 ), .Z(
        \MIXCOLUMNS[0].d/n187 ) );
  XOR \MIXCOLUMNS[0].d/U82  ( .A(n1103), .B(n489), .Z(\MIXCOLUMNS[0].d/n188 )
         );
  XOR \MIXCOLUMNS[0].d/U81  ( .A(n1103), .B(n488), .Z(\MIXCOLUMNS[0].d/n300 )
         );
  XOR \MIXCOLUMNS[0].d/U80  ( .A(\MIXCOLUMNS[0].d/n190 ), .B(
        \MIXCOLUMNS[0].d/n189 ), .Z(\w0[1][102] ) );
  XOR \MIXCOLUMNS[0].d/U79  ( .A(\MIXCOLUMNS[0].d/n300 ), .B(
        \MIXCOLUMNS[0].d/n191 ), .Z(\MIXCOLUMNS[0].d/n189 ) );
  XOR \MIXCOLUMNS[0].d/U78  ( .A(n1102), .B(\MIXCOLUMNS[0].d/n287 ), .Z(
        \MIXCOLUMNS[0].d/n190 ) );
  XOR \MIXCOLUMNS[0].d/U77  ( .A(n1101), .B(n487), .Z(\MIXCOLUMNS[0].d/n191 )
         );
  XOR \MIXCOLUMNS[0].d/U76  ( .A(n1101), .B(n486), .Z(\MIXCOLUMNS[0].d/n302 )
         );
  XOR \MIXCOLUMNS[0].d/U75  ( .A(\MIXCOLUMNS[0].d/n302 ), .B(
        \MIXCOLUMNS[0].d/n192 ), .Z(\w0[1][103] ) );
  XOR \MIXCOLUMNS[0].d/U74  ( .A(n485), .B(\MIXCOLUMNS[0].d/n287 ), .Z(
        \MIXCOLUMNS[0].d/n192 ) );
  XOR \MIXCOLUMNS[0].d/U73  ( .A(n496), .B(n1112), .Z(\MIXCOLUMNS[0].d/n291 )
         );
  XOR \MIXCOLUMNS[0].d/U72  ( .A(\MIXCOLUMNS[0].d/n291 ), .B(
        \MIXCOLUMNS[0].d/n193 ), .Z(\w0[1][104] ) );
  XOR \MIXCOLUMNS[0].d/U71  ( .A(n495), .B(\MIXCOLUMNS[0].d/n304 ), .Z(
        \MIXCOLUMNS[0].d/n193 ) );
  XOR \MIXCOLUMNS[0].d/U70  ( .A(\w3[0][106] ), .B(\w3[0][98] ), .Z(
        \MIXCOLUMNS[0].d/n293 ) );
  XOR \MIXCOLUMNS[0].d/U69  ( .A(\MIXCOLUMNS[0].d/n293 ), .B(
        \MIXCOLUMNS[0].d/n194 ), .Z(\w0[1][105] ) );
  XOR \MIXCOLUMNS[0].d/U68  ( .A(n1112), .B(\MIXCOLUMNS[0].d/n289 ), .Z(
        \MIXCOLUMNS[0].d/n194 ) );
  XOR \MIXCOLUMNS[0].d/U67  ( .A(n493), .B(n1110), .Z(\MIXCOLUMNS[0].d/n295 )
         );
  XOR \MIXCOLUMNS[0].d/U66  ( .A(\MIXCOLUMNS[0].d/n295 ), .B(
        \MIXCOLUMNS[0].d/n195 ), .Z(\w0[1][106] ) );
  XOR \MIXCOLUMNS[0].d/U65  ( .A(\w3[0][98] ), .B(\MIXCOLUMNS[0].d/n292 ), .Z(
        \MIXCOLUMNS[0].d/n195 ) );
  XOR \MIXCOLUMNS[0].d/U64  ( .A(n33), .B(n495), .Z(\MIXCOLUMNS[0].d/n290 ) );
  XOR \MIXCOLUMNS[0].d/U63  ( .A(n491), .B(n1108), .Z(\MIXCOLUMNS[0].d/n297 )
         );
  XOR \MIXCOLUMNS[0].d/U62  ( .A(\MIXCOLUMNS[0].d/n197 ), .B(
        \MIXCOLUMNS[0].d/n196 ), .Z(\w0[1][107] ) );
  XOR \MIXCOLUMNS[0].d/U61  ( .A(\MIXCOLUMNS[0].d/n294 ), .B(
        \MIXCOLUMNS[0].d/n297 ), .Z(\MIXCOLUMNS[0].d/n196 ) );
  XOR \MIXCOLUMNS[0].d/U60  ( .A(n1110), .B(\MIXCOLUMNS[0].d/n290 ), .Z(
        \MIXCOLUMNS[0].d/n197 ) );
  XOR \MIXCOLUMNS[0].d/U59  ( .A(n489), .B(n1106), .Z(\MIXCOLUMNS[0].d/n299 )
         );
  XOR \MIXCOLUMNS[0].d/U58  ( .A(\MIXCOLUMNS[0].d/n199 ), .B(
        \MIXCOLUMNS[0].d/n198 ), .Z(\w0[1][108] ) );
  XOR \MIXCOLUMNS[0].d/U57  ( .A(\MIXCOLUMNS[0].d/n296 ), .B(
        \MIXCOLUMNS[0].d/n299 ), .Z(\MIXCOLUMNS[0].d/n198 ) );
  XOR \MIXCOLUMNS[0].d/U56  ( .A(n1108), .B(\MIXCOLUMNS[0].d/n290 ), .Z(
        \MIXCOLUMNS[0].d/n199 ) );
  XOR \MIXCOLUMNS[0].d/U55  ( .A(n487), .B(n1104), .Z(\MIXCOLUMNS[0].d/n301 )
         );
  XOR \MIXCOLUMNS[0].d/U54  ( .A(\MIXCOLUMNS[0].d/n301 ), .B(
        \MIXCOLUMNS[0].d/n200 ), .Z(\w0[1][109] ) );
  XOR \MIXCOLUMNS[0].d/U53  ( .A(n1106), .B(\MIXCOLUMNS[0].d/n298 ), .Z(
        \MIXCOLUMNS[0].d/n200 ) );
  XOR \MIXCOLUMNS[0].d/U52  ( .A(n485), .B(n1102), .Z(\MIXCOLUMNS[0].d/n303 )
         );
  XOR \MIXCOLUMNS[0].d/U51  ( .A(\MIXCOLUMNS[0].d/n202 ), .B(
        \MIXCOLUMNS[0].d/n201 ), .Z(\w0[1][110] ) );
  XOR \MIXCOLUMNS[0].d/U50  ( .A(\MIXCOLUMNS[0].d/n300 ), .B(
        \MIXCOLUMNS[0].d/n303 ), .Z(\MIXCOLUMNS[0].d/n201 ) );
  XOR \MIXCOLUMNS[0].d/U49  ( .A(n1104), .B(\MIXCOLUMNS[0].d/n290 ), .Z(
        \MIXCOLUMNS[0].d/n202 ) );
  XOR \MIXCOLUMNS[0].d/U48  ( .A(\MIXCOLUMNS[0].d/n302 ), .B(
        \MIXCOLUMNS[0].d/n203 ), .Z(\w0[1][111] ) );
  XOR \MIXCOLUMNS[0].d/U47  ( .A(n1102), .B(\MIXCOLUMNS[0].d/n290 ), .Z(
        \MIXCOLUMNS[0].d/n203 ) );
  XOR \MIXCOLUMNS[0].d/U46  ( .A(\MIXCOLUMNS[0].d/n205 ), .B(
        \MIXCOLUMNS[0].d/n204 ), .Z(\w0[1][112] ) );
  XOR \MIXCOLUMNS[0].d/U45  ( .A(n496), .B(\MIXCOLUMNS[0].d/n290 ), .Z(
        \MIXCOLUMNS[0].d/n204 ) );
  XOR \MIXCOLUMNS[0].d/U44  ( .A(n1113), .B(n497), .Z(\MIXCOLUMNS[0].d/n205 )
         );
  XOR \MIXCOLUMNS[0].d/U43  ( .A(\MIXCOLUMNS[0].d/n207 ), .B(
        \MIXCOLUMNS[0].d/n206 ), .Z(\w0[1][113] ) );
  XOR \MIXCOLUMNS[0].d/U42  ( .A(\w3[0][106] ), .B(\MIXCOLUMNS[0].d/n291 ), 
        .Z(\MIXCOLUMNS[0].d/n206 ) );
  XOR \MIXCOLUMNS[0].d/U41  ( .A(n1111), .B(\w3[0][114] ), .Z(
        \MIXCOLUMNS[0].d/n207 ) );
  XOR \MIXCOLUMNS[0].d/U40  ( .A(\MIXCOLUMNS[0].d/n209 ), .B(
        \MIXCOLUMNS[0].d/n208 ), .Z(\w0[1][114] ) );
  XOR \MIXCOLUMNS[0].d/U39  ( .A(n493), .B(\MIXCOLUMNS[0].d/n293 ), .Z(
        \MIXCOLUMNS[0].d/n208 ) );
  XOR \MIXCOLUMNS[0].d/U38  ( .A(\w3[0][122] ), .B(n494), .Z(
        \MIXCOLUMNS[0].d/n209 ) );
  XOR \MIXCOLUMNS[0].d/U37  ( .A(n498), .B(n33), .Z(\MIXCOLUMNS[0].d/n288 ) );
  XOR \MIXCOLUMNS[0].d/U36  ( .A(\MIXCOLUMNS[0].d/n211 ), .B(
        \MIXCOLUMNS[0].d/n210 ), .Z(\w0[1][115] ) );
  XOR \MIXCOLUMNS[0].d/U35  ( .A(\MIXCOLUMNS[0].d/n295 ), .B(
        \MIXCOLUMNS[0].d/n212 ), .Z(\MIXCOLUMNS[0].d/n210 ) );
  XOR \MIXCOLUMNS[0].d/U34  ( .A(n491), .B(\MIXCOLUMNS[0].d/n288 ), .Z(
        \MIXCOLUMNS[0].d/n211 ) );
  XOR \MIXCOLUMNS[0].d/U33  ( .A(n1109), .B(n492), .Z(\MIXCOLUMNS[0].d/n212 )
         );
  XOR \MIXCOLUMNS[0].d/U32  ( .A(\MIXCOLUMNS[0].d/n214 ), .B(
        \MIXCOLUMNS[0].d/n213 ), .Z(\w0[1][116] ) );
  XOR \MIXCOLUMNS[0].d/U31  ( .A(\MIXCOLUMNS[0].d/n297 ), .B(
        \MIXCOLUMNS[0].d/n215 ), .Z(\MIXCOLUMNS[0].d/n213 ) );
  XOR \MIXCOLUMNS[0].d/U30  ( .A(n489), .B(\MIXCOLUMNS[0].d/n288 ), .Z(
        \MIXCOLUMNS[0].d/n214 ) );
  XOR \MIXCOLUMNS[0].d/U29  ( .A(n1107), .B(n490), .Z(\MIXCOLUMNS[0].d/n215 )
         );
  XOR \MIXCOLUMNS[0].d/U28  ( .A(\MIXCOLUMNS[0].d/n217 ), .B(
        \MIXCOLUMNS[0].d/n216 ), .Z(\w0[1][117] ) );
  XOR \MIXCOLUMNS[0].d/U27  ( .A(n487), .B(\MIXCOLUMNS[0].d/n299 ), .Z(
        \MIXCOLUMNS[0].d/n216 ) );
  XOR \MIXCOLUMNS[0].d/U26  ( .A(n1105), .B(n488), .Z(\MIXCOLUMNS[0].d/n217 )
         );
  XOR \MIXCOLUMNS[0].d/U25  ( .A(\MIXCOLUMNS[0].d/n219 ), .B(
        \MIXCOLUMNS[0].d/n218 ), .Z(\w0[1][118] ) );
  XOR \MIXCOLUMNS[0].d/U24  ( .A(\MIXCOLUMNS[0].d/n301 ), .B(
        \MIXCOLUMNS[0].d/n220 ), .Z(\MIXCOLUMNS[0].d/n218 ) );
  XOR \MIXCOLUMNS[0].d/U23  ( .A(n485), .B(\MIXCOLUMNS[0].d/n288 ), .Z(
        \MIXCOLUMNS[0].d/n219 ) );
  XOR \MIXCOLUMNS[0].d/U22  ( .A(n1103), .B(n486), .Z(\MIXCOLUMNS[0].d/n220 )
         );
  XOR \MIXCOLUMNS[0].d/U21  ( .A(\MIXCOLUMNS[0].d/n303 ), .B(
        \MIXCOLUMNS[0].d/n221 ), .Z(\w0[1][119] ) );
  XOR \MIXCOLUMNS[0].d/U20  ( .A(n1101), .B(\MIXCOLUMNS[0].d/n288 ), .Z(
        \MIXCOLUMNS[0].d/n221 ) );
  XOR \MIXCOLUMNS[0].d/U19  ( .A(\MIXCOLUMNS[0].d/n289 ), .B(
        \MIXCOLUMNS[0].d/n222 ), .Z(\w0[1][120] ) );
  XOR \MIXCOLUMNS[0].d/U18  ( .A(n498), .B(\MIXCOLUMNS[0].d/n290 ), .Z(
        \MIXCOLUMNS[0].d/n222 ) );
  XOR \MIXCOLUMNS[0].d/U17  ( .A(\MIXCOLUMNS[0].d/n291 ), .B(
        \MIXCOLUMNS[0].d/n223 ), .Z(\w0[1][121] ) );
  XOR \MIXCOLUMNS[0].d/U16  ( .A(n497), .B(\MIXCOLUMNS[0].d/n292 ), .Z(
        \MIXCOLUMNS[0].d/n223 ) );
  XOR \MIXCOLUMNS[0].d/U15  ( .A(\MIXCOLUMNS[0].d/n293 ), .B(
        \MIXCOLUMNS[0].d/n224 ), .Z(\w0[1][122] ) );
  XOR \MIXCOLUMNS[0].d/U14  ( .A(\w3[0][114] ), .B(\MIXCOLUMNS[0].d/n294 ), 
        .Z(\MIXCOLUMNS[0].d/n224 ) );
  XOR \MIXCOLUMNS[0].d/U13  ( .A(\MIXCOLUMNS[0].d/n226 ), .B(
        \MIXCOLUMNS[0].d/n225 ), .Z(\w0[1][123] ) );
  XOR \MIXCOLUMNS[0].d/U12  ( .A(\MIXCOLUMNS[0].d/n296 ), .B(
        \MIXCOLUMNS[0].d/n295 ), .Z(\MIXCOLUMNS[0].d/n225 ) );
  XOR \MIXCOLUMNS[0].d/U11  ( .A(n494), .B(\MIXCOLUMNS[0].d/n304 ), .Z(
        \MIXCOLUMNS[0].d/n226 ) );
  XOR \MIXCOLUMNS[0].d/U10  ( .A(\MIXCOLUMNS[0].d/n228 ), .B(
        \MIXCOLUMNS[0].d/n227 ), .Z(\w0[1][124] ) );
  XOR \MIXCOLUMNS[0].d/U9  ( .A(\MIXCOLUMNS[0].d/n298 ), .B(
        \MIXCOLUMNS[0].d/n297 ), .Z(\MIXCOLUMNS[0].d/n227 ) );
  XOR \MIXCOLUMNS[0].d/U8  ( .A(n492), .B(\MIXCOLUMNS[0].d/n304 ), .Z(
        \MIXCOLUMNS[0].d/n228 ) );
  XOR \MIXCOLUMNS[0].d/U7  ( .A(\MIXCOLUMNS[0].d/n299 ), .B(
        \MIXCOLUMNS[0].d/n229 ), .Z(\w0[1][125] ) );
  XOR \MIXCOLUMNS[0].d/U6  ( .A(n490), .B(\MIXCOLUMNS[0].d/n300 ), .Z(
        \MIXCOLUMNS[0].d/n229 ) );
  XOR \MIXCOLUMNS[0].d/U5  ( .A(\MIXCOLUMNS[0].d/n231 ), .B(
        \MIXCOLUMNS[0].d/n230 ), .Z(\w0[1][126] ) );
  XOR \MIXCOLUMNS[0].d/U4  ( .A(\MIXCOLUMNS[0].d/n302 ), .B(
        \MIXCOLUMNS[0].d/n301 ), .Z(\MIXCOLUMNS[0].d/n230 ) );
  XOR \MIXCOLUMNS[0].d/U3  ( .A(n488), .B(\MIXCOLUMNS[0].d/n304 ), .Z(
        \MIXCOLUMNS[0].d/n231 ) );
  XOR \MIXCOLUMNS[0].d/U2  ( .A(\MIXCOLUMNS[0].d/n303 ), .B(
        \MIXCOLUMNS[0].d/n232 ), .Z(\w0[1][127] ) );
  XOR \MIXCOLUMNS[0].d/U1  ( .A(n486), .B(\MIXCOLUMNS[0].d/n304 ), .Z(
        \MIXCOLUMNS[0].d/n232 ) );
  XOR \SUBBYTES[9].a/U5649  ( .A(\SUBBYTES[9].a/w3390 ), .B(
        \SUBBYTES[9].a/w3391 ), .Z(n17145) );
  XOR \SUBBYTES[9].a/U5648  ( .A(n17145), .B(n16104), .Z(n17144) );
  XOR \SUBBYTES[9].a/U5647  ( .A(\SUBBYTES[9].a/w3383 ), .B(
        \SUBBYTES[9].a/w3400 ), .Z(n16104) );
  XOR \SUBBYTES[9].a/U5646  ( .A(n17144), .B(n16105), .Z(n17336) );
  XOR \SUBBYTES[9].a/U5645  ( .A(\SUBBYTES[9].a/w3382 ), .B(
        \SUBBYTES[9].a/w3397 ), .Z(n16105) );
  XOR \SUBBYTES[9].a/U5644  ( .A(n17145), .B(n16106), .Z(n17338) );
  XOR \SUBBYTES[9].a/U5643  ( .A(\SUBBYTES[9].a/w3397 ), .B(
        \SUBBYTES[9].a/w3398 ), .Z(n16106) );
  XOR \SUBBYTES[9].a/U5642  ( .A(\SUBBYTES[9].a/w3359 ), .B(n16107), .Z(n17147) );
  XOR \SUBBYTES[9].a/U5641  ( .A(\SUBBYTES[9].a/w3350 ), .B(
        \SUBBYTES[9].a/w3351 ), .Z(n16107) );
  XOR \SUBBYTES[9].a/U5640  ( .A(n17147), .B(n16108), .Z(n17337) );
  XOR \SUBBYTES[9].a/U5639  ( .A(\SUBBYTES[9].a/w3361 ), .B(n17338), .Z(n16108) );
  XOR \SUBBYTES[9].a/U5638  ( .A(n16110), .B(n16109), .Z(n17148) );
  XOR \SUBBYTES[9].a/U5637  ( .A(n16112), .B(n16111), .Z(n16109) );
  XOR \SUBBYTES[9].a/U5636  ( .A(\SUBBYTES[9].a/w3397 ), .B(
        \SUBBYTES[9].a/w3398 ), .Z(n16110) );
  XOR \SUBBYTES[9].a/U5635  ( .A(\SUBBYTES[9].a/w3361 ), .B(
        \SUBBYTES[9].a/w3385 ), .Z(n16111) );
  XOR \SUBBYTES[9].a/U5634  ( .A(\SUBBYTES[9].a/w3350 ), .B(
        \SUBBYTES[9].a/w3359 ), .Z(n16112) );
  XOR \SUBBYTES[9].a/U5633  ( .A(\SUBBYTES[9].a/w3382 ), .B(n16113), .Z(n17146) );
  XOR \SUBBYTES[9].a/U5632  ( .A(\SUBBYTES[9].a/w3365 ), .B(
        \SUBBYTES[9].a/w3368 ), .Z(n16113) );
  XOR \SUBBYTES[9].a/U5631  ( .A(n17146), .B(n16114), .Z(n17339) );
  XOR \SUBBYTES[9].a/U5630  ( .A(\SUBBYTES[9].a/w3353 ), .B(n17148), .Z(n16114) );
  XOR \SUBBYTES[9].a/U5629  ( .A(n17144), .B(n16115), .Z(n17340) );
  XOR \SUBBYTES[9].a/U5628  ( .A(\SUBBYTES[9].a/w3385 ), .B(
        \SUBBYTES[9].a/w3398 ), .Z(n16115) );
  XOR \SUBBYTES[9].a/U5627  ( .A(n16117), .B(n16116), .Z(n17341) );
  XOR \SUBBYTES[9].a/U5626  ( .A(n16119), .B(n16118), .Z(n16116) );
  XOR \SUBBYTES[9].a/U5625  ( .A(n16121), .B(n16120), .Z(n16117) );
  XOR \SUBBYTES[9].a/U5624  ( .A(\SUBBYTES[9].a/w3397 ), .B(
        \SUBBYTES[9].a/w3400 ), .Z(n16118) );
  XOR \SUBBYTES[9].a/U5623  ( .A(\SUBBYTES[9].a/w3390 ), .B(
        \SUBBYTES[9].a/w3393 ), .Z(n16119) );
  XOR \SUBBYTES[9].a/U5622  ( .A(\SUBBYTES[9].a/w3365 ), .B(
        \SUBBYTES[9].a/w3366 ), .Z(n16120) );
  XOR \SUBBYTES[9].a/U5621  ( .A(\SUBBYTES[9].a/w3350 ), .B(
        \SUBBYTES[9].a/w3353 ), .Z(n16121) );
  XOR \SUBBYTES[9].a/U5620  ( .A(n16123), .B(n16122), .Z(n17342) );
  XOR \SUBBYTES[9].a/U5619  ( .A(n17145), .B(n16124), .Z(n16122) );
  XOR \SUBBYTES[9].a/U5618  ( .A(n17147), .B(n17146), .Z(n16123) );
  XOR \SUBBYTES[9].a/U5617  ( .A(\SUBBYTES[9].a/w3358 ), .B(
        \SUBBYTES[9].a/w3385 ), .Z(n16124) );
  XOR \SUBBYTES[9].a/U5616  ( .A(n16126), .B(n16125), .Z(n17343) );
  XOR \SUBBYTES[9].a/U5615  ( .A(n17148), .B(n16127), .Z(n16125) );
  XOR \SUBBYTES[9].a/U5614  ( .A(\SUBBYTES[9].a/w3391 ), .B(
        \SUBBYTES[9].a/w3393 ), .Z(n16126) );
  XOR \SUBBYTES[9].a/U5613  ( .A(\SUBBYTES[9].a/w3351 ), .B(
        \SUBBYTES[9].a/w3383 ), .Z(n16127) );
  XOR \SUBBYTES[9].a/U5612  ( .A(\SUBBYTES[9].a/w3183 ), .B(
        \SUBBYTES[9].a/w3184 ), .Z(n17150) );
  XOR \SUBBYTES[9].a/U5611  ( .A(n17150), .B(n16128), .Z(n17149) );
  XOR \SUBBYTES[9].a/U5610  ( .A(\SUBBYTES[9].a/w3176 ), .B(
        \SUBBYTES[9].a/w3193 ), .Z(n16128) );
  XOR \SUBBYTES[9].a/U5609  ( .A(n17149), .B(n16129), .Z(n17344) );
  XOR \SUBBYTES[9].a/U5608  ( .A(\SUBBYTES[9].a/w3175 ), .B(
        \SUBBYTES[9].a/w3190 ), .Z(n16129) );
  XOR \SUBBYTES[9].a/U5607  ( .A(n17150), .B(n16130), .Z(n17346) );
  XOR \SUBBYTES[9].a/U5606  ( .A(\SUBBYTES[9].a/w3190 ), .B(
        \SUBBYTES[9].a/w3191 ), .Z(n16130) );
  XOR \SUBBYTES[9].a/U5605  ( .A(\SUBBYTES[9].a/w3152 ), .B(n16131), .Z(n17152) );
  XOR \SUBBYTES[9].a/U5604  ( .A(\SUBBYTES[9].a/w3143 ), .B(
        \SUBBYTES[9].a/w3144 ), .Z(n16131) );
  XOR \SUBBYTES[9].a/U5603  ( .A(n17152), .B(n16132), .Z(n17345) );
  XOR \SUBBYTES[9].a/U5602  ( .A(\SUBBYTES[9].a/w3154 ), .B(n17346), .Z(n16132) );
  XOR \SUBBYTES[9].a/U5601  ( .A(n16134), .B(n16133), .Z(n17153) );
  XOR \SUBBYTES[9].a/U5600  ( .A(n16136), .B(n16135), .Z(n16133) );
  XOR \SUBBYTES[9].a/U5599  ( .A(\SUBBYTES[9].a/w3190 ), .B(
        \SUBBYTES[9].a/w3191 ), .Z(n16134) );
  XOR \SUBBYTES[9].a/U5598  ( .A(\SUBBYTES[9].a/w3154 ), .B(
        \SUBBYTES[9].a/w3178 ), .Z(n16135) );
  XOR \SUBBYTES[9].a/U5597  ( .A(\SUBBYTES[9].a/w3143 ), .B(
        \SUBBYTES[9].a/w3152 ), .Z(n16136) );
  XOR \SUBBYTES[9].a/U5596  ( .A(\SUBBYTES[9].a/w3175 ), .B(n16137), .Z(n17151) );
  XOR \SUBBYTES[9].a/U5595  ( .A(\SUBBYTES[9].a/w3158 ), .B(
        \SUBBYTES[9].a/w3161 ), .Z(n16137) );
  XOR \SUBBYTES[9].a/U5594  ( .A(n17151), .B(n16138), .Z(n17347) );
  XOR \SUBBYTES[9].a/U5593  ( .A(\SUBBYTES[9].a/w3146 ), .B(n17153), .Z(n16138) );
  XOR \SUBBYTES[9].a/U5592  ( .A(n17149), .B(n16139), .Z(n17348) );
  XOR \SUBBYTES[9].a/U5591  ( .A(\SUBBYTES[9].a/w3178 ), .B(
        \SUBBYTES[9].a/w3191 ), .Z(n16139) );
  XOR \SUBBYTES[9].a/U5590  ( .A(n16141), .B(n16140), .Z(n17349) );
  XOR \SUBBYTES[9].a/U5589  ( .A(n16143), .B(n16142), .Z(n16140) );
  XOR \SUBBYTES[9].a/U5588  ( .A(n16145), .B(n16144), .Z(n16141) );
  XOR \SUBBYTES[9].a/U5587  ( .A(\SUBBYTES[9].a/w3190 ), .B(
        \SUBBYTES[9].a/w3193 ), .Z(n16142) );
  XOR \SUBBYTES[9].a/U5586  ( .A(\SUBBYTES[9].a/w3183 ), .B(
        \SUBBYTES[9].a/w3186 ), .Z(n16143) );
  XOR \SUBBYTES[9].a/U5585  ( .A(\SUBBYTES[9].a/w3158 ), .B(
        \SUBBYTES[9].a/w3159 ), .Z(n16144) );
  XOR \SUBBYTES[9].a/U5584  ( .A(\SUBBYTES[9].a/w3143 ), .B(
        \SUBBYTES[9].a/w3146 ), .Z(n16145) );
  XOR \SUBBYTES[9].a/U5583  ( .A(n16147), .B(n16146), .Z(n17350) );
  XOR \SUBBYTES[9].a/U5582  ( .A(n17150), .B(n16148), .Z(n16146) );
  XOR \SUBBYTES[9].a/U5581  ( .A(n17152), .B(n17151), .Z(n16147) );
  XOR \SUBBYTES[9].a/U5580  ( .A(\SUBBYTES[9].a/w3151 ), .B(
        \SUBBYTES[9].a/w3178 ), .Z(n16148) );
  XOR \SUBBYTES[9].a/U5579  ( .A(n16150), .B(n16149), .Z(n17351) );
  XOR \SUBBYTES[9].a/U5578  ( .A(n17153), .B(n16151), .Z(n16149) );
  XOR \SUBBYTES[9].a/U5577  ( .A(\SUBBYTES[9].a/w3184 ), .B(
        \SUBBYTES[9].a/w3186 ), .Z(n16150) );
  XOR \SUBBYTES[9].a/U5576  ( .A(\SUBBYTES[9].a/w3144 ), .B(
        \SUBBYTES[9].a/w3176 ), .Z(n16151) );
  XOR \SUBBYTES[9].a/U5575  ( .A(\SUBBYTES[9].a/w2976 ), .B(
        \SUBBYTES[9].a/w2977 ), .Z(n17155) );
  XOR \SUBBYTES[9].a/U5574  ( .A(n17155), .B(n16152), .Z(n17154) );
  XOR \SUBBYTES[9].a/U5573  ( .A(\SUBBYTES[9].a/w2969 ), .B(
        \SUBBYTES[9].a/w2986 ), .Z(n16152) );
  XOR \SUBBYTES[9].a/U5572  ( .A(n17154), .B(n16153), .Z(n17352) );
  XOR \SUBBYTES[9].a/U5571  ( .A(\SUBBYTES[9].a/w2968 ), .B(
        \SUBBYTES[9].a/w2983 ), .Z(n16153) );
  XOR \SUBBYTES[9].a/U5570  ( .A(n17155), .B(n16154), .Z(n17354) );
  XOR \SUBBYTES[9].a/U5569  ( .A(\SUBBYTES[9].a/w2983 ), .B(
        \SUBBYTES[9].a/w2984 ), .Z(n16154) );
  XOR \SUBBYTES[9].a/U5568  ( .A(\SUBBYTES[9].a/w2945 ), .B(n16155), .Z(n17157) );
  XOR \SUBBYTES[9].a/U5567  ( .A(\SUBBYTES[9].a/w2936 ), .B(
        \SUBBYTES[9].a/w2937 ), .Z(n16155) );
  XOR \SUBBYTES[9].a/U5566  ( .A(n17157), .B(n16156), .Z(n17353) );
  XOR \SUBBYTES[9].a/U5565  ( .A(\SUBBYTES[9].a/w2947 ), .B(n17354), .Z(n16156) );
  XOR \SUBBYTES[9].a/U5564  ( .A(n16158), .B(n16157), .Z(n17158) );
  XOR \SUBBYTES[9].a/U5563  ( .A(n16160), .B(n16159), .Z(n16157) );
  XOR \SUBBYTES[9].a/U5562  ( .A(\SUBBYTES[9].a/w2983 ), .B(
        \SUBBYTES[9].a/w2984 ), .Z(n16158) );
  XOR \SUBBYTES[9].a/U5561  ( .A(\SUBBYTES[9].a/w2947 ), .B(
        \SUBBYTES[9].a/w2971 ), .Z(n16159) );
  XOR \SUBBYTES[9].a/U5560  ( .A(\SUBBYTES[9].a/w2936 ), .B(
        \SUBBYTES[9].a/w2945 ), .Z(n16160) );
  XOR \SUBBYTES[9].a/U5559  ( .A(\SUBBYTES[9].a/w2968 ), .B(n16161), .Z(n17156) );
  XOR \SUBBYTES[9].a/U5558  ( .A(\SUBBYTES[9].a/w2951 ), .B(
        \SUBBYTES[9].a/w2954 ), .Z(n16161) );
  XOR \SUBBYTES[9].a/U5557  ( .A(n17156), .B(n16162), .Z(n17355) );
  XOR \SUBBYTES[9].a/U5556  ( .A(\SUBBYTES[9].a/w2939 ), .B(n17158), .Z(n16162) );
  XOR \SUBBYTES[9].a/U5555  ( .A(n17154), .B(n16163), .Z(n17356) );
  XOR \SUBBYTES[9].a/U5554  ( .A(\SUBBYTES[9].a/w2971 ), .B(
        \SUBBYTES[9].a/w2984 ), .Z(n16163) );
  XOR \SUBBYTES[9].a/U5553  ( .A(n16165), .B(n16164), .Z(n17357) );
  XOR \SUBBYTES[9].a/U5552  ( .A(n16167), .B(n16166), .Z(n16164) );
  XOR \SUBBYTES[9].a/U5551  ( .A(n16169), .B(n16168), .Z(n16165) );
  XOR \SUBBYTES[9].a/U5550  ( .A(\SUBBYTES[9].a/w2983 ), .B(
        \SUBBYTES[9].a/w2986 ), .Z(n16166) );
  XOR \SUBBYTES[9].a/U5549  ( .A(\SUBBYTES[9].a/w2976 ), .B(
        \SUBBYTES[9].a/w2979 ), .Z(n16167) );
  XOR \SUBBYTES[9].a/U5548  ( .A(\SUBBYTES[9].a/w2951 ), .B(
        \SUBBYTES[9].a/w2952 ), .Z(n16168) );
  XOR \SUBBYTES[9].a/U5547  ( .A(\SUBBYTES[9].a/w2936 ), .B(
        \SUBBYTES[9].a/w2939 ), .Z(n16169) );
  XOR \SUBBYTES[9].a/U5546  ( .A(n16171), .B(n16170), .Z(n17358) );
  XOR \SUBBYTES[9].a/U5545  ( .A(n17155), .B(n16172), .Z(n16170) );
  XOR \SUBBYTES[9].a/U5544  ( .A(n17157), .B(n17156), .Z(n16171) );
  XOR \SUBBYTES[9].a/U5543  ( .A(\SUBBYTES[9].a/w2944 ), .B(
        \SUBBYTES[9].a/w2971 ), .Z(n16172) );
  XOR \SUBBYTES[9].a/U5542  ( .A(n16174), .B(n16173), .Z(n17359) );
  XOR \SUBBYTES[9].a/U5541  ( .A(n17158), .B(n16175), .Z(n16173) );
  XOR \SUBBYTES[9].a/U5540  ( .A(\SUBBYTES[9].a/w2977 ), .B(
        \SUBBYTES[9].a/w2979 ), .Z(n16174) );
  XOR \SUBBYTES[9].a/U5539  ( .A(\SUBBYTES[9].a/w2937 ), .B(
        \SUBBYTES[9].a/w2969 ), .Z(n16175) );
  XOR \SUBBYTES[9].a/U5538  ( .A(\SUBBYTES[9].a/w2769 ), .B(
        \SUBBYTES[9].a/w2770 ), .Z(n17160) );
  XOR \SUBBYTES[9].a/U5537  ( .A(n17160), .B(n16176), .Z(n17159) );
  XOR \SUBBYTES[9].a/U5536  ( .A(\SUBBYTES[9].a/w2762 ), .B(
        \SUBBYTES[9].a/w2779 ), .Z(n16176) );
  XOR \SUBBYTES[9].a/U5535  ( .A(n17159), .B(n16177), .Z(n17360) );
  XOR \SUBBYTES[9].a/U5534  ( .A(\SUBBYTES[9].a/w2761 ), .B(
        \SUBBYTES[9].a/w2776 ), .Z(n16177) );
  XOR \SUBBYTES[9].a/U5533  ( .A(n17160), .B(n16178), .Z(n17362) );
  XOR \SUBBYTES[9].a/U5532  ( .A(\SUBBYTES[9].a/w2776 ), .B(
        \SUBBYTES[9].a/w2777 ), .Z(n16178) );
  XOR \SUBBYTES[9].a/U5531  ( .A(\SUBBYTES[9].a/w2738 ), .B(n16179), .Z(n17162) );
  XOR \SUBBYTES[9].a/U5530  ( .A(\SUBBYTES[9].a/w2729 ), .B(
        \SUBBYTES[9].a/w2730 ), .Z(n16179) );
  XOR \SUBBYTES[9].a/U5529  ( .A(n17162), .B(n16180), .Z(n17361) );
  XOR \SUBBYTES[9].a/U5528  ( .A(\SUBBYTES[9].a/w2740 ), .B(n17362), .Z(n16180) );
  XOR \SUBBYTES[9].a/U5527  ( .A(n16182), .B(n16181), .Z(n17163) );
  XOR \SUBBYTES[9].a/U5526  ( .A(n16184), .B(n16183), .Z(n16181) );
  XOR \SUBBYTES[9].a/U5525  ( .A(\SUBBYTES[9].a/w2776 ), .B(
        \SUBBYTES[9].a/w2777 ), .Z(n16182) );
  XOR \SUBBYTES[9].a/U5524  ( .A(\SUBBYTES[9].a/w2740 ), .B(
        \SUBBYTES[9].a/w2764 ), .Z(n16183) );
  XOR \SUBBYTES[9].a/U5523  ( .A(\SUBBYTES[9].a/w2729 ), .B(
        \SUBBYTES[9].a/w2738 ), .Z(n16184) );
  XOR \SUBBYTES[9].a/U5522  ( .A(\SUBBYTES[9].a/w2761 ), .B(n16185), .Z(n17161) );
  XOR \SUBBYTES[9].a/U5521  ( .A(\SUBBYTES[9].a/w2744 ), .B(
        \SUBBYTES[9].a/w2747 ), .Z(n16185) );
  XOR \SUBBYTES[9].a/U5520  ( .A(n17161), .B(n16186), .Z(n17363) );
  XOR \SUBBYTES[9].a/U5519  ( .A(\SUBBYTES[9].a/w2732 ), .B(n17163), .Z(n16186) );
  XOR \SUBBYTES[9].a/U5518  ( .A(n17159), .B(n16187), .Z(n17364) );
  XOR \SUBBYTES[9].a/U5517  ( .A(\SUBBYTES[9].a/w2764 ), .B(
        \SUBBYTES[9].a/w2777 ), .Z(n16187) );
  XOR \SUBBYTES[9].a/U5516  ( .A(n16189), .B(n16188), .Z(n17365) );
  XOR \SUBBYTES[9].a/U5515  ( .A(n16191), .B(n16190), .Z(n16188) );
  XOR \SUBBYTES[9].a/U5514  ( .A(n16193), .B(n16192), .Z(n16189) );
  XOR \SUBBYTES[9].a/U5513  ( .A(\SUBBYTES[9].a/w2776 ), .B(
        \SUBBYTES[9].a/w2779 ), .Z(n16190) );
  XOR \SUBBYTES[9].a/U5512  ( .A(\SUBBYTES[9].a/w2769 ), .B(
        \SUBBYTES[9].a/w2772 ), .Z(n16191) );
  XOR \SUBBYTES[9].a/U5511  ( .A(\SUBBYTES[9].a/w2744 ), .B(
        \SUBBYTES[9].a/w2745 ), .Z(n16192) );
  XOR \SUBBYTES[9].a/U5510  ( .A(\SUBBYTES[9].a/w2729 ), .B(
        \SUBBYTES[9].a/w2732 ), .Z(n16193) );
  XOR \SUBBYTES[9].a/U5509  ( .A(n16195), .B(n16194), .Z(n17366) );
  XOR \SUBBYTES[9].a/U5508  ( .A(n17160), .B(n16196), .Z(n16194) );
  XOR \SUBBYTES[9].a/U5507  ( .A(n17162), .B(n17161), .Z(n16195) );
  XOR \SUBBYTES[9].a/U5506  ( .A(\SUBBYTES[9].a/w2737 ), .B(
        \SUBBYTES[9].a/w2764 ), .Z(n16196) );
  XOR \SUBBYTES[9].a/U5505  ( .A(n16198), .B(n16197), .Z(n17367) );
  XOR \SUBBYTES[9].a/U5504  ( .A(n17163), .B(n16199), .Z(n16197) );
  XOR \SUBBYTES[9].a/U5503  ( .A(\SUBBYTES[9].a/w2770 ), .B(
        \SUBBYTES[9].a/w2772 ), .Z(n16198) );
  XOR \SUBBYTES[9].a/U5502  ( .A(\SUBBYTES[9].a/w2730 ), .B(
        \SUBBYTES[9].a/w2762 ), .Z(n16199) );
  XOR \SUBBYTES[9].a/U5501  ( .A(\SUBBYTES[9].a/w2562 ), .B(
        \SUBBYTES[9].a/w2563 ), .Z(n17165) );
  XOR \SUBBYTES[9].a/U5500  ( .A(n17165), .B(n16200), .Z(n17164) );
  XOR \SUBBYTES[9].a/U5499  ( .A(\SUBBYTES[9].a/w2555 ), .B(
        \SUBBYTES[9].a/w2572 ), .Z(n16200) );
  XOR \SUBBYTES[9].a/U5498  ( .A(n17164), .B(n16201), .Z(n17368) );
  XOR \SUBBYTES[9].a/U5497  ( .A(\SUBBYTES[9].a/w2554 ), .B(
        \SUBBYTES[9].a/w2569 ), .Z(n16201) );
  XOR \SUBBYTES[9].a/U5496  ( .A(n17165), .B(n16202), .Z(n17370) );
  XOR \SUBBYTES[9].a/U5495  ( .A(\SUBBYTES[9].a/w2569 ), .B(
        \SUBBYTES[9].a/w2570 ), .Z(n16202) );
  XOR \SUBBYTES[9].a/U5494  ( .A(\SUBBYTES[9].a/w2531 ), .B(n16203), .Z(n17167) );
  XOR \SUBBYTES[9].a/U5493  ( .A(\SUBBYTES[9].a/w2522 ), .B(
        \SUBBYTES[9].a/w2523 ), .Z(n16203) );
  XOR \SUBBYTES[9].a/U5492  ( .A(n17167), .B(n16204), .Z(n17369) );
  XOR \SUBBYTES[9].a/U5491  ( .A(\SUBBYTES[9].a/w2533 ), .B(n17370), .Z(n16204) );
  XOR \SUBBYTES[9].a/U5490  ( .A(n16206), .B(n16205), .Z(n17168) );
  XOR \SUBBYTES[9].a/U5489  ( .A(n16208), .B(n16207), .Z(n16205) );
  XOR \SUBBYTES[9].a/U5488  ( .A(\SUBBYTES[9].a/w2569 ), .B(
        \SUBBYTES[9].a/w2570 ), .Z(n16206) );
  XOR \SUBBYTES[9].a/U5487  ( .A(\SUBBYTES[9].a/w2533 ), .B(
        \SUBBYTES[9].a/w2557 ), .Z(n16207) );
  XOR \SUBBYTES[9].a/U5486  ( .A(\SUBBYTES[9].a/w2522 ), .B(
        \SUBBYTES[9].a/w2531 ), .Z(n16208) );
  XOR \SUBBYTES[9].a/U5485  ( .A(\SUBBYTES[9].a/w2554 ), .B(n16209), .Z(n17166) );
  XOR \SUBBYTES[9].a/U5484  ( .A(\SUBBYTES[9].a/w2537 ), .B(
        \SUBBYTES[9].a/w2540 ), .Z(n16209) );
  XOR \SUBBYTES[9].a/U5483  ( .A(n17166), .B(n16210), .Z(n17371) );
  XOR \SUBBYTES[9].a/U5482  ( .A(\SUBBYTES[9].a/w2525 ), .B(n17168), .Z(n16210) );
  XOR \SUBBYTES[9].a/U5481  ( .A(n17164), .B(n16211), .Z(n17372) );
  XOR \SUBBYTES[9].a/U5480  ( .A(\SUBBYTES[9].a/w2557 ), .B(
        \SUBBYTES[9].a/w2570 ), .Z(n16211) );
  XOR \SUBBYTES[9].a/U5479  ( .A(n16213), .B(n16212), .Z(n17373) );
  XOR \SUBBYTES[9].a/U5478  ( .A(n16215), .B(n16214), .Z(n16212) );
  XOR \SUBBYTES[9].a/U5477  ( .A(n16217), .B(n16216), .Z(n16213) );
  XOR \SUBBYTES[9].a/U5476  ( .A(\SUBBYTES[9].a/w2569 ), .B(
        \SUBBYTES[9].a/w2572 ), .Z(n16214) );
  XOR \SUBBYTES[9].a/U5475  ( .A(\SUBBYTES[9].a/w2562 ), .B(
        \SUBBYTES[9].a/w2565 ), .Z(n16215) );
  XOR \SUBBYTES[9].a/U5474  ( .A(\SUBBYTES[9].a/w2537 ), .B(
        \SUBBYTES[9].a/w2538 ), .Z(n16216) );
  XOR \SUBBYTES[9].a/U5473  ( .A(\SUBBYTES[9].a/w2522 ), .B(
        \SUBBYTES[9].a/w2525 ), .Z(n16217) );
  XOR \SUBBYTES[9].a/U5472  ( .A(n16219), .B(n16218), .Z(n17374) );
  XOR \SUBBYTES[9].a/U5471  ( .A(n17165), .B(n16220), .Z(n16218) );
  XOR \SUBBYTES[9].a/U5470  ( .A(n17167), .B(n17166), .Z(n16219) );
  XOR \SUBBYTES[9].a/U5469  ( .A(\SUBBYTES[9].a/w2530 ), .B(
        \SUBBYTES[9].a/w2557 ), .Z(n16220) );
  XOR \SUBBYTES[9].a/U5468  ( .A(n16222), .B(n16221), .Z(n17375) );
  XOR \SUBBYTES[9].a/U5467  ( .A(n17168), .B(n16223), .Z(n16221) );
  XOR \SUBBYTES[9].a/U5466  ( .A(\SUBBYTES[9].a/w2563 ), .B(
        \SUBBYTES[9].a/w2565 ), .Z(n16222) );
  XOR \SUBBYTES[9].a/U5465  ( .A(\SUBBYTES[9].a/w2523 ), .B(
        \SUBBYTES[9].a/w2555 ), .Z(n16223) );
  XOR \SUBBYTES[9].a/U5464  ( .A(\SUBBYTES[9].a/w2355 ), .B(
        \SUBBYTES[9].a/w2356 ), .Z(n17170) );
  XOR \SUBBYTES[9].a/U5463  ( .A(n17170), .B(n16224), .Z(n17169) );
  XOR \SUBBYTES[9].a/U5462  ( .A(\SUBBYTES[9].a/w2348 ), .B(
        \SUBBYTES[9].a/w2365 ), .Z(n16224) );
  XOR \SUBBYTES[9].a/U5461  ( .A(n17169), .B(n16225), .Z(n17376) );
  XOR \SUBBYTES[9].a/U5460  ( .A(\SUBBYTES[9].a/w2347 ), .B(
        \SUBBYTES[9].a/w2362 ), .Z(n16225) );
  XOR \SUBBYTES[9].a/U5459  ( .A(n17170), .B(n16226), .Z(n17378) );
  XOR \SUBBYTES[9].a/U5458  ( .A(\SUBBYTES[9].a/w2362 ), .B(
        \SUBBYTES[9].a/w2363 ), .Z(n16226) );
  XOR \SUBBYTES[9].a/U5457  ( .A(\SUBBYTES[9].a/w2324 ), .B(n16227), .Z(n17172) );
  XOR \SUBBYTES[9].a/U5456  ( .A(\SUBBYTES[9].a/w2315 ), .B(
        \SUBBYTES[9].a/w2316 ), .Z(n16227) );
  XOR \SUBBYTES[9].a/U5455  ( .A(n17172), .B(n16228), .Z(n17377) );
  XOR \SUBBYTES[9].a/U5454  ( .A(\SUBBYTES[9].a/w2326 ), .B(n17378), .Z(n16228) );
  XOR \SUBBYTES[9].a/U5453  ( .A(n16230), .B(n16229), .Z(n17173) );
  XOR \SUBBYTES[9].a/U5452  ( .A(n16232), .B(n16231), .Z(n16229) );
  XOR \SUBBYTES[9].a/U5451  ( .A(\SUBBYTES[9].a/w2362 ), .B(
        \SUBBYTES[9].a/w2363 ), .Z(n16230) );
  XOR \SUBBYTES[9].a/U5450  ( .A(\SUBBYTES[9].a/w2326 ), .B(
        \SUBBYTES[9].a/w2350 ), .Z(n16231) );
  XOR \SUBBYTES[9].a/U5449  ( .A(\SUBBYTES[9].a/w2315 ), .B(
        \SUBBYTES[9].a/w2324 ), .Z(n16232) );
  XOR \SUBBYTES[9].a/U5448  ( .A(\SUBBYTES[9].a/w2347 ), .B(n16233), .Z(n17171) );
  XOR \SUBBYTES[9].a/U5447  ( .A(\SUBBYTES[9].a/w2330 ), .B(
        \SUBBYTES[9].a/w2333 ), .Z(n16233) );
  XOR \SUBBYTES[9].a/U5446  ( .A(n17171), .B(n16234), .Z(n17379) );
  XOR \SUBBYTES[9].a/U5445  ( .A(\SUBBYTES[9].a/w2318 ), .B(n17173), .Z(n16234) );
  XOR \SUBBYTES[9].a/U5444  ( .A(n17169), .B(n16235), .Z(n17380) );
  XOR \SUBBYTES[9].a/U5443  ( .A(\SUBBYTES[9].a/w2350 ), .B(
        \SUBBYTES[9].a/w2363 ), .Z(n16235) );
  XOR \SUBBYTES[9].a/U5442  ( .A(n16237), .B(n16236), .Z(n17381) );
  XOR \SUBBYTES[9].a/U5441  ( .A(n16239), .B(n16238), .Z(n16236) );
  XOR \SUBBYTES[9].a/U5440  ( .A(n16241), .B(n16240), .Z(n16237) );
  XOR \SUBBYTES[9].a/U5439  ( .A(\SUBBYTES[9].a/w2362 ), .B(
        \SUBBYTES[9].a/w2365 ), .Z(n16238) );
  XOR \SUBBYTES[9].a/U5438  ( .A(\SUBBYTES[9].a/w2355 ), .B(
        \SUBBYTES[9].a/w2358 ), .Z(n16239) );
  XOR \SUBBYTES[9].a/U5437  ( .A(\SUBBYTES[9].a/w2330 ), .B(
        \SUBBYTES[9].a/w2331 ), .Z(n16240) );
  XOR \SUBBYTES[9].a/U5436  ( .A(\SUBBYTES[9].a/w2315 ), .B(
        \SUBBYTES[9].a/w2318 ), .Z(n16241) );
  XOR \SUBBYTES[9].a/U5435  ( .A(n16243), .B(n16242), .Z(n17382) );
  XOR \SUBBYTES[9].a/U5434  ( .A(n17170), .B(n16244), .Z(n16242) );
  XOR \SUBBYTES[9].a/U5433  ( .A(n17172), .B(n17171), .Z(n16243) );
  XOR \SUBBYTES[9].a/U5432  ( .A(\SUBBYTES[9].a/w2323 ), .B(
        \SUBBYTES[9].a/w2350 ), .Z(n16244) );
  XOR \SUBBYTES[9].a/U5431  ( .A(n16246), .B(n16245), .Z(n17383) );
  XOR \SUBBYTES[9].a/U5430  ( .A(n17173), .B(n16247), .Z(n16245) );
  XOR \SUBBYTES[9].a/U5429  ( .A(\SUBBYTES[9].a/w2356 ), .B(
        \SUBBYTES[9].a/w2358 ), .Z(n16246) );
  XOR \SUBBYTES[9].a/U5428  ( .A(\SUBBYTES[9].a/w2316 ), .B(
        \SUBBYTES[9].a/w2348 ), .Z(n16247) );
  XOR \SUBBYTES[9].a/U5427  ( .A(\SUBBYTES[9].a/w2148 ), .B(
        \SUBBYTES[9].a/w2149 ), .Z(n17175) );
  XOR \SUBBYTES[9].a/U5426  ( .A(n17175), .B(n16248), .Z(n17174) );
  XOR \SUBBYTES[9].a/U5425  ( .A(\SUBBYTES[9].a/w2141 ), .B(
        \SUBBYTES[9].a/w2158 ), .Z(n16248) );
  XOR \SUBBYTES[9].a/U5424  ( .A(n17174), .B(n16249), .Z(n17384) );
  XOR \SUBBYTES[9].a/U5423  ( .A(\SUBBYTES[9].a/w2140 ), .B(
        \SUBBYTES[9].a/w2155 ), .Z(n16249) );
  XOR \SUBBYTES[9].a/U5422  ( .A(n17175), .B(n16250), .Z(n17386) );
  XOR \SUBBYTES[9].a/U5421  ( .A(\SUBBYTES[9].a/w2155 ), .B(
        \SUBBYTES[9].a/w2156 ), .Z(n16250) );
  XOR \SUBBYTES[9].a/U5420  ( .A(\SUBBYTES[9].a/w2117 ), .B(n16251), .Z(n17177) );
  XOR \SUBBYTES[9].a/U5419  ( .A(\SUBBYTES[9].a/w2108 ), .B(
        \SUBBYTES[9].a/w2109 ), .Z(n16251) );
  XOR \SUBBYTES[9].a/U5418  ( .A(n17177), .B(n16252), .Z(n17385) );
  XOR \SUBBYTES[9].a/U5417  ( .A(\SUBBYTES[9].a/w2119 ), .B(n17386), .Z(n16252) );
  XOR \SUBBYTES[9].a/U5416  ( .A(n16254), .B(n16253), .Z(n17178) );
  XOR \SUBBYTES[9].a/U5415  ( .A(n16256), .B(n16255), .Z(n16253) );
  XOR \SUBBYTES[9].a/U5414  ( .A(\SUBBYTES[9].a/w2155 ), .B(
        \SUBBYTES[9].a/w2156 ), .Z(n16254) );
  XOR \SUBBYTES[9].a/U5413  ( .A(\SUBBYTES[9].a/w2119 ), .B(
        \SUBBYTES[9].a/w2143 ), .Z(n16255) );
  XOR \SUBBYTES[9].a/U5412  ( .A(\SUBBYTES[9].a/w2108 ), .B(
        \SUBBYTES[9].a/w2117 ), .Z(n16256) );
  XOR \SUBBYTES[9].a/U5411  ( .A(\SUBBYTES[9].a/w2140 ), .B(n16257), .Z(n17176) );
  XOR \SUBBYTES[9].a/U5410  ( .A(\SUBBYTES[9].a/w2123 ), .B(
        \SUBBYTES[9].a/w2126 ), .Z(n16257) );
  XOR \SUBBYTES[9].a/U5409  ( .A(n17176), .B(n16258), .Z(n17387) );
  XOR \SUBBYTES[9].a/U5408  ( .A(\SUBBYTES[9].a/w2111 ), .B(n17178), .Z(n16258) );
  XOR \SUBBYTES[9].a/U5407  ( .A(n17174), .B(n16259), .Z(n17388) );
  XOR \SUBBYTES[9].a/U5406  ( .A(\SUBBYTES[9].a/w2143 ), .B(
        \SUBBYTES[9].a/w2156 ), .Z(n16259) );
  XOR \SUBBYTES[9].a/U5405  ( .A(n16261), .B(n16260), .Z(n17389) );
  XOR \SUBBYTES[9].a/U5404  ( .A(n16263), .B(n16262), .Z(n16260) );
  XOR \SUBBYTES[9].a/U5403  ( .A(n16265), .B(n16264), .Z(n16261) );
  XOR \SUBBYTES[9].a/U5402  ( .A(\SUBBYTES[9].a/w2155 ), .B(
        \SUBBYTES[9].a/w2158 ), .Z(n16262) );
  XOR \SUBBYTES[9].a/U5401  ( .A(\SUBBYTES[9].a/w2148 ), .B(
        \SUBBYTES[9].a/w2151 ), .Z(n16263) );
  XOR \SUBBYTES[9].a/U5400  ( .A(\SUBBYTES[9].a/w2123 ), .B(
        \SUBBYTES[9].a/w2124 ), .Z(n16264) );
  XOR \SUBBYTES[9].a/U5399  ( .A(\SUBBYTES[9].a/w2108 ), .B(
        \SUBBYTES[9].a/w2111 ), .Z(n16265) );
  XOR \SUBBYTES[9].a/U5398  ( .A(n16267), .B(n16266), .Z(n17390) );
  XOR \SUBBYTES[9].a/U5397  ( .A(n17175), .B(n16268), .Z(n16266) );
  XOR \SUBBYTES[9].a/U5396  ( .A(n17177), .B(n17176), .Z(n16267) );
  XOR \SUBBYTES[9].a/U5395  ( .A(\SUBBYTES[9].a/w2116 ), .B(
        \SUBBYTES[9].a/w2143 ), .Z(n16268) );
  XOR \SUBBYTES[9].a/U5394  ( .A(n16270), .B(n16269), .Z(n17391) );
  XOR \SUBBYTES[9].a/U5393  ( .A(n17178), .B(n16271), .Z(n16269) );
  XOR \SUBBYTES[9].a/U5392  ( .A(\SUBBYTES[9].a/w2149 ), .B(
        \SUBBYTES[9].a/w2151 ), .Z(n16270) );
  XOR \SUBBYTES[9].a/U5391  ( .A(\SUBBYTES[9].a/w2109 ), .B(
        \SUBBYTES[9].a/w2141 ), .Z(n16271) );
  XOR \SUBBYTES[9].a/U5390  ( .A(\SUBBYTES[9].a/w1941 ), .B(
        \SUBBYTES[9].a/w1942 ), .Z(n17180) );
  XOR \SUBBYTES[9].a/U5389  ( .A(n17180), .B(n16272), .Z(n17179) );
  XOR \SUBBYTES[9].a/U5388  ( .A(\SUBBYTES[9].a/w1934 ), .B(
        \SUBBYTES[9].a/w1951 ), .Z(n16272) );
  XOR \SUBBYTES[9].a/U5387  ( .A(n17179), .B(n16273), .Z(n17392) );
  XOR \SUBBYTES[9].a/U5386  ( .A(\SUBBYTES[9].a/w1933 ), .B(
        \SUBBYTES[9].a/w1948 ), .Z(n16273) );
  XOR \SUBBYTES[9].a/U5385  ( .A(n17180), .B(n16274), .Z(n17394) );
  XOR \SUBBYTES[9].a/U5384  ( .A(\SUBBYTES[9].a/w1948 ), .B(
        \SUBBYTES[9].a/w1949 ), .Z(n16274) );
  XOR \SUBBYTES[9].a/U5383  ( .A(\SUBBYTES[9].a/w1910 ), .B(n16275), .Z(n17182) );
  XOR \SUBBYTES[9].a/U5382  ( .A(\SUBBYTES[9].a/w1901 ), .B(
        \SUBBYTES[9].a/w1902 ), .Z(n16275) );
  XOR \SUBBYTES[9].a/U5381  ( .A(n17182), .B(n16276), .Z(n17393) );
  XOR \SUBBYTES[9].a/U5380  ( .A(\SUBBYTES[9].a/w1912 ), .B(n17394), .Z(n16276) );
  XOR \SUBBYTES[9].a/U5379  ( .A(n16278), .B(n16277), .Z(n17183) );
  XOR \SUBBYTES[9].a/U5378  ( .A(n16280), .B(n16279), .Z(n16277) );
  XOR \SUBBYTES[9].a/U5377  ( .A(\SUBBYTES[9].a/w1948 ), .B(
        \SUBBYTES[9].a/w1949 ), .Z(n16278) );
  XOR \SUBBYTES[9].a/U5376  ( .A(\SUBBYTES[9].a/w1912 ), .B(
        \SUBBYTES[9].a/w1936 ), .Z(n16279) );
  XOR \SUBBYTES[9].a/U5375  ( .A(\SUBBYTES[9].a/w1901 ), .B(
        \SUBBYTES[9].a/w1910 ), .Z(n16280) );
  XOR \SUBBYTES[9].a/U5374  ( .A(\SUBBYTES[9].a/w1933 ), .B(n16281), .Z(n17181) );
  XOR \SUBBYTES[9].a/U5373  ( .A(\SUBBYTES[9].a/w1916 ), .B(
        \SUBBYTES[9].a/w1919 ), .Z(n16281) );
  XOR \SUBBYTES[9].a/U5372  ( .A(n17181), .B(n16282), .Z(n17395) );
  XOR \SUBBYTES[9].a/U5371  ( .A(\SUBBYTES[9].a/w1904 ), .B(n17183), .Z(n16282) );
  XOR \SUBBYTES[9].a/U5370  ( .A(n17179), .B(n16283), .Z(n17396) );
  XOR \SUBBYTES[9].a/U5369  ( .A(\SUBBYTES[9].a/w1936 ), .B(
        \SUBBYTES[9].a/w1949 ), .Z(n16283) );
  XOR \SUBBYTES[9].a/U5368  ( .A(n16285), .B(n16284), .Z(n17397) );
  XOR \SUBBYTES[9].a/U5367  ( .A(n16287), .B(n16286), .Z(n16284) );
  XOR \SUBBYTES[9].a/U5366  ( .A(n16289), .B(n16288), .Z(n16285) );
  XOR \SUBBYTES[9].a/U5365  ( .A(\SUBBYTES[9].a/w1948 ), .B(
        \SUBBYTES[9].a/w1951 ), .Z(n16286) );
  XOR \SUBBYTES[9].a/U5364  ( .A(\SUBBYTES[9].a/w1941 ), .B(
        \SUBBYTES[9].a/w1944 ), .Z(n16287) );
  XOR \SUBBYTES[9].a/U5363  ( .A(\SUBBYTES[9].a/w1916 ), .B(
        \SUBBYTES[9].a/w1917 ), .Z(n16288) );
  XOR \SUBBYTES[9].a/U5362  ( .A(\SUBBYTES[9].a/w1901 ), .B(
        \SUBBYTES[9].a/w1904 ), .Z(n16289) );
  XOR \SUBBYTES[9].a/U5361  ( .A(n16291), .B(n16290), .Z(n17398) );
  XOR \SUBBYTES[9].a/U5360  ( .A(n17180), .B(n16292), .Z(n16290) );
  XOR \SUBBYTES[9].a/U5359  ( .A(n17182), .B(n17181), .Z(n16291) );
  XOR \SUBBYTES[9].a/U5358  ( .A(\SUBBYTES[9].a/w1909 ), .B(
        \SUBBYTES[9].a/w1936 ), .Z(n16292) );
  XOR \SUBBYTES[9].a/U5357  ( .A(n16294), .B(n16293), .Z(n17399) );
  XOR \SUBBYTES[9].a/U5356  ( .A(n17183), .B(n16295), .Z(n16293) );
  XOR \SUBBYTES[9].a/U5355  ( .A(\SUBBYTES[9].a/w1942 ), .B(
        \SUBBYTES[9].a/w1944 ), .Z(n16294) );
  XOR \SUBBYTES[9].a/U5354  ( .A(\SUBBYTES[9].a/w1902 ), .B(
        \SUBBYTES[9].a/w1934 ), .Z(n16295) );
  XOR \SUBBYTES[9].a/U5353  ( .A(\SUBBYTES[9].a/w1734 ), .B(
        \SUBBYTES[9].a/w1735 ), .Z(n17185) );
  XOR \SUBBYTES[9].a/U5352  ( .A(n17185), .B(n16296), .Z(n17184) );
  XOR \SUBBYTES[9].a/U5351  ( .A(\SUBBYTES[9].a/w1727 ), .B(
        \SUBBYTES[9].a/w1744 ), .Z(n16296) );
  XOR \SUBBYTES[9].a/U5350  ( .A(n17184), .B(n16297), .Z(n17400) );
  XOR \SUBBYTES[9].a/U5349  ( .A(\SUBBYTES[9].a/w1726 ), .B(
        \SUBBYTES[9].a/w1741 ), .Z(n16297) );
  XOR \SUBBYTES[9].a/U5348  ( .A(n17185), .B(n16298), .Z(n17402) );
  XOR \SUBBYTES[9].a/U5347  ( .A(\SUBBYTES[9].a/w1741 ), .B(
        \SUBBYTES[9].a/w1742 ), .Z(n16298) );
  XOR \SUBBYTES[9].a/U5346  ( .A(\SUBBYTES[9].a/w1703 ), .B(n16299), .Z(n17187) );
  XOR \SUBBYTES[9].a/U5345  ( .A(\SUBBYTES[9].a/w1694 ), .B(
        \SUBBYTES[9].a/w1695 ), .Z(n16299) );
  XOR \SUBBYTES[9].a/U5344  ( .A(n17187), .B(n16300), .Z(n17401) );
  XOR \SUBBYTES[9].a/U5343  ( .A(\SUBBYTES[9].a/w1705 ), .B(n17402), .Z(n16300) );
  XOR \SUBBYTES[9].a/U5342  ( .A(n16302), .B(n16301), .Z(n17188) );
  XOR \SUBBYTES[9].a/U5341  ( .A(n16304), .B(n16303), .Z(n16301) );
  XOR \SUBBYTES[9].a/U5340  ( .A(\SUBBYTES[9].a/w1741 ), .B(
        \SUBBYTES[9].a/w1742 ), .Z(n16302) );
  XOR \SUBBYTES[9].a/U5339  ( .A(\SUBBYTES[9].a/w1705 ), .B(
        \SUBBYTES[9].a/w1729 ), .Z(n16303) );
  XOR \SUBBYTES[9].a/U5338  ( .A(\SUBBYTES[9].a/w1694 ), .B(
        \SUBBYTES[9].a/w1703 ), .Z(n16304) );
  XOR \SUBBYTES[9].a/U5337  ( .A(\SUBBYTES[9].a/w1726 ), .B(n16305), .Z(n17186) );
  XOR \SUBBYTES[9].a/U5336  ( .A(\SUBBYTES[9].a/w1709 ), .B(
        \SUBBYTES[9].a/w1712 ), .Z(n16305) );
  XOR \SUBBYTES[9].a/U5335  ( .A(n17186), .B(n16306), .Z(n17403) );
  XOR \SUBBYTES[9].a/U5334  ( .A(\SUBBYTES[9].a/w1697 ), .B(n17188), .Z(n16306) );
  XOR \SUBBYTES[9].a/U5333  ( .A(n17184), .B(n16307), .Z(n17404) );
  XOR \SUBBYTES[9].a/U5332  ( .A(\SUBBYTES[9].a/w1729 ), .B(
        \SUBBYTES[9].a/w1742 ), .Z(n16307) );
  XOR \SUBBYTES[9].a/U5331  ( .A(n16309), .B(n16308), .Z(n17405) );
  XOR \SUBBYTES[9].a/U5330  ( .A(n16311), .B(n16310), .Z(n16308) );
  XOR \SUBBYTES[9].a/U5329  ( .A(n16313), .B(n16312), .Z(n16309) );
  XOR \SUBBYTES[9].a/U5328  ( .A(\SUBBYTES[9].a/w1741 ), .B(
        \SUBBYTES[9].a/w1744 ), .Z(n16310) );
  XOR \SUBBYTES[9].a/U5327  ( .A(\SUBBYTES[9].a/w1734 ), .B(
        \SUBBYTES[9].a/w1737 ), .Z(n16311) );
  XOR \SUBBYTES[9].a/U5326  ( .A(\SUBBYTES[9].a/w1709 ), .B(
        \SUBBYTES[9].a/w1710 ), .Z(n16312) );
  XOR \SUBBYTES[9].a/U5325  ( .A(\SUBBYTES[9].a/w1694 ), .B(
        \SUBBYTES[9].a/w1697 ), .Z(n16313) );
  XOR \SUBBYTES[9].a/U5324  ( .A(n16315), .B(n16314), .Z(n17406) );
  XOR \SUBBYTES[9].a/U5323  ( .A(n17185), .B(n16316), .Z(n16314) );
  XOR \SUBBYTES[9].a/U5322  ( .A(n17187), .B(n17186), .Z(n16315) );
  XOR \SUBBYTES[9].a/U5321  ( .A(\SUBBYTES[9].a/w1702 ), .B(
        \SUBBYTES[9].a/w1729 ), .Z(n16316) );
  XOR \SUBBYTES[9].a/U5320  ( .A(n16318), .B(n16317), .Z(n17407) );
  XOR \SUBBYTES[9].a/U5319  ( .A(n17188), .B(n16319), .Z(n16317) );
  XOR \SUBBYTES[9].a/U5318  ( .A(\SUBBYTES[9].a/w1735 ), .B(
        \SUBBYTES[9].a/w1737 ), .Z(n16318) );
  XOR \SUBBYTES[9].a/U5317  ( .A(\SUBBYTES[9].a/w1695 ), .B(
        \SUBBYTES[9].a/w1727 ), .Z(n16319) );
  XOR \SUBBYTES[9].a/U5316  ( .A(\SUBBYTES[9].a/w1527 ), .B(
        \SUBBYTES[9].a/w1528 ), .Z(n17190) );
  XOR \SUBBYTES[9].a/U5315  ( .A(n17190), .B(n16320), .Z(n17189) );
  XOR \SUBBYTES[9].a/U5314  ( .A(\SUBBYTES[9].a/w1520 ), .B(
        \SUBBYTES[9].a/w1537 ), .Z(n16320) );
  XOR \SUBBYTES[9].a/U5313  ( .A(n17189), .B(n16321), .Z(n17408) );
  XOR \SUBBYTES[9].a/U5312  ( .A(\SUBBYTES[9].a/w1519 ), .B(
        \SUBBYTES[9].a/w1534 ), .Z(n16321) );
  XOR \SUBBYTES[9].a/U5311  ( .A(n17190), .B(n16322), .Z(n17410) );
  XOR \SUBBYTES[9].a/U5310  ( .A(\SUBBYTES[9].a/w1534 ), .B(
        \SUBBYTES[9].a/w1535 ), .Z(n16322) );
  XOR \SUBBYTES[9].a/U5309  ( .A(\SUBBYTES[9].a/w1496 ), .B(n16323), .Z(n17192) );
  XOR \SUBBYTES[9].a/U5308  ( .A(\SUBBYTES[9].a/w1487 ), .B(
        \SUBBYTES[9].a/w1488 ), .Z(n16323) );
  XOR \SUBBYTES[9].a/U5307  ( .A(n17192), .B(n16324), .Z(n17409) );
  XOR \SUBBYTES[9].a/U5306  ( .A(\SUBBYTES[9].a/w1498 ), .B(n17410), .Z(n16324) );
  XOR \SUBBYTES[9].a/U5305  ( .A(n16326), .B(n16325), .Z(n17193) );
  XOR \SUBBYTES[9].a/U5304  ( .A(n16328), .B(n16327), .Z(n16325) );
  XOR \SUBBYTES[9].a/U5303  ( .A(\SUBBYTES[9].a/w1534 ), .B(
        \SUBBYTES[9].a/w1535 ), .Z(n16326) );
  XOR \SUBBYTES[9].a/U5302  ( .A(\SUBBYTES[9].a/w1498 ), .B(
        \SUBBYTES[9].a/w1522 ), .Z(n16327) );
  XOR \SUBBYTES[9].a/U5301  ( .A(\SUBBYTES[9].a/w1487 ), .B(
        \SUBBYTES[9].a/w1496 ), .Z(n16328) );
  XOR \SUBBYTES[9].a/U5300  ( .A(\SUBBYTES[9].a/w1519 ), .B(n16329), .Z(n17191) );
  XOR \SUBBYTES[9].a/U5299  ( .A(\SUBBYTES[9].a/w1502 ), .B(
        \SUBBYTES[9].a/w1505 ), .Z(n16329) );
  XOR \SUBBYTES[9].a/U5298  ( .A(n17191), .B(n16330), .Z(n17411) );
  XOR \SUBBYTES[9].a/U5297  ( .A(\SUBBYTES[9].a/w1490 ), .B(n17193), .Z(n16330) );
  XOR \SUBBYTES[9].a/U5296  ( .A(n17189), .B(n16331), .Z(n17412) );
  XOR \SUBBYTES[9].a/U5295  ( .A(\SUBBYTES[9].a/w1522 ), .B(
        \SUBBYTES[9].a/w1535 ), .Z(n16331) );
  XOR \SUBBYTES[9].a/U5294  ( .A(n16333), .B(n16332), .Z(n17413) );
  XOR \SUBBYTES[9].a/U5293  ( .A(n16335), .B(n16334), .Z(n16332) );
  XOR \SUBBYTES[9].a/U5292  ( .A(n16337), .B(n16336), .Z(n16333) );
  XOR \SUBBYTES[9].a/U5291  ( .A(\SUBBYTES[9].a/w1534 ), .B(
        \SUBBYTES[9].a/w1537 ), .Z(n16334) );
  XOR \SUBBYTES[9].a/U5290  ( .A(\SUBBYTES[9].a/w1527 ), .B(
        \SUBBYTES[9].a/w1530 ), .Z(n16335) );
  XOR \SUBBYTES[9].a/U5289  ( .A(\SUBBYTES[9].a/w1502 ), .B(
        \SUBBYTES[9].a/w1503 ), .Z(n16336) );
  XOR \SUBBYTES[9].a/U5288  ( .A(\SUBBYTES[9].a/w1487 ), .B(
        \SUBBYTES[9].a/w1490 ), .Z(n16337) );
  XOR \SUBBYTES[9].a/U5287  ( .A(n16339), .B(n16338), .Z(n17414) );
  XOR \SUBBYTES[9].a/U5286  ( .A(n17190), .B(n16340), .Z(n16338) );
  XOR \SUBBYTES[9].a/U5285  ( .A(n17192), .B(n17191), .Z(n16339) );
  XOR \SUBBYTES[9].a/U5284  ( .A(\SUBBYTES[9].a/w1495 ), .B(
        \SUBBYTES[9].a/w1522 ), .Z(n16340) );
  XOR \SUBBYTES[9].a/U5283  ( .A(n16342), .B(n16341), .Z(n17415) );
  XOR \SUBBYTES[9].a/U5282  ( .A(n17193), .B(n16343), .Z(n16341) );
  XOR \SUBBYTES[9].a/U5281  ( .A(\SUBBYTES[9].a/w1528 ), .B(
        \SUBBYTES[9].a/w1530 ), .Z(n16342) );
  XOR \SUBBYTES[9].a/U5280  ( .A(\SUBBYTES[9].a/w1488 ), .B(
        \SUBBYTES[9].a/w1520 ), .Z(n16343) );
  XOR \SUBBYTES[9].a/U5279  ( .A(\SUBBYTES[9].a/w1320 ), .B(
        \SUBBYTES[9].a/w1321 ), .Z(n17195) );
  XOR \SUBBYTES[9].a/U5278  ( .A(n17195), .B(n16344), .Z(n17194) );
  XOR \SUBBYTES[9].a/U5277  ( .A(\SUBBYTES[9].a/w1313 ), .B(
        \SUBBYTES[9].a/w1330 ), .Z(n16344) );
  XOR \SUBBYTES[9].a/U5276  ( .A(n17194), .B(n16345), .Z(n17416) );
  XOR \SUBBYTES[9].a/U5275  ( .A(\SUBBYTES[9].a/w1312 ), .B(
        \SUBBYTES[9].a/w1327 ), .Z(n16345) );
  XOR \SUBBYTES[9].a/U5274  ( .A(n17195), .B(n16346), .Z(n17418) );
  XOR \SUBBYTES[9].a/U5273  ( .A(\SUBBYTES[9].a/w1327 ), .B(
        \SUBBYTES[9].a/w1328 ), .Z(n16346) );
  XOR \SUBBYTES[9].a/U5272  ( .A(\SUBBYTES[9].a/w1289 ), .B(n16347), .Z(n17197) );
  XOR \SUBBYTES[9].a/U5271  ( .A(\SUBBYTES[9].a/w1280 ), .B(
        \SUBBYTES[9].a/w1281 ), .Z(n16347) );
  XOR \SUBBYTES[9].a/U5270  ( .A(n17197), .B(n16348), .Z(n17417) );
  XOR \SUBBYTES[9].a/U5269  ( .A(\SUBBYTES[9].a/w1291 ), .B(n17418), .Z(n16348) );
  XOR \SUBBYTES[9].a/U5268  ( .A(n16350), .B(n16349), .Z(n17198) );
  XOR \SUBBYTES[9].a/U5267  ( .A(n16352), .B(n16351), .Z(n16349) );
  XOR \SUBBYTES[9].a/U5266  ( .A(\SUBBYTES[9].a/w1327 ), .B(
        \SUBBYTES[9].a/w1328 ), .Z(n16350) );
  XOR \SUBBYTES[9].a/U5265  ( .A(\SUBBYTES[9].a/w1291 ), .B(
        \SUBBYTES[9].a/w1315 ), .Z(n16351) );
  XOR \SUBBYTES[9].a/U5264  ( .A(\SUBBYTES[9].a/w1280 ), .B(
        \SUBBYTES[9].a/w1289 ), .Z(n16352) );
  XOR \SUBBYTES[9].a/U5263  ( .A(\SUBBYTES[9].a/w1312 ), .B(n16353), .Z(n17196) );
  XOR \SUBBYTES[9].a/U5262  ( .A(\SUBBYTES[9].a/w1295 ), .B(
        \SUBBYTES[9].a/w1298 ), .Z(n16353) );
  XOR \SUBBYTES[9].a/U5261  ( .A(n17196), .B(n16354), .Z(n17419) );
  XOR \SUBBYTES[9].a/U5260  ( .A(\SUBBYTES[9].a/w1283 ), .B(n17198), .Z(n16354) );
  XOR \SUBBYTES[9].a/U5259  ( .A(n17194), .B(n16355), .Z(n17420) );
  XOR \SUBBYTES[9].a/U5258  ( .A(\SUBBYTES[9].a/w1315 ), .B(
        \SUBBYTES[9].a/w1328 ), .Z(n16355) );
  XOR \SUBBYTES[9].a/U5257  ( .A(n16357), .B(n16356), .Z(n17421) );
  XOR \SUBBYTES[9].a/U5256  ( .A(n16359), .B(n16358), .Z(n16356) );
  XOR \SUBBYTES[9].a/U5255  ( .A(n16361), .B(n16360), .Z(n16357) );
  XOR \SUBBYTES[9].a/U5254  ( .A(\SUBBYTES[9].a/w1327 ), .B(
        \SUBBYTES[9].a/w1330 ), .Z(n16358) );
  XOR \SUBBYTES[9].a/U5253  ( .A(\SUBBYTES[9].a/w1320 ), .B(
        \SUBBYTES[9].a/w1323 ), .Z(n16359) );
  XOR \SUBBYTES[9].a/U5252  ( .A(\SUBBYTES[9].a/w1295 ), .B(
        \SUBBYTES[9].a/w1296 ), .Z(n16360) );
  XOR \SUBBYTES[9].a/U5251  ( .A(\SUBBYTES[9].a/w1280 ), .B(
        \SUBBYTES[9].a/w1283 ), .Z(n16361) );
  XOR \SUBBYTES[9].a/U5250  ( .A(n16363), .B(n16362), .Z(n17422) );
  XOR \SUBBYTES[9].a/U5249  ( .A(n17195), .B(n16364), .Z(n16362) );
  XOR \SUBBYTES[9].a/U5248  ( .A(n17197), .B(n17196), .Z(n16363) );
  XOR \SUBBYTES[9].a/U5247  ( .A(\SUBBYTES[9].a/w1288 ), .B(
        \SUBBYTES[9].a/w1315 ), .Z(n16364) );
  XOR \SUBBYTES[9].a/U5246  ( .A(n16366), .B(n16365), .Z(n17423) );
  XOR \SUBBYTES[9].a/U5245  ( .A(n17198), .B(n16367), .Z(n16365) );
  XOR \SUBBYTES[9].a/U5244  ( .A(\SUBBYTES[9].a/w1321 ), .B(
        \SUBBYTES[9].a/w1323 ), .Z(n16366) );
  XOR \SUBBYTES[9].a/U5243  ( .A(\SUBBYTES[9].a/w1281 ), .B(
        \SUBBYTES[9].a/w1313 ), .Z(n16367) );
  XOR \SUBBYTES[9].a/U5242  ( .A(\SUBBYTES[9].a/w1113 ), .B(
        \SUBBYTES[9].a/w1114 ), .Z(n17200) );
  XOR \SUBBYTES[9].a/U5241  ( .A(n17200), .B(n16368), .Z(n17199) );
  XOR \SUBBYTES[9].a/U5240  ( .A(\SUBBYTES[9].a/w1106 ), .B(
        \SUBBYTES[9].a/w1123 ), .Z(n16368) );
  XOR \SUBBYTES[9].a/U5239  ( .A(n17199), .B(n16369), .Z(n17424) );
  XOR \SUBBYTES[9].a/U5238  ( .A(\SUBBYTES[9].a/w1105 ), .B(
        \SUBBYTES[9].a/w1120 ), .Z(n16369) );
  XOR \SUBBYTES[9].a/U5237  ( .A(n17200), .B(n16370), .Z(n17426) );
  XOR \SUBBYTES[9].a/U5236  ( .A(\SUBBYTES[9].a/w1120 ), .B(
        \SUBBYTES[9].a/w1121 ), .Z(n16370) );
  XOR \SUBBYTES[9].a/U5235  ( .A(\SUBBYTES[9].a/w1082 ), .B(n16371), .Z(n17202) );
  XOR \SUBBYTES[9].a/U5234  ( .A(\SUBBYTES[9].a/w1073 ), .B(
        \SUBBYTES[9].a/w1074 ), .Z(n16371) );
  XOR \SUBBYTES[9].a/U5233  ( .A(n17202), .B(n16372), .Z(n17425) );
  XOR \SUBBYTES[9].a/U5232  ( .A(\SUBBYTES[9].a/w1084 ), .B(n17426), .Z(n16372) );
  XOR \SUBBYTES[9].a/U5231  ( .A(n16374), .B(n16373), .Z(n17203) );
  XOR \SUBBYTES[9].a/U5230  ( .A(n16376), .B(n16375), .Z(n16373) );
  XOR \SUBBYTES[9].a/U5229  ( .A(\SUBBYTES[9].a/w1120 ), .B(
        \SUBBYTES[9].a/w1121 ), .Z(n16374) );
  XOR \SUBBYTES[9].a/U5228  ( .A(\SUBBYTES[9].a/w1084 ), .B(
        \SUBBYTES[9].a/w1108 ), .Z(n16375) );
  XOR \SUBBYTES[9].a/U5227  ( .A(\SUBBYTES[9].a/w1073 ), .B(
        \SUBBYTES[9].a/w1082 ), .Z(n16376) );
  XOR \SUBBYTES[9].a/U5226  ( .A(\SUBBYTES[9].a/w1105 ), .B(n16377), .Z(n17201) );
  XOR \SUBBYTES[9].a/U5225  ( .A(\SUBBYTES[9].a/w1088 ), .B(
        \SUBBYTES[9].a/w1091 ), .Z(n16377) );
  XOR \SUBBYTES[9].a/U5224  ( .A(n17201), .B(n16378), .Z(n17427) );
  XOR \SUBBYTES[9].a/U5223  ( .A(\SUBBYTES[9].a/w1076 ), .B(n17203), .Z(n16378) );
  XOR \SUBBYTES[9].a/U5222  ( .A(n17199), .B(n16379), .Z(n17428) );
  XOR \SUBBYTES[9].a/U5221  ( .A(\SUBBYTES[9].a/w1108 ), .B(
        \SUBBYTES[9].a/w1121 ), .Z(n16379) );
  XOR \SUBBYTES[9].a/U5220  ( .A(n16381), .B(n16380), .Z(n17429) );
  XOR \SUBBYTES[9].a/U5219  ( .A(n16383), .B(n16382), .Z(n16380) );
  XOR \SUBBYTES[9].a/U5218  ( .A(n16385), .B(n16384), .Z(n16381) );
  XOR \SUBBYTES[9].a/U5217  ( .A(\SUBBYTES[9].a/w1120 ), .B(
        \SUBBYTES[9].a/w1123 ), .Z(n16382) );
  XOR \SUBBYTES[9].a/U5216  ( .A(\SUBBYTES[9].a/w1113 ), .B(
        \SUBBYTES[9].a/w1116 ), .Z(n16383) );
  XOR \SUBBYTES[9].a/U5215  ( .A(\SUBBYTES[9].a/w1088 ), .B(
        \SUBBYTES[9].a/w1089 ), .Z(n16384) );
  XOR \SUBBYTES[9].a/U5214  ( .A(\SUBBYTES[9].a/w1073 ), .B(
        \SUBBYTES[9].a/w1076 ), .Z(n16385) );
  XOR \SUBBYTES[9].a/U5213  ( .A(n16387), .B(n16386), .Z(n17430) );
  XOR \SUBBYTES[9].a/U5212  ( .A(n17200), .B(n16388), .Z(n16386) );
  XOR \SUBBYTES[9].a/U5211  ( .A(n17202), .B(n17201), .Z(n16387) );
  XOR \SUBBYTES[9].a/U5210  ( .A(\SUBBYTES[9].a/w1081 ), .B(
        \SUBBYTES[9].a/w1108 ), .Z(n16388) );
  XOR \SUBBYTES[9].a/U5209  ( .A(n16390), .B(n16389), .Z(n17431) );
  XOR \SUBBYTES[9].a/U5208  ( .A(n17203), .B(n16391), .Z(n16389) );
  XOR \SUBBYTES[9].a/U5207  ( .A(\SUBBYTES[9].a/w1114 ), .B(
        \SUBBYTES[9].a/w1116 ), .Z(n16390) );
  XOR \SUBBYTES[9].a/U5206  ( .A(\SUBBYTES[9].a/w1074 ), .B(
        \SUBBYTES[9].a/w1106 ), .Z(n16391) );
  XOR \SUBBYTES[9].a/U5205  ( .A(\SUBBYTES[9].a/w906 ), .B(
        \SUBBYTES[9].a/w907 ), .Z(n17205) );
  XOR \SUBBYTES[9].a/U5204  ( .A(n17205), .B(n16392), .Z(n17204) );
  XOR \SUBBYTES[9].a/U5203  ( .A(\SUBBYTES[9].a/w899 ), .B(
        \SUBBYTES[9].a/w916 ), .Z(n16392) );
  XOR \SUBBYTES[9].a/U5202  ( .A(n17204), .B(n16393), .Z(n17432) );
  XOR \SUBBYTES[9].a/U5201  ( .A(\SUBBYTES[9].a/w898 ), .B(
        \SUBBYTES[9].a/w913 ), .Z(n16393) );
  XOR \SUBBYTES[9].a/U5200  ( .A(n17205), .B(n16394), .Z(n17434) );
  XOR \SUBBYTES[9].a/U5199  ( .A(\SUBBYTES[9].a/w913 ), .B(
        \SUBBYTES[9].a/w914 ), .Z(n16394) );
  XOR \SUBBYTES[9].a/U5198  ( .A(\SUBBYTES[9].a/w875 ), .B(n16395), .Z(n17207)
         );
  XOR \SUBBYTES[9].a/U5197  ( .A(\SUBBYTES[9].a/w866 ), .B(
        \SUBBYTES[9].a/w867 ), .Z(n16395) );
  XOR \SUBBYTES[9].a/U5196  ( .A(n17207), .B(n16396), .Z(n17433) );
  XOR \SUBBYTES[9].a/U5195  ( .A(\SUBBYTES[9].a/w877 ), .B(n17434), .Z(n16396)
         );
  XOR \SUBBYTES[9].a/U5194  ( .A(n16398), .B(n16397), .Z(n17208) );
  XOR \SUBBYTES[9].a/U5193  ( .A(n16400), .B(n16399), .Z(n16397) );
  XOR \SUBBYTES[9].a/U5192  ( .A(\SUBBYTES[9].a/w913 ), .B(
        \SUBBYTES[9].a/w914 ), .Z(n16398) );
  XOR \SUBBYTES[9].a/U5191  ( .A(\SUBBYTES[9].a/w877 ), .B(
        \SUBBYTES[9].a/w901 ), .Z(n16399) );
  XOR \SUBBYTES[9].a/U5190  ( .A(\SUBBYTES[9].a/w866 ), .B(
        \SUBBYTES[9].a/w875 ), .Z(n16400) );
  XOR \SUBBYTES[9].a/U5189  ( .A(\SUBBYTES[9].a/w898 ), .B(n16401), .Z(n17206)
         );
  XOR \SUBBYTES[9].a/U5188  ( .A(\SUBBYTES[9].a/w881 ), .B(
        \SUBBYTES[9].a/w884 ), .Z(n16401) );
  XOR \SUBBYTES[9].a/U5187  ( .A(n17206), .B(n16402), .Z(n17435) );
  XOR \SUBBYTES[9].a/U5186  ( .A(\SUBBYTES[9].a/w869 ), .B(n17208), .Z(n16402)
         );
  XOR \SUBBYTES[9].a/U5185  ( .A(n17204), .B(n16403), .Z(n17436) );
  XOR \SUBBYTES[9].a/U5184  ( .A(\SUBBYTES[9].a/w901 ), .B(
        \SUBBYTES[9].a/w914 ), .Z(n16403) );
  XOR \SUBBYTES[9].a/U5183  ( .A(n16405), .B(n16404), .Z(n17437) );
  XOR \SUBBYTES[9].a/U5182  ( .A(n16407), .B(n16406), .Z(n16404) );
  XOR \SUBBYTES[9].a/U5181  ( .A(n16409), .B(n16408), .Z(n16405) );
  XOR \SUBBYTES[9].a/U5180  ( .A(\SUBBYTES[9].a/w913 ), .B(
        \SUBBYTES[9].a/w916 ), .Z(n16406) );
  XOR \SUBBYTES[9].a/U5179  ( .A(\SUBBYTES[9].a/w906 ), .B(
        \SUBBYTES[9].a/w909 ), .Z(n16407) );
  XOR \SUBBYTES[9].a/U5178  ( .A(\SUBBYTES[9].a/w881 ), .B(
        \SUBBYTES[9].a/w882 ), .Z(n16408) );
  XOR \SUBBYTES[9].a/U5177  ( .A(\SUBBYTES[9].a/w866 ), .B(
        \SUBBYTES[9].a/w869 ), .Z(n16409) );
  XOR \SUBBYTES[9].a/U5176  ( .A(n16411), .B(n16410), .Z(n17438) );
  XOR \SUBBYTES[9].a/U5175  ( .A(n17205), .B(n16412), .Z(n16410) );
  XOR \SUBBYTES[9].a/U5174  ( .A(n17207), .B(n17206), .Z(n16411) );
  XOR \SUBBYTES[9].a/U5173  ( .A(\SUBBYTES[9].a/w874 ), .B(
        \SUBBYTES[9].a/w901 ), .Z(n16412) );
  XOR \SUBBYTES[9].a/U5172  ( .A(n16414), .B(n16413), .Z(n17439) );
  XOR \SUBBYTES[9].a/U5171  ( .A(n17208), .B(n16415), .Z(n16413) );
  XOR \SUBBYTES[9].a/U5170  ( .A(\SUBBYTES[9].a/w907 ), .B(
        \SUBBYTES[9].a/w909 ), .Z(n16414) );
  XOR \SUBBYTES[9].a/U5169  ( .A(\SUBBYTES[9].a/w867 ), .B(
        \SUBBYTES[9].a/w899 ), .Z(n16415) );
  XOR \SUBBYTES[9].a/U5168  ( .A(\SUBBYTES[9].a/w699 ), .B(
        \SUBBYTES[9].a/w700 ), .Z(n17210) );
  XOR \SUBBYTES[9].a/U5167  ( .A(n17210), .B(n16416), .Z(n17209) );
  XOR \SUBBYTES[9].a/U5166  ( .A(\SUBBYTES[9].a/w692 ), .B(
        \SUBBYTES[9].a/w709 ), .Z(n16416) );
  XOR \SUBBYTES[9].a/U5165  ( .A(n17209), .B(n16417), .Z(n17440) );
  XOR \SUBBYTES[9].a/U5164  ( .A(\SUBBYTES[9].a/w691 ), .B(
        \SUBBYTES[9].a/w706 ), .Z(n16417) );
  XOR \SUBBYTES[9].a/U5163  ( .A(n17210), .B(n16418), .Z(n17442) );
  XOR \SUBBYTES[9].a/U5162  ( .A(\SUBBYTES[9].a/w706 ), .B(
        \SUBBYTES[9].a/w707 ), .Z(n16418) );
  XOR \SUBBYTES[9].a/U5161  ( .A(\SUBBYTES[9].a/w668 ), .B(n16419), .Z(n17212)
         );
  XOR \SUBBYTES[9].a/U5160  ( .A(\SUBBYTES[9].a/w659 ), .B(
        \SUBBYTES[9].a/w660 ), .Z(n16419) );
  XOR \SUBBYTES[9].a/U5159  ( .A(n17212), .B(n16420), .Z(n17441) );
  XOR \SUBBYTES[9].a/U5158  ( .A(\SUBBYTES[9].a/w670 ), .B(n17442), .Z(n16420)
         );
  XOR \SUBBYTES[9].a/U5157  ( .A(n16422), .B(n16421), .Z(n17213) );
  XOR \SUBBYTES[9].a/U5156  ( .A(n16424), .B(n16423), .Z(n16421) );
  XOR \SUBBYTES[9].a/U5155  ( .A(\SUBBYTES[9].a/w706 ), .B(
        \SUBBYTES[9].a/w707 ), .Z(n16422) );
  XOR \SUBBYTES[9].a/U5154  ( .A(\SUBBYTES[9].a/w670 ), .B(
        \SUBBYTES[9].a/w694 ), .Z(n16423) );
  XOR \SUBBYTES[9].a/U5153  ( .A(\SUBBYTES[9].a/w659 ), .B(
        \SUBBYTES[9].a/w668 ), .Z(n16424) );
  XOR \SUBBYTES[9].a/U5152  ( .A(\SUBBYTES[9].a/w691 ), .B(n16425), .Z(n17211)
         );
  XOR \SUBBYTES[9].a/U5151  ( .A(\SUBBYTES[9].a/w674 ), .B(
        \SUBBYTES[9].a/w677 ), .Z(n16425) );
  XOR \SUBBYTES[9].a/U5150  ( .A(n17211), .B(n16426), .Z(n17443) );
  XOR \SUBBYTES[9].a/U5149  ( .A(\SUBBYTES[9].a/w662 ), .B(n17213), .Z(n16426)
         );
  XOR \SUBBYTES[9].a/U5148  ( .A(n17209), .B(n16427), .Z(n17444) );
  XOR \SUBBYTES[9].a/U5147  ( .A(\SUBBYTES[9].a/w694 ), .B(
        \SUBBYTES[9].a/w707 ), .Z(n16427) );
  XOR \SUBBYTES[9].a/U5146  ( .A(n16429), .B(n16428), .Z(n17445) );
  XOR \SUBBYTES[9].a/U5145  ( .A(n16431), .B(n16430), .Z(n16428) );
  XOR \SUBBYTES[9].a/U5144  ( .A(n16433), .B(n16432), .Z(n16429) );
  XOR \SUBBYTES[9].a/U5143  ( .A(\SUBBYTES[9].a/w706 ), .B(
        \SUBBYTES[9].a/w709 ), .Z(n16430) );
  XOR \SUBBYTES[9].a/U5142  ( .A(\SUBBYTES[9].a/w699 ), .B(
        \SUBBYTES[9].a/w702 ), .Z(n16431) );
  XOR \SUBBYTES[9].a/U5141  ( .A(\SUBBYTES[9].a/w674 ), .B(
        \SUBBYTES[9].a/w675 ), .Z(n16432) );
  XOR \SUBBYTES[9].a/U5140  ( .A(\SUBBYTES[9].a/w659 ), .B(
        \SUBBYTES[9].a/w662 ), .Z(n16433) );
  XOR \SUBBYTES[9].a/U5139  ( .A(n16435), .B(n16434), .Z(n17446) );
  XOR \SUBBYTES[9].a/U5138  ( .A(n17210), .B(n16436), .Z(n16434) );
  XOR \SUBBYTES[9].a/U5137  ( .A(n17212), .B(n17211), .Z(n16435) );
  XOR \SUBBYTES[9].a/U5136  ( .A(\SUBBYTES[9].a/w667 ), .B(
        \SUBBYTES[9].a/w694 ), .Z(n16436) );
  XOR \SUBBYTES[9].a/U5135  ( .A(n16438), .B(n16437), .Z(n17447) );
  XOR \SUBBYTES[9].a/U5134  ( .A(n17213), .B(n16439), .Z(n16437) );
  XOR \SUBBYTES[9].a/U5133  ( .A(\SUBBYTES[9].a/w700 ), .B(
        \SUBBYTES[9].a/w702 ), .Z(n16438) );
  XOR \SUBBYTES[9].a/U5132  ( .A(\SUBBYTES[9].a/w660 ), .B(
        \SUBBYTES[9].a/w692 ), .Z(n16439) );
  XOR \SUBBYTES[9].a/U5131  ( .A(\SUBBYTES[9].a/w492 ), .B(
        \SUBBYTES[9].a/w493 ), .Z(n17215) );
  XOR \SUBBYTES[9].a/U5130  ( .A(n17215), .B(n16440), .Z(n17214) );
  XOR \SUBBYTES[9].a/U5129  ( .A(\SUBBYTES[9].a/w485 ), .B(
        \SUBBYTES[9].a/w502 ), .Z(n16440) );
  XOR \SUBBYTES[9].a/U5128  ( .A(n17214), .B(n16441), .Z(n17448) );
  XOR \SUBBYTES[9].a/U5127  ( .A(\SUBBYTES[9].a/w484 ), .B(
        \SUBBYTES[9].a/w499 ), .Z(n16441) );
  XOR \SUBBYTES[9].a/U5126  ( .A(n17215), .B(n16442), .Z(n17450) );
  XOR \SUBBYTES[9].a/U5125  ( .A(\SUBBYTES[9].a/w499 ), .B(
        \SUBBYTES[9].a/w500 ), .Z(n16442) );
  XOR \SUBBYTES[9].a/U5124  ( .A(\SUBBYTES[9].a/w461 ), .B(n16443), .Z(n17217)
         );
  XOR \SUBBYTES[9].a/U5123  ( .A(\SUBBYTES[9].a/w452 ), .B(
        \SUBBYTES[9].a/w453 ), .Z(n16443) );
  XOR \SUBBYTES[9].a/U5122  ( .A(n17217), .B(n16444), .Z(n17449) );
  XOR \SUBBYTES[9].a/U5121  ( .A(\SUBBYTES[9].a/w463 ), .B(n17450), .Z(n16444)
         );
  XOR \SUBBYTES[9].a/U5120  ( .A(n16446), .B(n16445), .Z(n17218) );
  XOR \SUBBYTES[9].a/U5119  ( .A(n16448), .B(n16447), .Z(n16445) );
  XOR \SUBBYTES[9].a/U5118  ( .A(\SUBBYTES[9].a/w499 ), .B(
        \SUBBYTES[9].a/w500 ), .Z(n16446) );
  XOR \SUBBYTES[9].a/U5117  ( .A(\SUBBYTES[9].a/w463 ), .B(
        \SUBBYTES[9].a/w487 ), .Z(n16447) );
  XOR \SUBBYTES[9].a/U5116  ( .A(\SUBBYTES[9].a/w452 ), .B(
        \SUBBYTES[9].a/w461 ), .Z(n16448) );
  XOR \SUBBYTES[9].a/U5115  ( .A(\SUBBYTES[9].a/w484 ), .B(n16449), .Z(n17216)
         );
  XOR \SUBBYTES[9].a/U5114  ( .A(\SUBBYTES[9].a/w467 ), .B(
        \SUBBYTES[9].a/w470 ), .Z(n16449) );
  XOR \SUBBYTES[9].a/U5113  ( .A(n17216), .B(n16450), .Z(n17451) );
  XOR \SUBBYTES[9].a/U5112  ( .A(\SUBBYTES[9].a/w455 ), .B(n17218), .Z(n16450)
         );
  XOR \SUBBYTES[9].a/U5111  ( .A(n17214), .B(n16451), .Z(n17452) );
  XOR \SUBBYTES[9].a/U5110  ( .A(\SUBBYTES[9].a/w487 ), .B(
        \SUBBYTES[9].a/w500 ), .Z(n16451) );
  XOR \SUBBYTES[9].a/U5109  ( .A(n16453), .B(n16452), .Z(n17453) );
  XOR \SUBBYTES[9].a/U5108  ( .A(n16455), .B(n16454), .Z(n16452) );
  XOR \SUBBYTES[9].a/U5107  ( .A(n16457), .B(n16456), .Z(n16453) );
  XOR \SUBBYTES[9].a/U5106  ( .A(\SUBBYTES[9].a/w499 ), .B(
        \SUBBYTES[9].a/w502 ), .Z(n16454) );
  XOR \SUBBYTES[9].a/U5105  ( .A(\SUBBYTES[9].a/w492 ), .B(
        \SUBBYTES[9].a/w495 ), .Z(n16455) );
  XOR \SUBBYTES[9].a/U5104  ( .A(\SUBBYTES[9].a/w467 ), .B(
        \SUBBYTES[9].a/w468 ), .Z(n16456) );
  XOR \SUBBYTES[9].a/U5103  ( .A(\SUBBYTES[9].a/w452 ), .B(
        \SUBBYTES[9].a/w455 ), .Z(n16457) );
  XOR \SUBBYTES[9].a/U5102  ( .A(n16459), .B(n16458), .Z(n17454) );
  XOR \SUBBYTES[9].a/U5101  ( .A(n17215), .B(n16460), .Z(n16458) );
  XOR \SUBBYTES[9].a/U5100  ( .A(n17217), .B(n17216), .Z(n16459) );
  XOR \SUBBYTES[9].a/U5099  ( .A(\SUBBYTES[9].a/w460 ), .B(
        \SUBBYTES[9].a/w487 ), .Z(n16460) );
  XOR \SUBBYTES[9].a/U5098  ( .A(n16462), .B(n16461), .Z(n17455) );
  XOR \SUBBYTES[9].a/U5097  ( .A(n17218), .B(n16463), .Z(n16461) );
  XOR \SUBBYTES[9].a/U5096  ( .A(\SUBBYTES[9].a/w493 ), .B(
        \SUBBYTES[9].a/w495 ), .Z(n16462) );
  XOR \SUBBYTES[9].a/U5095  ( .A(\SUBBYTES[9].a/w453 ), .B(
        \SUBBYTES[9].a/w485 ), .Z(n16463) );
  XOR \SUBBYTES[9].a/U5094  ( .A(\SUBBYTES[9].a/w285 ), .B(
        \SUBBYTES[9].a/w286 ), .Z(n17220) );
  XOR \SUBBYTES[9].a/U5093  ( .A(n17220), .B(n16464), .Z(n17219) );
  XOR \SUBBYTES[9].a/U5092  ( .A(\SUBBYTES[9].a/w278 ), .B(
        \SUBBYTES[9].a/w295 ), .Z(n16464) );
  XOR \SUBBYTES[9].a/U5091  ( .A(n17219), .B(n16465), .Z(n17456) );
  XOR \SUBBYTES[9].a/U5090  ( .A(\SUBBYTES[9].a/w277 ), .B(
        \SUBBYTES[9].a/w292 ), .Z(n16465) );
  XOR \SUBBYTES[9].a/U5089  ( .A(n17220), .B(n16466), .Z(n17458) );
  XOR \SUBBYTES[9].a/U5088  ( .A(\SUBBYTES[9].a/w292 ), .B(
        \SUBBYTES[9].a/w293 ), .Z(n16466) );
  XOR \SUBBYTES[9].a/U5087  ( .A(\SUBBYTES[9].a/w254 ), .B(n16467), .Z(n17222)
         );
  XOR \SUBBYTES[9].a/U5086  ( .A(\SUBBYTES[9].a/w245 ), .B(
        \SUBBYTES[9].a/w246 ), .Z(n16467) );
  XOR \SUBBYTES[9].a/U5085  ( .A(n17222), .B(n16468), .Z(n17457) );
  XOR \SUBBYTES[9].a/U5084  ( .A(\SUBBYTES[9].a/w256 ), .B(n17458), .Z(n16468)
         );
  XOR \SUBBYTES[9].a/U5083  ( .A(n16470), .B(n16469), .Z(n17223) );
  XOR \SUBBYTES[9].a/U5082  ( .A(n16472), .B(n16471), .Z(n16469) );
  XOR \SUBBYTES[9].a/U5081  ( .A(\SUBBYTES[9].a/w292 ), .B(
        \SUBBYTES[9].a/w293 ), .Z(n16470) );
  XOR \SUBBYTES[9].a/U5080  ( .A(\SUBBYTES[9].a/w256 ), .B(
        \SUBBYTES[9].a/w280 ), .Z(n16471) );
  XOR \SUBBYTES[9].a/U5079  ( .A(\SUBBYTES[9].a/w245 ), .B(
        \SUBBYTES[9].a/w254 ), .Z(n16472) );
  XOR \SUBBYTES[9].a/U5078  ( .A(\SUBBYTES[9].a/w277 ), .B(n16473), .Z(n17221)
         );
  XOR \SUBBYTES[9].a/U5077  ( .A(\SUBBYTES[9].a/w260 ), .B(
        \SUBBYTES[9].a/w263 ), .Z(n16473) );
  XOR \SUBBYTES[9].a/U5076  ( .A(n17221), .B(n16474), .Z(n17459) );
  XOR \SUBBYTES[9].a/U5075  ( .A(\SUBBYTES[9].a/w248 ), .B(n17223), .Z(n16474)
         );
  XOR \SUBBYTES[9].a/U5074  ( .A(n17219), .B(n16475), .Z(n17460) );
  XOR \SUBBYTES[9].a/U5073  ( .A(\SUBBYTES[9].a/w280 ), .B(
        \SUBBYTES[9].a/w293 ), .Z(n16475) );
  XOR \SUBBYTES[9].a/U5072  ( .A(n16477), .B(n16476), .Z(n17461) );
  XOR \SUBBYTES[9].a/U5071  ( .A(n16479), .B(n16478), .Z(n16476) );
  XOR \SUBBYTES[9].a/U5070  ( .A(n16481), .B(n16480), .Z(n16477) );
  XOR \SUBBYTES[9].a/U5069  ( .A(\SUBBYTES[9].a/w292 ), .B(
        \SUBBYTES[9].a/w295 ), .Z(n16478) );
  XOR \SUBBYTES[9].a/U5068  ( .A(\SUBBYTES[9].a/w285 ), .B(
        \SUBBYTES[9].a/w288 ), .Z(n16479) );
  XOR \SUBBYTES[9].a/U5067  ( .A(\SUBBYTES[9].a/w260 ), .B(
        \SUBBYTES[9].a/w261 ), .Z(n16480) );
  XOR \SUBBYTES[9].a/U5066  ( .A(\SUBBYTES[9].a/w245 ), .B(
        \SUBBYTES[9].a/w248 ), .Z(n16481) );
  XOR \SUBBYTES[9].a/U5065  ( .A(n16483), .B(n16482), .Z(n17462) );
  XOR \SUBBYTES[9].a/U5064  ( .A(n17220), .B(n16484), .Z(n16482) );
  XOR \SUBBYTES[9].a/U5063  ( .A(n17222), .B(n17221), .Z(n16483) );
  XOR \SUBBYTES[9].a/U5062  ( .A(\SUBBYTES[9].a/w253 ), .B(
        \SUBBYTES[9].a/w280 ), .Z(n16484) );
  XOR \SUBBYTES[9].a/U5061  ( .A(n16486), .B(n16485), .Z(n17463) );
  XOR \SUBBYTES[9].a/U5060  ( .A(n17223), .B(n16487), .Z(n16485) );
  XOR \SUBBYTES[9].a/U5059  ( .A(\SUBBYTES[9].a/w286 ), .B(
        \SUBBYTES[9].a/w288 ), .Z(n16486) );
  XOR \SUBBYTES[9].a/U5058  ( .A(\SUBBYTES[9].a/w246 ), .B(
        \SUBBYTES[9].a/w278 ), .Z(n16487) );
  XOR \SUBBYTES[9].a/U5057  ( .A(\w1[9][1] ), .B(n16488), .Z(n17224) );
  XOR \SUBBYTES[9].a/U5056  ( .A(\w1[9][3] ), .B(\w1[9][2] ), .Z(n16488) );
  XOR \SUBBYTES[9].a/U5055  ( .A(\w1[9][6] ), .B(n17224), .Z(
        \SUBBYTES[9].a/w3378 ) );
  XOR \SUBBYTES[9].a/U5054  ( .A(\w1[9][0] ), .B(\SUBBYTES[9].a/w3378 ), .Z(
        \SUBBYTES[9].a/w3265 ) );
  XOR \SUBBYTES[9].a/U5053  ( .A(\w1[9][0] ), .B(n16489), .Z(
        \SUBBYTES[9].a/w3266 ) );
  XOR \SUBBYTES[9].a/U5052  ( .A(\w1[9][6] ), .B(\w1[9][5] ), .Z(n16489) );
  XOR \SUBBYTES[9].a/U5051  ( .A(\w1[9][5] ), .B(n17224), .Z(
        \SUBBYTES[9].a/w3396 ) );
  XOR \SUBBYTES[9].a/U5050  ( .A(n16491), .B(n16490), .Z(\SUBBYTES[9].a/w3389 ) );
  XOR \SUBBYTES[9].a/U5049  ( .A(\w1[9][3] ), .B(\w1[9][1] ), .Z(n16490) );
  XOR \SUBBYTES[9].a/U5048  ( .A(\w1[9][7] ), .B(\w1[9][4] ), .Z(n16491) );
  XOR \SUBBYTES[9].a/U5047  ( .A(\w1[9][0] ), .B(\SUBBYTES[9].a/w3389 ), .Z(
        \SUBBYTES[9].a/w3268 ) );
  XOR \SUBBYTES[9].a/U5046  ( .A(n16493), .B(n16492), .Z(\SUBBYTES[9].a/w3376 ) );
  XOR \SUBBYTES[9].a/U5045  ( .A(\SUBBYTES[9].a/w3337 ), .B(n1100), .Z(n16492)
         );
  XOR \SUBBYTES[9].a/U5044  ( .A(\SUBBYTES[9].a/w3330 ), .B(
        \SUBBYTES[9].a/w3333 ), .Z(n16493) );
  XOR \SUBBYTES[9].a/U5043  ( .A(n16495), .B(n16494), .Z(\SUBBYTES[9].a/w3377 ) );
  XOR \SUBBYTES[9].a/U5042  ( .A(\SUBBYTES[9].a/w3337 ), .B(n16103), .Z(n16494) );
  XOR \SUBBYTES[9].a/U5041  ( .A(\SUBBYTES[9].a/w3330 ), .B(n16102), .Z(n16495) );
  XOR \SUBBYTES[9].a/U5040  ( .A(\SUBBYTES[9].a/w3389 ), .B(n16496), .Z(
        \SUBBYTES[9].a/w3379 ) );
  XOR \SUBBYTES[9].a/U5039  ( .A(\w1[9][6] ), .B(\w1[9][5] ), .Z(n16496) );
  XOR \SUBBYTES[9].a/U5038  ( .A(n16498), .B(n16497), .Z(\SUBBYTES[9].a/w3380 ) );
  XOR \SUBBYTES[9].a/U5037  ( .A(n16103), .B(n1100), .Z(n16497) );
  XOR \SUBBYTES[9].a/U5036  ( .A(n16102), .B(\SUBBYTES[9].a/w3333 ), .Z(n16498) );
  XOR \SUBBYTES[9].a/U5035  ( .A(\w1[9][7] ), .B(\w1[9][2] ), .Z(n17230) );
  XOR \SUBBYTES[9].a/U5034  ( .A(n17230), .B(n16499), .Z(\SUBBYTES[9].a/w3381 ) );
  XOR \SUBBYTES[9].a/U5033  ( .A(\w1[9][5] ), .B(\w1[9][4] ), .Z(n16499) );
  XOR \SUBBYTES[9].a/U5032  ( .A(\w1[9][7] ), .B(\SUBBYTES[9].a/w3266 ), .Z(
        \SUBBYTES[9].a/w3269 ) );
  XOR \SUBBYTES[9].a/U5031  ( .A(\w1[9][1] ), .B(\SUBBYTES[9].a/w3266 ), .Z(
        \SUBBYTES[9].a/w3270 ) );
  XOR \SUBBYTES[9].a/U5030  ( .A(\w1[9][4] ), .B(\SUBBYTES[9].a/w3266 ), .Z(
        \SUBBYTES[9].a/w3271 ) );
  XOR \SUBBYTES[9].a/U5029  ( .A(\SUBBYTES[9].a/w3270 ), .B(n17230), .Z(
        \SUBBYTES[9].a/w3272 ) );
  XOR \SUBBYTES[9].a/U5028  ( .A(n17230), .B(n16500), .Z(\SUBBYTES[9].a/w3357 ) );
  XOR \SUBBYTES[9].a/U5027  ( .A(\w1[9][4] ), .B(\w1[9][1] ), .Z(n16500) );
  XOR \SUBBYTES[9].a/U5026  ( .A(n16502), .B(n16501), .Z(n17227) );
  XOR \SUBBYTES[9].a/U5025  ( .A(\w1[9][4] ), .B(n16503), .Z(n16501) );
  XOR \SUBBYTES[9].a/U5024  ( .A(\SUBBYTES[9].a/w3322 ), .B(\w1[9][6] ), .Z(
        n16502) );
  XOR \SUBBYTES[9].a/U5023  ( .A(\SUBBYTES[9].a/w3296 ), .B(
        \SUBBYTES[9].a/w3303 ), .Z(n16503) );
  XOR \SUBBYTES[9].a/U5022  ( .A(n16505), .B(n16504), .Z(n17225) );
  XOR \SUBBYTES[9].a/U5021  ( .A(\w1[9][1] ), .B(n16506), .Z(n16504) );
  XOR \SUBBYTES[9].a/U5020  ( .A(\SUBBYTES[9].a/w3321 ), .B(\w1[9][5] ), .Z(
        n16505) );
  XOR \SUBBYTES[9].a/U5019  ( .A(\SUBBYTES[9].a/w3297 ), .B(
        \SUBBYTES[9].a/w3304 ), .Z(n16506) );
  XOR \SUBBYTES[9].a/U5018  ( .A(n17227), .B(n17225), .Z(\SUBBYTES[9].a/w3327 ) );
  XOR \SUBBYTES[9].a/U5017  ( .A(\w1[9][5] ), .B(n16507), .Z(n17228) );
  XOR \SUBBYTES[9].a/U5016  ( .A(\SUBBYTES[9].a/w3289 ), .B(
        \SUBBYTES[9].a/w3299 ), .Z(n16507) );
  XOR \SUBBYTES[9].a/U5015  ( .A(n16509), .B(n16508), .Z(\SUBBYTES[9].a/w3314 ) );
  XOR \SUBBYTES[9].a/U5014  ( .A(n17228), .B(n16510), .Z(n16508) );
  XOR \SUBBYTES[9].a/U5013  ( .A(\w1[9][4] ), .B(\SUBBYTES[9].a/w3378 ), .Z(
        n16509) );
  XOR \SUBBYTES[9].a/U5012  ( .A(\SUBBYTES[9].a/w3291 ), .B(
        \SUBBYTES[9].a/w3296 ), .Z(n16510) );
  XOR \SUBBYTES[9].a/U5011  ( .A(n16512), .B(n16511), .Z(n17226) );
  XOR \SUBBYTES[9].a/U5010  ( .A(\SUBBYTES[9].a/w3324 ), .B(\w1[9][7] ), .Z(
        n16511) );
  XOR \SUBBYTES[9].a/U5009  ( .A(\SUBBYTES[9].a/w3299 ), .B(
        \SUBBYTES[9].a/w3306 ), .Z(n16512) );
  XOR \SUBBYTES[9].a/U5008  ( .A(n17225), .B(n17226), .Z(\SUBBYTES[9].a/w3326 ) );
  XOR \SUBBYTES[9].a/U5007  ( .A(\w1[9][3] ), .B(n16513), .Z(n17229) );
  XOR \SUBBYTES[9].a/U5006  ( .A(\SUBBYTES[9].a/w3288 ), .B(
        \SUBBYTES[9].a/w3291 ), .Z(n16513) );
  XOR \SUBBYTES[9].a/U5005  ( .A(n16515), .B(n16514), .Z(\SUBBYTES[9].a/w3315 ) );
  XOR \SUBBYTES[9].a/U5004  ( .A(n17229), .B(n16516), .Z(n16514) );
  XOR \SUBBYTES[9].a/U5003  ( .A(\w1[9][6] ), .B(\SUBBYTES[9].a/w3357 ), .Z(
        n16515) );
  XOR \SUBBYTES[9].a/U5002  ( .A(\SUBBYTES[9].a/w3296 ), .B(
        \SUBBYTES[9].a/w3297 ), .Z(n16516) );
  XOR \SUBBYTES[9].a/U5001  ( .A(n17227), .B(n17226), .Z(\SUBBYTES[9].a/w3335 ) );
  XOR \SUBBYTES[9].a/U5000  ( .A(n16518), .B(n16517), .Z(\SUBBYTES[9].a/w3336 ) );
  XOR \SUBBYTES[9].a/U4999  ( .A(\w1[9][7] ), .B(n17228), .Z(n16517) );
  XOR \SUBBYTES[9].a/U4998  ( .A(\SUBBYTES[9].a/w3288 ), .B(
        \SUBBYTES[9].a/w3297 ), .Z(n16518) );
  XOR \SUBBYTES[9].a/U4997  ( .A(n16520), .B(n16519), .Z(\SUBBYTES[9].a/w3312 ) );
  XOR \SUBBYTES[9].a/U4996  ( .A(n16522), .B(n16521), .Z(n16519) );
  XOR \SUBBYTES[9].a/U4995  ( .A(\w1[9][7] ), .B(\SUBBYTES[9].a/w3396 ), .Z(
        n16520) );
  XOR \SUBBYTES[9].a/U4994  ( .A(\SUBBYTES[9].a/w3303 ), .B(
        \SUBBYTES[9].a/w3306 ), .Z(n16521) );
  XOR \SUBBYTES[9].a/U4993  ( .A(\SUBBYTES[9].a/w3289 ), .B(
        \SUBBYTES[9].a/w3291 ), .Z(n16522) );
  XOR \SUBBYTES[9].a/U4992  ( .A(n16524), .B(n16523), .Z(\SUBBYTES[9].a/w3313 ) );
  XOR \SUBBYTES[9].a/U4991  ( .A(n17229), .B(n16525), .Z(n16523) );
  XOR \SUBBYTES[9].a/U4990  ( .A(\w1[9][5] ), .B(n17230), .Z(n16524) );
  XOR \SUBBYTES[9].a/U4989  ( .A(\SUBBYTES[9].a/w3303 ), .B(
        \SUBBYTES[9].a/w3304 ), .Z(n16525) );
  XOR \SUBBYTES[9].a/U4988  ( .A(n16527), .B(n16526), .Z(\SUBBYTES[9].a/w3329 ) );
  XOR \SUBBYTES[9].a/U4987  ( .A(\w1[9][1] ), .B(n16528), .Z(n16526) );
  XOR \SUBBYTES[9].a/U4986  ( .A(\SUBBYTES[9].a/w3304 ), .B(
        \SUBBYTES[9].a/w3306 ), .Z(n16527) );
  XOR \SUBBYTES[9].a/U4985  ( .A(\SUBBYTES[9].a/w3288 ), .B(
        \SUBBYTES[9].a/w3289 ), .Z(n16528) );
  XOR \SUBBYTES[9].a/U4984  ( .A(\w1[9][9] ), .B(n16529), .Z(n17231) );
  XOR \SUBBYTES[9].a/U4983  ( .A(\w1[9][11] ), .B(\w1[9][10] ), .Z(n16529) );
  XOR \SUBBYTES[9].a/U4982  ( .A(\w1[9][14] ), .B(n17231), .Z(
        \SUBBYTES[9].a/w3171 ) );
  XOR \SUBBYTES[9].a/U4981  ( .A(\w1[9][8] ), .B(\SUBBYTES[9].a/w3171 ), .Z(
        \SUBBYTES[9].a/w3058 ) );
  XOR \SUBBYTES[9].a/U4980  ( .A(\w1[9][8] ), .B(n16530), .Z(
        \SUBBYTES[9].a/w3059 ) );
  XOR \SUBBYTES[9].a/U4979  ( .A(\w1[9][14] ), .B(\w1[9][13] ), .Z(n16530) );
  XOR \SUBBYTES[9].a/U4978  ( .A(\w1[9][13] ), .B(n17231), .Z(
        \SUBBYTES[9].a/w3189 ) );
  XOR \SUBBYTES[9].a/U4977  ( .A(n16532), .B(n16531), .Z(\SUBBYTES[9].a/w3182 ) );
  XOR \SUBBYTES[9].a/U4976  ( .A(\w1[9][11] ), .B(\w1[9][9] ), .Z(n16531) );
  XOR \SUBBYTES[9].a/U4975  ( .A(\w1[9][15] ), .B(\w1[9][12] ), .Z(n16532) );
  XOR \SUBBYTES[9].a/U4974  ( .A(\w1[9][8] ), .B(\SUBBYTES[9].a/w3182 ), .Z(
        \SUBBYTES[9].a/w3061 ) );
  XOR \SUBBYTES[9].a/U4973  ( .A(n16534), .B(n16533), .Z(\SUBBYTES[9].a/w3169 ) );
  XOR \SUBBYTES[9].a/U4972  ( .A(\SUBBYTES[9].a/w3130 ), .B(n1099), .Z(n16533)
         );
  XOR \SUBBYTES[9].a/U4971  ( .A(\SUBBYTES[9].a/w3123 ), .B(
        \SUBBYTES[9].a/w3126 ), .Z(n16534) );
  XOR \SUBBYTES[9].a/U4970  ( .A(n16536), .B(n16535), .Z(\SUBBYTES[9].a/w3170 ) );
  XOR \SUBBYTES[9].a/U4969  ( .A(\SUBBYTES[9].a/w3130 ), .B(n16101), .Z(n16535) );
  XOR \SUBBYTES[9].a/U4968  ( .A(\SUBBYTES[9].a/w3123 ), .B(n16100), .Z(n16536) );
  XOR \SUBBYTES[9].a/U4967  ( .A(\SUBBYTES[9].a/w3182 ), .B(n16537), .Z(
        \SUBBYTES[9].a/w3172 ) );
  XOR \SUBBYTES[9].a/U4966  ( .A(\w1[9][14] ), .B(\w1[9][13] ), .Z(n16537) );
  XOR \SUBBYTES[9].a/U4965  ( .A(n16539), .B(n16538), .Z(\SUBBYTES[9].a/w3173 ) );
  XOR \SUBBYTES[9].a/U4964  ( .A(n16101), .B(n1099), .Z(n16538) );
  XOR \SUBBYTES[9].a/U4963  ( .A(n16100), .B(\SUBBYTES[9].a/w3126 ), .Z(n16539) );
  XOR \SUBBYTES[9].a/U4962  ( .A(\w1[9][15] ), .B(\w1[9][10] ), .Z(n17237) );
  XOR \SUBBYTES[9].a/U4961  ( .A(n17237), .B(n16540), .Z(\SUBBYTES[9].a/w3174 ) );
  XOR \SUBBYTES[9].a/U4960  ( .A(\w1[9][13] ), .B(\w1[9][12] ), .Z(n16540) );
  XOR \SUBBYTES[9].a/U4959  ( .A(\w1[9][15] ), .B(\SUBBYTES[9].a/w3059 ), .Z(
        \SUBBYTES[9].a/w3062 ) );
  XOR \SUBBYTES[9].a/U4958  ( .A(\w1[9][9] ), .B(\SUBBYTES[9].a/w3059 ), .Z(
        \SUBBYTES[9].a/w3063 ) );
  XOR \SUBBYTES[9].a/U4957  ( .A(\w1[9][12] ), .B(\SUBBYTES[9].a/w3059 ), .Z(
        \SUBBYTES[9].a/w3064 ) );
  XOR \SUBBYTES[9].a/U4956  ( .A(\SUBBYTES[9].a/w3063 ), .B(n17237), .Z(
        \SUBBYTES[9].a/w3065 ) );
  XOR \SUBBYTES[9].a/U4955  ( .A(n17237), .B(n16541), .Z(\SUBBYTES[9].a/w3150 ) );
  XOR \SUBBYTES[9].a/U4954  ( .A(\w1[9][12] ), .B(\w1[9][9] ), .Z(n16541) );
  XOR \SUBBYTES[9].a/U4953  ( .A(n16543), .B(n16542), .Z(n17234) );
  XOR \SUBBYTES[9].a/U4952  ( .A(\w1[9][12] ), .B(n16544), .Z(n16542) );
  XOR \SUBBYTES[9].a/U4951  ( .A(\SUBBYTES[9].a/w3115 ), .B(\w1[9][14] ), .Z(
        n16543) );
  XOR \SUBBYTES[9].a/U4950  ( .A(\SUBBYTES[9].a/w3089 ), .B(
        \SUBBYTES[9].a/w3096 ), .Z(n16544) );
  XOR \SUBBYTES[9].a/U4949  ( .A(n16546), .B(n16545), .Z(n17232) );
  XOR \SUBBYTES[9].a/U4948  ( .A(\w1[9][9] ), .B(n16547), .Z(n16545) );
  XOR \SUBBYTES[9].a/U4947  ( .A(\SUBBYTES[9].a/w3114 ), .B(\w1[9][13] ), .Z(
        n16546) );
  XOR \SUBBYTES[9].a/U4946  ( .A(\SUBBYTES[9].a/w3090 ), .B(
        \SUBBYTES[9].a/w3097 ), .Z(n16547) );
  XOR \SUBBYTES[9].a/U4945  ( .A(n17234), .B(n17232), .Z(\SUBBYTES[9].a/w3120 ) );
  XOR \SUBBYTES[9].a/U4944  ( .A(\w1[9][13] ), .B(n16548), .Z(n17235) );
  XOR \SUBBYTES[9].a/U4943  ( .A(\SUBBYTES[9].a/w3082 ), .B(
        \SUBBYTES[9].a/w3092 ), .Z(n16548) );
  XOR \SUBBYTES[9].a/U4942  ( .A(n16550), .B(n16549), .Z(\SUBBYTES[9].a/w3107 ) );
  XOR \SUBBYTES[9].a/U4941  ( .A(n17235), .B(n16551), .Z(n16549) );
  XOR \SUBBYTES[9].a/U4940  ( .A(\w1[9][12] ), .B(\SUBBYTES[9].a/w3171 ), .Z(
        n16550) );
  XOR \SUBBYTES[9].a/U4939  ( .A(\SUBBYTES[9].a/w3084 ), .B(
        \SUBBYTES[9].a/w3089 ), .Z(n16551) );
  XOR \SUBBYTES[9].a/U4938  ( .A(n16553), .B(n16552), .Z(n17233) );
  XOR \SUBBYTES[9].a/U4937  ( .A(\SUBBYTES[9].a/w3117 ), .B(\w1[9][15] ), .Z(
        n16552) );
  XOR \SUBBYTES[9].a/U4936  ( .A(\SUBBYTES[9].a/w3092 ), .B(
        \SUBBYTES[9].a/w3099 ), .Z(n16553) );
  XOR \SUBBYTES[9].a/U4935  ( .A(n17232), .B(n17233), .Z(\SUBBYTES[9].a/w3119 ) );
  XOR \SUBBYTES[9].a/U4934  ( .A(\w1[9][11] ), .B(n16554), .Z(n17236) );
  XOR \SUBBYTES[9].a/U4933  ( .A(\SUBBYTES[9].a/w3081 ), .B(
        \SUBBYTES[9].a/w3084 ), .Z(n16554) );
  XOR \SUBBYTES[9].a/U4932  ( .A(n16556), .B(n16555), .Z(\SUBBYTES[9].a/w3108 ) );
  XOR \SUBBYTES[9].a/U4931  ( .A(n17236), .B(n16557), .Z(n16555) );
  XOR \SUBBYTES[9].a/U4930  ( .A(\w1[9][14] ), .B(\SUBBYTES[9].a/w3150 ), .Z(
        n16556) );
  XOR \SUBBYTES[9].a/U4929  ( .A(\SUBBYTES[9].a/w3089 ), .B(
        \SUBBYTES[9].a/w3090 ), .Z(n16557) );
  XOR \SUBBYTES[9].a/U4928  ( .A(n17234), .B(n17233), .Z(\SUBBYTES[9].a/w3128 ) );
  XOR \SUBBYTES[9].a/U4927  ( .A(n16559), .B(n16558), .Z(\SUBBYTES[9].a/w3129 ) );
  XOR \SUBBYTES[9].a/U4926  ( .A(\w1[9][15] ), .B(n17235), .Z(n16558) );
  XOR \SUBBYTES[9].a/U4925  ( .A(\SUBBYTES[9].a/w3081 ), .B(
        \SUBBYTES[9].a/w3090 ), .Z(n16559) );
  XOR \SUBBYTES[9].a/U4924  ( .A(n16561), .B(n16560), .Z(\SUBBYTES[9].a/w3105 ) );
  XOR \SUBBYTES[9].a/U4923  ( .A(n16563), .B(n16562), .Z(n16560) );
  XOR \SUBBYTES[9].a/U4922  ( .A(\w1[9][15] ), .B(\SUBBYTES[9].a/w3189 ), .Z(
        n16561) );
  XOR \SUBBYTES[9].a/U4921  ( .A(\SUBBYTES[9].a/w3096 ), .B(
        \SUBBYTES[9].a/w3099 ), .Z(n16562) );
  XOR \SUBBYTES[9].a/U4920  ( .A(\SUBBYTES[9].a/w3082 ), .B(
        \SUBBYTES[9].a/w3084 ), .Z(n16563) );
  XOR \SUBBYTES[9].a/U4919  ( .A(n16565), .B(n16564), .Z(\SUBBYTES[9].a/w3106 ) );
  XOR \SUBBYTES[9].a/U4918  ( .A(n17236), .B(n16566), .Z(n16564) );
  XOR \SUBBYTES[9].a/U4917  ( .A(\w1[9][13] ), .B(n17237), .Z(n16565) );
  XOR \SUBBYTES[9].a/U4916  ( .A(\SUBBYTES[9].a/w3096 ), .B(
        \SUBBYTES[9].a/w3097 ), .Z(n16566) );
  XOR \SUBBYTES[9].a/U4915  ( .A(n16568), .B(n16567), .Z(\SUBBYTES[9].a/w3122 ) );
  XOR \SUBBYTES[9].a/U4914  ( .A(\w1[9][9] ), .B(n16569), .Z(n16567) );
  XOR \SUBBYTES[9].a/U4913  ( .A(\SUBBYTES[9].a/w3097 ), .B(
        \SUBBYTES[9].a/w3099 ), .Z(n16568) );
  XOR \SUBBYTES[9].a/U4912  ( .A(\SUBBYTES[9].a/w3081 ), .B(
        \SUBBYTES[9].a/w3082 ), .Z(n16569) );
  XOR \SUBBYTES[9].a/U4911  ( .A(\w1[9][17] ), .B(n16570), .Z(n17238) );
  XOR \SUBBYTES[9].a/U4910  ( .A(\w1[9][19] ), .B(\w1[9][18] ), .Z(n16570) );
  XOR \SUBBYTES[9].a/U4909  ( .A(\w1[9][22] ), .B(n17238), .Z(
        \SUBBYTES[9].a/w2964 ) );
  XOR \SUBBYTES[9].a/U4908  ( .A(\w1[9][16] ), .B(\SUBBYTES[9].a/w2964 ), .Z(
        \SUBBYTES[9].a/w2851 ) );
  XOR \SUBBYTES[9].a/U4907  ( .A(\w1[9][16] ), .B(n16571), .Z(
        \SUBBYTES[9].a/w2852 ) );
  XOR \SUBBYTES[9].a/U4906  ( .A(\w1[9][22] ), .B(\w1[9][21] ), .Z(n16571) );
  XOR \SUBBYTES[9].a/U4905  ( .A(\w1[9][21] ), .B(n17238), .Z(
        \SUBBYTES[9].a/w2982 ) );
  XOR \SUBBYTES[9].a/U4904  ( .A(n16573), .B(n16572), .Z(\SUBBYTES[9].a/w2975 ) );
  XOR \SUBBYTES[9].a/U4903  ( .A(\w1[9][19] ), .B(\w1[9][17] ), .Z(n16572) );
  XOR \SUBBYTES[9].a/U4902  ( .A(\w1[9][23] ), .B(\w1[9][20] ), .Z(n16573) );
  XOR \SUBBYTES[9].a/U4901  ( .A(\w1[9][16] ), .B(\SUBBYTES[9].a/w2975 ), .Z(
        \SUBBYTES[9].a/w2854 ) );
  XOR \SUBBYTES[9].a/U4900  ( .A(n16575), .B(n16574), .Z(\SUBBYTES[9].a/w2962 ) );
  XOR \SUBBYTES[9].a/U4899  ( .A(\SUBBYTES[9].a/w2923 ), .B(n1098), .Z(n16574)
         );
  XOR \SUBBYTES[9].a/U4898  ( .A(\SUBBYTES[9].a/w2916 ), .B(
        \SUBBYTES[9].a/w2919 ), .Z(n16575) );
  XOR \SUBBYTES[9].a/U4897  ( .A(n16577), .B(n16576), .Z(\SUBBYTES[9].a/w2963 ) );
  XOR \SUBBYTES[9].a/U4896  ( .A(\SUBBYTES[9].a/w2923 ), .B(n16099), .Z(n16576) );
  XOR \SUBBYTES[9].a/U4895  ( .A(\SUBBYTES[9].a/w2916 ), .B(n16098), .Z(n16577) );
  XOR \SUBBYTES[9].a/U4894  ( .A(\SUBBYTES[9].a/w2975 ), .B(n16578), .Z(
        \SUBBYTES[9].a/w2965 ) );
  XOR \SUBBYTES[9].a/U4893  ( .A(\w1[9][22] ), .B(\w1[9][21] ), .Z(n16578) );
  XOR \SUBBYTES[9].a/U4892  ( .A(n16580), .B(n16579), .Z(\SUBBYTES[9].a/w2966 ) );
  XOR \SUBBYTES[9].a/U4891  ( .A(n16099), .B(n1098), .Z(n16579) );
  XOR \SUBBYTES[9].a/U4890  ( .A(n16098), .B(\SUBBYTES[9].a/w2919 ), .Z(n16580) );
  XOR \SUBBYTES[9].a/U4889  ( .A(\w1[9][23] ), .B(\w1[9][18] ), .Z(n17244) );
  XOR \SUBBYTES[9].a/U4888  ( .A(n17244), .B(n16581), .Z(\SUBBYTES[9].a/w2967 ) );
  XOR \SUBBYTES[9].a/U4887  ( .A(\w1[9][21] ), .B(\w1[9][20] ), .Z(n16581) );
  XOR \SUBBYTES[9].a/U4886  ( .A(\w1[9][23] ), .B(\SUBBYTES[9].a/w2852 ), .Z(
        \SUBBYTES[9].a/w2855 ) );
  XOR \SUBBYTES[9].a/U4885  ( .A(\w1[9][17] ), .B(\SUBBYTES[9].a/w2852 ), .Z(
        \SUBBYTES[9].a/w2856 ) );
  XOR \SUBBYTES[9].a/U4884  ( .A(\w1[9][20] ), .B(\SUBBYTES[9].a/w2852 ), .Z(
        \SUBBYTES[9].a/w2857 ) );
  XOR \SUBBYTES[9].a/U4883  ( .A(\SUBBYTES[9].a/w2856 ), .B(n17244), .Z(
        \SUBBYTES[9].a/w2858 ) );
  XOR \SUBBYTES[9].a/U4882  ( .A(n17244), .B(n16582), .Z(\SUBBYTES[9].a/w2943 ) );
  XOR \SUBBYTES[9].a/U4881  ( .A(\w1[9][20] ), .B(\w1[9][17] ), .Z(n16582) );
  XOR \SUBBYTES[9].a/U4880  ( .A(n16584), .B(n16583), .Z(n17241) );
  XOR \SUBBYTES[9].a/U4879  ( .A(\w1[9][20] ), .B(n16585), .Z(n16583) );
  XOR \SUBBYTES[9].a/U4878  ( .A(\SUBBYTES[9].a/w2908 ), .B(\w1[9][22] ), .Z(
        n16584) );
  XOR \SUBBYTES[9].a/U4877  ( .A(\SUBBYTES[9].a/w2882 ), .B(
        \SUBBYTES[9].a/w2889 ), .Z(n16585) );
  XOR \SUBBYTES[9].a/U4876  ( .A(n16587), .B(n16586), .Z(n17239) );
  XOR \SUBBYTES[9].a/U4875  ( .A(\w1[9][17] ), .B(n16588), .Z(n16586) );
  XOR \SUBBYTES[9].a/U4874  ( .A(\SUBBYTES[9].a/w2907 ), .B(\w1[9][21] ), .Z(
        n16587) );
  XOR \SUBBYTES[9].a/U4873  ( .A(\SUBBYTES[9].a/w2883 ), .B(
        \SUBBYTES[9].a/w2890 ), .Z(n16588) );
  XOR \SUBBYTES[9].a/U4872  ( .A(n17241), .B(n17239), .Z(\SUBBYTES[9].a/w2913 ) );
  XOR \SUBBYTES[9].a/U4871  ( .A(\w1[9][21] ), .B(n16589), .Z(n17242) );
  XOR \SUBBYTES[9].a/U4870  ( .A(\SUBBYTES[9].a/w2875 ), .B(
        \SUBBYTES[9].a/w2885 ), .Z(n16589) );
  XOR \SUBBYTES[9].a/U4869  ( .A(n16591), .B(n16590), .Z(\SUBBYTES[9].a/w2900 ) );
  XOR \SUBBYTES[9].a/U4868  ( .A(n17242), .B(n16592), .Z(n16590) );
  XOR \SUBBYTES[9].a/U4867  ( .A(\w1[9][20] ), .B(\SUBBYTES[9].a/w2964 ), .Z(
        n16591) );
  XOR \SUBBYTES[9].a/U4866  ( .A(\SUBBYTES[9].a/w2877 ), .B(
        \SUBBYTES[9].a/w2882 ), .Z(n16592) );
  XOR \SUBBYTES[9].a/U4865  ( .A(n16594), .B(n16593), .Z(n17240) );
  XOR \SUBBYTES[9].a/U4864  ( .A(\SUBBYTES[9].a/w2910 ), .B(\w1[9][23] ), .Z(
        n16593) );
  XOR \SUBBYTES[9].a/U4863  ( .A(\SUBBYTES[9].a/w2885 ), .B(
        \SUBBYTES[9].a/w2892 ), .Z(n16594) );
  XOR \SUBBYTES[9].a/U4862  ( .A(n17239), .B(n17240), .Z(\SUBBYTES[9].a/w2912 ) );
  XOR \SUBBYTES[9].a/U4861  ( .A(\w1[9][19] ), .B(n16595), .Z(n17243) );
  XOR \SUBBYTES[9].a/U4860  ( .A(\SUBBYTES[9].a/w2874 ), .B(
        \SUBBYTES[9].a/w2877 ), .Z(n16595) );
  XOR \SUBBYTES[9].a/U4859  ( .A(n16597), .B(n16596), .Z(\SUBBYTES[9].a/w2901 ) );
  XOR \SUBBYTES[9].a/U4858  ( .A(n17243), .B(n16598), .Z(n16596) );
  XOR \SUBBYTES[9].a/U4857  ( .A(\w1[9][22] ), .B(\SUBBYTES[9].a/w2943 ), .Z(
        n16597) );
  XOR \SUBBYTES[9].a/U4856  ( .A(\SUBBYTES[9].a/w2882 ), .B(
        \SUBBYTES[9].a/w2883 ), .Z(n16598) );
  XOR \SUBBYTES[9].a/U4855  ( .A(n17241), .B(n17240), .Z(\SUBBYTES[9].a/w2921 ) );
  XOR \SUBBYTES[9].a/U4854  ( .A(n16600), .B(n16599), .Z(\SUBBYTES[9].a/w2922 ) );
  XOR \SUBBYTES[9].a/U4853  ( .A(\w1[9][23] ), .B(n17242), .Z(n16599) );
  XOR \SUBBYTES[9].a/U4852  ( .A(\SUBBYTES[9].a/w2874 ), .B(
        \SUBBYTES[9].a/w2883 ), .Z(n16600) );
  XOR \SUBBYTES[9].a/U4851  ( .A(n16602), .B(n16601), .Z(\SUBBYTES[9].a/w2898 ) );
  XOR \SUBBYTES[9].a/U4850  ( .A(n16604), .B(n16603), .Z(n16601) );
  XOR \SUBBYTES[9].a/U4849  ( .A(\w1[9][23] ), .B(\SUBBYTES[9].a/w2982 ), .Z(
        n16602) );
  XOR \SUBBYTES[9].a/U4848  ( .A(\SUBBYTES[9].a/w2889 ), .B(
        \SUBBYTES[9].a/w2892 ), .Z(n16603) );
  XOR \SUBBYTES[9].a/U4847  ( .A(\SUBBYTES[9].a/w2875 ), .B(
        \SUBBYTES[9].a/w2877 ), .Z(n16604) );
  XOR \SUBBYTES[9].a/U4846  ( .A(n16606), .B(n16605), .Z(\SUBBYTES[9].a/w2899 ) );
  XOR \SUBBYTES[9].a/U4845  ( .A(n17243), .B(n16607), .Z(n16605) );
  XOR \SUBBYTES[9].a/U4844  ( .A(\w1[9][21] ), .B(n17244), .Z(n16606) );
  XOR \SUBBYTES[9].a/U4843  ( .A(\SUBBYTES[9].a/w2889 ), .B(
        \SUBBYTES[9].a/w2890 ), .Z(n16607) );
  XOR \SUBBYTES[9].a/U4842  ( .A(n16609), .B(n16608), .Z(\SUBBYTES[9].a/w2915 ) );
  XOR \SUBBYTES[9].a/U4841  ( .A(\w1[9][17] ), .B(n16610), .Z(n16608) );
  XOR \SUBBYTES[9].a/U4840  ( .A(\SUBBYTES[9].a/w2890 ), .B(
        \SUBBYTES[9].a/w2892 ), .Z(n16609) );
  XOR \SUBBYTES[9].a/U4839  ( .A(\SUBBYTES[9].a/w2874 ), .B(
        \SUBBYTES[9].a/w2875 ), .Z(n16610) );
  XOR \SUBBYTES[9].a/U4838  ( .A(\w1[9][25] ), .B(n16611), .Z(n17245) );
  XOR \SUBBYTES[9].a/U4837  ( .A(\w1[9][27] ), .B(\w1[9][26] ), .Z(n16611) );
  XOR \SUBBYTES[9].a/U4836  ( .A(\w1[9][30] ), .B(n17245), .Z(
        \SUBBYTES[9].a/w2757 ) );
  XOR \SUBBYTES[9].a/U4835  ( .A(\w1[9][24] ), .B(\SUBBYTES[9].a/w2757 ), .Z(
        \SUBBYTES[9].a/w2644 ) );
  XOR \SUBBYTES[9].a/U4834  ( .A(\w1[9][24] ), .B(n16612), .Z(
        \SUBBYTES[9].a/w2645 ) );
  XOR \SUBBYTES[9].a/U4833  ( .A(\w1[9][30] ), .B(\w1[9][29] ), .Z(n16612) );
  XOR \SUBBYTES[9].a/U4832  ( .A(\w1[9][29] ), .B(n17245), .Z(
        \SUBBYTES[9].a/w2775 ) );
  XOR \SUBBYTES[9].a/U4831  ( .A(n16614), .B(n16613), .Z(\SUBBYTES[9].a/w2768 ) );
  XOR \SUBBYTES[9].a/U4830  ( .A(\w1[9][27] ), .B(\w1[9][25] ), .Z(n16613) );
  XOR \SUBBYTES[9].a/U4829  ( .A(\w1[9][31] ), .B(\w1[9][28] ), .Z(n16614) );
  XOR \SUBBYTES[9].a/U4828  ( .A(\w1[9][24] ), .B(\SUBBYTES[9].a/w2768 ), .Z(
        \SUBBYTES[9].a/w2647 ) );
  XOR \SUBBYTES[9].a/U4827  ( .A(n16616), .B(n16615), .Z(\SUBBYTES[9].a/w2755 ) );
  XOR \SUBBYTES[9].a/U4826  ( .A(\SUBBYTES[9].a/w2716 ), .B(n1097), .Z(n16615)
         );
  XOR \SUBBYTES[9].a/U4825  ( .A(\SUBBYTES[9].a/w2709 ), .B(
        \SUBBYTES[9].a/w2712 ), .Z(n16616) );
  XOR \SUBBYTES[9].a/U4824  ( .A(n16618), .B(n16617), .Z(\SUBBYTES[9].a/w2756 ) );
  XOR \SUBBYTES[9].a/U4823  ( .A(\SUBBYTES[9].a/w2716 ), .B(n16097), .Z(n16617) );
  XOR \SUBBYTES[9].a/U4822  ( .A(\SUBBYTES[9].a/w2709 ), .B(n16096), .Z(n16618) );
  XOR \SUBBYTES[9].a/U4821  ( .A(\SUBBYTES[9].a/w2768 ), .B(n16619), .Z(
        \SUBBYTES[9].a/w2758 ) );
  XOR \SUBBYTES[9].a/U4820  ( .A(\w1[9][30] ), .B(\w1[9][29] ), .Z(n16619) );
  XOR \SUBBYTES[9].a/U4819  ( .A(n16621), .B(n16620), .Z(\SUBBYTES[9].a/w2759 ) );
  XOR \SUBBYTES[9].a/U4818  ( .A(n16097), .B(n1097), .Z(n16620) );
  XOR \SUBBYTES[9].a/U4817  ( .A(n16096), .B(\SUBBYTES[9].a/w2712 ), .Z(n16621) );
  XOR \SUBBYTES[9].a/U4816  ( .A(\w1[9][31] ), .B(\w1[9][26] ), .Z(n17251) );
  XOR \SUBBYTES[9].a/U4815  ( .A(n17251), .B(n16622), .Z(\SUBBYTES[9].a/w2760 ) );
  XOR \SUBBYTES[9].a/U4814  ( .A(\w1[9][29] ), .B(\w1[9][28] ), .Z(n16622) );
  XOR \SUBBYTES[9].a/U4813  ( .A(\w1[9][31] ), .B(\SUBBYTES[9].a/w2645 ), .Z(
        \SUBBYTES[9].a/w2648 ) );
  XOR \SUBBYTES[9].a/U4812  ( .A(\w1[9][25] ), .B(\SUBBYTES[9].a/w2645 ), .Z(
        \SUBBYTES[9].a/w2649 ) );
  XOR \SUBBYTES[9].a/U4811  ( .A(\w1[9][28] ), .B(\SUBBYTES[9].a/w2645 ), .Z(
        \SUBBYTES[9].a/w2650 ) );
  XOR \SUBBYTES[9].a/U4810  ( .A(\SUBBYTES[9].a/w2649 ), .B(n17251), .Z(
        \SUBBYTES[9].a/w2651 ) );
  XOR \SUBBYTES[9].a/U4809  ( .A(n17251), .B(n16623), .Z(\SUBBYTES[9].a/w2736 ) );
  XOR \SUBBYTES[9].a/U4808  ( .A(\w1[9][28] ), .B(\w1[9][25] ), .Z(n16623) );
  XOR \SUBBYTES[9].a/U4807  ( .A(n16625), .B(n16624), .Z(n17248) );
  XOR \SUBBYTES[9].a/U4806  ( .A(\w1[9][28] ), .B(n16626), .Z(n16624) );
  XOR \SUBBYTES[9].a/U4805  ( .A(\SUBBYTES[9].a/w2701 ), .B(\w1[9][30] ), .Z(
        n16625) );
  XOR \SUBBYTES[9].a/U4804  ( .A(\SUBBYTES[9].a/w2675 ), .B(
        \SUBBYTES[9].a/w2682 ), .Z(n16626) );
  XOR \SUBBYTES[9].a/U4803  ( .A(n16628), .B(n16627), .Z(n17246) );
  XOR \SUBBYTES[9].a/U4802  ( .A(\w1[9][25] ), .B(n16629), .Z(n16627) );
  XOR \SUBBYTES[9].a/U4801  ( .A(\SUBBYTES[9].a/w2700 ), .B(\w1[9][29] ), .Z(
        n16628) );
  XOR \SUBBYTES[9].a/U4800  ( .A(\SUBBYTES[9].a/w2676 ), .B(
        \SUBBYTES[9].a/w2683 ), .Z(n16629) );
  XOR \SUBBYTES[9].a/U4799  ( .A(n17248), .B(n17246), .Z(\SUBBYTES[9].a/w2706 ) );
  XOR \SUBBYTES[9].a/U4798  ( .A(\w1[9][29] ), .B(n16630), .Z(n17249) );
  XOR \SUBBYTES[9].a/U4797  ( .A(\SUBBYTES[9].a/w2668 ), .B(
        \SUBBYTES[9].a/w2678 ), .Z(n16630) );
  XOR \SUBBYTES[9].a/U4796  ( .A(n16632), .B(n16631), .Z(\SUBBYTES[9].a/w2693 ) );
  XOR \SUBBYTES[9].a/U4795  ( .A(n17249), .B(n16633), .Z(n16631) );
  XOR \SUBBYTES[9].a/U4794  ( .A(\w1[9][28] ), .B(\SUBBYTES[9].a/w2757 ), .Z(
        n16632) );
  XOR \SUBBYTES[9].a/U4793  ( .A(\SUBBYTES[9].a/w2670 ), .B(
        \SUBBYTES[9].a/w2675 ), .Z(n16633) );
  XOR \SUBBYTES[9].a/U4792  ( .A(n16635), .B(n16634), .Z(n17247) );
  XOR \SUBBYTES[9].a/U4791  ( .A(\SUBBYTES[9].a/w2703 ), .B(\w1[9][31] ), .Z(
        n16634) );
  XOR \SUBBYTES[9].a/U4790  ( .A(\SUBBYTES[9].a/w2678 ), .B(
        \SUBBYTES[9].a/w2685 ), .Z(n16635) );
  XOR \SUBBYTES[9].a/U4789  ( .A(n17246), .B(n17247), .Z(\SUBBYTES[9].a/w2705 ) );
  XOR \SUBBYTES[9].a/U4788  ( .A(\w1[9][27] ), .B(n16636), .Z(n17250) );
  XOR \SUBBYTES[9].a/U4787  ( .A(\SUBBYTES[9].a/w2667 ), .B(
        \SUBBYTES[9].a/w2670 ), .Z(n16636) );
  XOR \SUBBYTES[9].a/U4786  ( .A(n16638), .B(n16637), .Z(\SUBBYTES[9].a/w2694 ) );
  XOR \SUBBYTES[9].a/U4785  ( .A(n17250), .B(n16639), .Z(n16637) );
  XOR \SUBBYTES[9].a/U4784  ( .A(\w1[9][30] ), .B(\SUBBYTES[9].a/w2736 ), .Z(
        n16638) );
  XOR \SUBBYTES[9].a/U4783  ( .A(\SUBBYTES[9].a/w2675 ), .B(
        \SUBBYTES[9].a/w2676 ), .Z(n16639) );
  XOR \SUBBYTES[9].a/U4782  ( .A(n17248), .B(n17247), .Z(\SUBBYTES[9].a/w2714 ) );
  XOR \SUBBYTES[9].a/U4781  ( .A(n16641), .B(n16640), .Z(\SUBBYTES[9].a/w2715 ) );
  XOR \SUBBYTES[9].a/U4780  ( .A(\w1[9][31] ), .B(n17249), .Z(n16640) );
  XOR \SUBBYTES[9].a/U4779  ( .A(\SUBBYTES[9].a/w2667 ), .B(
        \SUBBYTES[9].a/w2676 ), .Z(n16641) );
  XOR \SUBBYTES[9].a/U4778  ( .A(n16643), .B(n16642), .Z(\SUBBYTES[9].a/w2691 ) );
  XOR \SUBBYTES[9].a/U4777  ( .A(n16645), .B(n16644), .Z(n16642) );
  XOR \SUBBYTES[9].a/U4776  ( .A(\w1[9][31] ), .B(\SUBBYTES[9].a/w2775 ), .Z(
        n16643) );
  XOR \SUBBYTES[9].a/U4775  ( .A(\SUBBYTES[9].a/w2682 ), .B(
        \SUBBYTES[9].a/w2685 ), .Z(n16644) );
  XOR \SUBBYTES[9].a/U4774  ( .A(\SUBBYTES[9].a/w2668 ), .B(
        \SUBBYTES[9].a/w2670 ), .Z(n16645) );
  XOR \SUBBYTES[9].a/U4773  ( .A(n16647), .B(n16646), .Z(\SUBBYTES[9].a/w2692 ) );
  XOR \SUBBYTES[9].a/U4772  ( .A(n17250), .B(n16648), .Z(n16646) );
  XOR \SUBBYTES[9].a/U4771  ( .A(\w1[9][29] ), .B(n17251), .Z(n16647) );
  XOR \SUBBYTES[9].a/U4770  ( .A(\SUBBYTES[9].a/w2682 ), .B(
        \SUBBYTES[9].a/w2683 ), .Z(n16648) );
  XOR \SUBBYTES[9].a/U4769  ( .A(n16650), .B(n16649), .Z(\SUBBYTES[9].a/w2708 ) );
  XOR \SUBBYTES[9].a/U4768  ( .A(\w1[9][25] ), .B(n16651), .Z(n16649) );
  XOR \SUBBYTES[9].a/U4767  ( .A(\SUBBYTES[9].a/w2683 ), .B(
        \SUBBYTES[9].a/w2685 ), .Z(n16650) );
  XOR \SUBBYTES[9].a/U4766  ( .A(\SUBBYTES[9].a/w2667 ), .B(
        \SUBBYTES[9].a/w2668 ), .Z(n16651) );
  XOR \SUBBYTES[9].a/U4765  ( .A(\w1[9][33] ), .B(n16652), .Z(n17252) );
  XOR \SUBBYTES[9].a/U4764  ( .A(\w1[9][35] ), .B(\w1[9][34] ), .Z(n16652) );
  XOR \SUBBYTES[9].a/U4763  ( .A(\w1[9][38] ), .B(n17252), .Z(
        \SUBBYTES[9].a/w2550 ) );
  XOR \SUBBYTES[9].a/U4762  ( .A(\w1[9][32] ), .B(\SUBBYTES[9].a/w2550 ), .Z(
        \SUBBYTES[9].a/w2437 ) );
  XOR \SUBBYTES[9].a/U4761  ( .A(\w1[9][32] ), .B(n16653), .Z(
        \SUBBYTES[9].a/w2438 ) );
  XOR \SUBBYTES[9].a/U4760  ( .A(\w1[9][38] ), .B(\w1[9][37] ), .Z(n16653) );
  XOR \SUBBYTES[9].a/U4759  ( .A(\w1[9][37] ), .B(n17252), .Z(
        \SUBBYTES[9].a/w2568 ) );
  XOR \SUBBYTES[9].a/U4758  ( .A(n16655), .B(n16654), .Z(\SUBBYTES[9].a/w2561 ) );
  XOR \SUBBYTES[9].a/U4757  ( .A(\w1[9][35] ), .B(\w1[9][33] ), .Z(n16654) );
  XOR \SUBBYTES[9].a/U4756  ( .A(\w1[9][39] ), .B(\w1[9][36] ), .Z(n16655) );
  XOR \SUBBYTES[9].a/U4755  ( .A(\w1[9][32] ), .B(\SUBBYTES[9].a/w2561 ), .Z(
        \SUBBYTES[9].a/w2440 ) );
  XOR \SUBBYTES[9].a/U4754  ( .A(n16657), .B(n16656), .Z(\SUBBYTES[9].a/w2548 ) );
  XOR \SUBBYTES[9].a/U4753  ( .A(\SUBBYTES[9].a/w2509 ), .B(n1096), .Z(n16656)
         );
  XOR \SUBBYTES[9].a/U4752  ( .A(\SUBBYTES[9].a/w2502 ), .B(
        \SUBBYTES[9].a/w2505 ), .Z(n16657) );
  XOR \SUBBYTES[9].a/U4751  ( .A(n16659), .B(n16658), .Z(\SUBBYTES[9].a/w2549 ) );
  XOR \SUBBYTES[9].a/U4750  ( .A(\SUBBYTES[9].a/w2509 ), .B(n16095), .Z(n16658) );
  XOR \SUBBYTES[9].a/U4749  ( .A(\SUBBYTES[9].a/w2502 ), .B(n16094), .Z(n16659) );
  XOR \SUBBYTES[9].a/U4748  ( .A(\SUBBYTES[9].a/w2561 ), .B(n16660), .Z(
        \SUBBYTES[9].a/w2551 ) );
  XOR \SUBBYTES[9].a/U4747  ( .A(\w1[9][38] ), .B(\w1[9][37] ), .Z(n16660) );
  XOR \SUBBYTES[9].a/U4746  ( .A(n16662), .B(n16661), .Z(\SUBBYTES[9].a/w2552 ) );
  XOR \SUBBYTES[9].a/U4745  ( .A(n16095), .B(n1096), .Z(n16661) );
  XOR \SUBBYTES[9].a/U4744  ( .A(n16094), .B(\SUBBYTES[9].a/w2505 ), .Z(n16662) );
  XOR \SUBBYTES[9].a/U4743  ( .A(\w1[9][39] ), .B(\w1[9][34] ), .Z(n17258) );
  XOR \SUBBYTES[9].a/U4742  ( .A(n17258), .B(n16663), .Z(\SUBBYTES[9].a/w2553 ) );
  XOR \SUBBYTES[9].a/U4741  ( .A(\w1[9][37] ), .B(\w1[9][36] ), .Z(n16663) );
  XOR \SUBBYTES[9].a/U4740  ( .A(\w1[9][39] ), .B(\SUBBYTES[9].a/w2438 ), .Z(
        \SUBBYTES[9].a/w2441 ) );
  XOR \SUBBYTES[9].a/U4739  ( .A(\w1[9][33] ), .B(\SUBBYTES[9].a/w2438 ), .Z(
        \SUBBYTES[9].a/w2442 ) );
  XOR \SUBBYTES[9].a/U4738  ( .A(\w1[9][36] ), .B(\SUBBYTES[9].a/w2438 ), .Z(
        \SUBBYTES[9].a/w2443 ) );
  XOR \SUBBYTES[9].a/U4737  ( .A(\SUBBYTES[9].a/w2442 ), .B(n17258), .Z(
        \SUBBYTES[9].a/w2444 ) );
  XOR \SUBBYTES[9].a/U4736  ( .A(n17258), .B(n16664), .Z(\SUBBYTES[9].a/w2529 ) );
  XOR \SUBBYTES[9].a/U4735  ( .A(\w1[9][36] ), .B(\w1[9][33] ), .Z(n16664) );
  XOR \SUBBYTES[9].a/U4734  ( .A(n16666), .B(n16665), .Z(n17255) );
  XOR \SUBBYTES[9].a/U4733  ( .A(\w1[9][36] ), .B(n16667), .Z(n16665) );
  XOR \SUBBYTES[9].a/U4732  ( .A(\SUBBYTES[9].a/w2494 ), .B(\w1[9][38] ), .Z(
        n16666) );
  XOR \SUBBYTES[9].a/U4731  ( .A(\SUBBYTES[9].a/w2468 ), .B(
        \SUBBYTES[9].a/w2475 ), .Z(n16667) );
  XOR \SUBBYTES[9].a/U4730  ( .A(n16669), .B(n16668), .Z(n17253) );
  XOR \SUBBYTES[9].a/U4729  ( .A(\w1[9][33] ), .B(n16670), .Z(n16668) );
  XOR \SUBBYTES[9].a/U4728  ( .A(\SUBBYTES[9].a/w2493 ), .B(\w1[9][37] ), .Z(
        n16669) );
  XOR \SUBBYTES[9].a/U4727  ( .A(\SUBBYTES[9].a/w2469 ), .B(
        \SUBBYTES[9].a/w2476 ), .Z(n16670) );
  XOR \SUBBYTES[9].a/U4726  ( .A(n17255), .B(n17253), .Z(\SUBBYTES[9].a/w2499 ) );
  XOR \SUBBYTES[9].a/U4725  ( .A(\w1[9][37] ), .B(n16671), .Z(n17256) );
  XOR \SUBBYTES[9].a/U4724  ( .A(\SUBBYTES[9].a/w2461 ), .B(
        \SUBBYTES[9].a/w2471 ), .Z(n16671) );
  XOR \SUBBYTES[9].a/U4723  ( .A(n16673), .B(n16672), .Z(\SUBBYTES[9].a/w2486 ) );
  XOR \SUBBYTES[9].a/U4722  ( .A(n17256), .B(n16674), .Z(n16672) );
  XOR \SUBBYTES[9].a/U4721  ( .A(\w1[9][36] ), .B(\SUBBYTES[9].a/w2550 ), .Z(
        n16673) );
  XOR \SUBBYTES[9].a/U4720  ( .A(\SUBBYTES[9].a/w2463 ), .B(
        \SUBBYTES[9].a/w2468 ), .Z(n16674) );
  XOR \SUBBYTES[9].a/U4719  ( .A(n16676), .B(n16675), .Z(n17254) );
  XOR \SUBBYTES[9].a/U4718  ( .A(\SUBBYTES[9].a/w2496 ), .B(\w1[9][39] ), .Z(
        n16675) );
  XOR \SUBBYTES[9].a/U4717  ( .A(\SUBBYTES[9].a/w2471 ), .B(
        \SUBBYTES[9].a/w2478 ), .Z(n16676) );
  XOR \SUBBYTES[9].a/U4716  ( .A(n17253), .B(n17254), .Z(\SUBBYTES[9].a/w2498 ) );
  XOR \SUBBYTES[9].a/U4715  ( .A(\w1[9][35] ), .B(n16677), .Z(n17257) );
  XOR \SUBBYTES[9].a/U4714  ( .A(\SUBBYTES[9].a/w2460 ), .B(
        \SUBBYTES[9].a/w2463 ), .Z(n16677) );
  XOR \SUBBYTES[9].a/U4713  ( .A(n16679), .B(n16678), .Z(\SUBBYTES[9].a/w2487 ) );
  XOR \SUBBYTES[9].a/U4712  ( .A(n17257), .B(n16680), .Z(n16678) );
  XOR \SUBBYTES[9].a/U4711  ( .A(\w1[9][38] ), .B(\SUBBYTES[9].a/w2529 ), .Z(
        n16679) );
  XOR \SUBBYTES[9].a/U4710  ( .A(\SUBBYTES[9].a/w2468 ), .B(
        \SUBBYTES[9].a/w2469 ), .Z(n16680) );
  XOR \SUBBYTES[9].a/U4709  ( .A(n17255), .B(n17254), .Z(\SUBBYTES[9].a/w2507 ) );
  XOR \SUBBYTES[9].a/U4708  ( .A(n16682), .B(n16681), .Z(\SUBBYTES[9].a/w2508 ) );
  XOR \SUBBYTES[9].a/U4707  ( .A(\w1[9][39] ), .B(n17256), .Z(n16681) );
  XOR \SUBBYTES[9].a/U4706  ( .A(\SUBBYTES[9].a/w2460 ), .B(
        \SUBBYTES[9].a/w2469 ), .Z(n16682) );
  XOR \SUBBYTES[9].a/U4705  ( .A(n16684), .B(n16683), .Z(\SUBBYTES[9].a/w2484 ) );
  XOR \SUBBYTES[9].a/U4704  ( .A(n16686), .B(n16685), .Z(n16683) );
  XOR \SUBBYTES[9].a/U4703  ( .A(\w1[9][39] ), .B(\SUBBYTES[9].a/w2568 ), .Z(
        n16684) );
  XOR \SUBBYTES[9].a/U4702  ( .A(\SUBBYTES[9].a/w2475 ), .B(
        \SUBBYTES[9].a/w2478 ), .Z(n16685) );
  XOR \SUBBYTES[9].a/U4701  ( .A(\SUBBYTES[9].a/w2461 ), .B(
        \SUBBYTES[9].a/w2463 ), .Z(n16686) );
  XOR \SUBBYTES[9].a/U4700  ( .A(n16688), .B(n16687), .Z(\SUBBYTES[9].a/w2485 ) );
  XOR \SUBBYTES[9].a/U4699  ( .A(n17257), .B(n16689), .Z(n16687) );
  XOR \SUBBYTES[9].a/U4698  ( .A(\w1[9][37] ), .B(n17258), .Z(n16688) );
  XOR \SUBBYTES[9].a/U4697  ( .A(\SUBBYTES[9].a/w2475 ), .B(
        \SUBBYTES[9].a/w2476 ), .Z(n16689) );
  XOR \SUBBYTES[9].a/U4696  ( .A(n16691), .B(n16690), .Z(\SUBBYTES[9].a/w2501 ) );
  XOR \SUBBYTES[9].a/U4695  ( .A(\w1[9][33] ), .B(n16692), .Z(n16690) );
  XOR \SUBBYTES[9].a/U4694  ( .A(\SUBBYTES[9].a/w2476 ), .B(
        \SUBBYTES[9].a/w2478 ), .Z(n16691) );
  XOR \SUBBYTES[9].a/U4693  ( .A(\SUBBYTES[9].a/w2460 ), .B(
        \SUBBYTES[9].a/w2461 ), .Z(n16692) );
  XOR \SUBBYTES[9].a/U4692  ( .A(\w1[9][41] ), .B(n16693), .Z(n17259) );
  XOR \SUBBYTES[9].a/U4691  ( .A(\w1[9][43] ), .B(\w1[9][42] ), .Z(n16693) );
  XOR \SUBBYTES[9].a/U4690  ( .A(\w1[9][46] ), .B(n17259), .Z(
        \SUBBYTES[9].a/w2343 ) );
  XOR \SUBBYTES[9].a/U4689  ( .A(\w1[9][40] ), .B(\SUBBYTES[9].a/w2343 ), .Z(
        \SUBBYTES[9].a/w2230 ) );
  XOR \SUBBYTES[9].a/U4688  ( .A(\w1[9][40] ), .B(n16694), .Z(
        \SUBBYTES[9].a/w2231 ) );
  XOR \SUBBYTES[9].a/U4687  ( .A(\w1[9][46] ), .B(\w1[9][45] ), .Z(n16694) );
  XOR \SUBBYTES[9].a/U4686  ( .A(\w1[9][45] ), .B(n17259), .Z(
        \SUBBYTES[9].a/w2361 ) );
  XOR \SUBBYTES[9].a/U4685  ( .A(n16696), .B(n16695), .Z(\SUBBYTES[9].a/w2354 ) );
  XOR \SUBBYTES[9].a/U4684  ( .A(\w1[9][43] ), .B(\w1[9][41] ), .Z(n16695) );
  XOR \SUBBYTES[9].a/U4683  ( .A(\w1[9][47] ), .B(\w1[9][44] ), .Z(n16696) );
  XOR \SUBBYTES[9].a/U4682  ( .A(\w1[9][40] ), .B(\SUBBYTES[9].a/w2354 ), .Z(
        \SUBBYTES[9].a/w2233 ) );
  XOR \SUBBYTES[9].a/U4681  ( .A(n16698), .B(n16697), .Z(\SUBBYTES[9].a/w2341 ) );
  XOR \SUBBYTES[9].a/U4680  ( .A(\SUBBYTES[9].a/w2302 ), .B(n1095), .Z(n16697)
         );
  XOR \SUBBYTES[9].a/U4679  ( .A(\SUBBYTES[9].a/w2295 ), .B(
        \SUBBYTES[9].a/w2298 ), .Z(n16698) );
  XOR \SUBBYTES[9].a/U4678  ( .A(n16700), .B(n16699), .Z(\SUBBYTES[9].a/w2342 ) );
  XOR \SUBBYTES[9].a/U4677  ( .A(\SUBBYTES[9].a/w2302 ), .B(n16093), .Z(n16699) );
  XOR \SUBBYTES[9].a/U4676  ( .A(\SUBBYTES[9].a/w2295 ), .B(n16092), .Z(n16700) );
  XOR \SUBBYTES[9].a/U4675  ( .A(\SUBBYTES[9].a/w2354 ), .B(n16701), .Z(
        \SUBBYTES[9].a/w2344 ) );
  XOR \SUBBYTES[9].a/U4674  ( .A(\w1[9][46] ), .B(\w1[9][45] ), .Z(n16701) );
  XOR \SUBBYTES[9].a/U4673  ( .A(n16703), .B(n16702), .Z(\SUBBYTES[9].a/w2345 ) );
  XOR \SUBBYTES[9].a/U4672  ( .A(n16093), .B(n1095), .Z(n16702) );
  XOR \SUBBYTES[9].a/U4671  ( .A(n16092), .B(\SUBBYTES[9].a/w2298 ), .Z(n16703) );
  XOR \SUBBYTES[9].a/U4670  ( .A(\w1[9][47] ), .B(\w1[9][42] ), .Z(n17265) );
  XOR \SUBBYTES[9].a/U4669  ( .A(n17265), .B(n16704), .Z(\SUBBYTES[9].a/w2346 ) );
  XOR \SUBBYTES[9].a/U4668  ( .A(\w1[9][45] ), .B(\w1[9][44] ), .Z(n16704) );
  XOR \SUBBYTES[9].a/U4667  ( .A(\w1[9][47] ), .B(\SUBBYTES[9].a/w2231 ), .Z(
        \SUBBYTES[9].a/w2234 ) );
  XOR \SUBBYTES[9].a/U4666  ( .A(\w1[9][41] ), .B(\SUBBYTES[9].a/w2231 ), .Z(
        \SUBBYTES[9].a/w2235 ) );
  XOR \SUBBYTES[9].a/U4665  ( .A(\w1[9][44] ), .B(\SUBBYTES[9].a/w2231 ), .Z(
        \SUBBYTES[9].a/w2236 ) );
  XOR \SUBBYTES[9].a/U4664  ( .A(\SUBBYTES[9].a/w2235 ), .B(n17265), .Z(
        \SUBBYTES[9].a/w2237 ) );
  XOR \SUBBYTES[9].a/U4663  ( .A(n17265), .B(n16705), .Z(\SUBBYTES[9].a/w2322 ) );
  XOR \SUBBYTES[9].a/U4662  ( .A(\w1[9][44] ), .B(\w1[9][41] ), .Z(n16705) );
  XOR \SUBBYTES[9].a/U4661  ( .A(n16707), .B(n16706), .Z(n17262) );
  XOR \SUBBYTES[9].a/U4660  ( .A(\w1[9][44] ), .B(n16708), .Z(n16706) );
  XOR \SUBBYTES[9].a/U4659  ( .A(\SUBBYTES[9].a/w2287 ), .B(\w1[9][46] ), .Z(
        n16707) );
  XOR \SUBBYTES[9].a/U4658  ( .A(\SUBBYTES[9].a/w2261 ), .B(
        \SUBBYTES[9].a/w2268 ), .Z(n16708) );
  XOR \SUBBYTES[9].a/U4657  ( .A(n16710), .B(n16709), .Z(n17260) );
  XOR \SUBBYTES[9].a/U4656  ( .A(\w1[9][41] ), .B(n16711), .Z(n16709) );
  XOR \SUBBYTES[9].a/U4655  ( .A(\SUBBYTES[9].a/w2286 ), .B(\w1[9][45] ), .Z(
        n16710) );
  XOR \SUBBYTES[9].a/U4654  ( .A(\SUBBYTES[9].a/w2262 ), .B(
        \SUBBYTES[9].a/w2269 ), .Z(n16711) );
  XOR \SUBBYTES[9].a/U4653  ( .A(n17262), .B(n17260), .Z(\SUBBYTES[9].a/w2292 ) );
  XOR \SUBBYTES[9].a/U4652  ( .A(\w1[9][45] ), .B(n16712), .Z(n17263) );
  XOR \SUBBYTES[9].a/U4651  ( .A(\SUBBYTES[9].a/w2254 ), .B(
        \SUBBYTES[9].a/w2264 ), .Z(n16712) );
  XOR \SUBBYTES[9].a/U4650  ( .A(n16714), .B(n16713), .Z(\SUBBYTES[9].a/w2279 ) );
  XOR \SUBBYTES[9].a/U4649  ( .A(n17263), .B(n16715), .Z(n16713) );
  XOR \SUBBYTES[9].a/U4648  ( .A(\w1[9][44] ), .B(\SUBBYTES[9].a/w2343 ), .Z(
        n16714) );
  XOR \SUBBYTES[9].a/U4647  ( .A(\SUBBYTES[9].a/w2256 ), .B(
        \SUBBYTES[9].a/w2261 ), .Z(n16715) );
  XOR \SUBBYTES[9].a/U4646  ( .A(n16717), .B(n16716), .Z(n17261) );
  XOR \SUBBYTES[9].a/U4645  ( .A(\SUBBYTES[9].a/w2289 ), .B(\w1[9][47] ), .Z(
        n16716) );
  XOR \SUBBYTES[9].a/U4644  ( .A(\SUBBYTES[9].a/w2264 ), .B(
        \SUBBYTES[9].a/w2271 ), .Z(n16717) );
  XOR \SUBBYTES[9].a/U4643  ( .A(n17260), .B(n17261), .Z(\SUBBYTES[9].a/w2291 ) );
  XOR \SUBBYTES[9].a/U4642  ( .A(\w1[9][43] ), .B(n16718), .Z(n17264) );
  XOR \SUBBYTES[9].a/U4641  ( .A(\SUBBYTES[9].a/w2253 ), .B(
        \SUBBYTES[9].a/w2256 ), .Z(n16718) );
  XOR \SUBBYTES[9].a/U4640  ( .A(n16720), .B(n16719), .Z(\SUBBYTES[9].a/w2280 ) );
  XOR \SUBBYTES[9].a/U4639  ( .A(n17264), .B(n16721), .Z(n16719) );
  XOR \SUBBYTES[9].a/U4638  ( .A(\w1[9][46] ), .B(\SUBBYTES[9].a/w2322 ), .Z(
        n16720) );
  XOR \SUBBYTES[9].a/U4637  ( .A(\SUBBYTES[9].a/w2261 ), .B(
        \SUBBYTES[9].a/w2262 ), .Z(n16721) );
  XOR \SUBBYTES[9].a/U4636  ( .A(n17262), .B(n17261), .Z(\SUBBYTES[9].a/w2300 ) );
  XOR \SUBBYTES[9].a/U4635  ( .A(n16723), .B(n16722), .Z(\SUBBYTES[9].a/w2301 ) );
  XOR \SUBBYTES[9].a/U4634  ( .A(\w1[9][47] ), .B(n17263), .Z(n16722) );
  XOR \SUBBYTES[9].a/U4633  ( .A(\SUBBYTES[9].a/w2253 ), .B(
        \SUBBYTES[9].a/w2262 ), .Z(n16723) );
  XOR \SUBBYTES[9].a/U4632  ( .A(n16725), .B(n16724), .Z(\SUBBYTES[9].a/w2277 ) );
  XOR \SUBBYTES[9].a/U4631  ( .A(n16727), .B(n16726), .Z(n16724) );
  XOR \SUBBYTES[9].a/U4630  ( .A(\w1[9][47] ), .B(\SUBBYTES[9].a/w2361 ), .Z(
        n16725) );
  XOR \SUBBYTES[9].a/U4629  ( .A(\SUBBYTES[9].a/w2268 ), .B(
        \SUBBYTES[9].a/w2271 ), .Z(n16726) );
  XOR \SUBBYTES[9].a/U4628  ( .A(\SUBBYTES[9].a/w2254 ), .B(
        \SUBBYTES[9].a/w2256 ), .Z(n16727) );
  XOR \SUBBYTES[9].a/U4627  ( .A(n16729), .B(n16728), .Z(\SUBBYTES[9].a/w2278 ) );
  XOR \SUBBYTES[9].a/U4626  ( .A(n17264), .B(n16730), .Z(n16728) );
  XOR \SUBBYTES[9].a/U4625  ( .A(\w1[9][45] ), .B(n17265), .Z(n16729) );
  XOR \SUBBYTES[9].a/U4624  ( .A(\SUBBYTES[9].a/w2268 ), .B(
        \SUBBYTES[9].a/w2269 ), .Z(n16730) );
  XOR \SUBBYTES[9].a/U4623  ( .A(n16732), .B(n16731), .Z(\SUBBYTES[9].a/w2294 ) );
  XOR \SUBBYTES[9].a/U4622  ( .A(\w1[9][41] ), .B(n16733), .Z(n16731) );
  XOR \SUBBYTES[9].a/U4621  ( .A(\SUBBYTES[9].a/w2269 ), .B(
        \SUBBYTES[9].a/w2271 ), .Z(n16732) );
  XOR \SUBBYTES[9].a/U4620  ( .A(\SUBBYTES[9].a/w2253 ), .B(
        \SUBBYTES[9].a/w2254 ), .Z(n16733) );
  XOR \SUBBYTES[9].a/U4619  ( .A(\w1[9][49] ), .B(n16734), .Z(n17266) );
  XOR \SUBBYTES[9].a/U4618  ( .A(\w1[9][51] ), .B(\w1[9][50] ), .Z(n16734) );
  XOR \SUBBYTES[9].a/U4617  ( .A(\w1[9][54] ), .B(n17266), .Z(
        \SUBBYTES[9].a/w2136 ) );
  XOR \SUBBYTES[9].a/U4616  ( .A(\w1[9][48] ), .B(\SUBBYTES[9].a/w2136 ), .Z(
        \SUBBYTES[9].a/w2023 ) );
  XOR \SUBBYTES[9].a/U4615  ( .A(\w1[9][48] ), .B(n16735), .Z(
        \SUBBYTES[9].a/w2024 ) );
  XOR \SUBBYTES[9].a/U4614  ( .A(\w1[9][54] ), .B(\w1[9][53] ), .Z(n16735) );
  XOR \SUBBYTES[9].a/U4613  ( .A(\w1[9][53] ), .B(n17266), .Z(
        \SUBBYTES[9].a/w2154 ) );
  XOR \SUBBYTES[9].a/U4612  ( .A(n16737), .B(n16736), .Z(\SUBBYTES[9].a/w2147 ) );
  XOR \SUBBYTES[9].a/U4611  ( .A(\w1[9][51] ), .B(\w1[9][49] ), .Z(n16736) );
  XOR \SUBBYTES[9].a/U4610  ( .A(\w1[9][55] ), .B(\w1[9][52] ), .Z(n16737) );
  XOR \SUBBYTES[9].a/U4609  ( .A(\w1[9][48] ), .B(\SUBBYTES[9].a/w2147 ), .Z(
        \SUBBYTES[9].a/w2026 ) );
  XOR \SUBBYTES[9].a/U4608  ( .A(n16739), .B(n16738), .Z(\SUBBYTES[9].a/w2134 ) );
  XOR \SUBBYTES[9].a/U4607  ( .A(\SUBBYTES[9].a/w2095 ), .B(n1094), .Z(n16738)
         );
  XOR \SUBBYTES[9].a/U4606  ( .A(\SUBBYTES[9].a/w2088 ), .B(
        \SUBBYTES[9].a/w2091 ), .Z(n16739) );
  XOR \SUBBYTES[9].a/U4605  ( .A(n16741), .B(n16740), .Z(\SUBBYTES[9].a/w2135 ) );
  XOR \SUBBYTES[9].a/U4604  ( .A(\SUBBYTES[9].a/w2095 ), .B(n16091), .Z(n16740) );
  XOR \SUBBYTES[9].a/U4603  ( .A(\SUBBYTES[9].a/w2088 ), .B(n16090), .Z(n16741) );
  XOR \SUBBYTES[9].a/U4602  ( .A(\SUBBYTES[9].a/w2147 ), .B(n16742), .Z(
        \SUBBYTES[9].a/w2137 ) );
  XOR \SUBBYTES[9].a/U4601  ( .A(\w1[9][54] ), .B(\w1[9][53] ), .Z(n16742) );
  XOR \SUBBYTES[9].a/U4600  ( .A(n16744), .B(n16743), .Z(\SUBBYTES[9].a/w2138 ) );
  XOR \SUBBYTES[9].a/U4599  ( .A(n16091), .B(n1094), .Z(n16743) );
  XOR \SUBBYTES[9].a/U4598  ( .A(n16090), .B(\SUBBYTES[9].a/w2091 ), .Z(n16744) );
  XOR \SUBBYTES[9].a/U4597  ( .A(\w1[9][55] ), .B(\w1[9][50] ), .Z(n17272) );
  XOR \SUBBYTES[9].a/U4596  ( .A(n17272), .B(n16745), .Z(\SUBBYTES[9].a/w2139 ) );
  XOR \SUBBYTES[9].a/U4595  ( .A(\w1[9][53] ), .B(\w1[9][52] ), .Z(n16745) );
  XOR \SUBBYTES[9].a/U4594  ( .A(\w1[9][55] ), .B(\SUBBYTES[9].a/w2024 ), .Z(
        \SUBBYTES[9].a/w2027 ) );
  XOR \SUBBYTES[9].a/U4593  ( .A(\w1[9][49] ), .B(\SUBBYTES[9].a/w2024 ), .Z(
        \SUBBYTES[9].a/w2028 ) );
  XOR \SUBBYTES[9].a/U4592  ( .A(\w1[9][52] ), .B(\SUBBYTES[9].a/w2024 ), .Z(
        \SUBBYTES[9].a/w2029 ) );
  XOR \SUBBYTES[9].a/U4591  ( .A(\SUBBYTES[9].a/w2028 ), .B(n17272), .Z(
        \SUBBYTES[9].a/w2030 ) );
  XOR \SUBBYTES[9].a/U4590  ( .A(n17272), .B(n16746), .Z(\SUBBYTES[9].a/w2115 ) );
  XOR \SUBBYTES[9].a/U4589  ( .A(\w1[9][52] ), .B(\w1[9][49] ), .Z(n16746) );
  XOR \SUBBYTES[9].a/U4588  ( .A(n16748), .B(n16747), .Z(n17269) );
  XOR \SUBBYTES[9].a/U4587  ( .A(\w1[9][52] ), .B(n16749), .Z(n16747) );
  XOR \SUBBYTES[9].a/U4586  ( .A(\SUBBYTES[9].a/w2080 ), .B(\w1[9][54] ), .Z(
        n16748) );
  XOR \SUBBYTES[9].a/U4585  ( .A(\SUBBYTES[9].a/w2054 ), .B(
        \SUBBYTES[9].a/w2061 ), .Z(n16749) );
  XOR \SUBBYTES[9].a/U4584  ( .A(n16751), .B(n16750), .Z(n17267) );
  XOR \SUBBYTES[9].a/U4583  ( .A(\w1[9][49] ), .B(n16752), .Z(n16750) );
  XOR \SUBBYTES[9].a/U4582  ( .A(\SUBBYTES[9].a/w2079 ), .B(\w1[9][53] ), .Z(
        n16751) );
  XOR \SUBBYTES[9].a/U4581  ( .A(\SUBBYTES[9].a/w2055 ), .B(
        \SUBBYTES[9].a/w2062 ), .Z(n16752) );
  XOR \SUBBYTES[9].a/U4580  ( .A(n17269), .B(n17267), .Z(\SUBBYTES[9].a/w2085 ) );
  XOR \SUBBYTES[9].a/U4579  ( .A(\w1[9][53] ), .B(n16753), .Z(n17270) );
  XOR \SUBBYTES[9].a/U4578  ( .A(\SUBBYTES[9].a/w2047 ), .B(
        \SUBBYTES[9].a/w2057 ), .Z(n16753) );
  XOR \SUBBYTES[9].a/U4577  ( .A(n16755), .B(n16754), .Z(\SUBBYTES[9].a/w2072 ) );
  XOR \SUBBYTES[9].a/U4576  ( .A(n17270), .B(n16756), .Z(n16754) );
  XOR \SUBBYTES[9].a/U4575  ( .A(\w1[9][52] ), .B(\SUBBYTES[9].a/w2136 ), .Z(
        n16755) );
  XOR \SUBBYTES[9].a/U4574  ( .A(\SUBBYTES[9].a/w2049 ), .B(
        \SUBBYTES[9].a/w2054 ), .Z(n16756) );
  XOR \SUBBYTES[9].a/U4573  ( .A(n16758), .B(n16757), .Z(n17268) );
  XOR \SUBBYTES[9].a/U4572  ( .A(\SUBBYTES[9].a/w2082 ), .B(\w1[9][55] ), .Z(
        n16757) );
  XOR \SUBBYTES[9].a/U4571  ( .A(\SUBBYTES[9].a/w2057 ), .B(
        \SUBBYTES[9].a/w2064 ), .Z(n16758) );
  XOR \SUBBYTES[9].a/U4570  ( .A(n17267), .B(n17268), .Z(\SUBBYTES[9].a/w2084 ) );
  XOR \SUBBYTES[9].a/U4569  ( .A(\w1[9][51] ), .B(n16759), .Z(n17271) );
  XOR \SUBBYTES[9].a/U4568  ( .A(\SUBBYTES[9].a/w2046 ), .B(
        \SUBBYTES[9].a/w2049 ), .Z(n16759) );
  XOR \SUBBYTES[9].a/U4567  ( .A(n16761), .B(n16760), .Z(\SUBBYTES[9].a/w2073 ) );
  XOR \SUBBYTES[9].a/U4566  ( .A(n17271), .B(n16762), .Z(n16760) );
  XOR \SUBBYTES[9].a/U4565  ( .A(\w1[9][54] ), .B(\SUBBYTES[9].a/w2115 ), .Z(
        n16761) );
  XOR \SUBBYTES[9].a/U4564  ( .A(\SUBBYTES[9].a/w2054 ), .B(
        \SUBBYTES[9].a/w2055 ), .Z(n16762) );
  XOR \SUBBYTES[9].a/U4563  ( .A(n17269), .B(n17268), .Z(\SUBBYTES[9].a/w2093 ) );
  XOR \SUBBYTES[9].a/U4562  ( .A(n16764), .B(n16763), .Z(\SUBBYTES[9].a/w2094 ) );
  XOR \SUBBYTES[9].a/U4561  ( .A(\w1[9][55] ), .B(n17270), .Z(n16763) );
  XOR \SUBBYTES[9].a/U4560  ( .A(\SUBBYTES[9].a/w2046 ), .B(
        \SUBBYTES[9].a/w2055 ), .Z(n16764) );
  XOR \SUBBYTES[9].a/U4559  ( .A(n16766), .B(n16765), .Z(\SUBBYTES[9].a/w2070 ) );
  XOR \SUBBYTES[9].a/U4558  ( .A(n16768), .B(n16767), .Z(n16765) );
  XOR \SUBBYTES[9].a/U4557  ( .A(\w1[9][55] ), .B(\SUBBYTES[9].a/w2154 ), .Z(
        n16766) );
  XOR \SUBBYTES[9].a/U4556  ( .A(\SUBBYTES[9].a/w2061 ), .B(
        \SUBBYTES[9].a/w2064 ), .Z(n16767) );
  XOR \SUBBYTES[9].a/U4555  ( .A(\SUBBYTES[9].a/w2047 ), .B(
        \SUBBYTES[9].a/w2049 ), .Z(n16768) );
  XOR \SUBBYTES[9].a/U4554  ( .A(n16770), .B(n16769), .Z(\SUBBYTES[9].a/w2071 ) );
  XOR \SUBBYTES[9].a/U4553  ( .A(n17271), .B(n16771), .Z(n16769) );
  XOR \SUBBYTES[9].a/U4552  ( .A(\w1[9][53] ), .B(n17272), .Z(n16770) );
  XOR \SUBBYTES[9].a/U4551  ( .A(\SUBBYTES[9].a/w2061 ), .B(
        \SUBBYTES[9].a/w2062 ), .Z(n16771) );
  XOR \SUBBYTES[9].a/U4550  ( .A(n16773), .B(n16772), .Z(\SUBBYTES[9].a/w2087 ) );
  XOR \SUBBYTES[9].a/U4549  ( .A(\w1[9][49] ), .B(n16774), .Z(n16772) );
  XOR \SUBBYTES[9].a/U4548  ( .A(\SUBBYTES[9].a/w2062 ), .B(
        \SUBBYTES[9].a/w2064 ), .Z(n16773) );
  XOR \SUBBYTES[9].a/U4547  ( .A(\SUBBYTES[9].a/w2046 ), .B(
        \SUBBYTES[9].a/w2047 ), .Z(n16774) );
  XOR \SUBBYTES[9].a/U4546  ( .A(\w1[9][57] ), .B(n16775), .Z(n17273) );
  XOR \SUBBYTES[9].a/U4545  ( .A(\w1[9][59] ), .B(\w1[9][58] ), .Z(n16775) );
  XOR \SUBBYTES[9].a/U4544  ( .A(\w1[9][62] ), .B(n17273), .Z(
        \SUBBYTES[9].a/w1929 ) );
  XOR \SUBBYTES[9].a/U4543  ( .A(\w1[9][56] ), .B(\SUBBYTES[9].a/w1929 ), .Z(
        \SUBBYTES[9].a/w1816 ) );
  XOR \SUBBYTES[9].a/U4542  ( .A(\w1[9][56] ), .B(n16776), .Z(
        \SUBBYTES[9].a/w1817 ) );
  XOR \SUBBYTES[9].a/U4541  ( .A(\w1[9][62] ), .B(\w1[9][61] ), .Z(n16776) );
  XOR \SUBBYTES[9].a/U4540  ( .A(\w1[9][61] ), .B(n17273), .Z(
        \SUBBYTES[9].a/w1947 ) );
  XOR \SUBBYTES[9].a/U4539  ( .A(n16778), .B(n16777), .Z(\SUBBYTES[9].a/w1940 ) );
  XOR \SUBBYTES[9].a/U4538  ( .A(\w1[9][59] ), .B(\w1[9][57] ), .Z(n16777) );
  XOR \SUBBYTES[9].a/U4537  ( .A(\w1[9][63] ), .B(\w1[9][60] ), .Z(n16778) );
  XOR \SUBBYTES[9].a/U4536  ( .A(\w1[9][56] ), .B(\SUBBYTES[9].a/w1940 ), .Z(
        \SUBBYTES[9].a/w1819 ) );
  XOR \SUBBYTES[9].a/U4535  ( .A(n16780), .B(n16779), .Z(\SUBBYTES[9].a/w1927 ) );
  XOR \SUBBYTES[9].a/U4534  ( .A(\SUBBYTES[9].a/w1888 ), .B(n1093), .Z(n16779)
         );
  XOR \SUBBYTES[9].a/U4533  ( .A(\SUBBYTES[9].a/w1881 ), .B(
        \SUBBYTES[9].a/w1884 ), .Z(n16780) );
  XOR \SUBBYTES[9].a/U4532  ( .A(n16782), .B(n16781), .Z(\SUBBYTES[9].a/w1928 ) );
  XOR \SUBBYTES[9].a/U4531  ( .A(\SUBBYTES[9].a/w1888 ), .B(n16089), .Z(n16781) );
  XOR \SUBBYTES[9].a/U4530  ( .A(\SUBBYTES[9].a/w1881 ), .B(n16088), .Z(n16782) );
  XOR \SUBBYTES[9].a/U4529  ( .A(\SUBBYTES[9].a/w1940 ), .B(n16783), .Z(
        \SUBBYTES[9].a/w1930 ) );
  XOR \SUBBYTES[9].a/U4528  ( .A(\w1[9][62] ), .B(\w1[9][61] ), .Z(n16783) );
  XOR \SUBBYTES[9].a/U4527  ( .A(n16785), .B(n16784), .Z(\SUBBYTES[9].a/w1931 ) );
  XOR \SUBBYTES[9].a/U4526  ( .A(n16089), .B(n1093), .Z(n16784) );
  XOR \SUBBYTES[9].a/U4525  ( .A(n16088), .B(\SUBBYTES[9].a/w1884 ), .Z(n16785) );
  XOR \SUBBYTES[9].a/U4524  ( .A(\w1[9][63] ), .B(\w1[9][58] ), .Z(n17279) );
  XOR \SUBBYTES[9].a/U4523  ( .A(n17279), .B(n16786), .Z(\SUBBYTES[9].a/w1932 ) );
  XOR \SUBBYTES[9].a/U4522  ( .A(\w1[9][61] ), .B(\w1[9][60] ), .Z(n16786) );
  XOR \SUBBYTES[9].a/U4521  ( .A(\w1[9][63] ), .B(\SUBBYTES[9].a/w1817 ), .Z(
        \SUBBYTES[9].a/w1820 ) );
  XOR \SUBBYTES[9].a/U4520  ( .A(\w1[9][57] ), .B(\SUBBYTES[9].a/w1817 ), .Z(
        \SUBBYTES[9].a/w1821 ) );
  XOR \SUBBYTES[9].a/U4519  ( .A(\w1[9][60] ), .B(\SUBBYTES[9].a/w1817 ), .Z(
        \SUBBYTES[9].a/w1822 ) );
  XOR \SUBBYTES[9].a/U4518  ( .A(\SUBBYTES[9].a/w1821 ), .B(n17279), .Z(
        \SUBBYTES[9].a/w1823 ) );
  XOR \SUBBYTES[9].a/U4517  ( .A(n17279), .B(n16787), .Z(\SUBBYTES[9].a/w1908 ) );
  XOR \SUBBYTES[9].a/U4516  ( .A(\w1[9][60] ), .B(\w1[9][57] ), .Z(n16787) );
  XOR \SUBBYTES[9].a/U4515  ( .A(n16789), .B(n16788), .Z(n17276) );
  XOR \SUBBYTES[9].a/U4514  ( .A(\w1[9][60] ), .B(n16790), .Z(n16788) );
  XOR \SUBBYTES[9].a/U4513  ( .A(\SUBBYTES[9].a/w1873 ), .B(\w1[9][62] ), .Z(
        n16789) );
  XOR \SUBBYTES[9].a/U4512  ( .A(\SUBBYTES[9].a/w1847 ), .B(
        \SUBBYTES[9].a/w1854 ), .Z(n16790) );
  XOR \SUBBYTES[9].a/U4511  ( .A(n16792), .B(n16791), .Z(n17274) );
  XOR \SUBBYTES[9].a/U4510  ( .A(\w1[9][57] ), .B(n16793), .Z(n16791) );
  XOR \SUBBYTES[9].a/U4509  ( .A(\SUBBYTES[9].a/w1872 ), .B(\w1[9][61] ), .Z(
        n16792) );
  XOR \SUBBYTES[9].a/U4508  ( .A(\SUBBYTES[9].a/w1848 ), .B(
        \SUBBYTES[9].a/w1855 ), .Z(n16793) );
  XOR \SUBBYTES[9].a/U4507  ( .A(n17276), .B(n17274), .Z(\SUBBYTES[9].a/w1878 ) );
  XOR \SUBBYTES[9].a/U4506  ( .A(\w1[9][61] ), .B(n16794), .Z(n17277) );
  XOR \SUBBYTES[9].a/U4505  ( .A(\SUBBYTES[9].a/w1840 ), .B(
        \SUBBYTES[9].a/w1850 ), .Z(n16794) );
  XOR \SUBBYTES[9].a/U4504  ( .A(n16796), .B(n16795), .Z(\SUBBYTES[9].a/w1865 ) );
  XOR \SUBBYTES[9].a/U4503  ( .A(n17277), .B(n16797), .Z(n16795) );
  XOR \SUBBYTES[9].a/U4502  ( .A(\w1[9][60] ), .B(\SUBBYTES[9].a/w1929 ), .Z(
        n16796) );
  XOR \SUBBYTES[9].a/U4501  ( .A(\SUBBYTES[9].a/w1842 ), .B(
        \SUBBYTES[9].a/w1847 ), .Z(n16797) );
  XOR \SUBBYTES[9].a/U4500  ( .A(n16799), .B(n16798), .Z(n17275) );
  XOR \SUBBYTES[9].a/U4499  ( .A(\SUBBYTES[9].a/w1875 ), .B(\w1[9][63] ), .Z(
        n16798) );
  XOR \SUBBYTES[9].a/U4498  ( .A(\SUBBYTES[9].a/w1850 ), .B(
        \SUBBYTES[9].a/w1857 ), .Z(n16799) );
  XOR \SUBBYTES[9].a/U4497  ( .A(n17274), .B(n17275), .Z(\SUBBYTES[9].a/w1877 ) );
  XOR \SUBBYTES[9].a/U4496  ( .A(\w1[9][59] ), .B(n16800), .Z(n17278) );
  XOR \SUBBYTES[9].a/U4495  ( .A(\SUBBYTES[9].a/w1839 ), .B(
        \SUBBYTES[9].a/w1842 ), .Z(n16800) );
  XOR \SUBBYTES[9].a/U4494  ( .A(n16802), .B(n16801), .Z(\SUBBYTES[9].a/w1866 ) );
  XOR \SUBBYTES[9].a/U4493  ( .A(n17278), .B(n16803), .Z(n16801) );
  XOR \SUBBYTES[9].a/U4492  ( .A(\w1[9][62] ), .B(\SUBBYTES[9].a/w1908 ), .Z(
        n16802) );
  XOR \SUBBYTES[9].a/U4491  ( .A(\SUBBYTES[9].a/w1847 ), .B(
        \SUBBYTES[9].a/w1848 ), .Z(n16803) );
  XOR \SUBBYTES[9].a/U4490  ( .A(n17276), .B(n17275), .Z(\SUBBYTES[9].a/w1886 ) );
  XOR \SUBBYTES[9].a/U4489  ( .A(n16805), .B(n16804), .Z(\SUBBYTES[9].a/w1887 ) );
  XOR \SUBBYTES[9].a/U4488  ( .A(\w1[9][63] ), .B(n17277), .Z(n16804) );
  XOR \SUBBYTES[9].a/U4487  ( .A(\SUBBYTES[9].a/w1839 ), .B(
        \SUBBYTES[9].a/w1848 ), .Z(n16805) );
  XOR \SUBBYTES[9].a/U4486  ( .A(n16807), .B(n16806), .Z(\SUBBYTES[9].a/w1863 ) );
  XOR \SUBBYTES[9].a/U4485  ( .A(n16809), .B(n16808), .Z(n16806) );
  XOR \SUBBYTES[9].a/U4484  ( .A(\w1[9][63] ), .B(\SUBBYTES[9].a/w1947 ), .Z(
        n16807) );
  XOR \SUBBYTES[9].a/U4483  ( .A(\SUBBYTES[9].a/w1854 ), .B(
        \SUBBYTES[9].a/w1857 ), .Z(n16808) );
  XOR \SUBBYTES[9].a/U4482  ( .A(\SUBBYTES[9].a/w1840 ), .B(
        \SUBBYTES[9].a/w1842 ), .Z(n16809) );
  XOR \SUBBYTES[9].a/U4481  ( .A(n16811), .B(n16810), .Z(\SUBBYTES[9].a/w1864 ) );
  XOR \SUBBYTES[9].a/U4480  ( .A(n17278), .B(n16812), .Z(n16810) );
  XOR \SUBBYTES[9].a/U4479  ( .A(\w1[9][61] ), .B(n17279), .Z(n16811) );
  XOR \SUBBYTES[9].a/U4478  ( .A(\SUBBYTES[9].a/w1854 ), .B(
        \SUBBYTES[9].a/w1855 ), .Z(n16812) );
  XOR \SUBBYTES[9].a/U4477  ( .A(n16814), .B(n16813), .Z(\SUBBYTES[9].a/w1880 ) );
  XOR \SUBBYTES[9].a/U4476  ( .A(\w1[9][57] ), .B(n16815), .Z(n16813) );
  XOR \SUBBYTES[9].a/U4475  ( .A(\SUBBYTES[9].a/w1855 ), .B(
        \SUBBYTES[9].a/w1857 ), .Z(n16814) );
  XOR \SUBBYTES[9].a/U4474  ( .A(\SUBBYTES[9].a/w1839 ), .B(
        \SUBBYTES[9].a/w1840 ), .Z(n16815) );
  XOR \SUBBYTES[9].a/U4473  ( .A(\w1[9][65] ), .B(n16816), .Z(n17280) );
  XOR \SUBBYTES[9].a/U4472  ( .A(\w1[9][67] ), .B(\w1[9][66] ), .Z(n16816) );
  XOR \SUBBYTES[9].a/U4471  ( .A(\w1[9][70] ), .B(n17280), .Z(
        \SUBBYTES[9].a/w1722 ) );
  XOR \SUBBYTES[9].a/U4470  ( .A(\w1[9][64] ), .B(\SUBBYTES[9].a/w1722 ), .Z(
        \SUBBYTES[9].a/w1609 ) );
  XOR \SUBBYTES[9].a/U4469  ( .A(\w1[9][64] ), .B(n16817), .Z(
        \SUBBYTES[9].a/w1610 ) );
  XOR \SUBBYTES[9].a/U4468  ( .A(\w1[9][70] ), .B(\w1[9][69] ), .Z(n16817) );
  XOR \SUBBYTES[9].a/U4467  ( .A(\w1[9][69] ), .B(n17280), .Z(
        \SUBBYTES[9].a/w1740 ) );
  XOR \SUBBYTES[9].a/U4466  ( .A(n16819), .B(n16818), .Z(\SUBBYTES[9].a/w1733 ) );
  XOR \SUBBYTES[9].a/U4465  ( .A(\w1[9][67] ), .B(\w1[9][65] ), .Z(n16818) );
  XOR \SUBBYTES[9].a/U4464  ( .A(\w1[9][71] ), .B(\w1[9][68] ), .Z(n16819) );
  XOR \SUBBYTES[9].a/U4463  ( .A(\w1[9][64] ), .B(\SUBBYTES[9].a/w1733 ), .Z(
        \SUBBYTES[9].a/w1612 ) );
  XOR \SUBBYTES[9].a/U4462  ( .A(n16821), .B(n16820), .Z(\SUBBYTES[9].a/w1720 ) );
  XOR \SUBBYTES[9].a/U4461  ( .A(\SUBBYTES[9].a/w1681 ), .B(n1092), .Z(n16820)
         );
  XOR \SUBBYTES[9].a/U4460  ( .A(\SUBBYTES[9].a/w1674 ), .B(
        \SUBBYTES[9].a/w1677 ), .Z(n16821) );
  XOR \SUBBYTES[9].a/U4459  ( .A(n16823), .B(n16822), .Z(\SUBBYTES[9].a/w1721 ) );
  XOR \SUBBYTES[9].a/U4458  ( .A(\SUBBYTES[9].a/w1681 ), .B(n16087), .Z(n16822) );
  XOR \SUBBYTES[9].a/U4457  ( .A(\SUBBYTES[9].a/w1674 ), .B(n16086), .Z(n16823) );
  XOR \SUBBYTES[9].a/U4456  ( .A(\SUBBYTES[9].a/w1733 ), .B(n16824), .Z(
        \SUBBYTES[9].a/w1723 ) );
  XOR \SUBBYTES[9].a/U4455  ( .A(\w1[9][70] ), .B(\w1[9][69] ), .Z(n16824) );
  XOR \SUBBYTES[9].a/U4454  ( .A(n16826), .B(n16825), .Z(\SUBBYTES[9].a/w1724 ) );
  XOR \SUBBYTES[9].a/U4453  ( .A(n16087), .B(n1092), .Z(n16825) );
  XOR \SUBBYTES[9].a/U4452  ( .A(n16086), .B(\SUBBYTES[9].a/w1677 ), .Z(n16826) );
  XOR \SUBBYTES[9].a/U4451  ( .A(\w1[9][71] ), .B(\w1[9][66] ), .Z(n17286) );
  XOR \SUBBYTES[9].a/U4450  ( .A(n17286), .B(n16827), .Z(\SUBBYTES[9].a/w1725 ) );
  XOR \SUBBYTES[9].a/U4449  ( .A(\w1[9][69] ), .B(\w1[9][68] ), .Z(n16827) );
  XOR \SUBBYTES[9].a/U4448  ( .A(\w1[9][71] ), .B(\SUBBYTES[9].a/w1610 ), .Z(
        \SUBBYTES[9].a/w1613 ) );
  XOR \SUBBYTES[9].a/U4447  ( .A(\w1[9][65] ), .B(\SUBBYTES[9].a/w1610 ), .Z(
        \SUBBYTES[9].a/w1614 ) );
  XOR \SUBBYTES[9].a/U4446  ( .A(\w1[9][68] ), .B(\SUBBYTES[9].a/w1610 ), .Z(
        \SUBBYTES[9].a/w1615 ) );
  XOR \SUBBYTES[9].a/U4445  ( .A(\SUBBYTES[9].a/w1614 ), .B(n17286), .Z(
        \SUBBYTES[9].a/w1616 ) );
  XOR \SUBBYTES[9].a/U4444  ( .A(n17286), .B(n16828), .Z(\SUBBYTES[9].a/w1701 ) );
  XOR \SUBBYTES[9].a/U4443  ( .A(\w1[9][68] ), .B(\w1[9][65] ), .Z(n16828) );
  XOR \SUBBYTES[9].a/U4442  ( .A(n16830), .B(n16829), .Z(n17283) );
  XOR \SUBBYTES[9].a/U4441  ( .A(\w1[9][68] ), .B(n16831), .Z(n16829) );
  XOR \SUBBYTES[9].a/U4440  ( .A(\SUBBYTES[9].a/w1666 ), .B(\w1[9][70] ), .Z(
        n16830) );
  XOR \SUBBYTES[9].a/U4439  ( .A(\SUBBYTES[9].a/w1640 ), .B(
        \SUBBYTES[9].a/w1647 ), .Z(n16831) );
  XOR \SUBBYTES[9].a/U4438  ( .A(n16833), .B(n16832), .Z(n17281) );
  XOR \SUBBYTES[9].a/U4437  ( .A(\w1[9][65] ), .B(n16834), .Z(n16832) );
  XOR \SUBBYTES[9].a/U4436  ( .A(\SUBBYTES[9].a/w1665 ), .B(\w1[9][69] ), .Z(
        n16833) );
  XOR \SUBBYTES[9].a/U4435  ( .A(\SUBBYTES[9].a/w1641 ), .B(
        \SUBBYTES[9].a/w1648 ), .Z(n16834) );
  XOR \SUBBYTES[9].a/U4434  ( .A(n17283), .B(n17281), .Z(\SUBBYTES[9].a/w1671 ) );
  XOR \SUBBYTES[9].a/U4433  ( .A(\w1[9][69] ), .B(n16835), .Z(n17284) );
  XOR \SUBBYTES[9].a/U4432  ( .A(\SUBBYTES[9].a/w1633 ), .B(
        \SUBBYTES[9].a/w1643 ), .Z(n16835) );
  XOR \SUBBYTES[9].a/U4431  ( .A(n16837), .B(n16836), .Z(\SUBBYTES[9].a/w1658 ) );
  XOR \SUBBYTES[9].a/U4430  ( .A(n17284), .B(n16838), .Z(n16836) );
  XOR \SUBBYTES[9].a/U4429  ( .A(\w1[9][68] ), .B(\SUBBYTES[9].a/w1722 ), .Z(
        n16837) );
  XOR \SUBBYTES[9].a/U4428  ( .A(\SUBBYTES[9].a/w1635 ), .B(
        \SUBBYTES[9].a/w1640 ), .Z(n16838) );
  XOR \SUBBYTES[9].a/U4427  ( .A(n16840), .B(n16839), .Z(n17282) );
  XOR \SUBBYTES[9].a/U4426  ( .A(\SUBBYTES[9].a/w1668 ), .B(\w1[9][71] ), .Z(
        n16839) );
  XOR \SUBBYTES[9].a/U4425  ( .A(\SUBBYTES[9].a/w1643 ), .B(
        \SUBBYTES[9].a/w1650 ), .Z(n16840) );
  XOR \SUBBYTES[9].a/U4424  ( .A(n17281), .B(n17282), .Z(\SUBBYTES[9].a/w1670 ) );
  XOR \SUBBYTES[9].a/U4423  ( .A(\w1[9][67] ), .B(n16841), .Z(n17285) );
  XOR \SUBBYTES[9].a/U4422  ( .A(\SUBBYTES[9].a/w1632 ), .B(
        \SUBBYTES[9].a/w1635 ), .Z(n16841) );
  XOR \SUBBYTES[9].a/U4421  ( .A(n16843), .B(n16842), .Z(\SUBBYTES[9].a/w1659 ) );
  XOR \SUBBYTES[9].a/U4420  ( .A(n17285), .B(n16844), .Z(n16842) );
  XOR \SUBBYTES[9].a/U4419  ( .A(\w1[9][70] ), .B(\SUBBYTES[9].a/w1701 ), .Z(
        n16843) );
  XOR \SUBBYTES[9].a/U4418  ( .A(\SUBBYTES[9].a/w1640 ), .B(
        \SUBBYTES[9].a/w1641 ), .Z(n16844) );
  XOR \SUBBYTES[9].a/U4417  ( .A(n17283), .B(n17282), .Z(\SUBBYTES[9].a/w1679 ) );
  XOR \SUBBYTES[9].a/U4416  ( .A(n16846), .B(n16845), .Z(\SUBBYTES[9].a/w1680 ) );
  XOR \SUBBYTES[9].a/U4415  ( .A(\w1[9][71] ), .B(n17284), .Z(n16845) );
  XOR \SUBBYTES[9].a/U4414  ( .A(\SUBBYTES[9].a/w1632 ), .B(
        \SUBBYTES[9].a/w1641 ), .Z(n16846) );
  XOR \SUBBYTES[9].a/U4413  ( .A(n16848), .B(n16847), .Z(\SUBBYTES[9].a/w1656 ) );
  XOR \SUBBYTES[9].a/U4412  ( .A(n16850), .B(n16849), .Z(n16847) );
  XOR \SUBBYTES[9].a/U4411  ( .A(\w1[9][71] ), .B(\SUBBYTES[9].a/w1740 ), .Z(
        n16848) );
  XOR \SUBBYTES[9].a/U4410  ( .A(\SUBBYTES[9].a/w1647 ), .B(
        \SUBBYTES[9].a/w1650 ), .Z(n16849) );
  XOR \SUBBYTES[9].a/U4409  ( .A(\SUBBYTES[9].a/w1633 ), .B(
        \SUBBYTES[9].a/w1635 ), .Z(n16850) );
  XOR \SUBBYTES[9].a/U4408  ( .A(n16852), .B(n16851), .Z(\SUBBYTES[9].a/w1657 ) );
  XOR \SUBBYTES[9].a/U4407  ( .A(n17285), .B(n16853), .Z(n16851) );
  XOR \SUBBYTES[9].a/U4406  ( .A(\w1[9][69] ), .B(n17286), .Z(n16852) );
  XOR \SUBBYTES[9].a/U4405  ( .A(\SUBBYTES[9].a/w1647 ), .B(
        \SUBBYTES[9].a/w1648 ), .Z(n16853) );
  XOR \SUBBYTES[9].a/U4404  ( .A(n16855), .B(n16854), .Z(\SUBBYTES[9].a/w1673 ) );
  XOR \SUBBYTES[9].a/U4403  ( .A(\w1[9][65] ), .B(n16856), .Z(n16854) );
  XOR \SUBBYTES[9].a/U4402  ( .A(\SUBBYTES[9].a/w1648 ), .B(
        \SUBBYTES[9].a/w1650 ), .Z(n16855) );
  XOR \SUBBYTES[9].a/U4401  ( .A(\SUBBYTES[9].a/w1632 ), .B(
        \SUBBYTES[9].a/w1633 ), .Z(n16856) );
  XOR \SUBBYTES[9].a/U4400  ( .A(\w1[9][73] ), .B(n16857), .Z(n17287) );
  XOR \SUBBYTES[9].a/U4399  ( .A(\w1[9][75] ), .B(\w1[9][74] ), .Z(n16857) );
  XOR \SUBBYTES[9].a/U4398  ( .A(\w1[9][78] ), .B(n17287), .Z(
        \SUBBYTES[9].a/w1515 ) );
  XOR \SUBBYTES[9].a/U4397  ( .A(\w1[9][72] ), .B(\SUBBYTES[9].a/w1515 ), .Z(
        \SUBBYTES[9].a/w1402 ) );
  XOR \SUBBYTES[9].a/U4396  ( .A(\w1[9][72] ), .B(n16858), .Z(
        \SUBBYTES[9].a/w1403 ) );
  XOR \SUBBYTES[9].a/U4395  ( .A(\w1[9][78] ), .B(\w1[9][77] ), .Z(n16858) );
  XOR \SUBBYTES[9].a/U4394  ( .A(\w1[9][77] ), .B(n17287), .Z(
        \SUBBYTES[9].a/w1533 ) );
  XOR \SUBBYTES[9].a/U4393  ( .A(n16860), .B(n16859), .Z(\SUBBYTES[9].a/w1526 ) );
  XOR \SUBBYTES[9].a/U4392  ( .A(\w1[9][75] ), .B(\w1[9][73] ), .Z(n16859) );
  XOR \SUBBYTES[9].a/U4391  ( .A(\w1[9][79] ), .B(\w1[9][76] ), .Z(n16860) );
  XOR \SUBBYTES[9].a/U4390  ( .A(\w1[9][72] ), .B(\SUBBYTES[9].a/w1526 ), .Z(
        \SUBBYTES[9].a/w1405 ) );
  XOR \SUBBYTES[9].a/U4389  ( .A(n16862), .B(n16861), .Z(\SUBBYTES[9].a/w1513 ) );
  XOR \SUBBYTES[9].a/U4388  ( .A(\SUBBYTES[9].a/w1474 ), .B(n1091), .Z(n16861)
         );
  XOR \SUBBYTES[9].a/U4387  ( .A(\SUBBYTES[9].a/w1467 ), .B(
        \SUBBYTES[9].a/w1470 ), .Z(n16862) );
  XOR \SUBBYTES[9].a/U4386  ( .A(n16864), .B(n16863), .Z(\SUBBYTES[9].a/w1514 ) );
  XOR \SUBBYTES[9].a/U4385  ( .A(\SUBBYTES[9].a/w1474 ), .B(n16085), .Z(n16863) );
  XOR \SUBBYTES[9].a/U4384  ( .A(\SUBBYTES[9].a/w1467 ), .B(n16084), .Z(n16864) );
  XOR \SUBBYTES[9].a/U4383  ( .A(\SUBBYTES[9].a/w1526 ), .B(n16865), .Z(
        \SUBBYTES[9].a/w1516 ) );
  XOR \SUBBYTES[9].a/U4382  ( .A(\w1[9][78] ), .B(\w1[9][77] ), .Z(n16865) );
  XOR \SUBBYTES[9].a/U4381  ( .A(n16867), .B(n16866), .Z(\SUBBYTES[9].a/w1517 ) );
  XOR \SUBBYTES[9].a/U4380  ( .A(n16085), .B(n1091), .Z(n16866) );
  XOR \SUBBYTES[9].a/U4379  ( .A(n16084), .B(\SUBBYTES[9].a/w1470 ), .Z(n16867) );
  XOR \SUBBYTES[9].a/U4378  ( .A(\w1[9][79] ), .B(\w1[9][74] ), .Z(n17293) );
  XOR \SUBBYTES[9].a/U4377  ( .A(n17293), .B(n16868), .Z(\SUBBYTES[9].a/w1518 ) );
  XOR \SUBBYTES[9].a/U4376  ( .A(\w1[9][77] ), .B(\w1[9][76] ), .Z(n16868) );
  XOR \SUBBYTES[9].a/U4375  ( .A(\w1[9][79] ), .B(\SUBBYTES[9].a/w1403 ), .Z(
        \SUBBYTES[9].a/w1406 ) );
  XOR \SUBBYTES[9].a/U4374  ( .A(\w1[9][73] ), .B(\SUBBYTES[9].a/w1403 ), .Z(
        \SUBBYTES[9].a/w1407 ) );
  XOR \SUBBYTES[9].a/U4373  ( .A(\w1[9][76] ), .B(\SUBBYTES[9].a/w1403 ), .Z(
        \SUBBYTES[9].a/w1408 ) );
  XOR \SUBBYTES[9].a/U4372  ( .A(\SUBBYTES[9].a/w1407 ), .B(n17293), .Z(
        \SUBBYTES[9].a/w1409 ) );
  XOR \SUBBYTES[9].a/U4371  ( .A(n17293), .B(n16869), .Z(\SUBBYTES[9].a/w1494 ) );
  XOR \SUBBYTES[9].a/U4370  ( .A(\w1[9][76] ), .B(\w1[9][73] ), .Z(n16869) );
  XOR \SUBBYTES[9].a/U4369  ( .A(n16871), .B(n16870), .Z(n17290) );
  XOR \SUBBYTES[9].a/U4368  ( .A(\w1[9][76] ), .B(n16872), .Z(n16870) );
  XOR \SUBBYTES[9].a/U4367  ( .A(\SUBBYTES[9].a/w1459 ), .B(\w1[9][78] ), .Z(
        n16871) );
  XOR \SUBBYTES[9].a/U4366  ( .A(\SUBBYTES[9].a/w1433 ), .B(
        \SUBBYTES[9].a/w1440 ), .Z(n16872) );
  XOR \SUBBYTES[9].a/U4365  ( .A(n16874), .B(n16873), .Z(n17288) );
  XOR \SUBBYTES[9].a/U4364  ( .A(\w1[9][73] ), .B(n16875), .Z(n16873) );
  XOR \SUBBYTES[9].a/U4363  ( .A(\SUBBYTES[9].a/w1458 ), .B(\w1[9][77] ), .Z(
        n16874) );
  XOR \SUBBYTES[9].a/U4362  ( .A(\SUBBYTES[9].a/w1434 ), .B(
        \SUBBYTES[9].a/w1441 ), .Z(n16875) );
  XOR \SUBBYTES[9].a/U4361  ( .A(n17290), .B(n17288), .Z(\SUBBYTES[9].a/w1464 ) );
  XOR \SUBBYTES[9].a/U4360  ( .A(\w1[9][77] ), .B(n16876), .Z(n17291) );
  XOR \SUBBYTES[9].a/U4359  ( .A(\SUBBYTES[9].a/w1426 ), .B(
        \SUBBYTES[9].a/w1436 ), .Z(n16876) );
  XOR \SUBBYTES[9].a/U4358  ( .A(n16878), .B(n16877), .Z(\SUBBYTES[9].a/w1451 ) );
  XOR \SUBBYTES[9].a/U4357  ( .A(n17291), .B(n16879), .Z(n16877) );
  XOR \SUBBYTES[9].a/U4356  ( .A(\w1[9][76] ), .B(\SUBBYTES[9].a/w1515 ), .Z(
        n16878) );
  XOR \SUBBYTES[9].a/U4355  ( .A(\SUBBYTES[9].a/w1428 ), .B(
        \SUBBYTES[9].a/w1433 ), .Z(n16879) );
  XOR \SUBBYTES[9].a/U4354  ( .A(n16881), .B(n16880), .Z(n17289) );
  XOR \SUBBYTES[9].a/U4353  ( .A(\SUBBYTES[9].a/w1461 ), .B(\w1[9][79] ), .Z(
        n16880) );
  XOR \SUBBYTES[9].a/U4352  ( .A(\SUBBYTES[9].a/w1436 ), .B(
        \SUBBYTES[9].a/w1443 ), .Z(n16881) );
  XOR \SUBBYTES[9].a/U4351  ( .A(n17288), .B(n17289), .Z(\SUBBYTES[9].a/w1463 ) );
  XOR \SUBBYTES[9].a/U4350  ( .A(\w1[9][75] ), .B(n16882), .Z(n17292) );
  XOR \SUBBYTES[9].a/U4349  ( .A(\SUBBYTES[9].a/w1425 ), .B(
        \SUBBYTES[9].a/w1428 ), .Z(n16882) );
  XOR \SUBBYTES[9].a/U4348  ( .A(n16884), .B(n16883), .Z(\SUBBYTES[9].a/w1452 ) );
  XOR \SUBBYTES[9].a/U4347  ( .A(n17292), .B(n16885), .Z(n16883) );
  XOR \SUBBYTES[9].a/U4346  ( .A(\w1[9][78] ), .B(\SUBBYTES[9].a/w1494 ), .Z(
        n16884) );
  XOR \SUBBYTES[9].a/U4345  ( .A(\SUBBYTES[9].a/w1433 ), .B(
        \SUBBYTES[9].a/w1434 ), .Z(n16885) );
  XOR \SUBBYTES[9].a/U4344  ( .A(n17290), .B(n17289), .Z(\SUBBYTES[9].a/w1472 ) );
  XOR \SUBBYTES[9].a/U4343  ( .A(n16887), .B(n16886), .Z(\SUBBYTES[9].a/w1473 ) );
  XOR \SUBBYTES[9].a/U4342  ( .A(\w1[9][79] ), .B(n17291), .Z(n16886) );
  XOR \SUBBYTES[9].a/U4341  ( .A(\SUBBYTES[9].a/w1425 ), .B(
        \SUBBYTES[9].a/w1434 ), .Z(n16887) );
  XOR \SUBBYTES[9].a/U4340  ( .A(n16889), .B(n16888), .Z(\SUBBYTES[9].a/w1449 ) );
  XOR \SUBBYTES[9].a/U4339  ( .A(n16891), .B(n16890), .Z(n16888) );
  XOR \SUBBYTES[9].a/U4338  ( .A(\w1[9][79] ), .B(\SUBBYTES[9].a/w1533 ), .Z(
        n16889) );
  XOR \SUBBYTES[9].a/U4337  ( .A(\SUBBYTES[9].a/w1440 ), .B(
        \SUBBYTES[9].a/w1443 ), .Z(n16890) );
  XOR \SUBBYTES[9].a/U4336  ( .A(\SUBBYTES[9].a/w1426 ), .B(
        \SUBBYTES[9].a/w1428 ), .Z(n16891) );
  XOR \SUBBYTES[9].a/U4335  ( .A(n16893), .B(n16892), .Z(\SUBBYTES[9].a/w1450 ) );
  XOR \SUBBYTES[9].a/U4334  ( .A(n17292), .B(n16894), .Z(n16892) );
  XOR \SUBBYTES[9].a/U4333  ( .A(\w1[9][77] ), .B(n17293), .Z(n16893) );
  XOR \SUBBYTES[9].a/U4332  ( .A(\SUBBYTES[9].a/w1440 ), .B(
        \SUBBYTES[9].a/w1441 ), .Z(n16894) );
  XOR \SUBBYTES[9].a/U4331  ( .A(n16896), .B(n16895), .Z(\SUBBYTES[9].a/w1466 ) );
  XOR \SUBBYTES[9].a/U4330  ( .A(\w1[9][73] ), .B(n16897), .Z(n16895) );
  XOR \SUBBYTES[9].a/U4329  ( .A(\SUBBYTES[9].a/w1441 ), .B(
        \SUBBYTES[9].a/w1443 ), .Z(n16896) );
  XOR \SUBBYTES[9].a/U4328  ( .A(\SUBBYTES[9].a/w1425 ), .B(
        \SUBBYTES[9].a/w1426 ), .Z(n16897) );
  XOR \SUBBYTES[9].a/U4327  ( .A(\w1[9][81] ), .B(n16898), .Z(n17294) );
  XOR \SUBBYTES[9].a/U4326  ( .A(\w1[9][83] ), .B(\w1[9][82] ), .Z(n16898) );
  XOR \SUBBYTES[9].a/U4325  ( .A(\w1[9][86] ), .B(n17294), .Z(
        \SUBBYTES[9].a/w1308 ) );
  XOR \SUBBYTES[9].a/U4324  ( .A(\w1[9][80] ), .B(\SUBBYTES[9].a/w1308 ), .Z(
        \SUBBYTES[9].a/w1195 ) );
  XOR \SUBBYTES[9].a/U4323  ( .A(\w1[9][80] ), .B(n16899), .Z(
        \SUBBYTES[9].a/w1196 ) );
  XOR \SUBBYTES[9].a/U4322  ( .A(\w1[9][86] ), .B(\w1[9][85] ), .Z(n16899) );
  XOR \SUBBYTES[9].a/U4321  ( .A(\w1[9][85] ), .B(n17294), .Z(
        \SUBBYTES[9].a/w1326 ) );
  XOR \SUBBYTES[9].a/U4320  ( .A(n16901), .B(n16900), .Z(\SUBBYTES[9].a/w1319 ) );
  XOR \SUBBYTES[9].a/U4319  ( .A(\w1[9][83] ), .B(\w1[9][81] ), .Z(n16900) );
  XOR \SUBBYTES[9].a/U4318  ( .A(\w1[9][87] ), .B(\w1[9][84] ), .Z(n16901) );
  XOR \SUBBYTES[9].a/U4317  ( .A(\w1[9][80] ), .B(\SUBBYTES[9].a/w1319 ), .Z(
        \SUBBYTES[9].a/w1198 ) );
  XOR \SUBBYTES[9].a/U4316  ( .A(n16903), .B(n16902), .Z(\SUBBYTES[9].a/w1306 ) );
  XOR \SUBBYTES[9].a/U4315  ( .A(\SUBBYTES[9].a/w1267 ), .B(n1090), .Z(n16902)
         );
  XOR \SUBBYTES[9].a/U4314  ( .A(\SUBBYTES[9].a/w1260 ), .B(
        \SUBBYTES[9].a/w1263 ), .Z(n16903) );
  XOR \SUBBYTES[9].a/U4313  ( .A(n16905), .B(n16904), .Z(\SUBBYTES[9].a/w1307 ) );
  XOR \SUBBYTES[9].a/U4312  ( .A(\SUBBYTES[9].a/w1267 ), .B(n16083), .Z(n16904) );
  XOR \SUBBYTES[9].a/U4311  ( .A(\SUBBYTES[9].a/w1260 ), .B(n16082), .Z(n16905) );
  XOR \SUBBYTES[9].a/U4310  ( .A(\SUBBYTES[9].a/w1319 ), .B(n16906), .Z(
        \SUBBYTES[9].a/w1309 ) );
  XOR \SUBBYTES[9].a/U4309  ( .A(\w1[9][86] ), .B(\w1[9][85] ), .Z(n16906) );
  XOR \SUBBYTES[9].a/U4308  ( .A(n16908), .B(n16907), .Z(\SUBBYTES[9].a/w1310 ) );
  XOR \SUBBYTES[9].a/U4307  ( .A(n16083), .B(n1090), .Z(n16907) );
  XOR \SUBBYTES[9].a/U4306  ( .A(n16082), .B(\SUBBYTES[9].a/w1263 ), .Z(n16908) );
  XOR \SUBBYTES[9].a/U4305  ( .A(\w1[9][87] ), .B(\w1[9][82] ), .Z(n17300) );
  XOR \SUBBYTES[9].a/U4304  ( .A(n17300), .B(n16909), .Z(\SUBBYTES[9].a/w1311 ) );
  XOR \SUBBYTES[9].a/U4303  ( .A(\w1[9][85] ), .B(\w1[9][84] ), .Z(n16909) );
  XOR \SUBBYTES[9].a/U4302  ( .A(\w1[9][87] ), .B(\SUBBYTES[9].a/w1196 ), .Z(
        \SUBBYTES[9].a/w1199 ) );
  XOR \SUBBYTES[9].a/U4301  ( .A(\w1[9][81] ), .B(\SUBBYTES[9].a/w1196 ), .Z(
        \SUBBYTES[9].a/w1200 ) );
  XOR \SUBBYTES[9].a/U4300  ( .A(\w1[9][84] ), .B(\SUBBYTES[9].a/w1196 ), .Z(
        \SUBBYTES[9].a/w1201 ) );
  XOR \SUBBYTES[9].a/U4299  ( .A(\SUBBYTES[9].a/w1200 ), .B(n17300), .Z(
        \SUBBYTES[9].a/w1202 ) );
  XOR \SUBBYTES[9].a/U4298  ( .A(n17300), .B(n16910), .Z(\SUBBYTES[9].a/w1287 ) );
  XOR \SUBBYTES[9].a/U4297  ( .A(\w1[9][84] ), .B(\w1[9][81] ), .Z(n16910) );
  XOR \SUBBYTES[9].a/U4296  ( .A(n16912), .B(n16911), .Z(n17297) );
  XOR \SUBBYTES[9].a/U4295  ( .A(\w1[9][84] ), .B(n16913), .Z(n16911) );
  XOR \SUBBYTES[9].a/U4294  ( .A(\SUBBYTES[9].a/w1252 ), .B(\w1[9][86] ), .Z(
        n16912) );
  XOR \SUBBYTES[9].a/U4293  ( .A(\SUBBYTES[9].a/w1226 ), .B(
        \SUBBYTES[9].a/w1233 ), .Z(n16913) );
  XOR \SUBBYTES[9].a/U4292  ( .A(n16915), .B(n16914), .Z(n17295) );
  XOR \SUBBYTES[9].a/U4291  ( .A(\w1[9][81] ), .B(n16916), .Z(n16914) );
  XOR \SUBBYTES[9].a/U4290  ( .A(\SUBBYTES[9].a/w1251 ), .B(\w1[9][85] ), .Z(
        n16915) );
  XOR \SUBBYTES[9].a/U4289  ( .A(\SUBBYTES[9].a/w1227 ), .B(
        \SUBBYTES[9].a/w1234 ), .Z(n16916) );
  XOR \SUBBYTES[9].a/U4288  ( .A(n17297), .B(n17295), .Z(\SUBBYTES[9].a/w1257 ) );
  XOR \SUBBYTES[9].a/U4287  ( .A(\w1[9][85] ), .B(n16917), .Z(n17298) );
  XOR \SUBBYTES[9].a/U4286  ( .A(\SUBBYTES[9].a/w1219 ), .B(
        \SUBBYTES[9].a/w1229 ), .Z(n16917) );
  XOR \SUBBYTES[9].a/U4285  ( .A(n16919), .B(n16918), .Z(\SUBBYTES[9].a/w1244 ) );
  XOR \SUBBYTES[9].a/U4284  ( .A(n17298), .B(n16920), .Z(n16918) );
  XOR \SUBBYTES[9].a/U4283  ( .A(\w1[9][84] ), .B(\SUBBYTES[9].a/w1308 ), .Z(
        n16919) );
  XOR \SUBBYTES[9].a/U4282  ( .A(\SUBBYTES[9].a/w1221 ), .B(
        \SUBBYTES[9].a/w1226 ), .Z(n16920) );
  XOR \SUBBYTES[9].a/U4281  ( .A(n16922), .B(n16921), .Z(n17296) );
  XOR \SUBBYTES[9].a/U4280  ( .A(\SUBBYTES[9].a/w1254 ), .B(\w1[9][87] ), .Z(
        n16921) );
  XOR \SUBBYTES[9].a/U4279  ( .A(\SUBBYTES[9].a/w1229 ), .B(
        \SUBBYTES[9].a/w1236 ), .Z(n16922) );
  XOR \SUBBYTES[9].a/U4278  ( .A(n17295), .B(n17296), .Z(\SUBBYTES[9].a/w1256 ) );
  XOR \SUBBYTES[9].a/U4277  ( .A(\w1[9][83] ), .B(n16923), .Z(n17299) );
  XOR \SUBBYTES[9].a/U4276  ( .A(\SUBBYTES[9].a/w1218 ), .B(
        \SUBBYTES[9].a/w1221 ), .Z(n16923) );
  XOR \SUBBYTES[9].a/U4275  ( .A(n16925), .B(n16924), .Z(\SUBBYTES[9].a/w1245 ) );
  XOR \SUBBYTES[9].a/U4274  ( .A(n17299), .B(n16926), .Z(n16924) );
  XOR \SUBBYTES[9].a/U4273  ( .A(\w1[9][86] ), .B(\SUBBYTES[9].a/w1287 ), .Z(
        n16925) );
  XOR \SUBBYTES[9].a/U4272  ( .A(\SUBBYTES[9].a/w1226 ), .B(
        \SUBBYTES[9].a/w1227 ), .Z(n16926) );
  XOR \SUBBYTES[9].a/U4271  ( .A(n17297), .B(n17296), .Z(\SUBBYTES[9].a/w1265 ) );
  XOR \SUBBYTES[9].a/U4270  ( .A(n16928), .B(n16927), .Z(\SUBBYTES[9].a/w1266 ) );
  XOR \SUBBYTES[9].a/U4269  ( .A(\w1[9][87] ), .B(n17298), .Z(n16927) );
  XOR \SUBBYTES[9].a/U4268  ( .A(\SUBBYTES[9].a/w1218 ), .B(
        \SUBBYTES[9].a/w1227 ), .Z(n16928) );
  XOR \SUBBYTES[9].a/U4267  ( .A(n16930), .B(n16929), .Z(\SUBBYTES[9].a/w1242 ) );
  XOR \SUBBYTES[9].a/U4266  ( .A(n16932), .B(n16931), .Z(n16929) );
  XOR \SUBBYTES[9].a/U4265  ( .A(\w1[9][87] ), .B(\SUBBYTES[9].a/w1326 ), .Z(
        n16930) );
  XOR \SUBBYTES[9].a/U4264  ( .A(\SUBBYTES[9].a/w1233 ), .B(
        \SUBBYTES[9].a/w1236 ), .Z(n16931) );
  XOR \SUBBYTES[9].a/U4263  ( .A(\SUBBYTES[9].a/w1219 ), .B(
        \SUBBYTES[9].a/w1221 ), .Z(n16932) );
  XOR \SUBBYTES[9].a/U4262  ( .A(n16934), .B(n16933), .Z(\SUBBYTES[9].a/w1243 ) );
  XOR \SUBBYTES[9].a/U4261  ( .A(n17299), .B(n16935), .Z(n16933) );
  XOR \SUBBYTES[9].a/U4260  ( .A(\w1[9][85] ), .B(n17300), .Z(n16934) );
  XOR \SUBBYTES[9].a/U4259  ( .A(\SUBBYTES[9].a/w1233 ), .B(
        \SUBBYTES[9].a/w1234 ), .Z(n16935) );
  XOR \SUBBYTES[9].a/U4258  ( .A(n16937), .B(n16936), .Z(\SUBBYTES[9].a/w1259 ) );
  XOR \SUBBYTES[9].a/U4257  ( .A(\w1[9][81] ), .B(n16938), .Z(n16936) );
  XOR \SUBBYTES[9].a/U4256  ( .A(\SUBBYTES[9].a/w1234 ), .B(
        \SUBBYTES[9].a/w1236 ), .Z(n16937) );
  XOR \SUBBYTES[9].a/U4255  ( .A(\SUBBYTES[9].a/w1218 ), .B(
        \SUBBYTES[9].a/w1219 ), .Z(n16938) );
  XOR \SUBBYTES[9].a/U4254  ( .A(\w1[9][89] ), .B(n16939), .Z(n17301) );
  XOR \SUBBYTES[9].a/U4253  ( .A(\w1[9][91] ), .B(\w1[9][90] ), .Z(n16939) );
  XOR \SUBBYTES[9].a/U4252  ( .A(\w1[9][94] ), .B(n17301), .Z(
        \SUBBYTES[9].a/w1101 ) );
  XOR \SUBBYTES[9].a/U4251  ( .A(\w1[9][88] ), .B(\SUBBYTES[9].a/w1101 ), .Z(
        \SUBBYTES[9].a/w988 ) );
  XOR \SUBBYTES[9].a/U4250  ( .A(\w1[9][88] ), .B(n16940), .Z(
        \SUBBYTES[9].a/w989 ) );
  XOR \SUBBYTES[9].a/U4249  ( .A(\w1[9][94] ), .B(\w1[9][93] ), .Z(n16940) );
  XOR \SUBBYTES[9].a/U4248  ( .A(\w1[9][93] ), .B(n17301), .Z(
        \SUBBYTES[9].a/w1119 ) );
  XOR \SUBBYTES[9].a/U4247  ( .A(n16942), .B(n16941), .Z(\SUBBYTES[9].a/w1112 ) );
  XOR \SUBBYTES[9].a/U4246  ( .A(\w1[9][91] ), .B(\w1[9][89] ), .Z(n16941) );
  XOR \SUBBYTES[9].a/U4245  ( .A(\w1[9][95] ), .B(\w1[9][92] ), .Z(n16942) );
  XOR \SUBBYTES[9].a/U4244  ( .A(\w1[9][88] ), .B(\SUBBYTES[9].a/w1112 ), .Z(
        \SUBBYTES[9].a/w991 ) );
  XOR \SUBBYTES[9].a/U4243  ( .A(n16944), .B(n16943), .Z(\SUBBYTES[9].a/w1099 ) );
  XOR \SUBBYTES[9].a/U4242  ( .A(\SUBBYTES[9].a/w1060 ), .B(n1089), .Z(n16943)
         );
  XOR \SUBBYTES[9].a/U4241  ( .A(\SUBBYTES[9].a/w1053 ), .B(
        \SUBBYTES[9].a/w1056 ), .Z(n16944) );
  XOR \SUBBYTES[9].a/U4240  ( .A(n16946), .B(n16945), .Z(\SUBBYTES[9].a/w1100 ) );
  XOR \SUBBYTES[9].a/U4239  ( .A(\SUBBYTES[9].a/w1060 ), .B(n16081), .Z(n16945) );
  XOR \SUBBYTES[9].a/U4238  ( .A(\SUBBYTES[9].a/w1053 ), .B(n16080), .Z(n16946) );
  XOR \SUBBYTES[9].a/U4237  ( .A(\SUBBYTES[9].a/w1112 ), .B(n16947), .Z(
        \SUBBYTES[9].a/w1102 ) );
  XOR \SUBBYTES[9].a/U4236  ( .A(\w1[9][94] ), .B(\w1[9][93] ), .Z(n16947) );
  XOR \SUBBYTES[9].a/U4235  ( .A(n16949), .B(n16948), .Z(\SUBBYTES[9].a/w1103 ) );
  XOR \SUBBYTES[9].a/U4234  ( .A(n16081), .B(n1089), .Z(n16948) );
  XOR \SUBBYTES[9].a/U4233  ( .A(n16080), .B(\SUBBYTES[9].a/w1056 ), .Z(n16949) );
  XOR \SUBBYTES[9].a/U4232  ( .A(\w1[9][95] ), .B(\w1[9][90] ), .Z(n17307) );
  XOR \SUBBYTES[9].a/U4231  ( .A(n17307), .B(n16950), .Z(\SUBBYTES[9].a/w1104 ) );
  XOR \SUBBYTES[9].a/U4230  ( .A(\w1[9][93] ), .B(\w1[9][92] ), .Z(n16950) );
  XOR \SUBBYTES[9].a/U4229  ( .A(\w1[9][95] ), .B(\SUBBYTES[9].a/w989 ), .Z(
        \SUBBYTES[9].a/w992 ) );
  XOR \SUBBYTES[9].a/U4228  ( .A(\w1[9][89] ), .B(\SUBBYTES[9].a/w989 ), .Z(
        \SUBBYTES[9].a/w993 ) );
  XOR \SUBBYTES[9].a/U4227  ( .A(\w1[9][92] ), .B(\SUBBYTES[9].a/w989 ), .Z(
        \SUBBYTES[9].a/w994 ) );
  XOR \SUBBYTES[9].a/U4226  ( .A(\SUBBYTES[9].a/w993 ), .B(n17307), .Z(
        \SUBBYTES[9].a/w995 ) );
  XOR \SUBBYTES[9].a/U4225  ( .A(n17307), .B(n16951), .Z(\SUBBYTES[9].a/w1080 ) );
  XOR \SUBBYTES[9].a/U4224  ( .A(\w1[9][92] ), .B(\w1[9][89] ), .Z(n16951) );
  XOR \SUBBYTES[9].a/U4223  ( .A(n16953), .B(n16952), .Z(n17304) );
  XOR \SUBBYTES[9].a/U4222  ( .A(\w1[9][92] ), .B(n16954), .Z(n16952) );
  XOR \SUBBYTES[9].a/U4221  ( .A(\SUBBYTES[9].a/w1045 ), .B(\w1[9][94] ), .Z(
        n16953) );
  XOR \SUBBYTES[9].a/U4220  ( .A(\SUBBYTES[9].a/w1019 ), .B(
        \SUBBYTES[9].a/w1026 ), .Z(n16954) );
  XOR \SUBBYTES[9].a/U4219  ( .A(n16956), .B(n16955), .Z(n17302) );
  XOR \SUBBYTES[9].a/U4218  ( .A(\w1[9][89] ), .B(n16957), .Z(n16955) );
  XOR \SUBBYTES[9].a/U4217  ( .A(\SUBBYTES[9].a/w1044 ), .B(\w1[9][93] ), .Z(
        n16956) );
  XOR \SUBBYTES[9].a/U4216  ( .A(\SUBBYTES[9].a/w1020 ), .B(
        \SUBBYTES[9].a/w1027 ), .Z(n16957) );
  XOR \SUBBYTES[9].a/U4215  ( .A(n17304), .B(n17302), .Z(\SUBBYTES[9].a/w1050 ) );
  XOR \SUBBYTES[9].a/U4214  ( .A(\w1[9][93] ), .B(n16958), .Z(n17305) );
  XOR \SUBBYTES[9].a/U4213  ( .A(\SUBBYTES[9].a/w1012 ), .B(
        \SUBBYTES[9].a/w1022 ), .Z(n16958) );
  XOR \SUBBYTES[9].a/U4212  ( .A(n16960), .B(n16959), .Z(\SUBBYTES[9].a/w1037 ) );
  XOR \SUBBYTES[9].a/U4211  ( .A(n17305), .B(n16961), .Z(n16959) );
  XOR \SUBBYTES[9].a/U4210  ( .A(\w1[9][92] ), .B(\SUBBYTES[9].a/w1101 ), .Z(
        n16960) );
  XOR \SUBBYTES[9].a/U4209  ( .A(\SUBBYTES[9].a/w1014 ), .B(
        \SUBBYTES[9].a/w1019 ), .Z(n16961) );
  XOR \SUBBYTES[9].a/U4208  ( .A(n16963), .B(n16962), .Z(n17303) );
  XOR \SUBBYTES[9].a/U4207  ( .A(\SUBBYTES[9].a/w1047 ), .B(\w1[9][95] ), .Z(
        n16962) );
  XOR \SUBBYTES[9].a/U4206  ( .A(\SUBBYTES[9].a/w1022 ), .B(
        \SUBBYTES[9].a/w1029 ), .Z(n16963) );
  XOR \SUBBYTES[9].a/U4205  ( .A(n17302), .B(n17303), .Z(\SUBBYTES[9].a/w1049 ) );
  XOR \SUBBYTES[9].a/U4204  ( .A(\w1[9][91] ), .B(n16964), .Z(n17306) );
  XOR \SUBBYTES[9].a/U4203  ( .A(\SUBBYTES[9].a/w1011 ), .B(
        \SUBBYTES[9].a/w1014 ), .Z(n16964) );
  XOR \SUBBYTES[9].a/U4202  ( .A(n16966), .B(n16965), .Z(\SUBBYTES[9].a/w1038 ) );
  XOR \SUBBYTES[9].a/U4201  ( .A(n17306), .B(n16967), .Z(n16965) );
  XOR \SUBBYTES[9].a/U4200  ( .A(\w1[9][94] ), .B(\SUBBYTES[9].a/w1080 ), .Z(
        n16966) );
  XOR \SUBBYTES[9].a/U4199  ( .A(\SUBBYTES[9].a/w1019 ), .B(
        \SUBBYTES[9].a/w1020 ), .Z(n16967) );
  XOR \SUBBYTES[9].a/U4198  ( .A(n17304), .B(n17303), .Z(\SUBBYTES[9].a/w1058 ) );
  XOR \SUBBYTES[9].a/U4197  ( .A(n16969), .B(n16968), .Z(\SUBBYTES[9].a/w1059 ) );
  XOR \SUBBYTES[9].a/U4196  ( .A(\w1[9][95] ), .B(n17305), .Z(n16968) );
  XOR \SUBBYTES[9].a/U4195  ( .A(\SUBBYTES[9].a/w1011 ), .B(
        \SUBBYTES[9].a/w1020 ), .Z(n16969) );
  XOR \SUBBYTES[9].a/U4194  ( .A(n16971), .B(n16970), .Z(\SUBBYTES[9].a/w1035 ) );
  XOR \SUBBYTES[9].a/U4193  ( .A(n16973), .B(n16972), .Z(n16970) );
  XOR \SUBBYTES[9].a/U4192  ( .A(\w1[9][95] ), .B(\SUBBYTES[9].a/w1119 ), .Z(
        n16971) );
  XOR \SUBBYTES[9].a/U4191  ( .A(\SUBBYTES[9].a/w1026 ), .B(
        \SUBBYTES[9].a/w1029 ), .Z(n16972) );
  XOR \SUBBYTES[9].a/U4190  ( .A(\SUBBYTES[9].a/w1012 ), .B(
        \SUBBYTES[9].a/w1014 ), .Z(n16973) );
  XOR \SUBBYTES[9].a/U4189  ( .A(n16975), .B(n16974), .Z(\SUBBYTES[9].a/w1036 ) );
  XOR \SUBBYTES[9].a/U4188  ( .A(n17306), .B(n16976), .Z(n16974) );
  XOR \SUBBYTES[9].a/U4187  ( .A(\w1[9][93] ), .B(n17307), .Z(n16975) );
  XOR \SUBBYTES[9].a/U4186  ( .A(\SUBBYTES[9].a/w1026 ), .B(
        \SUBBYTES[9].a/w1027 ), .Z(n16976) );
  XOR \SUBBYTES[9].a/U4185  ( .A(n16978), .B(n16977), .Z(\SUBBYTES[9].a/w1052 ) );
  XOR \SUBBYTES[9].a/U4184  ( .A(\w1[9][89] ), .B(n16979), .Z(n16977) );
  XOR \SUBBYTES[9].a/U4183  ( .A(\SUBBYTES[9].a/w1027 ), .B(
        \SUBBYTES[9].a/w1029 ), .Z(n16978) );
  XOR \SUBBYTES[9].a/U4182  ( .A(\SUBBYTES[9].a/w1011 ), .B(
        \SUBBYTES[9].a/w1012 ), .Z(n16979) );
  XOR \SUBBYTES[9].a/U4181  ( .A(\w1[9][97] ), .B(n16980), .Z(n17308) );
  XOR \SUBBYTES[9].a/U4180  ( .A(\w1[9][99] ), .B(\w1[9][98] ), .Z(n16980) );
  XOR \SUBBYTES[9].a/U4179  ( .A(\w1[9][102] ), .B(n17308), .Z(
        \SUBBYTES[9].a/w894 ) );
  XOR \SUBBYTES[9].a/U4178  ( .A(\w1[9][96] ), .B(\SUBBYTES[9].a/w894 ), .Z(
        \SUBBYTES[9].a/w781 ) );
  XOR \SUBBYTES[9].a/U4177  ( .A(\w1[9][96] ), .B(n16981), .Z(
        \SUBBYTES[9].a/w782 ) );
  XOR \SUBBYTES[9].a/U4176  ( .A(\w1[9][102] ), .B(\w1[9][101] ), .Z(n16981)
         );
  XOR \SUBBYTES[9].a/U4175  ( .A(\w1[9][101] ), .B(n17308), .Z(
        \SUBBYTES[9].a/w912 ) );
  XOR \SUBBYTES[9].a/U4174  ( .A(n16983), .B(n16982), .Z(\SUBBYTES[9].a/w905 )
         );
  XOR \SUBBYTES[9].a/U4173  ( .A(\w1[9][99] ), .B(\w1[9][97] ), .Z(n16982) );
  XOR \SUBBYTES[9].a/U4172  ( .A(\w1[9][103] ), .B(\w1[9][100] ), .Z(n16983)
         );
  XOR \SUBBYTES[9].a/U4171  ( .A(\w1[9][96] ), .B(\SUBBYTES[9].a/w905 ), .Z(
        \SUBBYTES[9].a/w784 ) );
  XOR \SUBBYTES[9].a/U4170  ( .A(n16985), .B(n16984), .Z(\SUBBYTES[9].a/w892 )
         );
  XOR \SUBBYTES[9].a/U4169  ( .A(\SUBBYTES[9].a/w853 ), .B(n1088), .Z(n16984)
         );
  XOR \SUBBYTES[9].a/U4168  ( .A(\SUBBYTES[9].a/w846 ), .B(
        \SUBBYTES[9].a/w849 ), .Z(n16985) );
  XOR \SUBBYTES[9].a/U4167  ( .A(n16987), .B(n16986), .Z(\SUBBYTES[9].a/w893 )
         );
  XOR \SUBBYTES[9].a/U4166  ( .A(\SUBBYTES[9].a/w853 ), .B(n16079), .Z(n16986)
         );
  XOR \SUBBYTES[9].a/U4165  ( .A(\SUBBYTES[9].a/w846 ), .B(n16078), .Z(n16987)
         );
  XOR \SUBBYTES[9].a/U4164  ( .A(\SUBBYTES[9].a/w905 ), .B(n16988), .Z(
        \SUBBYTES[9].a/w895 ) );
  XOR \SUBBYTES[9].a/U4163  ( .A(\w1[9][102] ), .B(\w1[9][101] ), .Z(n16988)
         );
  XOR \SUBBYTES[9].a/U4162  ( .A(n16990), .B(n16989), .Z(\SUBBYTES[9].a/w896 )
         );
  XOR \SUBBYTES[9].a/U4161  ( .A(n16079), .B(n1088), .Z(n16989) );
  XOR \SUBBYTES[9].a/U4160  ( .A(n16078), .B(\SUBBYTES[9].a/w849 ), .Z(n16990)
         );
  XOR \SUBBYTES[9].a/U4159  ( .A(\w1[9][103] ), .B(\w1[9][98] ), .Z(n17314) );
  XOR \SUBBYTES[9].a/U4158  ( .A(n17314), .B(n16991), .Z(\SUBBYTES[9].a/w897 )
         );
  XOR \SUBBYTES[9].a/U4157  ( .A(\w1[9][101] ), .B(\w1[9][100] ), .Z(n16991)
         );
  XOR \SUBBYTES[9].a/U4156  ( .A(\w1[9][103] ), .B(\SUBBYTES[9].a/w782 ), .Z(
        \SUBBYTES[9].a/w785 ) );
  XOR \SUBBYTES[9].a/U4155  ( .A(\w1[9][97] ), .B(\SUBBYTES[9].a/w782 ), .Z(
        \SUBBYTES[9].a/w786 ) );
  XOR \SUBBYTES[9].a/U4154  ( .A(\w1[9][100] ), .B(\SUBBYTES[9].a/w782 ), .Z(
        \SUBBYTES[9].a/w787 ) );
  XOR \SUBBYTES[9].a/U4153  ( .A(\SUBBYTES[9].a/w786 ), .B(n17314), .Z(
        \SUBBYTES[9].a/w788 ) );
  XOR \SUBBYTES[9].a/U4152  ( .A(n17314), .B(n16992), .Z(\SUBBYTES[9].a/w873 )
         );
  XOR \SUBBYTES[9].a/U4151  ( .A(\w1[9][100] ), .B(\w1[9][97] ), .Z(n16992) );
  XOR \SUBBYTES[9].a/U4150  ( .A(n16994), .B(n16993), .Z(n17311) );
  XOR \SUBBYTES[9].a/U4149  ( .A(\w1[9][100] ), .B(n16995), .Z(n16993) );
  XOR \SUBBYTES[9].a/U4148  ( .A(\SUBBYTES[9].a/w838 ), .B(\w1[9][102] ), .Z(
        n16994) );
  XOR \SUBBYTES[9].a/U4147  ( .A(\SUBBYTES[9].a/w812 ), .B(
        \SUBBYTES[9].a/w819 ), .Z(n16995) );
  XOR \SUBBYTES[9].a/U4146  ( .A(n16997), .B(n16996), .Z(n17309) );
  XOR \SUBBYTES[9].a/U4145  ( .A(\w1[9][97] ), .B(n16998), .Z(n16996) );
  XOR \SUBBYTES[9].a/U4144  ( .A(\SUBBYTES[9].a/w837 ), .B(\w1[9][101] ), .Z(
        n16997) );
  XOR \SUBBYTES[9].a/U4143  ( .A(\SUBBYTES[9].a/w813 ), .B(
        \SUBBYTES[9].a/w820 ), .Z(n16998) );
  XOR \SUBBYTES[9].a/U4142  ( .A(n17311), .B(n17309), .Z(\SUBBYTES[9].a/w843 )
         );
  XOR \SUBBYTES[9].a/U4141  ( .A(\w1[9][101] ), .B(n16999), .Z(n17312) );
  XOR \SUBBYTES[9].a/U4140  ( .A(\SUBBYTES[9].a/w805 ), .B(
        \SUBBYTES[9].a/w815 ), .Z(n16999) );
  XOR \SUBBYTES[9].a/U4139  ( .A(n17001), .B(n17000), .Z(\SUBBYTES[9].a/w830 )
         );
  XOR \SUBBYTES[9].a/U4138  ( .A(n17312), .B(n17002), .Z(n17000) );
  XOR \SUBBYTES[9].a/U4137  ( .A(\w1[9][100] ), .B(\SUBBYTES[9].a/w894 ), .Z(
        n17001) );
  XOR \SUBBYTES[9].a/U4136  ( .A(\SUBBYTES[9].a/w807 ), .B(
        \SUBBYTES[9].a/w812 ), .Z(n17002) );
  XOR \SUBBYTES[9].a/U4135  ( .A(n17004), .B(n17003), .Z(n17310) );
  XOR \SUBBYTES[9].a/U4134  ( .A(\SUBBYTES[9].a/w840 ), .B(\w1[9][103] ), .Z(
        n17003) );
  XOR \SUBBYTES[9].a/U4133  ( .A(\SUBBYTES[9].a/w815 ), .B(
        \SUBBYTES[9].a/w822 ), .Z(n17004) );
  XOR \SUBBYTES[9].a/U4132  ( .A(n17309), .B(n17310), .Z(\SUBBYTES[9].a/w842 )
         );
  XOR \SUBBYTES[9].a/U4131  ( .A(\w1[9][99] ), .B(n17005), .Z(n17313) );
  XOR \SUBBYTES[9].a/U4130  ( .A(\SUBBYTES[9].a/w804 ), .B(
        \SUBBYTES[9].a/w807 ), .Z(n17005) );
  XOR \SUBBYTES[9].a/U4129  ( .A(n17007), .B(n17006), .Z(\SUBBYTES[9].a/w831 )
         );
  XOR \SUBBYTES[9].a/U4128  ( .A(n17313), .B(n17008), .Z(n17006) );
  XOR \SUBBYTES[9].a/U4127  ( .A(\w1[9][102] ), .B(\SUBBYTES[9].a/w873 ), .Z(
        n17007) );
  XOR \SUBBYTES[9].a/U4126  ( .A(\SUBBYTES[9].a/w812 ), .B(
        \SUBBYTES[9].a/w813 ), .Z(n17008) );
  XOR \SUBBYTES[9].a/U4125  ( .A(n17311), .B(n17310), .Z(\SUBBYTES[9].a/w851 )
         );
  XOR \SUBBYTES[9].a/U4124  ( .A(n17010), .B(n17009), .Z(\SUBBYTES[9].a/w852 )
         );
  XOR \SUBBYTES[9].a/U4123  ( .A(\w1[9][103] ), .B(n17312), .Z(n17009) );
  XOR \SUBBYTES[9].a/U4122  ( .A(\SUBBYTES[9].a/w804 ), .B(
        \SUBBYTES[9].a/w813 ), .Z(n17010) );
  XOR \SUBBYTES[9].a/U4121  ( .A(n17012), .B(n17011), .Z(\SUBBYTES[9].a/w828 )
         );
  XOR \SUBBYTES[9].a/U4120  ( .A(n17014), .B(n17013), .Z(n17011) );
  XOR \SUBBYTES[9].a/U4119  ( .A(\w1[9][103] ), .B(\SUBBYTES[9].a/w912 ), .Z(
        n17012) );
  XOR \SUBBYTES[9].a/U4118  ( .A(\SUBBYTES[9].a/w819 ), .B(
        \SUBBYTES[9].a/w822 ), .Z(n17013) );
  XOR \SUBBYTES[9].a/U4117  ( .A(\SUBBYTES[9].a/w805 ), .B(
        \SUBBYTES[9].a/w807 ), .Z(n17014) );
  XOR \SUBBYTES[9].a/U4116  ( .A(n17016), .B(n17015), .Z(\SUBBYTES[9].a/w829 )
         );
  XOR \SUBBYTES[9].a/U4115  ( .A(n17313), .B(n17017), .Z(n17015) );
  XOR \SUBBYTES[9].a/U4114  ( .A(\w1[9][101] ), .B(n17314), .Z(n17016) );
  XOR \SUBBYTES[9].a/U4113  ( .A(\SUBBYTES[9].a/w819 ), .B(
        \SUBBYTES[9].a/w820 ), .Z(n17017) );
  XOR \SUBBYTES[9].a/U4112  ( .A(n17019), .B(n17018), .Z(\SUBBYTES[9].a/w845 )
         );
  XOR \SUBBYTES[9].a/U4111  ( .A(\w1[9][97] ), .B(n17020), .Z(n17018) );
  XOR \SUBBYTES[9].a/U4110  ( .A(\SUBBYTES[9].a/w820 ), .B(
        \SUBBYTES[9].a/w822 ), .Z(n17019) );
  XOR \SUBBYTES[9].a/U4109  ( .A(\SUBBYTES[9].a/w804 ), .B(
        \SUBBYTES[9].a/w805 ), .Z(n17020) );
  XOR \SUBBYTES[9].a/U4108  ( .A(\w1[9][105] ), .B(n17021), .Z(n17315) );
  XOR \SUBBYTES[9].a/U4107  ( .A(\w1[9][107] ), .B(\w1[9][106] ), .Z(n17021)
         );
  XOR \SUBBYTES[9].a/U4106  ( .A(\w1[9][110] ), .B(n17315), .Z(
        \SUBBYTES[9].a/w687 ) );
  XOR \SUBBYTES[9].a/U4105  ( .A(\w1[9][104] ), .B(\SUBBYTES[9].a/w687 ), .Z(
        \SUBBYTES[9].a/w574 ) );
  XOR \SUBBYTES[9].a/U4104  ( .A(\w1[9][104] ), .B(n17022), .Z(
        \SUBBYTES[9].a/w575 ) );
  XOR \SUBBYTES[9].a/U4103  ( .A(\w1[9][110] ), .B(\w1[9][109] ), .Z(n17022)
         );
  XOR \SUBBYTES[9].a/U4102  ( .A(\w1[9][109] ), .B(n17315), .Z(
        \SUBBYTES[9].a/w705 ) );
  XOR \SUBBYTES[9].a/U4101  ( .A(n17024), .B(n17023), .Z(\SUBBYTES[9].a/w698 )
         );
  XOR \SUBBYTES[9].a/U4100  ( .A(\w1[9][107] ), .B(\w1[9][105] ), .Z(n17023)
         );
  XOR \SUBBYTES[9].a/U4099  ( .A(\w1[9][111] ), .B(\w1[9][108] ), .Z(n17024)
         );
  XOR \SUBBYTES[9].a/U4098  ( .A(\w1[9][104] ), .B(\SUBBYTES[9].a/w698 ), .Z(
        \SUBBYTES[9].a/w577 ) );
  XOR \SUBBYTES[9].a/U4097  ( .A(n17026), .B(n17025), .Z(\SUBBYTES[9].a/w685 )
         );
  XOR \SUBBYTES[9].a/U4096  ( .A(\SUBBYTES[9].a/w646 ), .B(n1087), .Z(n17025)
         );
  XOR \SUBBYTES[9].a/U4095  ( .A(\SUBBYTES[9].a/w639 ), .B(
        \SUBBYTES[9].a/w642 ), .Z(n17026) );
  XOR \SUBBYTES[9].a/U4094  ( .A(n17028), .B(n17027), .Z(\SUBBYTES[9].a/w686 )
         );
  XOR \SUBBYTES[9].a/U4093  ( .A(\SUBBYTES[9].a/w646 ), .B(n16077), .Z(n17027)
         );
  XOR \SUBBYTES[9].a/U4092  ( .A(\SUBBYTES[9].a/w639 ), .B(n16076), .Z(n17028)
         );
  XOR \SUBBYTES[9].a/U4091  ( .A(\SUBBYTES[9].a/w698 ), .B(n17029), .Z(
        \SUBBYTES[9].a/w688 ) );
  XOR \SUBBYTES[9].a/U4090  ( .A(\w1[9][110] ), .B(\w1[9][109] ), .Z(n17029)
         );
  XOR \SUBBYTES[9].a/U4089  ( .A(n17031), .B(n17030), .Z(\SUBBYTES[9].a/w689 )
         );
  XOR \SUBBYTES[9].a/U4088  ( .A(n16077), .B(n1087), .Z(n17030) );
  XOR \SUBBYTES[9].a/U4087  ( .A(n16076), .B(\SUBBYTES[9].a/w642 ), .Z(n17031)
         );
  XOR \SUBBYTES[9].a/U4086  ( .A(\w1[9][111] ), .B(\w1[9][106] ), .Z(n17321)
         );
  XOR \SUBBYTES[9].a/U4085  ( .A(n17321), .B(n17032), .Z(\SUBBYTES[9].a/w690 )
         );
  XOR \SUBBYTES[9].a/U4084  ( .A(\w1[9][109] ), .B(\w1[9][108] ), .Z(n17032)
         );
  XOR \SUBBYTES[9].a/U4083  ( .A(\w1[9][111] ), .B(\SUBBYTES[9].a/w575 ), .Z(
        \SUBBYTES[9].a/w578 ) );
  XOR \SUBBYTES[9].a/U4082  ( .A(\w1[9][105] ), .B(\SUBBYTES[9].a/w575 ), .Z(
        \SUBBYTES[9].a/w579 ) );
  XOR \SUBBYTES[9].a/U4081  ( .A(\w1[9][108] ), .B(\SUBBYTES[9].a/w575 ), .Z(
        \SUBBYTES[9].a/w580 ) );
  XOR \SUBBYTES[9].a/U4080  ( .A(\SUBBYTES[9].a/w579 ), .B(n17321), .Z(
        \SUBBYTES[9].a/w581 ) );
  XOR \SUBBYTES[9].a/U4079  ( .A(n17321), .B(n17033), .Z(\SUBBYTES[9].a/w666 )
         );
  XOR \SUBBYTES[9].a/U4078  ( .A(\w1[9][108] ), .B(\w1[9][105] ), .Z(n17033)
         );
  XOR \SUBBYTES[9].a/U4077  ( .A(n17035), .B(n17034), .Z(n17318) );
  XOR \SUBBYTES[9].a/U4076  ( .A(\w1[9][108] ), .B(n17036), .Z(n17034) );
  XOR \SUBBYTES[9].a/U4075  ( .A(\SUBBYTES[9].a/w631 ), .B(\w1[9][110] ), .Z(
        n17035) );
  XOR \SUBBYTES[9].a/U4074  ( .A(\SUBBYTES[9].a/w605 ), .B(
        \SUBBYTES[9].a/w612 ), .Z(n17036) );
  XOR \SUBBYTES[9].a/U4073  ( .A(n17038), .B(n17037), .Z(n17316) );
  XOR \SUBBYTES[9].a/U4072  ( .A(\w1[9][105] ), .B(n17039), .Z(n17037) );
  XOR \SUBBYTES[9].a/U4071  ( .A(\SUBBYTES[9].a/w630 ), .B(\w1[9][109] ), .Z(
        n17038) );
  XOR \SUBBYTES[9].a/U4070  ( .A(\SUBBYTES[9].a/w606 ), .B(
        \SUBBYTES[9].a/w613 ), .Z(n17039) );
  XOR \SUBBYTES[9].a/U4069  ( .A(n17318), .B(n17316), .Z(\SUBBYTES[9].a/w636 )
         );
  XOR \SUBBYTES[9].a/U4068  ( .A(\w1[9][109] ), .B(n17040), .Z(n17319) );
  XOR \SUBBYTES[9].a/U4067  ( .A(\SUBBYTES[9].a/w598 ), .B(
        \SUBBYTES[9].a/w608 ), .Z(n17040) );
  XOR \SUBBYTES[9].a/U4066  ( .A(n17042), .B(n17041), .Z(\SUBBYTES[9].a/w623 )
         );
  XOR \SUBBYTES[9].a/U4065  ( .A(n17319), .B(n17043), .Z(n17041) );
  XOR \SUBBYTES[9].a/U4064  ( .A(\w1[9][108] ), .B(\SUBBYTES[9].a/w687 ), .Z(
        n17042) );
  XOR \SUBBYTES[9].a/U4063  ( .A(\SUBBYTES[9].a/w600 ), .B(
        \SUBBYTES[9].a/w605 ), .Z(n17043) );
  XOR \SUBBYTES[9].a/U4062  ( .A(n17045), .B(n17044), .Z(n17317) );
  XOR \SUBBYTES[9].a/U4061  ( .A(\SUBBYTES[9].a/w633 ), .B(\w1[9][111] ), .Z(
        n17044) );
  XOR \SUBBYTES[9].a/U4060  ( .A(\SUBBYTES[9].a/w608 ), .B(
        \SUBBYTES[9].a/w615 ), .Z(n17045) );
  XOR \SUBBYTES[9].a/U4059  ( .A(n17316), .B(n17317), .Z(\SUBBYTES[9].a/w635 )
         );
  XOR \SUBBYTES[9].a/U4058  ( .A(\w1[9][107] ), .B(n17046), .Z(n17320) );
  XOR \SUBBYTES[9].a/U4057  ( .A(\SUBBYTES[9].a/w597 ), .B(
        \SUBBYTES[9].a/w600 ), .Z(n17046) );
  XOR \SUBBYTES[9].a/U4056  ( .A(n17048), .B(n17047), .Z(\SUBBYTES[9].a/w624 )
         );
  XOR \SUBBYTES[9].a/U4055  ( .A(n17320), .B(n17049), .Z(n17047) );
  XOR \SUBBYTES[9].a/U4054  ( .A(\w1[9][110] ), .B(\SUBBYTES[9].a/w666 ), .Z(
        n17048) );
  XOR \SUBBYTES[9].a/U4053  ( .A(\SUBBYTES[9].a/w605 ), .B(
        \SUBBYTES[9].a/w606 ), .Z(n17049) );
  XOR \SUBBYTES[9].a/U4052  ( .A(n17318), .B(n17317), .Z(\SUBBYTES[9].a/w644 )
         );
  XOR \SUBBYTES[9].a/U4051  ( .A(n17051), .B(n17050), .Z(\SUBBYTES[9].a/w645 )
         );
  XOR \SUBBYTES[9].a/U4050  ( .A(\w1[9][111] ), .B(n17319), .Z(n17050) );
  XOR \SUBBYTES[9].a/U4049  ( .A(\SUBBYTES[9].a/w597 ), .B(
        \SUBBYTES[9].a/w606 ), .Z(n17051) );
  XOR \SUBBYTES[9].a/U4048  ( .A(n17053), .B(n17052), .Z(\SUBBYTES[9].a/w621 )
         );
  XOR \SUBBYTES[9].a/U4047  ( .A(n17055), .B(n17054), .Z(n17052) );
  XOR \SUBBYTES[9].a/U4046  ( .A(\w1[9][111] ), .B(\SUBBYTES[9].a/w705 ), .Z(
        n17053) );
  XOR \SUBBYTES[9].a/U4045  ( .A(\SUBBYTES[9].a/w612 ), .B(
        \SUBBYTES[9].a/w615 ), .Z(n17054) );
  XOR \SUBBYTES[9].a/U4044  ( .A(\SUBBYTES[9].a/w598 ), .B(
        \SUBBYTES[9].a/w600 ), .Z(n17055) );
  XOR \SUBBYTES[9].a/U4043  ( .A(n17057), .B(n17056), .Z(\SUBBYTES[9].a/w622 )
         );
  XOR \SUBBYTES[9].a/U4042  ( .A(n17320), .B(n17058), .Z(n17056) );
  XOR \SUBBYTES[9].a/U4041  ( .A(\w1[9][109] ), .B(n17321), .Z(n17057) );
  XOR \SUBBYTES[9].a/U4040  ( .A(\SUBBYTES[9].a/w612 ), .B(
        \SUBBYTES[9].a/w613 ), .Z(n17058) );
  XOR \SUBBYTES[9].a/U4039  ( .A(n17060), .B(n17059), .Z(\SUBBYTES[9].a/w638 )
         );
  XOR \SUBBYTES[9].a/U4038  ( .A(\w1[9][105] ), .B(n17061), .Z(n17059) );
  XOR \SUBBYTES[9].a/U4037  ( .A(\SUBBYTES[9].a/w613 ), .B(
        \SUBBYTES[9].a/w615 ), .Z(n17060) );
  XOR \SUBBYTES[9].a/U4036  ( .A(\SUBBYTES[9].a/w597 ), .B(
        \SUBBYTES[9].a/w598 ), .Z(n17061) );
  XOR \SUBBYTES[9].a/U4035  ( .A(\w1[9][113] ), .B(n17062), .Z(n17322) );
  XOR \SUBBYTES[9].a/U4034  ( .A(\w1[9][115] ), .B(\w1[9][114] ), .Z(n17062)
         );
  XOR \SUBBYTES[9].a/U4033  ( .A(\w1[9][118] ), .B(n17322), .Z(
        \SUBBYTES[9].a/w480 ) );
  XOR \SUBBYTES[9].a/U4032  ( .A(\w1[9][112] ), .B(\SUBBYTES[9].a/w480 ), .Z(
        \SUBBYTES[9].a/w367 ) );
  XOR \SUBBYTES[9].a/U4031  ( .A(\w1[9][112] ), .B(n17063), .Z(
        \SUBBYTES[9].a/w368 ) );
  XOR \SUBBYTES[9].a/U4030  ( .A(\w1[9][118] ), .B(\w1[9][117] ), .Z(n17063)
         );
  XOR \SUBBYTES[9].a/U4029  ( .A(\w1[9][117] ), .B(n17322), .Z(
        \SUBBYTES[9].a/w498 ) );
  XOR \SUBBYTES[9].a/U4028  ( .A(n17065), .B(n17064), .Z(\SUBBYTES[9].a/w491 )
         );
  XOR \SUBBYTES[9].a/U4027  ( .A(\w1[9][115] ), .B(\w1[9][113] ), .Z(n17064)
         );
  XOR \SUBBYTES[9].a/U4026  ( .A(\w1[9][119] ), .B(\w1[9][116] ), .Z(n17065)
         );
  XOR \SUBBYTES[9].a/U4025  ( .A(\w1[9][112] ), .B(\SUBBYTES[9].a/w491 ), .Z(
        \SUBBYTES[9].a/w370 ) );
  XOR \SUBBYTES[9].a/U4024  ( .A(n17067), .B(n17066), .Z(\SUBBYTES[9].a/w478 )
         );
  XOR \SUBBYTES[9].a/U4023  ( .A(\SUBBYTES[9].a/w439 ), .B(n1086), .Z(n17066)
         );
  XOR \SUBBYTES[9].a/U4022  ( .A(\SUBBYTES[9].a/w432 ), .B(
        \SUBBYTES[9].a/w435 ), .Z(n17067) );
  XOR \SUBBYTES[9].a/U4021  ( .A(n17069), .B(n17068), .Z(\SUBBYTES[9].a/w479 )
         );
  XOR \SUBBYTES[9].a/U4020  ( .A(\SUBBYTES[9].a/w439 ), .B(n16075), .Z(n17068)
         );
  XOR \SUBBYTES[9].a/U4019  ( .A(\SUBBYTES[9].a/w432 ), .B(n16074), .Z(n17069)
         );
  XOR \SUBBYTES[9].a/U4018  ( .A(\SUBBYTES[9].a/w491 ), .B(n17070), .Z(
        \SUBBYTES[9].a/w481 ) );
  XOR \SUBBYTES[9].a/U4017  ( .A(\w1[9][118] ), .B(\w1[9][117] ), .Z(n17070)
         );
  XOR \SUBBYTES[9].a/U4016  ( .A(n17072), .B(n17071), .Z(\SUBBYTES[9].a/w482 )
         );
  XOR \SUBBYTES[9].a/U4015  ( .A(n16075), .B(n1086), .Z(n17071) );
  XOR \SUBBYTES[9].a/U4014  ( .A(n16074), .B(\SUBBYTES[9].a/w435 ), .Z(n17072)
         );
  XOR \SUBBYTES[9].a/U4013  ( .A(\w1[9][119] ), .B(\w1[9][114] ), .Z(n17328)
         );
  XOR \SUBBYTES[9].a/U4012  ( .A(n17328), .B(n17073), .Z(\SUBBYTES[9].a/w483 )
         );
  XOR \SUBBYTES[9].a/U4011  ( .A(\w1[9][117] ), .B(\w1[9][116] ), .Z(n17073)
         );
  XOR \SUBBYTES[9].a/U4010  ( .A(\w1[9][119] ), .B(\SUBBYTES[9].a/w368 ), .Z(
        \SUBBYTES[9].a/w371 ) );
  XOR \SUBBYTES[9].a/U4009  ( .A(\w1[9][113] ), .B(\SUBBYTES[9].a/w368 ), .Z(
        \SUBBYTES[9].a/w372 ) );
  XOR \SUBBYTES[9].a/U4008  ( .A(\w1[9][116] ), .B(\SUBBYTES[9].a/w368 ), .Z(
        \SUBBYTES[9].a/w373 ) );
  XOR \SUBBYTES[9].a/U4007  ( .A(\SUBBYTES[9].a/w372 ), .B(n17328), .Z(
        \SUBBYTES[9].a/w374 ) );
  XOR \SUBBYTES[9].a/U4006  ( .A(n17328), .B(n17074), .Z(\SUBBYTES[9].a/w459 )
         );
  XOR \SUBBYTES[9].a/U4005  ( .A(\w1[9][116] ), .B(\w1[9][113] ), .Z(n17074)
         );
  XOR \SUBBYTES[9].a/U4004  ( .A(n17076), .B(n17075), .Z(n17325) );
  XOR \SUBBYTES[9].a/U4003  ( .A(\w1[9][116] ), .B(n17077), .Z(n17075) );
  XOR \SUBBYTES[9].a/U4002  ( .A(\SUBBYTES[9].a/w424 ), .B(\w1[9][118] ), .Z(
        n17076) );
  XOR \SUBBYTES[9].a/U4001  ( .A(\SUBBYTES[9].a/w398 ), .B(
        \SUBBYTES[9].a/w405 ), .Z(n17077) );
  XOR \SUBBYTES[9].a/U4000  ( .A(n17079), .B(n17078), .Z(n17323) );
  XOR \SUBBYTES[9].a/U3999  ( .A(\w1[9][113] ), .B(n17080), .Z(n17078) );
  XOR \SUBBYTES[9].a/U3998  ( .A(\SUBBYTES[9].a/w423 ), .B(\w1[9][117] ), .Z(
        n17079) );
  XOR \SUBBYTES[9].a/U3997  ( .A(\SUBBYTES[9].a/w399 ), .B(
        \SUBBYTES[9].a/w406 ), .Z(n17080) );
  XOR \SUBBYTES[9].a/U3996  ( .A(n17325), .B(n17323), .Z(\SUBBYTES[9].a/w429 )
         );
  XOR \SUBBYTES[9].a/U3995  ( .A(\w1[9][117] ), .B(n17081), .Z(n17326) );
  XOR \SUBBYTES[9].a/U3994  ( .A(\SUBBYTES[9].a/w391 ), .B(
        \SUBBYTES[9].a/w401 ), .Z(n17081) );
  XOR \SUBBYTES[9].a/U3993  ( .A(n17083), .B(n17082), .Z(\SUBBYTES[9].a/w416 )
         );
  XOR \SUBBYTES[9].a/U3992  ( .A(n17326), .B(n17084), .Z(n17082) );
  XOR \SUBBYTES[9].a/U3991  ( .A(\w1[9][116] ), .B(\SUBBYTES[9].a/w480 ), .Z(
        n17083) );
  XOR \SUBBYTES[9].a/U3990  ( .A(\SUBBYTES[9].a/w393 ), .B(
        \SUBBYTES[9].a/w398 ), .Z(n17084) );
  XOR \SUBBYTES[9].a/U3989  ( .A(n17086), .B(n17085), .Z(n17324) );
  XOR \SUBBYTES[9].a/U3988  ( .A(\SUBBYTES[9].a/w426 ), .B(\w1[9][119] ), .Z(
        n17085) );
  XOR \SUBBYTES[9].a/U3987  ( .A(\SUBBYTES[9].a/w401 ), .B(
        \SUBBYTES[9].a/w408 ), .Z(n17086) );
  XOR \SUBBYTES[9].a/U3986  ( .A(n17323), .B(n17324), .Z(\SUBBYTES[9].a/w428 )
         );
  XOR \SUBBYTES[9].a/U3985  ( .A(\w1[9][115] ), .B(n17087), .Z(n17327) );
  XOR \SUBBYTES[9].a/U3984  ( .A(\SUBBYTES[9].a/w390 ), .B(
        \SUBBYTES[9].a/w393 ), .Z(n17087) );
  XOR \SUBBYTES[9].a/U3983  ( .A(n17089), .B(n17088), .Z(\SUBBYTES[9].a/w417 )
         );
  XOR \SUBBYTES[9].a/U3982  ( .A(n17327), .B(n17090), .Z(n17088) );
  XOR \SUBBYTES[9].a/U3981  ( .A(\w1[9][118] ), .B(\SUBBYTES[9].a/w459 ), .Z(
        n17089) );
  XOR \SUBBYTES[9].a/U3980  ( .A(\SUBBYTES[9].a/w398 ), .B(
        \SUBBYTES[9].a/w399 ), .Z(n17090) );
  XOR \SUBBYTES[9].a/U3979  ( .A(n17325), .B(n17324), .Z(\SUBBYTES[9].a/w437 )
         );
  XOR \SUBBYTES[9].a/U3978  ( .A(n17092), .B(n17091), .Z(\SUBBYTES[9].a/w438 )
         );
  XOR \SUBBYTES[9].a/U3977  ( .A(\w1[9][119] ), .B(n17326), .Z(n17091) );
  XOR \SUBBYTES[9].a/U3976  ( .A(\SUBBYTES[9].a/w390 ), .B(
        \SUBBYTES[9].a/w399 ), .Z(n17092) );
  XOR \SUBBYTES[9].a/U3975  ( .A(n17094), .B(n17093), .Z(\SUBBYTES[9].a/w414 )
         );
  XOR \SUBBYTES[9].a/U3974  ( .A(n17096), .B(n17095), .Z(n17093) );
  XOR \SUBBYTES[9].a/U3973  ( .A(\w1[9][119] ), .B(\SUBBYTES[9].a/w498 ), .Z(
        n17094) );
  XOR \SUBBYTES[9].a/U3972  ( .A(\SUBBYTES[9].a/w405 ), .B(
        \SUBBYTES[9].a/w408 ), .Z(n17095) );
  XOR \SUBBYTES[9].a/U3971  ( .A(\SUBBYTES[9].a/w391 ), .B(
        \SUBBYTES[9].a/w393 ), .Z(n17096) );
  XOR \SUBBYTES[9].a/U3970  ( .A(n17098), .B(n17097), .Z(\SUBBYTES[9].a/w415 )
         );
  XOR \SUBBYTES[9].a/U3969  ( .A(n17327), .B(n17099), .Z(n17097) );
  XOR \SUBBYTES[9].a/U3968  ( .A(\w1[9][117] ), .B(n17328), .Z(n17098) );
  XOR \SUBBYTES[9].a/U3967  ( .A(\SUBBYTES[9].a/w405 ), .B(
        \SUBBYTES[9].a/w406 ), .Z(n17099) );
  XOR \SUBBYTES[9].a/U3966  ( .A(n17101), .B(n17100), .Z(\SUBBYTES[9].a/w431 )
         );
  XOR \SUBBYTES[9].a/U3965  ( .A(\w1[9][113] ), .B(n17102), .Z(n17100) );
  XOR \SUBBYTES[9].a/U3964  ( .A(\SUBBYTES[9].a/w406 ), .B(
        \SUBBYTES[9].a/w408 ), .Z(n17101) );
  XOR \SUBBYTES[9].a/U3963  ( .A(\SUBBYTES[9].a/w390 ), .B(
        \SUBBYTES[9].a/w391 ), .Z(n17102) );
  XOR \SUBBYTES[9].a/U3962  ( .A(\w1[9][121] ), .B(n17103), .Z(n17329) );
  XOR \SUBBYTES[9].a/U3961  ( .A(\w1[9][123] ), .B(\w1[9][122] ), .Z(n17103)
         );
  XOR \SUBBYTES[9].a/U3960  ( .A(\w1[9][126] ), .B(n17329), .Z(
        \SUBBYTES[9].a/w273 ) );
  XOR \SUBBYTES[9].a/U3959  ( .A(\w1[9][120] ), .B(\SUBBYTES[9].a/w273 ), .Z(
        \SUBBYTES[9].a/w160 ) );
  XOR \SUBBYTES[9].a/U3958  ( .A(\w1[9][120] ), .B(n17104), .Z(
        \SUBBYTES[9].a/w161 ) );
  XOR \SUBBYTES[9].a/U3957  ( .A(\w1[9][126] ), .B(\w1[9][125] ), .Z(n17104)
         );
  XOR \SUBBYTES[9].a/U3956  ( .A(\w1[9][125] ), .B(n17329), .Z(
        \SUBBYTES[9].a/w291 ) );
  XOR \SUBBYTES[9].a/U3955  ( .A(n17106), .B(n17105), .Z(\SUBBYTES[9].a/w284 )
         );
  XOR \SUBBYTES[9].a/U3954  ( .A(\w1[9][123] ), .B(\w1[9][121] ), .Z(n17105)
         );
  XOR \SUBBYTES[9].a/U3953  ( .A(\w1[9][127] ), .B(\w1[9][124] ), .Z(n17106)
         );
  XOR \SUBBYTES[9].a/U3952  ( .A(\w1[9][120] ), .B(\SUBBYTES[9].a/w284 ), .Z(
        \SUBBYTES[9].a/w163 ) );
  XOR \SUBBYTES[9].a/U3951  ( .A(n17108), .B(n17107), .Z(\SUBBYTES[9].a/w271 )
         );
  XOR \SUBBYTES[9].a/U3950  ( .A(\SUBBYTES[9].a/w232 ), .B(n1085), .Z(n17107)
         );
  XOR \SUBBYTES[9].a/U3949  ( .A(\SUBBYTES[9].a/w225 ), .B(
        \SUBBYTES[9].a/w228 ), .Z(n17108) );
  XOR \SUBBYTES[9].a/U3948  ( .A(n17110), .B(n17109), .Z(\SUBBYTES[9].a/w272 )
         );
  XOR \SUBBYTES[9].a/U3947  ( .A(\SUBBYTES[9].a/w232 ), .B(n16073), .Z(n17109)
         );
  XOR \SUBBYTES[9].a/U3946  ( .A(\SUBBYTES[9].a/w225 ), .B(n16072), .Z(n17110)
         );
  XOR \SUBBYTES[9].a/U3945  ( .A(\SUBBYTES[9].a/w284 ), .B(n17111), .Z(
        \SUBBYTES[9].a/w274 ) );
  XOR \SUBBYTES[9].a/U3944  ( .A(\w1[9][126] ), .B(\w1[9][125] ), .Z(n17111)
         );
  XOR \SUBBYTES[9].a/U3943  ( .A(n17113), .B(n17112), .Z(\SUBBYTES[9].a/w275 )
         );
  XOR \SUBBYTES[9].a/U3942  ( .A(n16073), .B(n1085), .Z(n17112) );
  XOR \SUBBYTES[9].a/U3941  ( .A(n16072), .B(\SUBBYTES[9].a/w228 ), .Z(n17113)
         );
  XOR \SUBBYTES[9].a/U3940  ( .A(\w1[9][127] ), .B(\w1[9][122] ), .Z(n17335)
         );
  XOR \SUBBYTES[9].a/U3939  ( .A(n17335), .B(n17114), .Z(\SUBBYTES[9].a/w276 )
         );
  XOR \SUBBYTES[9].a/U3938  ( .A(\w1[9][125] ), .B(\w1[9][124] ), .Z(n17114)
         );
  XOR \SUBBYTES[9].a/U3937  ( .A(\w1[9][127] ), .B(\SUBBYTES[9].a/w161 ), .Z(
        \SUBBYTES[9].a/w164 ) );
  XOR \SUBBYTES[9].a/U3936  ( .A(\w1[9][121] ), .B(\SUBBYTES[9].a/w161 ), .Z(
        \SUBBYTES[9].a/w165 ) );
  XOR \SUBBYTES[9].a/U3935  ( .A(\w1[9][124] ), .B(\SUBBYTES[9].a/w161 ), .Z(
        \SUBBYTES[9].a/w166 ) );
  XOR \SUBBYTES[9].a/U3934  ( .A(\SUBBYTES[9].a/w165 ), .B(n17335), .Z(
        \SUBBYTES[9].a/w167 ) );
  XOR \SUBBYTES[9].a/U3933  ( .A(n17335), .B(n17115), .Z(\SUBBYTES[9].a/w252 )
         );
  XOR \SUBBYTES[9].a/U3932  ( .A(\w1[9][124] ), .B(\w1[9][121] ), .Z(n17115)
         );
  XOR \SUBBYTES[9].a/U3931  ( .A(n17117), .B(n17116), .Z(n17332) );
  XOR \SUBBYTES[9].a/U3930  ( .A(\w1[9][124] ), .B(n17118), .Z(n17116) );
  XOR \SUBBYTES[9].a/U3929  ( .A(\SUBBYTES[9].a/w217 ), .B(\w1[9][126] ), .Z(
        n17117) );
  XOR \SUBBYTES[9].a/U3928  ( .A(\SUBBYTES[9].a/w191 ), .B(
        \SUBBYTES[9].a/w198 ), .Z(n17118) );
  XOR \SUBBYTES[9].a/U3927  ( .A(n17120), .B(n17119), .Z(n17330) );
  XOR \SUBBYTES[9].a/U3926  ( .A(\w1[9][121] ), .B(n17121), .Z(n17119) );
  XOR \SUBBYTES[9].a/U3925  ( .A(\SUBBYTES[9].a/w216 ), .B(\w1[9][125] ), .Z(
        n17120) );
  XOR \SUBBYTES[9].a/U3924  ( .A(\SUBBYTES[9].a/w192 ), .B(
        \SUBBYTES[9].a/w199 ), .Z(n17121) );
  XOR \SUBBYTES[9].a/U3923  ( .A(n17332), .B(n17330), .Z(\SUBBYTES[9].a/w222 )
         );
  XOR \SUBBYTES[9].a/U3922  ( .A(\w1[9][125] ), .B(n17122), .Z(n17333) );
  XOR \SUBBYTES[9].a/U3921  ( .A(\SUBBYTES[9].a/w184 ), .B(
        \SUBBYTES[9].a/w194 ), .Z(n17122) );
  XOR \SUBBYTES[9].a/U3920  ( .A(n17124), .B(n17123), .Z(\SUBBYTES[9].a/w209 )
         );
  XOR \SUBBYTES[9].a/U3919  ( .A(n17333), .B(n17125), .Z(n17123) );
  XOR \SUBBYTES[9].a/U3918  ( .A(\w1[9][124] ), .B(\SUBBYTES[9].a/w273 ), .Z(
        n17124) );
  XOR \SUBBYTES[9].a/U3917  ( .A(\SUBBYTES[9].a/w186 ), .B(
        \SUBBYTES[9].a/w191 ), .Z(n17125) );
  XOR \SUBBYTES[9].a/U3916  ( .A(n17127), .B(n17126), .Z(n17331) );
  XOR \SUBBYTES[9].a/U3915  ( .A(\SUBBYTES[9].a/w219 ), .B(\w1[9][127] ), .Z(
        n17126) );
  XOR \SUBBYTES[9].a/U3914  ( .A(\SUBBYTES[9].a/w194 ), .B(
        \SUBBYTES[9].a/w201 ), .Z(n17127) );
  XOR \SUBBYTES[9].a/U3913  ( .A(n17330), .B(n17331), .Z(\SUBBYTES[9].a/w221 )
         );
  XOR \SUBBYTES[9].a/U3912  ( .A(\w1[9][123] ), .B(n17128), .Z(n17334) );
  XOR \SUBBYTES[9].a/U3911  ( .A(\SUBBYTES[9].a/w183 ), .B(
        \SUBBYTES[9].a/w186 ), .Z(n17128) );
  XOR \SUBBYTES[9].a/U3910  ( .A(n17130), .B(n17129), .Z(\SUBBYTES[9].a/w210 )
         );
  XOR \SUBBYTES[9].a/U3909  ( .A(n17334), .B(n17131), .Z(n17129) );
  XOR \SUBBYTES[9].a/U3908  ( .A(\w1[9][126] ), .B(\SUBBYTES[9].a/w252 ), .Z(
        n17130) );
  XOR \SUBBYTES[9].a/U3907  ( .A(\SUBBYTES[9].a/w191 ), .B(
        \SUBBYTES[9].a/w192 ), .Z(n17131) );
  XOR \SUBBYTES[9].a/U3906  ( .A(n17332), .B(n17331), .Z(\SUBBYTES[9].a/w230 )
         );
  XOR \SUBBYTES[9].a/U3905  ( .A(n17133), .B(n17132), .Z(\SUBBYTES[9].a/w231 )
         );
  XOR \SUBBYTES[9].a/U3904  ( .A(\w1[9][127] ), .B(n17333), .Z(n17132) );
  XOR \SUBBYTES[9].a/U3903  ( .A(\SUBBYTES[9].a/w183 ), .B(
        \SUBBYTES[9].a/w192 ), .Z(n17133) );
  XOR \SUBBYTES[9].a/U3902  ( .A(n17135), .B(n17134), .Z(\SUBBYTES[9].a/w207 )
         );
  XOR \SUBBYTES[9].a/U3901  ( .A(n17137), .B(n17136), .Z(n17134) );
  XOR \SUBBYTES[9].a/U3900  ( .A(\w1[9][127] ), .B(\SUBBYTES[9].a/w291 ), .Z(
        n17135) );
  XOR \SUBBYTES[9].a/U3899  ( .A(\SUBBYTES[9].a/w198 ), .B(
        \SUBBYTES[9].a/w201 ), .Z(n17136) );
  XOR \SUBBYTES[9].a/U3898  ( .A(\SUBBYTES[9].a/w184 ), .B(
        \SUBBYTES[9].a/w186 ), .Z(n17137) );
  XOR \SUBBYTES[9].a/U3897  ( .A(n17139), .B(n17138), .Z(\SUBBYTES[9].a/w208 )
         );
  XOR \SUBBYTES[9].a/U3896  ( .A(n17334), .B(n17140), .Z(n17138) );
  XOR \SUBBYTES[9].a/U3895  ( .A(\w1[9][125] ), .B(n17335), .Z(n17139) );
  XOR \SUBBYTES[9].a/U3894  ( .A(\SUBBYTES[9].a/w198 ), .B(
        \SUBBYTES[9].a/w199 ), .Z(n17140) );
  XOR \SUBBYTES[9].a/U3893  ( .A(n17142), .B(n17141), .Z(\SUBBYTES[9].a/w224 )
         );
  XOR \SUBBYTES[9].a/U3892  ( .A(\w1[9][121] ), .B(n17143), .Z(n17141) );
  XOR \SUBBYTES[9].a/U3891  ( .A(\SUBBYTES[9].a/w199 ), .B(
        \SUBBYTES[9].a/w201 ), .Z(n17142) );
  XOR \SUBBYTES[9].a/U3890  ( .A(\SUBBYTES[9].a/w183 ), .B(
        \SUBBYTES[9].a/w184 ), .Z(n17143) );
  XOR \SUBBYTES[8].a/U5649  ( .A(\SUBBYTES[8].a/w3390 ), .B(
        \SUBBYTES[8].a/w3391 ), .Z(n15865) );
  XOR \SUBBYTES[8].a/U5648  ( .A(n15865), .B(n14824), .Z(n15864) );
  XOR \SUBBYTES[8].a/U5647  ( .A(\SUBBYTES[8].a/w3383 ), .B(
        \SUBBYTES[8].a/w3400 ), .Z(n14824) );
  XOR \SUBBYTES[8].a/U5645  ( .A(\SUBBYTES[8].a/w3382 ), .B(
        \SUBBYTES[8].a/w3397 ), .Z(n14825) );
  XOR \SUBBYTES[8].a/U5644  ( .A(n15865), .B(n14826), .Z(n16056) );
  XOR \SUBBYTES[8].a/U5643  ( .A(\SUBBYTES[8].a/w3397 ), .B(
        \SUBBYTES[8].a/w3398 ), .Z(n14826) );
  XOR \SUBBYTES[8].a/U5642  ( .A(\SUBBYTES[8].a/w3359 ), .B(n14827), .Z(n15867) );
  XOR \SUBBYTES[8].a/U5641  ( .A(\SUBBYTES[8].a/w3350 ), .B(
        \SUBBYTES[8].a/w3351 ), .Z(n14827) );
  XOR \SUBBYTES[8].a/U5639  ( .A(\SUBBYTES[8].a/w3361 ), .B(n16056), .Z(n14828) );
  XOR \SUBBYTES[8].a/U5638  ( .A(n14830), .B(n14829), .Z(n15868) );
  XOR \SUBBYTES[8].a/U5637  ( .A(n14832), .B(n14831), .Z(n14829) );
  XOR \SUBBYTES[8].a/U5636  ( .A(\SUBBYTES[8].a/w3397 ), .B(
        \SUBBYTES[8].a/w3398 ), .Z(n14830) );
  XOR \SUBBYTES[8].a/U5635  ( .A(\SUBBYTES[8].a/w3361 ), .B(
        \SUBBYTES[8].a/w3385 ), .Z(n14831) );
  XOR \SUBBYTES[8].a/U5634  ( .A(\SUBBYTES[8].a/w3350 ), .B(
        \SUBBYTES[8].a/w3359 ), .Z(n14832) );
  XOR \SUBBYTES[8].a/U5633  ( .A(\SUBBYTES[8].a/w3382 ), .B(n14833), .Z(n15866) );
  XOR \SUBBYTES[8].a/U5632  ( .A(\SUBBYTES[8].a/w3365 ), .B(
        \SUBBYTES[8].a/w3368 ), .Z(n14833) );
  XOR \SUBBYTES[8].a/U5630  ( .A(\SUBBYTES[8].a/w3353 ), .B(n15868), .Z(n14834) );
  XOR \SUBBYTES[8].a/U5628  ( .A(\SUBBYTES[8].a/w3385 ), .B(
        \SUBBYTES[8].a/w3398 ), .Z(n14835) );
  XOR \SUBBYTES[8].a/U5626  ( .A(n14839), .B(n14838), .Z(n14836) );
  XOR \SUBBYTES[8].a/U5625  ( .A(n14841), .B(n14840), .Z(n14837) );
  XOR \SUBBYTES[8].a/U5624  ( .A(\SUBBYTES[8].a/w3397 ), .B(
        \SUBBYTES[8].a/w3400 ), .Z(n14838) );
  XOR \SUBBYTES[8].a/U5623  ( .A(\SUBBYTES[8].a/w3390 ), .B(
        \SUBBYTES[8].a/w3393 ), .Z(n14839) );
  XOR \SUBBYTES[8].a/U5622  ( .A(\SUBBYTES[8].a/w3365 ), .B(
        \SUBBYTES[8].a/w3366 ), .Z(n14840) );
  XOR \SUBBYTES[8].a/U5621  ( .A(\SUBBYTES[8].a/w3350 ), .B(
        \SUBBYTES[8].a/w3353 ), .Z(n14841) );
  XOR \SUBBYTES[8].a/U5619  ( .A(n15865), .B(n14844), .Z(n14842) );
  XOR \SUBBYTES[8].a/U5618  ( .A(n15867), .B(n15866), .Z(n14843) );
  XOR \SUBBYTES[8].a/U5617  ( .A(\SUBBYTES[8].a/w3358 ), .B(
        \SUBBYTES[8].a/w3385 ), .Z(n14844) );
  XOR \SUBBYTES[8].a/U5615  ( .A(n15868), .B(n14847), .Z(n14845) );
  XOR \SUBBYTES[8].a/U5614  ( .A(\SUBBYTES[8].a/w3391 ), .B(
        \SUBBYTES[8].a/w3393 ), .Z(n14846) );
  XOR \SUBBYTES[8].a/U5613  ( .A(\SUBBYTES[8].a/w3351 ), .B(
        \SUBBYTES[8].a/w3383 ), .Z(n14847) );
  XOR \SUBBYTES[8].a/U5612  ( .A(\SUBBYTES[8].a/w3183 ), .B(
        \SUBBYTES[8].a/w3184 ), .Z(n15870) );
  XOR \SUBBYTES[8].a/U5611  ( .A(n15870), .B(n14848), .Z(n15869) );
  XOR \SUBBYTES[8].a/U5610  ( .A(\SUBBYTES[8].a/w3176 ), .B(
        \SUBBYTES[8].a/w3193 ), .Z(n14848) );
  XOR \SUBBYTES[8].a/U5608  ( .A(\SUBBYTES[8].a/w3175 ), .B(
        \SUBBYTES[8].a/w3190 ), .Z(n14849) );
  XOR \SUBBYTES[8].a/U5607  ( .A(n15870), .B(n14850), .Z(n16057) );
  XOR \SUBBYTES[8].a/U5606  ( .A(\SUBBYTES[8].a/w3190 ), .B(
        \SUBBYTES[8].a/w3191 ), .Z(n14850) );
  XOR \SUBBYTES[8].a/U5605  ( .A(\SUBBYTES[8].a/w3152 ), .B(n14851), .Z(n15872) );
  XOR \SUBBYTES[8].a/U5604  ( .A(\SUBBYTES[8].a/w3143 ), .B(
        \SUBBYTES[8].a/w3144 ), .Z(n14851) );
  XOR \SUBBYTES[8].a/U5602  ( .A(\SUBBYTES[8].a/w3154 ), .B(n16057), .Z(n14852) );
  XOR \SUBBYTES[8].a/U5601  ( .A(n14854), .B(n14853), .Z(n15873) );
  XOR \SUBBYTES[8].a/U5600  ( .A(n14856), .B(n14855), .Z(n14853) );
  XOR \SUBBYTES[8].a/U5599  ( .A(\SUBBYTES[8].a/w3190 ), .B(
        \SUBBYTES[8].a/w3191 ), .Z(n14854) );
  XOR \SUBBYTES[8].a/U5598  ( .A(\SUBBYTES[8].a/w3154 ), .B(
        \SUBBYTES[8].a/w3178 ), .Z(n14855) );
  XOR \SUBBYTES[8].a/U5597  ( .A(\SUBBYTES[8].a/w3143 ), .B(
        \SUBBYTES[8].a/w3152 ), .Z(n14856) );
  XOR \SUBBYTES[8].a/U5596  ( .A(\SUBBYTES[8].a/w3175 ), .B(n14857), .Z(n15871) );
  XOR \SUBBYTES[8].a/U5595  ( .A(\SUBBYTES[8].a/w3158 ), .B(
        \SUBBYTES[8].a/w3161 ), .Z(n14857) );
  XOR \SUBBYTES[8].a/U5593  ( .A(\SUBBYTES[8].a/w3146 ), .B(n15873), .Z(n14858) );
  XOR \SUBBYTES[8].a/U5591  ( .A(\SUBBYTES[8].a/w3178 ), .B(
        \SUBBYTES[8].a/w3191 ), .Z(n14859) );
  XOR \SUBBYTES[8].a/U5589  ( .A(n14863), .B(n14862), .Z(n14860) );
  XOR \SUBBYTES[8].a/U5588  ( .A(n14865), .B(n14864), .Z(n14861) );
  XOR \SUBBYTES[8].a/U5587  ( .A(\SUBBYTES[8].a/w3190 ), .B(
        \SUBBYTES[8].a/w3193 ), .Z(n14862) );
  XOR \SUBBYTES[8].a/U5586  ( .A(\SUBBYTES[8].a/w3183 ), .B(
        \SUBBYTES[8].a/w3186 ), .Z(n14863) );
  XOR \SUBBYTES[8].a/U5585  ( .A(\SUBBYTES[8].a/w3158 ), .B(
        \SUBBYTES[8].a/w3159 ), .Z(n14864) );
  XOR \SUBBYTES[8].a/U5584  ( .A(\SUBBYTES[8].a/w3143 ), .B(
        \SUBBYTES[8].a/w3146 ), .Z(n14865) );
  XOR \SUBBYTES[8].a/U5582  ( .A(n15870), .B(n14868), .Z(n14866) );
  XOR \SUBBYTES[8].a/U5581  ( .A(n15872), .B(n15871), .Z(n14867) );
  XOR \SUBBYTES[8].a/U5580  ( .A(\SUBBYTES[8].a/w3151 ), .B(
        \SUBBYTES[8].a/w3178 ), .Z(n14868) );
  XOR \SUBBYTES[8].a/U5578  ( .A(n15873), .B(n14871), .Z(n14869) );
  XOR \SUBBYTES[8].a/U5577  ( .A(\SUBBYTES[8].a/w3184 ), .B(
        \SUBBYTES[8].a/w3186 ), .Z(n14870) );
  XOR \SUBBYTES[8].a/U5576  ( .A(\SUBBYTES[8].a/w3144 ), .B(
        \SUBBYTES[8].a/w3176 ), .Z(n14871) );
  XOR \SUBBYTES[8].a/U5575  ( .A(\SUBBYTES[8].a/w2976 ), .B(
        \SUBBYTES[8].a/w2977 ), .Z(n15875) );
  XOR \SUBBYTES[8].a/U5574  ( .A(n15875), .B(n14872), .Z(n15874) );
  XOR \SUBBYTES[8].a/U5573  ( .A(\SUBBYTES[8].a/w2969 ), .B(
        \SUBBYTES[8].a/w2986 ), .Z(n14872) );
  XOR \SUBBYTES[8].a/U5571  ( .A(\SUBBYTES[8].a/w2968 ), .B(
        \SUBBYTES[8].a/w2983 ), .Z(n14873) );
  XOR \SUBBYTES[8].a/U5570  ( .A(n15875), .B(n14874), .Z(n16058) );
  XOR \SUBBYTES[8].a/U5569  ( .A(\SUBBYTES[8].a/w2983 ), .B(
        \SUBBYTES[8].a/w2984 ), .Z(n14874) );
  XOR \SUBBYTES[8].a/U5568  ( .A(\SUBBYTES[8].a/w2945 ), .B(n14875), .Z(n15877) );
  XOR \SUBBYTES[8].a/U5567  ( .A(\SUBBYTES[8].a/w2936 ), .B(
        \SUBBYTES[8].a/w2937 ), .Z(n14875) );
  XOR \SUBBYTES[8].a/U5565  ( .A(\SUBBYTES[8].a/w2947 ), .B(n16058), .Z(n14876) );
  XOR \SUBBYTES[8].a/U5564  ( .A(n14878), .B(n14877), .Z(n15878) );
  XOR \SUBBYTES[8].a/U5563  ( .A(n14880), .B(n14879), .Z(n14877) );
  XOR \SUBBYTES[8].a/U5562  ( .A(\SUBBYTES[8].a/w2983 ), .B(
        \SUBBYTES[8].a/w2984 ), .Z(n14878) );
  XOR \SUBBYTES[8].a/U5561  ( .A(\SUBBYTES[8].a/w2947 ), .B(
        \SUBBYTES[8].a/w2971 ), .Z(n14879) );
  XOR \SUBBYTES[8].a/U5560  ( .A(\SUBBYTES[8].a/w2936 ), .B(
        \SUBBYTES[8].a/w2945 ), .Z(n14880) );
  XOR \SUBBYTES[8].a/U5559  ( .A(\SUBBYTES[8].a/w2968 ), .B(n14881), .Z(n15876) );
  XOR \SUBBYTES[8].a/U5558  ( .A(\SUBBYTES[8].a/w2951 ), .B(
        \SUBBYTES[8].a/w2954 ), .Z(n14881) );
  XOR \SUBBYTES[8].a/U5556  ( .A(\SUBBYTES[8].a/w2939 ), .B(n15878), .Z(n14882) );
  XOR \SUBBYTES[8].a/U5554  ( .A(\SUBBYTES[8].a/w2971 ), .B(
        \SUBBYTES[8].a/w2984 ), .Z(n14883) );
  XOR \SUBBYTES[8].a/U5552  ( .A(n14887), .B(n14886), .Z(n14884) );
  XOR \SUBBYTES[8].a/U5551  ( .A(n14889), .B(n14888), .Z(n14885) );
  XOR \SUBBYTES[8].a/U5550  ( .A(\SUBBYTES[8].a/w2983 ), .B(
        \SUBBYTES[8].a/w2986 ), .Z(n14886) );
  XOR \SUBBYTES[8].a/U5549  ( .A(\SUBBYTES[8].a/w2976 ), .B(
        \SUBBYTES[8].a/w2979 ), .Z(n14887) );
  XOR \SUBBYTES[8].a/U5548  ( .A(\SUBBYTES[8].a/w2951 ), .B(
        \SUBBYTES[8].a/w2952 ), .Z(n14888) );
  XOR \SUBBYTES[8].a/U5547  ( .A(\SUBBYTES[8].a/w2936 ), .B(
        \SUBBYTES[8].a/w2939 ), .Z(n14889) );
  XOR \SUBBYTES[8].a/U5545  ( .A(n15875), .B(n14892), .Z(n14890) );
  XOR \SUBBYTES[8].a/U5544  ( .A(n15877), .B(n15876), .Z(n14891) );
  XOR \SUBBYTES[8].a/U5543  ( .A(\SUBBYTES[8].a/w2944 ), .B(
        \SUBBYTES[8].a/w2971 ), .Z(n14892) );
  XOR \SUBBYTES[8].a/U5541  ( .A(n15878), .B(n14895), .Z(n14893) );
  XOR \SUBBYTES[8].a/U5540  ( .A(\SUBBYTES[8].a/w2977 ), .B(
        \SUBBYTES[8].a/w2979 ), .Z(n14894) );
  XOR \SUBBYTES[8].a/U5539  ( .A(\SUBBYTES[8].a/w2937 ), .B(
        \SUBBYTES[8].a/w2969 ), .Z(n14895) );
  XOR \SUBBYTES[8].a/U5538  ( .A(\SUBBYTES[8].a/w2769 ), .B(
        \SUBBYTES[8].a/w2770 ), .Z(n15880) );
  XOR \SUBBYTES[8].a/U5537  ( .A(n15880), .B(n14896), .Z(n15879) );
  XOR \SUBBYTES[8].a/U5536  ( .A(\SUBBYTES[8].a/w2762 ), .B(
        \SUBBYTES[8].a/w2779 ), .Z(n14896) );
  XOR \SUBBYTES[8].a/U5534  ( .A(\SUBBYTES[8].a/w2761 ), .B(
        \SUBBYTES[8].a/w2776 ), .Z(n14897) );
  XOR \SUBBYTES[8].a/U5533  ( .A(n15880), .B(n14898), .Z(n16059) );
  XOR \SUBBYTES[8].a/U5532  ( .A(\SUBBYTES[8].a/w2776 ), .B(
        \SUBBYTES[8].a/w2777 ), .Z(n14898) );
  XOR \SUBBYTES[8].a/U5531  ( .A(\SUBBYTES[8].a/w2738 ), .B(n14899), .Z(n15882) );
  XOR \SUBBYTES[8].a/U5530  ( .A(\SUBBYTES[8].a/w2729 ), .B(
        \SUBBYTES[8].a/w2730 ), .Z(n14899) );
  XOR \SUBBYTES[8].a/U5528  ( .A(\SUBBYTES[8].a/w2740 ), .B(n16059), .Z(n14900) );
  XOR \SUBBYTES[8].a/U5527  ( .A(n14902), .B(n14901), .Z(n15883) );
  XOR \SUBBYTES[8].a/U5526  ( .A(n14904), .B(n14903), .Z(n14901) );
  XOR \SUBBYTES[8].a/U5525  ( .A(\SUBBYTES[8].a/w2776 ), .B(
        \SUBBYTES[8].a/w2777 ), .Z(n14902) );
  XOR \SUBBYTES[8].a/U5524  ( .A(\SUBBYTES[8].a/w2740 ), .B(
        \SUBBYTES[8].a/w2764 ), .Z(n14903) );
  XOR \SUBBYTES[8].a/U5523  ( .A(\SUBBYTES[8].a/w2729 ), .B(
        \SUBBYTES[8].a/w2738 ), .Z(n14904) );
  XOR \SUBBYTES[8].a/U5522  ( .A(\SUBBYTES[8].a/w2761 ), .B(n14905), .Z(n15881) );
  XOR \SUBBYTES[8].a/U5521  ( .A(\SUBBYTES[8].a/w2744 ), .B(
        \SUBBYTES[8].a/w2747 ), .Z(n14905) );
  XOR \SUBBYTES[8].a/U5519  ( .A(\SUBBYTES[8].a/w2732 ), .B(n15883), .Z(n14906) );
  XOR \SUBBYTES[8].a/U5517  ( .A(\SUBBYTES[8].a/w2764 ), .B(
        \SUBBYTES[8].a/w2777 ), .Z(n14907) );
  XOR \SUBBYTES[8].a/U5515  ( .A(n14911), .B(n14910), .Z(n14908) );
  XOR \SUBBYTES[8].a/U5514  ( .A(n14913), .B(n14912), .Z(n14909) );
  XOR \SUBBYTES[8].a/U5513  ( .A(\SUBBYTES[8].a/w2776 ), .B(
        \SUBBYTES[8].a/w2779 ), .Z(n14910) );
  XOR \SUBBYTES[8].a/U5512  ( .A(\SUBBYTES[8].a/w2769 ), .B(
        \SUBBYTES[8].a/w2772 ), .Z(n14911) );
  XOR \SUBBYTES[8].a/U5511  ( .A(\SUBBYTES[8].a/w2744 ), .B(
        \SUBBYTES[8].a/w2745 ), .Z(n14912) );
  XOR \SUBBYTES[8].a/U5510  ( .A(\SUBBYTES[8].a/w2729 ), .B(
        \SUBBYTES[8].a/w2732 ), .Z(n14913) );
  XOR \SUBBYTES[8].a/U5508  ( .A(n15880), .B(n14916), .Z(n14914) );
  XOR \SUBBYTES[8].a/U5507  ( .A(n15882), .B(n15881), .Z(n14915) );
  XOR \SUBBYTES[8].a/U5506  ( .A(\SUBBYTES[8].a/w2737 ), .B(
        \SUBBYTES[8].a/w2764 ), .Z(n14916) );
  XOR \SUBBYTES[8].a/U5504  ( .A(n15883), .B(n14919), .Z(n14917) );
  XOR \SUBBYTES[8].a/U5503  ( .A(\SUBBYTES[8].a/w2770 ), .B(
        \SUBBYTES[8].a/w2772 ), .Z(n14918) );
  XOR \SUBBYTES[8].a/U5502  ( .A(\SUBBYTES[8].a/w2730 ), .B(
        \SUBBYTES[8].a/w2762 ), .Z(n14919) );
  XOR \SUBBYTES[8].a/U5501  ( .A(\SUBBYTES[8].a/w2562 ), .B(
        \SUBBYTES[8].a/w2563 ), .Z(n15885) );
  XOR \SUBBYTES[8].a/U5500  ( .A(n15885), .B(n14920), .Z(n15884) );
  XOR \SUBBYTES[8].a/U5499  ( .A(\SUBBYTES[8].a/w2555 ), .B(
        \SUBBYTES[8].a/w2572 ), .Z(n14920) );
  XOR \SUBBYTES[8].a/U5497  ( .A(\SUBBYTES[8].a/w2554 ), .B(
        \SUBBYTES[8].a/w2569 ), .Z(n14921) );
  XOR \SUBBYTES[8].a/U5496  ( .A(n15885), .B(n14922), .Z(n16060) );
  XOR \SUBBYTES[8].a/U5495  ( .A(\SUBBYTES[8].a/w2569 ), .B(
        \SUBBYTES[8].a/w2570 ), .Z(n14922) );
  XOR \SUBBYTES[8].a/U5494  ( .A(\SUBBYTES[8].a/w2531 ), .B(n14923), .Z(n15887) );
  XOR \SUBBYTES[8].a/U5493  ( .A(\SUBBYTES[8].a/w2522 ), .B(
        \SUBBYTES[8].a/w2523 ), .Z(n14923) );
  XOR \SUBBYTES[8].a/U5491  ( .A(\SUBBYTES[8].a/w2533 ), .B(n16060), .Z(n14924) );
  XOR \SUBBYTES[8].a/U5490  ( .A(n14926), .B(n14925), .Z(n15888) );
  XOR \SUBBYTES[8].a/U5489  ( .A(n14928), .B(n14927), .Z(n14925) );
  XOR \SUBBYTES[8].a/U5488  ( .A(\SUBBYTES[8].a/w2569 ), .B(
        \SUBBYTES[8].a/w2570 ), .Z(n14926) );
  XOR \SUBBYTES[8].a/U5487  ( .A(\SUBBYTES[8].a/w2533 ), .B(
        \SUBBYTES[8].a/w2557 ), .Z(n14927) );
  XOR \SUBBYTES[8].a/U5486  ( .A(\SUBBYTES[8].a/w2522 ), .B(
        \SUBBYTES[8].a/w2531 ), .Z(n14928) );
  XOR \SUBBYTES[8].a/U5485  ( .A(\SUBBYTES[8].a/w2554 ), .B(n14929), .Z(n15886) );
  XOR \SUBBYTES[8].a/U5484  ( .A(\SUBBYTES[8].a/w2537 ), .B(
        \SUBBYTES[8].a/w2540 ), .Z(n14929) );
  XOR \SUBBYTES[8].a/U5482  ( .A(\SUBBYTES[8].a/w2525 ), .B(n15888), .Z(n14930) );
  XOR \SUBBYTES[8].a/U5480  ( .A(\SUBBYTES[8].a/w2557 ), .B(
        \SUBBYTES[8].a/w2570 ), .Z(n14931) );
  XOR \SUBBYTES[8].a/U5478  ( .A(n14935), .B(n14934), .Z(n14932) );
  XOR \SUBBYTES[8].a/U5477  ( .A(n14937), .B(n14936), .Z(n14933) );
  XOR \SUBBYTES[8].a/U5476  ( .A(\SUBBYTES[8].a/w2569 ), .B(
        \SUBBYTES[8].a/w2572 ), .Z(n14934) );
  XOR \SUBBYTES[8].a/U5475  ( .A(\SUBBYTES[8].a/w2562 ), .B(
        \SUBBYTES[8].a/w2565 ), .Z(n14935) );
  XOR \SUBBYTES[8].a/U5474  ( .A(\SUBBYTES[8].a/w2537 ), .B(
        \SUBBYTES[8].a/w2538 ), .Z(n14936) );
  XOR \SUBBYTES[8].a/U5473  ( .A(\SUBBYTES[8].a/w2522 ), .B(
        \SUBBYTES[8].a/w2525 ), .Z(n14937) );
  XOR \SUBBYTES[8].a/U5471  ( .A(n15885), .B(n14940), .Z(n14938) );
  XOR \SUBBYTES[8].a/U5470  ( .A(n15887), .B(n15886), .Z(n14939) );
  XOR \SUBBYTES[8].a/U5469  ( .A(\SUBBYTES[8].a/w2530 ), .B(
        \SUBBYTES[8].a/w2557 ), .Z(n14940) );
  XOR \SUBBYTES[8].a/U5467  ( .A(n15888), .B(n14943), .Z(n14941) );
  XOR \SUBBYTES[8].a/U5466  ( .A(\SUBBYTES[8].a/w2563 ), .B(
        \SUBBYTES[8].a/w2565 ), .Z(n14942) );
  XOR \SUBBYTES[8].a/U5465  ( .A(\SUBBYTES[8].a/w2523 ), .B(
        \SUBBYTES[8].a/w2555 ), .Z(n14943) );
  XOR \SUBBYTES[8].a/U5464  ( .A(\SUBBYTES[8].a/w2355 ), .B(
        \SUBBYTES[8].a/w2356 ), .Z(n15890) );
  XOR \SUBBYTES[8].a/U5463  ( .A(n15890), .B(n14944), .Z(n15889) );
  XOR \SUBBYTES[8].a/U5462  ( .A(\SUBBYTES[8].a/w2348 ), .B(
        \SUBBYTES[8].a/w2365 ), .Z(n14944) );
  XOR \SUBBYTES[8].a/U5460  ( .A(\SUBBYTES[8].a/w2347 ), .B(
        \SUBBYTES[8].a/w2362 ), .Z(n14945) );
  XOR \SUBBYTES[8].a/U5459  ( .A(n15890), .B(n14946), .Z(n16061) );
  XOR \SUBBYTES[8].a/U5458  ( .A(\SUBBYTES[8].a/w2362 ), .B(
        \SUBBYTES[8].a/w2363 ), .Z(n14946) );
  XOR \SUBBYTES[8].a/U5457  ( .A(\SUBBYTES[8].a/w2324 ), .B(n14947), .Z(n15892) );
  XOR \SUBBYTES[8].a/U5456  ( .A(\SUBBYTES[8].a/w2315 ), .B(
        \SUBBYTES[8].a/w2316 ), .Z(n14947) );
  XOR \SUBBYTES[8].a/U5454  ( .A(\SUBBYTES[8].a/w2326 ), .B(n16061), .Z(n14948) );
  XOR \SUBBYTES[8].a/U5453  ( .A(n14950), .B(n14949), .Z(n15893) );
  XOR \SUBBYTES[8].a/U5452  ( .A(n14952), .B(n14951), .Z(n14949) );
  XOR \SUBBYTES[8].a/U5451  ( .A(\SUBBYTES[8].a/w2362 ), .B(
        \SUBBYTES[8].a/w2363 ), .Z(n14950) );
  XOR \SUBBYTES[8].a/U5450  ( .A(\SUBBYTES[8].a/w2326 ), .B(
        \SUBBYTES[8].a/w2350 ), .Z(n14951) );
  XOR \SUBBYTES[8].a/U5449  ( .A(\SUBBYTES[8].a/w2315 ), .B(
        \SUBBYTES[8].a/w2324 ), .Z(n14952) );
  XOR \SUBBYTES[8].a/U5448  ( .A(\SUBBYTES[8].a/w2347 ), .B(n14953), .Z(n15891) );
  XOR \SUBBYTES[8].a/U5447  ( .A(\SUBBYTES[8].a/w2330 ), .B(
        \SUBBYTES[8].a/w2333 ), .Z(n14953) );
  XOR \SUBBYTES[8].a/U5445  ( .A(\SUBBYTES[8].a/w2318 ), .B(n15893), .Z(n14954) );
  XOR \SUBBYTES[8].a/U5443  ( .A(\SUBBYTES[8].a/w2350 ), .B(
        \SUBBYTES[8].a/w2363 ), .Z(n14955) );
  XOR \SUBBYTES[8].a/U5441  ( .A(n14959), .B(n14958), .Z(n14956) );
  XOR \SUBBYTES[8].a/U5440  ( .A(n14961), .B(n14960), .Z(n14957) );
  XOR \SUBBYTES[8].a/U5439  ( .A(\SUBBYTES[8].a/w2362 ), .B(
        \SUBBYTES[8].a/w2365 ), .Z(n14958) );
  XOR \SUBBYTES[8].a/U5438  ( .A(\SUBBYTES[8].a/w2355 ), .B(
        \SUBBYTES[8].a/w2358 ), .Z(n14959) );
  XOR \SUBBYTES[8].a/U5437  ( .A(\SUBBYTES[8].a/w2330 ), .B(
        \SUBBYTES[8].a/w2331 ), .Z(n14960) );
  XOR \SUBBYTES[8].a/U5436  ( .A(\SUBBYTES[8].a/w2315 ), .B(
        \SUBBYTES[8].a/w2318 ), .Z(n14961) );
  XOR \SUBBYTES[8].a/U5434  ( .A(n15890), .B(n14964), .Z(n14962) );
  XOR \SUBBYTES[8].a/U5433  ( .A(n15892), .B(n15891), .Z(n14963) );
  XOR \SUBBYTES[8].a/U5432  ( .A(\SUBBYTES[8].a/w2323 ), .B(
        \SUBBYTES[8].a/w2350 ), .Z(n14964) );
  XOR \SUBBYTES[8].a/U5430  ( .A(n15893), .B(n14967), .Z(n14965) );
  XOR \SUBBYTES[8].a/U5429  ( .A(\SUBBYTES[8].a/w2356 ), .B(
        \SUBBYTES[8].a/w2358 ), .Z(n14966) );
  XOR \SUBBYTES[8].a/U5428  ( .A(\SUBBYTES[8].a/w2316 ), .B(
        \SUBBYTES[8].a/w2348 ), .Z(n14967) );
  XOR \SUBBYTES[8].a/U5427  ( .A(\SUBBYTES[8].a/w2148 ), .B(
        \SUBBYTES[8].a/w2149 ), .Z(n15895) );
  XOR \SUBBYTES[8].a/U5426  ( .A(n15895), .B(n14968), .Z(n15894) );
  XOR \SUBBYTES[8].a/U5425  ( .A(\SUBBYTES[8].a/w2141 ), .B(
        \SUBBYTES[8].a/w2158 ), .Z(n14968) );
  XOR \SUBBYTES[8].a/U5423  ( .A(\SUBBYTES[8].a/w2140 ), .B(
        \SUBBYTES[8].a/w2155 ), .Z(n14969) );
  XOR \SUBBYTES[8].a/U5422  ( .A(n15895), .B(n14970), .Z(n16062) );
  XOR \SUBBYTES[8].a/U5421  ( .A(\SUBBYTES[8].a/w2155 ), .B(
        \SUBBYTES[8].a/w2156 ), .Z(n14970) );
  XOR \SUBBYTES[8].a/U5420  ( .A(\SUBBYTES[8].a/w2117 ), .B(n14971), .Z(n15897) );
  XOR \SUBBYTES[8].a/U5419  ( .A(\SUBBYTES[8].a/w2108 ), .B(
        \SUBBYTES[8].a/w2109 ), .Z(n14971) );
  XOR \SUBBYTES[8].a/U5417  ( .A(\SUBBYTES[8].a/w2119 ), .B(n16062), .Z(n14972) );
  XOR \SUBBYTES[8].a/U5416  ( .A(n14974), .B(n14973), .Z(n15898) );
  XOR \SUBBYTES[8].a/U5415  ( .A(n14976), .B(n14975), .Z(n14973) );
  XOR \SUBBYTES[8].a/U5414  ( .A(\SUBBYTES[8].a/w2155 ), .B(
        \SUBBYTES[8].a/w2156 ), .Z(n14974) );
  XOR \SUBBYTES[8].a/U5413  ( .A(\SUBBYTES[8].a/w2119 ), .B(
        \SUBBYTES[8].a/w2143 ), .Z(n14975) );
  XOR \SUBBYTES[8].a/U5412  ( .A(\SUBBYTES[8].a/w2108 ), .B(
        \SUBBYTES[8].a/w2117 ), .Z(n14976) );
  XOR \SUBBYTES[8].a/U5411  ( .A(\SUBBYTES[8].a/w2140 ), .B(n14977), .Z(n15896) );
  XOR \SUBBYTES[8].a/U5410  ( .A(\SUBBYTES[8].a/w2123 ), .B(
        \SUBBYTES[8].a/w2126 ), .Z(n14977) );
  XOR \SUBBYTES[8].a/U5408  ( .A(\SUBBYTES[8].a/w2111 ), .B(n15898), .Z(n14978) );
  XOR \SUBBYTES[8].a/U5406  ( .A(\SUBBYTES[8].a/w2143 ), .B(
        \SUBBYTES[8].a/w2156 ), .Z(n14979) );
  XOR \SUBBYTES[8].a/U5404  ( .A(n14983), .B(n14982), .Z(n14980) );
  XOR \SUBBYTES[8].a/U5403  ( .A(n14985), .B(n14984), .Z(n14981) );
  XOR \SUBBYTES[8].a/U5402  ( .A(\SUBBYTES[8].a/w2155 ), .B(
        \SUBBYTES[8].a/w2158 ), .Z(n14982) );
  XOR \SUBBYTES[8].a/U5401  ( .A(\SUBBYTES[8].a/w2148 ), .B(
        \SUBBYTES[8].a/w2151 ), .Z(n14983) );
  XOR \SUBBYTES[8].a/U5400  ( .A(\SUBBYTES[8].a/w2123 ), .B(
        \SUBBYTES[8].a/w2124 ), .Z(n14984) );
  XOR \SUBBYTES[8].a/U5399  ( .A(\SUBBYTES[8].a/w2108 ), .B(
        \SUBBYTES[8].a/w2111 ), .Z(n14985) );
  XOR \SUBBYTES[8].a/U5397  ( .A(n15895), .B(n14988), .Z(n14986) );
  XOR \SUBBYTES[8].a/U5396  ( .A(n15897), .B(n15896), .Z(n14987) );
  XOR \SUBBYTES[8].a/U5395  ( .A(\SUBBYTES[8].a/w2116 ), .B(
        \SUBBYTES[8].a/w2143 ), .Z(n14988) );
  XOR \SUBBYTES[8].a/U5393  ( .A(n15898), .B(n14991), .Z(n14989) );
  XOR \SUBBYTES[8].a/U5392  ( .A(\SUBBYTES[8].a/w2149 ), .B(
        \SUBBYTES[8].a/w2151 ), .Z(n14990) );
  XOR \SUBBYTES[8].a/U5391  ( .A(\SUBBYTES[8].a/w2109 ), .B(
        \SUBBYTES[8].a/w2141 ), .Z(n14991) );
  XOR \SUBBYTES[8].a/U5390  ( .A(\SUBBYTES[8].a/w1941 ), .B(
        \SUBBYTES[8].a/w1942 ), .Z(n15900) );
  XOR \SUBBYTES[8].a/U5389  ( .A(n15900), .B(n14992), .Z(n15899) );
  XOR \SUBBYTES[8].a/U5388  ( .A(\SUBBYTES[8].a/w1934 ), .B(
        \SUBBYTES[8].a/w1951 ), .Z(n14992) );
  XOR \SUBBYTES[8].a/U5386  ( .A(\SUBBYTES[8].a/w1933 ), .B(
        \SUBBYTES[8].a/w1948 ), .Z(n14993) );
  XOR \SUBBYTES[8].a/U5385  ( .A(n15900), .B(n14994), .Z(n16063) );
  XOR \SUBBYTES[8].a/U5384  ( .A(\SUBBYTES[8].a/w1948 ), .B(
        \SUBBYTES[8].a/w1949 ), .Z(n14994) );
  XOR \SUBBYTES[8].a/U5383  ( .A(\SUBBYTES[8].a/w1910 ), .B(n14995), .Z(n15902) );
  XOR \SUBBYTES[8].a/U5382  ( .A(\SUBBYTES[8].a/w1901 ), .B(
        \SUBBYTES[8].a/w1902 ), .Z(n14995) );
  XOR \SUBBYTES[8].a/U5380  ( .A(\SUBBYTES[8].a/w1912 ), .B(n16063), .Z(n14996) );
  XOR \SUBBYTES[8].a/U5379  ( .A(n14998), .B(n14997), .Z(n15903) );
  XOR \SUBBYTES[8].a/U5378  ( .A(n15000), .B(n14999), .Z(n14997) );
  XOR \SUBBYTES[8].a/U5377  ( .A(\SUBBYTES[8].a/w1948 ), .B(
        \SUBBYTES[8].a/w1949 ), .Z(n14998) );
  XOR \SUBBYTES[8].a/U5376  ( .A(\SUBBYTES[8].a/w1912 ), .B(
        \SUBBYTES[8].a/w1936 ), .Z(n14999) );
  XOR \SUBBYTES[8].a/U5375  ( .A(\SUBBYTES[8].a/w1901 ), .B(
        \SUBBYTES[8].a/w1910 ), .Z(n15000) );
  XOR \SUBBYTES[8].a/U5374  ( .A(\SUBBYTES[8].a/w1933 ), .B(n15001), .Z(n15901) );
  XOR \SUBBYTES[8].a/U5373  ( .A(\SUBBYTES[8].a/w1916 ), .B(
        \SUBBYTES[8].a/w1919 ), .Z(n15001) );
  XOR \SUBBYTES[8].a/U5371  ( .A(\SUBBYTES[8].a/w1904 ), .B(n15903), .Z(n15002) );
  XOR \SUBBYTES[8].a/U5369  ( .A(\SUBBYTES[8].a/w1936 ), .B(
        \SUBBYTES[8].a/w1949 ), .Z(n15003) );
  XOR \SUBBYTES[8].a/U5367  ( .A(n15007), .B(n15006), .Z(n15004) );
  XOR \SUBBYTES[8].a/U5366  ( .A(n15009), .B(n15008), .Z(n15005) );
  XOR \SUBBYTES[8].a/U5365  ( .A(\SUBBYTES[8].a/w1948 ), .B(
        \SUBBYTES[8].a/w1951 ), .Z(n15006) );
  XOR \SUBBYTES[8].a/U5364  ( .A(\SUBBYTES[8].a/w1941 ), .B(
        \SUBBYTES[8].a/w1944 ), .Z(n15007) );
  XOR \SUBBYTES[8].a/U5363  ( .A(\SUBBYTES[8].a/w1916 ), .B(
        \SUBBYTES[8].a/w1917 ), .Z(n15008) );
  XOR \SUBBYTES[8].a/U5362  ( .A(\SUBBYTES[8].a/w1901 ), .B(
        \SUBBYTES[8].a/w1904 ), .Z(n15009) );
  XOR \SUBBYTES[8].a/U5360  ( .A(n15900), .B(n15012), .Z(n15010) );
  XOR \SUBBYTES[8].a/U5359  ( .A(n15902), .B(n15901), .Z(n15011) );
  XOR \SUBBYTES[8].a/U5358  ( .A(\SUBBYTES[8].a/w1909 ), .B(
        \SUBBYTES[8].a/w1936 ), .Z(n15012) );
  XOR \SUBBYTES[8].a/U5356  ( .A(n15903), .B(n15015), .Z(n15013) );
  XOR \SUBBYTES[8].a/U5355  ( .A(\SUBBYTES[8].a/w1942 ), .B(
        \SUBBYTES[8].a/w1944 ), .Z(n15014) );
  XOR \SUBBYTES[8].a/U5354  ( .A(\SUBBYTES[8].a/w1902 ), .B(
        \SUBBYTES[8].a/w1934 ), .Z(n15015) );
  XOR \SUBBYTES[8].a/U5353  ( .A(\SUBBYTES[8].a/w1734 ), .B(
        \SUBBYTES[8].a/w1735 ), .Z(n15905) );
  XOR \SUBBYTES[8].a/U5352  ( .A(n15905), .B(n15016), .Z(n15904) );
  XOR \SUBBYTES[8].a/U5351  ( .A(\SUBBYTES[8].a/w1727 ), .B(
        \SUBBYTES[8].a/w1744 ), .Z(n15016) );
  XOR \SUBBYTES[8].a/U5349  ( .A(\SUBBYTES[8].a/w1726 ), .B(
        \SUBBYTES[8].a/w1741 ), .Z(n15017) );
  XOR \SUBBYTES[8].a/U5348  ( .A(n15905), .B(n15018), .Z(n16064) );
  XOR \SUBBYTES[8].a/U5347  ( .A(\SUBBYTES[8].a/w1741 ), .B(
        \SUBBYTES[8].a/w1742 ), .Z(n15018) );
  XOR \SUBBYTES[8].a/U5346  ( .A(\SUBBYTES[8].a/w1703 ), .B(n15019), .Z(n15907) );
  XOR \SUBBYTES[8].a/U5345  ( .A(\SUBBYTES[8].a/w1694 ), .B(
        \SUBBYTES[8].a/w1695 ), .Z(n15019) );
  XOR \SUBBYTES[8].a/U5343  ( .A(\SUBBYTES[8].a/w1705 ), .B(n16064), .Z(n15020) );
  XOR \SUBBYTES[8].a/U5342  ( .A(n15022), .B(n15021), .Z(n15908) );
  XOR \SUBBYTES[8].a/U5341  ( .A(n15024), .B(n15023), .Z(n15021) );
  XOR \SUBBYTES[8].a/U5340  ( .A(\SUBBYTES[8].a/w1741 ), .B(
        \SUBBYTES[8].a/w1742 ), .Z(n15022) );
  XOR \SUBBYTES[8].a/U5339  ( .A(\SUBBYTES[8].a/w1705 ), .B(
        \SUBBYTES[8].a/w1729 ), .Z(n15023) );
  XOR \SUBBYTES[8].a/U5338  ( .A(\SUBBYTES[8].a/w1694 ), .B(
        \SUBBYTES[8].a/w1703 ), .Z(n15024) );
  XOR \SUBBYTES[8].a/U5337  ( .A(\SUBBYTES[8].a/w1726 ), .B(n15025), .Z(n15906) );
  XOR \SUBBYTES[8].a/U5336  ( .A(\SUBBYTES[8].a/w1709 ), .B(
        \SUBBYTES[8].a/w1712 ), .Z(n15025) );
  XOR \SUBBYTES[8].a/U5334  ( .A(\SUBBYTES[8].a/w1697 ), .B(n15908), .Z(n15026) );
  XOR \SUBBYTES[8].a/U5332  ( .A(\SUBBYTES[8].a/w1729 ), .B(
        \SUBBYTES[8].a/w1742 ), .Z(n15027) );
  XOR \SUBBYTES[8].a/U5330  ( .A(n15031), .B(n15030), .Z(n15028) );
  XOR \SUBBYTES[8].a/U5329  ( .A(n15033), .B(n15032), .Z(n15029) );
  XOR \SUBBYTES[8].a/U5328  ( .A(\SUBBYTES[8].a/w1741 ), .B(
        \SUBBYTES[8].a/w1744 ), .Z(n15030) );
  XOR \SUBBYTES[8].a/U5327  ( .A(\SUBBYTES[8].a/w1734 ), .B(
        \SUBBYTES[8].a/w1737 ), .Z(n15031) );
  XOR \SUBBYTES[8].a/U5326  ( .A(\SUBBYTES[8].a/w1709 ), .B(
        \SUBBYTES[8].a/w1710 ), .Z(n15032) );
  XOR \SUBBYTES[8].a/U5325  ( .A(\SUBBYTES[8].a/w1694 ), .B(
        \SUBBYTES[8].a/w1697 ), .Z(n15033) );
  XOR \SUBBYTES[8].a/U5323  ( .A(n15905), .B(n15036), .Z(n15034) );
  XOR \SUBBYTES[8].a/U5322  ( .A(n15907), .B(n15906), .Z(n15035) );
  XOR \SUBBYTES[8].a/U5321  ( .A(\SUBBYTES[8].a/w1702 ), .B(
        \SUBBYTES[8].a/w1729 ), .Z(n15036) );
  XOR \SUBBYTES[8].a/U5319  ( .A(n15908), .B(n15039), .Z(n15037) );
  XOR \SUBBYTES[8].a/U5318  ( .A(\SUBBYTES[8].a/w1735 ), .B(
        \SUBBYTES[8].a/w1737 ), .Z(n15038) );
  XOR \SUBBYTES[8].a/U5317  ( .A(\SUBBYTES[8].a/w1695 ), .B(
        \SUBBYTES[8].a/w1727 ), .Z(n15039) );
  XOR \SUBBYTES[8].a/U5316  ( .A(\SUBBYTES[8].a/w1527 ), .B(
        \SUBBYTES[8].a/w1528 ), .Z(n15910) );
  XOR \SUBBYTES[8].a/U5315  ( .A(n15910), .B(n15040), .Z(n15909) );
  XOR \SUBBYTES[8].a/U5314  ( .A(\SUBBYTES[8].a/w1520 ), .B(
        \SUBBYTES[8].a/w1537 ), .Z(n15040) );
  XOR \SUBBYTES[8].a/U5312  ( .A(\SUBBYTES[8].a/w1519 ), .B(
        \SUBBYTES[8].a/w1534 ), .Z(n15041) );
  XOR \SUBBYTES[8].a/U5311  ( .A(n15910), .B(n15042), .Z(n16065) );
  XOR \SUBBYTES[8].a/U5310  ( .A(\SUBBYTES[8].a/w1534 ), .B(
        \SUBBYTES[8].a/w1535 ), .Z(n15042) );
  XOR \SUBBYTES[8].a/U5309  ( .A(\SUBBYTES[8].a/w1496 ), .B(n15043), .Z(n15912) );
  XOR \SUBBYTES[8].a/U5308  ( .A(\SUBBYTES[8].a/w1487 ), .B(
        \SUBBYTES[8].a/w1488 ), .Z(n15043) );
  XOR \SUBBYTES[8].a/U5306  ( .A(\SUBBYTES[8].a/w1498 ), .B(n16065), .Z(n15044) );
  XOR \SUBBYTES[8].a/U5305  ( .A(n15046), .B(n15045), .Z(n15913) );
  XOR \SUBBYTES[8].a/U5304  ( .A(n15048), .B(n15047), .Z(n15045) );
  XOR \SUBBYTES[8].a/U5303  ( .A(\SUBBYTES[8].a/w1534 ), .B(
        \SUBBYTES[8].a/w1535 ), .Z(n15046) );
  XOR \SUBBYTES[8].a/U5302  ( .A(\SUBBYTES[8].a/w1498 ), .B(
        \SUBBYTES[8].a/w1522 ), .Z(n15047) );
  XOR \SUBBYTES[8].a/U5301  ( .A(\SUBBYTES[8].a/w1487 ), .B(
        \SUBBYTES[8].a/w1496 ), .Z(n15048) );
  XOR \SUBBYTES[8].a/U5300  ( .A(\SUBBYTES[8].a/w1519 ), .B(n15049), .Z(n15911) );
  XOR \SUBBYTES[8].a/U5299  ( .A(\SUBBYTES[8].a/w1502 ), .B(
        \SUBBYTES[8].a/w1505 ), .Z(n15049) );
  XOR \SUBBYTES[8].a/U5297  ( .A(\SUBBYTES[8].a/w1490 ), .B(n15913), .Z(n15050) );
  XOR \SUBBYTES[8].a/U5295  ( .A(\SUBBYTES[8].a/w1522 ), .B(
        \SUBBYTES[8].a/w1535 ), .Z(n15051) );
  XOR \SUBBYTES[8].a/U5293  ( .A(n15055), .B(n15054), .Z(n15052) );
  XOR \SUBBYTES[8].a/U5292  ( .A(n15057), .B(n15056), .Z(n15053) );
  XOR \SUBBYTES[8].a/U5291  ( .A(\SUBBYTES[8].a/w1534 ), .B(
        \SUBBYTES[8].a/w1537 ), .Z(n15054) );
  XOR \SUBBYTES[8].a/U5290  ( .A(\SUBBYTES[8].a/w1527 ), .B(
        \SUBBYTES[8].a/w1530 ), .Z(n15055) );
  XOR \SUBBYTES[8].a/U5289  ( .A(\SUBBYTES[8].a/w1502 ), .B(
        \SUBBYTES[8].a/w1503 ), .Z(n15056) );
  XOR \SUBBYTES[8].a/U5288  ( .A(\SUBBYTES[8].a/w1487 ), .B(
        \SUBBYTES[8].a/w1490 ), .Z(n15057) );
  XOR \SUBBYTES[8].a/U5286  ( .A(n15910), .B(n15060), .Z(n15058) );
  XOR \SUBBYTES[8].a/U5285  ( .A(n15912), .B(n15911), .Z(n15059) );
  XOR \SUBBYTES[8].a/U5284  ( .A(\SUBBYTES[8].a/w1495 ), .B(
        \SUBBYTES[8].a/w1522 ), .Z(n15060) );
  XOR \SUBBYTES[8].a/U5282  ( .A(n15913), .B(n15063), .Z(n15061) );
  XOR \SUBBYTES[8].a/U5281  ( .A(\SUBBYTES[8].a/w1528 ), .B(
        \SUBBYTES[8].a/w1530 ), .Z(n15062) );
  XOR \SUBBYTES[8].a/U5280  ( .A(\SUBBYTES[8].a/w1488 ), .B(
        \SUBBYTES[8].a/w1520 ), .Z(n15063) );
  XOR \SUBBYTES[8].a/U5279  ( .A(\SUBBYTES[8].a/w1320 ), .B(
        \SUBBYTES[8].a/w1321 ), .Z(n15915) );
  XOR \SUBBYTES[8].a/U5278  ( .A(n15915), .B(n15064), .Z(n15914) );
  XOR \SUBBYTES[8].a/U5277  ( .A(\SUBBYTES[8].a/w1313 ), .B(
        \SUBBYTES[8].a/w1330 ), .Z(n15064) );
  XOR \SUBBYTES[8].a/U5275  ( .A(\SUBBYTES[8].a/w1312 ), .B(
        \SUBBYTES[8].a/w1327 ), .Z(n15065) );
  XOR \SUBBYTES[8].a/U5274  ( .A(n15915), .B(n15066), .Z(n16066) );
  XOR \SUBBYTES[8].a/U5273  ( .A(\SUBBYTES[8].a/w1327 ), .B(
        \SUBBYTES[8].a/w1328 ), .Z(n15066) );
  XOR \SUBBYTES[8].a/U5272  ( .A(\SUBBYTES[8].a/w1289 ), .B(n15067), .Z(n15917) );
  XOR \SUBBYTES[8].a/U5271  ( .A(\SUBBYTES[8].a/w1280 ), .B(
        \SUBBYTES[8].a/w1281 ), .Z(n15067) );
  XOR \SUBBYTES[8].a/U5269  ( .A(\SUBBYTES[8].a/w1291 ), .B(n16066), .Z(n15068) );
  XOR \SUBBYTES[8].a/U5268  ( .A(n15070), .B(n15069), .Z(n15918) );
  XOR \SUBBYTES[8].a/U5267  ( .A(n15072), .B(n15071), .Z(n15069) );
  XOR \SUBBYTES[8].a/U5266  ( .A(\SUBBYTES[8].a/w1327 ), .B(
        \SUBBYTES[8].a/w1328 ), .Z(n15070) );
  XOR \SUBBYTES[8].a/U5265  ( .A(\SUBBYTES[8].a/w1291 ), .B(
        \SUBBYTES[8].a/w1315 ), .Z(n15071) );
  XOR \SUBBYTES[8].a/U5264  ( .A(\SUBBYTES[8].a/w1280 ), .B(
        \SUBBYTES[8].a/w1289 ), .Z(n15072) );
  XOR \SUBBYTES[8].a/U5263  ( .A(\SUBBYTES[8].a/w1312 ), .B(n15073), .Z(n15916) );
  XOR \SUBBYTES[8].a/U5262  ( .A(\SUBBYTES[8].a/w1295 ), .B(
        \SUBBYTES[8].a/w1298 ), .Z(n15073) );
  XOR \SUBBYTES[8].a/U5260  ( .A(\SUBBYTES[8].a/w1283 ), .B(n15918), .Z(n15074) );
  XOR \SUBBYTES[8].a/U5258  ( .A(\SUBBYTES[8].a/w1315 ), .B(
        \SUBBYTES[8].a/w1328 ), .Z(n15075) );
  XOR \SUBBYTES[8].a/U5256  ( .A(n15079), .B(n15078), .Z(n15076) );
  XOR \SUBBYTES[8].a/U5255  ( .A(n15081), .B(n15080), .Z(n15077) );
  XOR \SUBBYTES[8].a/U5254  ( .A(\SUBBYTES[8].a/w1327 ), .B(
        \SUBBYTES[8].a/w1330 ), .Z(n15078) );
  XOR \SUBBYTES[8].a/U5253  ( .A(\SUBBYTES[8].a/w1320 ), .B(
        \SUBBYTES[8].a/w1323 ), .Z(n15079) );
  XOR \SUBBYTES[8].a/U5252  ( .A(\SUBBYTES[8].a/w1295 ), .B(
        \SUBBYTES[8].a/w1296 ), .Z(n15080) );
  XOR \SUBBYTES[8].a/U5251  ( .A(\SUBBYTES[8].a/w1280 ), .B(
        \SUBBYTES[8].a/w1283 ), .Z(n15081) );
  XOR \SUBBYTES[8].a/U5249  ( .A(n15915), .B(n15084), .Z(n15082) );
  XOR \SUBBYTES[8].a/U5248  ( .A(n15917), .B(n15916), .Z(n15083) );
  XOR \SUBBYTES[8].a/U5247  ( .A(\SUBBYTES[8].a/w1288 ), .B(
        \SUBBYTES[8].a/w1315 ), .Z(n15084) );
  XOR \SUBBYTES[8].a/U5245  ( .A(n15918), .B(n15087), .Z(n15085) );
  XOR \SUBBYTES[8].a/U5244  ( .A(\SUBBYTES[8].a/w1321 ), .B(
        \SUBBYTES[8].a/w1323 ), .Z(n15086) );
  XOR \SUBBYTES[8].a/U5243  ( .A(\SUBBYTES[8].a/w1281 ), .B(
        \SUBBYTES[8].a/w1313 ), .Z(n15087) );
  XOR \SUBBYTES[8].a/U5242  ( .A(\SUBBYTES[8].a/w1113 ), .B(
        \SUBBYTES[8].a/w1114 ), .Z(n15920) );
  XOR \SUBBYTES[8].a/U5241  ( .A(n15920), .B(n15088), .Z(n15919) );
  XOR \SUBBYTES[8].a/U5240  ( .A(\SUBBYTES[8].a/w1106 ), .B(
        \SUBBYTES[8].a/w1123 ), .Z(n15088) );
  XOR \SUBBYTES[8].a/U5238  ( .A(\SUBBYTES[8].a/w1105 ), .B(
        \SUBBYTES[8].a/w1120 ), .Z(n15089) );
  XOR \SUBBYTES[8].a/U5237  ( .A(n15920), .B(n15090), .Z(n16067) );
  XOR \SUBBYTES[8].a/U5236  ( .A(\SUBBYTES[8].a/w1120 ), .B(
        \SUBBYTES[8].a/w1121 ), .Z(n15090) );
  XOR \SUBBYTES[8].a/U5235  ( .A(\SUBBYTES[8].a/w1082 ), .B(n15091), .Z(n15922) );
  XOR \SUBBYTES[8].a/U5234  ( .A(\SUBBYTES[8].a/w1073 ), .B(
        \SUBBYTES[8].a/w1074 ), .Z(n15091) );
  XOR \SUBBYTES[8].a/U5232  ( .A(\SUBBYTES[8].a/w1084 ), .B(n16067), .Z(n15092) );
  XOR \SUBBYTES[8].a/U5231  ( .A(n15094), .B(n15093), .Z(n15923) );
  XOR \SUBBYTES[8].a/U5230  ( .A(n15096), .B(n15095), .Z(n15093) );
  XOR \SUBBYTES[8].a/U5229  ( .A(\SUBBYTES[8].a/w1120 ), .B(
        \SUBBYTES[8].a/w1121 ), .Z(n15094) );
  XOR \SUBBYTES[8].a/U5228  ( .A(\SUBBYTES[8].a/w1084 ), .B(
        \SUBBYTES[8].a/w1108 ), .Z(n15095) );
  XOR \SUBBYTES[8].a/U5227  ( .A(\SUBBYTES[8].a/w1073 ), .B(
        \SUBBYTES[8].a/w1082 ), .Z(n15096) );
  XOR \SUBBYTES[8].a/U5226  ( .A(\SUBBYTES[8].a/w1105 ), .B(n15097), .Z(n15921) );
  XOR \SUBBYTES[8].a/U5225  ( .A(\SUBBYTES[8].a/w1088 ), .B(
        \SUBBYTES[8].a/w1091 ), .Z(n15097) );
  XOR \SUBBYTES[8].a/U5223  ( .A(\SUBBYTES[8].a/w1076 ), .B(n15923), .Z(n15098) );
  XOR \SUBBYTES[8].a/U5221  ( .A(\SUBBYTES[8].a/w1108 ), .B(
        \SUBBYTES[8].a/w1121 ), .Z(n15099) );
  XOR \SUBBYTES[8].a/U5219  ( .A(n15103), .B(n15102), .Z(n15100) );
  XOR \SUBBYTES[8].a/U5218  ( .A(n15105), .B(n15104), .Z(n15101) );
  XOR \SUBBYTES[8].a/U5217  ( .A(\SUBBYTES[8].a/w1120 ), .B(
        \SUBBYTES[8].a/w1123 ), .Z(n15102) );
  XOR \SUBBYTES[8].a/U5216  ( .A(\SUBBYTES[8].a/w1113 ), .B(
        \SUBBYTES[8].a/w1116 ), .Z(n15103) );
  XOR \SUBBYTES[8].a/U5215  ( .A(\SUBBYTES[8].a/w1088 ), .B(
        \SUBBYTES[8].a/w1089 ), .Z(n15104) );
  XOR \SUBBYTES[8].a/U5214  ( .A(\SUBBYTES[8].a/w1073 ), .B(
        \SUBBYTES[8].a/w1076 ), .Z(n15105) );
  XOR \SUBBYTES[8].a/U5212  ( .A(n15920), .B(n15108), .Z(n15106) );
  XOR \SUBBYTES[8].a/U5211  ( .A(n15922), .B(n15921), .Z(n15107) );
  XOR \SUBBYTES[8].a/U5210  ( .A(\SUBBYTES[8].a/w1081 ), .B(
        \SUBBYTES[8].a/w1108 ), .Z(n15108) );
  XOR \SUBBYTES[8].a/U5208  ( .A(n15923), .B(n15111), .Z(n15109) );
  XOR \SUBBYTES[8].a/U5207  ( .A(\SUBBYTES[8].a/w1114 ), .B(
        \SUBBYTES[8].a/w1116 ), .Z(n15110) );
  XOR \SUBBYTES[8].a/U5206  ( .A(\SUBBYTES[8].a/w1074 ), .B(
        \SUBBYTES[8].a/w1106 ), .Z(n15111) );
  XOR \SUBBYTES[8].a/U5205  ( .A(\SUBBYTES[8].a/w906 ), .B(
        \SUBBYTES[8].a/w907 ), .Z(n15925) );
  XOR \SUBBYTES[8].a/U5204  ( .A(n15925), .B(n15112), .Z(n15924) );
  XOR \SUBBYTES[8].a/U5203  ( .A(\SUBBYTES[8].a/w899 ), .B(
        \SUBBYTES[8].a/w916 ), .Z(n15112) );
  XOR \SUBBYTES[8].a/U5201  ( .A(\SUBBYTES[8].a/w898 ), .B(
        \SUBBYTES[8].a/w913 ), .Z(n15113) );
  XOR \SUBBYTES[8].a/U5200  ( .A(n15925), .B(n15114), .Z(n16068) );
  XOR \SUBBYTES[8].a/U5199  ( .A(\SUBBYTES[8].a/w913 ), .B(
        \SUBBYTES[8].a/w914 ), .Z(n15114) );
  XOR \SUBBYTES[8].a/U5198  ( .A(\SUBBYTES[8].a/w875 ), .B(n15115), .Z(n15927)
         );
  XOR \SUBBYTES[8].a/U5197  ( .A(\SUBBYTES[8].a/w866 ), .B(
        \SUBBYTES[8].a/w867 ), .Z(n15115) );
  XOR \SUBBYTES[8].a/U5195  ( .A(\SUBBYTES[8].a/w877 ), .B(n16068), .Z(n15116)
         );
  XOR \SUBBYTES[8].a/U5194  ( .A(n15118), .B(n15117), .Z(n15928) );
  XOR \SUBBYTES[8].a/U5193  ( .A(n15120), .B(n15119), .Z(n15117) );
  XOR \SUBBYTES[8].a/U5192  ( .A(\SUBBYTES[8].a/w913 ), .B(
        \SUBBYTES[8].a/w914 ), .Z(n15118) );
  XOR \SUBBYTES[8].a/U5191  ( .A(\SUBBYTES[8].a/w877 ), .B(
        \SUBBYTES[8].a/w901 ), .Z(n15119) );
  XOR \SUBBYTES[8].a/U5190  ( .A(\SUBBYTES[8].a/w866 ), .B(
        \SUBBYTES[8].a/w875 ), .Z(n15120) );
  XOR \SUBBYTES[8].a/U5189  ( .A(\SUBBYTES[8].a/w898 ), .B(n15121), .Z(n15926)
         );
  XOR \SUBBYTES[8].a/U5188  ( .A(\SUBBYTES[8].a/w881 ), .B(
        \SUBBYTES[8].a/w884 ), .Z(n15121) );
  XOR \SUBBYTES[8].a/U5186  ( .A(\SUBBYTES[8].a/w869 ), .B(n15928), .Z(n15122)
         );
  XOR \SUBBYTES[8].a/U5184  ( .A(\SUBBYTES[8].a/w901 ), .B(
        \SUBBYTES[8].a/w914 ), .Z(n15123) );
  XOR \SUBBYTES[8].a/U5182  ( .A(n15127), .B(n15126), .Z(n15124) );
  XOR \SUBBYTES[8].a/U5181  ( .A(n15129), .B(n15128), .Z(n15125) );
  XOR \SUBBYTES[8].a/U5180  ( .A(\SUBBYTES[8].a/w913 ), .B(
        \SUBBYTES[8].a/w916 ), .Z(n15126) );
  XOR \SUBBYTES[8].a/U5179  ( .A(\SUBBYTES[8].a/w906 ), .B(
        \SUBBYTES[8].a/w909 ), .Z(n15127) );
  XOR \SUBBYTES[8].a/U5178  ( .A(\SUBBYTES[8].a/w881 ), .B(
        \SUBBYTES[8].a/w882 ), .Z(n15128) );
  XOR \SUBBYTES[8].a/U5177  ( .A(\SUBBYTES[8].a/w866 ), .B(
        \SUBBYTES[8].a/w869 ), .Z(n15129) );
  XOR \SUBBYTES[8].a/U5175  ( .A(n15925), .B(n15132), .Z(n15130) );
  XOR \SUBBYTES[8].a/U5174  ( .A(n15927), .B(n15926), .Z(n15131) );
  XOR \SUBBYTES[8].a/U5173  ( .A(\SUBBYTES[8].a/w874 ), .B(
        \SUBBYTES[8].a/w901 ), .Z(n15132) );
  XOR \SUBBYTES[8].a/U5171  ( .A(n15928), .B(n15135), .Z(n15133) );
  XOR \SUBBYTES[8].a/U5170  ( .A(\SUBBYTES[8].a/w907 ), .B(
        \SUBBYTES[8].a/w909 ), .Z(n15134) );
  XOR \SUBBYTES[8].a/U5169  ( .A(\SUBBYTES[8].a/w867 ), .B(
        \SUBBYTES[8].a/w899 ), .Z(n15135) );
  XOR \SUBBYTES[8].a/U5168  ( .A(\SUBBYTES[8].a/w699 ), .B(
        \SUBBYTES[8].a/w700 ), .Z(n15930) );
  XOR \SUBBYTES[8].a/U5167  ( .A(n15930), .B(n15136), .Z(n15929) );
  XOR \SUBBYTES[8].a/U5166  ( .A(\SUBBYTES[8].a/w692 ), .B(
        \SUBBYTES[8].a/w709 ), .Z(n15136) );
  XOR \SUBBYTES[8].a/U5164  ( .A(\SUBBYTES[8].a/w691 ), .B(
        \SUBBYTES[8].a/w706 ), .Z(n15137) );
  XOR \SUBBYTES[8].a/U5163  ( .A(n15930), .B(n15138), .Z(n16069) );
  XOR \SUBBYTES[8].a/U5162  ( .A(\SUBBYTES[8].a/w706 ), .B(
        \SUBBYTES[8].a/w707 ), .Z(n15138) );
  XOR \SUBBYTES[8].a/U5161  ( .A(\SUBBYTES[8].a/w668 ), .B(n15139), .Z(n15932)
         );
  XOR \SUBBYTES[8].a/U5160  ( .A(\SUBBYTES[8].a/w659 ), .B(
        \SUBBYTES[8].a/w660 ), .Z(n15139) );
  XOR \SUBBYTES[8].a/U5158  ( .A(\SUBBYTES[8].a/w670 ), .B(n16069), .Z(n15140)
         );
  XOR \SUBBYTES[8].a/U5157  ( .A(n15142), .B(n15141), .Z(n15933) );
  XOR \SUBBYTES[8].a/U5156  ( .A(n15144), .B(n15143), .Z(n15141) );
  XOR \SUBBYTES[8].a/U5155  ( .A(\SUBBYTES[8].a/w706 ), .B(
        \SUBBYTES[8].a/w707 ), .Z(n15142) );
  XOR \SUBBYTES[8].a/U5154  ( .A(\SUBBYTES[8].a/w670 ), .B(
        \SUBBYTES[8].a/w694 ), .Z(n15143) );
  XOR \SUBBYTES[8].a/U5153  ( .A(\SUBBYTES[8].a/w659 ), .B(
        \SUBBYTES[8].a/w668 ), .Z(n15144) );
  XOR \SUBBYTES[8].a/U5152  ( .A(\SUBBYTES[8].a/w691 ), .B(n15145), .Z(n15931)
         );
  XOR \SUBBYTES[8].a/U5151  ( .A(\SUBBYTES[8].a/w674 ), .B(
        \SUBBYTES[8].a/w677 ), .Z(n15145) );
  XOR \SUBBYTES[8].a/U5149  ( .A(\SUBBYTES[8].a/w662 ), .B(n15933), .Z(n15146)
         );
  XOR \SUBBYTES[8].a/U5147  ( .A(\SUBBYTES[8].a/w694 ), .B(
        \SUBBYTES[8].a/w707 ), .Z(n15147) );
  XOR \SUBBYTES[8].a/U5145  ( .A(n15151), .B(n15150), .Z(n15148) );
  XOR \SUBBYTES[8].a/U5144  ( .A(n15153), .B(n15152), .Z(n15149) );
  XOR \SUBBYTES[8].a/U5143  ( .A(\SUBBYTES[8].a/w706 ), .B(
        \SUBBYTES[8].a/w709 ), .Z(n15150) );
  XOR \SUBBYTES[8].a/U5142  ( .A(\SUBBYTES[8].a/w699 ), .B(
        \SUBBYTES[8].a/w702 ), .Z(n15151) );
  XOR \SUBBYTES[8].a/U5141  ( .A(\SUBBYTES[8].a/w674 ), .B(
        \SUBBYTES[8].a/w675 ), .Z(n15152) );
  XOR \SUBBYTES[8].a/U5140  ( .A(\SUBBYTES[8].a/w659 ), .B(
        \SUBBYTES[8].a/w662 ), .Z(n15153) );
  XOR \SUBBYTES[8].a/U5138  ( .A(n15930), .B(n15156), .Z(n15154) );
  XOR \SUBBYTES[8].a/U5137  ( .A(n15932), .B(n15931), .Z(n15155) );
  XOR \SUBBYTES[8].a/U5136  ( .A(\SUBBYTES[8].a/w667 ), .B(
        \SUBBYTES[8].a/w694 ), .Z(n15156) );
  XOR \SUBBYTES[8].a/U5134  ( .A(n15933), .B(n15159), .Z(n15157) );
  XOR \SUBBYTES[8].a/U5133  ( .A(\SUBBYTES[8].a/w700 ), .B(
        \SUBBYTES[8].a/w702 ), .Z(n15158) );
  XOR \SUBBYTES[8].a/U5132  ( .A(\SUBBYTES[8].a/w660 ), .B(
        \SUBBYTES[8].a/w692 ), .Z(n15159) );
  XOR \SUBBYTES[8].a/U5131  ( .A(\SUBBYTES[8].a/w492 ), .B(
        \SUBBYTES[8].a/w493 ), .Z(n15935) );
  XOR \SUBBYTES[8].a/U5130  ( .A(n15935), .B(n15160), .Z(n15934) );
  XOR \SUBBYTES[8].a/U5129  ( .A(\SUBBYTES[8].a/w485 ), .B(
        \SUBBYTES[8].a/w502 ), .Z(n15160) );
  XOR \SUBBYTES[8].a/U5127  ( .A(\SUBBYTES[8].a/w484 ), .B(
        \SUBBYTES[8].a/w499 ), .Z(n15161) );
  XOR \SUBBYTES[8].a/U5126  ( .A(n15935), .B(n15162), .Z(n16070) );
  XOR \SUBBYTES[8].a/U5125  ( .A(\SUBBYTES[8].a/w499 ), .B(
        \SUBBYTES[8].a/w500 ), .Z(n15162) );
  XOR \SUBBYTES[8].a/U5124  ( .A(\SUBBYTES[8].a/w461 ), .B(n15163), .Z(n15937)
         );
  XOR \SUBBYTES[8].a/U5123  ( .A(\SUBBYTES[8].a/w452 ), .B(
        \SUBBYTES[8].a/w453 ), .Z(n15163) );
  XOR \SUBBYTES[8].a/U5121  ( .A(\SUBBYTES[8].a/w463 ), .B(n16070), .Z(n15164)
         );
  XOR \SUBBYTES[8].a/U5120  ( .A(n15166), .B(n15165), .Z(n15938) );
  XOR \SUBBYTES[8].a/U5119  ( .A(n15168), .B(n15167), .Z(n15165) );
  XOR \SUBBYTES[8].a/U5118  ( .A(\SUBBYTES[8].a/w499 ), .B(
        \SUBBYTES[8].a/w500 ), .Z(n15166) );
  XOR \SUBBYTES[8].a/U5117  ( .A(\SUBBYTES[8].a/w463 ), .B(
        \SUBBYTES[8].a/w487 ), .Z(n15167) );
  XOR \SUBBYTES[8].a/U5116  ( .A(\SUBBYTES[8].a/w452 ), .B(
        \SUBBYTES[8].a/w461 ), .Z(n15168) );
  XOR \SUBBYTES[8].a/U5115  ( .A(\SUBBYTES[8].a/w484 ), .B(n15169), .Z(n15936)
         );
  XOR \SUBBYTES[8].a/U5114  ( .A(\SUBBYTES[8].a/w467 ), .B(
        \SUBBYTES[8].a/w470 ), .Z(n15169) );
  XOR \SUBBYTES[8].a/U5112  ( .A(\SUBBYTES[8].a/w455 ), .B(n15938), .Z(n15170)
         );
  XOR \SUBBYTES[8].a/U5110  ( .A(\SUBBYTES[8].a/w487 ), .B(
        \SUBBYTES[8].a/w500 ), .Z(n15171) );
  XOR \SUBBYTES[8].a/U5108  ( .A(n15175), .B(n15174), .Z(n15172) );
  XOR \SUBBYTES[8].a/U5107  ( .A(n15177), .B(n15176), .Z(n15173) );
  XOR \SUBBYTES[8].a/U5106  ( .A(\SUBBYTES[8].a/w499 ), .B(
        \SUBBYTES[8].a/w502 ), .Z(n15174) );
  XOR \SUBBYTES[8].a/U5105  ( .A(\SUBBYTES[8].a/w492 ), .B(
        \SUBBYTES[8].a/w495 ), .Z(n15175) );
  XOR \SUBBYTES[8].a/U5104  ( .A(\SUBBYTES[8].a/w467 ), .B(
        \SUBBYTES[8].a/w468 ), .Z(n15176) );
  XOR \SUBBYTES[8].a/U5103  ( .A(\SUBBYTES[8].a/w452 ), .B(
        \SUBBYTES[8].a/w455 ), .Z(n15177) );
  XOR \SUBBYTES[8].a/U5101  ( .A(n15935), .B(n15180), .Z(n15178) );
  XOR \SUBBYTES[8].a/U5100  ( .A(n15937), .B(n15936), .Z(n15179) );
  XOR \SUBBYTES[8].a/U5099  ( .A(\SUBBYTES[8].a/w460 ), .B(
        \SUBBYTES[8].a/w487 ), .Z(n15180) );
  XOR \SUBBYTES[8].a/U5097  ( .A(n15938), .B(n15183), .Z(n15181) );
  XOR \SUBBYTES[8].a/U5096  ( .A(\SUBBYTES[8].a/w493 ), .B(
        \SUBBYTES[8].a/w495 ), .Z(n15182) );
  XOR \SUBBYTES[8].a/U5095  ( .A(\SUBBYTES[8].a/w453 ), .B(
        \SUBBYTES[8].a/w485 ), .Z(n15183) );
  XOR \SUBBYTES[8].a/U5094  ( .A(\SUBBYTES[8].a/w285 ), .B(
        \SUBBYTES[8].a/w286 ), .Z(n15940) );
  XOR \SUBBYTES[8].a/U5093  ( .A(n15940), .B(n15184), .Z(n15939) );
  XOR \SUBBYTES[8].a/U5092  ( .A(\SUBBYTES[8].a/w278 ), .B(
        \SUBBYTES[8].a/w295 ), .Z(n15184) );
  XOR \SUBBYTES[8].a/U5090  ( .A(\SUBBYTES[8].a/w277 ), .B(
        \SUBBYTES[8].a/w292 ), .Z(n15185) );
  XOR \SUBBYTES[8].a/U5089  ( .A(n15940), .B(n15186), .Z(n16071) );
  XOR \SUBBYTES[8].a/U5088  ( .A(\SUBBYTES[8].a/w292 ), .B(
        \SUBBYTES[8].a/w293 ), .Z(n15186) );
  XOR \SUBBYTES[8].a/U5087  ( .A(\SUBBYTES[8].a/w254 ), .B(n15187), .Z(n15942)
         );
  XOR \SUBBYTES[8].a/U5086  ( .A(\SUBBYTES[8].a/w245 ), .B(
        \SUBBYTES[8].a/w246 ), .Z(n15187) );
  XOR \SUBBYTES[8].a/U5084  ( .A(\SUBBYTES[8].a/w256 ), .B(n16071), .Z(n15188)
         );
  XOR \SUBBYTES[8].a/U5083  ( .A(n15190), .B(n15189), .Z(n15943) );
  XOR \SUBBYTES[8].a/U5082  ( .A(n15192), .B(n15191), .Z(n15189) );
  XOR \SUBBYTES[8].a/U5081  ( .A(\SUBBYTES[8].a/w292 ), .B(
        \SUBBYTES[8].a/w293 ), .Z(n15190) );
  XOR \SUBBYTES[8].a/U5080  ( .A(\SUBBYTES[8].a/w256 ), .B(
        \SUBBYTES[8].a/w280 ), .Z(n15191) );
  XOR \SUBBYTES[8].a/U5079  ( .A(\SUBBYTES[8].a/w245 ), .B(
        \SUBBYTES[8].a/w254 ), .Z(n15192) );
  XOR \SUBBYTES[8].a/U5078  ( .A(\SUBBYTES[8].a/w277 ), .B(n15193), .Z(n15941)
         );
  XOR \SUBBYTES[8].a/U5077  ( .A(\SUBBYTES[8].a/w260 ), .B(
        \SUBBYTES[8].a/w263 ), .Z(n15193) );
  XOR \SUBBYTES[8].a/U5075  ( .A(\SUBBYTES[8].a/w248 ), .B(n15943), .Z(n15194)
         );
  XOR \SUBBYTES[8].a/U5073  ( .A(\SUBBYTES[8].a/w280 ), .B(
        \SUBBYTES[8].a/w293 ), .Z(n15195) );
  XOR \SUBBYTES[8].a/U5071  ( .A(n15199), .B(n15198), .Z(n15196) );
  XOR \SUBBYTES[8].a/U5070  ( .A(n15201), .B(n15200), .Z(n15197) );
  XOR \SUBBYTES[8].a/U5069  ( .A(\SUBBYTES[8].a/w292 ), .B(
        \SUBBYTES[8].a/w295 ), .Z(n15198) );
  XOR \SUBBYTES[8].a/U5068  ( .A(\SUBBYTES[8].a/w285 ), .B(
        \SUBBYTES[8].a/w288 ), .Z(n15199) );
  XOR \SUBBYTES[8].a/U5067  ( .A(\SUBBYTES[8].a/w260 ), .B(
        \SUBBYTES[8].a/w261 ), .Z(n15200) );
  XOR \SUBBYTES[8].a/U5066  ( .A(\SUBBYTES[8].a/w245 ), .B(
        \SUBBYTES[8].a/w248 ), .Z(n15201) );
  XOR \SUBBYTES[8].a/U5064  ( .A(n15940), .B(n15204), .Z(n15202) );
  XOR \SUBBYTES[8].a/U5063  ( .A(n15942), .B(n15941), .Z(n15203) );
  XOR \SUBBYTES[8].a/U5062  ( .A(\SUBBYTES[8].a/w253 ), .B(
        \SUBBYTES[8].a/w280 ), .Z(n15204) );
  XOR \SUBBYTES[8].a/U5060  ( .A(n15943), .B(n15207), .Z(n15205) );
  XOR \SUBBYTES[8].a/U5059  ( .A(\SUBBYTES[8].a/w286 ), .B(
        \SUBBYTES[8].a/w288 ), .Z(n15206) );
  XOR \SUBBYTES[8].a/U5058  ( .A(\SUBBYTES[8].a/w246 ), .B(
        \SUBBYTES[8].a/w278 ), .Z(n15207) );
  XOR \SUBBYTES[8].a/U5057  ( .A(\w1[8][1] ), .B(n15208), .Z(n15944) );
  XOR \SUBBYTES[8].a/U5056  ( .A(\w1[8][3] ), .B(\w1[8][2] ), .Z(n15208) );
  XOR \SUBBYTES[8].a/U5055  ( .A(\w1[8][6] ), .B(n15944), .Z(
        \SUBBYTES[8].a/w3378 ) );
  XOR \SUBBYTES[8].a/U5054  ( .A(\w1[8][0] ), .B(\SUBBYTES[8].a/w3378 ), .Z(
        \SUBBYTES[8].a/w3265 ) );
  XOR \SUBBYTES[8].a/U5053  ( .A(\w1[8][0] ), .B(n15209), .Z(
        \SUBBYTES[8].a/w3266 ) );
  XOR \SUBBYTES[8].a/U5052  ( .A(\w1[8][6] ), .B(\w1[8][5] ), .Z(n15209) );
  XOR \SUBBYTES[8].a/U5051  ( .A(\w1[8][5] ), .B(n15944), .Z(
        \SUBBYTES[8].a/w3396 ) );
  XOR \SUBBYTES[8].a/U5050  ( .A(n15211), .B(n15210), .Z(\SUBBYTES[8].a/w3389 ) );
  XOR \SUBBYTES[8].a/U5049  ( .A(\w1[8][3] ), .B(\w1[8][1] ), .Z(n15210) );
  XOR \SUBBYTES[8].a/U5048  ( .A(\w1[8][7] ), .B(\w1[8][4] ), .Z(n15211) );
  XOR \SUBBYTES[8].a/U5047  ( .A(\w1[8][0] ), .B(\SUBBYTES[8].a/w3389 ), .Z(
        \SUBBYTES[8].a/w3268 ) );
  XOR \SUBBYTES[8].a/U5046  ( .A(n15213), .B(n15212), .Z(\SUBBYTES[8].a/w3376 ) );
  XOR \SUBBYTES[8].a/U5045  ( .A(\SUBBYTES[8].a/w3337 ), .B(n1084), .Z(n15212)
         );
  XOR \SUBBYTES[8].a/U5044  ( .A(\SUBBYTES[8].a/w3330 ), .B(
        \SUBBYTES[8].a/w3333 ), .Z(n15213) );
  XOR \SUBBYTES[8].a/U5043  ( .A(n15215), .B(n15214), .Z(\SUBBYTES[8].a/w3377 ) );
  XOR \SUBBYTES[8].a/U5042  ( .A(\SUBBYTES[8].a/w3337 ), .B(n14823), .Z(n15214) );
  XOR \SUBBYTES[8].a/U5041  ( .A(\SUBBYTES[8].a/w3330 ), .B(n14822), .Z(n15215) );
  XOR \SUBBYTES[8].a/U5040  ( .A(\SUBBYTES[8].a/w3389 ), .B(n15216), .Z(
        \SUBBYTES[8].a/w3379 ) );
  XOR \SUBBYTES[8].a/U5039  ( .A(\w1[8][6] ), .B(\w1[8][5] ), .Z(n15216) );
  XOR \SUBBYTES[8].a/U5038  ( .A(n15218), .B(n15217), .Z(\SUBBYTES[8].a/w3380 ) );
  XOR \SUBBYTES[8].a/U5037  ( .A(n14823), .B(n1084), .Z(n15217) );
  XOR \SUBBYTES[8].a/U5036  ( .A(n14822), .B(\SUBBYTES[8].a/w3333 ), .Z(n15218) );
  XOR \SUBBYTES[8].a/U5035  ( .A(\w1[8][7] ), .B(\w1[8][2] ), .Z(n15950) );
  XOR \SUBBYTES[8].a/U5034  ( .A(n15950), .B(n15219), .Z(\SUBBYTES[8].a/w3381 ) );
  XOR \SUBBYTES[8].a/U5033  ( .A(\w1[8][5] ), .B(\w1[8][4] ), .Z(n15219) );
  XOR \SUBBYTES[8].a/U5032  ( .A(\w1[8][7] ), .B(\SUBBYTES[8].a/w3266 ), .Z(
        \SUBBYTES[8].a/w3269 ) );
  XOR \SUBBYTES[8].a/U5031  ( .A(\w1[8][1] ), .B(\SUBBYTES[8].a/w3266 ), .Z(
        \SUBBYTES[8].a/w3270 ) );
  XOR \SUBBYTES[8].a/U5030  ( .A(\w1[8][4] ), .B(\SUBBYTES[8].a/w3266 ), .Z(
        \SUBBYTES[8].a/w3271 ) );
  XOR \SUBBYTES[8].a/U5029  ( .A(\SUBBYTES[8].a/w3270 ), .B(n15950), .Z(
        \SUBBYTES[8].a/w3272 ) );
  XOR \SUBBYTES[8].a/U5028  ( .A(n15950), .B(n15220), .Z(\SUBBYTES[8].a/w3357 ) );
  XOR \SUBBYTES[8].a/U5027  ( .A(\w1[8][4] ), .B(\w1[8][1] ), .Z(n15220) );
  XOR \SUBBYTES[8].a/U5026  ( .A(n15222), .B(n15221), .Z(n15947) );
  XOR \SUBBYTES[8].a/U5025  ( .A(\w1[8][4] ), .B(n15223), .Z(n15221) );
  XOR \SUBBYTES[8].a/U5024  ( .A(\SUBBYTES[8].a/w3322 ), .B(\w1[8][6] ), .Z(
        n15222) );
  XOR \SUBBYTES[8].a/U5023  ( .A(\SUBBYTES[8].a/w3296 ), .B(
        \SUBBYTES[8].a/w3303 ), .Z(n15223) );
  XOR \SUBBYTES[8].a/U5022  ( .A(n15225), .B(n15224), .Z(n15945) );
  XOR \SUBBYTES[8].a/U5021  ( .A(\w1[8][1] ), .B(n15226), .Z(n15224) );
  XOR \SUBBYTES[8].a/U5020  ( .A(\SUBBYTES[8].a/w3321 ), .B(\w1[8][5] ), .Z(
        n15225) );
  XOR \SUBBYTES[8].a/U5019  ( .A(\SUBBYTES[8].a/w3297 ), .B(
        \SUBBYTES[8].a/w3304 ), .Z(n15226) );
  XOR \SUBBYTES[8].a/U5018  ( .A(n15947), .B(n15945), .Z(\SUBBYTES[8].a/w3327 ) );
  XOR \SUBBYTES[8].a/U5017  ( .A(\w1[8][5] ), .B(n15227), .Z(n15948) );
  XOR \SUBBYTES[8].a/U5016  ( .A(\SUBBYTES[8].a/w3289 ), .B(
        \SUBBYTES[8].a/w3299 ), .Z(n15227) );
  XOR \SUBBYTES[8].a/U5015  ( .A(n15229), .B(n15228), .Z(\SUBBYTES[8].a/w3314 ) );
  XOR \SUBBYTES[8].a/U5014  ( .A(n15948), .B(n15230), .Z(n15228) );
  XOR \SUBBYTES[8].a/U5013  ( .A(\w1[8][4] ), .B(\SUBBYTES[8].a/w3378 ), .Z(
        n15229) );
  XOR \SUBBYTES[8].a/U5012  ( .A(\SUBBYTES[8].a/w3291 ), .B(
        \SUBBYTES[8].a/w3296 ), .Z(n15230) );
  XOR \SUBBYTES[8].a/U5011  ( .A(n15232), .B(n15231), .Z(n15946) );
  XOR \SUBBYTES[8].a/U5010  ( .A(\SUBBYTES[8].a/w3324 ), .B(\w1[8][7] ), .Z(
        n15231) );
  XOR \SUBBYTES[8].a/U5009  ( .A(\SUBBYTES[8].a/w3299 ), .B(
        \SUBBYTES[8].a/w3306 ), .Z(n15232) );
  XOR \SUBBYTES[8].a/U5008  ( .A(n15945), .B(n15946), .Z(\SUBBYTES[8].a/w3326 ) );
  XOR \SUBBYTES[8].a/U5007  ( .A(\w1[8][3] ), .B(n15233), .Z(n15949) );
  XOR \SUBBYTES[8].a/U5006  ( .A(\SUBBYTES[8].a/w3288 ), .B(
        \SUBBYTES[8].a/w3291 ), .Z(n15233) );
  XOR \SUBBYTES[8].a/U5005  ( .A(n15235), .B(n15234), .Z(\SUBBYTES[8].a/w3315 ) );
  XOR \SUBBYTES[8].a/U5004  ( .A(n15949), .B(n15236), .Z(n15234) );
  XOR \SUBBYTES[8].a/U5003  ( .A(\w1[8][6] ), .B(\SUBBYTES[8].a/w3357 ), .Z(
        n15235) );
  XOR \SUBBYTES[8].a/U5002  ( .A(\SUBBYTES[8].a/w3296 ), .B(
        \SUBBYTES[8].a/w3297 ), .Z(n15236) );
  XOR \SUBBYTES[8].a/U5001  ( .A(n15947), .B(n15946), .Z(\SUBBYTES[8].a/w3335 ) );
  XOR \SUBBYTES[8].a/U5000  ( .A(n15238), .B(n15237), .Z(\SUBBYTES[8].a/w3336 ) );
  XOR \SUBBYTES[8].a/U4999  ( .A(\w1[8][7] ), .B(n15948), .Z(n15237) );
  XOR \SUBBYTES[8].a/U4998  ( .A(\SUBBYTES[8].a/w3288 ), .B(
        \SUBBYTES[8].a/w3297 ), .Z(n15238) );
  XOR \SUBBYTES[8].a/U4997  ( .A(n15240), .B(n15239), .Z(\SUBBYTES[8].a/w3312 ) );
  XOR \SUBBYTES[8].a/U4996  ( .A(n15242), .B(n15241), .Z(n15239) );
  XOR \SUBBYTES[8].a/U4995  ( .A(\w1[8][7] ), .B(\SUBBYTES[8].a/w3396 ), .Z(
        n15240) );
  XOR \SUBBYTES[8].a/U4994  ( .A(\SUBBYTES[8].a/w3303 ), .B(
        \SUBBYTES[8].a/w3306 ), .Z(n15241) );
  XOR \SUBBYTES[8].a/U4993  ( .A(\SUBBYTES[8].a/w3289 ), .B(
        \SUBBYTES[8].a/w3291 ), .Z(n15242) );
  XOR \SUBBYTES[8].a/U4992  ( .A(n15244), .B(n15243), .Z(\SUBBYTES[8].a/w3313 ) );
  XOR \SUBBYTES[8].a/U4991  ( .A(n15949), .B(n15245), .Z(n15243) );
  XOR \SUBBYTES[8].a/U4990  ( .A(\w1[8][5] ), .B(n15950), .Z(n15244) );
  XOR \SUBBYTES[8].a/U4989  ( .A(\SUBBYTES[8].a/w3303 ), .B(
        \SUBBYTES[8].a/w3304 ), .Z(n15245) );
  XOR \SUBBYTES[8].a/U4988  ( .A(n15247), .B(n15246), .Z(\SUBBYTES[8].a/w3329 ) );
  XOR \SUBBYTES[8].a/U4987  ( .A(\w1[8][1] ), .B(n15248), .Z(n15246) );
  XOR \SUBBYTES[8].a/U4986  ( .A(\SUBBYTES[8].a/w3304 ), .B(
        \SUBBYTES[8].a/w3306 ), .Z(n15247) );
  XOR \SUBBYTES[8].a/U4985  ( .A(\SUBBYTES[8].a/w3288 ), .B(
        \SUBBYTES[8].a/w3289 ), .Z(n15248) );
  XOR \SUBBYTES[8].a/U4984  ( .A(\w1[8][9] ), .B(n15249), .Z(n15951) );
  XOR \SUBBYTES[8].a/U4983  ( .A(\w1[8][11] ), .B(\w1[8][10] ), .Z(n15249) );
  XOR \SUBBYTES[8].a/U4982  ( .A(\w1[8][14] ), .B(n15951), .Z(
        \SUBBYTES[8].a/w3171 ) );
  XOR \SUBBYTES[8].a/U4981  ( .A(\w1[8][8] ), .B(\SUBBYTES[8].a/w3171 ), .Z(
        \SUBBYTES[8].a/w3058 ) );
  XOR \SUBBYTES[8].a/U4980  ( .A(\w1[8][8] ), .B(n15250), .Z(
        \SUBBYTES[8].a/w3059 ) );
  XOR \SUBBYTES[8].a/U4979  ( .A(\w1[8][14] ), .B(\w1[8][13] ), .Z(n15250) );
  XOR \SUBBYTES[8].a/U4978  ( .A(\w1[8][13] ), .B(n15951), .Z(
        \SUBBYTES[8].a/w3189 ) );
  XOR \SUBBYTES[8].a/U4977  ( .A(n15252), .B(n15251), .Z(\SUBBYTES[8].a/w3182 ) );
  XOR \SUBBYTES[8].a/U4976  ( .A(\w1[8][11] ), .B(\w1[8][9] ), .Z(n15251) );
  XOR \SUBBYTES[8].a/U4975  ( .A(\w1[8][15] ), .B(\w1[8][12] ), .Z(n15252) );
  XOR \SUBBYTES[8].a/U4974  ( .A(\w1[8][8] ), .B(\SUBBYTES[8].a/w3182 ), .Z(
        \SUBBYTES[8].a/w3061 ) );
  XOR \SUBBYTES[8].a/U4973  ( .A(n15254), .B(n15253), .Z(\SUBBYTES[8].a/w3169 ) );
  XOR \SUBBYTES[8].a/U4972  ( .A(\SUBBYTES[8].a/w3130 ), .B(n1083), .Z(n15253)
         );
  XOR \SUBBYTES[8].a/U4971  ( .A(\SUBBYTES[8].a/w3123 ), .B(
        \SUBBYTES[8].a/w3126 ), .Z(n15254) );
  XOR \SUBBYTES[8].a/U4970  ( .A(n15256), .B(n15255), .Z(\SUBBYTES[8].a/w3170 ) );
  XOR \SUBBYTES[8].a/U4969  ( .A(\SUBBYTES[8].a/w3130 ), .B(n14821), .Z(n15255) );
  XOR \SUBBYTES[8].a/U4968  ( .A(\SUBBYTES[8].a/w3123 ), .B(n14820), .Z(n15256) );
  XOR \SUBBYTES[8].a/U4967  ( .A(\SUBBYTES[8].a/w3182 ), .B(n15257), .Z(
        \SUBBYTES[8].a/w3172 ) );
  XOR \SUBBYTES[8].a/U4966  ( .A(\w1[8][14] ), .B(\w1[8][13] ), .Z(n15257) );
  XOR \SUBBYTES[8].a/U4965  ( .A(n15259), .B(n15258), .Z(\SUBBYTES[8].a/w3173 ) );
  XOR \SUBBYTES[8].a/U4964  ( .A(n14821), .B(n1083), .Z(n15258) );
  XOR \SUBBYTES[8].a/U4963  ( .A(n14820), .B(\SUBBYTES[8].a/w3126 ), .Z(n15259) );
  XOR \SUBBYTES[8].a/U4962  ( .A(\w1[8][15] ), .B(\w1[8][10] ), .Z(n15957) );
  XOR \SUBBYTES[8].a/U4961  ( .A(n15957), .B(n15260), .Z(\SUBBYTES[8].a/w3174 ) );
  XOR \SUBBYTES[8].a/U4960  ( .A(\w1[8][13] ), .B(\w1[8][12] ), .Z(n15260) );
  XOR \SUBBYTES[8].a/U4959  ( .A(\w1[8][15] ), .B(\SUBBYTES[8].a/w3059 ), .Z(
        \SUBBYTES[8].a/w3062 ) );
  XOR \SUBBYTES[8].a/U4958  ( .A(\w1[8][9] ), .B(\SUBBYTES[8].a/w3059 ), .Z(
        \SUBBYTES[8].a/w3063 ) );
  XOR \SUBBYTES[8].a/U4957  ( .A(\w1[8][12] ), .B(\SUBBYTES[8].a/w3059 ), .Z(
        \SUBBYTES[8].a/w3064 ) );
  XOR \SUBBYTES[8].a/U4956  ( .A(\SUBBYTES[8].a/w3063 ), .B(n15957), .Z(
        \SUBBYTES[8].a/w3065 ) );
  XOR \SUBBYTES[8].a/U4955  ( .A(n15957), .B(n15261), .Z(\SUBBYTES[8].a/w3150 ) );
  XOR \SUBBYTES[8].a/U4954  ( .A(\w1[8][12] ), .B(\w1[8][9] ), .Z(n15261) );
  XOR \SUBBYTES[8].a/U4953  ( .A(n15263), .B(n15262), .Z(n15954) );
  XOR \SUBBYTES[8].a/U4952  ( .A(\w1[8][12] ), .B(n15264), .Z(n15262) );
  XOR \SUBBYTES[8].a/U4951  ( .A(\SUBBYTES[8].a/w3115 ), .B(\w1[8][14] ), .Z(
        n15263) );
  XOR \SUBBYTES[8].a/U4950  ( .A(\SUBBYTES[8].a/w3089 ), .B(
        \SUBBYTES[8].a/w3096 ), .Z(n15264) );
  XOR \SUBBYTES[8].a/U4949  ( .A(n15266), .B(n15265), .Z(n15952) );
  XOR \SUBBYTES[8].a/U4948  ( .A(\w1[8][9] ), .B(n15267), .Z(n15265) );
  XOR \SUBBYTES[8].a/U4947  ( .A(\SUBBYTES[8].a/w3114 ), .B(\w1[8][13] ), .Z(
        n15266) );
  XOR \SUBBYTES[8].a/U4946  ( .A(\SUBBYTES[8].a/w3090 ), .B(
        \SUBBYTES[8].a/w3097 ), .Z(n15267) );
  XOR \SUBBYTES[8].a/U4945  ( .A(n15954), .B(n15952), .Z(\SUBBYTES[8].a/w3120 ) );
  XOR \SUBBYTES[8].a/U4944  ( .A(\w1[8][13] ), .B(n15268), .Z(n15955) );
  XOR \SUBBYTES[8].a/U4943  ( .A(\SUBBYTES[8].a/w3082 ), .B(
        \SUBBYTES[8].a/w3092 ), .Z(n15268) );
  XOR \SUBBYTES[8].a/U4942  ( .A(n15270), .B(n15269), .Z(\SUBBYTES[8].a/w3107 ) );
  XOR \SUBBYTES[8].a/U4941  ( .A(n15955), .B(n15271), .Z(n15269) );
  XOR \SUBBYTES[8].a/U4940  ( .A(\w1[8][12] ), .B(\SUBBYTES[8].a/w3171 ), .Z(
        n15270) );
  XOR \SUBBYTES[8].a/U4939  ( .A(\SUBBYTES[8].a/w3084 ), .B(
        \SUBBYTES[8].a/w3089 ), .Z(n15271) );
  XOR \SUBBYTES[8].a/U4938  ( .A(n15273), .B(n15272), .Z(n15953) );
  XOR \SUBBYTES[8].a/U4937  ( .A(\SUBBYTES[8].a/w3117 ), .B(\w1[8][15] ), .Z(
        n15272) );
  XOR \SUBBYTES[8].a/U4936  ( .A(\SUBBYTES[8].a/w3092 ), .B(
        \SUBBYTES[8].a/w3099 ), .Z(n15273) );
  XOR \SUBBYTES[8].a/U4935  ( .A(n15952), .B(n15953), .Z(\SUBBYTES[8].a/w3119 ) );
  XOR \SUBBYTES[8].a/U4934  ( .A(\w1[8][11] ), .B(n15274), .Z(n15956) );
  XOR \SUBBYTES[8].a/U4933  ( .A(\SUBBYTES[8].a/w3081 ), .B(
        \SUBBYTES[8].a/w3084 ), .Z(n15274) );
  XOR \SUBBYTES[8].a/U4932  ( .A(n15276), .B(n15275), .Z(\SUBBYTES[8].a/w3108 ) );
  XOR \SUBBYTES[8].a/U4931  ( .A(n15956), .B(n15277), .Z(n15275) );
  XOR \SUBBYTES[8].a/U4930  ( .A(\w1[8][14] ), .B(\SUBBYTES[8].a/w3150 ), .Z(
        n15276) );
  XOR \SUBBYTES[8].a/U4929  ( .A(\SUBBYTES[8].a/w3089 ), .B(
        \SUBBYTES[8].a/w3090 ), .Z(n15277) );
  XOR \SUBBYTES[8].a/U4928  ( .A(n15954), .B(n15953), .Z(\SUBBYTES[8].a/w3128 ) );
  XOR \SUBBYTES[8].a/U4927  ( .A(n15279), .B(n15278), .Z(\SUBBYTES[8].a/w3129 ) );
  XOR \SUBBYTES[8].a/U4926  ( .A(\w1[8][15] ), .B(n15955), .Z(n15278) );
  XOR \SUBBYTES[8].a/U4925  ( .A(\SUBBYTES[8].a/w3081 ), .B(
        \SUBBYTES[8].a/w3090 ), .Z(n15279) );
  XOR \SUBBYTES[8].a/U4924  ( .A(n15281), .B(n15280), .Z(\SUBBYTES[8].a/w3105 ) );
  XOR \SUBBYTES[8].a/U4923  ( .A(n15283), .B(n15282), .Z(n15280) );
  XOR \SUBBYTES[8].a/U4922  ( .A(\w1[8][15] ), .B(\SUBBYTES[8].a/w3189 ), .Z(
        n15281) );
  XOR \SUBBYTES[8].a/U4921  ( .A(\SUBBYTES[8].a/w3096 ), .B(
        \SUBBYTES[8].a/w3099 ), .Z(n15282) );
  XOR \SUBBYTES[8].a/U4920  ( .A(\SUBBYTES[8].a/w3082 ), .B(
        \SUBBYTES[8].a/w3084 ), .Z(n15283) );
  XOR \SUBBYTES[8].a/U4919  ( .A(n15285), .B(n15284), .Z(\SUBBYTES[8].a/w3106 ) );
  XOR \SUBBYTES[8].a/U4918  ( .A(n15956), .B(n15286), .Z(n15284) );
  XOR \SUBBYTES[8].a/U4917  ( .A(\w1[8][13] ), .B(n15957), .Z(n15285) );
  XOR \SUBBYTES[8].a/U4916  ( .A(\SUBBYTES[8].a/w3096 ), .B(
        \SUBBYTES[8].a/w3097 ), .Z(n15286) );
  XOR \SUBBYTES[8].a/U4915  ( .A(n15288), .B(n15287), .Z(\SUBBYTES[8].a/w3122 ) );
  XOR \SUBBYTES[8].a/U4914  ( .A(\w1[8][9] ), .B(n15289), .Z(n15287) );
  XOR \SUBBYTES[8].a/U4913  ( .A(\SUBBYTES[8].a/w3097 ), .B(
        \SUBBYTES[8].a/w3099 ), .Z(n15288) );
  XOR \SUBBYTES[8].a/U4912  ( .A(\SUBBYTES[8].a/w3081 ), .B(
        \SUBBYTES[8].a/w3082 ), .Z(n15289) );
  XOR \SUBBYTES[8].a/U4911  ( .A(\w1[8][17] ), .B(n15290), .Z(n15958) );
  XOR \SUBBYTES[8].a/U4910  ( .A(\w1[8][19] ), .B(\w1[8][18] ), .Z(n15290) );
  XOR \SUBBYTES[8].a/U4909  ( .A(\w1[8][22] ), .B(n15958), .Z(
        \SUBBYTES[8].a/w2964 ) );
  XOR \SUBBYTES[8].a/U4908  ( .A(\w1[8][16] ), .B(\SUBBYTES[8].a/w2964 ), .Z(
        \SUBBYTES[8].a/w2851 ) );
  XOR \SUBBYTES[8].a/U4907  ( .A(\w1[8][16] ), .B(n15291), .Z(
        \SUBBYTES[8].a/w2852 ) );
  XOR \SUBBYTES[8].a/U4906  ( .A(\w1[8][22] ), .B(\w1[8][21] ), .Z(n15291) );
  XOR \SUBBYTES[8].a/U4905  ( .A(\w1[8][21] ), .B(n15958), .Z(
        \SUBBYTES[8].a/w2982 ) );
  XOR \SUBBYTES[8].a/U4904  ( .A(n15293), .B(n15292), .Z(\SUBBYTES[8].a/w2975 ) );
  XOR \SUBBYTES[8].a/U4903  ( .A(\w1[8][19] ), .B(\w1[8][17] ), .Z(n15292) );
  XOR \SUBBYTES[8].a/U4902  ( .A(\w1[8][23] ), .B(\w1[8][20] ), .Z(n15293) );
  XOR \SUBBYTES[8].a/U4901  ( .A(\w1[8][16] ), .B(\SUBBYTES[8].a/w2975 ), .Z(
        \SUBBYTES[8].a/w2854 ) );
  XOR \SUBBYTES[8].a/U4900  ( .A(n15295), .B(n15294), .Z(\SUBBYTES[8].a/w2962 ) );
  XOR \SUBBYTES[8].a/U4899  ( .A(\SUBBYTES[8].a/w2923 ), .B(n1082), .Z(n15294)
         );
  XOR \SUBBYTES[8].a/U4898  ( .A(\SUBBYTES[8].a/w2916 ), .B(
        \SUBBYTES[8].a/w2919 ), .Z(n15295) );
  XOR \SUBBYTES[8].a/U4897  ( .A(n15297), .B(n15296), .Z(\SUBBYTES[8].a/w2963 ) );
  XOR \SUBBYTES[8].a/U4896  ( .A(\SUBBYTES[8].a/w2923 ), .B(n14819), .Z(n15296) );
  XOR \SUBBYTES[8].a/U4895  ( .A(\SUBBYTES[8].a/w2916 ), .B(n14818), .Z(n15297) );
  XOR \SUBBYTES[8].a/U4894  ( .A(\SUBBYTES[8].a/w2975 ), .B(n15298), .Z(
        \SUBBYTES[8].a/w2965 ) );
  XOR \SUBBYTES[8].a/U4893  ( .A(\w1[8][22] ), .B(\w1[8][21] ), .Z(n15298) );
  XOR \SUBBYTES[8].a/U4892  ( .A(n15300), .B(n15299), .Z(\SUBBYTES[8].a/w2966 ) );
  XOR \SUBBYTES[8].a/U4891  ( .A(n14819), .B(n1082), .Z(n15299) );
  XOR \SUBBYTES[8].a/U4890  ( .A(n14818), .B(\SUBBYTES[8].a/w2919 ), .Z(n15300) );
  XOR \SUBBYTES[8].a/U4889  ( .A(\w1[8][23] ), .B(\w1[8][18] ), .Z(n15964) );
  XOR \SUBBYTES[8].a/U4888  ( .A(n15964), .B(n15301), .Z(\SUBBYTES[8].a/w2967 ) );
  XOR \SUBBYTES[8].a/U4887  ( .A(\w1[8][21] ), .B(\w1[8][20] ), .Z(n15301) );
  XOR \SUBBYTES[8].a/U4886  ( .A(\w1[8][23] ), .B(\SUBBYTES[8].a/w2852 ), .Z(
        \SUBBYTES[8].a/w2855 ) );
  XOR \SUBBYTES[8].a/U4885  ( .A(\w1[8][17] ), .B(\SUBBYTES[8].a/w2852 ), .Z(
        \SUBBYTES[8].a/w2856 ) );
  XOR \SUBBYTES[8].a/U4884  ( .A(\w1[8][20] ), .B(\SUBBYTES[8].a/w2852 ), .Z(
        \SUBBYTES[8].a/w2857 ) );
  XOR \SUBBYTES[8].a/U4883  ( .A(\SUBBYTES[8].a/w2856 ), .B(n15964), .Z(
        \SUBBYTES[8].a/w2858 ) );
  XOR \SUBBYTES[8].a/U4882  ( .A(n15964), .B(n15302), .Z(\SUBBYTES[8].a/w2943 ) );
  XOR \SUBBYTES[8].a/U4881  ( .A(\w1[8][20] ), .B(\w1[8][17] ), .Z(n15302) );
  XOR \SUBBYTES[8].a/U4880  ( .A(n15304), .B(n15303), .Z(n15961) );
  XOR \SUBBYTES[8].a/U4879  ( .A(\w1[8][20] ), .B(n15305), .Z(n15303) );
  XOR \SUBBYTES[8].a/U4878  ( .A(\SUBBYTES[8].a/w2908 ), .B(\w1[8][22] ), .Z(
        n15304) );
  XOR \SUBBYTES[8].a/U4877  ( .A(\SUBBYTES[8].a/w2882 ), .B(
        \SUBBYTES[8].a/w2889 ), .Z(n15305) );
  XOR \SUBBYTES[8].a/U4876  ( .A(n15307), .B(n15306), .Z(n15959) );
  XOR \SUBBYTES[8].a/U4875  ( .A(\w1[8][17] ), .B(n15308), .Z(n15306) );
  XOR \SUBBYTES[8].a/U4874  ( .A(\SUBBYTES[8].a/w2907 ), .B(\w1[8][21] ), .Z(
        n15307) );
  XOR \SUBBYTES[8].a/U4873  ( .A(\SUBBYTES[8].a/w2883 ), .B(
        \SUBBYTES[8].a/w2890 ), .Z(n15308) );
  XOR \SUBBYTES[8].a/U4872  ( .A(n15961), .B(n15959), .Z(\SUBBYTES[8].a/w2913 ) );
  XOR \SUBBYTES[8].a/U4871  ( .A(\w1[8][21] ), .B(n15309), .Z(n15962) );
  XOR \SUBBYTES[8].a/U4870  ( .A(\SUBBYTES[8].a/w2875 ), .B(
        \SUBBYTES[8].a/w2885 ), .Z(n15309) );
  XOR \SUBBYTES[8].a/U4869  ( .A(n15311), .B(n15310), .Z(\SUBBYTES[8].a/w2900 ) );
  XOR \SUBBYTES[8].a/U4868  ( .A(n15962), .B(n15312), .Z(n15310) );
  XOR \SUBBYTES[8].a/U4867  ( .A(\w1[8][20] ), .B(\SUBBYTES[8].a/w2964 ), .Z(
        n15311) );
  XOR \SUBBYTES[8].a/U4866  ( .A(\SUBBYTES[8].a/w2877 ), .B(
        \SUBBYTES[8].a/w2882 ), .Z(n15312) );
  XOR \SUBBYTES[8].a/U4865  ( .A(n15314), .B(n15313), .Z(n15960) );
  XOR \SUBBYTES[8].a/U4864  ( .A(\SUBBYTES[8].a/w2910 ), .B(\w1[8][23] ), .Z(
        n15313) );
  XOR \SUBBYTES[8].a/U4863  ( .A(\SUBBYTES[8].a/w2885 ), .B(
        \SUBBYTES[8].a/w2892 ), .Z(n15314) );
  XOR \SUBBYTES[8].a/U4862  ( .A(n15959), .B(n15960), .Z(\SUBBYTES[8].a/w2912 ) );
  XOR \SUBBYTES[8].a/U4861  ( .A(\w1[8][19] ), .B(n15315), .Z(n15963) );
  XOR \SUBBYTES[8].a/U4860  ( .A(\SUBBYTES[8].a/w2874 ), .B(
        \SUBBYTES[8].a/w2877 ), .Z(n15315) );
  XOR \SUBBYTES[8].a/U4859  ( .A(n15317), .B(n15316), .Z(\SUBBYTES[8].a/w2901 ) );
  XOR \SUBBYTES[8].a/U4858  ( .A(n15963), .B(n15318), .Z(n15316) );
  XOR \SUBBYTES[8].a/U4857  ( .A(\w1[8][22] ), .B(\SUBBYTES[8].a/w2943 ), .Z(
        n15317) );
  XOR \SUBBYTES[8].a/U4856  ( .A(\SUBBYTES[8].a/w2882 ), .B(
        \SUBBYTES[8].a/w2883 ), .Z(n15318) );
  XOR \SUBBYTES[8].a/U4855  ( .A(n15961), .B(n15960), .Z(\SUBBYTES[8].a/w2921 ) );
  XOR \SUBBYTES[8].a/U4854  ( .A(n15320), .B(n15319), .Z(\SUBBYTES[8].a/w2922 ) );
  XOR \SUBBYTES[8].a/U4853  ( .A(\w1[8][23] ), .B(n15962), .Z(n15319) );
  XOR \SUBBYTES[8].a/U4852  ( .A(\SUBBYTES[8].a/w2874 ), .B(
        \SUBBYTES[8].a/w2883 ), .Z(n15320) );
  XOR \SUBBYTES[8].a/U4851  ( .A(n15322), .B(n15321), .Z(\SUBBYTES[8].a/w2898 ) );
  XOR \SUBBYTES[8].a/U4850  ( .A(n15324), .B(n15323), .Z(n15321) );
  XOR \SUBBYTES[8].a/U4849  ( .A(\w1[8][23] ), .B(\SUBBYTES[8].a/w2982 ), .Z(
        n15322) );
  XOR \SUBBYTES[8].a/U4848  ( .A(\SUBBYTES[8].a/w2889 ), .B(
        \SUBBYTES[8].a/w2892 ), .Z(n15323) );
  XOR \SUBBYTES[8].a/U4847  ( .A(\SUBBYTES[8].a/w2875 ), .B(
        \SUBBYTES[8].a/w2877 ), .Z(n15324) );
  XOR \SUBBYTES[8].a/U4846  ( .A(n15326), .B(n15325), .Z(\SUBBYTES[8].a/w2899 ) );
  XOR \SUBBYTES[8].a/U4845  ( .A(n15963), .B(n15327), .Z(n15325) );
  XOR \SUBBYTES[8].a/U4844  ( .A(\w1[8][21] ), .B(n15964), .Z(n15326) );
  XOR \SUBBYTES[8].a/U4843  ( .A(\SUBBYTES[8].a/w2889 ), .B(
        \SUBBYTES[8].a/w2890 ), .Z(n15327) );
  XOR \SUBBYTES[8].a/U4842  ( .A(n15329), .B(n15328), .Z(\SUBBYTES[8].a/w2915 ) );
  XOR \SUBBYTES[8].a/U4841  ( .A(\w1[8][17] ), .B(n15330), .Z(n15328) );
  XOR \SUBBYTES[8].a/U4840  ( .A(\SUBBYTES[8].a/w2890 ), .B(
        \SUBBYTES[8].a/w2892 ), .Z(n15329) );
  XOR \SUBBYTES[8].a/U4839  ( .A(\SUBBYTES[8].a/w2874 ), .B(
        \SUBBYTES[8].a/w2875 ), .Z(n15330) );
  XOR \SUBBYTES[8].a/U4838  ( .A(\w1[8][25] ), .B(n15331), .Z(n15965) );
  XOR \SUBBYTES[8].a/U4837  ( .A(\w1[8][27] ), .B(\w1[8][26] ), .Z(n15331) );
  XOR \SUBBYTES[8].a/U4836  ( .A(\w1[8][30] ), .B(n15965), .Z(
        \SUBBYTES[8].a/w2757 ) );
  XOR \SUBBYTES[8].a/U4835  ( .A(\w1[8][24] ), .B(\SUBBYTES[8].a/w2757 ), .Z(
        \SUBBYTES[8].a/w2644 ) );
  XOR \SUBBYTES[8].a/U4834  ( .A(\w1[8][24] ), .B(n15332), .Z(
        \SUBBYTES[8].a/w2645 ) );
  XOR \SUBBYTES[8].a/U4833  ( .A(\w1[8][30] ), .B(\w1[8][29] ), .Z(n15332) );
  XOR \SUBBYTES[8].a/U4832  ( .A(\w1[8][29] ), .B(n15965), .Z(
        \SUBBYTES[8].a/w2775 ) );
  XOR \SUBBYTES[8].a/U4831  ( .A(n15334), .B(n15333), .Z(\SUBBYTES[8].a/w2768 ) );
  XOR \SUBBYTES[8].a/U4830  ( .A(\w1[8][27] ), .B(\w1[8][25] ), .Z(n15333) );
  XOR \SUBBYTES[8].a/U4829  ( .A(\w1[8][31] ), .B(\w1[8][28] ), .Z(n15334) );
  XOR \SUBBYTES[8].a/U4828  ( .A(\w1[8][24] ), .B(\SUBBYTES[8].a/w2768 ), .Z(
        \SUBBYTES[8].a/w2647 ) );
  XOR \SUBBYTES[8].a/U4827  ( .A(n15336), .B(n15335), .Z(\SUBBYTES[8].a/w2755 ) );
  XOR \SUBBYTES[8].a/U4826  ( .A(\SUBBYTES[8].a/w2716 ), .B(n1081), .Z(n15335)
         );
  XOR \SUBBYTES[8].a/U4825  ( .A(\SUBBYTES[8].a/w2709 ), .B(
        \SUBBYTES[8].a/w2712 ), .Z(n15336) );
  XOR \SUBBYTES[8].a/U4824  ( .A(n15338), .B(n15337), .Z(\SUBBYTES[8].a/w2756 ) );
  XOR \SUBBYTES[8].a/U4823  ( .A(\SUBBYTES[8].a/w2716 ), .B(n14817), .Z(n15337) );
  XOR \SUBBYTES[8].a/U4822  ( .A(\SUBBYTES[8].a/w2709 ), .B(n14816), .Z(n15338) );
  XOR \SUBBYTES[8].a/U4821  ( .A(\SUBBYTES[8].a/w2768 ), .B(n15339), .Z(
        \SUBBYTES[8].a/w2758 ) );
  XOR \SUBBYTES[8].a/U4820  ( .A(\w1[8][30] ), .B(\w1[8][29] ), .Z(n15339) );
  XOR \SUBBYTES[8].a/U4819  ( .A(n15341), .B(n15340), .Z(\SUBBYTES[8].a/w2759 ) );
  XOR \SUBBYTES[8].a/U4818  ( .A(n14817), .B(n1081), .Z(n15340) );
  XOR \SUBBYTES[8].a/U4817  ( .A(n14816), .B(\SUBBYTES[8].a/w2712 ), .Z(n15341) );
  XOR \SUBBYTES[8].a/U4816  ( .A(\w1[8][31] ), .B(\w1[8][26] ), .Z(n15971) );
  XOR \SUBBYTES[8].a/U4815  ( .A(n15971), .B(n15342), .Z(\SUBBYTES[8].a/w2760 ) );
  XOR \SUBBYTES[8].a/U4814  ( .A(\w1[8][29] ), .B(\w1[8][28] ), .Z(n15342) );
  XOR \SUBBYTES[8].a/U4813  ( .A(\w1[8][31] ), .B(\SUBBYTES[8].a/w2645 ), .Z(
        \SUBBYTES[8].a/w2648 ) );
  XOR \SUBBYTES[8].a/U4812  ( .A(\w1[8][25] ), .B(\SUBBYTES[8].a/w2645 ), .Z(
        \SUBBYTES[8].a/w2649 ) );
  XOR \SUBBYTES[8].a/U4811  ( .A(\w1[8][28] ), .B(\SUBBYTES[8].a/w2645 ), .Z(
        \SUBBYTES[8].a/w2650 ) );
  XOR \SUBBYTES[8].a/U4810  ( .A(\SUBBYTES[8].a/w2649 ), .B(n15971), .Z(
        \SUBBYTES[8].a/w2651 ) );
  XOR \SUBBYTES[8].a/U4809  ( .A(n15971), .B(n15343), .Z(\SUBBYTES[8].a/w2736 ) );
  XOR \SUBBYTES[8].a/U4808  ( .A(\w1[8][28] ), .B(\w1[8][25] ), .Z(n15343) );
  XOR \SUBBYTES[8].a/U4807  ( .A(n15345), .B(n15344), .Z(n15968) );
  XOR \SUBBYTES[8].a/U4806  ( .A(\w1[8][28] ), .B(n15346), .Z(n15344) );
  XOR \SUBBYTES[8].a/U4805  ( .A(\SUBBYTES[8].a/w2701 ), .B(\w1[8][30] ), .Z(
        n15345) );
  XOR \SUBBYTES[8].a/U4804  ( .A(\SUBBYTES[8].a/w2675 ), .B(
        \SUBBYTES[8].a/w2682 ), .Z(n15346) );
  XOR \SUBBYTES[8].a/U4803  ( .A(n15348), .B(n15347), .Z(n15966) );
  XOR \SUBBYTES[8].a/U4802  ( .A(\w1[8][25] ), .B(n15349), .Z(n15347) );
  XOR \SUBBYTES[8].a/U4801  ( .A(\SUBBYTES[8].a/w2700 ), .B(\w1[8][29] ), .Z(
        n15348) );
  XOR \SUBBYTES[8].a/U4800  ( .A(\SUBBYTES[8].a/w2676 ), .B(
        \SUBBYTES[8].a/w2683 ), .Z(n15349) );
  XOR \SUBBYTES[8].a/U4799  ( .A(n15968), .B(n15966), .Z(\SUBBYTES[8].a/w2706 ) );
  XOR \SUBBYTES[8].a/U4798  ( .A(\w1[8][29] ), .B(n15350), .Z(n15969) );
  XOR \SUBBYTES[8].a/U4797  ( .A(\SUBBYTES[8].a/w2668 ), .B(
        \SUBBYTES[8].a/w2678 ), .Z(n15350) );
  XOR \SUBBYTES[8].a/U4796  ( .A(n15352), .B(n15351), .Z(\SUBBYTES[8].a/w2693 ) );
  XOR \SUBBYTES[8].a/U4795  ( .A(n15969), .B(n15353), .Z(n15351) );
  XOR \SUBBYTES[8].a/U4794  ( .A(\w1[8][28] ), .B(\SUBBYTES[8].a/w2757 ), .Z(
        n15352) );
  XOR \SUBBYTES[8].a/U4793  ( .A(\SUBBYTES[8].a/w2670 ), .B(
        \SUBBYTES[8].a/w2675 ), .Z(n15353) );
  XOR \SUBBYTES[8].a/U4792  ( .A(n15355), .B(n15354), .Z(n15967) );
  XOR \SUBBYTES[8].a/U4791  ( .A(\SUBBYTES[8].a/w2703 ), .B(\w1[8][31] ), .Z(
        n15354) );
  XOR \SUBBYTES[8].a/U4790  ( .A(\SUBBYTES[8].a/w2678 ), .B(
        \SUBBYTES[8].a/w2685 ), .Z(n15355) );
  XOR \SUBBYTES[8].a/U4789  ( .A(n15966), .B(n15967), .Z(\SUBBYTES[8].a/w2705 ) );
  XOR \SUBBYTES[8].a/U4788  ( .A(\w1[8][27] ), .B(n15356), .Z(n15970) );
  XOR \SUBBYTES[8].a/U4787  ( .A(\SUBBYTES[8].a/w2667 ), .B(
        \SUBBYTES[8].a/w2670 ), .Z(n15356) );
  XOR \SUBBYTES[8].a/U4786  ( .A(n15358), .B(n15357), .Z(\SUBBYTES[8].a/w2694 ) );
  XOR \SUBBYTES[8].a/U4785  ( .A(n15970), .B(n15359), .Z(n15357) );
  XOR \SUBBYTES[8].a/U4784  ( .A(\w1[8][30] ), .B(\SUBBYTES[8].a/w2736 ), .Z(
        n15358) );
  XOR \SUBBYTES[8].a/U4783  ( .A(\SUBBYTES[8].a/w2675 ), .B(
        \SUBBYTES[8].a/w2676 ), .Z(n15359) );
  XOR \SUBBYTES[8].a/U4782  ( .A(n15968), .B(n15967), .Z(\SUBBYTES[8].a/w2714 ) );
  XOR \SUBBYTES[8].a/U4781  ( .A(n15361), .B(n15360), .Z(\SUBBYTES[8].a/w2715 ) );
  XOR \SUBBYTES[8].a/U4780  ( .A(\w1[8][31] ), .B(n15969), .Z(n15360) );
  XOR \SUBBYTES[8].a/U4779  ( .A(\SUBBYTES[8].a/w2667 ), .B(
        \SUBBYTES[8].a/w2676 ), .Z(n15361) );
  XOR \SUBBYTES[8].a/U4778  ( .A(n15363), .B(n15362), .Z(\SUBBYTES[8].a/w2691 ) );
  XOR \SUBBYTES[8].a/U4777  ( .A(n15365), .B(n15364), .Z(n15362) );
  XOR \SUBBYTES[8].a/U4776  ( .A(\w1[8][31] ), .B(\SUBBYTES[8].a/w2775 ), .Z(
        n15363) );
  XOR \SUBBYTES[8].a/U4775  ( .A(\SUBBYTES[8].a/w2682 ), .B(
        \SUBBYTES[8].a/w2685 ), .Z(n15364) );
  XOR \SUBBYTES[8].a/U4774  ( .A(\SUBBYTES[8].a/w2668 ), .B(
        \SUBBYTES[8].a/w2670 ), .Z(n15365) );
  XOR \SUBBYTES[8].a/U4773  ( .A(n15367), .B(n15366), .Z(\SUBBYTES[8].a/w2692 ) );
  XOR \SUBBYTES[8].a/U4772  ( .A(n15970), .B(n15368), .Z(n15366) );
  XOR \SUBBYTES[8].a/U4771  ( .A(\w1[8][29] ), .B(n15971), .Z(n15367) );
  XOR \SUBBYTES[8].a/U4770  ( .A(\SUBBYTES[8].a/w2682 ), .B(
        \SUBBYTES[8].a/w2683 ), .Z(n15368) );
  XOR \SUBBYTES[8].a/U4769  ( .A(n15370), .B(n15369), .Z(\SUBBYTES[8].a/w2708 ) );
  XOR \SUBBYTES[8].a/U4768  ( .A(\w1[8][25] ), .B(n15371), .Z(n15369) );
  XOR \SUBBYTES[8].a/U4767  ( .A(\SUBBYTES[8].a/w2683 ), .B(
        \SUBBYTES[8].a/w2685 ), .Z(n15370) );
  XOR \SUBBYTES[8].a/U4766  ( .A(\SUBBYTES[8].a/w2667 ), .B(
        \SUBBYTES[8].a/w2668 ), .Z(n15371) );
  XOR \SUBBYTES[8].a/U4765  ( .A(\w1[8][33] ), .B(n15372), .Z(n15972) );
  XOR \SUBBYTES[8].a/U4764  ( .A(\w1[8][35] ), .B(\w1[8][34] ), .Z(n15372) );
  XOR \SUBBYTES[8].a/U4763  ( .A(\w1[8][38] ), .B(n15972), .Z(
        \SUBBYTES[8].a/w2550 ) );
  XOR \SUBBYTES[8].a/U4762  ( .A(\w1[8][32] ), .B(\SUBBYTES[8].a/w2550 ), .Z(
        \SUBBYTES[8].a/w2437 ) );
  XOR \SUBBYTES[8].a/U4761  ( .A(\w1[8][32] ), .B(n15373), .Z(
        \SUBBYTES[8].a/w2438 ) );
  XOR \SUBBYTES[8].a/U4760  ( .A(\w1[8][38] ), .B(\w1[8][37] ), .Z(n15373) );
  XOR \SUBBYTES[8].a/U4759  ( .A(\w1[8][37] ), .B(n15972), .Z(
        \SUBBYTES[8].a/w2568 ) );
  XOR \SUBBYTES[8].a/U4758  ( .A(n15375), .B(n15374), .Z(\SUBBYTES[8].a/w2561 ) );
  XOR \SUBBYTES[8].a/U4757  ( .A(\w1[8][35] ), .B(\w1[8][33] ), .Z(n15374) );
  XOR \SUBBYTES[8].a/U4756  ( .A(\w1[8][39] ), .B(\w1[8][36] ), .Z(n15375) );
  XOR \SUBBYTES[8].a/U4755  ( .A(\w1[8][32] ), .B(\SUBBYTES[8].a/w2561 ), .Z(
        \SUBBYTES[8].a/w2440 ) );
  XOR \SUBBYTES[8].a/U4754  ( .A(n15377), .B(n15376), .Z(\SUBBYTES[8].a/w2548 ) );
  XOR \SUBBYTES[8].a/U4753  ( .A(\SUBBYTES[8].a/w2509 ), .B(n1080), .Z(n15376)
         );
  XOR \SUBBYTES[8].a/U4752  ( .A(\SUBBYTES[8].a/w2502 ), .B(
        \SUBBYTES[8].a/w2505 ), .Z(n15377) );
  XOR \SUBBYTES[8].a/U4751  ( .A(n15379), .B(n15378), .Z(\SUBBYTES[8].a/w2549 ) );
  XOR \SUBBYTES[8].a/U4750  ( .A(\SUBBYTES[8].a/w2509 ), .B(n14815), .Z(n15378) );
  XOR \SUBBYTES[8].a/U4749  ( .A(\SUBBYTES[8].a/w2502 ), .B(n14814), .Z(n15379) );
  XOR \SUBBYTES[8].a/U4748  ( .A(\SUBBYTES[8].a/w2561 ), .B(n15380), .Z(
        \SUBBYTES[8].a/w2551 ) );
  XOR \SUBBYTES[8].a/U4747  ( .A(\w1[8][38] ), .B(\w1[8][37] ), .Z(n15380) );
  XOR \SUBBYTES[8].a/U4746  ( .A(n15382), .B(n15381), .Z(\SUBBYTES[8].a/w2552 ) );
  XOR \SUBBYTES[8].a/U4745  ( .A(n14815), .B(n1080), .Z(n15381) );
  XOR \SUBBYTES[8].a/U4744  ( .A(n14814), .B(\SUBBYTES[8].a/w2505 ), .Z(n15382) );
  XOR \SUBBYTES[8].a/U4743  ( .A(\w1[8][39] ), .B(\w1[8][34] ), .Z(n15978) );
  XOR \SUBBYTES[8].a/U4742  ( .A(n15978), .B(n15383), .Z(\SUBBYTES[8].a/w2553 ) );
  XOR \SUBBYTES[8].a/U4741  ( .A(\w1[8][37] ), .B(\w1[8][36] ), .Z(n15383) );
  XOR \SUBBYTES[8].a/U4740  ( .A(\w1[8][39] ), .B(\SUBBYTES[8].a/w2438 ), .Z(
        \SUBBYTES[8].a/w2441 ) );
  XOR \SUBBYTES[8].a/U4739  ( .A(\w1[8][33] ), .B(\SUBBYTES[8].a/w2438 ), .Z(
        \SUBBYTES[8].a/w2442 ) );
  XOR \SUBBYTES[8].a/U4738  ( .A(\w1[8][36] ), .B(\SUBBYTES[8].a/w2438 ), .Z(
        \SUBBYTES[8].a/w2443 ) );
  XOR \SUBBYTES[8].a/U4737  ( .A(\SUBBYTES[8].a/w2442 ), .B(n15978), .Z(
        \SUBBYTES[8].a/w2444 ) );
  XOR \SUBBYTES[8].a/U4736  ( .A(n15978), .B(n15384), .Z(\SUBBYTES[8].a/w2529 ) );
  XOR \SUBBYTES[8].a/U4735  ( .A(\w1[8][36] ), .B(\w1[8][33] ), .Z(n15384) );
  XOR \SUBBYTES[8].a/U4734  ( .A(n15386), .B(n15385), .Z(n15975) );
  XOR \SUBBYTES[8].a/U4733  ( .A(\w1[8][36] ), .B(n15387), .Z(n15385) );
  XOR \SUBBYTES[8].a/U4732  ( .A(\SUBBYTES[8].a/w2494 ), .B(\w1[8][38] ), .Z(
        n15386) );
  XOR \SUBBYTES[8].a/U4731  ( .A(\SUBBYTES[8].a/w2468 ), .B(
        \SUBBYTES[8].a/w2475 ), .Z(n15387) );
  XOR \SUBBYTES[8].a/U4730  ( .A(n15389), .B(n15388), .Z(n15973) );
  XOR \SUBBYTES[8].a/U4729  ( .A(\w1[8][33] ), .B(n15390), .Z(n15388) );
  XOR \SUBBYTES[8].a/U4728  ( .A(\SUBBYTES[8].a/w2493 ), .B(\w1[8][37] ), .Z(
        n15389) );
  XOR \SUBBYTES[8].a/U4727  ( .A(\SUBBYTES[8].a/w2469 ), .B(
        \SUBBYTES[8].a/w2476 ), .Z(n15390) );
  XOR \SUBBYTES[8].a/U4726  ( .A(n15975), .B(n15973), .Z(\SUBBYTES[8].a/w2499 ) );
  XOR \SUBBYTES[8].a/U4725  ( .A(\w1[8][37] ), .B(n15391), .Z(n15976) );
  XOR \SUBBYTES[8].a/U4724  ( .A(\SUBBYTES[8].a/w2461 ), .B(
        \SUBBYTES[8].a/w2471 ), .Z(n15391) );
  XOR \SUBBYTES[8].a/U4723  ( .A(n15393), .B(n15392), .Z(\SUBBYTES[8].a/w2486 ) );
  XOR \SUBBYTES[8].a/U4722  ( .A(n15976), .B(n15394), .Z(n15392) );
  XOR \SUBBYTES[8].a/U4721  ( .A(\w1[8][36] ), .B(\SUBBYTES[8].a/w2550 ), .Z(
        n15393) );
  XOR \SUBBYTES[8].a/U4720  ( .A(\SUBBYTES[8].a/w2463 ), .B(
        \SUBBYTES[8].a/w2468 ), .Z(n15394) );
  XOR \SUBBYTES[8].a/U4719  ( .A(n15396), .B(n15395), .Z(n15974) );
  XOR \SUBBYTES[8].a/U4718  ( .A(\SUBBYTES[8].a/w2496 ), .B(\w1[8][39] ), .Z(
        n15395) );
  XOR \SUBBYTES[8].a/U4717  ( .A(\SUBBYTES[8].a/w2471 ), .B(
        \SUBBYTES[8].a/w2478 ), .Z(n15396) );
  XOR \SUBBYTES[8].a/U4716  ( .A(n15973), .B(n15974), .Z(\SUBBYTES[8].a/w2498 ) );
  XOR \SUBBYTES[8].a/U4715  ( .A(\w1[8][35] ), .B(n15397), .Z(n15977) );
  XOR \SUBBYTES[8].a/U4714  ( .A(\SUBBYTES[8].a/w2460 ), .B(
        \SUBBYTES[8].a/w2463 ), .Z(n15397) );
  XOR \SUBBYTES[8].a/U4713  ( .A(n15399), .B(n15398), .Z(\SUBBYTES[8].a/w2487 ) );
  XOR \SUBBYTES[8].a/U4712  ( .A(n15977), .B(n15400), .Z(n15398) );
  XOR \SUBBYTES[8].a/U4711  ( .A(\w1[8][38] ), .B(\SUBBYTES[8].a/w2529 ), .Z(
        n15399) );
  XOR \SUBBYTES[8].a/U4710  ( .A(\SUBBYTES[8].a/w2468 ), .B(
        \SUBBYTES[8].a/w2469 ), .Z(n15400) );
  XOR \SUBBYTES[8].a/U4709  ( .A(n15975), .B(n15974), .Z(\SUBBYTES[8].a/w2507 ) );
  XOR \SUBBYTES[8].a/U4708  ( .A(n15402), .B(n15401), .Z(\SUBBYTES[8].a/w2508 ) );
  XOR \SUBBYTES[8].a/U4707  ( .A(\w1[8][39] ), .B(n15976), .Z(n15401) );
  XOR \SUBBYTES[8].a/U4706  ( .A(\SUBBYTES[8].a/w2460 ), .B(
        \SUBBYTES[8].a/w2469 ), .Z(n15402) );
  XOR \SUBBYTES[8].a/U4705  ( .A(n15404), .B(n15403), .Z(\SUBBYTES[8].a/w2484 ) );
  XOR \SUBBYTES[8].a/U4704  ( .A(n15406), .B(n15405), .Z(n15403) );
  XOR \SUBBYTES[8].a/U4703  ( .A(\w1[8][39] ), .B(\SUBBYTES[8].a/w2568 ), .Z(
        n15404) );
  XOR \SUBBYTES[8].a/U4702  ( .A(\SUBBYTES[8].a/w2475 ), .B(
        \SUBBYTES[8].a/w2478 ), .Z(n15405) );
  XOR \SUBBYTES[8].a/U4701  ( .A(\SUBBYTES[8].a/w2461 ), .B(
        \SUBBYTES[8].a/w2463 ), .Z(n15406) );
  XOR \SUBBYTES[8].a/U4700  ( .A(n15408), .B(n15407), .Z(\SUBBYTES[8].a/w2485 ) );
  XOR \SUBBYTES[8].a/U4699  ( .A(n15977), .B(n15409), .Z(n15407) );
  XOR \SUBBYTES[8].a/U4698  ( .A(\w1[8][37] ), .B(n15978), .Z(n15408) );
  XOR \SUBBYTES[8].a/U4697  ( .A(\SUBBYTES[8].a/w2475 ), .B(
        \SUBBYTES[8].a/w2476 ), .Z(n15409) );
  XOR \SUBBYTES[8].a/U4696  ( .A(n15411), .B(n15410), .Z(\SUBBYTES[8].a/w2501 ) );
  XOR \SUBBYTES[8].a/U4695  ( .A(\w1[8][33] ), .B(n15412), .Z(n15410) );
  XOR \SUBBYTES[8].a/U4694  ( .A(\SUBBYTES[8].a/w2476 ), .B(
        \SUBBYTES[8].a/w2478 ), .Z(n15411) );
  XOR \SUBBYTES[8].a/U4693  ( .A(\SUBBYTES[8].a/w2460 ), .B(
        \SUBBYTES[8].a/w2461 ), .Z(n15412) );
  XOR \SUBBYTES[8].a/U4692  ( .A(\w1[8][41] ), .B(n15413), .Z(n15979) );
  XOR \SUBBYTES[8].a/U4691  ( .A(\w1[8][43] ), .B(\w1[8][42] ), .Z(n15413) );
  XOR \SUBBYTES[8].a/U4690  ( .A(\w1[8][46] ), .B(n15979), .Z(
        \SUBBYTES[8].a/w2343 ) );
  XOR \SUBBYTES[8].a/U4689  ( .A(\w1[8][40] ), .B(\SUBBYTES[8].a/w2343 ), .Z(
        \SUBBYTES[8].a/w2230 ) );
  XOR \SUBBYTES[8].a/U4688  ( .A(\w1[8][40] ), .B(n15414), .Z(
        \SUBBYTES[8].a/w2231 ) );
  XOR \SUBBYTES[8].a/U4687  ( .A(\w1[8][46] ), .B(\w1[8][45] ), .Z(n15414) );
  XOR \SUBBYTES[8].a/U4686  ( .A(\w1[8][45] ), .B(n15979), .Z(
        \SUBBYTES[8].a/w2361 ) );
  XOR \SUBBYTES[8].a/U4685  ( .A(n15416), .B(n15415), .Z(\SUBBYTES[8].a/w2354 ) );
  XOR \SUBBYTES[8].a/U4684  ( .A(\w1[8][43] ), .B(\w1[8][41] ), .Z(n15415) );
  XOR \SUBBYTES[8].a/U4683  ( .A(\w1[8][47] ), .B(\w1[8][44] ), .Z(n15416) );
  XOR \SUBBYTES[8].a/U4682  ( .A(\w1[8][40] ), .B(\SUBBYTES[8].a/w2354 ), .Z(
        \SUBBYTES[8].a/w2233 ) );
  XOR \SUBBYTES[8].a/U4681  ( .A(n15418), .B(n15417), .Z(\SUBBYTES[8].a/w2341 ) );
  XOR \SUBBYTES[8].a/U4680  ( .A(\SUBBYTES[8].a/w2302 ), .B(n1079), .Z(n15417)
         );
  XOR \SUBBYTES[8].a/U4679  ( .A(\SUBBYTES[8].a/w2295 ), .B(
        \SUBBYTES[8].a/w2298 ), .Z(n15418) );
  XOR \SUBBYTES[8].a/U4678  ( .A(n15420), .B(n15419), .Z(\SUBBYTES[8].a/w2342 ) );
  XOR \SUBBYTES[8].a/U4677  ( .A(\SUBBYTES[8].a/w2302 ), .B(n14813), .Z(n15419) );
  XOR \SUBBYTES[8].a/U4676  ( .A(\SUBBYTES[8].a/w2295 ), .B(n14812), .Z(n15420) );
  XOR \SUBBYTES[8].a/U4675  ( .A(\SUBBYTES[8].a/w2354 ), .B(n15421), .Z(
        \SUBBYTES[8].a/w2344 ) );
  XOR \SUBBYTES[8].a/U4674  ( .A(\w1[8][46] ), .B(\w1[8][45] ), .Z(n15421) );
  XOR \SUBBYTES[8].a/U4673  ( .A(n15423), .B(n15422), .Z(\SUBBYTES[8].a/w2345 ) );
  XOR \SUBBYTES[8].a/U4672  ( .A(n14813), .B(n1079), .Z(n15422) );
  XOR \SUBBYTES[8].a/U4671  ( .A(n14812), .B(\SUBBYTES[8].a/w2298 ), .Z(n15423) );
  XOR \SUBBYTES[8].a/U4670  ( .A(\w1[8][47] ), .B(\w1[8][42] ), .Z(n15985) );
  XOR \SUBBYTES[8].a/U4669  ( .A(n15985), .B(n15424), .Z(\SUBBYTES[8].a/w2346 ) );
  XOR \SUBBYTES[8].a/U4668  ( .A(\w1[8][45] ), .B(\w1[8][44] ), .Z(n15424) );
  XOR \SUBBYTES[8].a/U4667  ( .A(\w1[8][47] ), .B(\SUBBYTES[8].a/w2231 ), .Z(
        \SUBBYTES[8].a/w2234 ) );
  XOR \SUBBYTES[8].a/U4666  ( .A(\w1[8][41] ), .B(\SUBBYTES[8].a/w2231 ), .Z(
        \SUBBYTES[8].a/w2235 ) );
  XOR \SUBBYTES[8].a/U4665  ( .A(\w1[8][44] ), .B(\SUBBYTES[8].a/w2231 ), .Z(
        \SUBBYTES[8].a/w2236 ) );
  XOR \SUBBYTES[8].a/U4664  ( .A(\SUBBYTES[8].a/w2235 ), .B(n15985), .Z(
        \SUBBYTES[8].a/w2237 ) );
  XOR \SUBBYTES[8].a/U4663  ( .A(n15985), .B(n15425), .Z(\SUBBYTES[8].a/w2322 ) );
  XOR \SUBBYTES[8].a/U4662  ( .A(\w1[8][44] ), .B(\w1[8][41] ), .Z(n15425) );
  XOR \SUBBYTES[8].a/U4661  ( .A(n15427), .B(n15426), .Z(n15982) );
  XOR \SUBBYTES[8].a/U4660  ( .A(\w1[8][44] ), .B(n15428), .Z(n15426) );
  XOR \SUBBYTES[8].a/U4659  ( .A(\SUBBYTES[8].a/w2287 ), .B(\w1[8][46] ), .Z(
        n15427) );
  XOR \SUBBYTES[8].a/U4658  ( .A(\SUBBYTES[8].a/w2261 ), .B(
        \SUBBYTES[8].a/w2268 ), .Z(n15428) );
  XOR \SUBBYTES[8].a/U4657  ( .A(n15430), .B(n15429), .Z(n15980) );
  XOR \SUBBYTES[8].a/U4656  ( .A(\w1[8][41] ), .B(n15431), .Z(n15429) );
  XOR \SUBBYTES[8].a/U4655  ( .A(\SUBBYTES[8].a/w2286 ), .B(\w1[8][45] ), .Z(
        n15430) );
  XOR \SUBBYTES[8].a/U4654  ( .A(\SUBBYTES[8].a/w2262 ), .B(
        \SUBBYTES[8].a/w2269 ), .Z(n15431) );
  XOR \SUBBYTES[8].a/U4653  ( .A(n15982), .B(n15980), .Z(\SUBBYTES[8].a/w2292 ) );
  XOR \SUBBYTES[8].a/U4652  ( .A(\w1[8][45] ), .B(n15432), .Z(n15983) );
  XOR \SUBBYTES[8].a/U4651  ( .A(\SUBBYTES[8].a/w2254 ), .B(
        \SUBBYTES[8].a/w2264 ), .Z(n15432) );
  XOR \SUBBYTES[8].a/U4650  ( .A(n15434), .B(n15433), .Z(\SUBBYTES[8].a/w2279 ) );
  XOR \SUBBYTES[8].a/U4649  ( .A(n15983), .B(n15435), .Z(n15433) );
  XOR \SUBBYTES[8].a/U4648  ( .A(\w1[8][44] ), .B(\SUBBYTES[8].a/w2343 ), .Z(
        n15434) );
  XOR \SUBBYTES[8].a/U4647  ( .A(\SUBBYTES[8].a/w2256 ), .B(
        \SUBBYTES[8].a/w2261 ), .Z(n15435) );
  XOR \SUBBYTES[8].a/U4646  ( .A(n15437), .B(n15436), .Z(n15981) );
  XOR \SUBBYTES[8].a/U4645  ( .A(\SUBBYTES[8].a/w2289 ), .B(\w1[8][47] ), .Z(
        n15436) );
  XOR \SUBBYTES[8].a/U4644  ( .A(\SUBBYTES[8].a/w2264 ), .B(
        \SUBBYTES[8].a/w2271 ), .Z(n15437) );
  XOR \SUBBYTES[8].a/U4643  ( .A(n15980), .B(n15981), .Z(\SUBBYTES[8].a/w2291 ) );
  XOR \SUBBYTES[8].a/U4642  ( .A(\w1[8][43] ), .B(n15438), .Z(n15984) );
  XOR \SUBBYTES[8].a/U4641  ( .A(\SUBBYTES[8].a/w2253 ), .B(
        \SUBBYTES[8].a/w2256 ), .Z(n15438) );
  XOR \SUBBYTES[8].a/U4640  ( .A(n15440), .B(n15439), .Z(\SUBBYTES[8].a/w2280 ) );
  XOR \SUBBYTES[8].a/U4639  ( .A(n15984), .B(n15441), .Z(n15439) );
  XOR \SUBBYTES[8].a/U4638  ( .A(\w1[8][46] ), .B(\SUBBYTES[8].a/w2322 ), .Z(
        n15440) );
  XOR \SUBBYTES[8].a/U4637  ( .A(\SUBBYTES[8].a/w2261 ), .B(
        \SUBBYTES[8].a/w2262 ), .Z(n15441) );
  XOR \SUBBYTES[8].a/U4636  ( .A(n15982), .B(n15981), .Z(\SUBBYTES[8].a/w2300 ) );
  XOR \SUBBYTES[8].a/U4635  ( .A(n15443), .B(n15442), .Z(\SUBBYTES[8].a/w2301 ) );
  XOR \SUBBYTES[8].a/U4634  ( .A(\w1[8][47] ), .B(n15983), .Z(n15442) );
  XOR \SUBBYTES[8].a/U4633  ( .A(\SUBBYTES[8].a/w2253 ), .B(
        \SUBBYTES[8].a/w2262 ), .Z(n15443) );
  XOR \SUBBYTES[8].a/U4632  ( .A(n15445), .B(n15444), .Z(\SUBBYTES[8].a/w2277 ) );
  XOR \SUBBYTES[8].a/U4631  ( .A(n15447), .B(n15446), .Z(n15444) );
  XOR \SUBBYTES[8].a/U4630  ( .A(\w1[8][47] ), .B(\SUBBYTES[8].a/w2361 ), .Z(
        n15445) );
  XOR \SUBBYTES[8].a/U4629  ( .A(\SUBBYTES[8].a/w2268 ), .B(
        \SUBBYTES[8].a/w2271 ), .Z(n15446) );
  XOR \SUBBYTES[8].a/U4628  ( .A(\SUBBYTES[8].a/w2254 ), .B(
        \SUBBYTES[8].a/w2256 ), .Z(n15447) );
  XOR \SUBBYTES[8].a/U4627  ( .A(n15449), .B(n15448), .Z(\SUBBYTES[8].a/w2278 ) );
  XOR \SUBBYTES[8].a/U4626  ( .A(n15984), .B(n15450), .Z(n15448) );
  XOR \SUBBYTES[8].a/U4625  ( .A(\w1[8][45] ), .B(n15985), .Z(n15449) );
  XOR \SUBBYTES[8].a/U4624  ( .A(\SUBBYTES[8].a/w2268 ), .B(
        \SUBBYTES[8].a/w2269 ), .Z(n15450) );
  XOR \SUBBYTES[8].a/U4623  ( .A(n15452), .B(n15451), .Z(\SUBBYTES[8].a/w2294 ) );
  XOR \SUBBYTES[8].a/U4622  ( .A(\w1[8][41] ), .B(n15453), .Z(n15451) );
  XOR \SUBBYTES[8].a/U4621  ( .A(\SUBBYTES[8].a/w2269 ), .B(
        \SUBBYTES[8].a/w2271 ), .Z(n15452) );
  XOR \SUBBYTES[8].a/U4620  ( .A(\SUBBYTES[8].a/w2253 ), .B(
        \SUBBYTES[8].a/w2254 ), .Z(n15453) );
  XOR \SUBBYTES[8].a/U4619  ( .A(\w1[8][49] ), .B(n15454), .Z(n15986) );
  XOR \SUBBYTES[8].a/U4618  ( .A(\w1[8][51] ), .B(\w1[8][50] ), .Z(n15454) );
  XOR \SUBBYTES[8].a/U4617  ( .A(\w1[8][54] ), .B(n15986), .Z(
        \SUBBYTES[8].a/w2136 ) );
  XOR \SUBBYTES[8].a/U4616  ( .A(\w1[8][48] ), .B(\SUBBYTES[8].a/w2136 ), .Z(
        \SUBBYTES[8].a/w2023 ) );
  XOR \SUBBYTES[8].a/U4615  ( .A(\w1[8][48] ), .B(n15455), .Z(
        \SUBBYTES[8].a/w2024 ) );
  XOR \SUBBYTES[8].a/U4614  ( .A(\w1[8][54] ), .B(\w1[8][53] ), .Z(n15455) );
  XOR \SUBBYTES[8].a/U4613  ( .A(\w1[8][53] ), .B(n15986), .Z(
        \SUBBYTES[8].a/w2154 ) );
  XOR \SUBBYTES[8].a/U4612  ( .A(n15457), .B(n15456), .Z(\SUBBYTES[8].a/w2147 ) );
  XOR \SUBBYTES[8].a/U4611  ( .A(\w1[8][51] ), .B(\w1[8][49] ), .Z(n15456) );
  XOR \SUBBYTES[8].a/U4610  ( .A(\w1[8][55] ), .B(\w1[8][52] ), .Z(n15457) );
  XOR \SUBBYTES[8].a/U4609  ( .A(\w1[8][48] ), .B(\SUBBYTES[8].a/w2147 ), .Z(
        \SUBBYTES[8].a/w2026 ) );
  XOR \SUBBYTES[8].a/U4608  ( .A(n15459), .B(n15458), .Z(\SUBBYTES[8].a/w2134 ) );
  XOR \SUBBYTES[8].a/U4607  ( .A(\SUBBYTES[8].a/w2095 ), .B(n1078), .Z(n15458)
         );
  XOR \SUBBYTES[8].a/U4606  ( .A(\SUBBYTES[8].a/w2088 ), .B(
        \SUBBYTES[8].a/w2091 ), .Z(n15459) );
  XOR \SUBBYTES[8].a/U4605  ( .A(n15461), .B(n15460), .Z(\SUBBYTES[8].a/w2135 ) );
  XOR \SUBBYTES[8].a/U4604  ( .A(\SUBBYTES[8].a/w2095 ), .B(n14811), .Z(n15460) );
  XOR \SUBBYTES[8].a/U4603  ( .A(\SUBBYTES[8].a/w2088 ), .B(n14810), .Z(n15461) );
  XOR \SUBBYTES[8].a/U4602  ( .A(\SUBBYTES[8].a/w2147 ), .B(n15462), .Z(
        \SUBBYTES[8].a/w2137 ) );
  XOR \SUBBYTES[8].a/U4601  ( .A(\w1[8][54] ), .B(\w1[8][53] ), .Z(n15462) );
  XOR \SUBBYTES[8].a/U4600  ( .A(n15464), .B(n15463), .Z(\SUBBYTES[8].a/w2138 ) );
  XOR \SUBBYTES[8].a/U4599  ( .A(n14811), .B(n1078), .Z(n15463) );
  XOR \SUBBYTES[8].a/U4598  ( .A(n14810), .B(\SUBBYTES[8].a/w2091 ), .Z(n15464) );
  XOR \SUBBYTES[8].a/U4597  ( .A(\w1[8][55] ), .B(\w1[8][50] ), .Z(n15992) );
  XOR \SUBBYTES[8].a/U4596  ( .A(n15992), .B(n15465), .Z(\SUBBYTES[8].a/w2139 ) );
  XOR \SUBBYTES[8].a/U4595  ( .A(\w1[8][53] ), .B(\w1[8][52] ), .Z(n15465) );
  XOR \SUBBYTES[8].a/U4594  ( .A(\w1[8][55] ), .B(\SUBBYTES[8].a/w2024 ), .Z(
        \SUBBYTES[8].a/w2027 ) );
  XOR \SUBBYTES[8].a/U4593  ( .A(\w1[8][49] ), .B(\SUBBYTES[8].a/w2024 ), .Z(
        \SUBBYTES[8].a/w2028 ) );
  XOR \SUBBYTES[8].a/U4592  ( .A(\w1[8][52] ), .B(\SUBBYTES[8].a/w2024 ), .Z(
        \SUBBYTES[8].a/w2029 ) );
  XOR \SUBBYTES[8].a/U4591  ( .A(\SUBBYTES[8].a/w2028 ), .B(n15992), .Z(
        \SUBBYTES[8].a/w2030 ) );
  XOR \SUBBYTES[8].a/U4590  ( .A(n15992), .B(n15466), .Z(\SUBBYTES[8].a/w2115 ) );
  XOR \SUBBYTES[8].a/U4589  ( .A(\w1[8][52] ), .B(\w1[8][49] ), .Z(n15466) );
  XOR \SUBBYTES[8].a/U4588  ( .A(n15468), .B(n15467), .Z(n15989) );
  XOR \SUBBYTES[8].a/U4587  ( .A(\w1[8][52] ), .B(n15469), .Z(n15467) );
  XOR \SUBBYTES[8].a/U4586  ( .A(\SUBBYTES[8].a/w2080 ), .B(\w1[8][54] ), .Z(
        n15468) );
  XOR \SUBBYTES[8].a/U4585  ( .A(\SUBBYTES[8].a/w2054 ), .B(
        \SUBBYTES[8].a/w2061 ), .Z(n15469) );
  XOR \SUBBYTES[8].a/U4584  ( .A(n15471), .B(n15470), .Z(n15987) );
  XOR \SUBBYTES[8].a/U4583  ( .A(\w1[8][49] ), .B(n15472), .Z(n15470) );
  XOR \SUBBYTES[8].a/U4582  ( .A(\SUBBYTES[8].a/w2079 ), .B(\w1[8][53] ), .Z(
        n15471) );
  XOR \SUBBYTES[8].a/U4581  ( .A(\SUBBYTES[8].a/w2055 ), .B(
        \SUBBYTES[8].a/w2062 ), .Z(n15472) );
  XOR \SUBBYTES[8].a/U4580  ( .A(n15989), .B(n15987), .Z(\SUBBYTES[8].a/w2085 ) );
  XOR \SUBBYTES[8].a/U4579  ( .A(\w1[8][53] ), .B(n15473), .Z(n15990) );
  XOR \SUBBYTES[8].a/U4578  ( .A(\SUBBYTES[8].a/w2047 ), .B(
        \SUBBYTES[8].a/w2057 ), .Z(n15473) );
  XOR \SUBBYTES[8].a/U4577  ( .A(n15475), .B(n15474), .Z(\SUBBYTES[8].a/w2072 ) );
  XOR \SUBBYTES[8].a/U4576  ( .A(n15990), .B(n15476), .Z(n15474) );
  XOR \SUBBYTES[8].a/U4575  ( .A(\w1[8][52] ), .B(\SUBBYTES[8].a/w2136 ), .Z(
        n15475) );
  XOR \SUBBYTES[8].a/U4574  ( .A(\SUBBYTES[8].a/w2049 ), .B(
        \SUBBYTES[8].a/w2054 ), .Z(n15476) );
  XOR \SUBBYTES[8].a/U4573  ( .A(n15478), .B(n15477), .Z(n15988) );
  XOR \SUBBYTES[8].a/U4572  ( .A(\SUBBYTES[8].a/w2082 ), .B(\w1[8][55] ), .Z(
        n15477) );
  XOR \SUBBYTES[8].a/U4571  ( .A(\SUBBYTES[8].a/w2057 ), .B(
        \SUBBYTES[8].a/w2064 ), .Z(n15478) );
  XOR \SUBBYTES[8].a/U4570  ( .A(n15987), .B(n15988), .Z(\SUBBYTES[8].a/w2084 ) );
  XOR \SUBBYTES[8].a/U4569  ( .A(\w1[8][51] ), .B(n15479), .Z(n15991) );
  XOR \SUBBYTES[8].a/U4568  ( .A(\SUBBYTES[8].a/w2046 ), .B(
        \SUBBYTES[8].a/w2049 ), .Z(n15479) );
  XOR \SUBBYTES[8].a/U4567  ( .A(n15481), .B(n15480), .Z(\SUBBYTES[8].a/w2073 ) );
  XOR \SUBBYTES[8].a/U4566  ( .A(n15991), .B(n15482), .Z(n15480) );
  XOR \SUBBYTES[8].a/U4565  ( .A(\w1[8][54] ), .B(\SUBBYTES[8].a/w2115 ), .Z(
        n15481) );
  XOR \SUBBYTES[8].a/U4564  ( .A(\SUBBYTES[8].a/w2054 ), .B(
        \SUBBYTES[8].a/w2055 ), .Z(n15482) );
  XOR \SUBBYTES[8].a/U4563  ( .A(n15989), .B(n15988), .Z(\SUBBYTES[8].a/w2093 ) );
  XOR \SUBBYTES[8].a/U4562  ( .A(n15484), .B(n15483), .Z(\SUBBYTES[8].a/w2094 ) );
  XOR \SUBBYTES[8].a/U4561  ( .A(\w1[8][55] ), .B(n15990), .Z(n15483) );
  XOR \SUBBYTES[8].a/U4560  ( .A(\SUBBYTES[8].a/w2046 ), .B(
        \SUBBYTES[8].a/w2055 ), .Z(n15484) );
  XOR \SUBBYTES[8].a/U4559  ( .A(n15486), .B(n15485), .Z(\SUBBYTES[8].a/w2070 ) );
  XOR \SUBBYTES[8].a/U4558  ( .A(n15488), .B(n15487), .Z(n15485) );
  XOR \SUBBYTES[8].a/U4557  ( .A(\w1[8][55] ), .B(\SUBBYTES[8].a/w2154 ), .Z(
        n15486) );
  XOR \SUBBYTES[8].a/U4556  ( .A(\SUBBYTES[8].a/w2061 ), .B(
        \SUBBYTES[8].a/w2064 ), .Z(n15487) );
  XOR \SUBBYTES[8].a/U4555  ( .A(\SUBBYTES[8].a/w2047 ), .B(
        \SUBBYTES[8].a/w2049 ), .Z(n15488) );
  XOR \SUBBYTES[8].a/U4554  ( .A(n15490), .B(n15489), .Z(\SUBBYTES[8].a/w2071 ) );
  XOR \SUBBYTES[8].a/U4553  ( .A(n15991), .B(n15491), .Z(n15489) );
  XOR \SUBBYTES[8].a/U4552  ( .A(\w1[8][53] ), .B(n15992), .Z(n15490) );
  XOR \SUBBYTES[8].a/U4551  ( .A(\SUBBYTES[8].a/w2061 ), .B(
        \SUBBYTES[8].a/w2062 ), .Z(n15491) );
  XOR \SUBBYTES[8].a/U4550  ( .A(n15493), .B(n15492), .Z(\SUBBYTES[8].a/w2087 ) );
  XOR \SUBBYTES[8].a/U4549  ( .A(\w1[8][49] ), .B(n15494), .Z(n15492) );
  XOR \SUBBYTES[8].a/U4548  ( .A(\SUBBYTES[8].a/w2062 ), .B(
        \SUBBYTES[8].a/w2064 ), .Z(n15493) );
  XOR \SUBBYTES[8].a/U4547  ( .A(\SUBBYTES[8].a/w2046 ), .B(
        \SUBBYTES[8].a/w2047 ), .Z(n15494) );
  XOR \SUBBYTES[8].a/U4546  ( .A(\w1[8][57] ), .B(n15495), .Z(n15993) );
  XOR \SUBBYTES[8].a/U4545  ( .A(\w1[8][59] ), .B(\w1[8][58] ), .Z(n15495) );
  XOR \SUBBYTES[8].a/U4544  ( .A(\w1[8][62] ), .B(n15993), .Z(
        \SUBBYTES[8].a/w1929 ) );
  XOR \SUBBYTES[8].a/U4543  ( .A(\w1[8][56] ), .B(\SUBBYTES[8].a/w1929 ), .Z(
        \SUBBYTES[8].a/w1816 ) );
  XOR \SUBBYTES[8].a/U4542  ( .A(\w1[8][56] ), .B(n15496), .Z(
        \SUBBYTES[8].a/w1817 ) );
  XOR \SUBBYTES[8].a/U4541  ( .A(\w1[8][62] ), .B(\w1[8][61] ), .Z(n15496) );
  XOR \SUBBYTES[8].a/U4540  ( .A(\w1[8][61] ), .B(n15993), .Z(
        \SUBBYTES[8].a/w1947 ) );
  XOR \SUBBYTES[8].a/U4539  ( .A(n15498), .B(n15497), .Z(\SUBBYTES[8].a/w1940 ) );
  XOR \SUBBYTES[8].a/U4538  ( .A(\w1[8][59] ), .B(\w1[8][57] ), .Z(n15497) );
  XOR \SUBBYTES[8].a/U4537  ( .A(\w1[8][63] ), .B(\w1[8][60] ), .Z(n15498) );
  XOR \SUBBYTES[8].a/U4536  ( .A(\w1[8][56] ), .B(\SUBBYTES[8].a/w1940 ), .Z(
        \SUBBYTES[8].a/w1819 ) );
  XOR \SUBBYTES[8].a/U4535  ( .A(n15500), .B(n15499), .Z(\SUBBYTES[8].a/w1927 ) );
  XOR \SUBBYTES[8].a/U4534  ( .A(\SUBBYTES[8].a/w1888 ), .B(n1077), .Z(n15499)
         );
  XOR \SUBBYTES[8].a/U4533  ( .A(\SUBBYTES[8].a/w1881 ), .B(
        \SUBBYTES[8].a/w1884 ), .Z(n15500) );
  XOR \SUBBYTES[8].a/U4532  ( .A(n15502), .B(n15501), .Z(\SUBBYTES[8].a/w1928 ) );
  XOR \SUBBYTES[8].a/U4531  ( .A(\SUBBYTES[8].a/w1888 ), .B(n14809), .Z(n15501) );
  XOR \SUBBYTES[8].a/U4530  ( .A(\SUBBYTES[8].a/w1881 ), .B(n14808), .Z(n15502) );
  XOR \SUBBYTES[8].a/U4529  ( .A(\SUBBYTES[8].a/w1940 ), .B(n15503), .Z(
        \SUBBYTES[8].a/w1930 ) );
  XOR \SUBBYTES[8].a/U4528  ( .A(\w1[8][62] ), .B(\w1[8][61] ), .Z(n15503) );
  XOR \SUBBYTES[8].a/U4527  ( .A(n15505), .B(n15504), .Z(\SUBBYTES[8].a/w1931 ) );
  XOR \SUBBYTES[8].a/U4526  ( .A(n14809), .B(n1077), .Z(n15504) );
  XOR \SUBBYTES[8].a/U4525  ( .A(n14808), .B(\SUBBYTES[8].a/w1884 ), .Z(n15505) );
  XOR \SUBBYTES[8].a/U4524  ( .A(\w1[8][63] ), .B(\w1[8][58] ), .Z(n15999) );
  XOR \SUBBYTES[8].a/U4523  ( .A(n15999), .B(n15506), .Z(\SUBBYTES[8].a/w1932 ) );
  XOR \SUBBYTES[8].a/U4522  ( .A(\w1[8][61] ), .B(\w1[8][60] ), .Z(n15506) );
  XOR \SUBBYTES[8].a/U4521  ( .A(\w1[8][63] ), .B(\SUBBYTES[8].a/w1817 ), .Z(
        \SUBBYTES[8].a/w1820 ) );
  XOR \SUBBYTES[8].a/U4520  ( .A(\w1[8][57] ), .B(\SUBBYTES[8].a/w1817 ), .Z(
        \SUBBYTES[8].a/w1821 ) );
  XOR \SUBBYTES[8].a/U4519  ( .A(\w1[8][60] ), .B(\SUBBYTES[8].a/w1817 ), .Z(
        \SUBBYTES[8].a/w1822 ) );
  XOR \SUBBYTES[8].a/U4518  ( .A(\SUBBYTES[8].a/w1821 ), .B(n15999), .Z(
        \SUBBYTES[8].a/w1823 ) );
  XOR \SUBBYTES[8].a/U4517  ( .A(n15999), .B(n15507), .Z(\SUBBYTES[8].a/w1908 ) );
  XOR \SUBBYTES[8].a/U4516  ( .A(\w1[8][60] ), .B(\w1[8][57] ), .Z(n15507) );
  XOR \SUBBYTES[8].a/U4515  ( .A(n15509), .B(n15508), .Z(n15996) );
  XOR \SUBBYTES[8].a/U4514  ( .A(\w1[8][60] ), .B(n15510), .Z(n15508) );
  XOR \SUBBYTES[8].a/U4513  ( .A(\SUBBYTES[8].a/w1873 ), .B(\w1[8][62] ), .Z(
        n15509) );
  XOR \SUBBYTES[8].a/U4512  ( .A(\SUBBYTES[8].a/w1847 ), .B(
        \SUBBYTES[8].a/w1854 ), .Z(n15510) );
  XOR \SUBBYTES[8].a/U4511  ( .A(n15512), .B(n15511), .Z(n15994) );
  XOR \SUBBYTES[8].a/U4510  ( .A(\w1[8][57] ), .B(n15513), .Z(n15511) );
  XOR \SUBBYTES[8].a/U4509  ( .A(\SUBBYTES[8].a/w1872 ), .B(\w1[8][61] ), .Z(
        n15512) );
  XOR \SUBBYTES[8].a/U4508  ( .A(\SUBBYTES[8].a/w1848 ), .B(
        \SUBBYTES[8].a/w1855 ), .Z(n15513) );
  XOR \SUBBYTES[8].a/U4507  ( .A(n15996), .B(n15994), .Z(\SUBBYTES[8].a/w1878 ) );
  XOR \SUBBYTES[8].a/U4506  ( .A(\w1[8][61] ), .B(n15514), .Z(n15997) );
  XOR \SUBBYTES[8].a/U4505  ( .A(\SUBBYTES[8].a/w1840 ), .B(
        \SUBBYTES[8].a/w1850 ), .Z(n15514) );
  XOR \SUBBYTES[8].a/U4504  ( .A(n15516), .B(n15515), .Z(\SUBBYTES[8].a/w1865 ) );
  XOR \SUBBYTES[8].a/U4503  ( .A(n15997), .B(n15517), .Z(n15515) );
  XOR \SUBBYTES[8].a/U4502  ( .A(\w1[8][60] ), .B(\SUBBYTES[8].a/w1929 ), .Z(
        n15516) );
  XOR \SUBBYTES[8].a/U4501  ( .A(\SUBBYTES[8].a/w1842 ), .B(
        \SUBBYTES[8].a/w1847 ), .Z(n15517) );
  XOR \SUBBYTES[8].a/U4500  ( .A(n15519), .B(n15518), .Z(n15995) );
  XOR \SUBBYTES[8].a/U4499  ( .A(\SUBBYTES[8].a/w1875 ), .B(\w1[8][63] ), .Z(
        n15518) );
  XOR \SUBBYTES[8].a/U4498  ( .A(\SUBBYTES[8].a/w1850 ), .B(
        \SUBBYTES[8].a/w1857 ), .Z(n15519) );
  XOR \SUBBYTES[8].a/U4497  ( .A(n15994), .B(n15995), .Z(\SUBBYTES[8].a/w1877 ) );
  XOR \SUBBYTES[8].a/U4496  ( .A(\w1[8][59] ), .B(n15520), .Z(n15998) );
  XOR \SUBBYTES[8].a/U4495  ( .A(\SUBBYTES[8].a/w1839 ), .B(
        \SUBBYTES[8].a/w1842 ), .Z(n15520) );
  XOR \SUBBYTES[8].a/U4494  ( .A(n15522), .B(n15521), .Z(\SUBBYTES[8].a/w1866 ) );
  XOR \SUBBYTES[8].a/U4493  ( .A(n15998), .B(n15523), .Z(n15521) );
  XOR \SUBBYTES[8].a/U4492  ( .A(\w1[8][62] ), .B(\SUBBYTES[8].a/w1908 ), .Z(
        n15522) );
  XOR \SUBBYTES[8].a/U4491  ( .A(\SUBBYTES[8].a/w1847 ), .B(
        \SUBBYTES[8].a/w1848 ), .Z(n15523) );
  XOR \SUBBYTES[8].a/U4490  ( .A(n15996), .B(n15995), .Z(\SUBBYTES[8].a/w1886 ) );
  XOR \SUBBYTES[8].a/U4489  ( .A(n15525), .B(n15524), .Z(\SUBBYTES[8].a/w1887 ) );
  XOR \SUBBYTES[8].a/U4488  ( .A(\w1[8][63] ), .B(n15997), .Z(n15524) );
  XOR \SUBBYTES[8].a/U4487  ( .A(\SUBBYTES[8].a/w1839 ), .B(
        \SUBBYTES[8].a/w1848 ), .Z(n15525) );
  XOR \SUBBYTES[8].a/U4486  ( .A(n15527), .B(n15526), .Z(\SUBBYTES[8].a/w1863 ) );
  XOR \SUBBYTES[8].a/U4485  ( .A(n15529), .B(n15528), .Z(n15526) );
  XOR \SUBBYTES[8].a/U4484  ( .A(\w1[8][63] ), .B(\SUBBYTES[8].a/w1947 ), .Z(
        n15527) );
  XOR \SUBBYTES[8].a/U4483  ( .A(\SUBBYTES[8].a/w1854 ), .B(
        \SUBBYTES[8].a/w1857 ), .Z(n15528) );
  XOR \SUBBYTES[8].a/U4482  ( .A(\SUBBYTES[8].a/w1840 ), .B(
        \SUBBYTES[8].a/w1842 ), .Z(n15529) );
  XOR \SUBBYTES[8].a/U4481  ( .A(n15531), .B(n15530), .Z(\SUBBYTES[8].a/w1864 ) );
  XOR \SUBBYTES[8].a/U4480  ( .A(n15998), .B(n15532), .Z(n15530) );
  XOR \SUBBYTES[8].a/U4479  ( .A(\w1[8][61] ), .B(n15999), .Z(n15531) );
  XOR \SUBBYTES[8].a/U4478  ( .A(\SUBBYTES[8].a/w1854 ), .B(
        \SUBBYTES[8].a/w1855 ), .Z(n15532) );
  XOR \SUBBYTES[8].a/U4477  ( .A(n15534), .B(n15533), .Z(\SUBBYTES[8].a/w1880 ) );
  XOR \SUBBYTES[8].a/U4476  ( .A(\w1[8][57] ), .B(n15535), .Z(n15533) );
  XOR \SUBBYTES[8].a/U4475  ( .A(\SUBBYTES[8].a/w1855 ), .B(
        \SUBBYTES[8].a/w1857 ), .Z(n15534) );
  XOR \SUBBYTES[8].a/U4474  ( .A(\SUBBYTES[8].a/w1839 ), .B(
        \SUBBYTES[8].a/w1840 ), .Z(n15535) );
  XOR \SUBBYTES[8].a/U4473  ( .A(\w1[8][65] ), .B(n15536), .Z(n16000) );
  XOR \SUBBYTES[8].a/U4472  ( .A(\w1[8][67] ), .B(\w1[8][66] ), .Z(n15536) );
  XOR \SUBBYTES[8].a/U4471  ( .A(\w1[8][70] ), .B(n16000), .Z(
        \SUBBYTES[8].a/w1722 ) );
  XOR \SUBBYTES[8].a/U4470  ( .A(\w1[8][64] ), .B(\SUBBYTES[8].a/w1722 ), .Z(
        \SUBBYTES[8].a/w1609 ) );
  XOR \SUBBYTES[8].a/U4469  ( .A(\w1[8][64] ), .B(n15537), .Z(
        \SUBBYTES[8].a/w1610 ) );
  XOR \SUBBYTES[8].a/U4468  ( .A(\w1[8][70] ), .B(\w1[8][69] ), .Z(n15537) );
  XOR \SUBBYTES[8].a/U4467  ( .A(\w1[8][69] ), .B(n16000), .Z(
        \SUBBYTES[8].a/w1740 ) );
  XOR \SUBBYTES[8].a/U4466  ( .A(n15539), .B(n15538), .Z(\SUBBYTES[8].a/w1733 ) );
  XOR \SUBBYTES[8].a/U4465  ( .A(\w1[8][67] ), .B(\w1[8][65] ), .Z(n15538) );
  XOR \SUBBYTES[8].a/U4464  ( .A(\w1[8][71] ), .B(\w1[8][68] ), .Z(n15539) );
  XOR \SUBBYTES[8].a/U4463  ( .A(\w1[8][64] ), .B(\SUBBYTES[8].a/w1733 ), .Z(
        \SUBBYTES[8].a/w1612 ) );
  XOR \SUBBYTES[8].a/U4462  ( .A(n15541), .B(n15540), .Z(\SUBBYTES[8].a/w1720 ) );
  XOR \SUBBYTES[8].a/U4461  ( .A(\SUBBYTES[8].a/w1681 ), .B(n1076), .Z(n15540)
         );
  XOR \SUBBYTES[8].a/U4460  ( .A(\SUBBYTES[8].a/w1674 ), .B(
        \SUBBYTES[8].a/w1677 ), .Z(n15541) );
  XOR \SUBBYTES[8].a/U4459  ( .A(n15543), .B(n15542), .Z(\SUBBYTES[8].a/w1721 ) );
  XOR \SUBBYTES[8].a/U4458  ( .A(\SUBBYTES[8].a/w1681 ), .B(n14807), .Z(n15542) );
  XOR \SUBBYTES[8].a/U4457  ( .A(\SUBBYTES[8].a/w1674 ), .B(n14806), .Z(n15543) );
  XOR \SUBBYTES[8].a/U4456  ( .A(\SUBBYTES[8].a/w1733 ), .B(n15544), .Z(
        \SUBBYTES[8].a/w1723 ) );
  XOR \SUBBYTES[8].a/U4455  ( .A(\w1[8][70] ), .B(\w1[8][69] ), .Z(n15544) );
  XOR \SUBBYTES[8].a/U4454  ( .A(n15546), .B(n15545), .Z(\SUBBYTES[8].a/w1724 ) );
  XOR \SUBBYTES[8].a/U4453  ( .A(n14807), .B(n1076), .Z(n15545) );
  XOR \SUBBYTES[8].a/U4452  ( .A(n14806), .B(\SUBBYTES[8].a/w1677 ), .Z(n15546) );
  XOR \SUBBYTES[8].a/U4451  ( .A(\w1[8][71] ), .B(\w1[8][66] ), .Z(n16006) );
  XOR \SUBBYTES[8].a/U4450  ( .A(n16006), .B(n15547), .Z(\SUBBYTES[8].a/w1725 ) );
  XOR \SUBBYTES[8].a/U4449  ( .A(\w1[8][69] ), .B(\w1[8][68] ), .Z(n15547) );
  XOR \SUBBYTES[8].a/U4448  ( .A(\w1[8][71] ), .B(\SUBBYTES[8].a/w1610 ), .Z(
        \SUBBYTES[8].a/w1613 ) );
  XOR \SUBBYTES[8].a/U4447  ( .A(\w1[8][65] ), .B(\SUBBYTES[8].a/w1610 ), .Z(
        \SUBBYTES[8].a/w1614 ) );
  XOR \SUBBYTES[8].a/U4446  ( .A(\w1[8][68] ), .B(\SUBBYTES[8].a/w1610 ), .Z(
        \SUBBYTES[8].a/w1615 ) );
  XOR \SUBBYTES[8].a/U4445  ( .A(\SUBBYTES[8].a/w1614 ), .B(n16006), .Z(
        \SUBBYTES[8].a/w1616 ) );
  XOR \SUBBYTES[8].a/U4444  ( .A(n16006), .B(n15548), .Z(\SUBBYTES[8].a/w1701 ) );
  XOR \SUBBYTES[8].a/U4443  ( .A(\w1[8][68] ), .B(\w1[8][65] ), .Z(n15548) );
  XOR \SUBBYTES[8].a/U4442  ( .A(n15550), .B(n15549), .Z(n16003) );
  XOR \SUBBYTES[8].a/U4441  ( .A(\w1[8][68] ), .B(n15551), .Z(n15549) );
  XOR \SUBBYTES[8].a/U4440  ( .A(\SUBBYTES[8].a/w1666 ), .B(\w1[8][70] ), .Z(
        n15550) );
  XOR \SUBBYTES[8].a/U4439  ( .A(\SUBBYTES[8].a/w1640 ), .B(
        \SUBBYTES[8].a/w1647 ), .Z(n15551) );
  XOR \SUBBYTES[8].a/U4438  ( .A(n15553), .B(n15552), .Z(n16001) );
  XOR \SUBBYTES[8].a/U4437  ( .A(\w1[8][65] ), .B(n15554), .Z(n15552) );
  XOR \SUBBYTES[8].a/U4436  ( .A(\SUBBYTES[8].a/w1665 ), .B(\w1[8][69] ), .Z(
        n15553) );
  XOR \SUBBYTES[8].a/U4435  ( .A(\SUBBYTES[8].a/w1641 ), .B(
        \SUBBYTES[8].a/w1648 ), .Z(n15554) );
  XOR \SUBBYTES[8].a/U4434  ( .A(n16003), .B(n16001), .Z(\SUBBYTES[8].a/w1671 ) );
  XOR \SUBBYTES[8].a/U4433  ( .A(\w1[8][69] ), .B(n15555), .Z(n16004) );
  XOR \SUBBYTES[8].a/U4432  ( .A(\SUBBYTES[8].a/w1633 ), .B(
        \SUBBYTES[8].a/w1643 ), .Z(n15555) );
  XOR \SUBBYTES[8].a/U4431  ( .A(n15557), .B(n15556), .Z(\SUBBYTES[8].a/w1658 ) );
  XOR \SUBBYTES[8].a/U4430  ( .A(n16004), .B(n15558), .Z(n15556) );
  XOR \SUBBYTES[8].a/U4429  ( .A(\w1[8][68] ), .B(\SUBBYTES[8].a/w1722 ), .Z(
        n15557) );
  XOR \SUBBYTES[8].a/U4428  ( .A(\SUBBYTES[8].a/w1635 ), .B(
        \SUBBYTES[8].a/w1640 ), .Z(n15558) );
  XOR \SUBBYTES[8].a/U4427  ( .A(n15560), .B(n15559), .Z(n16002) );
  XOR \SUBBYTES[8].a/U4426  ( .A(\SUBBYTES[8].a/w1668 ), .B(\w1[8][71] ), .Z(
        n15559) );
  XOR \SUBBYTES[8].a/U4425  ( .A(\SUBBYTES[8].a/w1643 ), .B(
        \SUBBYTES[8].a/w1650 ), .Z(n15560) );
  XOR \SUBBYTES[8].a/U4424  ( .A(n16001), .B(n16002), .Z(\SUBBYTES[8].a/w1670 ) );
  XOR \SUBBYTES[8].a/U4423  ( .A(\w1[8][67] ), .B(n15561), .Z(n16005) );
  XOR \SUBBYTES[8].a/U4422  ( .A(\SUBBYTES[8].a/w1632 ), .B(
        \SUBBYTES[8].a/w1635 ), .Z(n15561) );
  XOR \SUBBYTES[8].a/U4421  ( .A(n15563), .B(n15562), .Z(\SUBBYTES[8].a/w1659 ) );
  XOR \SUBBYTES[8].a/U4420  ( .A(n16005), .B(n15564), .Z(n15562) );
  XOR \SUBBYTES[8].a/U4419  ( .A(\w1[8][70] ), .B(\SUBBYTES[8].a/w1701 ), .Z(
        n15563) );
  XOR \SUBBYTES[8].a/U4418  ( .A(\SUBBYTES[8].a/w1640 ), .B(
        \SUBBYTES[8].a/w1641 ), .Z(n15564) );
  XOR \SUBBYTES[8].a/U4417  ( .A(n16003), .B(n16002), .Z(\SUBBYTES[8].a/w1679 ) );
  XOR \SUBBYTES[8].a/U4416  ( .A(n15566), .B(n15565), .Z(\SUBBYTES[8].a/w1680 ) );
  XOR \SUBBYTES[8].a/U4415  ( .A(\w1[8][71] ), .B(n16004), .Z(n15565) );
  XOR \SUBBYTES[8].a/U4414  ( .A(\SUBBYTES[8].a/w1632 ), .B(
        \SUBBYTES[8].a/w1641 ), .Z(n15566) );
  XOR \SUBBYTES[8].a/U4413  ( .A(n15568), .B(n15567), .Z(\SUBBYTES[8].a/w1656 ) );
  XOR \SUBBYTES[8].a/U4412  ( .A(n15570), .B(n15569), .Z(n15567) );
  XOR \SUBBYTES[8].a/U4411  ( .A(\w1[8][71] ), .B(\SUBBYTES[8].a/w1740 ), .Z(
        n15568) );
  XOR \SUBBYTES[8].a/U4410  ( .A(\SUBBYTES[8].a/w1647 ), .B(
        \SUBBYTES[8].a/w1650 ), .Z(n15569) );
  XOR \SUBBYTES[8].a/U4409  ( .A(\SUBBYTES[8].a/w1633 ), .B(
        \SUBBYTES[8].a/w1635 ), .Z(n15570) );
  XOR \SUBBYTES[8].a/U4408  ( .A(n15572), .B(n15571), .Z(\SUBBYTES[8].a/w1657 ) );
  XOR \SUBBYTES[8].a/U4407  ( .A(n16005), .B(n15573), .Z(n15571) );
  XOR \SUBBYTES[8].a/U4406  ( .A(\w1[8][69] ), .B(n16006), .Z(n15572) );
  XOR \SUBBYTES[8].a/U4405  ( .A(\SUBBYTES[8].a/w1647 ), .B(
        \SUBBYTES[8].a/w1648 ), .Z(n15573) );
  XOR \SUBBYTES[8].a/U4404  ( .A(n15575), .B(n15574), .Z(\SUBBYTES[8].a/w1673 ) );
  XOR \SUBBYTES[8].a/U4403  ( .A(\w1[8][65] ), .B(n15576), .Z(n15574) );
  XOR \SUBBYTES[8].a/U4402  ( .A(\SUBBYTES[8].a/w1648 ), .B(
        \SUBBYTES[8].a/w1650 ), .Z(n15575) );
  XOR \SUBBYTES[8].a/U4401  ( .A(\SUBBYTES[8].a/w1632 ), .B(
        \SUBBYTES[8].a/w1633 ), .Z(n15576) );
  XOR \SUBBYTES[8].a/U4400  ( .A(\w1[8][73] ), .B(n15577), .Z(n16007) );
  XOR \SUBBYTES[8].a/U4399  ( .A(\w1[8][75] ), .B(\w1[8][74] ), .Z(n15577) );
  XOR \SUBBYTES[8].a/U4398  ( .A(\w1[8][78] ), .B(n16007), .Z(
        \SUBBYTES[8].a/w1515 ) );
  XOR \SUBBYTES[8].a/U4397  ( .A(\w1[8][72] ), .B(\SUBBYTES[8].a/w1515 ), .Z(
        \SUBBYTES[8].a/w1402 ) );
  XOR \SUBBYTES[8].a/U4396  ( .A(\w1[8][72] ), .B(n15578), .Z(
        \SUBBYTES[8].a/w1403 ) );
  XOR \SUBBYTES[8].a/U4395  ( .A(\w1[8][78] ), .B(\w1[8][77] ), .Z(n15578) );
  XOR \SUBBYTES[8].a/U4394  ( .A(\w1[8][77] ), .B(n16007), .Z(
        \SUBBYTES[8].a/w1533 ) );
  XOR \SUBBYTES[8].a/U4393  ( .A(n15580), .B(n15579), .Z(\SUBBYTES[8].a/w1526 ) );
  XOR \SUBBYTES[8].a/U4392  ( .A(\w1[8][75] ), .B(\w1[8][73] ), .Z(n15579) );
  XOR \SUBBYTES[8].a/U4391  ( .A(\w1[8][79] ), .B(\w1[8][76] ), .Z(n15580) );
  XOR \SUBBYTES[8].a/U4390  ( .A(\w1[8][72] ), .B(\SUBBYTES[8].a/w1526 ), .Z(
        \SUBBYTES[8].a/w1405 ) );
  XOR \SUBBYTES[8].a/U4389  ( .A(n15582), .B(n15581), .Z(\SUBBYTES[8].a/w1513 ) );
  XOR \SUBBYTES[8].a/U4388  ( .A(\SUBBYTES[8].a/w1474 ), .B(n1075), .Z(n15581)
         );
  XOR \SUBBYTES[8].a/U4387  ( .A(\SUBBYTES[8].a/w1467 ), .B(
        \SUBBYTES[8].a/w1470 ), .Z(n15582) );
  XOR \SUBBYTES[8].a/U4386  ( .A(n15584), .B(n15583), .Z(\SUBBYTES[8].a/w1514 ) );
  XOR \SUBBYTES[8].a/U4385  ( .A(\SUBBYTES[8].a/w1474 ), .B(n14805), .Z(n15583) );
  XOR \SUBBYTES[8].a/U4384  ( .A(\SUBBYTES[8].a/w1467 ), .B(n14804), .Z(n15584) );
  XOR \SUBBYTES[8].a/U4383  ( .A(\SUBBYTES[8].a/w1526 ), .B(n15585), .Z(
        \SUBBYTES[8].a/w1516 ) );
  XOR \SUBBYTES[8].a/U4382  ( .A(\w1[8][78] ), .B(\w1[8][77] ), .Z(n15585) );
  XOR \SUBBYTES[8].a/U4381  ( .A(n15587), .B(n15586), .Z(\SUBBYTES[8].a/w1517 ) );
  XOR \SUBBYTES[8].a/U4380  ( .A(n14805), .B(n1075), .Z(n15586) );
  XOR \SUBBYTES[8].a/U4379  ( .A(n14804), .B(\SUBBYTES[8].a/w1470 ), .Z(n15587) );
  XOR \SUBBYTES[8].a/U4378  ( .A(\w1[8][79] ), .B(\w1[8][74] ), .Z(n16013) );
  XOR \SUBBYTES[8].a/U4377  ( .A(n16013), .B(n15588), .Z(\SUBBYTES[8].a/w1518 ) );
  XOR \SUBBYTES[8].a/U4376  ( .A(\w1[8][77] ), .B(\w1[8][76] ), .Z(n15588) );
  XOR \SUBBYTES[8].a/U4375  ( .A(\w1[8][79] ), .B(\SUBBYTES[8].a/w1403 ), .Z(
        \SUBBYTES[8].a/w1406 ) );
  XOR \SUBBYTES[8].a/U4374  ( .A(\w1[8][73] ), .B(\SUBBYTES[8].a/w1403 ), .Z(
        \SUBBYTES[8].a/w1407 ) );
  XOR \SUBBYTES[8].a/U4373  ( .A(\w1[8][76] ), .B(\SUBBYTES[8].a/w1403 ), .Z(
        \SUBBYTES[8].a/w1408 ) );
  XOR \SUBBYTES[8].a/U4372  ( .A(\SUBBYTES[8].a/w1407 ), .B(n16013), .Z(
        \SUBBYTES[8].a/w1409 ) );
  XOR \SUBBYTES[8].a/U4371  ( .A(n16013), .B(n15589), .Z(\SUBBYTES[8].a/w1494 ) );
  XOR \SUBBYTES[8].a/U4370  ( .A(\w1[8][76] ), .B(\w1[8][73] ), .Z(n15589) );
  XOR \SUBBYTES[8].a/U4369  ( .A(n15591), .B(n15590), .Z(n16010) );
  XOR \SUBBYTES[8].a/U4368  ( .A(\w1[8][76] ), .B(n15592), .Z(n15590) );
  XOR \SUBBYTES[8].a/U4367  ( .A(\SUBBYTES[8].a/w1459 ), .B(\w1[8][78] ), .Z(
        n15591) );
  XOR \SUBBYTES[8].a/U4366  ( .A(\SUBBYTES[8].a/w1433 ), .B(
        \SUBBYTES[8].a/w1440 ), .Z(n15592) );
  XOR \SUBBYTES[8].a/U4365  ( .A(n15594), .B(n15593), .Z(n16008) );
  XOR \SUBBYTES[8].a/U4364  ( .A(\w1[8][73] ), .B(n15595), .Z(n15593) );
  XOR \SUBBYTES[8].a/U4363  ( .A(\SUBBYTES[8].a/w1458 ), .B(\w1[8][77] ), .Z(
        n15594) );
  XOR \SUBBYTES[8].a/U4362  ( .A(\SUBBYTES[8].a/w1434 ), .B(
        \SUBBYTES[8].a/w1441 ), .Z(n15595) );
  XOR \SUBBYTES[8].a/U4361  ( .A(n16010), .B(n16008), .Z(\SUBBYTES[8].a/w1464 ) );
  XOR \SUBBYTES[8].a/U4360  ( .A(\w1[8][77] ), .B(n15596), .Z(n16011) );
  XOR \SUBBYTES[8].a/U4359  ( .A(\SUBBYTES[8].a/w1426 ), .B(
        \SUBBYTES[8].a/w1436 ), .Z(n15596) );
  XOR \SUBBYTES[8].a/U4358  ( .A(n15598), .B(n15597), .Z(\SUBBYTES[8].a/w1451 ) );
  XOR \SUBBYTES[8].a/U4357  ( .A(n16011), .B(n15599), .Z(n15597) );
  XOR \SUBBYTES[8].a/U4356  ( .A(\w1[8][76] ), .B(\SUBBYTES[8].a/w1515 ), .Z(
        n15598) );
  XOR \SUBBYTES[8].a/U4355  ( .A(\SUBBYTES[8].a/w1428 ), .B(
        \SUBBYTES[8].a/w1433 ), .Z(n15599) );
  XOR \SUBBYTES[8].a/U4354  ( .A(n15601), .B(n15600), .Z(n16009) );
  XOR \SUBBYTES[8].a/U4353  ( .A(\SUBBYTES[8].a/w1461 ), .B(\w1[8][79] ), .Z(
        n15600) );
  XOR \SUBBYTES[8].a/U4352  ( .A(\SUBBYTES[8].a/w1436 ), .B(
        \SUBBYTES[8].a/w1443 ), .Z(n15601) );
  XOR \SUBBYTES[8].a/U4351  ( .A(n16008), .B(n16009), .Z(\SUBBYTES[8].a/w1463 ) );
  XOR \SUBBYTES[8].a/U4350  ( .A(\w1[8][75] ), .B(n15602), .Z(n16012) );
  XOR \SUBBYTES[8].a/U4349  ( .A(\SUBBYTES[8].a/w1425 ), .B(
        \SUBBYTES[8].a/w1428 ), .Z(n15602) );
  XOR \SUBBYTES[8].a/U4348  ( .A(n15604), .B(n15603), .Z(\SUBBYTES[8].a/w1452 ) );
  XOR \SUBBYTES[8].a/U4347  ( .A(n16012), .B(n15605), .Z(n15603) );
  XOR \SUBBYTES[8].a/U4346  ( .A(\w1[8][78] ), .B(\SUBBYTES[8].a/w1494 ), .Z(
        n15604) );
  XOR \SUBBYTES[8].a/U4345  ( .A(\SUBBYTES[8].a/w1433 ), .B(
        \SUBBYTES[8].a/w1434 ), .Z(n15605) );
  XOR \SUBBYTES[8].a/U4344  ( .A(n16010), .B(n16009), .Z(\SUBBYTES[8].a/w1472 ) );
  XOR \SUBBYTES[8].a/U4343  ( .A(n15607), .B(n15606), .Z(\SUBBYTES[8].a/w1473 ) );
  XOR \SUBBYTES[8].a/U4342  ( .A(\w1[8][79] ), .B(n16011), .Z(n15606) );
  XOR \SUBBYTES[8].a/U4341  ( .A(\SUBBYTES[8].a/w1425 ), .B(
        \SUBBYTES[8].a/w1434 ), .Z(n15607) );
  XOR \SUBBYTES[8].a/U4340  ( .A(n15609), .B(n15608), .Z(\SUBBYTES[8].a/w1449 ) );
  XOR \SUBBYTES[8].a/U4339  ( .A(n15611), .B(n15610), .Z(n15608) );
  XOR \SUBBYTES[8].a/U4338  ( .A(\w1[8][79] ), .B(\SUBBYTES[8].a/w1533 ), .Z(
        n15609) );
  XOR \SUBBYTES[8].a/U4337  ( .A(\SUBBYTES[8].a/w1440 ), .B(
        \SUBBYTES[8].a/w1443 ), .Z(n15610) );
  XOR \SUBBYTES[8].a/U4336  ( .A(\SUBBYTES[8].a/w1426 ), .B(
        \SUBBYTES[8].a/w1428 ), .Z(n15611) );
  XOR \SUBBYTES[8].a/U4335  ( .A(n15613), .B(n15612), .Z(\SUBBYTES[8].a/w1450 ) );
  XOR \SUBBYTES[8].a/U4334  ( .A(n16012), .B(n15614), .Z(n15612) );
  XOR \SUBBYTES[8].a/U4333  ( .A(\w1[8][77] ), .B(n16013), .Z(n15613) );
  XOR \SUBBYTES[8].a/U4332  ( .A(\SUBBYTES[8].a/w1440 ), .B(
        \SUBBYTES[8].a/w1441 ), .Z(n15614) );
  XOR \SUBBYTES[8].a/U4331  ( .A(n15616), .B(n15615), .Z(\SUBBYTES[8].a/w1466 ) );
  XOR \SUBBYTES[8].a/U4330  ( .A(\w1[8][73] ), .B(n15617), .Z(n15615) );
  XOR \SUBBYTES[8].a/U4329  ( .A(\SUBBYTES[8].a/w1441 ), .B(
        \SUBBYTES[8].a/w1443 ), .Z(n15616) );
  XOR \SUBBYTES[8].a/U4328  ( .A(\SUBBYTES[8].a/w1425 ), .B(
        \SUBBYTES[8].a/w1426 ), .Z(n15617) );
  XOR \SUBBYTES[8].a/U4327  ( .A(\w1[8][81] ), .B(n15618), .Z(n16014) );
  XOR \SUBBYTES[8].a/U4326  ( .A(\w1[8][83] ), .B(\w1[8][82] ), .Z(n15618) );
  XOR \SUBBYTES[8].a/U4325  ( .A(\w1[8][86] ), .B(n16014), .Z(
        \SUBBYTES[8].a/w1308 ) );
  XOR \SUBBYTES[8].a/U4324  ( .A(\w1[8][80] ), .B(\SUBBYTES[8].a/w1308 ), .Z(
        \SUBBYTES[8].a/w1195 ) );
  XOR \SUBBYTES[8].a/U4323  ( .A(\w1[8][80] ), .B(n15619), .Z(
        \SUBBYTES[8].a/w1196 ) );
  XOR \SUBBYTES[8].a/U4322  ( .A(\w1[8][86] ), .B(\w1[8][85] ), .Z(n15619) );
  XOR \SUBBYTES[8].a/U4321  ( .A(\w1[8][85] ), .B(n16014), .Z(
        \SUBBYTES[8].a/w1326 ) );
  XOR \SUBBYTES[8].a/U4320  ( .A(n15621), .B(n15620), .Z(\SUBBYTES[8].a/w1319 ) );
  XOR \SUBBYTES[8].a/U4319  ( .A(\w1[8][83] ), .B(\w1[8][81] ), .Z(n15620) );
  XOR \SUBBYTES[8].a/U4318  ( .A(\w1[8][87] ), .B(\w1[8][84] ), .Z(n15621) );
  XOR \SUBBYTES[8].a/U4317  ( .A(\w1[8][80] ), .B(\SUBBYTES[8].a/w1319 ), .Z(
        \SUBBYTES[8].a/w1198 ) );
  XOR \SUBBYTES[8].a/U4316  ( .A(n15623), .B(n15622), .Z(\SUBBYTES[8].a/w1306 ) );
  XOR \SUBBYTES[8].a/U4315  ( .A(\SUBBYTES[8].a/w1267 ), .B(n1074), .Z(n15622)
         );
  XOR \SUBBYTES[8].a/U4314  ( .A(\SUBBYTES[8].a/w1260 ), .B(
        \SUBBYTES[8].a/w1263 ), .Z(n15623) );
  XOR \SUBBYTES[8].a/U4313  ( .A(n15625), .B(n15624), .Z(\SUBBYTES[8].a/w1307 ) );
  XOR \SUBBYTES[8].a/U4312  ( .A(\SUBBYTES[8].a/w1267 ), .B(n14803), .Z(n15624) );
  XOR \SUBBYTES[8].a/U4311  ( .A(\SUBBYTES[8].a/w1260 ), .B(n14802), .Z(n15625) );
  XOR \SUBBYTES[8].a/U4310  ( .A(\SUBBYTES[8].a/w1319 ), .B(n15626), .Z(
        \SUBBYTES[8].a/w1309 ) );
  XOR \SUBBYTES[8].a/U4309  ( .A(\w1[8][86] ), .B(\w1[8][85] ), .Z(n15626) );
  XOR \SUBBYTES[8].a/U4308  ( .A(n15628), .B(n15627), .Z(\SUBBYTES[8].a/w1310 ) );
  XOR \SUBBYTES[8].a/U4307  ( .A(n14803), .B(n1074), .Z(n15627) );
  XOR \SUBBYTES[8].a/U4306  ( .A(n14802), .B(\SUBBYTES[8].a/w1263 ), .Z(n15628) );
  XOR \SUBBYTES[8].a/U4305  ( .A(\w1[8][87] ), .B(\w1[8][82] ), .Z(n16020) );
  XOR \SUBBYTES[8].a/U4304  ( .A(n16020), .B(n15629), .Z(\SUBBYTES[8].a/w1311 ) );
  XOR \SUBBYTES[8].a/U4303  ( .A(\w1[8][85] ), .B(\w1[8][84] ), .Z(n15629) );
  XOR \SUBBYTES[8].a/U4302  ( .A(\w1[8][87] ), .B(\SUBBYTES[8].a/w1196 ), .Z(
        \SUBBYTES[8].a/w1199 ) );
  XOR \SUBBYTES[8].a/U4301  ( .A(\w1[8][81] ), .B(\SUBBYTES[8].a/w1196 ), .Z(
        \SUBBYTES[8].a/w1200 ) );
  XOR \SUBBYTES[8].a/U4300  ( .A(\w1[8][84] ), .B(\SUBBYTES[8].a/w1196 ), .Z(
        \SUBBYTES[8].a/w1201 ) );
  XOR \SUBBYTES[8].a/U4299  ( .A(\SUBBYTES[8].a/w1200 ), .B(n16020), .Z(
        \SUBBYTES[8].a/w1202 ) );
  XOR \SUBBYTES[8].a/U4298  ( .A(n16020), .B(n15630), .Z(\SUBBYTES[8].a/w1287 ) );
  XOR \SUBBYTES[8].a/U4297  ( .A(\w1[8][84] ), .B(\w1[8][81] ), .Z(n15630) );
  XOR \SUBBYTES[8].a/U4296  ( .A(n15632), .B(n15631), .Z(n16017) );
  XOR \SUBBYTES[8].a/U4295  ( .A(\w1[8][84] ), .B(n15633), .Z(n15631) );
  XOR \SUBBYTES[8].a/U4294  ( .A(\SUBBYTES[8].a/w1252 ), .B(\w1[8][86] ), .Z(
        n15632) );
  XOR \SUBBYTES[8].a/U4293  ( .A(\SUBBYTES[8].a/w1226 ), .B(
        \SUBBYTES[8].a/w1233 ), .Z(n15633) );
  XOR \SUBBYTES[8].a/U4292  ( .A(n15635), .B(n15634), .Z(n16015) );
  XOR \SUBBYTES[8].a/U4291  ( .A(\w1[8][81] ), .B(n15636), .Z(n15634) );
  XOR \SUBBYTES[8].a/U4290  ( .A(\SUBBYTES[8].a/w1251 ), .B(\w1[8][85] ), .Z(
        n15635) );
  XOR \SUBBYTES[8].a/U4289  ( .A(\SUBBYTES[8].a/w1227 ), .B(
        \SUBBYTES[8].a/w1234 ), .Z(n15636) );
  XOR \SUBBYTES[8].a/U4288  ( .A(n16017), .B(n16015), .Z(\SUBBYTES[8].a/w1257 ) );
  XOR \SUBBYTES[8].a/U4287  ( .A(\w1[8][85] ), .B(n15637), .Z(n16018) );
  XOR \SUBBYTES[8].a/U4286  ( .A(\SUBBYTES[8].a/w1219 ), .B(
        \SUBBYTES[8].a/w1229 ), .Z(n15637) );
  XOR \SUBBYTES[8].a/U4285  ( .A(n15639), .B(n15638), .Z(\SUBBYTES[8].a/w1244 ) );
  XOR \SUBBYTES[8].a/U4284  ( .A(n16018), .B(n15640), .Z(n15638) );
  XOR \SUBBYTES[8].a/U4283  ( .A(\w1[8][84] ), .B(\SUBBYTES[8].a/w1308 ), .Z(
        n15639) );
  XOR \SUBBYTES[8].a/U4282  ( .A(\SUBBYTES[8].a/w1221 ), .B(
        \SUBBYTES[8].a/w1226 ), .Z(n15640) );
  XOR \SUBBYTES[8].a/U4281  ( .A(n15642), .B(n15641), .Z(n16016) );
  XOR \SUBBYTES[8].a/U4280  ( .A(\SUBBYTES[8].a/w1254 ), .B(\w1[8][87] ), .Z(
        n15641) );
  XOR \SUBBYTES[8].a/U4279  ( .A(\SUBBYTES[8].a/w1229 ), .B(
        \SUBBYTES[8].a/w1236 ), .Z(n15642) );
  XOR \SUBBYTES[8].a/U4278  ( .A(n16015), .B(n16016), .Z(\SUBBYTES[8].a/w1256 ) );
  XOR \SUBBYTES[8].a/U4277  ( .A(\w1[8][83] ), .B(n15643), .Z(n16019) );
  XOR \SUBBYTES[8].a/U4276  ( .A(\SUBBYTES[8].a/w1218 ), .B(
        \SUBBYTES[8].a/w1221 ), .Z(n15643) );
  XOR \SUBBYTES[8].a/U4275  ( .A(n15645), .B(n15644), .Z(\SUBBYTES[8].a/w1245 ) );
  XOR \SUBBYTES[8].a/U4274  ( .A(n16019), .B(n15646), .Z(n15644) );
  XOR \SUBBYTES[8].a/U4273  ( .A(\w1[8][86] ), .B(\SUBBYTES[8].a/w1287 ), .Z(
        n15645) );
  XOR \SUBBYTES[8].a/U4272  ( .A(\SUBBYTES[8].a/w1226 ), .B(
        \SUBBYTES[8].a/w1227 ), .Z(n15646) );
  XOR \SUBBYTES[8].a/U4271  ( .A(n16017), .B(n16016), .Z(\SUBBYTES[8].a/w1265 ) );
  XOR \SUBBYTES[8].a/U4270  ( .A(n15648), .B(n15647), .Z(\SUBBYTES[8].a/w1266 ) );
  XOR \SUBBYTES[8].a/U4269  ( .A(\w1[8][87] ), .B(n16018), .Z(n15647) );
  XOR \SUBBYTES[8].a/U4268  ( .A(\SUBBYTES[8].a/w1218 ), .B(
        \SUBBYTES[8].a/w1227 ), .Z(n15648) );
  XOR \SUBBYTES[8].a/U4267  ( .A(n15650), .B(n15649), .Z(\SUBBYTES[8].a/w1242 ) );
  XOR \SUBBYTES[8].a/U4266  ( .A(n15652), .B(n15651), .Z(n15649) );
  XOR \SUBBYTES[8].a/U4265  ( .A(\w1[8][87] ), .B(\SUBBYTES[8].a/w1326 ), .Z(
        n15650) );
  XOR \SUBBYTES[8].a/U4264  ( .A(\SUBBYTES[8].a/w1233 ), .B(
        \SUBBYTES[8].a/w1236 ), .Z(n15651) );
  XOR \SUBBYTES[8].a/U4263  ( .A(\SUBBYTES[8].a/w1219 ), .B(
        \SUBBYTES[8].a/w1221 ), .Z(n15652) );
  XOR \SUBBYTES[8].a/U4262  ( .A(n15654), .B(n15653), .Z(\SUBBYTES[8].a/w1243 ) );
  XOR \SUBBYTES[8].a/U4261  ( .A(n16019), .B(n15655), .Z(n15653) );
  XOR \SUBBYTES[8].a/U4260  ( .A(\w1[8][85] ), .B(n16020), .Z(n15654) );
  XOR \SUBBYTES[8].a/U4259  ( .A(\SUBBYTES[8].a/w1233 ), .B(
        \SUBBYTES[8].a/w1234 ), .Z(n15655) );
  XOR \SUBBYTES[8].a/U4258  ( .A(n15657), .B(n15656), .Z(\SUBBYTES[8].a/w1259 ) );
  XOR \SUBBYTES[8].a/U4257  ( .A(\w1[8][81] ), .B(n15658), .Z(n15656) );
  XOR \SUBBYTES[8].a/U4256  ( .A(\SUBBYTES[8].a/w1234 ), .B(
        \SUBBYTES[8].a/w1236 ), .Z(n15657) );
  XOR \SUBBYTES[8].a/U4255  ( .A(\SUBBYTES[8].a/w1218 ), .B(
        \SUBBYTES[8].a/w1219 ), .Z(n15658) );
  XOR \SUBBYTES[8].a/U4254  ( .A(\w1[8][89] ), .B(n15659), .Z(n16021) );
  XOR \SUBBYTES[8].a/U4253  ( .A(\w1[8][91] ), .B(\w1[8][90] ), .Z(n15659) );
  XOR \SUBBYTES[8].a/U4252  ( .A(\w1[8][94] ), .B(n16021), .Z(
        \SUBBYTES[8].a/w1101 ) );
  XOR \SUBBYTES[8].a/U4251  ( .A(\w1[8][88] ), .B(\SUBBYTES[8].a/w1101 ), .Z(
        \SUBBYTES[8].a/w988 ) );
  XOR \SUBBYTES[8].a/U4250  ( .A(\w1[8][88] ), .B(n15660), .Z(
        \SUBBYTES[8].a/w989 ) );
  XOR \SUBBYTES[8].a/U4249  ( .A(\w1[8][94] ), .B(\w1[8][93] ), .Z(n15660) );
  XOR \SUBBYTES[8].a/U4248  ( .A(\w1[8][93] ), .B(n16021), .Z(
        \SUBBYTES[8].a/w1119 ) );
  XOR \SUBBYTES[8].a/U4247  ( .A(n15662), .B(n15661), .Z(\SUBBYTES[8].a/w1112 ) );
  XOR \SUBBYTES[8].a/U4246  ( .A(\w1[8][91] ), .B(\w1[8][89] ), .Z(n15661) );
  XOR \SUBBYTES[8].a/U4245  ( .A(\w1[8][95] ), .B(\w1[8][92] ), .Z(n15662) );
  XOR \SUBBYTES[8].a/U4244  ( .A(\w1[8][88] ), .B(\SUBBYTES[8].a/w1112 ), .Z(
        \SUBBYTES[8].a/w991 ) );
  XOR \SUBBYTES[8].a/U4243  ( .A(n15664), .B(n15663), .Z(\SUBBYTES[8].a/w1099 ) );
  XOR \SUBBYTES[8].a/U4242  ( .A(\SUBBYTES[8].a/w1060 ), .B(n1073), .Z(n15663)
         );
  XOR \SUBBYTES[8].a/U4241  ( .A(\SUBBYTES[8].a/w1053 ), .B(
        \SUBBYTES[8].a/w1056 ), .Z(n15664) );
  XOR \SUBBYTES[8].a/U4240  ( .A(n15666), .B(n15665), .Z(\SUBBYTES[8].a/w1100 ) );
  XOR \SUBBYTES[8].a/U4239  ( .A(\SUBBYTES[8].a/w1060 ), .B(n14801), .Z(n15665) );
  XOR \SUBBYTES[8].a/U4238  ( .A(\SUBBYTES[8].a/w1053 ), .B(n14800), .Z(n15666) );
  XOR \SUBBYTES[8].a/U4237  ( .A(\SUBBYTES[8].a/w1112 ), .B(n15667), .Z(
        \SUBBYTES[8].a/w1102 ) );
  XOR \SUBBYTES[8].a/U4236  ( .A(\w1[8][94] ), .B(\w1[8][93] ), .Z(n15667) );
  XOR \SUBBYTES[8].a/U4235  ( .A(n15669), .B(n15668), .Z(\SUBBYTES[8].a/w1103 ) );
  XOR \SUBBYTES[8].a/U4234  ( .A(n14801), .B(n1073), .Z(n15668) );
  XOR \SUBBYTES[8].a/U4233  ( .A(n14800), .B(\SUBBYTES[8].a/w1056 ), .Z(n15669) );
  XOR \SUBBYTES[8].a/U4232  ( .A(\w1[8][95] ), .B(\w1[8][90] ), .Z(n16027) );
  XOR \SUBBYTES[8].a/U4231  ( .A(n16027), .B(n15670), .Z(\SUBBYTES[8].a/w1104 ) );
  XOR \SUBBYTES[8].a/U4230  ( .A(\w1[8][93] ), .B(\w1[8][92] ), .Z(n15670) );
  XOR \SUBBYTES[8].a/U4229  ( .A(\w1[8][95] ), .B(\SUBBYTES[8].a/w989 ), .Z(
        \SUBBYTES[8].a/w992 ) );
  XOR \SUBBYTES[8].a/U4228  ( .A(\w1[8][89] ), .B(\SUBBYTES[8].a/w989 ), .Z(
        \SUBBYTES[8].a/w993 ) );
  XOR \SUBBYTES[8].a/U4227  ( .A(\w1[8][92] ), .B(\SUBBYTES[8].a/w989 ), .Z(
        \SUBBYTES[8].a/w994 ) );
  XOR \SUBBYTES[8].a/U4226  ( .A(\SUBBYTES[8].a/w993 ), .B(n16027), .Z(
        \SUBBYTES[8].a/w995 ) );
  XOR \SUBBYTES[8].a/U4225  ( .A(n16027), .B(n15671), .Z(\SUBBYTES[8].a/w1080 ) );
  XOR \SUBBYTES[8].a/U4224  ( .A(\w1[8][92] ), .B(\w1[8][89] ), .Z(n15671) );
  XOR \SUBBYTES[8].a/U4223  ( .A(n15673), .B(n15672), .Z(n16024) );
  XOR \SUBBYTES[8].a/U4222  ( .A(\w1[8][92] ), .B(n15674), .Z(n15672) );
  XOR \SUBBYTES[8].a/U4221  ( .A(\SUBBYTES[8].a/w1045 ), .B(\w1[8][94] ), .Z(
        n15673) );
  XOR \SUBBYTES[8].a/U4220  ( .A(\SUBBYTES[8].a/w1019 ), .B(
        \SUBBYTES[8].a/w1026 ), .Z(n15674) );
  XOR \SUBBYTES[8].a/U4219  ( .A(n15676), .B(n15675), .Z(n16022) );
  XOR \SUBBYTES[8].a/U4218  ( .A(\w1[8][89] ), .B(n15677), .Z(n15675) );
  XOR \SUBBYTES[8].a/U4217  ( .A(\SUBBYTES[8].a/w1044 ), .B(\w1[8][93] ), .Z(
        n15676) );
  XOR \SUBBYTES[8].a/U4216  ( .A(\SUBBYTES[8].a/w1020 ), .B(
        \SUBBYTES[8].a/w1027 ), .Z(n15677) );
  XOR \SUBBYTES[8].a/U4215  ( .A(n16024), .B(n16022), .Z(\SUBBYTES[8].a/w1050 ) );
  XOR \SUBBYTES[8].a/U4214  ( .A(\w1[8][93] ), .B(n15678), .Z(n16025) );
  XOR \SUBBYTES[8].a/U4213  ( .A(\SUBBYTES[8].a/w1012 ), .B(
        \SUBBYTES[8].a/w1022 ), .Z(n15678) );
  XOR \SUBBYTES[8].a/U4212  ( .A(n15680), .B(n15679), .Z(\SUBBYTES[8].a/w1037 ) );
  XOR \SUBBYTES[8].a/U4211  ( .A(n16025), .B(n15681), .Z(n15679) );
  XOR \SUBBYTES[8].a/U4210  ( .A(\w1[8][92] ), .B(\SUBBYTES[8].a/w1101 ), .Z(
        n15680) );
  XOR \SUBBYTES[8].a/U4209  ( .A(\SUBBYTES[8].a/w1014 ), .B(
        \SUBBYTES[8].a/w1019 ), .Z(n15681) );
  XOR \SUBBYTES[8].a/U4208  ( .A(n15683), .B(n15682), .Z(n16023) );
  XOR \SUBBYTES[8].a/U4207  ( .A(\SUBBYTES[8].a/w1047 ), .B(\w1[8][95] ), .Z(
        n15682) );
  XOR \SUBBYTES[8].a/U4206  ( .A(\SUBBYTES[8].a/w1022 ), .B(
        \SUBBYTES[8].a/w1029 ), .Z(n15683) );
  XOR \SUBBYTES[8].a/U4205  ( .A(n16022), .B(n16023), .Z(\SUBBYTES[8].a/w1049 ) );
  XOR \SUBBYTES[8].a/U4204  ( .A(\w1[8][91] ), .B(n15684), .Z(n16026) );
  XOR \SUBBYTES[8].a/U4203  ( .A(\SUBBYTES[8].a/w1011 ), .B(
        \SUBBYTES[8].a/w1014 ), .Z(n15684) );
  XOR \SUBBYTES[8].a/U4202  ( .A(n15686), .B(n15685), .Z(\SUBBYTES[8].a/w1038 ) );
  XOR \SUBBYTES[8].a/U4201  ( .A(n16026), .B(n15687), .Z(n15685) );
  XOR \SUBBYTES[8].a/U4200  ( .A(\w1[8][94] ), .B(\SUBBYTES[8].a/w1080 ), .Z(
        n15686) );
  XOR \SUBBYTES[8].a/U4199  ( .A(\SUBBYTES[8].a/w1019 ), .B(
        \SUBBYTES[8].a/w1020 ), .Z(n15687) );
  XOR \SUBBYTES[8].a/U4198  ( .A(n16024), .B(n16023), .Z(\SUBBYTES[8].a/w1058 ) );
  XOR \SUBBYTES[8].a/U4197  ( .A(n15689), .B(n15688), .Z(\SUBBYTES[8].a/w1059 ) );
  XOR \SUBBYTES[8].a/U4196  ( .A(\w1[8][95] ), .B(n16025), .Z(n15688) );
  XOR \SUBBYTES[8].a/U4195  ( .A(\SUBBYTES[8].a/w1011 ), .B(
        \SUBBYTES[8].a/w1020 ), .Z(n15689) );
  XOR \SUBBYTES[8].a/U4194  ( .A(n15691), .B(n15690), .Z(\SUBBYTES[8].a/w1035 ) );
  XOR \SUBBYTES[8].a/U4193  ( .A(n15693), .B(n15692), .Z(n15690) );
  XOR \SUBBYTES[8].a/U4192  ( .A(\w1[8][95] ), .B(\SUBBYTES[8].a/w1119 ), .Z(
        n15691) );
  XOR \SUBBYTES[8].a/U4191  ( .A(\SUBBYTES[8].a/w1026 ), .B(
        \SUBBYTES[8].a/w1029 ), .Z(n15692) );
  XOR \SUBBYTES[8].a/U4190  ( .A(\SUBBYTES[8].a/w1012 ), .B(
        \SUBBYTES[8].a/w1014 ), .Z(n15693) );
  XOR \SUBBYTES[8].a/U4189  ( .A(n15695), .B(n15694), .Z(\SUBBYTES[8].a/w1036 ) );
  XOR \SUBBYTES[8].a/U4188  ( .A(n16026), .B(n15696), .Z(n15694) );
  XOR \SUBBYTES[8].a/U4187  ( .A(\w1[8][93] ), .B(n16027), .Z(n15695) );
  XOR \SUBBYTES[8].a/U4186  ( .A(\SUBBYTES[8].a/w1026 ), .B(
        \SUBBYTES[8].a/w1027 ), .Z(n15696) );
  XOR \SUBBYTES[8].a/U4185  ( .A(n15698), .B(n15697), .Z(\SUBBYTES[8].a/w1052 ) );
  XOR \SUBBYTES[8].a/U4184  ( .A(\w1[8][89] ), .B(n15699), .Z(n15697) );
  XOR \SUBBYTES[8].a/U4183  ( .A(\SUBBYTES[8].a/w1027 ), .B(
        \SUBBYTES[8].a/w1029 ), .Z(n15698) );
  XOR \SUBBYTES[8].a/U4182  ( .A(\SUBBYTES[8].a/w1011 ), .B(
        \SUBBYTES[8].a/w1012 ), .Z(n15699) );
  XOR \SUBBYTES[8].a/U4181  ( .A(\w1[8][97] ), .B(n15700), .Z(n16028) );
  XOR \SUBBYTES[8].a/U4180  ( .A(\w1[8][99] ), .B(\w1[8][98] ), .Z(n15700) );
  XOR \SUBBYTES[8].a/U4179  ( .A(\w1[8][102] ), .B(n16028), .Z(
        \SUBBYTES[8].a/w894 ) );
  XOR \SUBBYTES[8].a/U4178  ( .A(\w1[8][96] ), .B(\SUBBYTES[8].a/w894 ), .Z(
        \SUBBYTES[8].a/w781 ) );
  XOR \SUBBYTES[8].a/U4177  ( .A(\w1[8][96] ), .B(n15701), .Z(
        \SUBBYTES[8].a/w782 ) );
  XOR \SUBBYTES[8].a/U4176  ( .A(\w1[8][102] ), .B(\w1[8][101] ), .Z(n15701)
         );
  XOR \SUBBYTES[8].a/U4175  ( .A(\w1[8][101] ), .B(n16028), .Z(
        \SUBBYTES[8].a/w912 ) );
  XOR \SUBBYTES[8].a/U4174  ( .A(n15703), .B(n15702), .Z(\SUBBYTES[8].a/w905 )
         );
  XOR \SUBBYTES[8].a/U4173  ( .A(\w1[8][99] ), .B(\w1[8][97] ), .Z(n15702) );
  XOR \SUBBYTES[8].a/U4172  ( .A(\w1[8][103] ), .B(\w1[8][100] ), .Z(n15703)
         );
  XOR \SUBBYTES[8].a/U4171  ( .A(\w1[8][96] ), .B(\SUBBYTES[8].a/w905 ), .Z(
        \SUBBYTES[8].a/w784 ) );
  XOR \SUBBYTES[8].a/U4170  ( .A(n15705), .B(n15704), .Z(\SUBBYTES[8].a/w892 )
         );
  XOR \SUBBYTES[8].a/U4169  ( .A(\SUBBYTES[8].a/w853 ), .B(n1072), .Z(n15704)
         );
  XOR \SUBBYTES[8].a/U4168  ( .A(\SUBBYTES[8].a/w846 ), .B(
        \SUBBYTES[8].a/w849 ), .Z(n15705) );
  XOR \SUBBYTES[8].a/U4167  ( .A(n15707), .B(n15706), .Z(\SUBBYTES[8].a/w893 )
         );
  XOR \SUBBYTES[8].a/U4166  ( .A(\SUBBYTES[8].a/w853 ), .B(n14799), .Z(n15706)
         );
  XOR \SUBBYTES[8].a/U4165  ( .A(\SUBBYTES[8].a/w846 ), .B(n14798), .Z(n15707)
         );
  XOR \SUBBYTES[8].a/U4164  ( .A(\SUBBYTES[8].a/w905 ), .B(n15708), .Z(
        \SUBBYTES[8].a/w895 ) );
  XOR \SUBBYTES[8].a/U4163  ( .A(\w1[8][102] ), .B(\w1[8][101] ), .Z(n15708)
         );
  XOR \SUBBYTES[8].a/U4162  ( .A(n15710), .B(n15709), .Z(\SUBBYTES[8].a/w896 )
         );
  XOR \SUBBYTES[8].a/U4161  ( .A(n14799), .B(n1072), .Z(n15709) );
  XOR \SUBBYTES[8].a/U4160  ( .A(n14798), .B(\SUBBYTES[8].a/w849 ), .Z(n15710)
         );
  XOR \SUBBYTES[8].a/U4159  ( .A(\w1[8][103] ), .B(\w1[8][98] ), .Z(n16034) );
  XOR \SUBBYTES[8].a/U4158  ( .A(n16034), .B(n15711), .Z(\SUBBYTES[8].a/w897 )
         );
  XOR \SUBBYTES[8].a/U4157  ( .A(\w1[8][101] ), .B(\w1[8][100] ), .Z(n15711)
         );
  XOR \SUBBYTES[8].a/U4156  ( .A(\w1[8][103] ), .B(\SUBBYTES[8].a/w782 ), .Z(
        \SUBBYTES[8].a/w785 ) );
  XOR \SUBBYTES[8].a/U4155  ( .A(\w1[8][97] ), .B(\SUBBYTES[8].a/w782 ), .Z(
        \SUBBYTES[8].a/w786 ) );
  XOR \SUBBYTES[8].a/U4154  ( .A(\w1[8][100] ), .B(\SUBBYTES[8].a/w782 ), .Z(
        \SUBBYTES[8].a/w787 ) );
  XOR \SUBBYTES[8].a/U4153  ( .A(\SUBBYTES[8].a/w786 ), .B(n16034), .Z(
        \SUBBYTES[8].a/w788 ) );
  XOR \SUBBYTES[8].a/U4152  ( .A(n16034), .B(n15712), .Z(\SUBBYTES[8].a/w873 )
         );
  XOR \SUBBYTES[8].a/U4151  ( .A(\w1[8][100] ), .B(\w1[8][97] ), .Z(n15712) );
  XOR \SUBBYTES[8].a/U4150  ( .A(n15714), .B(n15713), .Z(n16031) );
  XOR \SUBBYTES[8].a/U4149  ( .A(\w1[8][100] ), .B(n15715), .Z(n15713) );
  XOR \SUBBYTES[8].a/U4148  ( .A(\SUBBYTES[8].a/w838 ), .B(\w1[8][102] ), .Z(
        n15714) );
  XOR \SUBBYTES[8].a/U4147  ( .A(\SUBBYTES[8].a/w812 ), .B(
        \SUBBYTES[8].a/w819 ), .Z(n15715) );
  XOR \SUBBYTES[8].a/U4146  ( .A(n15717), .B(n15716), .Z(n16029) );
  XOR \SUBBYTES[8].a/U4145  ( .A(\w1[8][97] ), .B(n15718), .Z(n15716) );
  XOR \SUBBYTES[8].a/U4144  ( .A(\SUBBYTES[8].a/w837 ), .B(\w1[8][101] ), .Z(
        n15717) );
  XOR \SUBBYTES[8].a/U4143  ( .A(\SUBBYTES[8].a/w813 ), .B(
        \SUBBYTES[8].a/w820 ), .Z(n15718) );
  XOR \SUBBYTES[8].a/U4142  ( .A(n16031), .B(n16029), .Z(\SUBBYTES[8].a/w843 )
         );
  XOR \SUBBYTES[8].a/U4141  ( .A(\w1[8][101] ), .B(n15719), .Z(n16032) );
  XOR \SUBBYTES[8].a/U4140  ( .A(\SUBBYTES[8].a/w805 ), .B(
        \SUBBYTES[8].a/w815 ), .Z(n15719) );
  XOR \SUBBYTES[8].a/U4139  ( .A(n15721), .B(n15720), .Z(\SUBBYTES[8].a/w830 )
         );
  XOR \SUBBYTES[8].a/U4138  ( .A(n16032), .B(n15722), .Z(n15720) );
  XOR \SUBBYTES[8].a/U4137  ( .A(\w1[8][100] ), .B(\SUBBYTES[8].a/w894 ), .Z(
        n15721) );
  XOR \SUBBYTES[8].a/U4136  ( .A(\SUBBYTES[8].a/w807 ), .B(
        \SUBBYTES[8].a/w812 ), .Z(n15722) );
  XOR \SUBBYTES[8].a/U4135  ( .A(n15724), .B(n15723), .Z(n16030) );
  XOR \SUBBYTES[8].a/U4134  ( .A(\SUBBYTES[8].a/w840 ), .B(\w1[8][103] ), .Z(
        n15723) );
  XOR \SUBBYTES[8].a/U4133  ( .A(\SUBBYTES[8].a/w815 ), .B(
        \SUBBYTES[8].a/w822 ), .Z(n15724) );
  XOR \SUBBYTES[8].a/U4132  ( .A(n16029), .B(n16030), .Z(\SUBBYTES[8].a/w842 )
         );
  XOR \SUBBYTES[8].a/U4131  ( .A(\w1[8][99] ), .B(n15725), .Z(n16033) );
  XOR \SUBBYTES[8].a/U4130  ( .A(\SUBBYTES[8].a/w804 ), .B(
        \SUBBYTES[8].a/w807 ), .Z(n15725) );
  XOR \SUBBYTES[8].a/U4129  ( .A(n15727), .B(n15726), .Z(\SUBBYTES[8].a/w831 )
         );
  XOR \SUBBYTES[8].a/U4128  ( .A(n16033), .B(n15728), .Z(n15726) );
  XOR \SUBBYTES[8].a/U4127  ( .A(\w1[8][102] ), .B(\SUBBYTES[8].a/w873 ), .Z(
        n15727) );
  XOR \SUBBYTES[8].a/U4126  ( .A(\SUBBYTES[8].a/w812 ), .B(
        \SUBBYTES[8].a/w813 ), .Z(n15728) );
  XOR \SUBBYTES[8].a/U4125  ( .A(n16031), .B(n16030), .Z(\SUBBYTES[8].a/w851 )
         );
  XOR \SUBBYTES[8].a/U4124  ( .A(n15730), .B(n15729), .Z(\SUBBYTES[8].a/w852 )
         );
  XOR \SUBBYTES[8].a/U4123  ( .A(\w1[8][103] ), .B(n16032), .Z(n15729) );
  XOR \SUBBYTES[8].a/U4122  ( .A(\SUBBYTES[8].a/w804 ), .B(
        \SUBBYTES[8].a/w813 ), .Z(n15730) );
  XOR \SUBBYTES[8].a/U4121  ( .A(n15732), .B(n15731), .Z(\SUBBYTES[8].a/w828 )
         );
  XOR \SUBBYTES[8].a/U4120  ( .A(n15734), .B(n15733), .Z(n15731) );
  XOR \SUBBYTES[8].a/U4119  ( .A(\w1[8][103] ), .B(\SUBBYTES[8].a/w912 ), .Z(
        n15732) );
  XOR \SUBBYTES[8].a/U4118  ( .A(\SUBBYTES[8].a/w819 ), .B(
        \SUBBYTES[8].a/w822 ), .Z(n15733) );
  XOR \SUBBYTES[8].a/U4117  ( .A(\SUBBYTES[8].a/w805 ), .B(
        \SUBBYTES[8].a/w807 ), .Z(n15734) );
  XOR \SUBBYTES[8].a/U4116  ( .A(n15736), .B(n15735), .Z(\SUBBYTES[8].a/w829 )
         );
  XOR \SUBBYTES[8].a/U4115  ( .A(n16033), .B(n15737), .Z(n15735) );
  XOR \SUBBYTES[8].a/U4114  ( .A(\w1[8][101] ), .B(n16034), .Z(n15736) );
  XOR \SUBBYTES[8].a/U4113  ( .A(\SUBBYTES[8].a/w819 ), .B(
        \SUBBYTES[8].a/w820 ), .Z(n15737) );
  XOR \SUBBYTES[8].a/U4112  ( .A(n15739), .B(n15738), .Z(\SUBBYTES[8].a/w845 )
         );
  XOR \SUBBYTES[8].a/U4111  ( .A(\w1[8][97] ), .B(n15740), .Z(n15738) );
  XOR \SUBBYTES[8].a/U4110  ( .A(\SUBBYTES[8].a/w820 ), .B(
        \SUBBYTES[8].a/w822 ), .Z(n15739) );
  XOR \SUBBYTES[8].a/U4109  ( .A(\SUBBYTES[8].a/w804 ), .B(
        \SUBBYTES[8].a/w805 ), .Z(n15740) );
  XOR \SUBBYTES[8].a/U4108  ( .A(\w1[8][105] ), .B(n15741), .Z(n16035) );
  XOR \SUBBYTES[8].a/U4107  ( .A(\w1[8][107] ), .B(\w1[8][106] ), .Z(n15741)
         );
  XOR \SUBBYTES[8].a/U4106  ( .A(\w1[8][110] ), .B(n16035), .Z(
        \SUBBYTES[8].a/w687 ) );
  XOR \SUBBYTES[8].a/U4105  ( .A(\w1[8][104] ), .B(\SUBBYTES[8].a/w687 ), .Z(
        \SUBBYTES[8].a/w574 ) );
  XOR \SUBBYTES[8].a/U4104  ( .A(\w1[8][104] ), .B(n15742), .Z(
        \SUBBYTES[8].a/w575 ) );
  XOR \SUBBYTES[8].a/U4103  ( .A(\w1[8][110] ), .B(\w1[8][109] ), .Z(n15742)
         );
  XOR \SUBBYTES[8].a/U4102  ( .A(\w1[8][109] ), .B(n16035), .Z(
        \SUBBYTES[8].a/w705 ) );
  XOR \SUBBYTES[8].a/U4101  ( .A(n15744), .B(n15743), .Z(\SUBBYTES[8].a/w698 )
         );
  XOR \SUBBYTES[8].a/U4100  ( .A(\w1[8][107] ), .B(\w1[8][105] ), .Z(n15743)
         );
  XOR \SUBBYTES[8].a/U4099  ( .A(\w1[8][111] ), .B(\w1[8][108] ), .Z(n15744)
         );
  XOR \SUBBYTES[8].a/U4098  ( .A(\w1[8][104] ), .B(\SUBBYTES[8].a/w698 ), .Z(
        \SUBBYTES[8].a/w577 ) );
  XOR \SUBBYTES[8].a/U4097  ( .A(n15746), .B(n15745), .Z(\SUBBYTES[8].a/w685 )
         );
  XOR \SUBBYTES[8].a/U4096  ( .A(\SUBBYTES[8].a/w646 ), .B(n1071), .Z(n15745)
         );
  XOR \SUBBYTES[8].a/U4095  ( .A(\SUBBYTES[8].a/w639 ), .B(
        \SUBBYTES[8].a/w642 ), .Z(n15746) );
  XOR \SUBBYTES[8].a/U4094  ( .A(n15748), .B(n15747), .Z(\SUBBYTES[8].a/w686 )
         );
  XOR \SUBBYTES[8].a/U4093  ( .A(\SUBBYTES[8].a/w646 ), .B(n14797), .Z(n15747)
         );
  XOR \SUBBYTES[8].a/U4092  ( .A(\SUBBYTES[8].a/w639 ), .B(n14796), .Z(n15748)
         );
  XOR \SUBBYTES[8].a/U4091  ( .A(\SUBBYTES[8].a/w698 ), .B(n15749), .Z(
        \SUBBYTES[8].a/w688 ) );
  XOR \SUBBYTES[8].a/U4090  ( .A(\w1[8][110] ), .B(\w1[8][109] ), .Z(n15749)
         );
  XOR \SUBBYTES[8].a/U4089  ( .A(n15751), .B(n15750), .Z(\SUBBYTES[8].a/w689 )
         );
  XOR \SUBBYTES[8].a/U4088  ( .A(n14797), .B(n1071), .Z(n15750) );
  XOR \SUBBYTES[8].a/U4087  ( .A(n14796), .B(\SUBBYTES[8].a/w642 ), .Z(n15751)
         );
  XOR \SUBBYTES[8].a/U4086  ( .A(\w1[8][111] ), .B(\w1[8][106] ), .Z(n16041)
         );
  XOR \SUBBYTES[8].a/U4085  ( .A(n16041), .B(n15752), .Z(\SUBBYTES[8].a/w690 )
         );
  XOR \SUBBYTES[8].a/U4084  ( .A(\w1[8][109] ), .B(\w1[8][108] ), .Z(n15752)
         );
  XOR \SUBBYTES[8].a/U4083  ( .A(\w1[8][111] ), .B(\SUBBYTES[8].a/w575 ), .Z(
        \SUBBYTES[8].a/w578 ) );
  XOR \SUBBYTES[8].a/U4082  ( .A(\w1[8][105] ), .B(\SUBBYTES[8].a/w575 ), .Z(
        \SUBBYTES[8].a/w579 ) );
  XOR \SUBBYTES[8].a/U4081  ( .A(\w1[8][108] ), .B(\SUBBYTES[8].a/w575 ), .Z(
        \SUBBYTES[8].a/w580 ) );
  XOR \SUBBYTES[8].a/U4080  ( .A(\SUBBYTES[8].a/w579 ), .B(n16041), .Z(
        \SUBBYTES[8].a/w581 ) );
  XOR \SUBBYTES[8].a/U4079  ( .A(n16041), .B(n15753), .Z(\SUBBYTES[8].a/w666 )
         );
  XOR \SUBBYTES[8].a/U4078  ( .A(\w1[8][108] ), .B(\w1[8][105] ), .Z(n15753)
         );
  XOR \SUBBYTES[8].a/U4077  ( .A(n15755), .B(n15754), .Z(n16038) );
  XOR \SUBBYTES[8].a/U4076  ( .A(\w1[8][108] ), .B(n15756), .Z(n15754) );
  XOR \SUBBYTES[8].a/U4075  ( .A(\SUBBYTES[8].a/w631 ), .B(\w1[8][110] ), .Z(
        n15755) );
  XOR \SUBBYTES[8].a/U4074  ( .A(\SUBBYTES[8].a/w605 ), .B(
        \SUBBYTES[8].a/w612 ), .Z(n15756) );
  XOR \SUBBYTES[8].a/U4073  ( .A(n15758), .B(n15757), .Z(n16036) );
  XOR \SUBBYTES[8].a/U4072  ( .A(\w1[8][105] ), .B(n15759), .Z(n15757) );
  XOR \SUBBYTES[8].a/U4071  ( .A(\SUBBYTES[8].a/w630 ), .B(\w1[8][109] ), .Z(
        n15758) );
  XOR \SUBBYTES[8].a/U4070  ( .A(\SUBBYTES[8].a/w606 ), .B(
        \SUBBYTES[8].a/w613 ), .Z(n15759) );
  XOR \SUBBYTES[8].a/U4069  ( .A(n16038), .B(n16036), .Z(\SUBBYTES[8].a/w636 )
         );
  XOR \SUBBYTES[8].a/U4068  ( .A(\w1[8][109] ), .B(n15760), .Z(n16039) );
  XOR \SUBBYTES[8].a/U4067  ( .A(\SUBBYTES[8].a/w598 ), .B(
        \SUBBYTES[8].a/w608 ), .Z(n15760) );
  XOR \SUBBYTES[8].a/U4066  ( .A(n15762), .B(n15761), .Z(\SUBBYTES[8].a/w623 )
         );
  XOR \SUBBYTES[8].a/U4065  ( .A(n16039), .B(n15763), .Z(n15761) );
  XOR \SUBBYTES[8].a/U4064  ( .A(\w1[8][108] ), .B(\SUBBYTES[8].a/w687 ), .Z(
        n15762) );
  XOR \SUBBYTES[8].a/U4063  ( .A(\SUBBYTES[8].a/w600 ), .B(
        \SUBBYTES[8].a/w605 ), .Z(n15763) );
  XOR \SUBBYTES[8].a/U4062  ( .A(n15765), .B(n15764), .Z(n16037) );
  XOR \SUBBYTES[8].a/U4061  ( .A(\SUBBYTES[8].a/w633 ), .B(\w1[8][111] ), .Z(
        n15764) );
  XOR \SUBBYTES[8].a/U4060  ( .A(\SUBBYTES[8].a/w608 ), .B(
        \SUBBYTES[8].a/w615 ), .Z(n15765) );
  XOR \SUBBYTES[8].a/U4059  ( .A(n16036), .B(n16037), .Z(\SUBBYTES[8].a/w635 )
         );
  XOR \SUBBYTES[8].a/U4058  ( .A(\w1[8][107] ), .B(n15766), .Z(n16040) );
  XOR \SUBBYTES[8].a/U4057  ( .A(\SUBBYTES[8].a/w597 ), .B(
        \SUBBYTES[8].a/w600 ), .Z(n15766) );
  XOR \SUBBYTES[8].a/U4056  ( .A(n15768), .B(n15767), .Z(\SUBBYTES[8].a/w624 )
         );
  XOR \SUBBYTES[8].a/U4055  ( .A(n16040), .B(n15769), .Z(n15767) );
  XOR \SUBBYTES[8].a/U4054  ( .A(\w1[8][110] ), .B(\SUBBYTES[8].a/w666 ), .Z(
        n15768) );
  XOR \SUBBYTES[8].a/U4053  ( .A(\SUBBYTES[8].a/w605 ), .B(
        \SUBBYTES[8].a/w606 ), .Z(n15769) );
  XOR \SUBBYTES[8].a/U4052  ( .A(n16038), .B(n16037), .Z(\SUBBYTES[8].a/w644 )
         );
  XOR \SUBBYTES[8].a/U4051  ( .A(n15771), .B(n15770), .Z(\SUBBYTES[8].a/w645 )
         );
  XOR \SUBBYTES[8].a/U4050  ( .A(\w1[8][111] ), .B(n16039), .Z(n15770) );
  XOR \SUBBYTES[8].a/U4049  ( .A(\SUBBYTES[8].a/w597 ), .B(
        \SUBBYTES[8].a/w606 ), .Z(n15771) );
  XOR \SUBBYTES[8].a/U4048  ( .A(n15773), .B(n15772), .Z(\SUBBYTES[8].a/w621 )
         );
  XOR \SUBBYTES[8].a/U4047  ( .A(n15775), .B(n15774), .Z(n15772) );
  XOR \SUBBYTES[8].a/U4046  ( .A(\w1[8][111] ), .B(\SUBBYTES[8].a/w705 ), .Z(
        n15773) );
  XOR \SUBBYTES[8].a/U4045  ( .A(\SUBBYTES[8].a/w612 ), .B(
        \SUBBYTES[8].a/w615 ), .Z(n15774) );
  XOR \SUBBYTES[8].a/U4044  ( .A(\SUBBYTES[8].a/w598 ), .B(
        \SUBBYTES[8].a/w600 ), .Z(n15775) );
  XOR \SUBBYTES[8].a/U4043  ( .A(n15777), .B(n15776), .Z(\SUBBYTES[8].a/w622 )
         );
  XOR \SUBBYTES[8].a/U4042  ( .A(n16040), .B(n15778), .Z(n15776) );
  XOR \SUBBYTES[8].a/U4041  ( .A(\w1[8][109] ), .B(n16041), .Z(n15777) );
  XOR \SUBBYTES[8].a/U4040  ( .A(\SUBBYTES[8].a/w612 ), .B(
        \SUBBYTES[8].a/w613 ), .Z(n15778) );
  XOR \SUBBYTES[8].a/U4039  ( .A(n15780), .B(n15779), .Z(\SUBBYTES[8].a/w638 )
         );
  XOR \SUBBYTES[8].a/U4038  ( .A(\w1[8][105] ), .B(n15781), .Z(n15779) );
  XOR \SUBBYTES[8].a/U4037  ( .A(\SUBBYTES[8].a/w613 ), .B(
        \SUBBYTES[8].a/w615 ), .Z(n15780) );
  XOR \SUBBYTES[8].a/U4036  ( .A(\SUBBYTES[8].a/w597 ), .B(
        \SUBBYTES[8].a/w598 ), .Z(n15781) );
  XOR \SUBBYTES[8].a/U4035  ( .A(\w1[8][113] ), .B(n15782), .Z(n16042) );
  XOR \SUBBYTES[8].a/U4034  ( .A(\w1[8][115] ), .B(\w1[8][114] ), .Z(n15782)
         );
  XOR \SUBBYTES[8].a/U4033  ( .A(\w1[8][118] ), .B(n16042), .Z(
        \SUBBYTES[8].a/w480 ) );
  XOR \SUBBYTES[8].a/U4032  ( .A(\w1[8][112] ), .B(\SUBBYTES[8].a/w480 ), .Z(
        \SUBBYTES[8].a/w367 ) );
  XOR \SUBBYTES[8].a/U4031  ( .A(\w1[8][112] ), .B(n15783), .Z(
        \SUBBYTES[8].a/w368 ) );
  XOR \SUBBYTES[8].a/U4030  ( .A(\w1[8][118] ), .B(\w1[8][117] ), .Z(n15783)
         );
  XOR \SUBBYTES[8].a/U4029  ( .A(\w1[8][117] ), .B(n16042), .Z(
        \SUBBYTES[8].a/w498 ) );
  XOR \SUBBYTES[8].a/U4028  ( .A(n15785), .B(n15784), .Z(\SUBBYTES[8].a/w491 )
         );
  XOR \SUBBYTES[8].a/U4027  ( .A(\w1[8][115] ), .B(\w1[8][113] ), .Z(n15784)
         );
  XOR \SUBBYTES[8].a/U4026  ( .A(\w1[8][119] ), .B(\w1[8][116] ), .Z(n15785)
         );
  XOR \SUBBYTES[8].a/U4025  ( .A(\w1[8][112] ), .B(\SUBBYTES[8].a/w491 ), .Z(
        \SUBBYTES[8].a/w370 ) );
  XOR \SUBBYTES[8].a/U4024  ( .A(n15787), .B(n15786), .Z(\SUBBYTES[8].a/w478 )
         );
  XOR \SUBBYTES[8].a/U4023  ( .A(\SUBBYTES[8].a/w439 ), .B(n1070), .Z(n15786)
         );
  XOR \SUBBYTES[8].a/U4022  ( .A(\SUBBYTES[8].a/w432 ), .B(
        \SUBBYTES[8].a/w435 ), .Z(n15787) );
  XOR \SUBBYTES[8].a/U4021  ( .A(n15789), .B(n15788), .Z(\SUBBYTES[8].a/w479 )
         );
  XOR \SUBBYTES[8].a/U4020  ( .A(\SUBBYTES[8].a/w439 ), .B(n14795), .Z(n15788)
         );
  XOR \SUBBYTES[8].a/U4019  ( .A(\SUBBYTES[8].a/w432 ), .B(n14794), .Z(n15789)
         );
  XOR \SUBBYTES[8].a/U4018  ( .A(\SUBBYTES[8].a/w491 ), .B(n15790), .Z(
        \SUBBYTES[8].a/w481 ) );
  XOR \SUBBYTES[8].a/U4017  ( .A(\w1[8][118] ), .B(\w1[8][117] ), .Z(n15790)
         );
  XOR \SUBBYTES[8].a/U4016  ( .A(n15792), .B(n15791), .Z(\SUBBYTES[8].a/w482 )
         );
  XOR \SUBBYTES[8].a/U4015  ( .A(n14795), .B(n1070), .Z(n15791) );
  XOR \SUBBYTES[8].a/U4014  ( .A(n14794), .B(\SUBBYTES[8].a/w435 ), .Z(n15792)
         );
  XOR \SUBBYTES[8].a/U4013  ( .A(\w1[8][119] ), .B(\w1[8][114] ), .Z(n16048)
         );
  XOR \SUBBYTES[8].a/U4012  ( .A(n16048), .B(n15793), .Z(\SUBBYTES[8].a/w483 )
         );
  XOR \SUBBYTES[8].a/U4011  ( .A(\w1[8][117] ), .B(\w1[8][116] ), .Z(n15793)
         );
  XOR \SUBBYTES[8].a/U4010  ( .A(\w1[8][119] ), .B(\SUBBYTES[8].a/w368 ), .Z(
        \SUBBYTES[8].a/w371 ) );
  XOR \SUBBYTES[8].a/U4009  ( .A(\w1[8][113] ), .B(\SUBBYTES[8].a/w368 ), .Z(
        \SUBBYTES[8].a/w372 ) );
  XOR \SUBBYTES[8].a/U4008  ( .A(\w1[8][116] ), .B(\SUBBYTES[8].a/w368 ), .Z(
        \SUBBYTES[8].a/w373 ) );
  XOR \SUBBYTES[8].a/U4007  ( .A(\SUBBYTES[8].a/w372 ), .B(n16048), .Z(
        \SUBBYTES[8].a/w374 ) );
  XOR \SUBBYTES[8].a/U4006  ( .A(n16048), .B(n15794), .Z(\SUBBYTES[8].a/w459 )
         );
  XOR \SUBBYTES[8].a/U4005  ( .A(\w1[8][116] ), .B(\w1[8][113] ), .Z(n15794)
         );
  XOR \SUBBYTES[8].a/U4004  ( .A(n15796), .B(n15795), .Z(n16045) );
  XOR \SUBBYTES[8].a/U4003  ( .A(\w1[8][116] ), .B(n15797), .Z(n15795) );
  XOR \SUBBYTES[8].a/U4002  ( .A(\SUBBYTES[8].a/w424 ), .B(\w1[8][118] ), .Z(
        n15796) );
  XOR \SUBBYTES[8].a/U4001  ( .A(\SUBBYTES[8].a/w398 ), .B(
        \SUBBYTES[8].a/w405 ), .Z(n15797) );
  XOR \SUBBYTES[8].a/U4000  ( .A(n15799), .B(n15798), .Z(n16043) );
  XOR \SUBBYTES[8].a/U3999  ( .A(\w1[8][113] ), .B(n15800), .Z(n15798) );
  XOR \SUBBYTES[8].a/U3998  ( .A(\SUBBYTES[8].a/w423 ), .B(\w1[8][117] ), .Z(
        n15799) );
  XOR \SUBBYTES[8].a/U3997  ( .A(\SUBBYTES[8].a/w399 ), .B(
        \SUBBYTES[8].a/w406 ), .Z(n15800) );
  XOR \SUBBYTES[8].a/U3996  ( .A(n16045), .B(n16043), .Z(\SUBBYTES[8].a/w429 )
         );
  XOR \SUBBYTES[8].a/U3995  ( .A(\w1[8][117] ), .B(n15801), .Z(n16046) );
  XOR \SUBBYTES[8].a/U3994  ( .A(\SUBBYTES[8].a/w391 ), .B(
        \SUBBYTES[8].a/w401 ), .Z(n15801) );
  XOR \SUBBYTES[8].a/U3993  ( .A(n15803), .B(n15802), .Z(\SUBBYTES[8].a/w416 )
         );
  XOR \SUBBYTES[8].a/U3992  ( .A(n16046), .B(n15804), .Z(n15802) );
  XOR \SUBBYTES[8].a/U3991  ( .A(\w1[8][116] ), .B(\SUBBYTES[8].a/w480 ), .Z(
        n15803) );
  XOR \SUBBYTES[8].a/U3990  ( .A(\SUBBYTES[8].a/w393 ), .B(
        \SUBBYTES[8].a/w398 ), .Z(n15804) );
  XOR \SUBBYTES[8].a/U3989  ( .A(n15806), .B(n15805), .Z(n16044) );
  XOR \SUBBYTES[8].a/U3988  ( .A(\SUBBYTES[8].a/w426 ), .B(\w1[8][119] ), .Z(
        n15805) );
  XOR \SUBBYTES[8].a/U3987  ( .A(\SUBBYTES[8].a/w401 ), .B(
        \SUBBYTES[8].a/w408 ), .Z(n15806) );
  XOR \SUBBYTES[8].a/U3986  ( .A(n16043), .B(n16044), .Z(\SUBBYTES[8].a/w428 )
         );
  XOR \SUBBYTES[8].a/U3985  ( .A(\w1[8][115] ), .B(n15807), .Z(n16047) );
  XOR \SUBBYTES[8].a/U3984  ( .A(\SUBBYTES[8].a/w390 ), .B(
        \SUBBYTES[8].a/w393 ), .Z(n15807) );
  XOR \SUBBYTES[8].a/U3983  ( .A(n15809), .B(n15808), .Z(\SUBBYTES[8].a/w417 )
         );
  XOR \SUBBYTES[8].a/U3982  ( .A(n16047), .B(n15810), .Z(n15808) );
  XOR \SUBBYTES[8].a/U3981  ( .A(\w1[8][118] ), .B(\SUBBYTES[8].a/w459 ), .Z(
        n15809) );
  XOR \SUBBYTES[8].a/U3980  ( .A(\SUBBYTES[8].a/w398 ), .B(
        \SUBBYTES[8].a/w399 ), .Z(n15810) );
  XOR \SUBBYTES[8].a/U3979  ( .A(n16045), .B(n16044), .Z(\SUBBYTES[8].a/w437 )
         );
  XOR \SUBBYTES[8].a/U3978  ( .A(n15812), .B(n15811), .Z(\SUBBYTES[8].a/w438 )
         );
  XOR \SUBBYTES[8].a/U3977  ( .A(\w1[8][119] ), .B(n16046), .Z(n15811) );
  XOR \SUBBYTES[8].a/U3976  ( .A(\SUBBYTES[8].a/w390 ), .B(
        \SUBBYTES[8].a/w399 ), .Z(n15812) );
  XOR \SUBBYTES[8].a/U3975  ( .A(n15814), .B(n15813), .Z(\SUBBYTES[8].a/w414 )
         );
  XOR \SUBBYTES[8].a/U3974  ( .A(n15816), .B(n15815), .Z(n15813) );
  XOR \SUBBYTES[8].a/U3973  ( .A(\w1[8][119] ), .B(\SUBBYTES[8].a/w498 ), .Z(
        n15814) );
  XOR \SUBBYTES[8].a/U3972  ( .A(\SUBBYTES[8].a/w405 ), .B(
        \SUBBYTES[8].a/w408 ), .Z(n15815) );
  XOR \SUBBYTES[8].a/U3971  ( .A(\SUBBYTES[8].a/w391 ), .B(
        \SUBBYTES[8].a/w393 ), .Z(n15816) );
  XOR \SUBBYTES[8].a/U3970  ( .A(n15818), .B(n15817), .Z(\SUBBYTES[8].a/w415 )
         );
  XOR \SUBBYTES[8].a/U3969  ( .A(n16047), .B(n15819), .Z(n15817) );
  XOR \SUBBYTES[8].a/U3968  ( .A(\w1[8][117] ), .B(n16048), .Z(n15818) );
  XOR \SUBBYTES[8].a/U3967  ( .A(\SUBBYTES[8].a/w405 ), .B(
        \SUBBYTES[8].a/w406 ), .Z(n15819) );
  XOR \SUBBYTES[8].a/U3966  ( .A(n15821), .B(n15820), .Z(\SUBBYTES[8].a/w431 )
         );
  XOR \SUBBYTES[8].a/U3965  ( .A(\w1[8][113] ), .B(n15822), .Z(n15820) );
  XOR \SUBBYTES[8].a/U3964  ( .A(\SUBBYTES[8].a/w406 ), .B(
        \SUBBYTES[8].a/w408 ), .Z(n15821) );
  XOR \SUBBYTES[8].a/U3963  ( .A(\SUBBYTES[8].a/w390 ), .B(
        \SUBBYTES[8].a/w391 ), .Z(n15822) );
  XOR \SUBBYTES[8].a/U3962  ( .A(\w1[8][121] ), .B(n15823), .Z(n16049) );
  XOR \SUBBYTES[8].a/U3961  ( .A(\w1[8][123] ), .B(\w1[8][122] ), .Z(n15823)
         );
  XOR \SUBBYTES[8].a/U3960  ( .A(\w1[8][126] ), .B(n16049), .Z(
        \SUBBYTES[8].a/w273 ) );
  XOR \SUBBYTES[8].a/U3959  ( .A(\w1[8][120] ), .B(\SUBBYTES[8].a/w273 ), .Z(
        \SUBBYTES[8].a/w160 ) );
  XOR \SUBBYTES[8].a/U3958  ( .A(\w1[8][120] ), .B(n15824), .Z(
        \SUBBYTES[8].a/w161 ) );
  XOR \SUBBYTES[8].a/U3957  ( .A(\w1[8][126] ), .B(\w1[8][125] ), .Z(n15824)
         );
  XOR \SUBBYTES[8].a/U3956  ( .A(\w1[8][125] ), .B(n16049), .Z(
        \SUBBYTES[8].a/w291 ) );
  XOR \SUBBYTES[8].a/U3955  ( .A(n15826), .B(n15825), .Z(\SUBBYTES[8].a/w284 )
         );
  XOR \SUBBYTES[8].a/U3954  ( .A(\w1[8][123] ), .B(\w1[8][121] ), .Z(n15825)
         );
  XOR \SUBBYTES[8].a/U3953  ( .A(\w1[8][127] ), .B(\w1[8][124] ), .Z(n15826)
         );
  XOR \SUBBYTES[8].a/U3952  ( .A(\w1[8][120] ), .B(\SUBBYTES[8].a/w284 ), .Z(
        \SUBBYTES[8].a/w163 ) );
  XOR \SUBBYTES[8].a/U3951  ( .A(n15828), .B(n15827), .Z(\SUBBYTES[8].a/w271 )
         );
  XOR \SUBBYTES[8].a/U3950  ( .A(\SUBBYTES[8].a/w232 ), .B(n1069), .Z(n15827)
         );
  XOR \SUBBYTES[8].a/U3949  ( .A(\SUBBYTES[8].a/w225 ), .B(
        \SUBBYTES[8].a/w228 ), .Z(n15828) );
  XOR \SUBBYTES[8].a/U3948  ( .A(n15830), .B(n15829), .Z(\SUBBYTES[8].a/w272 )
         );
  XOR \SUBBYTES[8].a/U3947  ( .A(\SUBBYTES[8].a/w232 ), .B(n14793), .Z(n15829)
         );
  XOR \SUBBYTES[8].a/U3946  ( .A(\SUBBYTES[8].a/w225 ), .B(n14792), .Z(n15830)
         );
  XOR \SUBBYTES[8].a/U3945  ( .A(\SUBBYTES[8].a/w284 ), .B(n15831), .Z(
        \SUBBYTES[8].a/w274 ) );
  XOR \SUBBYTES[8].a/U3944  ( .A(\w1[8][126] ), .B(\w1[8][125] ), .Z(n15831)
         );
  XOR \SUBBYTES[8].a/U3943  ( .A(n15833), .B(n15832), .Z(\SUBBYTES[8].a/w275 )
         );
  XOR \SUBBYTES[8].a/U3942  ( .A(n14793), .B(n1069), .Z(n15832) );
  XOR \SUBBYTES[8].a/U3941  ( .A(n14792), .B(\SUBBYTES[8].a/w228 ), .Z(n15833)
         );
  XOR \SUBBYTES[8].a/U3940  ( .A(\w1[8][127] ), .B(\w1[8][122] ), .Z(n16055)
         );
  XOR \SUBBYTES[8].a/U3939  ( .A(n16055), .B(n15834), .Z(\SUBBYTES[8].a/w276 )
         );
  XOR \SUBBYTES[8].a/U3938  ( .A(\w1[8][125] ), .B(\w1[8][124] ), .Z(n15834)
         );
  XOR \SUBBYTES[8].a/U3937  ( .A(\w1[8][127] ), .B(\SUBBYTES[8].a/w161 ), .Z(
        \SUBBYTES[8].a/w164 ) );
  XOR \SUBBYTES[8].a/U3936  ( .A(\w1[8][121] ), .B(\SUBBYTES[8].a/w161 ), .Z(
        \SUBBYTES[8].a/w165 ) );
  XOR \SUBBYTES[8].a/U3935  ( .A(\w1[8][124] ), .B(\SUBBYTES[8].a/w161 ), .Z(
        \SUBBYTES[8].a/w166 ) );
  XOR \SUBBYTES[8].a/U3934  ( .A(\SUBBYTES[8].a/w165 ), .B(n16055), .Z(
        \SUBBYTES[8].a/w167 ) );
  XOR \SUBBYTES[8].a/U3933  ( .A(n16055), .B(n15835), .Z(\SUBBYTES[8].a/w252 )
         );
  XOR \SUBBYTES[8].a/U3932  ( .A(\w1[8][124] ), .B(\w1[8][121] ), .Z(n15835)
         );
  XOR \SUBBYTES[8].a/U3931  ( .A(n15837), .B(n15836), .Z(n16052) );
  XOR \SUBBYTES[8].a/U3930  ( .A(\w1[8][124] ), .B(n15838), .Z(n15836) );
  XOR \SUBBYTES[8].a/U3929  ( .A(\SUBBYTES[8].a/w217 ), .B(\w1[8][126] ), .Z(
        n15837) );
  XOR \SUBBYTES[8].a/U3928  ( .A(\SUBBYTES[8].a/w191 ), .B(
        \SUBBYTES[8].a/w198 ), .Z(n15838) );
  XOR \SUBBYTES[8].a/U3927  ( .A(n15840), .B(n15839), .Z(n16050) );
  XOR \SUBBYTES[8].a/U3926  ( .A(\w1[8][121] ), .B(n15841), .Z(n15839) );
  XOR \SUBBYTES[8].a/U3925  ( .A(\SUBBYTES[8].a/w216 ), .B(\w1[8][125] ), .Z(
        n15840) );
  XOR \SUBBYTES[8].a/U3924  ( .A(\SUBBYTES[8].a/w192 ), .B(
        \SUBBYTES[8].a/w199 ), .Z(n15841) );
  XOR \SUBBYTES[8].a/U3923  ( .A(n16052), .B(n16050), .Z(\SUBBYTES[8].a/w222 )
         );
  XOR \SUBBYTES[8].a/U3922  ( .A(\w1[8][125] ), .B(n15842), .Z(n16053) );
  XOR \SUBBYTES[8].a/U3921  ( .A(\SUBBYTES[8].a/w184 ), .B(
        \SUBBYTES[8].a/w194 ), .Z(n15842) );
  XOR \SUBBYTES[8].a/U3920  ( .A(n15844), .B(n15843), .Z(\SUBBYTES[8].a/w209 )
         );
  XOR \SUBBYTES[8].a/U3919  ( .A(n16053), .B(n15845), .Z(n15843) );
  XOR \SUBBYTES[8].a/U3918  ( .A(\w1[8][124] ), .B(\SUBBYTES[8].a/w273 ), .Z(
        n15844) );
  XOR \SUBBYTES[8].a/U3917  ( .A(\SUBBYTES[8].a/w186 ), .B(
        \SUBBYTES[8].a/w191 ), .Z(n15845) );
  XOR \SUBBYTES[8].a/U3916  ( .A(n15847), .B(n15846), .Z(n16051) );
  XOR \SUBBYTES[8].a/U3915  ( .A(\SUBBYTES[8].a/w219 ), .B(\w1[8][127] ), .Z(
        n15846) );
  XOR \SUBBYTES[8].a/U3914  ( .A(\SUBBYTES[8].a/w194 ), .B(
        \SUBBYTES[8].a/w201 ), .Z(n15847) );
  XOR \SUBBYTES[8].a/U3913  ( .A(n16050), .B(n16051), .Z(\SUBBYTES[8].a/w221 )
         );
  XOR \SUBBYTES[8].a/U3912  ( .A(\w1[8][123] ), .B(n15848), .Z(n16054) );
  XOR \SUBBYTES[8].a/U3911  ( .A(\SUBBYTES[8].a/w183 ), .B(
        \SUBBYTES[8].a/w186 ), .Z(n15848) );
  XOR \SUBBYTES[8].a/U3910  ( .A(n15850), .B(n15849), .Z(\SUBBYTES[8].a/w210 )
         );
  XOR \SUBBYTES[8].a/U3909  ( .A(n16054), .B(n15851), .Z(n15849) );
  XOR \SUBBYTES[8].a/U3908  ( .A(\w1[8][126] ), .B(\SUBBYTES[8].a/w252 ), .Z(
        n15850) );
  XOR \SUBBYTES[8].a/U3907  ( .A(\SUBBYTES[8].a/w191 ), .B(
        \SUBBYTES[8].a/w192 ), .Z(n15851) );
  XOR \SUBBYTES[8].a/U3906  ( .A(n16052), .B(n16051), .Z(\SUBBYTES[8].a/w230 )
         );
  XOR \SUBBYTES[8].a/U3905  ( .A(n15853), .B(n15852), .Z(\SUBBYTES[8].a/w231 )
         );
  XOR \SUBBYTES[8].a/U3904  ( .A(\w1[8][127] ), .B(n16053), .Z(n15852) );
  XOR \SUBBYTES[8].a/U3903  ( .A(\SUBBYTES[8].a/w183 ), .B(
        \SUBBYTES[8].a/w192 ), .Z(n15853) );
  XOR \SUBBYTES[8].a/U3902  ( .A(n15855), .B(n15854), .Z(\SUBBYTES[8].a/w207 )
         );
  XOR \SUBBYTES[8].a/U3901  ( .A(n15857), .B(n15856), .Z(n15854) );
  XOR \SUBBYTES[8].a/U3900  ( .A(\w1[8][127] ), .B(\SUBBYTES[8].a/w291 ), .Z(
        n15855) );
  XOR \SUBBYTES[8].a/U3899  ( .A(\SUBBYTES[8].a/w198 ), .B(
        \SUBBYTES[8].a/w201 ), .Z(n15856) );
  XOR \SUBBYTES[8].a/U3898  ( .A(\SUBBYTES[8].a/w184 ), .B(
        \SUBBYTES[8].a/w186 ), .Z(n15857) );
  XOR \SUBBYTES[8].a/U3897  ( .A(n15859), .B(n15858), .Z(\SUBBYTES[8].a/w208 )
         );
  XOR \SUBBYTES[8].a/U3896  ( .A(n16054), .B(n15860), .Z(n15858) );
  XOR \SUBBYTES[8].a/U3895  ( .A(\w1[8][125] ), .B(n16055), .Z(n15859) );
  XOR \SUBBYTES[8].a/U3894  ( .A(\SUBBYTES[8].a/w198 ), .B(
        \SUBBYTES[8].a/w199 ), .Z(n15860) );
  XOR \SUBBYTES[8].a/U3893  ( .A(n15862), .B(n15861), .Z(\SUBBYTES[8].a/w224 )
         );
  XOR \SUBBYTES[8].a/U3892  ( .A(\w1[8][121] ), .B(n15863), .Z(n15861) );
  XOR \SUBBYTES[8].a/U3891  ( .A(\SUBBYTES[8].a/w199 ), .B(
        \SUBBYTES[8].a/w201 ), .Z(n15862) );
  XOR \SUBBYTES[8].a/U3890  ( .A(\SUBBYTES[8].a/w183 ), .B(
        \SUBBYTES[8].a/w184 ), .Z(n15863) );
  XOR \SUBBYTES[7].a/U5649  ( .A(\SUBBYTES[7].a/w3390 ), .B(
        \SUBBYTES[7].a/w3391 ), .Z(n14585) );
  XOR \SUBBYTES[7].a/U5648  ( .A(n14585), .B(n13544), .Z(n14584) );
  XOR \SUBBYTES[7].a/U5647  ( .A(\SUBBYTES[7].a/w3383 ), .B(
        \SUBBYTES[7].a/w3400 ), .Z(n13544) );
  XOR \SUBBYTES[7].a/U5645  ( .A(\SUBBYTES[7].a/w3382 ), .B(
        \SUBBYTES[7].a/w3397 ), .Z(n13545) );
  XOR \SUBBYTES[7].a/U5644  ( .A(n14585), .B(n13546), .Z(n14776) );
  XOR \SUBBYTES[7].a/U5643  ( .A(\SUBBYTES[7].a/w3397 ), .B(
        \SUBBYTES[7].a/w3398 ), .Z(n13546) );
  XOR \SUBBYTES[7].a/U5642  ( .A(\SUBBYTES[7].a/w3359 ), .B(n13547), .Z(n14587) );
  XOR \SUBBYTES[7].a/U5641  ( .A(\SUBBYTES[7].a/w3350 ), .B(
        \SUBBYTES[7].a/w3351 ), .Z(n13547) );
  XOR \SUBBYTES[7].a/U5639  ( .A(\SUBBYTES[7].a/w3361 ), .B(n14776), .Z(n13548) );
  XOR \SUBBYTES[7].a/U5638  ( .A(n13550), .B(n13549), .Z(n14588) );
  XOR \SUBBYTES[7].a/U5637  ( .A(n13552), .B(n13551), .Z(n13549) );
  XOR \SUBBYTES[7].a/U5636  ( .A(\SUBBYTES[7].a/w3397 ), .B(
        \SUBBYTES[7].a/w3398 ), .Z(n13550) );
  XOR \SUBBYTES[7].a/U5635  ( .A(\SUBBYTES[7].a/w3361 ), .B(
        \SUBBYTES[7].a/w3385 ), .Z(n13551) );
  XOR \SUBBYTES[7].a/U5634  ( .A(\SUBBYTES[7].a/w3350 ), .B(
        \SUBBYTES[7].a/w3359 ), .Z(n13552) );
  XOR \SUBBYTES[7].a/U5633  ( .A(\SUBBYTES[7].a/w3382 ), .B(n13553), .Z(n14586) );
  XOR \SUBBYTES[7].a/U5632  ( .A(\SUBBYTES[7].a/w3365 ), .B(
        \SUBBYTES[7].a/w3368 ), .Z(n13553) );
  XOR \SUBBYTES[7].a/U5630  ( .A(\SUBBYTES[7].a/w3353 ), .B(n14588), .Z(n13554) );
  XOR \SUBBYTES[7].a/U5628  ( .A(\SUBBYTES[7].a/w3385 ), .B(
        \SUBBYTES[7].a/w3398 ), .Z(n13555) );
  XOR \SUBBYTES[7].a/U5626  ( .A(n13559), .B(n13558), .Z(n13556) );
  XOR \SUBBYTES[7].a/U5625  ( .A(n13561), .B(n13560), .Z(n13557) );
  XOR \SUBBYTES[7].a/U5624  ( .A(\SUBBYTES[7].a/w3397 ), .B(
        \SUBBYTES[7].a/w3400 ), .Z(n13558) );
  XOR \SUBBYTES[7].a/U5623  ( .A(\SUBBYTES[7].a/w3390 ), .B(
        \SUBBYTES[7].a/w3393 ), .Z(n13559) );
  XOR \SUBBYTES[7].a/U5622  ( .A(\SUBBYTES[7].a/w3365 ), .B(
        \SUBBYTES[7].a/w3366 ), .Z(n13560) );
  XOR \SUBBYTES[7].a/U5621  ( .A(\SUBBYTES[7].a/w3350 ), .B(
        \SUBBYTES[7].a/w3353 ), .Z(n13561) );
  XOR \SUBBYTES[7].a/U5619  ( .A(n14585), .B(n13564), .Z(n13562) );
  XOR \SUBBYTES[7].a/U5618  ( .A(n14587), .B(n14586), .Z(n13563) );
  XOR \SUBBYTES[7].a/U5617  ( .A(\SUBBYTES[7].a/w3358 ), .B(
        \SUBBYTES[7].a/w3385 ), .Z(n13564) );
  XOR \SUBBYTES[7].a/U5615  ( .A(n14588), .B(n13567), .Z(n13565) );
  XOR \SUBBYTES[7].a/U5614  ( .A(\SUBBYTES[7].a/w3391 ), .B(
        \SUBBYTES[7].a/w3393 ), .Z(n13566) );
  XOR \SUBBYTES[7].a/U5613  ( .A(\SUBBYTES[7].a/w3351 ), .B(
        \SUBBYTES[7].a/w3383 ), .Z(n13567) );
  XOR \SUBBYTES[7].a/U5612  ( .A(\SUBBYTES[7].a/w3183 ), .B(
        \SUBBYTES[7].a/w3184 ), .Z(n14590) );
  XOR \SUBBYTES[7].a/U5611  ( .A(n14590), .B(n13568), .Z(n14589) );
  XOR \SUBBYTES[7].a/U5610  ( .A(\SUBBYTES[7].a/w3176 ), .B(
        \SUBBYTES[7].a/w3193 ), .Z(n13568) );
  XOR \SUBBYTES[7].a/U5608  ( .A(\SUBBYTES[7].a/w3175 ), .B(
        \SUBBYTES[7].a/w3190 ), .Z(n13569) );
  XOR \SUBBYTES[7].a/U5607  ( .A(n14590), .B(n13570), .Z(n14777) );
  XOR \SUBBYTES[7].a/U5606  ( .A(\SUBBYTES[7].a/w3190 ), .B(
        \SUBBYTES[7].a/w3191 ), .Z(n13570) );
  XOR \SUBBYTES[7].a/U5605  ( .A(\SUBBYTES[7].a/w3152 ), .B(n13571), .Z(n14592) );
  XOR \SUBBYTES[7].a/U5604  ( .A(\SUBBYTES[7].a/w3143 ), .B(
        \SUBBYTES[7].a/w3144 ), .Z(n13571) );
  XOR \SUBBYTES[7].a/U5602  ( .A(\SUBBYTES[7].a/w3154 ), .B(n14777), .Z(n13572) );
  XOR \SUBBYTES[7].a/U5601  ( .A(n13574), .B(n13573), .Z(n14593) );
  XOR \SUBBYTES[7].a/U5600  ( .A(n13576), .B(n13575), .Z(n13573) );
  XOR \SUBBYTES[7].a/U5599  ( .A(\SUBBYTES[7].a/w3190 ), .B(
        \SUBBYTES[7].a/w3191 ), .Z(n13574) );
  XOR \SUBBYTES[7].a/U5598  ( .A(\SUBBYTES[7].a/w3154 ), .B(
        \SUBBYTES[7].a/w3178 ), .Z(n13575) );
  XOR \SUBBYTES[7].a/U5597  ( .A(\SUBBYTES[7].a/w3143 ), .B(
        \SUBBYTES[7].a/w3152 ), .Z(n13576) );
  XOR \SUBBYTES[7].a/U5596  ( .A(\SUBBYTES[7].a/w3175 ), .B(n13577), .Z(n14591) );
  XOR \SUBBYTES[7].a/U5595  ( .A(\SUBBYTES[7].a/w3158 ), .B(
        \SUBBYTES[7].a/w3161 ), .Z(n13577) );
  XOR \SUBBYTES[7].a/U5593  ( .A(\SUBBYTES[7].a/w3146 ), .B(n14593), .Z(n13578) );
  XOR \SUBBYTES[7].a/U5591  ( .A(\SUBBYTES[7].a/w3178 ), .B(
        \SUBBYTES[7].a/w3191 ), .Z(n13579) );
  XOR \SUBBYTES[7].a/U5589  ( .A(n13583), .B(n13582), .Z(n13580) );
  XOR \SUBBYTES[7].a/U5588  ( .A(n13585), .B(n13584), .Z(n13581) );
  XOR \SUBBYTES[7].a/U5587  ( .A(\SUBBYTES[7].a/w3190 ), .B(
        \SUBBYTES[7].a/w3193 ), .Z(n13582) );
  XOR \SUBBYTES[7].a/U5586  ( .A(\SUBBYTES[7].a/w3183 ), .B(
        \SUBBYTES[7].a/w3186 ), .Z(n13583) );
  XOR \SUBBYTES[7].a/U5585  ( .A(\SUBBYTES[7].a/w3158 ), .B(
        \SUBBYTES[7].a/w3159 ), .Z(n13584) );
  XOR \SUBBYTES[7].a/U5584  ( .A(\SUBBYTES[7].a/w3143 ), .B(
        \SUBBYTES[7].a/w3146 ), .Z(n13585) );
  XOR \SUBBYTES[7].a/U5582  ( .A(n14590), .B(n13588), .Z(n13586) );
  XOR \SUBBYTES[7].a/U5581  ( .A(n14592), .B(n14591), .Z(n13587) );
  XOR \SUBBYTES[7].a/U5580  ( .A(\SUBBYTES[7].a/w3151 ), .B(
        \SUBBYTES[7].a/w3178 ), .Z(n13588) );
  XOR \SUBBYTES[7].a/U5578  ( .A(n14593), .B(n13591), .Z(n13589) );
  XOR \SUBBYTES[7].a/U5577  ( .A(\SUBBYTES[7].a/w3184 ), .B(
        \SUBBYTES[7].a/w3186 ), .Z(n13590) );
  XOR \SUBBYTES[7].a/U5576  ( .A(\SUBBYTES[7].a/w3144 ), .B(
        \SUBBYTES[7].a/w3176 ), .Z(n13591) );
  XOR \SUBBYTES[7].a/U5575  ( .A(\SUBBYTES[7].a/w2976 ), .B(
        \SUBBYTES[7].a/w2977 ), .Z(n14595) );
  XOR \SUBBYTES[7].a/U5574  ( .A(n14595), .B(n13592), .Z(n14594) );
  XOR \SUBBYTES[7].a/U5573  ( .A(\SUBBYTES[7].a/w2969 ), .B(
        \SUBBYTES[7].a/w2986 ), .Z(n13592) );
  XOR \SUBBYTES[7].a/U5571  ( .A(\SUBBYTES[7].a/w2968 ), .B(
        \SUBBYTES[7].a/w2983 ), .Z(n13593) );
  XOR \SUBBYTES[7].a/U5570  ( .A(n14595), .B(n13594), .Z(n14778) );
  XOR \SUBBYTES[7].a/U5569  ( .A(\SUBBYTES[7].a/w2983 ), .B(
        \SUBBYTES[7].a/w2984 ), .Z(n13594) );
  XOR \SUBBYTES[7].a/U5568  ( .A(\SUBBYTES[7].a/w2945 ), .B(n13595), .Z(n14597) );
  XOR \SUBBYTES[7].a/U5567  ( .A(\SUBBYTES[7].a/w2936 ), .B(
        \SUBBYTES[7].a/w2937 ), .Z(n13595) );
  XOR \SUBBYTES[7].a/U5565  ( .A(\SUBBYTES[7].a/w2947 ), .B(n14778), .Z(n13596) );
  XOR \SUBBYTES[7].a/U5564  ( .A(n13598), .B(n13597), .Z(n14598) );
  XOR \SUBBYTES[7].a/U5563  ( .A(n13600), .B(n13599), .Z(n13597) );
  XOR \SUBBYTES[7].a/U5562  ( .A(\SUBBYTES[7].a/w2983 ), .B(
        \SUBBYTES[7].a/w2984 ), .Z(n13598) );
  XOR \SUBBYTES[7].a/U5561  ( .A(\SUBBYTES[7].a/w2947 ), .B(
        \SUBBYTES[7].a/w2971 ), .Z(n13599) );
  XOR \SUBBYTES[7].a/U5560  ( .A(\SUBBYTES[7].a/w2936 ), .B(
        \SUBBYTES[7].a/w2945 ), .Z(n13600) );
  XOR \SUBBYTES[7].a/U5559  ( .A(\SUBBYTES[7].a/w2968 ), .B(n13601), .Z(n14596) );
  XOR \SUBBYTES[7].a/U5558  ( .A(\SUBBYTES[7].a/w2951 ), .B(
        \SUBBYTES[7].a/w2954 ), .Z(n13601) );
  XOR \SUBBYTES[7].a/U5556  ( .A(\SUBBYTES[7].a/w2939 ), .B(n14598), .Z(n13602) );
  XOR \SUBBYTES[7].a/U5554  ( .A(\SUBBYTES[7].a/w2971 ), .B(
        \SUBBYTES[7].a/w2984 ), .Z(n13603) );
  XOR \SUBBYTES[7].a/U5552  ( .A(n13607), .B(n13606), .Z(n13604) );
  XOR \SUBBYTES[7].a/U5551  ( .A(n13609), .B(n13608), .Z(n13605) );
  XOR \SUBBYTES[7].a/U5550  ( .A(\SUBBYTES[7].a/w2983 ), .B(
        \SUBBYTES[7].a/w2986 ), .Z(n13606) );
  XOR \SUBBYTES[7].a/U5549  ( .A(\SUBBYTES[7].a/w2976 ), .B(
        \SUBBYTES[7].a/w2979 ), .Z(n13607) );
  XOR \SUBBYTES[7].a/U5548  ( .A(\SUBBYTES[7].a/w2951 ), .B(
        \SUBBYTES[7].a/w2952 ), .Z(n13608) );
  XOR \SUBBYTES[7].a/U5547  ( .A(\SUBBYTES[7].a/w2936 ), .B(
        \SUBBYTES[7].a/w2939 ), .Z(n13609) );
  XOR \SUBBYTES[7].a/U5545  ( .A(n14595), .B(n13612), .Z(n13610) );
  XOR \SUBBYTES[7].a/U5544  ( .A(n14597), .B(n14596), .Z(n13611) );
  XOR \SUBBYTES[7].a/U5543  ( .A(\SUBBYTES[7].a/w2944 ), .B(
        \SUBBYTES[7].a/w2971 ), .Z(n13612) );
  XOR \SUBBYTES[7].a/U5541  ( .A(n14598), .B(n13615), .Z(n13613) );
  XOR \SUBBYTES[7].a/U5540  ( .A(\SUBBYTES[7].a/w2977 ), .B(
        \SUBBYTES[7].a/w2979 ), .Z(n13614) );
  XOR \SUBBYTES[7].a/U5539  ( .A(\SUBBYTES[7].a/w2937 ), .B(
        \SUBBYTES[7].a/w2969 ), .Z(n13615) );
  XOR \SUBBYTES[7].a/U5538  ( .A(\SUBBYTES[7].a/w2769 ), .B(
        \SUBBYTES[7].a/w2770 ), .Z(n14600) );
  XOR \SUBBYTES[7].a/U5537  ( .A(n14600), .B(n13616), .Z(n14599) );
  XOR \SUBBYTES[7].a/U5536  ( .A(\SUBBYTES[7].a/w2762 ), .B(
        \SUBBYTES[7].a/w2779 ), .Z(n13616) );
  XOR \SUBBYTES[7].a/U5534  ( .A(\SUBBYTES[7].a/w2761 ), .B(
        \SUBBYTES[7].a/w2776 ), .Z(n13617) );
  XOR \SUBBYTES[7].a/U5533  ( .A(n14600), .B(n13618), .Z(n14779) );
  XOR \SUBBYTES[7].a/U5532  ( .A(\SUBBYTES[7].a/w2776 ), .B(
        \SUBBYTES[7].a/w2777 ), .Z(n13618) );
  XOR \SUBBYTES[7].a/U5531  ( .A(\SUBBYTES[7].a/w2738 ), .B(n13619), .Z(n14602) );
  XOR \SUBBYTES[7].a/U5530  ( .A(\SUBBYTES[7].a/w2729 ), .B(
        \SUBBYTES[7].a/w2730 ), .Z(n13619) );
  XOR \SUBBYTES[7].a/U5528  ( .A(\SUBBYTES[7].a/w2740 ), .B(n14779), .Z(n13620) );
  XOR \SUBBYTES[7].a/U5527  ( .A(n13622), .B(n13621), .Z(n14603) );
  XOR \SUBBYTES[7].a/U5526  ( .A(n13624), .B(n13623), .Z(n13621) );
  XOR \SUBBYTES[7].a/U5525  ( .A(\SUBBYTES[7].a/w2776 ), .B(
        \SUBBYTES[7].a/w2777 ), .Z(n13622) );
  XOR \SUBBYTES[7].a/U5524  ( .A(\SUBBYTES[7].a/w2740 ), .B(
        \SUBBYTES[7].a/w2764 ), .Z(n13623) );
  XOR \SUBBYTES[7].a/U5523  ( .A(\SUBBYTES[7].a/w2729 ), .B(
        \SUBBYTES[7].a/w2738 ), .Z(n13624) );
  XOR \SUBBYTES[7].a/U5522  ( .A(\SUBBYTES[7].a/w2761 ), .B(n13625), .Z(n14601) );
  XOR \SUBBYTES[7].a/U5521  ( .A(\SUBBYTES[7].a/w2744 ), .B(
        \SUBBYTES[7].a/w2747 ), .Z(n13625) );
  XOR \SUBBYTES[7].a/U5519  ( .A(\SUBBYTES[7].a/w2732 ), .B(n14603), .Z(n13626) );
  XOR \SUBBYTES[7].a/U5517  ( .A(\SUBBYTES[7].a/w2764 ), .B(
        \SUBBYTES[7].a/w2777 ), .Z(n13627) );
  XOR \SUBBYTES[7].a/U5515  ( .A(n13631), .B(n13630), .Z(n13628) );
  XOR \SUBBYTES[7].a/U5514  ( .A(n13633), .B(n13632), .Z(n13629) );
  XOR \SUBBYTES[7].a/U5513  ( .A(\SUBBYTES[7].a/w2776 ), .B(
        \SUBBYTES[7].a/w2779 ), .Z(n13630) );
  XOR \SUBBYTES[7].a/U5512  ( .A(\SUBBYTES[7].a/w2769 ), .B(
        \SUBBYTES[7].a/w2772 ), .Z(n13631) );
  XOR \SUBBYTES[7].a/U5511  ( .A(\SUBBYTES[7].a/w2744 ), .B(
        \SUBBYTES[7].a/w2745 ), .Z(n13632) );
  XOR \SUBBYTES[7].a/U5510  ( .A(\SUBBYTES[7].a/w2729 ), .B(
        \SUBBYTES[7].a/w2732 ), .Z(n13633) );
  XOR \SUBBYTES[7].a/U5508  ( .A(n14600), .B(n13636), .Z(n13634) );
  XOR \SUBBYTES[7].a/U5507  ( .A(n14602), .B(n14601), .Z(n13635) );
  XOR \SUBBYTES[7].a/U5506  ( .A(\SUBBYTES[7].a/w2737 ), .B(
        \SUBBYTES[7].a/w2764 ), .Z(n13636) );
  XOR \SUBBYTES[7].a/U5504  ( .A(n14603), .B(n13639), .Z(n13637) );
  XOR \SUBBYTES[7].a/U5503  ( .A(\SUBBYTES[7].a/w2770 ), .B(
        \SUBBYTES[7].a/w2772 ), .Z(n13638) );
  XOR \SUBBYTES[7].a/U5502  ( .A(\SUBBYTES[7].a/w2730 ), .B(
        \SUBBYTES[7].a/w2762 ), .Z(n13639) );
  XOR \SUBBYTES[7].a/U5501  ( .A(\SUBBYTES[7].a/w2562 ), .B(
        \SUBBYTES[7].a/w2563 ), .Z(n14605) );
  XOR \SUBBYTES[7].a/U5500  ( .A(n14605), .B(n13640), .Z(n14604) );
  XOR \SUBBYTES[7].a/U5499  ( .A(\SUBBYTES[7].a/w2555 ), .B(
        \SUBBYTES[7].a/w2572 ), .Z(n13640) );
  XOR \SUBBYTES[7].a/U5497  ( .A(\SUBBYTES[7].a/w2554 ), .B(
        \SUBBYTES[7].a/w2569 ), .Z(n13641) );
  XOR \SUBBYTES[7].a/U5496  ( .A(n14605), .B(n13642), .Z(n14780) );
  XOR \SUBBYTES[7].a/U5495  ( .A(\SUBBYTES[7].a/w2569 ), .B(
        \SUBBYTES[7].a/w2570 ), .Z(n13642) );
  XOR \SUBBYTES[7].a/U5494  ( .A(\SUBBYTES[7].a/w2531 ), .B(n13643), .Z(n14607) );
  XOR \SUBBYTES[7].a/U5493  ( .A(\SUBBYTES[7].a/w2522 ), .B(
        \SUBBYTES[7].a/w2523 ), .Z(n13643) );
  XOR \SUBBYTES[7].a/U5491  ( .A(\SUBBYTES[7].a/w2533 ), .B(n14780), .Z(n13644) );
  XOR \SUBBYTES[7].a/U5490  ( .A(n13646), .B(n13645), .Z(n14608) );
  XOR \SUBBYTES[7].a/U5489  ( .A(n13648), .B(n13647), .Z(n13645) );
  XOR \SUBBYTES[7].a/U5488  ( .A(\SUBBYTES[7].a/w2569 ), .B(
        \SUBBYTES[7].a/w2570 ), .Z(n13646) );
  XOR \SUBBYTES[7].a/U5487  ( .A(\SUBBYTES[7].a/w2533 ), .B(
        \SUBBYTES[7].a/w2557 ), .Z(n13647) );
  XOR \SUBBYTES[7].a/U5486  ( .A(\SUBBYTES[7].a/w2522 ), .B(
        \SUBBYTES[7].a/w2531 ), .Z(n13648) );
  XOR \SUBBYTES[7].a/U5485  ( .A(\SUBBYTES[7].a/w2554 ), .B(n13649), .Z(n14606) );
  XOR \SUBBYTES[7].a/U5484  ( .A(\SUBBYTES[7].a/w2537 ), .B(
        \SUBBYTES[7].a/w2540 ), .Z(n13649) );
  XOR \SUBBYTES[7].a/U5482  ( .A(\SUBBYTES[7].a/w2525 ), .B(n14608), .Z(n13650) );
  XOR \SUBBYTES[7].a/U5480  ( .A(\SUBBYTES[7].a/w2557 ), .B(
        \SUBBYTES[7].a/w2570 ), .Z(n13651) );
  XOR \SUBBYTES[7].a/U5478  ( .A(n13655), .B(n13654), .Z(n13652) );
  XOR \SUBBYTES[7].a/U5477  ( .A(n13657), .B(n13656), .Z(n13653) );
  XOR \SUBBYTES[7].a/U5476  ( .A(\SUBBYTES[7].a/w2569 ), .B(
        \SUBBYTES[7].a/w2572 ), .Z(n13654) );
  XOR \SUBBYTES[7].a/U5475  ( .A(\SUBBYTES[7].a/w2562 ), .B(
        \SUBBYTES[7].a/w2565 ), .Z(n13655) );
  XOR \SUBBYTES[7].a/U5474  ( .A(\SUBBYTES[7].a/w2537 ), .B(
        \SUBBYTES[7].a/w2538 ), .Z(n13656) );
  XOR \SUBBYTES[7].a/U5473  ( .A(\SUBBYTES[7].a/w2522 ), .B(
        \SUBBYTES[7].a/w2525 ), .Z(n13657) );
  XOR \SUBBYTES[7].a/U5471  ( .A(n14605), .B(n13660), .Z(n13658) );
  XOR \SUBBYTES[7].a/U5470  ( .A(n14607), .B(n14606), .Z(n13659) );
  XOR \SUBBYTES[7].a/U5469  ( .A(\SUBBYTES[7].a/w2530 ), .B(
        \SUBBYTES[7].a/w2557 ), .Z(n13660) );
  XOR \SUBBYTES[7].a/U5467  ( .A(n14608), .B(n13663), .Z(n13661) );
  XOR \SUBBYTES[7].a/U5466  ( .A(\SUBBYTES[7].a/w2563 ), .B(
        \SUBBYTES[7].a/w2565 ), .Z(n13662) );
  XOR \SUBBYTES[7].a/U5465  ( .A(\SUBBYTES[7].a/w2523 ), .B(
        \SUBBYTES[7].a/w2555 ), .Z(n13663) );
  XOR \SUBBYTES[7].a/U5464  ( .A(\SUBBYTES[7].a/w2355 ), .B(
        \SUBBYTES[7].a/w2356 ), .Z(n14610) );
  XOR \SUBBYTES[7].a/U5463  ( .A(n14610), .B(n13664), .Z(n14609) );
  XOR \SUBBYTES[7].a/U5462  ( .A(\SUBBYTES[7].a/w2348 ), .B(
        \SUBBYTES[7].a/w2365 ), .Z(n13664) );
  XOR \SUBBYTES[7].a/U5460  ( .A(\SUBBYTES[7].a/w2347 ), .B(
        \SUBBYTES[7].a/w2362 ), .Z(n13665) );
  XOR \SUBBYTES[7].a/U5459  ( .A(n14610), .B(n13666), .Z(n14781) );
  XOR \SUBBYTES[7].a/U5458  ( .A(\SUBBYTES[7].a/w2362 ), .B(
        \SUBBYTES[7].a/w2363 ), .Z(n13666) );
  XOR \SUBBYTES[7].a/U5457  ( .A(\SUBBYTES[7].a/w2324 ), .B(n13667), .Z(n14612) );
  XOR \SUBBYTES[7].a/U5456  ( .A(\SUBBYTES[7].a/w2315 ), .B(
        \SUBBYTES[7].a/w2316 ), .Z(n13667) );
  XOR \SUBBYTES[7].a/U5454  ( .A(\SUBBYTES[7].a/w2326 ), .B(n14781), .Z(n13668) );
  XOR \SUBBYTES[7].a/U5453  ( .A(n13670), .B(n13669), .Z(n14613) );
  XOR \SUBBYTES[7].a/U5452  ( .A(n13672), .B(n13671), .Z(n13669) );
  XOR \SUBBYTES[7].a/U5451  ( .A(\SUBBYTES[7].a/w2362 ), .B(
        \SUBBYTES[7].a/w2363 ), .Z(n13670) );
  XOR \SUBBYTES[7].a/U5450  ( .A(\SUBBYTES[7].a/w2326 ), .B(
        \SUBBYTES[7].a/w2350 ), .Z(n13671) );
  XOR \SUBBYTES[7].a/U5449  ( .A(\SUBBYTES[7].a/w2315 ), .B(
        \SUBBYTES[7].a/w2324 ), .Z(n13672) );
  XOR \SUBBYTES[7].a/U5448  ( .A(\SUBBYTES[7].a/w2347 ), .B(n13673), .Z(n14611) );
  XOR \SUBBYTES[7].a/U5447  ( .A(\SUBBYTES[7].a/w2330 ), .B(
        \SUBBYTES[7].a/w2333 ), .Z(n13673) );
  XOR \SUBBYTES[7].a/U5445  ( .A(\SUBBYTES[7].a/w2318 ), .B(n14613), .Z(n13674) );
  XOR \SUBBYTES[7].a/U5443  ( .A(\SUBBYTES[7].a/w2350 ), .B(
        \SUBBYTES[7].a/w2363 ), .Z(n13675) );
  XOR \SUBBYTES[7].a/U5441  ( .A(n13679), .B(n13678), .Z(n13676) );
  XOR \SUBBYTES[7].a/U5440  ( .A(n13681), .B(n13680), .Z(n13677) );
  XOR \SUBBYTES[7].a/U5439  ( .A(\SUBBYTES[7].a/w2362 ), .B(
        \SUBBYTES[7].a/w2365 ), .Z(n13678) );
  XOR \SUBBYTES[7].a/U5438  ( .A(\SUBBYTES[7].a/w2355 ), .B(
        \SUBBYTES[7].a/w2358 ), .Z(n13679) );
  XOR \SUBBYTES[7].a/U5437  ( .A(\SUBBYTES[7].a/w2330 ), .B(
        \SUBBYTES[7].a/w2331 ), .Z(n13680) );
  XOR \SUBBYTES[7].a/U5436  ( .A(\SUBBYTES[7].a/w2315 ), .B(
        \SUBBYTES[7].a/w2318 ), .Z(n13681) );
  XOR \SUBBYTES[7].a/U5434  ( .A(n14610), .B(n13684), .Z(n13682) );
  XOR \SUBBYTES[7].a/U5433  ( .A(n14612), .B(n14611), .Z(n13683) );
  XOR \SUBBYTES[7].a/U5432  ( .A(\SUBBYTES[7].a/w2323 ), .B(
        \SUBBYTES[7].a/w2350 ), .Z(n13684) );
  XOR \SUBBYTES[7].a/U5430  ( .A(n14613), .B(n13687), .Z(n13685) );
  XOR \SUBBYTES[7].a/U5429  ( .A(\SUBBYTES[7].a/w2356 ), .B(
        \SUBBYTES[7].a/w2358 ), .Z(n13686) );
  XOR \SUBBYTES[7].a/U5428  ( .A(\SUBBYTES[7].a/w2316 ), .B(
        \SUBBYTES[7].a/w2348 ), .Z(n13687) );
  XOR \SUBBYTES[7].a/U5427  ( .A(\SUBBYTES[7].a/w2148 ), .B(
        \SUBBYTES[7].a/w2149 ), .Z(n14615) );
  XOR \SUBBYTES[7].a/U5426  ( .A(n14615), .B(n13688), .Z(n14614) );
  XOR \SUBBYTES[7].a/U5425  ( .A(\SUBBYTES[7].a/w2141 ), .B(
        \SUBBYTES[7].a/w2158 ), .Z(n13688) );
  XOR \SUBBYTES[7].a/U5423  ( .A(\SUBBYTES[7].a/w2140 ), .B(
        \SUBBYTES[7].a/w2155 ), .Z(n13689) );
  XOR \SUBBYTES[7].a/U5422  ( .A(n14615), .B(n13690), .Z(n14782) );
  XOR \SUBBYTES[7].a/U5421  ( .A(\SUBBYTES[7].a/w2155 ), .B(
        \SUBBYTES[7].a/w2156 ), .Z(n13690) );
  XOR \SUBBYTES[7].a/U5420  ( .A(\SUBBYTES[7].a/w2117 ), .B(n13691), .Z(n14617) );
  XOR \SUBBYTES[7].a/U5419  ( .A(\SUBBYTES[7].a/w2108 ), .B(
        \SUBBYTES[7].a/w2109 ), .Z(n13691) );
  XOR \SUBBYTES[7].a/U5417  ( .A(\SUBBYTES[7].a/w2119 ), .B(n14782), .Z(n13692) );
  XOR \SUBBYTES[7].a/U5416  ( .A(n13694), .B(n13693), .Z(n14618) );
  XOR \SUBBYTES[7].a/U5415  ( .A(n13696), .B(n13695), .Z(n13693) );
  XOR \SUBBYTES[7].a/U5414  ( .A(\SUBBYTES[7].a/w2155 ), .B(
        \SUBBYTES[7].a/w2156 ), .Z(n13694) );
  XOR \SUBBYTES[7].a/U5413  ( .A(\SUBBYTES[7].a/w2119 ), .B(
        \SUBBYTES[7].a/w2143 ), .Z(n13695) );
  XOR \SUBBYTES[7].a/U5412  ( .A(\SUBBYTES[7].a/w2108 ), .B(
        \SUBBYTES[7].a/w2117 ), .Z(n13696) );
  XOR \SUBBYTES[7].a/U5411  ( .A(\SUBBYTES[7].a/w2140 ), .B(n13697), .Z(n14616) );
  XOR \SUBBYTES[7].a/U5410  ( .A(\SUBBYTES[7].a/w2123 ), .B(
        \SUBBYTES[7].a/w2126 ), .Z(n13697) );
  XOR \SUBBYTES[7].a/U5408  ( .A(\SUBBYTES[7].a/w2111 ), .B(n14618), .Z(n13698) );
  XOR \SUBBYTES[7].a/U5406  ( .A(\SUBBYTES[7].a/w2143 ), .B(
        \SUBBYTES[7].a/w2156 ), .Z(n13699) );
  XOR \SUBBYTES[7].a/U5404  ( .A(n13703), .B(n13702), .Z(n13700) );
  XOR \SUBBYTES[7].a/U5403  ( .A(n13705), .B(n13704), .Z(n13701) );
  XOR \SUBBYTES[7].a/U5402  ( .A(\SUBBYTES[7].a/w2155 ), .B(
        \SUBBYTES[7].a/w2158 ), .Z(n13702) );
  XOR \SUBBYTES[7].a/U5401  ( .A(\SUBBYTES[7].a/w2148 ), .B(
        \SUBBYTES[7].a/w2151 ), .Z(n13703) );
  XOR \SUBBYTES[7].a/U5400  ( .A(\SUBBYTES[7].a/w2123 ), .B(
        \SUBBYTES[7].a/w2124 ), .Z(n13704) );
  XOR \SUBBYTES[7].a/U5399  ( .A(\SUBBYTES[7].a/w2108 ), .B(
        \SUBBYTES[7].a/w2111 ), .Z(n13705) );
  XOR \SUBBYTES[7].a/U5397  ( .A(n14615), .B(n13708), .Z(n13706) );
  XOR \SUBBYTES[7].a/U5396  ( .A(n14617), .B(n14616), .Z(n13707) );
  XOR \SUBBYTES[7].a/U5395  ( .A(\SUBBYTES[7].a/w2116 ), .B(
        \SUBBYTES[7].a/w2143 ), .Z(n13708) );
  XOR \SUBBYTES[7].a/U5393  ( .A(n14618), .B(n13711), .Z(n13709) );
  XOR \SUBBYTES[7].a/U5392  ( .A(\SUBBYTES[7].a/w2149 ), .B(
        \SUBBYTES[7].a/w2151 ), .Z(n13710) );
  XOR \SUBBYTES[7].a/U5391  ( .A(\SUBBYTES[7].a/w2109 ), .B(
        \SUBBYTES[7].a/w2141 ), .Z(n13711) );
  XOR \SUBBYTES[7].a/U5390  ( .A(\SUBBYTES[7].a/w1941 ), .B(
        \SUBBYTES[7].a/w1942 ), .Z(n14620) );
  XOR \SUBBYTES[7].a/U5389  ( .A(n14620), .B(n13712), .Z(n14619) );
  XOR \SUBBYTES[7].a/U5388  ( .A(\SUBBYTES[7].a/w1934 ), .B(
        \SUBBYTES[7].a/w1951 ), .Z(n13712) );
  XOR \SUBBYTES[7].a/U5386  ( .A(\SUBBYTES[7].a/w1933 ), .B(
        \SUBBYTES[7].a/w1948 ), .Z(n13713) );
  XOR \SUBBYTES[7].a/U5385  ( .A(n14620), .B(n13714), .Z(n14783) );
  XOR \SUBBYTES[7].a/U5384  ( .A(\SUBBYTES[7].a/w1948 ), .B(
        \SUBBYTES[7].a/w1949 ), .Z(n13714) );
  XOR \SUBBYTES[7].a/U5383  ( .A(\SUBBYTES[7].a/w1910 ), .B(n13715), .Z(n14622) );
  XOR \SUBBYTES[7].a/U5382  ( .A(\SUBBYTES[7].a/w1901 ), .B(
        \SUBBYTES[7].a/w1902 ), .Z(n13715) );
  XOR \SUBBYTES[7].a/U5380  ( .A(\SUBBYTES[7].a/w1912 ), .B(n14783), .Z(n13716) );
  XOR \SUBBYTES[7].a/U5379  ( .A(n13718), .B(n13717), .Z(n14623) );
  XOR \SUBBYTES[7].a/U5378  ( .A(n13720), .B(n13719), .Z(n13717) );
  XOR \SUBBYTES[7].a/U5377  ( .A(\SUBBYTES[7].a/w1948 ), .B(
        \SUBBYTES[7].a/w1949 ), .Z(n13718) );
  XOR \SUBBYTES[7].a/U5376  ( .A(\SUBBYTES[7].a/w1912 ), .B(
        \SUBBYTES[7].a/w1936 ), .Z(n13719) );
  XOR \SUBBYTES[7].a/U5375  ( .A(\SUBBYTES[7].a/w1901 ), .B(
        \SUBBYTES[7].a/w1910 ), .Z(n13720) );
  XOR \SUBBYTES[7].a/U5374  ( .A(\SUBBYTES[7].a/w1933 ), .B(n13721), .Z(n14621) );
  XOR \SUBBYTES[7].a/U5373  ( .A(\SUBBYTES[7].a/w1916 ), .B(
        \SUBBYTES[7].a/w1919 ), .Z(n13721) );
  XOR \SUBBYTES[7].a/U5371  ( .A(\SUBBYTES[7].a/w1904 ), .B(n14623), .Z(n13722) );
  XOR \SUBBYTES[7].a/U5369  ( .A(\SUBBYTES[7].a/w1936 ), .B(
        \SUBBYTES[7].a/w1949 ), .Z(n13723) );
  XOR \SUBBYTES[7].a/U5367  ( .A(n13727), .B(n13726), .Z(n13724) );
  XOR \SUBBYTES[7].a/U5366  ( .A(n13729), .B(n13728), .Z(n13725) );
  XOR \SUBBYTES[7].a/U5365  ( .A(\SUBBYTES[7].a/w1948 ), .B(
        \SUBBYTES[7].a/w1951 ), .Z(n13726) );
  XOR \SUBBYTES[7].a/U5364  ( .A(\SUBBYTES[7].a/w1941 ), .B(
        \SUBBYTES[7].a/w1944 ), .Z(n13727) );
  XOR \SUBBYTES[7].a/U5363  ( .A(\SUBBYTES[7].a/w1916 ), .B(
        \SUBBYTES[7].a/w1917 ), .Z(n13728) );
  XOR \SUBBYTES[7].a/U5362  ( .A(\SUBBYTES[7].a/w1901 ), .B(
        \SUBBYTES[7].a/w1904 ), .Z(n13729) );
  XOR \SUBBYTES[7].a/U5360  ( .A(n14620), .B(n13732), .Z(n13730) );
  XOR \SUBBYTES[7].a/U5359  ( .A(n14622), .B(n14621), .Z(n13731) );
  XOR \SUBBYTES[7].a/U5358  ( .A(\SUBBYTES[7].a/w1909 ), .B(
        \SUBBYTES[7].a/w1936 ), .Z(n13732) );
  XOR \SUBBYTES[7].a/U5356  ( .A(n14623), .B(n13735), .Z(n13733) );
  XOR \SUBBYTES[7].a/U5355  ( .A(\SUBBYTES[7].a/w1942 ), .B(
        \SUBBYTES[7].a/w1944 ), .Z(n13734) );
  XOR \SUBBYTES[7].a/U5354  ( .A(\SUBBYTES[7].a/w1902 ), .B(
        \SUBBYTES[7].a/w1934 ), .Z(n13735) );
  XOR \SUBBYTES[7].a/U5353  ( .A(\SUBBYTES[7].a/w1734 ), .B(
        \SUBBYTES[7].a/w1735 ), .Z(n14625) );
  XOR \SUBBYTES[7].a/U5352  ( .A(n14625), .B(n13736), .Z(n14624) );
  XOR \SUBBYTES[7].a/U5351  ( .A(\SUBBYTES[7].a/w1727 ), .B(
        \SUBBYTES[7].a/w1744 ), .Z(n13736) );
  XOR \SUBBYTES[7].a/U5349  ( .A(\SUBBYTES[7].a/w1726 ), .B(
        \SUBBYTES[7].a/w1741 ), .Z(n13737) );
  XOR \SUBBYTES[7].a/U5348  ( .A(n14625), .B(n13738), .Z(n14784) );
  XOR \SUBBYTES[7].a/U5347  ( .A(\SUBBYTES[7].a/w1741 ), .B(
        \SUBBYTES[7].a/w1742 ), .Z(n13738) );
  XOR \SUBBYTES[7].a/U5346  ( .A(\SUBBYTES[7].a/w1703 ), .B(n13739), .Z(n14627) );
  XOR \SUBBYTES[7].a/U5345  ( .A(\SUBBYTES[7].a/w1694 ), .B(
        \SUBBYTES[7].a/w1695 ), .Z(n13739) );
  XOR \SUBBYTES[7].a/U5343  ( .A(\SUBBYTES[7].a/w1705 ), .B(n14784), .Z(n13740) );
  XOR \SUBBYTES[7].a/U5342  ( .A(n13742), .B(n13741), .Z(n14628) );
  XOR \SUBBYTES[7].a/U5341  ( .A(n13744), .B(n13743), .Z(n13741) );
  XOR \SUBBYTES[7].a/U5340  ( .A(\SUBBYTES[7].a/w1741 ), .B(
        \SUBBYTES[7].a/w1742 ), .Z(n13742) );
  XOR \SUBBYTES[7].a/U5339  ( .A(\SUBBYTES[7].a/w1705 ), .B(
        \SUBBYTES[7].a/w1729 ), .Z(n13743) );
  XOR \SUBBYTES[7].a/U5338  ( .A(\SUBBYTES[7].a/w1694 ), .B(
        \SUBBYTES[7].a/w1703 ), .Z(n13744) );
  XOR \SUBBYTES[7].a/U5337  ( .A(\SUBBYTES[7].a/w1726 ), .B(n13745), .Z(n14626) );
  XOR \SUBBYTES[7].a/U5336  ( .A(\SUBBYTES[7].a/w1709 ), .B(
        \SUBBYTES[7].a/w1712 ), .Z(n13745) );
  XOR \SUBBYTES[7].a/U5334  ( .A(\SUBBYTES[7].a/w1697 ), .B(n14628), .Z(n13746) );
  XOR \SUBBYTES[7].a/U5332  ( .A(\SUBBYTES[7].a/w1729 ), .B(
        \SUBBYTES[7].a/w1742 ), .Z(n13747) );
  XOR \SUBBYTES[7].a/U5330  ( .A(n13751), .B(n13750), .Z(n13748) );
  XOR \SUBBYTES[7].a/U5329  ( .A(n13753), .B(n13752), .Z(n13749) );
  XOR \SUBBYTES[7].a/U5328  ( .A(\SUBBYTES[7].a/w1741 ), .B(
        \SUBBYTES[7].a/w1744 ), .Z(n13750) );
  XOR \SUBBYTES[7].a/U5327  ( .A(\SUBBYTES[7].a/w1734 ), .B(
        \SUBBYTES[7].a/w1737 ), .Z(n13751) );
  XOR \SUBBYTES[7].a/U5326  ( .A(\SUBBYTES[7].a/w1709 ), .B(
        \SUBBYTES[7].a/w1710 ), .Z(n13752) );
  XOR \SUBBYTES[7].a/U5325  ( .A(\SUBBYTES[7].a/w1694 ), .B(
        \SUBBYTES[7].a/w1697 ), .Z(n13753) );
  XOR \SUBBYTES[7].a/U5323  ( .A(n14625), .B(n13756), .Z(n13754) );
  XOR \SUBBYTES[7].a/U5322  ( .A(n14627), .B(n14626), .Z(n13755) );
  XOR \SUBBYTES[7].a/U5321  ( .A(\SUBBYTES[7].a/w1702 ), .B(
        \SUBBYTES[7].a/w1729 ), .Z(n13756) );
  XOR \SUBBYTES[7].a/U5319  ( .A(n14628), .B(n13759), .Z(n13757) );
  XOR \SUBBYTES[7].a/U5318  ( .A(\SUBBYTES[7].a/w1735 ), .B(
        \SUBBYTES[7].a/w1737 ), .Z(n13758) );
  XOR \SUBBYTES[7].a/U5317  ( .A(\SUBBYTES[7].a/w1695 ), .B(
        \SUBBYTES[7].a/w1727 ), .Z(n13759) );
  XOR \SUBBYTES[7].a/U5316  ( .A(\SUBBYTES[7].a/w1527 ), .B(
        \SUBBYTES[7].a/w1528 ), .Z(n14630) );
  XOR \SUBBYTES[7].a/U5315  ( .A(n14630), .B(n13760), .Z(n14629) );
  XOR \SUBBYTES[7].a/U5314  ( .A(\SUBBYTES[7].a/w1520 ), .B(
        \SUBBYTES[7].a/w1537 ), .Z(n13760) );
  XOR \SUBBYTES[7].a/U5312  ( .A(\SUBBYTES[7].a/w1519 ), .B(
        \SUBBYTES[7].a/w1534 ), .Z(n13761) );
  XOR \SUBBYTES[7].a/U5311  ( .A(n14630), .B(n13762), .Z(n14785) );
  XOR \SUBBYTES[7].a/U5310  ( .A(\SUBBYTES[7].a/w1534 ), .B(
        \SUBBYTES[7].a/w1535 ), .Z(n13762) );
  XOR \SUBBYTES[7].a/U5309  ( .A(\SUBBYTES[7].a/w1496 ), .B(n13763), .Z(n14632) );
  XOR \SUBBYTES[7].a/U5308  ( .A(\SUBBYTES[7].a/w1487 ), .B(
        \SUBBYTES[7].a/w1488 ), .Z(n13763) );
  XOR \SUBBYTES[7].a/U5306  ( .A(\SUBBYTES[7].a/w1498 ), .B(n14785), .Z(n13764) );
  XOR \SUBBYTES[7].a/U5305  ( .A(n13766), .B(n13765), .Z(n14633) );
  XOR \SUBBYTES[7].a/U5304  ( .A(n13768), .B(n13767), .Z(n13765) );
  XOR \SUBBYTES[7].a/U5303  ( .A(\SUBBYTES[7].a/w1534 ), .B(
        \SUBBYTES[7].a/w1535 ), .Z(n13766) );
  XOR \SUBBYTES[7].a/U5302  ( .A(\SUBBYTES[7].a/w1498 ), .B(
        \SUBBYTES[7].a/w1522 ), .Z(n13767) );
  XOR \SUBBYTES[7].a/U5301  ( .A(\SUBBYTES[7].a/w1487 ), .B(
        \SUBBYTES[7].a/w1496 ), .Z(n13768) );
  XOR \SUBBYTES[7].a/U5300  ( .A(\SUBBYTES[7].a/w1519 ), .B(n13769), .Z(n14631) );
  XOR \SUBBYTES[7].a/U5299  ( .A(\SUBBYTES[7].a/w1502 ), .B(
        \SUBBYTES[7].a/w1505 ), .Z(n13769) );
  XOR \SUBBYTES[7].a/U5297  ( .A(\SUBBYTES[7].a/w1490 ), .B(n14633), .Z(n13770) );
  XOR \SUBBYTES[7].a/U5295  ( .A(\SUBBYTES[7].a/w1522 ), .B(
        \SUBBYTES[7].a/w1535 ), .Z(n13771) );
  XOR \SUBBYTES[7].a/U5293  ( .A(n13775), .B(n13774), .Z(n13772) );
  XOR \SUBBYTES[7].a/U5292  ( .A(n13777), .B(n13776), .Z(n13773) );
  XOR \SUBBYTES[7].a/U5291  ( .A(\SUBBYTES[7].a/w1534 ), .B(
        \SUBBYTES[7].a/w1537 ), .Z(n13774) );
  XOR \SUBBYTES[7].a/U5290  ( .A(\SUBBYTES[7].a/w1527 ), .B(
        \SUBBYTES[7].a/w1530 ), .Z(n13775) );
  XOR \SUBBYTES[7].a/U5289  ( .A(\SUBBYTES[7].a/w1502 ), .B(
        \SUBBYTES[7].a/w1503 ), .Z(n13776) );
  XOR \SUBBYTES[7].a/U5288  ( .A(\SUBBYTES[7].a/w1487 ), .B(
        \SUBBYTES[7].a/w1490 ), .Z(n13777) );
  XOR \SUBBYTES[7].a/U5286  ( .A(n14630), .B(n13780), .Z(n13778) );
  XOR \SUBBYTES[7].a/U5285  ( .A(n14632), .B(n14631), .Z(n13779) );
  XOR \SUBBYTES[7].a/U5284  ( .A(\SUBBYTES[7].a/w1495 ), .B(
        \SUBBYTES[7].a/w1522 ), .Z(n13780) );
  XOR \SUBBYTES[7].a/U5282  ( .A(n14633), .B(n13783), .Z(n13781) );
  XOR \SUBBYTES[7].a/U5281  ( .A(\SUBBYTES[7].a/w1528 ), .B(
        \SUBBYTES[7].a/w1530 ), .Z(n13782) );
  XOR \SUBBYTES[7].a/U5280  ( .A(\SUBBYTES[7].a/w1488 ), .B(
        \SUBBYTES[7].a/w1520 ), .Z(n13783) );
  XOR \SUBBYTES[7].a/U5279  ( .A(\SUBBYTES[7].a/w1320 ), .B(
        \SUBBYTES[7].a/w1321 ), .Z(n14635) );
  XOR \SUBBYTES[7].a/U5278  ( .A(n14635), .B(n13784), .Z(n14634) );
  XOR \SUBBYTES[7].a/U5277  ( .A(\SUBBYTES[7].a/w1313 ), .B(
        \SUBBYTES[7].a/w1330 ), .Z(n13784) );
  XOR \SUBBYTES[7].a/U5275  ( .A(\SUBBYTES[7].a/w1312 ), .B(
        \SUBBYTES[7].a/w1327 ), .Z(n13785) );
  XOR \SUBBYTES[7].a/U5274  ( .A(n14635), .B(n13786), .Z(n14786) );
  XOR \SUBBYTES[7].a/U5273  ( .A(\SUBBYTES[7].a/w1327 ), .B(
        \SUBBYTES[7].a/w1328 ), .Z(n13786) );
  XOR \SUBBYTES[7].a/U5272  ( .A(\SUBBYTES[7].a/w1289 ), .B(n13787), .Z(n14637) );
  XOR \SUBBYTES[7].a/U5271  ( .A(\SUBBYTES[7].a/w1280 ), .B(
        \SUBBYTES[7].a/w1281 ), .Z(n13787) );
  XOR \SUBBYTES[7].a/U5269  ( .A(\SUBBYTES[7].a/w1291 ), .B(n14786), .Z(n13788) );
  XOR \SUBBYTES[7].a/U5268  ( .A(n13790), .B(n13789), .Z(n14638) );
  XOR \SUBBYTES[7].a/U5267  ( .A(n13792), .B(n13791), .Z(n13789) );
  XOR \SUBBYTES[7].a/U5266  ( .A(\SUBBYTES[7].a/w1327 ), .B(
        \SUBBYTES[7].a/w1328 ), .Z(n13790) );
  XOR \SUBBYTES[7].a/U5265  ( .A(\SUBBYTES[7].a/w1291 ), .B(
        \SUBBYTES[7].a/w1315 ), .Z(n13791) );
  XOR \SUBBYTES[7].a/U5264  ( .A(\SUBBYTES[7].a/w1280 ), .B(
        \SUBBYTES[7].a/w1289 ), .Z(n13792) );
  XOR \SUBBYTES[7].a/U5263  ( .A(\SUBBYTES[7].a/w1312 ), .B(n13793), .Z(n14636) );
  XOR \SUBBYTES[7].a/U5262  ( .A(\SUBBYTES[7].a/w1295 ), .B(
        \SUBBYTES[7].a/w1298 ), .Z(n13793) );
  XOR \SUBBYTES[7].a/U5260  ( .A(\SUBBYTES[7].a/w1283 ), .B(n14638), .Z(n13794) );
  XOR \SUBBYTES[7].a/U5258  ( .A(\SUBBYTES[7].a/w1315 ), .B(
        \SUBBYTES[7].a/w1328 ), .Z(n13795) );
  XOR \SUBBYTES[7].a/U5256  ( .A(n13799), .B(n13798), .Z(n13796) );
  XOR \SUBBYTES[7].a/U5255  ( .A(n13801), .B(n13800), .Z(n13797) );
  XOR \SUBBYTES[7].a/U5254  ( .A(\SUBBYTES[7].a/w1327 ), .B(
        \SUBBYTES[7].a/w1330 ), .Z(n13798) );
  XOR \SUBBYTES[7].a/U5253  ( .A(\SUBBYTES[7].a/w1320 ), .B(
        \SUBBYTES[7].a/w1323 ), .Z(n13799) );
  XOR \SUBBYTES[7].a/U5252  ( .A(\SUBBYTES[7].a/w1295 ), .B(
        \SUBBYTES[7].a/w1296 ), .Z(n13800) );
  XOR \SUBBYTES[7].a/U5251  ( .A(\SUBBYTES[7].a/w1280 ), .B(
        \SUBBYTES[7].a/w1283 ), .Z(n13801) );
  XOR \SUBBYTES[7].a/U5249  ( .A(n14635), .B(n13804), .Z(n13802) );
  XOR \SUBBYTES[7].a/U5248  ( .A(n14637), .B(n14636), .Z(n13803) );
  XOR \SUBBYTES[7].a/U5247  ( .A(\SUBBYTES[7].a/w1288 ), .B(
        \SUBBYTES[7].a/w1315 ), .Z(n13804) );
  XOR \SUBBYTES[7].a/U5245  ( .A(n14638), .B(n13807), .Z(n13805) );
  XOR \SUBBYTES[7].a/U5244  ( .A(\SUBBYTES[7].a/w1321 ), .B(
        \SUBBYTES[7].a/w1323 ), .Z(n13806) );
  XOR \SUBBYTES[7].a/U5243  ( .A(\SUBBYTES[7].a/w1281 ), .B(
        \SUBBYTES[7].a/w1313 ), .Z(n13807) );
  XOR \SUBBYTES[7].a/U5242  ( .A(\SUBBYTES[7].a/w1113 ), .B(
        \SUBBYTES[7].a/w1114 ), .Z(n14640) );
  XOR \SUBBYTES[7].a/U5241  ( .A(n14640), .B(n13808), .Z(n14639) );
  XOR \SUBBYTES[7].a/U5240  ( .A(\SUBBYTES[7].a/w1106 ), .B(
        \SUBBYTES[7].a/w1123 ), .Z(n13808) );
  XOR \SUBBYTES[7].a/U5238  ( .A(\SUBBYTES[7].a/w1105 ), .B(
        \SUBBYTES[7].a/w1120 ), .Z(n13809) );
  XOR \SUBBYTES[7].a/U5237  ( .A(n14640), .B(n13810), .Z(n14787) );
  XOR \SUBBYTES[7].a/U5236  ( .A(\SUBBYTES[7].a/w1120 ), .B(
        \SUBBYTES[7].a/w1121 ), .Z(n13810) );
  XOR \SUBBYTES[7].a/U5235  ( .A(\SUBBYTES[7].a/w1082 ), .B(n13811), .Z(n14642) );
  XOR \SUBBYTES[7].a/U5234  ( .A(\SUBBYTES[7].a/w1073 ), .B(
        \SUBBYTES[7].a/w1074 ), .Z(n13811) );
  XOR \SUBBYTES[7].a/U5232  ( .A(\SUBBYTES[7].a/w1084 ), .B(n14787), .Z(n13812) );
  XOR \SUBBYTES[7].a/U5231  ( .A(n13814), .B(n13813), .Z(n14643) );
  XOR \SUBBYTES[7].a/U5230  ( .A(n13816), .B(n13815), .Z(n13813) );
  XOR \SUBBYTES[7].a/U5229  ( .A(\SUBBYTES[7].a/w1120 ), .B(
        \SUBBYTES[7].a/w1121 ), .Z(n13814) );
  XOR \SUBBYTES[7].a/U5228  ( .A(\SUBBYTES[7].a/w1084 ), .B(
        \SUBBYTES[7].a/w1108 ), .Z(n13815) );
  XOR \SUBBYTES[7].a/U5227  ( .A(\SUBBYTES[7].a/w1073 ), .B(
        \SUBBYTES[7].a/w1082 ), .Z(n13816) );
  XOR \SUBBYTES[7].a/U5226  ( .A(\SUBBYTES[7].a/w1105 ), .B(n13817), .Z(n14641) );
  XOR \SUBBYTES[7].a/U5225  ( .A(\SUBBYTES[7].a/w1088 ), .B(
        \SUBBYTES[7].a/w1091 ), .Z(n13817) );
  XOR \SUBBYTES[7].a/U5223  ( .A(\SUBBYTES[7].a/w1076 ), .B(n14643), .Z(n13818) );
  XOR \SUBBYTES[7].a/U5221  ( .A(\SUBBYTES[7].a/w1108 ), .B(
        \SUBBYTES[7].a/w1121 ), .Z(n13819) );
  XOR \SUBBYTES[7].a/U5219  ( .A(n13823), .B(n13822), .Z(n13820) );
  XOR \SUBBYTES[7].a/U5218  ( .A(n13825), .B(n13824), .Z(n13821) );
  XOR \SUBBYTES[7].a/U5217  ( .A(\SUBBYTES[7].a/w1120 ), .B(
        \SUBBYTES[7].a/w1123 ), .Z(n13822) );
  XOR \SUBBYTES[7].a/U5216  ( .A(\SUBBYTES[7].a/w1113 ), .B(
        \SUBBYTES[7].a/w1116 ), .Z(n13823) );
  XOR \SUBBYTES[7].a/U5215  ( .A(\SUBBYTES[7].a/w1088 ), .B(
        \SUBBYTES[7].a/w1089 ), .Z(n13824) );
  XOR \SUBBYTES[7].a/U5214  ( .A(\SUBBYTES[7].a/w1073 ), .B(
        \SUBBYTES[7].a/w1076 ), .Z(n13825) );
  XOR \SUBBYTES[7].a/U5212  ( .A(n14640), .B(n13828), .Z(n13826) );
  XOR \SUBBYTES[7].a/U5211  ( .A(n14642), .B(n14641), .Z(n13827) );
  XOR \SUBBYTES[7].a/U5210  ( .A(\SUBBYTES[7].a/w1081 ), .B(
        \SUBBYTES[7].a/w1108 ), .Z(n13828) );
  XOR \SUBBYTES[7].a/U5208  ( .A(n14643), .B(n13831), .Z(n13829) );
  XOR \SUBBYTES[7].a/U5207  ( .A(\SUBBYTES[7].a/w1114 ), .B(
        \SUBBYTES[7].a/w1116 ), .Z(n13830) );
  XOR \SUBBYTES[7].a/U5206  ( .A(\SUBBYTES[7].a/w1074 ), .B(
        \SUBBYTES[7].a/w1106 ), .Z(n13831) );
  XOR \SUBBYTES[7].a/U5205  ( .A(\SUBBYTES[7].a/w906 ), .B(
        \SUBBYTES[7].a/w907 ), .Z(n14645) );
  XOR \SUBBYTES[7].a/U5204  ( .A(n14645), .B(n13832), .Z(n14644) );
  XOR \SUBBYTES[7].a/U5203  ( .A(\SUBBYTES[7].a/w899 ), .B(
        \SUBBYTES[7].a/w916 ), .Z(n13832) );
  XOR \SUBBYTES[7].a/U5201  ( .A(\SUBBYTES[7].a/w898 ), .B(
        \SUBBYTES[7].a/w913 ), .Z(n13833) );
  XOR \SUBBYTES[7].a/U5200  ( .A(n14645), .B(n13834), .Z(n14788) );
  XOR \SUBBYTES[7].a/U5199  ( .A(\SUBBYTES[7].a/w913 ), .B(
        \SUBBYTES[7].a/w914 ), .Z(n13834) );
  XOR \SUBBYTES[7].a/U5198  ( .A(\SUBBYTES[7].a/w875 ), .B(n13835), .Z(n14647)
         );
  XOR \SUBBYTES[7].a/U5197  ( .A(\SUBBYTES[7].a/w866 ), .B(
        \SUBBYTES[7].a/w867 ), .Z(n13835) );
  XOR \SUBBYTES[7].a/U5195  ( .A(\SUBBYTES[7].a/w877 ), .B(n14788), .Z(n13836)
         );
  XOR \SUBBYTES[7].a/U5194  ( .A(n13838), .B(n13837), .Z(n14648) );
  XOR \SUBBYTES[7].a/U5193  ( .A(n13840), .B(n13839), .Z(n13837) );
  XOR \SUBBYTES[7].a/U5192  ( .A(\SUBBYTES[7].a/w913 ), .B(
        \SUBBYTES[7].a/w914 ), .Z(n13838) );
  XOR \SUBBYTES[7].a/U5191  ( .A(\SUBBYTES[7].a/w877 ), .B(
        \SUBBYTES[7].a/w901 ), .Z(n13839) );
  XOR \SUBBYTES[7].a/U5190  ( .A(\SUBBYTES[7].a/w866 ), .B(
        \SUBBYTES[7].a/w875 ), .Z(n13840) );
  XOR \SUBBYTES[7].a/U5189  ( .A(\SUBBYTES[7].a/w898 ), .B(n13841), .Z(n14646)
         );
  XOR \SUBBYTES[7].a/U5188  ( .A(\SUBBYTES[7].a/w881 ), .B(
        \SUBBYTES[7].a/w884 ), .Z(n13841) );
  XOR \SUBBYTES[7].a/U5186  ( .A(\SUBBYTES[7].a/w869 ), .B(n14648), .Z(n13842)
         );
  XOR \SUBBYTES[7].a/U5184  ( .A(\SUBBYTES[7].a/w901 ), .B(
        \SUBBYTES[7].a/w914 ), .Z(n13843) );
  XOR \SUBBYTES[7].a/U5182  ( .A(n13847), .B(n13846), .Z(n13844) );
  XOR \SUBBYTES[7].a/U5181  ( .A(n13849), .B(n13848), .Z(n13845) );
  XOR \SUBBYTES[7].a/U5180  ( .A(\SUBBYTES[7].a/w913 ), .B(
        \SUBBYTES[7].a/w916 ), .Z(n13846) );
  XOR \SUBBYTES[7].a/U5179  ( .A(\SUBBYTES[7].a/w906 ), .B(
        \SUBBYTES[7].a/w909 ), .Z(n13847) );
  XOR \SUBBYTES[7].a/U5178  ( .A(\SUBBYTES[7].a/w881 ), .B(
        \SUBBYTES[7].a/w882 ), .Z(n13848) );
  XOR \SUBBYTES[7].a/U5177  ( .A(\SUBBYTES[7].a/w866 ), .B(
        \SUBBYTES[7].a/w869 ), .Z(n13849) );
  XOR \SUBBYTES[7].a/U5175  ( .A(n14645), .B(n13852), .Z(n13850) );
  XOR \SUBBYTES[7].a/U5174  ( .A(n14647), .B(n14646), .Z(n13851) );
  XOR \SUBBYTES[7].a/U5173  ( .A(\SUBBYTES[7].a/w874 ), .B(
        \SUBBYTES[7].a/w901 ), .Z(n13852) );
  XOR \SUBBYTES[7].a/U5171  ( .A(n14648), .B(n13855), .Z(n13853) );
  XOR \SUBBYTES[7].a/U5170  ( .A(\SUBBYTES[7].a/w907 ), .B(
        \SUBBYTES[7].a/w909 ), .Z(n13854) );
  XOR \SUBBYTES[7].a/U5169  ( .A(\SUBBYTES[7].a/w867 ), .B(
        \SUBBYTES[7].a/w899 ), .Z(n13855) );
  XOR \SUBBYTES[7].a/U5168  ( .A(\SUBBYTES[7].a/w699 ), .B(
        \SUBBYTES[7].a/w700 ), .Z(n14650) );
  XOR \SUBBYTES[7].a/U5167  ( .A(n14650), .B(n13856), .Z(n14649) );
  XOR \SUBBYTES[7].a/U5166  ( .A(\SUBBYTES[7].a/w692 ), .B(
        \SUBBYTES[7].a/w709 ), .Z(n13856) );
  XOR \SUBBYTES[7].a/U5164  ( .A(\SUBBYTES[7].a/w691 ), .B(
        \SUBBYTES[7].a/w706 ), .Z(n13857) );
  XOR \SUBBYTES[7].a/U5163  ( .A(n14650), .B(n13858), .Z(n14789) );
  XOR \SUBBYTES[7].a/U5162  ( .A(\SUBBYTES[7].a/w706 ), .B(
        \SUBBYTES[7].a/w707 ), .Z(n13858) );
  XOR \SUBBYTES[7].a/U5161  ( .A(\SUBBYTES[7].a/w668 ), .B(n13859), .Z(n14652)
         );
  XOR \SUBBYTES[7].a/U5160  ( .A(\SUBBYTES[7].a/w659 ), .B(
        \SUBBYTES[7].a/w660 ), .Z(n13859) );
  XOR \SUBBYTES[7].a/U5158  ( .A(\SUBBYTES[7].a/w670 ), .B(n14789), .Z(n13860)
         );
  XOR \SUBBYTES[7].a/U5157  ( .A(n13862), .B(n13861), .Z(n14653) );
  XOR \SUBBYTES[7].a/U5156  ( .A(n13864), .B(n13863), .Z(n13861) );
  XOR \SUBBYTES[7].a/U5155  ( .A(\SUBBYTES[7].a/w706 ), .B(
        \SUBBYTES[7].a/w707 ), .Z(n13862) );
  XOR \SUBBYTES[7].a/U5154  ( .A(\SUBBYTES[7].a/w670 ), .B(
        \SUBBYTES[7].a/w694 ), .Z(n13863) );
  XOR \SUBBYTES[7].a/U5153  ( .A(\SUBBYTES[7].a/w659 ), .B(
        \SUBBYTES[7].a/w668 ), .Z(n13864) );
  XOR \SUBBYTES[7].a/U5152  ( .A(\SUBBYTES[7].a/w691 ), .B(n13865), .Z(n14651)
         );
  XOR \SUBBYTES[7].a/U5151  ( .A(\SUBBYTES[7].a/w674 ), .B(
        \SUBBYTES[7].a/w677 ), .Z(n13865) );
  XOR \SUBBYTES[7].a/U5149  ( .A(\SUBBYTES[7].a/w662 ), .B(n14653), .Z(n13866)
         );
  XOR \SUBBYTES[7].a/U5147  ( .A(\SUBBYTES[7].a/w694 ), .B(
        \SUBBYTES[7].a/w707 ), .Z(n13867) );
  XOR \SUBBYTES[7].a/U5145  ( .A(n13871), .B(n13870), .Z(n13868) );
  XOR \SUBBYTES[7].a/U5144  ( .A(n13873), .B(n13872), .Z(n13869) );
  XOR \SUBBYTES[7].a/U5143  ( .A(\SUBBYTES[7].a/w706 ), .B(
        \SUBBYTES[7].a/w709 ), .Z(n13870) );
  XOR \SUBBYTES[7].a/U5142  ( .A(\SUBBYTES[7].a/w699 ), .B(
        \SUBBYTES[7].a/w702 ), .Z(n13871) );
  XOR \SUBBYTES[7].a/U5141  ( .A(\SUBBYTES[7].a/w674 ), .B(
        \SUBBYTES[7].a/w675 ), .Z(n13872) );
  XOR \SUBBYTES[7].a/U5140  ( .A(\SUBBYTES[7].a/w659 ), .B(
        \SUBBYTES[7].a/w662 ), .Z(n13873) );
  XOR \SUBBYTES[7].a/U5138  ( .A(n14650), .B(n13876), .Z(n13874) );
  XOR \SUBBYTES[7].a/U5137  ( .A(n14652), .B(n14651), .Z(n13875) );
  XOR \SUBBYTES[7].a/U5136  ( .A(\SUBBYTES[7].a/w667 ), .B(
        \SUBBYTES[7].a/w694 ), .Z(n13876) );
  XOR \SUBBYTES[7].a/U5134  ( .A(n14653), .B(n13879), .Z(n13877) );
  XOR \SUBBYTES[7].a/U5133  ( .A(\SUBBYTES[7].a/w700 ), .B(
        \SUBBYTES[7].a/w702 ), .Z(n13878) );
  XOR \SUBBYTES[7].a/U5132  ( .A(\SUBBYTES[7].a/w660 ), .B(
        \SUBBYTES[7].a/w692 ), .Z(n13879) );
  XOR \SUBBYTES[7].a/U5131  ( .A(\SUBBYTES[7].a/w492 ), .B(
        \SUBBYTES[7].a/w493 ), .Z(n14655) );
  XOR \SUBBYTES[7].a/U5130  ( .A(n14655), .B(n13880), .Z(n14654) );
  XOR \SUBBYTES[7].a/U5129  ( .A(\SUBBYTES[7].a/w485 ), .B(
        \SUBBYTES[7].a/w502 ), .Z(n13880) );
  XOR \SUBBYTES[7].a/U5127  ( .A(\SUBBYTES[7].a/w484 ), .B(
        \SUBBYTES[7].a/w499 ), .Z(n13881) );
  XOR \SUBBYTES[7].a/U5126  ( .A(n14655), .B(n13882), .Z(n14790) );
  XOR \SUBBYTES[7].a/U5125  ( .A(\SUBBYTES[7].a/w499 ), .B(
        \SUBBYTES[7].a/w500 ), .Z(n13882) );
  XOR \SUBBYTES[7].a/U5124  ( .A(\SUBBYTES[7].a/w461 ), .B(n13883), .Z(n14657)
         );
  XOR \SUBBYTES[7].a/U5123  ( .A(\SUBBYTES[7].a/w452 ), .B(
        \SUBBYTES[7].a/w453 ), .Z(n13883) );
  XOR \SUBBYTES[7].a/U5121  ( .A(\SUBBYTES[7].a/w463 ), .B(n14790), .Z(n13884)
         );
  XOR \SUBBYTES[7].a/U5120  ( .A(n13886), .B(n13885), .Z(n14658) );
  XOR \SUBBYTES[7].a/U5119  ( .A(n13888), .B(n13887), .Z(n13885) );
  XOR \SUBBYTES[7].a/U5118  ( .A(\SUBBYTES[7].a/w499 ), .B(
        \SUBBYTES[7].a/w500 ), .Z(n13886) );
  XOR \SUBBYTES[7].a/U5117  ( .A(\SUBBYTES[7].a/w463 ), .B(
        \SUBBYTES[7].a/w487 ), .Z(n13887) );
  XOR \SUBBYTES[7].a/U5116  ( .A(\SUBBYTES[7].a/w452 ), .B(
        \SUBBYTES[7].a/w461 ), .Z(n13888) );
  XOR \SUBBYTES[7].a/U5115  ( .A(\SUBBYTES[7].a/w484 ), .B(n13889), .Z(n14656)
         );
  XOR \SUBBYTES[7].a/U5114  ( .A(\SUBBYTES[7].a/w467 ), .B(
        \SUBBYTES[7].a/w470 ), .Z(n13889) );
  XOR \SUBBYTES[7].a/U5112  ( .A(\SUBBYTES[7].a/w455 ), .B(n14658), .Z(n13890)
         );
  XOR \SUBBYTES[7].a/U5110  ( .A(\SUBBYTES[7].a/w487 ), .B(
        \SUBBYTES[7].a/w500 ), .Z(n13891) );
  XOR \SUBBYTES[7].a/U5108  ( .A(n13895), .B(n13894), .Z(n13892) );
  XOR \SUBBYTES[7].a/U5107  ( .A(n13897), .B(n13896), .Z(n13893) );
  XOR \SUBBYTES[7].a/U5106  ( .A(\SUBBYTES[7].a/w499 ), .B(
        \SUBBYTES[7].a/w502 ), .Z(n13894) );
  XOR \SUBBYTES[7].a/U5105  ( .A(\SUBBYTES[7].a/w492 ), .B(
        \SUBBYTES[7].a/w495 ), .Z(n13895) );
  XOR \SUBBYTES[7].a/U5104  ( .A(\SUBBYTES[7].a/w467 ), .B(
        \SUBBYTES[7].a/w468 ), .Z(n13896) );
  XOR \SUBBYTES[7].a/U5103  ( .A(\SUBBYTES[7].a/w452 ), .B(
        \SUBBYTES[7].a/w455 ), .Z(n13897) );
  XOR \SUBBYTES[7].a/U5101  ( .A(n14655), .B(n13900), .Z(n13898) );
  XOR \SUBBYTES[7].a/U5100  ( .A(n14657), .B(n14656), .Z(n13899) );
  XOR \SUBBYTES[7].a/U5099  ( .A(\SUBBYTES[7].a/w460 ), .B(
        \SUBBYTES[7].a/w487 ), .Z(n13900) );
  XOR \SUBBYTES[7].a/U5097  ( .A(n14658), .B(n13903), .Z(n13901) );
  XOR \SUBBYTES[7].a/U5096  ( .A(\SUBBYTES[7].a/w493 ), .B(
        \SUBBYTES[7].a/w495 ), .Z(n13902) );
  XOR \SUBBYTES[7].a/U5095  ( .A(\SUBBYTES[7].a/w453 ), .B(
        \SUBBYTES[7].a/w485 ), .Z(n13903) );
  XOR \SUBBYTES[7].a/U5094  ( .A(\SUBBYTES[7].a/w285 ), .B(
        \SUBBYTES[7].a/w286 ), .Z(n14660) );
  XOR \SUBBYTES[7].a/U5093  ( .A(n14660), .B(n13904), .Z(n14659) );
  XOR \SUBBYTES[7].a/U5092  ( .A(\SUBBYTES[7].a/w278 ), .B(
        \SUBBYTES[7].a/w295 ), .Z(n13904) );
  XOR \SUBBYTES[7].a/U5090  ( .A(\SUBBYTES[7].a/w277 ), .B(
        \SUBBYTES[7].a/w292 ), .Z(n13905) );
  XOR \SUBBYTES[7].a/U5089  ( .A(n14660), .B(n13906), .Z(n14791) );
  XOR \SUBBYTES[7].a/U5088  ( .A(\SUBBYTES[7].a/w292 ), .B(
        \SUBBYTES[7].a/w293 ), .Z(n13906) );
  XOR \SUBBYTES[7].a/U5087  ( .A(\SUBBYTES[7].a/w254 ), .B(n13907), .Z(n14662)
         );
  XOR \SUBBYTES[7].a/U5086  ( .A(\SUBBYTES[7].a/w245 ), .B(
        \SUBBYTES[7].a/w246 ), .Z(n13907) );
  XOR \SUBBYTES[7].a/U5084  ( .A(\SUBBYTES[7].a/w256 ), .B(n14791), .Z(n13908)
         );
  XOR \SUBBYTES[7].a/U5083  ( .A(n13910), .B(n13909), .Z(n14663) );
  XOR \SUBBYTES[7].a/U5082  ( .A(n13912), .B(n13911), .Z(n13909) );
  XOR \SUBBYTES[7].a/U5081  ( .A(\SUBBYTES[7].a/w292 ), .B(
        \SUBBYTES[7].a/w293 ), .Z(n13910) );
  XOR \SUBBYTES[7].a/U5080  ( .A(\SUBBYTES[7].a/w256 ), .B(
        \SUBBYTES[7].a/w280 ), .Z(n13911) );
  XOR \SUBBYTES[7].a/U5079  ( .A(\SUBBYTES[7].a/w245 ), .B(
        \SUBBYTES[7].a/w254 ), .Z(n13912) );
  XOR \SUBBYTES[7].a/U5078  ( .A(\SUBBYTES[7].a/w277 ), .B(n13913), .Z(n14661)
         );
  XOR \SUBBYTES[7].a/U5077  ( .A(\SUBBYTES[7].a/w260 ), .B(
        \SUBBYTES[7].a/w263 ), .Z(n13913) );
  XOR \SUBBYTES[7].a/U5075  ( .A(\SUBBYTES[7].a/w248 ), .B(n14663), .Z(n13914)
         );
  XOR \SUBBYTES[7].a/U5073  ( .A(\SUBBYTES[7].a/w280 ), .B(
        \SUBBYTES[7].a/w293 ), .Z(n13915) );
  XOR \SUBBYTES[7].a/U5071  ( .A(n13919), .B(n13918), .Z(n13916) );
  XOR \SUBBYTES[7].a/U5070  ( .A(n13921), .B(n13920), .Z(n13917) );
  XOR \SUBBYTES[7].a/U5069  ( .A(\SUBBYTES[7].a/w292 ), .B(
        \SUBBYTES[7].a/w295 ), .Z(n13918) );
  XOR \SUBBYTES[7].a/U5068  ( .A(\SUBBYTES[7].a/w285 ), .B(
        \SUBBYTES[7].a/w288 ), .Z(n13919) );
  XOR \SUBBYTES[7].a/U5067  ( .A(\SUBBYTES[7].a/w260 ), .B(
        \SUBBYTES[7].a/w261 ), .Z(n13920) );
  XOR \SUBBYTES[7].a/U5066  ( .A(\SUBBYTES[7].a/w245 ), .B(
        \SUBBYTES[7].a/w248 ), .Z(n13921) );
  XOR \SUBBYTES[7].a/U5064  ( .A(n14660), .B(n13924), .Z(n13922) );
  XOR \SUBBYTES[7].a/U5063  ( .A(n14662), .B(n14661), .Z(n13923) );
  XOR \SUBBYTES[7].a/U5062  ( .A(\SUBBYTES[7].a/w253 ), .B(
        \SUBBYTES[7].a/w280 ), .Z(n13924) );
  XOR \SUBBYTES[7].a/U5060  ( .A(n14663), .B(n13927), .Z(n13925) );
  XOR \SUBBYTES[7].a/U5059  ( .A(\SUBBYTES[7].a/w286 ), .B(
        \SUBBYTES[7].a/w288 ), .Z(n13926) );
  XOR \SUBBYTES[7].a/U5058  ( .A(\SUBBYTES[7].a/w246 ), .B(
        \SUBBYTES[7].a/w278 ), .Z(n13927) );
  XOR \SUBBYTES[7].a/U5057  ( .A(\w1[7][1] ), .B(n13928), .Z(n14664) );
  XOR \SUBBYTES[7].a/U5056  ( .A(\w1[7][3] ), .B(\w1[7][2] ), .Z(n13928) );
  XOR \SUBBYTES[7].a/U5055  ( .A(\w1[7][6] ), .B(n14664), .Z(
        \SUBBYTES[7].a/w3378 ) );
  XOR \SUBBYTES[7].a/U5054  ( .A(\w1[7][0] ), .B(\SUBBYTES[7].a/w3378 ), .Z(
        \SUBBYTES[7].a/w3265 ) );
  XOR \SUBBYTES[7].a/U5053  ( .A(\w1[7][0] ), .B(n13929), .Z(
        \SUBBYTES[7].a/w3266 ) );
  XOR \SUBBYTES[7].a/U5052  ( .A(\w1[7][6] ), .B(\w1[7][5] ), .Z(n13929) );
  XOR \SUBBYTES[7].a/U5051  ( .A(\w1[7][5] ), .B(n14664), .Z(
        \SUBBYTES[7].a/w3396 ) );
  XOR \SUBBYTES[7].a/U5050  ( .A(n13931), .B(n13930), .Z(\SUBBYTES[7].a/w3389 ) );
  XOR \SUBBYTES[7].a/U5049  ( .A(\w1[7][3] ), .B(\w1[7][1] ), .Z(n13930) );
  XOR \SUBBYTES[7].a/U5048  ( .A(\w1[7][7] ), .B(\w1[7][4] ), .Z(n13931) );
  XOR \SUBBYTES[7].a/U5047  ( .A(\w1[7][0] ), .B(\SUBBYTES[7].a/w3389 ), .Z(
        \SUBBYTES[7].a/w3268 ) );
  XOR \SUBBYTES[7].a/U5046  ( .A(n13933), .B(n13932), .Z(\SUBBYTES[7].a/w3376 ) );
  XOR \SUBBYTES[7].a/U5045  ( .A(\SUBBYTES[7].a/w3337 ), .B(n1068), .Z(n13932)
         );
  XOR \SUBBYTES[7].a/U5044  ( .A(\SUBBYTES[7].a/w3330 ), .B(
        \SUBBYTES[7].a/w3333 ), .Z(n13933) );
  XOR \SUBBYTES[7].a/U5043  ( .A(n13935), .B(n13934), .Z(\SUBBYTES[7].a/w3377 ) );
  XOR \SUBBYTES[7].a/U5042  ( .A(\SUBBYTES[7].a/w3337 ), .B(n13543), .Z(n13934) );
  XOR \SUBBYTES[7].a/U5041  ( .A(\SUBBYTES[7].a/w3330 ), .B(n13542), .Z(n13935) );
  XOR \SUBBYTES[7].a/U5040  ( .A(\SUBBYTES[7].a/w3389 ), .B(n13936), .Z(
        \SUBBYTES[7].a/w3379 ) );
  XOR \SUBBYTES[7].a/U5039  ( .A(\w1[7][6] ), .B(\w1[7][5] ), .Z(n13936) );
  XOR \SUBBYTES[7].a/U5038  ( .A(n13938), .B(n13937), .Z(\SUBBYTES[7].a/w3380 ) );
  XOR \SUBBYTES[7].a/U5037  ( .A(n13543), .B(n1068), .Z(n13937) );
  XOR \SUBBYTES[7].a/U5036  ( .A(n13542), .B(\SUBBYTES[7].a/w3333 ), .Z(n13938) );
  XOR \SUBBYTES[7].a/U5035  ( .A(\w1[7][7] ), .B(\w1[7][2] ), .Z(n14670) );
  XOR \SUBBYTES[7].a/U5034  ( .A(n14670), .B(n13939), .Z(\SUBBYTES[7].a/w3381 ) );
  XOR \SUBBYTES[7].a/U5033  ( .A(\w1[7][5] ), .B(\w1[7][4] ), .Z(n13939) );
  XOR \SUBBYTES[7].a/U5032  ( .A(\w1[7][7] ), .B(\SUBBYTES[7].a/w3266 ), .Z(
        \SUBBYTES[7].a/w3269 ) );
  XOR \SUBBYTES[7].a/U5031  ( .A(\w1[7][1] ), .B(\SUBBYTES[7].a/w3266 ), .Z(
        \SUBBYTES[7].a/w3270 ) );
  XOR \SUBBYTES[7].a/U5030  ( .A(\w1[7][4] ), .B(\SUBBYTES[7].a/w3266 ), .Z(
        \SUBBYTES[7].a/w3271 ) );
  XOR \SUBBYTES[7].a/U5029  ( .A(\SUBBYTES[7].a/w3270 ), .B(n14670), .Z(
        \SUBBYTES[7].a/w3272 ) );
  XOR \SUBBYTES[7].a/U5028  ( .A(n14670), .B(n13940), .Z(\SUBBYTES[7].a/w3357 ) );
  XOR \SUBBYTES[7].a/U5027  ( .A(\w1[7][4] ), .B(\w1[7][1] ), .Z(n13940) );
  XOR \SUBBYTES[7].a/U5026  ( .A(n13942), .B(n13941), .Z(n14667) );
  XOR \SUBBYTES[7].a/U5025  ( .A(\w1[7][4] ), .B(n13943), .Z(n13941) );
  XOR \SUBBYTES[7].a/U5024  ( .A(\SUBBYTES[7].a/w3322 ), .B(\w1[7][6] ), .Z(
        n13942) );
  XOR \SUBBYTES[7].a/U5023  ( .A(\SUBBYTES[7].a/w3296 ), .B(
        \SUBBYTES[7].a/w3303 ), .Z(n13943) );
  XOR \SUBBYTES[7].a/U5022  ( .A(n13945), .B(n13944), .Z(n14665) );
  XOR \SUBBYTES[7].a/U5021  ( .A(\w1[7][1] ), .B(n13946), .Z(n13944) );
  XOR \SUBBYTES[7].a/U5020  ( .A(\SUBBYTES[7].a/w3321 ), .B(\w1[7][5] ), .Z(
        n13945) );
  XOR \SUBBYTES[7].a/U5019  ( .A(\SUBBYTES[7].a/w3297 ), .B(
        \SUBBYTES[7].a/w3304 ), .Z(n13946) );
  XOR \SUBBYTES[7].a/U5018  ( .A(n14667), .B(n14665), .Z(\SUBBYTES[7].a/w3327 ) );
  XOR \SUBBYTES[7].a/U5017  ( .A(\w1[7][5] ), .B(n13947), .Z(n14668) );
  XOR \SUBBYTES[7].a/U5016  ( .A(\SUBBYTES[7].a/w3289 ), .B(
        \SUBBYTES[7].a/w3299 ), .Z(n13947) );
  XOR \SUBBYTES[7].a/U5015  ( .A(n13949), .B(n13948), .Z(\SUBBYTES[7].a/w3314 ) );
  XOR \SUBBYTES[7].a/U5014  ( .A(n14668), .B(n13950), .Z(n13948) );
  XOR \SUBBYTES[7].a/U5013  ( .A(\w1[7][4] ), .B(\SUBBYTES[7].a/w3378 ), .Z(
        n13949) );
  XOR \SUBBYTES[7].a/U5012  ( .A(\SUBBYTES[7].a/w3291 ), .B(
        \SUBBYTES[7].a/w3296 ), .Z(n13950) );
  XOR \SUBBYTES[7].a/U5011  ( .A(n13952), .B(n13951), .Z(n14666) );
  XOR \SUBBYTES[7].a/U5010  ( .A(\SUBBYTES[7].a/w3324 ), .B(\w1[7][7] ), .Z(
        n13951) );
  XOR \SUBBYTES[7].a/U5009  ( .A(\SUBBYTES[7].a/w3299 ), .B(
        \SUBBYTES[7].a/w3306 ), .Z(n13952) );
  XOR \SUBBYTES[7].a/U5008  ( .A(n14665), .B(n14666), .Z(\SUBBYTES[7].a/w3326 ) );
  XOR \SUBBYTES[7].a/U5007  ( .A(\w1[7][3] ), .B(n13953), .Z(n14669) );
  XOR \SUBBYTES[7].a/U5006  ( .A(\SUBBYTES[7].a/w3288 ), .B(
        \SUBBYTES[7].a/w3291 ), .Z(n13953) );
  XOR \SUBBYTES[7].a/U5005  ( .A(n13955), .B(n13954), .Z(\SUBBYTES[7].a/w3315 ) );
  XOR \SUBBYTES[7].a/U5004  ( .A(n14669), .B(n13956), .Z(n13954) );
  XOR \SUBBYTES[7].a/U5003  ( .A(\w1[7][6] ), .B(\SUBBYTES[7].a/w3357 ), .Z(
        n13955) );
  XOR \SUBBYTES[7].a/U5002  ( .A(\SUBBYTES[7].a/w3296 ), .B(
        \SUBBYTES[7].a/w3297 ), .Z(n13956) );
  XOR \SUBBYTES[7].a/U5001  ( .A(n14667), .B(n14666), .Z(\SUBBYTES[7].a/w3335 ) );
  XOR \SUBBYTES[7].a/U5000  ( .A(n13958), .B(n13957), .Z(\SUBBYTES[7].a/w3336 ) );
  XOR \SUBBYTES[7].a/U4999  ( .A(\w1[7][7] ), .B(n14668), .Z(n13957) );
  XOR \SUBBYTES[7].a/U4998  ( .A(\SUBBYTES[7].a/w3288 ), .B(
        \SUBBYTES[7].a/w3297 ), .Z(n13958) );
  XOR \SUBBYTES[7].a/U4997  ( .A(n13960), .B(n13959), .Z(\SUBBYTES[7].a/w3312 ) );
  XOR \SUBBYTES[7].a/U4996  ( .A(n13962), .B(n13961), .Z(n13959) );
  XOR \SUBBYTES[7].a/U4995  ( .A(\w1[7][7] ), .B(\SUBBYTES[7].a/w3396 ), .Z(
        n13960) );
  XOR \SUBBYTES[7].a/U4994  ( .A(\SUBBYTES[7].a/w3303 ), .B(
        \SUBBYTES[7].a/w3306 ), .Z(n13961) );
  XOR \SUBBYTES[7].a/U4993  ( .A(\SUBBYTES[7].a/w3289 ), .B(
        \SUBBYTES[7].a/w3291 ), .Z(n13962) );
  XOR \SUBBYTES[7].a/U4992  ( .A(n13964), .B(n13963), .Z(\SUBBYTES[7].a/w3313 ) );
  XOR \SUBBYTES[7].a/U4991  ( .A(n14669), .B(n13965), .Z(n13963) );
  XOR \SUBBYTES[7].a/U4990  ( .A(\w1[7][5] ), .B(n14670), .Z(n13964) );
  XOR \SUBBYTES[7].a/U4989  ( .A(\SUBBYTES[7].a/w3303 ), .B(
        \SUBBYTES[7].a/w3304 ), .Z(n13965) );
  XOR \SUBBYTES[7].a/U4988  ( .A(n13967), .B(n13966), .Z(\SUBBYTES[7].a/w3329 ) );
  XOR \SUBBYTES[7].a/U4987  ( .A(\w1[7][1] ), .B(n13968), .Z(n13966) );
  XOR \SUBBYTES[7].a/U4986  ( .A(\SUBBYTES[7].a/w3304 ), .B(
        \SUBBYTES[7].a/w3306 ), .Z(n13967) );
  XOR \SUBBYTES[7].a/U4985  ( .A(\SUBBYTES[7].a/w3288 ), .B(
        \SUBBYTES[7].a/w3289 ), .Z(n13968) );
  XOR \SUBBYTES[7].a/U4984  ( .A(\w1[7][9] ), .B(n13969), .Z(n14671) );
  XOR \SUBBYTES[7].a/U4983  ( .A(\w1[7][11] ), .B(\w1[7][10] ), .Z(n13969) );
  XOR \SUBBYTES[7].a/U4982  ( .A(\w1[7][14] ), .B(n14671), .Z(
        \SUBBYTES[7].a/w3171 ) );
  XOR \SUBBYTES[7].a/U4981  ( .A(\w1[7][8] ), .B(\SUBBYTES[7].a/w3171 ), .Z(
        \SUBBYTES[7].a/w3058 ) );
  XOR \SUBBYTES[7].a/U4980  ( .A(\w1[7][8] ), .B(n13970), .Z(
        \SUBBYTES[7].a/w3059 ) );
  XOR \SUBBYTES[7].a/U4979  ( .A(\w1[7][14] ), .B(\w1[7][13] ), .Z(n13970) );
  XOR \SUBBYTES[7].a/U4978  ( .A(\w1[7][13] ), .B(n14671), .Z(
        \SUBBYTES[7].a/w3189 ) );
  XOR \SUBBYTES[7].a/U4977  ( .A(n13972), .B(n13971), .Z(\SUBBYTES[7].a/w3182 ) );
  XOR \SUBBYTES[7].a/U4976  ( .A(\w1[7][11] ), .B(\w1[7][9] ), .Z(n13971) );
  XOR \SUBBYTES[7].a/U4975  ( .A(\w1[7][15] ), .B(\w1[7][12] ), .Z(n13972) );
  XOR \SUBBYTES[7].a/U4974  ( .A(\w1[7][8] ), .B(\SUBBYTES[7].a/w3182 ), .Z(
        \SUBBYTES[7].a/w3061 ) );
  XOR \SUBBYTES[7].a/U4973  ( .A(n13974), .B(n13973), .Z(\SUBBYTES[7].a/w3169 ) );
  XOR \SUBBYTES[7].a/U4972  ( .A(\SUBBYTES[7].a/w3130 ), .B(n1067), .Z(n13973)
         );
  XOR \SUBBYTES[7].a/U4971  ( .A(\SUBBYTES[7].a/w3123 ), .B(
        \SUBBYTES[7].a/w3126 ), .Z(n13974) );
  XOR \SUBBYTES[7].a/U4970  ( .A(n13976), .B(n13975), .Z(\SUBBYTES[7].a/w3170 ) );
  XOR \SUBBYTES[7].a/U4969  ( .A(\SUBBYTES[7].a/w3130 ), .B(n13541), .Z(n13975) );
  XOR \SUBBYTES[7].a/U4968  ( .A(\SUBBYTES[7].a/w3123 ), .B(n13540), .Z(n13976) );
  XOR \SUBBYTES[7].a/U4967  ( .A(\SUBBYTES[7].a/w3182 ), .B(n13977), .Z(
        \SUBBYTES[7].a/w3172 ) );
  XOR \SUBBYTES[7].a/U4966  ( .A(\w1[7][14] ), .B(\w1[7][13] ), .Z(n13977) );
  XOR \SUBBYTES[7].a/U4965  ( .A(n13979), .B(n13978), .Z(\SUBBYTES[7].a/w3173 ) );
  XOR \SUBBYTES[7].a/U4964  ( .A(n13541), .B(n1067), .Z(n13978) );
  XOR \SUBBYTES[7].a/U4963  ( .A(n13540), .B(\SUBBYTES[7].a/w3126 ), .Z(n13979) );
  XOR \SUBBYTES[7].a/U4962  ( .A(\w1[7][15] ), .B(\w1[7][10] ), .Z(n14677) );
  XOR \SUBBYTES[7].a/U4961  ( .A(n14677), .B(n13980), .Z(\SUBBYTES[7].a/w3174 ) );
  XOR \SUBBYTES[7].a/U4960  ( .A(\w1[7][13] ), .B(\w1[7][12] ), .Z(n13980) );
  XOR \SUBBYTES[7].a/U4959  ( .A(\w1[7][15] ), .B(\SUBBYTES[7].a/w3059 ), .Z(
        \SUBBYTES[7].a/w3062 ) );
  XOR \SUBBYTES[7].a/U4958  ( .A(\w1[7][9] ), .B(\SUBBYTES[7].a/w3059 ), .Z(
        \SUBBYTES[7].a/w3063 ) );
  XOR \SUBBYTES[7].a/U4957  ( .A(\w1[7][12] ), .B(\SUBBYTES[7].a/w3059 ), .Z(
        \SUBBYTES[7].a/w3064 ) );
  XOR \SUBBYTES[7].a/U4956  ( .A(\SUBBYTES[7].a/w3063 ), .B(n14677), .Z(
        \SUBBYTES[7].a/w3065 ) );
  XOR \SUBBYTES[7].a/U4955  ( .A(n14677), .B(n13981), .Z(\SUBBYTES[7].a/w3150 ) );
  XOR \SUBBYTES[7].a/U4954  ( .A(\w1[7][12] ), .B(\w1[7][9] ), .Z(n13981) );
  XOR \SUBBYTES[7].a/U4953  ( .A(n13983), .B(n13982), .Z(n14674) );
  XOR \SUBBYTES[7].a/U4952  ( .A(\w1[7][12] ), .B(n13984), .Z(n13982) );
  XOR \SUBBYTES[7].a/U4951  ( .A(\SUBBYTES[7].a/w3115 ), .B(\w1[7][14] ), .Z(
        n13983) );
  XOR \SUBBYTES[7].a/U4950  ( .A(\SUBBYTES[7].a/w3089 ), .B(
        \SUBBYTES[7].a/w3096 ), .Z(n13984) );
  XOR \SUBBYTES[7].a/U4949  ( .A(n13986), .B(n13985), .Z(n14672) );
  XOR \SUBBYTES[7].a/U4948  ( .A(\w1[7][9] ), .B(n13987), .Z(n13985) );
  XOR \SUBBYTES[7].a/U4947  ( .A(\SUBBYTES[7].a/w3114 ), .B(\w1[7][13] ), .Z(
        n13986) );
  XOR \SUBBYTES[7].a/U4946  ( .A(\SUBBYTES[7].a/w3090 ), .B(
        \SUBBYTES[7].a/w3097 ), .Z(n13987) );
  XOR \SUBBYTES[7].a/U4945  ( .A(n14674), .B(n14672), .Z(\SUBBYTES[7].a/w3120 ) );
  XOR \SUBBYTES[7].a/U4944  ( .A(\w1[7][13] ), .B(n13988), .Z(n14675) );
  XOR \SUBBYTES[7].a/U4943  ( .A(\SUBBYTES[7].a/w3082 ), .B(
        \SUBBYTES[7].a/w3092 ), .Z(n13988) );
  XOR \SUBBYTES[7].a/U4942  ( .A(n13990), .B(n13989), .Z(\SUBBYTES[7].a/w3107 ) );
  XOR \SUBBYTES[7].a/U4941  ( .A(n14675), .B(n13991), .Z(n13989) );
  XOR \SUBBYTES[7].a/U4940  ( .A(\w1[7][12] ), .B(\SUBBYTES[7].a/w3171 ), .Z(
        n13990) );
  XOR \SUBBYTES[7].a/U4939  ( .A(\SUBBYTES[7].a/w3084 ), .B(
        \SUBBYTES[7].a/w3089 ), .Z(n13991) );
  XOR \SUBBYTES[7].a/U4938  ( .A(n13993), .B(n13992), .Z(n14673) );
  XOR \SUBBYTES[7].a/U4937  ( .A(\SUBBYTES[7].a/w3117 ), .B(\w1[7][15] ), .Z(
        n13992) );
  XOR \SUBBYTES[7].a/U4936  ( .A(\SUBBYTES[7].a/w3092 ), .B(
        \SUBBYTES[7].a/w3099 ), .Z(n13993) );
  XOR \SUBBYTES[7].a/U4935  ( .A(n14672), .B(n14673), .Z(\SUBBYTES[7].a/w3119 ) );
  XOR \SUBBYTES[7].a/U4934  ( .A(\w1[7][11] ), .B(n13994), .Z(n14676) );
  XOR \SUBBYTES[7].a/U4933  ( .A(\SUBBYTES[7].a/w3081 ), .B(
        \SUBBYTES[7].a/w3084 ), .Z(n13994) );
  XOR \SUBBYTES[7].a/U4932  ( .A(n13996), .B(n13995), .Z(\SUBBYTES[7].a/w3108 ) );
  XOR \SUBBYTES[7].a/U4931  ( .A(n14676), .B(n13997), .Z(n13995) );
  XOR \SUBBYTES[7].a/U4930  ( .A(\w1[7][14] ), .B(\SUBBYTES[7].a/w3150 ), .Z(
        n13996) );
  XOR \SUBBYTES[7].a/U4929  ( .A(\SUBBYTES[7].a/w3089 ), .B(
        \SUBBYTES[7].a/w3090 ), .Z(n13997) );
  XOR \SUBBYTES[7].a/U4928  ( .A(n14674), .B(n14673), .Z(\SUBBYTES[7].a/w3128 ) );
  XOR \SUBBYTES[7].a/U4927  ( .A(n13999), .B(n13998), .Z(\SUBBYTES[7].a/w3129 ) );
  XOR \SUBBYTES[7].a/U4926  ( .A(\w1[7][15] ), .B(n14675), .Z(n13998) );
  XOR \SUBBYTES[7].a/U4925  ( .A(\SUBBYTES[7].a/w3081 ), .B(
        \SUBBYTES[7].a/w3090 ), .Z(n13999) );
  XOR \SUBBYTES[7].a/U4924  ( .A(n14001), .B(n14000), .Z(\SUBBYTES[7].a/w3105 ) );
  XOR \SUBBYTES[7].a/U4923  ( .A(n14003), .B(n14002), .Z(n14000) );
  XOR \SUBBYTES[7].a/U4922  ( .A(\w1[7][15] ), .B(\SUBBYTES[7].a/w3189 ), .Z(
        n14001) );
  XOR \SUBBYTES[7].a/U4921  ( .A(\SUBBYTES[7].a/w3096 ), .B(
        \SUBBYTES[7].a/w3099 ), .Z(n14002) );
  XOR \SUBBYTES[7].a/U4920  ( .A(\SUBBYTES[7].a/w3082 ), .B(
        \SUBBYTES[7].a/w3084 ), .Z(n14003) );
  XOR \SUBBYTES[7].a/U4919  ( .A(n14005), .B(n14004), .Z(\SUBBYTES[7].a/w3106 ) );
  XOR \SUBBYTES[7].a/U4918  ( .A(n14676), .B(n14006), .Z(n14004) );
  XOR \SUBBYTES[7].a/U4917  ( .A(\w1[7][13] ), .B(n14677), .Z(n14005) );
  XOR \SUBBYTES[7].a/U4916  ( .A(\SUBBYTES[7].a/w3096 ), .B(
        \SUBBYTES[7].a/w3097 ), .Z(n14006) );
  XOR \SUBBYTES[7].a/U4915  ( .A(n14008), .B(n14007), .Z(\SUBBYTES[7].a/w3122 ) );
  XOR \SUBBYTES[7].a/U4914  ( .A(\w1[7][9] ), .B(n14009), .Z(n14007) );
  XOR \SUBBYTES[7].a/U4913  ( .A(\SUBBYTES[7].a/w3097 ), .B(
        \SUBBYTES[7].a/w3099 ), .Z(n14008) );
  XOR \SUBBYTES[7].a/U4912  ( .A(\SUBBYTES[7].a/w3081 ), .B(
        \SUBBYTES[7].a/w3082 ), .Z(n14009) );
  XOR \SUBBYTES[7].a/U4911  ( .A(\w1[7][17] ), .B(n14010), .Z(n14678) );
  XOR \SUBBYTES[7].a/U4910  ( .A(\w1[7][19] ), .B(\w1[7][18] ), .Z(n14010) );
  XOR \SUBBYTES[7].a/U4909  ( .A(\w1[7][22] ), .B(n14678), .Z(
        \SUBBYTES[7].a/w2964 ) );
  XOR \SUBBYTES[7].a/U4908  ( .A(\w1[7][16] ), .B(\SUBBYTES[7].a/w2964 ), .Z(
        \SUBBYTES[7].a/w2851 ) );
  XOR \SUBBYTES[7].a/U4907  ( .A(\w1[7][16] ), .B(n14011), .Z(
        \SUBBYTES[7].a/w2852 ) );
  XOR \SUBBYTES[7].a/U4906  ( .A(\w1[7][22] ), .B(\w1[7][21] ), .Z(n14011) );
  XOR \SUBBYTES[7].a/U4905  ( .A(\w1[7][21] ), .B(n14678), .Z(
        \SUBBYTES[7].a/w2982 ) );
  XOR \SUBBYTES[7].a/U4904  ( .A(n14013), .B(n14012), .Z(\SUBBYTES[7].a/w2975 ) );
  XOR \SUBBYTES[7].a/U4903  ( .A(\w1[7][19] ), .B(\w1[7][17] ), .Z(n14012) );
  XOR \SUBBYTES[7].a/U4902  ( .A(\w1[7][23] ), .B(\w1[7][20] ), .Z(n14013) );
  XOR \SUBBYTES[7].a/U4901  ( .A(\w1[7][16] ), .B(\SUBBYTES[7].a/w2975 ), .Z(
        \SUBBYTES[7].a/w2854 ) );
  XOR \SUBBYTES[7].a/U4900  ( .A(n14015), .B(n14014), .Z(\SUBBYTES[7].a/w2962 ) );
  XOR \SUBBYTES[7].a/U4899  ( .A(\SUBBYTES[7].a/w2923 ), .B(n1066), .Z(n14014)
         );
  XOR \SUBBYTES[7].a/U4898  ( .A(\SUBBYTES[7].a/w2916 ), .B(
        \SUBBYTES[7].a/w2919 ), .Z(n14015) );
  XOR \SUBBYTES[7].a/U4897  ( .A(n14017), .B(n14016), .Z(\SUBBYTES[7].a/w2963 ) );
  XOR \SUBBYTES[7].a/U4896  ( .A(\SUBBYTES[7].a/w2923 ), .B(n13539), .Z(n14016) );
  XOR \SUBBYTES[7].a/U4895  ( .A(\SUBBYTES[7].a/w2916 ), .B(n13538), .Z(n14017) );
  XOR \SUBBYTES[7].a/U4894  ( .A(\SUBBYTES[7].a/w2975 ), .B(n14018), .Z(
        \SUBBYTES[7].a/w2965 ) );
  XOR \SUBBYTES[7].a/U4893  ( .A(\w1[7][22] ), .B(\w1[7][21] ), .Z(n14018) );
  XOR \SUBBYTES[7].a/U4892  ( .A(n14020), .B(n14019), .Z(\SUBBYTES[7].a/w2966 ) );
  XOR \SUBBYTES[7].a/U4891  ( .A(n13539), .B(n1066), .Z(n14019) );
  XOR \SUBBYTES[7].a/U4890  ( .A(n13538), .B(\SUBBYTES[7].a/w2919 ), .Z(n14020) );
  XOR \SUBBYTES[7].a/U4889  ( .A(\w1[7][23] ), .B(\w1[7][18] ), .Z(n14684) );
  XOR \SUBBYTES[7].a/U4888  ( .A(n14684), .B(n14021), .Z(\SUBBYTES[7].a/w2967 ) );
  XOR \SUBBYTES[7].a/U4887  ( .A(\w1[7][21] ), .B(\w1[7][20] ), .Z(n14021) );
  XOR \SUBBYTES[7].a/U4886  ( .A(\w1[7][23] ), .B(\SUBBYTES[7].a/w2852 ), .Z(
        \SUBBYTES[7].a/w2855 ) );
  XOR \SUBBYTES[7].a/U4885  ( .A(\w1[7][17] ), .B(\SUBBYTES[7].a/w2852 ), .Z(
        \SUBBYTES[7].a/w2856 ) );
  XOR \SUBBYTES[7].a/U4884  ( .A(\w1[7][20] ), .B(\SUBBYTES[7].a/w2852 ), .Z(
        \SUBBYTES[7].a/w2857 ) );
  XOR \SUBBYTES[7].a/U4883  ( .A(\SUBBYTES[7].a/w2856 ), .B(n14684), .Z(
        \SUBBYTES[7].a/w2858 ) );
  XOR \SUBBYTES[7].a/U4882  ( .A(n14684), .B(n14022), .Z(\SUBBYTES[7].a/w2943 ) );
  XOR \SUBBYTES[7].a/U4881  ( .A(\w1[7][20] ), .B(\w1[7][17] ), .Z(n14022) );
  XOR \SUBBYTES[7].a/U4880  ( .A(n14024), .B(n14023), .Z(n14681) );
  XOR \SUBBYTES[7].a/U4879  ( .A(\w1[7][20] ), .B(n14025), .Z(n14023) );
  XOR \SUBBYTES[7].a/U4878  ( .A(\SUBBYTES[7].a/w2908 ), .B(\w1[7][22] ), .Z(
        n14024) );
  XOR \SUBBYTES[7].a/U4877  ( .A(\SUBBYTES[7].a/w2882 ), .B(
        \SUBBYTES[7].a/w2889 ), .Z(n14025) );
  XOR \SUBBYTES[7].a/U4876  ( .A(n14027), .B(n14026), .Z(n14679) );
  XOR \SUBBYTES[7].a/U4875  ( .A(\w1[7][17] ), .B(n14028), .Z(n14026) );
  XOR \SUBBYTES[7].a/U4874  ( .A(\SUBBYTES[7].a/w2907 ), .B(\w1[7][21] ), .Z(
        n14027) );
  XOR \SUBBYTES[7].a/U4873  ( .A(\SUBBYTES[7].a/w2883 ), .B(
        \SUBBYTES[7].a/w2890 ), .Z(n14028) );
  XOR \SUBBYTES[7].a/U4872  ( .A(n14681), .B(n14679), .Z(\SUBBYTES[7].a/w2913 ) );
  XOR \SUBBYTES[7].a/U4871  ( .A(\w1[7][21] ), .B(n14029), .Z(n14682) );
  XOR \SUBBYTES[7].a/U4870  ( .A(\SUBBYTES[7].a/w2875 ), .B(
        \SUBBYTES[7].a/w2885 ), .Z(n14029) );
  XOR \SUBBYTES[7].a/U4869  ( .A(n14031), .B(n14030), .Z(\SUBBYTES[7].a/w2900 ) );
  XOR \SUBBYTES[7].a/U4868  ( .A(n14682), .B(n14032), .Z(n14030) );
  XOR \SUBBYTES[7].a/U4867  ( .A(\w1[7][20] ), .B(\SUBBYTES[7].a/w2964 ), .Z(
        n14031) );
  XOR \SUBBYTES[7].a/U4866  ( .A(\SUBBYTES[7].a/w2877 ), .B(
        \SUBBYTES[7].a/w2882 ), .Z(n14032) );
  XOR \SUBBYTES[7].a/U4865  ( .A(n14034), .B(n14033), .Z(n14680) );
  XOR \SUBBYTES[7].a/U4864  ( .A(\SUBBYTES[7].a/w2910 ), .B(\w1[7][23] ), .Z(
        n14033) );
  XOR \SUBBYTES[7].a/U4863  ( .A(\SUBBYTES[7].a/w2885 ), .B(
        \SUBBYTES[7].a/w2892 ), .Z(n14034) );
  XOR \SUBBYTES[7].a/U4862  ( .A(n14679), .B(n14680), .Z(\SUBBYTES[7].a/w2912 ) );
  XOR \SUBBYTES[7].a/U4861  ( .A(\w1[7][19] ), .B(n14035), .Z(n14683) );
  XOR \SUBBYTES[7].a/U4860  ( .A(\SUBBYTES[7].a/w2874 ), .B(
        \SUBBYTES[7].a/w2877 ), .Z(n14035) );
  XOR \SUBBYTES[7].a/U4859  ( .A(n14037), .B(n14036), .Z(\SUBBYTES[7].a/w2901 ) );
  XOR \SUBBYTES[7].a/U4858  ( .A(n14683), .B(n14038), .Z(n14036) );
  XOR \SUBBYTES[7].a/U4857  ( .A(\w1[7][22] ), .B(\SUBBYTES[7].a/w2943 ), .Z(
        n14037) );
  XOR \SUBBYTES[7].a/U4856  ( .A(\SUBBYTES[7].a/w2882 ), .B(
        \SUBBYTES[7].a/w2883 ), .Z(n14038) );
  XOR \SUBBYTES[7].a/U4855  ( .A(n14681), .B(n14680), .Z(\SUBBYTES[7].a/w2921 ) );
  XOR \SUBBYTES[7].a/U4854  ( .A(n14040), .B(n14039), .Z(\SUBBYTES[7].a/w2922 ) );
  XOR \SUBBYTES[7].a/U4853  ( .A(\w1[7][23] ), .B(n14682), .Z(n14039) );
  XOR \SUBBYTES[7].a/U4852  ( .A(\SUBBYTES[7].a/w2874 ), .B(
        \SUBBYTES[7].a/w2883 ), .Z(n14040) );
  XOR \SUBBYTES[7].a/U4851  ( .A(n14042), .B(n14041), .Z(\SUBBYTES[7].a/w2898 ) );
  XOR \SUBBYTES[7].a/U4850  ( .A(n14044), .B(n14043), .Z(n14041) );
  XOR \SUBBYTES[7].a/U4849  ( .A(\w1[7][23] ), .B(\SUBBYTES[7].a/w2982 ), .Z(
        n14042) );
  XOR \SUBBYTES[7].a/U4848  ( .A(\SUBBYTES[7].a/w2889 ), .B(
        \SUBBYTES[7].a/w2892 ), .Z(n14043) );
  XOR \SUBBYTES[7].a/U4847  ( .A(\SUBBYTES[7].a/w2875 ), .B(
        \SUBBYTES[7].a/w2877 ), .Z(n14044) );
  XOR \SUBBYTES[7].a/U4846  ( .A(n14046), .B(n14045), .Z(\SUBBYTES[7].a/w2899 ) );
  XOR \SUBBYTES[7].a/U4845  ( .A(n14683), .B(n14047), .Z(n14045) );
  XOR \SUBBYTES[7].a/U4844  ( .A(\w1[7][21] ), .B(n14684), .Z(n14046) );
  XOR \SUBBYTES[7].a/U4843  ( .A(\SUBBYTES[7].a/w2889 ), .B(
        \SUBBYTES[7].a/w2890 ), .Z(n14047) );
  XOR \SUBBYTES[7].a/U4842  ( .A(n14049), .B(n14048), .Z(\SUBBYTES[7].a/w2915 ) );
  XOR \SUBBYTES[7].a/U4841  ( .A(\w1[7][17] ), .B(n14050), .Z(n14048) );
  XOR \SUBBYTES[7].a/U4840  ( .A(\SUBBYTES[7].a/w2890 ), .B(
        \SUBBYTES[7].a/w2892 ), .Z(n14049) );
  XOR \SUBBYTES[7].a/U4839  ( .A(\SUBBYTES[7].a/w2874 ), .B(
        \SUBBYTES[7].a/w2875 ), .Z(n14050) );
  XOR \SUBBYTES[7].a/U4838  ( .A(\w1[7][25] ), .B(n14051), .Z(n14685) );
  XOR \SUBBYTES[7].a/U4837  ( .A(\w1[7][27] ), .B(\w1[7][26] ), .Z(n14051) );
  XOR \SUBBYTES[7].a/U4836  ( .A(\w1[7][30] ), .B(n14685), .Z(
        \SUBBYTES[7].a/w2757 ) );
  XOR \SUBBYTES[7].a/U4835  ( .A(\w1[7][24] ), .B(\SUBBYTES[7].a/w2757 ), .Z(
        \SUBBYTES[7].a/w2644 ) );
  XOR \SUBBYTES[7].a/U4834  ( .A(\w1[7][24] ), .B(n14052), .Z(
        \SUBBYTES[7].a/w2645 ) );
  XOR \SUBBYTES[7].a/U4833  ( .A(\w1[7][30] ), .B(\w1[7][29] ), .Z(n14052) );
  XOR \SUBBYTES[7].a/U4832  ( .A(\w1[7][29] ), .B(n14685), .Z(
        \SUBBYTES[7].a/w2775 ) );
  XOR \SUBBYTES[7].a/U4831  ( .A(n14054), .B(n14053), .Z(\SUBBYTES[7].a/w2768 ) );
  XOR \SUBBYTES[7].a/U4830  ( .A(\w1[7][27] ), .B(\w1[7][25] ), .Z(n14053) );
  XOR \SUBBYTES[7].a/U4829  ( .A(\w1[7][31] ), .B(\w1[7][28] ), .Z(n14054) );
  XOR \SUBBYTES[7].a/U4828  ( .A(\w1[7][24] ), .B(\SUBBYTES[7].a/w2768 ), .Z(
        \SUBBYTES[7].a/w2647 ) );
  XOR \SUBBYTES[7].a/U4827  ( .A(n14056), .B(n14055), .Z(\SUBBYTES[7].a/w2755 ) );
  XOR \SUBBYTES[7].a/U4826  ( .A(\SUBBYTES[7].a/w2716 ), .B(n1065), .Z(n14055)
         );
  XOR \SUBBYTES[7].a/U4825  ( .A(\SUBBYTES[7].a/w2709 ), .B(
        \SUBBYTES[7].a/w2712 ), .Z(n14056) );
  XOR \SUBBYTES[7].a/U4824  ( .A(n14058), .B(n14057), .Z(\SUBBYTES[7].a/w2756 ) );
  XOR \SUBBYTES[7].a/U4823  ( .A(\SUBBYTES[7].a/w2716 ), .B(n13537), .Z(n14057) );
  XOR \SUBBYTES[7].a/U4822  ( .A(\SUBBYTES[7].a/w2709 ), .B(n13536), .Z(n14058) );
  XOR \SUBBYTES[7].a/U4821  ( .A(\SUBBYTES[7].a/w2768 ), .B(n14059), .Z(
        \SUBBYTES[7].a/w2758 ) );
  XOR \SUBBYTES[7].a/U4820  ( .A(\w1[7][30] ), .B(\w1[7][29] ), .Z(n14059) );
  XOR \SUBBYTES[7].a/U4819  ( .A(n14061), .B(n14060), .Z(\SUBBYTES[7].a/w2759 ) );
  XOR \SUBBYTES[7].a/U4818  ( .A(n13537), .B(n1065), .Z(n14060) );
  XOR \SUBBYTES[7].a/U4817  ( .A(n13536), .B(\SUBBYTES[7].a/w2712 ), .Z(n14061) );
  XOR \SUBBYTES[7].a/U4816  ( .A(\w1[7][31] ), .B(\w1[7][26] ), .Z(n14691) );
  XOR \SUBBYTES[7].a/U4815  ( .A(n14691), .B(n14062), .Z(\SUBBYTES[7].a/w2760 ) );
  XOR \SUBBYTES[7].a/U4814  ( .A(\w1[7][29] ), .B(\w1[7][28] ), .Z(n14062) );
  XOR \SUBBYTES[7].a/U4813  ( .A(\w1[7][31] ), .B(\SUBBYTES[7].a/w2645 ), .Z(
        \SUBBYTES[7].a/w2648 ) );
  XOR \SUBBYTES[7].a/U4812  ( .A(\w1[7][25] ), .B(\SUBBYTES[7].a/w2645 ), .Z(
        \SUBBYTES[7].a/w2649 ) );
  XOR \SUBBYTES[7].a/U4811  ( .A(\w1[7][28] ), .B(\SUBBYTES[7].a/w2645 ), .Z(
        \SUBBYTES[7].a/w2650 ) );
  XOR \SUBBYTES[7].a/U4810  ( .A(\SUBBYTES[7].a/w2649 ), .B(n14691), .Z(
        \SUBBYTES[7].a/w2651 ) );
  XOR \SUBBYTES[7].a/U4809  ( .A(n14691), .B(n14063), .Z(\SUBBYTES[7].a/w2736 ) );
  XOR \SUBBYTES[7].a/U4808  ( .A(\w1[7][28] ), .B(\w1[7][25] ), .Z(n14063) );
  XOR \SUBBYTES[7].a/U4807  ( .A(n14065), .B(n14064), .Z(n14688) );
  XOR \SUBBYTES[7].a/U4806  ( .A(\w1[7][28] ), .B(n14066), .Z(n14064) );
  XOR \SUBBYTES[7].a/U4805  ( .A(\SUBBYTES[7].a/w2701 ), .B(\w1[7][30] ), .Z(
        n14065) );
  XOR \SUBBYTES[7].a/U4804  ( .A(\SUBBYTES[7].a/w2675 ), .B(
        \SUBBYTES[7].a/w2682 ), .Z(n14066) );
  XOR \SUBBYTES[7].a/U4803  ( .A(n14068), .B(n14067), .Z(n14686) );
  XOR \SUBBYTES[7].a/U4802  ( .A(\w1[7][25] ), .B(n14069), .Z(n14067) );
  XOR \SUBBYTES[7].a/U4801  ( .A(\SUBBYTES[7].a/w2700 ), .B(\w1[7][29] ), .Z(
        n14068) );
  XOR \SUBBYTES[7].a/U4800  ( .A(\SUBBYTES[7].a/w2676 ), .B(
        \SUBBYTES[7].a/w2683 ), .Z(n14069) );
  XOR \SUBBYTES[7].a/U4799  ( .A(n14688), .B(n14686), .Z(\SUBBYTES[7].a/w2706 ) );
  XOR \SUBBYTES[7].a/U4798  ( .A(\w1[7][29] ), .B(n14070), .Z(n14689) );
  XOR \SUBBYTES[7].a/U4797  ( .A(\SUBBYTES[7].a/w2668 ), .B(
        \SUBBYTES[7].a/w2678 ), .Z(n14070) );
  XOR \SUBBYTES[7].a/U4796  ( .A(n14072), .B(n14071), .Z(\SUBBYTES[7].a/w2693 ) );
  XOR \SUBBYTES[7].a/U4795  ( .A(n14689), .B(n14073), .Z(n14071) );
  XOR \SUBBYTES[7].a/U4794  ( .A(\w1[7][28] ), .B(\SUBBYTES[7].a/w2757 ), .Z(
        n14072) );
  XOR \SUBBYTES[7].a/U4793  ( .A(\SUBBYTES[7].a/w2670 ), .B(
        \SUBBYTES[7].a/w2675 ), .Z(n14073) );
  XOR \SUBBYTES[7].a/U4792  ( .A(n14075), .B(n14074), .Z(n14687) );
  XOR \SUBBYTES[7].a/U4791  ( .A(\SUBBYTES[7].a/w2703 ), .B(\w1[7][31] ), .Z(
        n14074) );
  XOR \SUBBYTES[7].a/U4790  ( .A(\SUBBYTES[7].a/w2678 ), .B(
        \SUBBYTES[7].a/w2685 ), .Z(n14075) );
  XOR \SUBBYTES[7].a/U4789  ( .A(n14686), .B(n14687), .Z(\SUBBYTES[7].a/w2705 ) );
  XOR \SUBBYTES[7].a/U4788  ( .A(\w1[7][27] ), .B(n14076), .Z(n14690) );
  XOR \SUBBYTES[7].a/U4787  ( .A(\SUBBYTES[7].a/w2667 ), .B(
        \SUBBYTES[7].a/w2670 ), .Z(n14076) );
  XOR \SUBBYTES[7].a/U4786  ( .A(n14078), .B(n14077), .Z(\SUBBYTES[7].a/w2694 ) );
  XOR \SUBBYTES[7].a/U4785  ( .A(n14690), .B(n14079), .Z(n14077) );
  XOR \SUBBYTES[7].a/U4784  ( .A(\w1[7][30] ), .B(\SUBBYTES[7].a/w2736 ), .Z(
        n14078) );
  XOR \SUBBYTES[7].a/U4783  ( .A(\SUBBYTES[7].a/w2675 ), .B(
        \SUBBYTES[7].a/w2676 ), .Z(n14079) );
  XOR \SUBBYTES[7].a/U4782  ( .A(n14688), .B(n14687), .Z(\SUBBYTES[7].a/w2714 ) );
  XOR \SUBBYTES[7].a/U4781  ( .A(n14081), .B(n14080), .Z(\SUBBYTES[7].a/w2715 ) );
  XOR \SUBBYTES[7].a/U4780  ( .A(\w1[7][31] ), .B(n14689), .Z(n14080) );
  XOR \SUBBYTES[7].a/U4779  ( .A(\SUBBYTES[7].a/w2667 ), .B(
        \SUBBYTES[7].a/w2676 ), .Z(n14081) );
  XOR \SUBBYTES[7].a/U4778  ( .A(n14083), .B(n14082), .Z(\SUBBYTES[7].a/w2691 ) );
  XOR \SUBBYTES[7].a/U4777  ( .A(n14085), .B(n14084), .Z(n14082) );
  XOR \SUBBYTES[7].a/U4776  ( .A(\w1[7][31] ), .B(\SUBBYTES[7].a/w2775 ), .Z(
        n14083) );
  XOR \SUBBYTES[7].a/U4775  ( .A(\SUBBYTES[7].a/w2682 ), .B(
        \SUBBYTES[7].a/w2685 ), .Z(n14084) );
  XOR \SUBBYTES[7].a/U4774  ( .A(\SUBBYTES[7].a/w2668 ), .B(
        \SUBBYTES[7].a/w2670 ), .Z(n14085) );
  XOR \SUBBYTES[7].a/U4773  ( .A(n14087), .B(n14086), .Z(\SUBBYTES[7].a/w2692 ) );
  XOR \SUBBYTES[7].a/U4772  ( .A(n14690), .B(n14088), .Z(n14086) );
  XOR \SUBBYTES[7].a/U4771  ( .A(\w1[7][29] ), .B(n14691), .Z(n14087) );
  XOR \SUBBYTES[7].a/U4770  ( .A(\SUBBYTES[7].a/w2682 ), .B(
        \SUBBYTES[7].a/w2683 ), .Z(n14088) );
  XOR \SUBBYTES[7].a/U4769  ( .A(n14090), .B(n14089), .Z(\SUBBYTES[7].a/w2708 ) );
  XOR \SUBBYTES[7].a/U4768  ( .A(\w1[7][25] ), .B(n14091), .Z(n14089) );
  XOR \SUBBYTES[7].a/U4767  ( .A(\SUBBYTES[7].a/w2683 ), .B(
        \SUBBYTES[7].a/w2685 ), .Z(n14090) );
  XOR \SUBBYTES[7].a/U4766  ( .A(\SUBBYTES[7].a/w2667 ), .B(
        \SUBBYTES[7].a/w2668 ), .Z(n14091) );
  XOR \SUBBYTES[7].a/U4765  ( .A(\w1[7][33] ), .B(n14092), .Z(n14692) );
  XOR \SUBBYTES[7].a/U4764  ( .A(\w1[7][35] ), .B(\w1[7][34] ), .Z(n14092) );
  XOR \SUBBYTES[7].a/U4763  ( .A(\w1[7][38] ), .B(n14692), .Z(
        \SUBBYTES[7].a/w2550 ) );
  XOR \SUBBYTES[7].a/U4762  ( .A(\w1[7][32] ), .B(\SUBBYTES[7].a/w2550 ), .Z(
        \SUBBYTES[7].a/w2437 ) );
  XOR \SUBBYTES[7].a/U4761  ( .A(\w1[7][32] ), .B(n14093), .Z(
        \SUBBYTES[7].a/w2438 ) );
  XOR \SUBBYTES[7].a/U4760  ( .A(\w1[7][38] ), .B(\w1[7][37] ), .Z(n14093) );
  XOR \SUBBYTES[7].a/U4759  ( .A(\w1[7][37] ), .B(n14692), .Z(
        \SUBBYTES[7].a/w2568 ) );
  XOR \SUBBYTES[7].a/U4758  ( .A(n14095), .B(n14094), .Z(\SUBBYTES[7].a/w2561 ) );
  XOR \SUBBYTES[7].a/U4757  ( .A(\w1[7][35] ), .B(\w1[7][33] ), .Z(n14094) );
  XOR \SUBBYTES[7].a/U4756  ( .A(\w1[7][39] ), .B(\w1[7][36] ), .Z(n14095) );
  XOR \SUBBYTES[7].a/U4755  ( .A(\w1[7][32] ), .B(\SUBBYTES[7].a/w2561 ), .Z(
        \SUBBYTES[7].a/w2440 ) );
  XOR \SUBBYTES[7].a/U4754  ( .A(n14097), .B(n14096), .Z(\SUBBYTES[7].a/w2548 ) );
  XOR \SUBBYTES[7].a/U4753  ( .A(\SUBBYTES[7].a/w2509 ), .B(n1064), .Z(n14096)
         );
  XOR \SUBBYTES[7].a/U4752  ( .A(\SUBBYTES[7].a/w2502 ), .B(
        \SUBBYTES[7].a/w2505 ), .Z(n14097) );
  XOR \SUBBYTES[7].a/U4751  ( .A(n14099), .B(n14098), .Z(\SUBBYTES[7].a/w2549 ) );
  XOR \SUBBYTES[7].a/U4750  ( .A(\SUBBYTES[7].a/w2509 ), .B(n13535), .Z(n14098) );
  XOR \SUBBYTES[7].a/U4749  ( .A(\SUBBYTES[7].a/w2502 ), .B(n13534), .Z(n14099) );
  XOR \SUBBYTES[7].a/U4748  ( .A(\SUBBYTES[7].a/w2561 ), .B(n14100), .Z(
        \SUBBYTES[7].a/w2551 ) );
  XOR \SUBBYTES[7].a/U4747  ( .A(\w1[7][38] ), .B(\w1[7][37] ), .Z(n14100) );
  XOR \SUBBYTES[7].a/U4746  ( .A(n14102), .B(n14101), .Z(\SUBBYTES[7].a/w2552 ) );
  XOR \SUBBYTES[7].a/U4745  ( .A(n13535), .B(n1064), .Z(n14101) );
  XOR \SUBBYTES[7].a/U4744  ( .A(n13534), .B(\SUBBYTES[7].a/w2505 ), .Z(n14102) );
  XOR \SUBBYTES[7].a/U4743  ( .A(\w1[7][39] ), .B(\w1[7][34] ), .Z(n14698) );
  XOR \SUBBYTES[7].a/U4742  ( .A(n14698), .B(n14103), .Z(\SUBBYTES[7].a/w2553 ) );
  XOR \SUBBYTES[7].a/U4741  ( .A(\w1[7][37] ), .B(\w1[7][36] ), .Z(n14103) );
  XOR \SUBBYTES[7].a/U4740  ( .A(\w1[7][39] ), .B(\SUBBYTES[7].a/w2438 ), .Z(
        \SUBBYTES[7].a/w2441 ) );
  XOR \SUBBYTES[7].a/U4739  ( .A(\w1[7][33] ), .B(\SUBBYTES[7].a/w2438 ), .Z(
        \SUBBYTES[7].a/w2442 ) );
  XOR \SUBBYTES[7].a/U4738  ( .A(\w1[7][36] ), .B(\SUBBYTES[7].a/w2438 ), .Z(
        \SUBBYTES[7].a/w2443 ) );
  XOR \SUBBYTES[7].a/U4737  ( .A(\SUBBYTES[7].a/w2442 ), .B(n14698), .Z(
        \SUBBYTES[7].a/w2444 ) );
  XOR \SUBBYTES[7].a/U4736  ( .A(n14698), .B(n14104), .Z(\SUBBYTES[7].a/w2529 ) );
  XOR \SUBBYTES[7].a/U4735  ( .A(\w1[7][36] ), .B(\w1[7][33] ), .Z(n14104) );
  XOR \SUBBYTES[7].a/U4734  ( .A(n14106), .B(n14105), .Z(n14695) );
  XOR \SUBBYTES[7].a/U4733  ( .A(\w1[7][36] ), .B(n14107), .Z(n14105) );
  XOR \SUBBYTES[7].a/U4732  ( .A(\SUBBYTES[7].a/w2494 ), .B(\w1[7][38] ), .Z(
        n14106) );
  XOR \SUBBYTES[7].a/U4731  ( .A(\SUBBYTES[7].a/w2468 ), .B(
        \SUBBYTES[7].a/w2475 ), .Z(n14107) );
  XOR \SUBBYTES[7].a/U4730  ( .A(n14109), .B(n14108), .Z(n14693) );
  XOR \SUBBYTES[7].a/U4729  ( .A(\w1[7][33] ), .B(n14110), .Z(n14108) );
  XOR \SUBBYTES[7].a/U4728  ( .A(\SUBBYTES[7].a/w2493 ), .B(\w1[7][37] ), .Z(
        n14109) );
  XOR \SUBBYTES[7].a/U4727  ( .A(\SUBBYTES[7].a/w2469 ), .B(
        \SUBBYTES[7].a/w2476 ), .Z(n14110) );
  XOR \SUBBYTES[7].a/U4726  ( .A(n14695), .B(n14693), .Z(\SUBBYTES[7].a/w2499 ) );
  XOR \SUBBYTES[7].a/U4725  ( .A(\w1[7][37] ), .B(n14111), .Z(n14696) );
  XOR \SUBBYTES[7].a/U4724  ( .A(\SUBBYTES[7].a/w2461 ), .B(
        \SUBBYTES[7].a/w2471 ), .Z(n14111) );
  XOR \SUBBYTES[7].a/U4723  ( .A(n14113), .B(n14112), .Z(\SUBBYTES[7].a/w2486 ) );
  XOR \SUBBYTES[7].a/U4722  ( .A(n14696), .B(n14114), .Z(n14112) );
  XOR \SUBBYTES[7].a/U4721  ( .A(\w1[7][36] ), .B(\SUBBYTES[7].a/w2550 ), .Z(
        n14113) );
  XOR \SUBBYTES[7].a/U4720  ( .A(\SUBBYTES[7].a/w2463 ), .B(
        \SUBBYTES[7].a/w2468 ), .Z(n14114) );
  XOR \SUBBYTES[7].a/U4719  ( .A(n14116), .B(n14115), .Z(n14694) );
  XOR \SUBBYTES[7].a/U4718  ( .A(\SUBBYTES[7].a/w2496 ), .B(\w1[7][39] ), .Z(
        n14115) );
  XOR \SUBBYTES[7].a/U4717  ( .A(\SUBBYTES[7].a/w2471 ), .B(
        \SUBBYTES[7].a/w2478 ), .Z(n14116) );
  XOR \SUBBYTES[7].a/U4716  ( .A(n14693), .B(n14694), .Z(\SUBBYTES[7].a/w2498 ) );
  XOR \SUBBYTES[7].a/U4715  ( .A(\w1[7][35] ), .B(n14117), .Z(n14697) );
  XOR \SUBBYTES[7].a/U4714  ( .A(\SUBBYTES[7].a/w2460 ), .B(
        \SUBBYTES[7].a/w2463 ), .Z(n14117) );
  XOR \SUBBYTES[7].a/U4713  ( .A(n14119), .B(n14118), .Z(\SUBBYTES[7].a/w2487 ) );
  XOR \SUBBYTES[7].a/U4712  ( .A(n14697), .B(n14120), .Z(n14118) );
  XOR \SUBBYTES[7].a/U4711  ( .A(\w1[7][38] ), .B(\SUBBYTES[7].a/w2529 ), .Z(
        n14119) );
  XOR \SUBBYTES[7].a/U4710  ( .A(\SUBBYTES[7].a/w2468 ), .B(
        \SUBBYTES[7].a/w2469 ), .Z(n14120) );
  XOR \SUBBYTES[7].a/U4709  ( .A(n14695), .B(n14694), .Z(\SUBBYTES[7].a/w2507 ) );
  XOR \SUBBYTES[7].a/U4708  ( .A(n14122), .B(n14121), .Z(\SUBBYTES[7].a/w2508 ) );
  XOR \SUBBYTES[7].a/U4707  ( .A(\w1[7][39] ), .B(n14696), .Z(n14121) );
  XOR \SUBBYTES[7].a/U4706  ( .A(\SUBBYTES[7].a/w2460 ), .B(
        \SUBBYTES[7].a/w2469 ), .Z(n14122) );
  XOR \SUBBYTES[7].a/U4705  ( .A(n14124), .B(n14123), .Z(\SUBBYTES[7].a/w2484 ) );
  XOR \SUBBYTES[7].a/U4704  ( .A(n14126), .B(n14125), .Z(n14123) );
  XOR \SUBBYTES[7].a/U4703  ( .A(\w1[7][39] ), .B(\SUBBYTES[7].a/w2568 ), .Z(
        n14124) );
  XOR \SUBBYTES[7].a/U4702  ( .A(\SUBBYTES[7].a/w2475 ), .B(
        \SUBBYTES[7].a/w2478 ), .Z(n14125) );
  XOR \SUBBYTES[7].a/U4701  ( .A(\SUBBYTES[7].a/w2461 ), .B(
        \SUBBYTES[7].a/w2463 ), .Z(n14126) );
  XOR \SUBBYTES[7].a/U4700  ( .A(n14128), .B(n14127), .Z(\SUBBYTES[7].a/w2485 ) );
  XOR \SUBBYTES[7].a/U4699  ( .A(n14697), .B(n14129), .Z(n14127) );
  XOR \SUBBYTES[7].a/U4698  ( .A(\w1[7][37] ), .B(n14698), .Z(n14128) );
  XOR \SUBBYTES[7].a/U4697  ( .A(\SUBBYTES[7].a/w2475 ), .B(
        \SUBBYTES[7].a/w2476 ), .Z(n14129) );
  XOR \SUBBYTES[7].a/U4696  ( .A(n14131), .B(n14130), .Z(\SUBBYTES[7].a/w2501 ) );
  XOR \SUBBYTES[7].a/U4695  ( .A(\w1[7][33] ), .B(n14132), .Z(n14130) );
  XOR \SUBBYTES[7].a/U4694  ( .A(\SUBBYTES[7].a/w2476 ), .B(
        \SUBBYTES[7].a/w2478 ), .Z(n14131) );
  XOR \SUBBYTES[7].a/U4693  ( .A(\SUBBYTES[7].a/w2460 ), .B(
        \SUBBYTES[7].a/w2461 ), .Z(n14132) );
  XOR \SUBBYTES[7].a/U4692  ( .A(\w1[7][41] ), .B(n14133), .Z(n14699) );
  XOR \SUBBYTES[7].a/U4691  ( .A(\w1[7][43] ), .B(\w1[7][42] ), .Z(n14133) );
  XOR \SUBBYTES[7].a/U4690  ( .A(\w1[7][46] ), .B(n14699), .Z(
        \SUBBYTES[7].a/w2343 ) );
  XOR \SUBBYTES[7].a/U4689  ( .A(\w1[7][40] ), .B(\SUBBYTES[7].a/w2343 ), .Z(
        \SUBBYTES[7].a/w2230 ) );
  XOR \SUBBYTES[7].a/U4688  ( .A(\w1[7][40] ), .B(n14134), .Z(
        \SUBBYTES[7].a/w2231 ) );
  XOR \SUBBYTES[7].a/U4687  ( .A(\w1[7][46] ), .B(\w1[7][45] ), .Z(n14134) );
  XOR \SUBBYTES[7].a/U4686  ( .A(\w1[7][45] ), .B(n14699), .Z(
        \SUBBYTES[7].a/w2361 ) );
  XOR \SUBBYTES[7].a/U4685  ( .A(n14136), .B(n14135), .Z(\SUBBYTES[7].a/w2354 ) );
  XOR \SUBBYTES[7].a/U4684  ( .A(\w1[7][43] ), .B(\w1[7][41] ), .Z(n14135) );
  XOR \SUBBYTES[7].a/U4683  ( .A(\w1[7][47] ), .B(\w1[7][44] ), .Z(n14136) );
  XOR \SUBBYTES[7].a/U4682  ( .A(\w1[7][40] ), .B(\SUBBYTES[7].a/w2354 ), .Z(
        \SUBBYTES[7].a/w2233 ) );
  XOR \SUBBYTES[7].a/U4681  ( .A(n14138), .B(n14137), .Z(\SUBBYTES[7].a/w2341 ) );
  XOR \SUBBYTES[7].a/U4680  ( .A(\SUBBYTES[7].a/w2302 ), .B(n1063), .Z(n14137)
         );
  XOR \SUBBYTES[7].a/U4679  ( .A(\SUBBYTES[7].a/w2295 ), .B(
        \SUBBYTES[7].a/w2298 ), .Z(n14138) );
  XOR \SUBBYTES[7].a/U4678  ( .A(n14140), .B(n14139), .Z(\SUBBYTES[7].a/w2342 ) );
  XOR \SUBBYTES[7].a/U4677  ( .A(\SUBBYTES[7].a/w2302 ), .B(n13533), .Z(n14139) );
  XOR \SUBBYTES[7].a/U4676  ( .A(\SUBBYTES[7].a/w2295 ), .B(n13532), .Z(n14140) );
  XOR \SUBBYTES[7].a/U4675  ( .A(\SUBBYTES[7].a/w2354 ), .B(n14141), .Z(
        \SUBBYTES[7].a/w2344 ) );
  XOR \SUBBYTES[7].a/U4674  ( .A(\w1[7][46] ), .B(\w1[7][45] ), .Z(n14141) );
  XOR \SUBBYTES[7].a/U4673  ( .A(n14143), .B(n14142), .Z(\SUBBYTES[7].a/w2345 ) );
  XOR \SUBBYTES[7].a/U4672  ( .A(n13533), .B(n1063), .Z(n14142) );
  XOR \SUBBYTES[7].a/U4671  ( .A(n13532), .B(\SUBBYTES[7].a/w2298 ), .Z(n14143) );
  XOR \SUBBYTES[7].a/U4670  ( .A(\w1[7][47] ), .B(\w1[7][42] ), .Z(n14705) );
  XOR \SUBBYTES[7].a/U4669  ( .A(n14705), .B(n14144), .Z(\SUBBYTES[7].a/w2346 ) );
  XOR \SUBBYTES[7].a/U4668  ( .A(\w1[7][45] ), .B(\w1[7][44] ), .Z(n14144) );
  XOR \SUBBYTES[7].a/U4667  ( .A(\w1[7][47] ), .B(\SUBBYTES[7].a/w2231 ), .Z(
        \SUBBYTES[7].a/w2234 ) );
  XOR \SUBBYTES[7].a/U4666  ( .A(\w1[7][41] ), .B(\SUBBYTES[7].a/w2231 ), .Z(
        \SUBBYTES[7].a/w2235 ) );
  XOR \SUBBYTES[7].a/U4665  ( .A(\w1[7][44] ), .B(\SUBBYTES[7].a/w2231 ), .Z(
        \SUBBYTES[7].a/w2236 ) );
  XOR \SUBBYTES[7].a/U4664  ( .A(\SUBBYTES[7].a/w2235 ), .B(n14705), .Z(
        \SUBBYTES[7].a/w2237 ) );
  XOR \SUBBYTES[7].a/U4663  ( .A(n14705), .B(n14145), .Z(\SUBBYTES[7].a/w2322 ) );
  XOR \SUBBYTES[7].a/U4662  ( .A(\w1[7][44] ), .B(\w1[7][41] ), .Z(n14145) );
  XOR \SUBBYTES[7].a/U4661  ( .A(n14147), .B(n14146), .Z(n14702) );
  XOR \SUBBYTES[7].a/U4660  ( .A(\w1[7][44] ), .B(n14148), .Z(n14146) );
  XOR \SUBBYTES[7].a/U4659  ( .A(\SUBBYTES[7].a/w2287 ), .B(\w1[7][46] ), .Z(
        n14147) );
  XOR \SUBBYTES[7].a/U4658  ( .A(\SUBBYTES[7].a/w2261 ), .B(
        \SUBBYTES[7].a/w2268 ), .Z(n14148) );
  XOR \SUBBYTES[7].a/U4657  ( .A(n14150), .B(n14149), .Z(n14700) );
  XOR \SUBBYTES[7].a/U4656  ( .A(\w1[7][41] ), .B(n14151), .Z(n14149) );
  XOR \SUBBYTES[7].a/U4655  ( .A(\SUBBYTES[7].a/w2286 ), .B(\w1[7][45] ), .Z(
        n14150) );
  XOR \SUBBYTES[7].a/U4654  ( .A(\SUBBYTES[7].a/w2262 ), .B(
        \SUBBYTES[7].a/w2269 ), .Z(n14151) );
  XOR \SUBBYTES[7].a/U4653  ( .A(n14702), .B(n14700), .Z(\SUBBYTES[7].a/w2292 ) );
  XOR \SUBBYTES[7].a/U4652  ( .A(\w1[7][45] ), .B(n14152), .Z(n14703) );
  XOR \SUBBYTES[7].a/U4651  ( .A(\SUBBYTES[7].a/w2254 ), .B(
        \SUBBYTES[7].a/w2264 ), .Z(n14152) );
  XOR \SUBBYTES[7].a/U4650  ( .A(n14154), .B(n14153), .Z(\SUBBYTES[7].a/w2279 ) );
  XOR \SUBBYTES[7].a/U4649  ( .A(n14703), .B(n14155), .Z(n14153) );
  XOR \SUBBYTES[7].a/U4648  ( .A(\w1[7][44] ), .B(\SUBBYTES[7].a/w2343 ), .Z(
        n14154) );
  XOR \SUBBYTES[7].a/U4647  ( .A(\SUBBYTES[7].a/w2256 ), .B(
        \SUBBYTES[7].a/w2261 ), .Z(n14155) );
  XOR \SUBBYTES[7].a/U4646  ( .A(n14157), .B(n14156), .Z(n14701) );
  XOR \SUBBYTES[7].a/U4645  ( .A(\SUBBYTES[7].a/w2289 ), .B(\w1[7][47] ), .Z(
        n14156) );
  XOR \SUBBYTES[7].a/U4644  ( .A(\SUBBYTES[7].a/w2264 ), .B(
        \SUBBYTES[7].a/w2271 ), .Z(n14157) );
  XOR \SUBBYTES[7].a/U4643  ( .A(n14700), .B(n14701), .Z(\SUBBYTES[7].a/w2291 ) );
  XOR \SUBBYTES[7].a/U4642  ( .A(\w1[7][43] ), .B(n14158), .Z(n14704) );
  XOR \SUBBYTES[7].a/U4641  ( .A(\SUBBYTES[7].a/w2253 ), .B(
        \SUBBYTES[7].a/w2256 ), .Z(n14158) );
  XOR \SUBBYTES[7].a/U4640  ( .A(n14160), .B(n14159), .Z(\SUBBYTES[7].a/w2280 ) );
  XOR \SUBBYTES[7].a/U4639  ( .A(n14704), .B(n14161), .Z(n14159) );
  XOR \SUBBYTES[7].a/U4638  ( .A(\w1[7][46] ), .B(\SUBBYTES[7].a/w2322 ), .Z(
        n14160) );
  XOR \SUBBYTES[7].a/U4637  ( .A(\SUBBYTES[7].a/w2261 ), .B(
        \SUBBYTES[7].a/w2262 ), .Z(n14161) );
  XOR \SUBBYTES[7].a/U4636  ( .A(n14702), .B(n14701), .Z(\SUBBYTES[7].a/w2300 ) );
  XOR \SUBBYTES[7].a/U4635  ( .A(n14163), .B(n14162), .Z(\SUBBYTES[7].a/w2301 ) );
  XOR \SUBBYTES[7].a/U4634  ( .A(\w1[7][47] ), .B(n14703), .Z(n14162) );
  XOR \SUBBYTES[7].a/U4633  ( .A(\SUBBYTES[7].a/w2253 ), .B(
        \SUBBYTES[7].a/w2262 ), .Z(n14163) );
  XOR \SUBBYTES[7].a/U4632  ( .A(n14165), .B(n14164), .Z(\SUBBYTES[7].a/w2277 ) );
  XOR \SUBBYTES[7].a/U4631  ( .A(n14167), .B(n14166), .Z(n14164) );
  XOR \SUBBYTES[7].a/U4630  ( .A(\w1[7][47] ), .B(\SUBBYTES[7].a/w2361 ), .Z(
        n14165) );
  XOR \SUBBYTES[7].a/U4629  ( .A(\SUBBYTES[7].a/w2268 ), .B(
        \SUBBYTES[7].a/w2271 ), .Z(n14166) );
  XOR \SUBBYTES[7].a/U4628  ( .A(\SUBBYTES[7].a/w2254 ), .B(
        \SUBBYTES[7].a/w2256 ), .Z(n14167) );
  XOR \SUBBYTES[7].a/U4627  ( .A(n14169), .B(n14168), .Z(\SUBBYTES[7].a/w2278 ) );
  XOR \SUBBYTES[7].a/U4626  ( .A(n14704), .B(n14170), .Z(n14168) );
  XOR \SUBBYTES[7].a/U4625  ( .A(\w1[7][45] ), .B(n14705), .Z(n14169) );
  XOR \SUBBYTES[7].a/U4624  ( .A(\SUBBYTES[7].a/w2268 ), .B(
        \SUBBYTES[7].a/w2269 ), .Z(n14170) );
  XOR \SUBBYTES[7].a/U4623  ( .A(n14172), .B(n14171), .Z(\SUBBYTES[7].a/w2294 ) );
  XOR \SUBBYTES[7].a/U4622  ( .A(\w1[7][41] ), .B(n14173), .Z(n14171) );
  XOR \SUBBYTES[7].a/U4621  ( .A(\SUBBYTES[7].a/w2269 ), .B(
        \SUBBYTES[7].a/w2271 ), .Z(n14172) );
  XOR \SUBBYTES[7].a/U4620  ( .A(\SUBBYTES[7].a/w2253 ), .B(
        \SUBBYTES[7].a/w2254 ), .Z(n14173) );
  XOR \SUBBYTES[7].a/U4619  ( .A(\w1[7][49] ), .B(n14174), .Z(n14706) );
  XOR \SUBBYTES[7].a/U4618  ( .A(\w1[7][51] ), .B(\w1[7][50] ), .Z(n14174) );
  XOR \SUBBYTES[7].a/U4617  ( .A(\w1[7][54] ), .B(n14706), .Z(
        \SUBBYTES[7].a/w2136 ) );
  XOR \SUBBYTES[7].a/U4616  ( .A(\w1[7][48] ), .B(\SUBBYTES[7].a/w2136 ), .Z(
        \SUBBYTES[7].a/w2023 ) );
  XOR \SUBBYTES[7].a/U4615  ( .A(\w1[7][48] ), .B(n14175), .Z(
        \SUBBYTES[7].a/w2024 ) );
  XOR \SUBBYTES[7].a/U4614  ( .A(\w1[7][54] ), .B(\w1[7][53] ), .Z(n14175) );
  XOR \SUBBYTES[7].a/U4613  ( .A(\w1[7][53] ), .B(n14706), .Z(
        \SUBBYTES[7].a/w2154 ) );
  XOR \SUBBYTES[7].a/U4612  ( .A(n14177), .B(n14176), .Z(\SUBBYTES[7].a/w2147 ) );
  XOR \SUBBYTES[7].a/U4611  ( .A(\w1[7][51] ), .B(\w1[7][49] ), .Z(n14176) );
  XOR \SUBBYTES[7].a/U4610  ( .A(\w1[7][55] ), .B(\w1[7][52] ), .Z(n14177) );
  XOR \SUBBYTES[7].a/U4609  ( .A(\w1[7][48] ), .B(\SUBBYTES[7].a/w2147 ), .Z(
        \SUBBYTES[7].a/w2026 ) );
  XOR \SUBBYTES[7].a/U4608  ( .A(n14179), .B(n14178), .Z(\SUBBYTES[7].a/w2134 ) );
  XOR \SUBBYTES[7].a/U4607  ( .A(\SUBBYTES[7].a/w2095 ), .B(n1062), .Z(n14178)
         );
  XOR \SUBBYTES[7].a/U4606  ( .A(\SUBBYTES[7].a/w2088 ), .B(
        \SUBBYTES[7].a/w2091 ), .Z(n14179) );
  XOR \SUBBYTES[7].a/U4605  ( .A(n14181), .B(n14180), .Z(\SUBBYTES[7].a/w2135 ) );
  XOR \SUBBYTES[7].a/U4604  ( .A(\SUBBYTES[7].a/w2095 ), .B(n13531), .Z(n14180) );
  XOR \SUBBYTES[7].a/U4603  ( .A(\SUBBYTES[7].a/w2088 ), .B(n13530), .Z(n14181) );
  XOR \SUBBYTES[7].a/U4602  ( .A(\SUBBYTES[7].a/w2147 ), .B(n14182), .Z(
        \SUBBYTES[7].a/w2137 ) );
  XOR \SUBBYTES[7].a/U4601  ( .A(\w1[7][54] ), .B(\w1[7][53] ), .Z(n14182) );
  XOR \SUBBYTES[7].a/U4600  ( .A(n14184), .B(n14183), .Z(\SUBBYTES[7].a/w2138 ) );
  XOR \SUBBYTES[7].a/U4599  ( .A(n13531), .B(n1062), .Z(n14183) );
  XOR \SUBBYTES[7].a/U4598  ( .A(n13530), .B(\SUBBYTES[7].a/w2091 ), .Z(n14184) );
  XOR \SUBBYTES[7].a/U4597  ( .A(\w1[7][55] ), .B(\w1[7][50] ), .Z(n14712) );
  XOR \SUBBYTES[7].a/U4596  ( .A(n14712), .B(n14185), .Z(\SUBBYTES[7].a/w2139 ) );
  XOR \SUBBYTES[7].a/U4595  ( .A(\w1[7][53] ), .B(\w1[7][52] ), .Z(n14185) );
  XOR \SUBBYTES[7].a/U4594  ( .A(\w1[7][55] ), .B(\SUBBYTES[7].a/w2024 ), .Z(
        \SUBBYTES[7].a/w2027 ) );
  XOR \SUBBYTES[7].a/U4593  ( .A(\w1[7][49] ), .B(\SUBBYTES[7].a/w2024 ), .Z(
        \SUBBYTES[7].a/w2028 ) );
  XOR \SUBBYTES[7].a/U4592  ( .A(\w1[7][52] ), .B(\SUBBYTES[7].a/w2024 ), .Z(
        \SUBBYTES[7].a/w2029 ) );
  XOR \SUBBYTES[7].a/U4591  ( .A(\SUBBYTES[7].a/w2028 ), .B(n14712), .Z(
        \SUBBYTES[7].a/w2030 ) );
  XOR \SUBBYTES[7].a/U4590  ( .A(n14712), .B(n14186), .Z(\SUBBYTES[7].a/w2115 ) );
  XOR \SUBBYTES[7].a/U4589  ( .A(\w1[7][52] ), .B(\w1[7][49] ), .Z(n14186) );
  XOR \SUBBYTES[7].a/U4588  ( .A(n14188), .B(n14187), .Z(n14709) );
  XOR \SUBBYTES[7].a/U4587  ( .A(\w1[7][52] ), .B(n14189), .Z(n14187) );
  XOR \SUBBYTES[7].a/U4586  ( .A(\SUBBYTES[7].a/w2080 ), .B(\w1[7][54] ), .Z(
        n14188) );
  XOR \SUBBYTES[7].a/U4585  ( .A(\SUBBYTES[7].a/w2054 ), .B(
        \SUBBYTES[7].a/w2061 ), .Z(n14189) );
  XOR \SUBBYTES[7].a/U4584  ( .A(n14191), .B(n14190), .Z(n14707) );
  XOR \SUBBYTES[7].a/U4583  ( .A(\w1[7][49] ), .B(n14192), .Z(n14190) );
  XOR \SUBBYTES[7].a/U4582  ( .A(\SUBBYTES[7].a/w2079 ), .B(\w1[7][53] ), .Z(
        n14191) );
  XOR \SUBBYTES[7].a/U4581  ( .A(\SUBBYTES[7].a/w2055 ), .B(
        \SUBBYTES[7].a/w2062 ), .Z(n14192) );
  XOR \SUBBYTES[7].a/U4580  ( .A(n14709), .B(n14707), .Z(\SUBBYTES[7].a/w2085 ) );
  XOR \SUBBYTES[7].a/U4579  ( .A(\w1[7][53] ), .B(n14193), .Z(n14710) );
  XOR \SUBBYTES[7].a/U4578  ( .A(\SUBBYTES[7].a/w2047 ), .B(
        \SUBBYTES[7].a/w2057 ), .Z(n14193) );
  XOR \SUBBYTES[7].a/U4577  ( .A(n14195), .B(n14194), .Z(\SUBBYTES[7].a/w2072 ) );
  XOR \SUBBYTES[7].a/U4576  ( .A(n14710), .B(n14196), .Z(n14194) );
  XOR \SUBBYTES[7].a/U4575  ( .A(\w1[7][52] ), .B(\SUBBYTES[7].a/w2136 ), .Z(
        n14195) );
  XOR \SUBBYTES[7].a/U4574  ( .A(\SUBBYTES[7].a/w2049 ), .B(
        \SUBBYTES[7].a/w2054 ), .Z(n14196) );
  XOR \SUBBYTES[7].a/U4573  ( .A(n14198), .B(n14197), .Z(n14708) );
  XOR \SUBBYTES[7].a/U4572  ( .A(\SUBBYTES[7].a/w2082 ), .B(\w1[7][55] ), .Z(
        n14197) );
  XOR \SUBBYTES[7].a/U4571  ( .A(\SUBBYTES[7].a/w2057 ), .B(
        \SUBBYTES[7].a/w2064 ), .Z(n14198) );
  XOR \SUBBYTES[7].a/U4570  ( .A(n14707), .B(n14708), .Z(\SUBBYTES[7].a/w2084 ) );
  XOR \SUBBYTES[7].a/U4569  ( .A(\w1[7][51] ), .B(n14199), .Z(n14711) );
  XOR \SUBBYTES[7].a/U4568  ( .A(\SUBBYTES[7].a/w2046 ), .B(
        \SUBBYTES[7].a/w2049 ), .Z(n14199) );
  XOR \SUBBYTES[7].a/U4567  ( .A(n14201), .B(n14200), .Z(\SUBBYTES[7].a/w2073 ) );
  XOR \SUBBYTES[7].a/U4566  ( .A(n14711), .B(n14202), .Z(n14200) );
  XOR \SUBBYTES[7].a/U4565  ( .A(\w1[7][54] ), .B(\SUBBYTES[7].a/w2115 ), .Z(
        n14201) );
  XOR \SUBBYTES[7].a/U4564  ( .A(\SUBBYTES[7].a/w2054 ), .B(
        \SUBBYTES[7].a/w2055 ), .Z(n14202) );
  XOR \SUBBYTES[7].a/U4563  ( .A(n14709), .B(n14708), .Z(\SUBBYTES[7].a/w2093 ) );
  XOR \SUBBYTES[7].a/U4562  ( .A(n14204), .B(n14203), .Z(\SUBBYTES[7].a/w2094 ) );
  XOR \SUBBYTES[7].a/U4561  ( .A(\w1[7][55] ), .B(n14710), .Z(n14203) );
  XOR \SUBBYTES[7].a/U4560  ( .A(\SUBBYTES[7].a/w2046 ), .B(
        \SUBBYTES[7].a/w2055 ), .Z(n14204) );
  XOR \SUBBYTES[7].a/U4559  ( .A(n14206), .B(n14205), .Z(\SUBBYTES[7].a/w2070 ) );
  XOR \SUBBYTES[7].a/U4558  ( .A(n14208), .B(n14207), .Z(n14205) );
  XOR \SUBBYTES[7].a/U4557  ( .A(\w1[7][55] ), .B(\SUBBYTES[7].a/w2154 ), .Z(
        n14206) );
  XOR \SUBBYTES[7].a/U4556  ( .A(\SUBBYTES[7].a/w2061 ), .B(
        \SUBBYTES[7].a/w2064 ), .Z(n14207) );
  XOR \SUBBYTES[7].a/U4555  ( .A(\SUBBYTES[7].a/w2047 ), .B(
        \SUBBYTES[7].a/w2049 ), .Z(n14208) );
  XOR \SUBBYTES[7].a/U4554  ( .A(n14210), .B(n14209), .Z(\SUBBYTES[7].a/w2071 ) );
  XOR \SUBBYTES[7].a/U4553  ( .A(n14711), .B(n14211), .Z(n14209) );
  XOR \SUBBYTES[7].a/U4552  ( .A(\w1[7][53] ), .B(n14712), .Z(n14210) );
  XOR \SUBBYTES[7].a/U4551  ( .A(\SUBBYTES[7].a/w2061 ), .B(
        \SUBBYTES[7].a/w2062 ), .Z(n14211) );
  XOR \SUBBYTES[7].a/U4550  ( .A(n14213), .B(n14212), .Z(\SUBBYTES[7].a/w2087 ) );
  XOR \SUBBYTES[7].a/U4549  ( .A(\w1[7][49] ), .B(n14214), .Z(n14212) );
  XOR \SUBBYTES[7].a/U4548  ( .A(\SUBBYTES[7].a/w2062 ), .B(
        \SUBBYTES[7].a/w2064 ), .Z(n14213) );
  XOR \SUBBYTES[7].a/U4547  ( .A(\SUBBYTES[7].a/w2046 ), .B(
        \SUBBYTES[7].a/w2047 ), .Z(n14214) );
  XOR \SUBBYTES[7].a/U4546  ( .A(\w1[7][57] ), .B(n14215), .Z(n14713) );
  XOR \SUBBYTES[7].a/U4545  ( .A(\w1[7][59] ), .B(\w1[7][58] ), .Z(n14215) );
  XOR \SUBBYTES[7].a/U4544  ( .A(\w1[7][62] ), .B(n14713), .Z(
        \SUBBYTES[7].a/w1929 ) );
  XOR \SUBBYTES[7].a/U4543  ( .A(\w1[7][56] ), .B(\SUBBYTES[7].a/w1929 ), .Z(
        \SUBBYTES[7].a/w1816 ) );
  XOR \SUBBYTES[7].a/U4542  ( .A(\w1[7][56] ), .B(n14216), .Z(
        \SUBBYTES[7].a/w1817 ) );
  XOR \SUBBYTES[7].a/U4541  ( .A(\w1[7][62] ), .B(\w1[7][61] ), .Z(n14216) );
  XOR \SUBBYTES[7].a/U4540  ( .A(\w1[7][61] ), .B(n14713), .Z(
        \SUBBYTES[7].a/w1947 ) );
  XOR \SUBBYTES[7].a/U4539  ( .A(n14218), .B(n14217), .Z(\SUBBYTES[7].a/w1940 ) );
  XOR \SUBBYTES[7].a/U4538  ( .A(\w1[7][59] ), .B(\w1[7][57] ), .Z(n14217) );
  XOR \SUBBYTES[7].a/U4537  ( .A(\w1[7][63] ), .B(\w1[7][60] ), .Z(n14218) );
  XOR \SUBBYTES[7].a/U4536  ( .A(\w1[7][56] ), .B(\SUBBYTES[7].a/w1940 ), .Z(
        \SUBBYTES[7].a/w1819 ) );
  XOR \SUBBYTES[7].a/U4535  ( .A(n14220), .B(n14219), .Z(\SUBBYTES[7].a/w1927 ) );
  XOR \SUBBYTES[7].a/U4534  ( .A(\SUBBYTES[7].a/w1888 ), .B(n1061), .Z(n14219)
         );
  XOR \SUBBYTES[7].a/U4533  ( .A(\SUBBYTES[7].a/w1881 ), .B(
        \SUBBYTES[7].a/w1884 ), .Z(n14220) );
  XOR \SUBBYTES[7].a/U4532  ( .A(n14222), .B(n14221), .Z(\SUBBYTES[7].a/w1928 ) );
  XOR \SUBBYTES[7].a/U4531  ( .A(\SUBBYTES[7].a/w1888 ), .B(n13529), .Z(n14221) );
  XOR \SUBBYTES[7].a/U4530  ( .A(\SUBBYTES[7].a/w1881 ), .B(n13528), .Z(n14222) );
  XOR \SUBBYTES[7].a/U4529  ( .A(\SUBBYTES[7].a/w1940 ), .B(n14223), .Z(
        \SUBBYTES[7].a/w1930 ) );
  XOR \SUBBYTES[7].a/U4528  ( .A(\w1[7][62] ), .B(\w1[7][61] ), .Z(n14223) );
  XOR \SUBBYTES[7].a/U4527  ( .A(n14225), .B(n14224), .Z(\SUBBYTES[7].a/w1931 ) );
  XOR \SUBBYTES[7].a/U4526  ( .A(n13529), .B(n1061), .Z(n14224) );
  XOR \SUBBYTES[7].a/U4525  ( .A(n13528), .B(\SUBBYTES[7].a/w1884 ), .Z(n14225) );
  XOR \SUBBYTES[7].a/U4524  ( .A(\w1[7][63] ), .B(\w1[7][58] ), .Z(n14719) );
  XOR \SUBBYTES[7].a/U4523  ( .A(n14719), .B(n14226), .Z(\SUBBYTES[7].a/w1932 ) );
  XOR \SUBBYTES[7].a/U4522  ( .A(\w1[7][61] ), .B(\w1[7][60] ), .Z(n14226) );
  XOR \SUBBYTES[7].a/U4521  ( .A(\w1[7][63] ), .B(\SUBBYTES[7].a/w1817 ), .Z(
        \SUBBYTES[7].a/w1820 ) );
  XOR \SUBBYTES[7].a/U4520  ( .A(\w1[7][57] ), .B(\SUBBYTES[7].a/w1817 ), .Z(
        \SUBBYTES[7].a/w1821 ) );
  XOR \SUBBYTES[7].a/U4519  ( .A(\w1[7][60] ), .B(\SUBBYTES[7].a/w1817 ), .Z(
        \SUBBYTES[7].a/w1822 ) );
  XOR \SUBBYTES[7].a/U4518  ( .A(\SUBBYTES[7].a/w1821 ), .B(n14719), .Z(
        \SUBBYTES[7].a/w1823 ) );
  XOR \SUBBYTES[7].a/U4517  ( .A(n14719), .B(n14227), .Z(\SUBBYTES[7].a/w1908 ) );
  XOR \SUBBYTES[7].a/U4516  ( .A(\w1[7][60] ), .B(\w1[7][57] ), .Z(n14227) );
  XOR \SUBBYTES[7].a/U4515  ( .A(n14229), .B(n14228), .Z(n14716) );
  XOR \SUBBYTES[7].a/U4514  ( .A(\w1[7][60] ), .B(n14230), .Z(n14228) );
  XOR \SUBBYTES[7].a/U4513  ( .A(\SUBBYTES[7].a/w1873 ), .B(\w1[7][62] ), .Z(
        n14229) );
  XOR \SUBBYTES[7].a/U4512  ( .A(\SUBBYTES[7].a/w1847 ), .B(
        \SUBBYTES[7].a/w1854 ), .Z(n14230) );
  XOR \SUBBYTES[7].a/U4511  ( .A(n14232), .B(n14231), .Z(n14714) );
  XOR \SUBBYTES[7].a/U4510  ( .A(\w1[7][57] ), .B(n14233), .Z(n14231) );
  XOR \SUBBYTES[7].a/U4509  ( .A(\SUBBYTES[7].a/w1872 ), .B(\w1[7][61] ), .Z(
        n14232) );
  XOR \SUBBYTES[7].a/U4508  ( .A(\SUBBYTES[7].a/w1848 ), .B(
        \SUBBYTES[7].a/w1855 ), .Z(n14233) );
  XOR \SUBBYTES[7].a/U4507  ( .A(n14716), .B(n14714), .Z(\SUBBYTES[7].a/w1878 ) );
  XOR \SUBBYTES[7].a/U4506  ( .A(\w1[7][61] ), .B(n14234), .Z(n14717) );
  XOR \SUBBYTES[7].a/U4505  ( .A(\SUBBYTES[7].a/w1840 ), .B(
        \SUBBYTES[7].a/w1850 ), .Z(n14234) );
  XOR \SUBBYTES[7].a/U4504  ( .A(n14236), .B(n14235), .Z(\SUBBYTES[7].a/w1865 ) );
  XOR \SUBBYTES[7].a/U4503  ( .A(n14717), .B(n14237), .Z(n14235) );
  XOR \SUBBYTES[7].a/U4502  ( .A(\w1[7][60] ), .B(\SUBBYTES[7].a/w1929 ), .Z(
        n14236) );
  XOR \SUBBYTES[7].a/U4501  ( .A(\SUBBYTES[7].a/w1842 ), .B(
        \SUBBYTES[7].a/w1847 ), .Z(n14237) );
  XOR \SUBBYTES[7].a/U4500  ( .A(n14239), .B(n14238), .Z(n14715) );
  XOR \SUBBYTES[7].a/U4499  ( .A(\SUBBYTES[7].a/w1875 ), .B(\w1[7][63] ), .Z(
        n14238) );
  XOR \SUBBYTES[7].a/U4498  ( .A(\SUBBYTES[7].a/w1850 ), .B(
        \SUBBYTES[7].a/w1857 ), .Z(n14239) );
  XOR \SUBBYTES[7].a/U4497  ( .A(n14714), .B(n14715), .Z(\SUBBYTES[7].a/w1877 ) );
  XOR \SUBBYTES[7].a/U4496  ( .A(\w1[7][59] ), .B(n14240), .Z(n14718) );
  XOR \SUBBYTES[7].a/U4495  ( .A(\SUBBYTES[7].a/w1839 ), .B(
        \SUBBYTES[7].a/w1842 ), .Z(n14240) );
  XOR \SUBBYTES[7].a/U4494  ( .A(n14242), .B(n14241), .Z(\SUBBYTES[7].a/w1866 ) );
  XOR \SUBBYTES[7].a/U4493  ( .A(n14718), .B(n14243), .Z(n14241) );
  XOR \SUBBYTES[7].a/U4492  ( .A(\w1[7][62] ), .B(\SUBBYTES[7].a/w1908 ), .Z(
        n14242) );
  XOR \SUBBYTES[7].a/U4491  ( .A(\SUBBYTES[7].a/w1847 ), .B(
        \SUBBYTES[7].a/w1848 ), .Z(n14243) );
  XOR \SUBBYTES[7].a/U4490  ( .A(n14716), .B(n14715), .Z(\SUBBYTES[7].a/w1886 ) );
  XOR \SUBBYTES[7].a/U4489  ( .A(n14245), .B(n14244), .Z(\SUBBYTES[7].a/w1887 ) );
  XOR \SUBBYTES[7].a/U4488  ( .A(\w1[7][63] ), .B(n14717), .Z(n14244) );
  XOR \SUBBYTES[7].a/U4487  ( .A(\SUBBYTES[7].a/w1839 ), .B(
        \SUBBYTES[7].a/w1848 ), .Z(n14245) );
  XOR \SUBBYTES[7].a/U4486  ( .A(n14247), .B(n14246), .Z(\SUBBYTES[7].a/w1863 ) );
  XOR \SUBBYTES[7].a/U4485  ( .A(n14249), .B(n14248), .Z(n14246) );
  XOR \SUBBYTES[7].a/U4484  ( .A(\w1[7][63] ), .B(\SUBBYTES[7].a/w1947 ), .Z(
        n14247) );
  XOR \SUBBYTES[7].a/U4483  ( .A(\SUBBYTES[7].a/w1854 ), .B(
        \SUBBYTES[7].a/w1857 ), .Z(n14248) );
  XOR \SUBBYTES[7].a/U4482  ( .A(\SUBBYTES[7].a/w1840 ), .B(
        \SUBBYTES[7].a/w1842 ), .Z(n14249) );
  XOR \SUBBYTES[7].a/U4481  ( .A(n14251), .B(n14250), .Z(\SUBBYTES[7].a/w1864 ) );
  XOR \SUBBYTES[7].a/U4480  ( .A(n14718), .B(n14252), .Z(n14250) );
  XOR \SUBBYTES[7].a/U4479  ( .A(\w1[7][61] ), .B(n14719), .Z(n14251) );
  XOR \SUBBYTES[7].a/U4478  ( .A(\SUBBYTES[7].a/w1854 ), .B(
        \SUBBYTES[7].a/w1855 ), .Z(n14252) );
  XOR \SUBBYTES[7].a/U4477  ( .A(n14254), .B(n14253), .Z(\SUBBYTES[7].a/w1880 ) );
  XOR \SUBBYTES[7].a/U4476  ( .A(\w1[7][57] ), .B(n14255), .Z(n14253) );
  XOR \SUBBYTES[7].a/U4475  ( .A(\SUBBYTES[7].a/w1855 ), .B(
        \SUBBYTES[7].a/w1857 ), .Z(n14254) );
  XOR \SUBBYTES[7].a/U4474  ( .A(\SUBBYTES[7].a/w1839 ), .B(
        \SUBBYTES[7].a/w1840 ), .Z(n14255) );
  XOR \SUBBYTES[7].a/U4473  ( .A(\w1[7][65] ), .B(n14256), .Z(n14720) );
  XOR \SUBBYTES[7].a/U4472  ( .A(\w1[7][67] ), .B(\w1[7][66] ), .Z(n14256) );
  XOR \SUBBYTES[7].a/U4471  ( .A(\w1[7][70] ), .B(n14720), .Z(
        \SUBBYTES[7].a/w1722 ) );
  XOR \SUBBYTES[7].a/U4470  ( .A(\w1[7][64] ), .B(\SUBBYTES[7].a/w1722 ), .Z(
        \SUBBYTES[7].a/w1609 ) );
  XOR \SUBBYTES[7].a/U4469  ( .A(\w1[7][64] ), .B(n14257), .Z(
        \SUBBYTES[7].a/w1610 ) );
  XOR \SUBBYTES[7].a/U4468  ( .A(\w1[7][70] ), .B(\w1[7][69] ), .Z(n14257) );
  XOR \SUBBYTES[7].a/U4467  ( .A(\w1[7][69] ), .B(n14720), .Z(
        \SUBBYTES[7].a/w1740 ) );
  XOR \SUBBYTES[7].a/U4466  ( .A(n14259), .B(n14258), .Z(\SUBBYTES[7].a/w1733 ) );
  XOR \SUBBYTES[7].a/U4465  ( .A(\w1[7][67] ), .B(\w1[7][65] ), .Z(n14258) );
  XOR \SUBBYTES[7].a/U4464  ( .A(\w1[7][71] ), .B(\w1[7][68] ), .Z(n14259) );
  XOR \SUBBYTES[7].a/U4463  ( .A(\w1[7][64] ), .B(\SUBBYTES[7].a/w1733 ), .Z(
        \SUBBYTES[7].a/w1612 ) );
  XOR \SUBBYTES[7].a/U4462  ( .A(n14261), .B(n14260), .Z(\SUBBYTES[7].a/w1720 ) );
  XOR \SUBBYTES[7].a/U4461  ( .A(\SUBBYTES[7].a/w1681 ), .B(n1060), .Z(n14260)
         );
  XOR \SUBBYTES[7].a/U4460  ( .A(\SUBBYTES[7].a/w1674 ), .B(
        \SUBBYTES[7].a/w1677 ), .Z(n14261) );
  XOR \SUBBYTES[7].a/U4459  ( .A(n14263), .B(n14262), .Z(\SUBBYTES[7].a/w1721 ) );
  XOR \SUBBYTES[7].a/U4458  ( .A(\SUBBYTES[7].a/w1681 ), .B(n13527), .Z(n14262) );
  XOR \SUBBYTES[7].a/U4457  ( .A(\SUBBYTES[7].a/w1674 ), .B(n13526), .Z(n14263) );
  XOR \SUBBYTES[7].a/U4456  ( .A(\SUBBYTES[7].a/w1733 ), .B(n14264), .Z(
        \SUBBYTES[7].a/w1723 ) );
  XOR \SUBBYTES[7].a/U4455  ( .A(\w1[7][70] ), .B(\w1[7][69] ), .Z(n14264) );
  XOR \SUBBYTES[7].a/U4454  ( .A(n14266), .B(n14265), .Z(\SUBBYTES[7].a/w1724 ) );
  XOR \SUBBYTES[7].a/U4453  ( .A(n13527), .B(n1060), .Z(n14265) );
  XOR \SUBBYTES[7].a/U4452  ( .A(n13526), .B(\SUBBYTES[7].a/w1677 ), .Z(n14266) );
  XOR \SUBBYTES[7].a/U4451  ( .A(\w1[7][71] ), .B(\w1[7][66] ), .Z(n14726) );
  XOR \SUBBYTES[7].a/U4450  ( .A(n14726), .B(n14267), .Z(\SUBBYTES[7].a/w1725 ) );
  XOR \SUBBYTES[7].a/U4449  ( .A(\w1[7][69] ), .B(\w1[7][68] ), .Z(n14267) );
  XOR \SUBBYTES[7].a/U4448  ( .A(\w1[7][71] ), .B(\SUBBYTES[7].a/w1610 ), .Z(
        \SUBBYTES[7].a/w1613 ) );
  XOR \SUBBYTES[7].a/U4447  ( .A(\w1[7][65] ), .B(\SUBBYTES[7].a/w1610 ), .Z(
        \SUBBYTES[7].a/w1614 ) );
  XOR \SUBBYTES[7].a/U4446  ( .A(\w1[7][68] ), .B(\SUBBYTES[7].a/w1610 ), .Z(
        \SUBBYTES[7].a/w1615 ) );
  XOR \SUBBYTES[7].a/U4445  ( .A(\SUBBYTES[7].a/w1614 ), .B(n14726), .Z(
        \SUBBYTES[7].a/w1616 ) );
  XOR \SUBBYTES[7].a/U4444  ( .A(n14726), .B(n14268), .Z(\SUBBYTES[7].a/w1701 ) );
  XOR \SUBBYTES[7].a/U4443  ( .A(\w1[7][68] ), .B(\w1[7][65] ), .Z(n14268) );
  XOR \SUBBYTES[7].a/U4442  ( .A(n14270), .B(n14269), .Z(n14723) );
  XOR \SUBBYTES[7].a/U4441  ( .A(\w1[7][68] ), .B(n14271), .Z(n14269) );
  XOR \SUBBYTES[7].a/U4440  ( .A(\SUBBYTES[7].a/w1666 ), .B(\w1[7][70] ), .Z(
        n14270) );
  XOR \SUBBYTES[7].a/U4439  ( .A(\SUBBYTES[7].a/w1640 ), .B(
        \SUBBYTES[7].a/w1647 ), .Z(n14271) );
  XOR \SUBBYTES[7].a/U4438  ( .A(n14273), .B(n14272), .Z(n14721) );
  XOR \SUBBYTES[7].a/U4437  ( .A(\w1[7][65] ), .B(n14274), .Z(n14272) );
  XOR \SUBBYTES[7].a/U4436  ( .A(\SUBBYTES[7].a/w1665 ), .B(\w1[7][69] ), .Z(
        n14273) );
  XOR \SUBBYTES[7].a/U4435  ( .A(\SUBBYTES[7].a/w1641 ), .B(
        \SUBBYTES[7].a/w1648 ), .Z(n14274) );
  XOR \SUBBYTES[7].a/U4434  ( .A(n14723), .B(n14721), .Z(\SUBBYTES[7].a/w1671 ) );
  XOR \SUBBYTES[7].a/U4433  ( .A(\w1[7][69] ), .B(n14275), .Z(n14724) );
  XOR \SUBBYTES[7].a/U4432  ( .A(\SUBBYTES[7].a/w1633 ), .B(
        \SUBBYTES[7].a/w1643 ), .Z(n14275) );
  XOR \SUBBYTES[7].a/U4431  ( .A(n14277), .B(n14276), .Z(\SUBBYTES[7].a/w1658 ) );
  XOR \SUBBYTES[7].a/U4430  ( .A(n14724), .B(n14278), .Z(n14276) );
  XOR \SUBBYTES[7].a/U4429  ( .A(\w1[7][68] ), .B(\SUBBYTES[7].a/w1722 ), .Z(
        n14277) );
  XOR \SUBBYTES[7].a/U4428  ( .A(\SUBBYTES[7].a/w1635 ), .B(
        \SUBBYTES[7].a/w1640 ), .Z(n14278) );
  XOR \SUBBYTES[7].a/U4427  ( .A(n14280), .B(n14279), .Z(n14722) );
  XOR \SUBBYTES[7].a/U4426  ( .A(\SUBBYTES[7].a/w1668 ), .B(\w1[7][71] ), .Z(
        n14279) );
  XOR \SUBBYTES[7].a/U4425  ( .A(\SUBBYTES[7].a/w1643 ), .B(
        \SUBBYTES[7].a/w1650 ), .Z(n14280) );
  XOR \SUBBYTES[7].a/U4424  ( .A(n14721), .B(n14722), .Z(\SUBBYTES[7].a/w1670 ) );
  XOR \SUBBYTES[7].a/U4423  ( .A(\w1[7][67] ), .B(n14281), .Z(n14725) );
  XOR \SUBBYTES[7].a/U4422  ( .A(\SUBBYTES[7].a/w1632 ), .B(
        \SUBBYTES[7].a/w1635 ), .Z(n14281) );
  XOR \SUBBYTES[7].a/U4421  ( .A(n14283), .B(n14282), .Z(\SUBBYTES[7].a/w1659 ) );
  XOR \SUBBYTES[7].a/U4420  ( .A(n14725), .B(n14284), .Z(n14282) );
  XOR \SUBBYTES[7].a/U4419  ( .A(\w1[7][70] ), .B(\SUBBYTES[7].a/w1701 ), .Z(
        n14283) );
  XOR \SUBBYTES[7].a/U4418  ( .A(\SUBBYTES[7].a/w1640 ), .B(
        \SUBBYTES[7].a/w1641 ), .Z(n14284) );
  XOR \SUBBYTES[7].a/U4417  ( .A(n14723), .B(n14722), .Z(\SUBBYTES[7].a/w1679 ) );
  XOR \SUBBYTES[7].a/U4416  ( .A(n14286), .B(n14285), .Z(\SUBBYTES[7].a/w1680 ) );
  XOR \SUBBYTES[7].a/U4415  ( .A(\w1[7][71] ), .B(n14724), .Z(n14285) );
  XOR \SUBBYTES[7].a/U4414  ( .A(\SUBBYTES[7].a/w1632 ), .B(
        \SUBBYTES[7].a/w1641 ), .Z(n14286) );
  XOR \SUBBYTES[7].a/U4413  ( .A(n14288), .B(n14287), .Z(\SUBBYTES[7].a/w1656 ) );
  XOR \SUBBYTES[7].a/U4412  ( .A(n14290), .B(n14289), .Z(n14287) );
  XOR \SUBBYTES[7].a/U4411  ( .A(\w1[7][71] ), .B(\SUBBYTES[7].a/w1740 ), .Z(
        n14288) );
  XOR \SUBBYTES[7].a/U4410  ( .A(\SUBBYTES[7].a/w1647 ), .B(
        \SUBBYTES[7].a/w1650 ), .Z(n14289) );
  XOR \SUBBYTES[7].a/U4409  ( .A(\SUBBYTES[7].a/w1633 ), .B(
        \SUBBYTES[7].a/w1635 ), .Z(n14290) );
  XOR \SUBBYTES[7].a/U4408  ( .A(n14292), .B(n14291), .Z(\SUBBYTES[7].a/w1657 ) );
  XOR \SUBBYTES[7].a/U4407  ( .A(n14725), .B(n14293), .Z(n14291) );
  XOR \SUBBYTES[7].a/U4406  ( .A(\w1[7][69] ), .B(n14726), .Z(n14292) );
  XOR \SUBBYTES[7].a/U4405  ( .A(\SUBBYTES[7].a/w1647 ), .B(
        \SUBBYTES[7].a/w1648 ), .Z(n14293) );
  XOR \SUBBYTES[7].a/U4404  ( .A(n14295), .B(n14294), .Z(\SUBBYTES[7].a/w1673 ) );
  XOR \SUBBYTES[7].a/U4403  ( .A(\w1[7][65] ), .B(n14296), .Z(n14294) );
  XOR \SUBBYTES[7].a/U4402  ( .A(\SUBBYTES[7].a/w1648 ), .B(
        \SUBBYTES[7].a/w1650 ), .Z(n14295) );
  XOR \SUBBYTES[7].a/U4401  ( .A(\SUBBYTES[7].a/w1632 ), .B(
        \SUBBYTES[7].a/w1633 ), .Z(n14296) );
  XOR \SUBBYTES[7].a/U4400  ( .A(\w1[7][73] ), .B(n14297), .Z(n14727) );
  XOR \SUBBYTES[7].a/U4399  ( .A(\w1[7][75] ), .B(\w1[7][74] ), .Z(n14297) );
  XOR \SUBBYTES[7].a/U4398  ( .A(\w1[7][78] ), .B(n14727), .Z(
        \SUBBYTES[7].a/w1515 ) );
  XOR \SUBBYTES[7].a/U4397  ( .A(\w1[7][72] ), .B(\SUBBYTES[7].a/w1515 ), .Z(
        \SUBBYTES[7].a/w1402 ) );
  XOR \SUBBYTES[7].a/U4396  ( .A(\w1[7][72] ), .B(n14298), .Z(
        \SUBBYTES[7].a/w1403 ) );
  XOR \SUBBYTES[7].a/U4395  ( .A(\w1[7][78] ), .B(\w1[7][77] ), .Z(n14298) );
  XOR \SUBBYTES[7].a/U4394  ( .A(\w1[7][77] ), .B(n14727), .Z(
        \SUBBYTES[7].a/w1533 ) );
  XOR \SUBBYTES[7].a/U4393  ( .A(n14300), .B(n14299), .Z(\SUBBYTES[7].a/w1526 ) );
  XOR \SUBBYTES[7].a/U4392  ( .A(\w1[7][75] ), .B(\w1[7][73] ), .Z(n14299) );
  XOR \SUBBYTES[7].a/U4391  ( .A(\w1[7][79] ), .B(\w1[7][76] ), .Z(n14300) );
  XOR \SUBBYTES[7].a/U4390  ( .A(\w1[7][72] ), .B(\SUBBYTES[7].a/w1526 ), .Z(
        \SUBBYTES[7].a/w1405 ) );
  XOR \SUBBYTES[7].a/U4389  ( .A(n14302), .B(n14301), .Z(\SUBBYTES[7].a/w1513 ) );
  XOR \SUBBYTES[7].a/U4388  ( .A(\SUBBYTES[7].a/w1474 ), .B(n1059), .Z(n14301)
         );
  XOR \SUBBYTES[7].a/U4387  ( .A(\SUBBYTES[7].a/w1467 ), .B(
        \SUBBYTES[7].a/w1470 ), .Z(n14302) );
  XOR \SUBBYTES[7].a/U4386  ( .A(n14304), .B(n14303), .Z(\SUBBYTES[7].a/w1514 ) );
  XOR \SUBBYTES[7].a/U4385  ( .A(\SUBBYTES[7].a/w1474 ), .B(n13525), .Z(n14303) );
  XOR \SUBBYTES[7].a/U4384  ( .A(\SUBBYTES[7].a/w1467 ), .B(n13524), .Z(n14304) );
  XOR \SUBBYTES[7].a/U4383  ( .A(\SUBBYTES[7].a/w1526 ), .B(n14305), .Z(
        \SUBBYTES[7].a/w1516 ) );
  XOR \SUBBYTES[7].a/U4382  ( .A(\w1[7][78] ), .B(\w1[7][77] ), .Z(n14305) );
  XOR \SUBBYTES[7].a/U4381  ( .A(n14307), .B(n14306), .Z(\SUBBYTES[7].a/w1517 ) );
  XOR \SUBBYTES[7].a/U4380  ( .A(n13525), .B(n1059), .Z(n14306) );
  XOR \SUBBYTES[7].a/U4379  ( .A(n13524), .B(\SUBBYTES[7].a/w1470 ), .Z(n14307) );
  XOR \SUBBYTES[7].a/U4378  ( .A(\w1[7][79] ), .B(\w1[7][74] ), .Z(n14733) );
  XOR \SUBBYTES[7].a/U4377  ( .A(n14733), .B(n14308), .Z(\SUBBYTES[7].a/w1518 ) );
  XOR \SUBBYTES[7].a/U4376  ( .A(\w1[7][77] ), .B(\w1[7][76] ), .Z(n14308) );
  XOR \SUBBYTES[7].a/U4375  ( .A(\w1[7][79] ), .B(\SUBBYTES[7].a/w1403 ), .Z(
        \SUBBYTES[7].a/w1406 ) );
  XOR \SUBBYTES[7].a/U4374  ( .A(\w1[7][73] ), .B(\SUBBYTES[7].a/w1403 ), .Z(
        \SUBBYTES[7].a/w1407 ) );
  XOR \SUBBYTES[7].a/U4373  ( .A(\w1[7][76] ), .B(\SUBBYTES[7].a/w1403 ), .Z(
        \SUBBYTES[7].a/w1408 ) );
  XOR \SUBBYTES[7].a/U4372  ( .A(\SUBBYTES[7].a/w1407 ), .B(n14733), .Z(
        \SUBBYTES[7].a/w1409 ) );
  XOR \SUBBYTES[7].a/U4371  ( .A(n14733), .B(n14309), .Z(\SUBBYTES[7].a/w1494 ) );
  XOR \SUBBYTES[7].a/U4370  ( .A(\w1[7][76] ), .B(\w1[7][73] ), .Z(n14309) );
  XOR \SUBBYTES[7].a/U4369  ( .A(n14311), .B(n14310), .Z(n14730) );
  XOR \SUBBYTES[7].a/U4368  ( .A(\w1[7][76] ), .B(n14312), .Z(n14310) );
  XOR \SUBBYTES[7].a/U4367  ( .A(\SUBBYTES[7].a/w1459 ), .B(\w1[7][78] ), .Z(
        n14311) );
  XOR \SUBBYTES[7].a/U4366  ( .A(\SUBBYTES[7].a/w1433 ), .B(
        \SUBBYTES[7].a/w1440 ), .Z(n14312) );
  XOR \SUBBYTES[7].a/U4365  ( .A(n14314), .B(n14313), .Z(n14728) );
  XOR \SUBBYTES[7].a/U4364  ( .A(\w1[7][73] ), .B(n14315), .Z(n14313) );
  XOR \SUBBYTES[7].a/U4363  ( .A(\SUBBYTES[7].a/w1458 ), .B(\w1[7][77] ), .Z(
        n14314) );
  XOR \SUBBYTES[7].a/U4362  ( .A(\SUBBYTES[7].a/w1434 ), .B(
        \SUBBYTES[7].a/w1441 ), .Z(n14315) );
  XOR \SUBBYTES[7].a/U4361  ( .A(n14730), .B(n14728), .Z(\SUBBYTES[7].a/w1464 ) );
  XOR \SUBBYTES[7].a/U4360  ( .A(\w1[7][77] ), .B(n14316), .Z(n14731) );
  XOR \SUBBYTES[7].a/U4359  ( .A(\SUBBYTES[7].a/w1426 ), .B(
        \SUBBYTES[7].a/w1436 ), .Z(n14316) );
  XOR \SUBBYTES[7].a/U4358  ( .A(n14318), .B(n14317), .Z(\SUBBYTES[7].a/w1451 ) );
  XOR \SUBBYTES[7].a/U4357  ( .A(n14731), .B(n14319), .Z(n14317) );
  XOR \SUBBYTES[7].a/U4356  ( .A(\w1[7][76] ), .B(\SUBBYTES[7].a/w1515 ), .Z(
        n14318) );
  XOR \SUBBYTES[7].a/U4355  ( .A(\SUBBYTES[7].a/w1428 ), .B(
        \SUBBYTES[7].a/w1433 ), .Z(n14319) );
  XOR \SUBBYTES[7].a/U4354  ( .A(n14321), .B(n14320), .Z(n14729) );
  XOR \SUBBYTES[7].a/U4353  ( .A(\SUBBYTES[7].a/w1461 ), .B(\w1[7][79] ), .Z(
        n14320) );
  XOR \SUBBYTES[7].a/U4352  ( .A(\SUBBYTES[7].a/w1436 ), .B(
        \SUBBYTES[7].a/w1443 ), .Z(n14321) );
  XOR \SUBBYTES[7].a/U4351  ( .A(n14728), .B(n14729), .Z(\SUBBYTES[7].a/w1463 ) );
  XOR \SUBBYTES[7].a/U4350  ( .A(\w1[7][75] ), .B(n14322), .Z(n14732) );
  XOR \SUBBYTES[7].a/U4349  ( .A(\SUBBYTES[7].a/w1425 ), .B(
        \SUBBYTES[7].a/w1428 ), .Z(n14322) );
  XOR \SUBBYTES[7].a/U4348  ( .A(n14324), .B(n14323), .Z(\SUBBYTES[7].a/w1452 ) );
  XOR \SUBBYTES[7].a/U4347  ( .A(n14732), .B(n14325), .Z(n14323) );
  XOR \SUBBYTES[7].a/U4346  ( .A(\w1[7][78] ), .B(\SUBBYTES[7].a/w1494 ), .Z(
        n14324) );
  XOR \SUBBYTES[7].a/U4345  ( .A(\SUBBYTES[7].a/w1433 ), .B(
        \SUBBYTES[7].a/w1434 ), .Z(n14325) );
  XOR \SUBBYTES[7].a/U4344  ( .A(n14730), .B(n14729), .Z(\SUBBYTES[7].a/w1472 ) );
  XOR \SUBBYTES[7].a/U4343  ( .A(n14327), .B(n14326), .Z(\SUBBYTES[7].a/w1473 ) );
  XOR \SUBBYTES[7].a/U4342  ( .A(\w1[7][79] ), .B(n14731), .Z(n14326) );
  XOR \SUBBYTES[7].a/U4341  ( .A(\SUBBYTES[7].a/w1425 ), .B(
        \SUBBYTES[7].a/w1434 ), .Z(n14327) );
  XOR \SUBBYTES[7].a/U4340  ( .A(n14329), .B(n14328), .Z(\SUBBYTES[7].a/w1449 ) );
  XOR \SUBBYTES[7].a/U4339  ( .A(n14331), .B(n14330), .Z(n14328) );
  XOR \SUBBYTES[7].a/U4338  ( .A(\w1[7][79] ), .B(\SUBBYTES[7].a/w1533 ), .Z(
        n14329) );
  XOR \SUBBYTES[7].a/U4337  ( .A(\SUBBYTES[7].a/w1440 ), .B(
        \SUBBYTES[7].a/w1443 ), .Z(n14330) );
  XOR \SUBBYTES[7].a/U4336  ( .A(\SUBBYTES[7].a/w1426 ), .B(
        \SUBBYTES[7].a/w1428 ), .Z(n14331) );
  XOR \SUBBYTES[7].a/U4335  ( .A(n14333), .B(n14332), .Z(\SUBBYTES[7].a/w1450 ) );
  XOR \SUBBYTES[7].a/U4334  ( .A(n14732), .B(n14334), .Z(n14332) );
  XOR \SUBBYTES[7].a/U4333  ( .A(\w1[7][77] ), .B(n14733), .Z(n14333) );
  XOR \SUBBYTES[7].a/U4332  ( .A(\SUBBYTES[7].a/w1440 ), .B(
        \SUBBYTES[7].a/w1441 ), .Z(n14334) );
  XOR \SUBBYTES[7].a/U4331  ( .A(n14336), .B(n14335), .Z(\SUBBYTES[7].a/w1466 ) );
  XOR \SUBBYTES[7].a/U4330  ( .A(\w1[7][73] ), .B(n14337), .Z(n14335) );
  XOR \SUBBYTES[7].a/U4329  ( .A(\SUBBYTES[7].a/w1441 ), .B(
        \SUBBYTES[7].a/w1443 ), .Z(n14336) );
  XOR \SUBBYTES[7].a/U4328  ( .A(\SUBBYTES[7].a/w1425 ), .B(
        \SUBBYTES[7].a/w1426 ), .Z(n14337) );
  XOR \SUBBYTES[7].a/U4327  ( .A(\w1[7][81] ), .B(n14338), .Z(n14734) );
  XOR \SUBBYTES[7].a/U4326  ( .A(\w1[7][83] ), .B(\w1[7][82] ), .Z(n14338) );
  XOR \SUBBYTES[7].a/U4325  ( .A(\w1[7][86] ), .B(n14734), .Z(
        \SUBBYTES[7].a/w1308 ) );
  XOR \SUBBYTES[7].a/U4324  ( .A(\w1[7][80] ), .B(\SUBBYTES[7].a/w1308 ), .Z(
        \SUBBYTES[7].a/w1195 ) );
  XOR \SUBBYTES[7].a/U4323  ( .A(\w1[7][80] ), .B(n14339), .Z(
        \SUBBYTES[7].a/w1196 ) );
  XOR \SUBBYTES[7].a/U4322  ( .A(\w1[7][86] ), .B(\w1[7][85] ), .Z(n14339) );
  XOR \SUBBYTES[7].a/U4321  ( .A(\w1[7][85] ), .B(n14734), .Z(
        \SUBBYTES[7].a/w1326 ) );
  XOR \SUBBYTES[7].a/U4320  ( .A(n14341), .B(n14340), .Z(\SUBBYTES[7].a/w1319 ) );
  XOR \SUBBYTES[7].a/U4319  ( .A(\w1[7][83] ), .B(\w1[7][81] ), .Z(n14340) );
  XOR \SUBBYTES[7].a/U4318  ( .A(\w1[7][87] ), .B(\w1[7][84] ), .Z(n14341) );
  XOR \SUBBYTES[7].a/U4317  ( .A(\w1[7][80] ), .B(\SUBBYTES[7].a/w1319 ), .Z(
        \SUBBYTES[7].a/w1198 ) );
  XOR \SUBBYTES[7].a/U4316  ( .A(n14343), .B(n14342), .Z(\SUBBYTES[7].a/w1306 ) );
  XOR \SUBBYTES[7].a/U4315  ( .A(\SUBBYTES[7].a/w1267 ), .B(n1058), .Z(n14342)
         );
  XOR \SUBBYTES[7].a/U4314  ( .A(\SUBBYTES[7].a/w1260 ), .B(
        \SUBBYTES[7].a/w1263 ), .Z(n14343) );
  XOR \SUBBYTES[7].a/U4313  ( .A(n14345), .B(n14344), .Z(\SUBBYTES[7].a/w1307 ) );
  XOR \SUBBYTES[7].a/U4312  ( .A(\SUBBYTES[7].a/w1267 ), .B(n13523), .Z(n14344) );
  XOR \SUBBYTES[7].a/U4311  ( .A(\SUBBYTES[7].a/w1260 ), .B(n13522), .Z(n14345) );
  XOR \SUBBYTES[7].a/U4310  ( .A(\SUBBYTES[7].a/w1319 ), .B(n14346), .Z(
        \SUBBYTES[7].a/w1309 ) );
  XOR \SUBBYTES[7].a/U4309  ( .A(\w1[7][86] ), .B(\w1[7][85] ), .Z(n14346) );
  XOR \SUBBYTES[7].a/U4308  ( .A(n14348), .B(n14347), .Z(\SUBBYTES[7].a/w1310 ) );
  XOR \SUBBYTES[7].a/U4307  ( .A(n13523), .B(n1058), .Z(n14347) );
  XOR \SUBBYTES[7].a/U4306  ( .A(n13522), .B(\SUBBYTES[7].a/w1263 ), .Z(n14348) );
  XOR \SUBBYTES[7].a/U4305  ( .A(\w1[7][87] ), .B(\w1[7][82] ), .Z(n14740) );
  XOR \SUBBYTES[7].a/U4304  ( .A(n14740), .B(n14349), .Z(\SUBBYTES[7].a/w1311 ) );
  XOR \SUBBYTES[7].a/U4303  ( .A(\w1[7][85] ), .B(\w1[7][84] ), .Z(n14349) );
  XOR \SUBBYTES[7].a/U4302  ( .A(\w1[7][87] ), .B(\SUBBYTES[7].a/w1196 ), .Z(
        \SUBBYTES[7].a/w1199 ) );
  XOR \SUBBYTES[7].a/U4301  ( .A(\w1[7][81] ), .B(\SUBBYTES[7].a/w1196 ), .Z(
        \SUBBYTES[7].a/w1200 ) );
  XOR \SUBBYTES[7].a/U4300  ( .A(\w1[7][84] ), .B(\SUBBYTES[7].a/w1196 ), .Z(
        \SUBBYTES[7].a/w1201 ) );
  XOR \SUBBYTES[7].a/U4299  ( .A(\SUBBYTES[7].a/w1200 ), .B(n14740), .Z(
        \SUBBYTES[7].a/w1202 ) );
  XOR \SUBBYTES[7].a/U4298  ( .A(n14740), .B(n14350), .Z(\SUBBYTES[7].a/w1287 ) );
  XOR \SUBBYTES[7].a/U4297  ( .A(\w1[7][84] ), .B(\w1[7][81] ), .Z(n14350) );
  XOR \SUBBYTES[7].a/U4296  ( .A(n14352), .B(n14351), .Z(n14737) );
  XOR \SUBBYTES[7].a/U4295  ( .A(\w1[7][84] ), .B(n14353), .Z(n14351) );
  XOR \SUBBYTES[7].a/U4294  ( .A(\SUBBYTES[7].a/w1252 ), .B(\w1[7][86] ), .Z(
        n14352) );
  XOR \SUBBYTES[7].a/U4293  ( .A(\SUBBYTES[7].a/w1226 ), .B(
        \SUBBYTES[7].a/w1233 ), .Z(n14353) );
  XOR \SUBBYTES[7].a/U4292  ( .A(n14355), .B(n14354), .Z(n14735) );
  XOR \SUBBYTES[7].a/U4291  ( .A(\w1[7][81] ), .B(n14356), .Z(n14354) );
  XOR \SUBBYTES[7].a/U4290  ( .A(\SUBBYTES[7].a/w1251 ), .B(\w1[7][85] ), .Z(
        n14355) );
  XOR \SUBBYTES[7].a/U4289  ( .A(\SUBBYTES[7].a/w1227 ), .B(
        \SUBBYTES[7].a/w1234 ), .Z(n14356) );
  XOR \SUBBYTES[7].a/U4288  ( .A(n14737), .B(n14735), .Z(\SUBBYTES[7].a/w1257 ) );
  XOR \SUBBYTES[7].a/U4287  ( .A(\w1[7][85] ), .B(n14357), .Z(n14738) );
  XOR \SUBBYTES[7].a/U4286  ( .A(\SUBBYTES[7].a/w1219 ), .B(
        \SUBBYTES[7].a/w1229 ), .Z(n14357) );
  XOR \SUBBYTES[7].a/U4285  ( .A(n14359), .B(n14358), .Z(\SUBBYTES[7].a/w1244 ) );
  XOR \SUBBYTES[7].a/U4284  ( .A(n14738), .B(n14360), .Z(n14358) );
  XOR \SUBBYTES[7].a/U4283  ( .A(\w1[7][84] ), .B(\SUBBYTES[7].a/w1308 ), .Z(
        n14359) );
  XOR \SUBBYTES[7].a/U4282  ( .A(\SUBBYTES[7].a/w1221 ), .B(
        \SUBBYTES[7].a/w1226 ), .Z(n14360) );
  XOR \SUBBYTES[7].a/U4281  ( .A(n14362), .B(n14361), .Z(n14736) );
  XOR \SUBBYTES[7].a/U4280  ( .A(\SUBBYTES[7].a/w1254 ), .B(\w1[7][87] ), .Z(
        n14361) );
  XOR \SUBBYTES[7].a/U4279  ( .A(\SUBBYTES[7].a/w1229 ), .B(
        \SUBBYTES[7].a/w1236 ), .Z(n14362) );
  XOR \SUBBYTES[7].a/U4278  ( .A(n14735), .B(n14736), .Z(\SUBBYTES[7].a/w1256 ) );
  XOR \SUBBYTES[7].a/U4277  ( .A(\w1[7][83] ), .B(n14363), .Z(n14739) );
  XOR \SUBBYTES[7].a/U4276  ( .A(\SUBBYTES[7].a/w1218 ), .B(
        \SUBBYTES[7].a/w1221 ), .Z(n14363) );
  XOR \SUBBYTES[7].a/U4275  ( .A(n14365), .B(n14364), .Z(\SUBBYTES[7].a/w1245 ) );
  XOR \SUBBYTES[7].a/U4274  ( .A(n14739), .B(n14366), .Z(n14364) );
  XOR \SUBBYTES[7].a/U4273  ( .A(\w1[7][86] ), .B(\SUBBYTES[7].a/w1287 ), .Z(
        n14365) );
  XOR \SUBBYTES[7].a/U4272  ( .A(\SUBBYTES[7].a/w1226 ), .B(
        \SUBBYTES[7].a/w1227 ), .Z(n14366) );
  XOR \SUBBYTES[7].a/U4271  ( .A(n14737), .B(n14736), .Z(\SUBBYTES[7].a/w1265 ) );
  XOR \SUBBYTES[7].a/U4270  ( .A(n14368), .B(n14367), .Z(\SUBBYTES[7].a/w1266 ) );
  XOR \SUBBYTES[7].a/U4269  ( .A(\w1[7][87] ), .B(n14738), .Z(n14367) );
  XOR \SUBBYTES[7].a/U4268  ( .A(\SUBBYTES[7].a/w1218 ), .B(
        \SUBBYTES[7].a/w1227 ), .Z(n14368) );
  XOR \SUBBYTES[7].a/U4267  ( .A(n14370), .B(n14369), .Z(\SUBBYTES[7].a/w1242 ) );
  XOR \SUBBYTES[7].a/U4266  ( .A(n14372), .B(n14371), .Z(n14369) );
  XOR \SUBBYTES[7].a/U4265  ( .A(\w1[7][87] ), .B(\SUBBYTES[7].a/w1326 ), .Z(
        n14370) );
  XOR \SUBBYTES[7].a/U4264  ( .A(\SUBBYTES[7].a/w1233 ), .B(
        \SUBBYTES[7].a/w1236 ), .Z(n14371) );
  XOR \SUBBYTES[7].a/U4263  ( .A(\SUBBYTES[7].a/w1219 ), .B(
        \SUBBYTES[7].a/w1221 ), .Z(n14372) );
  XOR \SUBBYTES[7].a/U4262  ( .A(n14374), .B(n14373), .Z(\SUBBYTES[7].a/w1243 ) );
  XOR \SUBBYTES[7].a/U4261  ( .A(n14739), .B(n14375), .Z(n14373) );
  XOR \SUBBYTES[7].a/U4260  ( .A(\w1[7][85] ), .B(n14740), .Z(n14374) );
  XOR \SUBBYTES[7].a/U4259  ( .A(\SUBBYTES[7].a/w1233 ), .B(
        \SUBBYTES[7].a/w1234 ), .Z(n14375) );
  XOR \SUBBYTES[7].a/U4258  ( .A(n14377), .B(n14376), .Z(\SUBBYTES[7].a/w1259 ) );
  XOR \SUBBYTES[7].a/U4257  ( .A(\w1[7][81] ), .B(n14378), .Z(n14376) );
  XOR \SUBBYTES[7].a/U4256  ( .A(\SUBBYTES[7].a/w1234 ), .B(
        \SUBBYTES[7].a/w1236 ), .Z(n14377) );
  XOR \SUBBYTES[7].a/U4255  ( .A(\SUBBYTES[7].a/w1218 ), .B(
        \SUBBYTES[7].a/w1219 ), .Z(n14378) );
  XOR \SUBBYTES[7].a/U4254  ( .A(\w1[7][89] ), .B(n14379), .Z(n14741) );
  XOR \SUBBYTES[7].a/U4253  ( .A(\w1[7][91] ), .B(\w1[7][90] ), .Z(n14379) );
  XOR \SUBBYTES[7].a/U4252  ( .A(\w1[7][94] ), .B(n14741), .Z(
        \SUBBYTES[7].a/w1101 ) );
  XOR \SUBBYTES[7].a/U4251  ( .A(\w1[7][88] ), .B(\SUBBYTES[7].a/w1101 ), .Z(
        \SUBBYTES[7].a/w988 ) );
  XOR \SUBBYTES[7].a/U4250  ( .A(\w1[7][88] ), .B(n14380), .Z(
        \SUBBYTES[7].a/w989 ) );
  XOR \SUBBYTES[7].a/U4249  ( .A(\w1[7][94] ), .B(\w1[7][93] ), .Z(n14380) );
  XOR \SUBBYTES[7].a/U4248  ( .A(\w1[7][93] ), .B(n14741), .Z(
        \SUBBYTES[7].a/w1119 ) );
  XOR \SUBBYTES[7].a/U4247  ( .A(n14382), .B(n14381), .Z(\SUBBYTES[7].a/w1112 ) );
  XOR \SUBBYTES[7].a/U4246  ( .A(\w1[7][91] ), .B(\w1[7][89] ), .Z(n14381) );
  XOR \SUBBYTES[7].a/U4245  ( .A(\w1[7][95] ), .B(\w1[7][92] ), .Z(n14382) );
  XOR \SUBBYTES[7].a/U4244  ( .A(\w1[7][88] ), .B(\SUBBYTES[7].a/w1112 ), .Z(
        \SUBBYTES[7].a/w991 ) );
  XOR \SUBBYTES[7].a/U4243  ( .A(n14384), .B(n14383), .Z(\SUBBYTES[7].a/w1099 ) );
  XOR \SUBBYTES[7].a/U4242  ( .A(\SUBBYTES[7].a/w1060 ), .B(n1057), .Z(n14383)
         );
  XOR \SUBBYTES[7].a/U4241  ( .A(\SUBBYTES[7].a/w1053 ), .B(
        \SUBBYTES[7].a/w1056 ), .Z(n14384) );
  XOR \SUBBYTES[7].a/U4240  ( .A(n14386), .B(n14385), .Z(\SUBBYTES[7].a/w1100 ) );
  XOR \SUBBYTES[7].a/U4239  ( .A(\SUBBYTES[7].a/w1060 ), .B(n13521), .Z(n14385) );
  XOR \SUBBYTES[7].a/U4238  ( .A(\SUBBYTES[7].a/w1053 ), .B(n13520), .Z(n14386) );
  XOR \SUBBYTES[7].a/U4237  ( .A(\SUBBYTES[7].a/w1112 ), .B(n14387), .Z(
        \SUBBYTES[7].a/w1102 ) );
  XOR \SUBBYTES[7].a/U4236  ( .A(\w1[7][94] ), .B(\w1[7][93] ), .Z(n14387) );
  XOR \SUBBYTES[7].a/U4235  ( .A(n14389), .B(n14388), .Z(\SUBBYTES[7].a/w1103 ) );
  XOR \SUBBYTES[7].a/U4234  ( .A(n13521), .B(n1057), .Z(n14388) );
  XOR \SUBBYTES[7].a/U4233  ( .A(n13520), .B(\SUBBYTES[7].a/w1056 ), .Z(n14389) );
  XOR \SUBBYTES[7].a/U4232  ( .A(\w1[7][95] ), .B(\w1[7][90] ), .Z(n14747) );
  XOR \SUBBYTES[7].a/U4231  ( .A(n14747), .B(n14390), .Z(\SUBBYTES[7].a/w1104 ) );
  XOR \SUBBYTES[7].a/U4230  ( .A(\w1[7][93] ), .B(\w1[7][92] ), .Z(n14390) );
  XOR \SUBBYTES[7].a/U4229  ( .A(\w1[7][95] ), .B(\SUBBYTES[7].a/w989 ), .Z(
        \SUBBYTES[7].a/w992 ) );
  XOR \SUBBYTES[7].a/U4228  ( .A(\w1[7][89] ), .B(\SUBBYTES[7].a/w989 ), .Z(
        \SUBBYTES[7].a/w993 ) );
  XOR \SUBBYTES[7].a/U4227  ( .A(\w1[7][92] ), .B(\SUBBYTES[7].a/w989 ), .Z(
        \SUBBYTES[7].a/w994 ) );
  XOR \SUBBYTES[7].a/U4226  ( .A(\SUBBYTES[7].a/w993 ), .B(n14747), .Z(
        \SUBBYTES[7].a/w995 ) );
  XOR \SUBBYTES[7].a/U4225  ( .A(n14747), .B(n14391), .Z(\SUBBYTES[7].a/w1080 ) );
  XOR \SUBBYTES[7].a/U4224  ( .A(\w1[7][92] ), .B(\w1[7][89] ), .Z(n14391) );
  XOR \SUBBYTES[7].a/U4223  ( .A(n14393), .B(n14392), .Z(n14744) );
  XOR \SUBBYTES[7].a/U4222  ( .A(\w1[7][92] ), .B(n14394), .Z(n14392) );
  XOR \SUBBYTES[7].a/U4221  ( .A(\SUBBYTES[7].a/w1045 ), .B(\w1[7][94] ), .Z(
        n14393) );
  XOR \SUBBYTES[7].a/U4220  ( .A(\SUBBYTES[7].a/w1019 ), .B(
        \SUBBYTES[7].a/w1026 ), .Z(n14394) );
  XOR \SUBBYTES[7].a/U4219  ( .A(n14396), .B(n14395), .Z(n14742) );
  XOR \SUBBYTES[7].a/U4218  ( .A(\w1[7][89] ), .B(n14397), .Z(n14395) );
  XOR \SUBBYTES[7].a/U4217  ( .A(\SUBBYTES[7].a/w1044 ), .B(\w1[7][93] ), .Z(
        n14396) );
  XOR \SUBBYTES[7].a/U4216  ( .A(\SUBBYTES[7].a/w1020 ), .B(
        \SUBBYTES[7].a/w1027 ), .Z(n14397) );
  XOR \SUBBYTES[7].a/U4215  ( .A(n14744), .B(n14742), .Z(\SUBBYTES[7].a/w1050 ) );
  XOR \SUBBYTES[7].a/U4214  ( .A(\w1[7][93] ), .B(n14398), .Z(n14745) );
  XOR \SUBBYTES[7].a/U4213  ( .A(\SUBBYTES[7].a/w1012 ), .B(
        \SUBBYTES[7].a/w1022 ), .Z(n14398) );
  XOR \SUBBYTES[7].a/U4212  ( .A(n14400), .B(n14399), .Z(\SUBBYTES[7].a/w1037 ) );
  XOR \SUBBYTES[7].a/U4211  ( .A(n14745), .B(n14401), .Z(n14399) );
  XOR \SUBBYTES[7].a/U4210  ( .A(\w1[7][92] ), .B(\SUBBYTES[7].a/w1101 ), .Z(
        n14400) );
  XOR \SUBBYTES[7].a/U4209  ( .A(\SUBBYTES[7].a/w1014 ), .B(
        \SUBBYTES[7].a/w1019 ), .Z(n14401) );
  XOR \SUBBYTES[7].a/U4208  ( .A(n14403), .B(n14402), .Z(n14743) );
  XOR \SUBBYTES[7].a/U4207  ( .A(\SUBBYTES[7].a/w1047 ), .B(\w1[7][95] ), .Z(
        n14402) );
  XOR \SUBBYTES[7].a/U4206  ( .A(\SUBBYTES[7].a/w1022 ), .B(
        \SUBBYTES[7].a/w1029 ), .Z(n14403) );
  XOR \SUBBYTES[7].a/U4205  ( .A(n14742), .B(n14743), .Z(\SUBBYTES[7].a/w1049 ) );
  XOR \SUBBYTES[7].a/U4204  ( .A(\w1[7][91] ), .B(n14404), .Z(n14746) );
  XOR \SUBBYTES[7].a/U4203  ( .A(\SUBBYTES[7].a/w1011 ), .B(
        \SUBBYTES[7].a/w1014 ), .Z(n14404) );
  XOR \SUBBYTES[7].a/U4202  ( .A(n14406), .B(n14405), .Z(\SUBBYTES[7].a/w1038 ) );
  XOR \SUBBYTES[7].a/U4201  ( .A(n14746), .B(n14407), .Z(n14405) );
  XOR \SUBBYTES[7].a/U4200  ( .A(\w1[7][94] ), .B(\SUBBYTES[7].a/w1080 ), .Z(
        n14406) );
  XOR \SUBBYTES[7].a/U4199  ( .A(\SUBBYTES[7].a/w1019 ), .B(
        \SUBBYTES[7].a/w1020 ), .Z(n14407) );
  XOR \SUBBYTES[7].a/U4198  ( .A(n14744), .B(n14743), .Z(\SUBBYTES[7].a/w1058 ) );
  XOR \SUBBYTES[7].a/U4197  ( .A(n14409), .B(n14408), .Z(\SUBBYTES[7].a/w1059 ) );
  XOR \SUBBYTES[7].a/U4196  ( .A(\w1[7][95] ), .B(n14745), .Z(n14408) );
  XOR \SUBBYTES[7].a/U4195  ( .A(\SUBBYTES[7].a/w1011 ), .B(
        \SUBBYTES[7].a/w1020 ), .Z(n14409) );
  XOR \SUBBYTES[7].a/U4194  ( .A(n14411), .B(n14410), .Z(\SUBBYTES[7].a/w1035 ) );
  XOR \SUBBYTES[7].a/U4193  ( .A(n14413), .B(n14412), .Z(n14410) );
  XOR \SUBBYTES[7].a/U4192  ( .A(\w1[7][95] ), .B(\SUBBYTES[7].a/w1119 ), .Z(
        n14411) );
  XOR \SUBBYTES[7].a/U4191  ( .A(\SUBBYTES[7].a/w1026 ), .B(
        \SUBBYTES[7].a/w1029 ), .Z(n14412) );
  XOR \SUBBYTES[7].a/U4190  ( .A(\SUBBYTES[7].a/w1012 ), .B(
        \SUBBYTES[7].a/w1014 ), .Z(n14413) );
  XOR \SUBBYTES[7].a/U4189  ( .A(n14415), .B(n14414), .Z(\SUBBYTES[7].a/w1036 ) );
  XOR \SUBBYTES[7].a/U4188  ( .A(n14746), .B(n14416), .Z(n14414) );
  XOR \SUBBYTES[7].a/U4187  ( .A(\w1[7][93] ), .B(n14747), .Z(n14415) );
  XOR \SUBBYTES[7].a/U4186  ( .A(\SUBBYTES[7].a/w1026 ), .B(
        \SUBBYTES[7].a/w1027 ), .Z(n14416) );
  XOR \SUBBYTES[7].a/U4185  ( .A(n14418), .B(n14417), .Z(\SUBBYTES[7].a/w1052 ) );
  XOR \SUBBYTES[7].a/U4184  ( .A(\w1[7][89] ), .B(n14419), .Z(n14417) );
  XOR \SUBBYTES[7].a/U4183  ( .A(\SUBBYTES[7].a/w1027 ), .B(
        \SUBBYTES[7].a/w1029 ), .Z(n14418) );
  XOR \SUBBYTES[7].a/U4182  ( .A(\SUBBYTES[7].a/w1011 ), .B(
        \SUBBYTES[7].a/w1012 ), .Z(n14419) );
  XOR \SUBBYTES[7].a/U4181  ( .A(\w1[7][97] ), .B(n14420), .Z(n14748) );
  XOR \SUBBYTES[7].a/U4180  ( .A(\w1[7][99] ), .B(\w1[7][98] ), .Z(n14420) );
  XOR \SUBBYTES[7].a/U4179  ( .A(\w1[7][102] ), .B(n14748), .Z(
        \SUBBYTES[7].a/w894 ) );
  XOR \SUBBYTES[7].a/U4178  ( .A(\w1[7][96] ), .B(\SUBBYTES[7].a/w894 ), .Z(
        \SUBBYTES[7].a/w781 ) );
  XOR \SUBBYTES[7].a/U4177  ( .A(\w1[7][96] ), .B(n14421), .Z(
        \SUBBYTES[7].a/w782 ) );
  XOR \SUBBYTES[7].a/U4176  ( .A(\w1[7][102] ), .B(\w1[7][101] ), .Z(n14421)
         );
  XOR \SUBBYTES[7].a/U4175  ( .A(\w1[7][101] ), .B(n14748), .Z(
        \SUBBYTES[7].a/w912 ) );
  XOR \SUBBYTES[7].a/U4174  ( .A(n14423), .B(n14422), .Z(\SUBBYTES[7].a/w905 )
         );
  XOR \SUBBYTES[7].a/U4173  ( .A(\w1[7][99] ), .B(\w1[7][97] ), .Z(n14422) );
  XOR \SUBBYTES[7].a/U4172  ( .A(\w1[7][103] ), .B(\w1[7][100] ), .Z(n14423)
         );
  XOR \SUBBYTES[7].a/U4171  ( .A(\w1[7][96] ), .B(\SUBBYTES[7].a/w905 ), .Z(
        \SUBBYTES[7].a/w784 ) );
  XOR \SUBBYTES[7].a/U4170  ( .A(n14425), .B(n14424), .Z(\SUBBYTES[7].a/w892 )
         );
  XOR \SUBBYTES[7].a/U4169  ( .A(\SUBBYTES[7].a/w853 ), .B(n1056), .Z(n14424)
         );
  XOR \SUBBYTES[7].a/U4168  ( .A(\SUBBYTES[7].a/w846 ), .B(
        \SUBBYTES[7].a/w849 ), .Z(n14425) );
  XOR \SUBBYTES[7].a/U4167  ( .A(n14427), .B(n14426), .Z(\SUBBYTES[7].a/w893 )
         );
  XOR \SUBBYTES[7].a/U4166  ( .A(\SUBBYTES[7].a/w853 ), .B(n13519), .Z(n14426)
         );
  XOR \SUBBYTES[7].a/U4165  ( .A(\SUBBYTES[7].a/w846 ), .B(n13518), .Z(n14427)
         );
  XOR \SUBBYTES[7].a/U4164  ( .A(\SUBBYTES[7].a/w905 ), .B(n14428), .Z(
        \SUBBYTES[7].a/w895 ) );
  XOR \SUBBYTES[7].a/U4163  ( .A(\w1[7][102] ), .B(\w1[7][101] ), .Z(n14428)
         );
  XOR \SUBBYTES[7].a/U4162  ( .A(n14430), .B(n14429), .Z(\SUBBYTES[7].a/w896 )
         );
  XOR \SUBBYTES[7].a/U4161  ( .A(n13519), .B(n1056), .Z(n14429) );
  XOR \SUBBYTES[7].a/U4160  ( .A(n13518), .B(\SUBBYTES[7].a/w849 ), .Z(n14430)
         );
  XOR \SUBBYTES[7].a/U4159  ( .A(\w1[7][103] ), .B(\w1[7][98] ), .Z(n14754) );
  XOR \SUBBYTES[7].a/U4158  ( .A(n14754), .B(n14431), .Z(\SUBBYTES[7].a/w897 )
         );
  XOR \SUBBYTES[7].a/U4157  ( .A(\w1[7][101] ), .B(\w1[7][100] ), .Z(n14431)
         );
  XOR \SUBBYTES[7].a/U4156  ( .A(\w1[7][103] ), .B(\SUBBYTES[7].a/w782 ), .Z(
        \SUBBYTES[7].a/w785 ) );
  XOR \SUBBYTES[7].a/U4155  ( .A(\w1[7][97] ), .B(\SUBBYTES[7].a/w782 ), .Z(
        \SUBBYTES[7].a/w786 ) );
  XOR \SUBBYTES[7].a/U4154  ( .A(\w1[7][100] ), .B(\SUBBYTES[7].a/w782 ), .Z(
        \SUBBYTES[7].a/w787 ) );
  XOR \SUBBYTES[7].a/U4153  ( .A(\SUBBYTES[7].a/w786 ), .B(n14754), .Z(
        \SUBBYTES[7].a/w788 ) );
  XOR \SUBBYTES[7].a/U4152  ( .A(n14754), .B(n14432), .Z(\SUBBYTES[7].a/w873 )
         );
  XOR \SUBBYTES[7].a/U4151  ( .A(\w1[7][100] ), .B(\w1[7][97] ), .Z(n14432) );
  XOR \SUBBYTES[7].a/U4150  ( .A(n14434), .B(n14433), .Z(n14751) );
  XOR \SUBBYTES[7].a/U4149  ( .A(\w1[7][100] ), .B(n14435), .Z(n14433) );
  XOR \SUBBYTES[7].a/U4148  ( .A(\SUBBYTES[7].a/w838 ), .B(\w1[7][102] ), .Z(
        n14434) );
  XOR \SUBBYTES[7].a/U4147  ( .A(\SUBBYTES[7].a/w812 ), .B(
        \SUBBYTES[7].a/w819 ), .Z(n14435) );
  XOR \SUBBYTES[7].a/U4146  ( .A(n14437), .B(n14436), .Z(n14749) );
  XOR \SUBBYTES[7].a/U4145  ( .A(\w1[7][97] ), .B(n14438), .Z(n14436) );
  XOR \SUBBYTES[7].a/U4144  ( .A(\SUBBYTES[7].a/w837 ), .B(\w1[7][101] ), .Z(
        n14437) );
  XOR \SUBBYTES[7].a/U4143  ( .A(\SUBBYTES[7].a/w813 ), .B(
        \SUBBYTES[7].a/w820 ), .Z(n14438) );
  XOR \SUBBYTES[7].a/U4142  ( .A(n14751), .B(n14749), .Z(\SUBBYTES[7].a/w843 )
         );
  XOR \SUBBYTES[7].a/U4141  ( .A(\w1[7][101] ), .B(n14439), .Z(n14752) );
  XOR \SUBBYTES[7].a/U4140  ( .A(\SUBBYTES[7].a/w805 ), .B(
        \SUBBYTES[7].a/w815 ), .Z(n14439) );
  XOR \SUBBYTES[7].a/U4139  ( .A(n14441), .B(n14440), .Z(\SUBBYTES[7].a/w830 )
         );
  XOR \SUBBYTES[7].a/U4138  ( .A(n14752), .B(n14442), .Z(n14440) );
  XOR \SUBBYTES[7].a/U4137  ( .A(\w1[7][100] ), .B(\SUBBYTES[7].a/w894 ), .Z(
        n14441) );
  XOR \SUBBYTES[7].a/U4136  ( .A(\SUBBYTES[7].a/w807 ), .B(
        \SUBBYTES[7].a/w812 ), .Z(n14442) );
  XOR \SUBBYTES[7].a/U4135  ( .A(n14444), .B(n14443), .Z(n14750) );
  XOR \SUBBYTES[7].a/U4134  ( .A(\SUBBYTES[7].a/w840 ), .B(\w1[7][103] ), .Z(
        n14443) );
  XOR \SUBBYTES[7].a/U4133  ( .A(\SUBBYTES[7].a/w815 ), .B(
        \SUBBYTES[7].a/w822 ), .Z(n14444) );
  XOR \SUBBYTES[7].a/U4132  ( .A(n14749), .B(n14750), .Z(\SUBBYTES[7].a/w842 )
         );
  XOR \SUBBYTES[7].a/U4131  ( .A(\w1[7][99] ), .B(n14445), .Z(n14753) );
  XOR \SUBBYTES[7].a/U4130  ( .A(\SUBBYTES[7].a/w804 ), .B(
        \SUBBYTES[7].a/w807 ), .Z(n14445) );
  XOR \SUBBYTES[7].a/U4129  ( .A(n14447), .B(n14446), .Z(\SUBBYTES[7].a/w831 )
         );
  XOR \SUBBYTES[7].a/U4128  ( .A(n14753), .B(n14448), .Z(n14446) );
  XOR \SUBBYTES[7].a/U4127  ( .A(\w1[7][102] ), .B(\SUBBYTES[7].a/w873 ), .Z(
        n14447) );
  XOR \SUBBYTES[7].a/U4126  ( .A(\SUBBYTES[7].a/w812 ), .B(
        \SUBBYTES[7].a/w813 ), .Z(n14448) );
  XOR \SUBBYTES[7].a/U4125  ( .A(n14751), .B(n14750), .Z(\SUBBYTES[7].a/w851 )
         );
  XOR \SUBBYTES[7].a/U4124  ( .A(n14450), .B(n14449), .Z(\SUBBYTES[7].a/w852 )
         );
  XOR \SUBBYTES[7].a/U4123  ( .A(\w1[7][103] ), .B(n14752), .Z(n14449) );
  XOR \SUBBYTES[7].a/U4122  ( .A(\SUBBYTES[7].a/w804 ), .B(
        \SUBBYTES[7].a/w813 ), .Z(n14450) );
  XOR \SUBBYTES[7].a/U4121  ( .A(n14452), .B(n14451), .Z(\SUBBYTES[7].a/w828 )
         );
  XOR \SUBBYTES[7].a/U4120  ( .A(n14454), .B(n14453), .Z(n14451) );
  XOR \SUBBYTES[7].a/U4119  ( .A(\w1[7][103] ), .B(\SUBBYTES[7].a/w912 ), .Z(
        n14452) );
  XOR \SUBBYTES[7].a/U4118  ( .A(\SUBBYTES[7].a/w819 ), .B(
        \SUBBYTES[7].a/w822 ), .Z(n14453) );
  XOR \SUBBYTES[7].a/U4117  ( .A(\SUBBYTES[7].a/w805 ), .B(
        \SUBBYTES[7].a/w807 ), .Z(n14454) );
  XOR \SUBBYTES[7].a/U4116  ( .A(n14456), .B(n14455), .Z(\SUBBYTES[7].a/w829 )
         );
  XOR \SUBBYTES[7].a/U4115  ( .A(n14753), .B(n14457), .Z(n14455) );
  XOR \SUBBYTES[7].a/U4114  ( .A(\w1[7][101] ), .B(n14754), .Z(n14456) );
  XOR \SUBBYTES[7].a/U4113  ( .A(\SUBBYTES[7].a/w819 ), .B(
        \SUBBYTES[7].a/w820 ), .Z(n14457) );
  XOR \SUBBYTES[7].a/U4112  ( .A(n14459), .B(n14458), .Z(\SUBBYTES[7].a/w845 )
         );
  XOR \SUBBYTES[7].a/U4111  ( .A(\w1[7][97] ), .B(n14460), .Z(n14458) );
  XOR \SUBBYTES[7].a/U4110  ( .A(\SUBBYTES[7].a/w820 ), .B(
        \SUBBYTES[7].a/w822 ), .Z(n14459) );
  XOR \SUBBYTES[7].a/U4109  ( .A(\SUBBYTES[7].a/w804 ), .B(
        \SUBBYTES[7].a/w805 ), .Z(n14460) );
  XOR \SUBBYTES[7].a/U4108  ( .A(\w1[7][105] ), .B(n14461), .Z(n14755) );
  XOR \SUBBYTES[7].a/U4107  ( .A(\w1[7][107] ), .B(\w1[7][106] ), .Z(n14461)
         );
  XOR \SUBBYTES[7].a/U4106  ( .A(\w1[7][110] ), .B(n14755), .Z(
        \SUBBYTES[7].a/w687 ) );
  XOR \SUBBYTES[7].a/U4105  ( .A(\w1[7][104] ), .B(\SUBBYTES[7].a/w687 ), .Z(
        \SUBBYTES[7].a/w574 ) );
  XOR \SUBBYTES[7].a/U4104  ( .A(\w1[7][104] ), .B(n14462), .Z(
        \SUBBYTES[7].a/w575 ) );
  XOR \SUBBYTES[7].a/U4103  ( .A(\w1[7][110] ), .B(\w1[7][109] ), .Z(n14462)
         );
  XOR \SUBBYTES[7].a/U4102  ( .A(\w1[7][109] ), .B(n14755), .Z(
        \SUBBYTES[7].a/w705 ) );
  XOR \SUBBYTES[7].a/U4101  ( .A(n14464), .B(n14463), .Z(\SUBBYTES[7].a/w698 )
         );
  XOR \SUBBYTES[7].a/U4100  ( .A(\w1[7][107] ), .B(\w1[7][105] ), .Z(n14463)
         );
  XOR \SUBBYTES[7].a/U4099  ( .A(\w1[7][111] ), .B(\w1[7][108] ), .Z(n14464)
         );
  XOR \SUBBYTES[7].a/U4098  ( .A(\w1[7][104] ), .B(\SUBBYTES[7].a/w698 ), .Z(
        \SUBBYTES[7].a/w577 ) );
  XOR \SUBBYTES[7].a/U4097  ( .A(n14466), .B(n14465), .Z(\SUBBYTES[7].a/w685 )
         );
  XOR \SUBBYTES[7].a/U4096  ( .A(\SUBBYTES[7].a/w646 ), .B(n1055), .Z(n14465)
         );
  XOR \SUBBYTES[7].a/U4095  ( .A(\SUBBYTES[7].a/w639 ), .B(
        \SUBBYTES[7].a/w642 ), .Z(n14466) );
  XOR \SUBBYTES[7].a/U4094  ( .A(n14468), .B(n14467), .Z(\SUBBYTES[7].a/w686 )
         );
  XOR \SUBBYTES[7].a/U4093  ( .A(\SUBBYTES[7].a/w646 ), .B(n13517), .Z(n14467)
         );
  XOR \SUBBYTES[7].a/U4092  ( .A(\SUBBYTES[7].a/w639 ), .B(n13516), .Z(n14468)
         );
  XOR \SUBBYTES[7].a/U4091  ( .A(\SUBBYTES[7].a/w698 ), .B(n14469), .Z(
        \SUBBYTES[7].a/w688 ) );
  XOR \SUBBYTES[7].a/U4090  ( .A(\w1[7][110] ), .B(\w1[7][109] ), .Z(n14469)
         );
  XOR \SUBBYTES[7].a/U4089  ( .A(n14471), .B(n14470), .Z(\SUBBYTES[7].a/w689 )
         );
  XOR \SUBBYTES[7].a/U4088  ( .A(n13517), .B(n1055), .Z(n14470) );
  XOR \SUBBYTES[7].a/U4087  ( .A(n13516), .B(\SUBBYTES[7].a/w642 ), .Z(n14471)
         );
  XOR \SUBBYTES[7].a/U4086  ( .A(\w1[7][111] ), .B(\w1[7][106] ), .Z(n14761)
         );
  XOR \SUBBYTES[7].a/U4085  ( .A(n14761), .B(n14472), .Z(\SUBBYTES[7].a/w690 )
         );
  XOR \SUBBYTES[7].a/U4084  ( .A(\w1[7][109] ), .B(\w1[7][108] ), .Z(n14472)
         );
  XOR \SUBBYTES[7].a/U4083  ( .A(\w1[7][111] ), .B(\SUBBYTES[7].a/w575 ), .Z(
        \SUBBYTES[7].a/w578 ) );
  XOR \SUBBYTES[7].a/U4082  ( .A(\w1[7][105] ), .B(\SUBBYTES[7].a/w575 ), .Z(
        \SUBBYTES[7].a/w579 ) );
  XOR \SUBBYTES[7].a/U4081  ( .A(\w1[7][108] ), .B(\SUBBYTES[7].a/w575 ), .Z(
        \SUBBYTES[7].a/w580 ) );
  XOR \SUBBYTES[7].a/U4080  ( .A(\SUBBYTES[7].a/w579 ), .B(n14761), .Z(
        \SUBBYTES[7].a/w581 ) );
  XOR \SUBBYTES[7].a/U4079  ( .A(n14761), .B(n14473), .Z(\SUBBYTES[7].a/w666 )
         );
  XOR \SUBBYTES[7].a/U4078  ( .A(\w1[7][108] ), .B(\w1[7][105] ), .Z(n14473)
         );
  XOR \SUBBYTES[7].a/U4077  ( .A(n14475), .B(n14474), .Z(n14758) );
  XOR \SUBBYTES[7].a/U4076  ( .A(\w1[7][108] ), .B(n14476), .Z(n14474) );
  XOR \SUBBYTES[7].a/U4075  ( .A(\SUBBYTES[7].a/w631 ), .B(\w1[7][110] ), .Z(
        n14475) );
  XOR \SUBBYTES[7].a/U4074  ( .A(\SUBBYTES[7].a/w605 ), .B(
        \SUBBYTES[7].a/w612 ), .Z(n14476) );
  XOR \SUBBYTES[7].a/U4073  ( .A(n14478), .B(n14477), .Z(n14756) );
  XOR \SUBBYTES[7].a/U4072  ( .A(\w1[7][105] ), .B(n14479), .Z(n14477) );
  XOR \SUBBYTES[7].a/U4071  ( .A(\SUBBYTES[7].a/w630 ), .B(\w1[7][109] ), .Z(
        n14478) );
  XOR \SUBBYTES[7].a/U4070  ( .A(\SUBBYTES[7].a/w606 ), .B(
        \SUBBYTES[7].a/w613 ), .Z(n14479) );
  XOR \SUBBYTES[7].a/U4069  ( .A(n14758), .B(n14756), .Z(\SUBBYTES[7].a/w636 )
         );
  XOR \SUBBYTES[7].a/U4068  ( .A(\w1[7][109] ), .B(n14480), .Z(n14759) );
  XOR \SUBBYTES[7].a/U4067  ( .A(\SUBBYTES[7].a/w598 ), .B(
        \SUBBYTES[7].a/w608 ), .Z(n14480) );
  XOR \SUBBYTES[7].a/U4066  ( .A(n14482), .B(n14481), .Z(\SUBBYTES[7].a/w623 )
         );
  XOR \SUBBYTES[7].a/U4065  ( .A(n14759), .B(n14483), .Z(n14481) );
  XOR \SUBBYTES[7].a/U4064  ( .A(\w1[7][108] ), .B(\SUBBYTES[7].a/w687 ), .Z(
        n14482) );
  XOR \SUBBYTES[7].a/U4063  ( .A(\SUBBYTES[7].a/w600 ), .B(
        \SUBBYTES[7].a/w605 ), .Z(n14483) );
  XOR \SUBBYTES[7].a/U4062  ( .A(n14485), .B(n14484), .Z(n14757) );
  XOR \SUBBYTES[7].a/U4061  ( .A(\SUBBYTES[7].a/w633 ), .B(\w1[7][111] ), .Z(
        n14484) );
  XOR \SUBBYTES[7].a/U4060  ( .A(\SUBBYTES[7].a/w608 ), .B(
        \SUBBYTES[7].a/w615 ), .Z(n14485) );
  XOR \SUBBYTES[7].a/U4059  ( .A(n14756), .B(n14757), .Z(\SUBBYTES[7].a/w635 )
         );
  XOR \SUBBYTES[7].a/U4058  ( .A(\w1[7][107] ), .B(n14486), .Z(n14760) );
  XOR \SUBBYTES[7].a/U4057  ( .A(\SUBBYTES[7].a/w597 ), .B(
        \SUBBYTES[7].a/w600 ), .Z(n14486) );
  XOR \SUBBYTES[7].a/U4056  ( .A(n14488), .B(n14487), .Z(\SUBBYTES[7].a/w624 )
         );
  XOR \SUBBYTES[7].a/U4055  ( .A(n14760), .B(n14489), .Z(n14487) );
  XOR \SUBBYTES[7].a/U4054  ( .A(\w1[7][110] ), .B(\SUBBYTES[7].a/w666 ), .Z(
        n14488) );
  XOR \SUBBYTES[7].a/U4053  ( .A(\SUBBYTES[7].a/w605 ), .B(
        \SUBBYTES[7].a/w606 ), .Z(n14489) );
  XOR \SUBBYTES[7].a/U4052  ( .A(n14758), .B(n14757), .Z(\SUBBYTES[7].a/w644 )
         );
  XOR \SUBBYTES[7].a/U4051  ( .A(n14491), .B(n14490), .Z(\SUBBYTES[7].a/w645 )
         );
  XOR \SUBBYTES[7].a/U4050  ( .A(\w1[7][111] ), .B(n14759), .Z(n14490) );
  XOR \SUBBYTES[7].a/U4049  ( .A(\SUBBYTES[7].a/w597 ), .B(
        \SUBBYTES[7].a/w606 ), .Z(n14491) );
  XOR \SUBBYTES[7].a/U4048  ( .A(n14493), .B(n14492), .Z(\SUBBYTES[7].a/w621 )
         );
  XOR \SUBBYTES[7].a/U4047  ( .A(n14495), .B(n14494), .Z(n14492) );
  XOR \SUBBYTES[7].a/U4046  ( .A(\w1[7][111] ), .B(\SUBBYTES[7].a/w705 ), .Z(
        n14493) );
  XOR \SUBBYTES[7].a/U4045  ( .A(\SUBBYTES[7].a/w612 ), .B(
        \SUBBYTES[7].a/w615 ), .Z(n14494) );
  XOR \SUBBYTES[7].a/U4044  ( .A(\SUBBYTES[7].a/w598 ), .B(
        \SUBBYTES[7].a/w600 ), .Z(n14495) );
  XOR \SUBBYTES[7].a/U4043  ( .A(n14497), .B(n14496), .Z(\SUBBYTES[7].a/w622 )
         );
  XOR \SUBBYTES[7].a/U4042  ( .A(n14760), .B(n14498), .Z(n14496) );
  XOR \SUBBYTES[7].a/U4041  ( .A(\w1[7][109] ), .B(n14761), .Z(n14497) );
  XOR \SUBBYTES[7].a/U4040  ( .A(\SUBBYTES[7].a/w612 ), .B(
        \SUBBYTES[7].a/w613 ), .Z(n14498) );
  XOR \SUBBYTES[7].a/U4039  ( .A(n14500), .B(n14499), .Z(\SUBBYTES[7].a/w638 )
         );
  XOR \SUBBYTES[7].a/U4038  ( .A(\w1[7][105] ), .B(n14501), .Z(n14499) );
  XOR \SUBBYTES[7].a/U4037  ( .A(\SUBBYTES[7].a/w613 ), .B(
        \SUBBYTES[7].a/w615 ), .Z(n14500) );
  XOR \SUBBYTES[7].a/U4036  ( .A(\SUBBYTES[7].a/w597 ), .B(
        \SUBBYTES[7].a/w598 ), .Z(n14501) );
  XOR \SUBBYTES[7].a/U4035  ( .A(\w1[7][113] ), .B(n14502), .Z(n14762) );
  XOR \SUBBYTES[7].a/U4034  ( .A(\w1[7][115] ), .B(\w1[7][114] ), .Z(n14502)
         );
  XOR \SUBBYTES[7].a/U4033  ( .A(\w1[7][118] ), .B(n14762), .Z(
        \SUBBYTES[7].a/w480 ) );
  XOR \SUBBYTES[7].a/U4032  ( .A(\w1[7][112] ), .B(\SUBBYTES[7].a/w480 ), .Z(
        \SUBBYTES[7].a/w367 ) );
  XOR \SUBBYTES[7].a/U4031  ( .A(\w1[7][112] ), .B(n14503), .Z(
        \SUBBYTES[7].a/w368 ) );
  XOR \SUBBYTES[7].a/U4030  ( .A(\w1[7][118] ), .B(\w1[7][117] ), .Z(n14503)
         );
  XOR \SUBBYTES[7].a/U4029  ( .A(\w1[7][117] ), .B(n14762), .Z(
        \SUBBYTES[7].a/w498 ) );
  XOR \SUBBYTES[7].a/U4028  ( .A(n14505), .B(n14504), .Z(\SUBBYTES[7].a/w491 )
         );
  XOR \SUBBYTES[7].a/U4027  ( .A(\w1[7][115] ), .B(\w1[7][113] ), .Z(n14504)
         );
  XOR \SUBBYTES[7].a/U4026  ( .A(\w1[7][119] ), .B(\w1[7][116] ), .Z(n14505)
         );
  XOR \SUBBYTES[7].a/U4025  ( .A(\w1[7][112] ), .B(\SUBBYTES[7].a/w491 ), .Z(
        \SUBBYTES[7].a/w370 ) );
  XOR \SUBBYTES[7].a/U4024  ( .A(n14507), .B(n14506), .Z(\SUBBYTES[7].a/w478 )
         );
  XOR \SUBBYTES[7].a/U4023  ( .A(\SUBBYTES[7].a/w439 ), .B(n1054), .Z(n14506)
         );
  XOR \SUBBYTES[7].a/U4022  ( .A(\SUBBYTES[7].a/w432 ), .B(
        \SUBBYTES[7].a/w435 ), .Z(n14507) );
  XOR \SUBBYTES[7].a/U4021  ( .A(n14509), .B(n14508), .Z(\SUBBYTES[7].a/w479 )
         );
  XOR \SUBBYTES[7].a/U4020  ( .A(\SUBBYTES[7].a/w439 ), .B(n13515), .Z(n14508)
         );
  XOR \SUBBYTES[7].a/U4019  ( .A(\SUBBYTES[7].a/w432 ), .B(n13514), .Z(n14509)
         );
  XOR \SUBBYTES[7].a/U4018  ( .A(\SUBBYTES[7].a/w491 ), .B(n14510), .Z(
        \SUBBYTES[7].a/w481 ) );
  XOR \SUBBYTES[7].a/U4017  ( .A(\w1[7][118] ), .B(\w1[7][117] ), .Z(n14510)
         );
  XOR \SUBBYTES[7].a/U4016  ( .A(n14512), .B(n14511), .Z(\SUBBYTES[7].a/w482 )
         );
  XOR \SUBBYTES[7].a/U4015  ( .A(n13515), .B(n1054), .Z(n14511) );
  XOR \SUBBYTES[7].a/U4014  ( .A(n13514), .B(\SUBBYTES[7].a/w435 ), .Z(n14512)
         );
  XOR \SUBBYTES[7].a/U4013  ( .A(\w1[7][119] ), .B(\w1[7][114] ), .Z(n14768)
         );
  XOR \SUBBYTES[7].a/U4012  ( .A(n14768), .B(n14513), .Z(\SUBBYTES[7].a/w483 )
         );
  XOR \SUBBYTES[7].a/U4011  ( .A(\w1[7][117] ), .B(\w1[7][116] ), .Z(n14513)
         );
  XOR \SUBBYTES[7].a/U4010  ( .A(\w1[7][119] ), .B(\SUBBYTES[7].a/w368 ), .Z(
        \SUBBYTES[7].a/w371 ) );
  XOR \SUBBYTES[7].a/U4009  ( .A(\w1[7][113] ), .B(\SUBBYTES[7].a/w368 ), .Z(
        \SUBBYTES[7].a/w372 ) );
  XOR \SUBBYTES[7].a/U4008  ( .A(\w1[7][116] ), .B(\SUBBYTES[7].a/w368 ), .Z(
        \SUBBYTES[7].a/w373 ) );
  XOR \SUBBYTES[7].a/U4007  ( .A(\SUBBYTES[7].a/w372 ), .B(n14768), .Z(
        \SUBBYTES[7].a/w374 ) );
  XOR \SUBBYTES[7].a/U4006  ( .A(n14768), .B(n14514), .Z(\SUBBYTES[7].a/w459 )
         );
  XOR \SUBBYTES[7].a/U4005  ( .A(\w1[7][116] ), .B(\w1[7][113] ), .Z(n14514)
         );
  XOR \SUBBYTES[7].a/U4004  ( .A(n14516), .B(n14515), .Z(n14765) );
  XOR \SUBBYTES[7].a/U4003  ( .A(\w1[7][116] ), .B(n14517), .Z(n14515) );
  XOR \SUBBYTES[7].a/U4002  ( .A(\SUBBYTES[7].a/w424 ), .B(\w1[7][118] ), .Z(
        n14516) );
  XOR \SUBBYTES[7].a/U4001  ( .A(\SUBBYTES[7].a/w398 ), .B(
        \SUBBYTES[7].a/w405 ), .Z(n14517) );
  XOR \SUBBYTES[7].a/U4000  ( .A(n14519), .B(n14518), .Z(n14763) );
  XOR \SUBBYTES[7].a/U3999  ( .A(\w1[7][113] ), .B(n14520), .Z(n14518) );
  XOR \SUBBYTES[7].a/U3998  ( .A(\SUBBYTES[7].a/w423 ), .B(\w1[7][117] ), .Z(
        n14519) );
  XOR \SUBBYTES[7].a/U3997  ( .A(\SUBBYTES[7].a/w399 ), .B(
        \SUBBYTES[7].a/w406 ), .Z(n14520) );
  XOR \SUBBYTES[7].a/U3996  ( .A(n14765), .B(n14763), .Z(\SUBBYTES[7].a/w429 )
         );
  XOR \SUBBYTES[7].a/U3995  ( .A(\w1[7][117] ), .B(n14521), .Z(n14766) );
  XOR \SUBBYTES[7].a/U3994  ( .A(\SUBBYTES[7].a/w391 ), .B(
        \SUBBYTES[7].a/w401 ), .Z(n14521) );
  XOR \SUBBYTES[7].a/U3993  ( .A(n14523), .B(n14522), .Z(\SUBBYTES[7].a/w416 )
         );
  XOR \SUBBYTES[7].a/U3992  ( .A(n14766), .B(n14524), .Z(n14522) );
  XOR \SUBBYTES[7].a/U3991  ( .A(\w1[7][116] ), .B(\SUBBYTES[7].a/w480 ), .Z(
        n14523) );
  XOR \SUBBYTES[7].a/U3990  ( .A(\SUBBYTES[7].a/w393 ), .B(
        \SUBBYTES[7].a/w398 ), .Z(n14524) );
  XOR \SUBBYTES[7].a/U3989  ( .A(n14526), .B(n14525), .Z(n14764) );
  XOR \SUBBYTES[7].a/U3988  ( .A(\SUBBYTES[7].a/w426 ), .B(\w1[7][119] ), .Z(
        n14525) );
  XOR \SUBBYTES[7].a/U3987  ( .A(\SUBBYTES[7].a/w401 ), .B(
        \SUBBYTES[7].a/w408 ), .Z(n14526) );
  XOR \SUBBYTES[7].a/U3986  ( .A(n14763), .B(n14764), .Z(\SUBBYTES[7].a/w428 )
         );
  XOR \SUBBYTES[7].a/U3985  ( .A(\w1[7][115] ), .B(n14527), .Z(n14767) );
  XOR \SUBBYTES[7].a/U3984  ( .A(\SUBBYTES[7].a/w390 ), .B(
        \SUBBYTES[7].a/w393 ), .Z(n14527) );
  XOR \SUBBYTES[7].a/U3983  ( .A(n14529), .B(n14528), .Z(\SUBBYTES[7].a/w417 )
         );
  XOR \SUBBYTES[7].a/U3982  ( .A(n14767), .B(n14530), .Z(n14528) );
  XOR \SUBBYTES[7].a/U3981  ( .A(\w1[7][118] ), .B(\SUBBYTES[7].a/w459 ), .Z(
        n14529) );
  XOR \SUBBYTES[7].a/U3980  ( .A(\SUBBYTES[7].a/w398 ), .B(
        \SUBBYTES[7].a/w399 ), .Z(n14530) );
  XOR \SUBBYTES[7].a/U3979  ( .A(n14765), .B(n14764), .Z(\SUBBYTES[7].a/w437 )
         );
  XOR \SUBBYTES[7].a/U3978  ( .A(n14532), .B(n14531), .Z(\SUBBYTES[7].a/w438 )
         );
  XOR \SUBBYTES[7].a/U3977  ( .A(\w1[7][119] ), .B(n14766), .Z(n14531) );
  XOR \SUBBYTES[7].a/U3976  ( .A(\SUBBYTES[7].a/w390 ), .B(
        \SUBBYTES[7].a/w399 ), .Z(n14532) );
  XOR \SUBBYTES[7].a/U3975  ( .A(n14534), .B(n14533), .Z(\SUBBYTES[7].a/w414 )
         );
  XOR \SUBBYTES[7].a/U3974  ( .A(n14536), .B(n14535), .Z(n14533) );
  XOR \SUBBYTES[7].a/U3973  ( .A(\w1[7][119] ), .B(\SUBBYTES[7].a/w498 ), .Z(
        n14534) );
  XOR \SUBBYTES[7].a/U3972  ( .A(\SUBBYTES[7].a/w405 ), .B(
        \SUBBYTES[7].a/w408 ), .Z(n14535) );
  XOR \SUBBYTES[7].a/U3971  ( .A(\SUBBYTES[7].a/w391 ), .B(
        \SUBBYTES[7].a/w393 ), .Z(n14536) );
  XOR \SUBBYTES[7].a/U3970  ( .A(n14538), .B(n14537), .Z(\SUBBYTES[7].a/w415 )
         );
  XOR \SUBBYTES[7].a/U3969  ( .A(n14767), .B(n14539), .Z(n14537) );
  XOR \SUBBYTES[7].a/U3968  ( .A(\w1[7][117] ), .B(n14768), .Z(n14538) );
  XOR \SUBBYTES[7].a/U3967  ( .A(\SUBBYTES[7].a/w405 ), .B(
        \SUBBYTES[7].a/w406 ), .Z(n14539) );
  XOR \SUBBYTES[7].a/U3966  ( .A(n14541), .B(n14540), .Z(\SUBBYTES[7].a/w431 )
         );
  XOR \SUBBYTES[7].a/U3965  ( .A(\w1[7][113] ), .B(n14542), .Z(n14540) );
  XOR \SUBBYTES[7].a/U3964  ( .A(\SUBBYTES[7].a/w406 ), .B(
        \SUBBYTES[7].a/w408 ), .Z(n14541) );
  XOR \SUBBYTES[7].a/U3963  ( .A(\SUBBYTES[7].a/w390 ), .B(
        \SUBBYTES[7].a/w391 ), .Z(n14542) );
  XOR \SUBBYTES[7].a/U3962  ( .A(\w1[7][121] ), .B(n14543), .Z(n14769) );
  XOR \SUBBYTES[7].a/U3961  ( .A(\w1[7][123] ), .B(\w1[7][122] ), .Z(n14543)
         );
  XOR \SUBBYTES[7].a/U3960  ( .A(\w1[7][126] ), .B(n14769), .Z(
        \SUBBYTES[7].a/w273 ) );
  XOR \SUBBYTES[7].a/U3959  ( .A(\w1[7][120] ), .B(\SUBBYTES[7].a/w273 ), .Z(
        \SUBBYTES[7].a/w160 ) );
  XOR \SUBBYTES[7].a/U3958  ( .A(\w1[7][120] ), .B(n14544), .Z(
        \SUBBYTES[7].a/w161 ) );
  XOR \SUBBYTES[7].a/U3957  ( .A(\w1[7][126] ), .B(\w1[7][125] ), .Z(n14544)
         );
  XOR \SUBBYTES[7].a/U3956  ( .A(\w1[7][125] ), .B(n14769), .Z(
        \SUBBYTES[7].a/w291 ) );
  XOR \SUBBYTES[7].a/U3955  ( .A(n14546), .B(n14545), .Z(\SUBBYTES[7].a/w284 )
         );
  XOR \SUBBYTES[7].a/U3954  ( .A(\w1[7][123] ), .B(\w1[7][121] ), .Z(n14545)
         );
  XOR \SUBBYTES[7].a/U3953  ( .A(\w1[7][127] ), .B(\w1[7][124] ), .Z(n14546)
         );
  XOR \SUBBYTES[7].a/U3952  ( .A(\w1[7][120] ), .B(\SUBBYTES[7].a/w284 ), .Z(
        \SUBBYTES[7].a/w163 ) );
  XOR \SUBBYTES[7].a/U3951  ( .A(n14548), .B(n14547), .Z(\SUBBYTES[7].a/w271 )
         );
  XOR \SUBBYTES[7].a/U3950  ( .A(\SUBBYTES[7].a/w232 ), .B(n1053), .Z(n14547)
         );
  XOR \SUBBYTES[7].a/U3949  ( .A(\SUBBYTES[7].a/w225 ), .B(
        \SUBBYTES[7].a/w228 ), .Z(n14548) );
  XOR \SUBBYTES[7].a/U3948  ( .A(n14550), .B(n14549), .Z(\SUBBYTES[7].a/w272 )
         );
  XOR \SUBBYTES[7].a/U3947  ( .A(\SUBBYTES[7].a/w232 ), .B(n13513), .Z(n14549)
         );
  XOR \SUBBYTES[7].a/U3946  ( .A(\SUBBYTES[7].a/w225 ), .B(n13512), .Z(n14550)
         );
  XOR \SUBBYTES[7].a/U3945  ( .A(\SUBBYTES[7].a/w284 ), .B(n14551), .Z(
        \SUBBYTES[7].a/w274 ) );
  XOR \SUBBYTES[7].a/U3944  ( .A(\w1[7][126] ), .B(\w1[7][125] ), .Z(n14551)
         );
  XOR \SUBBYTES[7].a/U3943  ( .A(n14553), .B(n14552), .Z(\SUBBYTES[7].a/w275 )
         );
  XOR \SUBBYTES[7].a/U3942  ( .A(n13513), .B(n1053), .Z(n14552) );
  XOR \SUBBYTES[7].a/U3941  ( .A(n13512), .B(\SUBBYTES[7].a/w228 ), .Z(n14553)
         );
  XOR \SUBBYTES[7].a/U3940  ( .A(\w1[7][127] ), .B(\w1[7][122] ), .Z(n14775)
         );
  XOR \SUBBYTES[7].a/U3939  ( .A(n14775), .B(n14554), .Z(\SUBBYTES[7].a/w276 )
         );
  XOR \SUBBYTES[7].a/U3938  ( .A(\w1[7][125] ), .B(\w1[7][124] ), .Z(n14554)
         );
  XOR \SUBBYTES[7].a/U3937  ( .A(\w1[7][127] ), .B(\SUBBYTES[7].a/w161 ), .Z(
        \SUBBYTES[7].a/w164 ) );
  XOR \SUBBYTES[7].a/U3936  ( .A(\w1[7][121] ), .B(\SUBBYTES[7].a/w161 ), .Z(
        \SUBBYTES[7].a/w165 ) );
  XOR \SUBBYTES[7].a/U3935  ( .A(\w1[7][124] ), .B(\SUBBYTES[7].a/w161 ), .Z(
        \SUBBYTES[7].a/w166 ) );
  XOR \SUBBYTES[7].a/U3934  ( .A(\SUBBYTES[7].a/w165 ), .B(n14775), .Z(
        \SUBBYTES[7].a/w167 ) );
  XOR \SUBBYTES[7].a/U3933  ( .A(n14775), .B(n14555), .Z(\SUBBYTES[7].a/w252 )
         );
  XOR \SUBBYTES[7].a/U3932  ( .A(\w1[7][124] ), .B(\w1[7][121] ), .Z(n14555)
         );
  XOR \SUBBYTES[7].a/U3931  ( .A(n14557), .B(n14556), .Z(n14772) );
  XOR \SUBBYTES[7].a/U3930  ( .A(\w1[7][124] ), .B(n14558), .Z(n14556) );
  XOR \SUBBYTES[7].a/U3929  ( .A(\SUBBYTES[7].a/w217 ), .B(\w1[7][126] ), .Z(
        n14557) );
  XOR \SUBBYTES[7].a/U3928  ( .A(\SUBBYTES[7].a/w191 ), .B(
        \SUBBYTES[7].a/w198 ), .Z(n14558) );
  XOR \SUBBYTES[7].a/U3927  ( .A(n14560), .B(n14559), .Z(n14770) );
  XOR \SUBBYTES[7].a/U3926  ( .A(\w1[7][121] ), .B(n14561), .Z(n14559) );
  XOR \SUBBYTES[7].a/U3925  ( .A(\SUBBYTES[7].a/w216 ), .B(\w1[7][125] ), .Z(
        n14560) );
  XOR \SUBBYTES[7].a/U3924  ( .A(\SUBBYTES[7].a/w192 ), .B(
        \SUBBYTES[7].a/w199 ), .Z(n14561) );
  XOR \SUBBYTES[7].a/U3923  ( .A(n14772), .B(n14770), .Z(\SUBBYTES[7].a/w222 )
         );
  XOR \SUBBYTES[7].a/U3922  ( .A(\w1[7][125] ), .B(n14562), .Z(n14773) );
  XOR \SUBBYTES[7].a/U3921  ( .A(\SUBBYTES[7].a/w184 ), .B(
        \SUBBYTES[7].a/w194 ), .Z(n14562) );
  XOR \SUBBYTES[7].a/U3920  ( .A(n14564), .B(n14563), .Z(\SUBBYTES[7].a/w209 )
         );
  XOR \SUBBYTES[7].a/U3919  ( .A(n14773), .B(n14565), .Z(n14563) );
  XOR \SUBBYTES[7].a/U3918  ( .A(\w1[7][124] ), .B(\SUBBYTES[7].a/w273 ), .Z(
        n14564) );
  XOR \SUBBYTES[7].a/U3917  ( .A(\SUBBYTES[7].a/w186 ), .B(
        \SUBBYTES[7].a/w191 ), .Z(n14565) );
  XOR \SUBBYTES[7].a/U3916  ( .A(n14567), .B(n14566), .Z(n14771) );
  XOR \SUBBYTES[7].a/U3915  ( .A(\SUBBYTES[7].a/w219 ), .B(\w1[7][127] ), .Z(
        n14566) );
  XOR \SUBBYTES[7].a/U3914  ( .A(\SUBBYTES[7].a/w194 ), .B(
        \SUBBYTES[7].a/w201 ), .Z(n14567) );
  XOR \SUBBYTES[7].a/U3913  ( .A(n14770), .B(n14771), .Z(\SUBBYTES[7].a/w221 )
         );
  XOR \SUBBYTES[7].a/U3912  ( .A(\w1[7][123] ), .B(n14568), .Z(n14774) );
  XOR \SUBBYTES[7].a/U3911  ( .A(\SUBBYTES[7].a/w183 ), .B(
        \SUBBYTES[7].a/w186 ), .Z(n14568) );
  XOR \SUBBYTES[7].a/U3910  ( .A(n14570), .B(n14569), .Z(\SUBBYTES[7].a/w210 )
         );
  XOR \SUBBYTES[7].a/U3909  ( .A(n14774), .B(n14571), .Z(n14569) );
  XOR \SUBBYTES[7].a/U3908  ( .A(\w1[7][126] ), .B(\SUBBYTES[7].a/w252 ), .Z(
        n14570) );
  XOR \SUBBYTES[7].a/U3907  ( .A(\SUBBYTES[7].a/w191 ), .B(
        \SUBBYTES[7].a/w192 ), .Z(n14571) );
  XOR \SUBBYTES[7].a/U3906  ( .A(n14772), .B(n14771), .Z(\SUBBYTES[7].a/w230 )
         );
  XOR \SUBBYTES[7].a/U3905  ( .A(n14573), .B(n14572), .Z(\SUBBYTES[7].a/w231 )
         );
  XOR \SUBBYTES[7].a/U3904  ( .A(\w1[7][127] ), .B(n14773), .Z(n14572) );
  XOR \SUBBYTES[7].a/U3903  ( .A(\SUBBYTES[7].a/w183 ), .B(
        \SUBBYTES[7].a/w192 ), .Z(n14573) );
  XOR \SUBBYTES[7].a/U3902  ( .A(n14575), .B(n14574), .Z(\SUBBYTES[7].a/w207 )
         );
  XOR \SUBBYTES[7].a/U3901  ( .A(n14577), .B(n14576), .Z(n14574) );
  XOR \SUBBYTES[7].a/U3900  ( .A(\w1[7][127] ), .B(\SUBBYTES[7].a/w291 ), .Z(
        n14575) );
  XOR \SUBBYTES[7].a/U3899  ( .A(\SUBBYTES[7].a/w198 ), .B(
        \SUBBYTES[7].a/w201 ), .Z(n14576) );
  XOR \SUBBYTES[7].a/U3898  ( .A(\SUBBYTES[7].a/w184 ), .B(
        \SUBBYTES[7].a/w186 ), .Z(n14577) );
  XOR \SUBBYTES[7].a/U3897  ( .A(n14579), .B(n14578), .Z(\SUBBYTES[7].a/w208 )
         );
  XOR \SUBBYTES[7].a/U3896  ( .A(n14774), .B(n14580), .Z(n14578) );
  XOR \SUBBYTES[7].a/U3895  ( .A(\w1[7][125] ), .B(n14775), .Z(n14579) );
  XOR \SUBBYTES[7].a/U3894  ( .A(\SUBBYTES[7].a/w198 ), .B(
        \SUBBYTES[7].a/w199 ), .Z(n14580) );
  XOR \SUBBYTES[7].a/U3893  ( .A(n14582), .B(n14581), .Z(\SUBBYTES[7].a/w224 )
         );
  XOR \SUBBYTES[7].a/U3892  ( .A(\w1[7][121] ), .B(n14583), .Z(n14581) );
  XOR \SUBBYTES[7].a/U3891  ( .A(\SUBBYTES[7].a/w199 ), .B(
        \SUBBYTES[7].a/w201 ), .Z(n14582) );
  XOR \SUBBYTES[7].a/U3890  ( .A(\SUBBYTES[7].a/w183 ), .B(
        \SUBBYTES[7].a/w184 ), .Z(n14583) );
  XOR \SUBBYTES[6].a/U5649  ( .A(\SUBBYTES[6].a/w3390 ), .B(
        \SUBBYTES[6].a/w3391 ), .Z(n13305) );
  XOR \SUBBYTES[6].a/U5648  ( .A(n13305), .B(n12264), .Z(n13304) );
  XOR \SUBBYTES[6].a/U5647  ( .A(\SUBBYTES[6].a/w3383 ), .B(
        \SUBBYTES[6].a/w3400 ), .Z(n12264) );
  XOR \SUBBYTES[6].a/U5645  ( .A(\SUBBYTES[6].a/w3382 ), .B(
        \SUBBYTES[6].a/w3397 ), .Z(n12265) );
  XOR \SUBBYTES[6].a/U5644  ( .A(n13305), .B(n12266), .Z(n13496) );
  XOR \SUBBYTES[6].a/U5643  ( .A(\SUBBYTES[6].a/w3397 ), .B(
        \SUBBYTES[6].a/w3398 ), .Z(n12266) );
  XOR \SUBBYTES[6].a/U5642  ( .A(\SUBBYTES[6].a/w3359 ), .B(n12267), .Z(n13307) );
  XOR \SUBBYTES[6].a/U5641  ( .A(\SUBBYTES[6].a/w3350 ), .B(
        \SUBBYTES[6].a/w3351 ), .Z(n12267) );
  XOR \SUBBYTES[6].a/U5639  ( .A(\SUBBYTES[6].a/w3361 ), .B(n13496), .Z(n12268) );
  XOR \SUBBYTES[6].a/U5638  ( .A(n12270), .B(n12269), .Z(n13308) );
  XOR \SUBBYTES[6].a/U5637  ( .A(n12272), .B(n12271), .Z(n12269) );
  XOR \SUBBYTES[6].a/U5636  ( .A(\SUBBYTES[6].a/w3397 ), .B(
        \SUBBYTES[6].a/w3398 ), .Z(n12270) );
  XOR \SUBBYTES[6].a/U5635  ( .A(\SUBBYTES[6].a/w3361 ), .B(
        \SUBBYTES[6].a/w3385 ), .Z(n12271) );
  XOR \SUBBYTES[6].a/U5634  ( .A(\SUBBYTES[6].a/w3350 ), .B(
        \SUBBYTES[6].a/w3359 ), .Z(n12272) );
  XOR \SUBBYTES[6].a/U5633  ( .A(\SUBBYTES[6].a/w3382 ), .B(n12273), .Z(n13306) );
  XOR \SUBBYTES[6].a/U5632  ( .A(\SUBBYTES[6].a/w3365 ), .B(
        \SUBBYTES[6].a/w3368 ), .Z(n12273) );
  XOR \SUBBYTES[6].a/U5630  ( .A(\SUBBYTES[6].a/w3353 ), .B(n13308), .Z(n12274) );
  XOR \SUBBYTES[6].a/U5628  ( .A(\SUBBYTES[6].a/w3385 ), .B(
        \SUBBYTES[6].a/w3398 ), .Z(n12275) );
  XOR \SUBBYTES[6].a/U5626  ( .A(n12279), .B(n12278), .Z(n12276) );
  XOR \SUBBYTES[6].a/U5625  ( .A(n12281), .B(n12280), .Z(n12277) );
  XOR \SUBBYTES[6].a/U5624  ( .A(\SUBBYTES[6].a/w3397 ), .B(
        \SUBBYTES[6].a/w3400 ), .Z(n12278) );
  XOR \SUBBYTES[6].a/U5623  ( .A(\SUBBYTES[6].a/w3390 ), .B(
        \SUBBYTES[6].a/w3393 ), .Z(n12279) );
  XOR \SUBBYTES[6].a/U5622  ( .A(\SUBBYTES[6].a/w3365 ), .B(
        \SUBBYTES[6].a/w3366 ), .Z(n12280) );
  XOR \SUBBYTES[6].a/U5621  ( .A(\SUBBYTES[6].a/w3350 ), .B(
        \SUBBYTES[6].a/w3353 ), .Z(n12281) );
  XOR \SUBBYTES[6].a/U5619  ( .A(n13305), .B(n12284), .Z(n12282) );
  XOR \SUBBYTES[6].a/U5618  ( .A(n13307), .B(n13306), .Z(n12283) );
  XOR \SUBBYTES[6].a/U5617  ( .A(\SUBBYTES[6].a/w3358 ), .B(
        \SUBBYTES[6].a/w3385 ), .Z(n12284) );
  XOR \SUBBYTES[6].a/U5615  ( .A(n13308), .B(n12287), .Z(n12285) );
  XOR \SUBBYTES[6].a/U5614  ( .A(\SUBBYTES[6].a/w3391 ), .B(
        \SUBBYTES[6].a/w3393 ), .Z(n12286) );
  XOR \SUBBYTES[6].a/U5613  ( .A(\SUBBYTES[6].a/w3351 ), .B(
        \SUBBYTES[6].a/w3383 ), .Z(n12287) );
  XOR \SUBBYTES[6].a/U5612  ( .A(\SUBBYTES[6].a/w3183 ), .B(
        \SUBBYTES[6].a/w3184 ), .Z(n13310) );
  XOR \SUBBYTES[6].a/U5611  ( .A(n13310), .B(n12288), .Z(n13309) );
  XOR \SUBBYTES[6].a/U5610  ( .A(\SUBBYTES[6].a/w3176 ), .B(
        \SUBBYTES[6].a/w3193 ), .Z(n12288) );
  XOR \SUBBYTES[6].a/U5608  ( .A(\SUBBYTES[6].a/w3175 ), .B(
        \SUBBYTES[6].a/w3190 ), .Z(n12289) );
  XOR \SUBBYTES[6].a/U5607  ( .A(n13310), .B(n12290), .Z(n13497) );
  XOR \SUBBYTES[6].a/U5606  ( .A(\SUBBYTES[6].a/w3190 ), .B(
        \SUBBYTES[6].a/w3191 ), .Z(n12290) );
  XOR \SUBBYTES[6].a/U5605  ( .A(\SUBBYTES[6].a/w3152 ), .B(n12291), .Z(n13312) );
  XOR \SUBBYTES[6].a/U5604  ( .A(\SUBBYTES[6].a/w3143 ), .B(
        \SUBBYTES[6].a/w3144 ), .Z(n12291) );
  XOR \SUBBYTES[6].a/U5602  ( .A(\SUBBYTES[6].a/w3154 ), .B(n13497), .Z(n12292) );
  XOR \SUBBYTES[6].a/U5601  ( .A(n12294), .B(n12293), .Z(n13313) );
  XOR \SUBBYTES[6].a/U5600  ( .A(n12296), .B(n12295), .Z(n12293) );
  XOR \SUBBYTES[6].a/U5599  ( .A(\SUBBYTES[6].a/w3190 ), .B(
        \SUBBYTES[6].a/w3191 ), .Z(n12294) );
  XOR \SUBBYTES[6].a/U5598  ( .A(\SUBBYTES[6].a/w3154 ), .B(
        \SUBBYTES[6].a/w3178 ), .Z(n12295) );
  XOR \SUBBYTES[6].a/U5597  ( .A(\SUBBYTES[6].a/w3143 ), .B(
        \SUBBYTES[6].a/w3152 ), .Z(n12296) );
  XOR \SUBBYTES[6].a/U5596  ( .A(\SUBBYTES[6].a/w3175 ), .B(n12297), .Z(n13311) );
  XOR \SUBBYTES[6].a/U5595  ( .A(\SUBBYTES[6].a/w3158 ), .B(
        \SUBBYTES[6].a/w3161 ), .Z(n12297) );
  XOR \SUBBYTES[6].a/U5593  ( .A(\SUBBYTES[6].a/w3146 ), .B(n13313), .Z(n12298) );
  XOR \SUBBYTES[6].a/U5591  ( .A(\SUBBYTES[6].a/w3178 ), .B(
        \SUBBYTES[6].a/w3191 ), .Z(n12299) );
  XOR \SUBBYTES[6].a/U5589  ( .A(n12303), .B(n12302), .Z(n12300) );
  XOR \SUBBYTES[6].a/U5588  ( .A(n12305), .B(n12304), .Z(n12301) );
  XOR \SUBBYTES[6].a/U5587  ( .A(\SUBBYTES[6].a/w3190 ), .B(
        \SUBBYTES[6].a/w3193 ), .Z(n12302) );
  XOR \SUBBYTES[6].a/U5586  ( .A(\SUBBYTES[6].a/w3183 ), .B(
        \SUBBYTES[6].a/w3186 ), .Z(n12303) );
  XOR \SUBBYTES[6].a/U5585  ( .A(\SUBBYTES[6].a/w3158 ), .B(
        \SUBBYTES[6].a/w3159 ), .Z(n12304) );
  XOR \SUBBYTES[6].a/U5584  ( .A(\SUBBYTES[6].a/w3143 ), .B(
        \SUBBYTES[6].a/w3146 ), .Z(n12305) );
  XOR \SUBBYTES[6].a/U5582  ( .A(n13310), .B(n12308), .Z(n12306) );
  XOR \SUBBYTES[6].a/U5581  ( .A(n13312), .B(n13311), .Z(n12307) );
  XOR \SUBBYTES[6].a/U5580  ( .A(\SUBBYTES[6].a/w3151 ), .B(
        \SUBBYTES[6].a/w3178 ), .Z(n12308) );
  XOR \SUBBYTES[6].a/U5578  ( .A(n13313), .B(n12311), .Z(n12309) );
  XOR \SUBBYTES[6].a/U5577  ( .A(\SUBBYTES[6].a/w3184 ), .B(
        \SUBBYTES[6].a/w3186 ), .Z(n12310) );
  XOR \SUBBYTES[6].a/U5576  ( .A(\SUBBYTES[6].a/w3144 ), .B(
        \SUBBYTES[6].a/w3176 ), .Z(n12311) );
  XOR \SUBBYTES[6].a/U5575  ( .A(\SUBBYTES[6].a/w2976 ), .B(
        \SUBBYTES[6].a/w2977 ), .Z(n13315) );
  XOR \SUBBYTES[6].a/U5574  ( .A(n13315), .B(n12312), .Z(n13314) );
  XOR \SUBBYTES[6].a/U5573  ( .A(\SUBBYTES[6].a/w2969 ), .B(
        \SUBBYTES[6].a/w2986 ), .Z(n12312) );
  XOR \SUBBYTES[6].a/U5571  ( .A(\SUBBYTES[6].a/w2968 ), .B(
        \SUBBYTES[6].a/w2983 ), .Z(n12313) );
  XOR \SUBBYTES[6].a/U5570  ( .A(n13315), .B(n12314), .Z(n13498) );
  XOR \SUBBYTES[6].a/U5569  ( .A(\SUBBYTES[6].a/w2983 ), .B(
        \SUBBYTES[6].a/w2984 ), .Z(n12314) );
  XOR \SUBBYTES[6].a/U5568  ( .A(\SUBBYTES[6].a/w2945 ), .B(n12315), .Z(n13317) );
  XOR \SUBBYTES[6].a/U5567  ( .A(\SUBBYTES[6].a/w2936 ), .B(
        \SUBBYTES[6].a/w2937 ), .Z(n12315) );
  XOR \SUBBYTES[6].a/U5565  ( .A(\SUBBYTES[6].a/w2947 ), .B(n13498), .Z(n12316) );
  XOR \SUBBYTES[6].a/U5564  ( .A(n12318), .B(n12317), .Z(n13318) );
  XOR \SUBBYTES[6].a/U5563  ( .A(n12320), .B(n12319), .Z(n12317) );
  XOR \SUBBYTES[6].a/U5562  ( .A(\SUBBYTES[6].a/w2983 ), .B(
        \SUBBYTES[6].a/w2984 ), .Z(n12318) );
  XOR \SUBBYTES[6].a/U5561  ( .A(\SUBBYTES[6].a/w2947 ), .B(
        \SUBBYTES[6].a/w2971 ), .Z(n12319) );
  XOR \SUBBYTES[6].a/U5560  ( .A(\SUBBYTES[6].a/w2936 ), .B(
        \SUBBYTES[6].a/w2945 ), .Z(n12320) );
  XOR \SUBBYTES[6].a/U5559  ( .A(\SUBBYTES[6].a/w2968 ), .B(n12321), .Z(n13316) );
  XOR \SUBBYTES[6].a/U5558  ( .A(\SUBBYTES[6].a/w2951 ), .B(
        \SUBBYTES[6].a/w2954 ), .Z(n12321) );
  XOR \SUBBYTES[6].a/U5556  ( .A(\SUBBYTES[6].a/w2939 ), .B(n13318), .Z(n12322) );
  XOR \SUBBYTES[6].a/U5554  ( .A(\SUBBYTES[6].a/w2971 ), .B(
        \SUBBYTES[6].a/w2984 ), .Z(n12323) );
  XOR \SUBBYTES[6].a/U5552  ( .A(n12327), .B(n12326), .Z(n12324) );
  XOR \SUBBYTES[6].a/U5551  ( .A(n12329), .B(n12328), .Z(n12325) );
  XOR \SUBBYTES[6].a/U5550  ( .A(\SUBBYTES[6].a/w2983 ), .B(
        \SUBBYTES[6].a/w2986 ), .Z(n12326) );
  XOR \SUBBYTES[6].a/U5549  ( .A(\SUBBYTES[6].a/w2976 ), .B(
        \SUBBYTES[6].a/w2979 ), .Z(n12327) );
  XOR \SUBBYTES[6].a/U5548  ( .A(\SUBBYTES[6].a/w2951 ), .B(
        \SUBBYTES[6].a/w2952 ), .Z(n12328) );
  XOR \SUBBYTES[6].a/U5547  ( .A(\SUBBYTES[6].a/w2936 ), .B(
        \SUBBYTES[6].a/w2939 ), .Z(n12329) );
  XOR \SUBBYTES[6].a/U5545  ( .A(n13315), .B(n12332), .Z(n12330) );
  XOR \SUBBYTES[6].a/U5544  ( .A(n13317), .B(n13316), .Z(n12331) );
  XOR \SUBBYTES[6].a/U5543  ( .A(\SUBBYTES[6].a/w2944 ), .B(
        \SUBBYTES[6].a/w2971 ), .Z(n12332) );
  XOR \SUBBYTES[6].a/U5541  ( .A(n13318), .B(n12335), .Z(n12333) );
  XOR \SUBBYTES[6].a/U5540  ( .A(\SUBBYTES[6].a/w2977 ), .B(
        \SUBBYTES[6].a/w2979 ), .Z(n12334) );
  XOR \SUBBYTES[6].a/U5539  ( .A(\SUBBYTES[6].a/w2937 ), .B(
        \SUBBYTES[6].a/w2969 ), .Z(n12335) );
  XOR \SUBBYTES[6].a/U5538  ( .A(\SUBBYTES[6].a/w2769 ), .B(
        \SUBBYTES[6].a/w2770 ), .Z(n13320) );
  XOR \SUBBYTES[6].a/U5537  ( .A(n13320), .B(n12336), .Z(n13319) );
  XOR \SUBBYTES[6].a/U5536  ( .A(\SUBBYTES[6].a/w2762 ), .B(
        \SUBBYTES[6].a/w2779 ), .Z(n12336) );
  XOR \SUBBYTES[6].a/U5534  ( .A(\SUBBYTES[6].a/w2761 ), .B(
        \SUBBYTES[6].a/w2776 ), .Z(n12337) );
  XOR \SUBBYTES[6].a/U5533  ( .A(n13320), .B(n12338), .Z(n13499) );
  XOR \SUBBYTES[6].a/U5532  ( .A(\SUBBYTES[6].a/w2776 ), .B(
        \SUBBYTES[6].a/w2777 ), .Z(n12338) );
  XOR \SUBBYTES[6].a/U5531  ( .A(\SUBBYTES[6].a/w2738 ), .B(n12339), .Z(n13322) );
  XOR \SUBBYTES[6].a/U5530  ( .A(\SUBBYTES[6].a/w2729 ), .B(
        \SUBBYTES[6].a/w2730 ), .Z(n12339) );
  XOR \SUBBYTES[6].a/U5528  ( .A(\SUBBYTES[6].a/w2740 ), .B(n13499), .Z(n12340) );
  XOR \SUBBYTES[6].a/U5527  ( .A(n12342), .B(n12341), .Z(n13323) );
  XOR \SUBBYTES[6].a/U5526  ( .A(n12344), .B(n12343), .Z(n12341) );
  XOR \SUBBYTES[6].a/U5525  ( .A(\SUBBYTES[6].a/w2776 ), .B(
        \SUBBYTES[6].a/w2777 ), .Z(n12342) );
  XOR \SUBBYTES[6].a/U5524  ( .A(\SUBBYTES[6].a/w2740 ), .B(
        \SUBBYTES[6].a/w2764 ), .Z(n12343) );
  XOR \SUBBYTES[6].a/U5523  ( .A(\SUBBYTES[6].a/w2729 ), .B(
        \SUBBYTES[6].a/w2738 ), .Z(n12344) );
  XOR \SUBBYTES[6].a/U5522  ( .A(\SUBBYTES[6].a/w2761 ), .B(n12345), .Z(n13321) );
  XOR \SUBBYTES[6].a/U5521  ( .A(\SUBBYTES[6].a/w2744 ), .B(
        \SUBBYTES[6].a/w2747 ), .Z(n12345) );
  XOR \SUBBYTES[6].a/U5519  ( .A(\SUBBYTES[6].a/w2732 ), .B(n13323), .Z(n12346) );
  XOR \SUBBYTES[6].a/U5517  ( .A(\SUBBYTES[6].a/w2764 ), .B(
        \SUBBYTES[6].a/w2777 ), .Z(n12347) );
  XOR \SUBBYTES[6].a/U5515  ( .A(n12351), .B(n12350), .Z(n12348) );
  XOR \SUBBYTES[6].a/U5514  ( .A(n12353), .B(n12352), .Z(n12349) );
  XOR \SUBBYTES[6].a/U5513  ( .A(\SUBBYTES[6].a/w2776 ), .B(
        \SUBBYTES[6].a/w2779 ), .Z(n12350) );
  XOR \SUBBYTES[6].a/U5512  ( .A(\SUBBYTES[6].a/w2769 ), .B(
        \SUBBYTES[6].a/w2772 ), .Z(n12351) );
  XOR \SUBBYTES[6].a/U5511  ( .A(\SUBBYTES[6].a/w2744 ), .B(
        \SUBBYTES[6].a/w2745 ), .Z(n12352) );
  XOR \SUBBYTES[6].a/U5510  ( .A(\SUBBYTES[6].a/w2729 ), .B(
        \SUBBYTES[6].a/w2732 ), .Z(n12353) );
  XOR \SUBBYTES[6].a/U5508  ( .A(n13320), .B(n12356), .Z(n12354) );
  XOR \SUBBYTES[6].a/U5507  ( .A(n13322), .B(n13321), .Z(n12355) );
  XOR \SUBBYTES[6].a/U5506  ( .A(\SUBBYTES[6].a/w2737 ), .B(
        \SUBBYTES[6].a/w2764 ), .Z(n12356) );
  XOR \SUBBYTES[6].a/U5504  ( .A(n13323), .B(n12359), .Z(n12357) );
  XOR \SUBBYTES[6].a/U5503  ( .A(\SUBBYTES[6].a/w2770 ), .B(
        \SUBBYTES[6].a/w2772 ), .Z(n12358) );
  XOR \SUBBYTES[6].a/U5502  ( .A(\SUBBYTES[6].a/w2730 ), .B(
        \SUBBYTES[6].a/w2762 ), .Z(n12359) );
  XOR \SUBBYTES[6].a/U5501  ( .A(\SUBBYTES[6].a/w2562 ), .B(
        \SUBBYTES[6].a/w2563 ), .Z(n13325) );
  XOR \SUBBYTES[6].a/U5500  ( .A(n13325), .B(n12360), .Z(n13324) );
  XOR \SUBBYTES[6].a/U5499  ( .A(\SUBBYTES[6].a/w2555 ), .B(
        \SUBBYTES[6].a/w2572 ), .Z(n12360) );
  XOR \SUBBYTES[6].a/U5497  ( .A(\SUBBYTES[6].a/w2554 ), .B(
        \SUBBYTES[6].a/w2569 ), .Z(n12361) );
  XOR \SUBBYTES[6].a/U5496  ( .A(n13325), .B(n12362), .Z(n13500) );
  XOR \SUBBYTES[6].a/U5495  ( .A(\SUBBYTES[6].a/w2569 ), .B(
        \SUBBYTES[6].a/w2570 ), .Z(n12362) );
  XOR \SUBBYTES[6].a/U5494  ( .A(\SUBBYTES[6].a/w2531 ), .B(n12363), .Z(n13327) );
  XOR \SUBBYTES[6].a/U5493  ( .A(\SUBBYTES[6].a/w2522 ), .B(
        \SUBBYTES[6].a/w2523 ), .Z(n12363) );
  XOR \SUBBYTES[6].a/U5491  ( .A(\SUBBYTES[6].a/w2533 ), .B(n13500), .Z(n12364) );
  XOR \SUBBYTES[6].a/U5490  ( .A(n12366), .B(n12365), .Z(n13328) );
  XOR \SUBBYTES[6].a/U5489  ( .A(n12368), .B(n12367), .Z(n12365) );
  XOR \SUBBYTES[6].a/U5488  ( .A(\SUBBYTES[6].a/w2569 ), .B(
        \SUBBYTES[6].a/w2570 ), .Z(n12366) );
  XOR \SUBBYTES[6].a/U5487  ( .A(\SUBBYTES[6].a/w2533 ), .B(
        \SUBBYTES[6].a/w2557 ), .Z(n12367) );
  XOR \SUBBYTES[6].a/U5486  ( .A(\SUBBYTES[6].a/w2522 ), .B(
        \SUBBYTES[6].a/w2531 ), .Z(n12368) );
  XOR \SUBBYTES[6].a/U5485  ( .A(\SUBBYTES[6].a/w2554 ), .B(n12369), .Z(n13326) );
  XOR \SUBBYTES[6].a/U5484  ( .A(\SUBBYTES[6].a/w2537 ), .B(
        \SUBBYTES[6].a/w2540 ), .Z(n12369) );
  XOR \SUBBYTES[6].a/U5482  ( .A(\SUBBYTES[6].a/w2525 ), .B(n13328), .Z(n12370) );
  XOR \SUBBYTES[6].a/U5480  ( .A(\SUBBYTES[6].a/w2557 ), .B(
        \SUBBYTES[6].a/w2570 ), .Z(n12371) );
  XOR \SUBBYTES[6].a/U5478  ( .A(n12375), .B(n12374), .Z(n12372) );
  XOR \SUBBYTES[6].a/U5477  ( .A(n12377), .B(n12376), .Z(n12373) );
  XOR \SUBBYTES[6].a/U5476  ( .A(\SUBBYTES[6].a/w2569 ), .B(
        \SUBBYTES[6].a/w2572 ), .Z(n12374) );
  XOR \SUBBYTES[6].a/U5475  ( .A(\SUBBYTES[6].a/w2562 ), .B(
        \SUBBYTES[6].a/w2565 ), .Z(n12375) );
  XOR \SUBBYTES[6].a/U5474  ( .A(\SUBBYTES[6].a/w2537 ), .B(
        \SUBBYTES[6].a/w2538 ), .Z(n12376) );
  XOR \SUBBYTES[6].a/U5473  ( .A(\SUBBYTES[6].a/w2522 ), .B(
        \SUBBYTES[6].a/w2525 ), .Z(n12377) );
  XOR \SUBBYTES[6].a/U5471  ( .A(n13325), .B(n12380), .Z(n12378) );
  XOR \SUBBYTES[6].a/U5470  ( .A(n13327), .B(n13326), .Z(n12379) );
  XOR \SUBBYTES[6].a/U5469  ( .A(\SUBBYTES[6].a/w2530 ), .B(
        \SUBBYTES[6].a/w2557 ), .Z(n12380) );
  XOR \SUBBYTES[6].a/U5467  ( .A(n13328), .B(n12383), .Z(n12381) );
  XOR \SUBBYTES[6].a/U5466  ( .A(\SUBBYTES[6].a/w2563 ), .B(
        \SUBBYTES[6].a/w2565 ), .Z(n12382) );
  XOR \SUBBYTES[6].a/U5465  ( .A(\SUBBYTES[6].a/w2523 ), .B(
        \SUBBYTES[6].a/w2555 ), .Z(n12383) );
  XOR \SUBBYTES[6].a/U5464  ( .A(\SUBBYTES[6].a/w2355 ), .B(
        \SUBBYTES[6].a/w2356 ), .Z(n13330) );
  XOR \SUBBYTES[6].a/U5463  ( .A(n13330), .B(n12384), .Z(n13329) );
  XOR \SUBBYTES[6].a/U5462  ( .A(\SUBBYTES[6].a/w2348 ), .B(
        \SUBBYTES[6].a/w2365 ), .Z(n12384) );
  XOR \SUBBYTES[6].a/U5460  ( .A(\SUBBYTES[6].a/w2347 ), .B(
        \SUBBYTES[6].a/w2362 ), .Z(n12385) );
  XOR \SUBBYTES[6].a/U5459  ( .A(n13330), .B(n12386), .Z(n13501) );
  XOR \SUBBYTES[6].a/U5458  ( .A(\SUBBYTES[6].a/w2362 ), .B(
        \SUBBYTES[6].a/w2363 ), .Z(n12386) );
  XOR \SUBBYTES[6].a/U5457  ( .A(\SUBBYTES[6].a/w2324 ), .B(n12387), .Z(n13332) );
  XOR \SUBBYTES[6].a/U5456  ( .A(\SUBBYTES[6].a/w2315 ), .B(
        \SUBBYTES[6].a/w2316 ), .Z(n12387) );
  XOR \SUBBYTES[6].a/U5454  ( .A(\SUBBYTES[6].a/w2326 ), .B(n13501), .Z(n12388) );
  XOR \SUBBYTES[6].a/U5453  ( .A(n12390), .B(n12389), .Z(n13333) );
  XOR \SUBBYTES[6].a/U5452  ( .A(n12392), .B(n12391), .Z(n12389) );
  XOR \SUBBYTES[6].a/U5451  ( .A(\SUBBYTES[6].a/w2362 ), .B(
        \SUBBYTES[6].a/w2363 ), .Z(n12390) );
  XOR \SUBBYTES[6].a/U5450  ( .A(\SUBBYTES[6].a/w2326 ), .B(
        \SUBBYTES[6].a/w2350 ), .Z(n12391) );
  XOR \SUBBYTES[6].a/U5449  ( .A(\SUBBYTES[6].a/w2315 ), .B(
        \SUBBYTES[6].a/w2324 ), .Z(n12392) );
  XOR \SUBBYTES[6].a/U5448  ( .A(\SUBBYTES[6].a/w2347 ), .B(n12393), .Z(n13331) );
  XOR \SUBBYTES[6].a/U5447  ( .A(\SUBBYTES[6].a/w2330 ), .B(
        \SUBBYTES[6].a/w2333 ), .Z(n12393) );
  XOR \SUBBYTES[6].a/U5445  ( .A(\SUBBYTES[6].a/w2318 ), .B(n13333), .Z(n12394) );
  XOR \SUBBYTES[6].a/U5443  ( .A(\SUBBYTES[6].a/w2350 ), .B(
        \SUBBYTES[6].a/w2363 ), .Z(n12395) );
  XOR \SUBBYTES[6].a/U5441  ( .A(n12399), .B(n12398), .Z(n12396) );
  XOR \SUBBYTES[6].a/U5440  ( .A(n12401), .B(n12400), .Z(n12397) );
  XOR \SUBBYTES[6].a/U5439  ( .A(\SUBBYTES[6].a/w2362 ), .B(
        \SUBBYTES[6].a/w2365 ), .Z(n12398) );
  XOR \SUBBYTES[6].a/U5438  ( .A(\SUBBYTES[6].a/w2355 ), .B(
        \SUBBYTES[6].a/w2358 ), .Z(n12399) );
  XOR \SUBBYTES[6].a/U5437  ( .A(\SUBBYTES[6].a/w2330 ), .B(
        \SUBBYTES[6].a/w2331 ), .Z(n12400) );
  XOR \SUBBYTES[6].a/U5436  ( .A(\SUBBYTES[6].a/w2315 ), .B(
        \SUBBYTES[6].a/w2318 ), .Z(n12401) );
  XOR \SUBBYTES[6].a/U5434  ( .A(n13330), .B(n12404), .Z(n12402) );
  XOR \SUBBYTES[6].a/U5433  ( .A(n13332), .B(n13331), .Z(n12403) );
  XOR \SUBBYTES[6].a/U5432  ( .A(\SUBBYTES[6].a/w2323 ), .B(
        \SUBBYTES[6].a/w2350 ), .Z(n12404) );
  XOR \SUBBYTES[6].a/U5430  ( .A(n13333), .B(n12407), .Z(n12405) );
  XOR \SUBBYTES[6].a/U5429  ( .A(\SUBBYTES[6].a/w2356 ), .B(
        \SUBBYTES[6].a/w2358 ), .Z(n12406) );
  XOR \SUBBYTES[6].a/U5428  ( .A(\SUBBYTES[6].a/w2316 ), .B(
        \SUBBYTES[6].a/w2348 ), .Z(n12407) );
  XOR \SUBBYTES[6].a/U5427  ( .A(\SUBBYTES[6].a/w2148 ), .B(
        \SUBBYTES[6].a/w2149 ), .Z(n13335) );
  XOR \SUBBYTES[6].a/U5426  ( .A(n13335), .B(n12408), .Z(n13334) );
  XOR \SUBBYTES[6].a/U5425  ( .A(\SUBBYTES[6].a/w2141 ), .B(
        \SUBBYTES[6].a/w2158 ), .Z(n12408) );
  XOR \SUBBYTES[6].a/U5423  ( .A(\SUBBYTES[6].a/w2140 ), .B(
        \SUBBYTES[6].a/w2155 ), .Z(n12409) );
  XOR \SUBBYTES[6].a/U5422  ( .A(n13335), .B(n12410), .Z(n13502) );
  XOR \SUBBYTES[6].a/U5421  ( .A(\SUBBYTES[6].a/w2155 ), .B(
        \SUBBYTES[6].a/w2156 ), .Z(n12410) );
  XOR \SUBBYTES[6].a/U5420  ( .A(\SUBBYTES[6].a/w2117 ), .B(n12411), .Z(n13337) );
  XOR \SUBBYTES[6].a/U5419  ( .A(\SUBBYTES[6].a/w2108 ), .B(
        \SUBBYTES[6].a/w2109 ), .Z(n12411) );
  XOR \SUBBYTES[6].a/U5417  ( .A(\SUBBYTES[6].a/w2119 ), .B(n13502), .Z(n12412) );
  XOR \SUBBYTES[6].a/U5416  ( .A(n12414), .B(n12413), .Z(n13338) );
  XOR \SUBBYTES[6].a/U5415  ( .A(n12416), .B(n12415), .Z(n12413) );
  XOR \SUBBYTES[6].a/U5414  ( .A(\SUBBYTES[6].a/w2155 ), .B(
        \SUBBYTES[6].a/w2156 ), .Z(n12414) );
  XOR \SUBBYTES[6].a/U5413  ( .A(\SUBBYTES[6].a/w2119 ), .B(
        \SUBBYTES[6].a/w2143 ), .Z(n12415) );
  XOR \SUBBYTES[6].a/U5412  ( .A(\SUBBYTES[6].a/w2108 ), .B(
        \SUBBYTES[6].a/w2117 ), .Z(n12416) );
  XOR \SUBBYTES[6].a/U5411  ( .A(\SUBBYTES[6].a/w2140 ), .B(n12417), .Z(n13336) );
  XOR \SUBBYTES[6].a/U5410  ( .A(\SUBBYTES[6].a/w2123 ), .B(
        \SUBBYTES[6].a/w2126 ), .Z(n12417) );
  XOR \SUBBYTES[6].a/U5408  ( .A(\SUBBYTES[6].a/w2111 ), .B(n13338), .Z(n12418) );
  XOR \SUBBYTES[6].a/U5406  ( .A(\SUBBYTES[6].a/w2143 ), .B(
        \SUBBYTES[6].a/w2156 ), .Z(n12419) );
  XOR \SUBBYTES[6].a/U5404  ( .A(n12423), .B(n12422), .Z(n12420) );
  XOR \SUBBYTES[6].a/U5403  ( .A(n12425), .B(n12424), .Z(n12421) );
  XOR \SUBBYTES[6].a/U5402  ( .A(\SUBBYTES[6].a/w2155 ), .B(
        \SUBBYTES[6].a/w2158 ), .Z(n12422) );
  XOR \SUBBYTES[6].a/U5401  ( .A(\SUBBYTES[6].a/w2148 ), .B(
        \SUBBYTES[6].a/w2151 ), .Z(n12423) );
  XOR \SUBBYTES[6].a/U5400  ( .A(\SUBBYTES[6].a/w2123 ), .B(
        \SUBBYTES[6].a/w2124 ), .Z(n12424) );
  XOR \SUBBYTES[6].a/U5399  ( .A(\SUBBYTES[6].a/w2108 ), .B(
        \SUBBYTES[6].a/w2111 ), .Z(n12425) );
  XOR \SUBBYTES[6].a/U5397  ( .A(n13335), .B(n12428), .Z(n12426) );
  XOR \SUBBYTES[6].a/U5396  ( .A(n13337), .B(n13336), .Z(n12427) );
  XOR \SUBBYTES[6].a/U5395  ( .A(\SUBBYTES[6].a/w2116 ), .B(
        \SUBBYTES[6].a/w2143 ), .Z(n12428) );
  XOR \SUBBYTES[6].a/U5393  ( .A(n13338), .B(n12431), .Z(n12429) );
  XOR \SUBBYTES[6].a/U5392  ( .A(\SUBBYTES[6].a/w2149 ), .B(
        \SUBBYTES[6].a/w2151 ), .Z(n12430) );
  XOR \SUBBYTES[6].a/U5391  ( .A(\SUBBYTES[6].a/w2109 ), .B(
        \SUBBYTES[6].a/w2141 ), .Z(n12431) );
  XOR \SUBBYTES[6].a/U5390  ( .A(\SUBBYTES[6].a/w1941 ), .B(
        \SUBBYTES[6].a/w1942 ), .Z(n13340) );
  XOR \SUBBYTES[6].a/U5389  ( .A(n13340), .B(n12432), .Z(n13339) );
  XOR \SUBBYTES[6].a/U5388  ( .A(\SUBBYTES[6].a/w1934 ), .B(
        \SUBBYTES[6].a/w1951 ), .Z(n12432) );
  XOR \SUBBYTES[6].a/U5386  ( .A(\SUBBYTES[6].a/w1933 ), .B(
        \SUBBYTES[6].a/w1948 ), .Z(n12433) );
  XOR \SUBBYTES[6].a/U5385  ( .A(n13340), .B(n12434), .Z(n13503) );
  XOR \SUBBYTES[6].a/U5384  ( .A(\SUBBYTES[6].a/w1948 ), .B(
        \SUBBYTES[6].a/w1949 ), .Z(n12434) );
  XOR \SUBBYTES[6].a/U5383  ( .A(\SUBBYTES[6].a/w1910 ), .B(n12435), .Z(n13342) );
  XOR \SUBBYTES[6].a/U5382  ( .A(\SUBBYTES[6].a/w1901 ), .B(
        \SUBBYTES[6].a/w1902 ), .Z(n12435) );
  XOR \SUBBYTES[6].a/U5380  ( .A(\SUBBYTES[6].a/w1912 ), .B(n13503), .Z(n12436) );
  XOR \SUBBYTES[6].a/U5379  ( .A(n12438), .B(n12437), .Z(n13343) );
  XOR \SUBBYTES[6].a/U5378  ( .A(n12440), .B(n12439), .Z(n12437) );
  XOR \SUBBYTES[6].a/U5377  ( .A(\SUBBYTES[6].a/w1948 ), .B(
        \SUBBYTES[6].a/w1949 ), .Z(n12438) );
  XOR \SUBBYTES[6].a/U5376  ( .A(\SUBBYTES[6].a/w1912 ), .B(
        \SUBBYTES[6].a/w1936 ), .Z(n12439) );
  XOR \SUBBYTES[6].a/U5375  ( .A(\SUBBYTES[6].a/w1901 ), .B(
        \SUBBYTES[6].a/w1910 ), .Z(n12440) );
  XOR \SUBBYTES[6].a/U5374  ( .A(\SUBBYTES[6].a/w1933 ), .B(n12441), .Z(n13341) );
  XOR \SUBBYTES[6].a/U5373  ( .A(\SUBBYTES[6].a/w1916 ), .B(
        \SUBBYTES[6].a/w1919 ), .Z(n12441) );
  XOR \SUBBYTES[6].a/U5371  ( .A(\SUBBYTES[6].a/w1904 ), .B(n13343), .Z(n12442) );
  XOR \SUBBYTES[6].a/U5369  ( .A(\SUBBYTES[6].a/w1936 ), .B(
        \SUBBYTES[6].a/w1949 ), .Z(n12443) );
  XOR \SUBBYTES[6].a/U5367  ( .A(n12447), .B(n12446), .Z(n12444) );
  XOR \SUBBYTES[6].a/U5366  ( .A(n12449), .B(n12448), .Z(n12445) );
  XOR \SUBBYTES[6].a/U5365  ( .A(\SUBBYTES[6].a/w1948 ), .B(
        \SUBBYTES[6].a/w1951 ), .Z(n12446) );
  XOR \SUBBYTES[6].a/U5364  ( .A(\SUBBYTES[6].a/w1941 ), .B(
        \SUBBYTES[6].a/w1944 ), .Z(n12447) );
  XOR \SUBBYTES[6].a/U5363  ( .A(\SUBBYTES[6].a/w1916 ), .B(
        \SUBBYTES[6].a/w1917 ), .Z(n12448) );
  XOR \SUBBYTES[6].a/U5362  ( .A(\SUBBYTES[6].a/w1901 ), .B(
        \SUBBYTES[6].a/w1904 ), .Z(n12449) );
  XOR \SUBBYTES[6].a/U5360  ( .A(n13340), .B(n12452), .Z(n12450) );
  XOR \SUBBYTES[6].a/U5359  ( .A(n13342), .B(n13341), .Z(n12451) );
  XOR \SUBBYTES[6].a/U5358  ( .A(\SUBBYTES[6].a/w1909 ), .B(
        \SUBBYTES[6].a/w1936 ), .Z(n12452) );
  XOR \SUBBYTES[6].a/U5356  ( .A(n13343), .B(n12455), .Z(n12453) );
  XOR \SUBBYTES[6].a/U5355  ( .A(\SUBBYTES[6].a/w1942 ), .B(
        \SUBBYTES[6].a/w1944 ), .Z(n12454) );
  XOR \SUBBYTES[6].a/U5354  ( .A(\SUBBYTES[6].a/w1902 ), .B(
        \SUBBYTES[6].a/w1934 ), .Z(n12455) );
  XOR \SUBBYTES[6].a/U5353  ( .A(\SUBBYTES[6].a/w1734 ), .B(
        \SUBBYTES[6].a/w1735 ), .Z(n13345) );
  XOR \SUBBYTES[6].a/U5352  ( .A(n13345), .B(n12456), .Z(n13344) );
  XOR \SUBBYTES[6].a/U5351  ( .A(\SUBBYTES[6].a/w1727 ), .B(
        \SUBBYTES[6].a/w1744 ), .Z(n12456) );
  XOR \SUBBYTES[6].a/U5349  ( .A(\SUBBYTES[6].a/w1726 ), .B(
        \SUBBYTES[6].a/w1741 ), .Z(n12457) );
  XOR \SUBBYTES[6].a/U5348  ( .A(n13345), .B(n12458), .Z(n13504) );
  XOR \SUBBYTES[6].a/U5347  ( .A(\SUBBYTES[6].a/w1741 ), .B(
        \SUBBYTES[6].a/w1742 ), .Z(n12458) );
  XOR \SUBBYTES[6].a/U5346  ( .A(\SUBBYTES[6].a/w1703 ), .B(n12459), .Z(n13347) );
  XOR \SUBBYTES[6].a/U5345  ( .A(\SUBBYTES[6].a/w1694 ), .B(
        \SUBBYTES[6].a/w1695 ), .Z(n12459) );
  XOR \SUBBYTES[6].a/U5343  ( .A(\SUBBYTES[6].a/w1705 ), .B(n13504), .Z(n12460) );
  XOR \SUBBYTES[6].a/U5342  ( .A(n12462), .B(n12461), .Z(n13348) );
  XOR \SUBBYTES[6].a/U5341  ( .A(n12464), .B(n12463), .Z(n12461) );
  XOR \SUBBYTES[6].a/U5340  ( .A(\SUBBYTES[6].a/w1741 ), .B(
        \SUBBYTES[6].a/w1742 ), .Z(n12462) );
  XOR \SUBBYTES[6].a/U5339  ( .A(\SUBBYTES[6].a/w1705 ), .B(
        \SUBBYTES[6].a/w1729 ), .Z(n12463) );
  XOR \SUBBYTES[6].a/U5338  ( .A(\SUBBYTES[6].a/w1694 ), .B(
        \SUBBYTES[6].a/w1703 ), .Z(n12464) );
  XOR \SUBBYTES[6].a/U5337  ( .A(\SUBBYTES[6].a/w1726 ), .B(n12465), .Z(n13346) );
  XOR \SUBBYTES[6].a/U5336  ( .A(\SUBBYTES[6].a/w1709 ), .B(
        \SUBBYTES[6].a/w1712 ), .Z(n12465) );
  XOR \SUBBYTES[6].a/U5334  ( .A(\SUBBYTES[6].a/w1697 ), .B(n13348), .Z(n12466) );
  XOR \SUBBYTES[6].a/U5332  ( .A(\SUBBYTES[6].a/w1729 ), .B(
        \SUBBYTES[6].a/w1742 ), .Z(n12467) );
  XOR \SUBBYTES[6].a/U5330  ( .A(n12471), .B(n12470), .Z(n12468) );
  XOR \SUBBYTES[6].a/U5329  ( .A(n12473), .B(n12472), .Z(n12469) );
  XOR \SUBBYTES[6].a/U5328  ( .A(\SUBBYTES[6].a/w1741 ), .B(
        \SUBBYTES[6].a/w1744 ), .Z(n12470) );
  XOR \SUBBYTES[6].a/U5327  ( .A(\SUBBYTES[6].a/w1734 ), .B(
        \SUBBYTES[6].a/w1737 ), .Z(n12471) );
  XOR \SUBBYTES[6].a/U5326  ( .A(\SUBBYTES[6].a/w1709 ), .B(
        \SUBBYTES[6].a/w1710 ), .Z(n12472) );
  XOR \SUBBYTES[6].a/U5325  ( .A(\SUBBYTES[6].a/w1694 ), .B(
        \SUBBYTES[6].a/w1697 ), .Z(n12473) );
  XOR \SUBBYTES[6].a/U5323  ( .A(n13345), .B(n12476), .Z(n12474) );
  XOR \SUBBYTES[6].a/U5322  ( .A(n13347), .B(n13346), .Z(n12475) );
  XOR \SUBBYTES[6].a/U5321  ( .A(\SUBBYTES[6].a/w1702 ), .B(
        \SUBBYTES[6].a/w1729 ), .Z(n12476) );
  XOR \SUBBYTES[6].a/U5319  ( .A(n13348), .B(n12479), .Z(n12477) );
  XOR \SUBBYTES[6].a/U5318  ( .A(\SUBBYTES[6].a/w1735 ), .B(
        \SUBBYTES[6].a/w1737 ), .Z(n12478) );
  XOR \SUBBYTES[6].a/U5317  ( .A(\SUBBYTES[6].a/w1695 ), .B(
        \SUBBYTES[6].a/w1727 ), .Z(n12479) );
  XOR \SUBBYTES[6].a/U5316  ( .A(\SUBBYTES[6].a/w1527 ), .B(
        \SUBBYTES[6].a/w1528 ), .Z(n13350) );
  XOR \SUBBYTES[6].a/U5315  ( .A(n13350), .B(n12480), .Z(n13349) );
  XOR \SUBBYTES[6].a/U5314  ( .A(\SUBBYTES[6].a/w1520 ), .B(
        \SUBBYTES[6].a/w1537 ), .Z(n12480) );
  XOR \SUBBYTES[6].a/U5312  ( .A(\SUBBYTES[6].a/w1519 ), .B(
        \SUBBYTES[6].a/w1534 ), .Z(n12481) );
  XOR \SUBBYTES[6].a/U5311  ( .A(n13350), .B(n12482), .Z(n13505) );
  XOR \SUBBYTES[6].a/U5310  ( .A(\SUBBYTES[6].a/w1534 ), .B(
        \SUBBYTES[6].a/w1535 ), .Z(n12482) );
  XOR \SUBBYTES[6].a/U5309  ( .A(\SUBBYTES[6].a/w1496 ), .B(n12483), .Z(n13352) );
  XOR \SUBBYTES[6].a/U5308  ( .A(\SUBBYTES[6].a/w1487 ), .B(
        \SUBBYTES[6].a/w1488 ), .Z(n12483) );
  XOR \SUBBYTES[6].a/U5306  ( .A(\SUBBYTES[6].a/w1498 ), .B(n13505), .Z(n12484) );
  XOR \SUBBYTES[6].a/U5305  ( .A(n12486), .B(n12485), .Z(n13353) );
  XOR \SUBBYTES[6].a/U5304  ( .A(n12488), .B(n12487), .Z(n12485) );
  XOR \SUBBYTES[6].a/U5303  ( .A(\SUBBYTES[6].a/w1534 ), .B(
        \SUBBYTES[6].a/w1535 ), .Z(n12486) );
  XOR \SUBBYTES[6].a/U5302  ( .A(\SUBBYTES[6].a/w1498 ), .B(
        \SUBBYTES[6].a/w1522 ), .Z(n12487) );
  XOR \SUBBYTES[6].a/U5301  ( .A(\SUBBYTES[6].a/w1487 ), .B(
        \SUBBYTES[6].a/w1496 ), .Z(n12488) );
  XOR \SUBBYTES[6].a/U5300  ( .A(\SUBBYTES[6].a/w1519 ), .B(n12489), .Z(n13351) );
  XOR \SUBBYTES[6].a/U5299  ( .A(\SUBBYTES[6].a/w1502 ), .B(
        \SUBBYTES[6].a/w1505 ), .Z(n12489) );
  XOR \SUBBYTES[6].a/U5297  ( .A(\SUBBYTES[6].a/w1490 ), .B(n13353), .Z(n12490) );
  XOR \SUBBYTES[6].a/U5295  ( .A(\SUBBYTES[6].a/w1522 ), .B(
        \SUBBYTES[6].a/w1535 ), .Z(n12491) );
  XOR \SUBBYTES[6].a/U5293  ( .A(n12495), .B(n12494), .Z(n12492) );
  XOR \SUBBYTES[6].a/U5292  ( .A(n12497), .B(n12496), .Z(n12493) );
  XOR \SUBBYTES[6].a/U5291  ( .A(\SUBBYTES[6].a/w1534 ), .B(
        \SUBBYTES[6].a/w1537 ), .Z(n12494) );
  XOR \SUBBYTES[6].a/U5290  ( .A(\SUBBYTES[6].a/w1527 ), .B(
        \SUBBYTES[6].a/w1530 ), .Z(n12495) );
  XOR \SUBBYTES[6].a/U5289  ( .A(\SUBBYTES[6].a/w1502 ), .B(
        \SUBBYTES[6].a/w1503 ), .Z(n12496) );
  XOR \SUBBYTES[6].a/U5288  ( .A(\SUBBYTES[6].a/w1487 ), .B(
        \SUBBYTES[6].a/w1490 ), .Z(n12497) );
  XOR \SUBBYTES[6].a/U5286  ( .A(n13350), .B(n12500), .Z(n12498) );
  XOR \SUBBYTES[6].a/U5285  ( .A(n13352), .B(n13351), .Z(n12499) );
  XOR \SUBBYTES[6].a/U5284  ( .A(\SUBBYTES[6].a/w1495 ), .B(
        \SUBBYTES[6].a/w1522 ), .Z(n12500) );
  XOR \SUBBYTES[6].a/U5282  ( .A(n13353), .B(n12503), .Z(n12501) );
  XOR \SUBBYTES[6].a/U5281  ( .A(\SUBBYTES[6].a/w1528 ), .B(
        \SUBBYTES[6].a/w1530 ), .Z(n12502) );
  XOR \SUBBYTES[6].a/U5280  ( .A(\SUBBYTES[6].a/w1488 ), .B(
        \SUBBYTES[6].a/w1520 ), .Z(n12503) );
  XOR \SUBBYTES[6].a/U5279  ( .A(\SUBBYTES[6].a/w1320 ), .B(
        \SUBBYTES[6].a/w1321 ), .Z(n13355) );
  XOR \SUBBYTES[6].a/U5278  ( .A(n13355), .B(n12504), .Z(n13354) );
  XOR \SUBBYTES[6].a/U5277  ( .A(\SUBBYTES[6].a/w1313 ), .B(
        \SUBBYTES[6].a/w1330 ), .Z(n12504) );
  XOR \SUBBYTES[6].a/U5275  ( .A(\SUBBYTES[6].a/w1312 ), .B(
        \SUBBYTES[6].a/w1327 ), .Z(n12505) );
  XOR \SUBBYTES[6].a/U5274  ( .A(n13355), .B(n12506), .Z(n13506) );
  XOR \SUBBYTES[6].a/U5273  ( .A(\SUBBYTES[6].a/w1327 ), .B(
        \SUBBYTES[6].a/w1328 ), .Z(n12506) );
  XOR \SUBBYTES[6].a/U5272  ( .A(\SUBBYTES[6].a/w1289 ), .B(n12507), .Z(n13357) );
  XOR \SUBBYTES[6].a/U5271  ( .A(\SUBBYTES[6].a/w1280 ), .B(
        \SUBBYTES[6].a/w1281 ), .Z(n12507) );
  XOR \SUBBYTES[6].a/U5269  ( .A(\SUBBYTES[6].a/w1291 ), .B(n13506), .Z(n12508) );
  XOR \SUBBYTES[6].a/U5268  ( .A(n12510), .B(n12509), .Z(n13358) );
  XOR \SUBBYTES[6].a/U5267  ( .A(n12512), .B(n12511), .Z(n12509) );
  XOR \SUBBYTES[6].a/U5266  ( .A(\SUBBYTES[6].a/w1327 ), .B(
        \SUBBYTES[6].a/w1328 ), .Z(n12510) );
  XOR \SUBBYTES[6].a/U5265  ( .A(\SUBBYTES[6].a/w1291 ), .B(
        \SUBBYTES[6].a/w1315 ), .Z(n12511) );
  XOR \SUBBYTES[6].a/U5264  ( .A(\SUBBYTES[6].a/w1280 ), .B(
        \SUBBYTES[6].a/w1289 ), .Z(n12512) );
  XOR \SUBBYTES[6].a/U5263  ( .A(\SUBBYTES[6].a/w1312 ), .B(n12513), .Z(n13356) );
  XOR \SUBBYTES[6].a/U5262  ( .A(\SUBBYTES[6].a/w1295 ), .B(
        \SUBBYTES[6].a/w1298 ), .Z(n12513) );
  XOR \SUBBYTES[6].a/U5260  ( .A(\SUBBYTES[6].a/w1283 ), .B(n13358), .Z(n12514) );
  XOR \SUBBYTES[6].a/U5258  ( .A(\SUBBYTES[6].a/w1315 ), .B(
        \SUBBYTES[6].a/w1328 ), .Z(n12515) );
  XOR \SUBBYTES[6].a/U5256  ( .A(n12519), .B(n12518), .Z(n12516) );
  XOR \SUBBYTES[6].a/U5255  ( .A(n12521), .B(n12520), .Z(n12517) );
  XOR \SUBBYTES[6].a/U5254  ( .A(\SUBBYTES[6].a/w1327 ), .B(
        \SUBBYTES[6].a/w1330 ), .Z(n12518) );
  XOR \SUBBYTES[6].a/U5253  ( .A(\SUBBYTES[6].a/w1320 ), .B(
        \SUBBYTES[6].a/w1323 ), .Z(n12519) );
  XOR \SUBBYTES[6].a/U5252  ( .A(\SUBBYTES[6].a/w1295 ), .B(
        \SUBBYTES[6].a/w1296 ), .Z(n12520) );
  XOR \SUBBYTES[6].a/U5251  ( .A(\SUBBYTES[6].a/w1280 ), .B(
        \SUBBYTES[6].a/w1283 ), .Z(n12521) );
  XOR \SUBBYTES[6].a/U5249  ( .A(n13355), .B(n12524), .Z(n12522) );
  XOR \SUBBYTES[6].a/U5248  ( .A(n13357), .B(n13356), .Z(n12523) );
  XOR \SUBBYTES[6].a/U5247  ( .A(\SUBBYTES[6].a/w1288 ), .B(
        \SUBBYTES[6].a/w1315 ), .Z(n12524) );
  XOR \SUBBYTES[6].a/U5245  ( .A(n13358), .B(n12527), .Z(n12525) );
  XOR \SUBBYTES[6].a/U5244  ( .A(\SUBBYTES[6].a/w1321 ), .B(
        \SUBBYTES[6].a/w1323 ), .Z(n12526) );
  XOR \SUBBYTES[6].a/U5243  ( .A(\SUBBYTES[6].a/w1281 ), .B(
        \SUBBYTES[6].a/w1313 ), .Z(n12527) );
  XOR \SUBBYTES[6].a/U5242  ( .A(\SUBBYTES[6].a/w1113 ), .B(
        \SUBBYTES[6].a/w1114 ), .Z(n13360) );
  XOR \SUBBYTES[6].a/U5241  ( .A(n13360), .B(n12528), .Z(n13359) );
  XOR \SUBBYTES[6].a/U5240  ( .A(\SUBBYTES[6].a/w1106 ), .B(
        \SUBBYTES[6].a/w1123 ), .Z(n12528) );
  XOR \SUBBYTES[6].a/U5238  ( .A(\SUBBYTES[6].a/w1105 ), .B(
        \SUBBYTES[6].a/w1120 ), .Z(n12529) );
  XOR \SUBBYTES[6].a/U5237  ( .A(n13360), .B(n12530), .Z(n13507) );
  XOR \SUBBYTES[6].a/U5236  ( .A(\SUBBYTES[6].a/w1120 ), .B(
        \SUBBYTES[6].a/w1121 ), .Z(n12530) );
  XOR \SUBBYTES[6].a/U5235  ( .A(\SUBBYTES[6].a/w1082 ), .B(n12531), .Z(n13362) );
  XOR \SUBBYTES[6].a/U5234  ( .A(\SUBBYTES[6].a/w1073 ), .B(
        \SUBBYTES[6].a/w1074 ), .Z(n12531) );
  XOR \SUBBYTES[6].a/U5232  ( .A(\SUBBYTES[6].a/w1084 ), .B(n13507), .Z(n12532) );
  XOR \SUBBYTES[6].a/U5231  ( .A(n12534), .B(n12533), .Z(n13363) );
  XOR \SUBBYTES[6].a/U5230  ( .A(n12536), .B(n12535), .Z(n12533) );
  XOR \SUBBYTES[6].a/U5229  ( .A(\SUBBYTES[6].a/w1120 ), .B(
        \SUBBYTES[6].a/w1121 ), .Z(n12534) );
  XOR \SUBBYTES[6].a/U5228  ( .A(\SUBBYTES[6].a/w1084 ), .B(
        \SUBBYTES[6].a/w1108 ), .Z(n12535) );
  XOR \SUBBYTES[6].a/U5227  ( .A(\SUBBYTES[6].a/w1073 ), .B(
        \SUBBYTES[6].a/w1082 ), .Z(n12536) );
  XOR \SUBBYTES[6].a/U5226  ( .A(\SUBBYTES[6].a/w1105 ), .B(n12537), .Z(n13361) );
  XOR \SUBBYTES[6].a/U5225  ( .A(\SUBBYTES[6].a/w1088 ), .B(
        \SUBBYTES[6].a/w1091 ), .Z(n12537) );
  XOR \SUBBYTES[6].a/U5223  ( .A(\SUBBYTES[6].a/w1076 ), .B(n13363), .Z(n12538) );
  XOR \SUBBYTES[6].a/U5221  ( .A(\SUBBYTES[6].a/w1108 ), .B(
        \SUBBYTES[6].a/w1121 ), .Z(n12539) );
  XOR \SUBBYTES[6].a/U5219  ( .A(n12543), .B(n12542), .Z(n12540) );
  XOR \SUBBYTES[6].a/U5218  ( .A(n12545), .B(n12544), .Z(n12541) );
  XOR \SUBBYTES[6].a/U5217  ( .A(\SUBBYTES[6].a/w1120 ), .B(
        \SUBBYTES[6].a/w1123 ), .Z(n12542) );
  XOR \SUBBYTES[6].a/U5216  ( .A(\SUBBYTES[6].a/w1113 ), .B(
        \SUBBYTES[6].a/w1116 ), .Z(n12543) );
  XOR \SUBBYTES[6].a/U5215  ( .A(\SUBBYTES[6].a/w1088 ), .B(
        \SUBBYTES[6].a/w1089 ), .Z(n12544) );
  XOR \SUBBYTES[6].a/U5214  ( .A(\SUBBYTES[6].a/w1073 ), .B(
        \SUBBYTES[6].a/w1076 ), .Z(n12545) );
  XOR \SUBBYTES[6].a/U5212  ( .A(n13360), .B(n12548), .Z(n12546) );
  XOR \SUBBYTES[6].a/U5211  ( .A(n13362), .B(n13361), .Z(n12547) );
  XOR \SUBBYTES[6].a/U5210  ( .A(\SUBBYTES[6].a/w1081 ), .B(
        \SUBBYTES[6].a/w1108 ), .Z(n12548) );
  XOR \SUBBYTES[6].a/U5208  ( .A(n13363), .B(n12551), .Z(n12549) );
  XOR \SUBBYTES[6].a/U5207  ( .A(\SUBBYTES[6].a/w1114 ), .B(
        \SUBBYTES[6].a/w1116 ), .Z(n12550) );
  XOR \SUBBYTES[6].a/U5206  ( .A(\SUBBYTES[6].a/w1074 ), .B(
        \SUBBYTES[6].a/w1106 ), .Z(n12551) );
  XOR \SUBBYTES[6].a/U5205  ( .A(\SUBBYTES[6].a/w906 ), .B(
        \SUBBYTES[6].a/w907 ), .Z(n13365) );
  XOR \SUBBYTES[6].a/U5204  ( .A(n13365), .B(n12552), .Z(n13364) );
  XOR \SUBBYTES[6].a/U5203  ( .A(\SUBBYTES[6].a/w899 ), .B(
        \SUBBYTES[6].a/w916 ), .Z(n12552) );
  XOR \SUBBYTES[6].a/U5201  ( .A(\SUBBYTES[6].a/w898 ), .B(
        \SUBBYTES[6].a/w913 ), .Z(n12553) );
  XOR \SUBBYTES[6].a/U5200  ( .A(n13365), .B(n12554), .Z(n13508) );
  XOR \SUBBYTES[6].a/U5199  ( .A(\SUBBYTES[6].a/w913 ), .B(
        \SUBBYTES[6].a/w914 ), .Z(n12554) );
  XOR \SUBBYTES[6].a/U5198  ( .A(\SUBBYTES[6].a/w875 ), .B(n12555), .Z(n13367)
         );
  XOR \SUBBYTES[6].a/U5197  ( .A(\SUBBYTES[6].a/w866 ), .B(
        \SUBBYTES[6].a/w867 ), .Z(n12555) );
  XOR \SUBBYTES[6].a/U5195  ( .A(\SUBBYTES[6].a/w877 ), .B(n13508), .Z(n12556)
         );
  XOR \SUBBYTES[6].a/U5194  ( .A(n12558), .B(n12557), .Z(n13368) );
  XOR \SUBBYTES[6].a/U5193  ( .A(n12560), .B(n12559), .Z(n12557) );
  XOR \SUBBYTES[6].a/U5192  ( .A(\SUBBYTES[6].a/w913 ), .B(
        \SUBBYTES[6].a/w914 ), .Z(n12558) );
  XOR \SUBBYTES[6].a/U5191  ( .A(\SUBBYTES[6].a/w877 ), .B(
        \SUBBYTES[6].a/w901 ), .Z(n12559) );
  XOR \SUBBYTES[6].a/U5190  ( .A(\SUBBYTES[6].a/w866 ), .B(
        \SUBBYTES[6].a/w875 ), .Z(n12560) );
  XOR \SUBBYTES[6].a/U5189  ( .A(\SUBBYTES[6].a/w898 ), .B(n12561), .Z(n13366)
         );
  XOR \SUBBYTES[6].a/U5188  ( .A(\SUBBYTES[6].a/w881 ), .B(
        \SUBBYTES[6].a/w884 ), .Z(n12561) );
  XOR \SUBBYTES[6].a/U5186  ( .A(\SUBBYTES[6].a/w869 ), .B(n13368), .Z(n12562)
         );
  XOR \SUBBYTES[6].a/U5184  ( .A(\SUBBYTES[6].a/w901 ), .B(
        \SUBBYTES[6].a/w914 ), .Z(n12563) );
  XOR \SUBBYTES[6].a/U5182  ( .A(n12567), .B(n12566), .Z(n12564) );
  XOR \SUBBYTES[6].a/U5181  ( .A(n12569), .B(n12568), .Z(n12565) );
  XOR \SUBBYTES[6].a/U5180  ( .A(\SUBBYTES[6].a/w913 ), .B(
        \SUBBYTES[6].a/w916 ), .Z(n12566) );
  XOR \SUBBYTES[6].a/U5179  ( .A(\SUBBYTES[6].a/w906 ), .B(
        \SUBBYTES[6].a/w909 ), .Z(n12567) );
  XOR \SUBBYTES[6].a/U5178  ( .A(\SUBBYTES[6].a/w881 ), .B(
        \SUBBYTES[6].a/w882 ), .Z(n12568) );
  XOR \SUBBYTES[6].a/U5177  ( .A(\SUBBYTES[6].a/w866 ), .B(
        \SUBBYTES[6].a/w869 ), .Z(n12569) );
  XOR \SUBBYTES[6].a/U5175  ( .A(n13365), .B(n12572), .Z(n12570) );
  XOR \SUBBYTES[6].a/U5174  ( .A(n13367), .B(n13366), .Z(n12571) );
  XOR \SUBBYTES[6].a/U5173  ( .A(\SUBBYTES[6].a/w874 ), .B(
        \SUBBYTES[6].a/w901 ), .Z(n12572) );
  XOR \SUBBYTES[6].a/U5171  ( .A(n13368), .B(n12575), .Z(n12573) );
  XOR \SUBBYTES[6].a/U5170  ( .A(\SUBBYTES[6].a/w907 ), .B(
        \SUBBYTES[6].a/w909 ), .Z(n12574) );
  XOR \SUBBYTES[6].a/U5169  ( .A(\SUBBYTES[6].a/w867 ), .B(
        \SUBBYTES[6].a/w899 ), .Z(n12575) );
  XOR \SUBBYTES[6].a/U5168  ( .A(\SUBBYTES[6].a/w699 ), .B(
        \SUBBYTES[6].a/w700 ), .Z(n13370) );
  XOR \SUBBYTES[6].a/U5167  ( .A(n13370), .B(n12576), .Z(n13369) );
  XOR \SUBBYTES[6].a/U5166  ( .A(\SUBBYTES[6].a/w692 ), .B(
        \SUBBYTES[6].a/w709 ), .Z(n12576) );
  XOR \SUBBYTES[6].a/U5164  ( .A(\SUBBYTES[6].a/w691 ), .B(
        \SUBBYTES[6].a/w706 ), .Z(n12577) );
  XOR \SUBBYTES[6].a/U5163  ( .A(n13370), .B(n12578), .Z(n13509) );
  XOR \SUBBYTES[6].a/U5162  ( .A(\SUBBYTES[6].a/w706 ), .B(
        \SUBBYTES[6].a/w707 ), .Z(n12578) );
  XOR \SUBBYTES[6].a/U5161  ( .A(\SUBBYTES[6].a/w668 ), .B(n12579), .Z(n13372)
         );
  XOR \SUBBYTES[6].a/U5160  ( .A(\SUBBYTES[6].a/w659 ), .B(
        \SUBBYTES[6].a/w660 ), .Z(n12579) );
  XOR \SUBBYTES[6].a/U5158  ( .A(\SUBBYTES[6].a/w670 ), .B(n13509), .Z(n12580)
         );
  XOR \SUBBYTES[6].a/U5157  ( .A(n12582), .B(n12581), .Z(n13373) );
  XOR \SUBBYTES[6].a/U5156  ( .A(n12584), .B(n12583), .Z(n12581) );
  XOR \SUBBYTES[6].a/U5155  ( .A(\SUBBYTES[6].a/w706 ), .B(
        \SUBBYTES[6].a/w707 ), .Z(n12582) );
  XOR \SUBBYTES[6].a/U5154  ( .A(\SUBBYTES[6].a/w670 ), .B(
        \SUBBYTES[6].a/w694 ), .Z(n12583) );
  XOR \SUBBYTES[6].a/U5153  ( .A(\SUBBYTES[6].a/w659 ), .B(
        \SUBBYTES[6].a/w668 ), .Z(n12584) );
  XOR \SUBBYTES[6].a/U5152  ( .A(\SUBBYTES[6].a/w691 ), .B(n12585), .Z(n13371)
         );
  XOR \SUBBYTES[6].a/U5151  ( .A(\SUBBYTES[6].a/w674 ), .B(
        \SUBBYTES[6].a/w677 ), .Z(n12585) );
  XOR \SUBBYTES[6].a/U5149  ( .A(\SUBBYTES[6].a/w662 ), .B(n13373), .Z(n12586)
         );
  XOR \SUBBYTES[6].a/U5147  ( .A(\SUBBYTES[6].a/w694 ), .B(
        \SUBBYTES[6].a/w707 ), .Z(n12587) );
  XOR \SUBBYTES[6].a/U5145  ( .A(n12591), .B(n12590), .Z(n12588) );
  XOR \SUBBYTES[6].a/U5144  ( .A(n12593), .B(n12592), .Z(n12589) );
  XOR \SUBBYTES[6].a/U5143  ( .A(\SUBBYTES[6].a/w706 ), .B(
        \SUBBYTES[6].a/w709 ), .Z(n12590) );
  XOR \SUBBYTES[6].a/U5142  ( .A(\SUBBYTES[6].a/w699 ), .B(
        \SUBBYTES[6].a/w702 ), .Z(n12591) );
  XOR \SUBBYTES[6].a/U5141  ( .A(\SUBBYTES[6].a/w674 ), .B(
        \SUBBYTES[6].a/w675 ), .Z(n12592) );
  XOR \SUBBYTES[6].a/U5140  ( .A(\SUBBYTES[6].a/w659 ), .B(
        \SUBBYTES[6].a/w662 ), .Z(n12593) );
  XOR \SUBBYTES[6].a/U5138  ( .A(n13370), .B(n12596), .Z(n12594) );
  XOR \SUBBYTES[6].a/U5137  ( .A(n13372), .B(n13371), .Z(n12595) );
  XOR \SUBBYTES[6].a/U5136  ( .A(\SUBBYTES[6].a/w667 ), .B(
        \SUBBYTES[6].a/w694 ), .Z(n12596) );
  XOR \SUBBYTES[6].a/U5134  ( .A(n13373), .B(n12599), .Z(n12597) );
  XOR \SUBBYTES[6].a/U5133  ( .A(\SUBBYTES[6].a/w700 ), .B(
        \SUBBYTES[6].a/w702 ), .Z(n12598) );
  XOR \SUBBYTES[6].a/U5132  ( .A(\SUBBYTES[6].a/w660 ), .B(
        \SUBBYTES[6].a/w692 ), .Z(n12599) );
  XOR \SUBBYTES[6].a/U5131  ( .A(\SUBBYTES[6].a/w492 ), .B(
        \SUBBYTES[6].a/w493 ), .Z(n13375) );
  XOR \SUBBYTES[6].a/U5130  ( .A(n13375), .B(n12600), .Z(n13374) );
  XOR \SUBBYTES[6].a/U5129  ( .A(\SUBBYTES[6].a/w485 ), .B(
        \SUBBYTES[6].a/w502 ), .Z(n12600) );
  XOR \SUBBYTES[6].a/U5127  ( .A(\SUBBYTES[6].a/w484 ), .B(
        \SUBBYTES[6].a/w499 ), .Z(n12601) );
  XOR \SUBBYTES[6].a/U5126  ( .A(n13375), .B(n12602), .Z(n13510) );
  XOR \SUBBYTES[6].a/U5125  ( .A(\SUBBYTES[6].a/w499 ), .B(
        \SUBBYTES[6].a/w500 ), .Z(n12602) );
  XOR \SUBBYTES[6].a/U5124  ( .A(\SUBBYTES[6].a/w461 ), .B(n12603), .Z(n13377)
         );
  XOR \SUBBYTES[6].a/U5123  ( .A(\SUBBYTES[6].a/w452 ), .B(
        \SUBBYTES[6].a/w453 ), .Z(n12603) );
  XOR \SUBBYTES[6].a/U5121  ( .A(\SUBBYTES[6].a/w463 ), .B(n13510), .Z(n12604)
         );
  XOR \SUBBYTES[6].a/U5120  ( .A(n12606), .B(n12605), .Z(n13378) );
  XOR \SUBBYTES[6].a/U5119  ( .A(n12608), .B(n12607), .Z(n12605) );
  XOR \SUBBYTES[6].a/U5118  ( .A(\SUBBYTES[6].a/w499 ), .B(
        \SUBBYTES[6].a/w500 ), .Z(n12606) );
  XOR \SUBBYTES[6].a/U5117  ( .A(\SUBBYTES[6].a/w463 ), .B(
        \SUBBYTES[6].a/w487 ), .Z(n12607) );
  XOR \SUBBYTES[6].a/U5116  ( .A(\SUBBYTES[6].a/w452 ), .B(
        \SUBBYTES[6].a/w461 ), .Z(n12608) );
  XOR \SUBBYTES[6].a/U5115  ( .A(\SUBBYTES[6].a/w484 ), .B(n12609), .Z(n13376)
         );
  XOR \SUBBYTES[6].a/U5114  ( .A(\SUBBYTES[6].a/w467 ), .B(
        \SUBBYTES[6].a/w470 ), .Z(n12609) );
  XOR \SUBBYTES[6].a/U5112  ( .A(\SUBBYTES[6].a/w455 ), .B(n13378), .Z(n12610)
         );
  XOR \SUBBYTES[6].a/U5110  ( .A(\SUBBYTES[6].a/w487 ), .B(
        \SUBBYTES[6].a/w500 ), .Z(n12611) );
  XOR \SUBBYTES[6].a/U5108  ( .A(n12615), .B(n12614), .Z(n12612) );
  XOR \SUBBYTES[6].a/U5107  ( .A(n12617), .B(n12616), .Z(n12613) );
  XOR \SUBBYTES[6].a/U5106  ( .A(\SUBBYTES[6].a/w499 ), .B(
        \SUBBYTES[6].a/w502 ), .Z(n12614) );
  XOR \SUBBYTES[6].a/U5105  ( .A(\SUBBYTES[6].a/w492 ), .B(
        \SUBBYTES[6].a/w495 ), .Z(n12615) );
  XOR \SUBBYTES[6].a/U5104  ( .A(\SUBBYTES[6].a/w467 ), .B(
        \SUBBYTES[6].a/w468 ), .Z(n12616) );
  XOR \SUBBYTES[6].a/U5103  ( .A(\SUBBYTES[6].a/w452 ), .B(
        \SUBBYTES[6].a/w455 ), .Z(n12617) );
  XOR \SUBBYTES[6].a/U5101  ( .A(n13375), .B(n12620), .Z(n12618) );
  XOR \SUBBYTES[6].a/U5100  ( .A(n13377), .B(n13376), .Z(n12619) );
  XOR \SUBBYTES[6].a/U5099  ( .A(\SUBBYTES[6].a/w460 ), .B(
        \SUBBYTES[6].a/w487 ), .Z(n12620) );
  XOR \SUBBYTES[6].a/U5097  ( .A(n13378), .B(n12623), .Z(n12621) );
  XOR \SUBBYTES[6].a/U5096  ( .A(\SUBBYTES[6].a/w493 ), .B(
        \SUBBYTES[6].a/w495 ), .Z(n12622) );
  XOR \SUBBYTES[6].a/U5095  ( .A(\SUBBYTES[6].a/w453 ), .B(
        \SUBBYTES[6].a/w485 ), .Z(n12623) );
  XOR \SUBBYTES[6].a/U5094  ( .A(\SUBBYTES[6].a/w285 ), .B(
        \SUBBYTES[6].a/w286 ), .Z(n13380) );
  XOR \SUBBYTES[6].a/U5093  ( .A(n13380), .B(n12624), .Z(n13379) );
  XOR \SUBBYTES[6].a/U5092  ( .A(\SUBBYTES[6].a/w278 ), .B(
        \SUBBYTES[6].a/w295 ), .Z(n12624) );
  XOR \SUBBYTES[6].a/U5090  ( .A(\SUBBYTES[6].a/w277 ), .B(
        \SUBBYTES[6].a/w292 ), .Z(n12625) );
  XOR \SUBBYTES[6].a/U5089  ( .A(n13380), .B(n12626), .Z(n13511) );
  XOR \SUBBYTES[6].a/U5088  ( .A(\SUBBYTES[6].a/w292 ), .B(
        \SUBBYTES[6].a/w293 ), .Z(n12626) );
  XOR \SUBBYTES[6].a/U5087  ( .A(\SUBBYTES[6].a/w254 ), .B(n12627), .Z(n13382)
         );
  XOR \SUBBYTES[6].a/U5086  ( .A(\SUBBYTES[6].a/w245 ), .B(
        \SUBBYTES[6].a/w246 ), .Z(n12627) );
  XOR \SUBBYTES[6].a/U5084  ( .A(\SUBBYTES[6].a/w256 ), .B(n13511), .Z(n12628)
         );
  XOR \SUBBYTES[6].a/U5083  ( .A(n12630), .B(n12629), .Z(n13383) );
  XOR \SUBBYTES[6].a/U5082  ( .A(n12632), .B(n12631), .Z(n12629) );
  XOR \SUBBYTES[6].a/U5081  ( .A(\SUBBYTES[6].a/w292 ), .B(
        \SUBBYTES[6].a/w293 ), .Z(n12630) );
  XOR \SUBBYTES[6].a/U5080  ( .A(\SUBBYTES[6].a/w256 ), .B(
        \SUBBYTES[6].a/w280 ), .Z(n12631) );
  XOR \SUBBYTES[6].a/U5079  ( .A(\SUBBYTES[6].a/w245 ), .B(
        \SUBBYTES[6].a/w254 ), .Z(n12632) );
  XOR \SUBBYTES[6].a/U5078  ( .A(\SUBBYTES[6].a/w277 ), .B(n12633), .Z(n13381)
         );
  XOR \SUBBYTES[6].a/U5077  ( .A(\SUBBYTES[6].a/w260 ), .B(
        \SUBBYTES[6].a/w263 ), .Z(n12633) );
  XOR \SUBBYTES[6].a/U5075  ( .A(\SUBBYTES[6].a/w248 ), .B(n13383), .Z(n12634)
         );
  XOR \SUBBYTES[6].a/U5073  ( .A(\SUBBYTES[6].a/w280 ), .B(
        \SUBBYTES[6].a/w293 ), .Z(n12635) );
  XOR \SUBBYTES[6].a/U5071  ( .A(n12639), .B(n12638), .Z(n12636) );
  XOR \SUBBYTES[6].a/U5070  ( .A(n12641), .B(n12640), .Z(n12637) );
  XOR \SUBBYTES[6].a/U5069  ( .A(\SUBBYTES[6].a/w292 ), .B(
        \SUBBYTES[6].a/w295 ), .Z(n12638) );
  XOR \SUBBYTES[6].a/U5068  ( .A(\SUBBYTES[6].a/w285 ), .B(
        \SUBBYTES[6].a/w288 ), .Z(n12639) );
  XOR \SUBBYTES[6].a/U5067  ( .A(\SUBBYTES[6].a/w260 ), .B(
        \SUBBYTES[6].a/w261 ), .Z(n12640) );
  XOR \SUBBYTES[6].a/U5066  ( .A(\SUBBYTES[6].a/w245 ), .B(
        \SUBBYTES[6].a/w248 ), .Z(n12641) );
  XOR \SUBBYTES[6].a/U5064  ( .A(n13380), .B(n12644), .Z(n12642) );
  XOR \SUBBYTES[6].a/U5063  ( .A(n13382), .B(n13381), .Z(n12643) );
  XOR \SUBBYTES[6].a/U5062  ( .A(\SUBBYTES[6].a/w253 ), .B(
        \SUBBYTES[6].a/w280 ), .Z(n12644) );
  XOR \SUBBYTES[6].a/U5060  ( .A(n13383), .B(n12647), .Z(n12645) );
  XOR \SUBBYTES[6].a/U5059  ( .A(\SUBBYTES[6].a/w286 ), .B(
        \SUBBYTES[6].a/w288 ), .Z(n12646) );
  XOR \SUBBYTES[6].a/U5058  ( .A(\SUBBYTES[6].a/w246 ), .B(
        \SUBBYTES[6].a/w278 ), .Z(n12647) );
  XOR \SUBBYTES[6].a/U5057  ( .A(\w1[6][1] ), .B(n12648), .Z(n13384) );
  XOR \SUBBYTES[6].a/U5056  ( .A(\w1[6][3] ), .B(\w1[6][2] ), .Z(n12648) );
  XOR \SUBBYTES[6].a/U5055  ( .A(\w1[6][6] ), .B(n13384), .Z(
        \SUBBYTES[6].a/w3378 ) );
  XOR \SUBBYTES[6].a/U5054  ( .A(\w1[6][0] ), .B(\SUBBYTES[6].a/w3378 ), .Z(
        \SUBBYTES[6].a/w3265 ) );
  XOR \SUBBYTES[6].a/U5053  ( .A(\w1[6][0] ), .B(n12649), .Z(
        \SUBBYTES[6].a/w3266 ) );
  XOR \SUBBYTES[6].a/U5052  ( .A(\w1[6][6] ), .B(\w1[6][5] ), .Z(n12649) );
  XOR \SUBBYTES[6].a/U5051  ( .A(\w1[6][5] ), .B(n13384), .Z(
        \SUBBYTES[6].a/w3396 ) );
  XOR \SUBBYTES[6].a/U5050  ( .A(n12651), .B(n12650), .Z(\SUBBYTES[6].a/w3389 ) );
  XOR \SUBBYTES[6].a/U5049  ( .A(\w1[6][3] ), .B(\w1[6][1] ), .Z(n12650) );
  XOR \SUBBYTES[6].a/U5048  ( .A(\w1[6][7] ), .B(\w1[6][4] ), .Z(n12651) );
  XOR \SUBBYTES[6].a/U5047  ( .A(\w1[6][0] ), .B(\SUBBYTES[6].a/w3389 ), .Z(
        \SUBBYTES[6].a/w3268 ) );
  XOR \SUBBYTES[6].a/U5046  ( .A(n12653), .B(n12652), .Z(\SUBBYTES[6].a/w3376 ) );
  XOR \SUBBYTES[6].a/U5045  ( .A(\SUBBYTES[6].a/w3337 ), .B(n1052), .Z(n12652)
         );
  XOR \SUBBYTES[6].a/U5044  ( .A(\SUBBYTES[6].a/w3330 ), .B(
        \SUBBYTES[6].a/w3333 ), .Z(n12653) );
  XOR \SUBBYTES[6].a/U5043  ( .A(n12655), .B(n12654), .Z(\SUBBYTES[6].a/w3377 ) );
  XOR \SUBBYTES[6].a/U5042  ( .A(\SUBBYTES[6].a/w3337 ), .B(n12263), .Z(n12654) );
  XOR \SUBBYTES[6].a/U5041  ( .A(\SUBBYTES[6].a/w3330 ), .B(n12262), .Z(n12655) );
  XOR \SUBBYTES[6].a/U5040  ( .A(\SUBBYTES[6].a/w3389 ), .B(n12656), .Z(
        \SUBBYTES[6].a/w3379 ) );
  XOR \SUBBYTES[6].a/U5039  ( .A(\w1[6][6] ), .B(\w1[6][5] ), .Z(n12656) );
  XOR \SUBBYTES[6].a/U5038  ( .A(n12658), .B(n12657), .Z(\SUBBYTES[6].a/w3380 ) );
  XOR \SUBBYTES[6].a/U5037  ( .A(n12263), .B(n1052), .Z(n12657) );
  XOR \SUBBYTES[6].a/U5036  ( .A(n12262), .B(\SUBBYTES[6].a/w3333 ), .Z(n12658) );
  XOR \SUBBYTES[6].a/U5035  ( .A(\w1[6][7] ), .B(\w1[6][2] ), .Z(n13390) );
  XOR \SUBBYTES[6].a/U5034  ( .A(n13390), .B(n12659), .Z(\SUBBYTES[6].a/w3381 ) );
  XOR \SUBBYTES[6].a/U5033  ( .A(\w1[6][5] ), .B(\w1[6][4] ), .Z(n12659) );
  XOR \SUBBYTES[6].a/U5032  ( .A(\w1[6][7] ), .B(\SUBBYTES[6].a/w3266 ), .Z(
        \SUBBYTES[6].a/w3269 ) );
  XOR \SUBBYTES[6].a/U5031  ( .A(\w1[6][1] ), .B(\SUBBYTES[6].a/w3266 ), .Z(
        \SUBBYTES[6].a/w3270 ) );
  XOR \SUBBYTES[6].a/U5030  ( .A(\w1[6][4] ), .B(\SUBBYTES[6].a/w3266 ), .Z(
        \SUBBYTES[6].a/w3271 ) );
  XOR \SUBBYTES[6].a/U5029  ( .A(\SUBBYTES[6].a/w3270 ), .B(n13390), .Z(
        \SUBBYTES[6].a/w3272 ) );
  XOR \SUBBYTES[6].a/U5028  ( .A(n13390), .B(n12660), .Z(\SUBBYTES[6].a/w3357 ) );
  XOR \SUBBYTES[6].a/U5027  ( .A(\w1[6][4] ), .B(\w1[6][1] ), .Z(n12660) );
  XOR \SUBBYTES[6].a/U5026  ( .A(n12662), .B(n12661), .Z(n13387) );
  XOR \SUBBYTES[6].a/U5025  ( .A(\w1[6][4] ), .B(n12663), .Z(n12661) );
  XOR \SUBBYTES[6].a/U5024  ( .A(\SUBBYTES[6].a/w3322 ), .B(\w1[6][6] ), .Z(
        n12662) );
  XOR \SUBBYTES[6].a/U5023  ( .A(\SUBBYTES[6].a/w3296 ), .B(
        \SUBBYTES[6].a/w3303 ), .Z(n12663) );
  XOR \SUBBYTES[6].a/U5022  ( .A(n12665), .B(n12664), .Z(n13385) );
  XOR \SUBBYTES[6].a/U5021  ( .A(\w1[6][1] ), .B(n12666), .Z(n12664) );
  XOR \SUBBYTES[6].a/U5020  ( .A(\SUBBYTES[6].a/w3321 ), .B(\w1[6][5] ), .Z(
        n12665) );
  XOR \SUBBYTES[6].a/U5019  ( .A(\SUBBYTES[6].a/w3297 ), .B(
        \SUBBYTES[6].a/w3304 ), .Z(n12666) );
  XOR \SUBBYTES[6].a/U5018  ( .A(n13387), .B(n13385), .Z(\SUBBYTES[6].a/w3327 ) );
  XOR \SUBBYTES[6].a/U5017  ( .A(\w1[6][5] ), .B(n12667), .Z(n13388) );
  XOR \SUBBYTES[6].a/U5016  ( .A(\SUBBYTES[6].a/w3289 ), .B(
        \SUBBYTES[6].a/w3299 ), .Z(n12667) );
  XOR \SUBBYTES[6].a/U5015  ( .A(n12669), .B(n12668), .Z(\SUBBYTES[6].a/w3314 ) );
  XOR \SUBBYTES[6].a/U5014  ( .A(n13388), .B(n12670), .Z(n12668) );
  XOR \SUBBYTES[6].a/U5013  ( .A(\w1[6][4] ), .B(\SUBBYTES[6].a/w3378 ), .Z(
        n12669) );
  XOR \SUBBYTES[6].a/U5012  ( .A(\SUBBYTES[6].a/w3291 ), .B(
        \SUBBYTES[6].a/w3296 ), .Z(n12670) );
  XOR \SUBBYTES[6].a/U5011  ( .A(n12672), .B(n12671), .Z(n13386) );
  XOR \SUBBYTES[6].a/U5010  ( .A(\SUBBYTES[6].a/w3324 ), .B(\w1[6][7] ), .Z(
        n12671) );
  XOR \SUBBYTES[6].a/U5009  ( .A(\SUBBYTES[6].a/w3299 ), .B(
        \SUBBYTES[6].a/w3306 ), .Z(n12672) );
  XOR \SUBBYTES[6].a/U5008  ( .A(n13385), .B(n13386), .Z(\SUBBYTES[6].a/w3326 ) );
  XOR \SUBBYTES[6].a/U5007  ( .A(\w1[6][3] ), .B(n12673), .Z(n13389) );
  XOR \SUBBYTES[6].a/U5006  ( .A(\SUBBYTES[6].a/w3288 ), .B(
        \SUBBYTES[6].a/w3291 ), .Z(n12673) );
  XOR \SUBBYTES[6].a/U5005  ( .A(n12675), .B(n12674), .Z(\SUBBYTES[6].a/w3315 ) );
  XOR \SUBBYTES[6].a/U5004  ( .A(n13389), .B(n12676), .Z(n12674) );
  XOR \SUBBYTES[6].a/U5003  ( .A(\w1[6][6] ), .B(\SUBBYTES[6].a/w3357 ), .Z(
        n12675) );
  XOR \SUBBYTES[6].a/U5002  ( .A(\SUBBYTES[6].a/w3296 ), .B(
        \SUBBYTES[6].a/w3297 ), .Z(n12676) );
  XOR \SUBBYTES[6].a/U5001  ( .A(n13387), .B(n13386), .Z(\SUBBYTES[6].a/w3335 ) );
  XOR \SUBBYTES[6].a/U5000  ( .A(n12678), .B(n12677), .Z(\SUBBYTES[6].a/w3336 ) );
  XOR \SUBBYTES[6].a/U4999  ( .A(\w1[6][7] ), .B(n13388), .Z(n12677) );
  XOR \SUBBYTES[6].a/U4998  ( .A(\SUBBYTES[6].a/w3288 ), .B(
        \SUBBYTES[6].a/w3297 ), .Z(n12678) );
  XOR \SUBBYTES[6].a/U4997  ( .A(n12680), .B(n12679), .Z(\SUBBYTES[6].a/w3312 ) );
  XOR \SUBBYTES[6].a/U4996  ( .A(n12682), .B(n12681), .Z(n12679) );
  XOR \SUBBYTES[6].a/U4995  ( .A(\w1[6][7] ), .B(\SUBBYTES[6].a/w3396 ), .Z(
        n12680) );
  XOR \SUBBYTES[6].a/U4994  ( .A(\SUBBYTES[6].a/w3303 ), .B(
        \SUBBYTES[6].a/w3306 ), .Z(n12681) );
  XOR \SUBBYTES[6].a/U4993  ( .A(\SUBBYTES[6].a/w3289 ), .B(
        \SUBBYTES[6].a/w3291 ), .Z(n12682) );
  XOR \SUBBYTES[6].a/U4992  ( .A(n12684), .B(n12683), .Z(\SUBBYTES[6].a/w3313 ) );
  XOR \SUBBYTES[6].a/U4991  ( .A(n13389), .B(n12685), .Z(n12683) );
  XOR \SUBBYTES[6].a/U4990  ( .A(\w1[6][5] ), .B(n13390), .Z(n12684) );
  XOR \SUBBYTES[6].a/U4989  ( .A(\SUBBYTES[6].a/w3303 ), .B(
        \SUBBYTES[6].a/w3304 ), .Z(n12685) );
  XOR \SUBBYTES[6].a/U4988  ( .A(n12687), .B(n12686), .Z(\SUBBYTES[6].a/w3329 ) );
  XOR \SUBBYTES[6].a/U4987  ( .A(\w1[6][1] ), .B(n12688), .Z(n12686) );
  XOR \SUBBYTES[6].a/U4986  ( .A(\SUBBYTES[6].a/w3304 ), .B(
        \SUBBYTES[6].a/w3306 ), .Z(n12687) );
  XOR \SUBBYTES[6].a/U4985  ( .A(\SUBBYTES[6].a/w3288 ), .B(
        \SUBBYTES[6].a/w3289 ), .Z(n12688) );
  XOR \SUBBYTES[6].a/U4984  ( .A(\w1[6][9] ), .B(n12689), .Z(n13391) );
  XOR \SUBBYTES[6].a/U4983  ( .A(\w1[6][11] ), .B(\w1[6][10] ), .Z(n12689) );
  XOR \SUBBYTES[6].a/U4982  ( .A(\w1[6][14] ), .B(n13391), .Z(
        \SUBBYTES[6].a/w3171 ) );
  XOR \SUBBYTES[6].a/U4981  ( .A(\w1[6][8] ), .B(\SUBBYTES[6].a/w3171 ), .Z(
        \SUBBYTES[6].a/w3058 ) );
  XOR \SUBBYTES[6].a/U4980  ( .A(\w1[6][8] ), .B(n12690), .Z(
        \SUBBYTES[6].a/w3059 ) );
  XOR \SUBBYTES[6].a/U4979  ( .A(\w1[6][14] ), .B(\w1[6][13] ), .Z(n12690) );
  XOR \SUBBYTES[6].a/U4978  ( .A(\w1[6][13] ), .B(n13391), .Z(
        \SUBBYTES[6].a/w3189 ) );
  XOR \SUBBYTES[6].a/U4977  ( .A(n12692), .B(n12691), .Z(\SUBBYTES[6].a/w3182 ) );
  XOR \SUBBYTES[6].a/U4976  ( .A(\w1[6][11] ), .B(\w1[6][9] ), .Z(n12691) );
  XOR \SUBBYTES[6].a/U4975  ( .A(\w1[6][15] ), .B(\w1[6][12] ), .Z(n12692) );
  XOR \SUBBYTES[6].a/U4974  ( .A(\w1[6][8] ), .B(\SUBBYTES[6].a/w3182 ), .Z(
        \SUBBYTES[6].a/w3061 ) );
  XOR \SUBBYTES[6].a/U4973  ( .A(n12694), .B(n12693), .Z(\SUBBYTES[6].a/w3169 ) );
  XOR \SUBBYTES[6].a/U4972  ( .A(\SUBBYTES[6].a/w3130 ), .B(n1051), .Z(n12693)
         );
  XOR \SUBBYTES[6].a/U4971  ( .A(\SUBBYTES[6].a/w3123 ), .B(
        \SUBBYTES[6].a/w3126 ), .Z(n12694) );
  XOR \SUBBYTES[6].a/U4970  ( .A(n12696), .B(n12695), .Z(\SUBBYTES[6].a/w3170 ) );
  XOR \SUBBYTES[6].a/U4969  ( .A(\SUBBYTES[6].a/w3130 ), .B(n12261), .Z(n12695) );
  XOR \SUBBYTES[6].a/U4968  ( .A(\SUBBYTES[6].a/w3123 ), .B(n12260), .Z(n12696) );
  XOR \SUBBYTES[6].a/U4967  ( .A(\SUBBYTES[6].a/w3182 ), .B(n12697), .Z(
        \SUBBYTES[6].a/w3172 ) );
  XOR \SUBBYTES[6].a/U4966  ( .A(\w1[6][14] ), .B(\w1[6][13] ), .Z(n12697) );
  XOR \SUBBYTES[6].a/U4965  ( .A(n12699), .B(n12698), .Z(\SUBBYTES[6].a/w3173 ) );
  XOR \SUBBYTES[6].a/U4964  ( .A(n12261), .B(n1051), .Z(n12698) );
  XOR \SUBBYTES[6].a/U4963  ( .A(n12260), .B(\SUBBYTES[6].a/w3126 ), .Z(n12699) );
  XOR \SUBBYTES[6].a/U4962  ( .A(\w1[6][15] ), .B(\w1[6][10] ), .Z(n13397) );
  XOR \SUBBYTES[6].a/U4961  ( .A(n13397), .B(n12700), .Z(\SUBBYTES[6].a/w3174 ) );
  XOR \SUBBYTES[6].a/U4960  ( .A(\w1[6][13] ), .B(\w1[6][12] ), .Z(n12700) );
  XOR \SUBBYTES[6].a/U4959  ( .A(\w1[6][15] ), .B(\SUBBYTES[6].a/w3059 ), .Z(
        \SUBBYTES[6].a/w3062 ) );
  XOR \SUBBYTES[6].a/U4958  ( .A(\w1[6][9] ), .B(\SUBBYTES[6].a/w3059 ), .Z(
        \SUBBYTES[6].a/w3063 ) );
  XOR \SUBBYTES[6].a/U4957  ( .A(\w1[6][12] ), .B(\SUBBYTES[6].a/w3059 ), .Z(
        \SUBBYTES[6].a/w3064 ) );
  XOR \SUBBYTES[6].a/U4956  ( .A(\SUBBYTES[6].a/w3063 ), .B(n13397), .Z(
        \SUBBYTES[6].a/w3065 ) );
  XOR \SUBBYTES[6].a/U4955  ( .A(n13397), .B(n12701), .Z(\SUBBYTES[6].a/w3150 ) );
  XOR \SUBBYTES[6].a/U4954  ( .A(\w1[6][12] ), .B(\w1[6][9] ), .Z(n12701) );
  XOR \SUBBYTES[6].a/U4953  ( .A(n12703), .B(n12702), .Z(n13394) );
  XOR \SUBBYTES[6].a/U4952  ( .A(\w1[6][12] ), .B(n12704), .Z(n12702) );
  XOR \SUBBYTES[6].a/U4951  ( .A(\SUBBYTES[6].a/w3115 ), .B(\w1[6][14] ), .Z(
        n12703) );
  XOR \SUBBYTES[6].a/U4950  ( .A(\SUBBYTES[6].a/w3089 ), .B(
        \SUBBYTES[6].a/w3096 ), .Z(n12704) );
  XOR \SUBBYTES[6].a/U4949  ( .A(n12706), .B(n12705), .Z(n13392) );
  XOR \SUBBYTES[6].a/U4948  ( .A(\w1[6][9] ), .B(n12707), .Z(n12705) );
  XOR \SUBBYTES[6].a/U4947  ( .A(\SUBBYTES[6].a/w3114 ), .B(\w1[6][13] ), .Z(
        n12706) );
  XOR \SUBBYTES[6].a/U4946  ( .A(\SUBBYTES[6].a/w3090 ), .B(
        \SUBBYTES[6].a/w3097 ), .Z(n12707) );
  XOR \SUBBYTES[6].a/U4945  ( .A(n13394), .B(n13392), .Z(\SUBBYTES[6].a/w3120 ) );
  XOR \SUBBYTES[6].a/U4944  ( .A(\w1[6][13] ), .B(n12708), .Z(n13395) );
  XOR \SUBBYTES[6].a/U4943  ( .A(\SUBBYTES[6].a/w3082 ), .B(
        \SUBBYTES[6].a/w3092 ), .Z(n12708) );
  XOR \SUBBYTES[6].a/U4942  ( .A(n12710), .B(n12709), .Z(\SUBBYTES[6].a/w3107 ) );
  XOR \SUBBYTES[6].a/U4941  ( .A(n13395), .B(n12711), .Z(n12709) );
  XOR \SUBBYTES[6].a/U4940  ( .A(\w1[6][12] ), .B(\SUBBYTES[6].a/w3171 ), .Z(
        n12710) );
  XOR \SUBBYTES[6].a/U4939  ( .A(\SUBBYTES[6].a/w3084 ), .B(
        \SUBBYTES[6].a/w3089 ), .Z(n12711) );
  XOR \SUBBYTES[6].a/U4938  ( .A(n12713), .B(n12712), .Z(n13393) );
  XOR \SUBBYTES[6].a/U4937  ( .A(\SUBBYTES[6].a/w3117 ), .B(\w1[6][15] ), .Z(
        n12712) );
  XOR \SUBBYTES[6].a/U4936  ( .A(\SUBBYTES[6].a/w3092 ), .B(
        \SUBBYTES[6].a/w3099 ), .Z(n12713) );
  XOR \SUBBYTES[6].a/U4935  ( .A(n13392), .B(n13393), .Z(\SUBBYTES[6].a/w3119 ) );
  XOR \SUBBYTES[6].a/U4934  ( .A(\w1[6][11] ), .B(n12714), .Z(n13396) );
  XOR \SUBBYTES[6].a/U4933  ( .A(\SUBBYTES[6].a/w3081 ), .B(
        \SUBBYTES[6].a/w3084 ), .Z(n12714) );
  XOR \SUBBYTES[6].a/U4932  ( .A(n12716), .B(n12715), .Z(\SUBBYTES[6].a/w3108 ) );
  XOR \SUBBYTES[6].a/U4931  ( .A(n13396), .B(n12717), .Z(n12715) );
  XOR \SUBBYTES[6].a/U4930  ( .A(\w1[6][14] ), .B(\SUBBYTES[6].a/w3150 ), .Z(
        n12716) );
  XOR \SUBBYTES[6].a/U4929  ( .A(\SUBBYTES[6].a/w3089 ), .B(
        \SUBBYTES[6].a/w3090 ), .Z(n12717) );
  XOR \SUBBYTES[6].a/U4928  ( .A(n13394), .B(n13393), .Z(\SUBBYTES[6].a/w3128 ) );
  XOR \SUBBYTES[6].a/U4927  ( .A(n12719), .B(n12718), .Z(\SUBBYTES[6].a/w3129 ) );
  XOR \SUBBYTES[6].a/U4926  ( .A(\w1[6][15] ), .B(n13395), .Z(n12718) );
  XOR \SUBBYTES[6].a/U4925  ( .A(\SUBBYTES[6].a/w3081 ), .B(
        \SUBBYTES[6].a/w3090 ), .Z(n12719) );
  XOR \SUBBYTES[6].a/U4924  ( .A(n12721), .B(n12720), .Z(\SUBBYTES[6].a/w3105 ) );
  XOR \SUBBYTES[6].a/U4923  ( .A(n12723), .B(n12722), .Z(n12720) );
  XOR \SUBBYTES[6].a/U4922  ( .A(\w1[6][15] ), .B(\SUBBYTES[6].a/w3189 ), .Z(
        n12721) );
  XOR \SUBBYTES[6].a/U4921  ( .A(\SUBBYTES[6].a/w3096 ), .B(
        \SUBBYTES[6].a/w3099 ), .Z(n12722) );
  XOR \SUBBYTES[6].a/U4920  ( .A(\SUBBYTES[6].a/w3082 ), .B(
        \SUBBYTES[6].a/w3084 ), .Z(n12723) );
  XOR \SUBBYTES[6].a/U4919  ( .A(n12725), .B(n12724), .Z(\SUBBYTES[6].a/w3106 ) );
  XOR \SUBBYTES[6].a/U4918  ( .A(n13396), .B(n12726), .Z(n12724) );
  XOR \SUBBYTES[6].a/U4917  ( .A(\w1[6][13] ), .B(n13397), .Z(n12725) );
  XOR \SUBBYTES[6].a/U4916  ( .A(\SUBBYTES[6].a/w3096 ), .B(
        \SUBBYTES[6].a/w3097 ), .Z(n12726) );
  XOR \SUBBYTES[6].a/U4915  ( .A(n12728), .B(n12727), .Z(\SUBBYTES[6].a/w3122 ) );
  XOR \SUBBYTES[6].a/U4914  ( .A(\w1[6][9] ), .B(n12729), .Z(n12727) );
  XOR \SUBBYTES[6].a/U4913  ( .A(\SUBBYTES[6].a/w3097 ), .B(
        \SUBBYTES[6].a/w3099 ), .Z(n12728) );
  XOR \SUBBYTES[6].a/U4912  ( .A(\SUBBYTES[6].a/w3081 ), .B(
        \SUBBYTES[6].a/w3082 ), .Z(n12729) );
  XOR \SUBBYTES[6].a/U4911  ( .A(\w1[6][17] ), .B(n12730), .Z(n13398) );
  XOR \SUBBYTES[6].a/U4910  ( .A(\w1[6][19] ), .B(\w1[6][18] ), .Z(n12730) );
  XOR \SUBBYTES[6].a/U4909  ( .A(\w1[6][22] ), .B(n13398), .Z(
        \SUBBYTES[6].a/w2964 ) );
  XOR \SUBBYTES[6].a/U4908  ( .A(\w1[6][16] ), .B(\SUBBYTES[6].a/w2964 ), .Z(
        \SUBBYTES[6].a/w2851 ) );
  XOR \SUBBYTES[6].a/U4907  ( .A(\w1[6][16] ), .B(n12731), .Z(
        \SUBBYTES[6].a/w2852 ) );
  XOR \SUBBYTES[6].a/U4906  ( .A(\w1[6][22] ), .B(\w1[6][21] ), .Z(n12731) );
  XOR \SUBBYTES[6].a/U4905  ( .A(\w1[6][21] ), .B(n13398), .Z(
        \SUBBYTES[6].a/w2982 ) );
  XOR \SUBBYTES[6].a/U4904  ( .A(n12733), .B(n12732), .Z(\SUBBYTES[6].a/w2975 ) );
  XOR \SUBBYTES[6].a/U4903  ( .A(\w1[6][19] ), .B(\w1[6][17] ), .Z(n12732) );
  XOR \SUBBYTES[6].a/U4902  ( .A(\w1[6][23] ), .B(\w1[6][20] ), .Z(n12733) );
  XOR \SUBBYTES[6].a/U4901  ( .A(\w1[6][16] ), .B(\SUBBYTES[6].a/w2975 ), .Z(
        \SUBBYTES[6].a/w2854 ) );
  XOR \SUBBYTES[6].a/U4900  ( .A(n12735), .B(n12734), .Z(\SUBBYTES[6].a/w2962 ) );
  XOR \SUBBYTES[6].a/U4899  ( .A(\SUBBYTES[6].a/w2923 ), .B(n1050), .Z(n12734)
         );
  XOR \SUBBYTES[6].a/U4898  ( .A(\SUBBYTES[6].a/w2916 ), .B(
        \SUBBYTES[6].a/w2919 ), .Z(n12735) );
  XOR \SUBBYTES[6].a/U4897  ( .A(n12737), .B(n12736), .Z(\SUBBYTES[6].a/w2963 ) );
  XOR \SUBBYTES[6].a/U4896  ( .A(\SUBBYTES[6].a/w2923 ), .B(n12259), .Z(n12736) );
  XOR \SUBBYTES[6].a/U4895  ( .A(\SUBBYTES[6].a/w2916 ), .B(n12258), .Z(n12737) );
  XOR \SUBBYTES[6].a/U4894  ( .A(\SUBBYTES[6].a/w2975 ), .B(n12738), .Z(
        \SUBBYTES[6].a/w2965 ) );
  XOR \SUBBYTES[6].a/U4893  ( .A(\w1[6][22] ), .B(\w1[6][21] ), .Z(n12738) );
  XOR \SUBBYTES[6].a/U4892  ( .A(n12740), .B(n12739), .Z(\SUBBYTES[6].a/w2966 ) );
  XOR \SUBBYTES[6].a/U4891  ( .A(n12259), .B(n1050), .Z(n12739) );
  XOR \SUBBYTES[6].a/U4890  ( .A(n12258), .B(\SUBBYTES[6].a/w2919 ), .Z(n12740) );
  XOR \SUBBYTES[6].a/U4889  ( .A(\w1[6][23] ), .B(\w1[6][18] ), .Z(n13404) );
  XOR \SUBBYTES[6].a/U4888  ( .A(n13404), .B(n12741), .Z(\SUBBYTES[6].a/w2967 ) );
  XOR \SUBBYTES[6].a/U4887  ( .A(\w1[6][21] ), .B(\w1[6][20] ), .Z(n12741) );
  XOR \SUBBYTES[6].a/U4886  ( .A(\w1[6][23] ), .B(\SUBBYTES[6].a/w2852 ), .Z(
        \SUBBYTES[6].a/w2855 ) );
  XOR \SUBBYTES[6].a/U4885  ( .A(\w1[6][17] ), .B(\SUBBYTES[6].a/w2852 ), .Z(
        \SUBBYTES[6].a/w2856 ) );
  XOR \SUBBYTES[6].a/U4884  ( .A(\w1[6][20] ), .B(\SUBBYTES[6].a/w2852 ), .Z(
        \SUBBYTES[6].a/w2857 ) );
  XOR \SUBBYTES[6].a/U4883  ( .A(\SUBBYTES[6].a/w2856 ), .B(n13404), .Z(
        \SUBBYTES[6].a/w2858 ) );
  XOR \SUBBYTES[6].a/U4882  ( .A(n13404), .B(n12742), .Z(\SUBBYTES[6].a/w2943 ) );
  XOR \SUBBYTES[6].a/U4881  ( .A(\w1[6][20] ), .B(\w1[6][17] ), .Z(n12742) );
  XOR \SUBBYTES[6].a/U4880  ( .A(n12744), .B(n12743), .Z(n13401) );
  XOR \SUBBYTES[6].a/U4879  ( .A(\w1[6][20] ), .B(n12745), .Z(n12743) );
  XOR \SUBBYTES[6].a/U4878  ( .A(\SUBBYTES[6].a/w2908 ), .B(\w1[6][22] ), .Z(
        n12744) );
  XOR \SUBBYTES[6].a/U4877  ( .A(\SUBBYTES[6].a/w2882 ), .B(
        \SUBBYTES[6].a/w2889 ), .Z(n12745) );
  XOR \SUBBYTES[6].a/U4876  ( .A(n12747), .B(n12746), .Z(n13399) );
  XOR \SUBBYTES[6].a/U4875  ( .A(\w1[6][17] ), .B(n12748), .Z(n12746) );
  XOR \SUBBYTES[6].a/U4874  ( .A(\SUBBYTES[6].a/w2907 ), .B(\w1[6][21] ), .Z(
        n12747) );
  XOR \SUBBYTES[6].a/U4873  ( .A(\SUBBYTES[6].a/w2883 ), .B(
        \SUBBYTES[6].a/w2890 ), .Z(n12748) );
  XOR \SUBBYTES[6].a/U4872  ( .A(n13401), .B(n13399), .Z(\SUBBYTES[6].a/w2913 ) );
  XOR \SUBBYTES[6].a/U4871  ( .A(\w1[6][21] ), .B(n12749), .Z(n13402) );
  XOR \SUBBYTES[6].a/U4870  ( .A(\SUBBYTES[6].a/w2875 ), .B(
        \SUBBYTES[6].a/w2885 ), .Z(n12749) );
  XOR \SUBBYTES[6].a/U4869  ( .A(n12751), .B(n12750), .Z(\SUBBYTES[6].a/w2900 ) );
  XOR \SUBBYTES[6].a/U4868  ( .A(n13402), .B(n12752), .Z(n12750) );
  XOR \SUBBYTES[6].a/U4867  ( .A(\w1[6][20] ), .B(\SUBBYTES[6].a/w2964 ), .Z(
        n12751) );
  XOR \SUBBYTES[6].a/U4866  ( .A(\SUBBYTES[6].a/w2877 ), .B(
        \SUBBYTES[6].a/w2882 ), .Z(n12752) );
  XOR \SUBBYTES[6].a/U4865  ( .A(n12754), .B(n12753), .Z(n13400) );
  XOR \SUBBYTES[6].a/U4864  ( .A(\SUBBYTES[6].a/w2910 ), .B(\w1[6][23] ), .Z(
        n12753) );
  XOR \SUBBYTES[6].a/U4863  ( .A(\SUBBYTES[6].a/w2885 ), .B(
        \SUBBYTES[6].a/w2892 ), .Z(n12754) );
  XOR \SUBBYTES[6].a/U4862  ( .A(n13399), .B(n13400), .Z(\SUBBYTES[6].a/w2912 ) );
  XOR \SUBBYTES[6].a/U4861  ( .A(\w1[6][19] ), .B(n12755), .Z(n13403) );
  XOR \SUBBYTES[6].a/U4860  ( .A(\SUBBYTES[6].a/w2874 ), .B(
        \SUBBYTES[6].a/w2877 ), .Z(n12755) );
  XOR \SUBBYTES[6].a/U4859  ( .A(n12757), .B(n12756), .Z(\SUBBYTES[6].a/w2901 ) );
  XOR \SUBBYTES[6].a/U4858  ( .A(n13403), .B(n12758), .Z(n12756) );
  XOR \SUBBYTES[6].a/U4857  ( .A(\w1[6][22] ), .B(\SUBBYTES[6].a/w2943 ), .Z(
        n12757) );
  XOR \SUBBYTES[6].a/U4856  ( .A(\SUBBYTES[6].a/w2882 ), .B(
        \SUBBYTES[6].a/w2883 ), .Z(n12758) );
  XOR \SUBBYTES[6].a/U4855  ( .A(n13401), .B(n13400), .Z(\SUBBYTES[6].a/w2921 ) );
  XOR \SUBBYTES[6].a/U4854  ( .A(n12760), .B(n12759), .Z(\SUBBYTES[6].a/w2922 ) );
  XOR \SUBBYTES[6].a/U4853  ( .A(\w1[6][23] ), .B(n13402), .Z(n12759) );
  XOR \SUBBYTES[6].a/U4852  ( .A(\SUBBYTES[6].a/w2874 ), .B(
        \SUBBYTES[6].a/w2883 ), .Z(n12760) );
  XOR \SUBBYTES[6].a/U4851  ( .A(n12762), .B(n12761), .Z(\SUBBYTES[6].a/w2898 ) );
  XOR \SUBBYTES[6].a/U4850  ( .A(n12764), .B(n12763), .Z(n12761) );
  XOR \SUBBYTES[6].a/U4849  ( .A(\w1[6][23] ), .B(\SUBBYTES[6].a/w2982 ), .Z(
        n12762) );
  XOR \SUBBYTES[6].a/U4848  ( .A(\SUBBYTES[6].a/w2889 ), .B(
        \SUBBYTES[6].a/w2892 ), .Z(n12763) );
  XOR \SUBBYTES[6].a/U4847  ( .A(\SUBBYTES[6].a/w2875 ), .B(
        \SUBBYTES[6].a/w2877 ), .Z(n12764) );
  XOR \SUBBYTES[6].a/U4846  ( .A(n12766), .B(n12765), .Z(\SUBBYTES[6].a/w2899 ) );
  XOR \SUBBYTES[6].a/U4845  ( .A(n13403), .B(n12767), .Z(n12765) );
  XOR \SUBBYTES[6].a/U4844  ( .A(\w1[6][21] ), .B(n13404), .Z(n12766) );
  XOR \SUBBYTES[6].a/U4843  ( .A(\SUBBYTES[6].a/w2889 ), .B(
        \SUBBYTES[6].a/w2890 ), .Z(n12767) );
  XOR \SUBBYTES[6].a/U4842  ( .A(n12769), .B(n12768), .Z(\SUBBYTES[6].a/w2915 ) );
  XOR \SUBBYTES[6].a/U4841  ( .A(\w1[6][17] ), .B(n12770), .Z(n12768) );
  XOR \SUBBYTES[6].a/U4840  ( .A(\SUBBYTES[6].a/w2890 ), .B(
        \SUBBYTES[6].a/w2892 ), .Z(n12769) );
  XOR \SUBBYTES[6].a/U4839  ( .A(\SUBBYTES[6].a/w2874 ), .B(
        \SUBBYTES[6].a/w2875 ), .Z(n12770) );
  XOR \SUBBYTES[6].a/U4838  ( .A(\w1[6][25] ), .B(n12771), .Z(n13405) );
  XOR \SUBBYTES[6].a/U4837  ( .A(\w1[6][27] ), .B(\w1[6][26] ), .Z(n12771) );
  XOR \SUBBYTES[6].a/U4836  ( .A(\w1[6][30] ), .B(n13405), .Z(
        \SUBBYTES[6].a/w2757 ) );
  XOR \SUBBYTES[6].a/U4835  ( .A(\w1[6][24] ), .B(\SUBBYTES[6].a/w2757 ), .Z(
        \SUBBYTES[6].a/w2644 ) );
  XOR \SUBBYTES[6].a/U4834  ( .A(\w1[6][24] ), .B(n12772), .Z(
        \SUBBYTES[6].a/w2645 ) );
  XOR \SUBBYTES[6].a/U4833  ( .A(\w1[6][30] ), .B(\w1[6][29] ), .Z(n12772) );
  XOR \SUBBYTES[6].a/U4832  ( .A(\w1[6][29] ), .B(n13405), .Z(
        \SUBBYTES[6].a/w2775 ) );
  XOR \SUBBYTES[6].a/U4831  ( .A(n12774), .B(n12773), .Z(\SUBBYTES[6].a/w2768 ) );
  XOR \SUBBYTES[6].a/U4830  ( .A(\w1[6][27] ), .B(\w1[6][25] ), .Z(n12773) );
  XOR \SUBBYTES[6].a/U4829  ( .A(\w1[6][31] ), .B(\w1[6][28] ), .Z(n12774) );
  XOR \SUBBYTES[6].a/U4828  ( .A(\w1[6][24] ), .B(\SUBBYTES[6].a/w2768 ), .Z(
        \SUBBYTES[6].a/w2647 ) );
  XOR \SUBBYTES[6].a/U4827  ( .A(n12776), .B(n12775), .Z(\SUBBYTES[6].a/w2755 ) );
  XOR \SUBBYTES[6].a/U4826  ( .A(\SUBBYTES[6].a/w2716 ), .B(n1049), .Z(n12775)
         );
  XOR \SUBBYTES[6].a/U4825  ( .A(\SUBBYTES[6].a/w2709 ), .B(
        \SUBBYTES[6].a/w2712 ), .Z(n12776) );
  XOR \SUBBYTES[6].a/U4824  ( .A(n12778), .B(n12777), .Z(\SUBBYTES[6].a/w2756 ) );
  XOR \SUBBYTES[6].a/U4823  ( .A(\SUBBYTES[6].a/w2716 ), .B(n12257), .Z(n12777) );
  XOR \SUBBYTES[6].a/U4822  ( .A(\SUBBYTES[6].a/w2709 ), .B(n12256), .Z(n12778) );
  XOR \SUBBYTES[6].a/U4821  ( .A(\SUBBYTES[6].a/w2768 ), .B(n12779), .Z(
        \SUBBYTES[6].a/w2758 ) );
  XOR \SUBBYTES[6].a/U4820  ( .A(\w1[6][30] ), .B(\w1[6][29] ), .Z(n12779) );
  XOR \SUBBYTES[6].a/U4819  ( .A(n12781), .B(n12780), .Z(\SUBBYTES[6].a/w2759 ) );
  XOR \SUBBYTES[6].a/U4818  ( .A(n12257), .B(n1049), .Z(n12780) );
  XOR \SUBBYTES[6].a/U4817  ( .A(n12256), .B(\SUBBYTES[6].a/w2712 ), .Z(n12781) );
  XOR \SUBBYTES[6].a/U4816  ( .A(\w1[6][31] ), .B(\w1[6][26] ), .Z(n13411) );
  XOR \SUBBYTES[6].a/U4815  ( .A(n13411), .B(n12782), .Z(\SUBBYTES[6].a/w2760 ) );
  XOR \SUBBYTES[6].a/U4814  ( .A(\w1[6][29] ), .B(\w1[6][28] ), .Z(n12782) );
  XOR \SUBBYTES[6].a/U4813  ( .A(\w1[6][31] ), .B(\SUBBYTES[6].a/w2645 ), .Z(
        \SUBBYTES[6].a/w2648 ) );
  XOR \SUBBYTES[6].a/U4812  ( .A(\w1[6][25] ), .B(\SUBBYTES[6].a/w2645 ), .Z(
        \SUBBYTES[6].a/w2649 ) );
  XOR \SUBBYTES[6].a/U4811  ( .A(\w1[6][28] ), .B(\SUBBYTES[6].a/w2645 ), .Z(
        \SUBBYTES[6].a/w2650 ) );
  XOR \SUBBYTES[6].a/U4810  ( .A(\SUBBYTES[6].a/w2649 ), .B(n13411), .Z(
        \SUBBYTES[6].a/w2651 ) );
  XOR \SUBBYTES[6].a/U4809  ( .A(n13411), .B(n12783), .Z(\SUBBYTES[6].a/w2736 ) );
  XOR \SUBBYTES[6].a/U4808  ( .A(\w1[6][28] ), .B(\w1[6][25] ), .Z(n12783) );
  XOR \SUBBYTES[6].a/U4807  ( .A(n12785), .B(n12784), .Z(n13408) );
  XOR \SUBBYTES[6].a/U4806  ( .A(\w1[6][28] ), .B(n12786), .Z(n12784) );
  XOR \SUBBYTES[6].a/U4805  ( .A(\SUBBYTES[6].a/w2701 ), .B(\w1[6][30] ), .Z(
        n12785) );
  XOR \SUBBYTES[6].a/U4804  ( .A(\SUBBYTES[6].a/w2675 ), .B(
        \SUBBYTES[6].a/w2682 ), .Z(n12786) );
  XOR \SUBBYTES[6].a/U4803  ( .A(n12788), .B(n12787), .Z(n13406) );
  XOR \SUBBYTES[6].a/U4802  ( .A(\w1[6][25] ), .B(n12789), .Z(n12787) );
  XOR \SUBBYTES[6].a/U4801  ( .A(\SUBBYTES[6].a/w2700 ), .B(\w1[6][29] ), .Z(
        n12788) );
  XOR \SUBBYTES[6].a/U4800  ( .A(\SUBBYTES[6].a/w2676 ), .B(
        \SUBBYTES[6].a/w2683 ), .Z(n12789) );
  XOR \SUBBYTES[6].a/U4799  ( .A(n13408), .B(n13406), .Z(\SUBBYTES[6].a/w2706 ) );
  XOR \SUBBYTES[6].a/U4798  ( .A(\w1[6][29] ), .B(n12790), .Z(n13409) );
  XOR \SUBBYTES[6].a/U4797  ( .A(\SUBBYTES[6].a/w2668 ), .B(
        \SUBBYTES[6].a/w2678 ), .Z(n12790) );
  XOR \SUBBYTES[6].a/U4796  ( .A(n12792), .B(n12791), .Z(\SUBBYTES[6].a/w2693 ) );
  XOR \SUBBYTES[6].a/U4795  ( .A(n13409), .B(n12793), .Z(n12791) );
  XOR \SUBBYTES[6].a/U4794  ( .A(\w1[6][28] ), .B(\SUBBYTES[6].a/w2757 ), .Z(
        n12792) );
  XOR \SUBBYTES[6].a/U4793  ( .A(\SUBBYTES[6].a/w2670 ), .B(
        \SUBBYTES[6].a/w2675 ), .Z(n12793) );
  XOR \SUBBYTES[6].a/U4792  ( .A(n12795), .B(n12794), .Z(n13407) );
  XOR \SUBBYTES[6].a/U4791  ( .A(\SUBBYTES[6].a/w2703 ), .B(\w1[6][31] ), .Z(
        n12794) );
  XOR \SUBBYTES[6].a/U4790  ( .A(\SUBBYTES[6].a/w2678 ), .B(
        \SUBBYTES[6].a/w2685 ), .Z(n12795) );
  XOR \SUBBYTES[6].a/U4789  ( .A(n13406), .B(n13407), .Z(\SUBBYTES[6].a/w2705 ) );
  XOR \SUBBYTES[6].a/U4788  ( .A(\w1[6][27] ), .B(n12796), .Z(n13410) );
  XOR \SUBBYTES[6].a/U4787  ( .A(\SUBBYTES[6].a/w2667 ), .B(
        \SUBBYTES[6].a/w2670 ), .Z(n12796) );
  XOR \SUBBYTES[6].a/U4786  ( .A(n12798), .B(n12797), .Z(\SUBBYTES[6].a/w2694 ) );
  XOR \SUBBYTES[6].a/U4785  ( .A(n13410), .B(n12799), .Z(n12797) );
  XOR \SUBBYTES[6].a/U4784  ( .A(\w1[6][30] ), .B(\SUBBYTES[6].a/w2736 ), .Z(
        n12798) );
  XOR \SUBBYTES[6].a/U4783  ( .A(\SUBBYTES[6].a/w2675 ), .B(
        \SUBBYTES[6].a/w2676 ), .Z(n12799) );
  XOR \SUBBYTES[6].a/U4782  ( .A(n13408), .B(n13407), .Z(\SUBBYTES[6].a/w2714 ) );
  XOR \SUBBYTES[6].a/U4781  ( .A(n12801), .B(n12800), .Z(\SUBBYTES[6].a/w2715 ) );
  XOR \SUBBYTES[6].a/U4780  ( .A(\w1[6][31] ), .B(n13409), .Z(n12800) );
  XOR \SUBBYTES[6].a/U4779  ( .A(\SUBBYTES[6].a/w2667 ), .B(
        \SUBBYTES[6].a/w2676 ), .Z(n12801) );
  XOR \SUBBYTES[6].a/U4778  ( .A(n12803), .B(n12802), .Z(\SUBBYTES[6].a/w2691 ) );
  XOR \SUBBYTES[6].a/U4777  ( .A(n12805), .B(n12804), .Z(n12802) );
  XOR \SUBBYTES[6].a/U4776  ( .A(\w1[6][31] ), .B(\SUBBYTES[6].a/w2775 ), .Z(
        n12803) );
  XOR \SUBBYTES[6].a/U4775  ( .A(\SUBBYTES[6].a/w2682 ), .B(
        \SUBBYTES[6].a/w2685 ), .Z(n12804) );
  XOR \SUBBYTES[6].a/U4774  ( .A(\SUBBYTES[6].a/w2668 ), .B(
        \SUBBYTES[6].a/w2670 ), .Z(n12805) );
  XOR \SUBBYTES[6].a/U4773  ( .A(n12807), .B(n12806), .Z(\SUBBYTES[6].a/w2692 ) );
  XOR \SUBBYTES[6].a/U4772  ( .A(n13410), .B(n12808), .Z(n12806) );
  XOR \SUBBYTES[6].a/U4771  ( .A(\w1[6][29] ), .B(n13411), .Z(n12807) );
  XOR \SUBBYTES[6].a/U4770  ( .A(\SUBBYTES[6].a/w2682 ), .B(
        \SUBBYTES[6].a/w2683 ), .Z(n12808) );
  XOR \SUBBYTES[6].a/U4769  ( .A(n12810), .B(n12809), .Z(\SUBBYTES[6].a/w2708 ) );
  XOR \SUBBYTES[6].a/U4768  ( .A(\w1[6][25] ), .B(n12811), .Z(n12809) );
  XOR \SUBBYTES[6].a/U4767  ( .A(\SUBBYTES[6].a/w2683 ), .B(
        \SUBBYTES[6].a/w2685 ), .Z(n12810) );
  XOR \SUBBYTES[6].a/U4766  ( .A(\SUBBYTES[6].a/w2667 ), .B(
        \SUBBYTES[6].a/w2668 ), .Z(n12811) );
  XOR \SUBBYTES[6].a/U4765  ( .A(\w1[6][33] ), .B(n12812), .Z(n13412) );
  XOR \SUBBYTES[6].a/U4764  ( .A(\w1[6][35] ), .B(\w1[6][34] ), .Z(n12812) );
  XOR \SUBBYTES[6].a/U4763  ( .A(\w1[6][38] ), .B(n13412), .Z(
        \SUBBYTES[6].a/w2550 ) );
  XOR \SUBBYTES[6].a/U4762  ( .A(\w1[6][32] ), .B(\SUBBYTES[6].a/w2550 ), .Z(
        \SUBBYTES[6].a/w2437 ) );
  XOR \SUBBYTES[6].a/U4761  ( .A(\w1[6][32] ), .B(n12813), .Z(
        \SUBBYTES[6].a/w2438 ) );
  XOR \SUBBYTES[6].a/U4760  ( .A(\w1[6][38] ), .B(\w1[6][37] ), .Z(n12813) );
  XOR \SUBBYTES[6].a/U4759  ( .A(\w1[6][37] ), .B(n13412), .Z(
        \SUBBYTES[6].a/w2568 ) );
  XOR \SUBBYTES[6].a/U4758  ( .A(n12815), .B(n12814), .Z(\SUBBYTES[6].a/w2561 ) );
  XOR \SUBBYTES[6].a/U4757  ( .A(\w1[6][35] ), .B(\w1[6][33] ), .Z(n12814) );
  XOR \SUBBYTES[6].a/U4756  ( .A(\w1[6][39] ), .B(\w1[6][36] ), .Z(n12815) );
  XOR \SUBBYTES[6].a/U4755  ( .A(\w1[6][32] ), .B(\SUBBYTES[6].a/w2561 ), .Z(
        \SUBBYTES[6].a/w2440 ) );
  XOR \SUBBYTES[6].a/U4754  ( .A(n12817), .B(n12816), .Z(\SUBBYTES[6].a/w2548 ) );
  XOR \SUBBYTES[6].a/U4753  ( .A(\SUBBYTES[6].a/w2509 ), .B(n1048), .Z(n12816)
         );
  XOR \SUBBYTES[6].a/U4752  ( .A(\SUBBYTES[6].a/w2502 ), .B(
        \SUBBYTES[6].a/w2505 ), .Z(n12817) );
  XOR \SUBBYTES[6].a/U4751  ( .A(n12819), .B(n12818), .Z(\SUBBYTES[6].a/w2549 ) );
  XOR \SUBBYTES[6].a/U4750  ( .A(\SUBBYTES[6].a/w2509 ), .B(n12255), .Z(n12818) );
  XOR \SUBBYTES[6].a/U4749  ( .A(\SUBBYTES[6].a/w2502 ), .B(n12254), .Z(n12819) );
  XOR \SUBBYTES[6].a/U4748  ( .A(\SUBBYTES[6].a/w2561 ), .B(n12820), .Z(
        \SUBBYTES[6].a/w2551 ) );
  XOR \SUBBYTES[6].a/U4747  ( .A(\w1[6][38] ), .B(\w1[6][37] ), .Z(n12820) );
  XOR \SUBBYTES[6].a/U4746  ( .A(n12822), .B(n12821), .Z(\SUBBYTES[6].a/w2552 ) );
  XOR \SUBBYTES[6].a/U4745  ( .A(n12255), .B(n1048), .Z(n12821) );
  XOR \SUBBYTES[6].a/U4744  ( .A(n12254), .B(\SUBBYTES[6].a/w2505 ), .Z(n12822) );
  XOR \SUBBYTES[6].a/U4743  ( .A(\w1[6][39] ), .B(\w1[6][34] ), .Z(n13418) );
  XOR \SUBBYTES[6].a/U4742  ( .A(n13418), .B(n12823), .Z(\SUBBYTES[6].a/w2553 ) );
  XOR \SUBBYTES[6].a/U4741  ( .A(\w1[6][37] ), .B(\w1[6][36] ), .Z(n12823) );
  XOR \SUBBYTES[6].a/U4740  ( .A(\w1[6][39] ), .B(\SUBBYTES[6].a/w2438 ), .Z(
        \SUBBYTES[6].a/w2441 ) );
  XOR \SUBBYTES[6].a/U4739  ( .A(\w1[6][33] ), .B(\SUBBYTES[6].a/w2438 ), .Z(
        \SUBBYTES[6].a/w2442 ) );
  XOR \SUBBYTES[6].a/U4738  ( .A(\w1[6][36] ), .B(\SUBBYTES[6].a/w2438 ), .Z(
        \SUBBYTES[6].a/w2443 ) );
  XOR \SUBBYTES[6].a/U4737  ( .A(\SUBBYTES[6].a/w2442 ), .B(n13418), .Z(
        \SUBBYTES[6].a/w2444 ) );
  XOR \SUBBYTES[6].a/U4736  ( .A(n13418), .B(n12824), .Z(\SUBBYTES[6].a/w2529 ) );
  XOR \SUBBYTES[6].a/U4735  ( .A(\w1[6][36] ), .B(\w1[6][33] ), .Z(n12824) );
  XOR \SUBBYTES[6].a/U4734  ( .A(n12826), .B(n12825), .Z(n13415) );
  XOR \SUBBYTES[6].a/U4733  ( .A(\w1[6][36] ), .B(n12827), .Z(n12825) );
  XOR \SUBBYTES[6].a/U4732  ( .A(\SUBBYTES[6].a/w2494 ), .B(\w1[6][38] ), .Z(
        n12826) );
  XOR \SUBBYTES[6].a/U4731  ( .A(\SUBBYTES[6].a/w2468 ), .B(
        \SUBBYTES[6].a/w2475 ), .Z(n12827) );
  XOR \SUBBYTES[6].a/U4730  ( .A(n12829), .B(n12828), .Z(n13413) );
  XOR \SUBBYTES[6].a/U4729  ( .A(\w1[6][33] ), .B(n12830), .Z(n12828) );
  XOR \SUBBYTES[6].a/U4728  ( .A(\SUBBYTES[6].a/w2493 ), .B(\w1[6][37] ), .Z(
        n12829) );
  XOR \SUBBYTES[6].a/U4727  ( .A(\SUBBYTES[6].a/w2469 ), .B(
        \SUBBYTES[6].a/w2476 ), .Z(n12830) );
  XOR \SUBBYTES[6].a/U4726  ( .A(n13415), .B(n13413), .Z(\SUBBYTES[6].a/w2499 ) );
  XOR \SUBBYTES[6].a/U4725  ( .A(\w1[6][37] ), .B(n12831), .Z(n13416) );
  XOR \SUBBYTES[6].a/U4724  ( .A(\SUBBYTES[6].a/w2461 ), .B(
        \SUBBYTES[6].a/w2471 ), .Z(n12831) );
  XOR \SUBBYTES[6].a/U4723  ( .A(n12833), .B(n12832), .Z(\SUBBYTES[6].a/w2486 ) );
  XOR \SUBBYTES[6].a/U4722  ( .A(n13416), .B(n12834), .Z(n12832) );
  XOR \SUBBYTES[6].a/U4721  ( .A(\w1[6][36] ), .B(\SUBBYTES[6].a/w2550 ), .Z(
        n12833) );
  XOR \SUBBYTES[6].a/U4720  ( .A(\SUBBYTES[6].a/w2463 ), .B(
        \SUBBYTES[6].a/w2468 ), .Z(n12834) );
  XOR \SUBBYTES[6].a/U4719  ( .A(n12836), .B(n12835), .Z(n13414) );
  XOR \SUBBYTES[6].a/U4718  ( .A(\SUBBYTES[6].a/w2496 ), .B(\w1[6][39] ), .Z(
        n12835) );
  XOR \SUBBYTES[6].a/U4717  ( .A(\SUBBYTES[6].a/w2471 ), .B(
        \SUBBYTES[6].a/w2478 ), .Z(n12836) );
  XOR \SUBBYTES[6].a/U4716  ( .A(n13413), .B(n13414), .Z(\SUBBYTES[6].a/w2498 ) );
  XOR \SUBBYTES[6].a/U4715  ( .A(\w1[6][35] ), .B(n12837), .Z(n13417) );
  XOR \SUBBYTES[6].a/U4714  ( .A(\SUBBYTES[6].a/w2460 ), .B(
        \SUBBYTES[6].a/w2463 ), .Z(n12837) );
  XOR \SUBBYTES[6].a/U4713  ( .A(n12839), .B(n12838), .Z(\SUBBYTES[6].a/w2487 ) );
  XOR \SUBBYTES[6].a/U4712  ( .A(n13417), .B(n12840), .Z(n12838) );
  XOR \SUBBYTES[6].a/U4711  ( .A(\w1[6][38] ), .B(\SUBBYTES[6].a/w2529 ), .Z(
        n12839) );
  XOR \SUBBYTES[6].a/U4710  ( .A(\SUBBYTES[6].a/w2468 ), .B(
        \SUBBYTES[6].a/w2469 ), .Z(n12840) );
  XOR \SUBBYTES[6].a/U4709  ( .A(n13415), .B(n13414), .Z(\SUBBYTES[6].a/w2507 ) );
  XOR \SUBBYTES[6].a/U4708  ( .A(n12842), .B(n12841), .Z(\SUBBYTES[6].a/w2508 ) );
  XOR \SUBBYTES[6].a/U4707  ( .A(\w1[6][39] ), .B(n13416), .Z(n12841) );
  XOR \SUBBYTES[6].a/U4706  ( .A(\SUBBYTES[6].a/w2460 ), .B(
        \SUBBYTES[6].a/w2469 ), .Z(n12842) );
  XOR \SUBBYTES[6].a/U4705  ( .A(n12844), .B(n12843), .Z(\SUBBYTES[6].a/w2484 ) );
  XOR \SUBBYTES[6].a/U4704  ( .A(n12846), .B(n12845), .Z(n12843) );
  XOR \SUBBYTES[6].a/U4703  ( .A(\w1[6][39] ), .B(\SUBBYTES[6].a/w2568 ), .Z(
        n12844) );
  XOR \SUBBYTES[6].a/U4702  ( .A(\SUBBYTES[6].a/w2475 ), .B(
        \SUBBYTES[6].a/w2478 ), .Z(n12845) );
  XOR \SUBBYTES[6].a/U4701  ( .A(\SUBBYTES[6].a/w2461 ), .B(
        \SUBBYTES[6].a/w2463 ), .Z(n12846) );
  XOR \SUBBYTES[6].a/U4700  ( .A(n12848), .B(n12847), .Z(\SUBBYTES[6].a/w2485 ) );
  XOR \SUBBYTES[6].a/U4699  ( .A(n13417), .B(n12849), .Z(n12847) );
  XOR \SUBBYTES[6].a/U4698  ( .A(\w1[6][37] ), .B(n13418), .Z(n12848) );
  XOR \SUBBYTES[6].a/U4697  ( .A(\SUBBYTES[6].a/w2475 ), .B(
        \SUBBYTES[6].a/w2476 ), .Z(n12849) );
  XOR \SUBBYTES[6].a/U4696  ( .A(n12851), .B(n12850), .Z(\SUBBYTES[6].a/w2501 ) );
  XOR \SUBBYTES[6].a/U4695  ( .A(\w1[6][33] ), .B(n12852), .Z(n12850) );
  XOR \SUBBYTES[6].a/U4694  ( .A(\SUBBYTES[6].a/w2476 ), .B(
        \SUBBYTES[6].a/w2478 ), .Z(n12851) );
  XOR \SUBBYTES[6].a/U4693  ( .A(\SUBBYTES[6].a/w2460 ), .B(
        \SUBBYTES[6].a/w2461 ), .Z(n12852) );
  XOR \SUBBYTES[6].a/U4692  ( .A(\w1[6][41] ), .B(n12853), .Z(n13419) );
  XOR \SUBBYTES[6].a/U4691  ( .A(\w1[6][43] ), .B(\w1[6][42] ), .Z(n12853) );
  XOR \SUBBYTES[6].a/U4690  ( .A(\w1[6][46] ), .B(n13419), .Z(
        \SUBBYTES[6].a/w2343 ) );
  XOR \SUBBYTES[6].a/U4689  ( .A(\w1[6][40] ), .B(\SUBBYTES[6].a/w2343 ), .Z(
        \SUBBYTES[6].a/w2230 ) );
  XOR \SUBBYTES[6].a/U4688  ( .A(\w1[6][40] ), .B(n12854), .Z(
        \SUBBYTES[6].a/w2231 ) );
  XOR \SUBBYTES[6].a/U4687  ( .A(\w1[6][46] ), .B(\w1[6][45] ), .Z(n12854) );
  XOR \SUBBYTES[6].a/U4686  ( .A(\w1[6][45] ), .B(n13419), .Z(
        \SUBBYTES[6].a/w2361 ) );
  XOR \SUBBYTES[6].a/U4685  ( .A(n12856), .B(n12855), .Z(\SUBBYTES[6].a/w2354 ) );
  XOR \SUBBYTES[6].a/U4684  ( .A(\w1[6][43] ), .B(\w1[6][41] ), .Z(n12855) );
  XOR \SUBBYTES[6].a/U4683  ( .A(\w1[6][47] ), .B(\w1[6][44] ), .Z(n12856) );
  XOR \SUBBYTES[6].a/U4682  ( .A(\w1[6][40] ), .B(\SUBBYTES[6].a/w2354 ), .Z(
        \SUBBYTES[6].a/w2233 ) );
  XOR \SUBBYTES[6].a/U4681  ( .A(n12858), .B(n12857), .Z(\SUBBYTES[6].a/w2341 ) );
  XOR \SUBBYTES[6].a/U4680  ( .A(\SUBBYTES[6].a/w2302 ), .B(n1047), .Z(n12857)
         );
  XOR \SUBBYTES[6].a/U4679  ( .A(\SUBBYTES[6].a/w2295 ), .B(
        \SUBBYTES[6].a/w2298 ), .Z(n12858) );
  XOR \SUBBYTES[6].a/U4678  ( .A(n12860), .B(n12859), .Z(\SUBBYTES[6].a/w2342 ) );
  XOR \SUBBYTES[6].a/U4677  ( .A(\SUBBYTES[6].a/w2302 ), .B(n12253), .Z(n12859) );
  XOR \SUBBYTES[6].a/U4676  ( .A(\SUBBYTES[6].a/w2295 ), .B(n12252), .Z(n12860) );
  XOR \SUBBYTES[6].a/U4675  ( .A(\SUBBYTES[6].a/w2354 ), .B(n12861), .Z(
        \SUBBYTES[6].a/w2344 ) );
  XOR \SUBBYTES[6].a/U4674  ( .A(\w1[6][46] ), .B(\w1[6][45] ), .Z(n12861) );
  XOR \SUBBYTES[6].a/U4673  ( .A(n12863), .B(n12862), .Z(\SUBBYTES[6].a/w2345 ) );
  XOR \SUBBYTES[6].a/U4672  ( .A(n12253), .B(n1047), .Z(n12862) );
  XOR \SUBBYTES[6].a/U4671  ( .A(n12252), .B(\SUBBYTES[6].a/w2298 ), .Z(n12863) );
  XOR \SUBBYTES[6].a/U4670  ( .A(\w1[6][47] ), .B(\w1[6][42] ), .Z(n13425) );
  XOR \SUBBYTES[6].a/U4669  ( .A(n13425), .B(n12864), .Z(\SUBBYTES[6].a/w2346 ) );
  XOR \SUBBYTES[6].a/U4668  ( .A(\w1[6][45] ), .B(\w1[6][44] ), .Z(n12864) );
  XOR \SUBBYTES[6].a/U4667  ( .A(\w1[6][47] ), .B(\SUBBYTES[6].a/w2231 ), .Z(
        \SUBBYTES[6].a/w2234 ) );
  XOR \SUBBYTES[6].a/U4666  ( .A(\w1[6][41] ), .B(\SUBBYTES[6].a/w2231 ), .Z(
        \SUBBYTES[6].a/w2235 ) );
  XOR \SUBBYTES[6].a/U4665  ( .A(\w1[6][44] ), .B(\SUBBYTES[6].a/w2231 ), .Z(
        \SUBBYTES[6].a/w2236 ) );
  XOR \SUBBYTES[6].a/U4664  ( .A(\SUBBYTES[6].a/w2235 ), .B(n13425), .Z(
        \SUBBYTES[6].a/w2237 ) );
  XOR \SUBBYTES[6].a/U4663  ( .A(n13425), .B(n12865), .Z(\SUBBYTES[6].a/w2322 ) );
  XOR \SUBBYTES[6].a/U4662  ( .A(\w1[6][44] ), .B(\w1[6][41] ), .Z(n12865) );
  XOR \SUBBYTES[6].a/U4661  ( .A(n12867), .B(n12866), .Z(n13422) );
  XOR \SUBBYTES[6].a/U4660  ( .A(\w1[6][44] ), .B(n12868), .Z(n12866) );
  XOR \SUBBYTES[6].a/U4659  ( .A(\SUBBYTES[6].a/w2287 ), .B(\w1[6][46] ), .Z(
        n12867) );
  XOR \SUBBYTES[6].a/U4658  ( .A(\SUBBYTES[6].a/w2261 ), .B(
        \SUBBYTES[6].a/w2268 ), .Z(n12868) );
  XOR \SUBBYTES[6].a/U4657  ( .A(n12870), .B(n12869), .Z(n13420) );
  XOR \SUBBYTES[6].a/U4656  ( .A(\w1[6][41] ), .B(n12871), .Z(n12869) );
  XOR \SUBBYTES[6].a/U4655  ( .A(\SUBBYTES[6].a/w2286 ), .B(\w1[6][45] ), .Z(
        n12870) );
  XOR \SUBBYTES[6].a/U4654  ( .A(\SUBBYTES[6].a/w2262 ), .B(
        \SUBBYTES[6].a/w2269 ), .Z(n12871) );
  XOR \SUBBYTES[6].a/U4653  ( .A(n13422), .B(n13420), .Z(\SUBBYTES[6].a/w2292 ) );
  XOR \SUBBYTES[6].a/U4652  ( .A(\w1[6][45] ), .B(n12872), .Z(n13423) );
  XOR \SUBBYTES[6].a/U4651  ( .A(\SUBBYTES[6].a/w2254 ), .B(
        \SUBBYTES[6].a/w2264 ), .Z(n12872) );
  XOR \SUBBYTES[6].a/U4650  ( .A(n12874), .B(n12873), .Z(\SUBBYTES[6].a/w2279 ) );
  XOR \SUBBYTES[6].a/U4649  ( .A(n13423), .B(n12875), .Z(n12873) );
  XOR \SUBBYTES[6].a/U4648  ( .A(\w1[6][44] ), .B(\SUBBYTES[6].a/w2343 ), .Z(
        n12874) );
  XOR \SUBBYTES[6].a/U4647  ( .A(\SUBBYTES[6].a/w2256 ), .B(
        \SUBBYTES[6].a/w2261 ), .Z(n12875) );
  XOR \SUBBYTES[6].a/U4646  ( .A(n12877), .B(n12876), .Z(n13421) );
  XOR \SUBBYTES[6].a/U4645  ( .A(\SUBBYTES[6].a/w2289 ), .B(\w1[6][47] ), .Z(
        n12876) );
  XOR \SUBBYTES[6].a/U4644  ( .A(\SUBBYTES[6].a/w2264 ), .B(
        \SUBBYTES[6].a/w2271 ), .Z(n12877) );
  XOR \SUBBYTES[6].a/U4643  ( .A(n13420), .B(n13421), .Z(\SUBBYTES[6].a/w2291 ) );
  XOR \SUBBYTES[6].a/U4642  ( .A(\w1[6][43] ), .B(n12878), .Z(n13424) );
  XOR \SUBBYTES[6].a/U4641  ( .A(\SUBBYTES[6].a/w2253 ), .B(
        \SUBBYTES[6].a/w2256 ), .Z(n12878) );
  XOR \SUBBYTES[6].a/U4640  ( .A(n12880), .B(n12879), .Z(\SUBBYTES[6].a/w2280 ) );
  XOR \SUBBYTES[6].a/U4639  ( .A(n13424), .B(n12881), .Z(n12879) );
  XOR \SUBBYTES[6].a/U4638  ( .A(\w1[6][46] ), .B(\SUBBYTES[6].a/w2322 ), .Z(
        n12880) );
  XOR \SUBBYTES[6].a/U4637  ( .A(\SUBBYTES[6].a/w2261 ), .B(
        \SUBBYTES[6].a/w2262 ), .Z(n12881) );
  XOR \SUBBYTES[6].a/U4636  ( .A(n13422), .B(n13421), .Z(\SUBBYTES[6].a/w2300 ) );
  XOR \SUBBYTES[6].a/U4635  ( .A(n12883), .B(n12882), .Z(\SUBBYTES[6].a/w2301 ) );
  XOR \SUBBYTES[6].a/U4634  ( .A(\w1[6][47] ), .B(n13423), .Z(n12882) );
  XOR \SUBBYTES[6].a/U4633  ( .A(\SUBBYTES[6].a/w2253 ), .B(
        \SUBBYTES[6].a/w2262 ), .Z(n12883) );
  XOR \SUBBYTES[6].a/U4632  ( .A(n12885), .B(n12884), .Z(\SUBBYTES[6].a/w2277 ) );
  XOR \SUBBYTES[6].a/U4631  ( .A(n12887), .B(n12886), .Z(n12884) );
  XOR \SUBBYTES[6].a/U4630  ( .A(\w1[6][47] ), .B(\SUBBYTES[6].a/w2361 ), .Z(
        n12885) );
  XOR \SUBBYTES[6].a/U4629  ( .A(\SUBBYTES[6].a/w2268 ), .B(
        \SUBBYTES[6].a/w2271 ), .Z(n12886) );
  XOR \SUBBYTES[6].a/U4628  ( .A(\SUBBYTES[6].a/w2254 ), .B(
        \SUBBYTES[6].a/w2256 ), .Z(n12887) );
  XOR \SUBBYTES[6].a/U4627  ( .A(n12889), .B(n12888), .Z(\SUBBYTES[6].a/w2278 ) );
  XOR \SUBBYTES[6].a/U4626  ( .A(n13424), .B(n12890), .Z(n12888) );
  XOR \SUBBYTES[6].a/U4625  ( .A(\w1[6][45] ), .B(n13425), .Z(n12889) );
  XOR \SUBBYTES[6].a/U4624  ( .A(\SUBBYTES[6].a/w2268 ), .B(
        \SUBBYTES[6].a/w2269 ), .Z(n12890) );
  XOR \SUBBYTES[6].a/U4623  ( .A(n12892), .B(n12891), .Z(\SUBBYTES[6].a/w2294 ) );
  XOR \SUBBYTES[6].a/U4622  ( .A(\w1[6][41] ), .B(n12893), .Z(n12891) );
  XOR \SUBBYTES[6].a/U4621  ( .A(\SUBBYTES[6].a/w2269 ), .B(
        \SUBBYTES[6].a/w2271 ), .Z(n12892) );
  XOR \SUBBYTES[6].a/U4620  ( .A(\SUBBYTES[6].a/w2253 ), .B(
        \SUBBYTES[6].a/w2254 ), .Z(n12893) );
  XOR \SUBBYTES[6].a/U4619  ( .A(\w1[6][49] ), .B(n12894), .Z(n13426) );
  XOR \SUBBYTES[6].a/U4618  ( .A(\w1[6][51] ), .B(\w1[6][50] ), .Z(n12894) );
  XOR \SUBBYTES[6].a/U4617  ( .A(\w1[6][54] ), .B(n13426), .Z(
        \SUBBYTES[6].a/w2136 ) );
  XOR \SUBBYTES[6].a/U4616  ( .A(\w1[6][48] ), .B(\SUBBYTES[6].a/w2136 ), .Z(
        \SUBBYTES[6].a/w2023 ) );
  XOR \SUBBYTES[6].a/U4615  ( .A(\w1[6][48] ), .B(n12895), .Z(
        \SUBBYTES[6].a/w2024 ) );
  XOR \SUBBYTES[6].a/U4614  ( .A(\w1[6][54] ), .B(\w1[6][53] ), .Z(n12895) );
  XOR \SUBBYTES[6].a/U4613  ( .A(\w1[6][53] ), .B(n13426), .Z(
        \SUBBYTES[6].a/w2154 ) );
  XOR \SUBBYTES[6].a/U4612  ( .A(n12897), .B(n12896), .Z(\SUBBYTES[6].a/w2147 ) );
  XOR \SUBBYTES[6].a/U4611  ( .A(\w1[6][51] ), .B(\w1[6][49] ), .Z(n12896) );
  XOR \SUBBYTES[6].a/U4610  ( .A(\w1[6][55] ), .B(\w1[6][52] ), .Z(n12897) );
  XOR \SUBBYTES[6].a/U4609  ( .A(\w1[6][48] ), .B(\SUBBYTES[6].a/w2147 ), .Z(
        \SUBBYTES[6].a/w2026 ) );
  XOR \SUBBYTES[6].a/U4608  ( .A(n12899), .B(n12898), .Z(\SUBBYTES[6].a/w2134 ) );
  XOR \SUBBYTES[6].a/U4607  ( .A(\SUBBYTES[6].a/w2095 ), .B(n1046), .Z(n12898)
         );
  XOR \SUBBYTES[6].a/U4606  ( .A(\SUBBYTES[6].a/w2088 ), .B(
        \SUBBYTES[6].a/w2091 ), .Z(n12899) );
  XOR \SUBBYTES[6].a/U4605  ( .A(n12901), .B(n12900), .Z(\SUBBYTES[6].a/w2135 ) );
  XOR \SUBBYTES[6].a/U4604  ( .A(\SUBBYTES[6].a/w2095 ), .B(n12251), .Z(n12900) );
  XOR \SUBBYTES[6].a/U4603  ( .A(\SUBBYTES[6].a/w2088 ), .B(n12250), .Z(n12901) );
  XOR \SUBBYTES[6].a/U4602  ( .A(\SUBBYTES[6].a/w2147 ), .B(n12902), .Z(
        \SUBBYTES[6].a/w2137 ) );
  XOR \SUBBYTES[6].a/U4601  ( .A(\w1[6][54] ), .B(\w1[6][53] ), .Z(n12902) );
  XOR \SUBBYTES[6].a/U4600  ( .A(n12904), .B(n12903), .Z(\SUBBYTES[6].a/w2138 ) );
  XOR \SUBBYTES[6].a/U4599  ( .A(n12251), .B(n1046), .Z(n12903) );
  XOR \SUBBYTES[6].a/U4598  ( .A(n12250), .B(\SUBBYTES[6].a/w2091 ), .Z(n12904) );
  XOR \SUBBYTES[6].a/U4597  ( .A(\w1[6][55] ), .B(\w1[6][50] ), .Z(n13432) );
  XOR \SUBBYTES[6].a/U4596  ( .A(n13432), .B(n12905), .Z(\SUBBYTES[6].a/w2139 ) );
  XOR \SUBBYTES[6].a/U4595  ( .A(\w1[6][53] ), .B(\w1[6][52] ), .Z(n12905) );
  XOR \SUBBYTES[6].a/U4594  ( .A(\w1[6][55] ), .B(\SUBBYTES[6].a/w2024 ), .Z(
        \SUBBYTES[6].a/w2027 ) );
  XOR \SUBBYTES[6].a/U4593  ( .A(\w1[6][49] ), .B(\SUBBYTES[6].a/w2024 ), .Z(
        \SUBBYTES[6].a/w2028 ) );
  XOR \SUBBYTES[6].a/U4592  ( .A(\w1[6][52] ), .B(\SUBBYTES[6].a/w2024 ), .Z(
        \SUBBYTES[6].a/w2029 ) );
  XOR \SUBBYTES[6].a/U4591  ( .A(\SUBBYTES[6].a/w2028 ), .B(n13432), .Z(
        \SUBBYTES[6].a/w2030 ) );
  XOR \SUBBYTES[6].a/U4590  ( .A(n13432), .B(n12906), .Z(\SUBBYTES[6].a/w2115 ) );
  XOR \SUBBYTES[6].a/U4589  ( .A(\w1[6][52] ), .B(\w1[6][49] ), .Z(n12906) );
  XOR \SUBBYTES[6].a/U4588  ( .A(n12908), .B(n12907), .Z(n13429) );
  XOR \SUBBYTES[6].a/U4587  ( .A(\w1[6][52] ), .B(n12909), .Z(n12907) );
  XOR \SUBBYTES[6].a/U4586  ( .A(\SUBBYTES[6].a/w2080 ), .B(\w1[6][54] ), .Z(
        n12908) );
  XOR \SUBBYTES[6].a/U4585  ( .A(\SUBBYTES[6].a/w2054 ), .B(
        \SUBBYTES[6].a/w2061 ), .Z(n12909) );
  XOR \SUBBYTES[6].a/U4584  ( .A(n12911), .B(n12910), .Z(n13427) );
  XOR \SUBBYTES[6].a/U4583  ( .A(\w1[6][49] ), .B(n12912), .Z(n12910) );
  XOR \SUBBYTES[6].a/U4582  ( .A(\SUBBYTES[6].a/w2079 ), .B(\w1[6][53] ), .Z(
        n12911) );
  XOR \SUBBYTES[6].a/U4581  ( .A(\SUBBYTES[6].a/w2055 ), .B(
        \SUBBYTES[6].a/w2062 ), .Z(n12912) );
  XOR \SUBBYTES[6].a/U4580  ( .A(n13429), .B(n13427), .Z(\SUBBYTES[6].a/w2085 ) );
  XOR \SUBBYTES[6].a/U4579  ( .A(\w1[6][53] ), .B(n12913), .Z(n13430) );
  XOR \SUBBYTES[6].a/U4578  ( .A(\SUBBYTES[6].a/w2047 ), .B(
        \SUBBYTES[6].a/w2057 ), .Z(n12913) );
  XOR \SUBBYTES[6].a/U4577  ( .A(n12915), .B(n12914), .Z(\SUBBYTES[6].a/w2072 ) );
  XOR \SUBBYTES[6].a/U4576  ( .A(n13430), .B(n12916), .Z(n12914) );
  XOR \SUBBYTES[6].a/U4575  ( .A(\w1[6][52] ), .B(\SUBBYTES[6].a/w2136 ), .Z(
        n12915) );
  XOR \SUBBYTES[6].a/U4574  ( .A(\SUBBYTES[6].a/w2049 ), .B(
        \SUBBYTES[6].a/w2054 ), .Z(n12916) );
  XOR \SUBBYTES[6].a/U4573  ( .A(n12918), .B(n12917), .Z(n13428) );
  XOR \SUBBYTES[6].a/U4572  ( .A(\SUBBYTES[6].a/w2082 ), .B(\w1[6][55] ), .Z(
        n12917) );
  XOR \SUBBYTES[6].a/U4571  ( .A(\SUBBYTES[6].a/w2057 ), .B(
        \SUBBYTES[6].a/w2064 ), .Z(n12918) );
  XOR \SUBBYTES[6].a/U4570  ( .A(n13427), .B(n13428), .Z(\SUBBYTES[6].a/w2084 ) );
  XOR \SUBBYTES[6].a/U4569  ( .A(\w1[6][51] ), .B(n12919), .Z(n13431) );
  XOR \SUBBYTES[6].a/U4568  ( .A(\SUBBYTES[6].a/w2046 ), .B(
        \SUBBYTES[6].a/w2049 ), .Z(n12919) );
  XOR \SUBBYTES[6].a/U4567  ( .A(n12921), .B(n12920), .Z(\SUBBYTES[6].a/w2073 ) );
  XOR \SUBBYTES[6].a/U4566  ( .A(n13431), .B(n12922), .Z(n12920) );
  XOR \SUBBYTES[6].a/U4565  ( .A(\w1[6][54] ), .B(\SUBBYTES[6].a/w2115 ), .Z(
        n12921) );
  XOR \SUBBYTES[6].a/U4564  ( .A(\SUBBYTES[6].a/w2054 ), .B(
        \SUBBYTES[6].a/w2055 ), .Z(n12922) );
  XOR \SUBBYTES[6].a/U4563  ( .A(n13429), .B(n13428), .Z(\SUBBYTES[6].a/w2093 ) );
  XOR \SUBBYTES[6].a/U4562  ( .A(n12924), .B(n12923), .Z(\SUBBYTES[6].a/w2094 ) );
  XOR \SUBBYTES[6].a/U4561  ( .A(\w1[6][55] ), .B(n13430), .Z(n12923) );
  XOR \SUBBYTES[6].a/U4560  ( .A(\SUBBYTES[6].a/w2046 ), .B(
        \SUBBYTES[6].a/w2055 ), .Z(n12924) );
  XOR \SUBBYTES[6].a/U4559  ( .A(n12926), .B(n12925), .Z(\SUBBYTES[6].a/w2070 ) );
  XOR \SUBBYTES[6].a/U4558  ( .A(n12928), .B(n12927), .Z(n12925) );
  XOR \SUBBYTES[6].a/U4557  ( .A(\w1[6][55] ), .B(\SUBBYTES[6].a/w2154 ), .Z(
        n12926) );
  XOR \SUBBYTES[6].a/U4556  ( .A(\SUBBYTES[6].a/w2061 ), .B(
        \SUBBYTES[6].a/w2064 ), .Z(n12927) );
  XOR \SUBBYTES[6].a/U4555  ( .A(\SUBBYTES[6].a/w2047 ), .B(
        \SUBBYTES[6].a/w2049 ), .Z(n12928) );
  XOR \SUBBYTES[6].a/U4554  ( .A(n12930), .B(n12929), .Z(\SUBBYTES[6].a/w2071 ) );
  XOR \SUBBYTES[6].a/U4553  ( .A(n13431), .B(n12931), .Z(n12929) );
  XOR \SUBBYTES[6].a/U4552  ( .A(\w1[6][53] ), .B(n13432), .Z(n12930) );
  XOR \SUBBYTES[6].a/U4551  ( .A(\SUBBYTES[6].a/w2061 ), .B(
        \SUBBYTES[6].a/w2062 ), .Z(n12931) );
  XOR \SUBBYTES[6].a/U4550  ( .A(n12933), .B(n12932), .Z(\SUBBYTES[6].a/w2087 ) );
  XOR \SUBBYTES[6].a/U4549  ( .A(\w1[6][49] ), .B(n12934), .Z(n12932) );
  XOR \SUBBYTES[6].a/U4548  ( .A(\SUBBYTES[6].a/w2062 ), .B(
        \SUBBYTES[6].a/w2064 ), .Z(n12933) );
  XOR \SUBBYTES[6].a/U4547  ( .A(\SUBBYTES[6].a/w2046 ), .B(
        \SUBBYTES[6].a/w2047 ), .Z(n12934) );
  XOR \SUBBYTES[6].a/U4546  ( .A(\w1[6][57] ), .B(n12935), .Z(n13433) );
  XOR \SUBBYTES[6].a/U4545  ( .A(\w1[6][59] ), .B(\w1[6][58] ), .Z(n12935) );
  XOR \SUBBYTES[6].a/U4544  ( .A(\w1[6][62] ), .B(n13433), .Z(
        \SUBBYTES[6].a/w1929 ) );
  XOR \SUBBYTES[6].a/U4543  ( .A(\w1[6][56] ), .B(\SUBBYTES[6].a/w1929 ), .Z(
        \SUBBYTES[6].a/w1816 ) );
  XOR \SUBBYTES[6].a/U4542  ( .A(\w1[6][56] ), .B(n12936), .Z(
        \SUBBYTES[6].a/w1817 ) );
  XOR \SUBBYTES[6].a/U4541  ( .A(\w1[6][62] ), .B(\w1[6][61] ), .Z(n12936) );
  XOR \SUBBYTES[6].a/U4540  ( .A(\w1[6][61] ), .B(n13433), .Z(
        \SUBBYTES[6].a/w1947 ) );
  XOR \SUBBYTES[6].a/U4539  ( .A(n12938), .B(n12937), .Z(\SUBBYTES[6].a/w1940 ) );
  XOR \SUBBYTES[6].a/U4538  ( .A(\w1[6][59] ), .B(\w1[6][57] ), .Z(n12937) );
  XOR \SUBBYTES[6].a/U4537  ( .A(\w1[6][63] ), .B(\w1[6][60] ), .Z(n12938) );
  XOR \SUBBYTES[6].a/U4536  ( .A(\w1[6][56] ), .B(\SUBBYTES[6].a/w1940 ), .Z(
        \SUBBYTES[6].a/w1819 ) );
  XOR \SUBBYTES[6].a/U4535  ( .A(n12940), .B(n12939), .Z(\SUBBYTES[6].a/w1927 ) );
  XOR \SUBBYTES[6].a/U4534  ( .A(\SUBBYTES[6].a/w1888 ), .B(n1045), .Z(n12939)
         );
  XOR \SUBBYTES[6].a/U4533  ( .A(\SUBBYTES[6].a/w1881 ), .B(
        \SUBBYTES[6].a/w1884 ), .Z(n12940) );
  XOR \SUBBYTES[6].a/U4532  ( .A(n12942), .B(n12941), .Z(\SUBBYTES[6].a/w1928 ) );
  XOR \SUBBYTES[6].a/U4531  ( .A(\SUBBYTES[6].a/w1888 ), .B(n12249), .Z(n12941) );
  XOR \SUBBYTES[6].a/U4530  ( .A(\SUBBYTES[6].a/w1881 ), .B(n12248), .Z(n12942) );
  XOR \SUBBYTES[6].a/U4529  ( .A(\SUBBYTES[6].a/w1940 ), .B(n12943), .Z(
        \SUBBYTES[6].a/w1930 ) );
  XOR \SUBBYTES[6].a/U4528  ( .A(\w1[6][62] ), .B(\w1[6][61] ), .Z(n12943) );
  XOR \SUBBYTES[6].a/U4527  ( .A(n12945), .B(n12944), .Z(\SUBBYTES[6].a/w1931 ) );
  XOR \SUBBYTES[6].a/U4526  ( .A(n12249), .B(n1045), .Z(n12944) );
  XOR \SUBBYTES[6].a/U4525  ( .A(n12248), .B(\SUBBYTES[6].a/w1884 ), .Z(n12945) );
  XOR \SUBBYTES[6].a/U4524  ( .A(\w1[6][63] ), .B(\w1[6][58] ), .Z(n13439) );
  XOR \SUBBYTES[6].a/U4523  ( .A(n13439), .B(n12946), .Z(\SUBBYTES[6].a/w1932 ) );
  XOR \SUBBYTES[6].a/U4522  ( .A(\w1[6][61] ), .B(\w1[6][60] ), .Z(n12946) );
  XOR \SUBBYTES[6].a/U4521  ( .A(\w1[6][63] ), .B(\SUBBYTES[6].a/w1817 ), .Z(
        \SUBBYTES[6].a/w1820 ) );
  XOR \SUBBYTES[6].a/U4520  ( .A(\w1[6][57] ), .B(\SUBBYTES[6].a/w1817 ), .Z(
        \SUBBYTES[6].a/w1821 ) );
  XOR \SUBBYTES[6].a/U4519  ( .A(\w1[6][60] ), .B(\SUBBYTES[6].a/w1817 ), .Z(
        \SUBBYTES[6].a/w1822 ) );
  XOR \SUBBYTES[6].a/U4518  ( .A(\SUBBYTES[6].a/w1821 ), .B(n13439), .Z(
        \SUBBYTES[6].a/w1823 ) );
  XOR \SUBBYTES[6].a/U4517  ( .A(n13439), .B(n12947), .Z(\SUBBYTES[6].a/w1908 ) );
  XOR \SUBBYTES[6].a/U4516  ( .A(\w1[6][60] ), .B(\w1[6][57] ), .Z(n12947) );
  XOR \SUBBYTES[6].a/U4515  ( .A(n12949), .B(n12948), .Z(n13436) );
  XOR \SUBBYTES[6].a/U4514  ( .A(\w1[6][60] ), .B(n12950), .Z(n12948) );
  XOR \SUBBYTES[6].a/U4513  ( .A(\SUBBYTES[6].a/w1873 ), .B(\w1[6][62] ), .Z(
        n12949) );
  XOR \SUBBYTES[6].a/U4512  ( .A(\SUBBYTES[6].a/w1847 ), .B(
        \SUBBYTES[6].a/w1854 ), .Z(n12950) );
  XOR \SUBBYTES[6].a/U4511  ( .A(n12952), .B(n12951), .Z(n13434) );
  XOR \SUBBYTES[6].a/U4510  ( .A(\w1[6][57] ), .B(n12953), .Z(n12951) );
  XOR \SUBBYTES[6].a/U4509  ( .A(\SUBBYTES[6].a/w1872 ), .B(\w1[6][61] ), .Z(
        n12952) );
  XOR \SUBBYTES[6].a/U4508  ( .A(\SUBBYTES[6].a/w1848 ), .B(
        \SUBBYTES[6].a/w1855 ), .Z(n12953) );
  XOR \SUBBYTES[6].a/U4507  ( .A(n13436), .B(n13434), .Z(\SUBBYTES[6].a/w1878 ) );
  XOR \SUBBYTES[6].a/U4506  ( .A(\w1[6][61] ), .B(n12954), .Z(n13437) );
  XOR \SUBBYTES[6].a/U4505  ( .A(\SUBBYTES[6].a/w1840 ), .B(
        \SUBBYTES[6].a/w1850 ), .Z(n12954) );
  XOR \SUBBYTES[6].a/U4504  ( .A(n12956), .B(n12955), .Z(\SUBBYTES[6].a/w1865 ) );
  XOR \SUBBYTES[6].a/U4503  ( .A(n13437), .B(n12957), .Z(n12955) );
  XOR \SUBBYTES[6].a/U4502  ( .A(\w1[6][60] ), .B(\SUBBYTES[6].a/w1929 ), .Z(
        n12956) );
  XOR \SUBBYTES[6].a/U4501  ( .A(\SUBBYTES[6].a/w1842 ), .B(
        \SUBBYTES[6].a/w1847 ), .Z(n12957) );
  XOR \SUBBYTES[6].a/U4500  ( .A(n12959), .B(n12958), .Z(n13435) );
  XOR \SUBBYTES[6].a/U4499  ( .A(\SUBBYTES[6].a/w1875 ), .B(\w1[6][63] ), .Z(
        n12958) );
  XOR \SUBBYTES[6].a/U4498  ( .A(\SUBBYTES[6].a/w1850 ), .B(
        \SUBBYTES[6].a/w1857 ), .Z(n12959) );
  XOR \SUBBYTES[6].a/U4497  ( .A(n13434), .B(n13435), .Z(\SUBBYTES[6].a/w1877 ) );
  XOR \SUBBYTES[6].a/U4496  ( .A(\w1[6][59] ), .B(n12960), .Z(n13438) );
  XOR \SUBBYTES[6].a/U4495  ( .A(\SUBBYTES[6].a/w1839 ), .B(
        \SUBBYTES[6].a/w1842 ), .Z(n12960) );
  XOR \SUBBYTES[6].a/U4494  ( .A(n12962), .B(n12961), .Z(\SUBBYTES[6].a/w1866 ) );
  XOR \SUBBYTES[6].a/U4493  ( .A(n13438), .B(n12963), .Z(n12961) );
  XOR \SUBBYTES[6].a/U4492  ( .A(\w1[6][62] ), .B(\SUBBYTES[6].a/w1908 ), .Z(
        n12962) );
  XOR \SUBBYTES[6].a/U4491  ( .A(\SUBBYTES[6].a/w1847 ), .B(
        \SUBBYTES[6].a/w1848 ), .Z(n12963) );
  XOR \SUBBYTES[6].a/U4490  ( .A(n13436), .B(n13435), .Z(\SUBBYTES[6].a/w1886 ) );
  XOR \SUBBYTES[6].a/U4489  ( .A(n12965), .B(n12964), .Z(\SUBBYTES[6].a/w1887 ) );
  XOR \SUBBYTES[6].a/U4488  ( .A(\w1[6][63] ), .B(n13437), .Z(n12964) );
  XOR \SUBBYTES[6].a/U4487  ( .A(\SUBBYTES[6].a/w1839 ), .B(
        \SUBBYTES[6].a/w1848 ), .Z(n12965) );
  XOR \SUBBYTES[6].a/U4486  ( .A(n12967), .B(n12966), .Z(\SUBBYTES[6].a/w1863 ) );
  XOR \SUBBYTES[6].a/U4485  ( .A(n12969), .B(n12968), .Z(n12966) );
  XOR \SUBBYTES[6].a/U4484  ( .A(\w1[6][63] ), .B(\SUBBYTES[6].a/w1947 ), .Z(
        n12967) );
  XOR \SUBBYTES[6].a/U4483  ( .A(\SUBBYTES[6].a/w1854 ), .B(
        \SUBBYTES[6].a/w1857 ), .Z(n12968) );
  XOR \SUBBYTES[6].a/U4482  ( .A(\SUBBYTES[6].a/w1840 ), .B(
        \SUBBYTES[6].a/w1842 ), .Z(n12969) );
  XOR \SUBBYTES[6].a/U4481  ( .A(n12971), .B(n12970), .Z(\SUBBYTES[6].a/w1864 ) );
  XOR \SUBBYTES[6].a/U4480  ( .A(n13438), .B(n12972), .Z(n12970) );
  XOR \SUBBYTES[6].a/U4479  ( .A(\w1[6][61] ), .B(n13439), .Z(n12971) );
  XOR \SUBBYTES[6].a/U4478  ( .A(\SUBBYTES[6].a/w1854 ), .B(
        \SUBBYTES[6].a/w1855 ), .Z(n12972) );
  XOR \SUBBYTES[6].a/U4477  ( .A(n12974), .B(n12973), .Z(\SUBBYTES[6].a/w1880 ) );
  XOR \SUBBYTES[6].a/U4476  ( .A(\w1[6][57] ), .B(n12975), .Z(n12973) );
  XOR \SUBBYTES[6].a/U4475  ( .A(\SUBBYTES[6].a/w1855 ), .B(
        \SUBBYTES[6].a/w1857 ), .Z(n12974) );
  XOR \SUBBYTES[6].a/U4474  ( .A(\SUBBYTES[6].a/w1839 ), .B(
        \SUBBYTES[6].a/w1840 ), .Z(n12975) );
  XOR \SUBBYTES[6].a/U4473  ( .A(\w1[6][65] ), .B(n12976), .Z(n13440) );
  XOR \SUBBYTES[6].a/U4472  ( .A(\w1[6][67] ), .B(\w1[6][66] ), .Z(n12976) );
  XOR \SUBBYTES[6].a/U4471  ( .A(\w1[6][70] ), .B(n13440), .Z(
        \SUBBYTES[6].a/w1722 ) );
  XOR \SUBBYTES[6].a/U4470  ( .A(\w1[6][64] ), .B(\SUBBYTES[6].a/w1722 ), .Z(
        \SUBBYTES[6].a/w1609 ) );
  XOR \SUBBYTES[6].a/U4469  ( .A(\w1[6][64] ), .B(n12977), .Z(
        \SUBBYTES[6].a/w1610 ) );
  XOR \SUBBYTES[6].a/U4468  ( .A(\w1[6][70] ), .B(\w1[6][69] ), .Z(n12977) );
  XOR \SUBBYTES[6].a/U4467  ( .A(\w1[6][69] ), .B(n13440), .Z(
        \SUBBYTES[6].a/w1740 ) );
  XOR \SUBBYTES[6].a/U4466  ( .A(n12979), .B(n12978), .Z(\SUBBYTES[6].a/w1733 ) );
  XOR \SUBBYTES[6].a/U4465  ( .A(\w1[6][67] ), .B(\w1[6][65] ), .Z(n12978) );
  XOR \SUBBYTES[6].a/U4464  ( .A(\w1[6][71] ), .B(\w1[6][68] ), .Z(n12979) );
  XOR \SUBBYTES[6].a/U4463  ( .A(\w1[6][64] ), .B(\SUBBYTES[6].a/w1733 ), .Z(
        \SUBBYTES[6].a/w1612 ) );
  XOR \SUBBYTES[6].a/U4462  ( .A(n12981), .B(n12980), .Z(\SUBBYTES[6].a/w1720 ) );
  XOR \SUBBYTES[6].a/U4461  ( .A(\SUBBYTES[6].a/w1681 ), .B(n1044), .Z(n12980)
         );
  XOR \SUBBYTES[6].a/U4460  ( .A(\SUBBYTES[6].a/w1674 ), .B(
        \SUBBYTES[6].a/w1677 ), .Z(n12981) );
  XOR \SUBBYTES[6].a/U4459  ( .A(n12983), .B(n12982), .Z(\SUBBYTES[6].a/w1721 ) );
  XOR \SUBBYTES[6].a/U4458  ( .A(\SUBBYTES[6].a/w1681 ), .B(n12247), .Z(n12982) );
  XOR \SUBBYTES[6].a/U4457  ( .A(\SUBBYTES[6].a/w1674 ), .B(n12246), .Z(n12983) );
  XOR \SUBBYTES[6].a/U4456  ( .A(\SUBBYTES[6].a/w1733 ), .B(n12984), .Z(
        \SUBBYTES[6].a/w1723 ) );
  XOR \SUBBYTES[6].a/U4455  ( .A(\w1[6][70] ), .B(\w1[6][69] ), .Z(n12984) );
  XOR \SUBBYTES[6].a/U4454  ( .A(n12986), .B(n12985), .Z(\SUBBYTES[6].a/w1724 ) );
  XOR \SUBBYTES[6].a/U4453  ( .A(n12247), .B(n1044), .Z(n12985) );
  XOR \SUBBYTES[6].a/U4452  ( .A(n12246), .B(\SUBBYTES[6].a/w1677 ), .Z(n12986) );
  XOR \SUBBYTES[6].a/U4451  ( .A(\w1[6][71] ), .B(\w1[6][66] ), .Z(n13446) );
  XOR \SUBBYTES[6].a/U4450  ( .A(n13446), .B(n12987), .Z(\SUBBYTES[6].a/w1725 ) );
  XOR \SUBBYTES[6].a/U4449  ( .A(\w1[6][69] ), .B(\w1[6][68] ), .Z(n12987) );
  XOR \SUBBYTES[6].a/U4448  ( .A(\w1[6][71] ), .B(\SUBBYTES[6].a/w1610 ), .Z(
        \SUBBYTES[6].a/w1613 ) );
  XOR \SUBBYTES[6].a/U4447  ( .A(\w1[6][65] ), .B(\SUBBYTES[6].a/w1610 ), .Z(
        \SUBBYTES[6].a/w1614 ) );
  XOR \SUBBYTES[6].a/U4446  ( .A(\w1[6][68] ), .B(\SUBBYTES[6].a/w1610 ), .Z(
        \SUBBYTES[6].a/w1615 ) );
  XOR \SUBBYTES[6].a/U4445  ( .A(\SUBBYTES[6].a/w1614 ), .B(n13446), .Z(
        \SUBBYTES[6].a/w1616 ) );
  XOR \SUBBYTES[6].a/U4444  ( .A(n13446), .B(n12988), .Z(\SUBBYTES[6].a/w1701 ) );
  XOR \SUBBYTES[6].a/U4443  ( .A(\w1[6][68] ), .B(\w1[6][65] ), .Z(n12988) );
  XOR \SUBBYTES[6].a/U4442  ( .A(n12990), .B(n12989), .Z(n13443) );
  XOR \SUBBYTES[6].a/U4441  ( .A(\w1[6][68] ), .B(n12991), .Z(n12989) );
  XOR \SUBBYTES[6].a/U4440  ( .A(\SUBBYTES[6].a/w1666 ), .B(\w1[6][70] ), .Z(
        n12990) );
  XOR \SUBBYTES[6].a/U4439  ( .A(\SUBBYTES[6].a/w1640 ), .B(
        \SUBBYTES[6].a/w1647 ), .Z(n12991) );
  XOR \SUBBYTES[6].a/U4438  ( .A(n12993), .B(n12992), .Z(n13441) );
  XOR \SUBBYTES[6].a/U4437  ( .A(\w1[6][65] ), .B(n12994), .Z(n12992) );
  XOR \SUBBYTES[6].a/U4436  ( .A(\SUBBYTES[6].a/w1665 ), .B(\w1[6][69] ), .Z(
        n12993) );
  XOR \SUBBYTES[6].a/U4435  ( .A(\SUBBYTES[6].a/w1641 ), .B(
        \SUBBYTES[6].a/w1648 ), .Z(n12994) );
  XOR \SUBBYTES[6].a/U4434  ( .A(n13443), .B(n13441), .Z(\SUBBYTES[6].a/w1671 ) );
  XOR \SUBBYTES[6].a/U4433  ( .A(\w1[6][69] ), .B(n12995), .Z(n13444) );
  XOR \SUBBYTES[6].a/U4432  ( .A(\SUBBYTES[6].a/w1633 ), .B(
        \SUBBYTES[6].a/w1643 ), .Z(n12995) );
  XOR \SUBBYTES[6].a/U4431  ( .A(n12997), .B(n12996), .Z(\SUBBYTES[6].a/w1658 ) );
  XOR \SUBBYTES[6].a/U4430  ( .A(n13444), .B(n12998), .Z(n12996) );
  XOR \SUBBYTES[6].a/U4429  ( .A(\w1[6][68] ), .B(\SUBBYTES[6].a/w1722 ), .Z(
        n12997) );
  XOR \SUBBYTES[6].a/U4428  ( .A(\SUBBYTES[6].a/w1635 ), .B(
        \SUBBYTES[6].a/w1640 ), .Z(n12998) );
  XOR \SUBBYTES[6].a/U4427  ( .A(n13000), .B(n12999), .Z(n13442) );
  XOR \SUBBYTES[6].a/U4426  ( .A(\SUBBYTES[6].a/w1668 ), .B(\w1[6][71] ), .Z(
        n12999) );
  XOR \SUBBYTES[6].a/U4425  ( .A(\SUBBYTES[6].a/w1643 ), .B(
        \SUBBYTES[6].a/w1650 ), .Z(n13000) );
  XOR \SUBBYTES[6].a/U4424  ( .A(n13441), .B(n13442), .Z(\SUBBYTES[6].a/w1670 ) );
  XOR \SUBBYTES[6].a/U4423  ( .A(\w1[6][67] ), .B(n13001), .Z(n13445) );
  XOR \SUBBYTES[6].a/U4422  ( .A(\SUBBYTES[6].a/w1632 ), .B(
        \SUBBYTES[6].a/w1635 ), .Z(n13001) );
  XOR \SUBBYTES[6].a/U4421  ( .A(n13003), .B(n13002), .Z(\SUBBYTES[6].a/w1659 ) );
  XOR \SUBBYTES[6].a/U4420  ( .A(n13445), .B(n13004), .Z(n13002) );
  XOR \SUBBYTES[6].a/U4419  ( .A(\w1[6][70] ), .B(\SUBBYTES[6].a/w1701 ), .Z(
        n13003) );
  XOR \SUBBYTES[6].a/U4418  ( .A(\SUBBYTES[6].a/w1640 ), .B(
        \SUBBYTES[6].a/w1641 ), .Z(n13004) );
  XOR \SUBBYTES[6].a/U4417  ( .A(n13443), .B(n13442), .Z(\SUBBYTES[6].a/w1679 ) );
  XOR \SUBBYTES[6].a/U4416  ( .A(n13006), .B(n13005), .Z(\SUBBYTES[6].a/w1680 ) );
  XOR \SUBBYTES[6].a/U4415  ( .A(\w1[6][71] ), .B(n13444), .Z(n13005) );
  XOR \SUBBYTES[6].a/U4414  ( .A(\SUBBYTES[6].a/w1632 ), .B(
        \SUBBYTES[6].a/w1641 ), .Z(n13006) );
  XOR \SUBBYTES[6].a/U4413  ( .A(n13008), .B(n13007), .Z(\SUBBYTES[6].a/w1656 ) );
  XOR \SUBBYTES[6].a/U4412  ( .A(n13010), .B(n13009), .Z(n13007) );
  XOR \SUBBYTES[6].a/U4411  ( .A(\w1[6][71] ), .B(\SUBBYTES[6].a/w1740 ), .Z(
        n13008) );
  XOR \SUBBYTES[6].a/U4410  ( .A(\SUBBYTES[6].a/w1647 ), .B(
        \SUBBYTES[6].a/w1650 ), .Z(n13009) );
  XOR \SUBBYTES[6].a/U4409  ( .A(\SUBBYTES[6].a/w1633 ), .B(
        \SUBBYTES[6].a/w1635 ), .Z(n13010) );
  XOR \SUBBYTES[6].a/U4408  ( .A(n13012), .B(n13011), .Z(\SUBBYTES[6].a/w1657 ) );
  XOR \SUBBYTES[6].a/U4407  ( .A(n13445), .B(n13013), .Z(n13011) );
  XOR \SUBBYTES[6].a/U4406  ( .A(\w1[6][69] ), .B(n13446), .Z(n13012) );
  XOR \SUBBYTES[6].a/U4405  ( .A(\SUBBYTES[6].a/w1647 ), .B(
        \SUBBYTES[6].a/w1648 ), .Z(n13013) );
  XOR \SUBBYTES[6].a/U4404  ( .A(n13015), .B(n13014), .Z(\SUBBYTES[6].a/w1673 ) );
  XOR \SUBBYTES[6].a/U4403  ( .A(\w1[6][65] ), .B(n13016), .Z(n13014) );
  XOR \SUBBYTES[6].a/U4402  ( .A(\SUBBYTES[6].a/w1648 ), .B(
        \SUBBYTES[6].a/w1650 ), .Z(n13015) );
  XOR \SUBBYTES[6].a/U4401  ( .A(\SUBBYTES[6].a/w1632 ), .B(
        \SUBBYTES[6].a/w1633 ), .Z(n13016) );
  XOR \SUBBYTES[6].a/U4400  ( .A(\w1[6][73] ), .B(n13017), .Z(n13447) );
  XOR \SUBBYTES[6].a/U4399  ( .A(\w1[6][75] ), .B(\w1[6][74] ), .Z(n13017) );
  XOR \SUBBYTES[6].a/U4398  ( .A(\w1[6][78] ), .B(n13447), .Z(
        \SUBBYTES[6].a/w1515 ) );
  XOR \SUBBYTES[6].a/U4397  ( .A(\w1[6][72] ), .B(\SUBBYTES[6].a/w1515 ), .Z(
        \SUBBYTES[6].a/w1402 ) );
  XOR \SUBBYTES[6].a/U4396  ( .A(\w1[6][72] ), .B(n13018), .Z(
        \SUBBYTES[6].a/w1403 ) );
  XOR \SUBBYTES[6].a/U4395  ( .A(\w1[6][78] ), .B(\w1[6][77] ), .Z(n13018) );
  XOR \SUBBYTES[6].a/U4394  ( .A(\w1[6][77] ), .B(n13447), .Z(
        \SUBBYTES[6].a/w1533 ) );
  XOR \SUBBYTES[6].a/U4393  ( .A(n13020), .B(n13019), .Z(\SUBBYTES[6].a/w1526 ) );
  XOR \SUBBYTES[6].a/U4392  ( .A(\w1[6][75] ), .B(\w1[6][73] ), .Z(n13019) );
  XOR \SUBBYTES[6].a/U4391  ( .A(\w1[6][79] ), .B(\w1[6][76] ), .Z(n13020) );
  XOR \SUBBYTES[6].a/U4390  ( .A(\w1[6][72] ), .B(\SUBBYTES[6].a/w1526 ), .Z(
        \SUBBYTES[6].a/w1405 ) );
  XOR \SUBBYTES[6].a/U4389  ( .A(n13022), .B(n13021), .Z(\SUBBYTES[6].a/w1513 ) );
  XOR \SUBBYTES[6].a/U4388  ( .A(\SUBBYTES[6].a/w1474 ), .B(n1043), .Z(n13021)
         );
  XOR \SUBBYTES[6].a/U4387  ( .A(\SUBBYTES[6].a/w1467 ), .B(
        \SUBBYTES[6].a/w1470 ), .Z(n13022) );
  XOR \SUBBYTES[6].a/U4386  ( .A(n13024), .B(n13023), .Z(\SUBBYTES[6].a/w1514 ) );
  XOR \SUBBYTES[6].a/U4385  ( .A(\SUBBYTES[6].a/w1474 ), .B(n12245), .Z(n13023) );
  XOR \SUBBYTES[6].a/U4384  ( .A(\SUBBYTES[6].a/w1467 ), .B(n12244), .Z(n13024) );
  XOR \SUBBYTES[6].a/U4383  ( .A(\SUBBYTES[6].a/w1526 ), .B(n13025), .Z(
        \SUBBYTES[6].a/w1516 ) );
  XOR \SUBBYTES[6].a/U4382  ( .A(\w1[6][78] ), .B(\w1[6][77] ), .Z(n13025) );
  XOR \SUBBYTES[6].a/U4381  ( .A(n13027), .B(n13026), .Z(\SUBBYTES[6].a/w1517 ) );
  XOR \SUBBYTES[6].a/U4380  ( .A(n12245), .B(n1043), .Z(n13026) );
  XOR \SUBBYTES[6].a/U4379  ( .A(n12244), .B(\SUBBYTES[6].a/w1470 ), .Z(n13027) );
  XOR \SUBBYTES[6].a/U4378  ( .A(\w1[6][79] ), .B(\w1[6][74] ), .Z(n13453) );
  XOR \SUBBYTES[6].a/U4377  ( .A(n13453), .B(n13028), .Z(\SUBBYTES[6].a/w1518 ) );
  XOR \SUBBYTES[6].a/U4376  ( .A(\w1[6][77] ), .B(\w1[6][76] ), .Z(n13028) );
  XOR \SUBBYTES[6].a/U4375  ( .A(\w1[6][79] ), .B(\SUBBYTES[6].a/w1403 ), .Z(
        \SUBBYTES[6].a/w1406 ) );
  XOR \SUBBYTES[6].a/U4374  ( .A(\w1[6][73] ), .B(\SUBBYTES[6].a/w1403 ), .Z(
        \SUBBYTES[6].a/w1407 ) );
  XOR \SUBBYTES[6].a/U4373  ( .A(\w1[6][76] ), .B(\SUBBYTES[6].a/w1403 ), .Z(
        \SUBBYTES[6].a/w1408 ) );
  XOR \SUBBYTES[6].a/U4372  ( .A(\SUBBYTES[6].a/w1407 ), .B(n13453), .Z(
        \SUBBYTES[6].a/w1409 ) );
  XOR \SUBBYTES[6].a/U4371  ( .A(n13453), .B(n13029), .Z(\SUBBYTES[6].a/w1494 ) );
  XOR \SUBBYTES[6].a/U4370  ( .A(\w1[6][76] ), .B(\w1[6][73] ), .Z(n13029) );
  XOR \SUBBYTES[6].a/U4369  ( .A(n13031), .B(n13030), .Z(n13450) );
  XOR \SUBBYTES[6].a/U4368  ( .A(\w1[6][76] ), .B(n13032), .Z(n13030) );
  XOR \SUBBYTES[6].a/U4367  ( .A(\SUBBYTES[6].a/w1459 ), .B(\w1[6][78] ), .Z(
        n13031) );
  XOR \SUBBYTES[6].a/U4366  ( .A(\SUBBYTES[6].a/w1433 ), .B(
        \SUBBYTES[6].a/w1440 ), .Z(n13032) );
  XOR \SUBBYTES[6].a/U4365  ( .A(n13034), .B(n13033), .Z(n13448) );
  XOR \SUBBYTES[6].a/U4364  ( .A(\w1[6][73] ), .B(n13035), .Z(n13033) );
  XOR \SUBBYTES[6].a/U4363  ( .A(\SUBBYTES[6].a/w1458 ), .B(\w1[6][77] ), .Z(
        n13034) );
  XOR \SUBBYTES[6].a/U4362  ( .A(\SUBBYTES[6].a/w1434 ), .B(
        \SUBBYTES[6].a/w1441 ), .Z(n13035) );
  XOR \SUBBYTES[6].a/U4361  ( .A(n13450), .B(n13448), .Z(\SUBBYTES[6].a/w1464 ) );
  XOR \SUBBYTES[6].a/U4360  ( .A(\w1[6][77] ), .B(n13036), .Z(n13451) );
  XOR \SUBBYTES[6].a/U4359  ( .A(\SUBBYTES[6].a/w1426 ), .B(
        \SUBBYTES[6].a/w1436 ), .Z(n13036) );
  XOR \SUBBYTES[6].a/U4358  ( .A(n13038), .B(n13037), .Z(\SUBBYTES[6].a/w1451 ) );
  XOR \SUBBYTES[6].a/U4357  ( .A(n13451), .B(n13039), .Z(n13037) );
  XOR \SUBBYTES[6].a/U4356  ( .A(\w1[6][76] ), .B(\SUBBYTES[6].a/w1515 ), .Z(
        n13038) );
  XOR \SUBBYTES[6].a/U4355  ( .A(\SUBBYTES[6].a/w1428 ), .B(
        \SUBBYTES[6].a/w1433 ), .Z(n13039) );
  XOR \SUBBYTES[6].a/U4354  ( .A(n13041), .B(n13040), .Z(n13449) );
  XOR \SUBBYTES[6].a/U4353  ( .A(\SUBBYTES[6].a/w1461 ), .B(\w1[6][79] ), .Z(
        n13040) );
  XOR \SUBBYTES[6].a/U4352  ( .A(\SUBBYTES[6].a/w1436 ), .B(
        \SUBBYTES[6].a/w1443 ), .Z(n13041) );
  XOR \SUBBYTES[6].a/U4351  ( .A(n13448), .B(n13449), .Z(\SUBBYTES[6].a/w1463 ) );
  XOR \SUBBYTES[6].a/U4350  ( .A(\w1[6][75] ), .B(n13042), .Z(n13452) );
  XOR \SUBBYTES[6].a/U4349  ( .A(\SUBBYTES[6].a/w1425 ), .B(
        \SUBBYTES[6].a/w1428 ), .Z(n13042) );
  XOR \SUBBYTES[6].a/U4348  ( .A(n13044), .B(n13043), .Z(\SUBBYTES[6].a/w1452 ) );
  XOR \SUBBYTES[6].a/U4347  ( .A(n13452), .B(n13045), .Z(n13043) );
  XOR \SUBBYTES[6].a/U4346  ( .A(\w1[6][78] ), .B(\SUBBYTES[6].a/w1494 ), .Z(
        n13044) );
  XOR \SUBBYTES[6].a/U4345  ( .A(\SUBBYTES[6].a/w1433 ), .B(
        \SUBBYTES[6].a/w1434 ), .Z(n13045) );
  XOR \SUBBYTES[6].a/U4344  ( .A(n13450), .B(n13449), .Z(\SUBBYTES[6].a/w1472 ) );
  XOR \SUBBYTES[6].a/U4343  ( .A(n13047), .B(n13046), .Z(\SUBBYTES[6].a/w1473 ) );
  XOR \SUBBYTES[6].a/U4342  ( .A(\w1[6][79] ), .B(n13451), .Z(n13046) );
  XOR \SUBBYTES[6].a/U4341  ( .A(\SUBBYTES[6].a/w1425 ), .B(
        \SUBBYTES[6].a/w1434 ), .Z(n13047) );
  XOR \SUBBYTES[6].a/U4340  ( .A(n13049), .B(n13048), .Z(\SUBBYTES[6].a/w1449 ) );
  XOR \SUBBYTES[6].a/U4339  ( .A(n13051), .B(n13050), .Z(n13048) );
  XOR \SUBBYTES[6].a/U4338  ( .A(\w1[6][79] ), .B(\SUBBYTES[6].a/w1533 ), .Z(
        n13049) );
  XOR \SUBBYTES[6].a/U4337  ( .A(\SUBBYTES[6].a/w1440 ), .B(
        \SUBBYTES[6].a/w1443 ), .Z(n13050) );
  XOR \SUBBYTES[6].a/U4336  ( .A(\SUBBYTES[6].a/w1426 ), .B(
        \SUBBYTES[6].a/w1428 ), .Z(n13051) );
  XOR \SUBBYTES[6].a/U4335  ( .A(n13053), .B(n13052), .Z(\SUBBYTES[6].a/w1450 ) );
  XOR \SUBBYTES[6].a/U4334  ( .A(n13452), .B(n13054), .Z(n13052) );
  XOR \SUBBYTES[6].a/U4333  ( .A(\w1[6][77] ), .B(n13453), .Z(n13053) );
  XOR \SUBBYTES[6].a/U4332  ( .A(\SUBBYTES[6].a/w1440 ), .B(
        \SUBBYTES[6].a/w1441 ), .Z(n13054) );
  XOR \SUBBYTES[6].a/U4331  ( .A(n13056), .B(n13055), .Z(\SUBBYTES[6].a/w1466 ) );
  XOR \SUBBYTES[6].a/U4330  ( .A(\w1[6][73] ), .B(n13057), .Z(n13055) );
  XOR \SUBBYTES[6].a/U4329  ( .A(\SUBBYTES[6].a/w1441 ), .B(
        \SUBBYTES[6].a/w1443 ), .Z(n13056) );
  XOR \SUBBYTES[6].a/U4328  ( .A(\SUBBYTES[6].a/w1425 ), .B(
        \SUBBYTES[6].a/w1426 ), .Z(n13057) );
  XOR \SUBBYTES[6].a/U4327  ( .A(\w1[6][81] ), .B(n13058), .Z(n13454) );
  XOR \SUBBYTES[6].a/U4326  ( .A(\w1[6][83] ), .B(\w1[6][82] ), .Z(n13058) );
  XOR \SUBBYTES[6].a/U4325  ( .A(\w1[6][86] ), .B(n13454), .Z(
        \SUBBYTES[6].a/w1308 ) );
  XOR \SUBBYTES[6].a/U4324  ( .A(\w1[6][80] ), .B(\SUBBYTES[6].a/w1308 ), .Z(
        \SUBBYTES[6].a/w1195 ) );
  XOR \SUBBYTES[6].a/U4323  ( .A(\w1[6][80] ), .B(n13059), .Z(
        \SUBBYTES[6].a/w1196 ) );
  XOR \SUBBYTES[6].a/U4322  ( .A(\w1[6][86] ), .B(\w1[6][85] ), .Z(n13059) );
  XOR \SUBBYTES[6].a/U4321  ( .A(\w1[6][85] ), .B(n13454), .Z(
        \SUBBYTES[6].a/w1326 ) );
  XOR \SUBBYTES[6].a/U4320  ( .A(n13061), .B(n13060), .Z(\SUBBYTES[6].a/w1319 ) );
  XOR \SUBBYTES[6].a/U4319  ( .A(\w1[6][83] ), .B(\w1[6][81] ), .Z(n13060) );
  XOR \SUBBYTES[6].a/U4318  ( .A(\w1[6][87] ), .B(\w1[6][84] ), .Z(n13061) );
  XOR \SUBBYTES[6].a/U4317  ( .A(\w1[6][80] ), .B(\SUBBYTES[6].a/w1319 ), .Z(
        \SUBBYTES[6].a/w1198 ) );
  XOR \SUBBYTES[6].a/U4316  ( .A(n13063), .B(n13062), .Z(\SUBBYTES[6].a/w1306 ) );
  XOR \SUBBYTES[6].a/U4315  ( .A(\SUBBYTES[6].a/w1267 ), .B(n1042), .Z(n13062)
         );
  XOR \SUBBYTES[6].a/U4314  ( .A(\SUBBYTES[6].a/w1260 ), .B(
        \SUBBYTES[6].a/w1263 ), .Z(n13063) );
  XOR \SUBBYTES[6].a/U4313  ( .A(n13065), .B(n13064), .Z(\SUBBYTES[6].a/w1307 ) );
  XOR \SUBBYTES[6].a/U4312  ( .A(\SUBBYTES[6].a/w1267 ), .B(n12243), .Z(n13064) );
  XOR \SUBBYTES[6].a/U4311  ( .A(\SUBBYTES[6].a/w1260 ), .B(n12242), .Z(n13065) );
  XOR \SUBBYTES[6].a/U4310  ( .A(\SUBBYTES[6].a/w1319 ), .B(n13066), .Z(
        \SUBBYTES[6].a/w1309 ) );
  XOR \SUBBYTES[6].a/U4309  ( .A(\w1[6][86] ), .B(\w1[6][85] ), .Z(n13066) );
  XOR \SUBBYTES[6].a/U4308  ( .A(n13068), .B(n13067), .Z(\SUBBYTES[6].a/w1310 ) );
  XOR \SUBBYTES[6].a/U4307  ( .A(n12243), .B(n1042), .Z(n13067) );
  XOR \SUBBYTES[6].a/U4306  ( .A(n12242), .B(\SUBBYTES[6].a/w1263 ), .Z(n13068) );
  XOR \SUBBYTES[6].a/U4305  ( .A(\w1[6][87] ), .B(\w1[6][82] ), .Z(n13460) );
  XOR \SUBBYTES[6].a/U4304  ( .A(n13460), .B(n13069), .Z(\SUBBYTES[6].a/w1311 ) );
  XOR \SUBBYTES[6].a/U4303  ( .A(\w1[6][85] ), .B(\w1[6][84] ), .Z(n13069) );
  XOR \SUBBYTES[6].a/U4302  ( .A(\w1[6][87] ), .B(\SUBBYTES[6].a/w1196 ), .Z(
        \SUBBYTES[6].a/w1199 ) );
  XOR \SUBBYTES[6].a/U4301  ( .A(\w1[6][81] ), .B(\SUBBYTES[6].a/w1196 ), .Z(
        \SUBBYTES[6].a/w1200 ) );
  XOR \SUBBYTES[6].a/U4300  ( .A(\w1[6][84] ), .B(\SUBBYTES[6].a/w1196 ), .Z(
        \SUBBYTES[6].a/w1201 ) );
  XOR \SUBBYTES[6].a/U4299  ( .A(\SUBBYTES[6].a/w1200 ), .B(n13460), .Z(
        \SUBBYTES[6].a/w1202 ) );
  XOR \SUBBYTES[6].a/U4298  ( .A(n13460), .B(n13070), .Z(\SUBBYTES[6].a/w1287 ) );
  XOR \SUBBYTES[6].a/U4297  ( .A(\w1[6][84] ), .B(\w1[6][81] ), .Z(n13070) );
  XOR \SUBBYTES[6].a/U4296  ( .A(n13072), .B(n13071), .Z(n13457) );
  XOR \SUBBYTES[6].a/U4295  ( .A(\w1[6][84] ), .B(n13073), .Z(n13071) );
  XOR \SUBBYTES[6].a/U4294  ( .A(\SUBBYTES[6].a/w1252 ), .B(\w1[6][86] ), .Z(
        n13072) );
  XOR \SUBBYTES[6].a/U4293  ( .A(\SUBBYTES[6].a/w1226 ), .B(
        \SUBBYTES[6].a/w1233 ), .Z(n13073) );
  XOR \SUBBYTES[6].a/U4292  ( .A(n13075), .B(n13074), .Z(n13455) );
  XOR \SUBBYTES[6].a/U4291  ( .A(\w1[6][81] ), .B(n13076), .Z(n13074) );
  XOR \SUBBYTES[6].a/U4290  ( .A(\SUBBYTES[6].a/w1251 ), .B(\w1[6][85] ), .Z(
        n13075) );
  XOR \SUBBYTES[6].a/U4289  ( .A(\SUBBYTES[6].a/w1227 ), .B(
        \SUBBYTES[6].a/w1234 ), .Z(n13076) );
  XOR \SUBBYTES[6].a/U4288  ( .A(n13457), .B(n13455), .Z(\SUBBYTES[6].a/w1257 ) );
  XOR \SUBBYTES[6].a/U4287  ( .A(\w1[6][85] ), .B(n13077), .Z(n13458) );
  XOR \SUBBYTES[6].a/U4286  ( .A(\SUBBYTES[6].a/w1219 ), .B(
        \SUBBYTES[6].a/w1229 ), .Z(n13077) );
  XOR \SUBBYTES[6].a/U4285  ( .A(n13079), .B(n13078), .Z(\SUBBYTES[6].a/w1244 ) );
  XOR \SUBBYTES[6].a/U4284  ( .A(n13458), .B(n13080), .Z(n13078) );
  XOR \SUBBYTES[6].a/U4283  ( .A(\w1[6][84] ), .B(\SUBBYTES[6].a/w1308 ), .Z(
        n13079) );
  XOR \SUBBYTES[6].a/U4282  ( .A(\SUBBYTES[6].a/w1221 ), .B(
        \SUBBYTES[6].a/w1226 ), .Z(n13080) );
  XOR \SUBBYTES[6].a/U4281  ( .A(n13082), .B(n13081), .Z(n13456) );
  XOR \SUBBYTES[6].a/U4280  ( .A(\SUBBYTES[6].a/w1254 ), .B(\w1[6][87] ), .Z(
        n13081) );
  XOR \SUBBYTES[6].a/U4279  ( .A(\SUBBYTES[6].a/w1229 ), .B(
        \SUBBYTES[6].a/w1236 ), .Z(n13082) );
  XOR \SUBBYTES[6].a/U4278  ( .A(n13455), .B(n13456), .Z(\SUBBYTES[6].a/w1256 ) );
  XOR \SUBBYTES[6].a/U4277  ( .A(\w1[6][83] ), .B(n13083), .Z(n13459) );
  XOR \SUBBYTES[6].a/U4276  ( .A(\SUBBYTES[6].a/w1218 ), .B(
        \SUBBYTES[6].a/w1221 ), .Z(n13083) );
  XOR \SUBBYTES[6].a/U4275  ( .A(n13085), .B(n13084), .Z(\SUBBYTES[6].a/w1245 ) );
  XOR \SUBBYTES[6].a/U4274  ( .A(n13459), .B(n13086), .Z(n13084) );
  XOR \SUBBYTES[6].a/U4273  ( .A(\w1[6][86] ), .B(\SUBBYTES[6].a/w1287 ), .Z(
        n13085) );
  XOR \SUBBYTES[6].a/U4272  ( .A(\SUBBYTES[6].a/w1226 ), .B(
        \SUBBYTES[6].a/w1227 ), .Z(n13086) );
  XOR \SUBBYTES[6].a/U4271  ( .A(n13457), .B(n13456), .Z(\SUBBYTES[6].a/w1265 ) );
  XOR \SUBBYTES[6].a/U4270  ( .A(n13088), .B(n13087), .Z(\SUBBYTES[6].a/w1266 ) );
  XOR \SUBBYTES[6].a/U4269  ( .A(\w1[6][87] ), .B(n13458), .Z(n13087) );
  XOR \SUBBYTES[6].a/U4268  ( .A(\SUBBYTES[6].a/w1218 ), .B(
        \SUBBYTES[6].a/w1227 ), .Z(n13088) );
  XOR \SUBBYTES[6].a/U4267  ( .A(n13090), .B(n13089), .Z(\SUBBYTES[6].a/w1242 ) );
  XOR \SUBBYTES[6].a/U4266  ( .A(n13092), .B(n13091), .Z(n13089) );
  XOR \SUBBYTES[6].a/U4265  ( .A(\w1[6][87] ), .B(\SUBBYTES[6].a/w1326 ), .Z(
        n13090) );
  XOR \SUBBYTES[6].a/U4264  ( .A(\SUBBYTES[6].a/w1233 ), .B(
        \SUBBYTES[6].a/w1236 ), .Z(n13091) );
  XOR \SUBBYTES[6].a/U4263  ( .A(\SUBBYTES[6].a/w1219 ), .B(
        \SUBBYTES[6].a/w1221 ), .Z(n13092) );
  XOR \SUBBYTES[6].a/U4262  ( .A(n13094), .B(n13093), .Z(\SUBBYTES[6].a/w1243 ) );
  XOR \SUBBYTES[6].a/U4261  ( .A(n13459), .B(n13095), .Z(n13093) );
  XOR \SUBBYTES[6].a/U4260  ( .A(\w1[6][85] ), .B(n13460), .Z(n13094) );
  XOR \SUBBYTES[6].a/U4259  ( .A(\SUBBYTES[6].a/w1233 ), .B(
        \SUBBYTES[6].a/w1234 ), .Z(n13095) );
  XOR \SUBBYTES[6].a/U4258  ( .A(n13097), .B(n13096), .Z(\SUBBYTES[6].a/w1259 ) );
  XOR \SUBBYTES[6].a/U4257  ( .A(\w1[6][81] ), .B(n13098), .Z(n13096) );
  XOR \SUBBYTES[6].a/U4256  ( .A(\SUBBYTES[6].a/w1234 ), .B(
        \SUBBYTES[6].a/w1236 ), .Z(n13097) );
  XOR \SUBBYTES[6].a/U4255  ( .A(\SUBBYTES[6].a/w1218 ), .B(
        \SUBBYTES[6].a/w1219 ), .Z(n13098) );
  XOR \SUBBYTES[6].a/U4254  ( .A(\w1[6][89] ), .B(n13099), .Z(n13461) );
  XOR \SUBBYTES[6].a/U4253  ( .A(\w1[6][91] ), .B(\w1[6][90] ), .Z(n13099) );
  XOR \SUBBYTES[6].a/U4252  ( .A(\w1[6][94] ), .B(n13461), .Z(
        \SUBBYTES[6].a/w1101 ) );
  XOR \SUBBYTES[6].a/U4251  ( .A(\w1[6][88] ), .B(\SUBBYTES[6].a/w1101 ), .Z(
        \SUBBYTES[6].a/w988 ) );
  XOR \SUBBYTES[6].a/U4250  ( .A(\w1[6][88] ), .B(n13100), .Z(
        \SUBBYTES[6].a/w989 ) );
  XOR \SUBBYTES[6].a/U4249  ( .A(\w1[6][94] ), .B(\w1[6][93] ), .Z(n13100) );
  XOR \SUBBYTES[6].a/U4248  ( .A(\w1[6][93] ), .B(n13461), .Z(
        \SUBBYTES[6].a/w1119 ) );
  XOR \SUBBYTES[6].a/U4247  ( .A(n13102), .B(n13101), .Z(\SUBBYTES[6].a/w1112 ) );
  XOR \SUBBYTES[6].a/U4246  ( .A(\w1[6][91] ), .B(\w1[6][89] ), .Z(n13101) );
  XOR \SUBBYTES[6].a/U4245  ( .A(\w1[6][95] ), .B(\w1[6][92] ), .Z(n13102) );
  XOR \SUBBYTES[6].a/U4244  ( .A(\w1[6][88] ), .B(\SUBBYTES[6].a/w1112 ), .Z(
        \SUBBYTES[6].a/w991 ) );
  XOR \SUBBYTES[6].a/U4243  ( .A(n13104), .B(n13103), .Z(\SUBBYTES[6].a/w1099 ) );
  XOR \SUBBYTES[6].a/U4242  ( .A(\SUBBYTES[6].a/w1060 ), .B(n1041), .Z(n13103)
         );
  XOR \SUBBYTES[6].a/U4241  ( .A(\SUBBYTES[6].a/w1053 ), .B(
        \SUBBYTES[6].a/w1056 ), .Z(n13104) );
  XOR \SUBBYTES[6].a/U4240  ( .A(n13106), .B(n13105), .Z(\SUBBYTES[6].a/w1100 ) );
  XOR \SUBBYTES[6].a/U4239  ( .A(\SUBBYTES[6].a/w1060 ), .B(n12241), .Z(n13105) );
  XOR \SUBBYTES[6].a/U4238  ( .A(\SUBBYTES[6].a/w1053 ), .B(n12240), .Z(n13106) );
  XOR \SUBBYTES[6].a/U4237  ( .A(\SUBBYTES[6].a/w1112 ), .B(n13107), .Z(
        \SUBBYTES[6].a/w1102 ) );
  XOR \SUBBYTES[6].a/U4236  ( .A(\w1[6][94] ), .B(\w1[6][93] ), .Z(n13107) );
  XOR \SUBBYTES[6].a/U4235  ( .A(n13109), .B(n13108), .Z(\SUBBYTES[6].a/w1103 ) );
  XOR \SUBBYTES[6].a/U4234  ( .A(n12241), .B(n1041), .Z(n13108) );
  XOR \SUBBYTES[6].a/U4233  ( .A(n12240), .B(\SUBBYTES[6].a/w1056 ), .Z(n13109) );
  XOR \SUBBYTES[6].a/U4232  ( .A(\w1[6][95] ), .B(\w1[6][90] ), .Z(n13467) );
  XOR \SUBBYTES[6].a/U4231  ( .A(n13467), .B(n13110), .Z(\SUBBYTES[6].a/w1104 ) );
  XOR \SUBBYTES[6].a/U4230  ( .A(\w1[6][93] ), .B(\w1[6][92] ), .Z(n13110) );
  XOR \SUBBYTES[6].a/U4229  ( .A(\w1[6][95] ), .B(\SUBBYTES[6].a/w989 ), .Z(
        \SUBBYTES[6].a/w992 ) );
  XOR \SUBBYTES[6].a/U4228  ( .A(\w1[6][89] ), .B(\SUBBYTES[6].a/w989 ), .Z(
        \SUBBYTES[6].a/w993 ) );
  XOR \SUBBYTES[6].a/U4227  ( .A(\w1[6][92] ), .B(\SUBBYTES[6].a/w989 ), .Z(
        \SUBBYTES[6].a/w994 ) );
  XOR \SUBBYTES[6].a/U4226  ( .A(\SUBBYTES[6].a/w993 ), .B(n13467), .Z(
        \SUBBYTES[6].a/w995 ) );
  XOR \SUBBYTES[6].a/U4225  ( .A(n13467), .B(n13111), .Z(\SUBBYTES[6].a/w1080 ) );
  XOR \SUBBYTES[6].a/U4224  ( .A(\w1[6][92] ), .B(\w1[6][89] ), .Z(n13111) );
  XOR \SUBBYTES[6].a/U4223  ( .A(n13113), .B(n13112), .Z(n13464) );
  XOR \SUBBYTES[6].a/U4222  ( .A(\w1[6][92] ), .B(n13114), .Z(n13112) );
  XOR \SUBBYTES[6].a/U4221  ( .A(\SUBBYTES[6].a/w1045 ), .B(\w1[6][94] ), .Z(
        n13113) );
  XOR \SUBBYTES[6].a/U4220  ( .A(\SUBBYTES[6].a/w1019 ), .B(
        \SUBBYTES[6].a/w1026 ), .Z(n13114) );
  XOR \SUBBYTES[6].a/U4219  ( .A(n13116), .B(n13115), .Z(n13462) );
  XOR \SUBBYTES[6].a/U4218  ( .A(\w1[6][89] ), .B(n13117), .Z(n13115) );
  XOR \SUBBYTES[6].a/U4217  ( .A(\SUBBYTES[6].a/w1044 ), .B(\w1[6][93] ), .Z(
        n13116) );
  XOR \SUBBYTES[6].a/U4216  ( .A(\SUBBYTES[6].a/w1020 ), .B(
        \SUBBYTES[6].a/w1027 ), .Z(n13117) );
  XOR \SUBBYTES[6].a/U4215  ( .A(n13464), .B(n13462), .Z(\SUBBYTES[6].a/w1050 ) );
  XOR \SUBBYTES[6].a/U4214  ( .A(\w1[6][93] ), .B(n13118), .Z(n13465) );
  XOR \SUBBYTES[6].a/U4213  ( .A(\SUBBYTES[6].a/w1012 ), .B(
        \SUBBYTES[6].a/w1022 ), .Z(n13118) );
  XOR \SUBBYTES[6].a/U4212  ( .A(n13120), .B(n13119), .Z(\SUBBYTES[6].a/w1037 ) );
  XOR \SUBBYTES[6].a/U4211  ( .A(n13465), .B(n13121), .Z(n13119) );
  XOR \SUBBYTES[6].a/U4210  ( .A(\w1[6][92] ), .B(\SUBBYTES[6].a/w1101 ), .Z(
        n13120) );
  XOR \SUBBYTES[6].a/U4209  ( .A(\SUBBYTES[6].a/w1014 ), .B(
        \SUBBYTES[6].a/w1019 ), .Z(n13121) );
  XOR \SUBBYTES[6].a/U4208  ( .A(n13123), .B(n13122), .Z(n13463) );
  XOR \SUBBYTES[6].a/U4207  ( .A(\SUBBYTES[6].a/w1047 ), .B(\w1[6][95] ), .Z(
        n13122) );
  XOR \SUBBYTES[6].a/U4206  ( .A(\SUBBYTES[6].a/w1022 ), .B(
        \SUBBYTES[6].a/w1029 ), .Z(n13123) );
  XOR \SUBBYTES[6].a/U4205  ( .A(n13462), .B(n13463), .Z(\SUBBYTES[6].a/w1049 ) );
  XOR \SUBBYTES[6].a/U4204  ( .A(\w1[6][91] ), .B(n13124), .Z(n13466) );
  XOR \SUBBYTES[6].a/U4203  ( .A(\SUBBYTES[6].a/w1011 ), .B(
        \SUBBYTES[6].a/w1014 ), .Z(n13124) );
  XOR \SUBBYTES[6].a/U4202  ( .A(n13126), .B(n13125), .Z(\SUBBYTES[6].a/w1038 ) );
  XOR \SUBBYTES[6].a/U4201  ( .A(n13466), .B(n13127), .Z(n13125) );
  XOR \SUBBYTES[6].a/U4200  ( .A(\w1[6][94] ), .B(\SUBBYTES[6].a/w1080 ), .Z(
        n13126) );
  XOR \SUBBYTES[6].a/U4199  ( .A(\SUBBYTES[6].a/w1019 ), .B(
        \SUBBYTES[6].a/w1020 ), .Z(n13127) );
  XOR \SUBBYTES[6].a/U4198  ( .A(n13464), .B(n13463), .Z(\SUBBYTES[6].a/w1058 ) );
  XOR \SUBBYTES[6].a/U4197  ( .A(n13129), .B(n13128), .Z(\SUBBYTES[6].a/w1059 ) );
  XOR \SUBBYTES[6].a/U4196  ( .A(\w1[6][95] ), .B(n13465), .Z(n13128) );
  XOR \SUBBYTES[6].a/U4195  ( .A(\SUBBYTES[6].a/w1011 ), .B(
        \SUBBYTES[6].a/w1020 ), .Z(n13129) );
  XOR \SUBBYTES[6].a/U4194  ( .A(n13131), .B(n13130), .Z(\SUBBYTES[6].a/w1035 ) );
  XOR \SUBBYTES[6].a/U4193  ( .A(n13133), .B(n13132), .Z(n13130) );
  XOR \SUBBYTES[6].a/U4192  ( .A(\w1[6][95] ), .B(\SUBBYTES[6].a/w1119 ), .Z(
        n13131) );
  XOR \SUBBYTES[6].a/U4191  ( .A(\SUBBYTES[6].a/w1026 ), .B(
        \SUBBYTES[6].a/w1029 ), .Z(n13132) );
  XOR \SUBBYTES[6].a/U4190  ( .A(\SUBBYTES[6].a/w1012 ), .B(
        \SUBBYTES[6].a/w1014 ), .Z(n13133) );
  XOR \SUBBYTES[6].a/U4189  ( .A(n13135), .B(n13134), .Z(\SUBBYTES[6].a/w1036 ) );
  XOR \SUBBYTES[6].a/U4188  ( .A(n13466), .B(n13136), .Z(n13134) );
  XOR \SUBBYTES[6].a/U4187  ( .A(\w1[6][93] ), .B(n13467), .Z(n13135) );
  XOR \SUBBYTES[6].a/U4186  ( .A(\SUBBYTES[6].a/w1026 ), .B(
        \SUBBYTES[6].a/w1027 ), .Z(n13136) );
  XOR \SUBBYTES[6].a/U4185  ( .A(n13138), .B(n13137), .Z(\SUBBYTES[6].a/w1052 ) );
  XOR \SUBBYTES[6].a/U4184  ( .A(\w1[6][89] ), .B(n13139), .Z(n13137) );
  XOR \SUBBYTES[6].a/U4183  ( .A(\SUBBYTES[6].a/w1027 ), .B(
        \SUBBYTES[6].a/w1029 ), .Z(n13138) );
  XOR \SUBBYTES[6].a/U4182  ( .A(\SUBBYTES[6].a/w1011 ), .B(
        \SUBBYTES[6].a/w1012 ), .Z(n13139) );
  XOR \SUBBYTES[6].a/U4181  ( .A(\w1[6][97] ), .B(n13140), .Z(n13468) );
  XOR \SUBBYTES[6].a/U4180  ( .A(\w1[6][99] ), .B(\w1[6][98] ), .Z(n13140) );
  XOR \SUBBYTES[6].a/U4179  ( .A(\w1[6][102] ), .B(n13468), .Z(
        \SUBBYTES[6].a/w894 ) );
  XOR \SUBBYTES[6].a/U4178  ( .A(\w1[6][96] ), .B(\SUBBYTES[6].a/w894 ), .Z(
        \SUBBYTES[6].a/w781 ) );
  XOR \SUBBYTES[6].a/U4177  ( .A(\w1[6][96] ), .B(n13141), .Z(
        \SUBBYTES[6].a/w782 ) );
  XOR \SUBBYTES[6].a/U4176  ( .A(\w1[6][102] ), .B(\w1[6][101] ), .Z(n13141)
         );
  XOR \SUBBYTES[6].a/U4175  ( .A(\w1[6][101] ), .B(n13468), .Z(
        \SUBBYTES[6].a/w912 ) );
  XOR \SUBBYTES[6].a/U4174  ( .A(n13143), .B(n13142), .Z(\SUBBYTES[6].a/w905 )
         );
  XOR \SUBBYTES[6].a/U4173  ( .A(\w1[6][99] ), .B(\w1[6][97] ), .Z(n13142) );
  XOR \SUBBYTES[6].a/U4172  ( .A(\w1[6][103] ), .B(\w1[6][100] ), .Z(n13143)
         );
  XOR \SUBBYTES[6].a/U4171  ( .A(\w1[6][96] ), .B(\SUBBYTES[6].a/w905 ), .Z(
        \SUBBYTES[6].a/w784 ) );
  XOR \SUBBYTES[6].a/U4170  ( .A(n13145), .B(n13144), .Z(\SUBBYTES[6].a/w892 )
         );
  XOR \SUBBYTES[6].a/U4169  ( .A(\SUBBYTES[6].a/w853 ), .B(n1040), .Z(n13144)
         );
  XOR \SUBBYTES[6].a/U4168  ( .A(\SUBBYTES[6].a/w846 ), .B(
        \SUBBYTES[6].a/w849 ), .Z(n13145) );
  XOR \SUBBYTES[6].a/U4167  ( .A(n13147), .B(n13146), .Z(\SUBBYTES[6].a/w893 )
         );
  XOR \SUBBYTES[6].a/U4166  ( .A(\SUBBYTES[6].a/w853 ), .B(n12239), .Z(n13146)
         );
  XOR \SUBBYTES[6].a/U4165  ( .A(\SUBBYTES[6].a/w846 ), .B(n12238), .Z(n13147)
         );
  XOR \SUBBYTES[6].a/U4164  ( .A(\SUBBYTES[6].a/w905 ), .B(n13148), .Z(
        \SUBBYTES[6].a/w895 ) );
  XOR \SUBBYTES[6].a/U4163  ( .A(\w1[6][102] ), .B(\w1[6][101] ), .Z(n13148)
         );
  XOR \SUBBYTES[6].a/U4162  ( .A(n13150), .B(n13149), .Z(\SUBBYTES[6].a/w896 )
         );
  XOR \SUBBYTES[6].a/U4161  ( .A(n12239), .B(n1040), .Z(n13149) );
  XOR \SUBBYTES[6].a/U4160  ( .A(n12238), .B(\SUBBYTES[6].a/w849 ), .Z(n13150)
         );
  XOR \SUBBYTES[6].a/U4159  ( .A(\w1[6][103] ), .B(\w1[6][98] ), .Z(n13474) );
  XOR \SUBBYTES[6].a/U4158  ( .A(n13474), .B(n13151), .Z(\SUBBYTES[6].a/w897 )
         );
  XOR \SUBBYTES[6].a/U4157  ( .A(\w1[6][101] ), .B(\w1[6][100] ), .Z(n13151)
         );
  XOR \SUBBYTES[6].a/U4156  ( .A(\w1[6][103] ), .B(\SUBBYTES[6].a/w782 ), .Z(
        \SUBBYTES[6].a/w785 ) );
  XOR \SUBBYTES[6].a/U4155  ( .A(\w1[6][97] ), .B(\SUBBYTES[6].a/w782 ), .Z(
        \SUBBYTES[6].a/w786 ) );
  XOR \SUBBYTES[6].a/U4154  ( .A(\w1[6][100] ), .B(\SUBBYTES[6].a/w782 ), .Z(
        \SUBBYTES[6].a/w787 ) );
  XOR \SUBBYTES[6].a/U4153  ( .A(\SUBBYTES[6].a/w786 ), .B(n13474), .Z(
        \SUBBYTES[6].a/w788 ) );
  XOR \SUBBYTES[6].a/U4152  ( .A(n13474), .B(n13152), .Z(\SUBBYTES[6].a/w873 )
         );
  XOR \SUBBYTES[6].a/U4151  ( .A(\w1[6][100] ), .B(\w1[6][97] ), .Z(n13152) );
  XOR \SUBBYTES[6].a/U4150  ( .A(n13154), .B(n13153), .Z(n13471) );
  XOR \SUBBYTES[6].a/U4149  ( .A(\w1[6][100] ), .B(n13155), .Z(n13153) );
  XOR \SUBBYTES[6].a/U4148  ( .A(\SUBBYTES[6].a/w838 ), .B(\w1[6][102] ), .Z(
        n13154) );
  XOR \SUBBYTES[6].a/U4147  ( .A(\SUBBYTES[6].a/w812 ), .B(
        \SUBBYTES[6].a/w819 ), .Z(n13155) );
  XOR \SUBBYTES[6].a/U4146  ( .A(n13157), .B(n13156), .Z(n13469) );
  XOR \SUBBYTES[6].a/U4145  ( .A(\w1[6][97] ), .B(n13158), .Z(n13156) );
  XOR \SUBBYTES[6].a/U4144  ( .A(\SUBBYTES[6].a/w837 ), .B(\w1[6][101] ), .Z(
        n13157) );
  XOR \SUBBYTES[6].a/U4143  ( .A(\SUBBYTES[6].a/w813 ), .B(
        \SUBBYTES[6].a/w820 ), .Z(n13158) );
  XOR \SUBBYTES[6].a/U4142  ( .A(n13471), .B(n13469), .Z(\SUBBYTES[6].a/w843 )
         );
  XOR \SUBBYTES[6].a/U4141  ( .A(\w1[6][101] ), .B(n13159), .Z(n13472) );
  XOR \SUBBYTES[6].a/U4140  ( .A(\SUBBYTES[6].a/w805 ), .B(
        \SUBBYTES[6].a/w815 ), .Z(n13159) );
  XOR \SUBBYTES[6].a/U4139  ( .A(n13161), .B(n13160), .Z(\SUBBYTES[6].a/w830 )
         );
  XOR \SUBBYTES[6].a/U4138  ( .A(n13472), .B(n13162), .Z(n13160) );
  XOR \SUBBYTES[6].a/U4137  ( .A(\w1[6][100] ), .B(\SUBBYTES[6].a/w894 ), .Z(
        n13161) );
  XOR \SUBBYTES[6].a/U4136  ( .A(\SUBBYTES[6].a/w807 ), .B(
        \SUBBYTES[6].a/w812 ), .Z(n13162) );
  XOR \SUBBYTES[6].a/U4135  ( .A(n13164), .B(n13163), .Z(n13470) );
  XOR \SUBBYTES[6].a/U4134  ( .A(\SUBBYTES[6].a/w840 ), .B(\w1[6][103] ), .Z(
        n13163) );
  XOR \SUBBYTES[6].a/U4133  ( .A(\SUBBYTES[6].a/w815 ), .B(
        \SUBBYTES[6].a/w822 ), .Z(n13164) );
  XOR \SUBBYTES[6].a/U4132  ( .A(n13469), .B(n13470), .Z(\SUBBYTES[6].a/w842 )
         );
  XOR \SUBBYTES[6].a/U4131  ( .A(\w1[6][99] ), .B(n13165), .Z(n13473) );
  XOR \SUBBYTES[6].a/U4130  ( .A(\SUBBYTES[6].a/w804 ), .B(
        \SUBBYTES[6].a/w807 ), .Z(n13165) );
  XOR \SUBBYTES[6].a/U4129  ( .A(n13167), .B(n13166), .Z(\SUBBYTES[6].a/w831 )
         );
  XOR \SUBBYTES[6].a/U4128  ( .A(n13473), .B(n13168), .Z(n13166) );
  XOR \SUBBYTES[6].a/U4127  ( .A(\w1[6][102] ), .B(\SUBBYTES[6].a/w873 ), .Z(
        n13167) );
  XOR \SUBBYTES[6].a/U4126  ( .A(\SUBBYTES[6].a/w812 ), .B(
        \SUBBYTES[6].a/w813 ), .Z(n13168) );
  XOR \SUBBYTES[6].a/U4125  ( .A(n13471), .B(n13470), .Z(\SUBBYTES[6].a/w851 )
         );
  XOR \SUBBYTES[6].a/U4124  ( .A(n13170), .B(n13169), .Z(\SUBBYTES[6].a/w852 )
         );
  XOR \SUBBYTES[6].a/U4123  ( .A(\w1[6][103] ), .B(n13472), .Z(n13169) );
  XOR \SUBBYTES[6].a/U4122  ( .A(\SUBBYTES[6].a/w804 ), .B(
        \SUBBYTES[6].a/w813 ), .Z(n13170) );
  XOR \SUBBYTES[6].a/U4121  ( .A(n13172), .B(n13171), .Z(\SUBBYTES[6].a/w828 )
         );
  XOR \SUBBYTES[6].a/U4120  ( .A(n13174), .B(n13173), .Z(n13171) );
  XOR \SUBBYTES[6].a/U4119  ( .A(\w1[6][103] ), .B(\SUBBYTES[6].a/w912 ), .Z(
        n13172) );
  XOR \SUBBYTES[6].a/U4118  ( .A(\SUBBYTES[6].a/w819 ), .B(
        \SUBBYTES[6].a/w822 ), .Z(n13173) );
  XOR \SUBBYTES[6].a/U4117  ( .A(\SUBBYTES[6].a/w805 ), .B(
        \SUBBYTES[6].a/w807 ), .Z(n13174) );
  XOR \SUBBYTES[6].a/U4116  ( .A(n13176), .B(n13175), .Z(\SUBBYTES[6].a/w829 )
         );
  XOR \SUBBYTES[6].a/U4115  ( .A(n13473), .B(n13177), .Z(n13175) );
  XOR \SUBBYTES[6].a/U4114  ( .A(\w1[6][101] ), .B(n13474), .Z(n13176) );
  XOR \SUBBYTES[6].a/U4113  ( .A(\SUBBYTES[6].a/w819 ), .B(
        \SUBBYTES[6].a/w820 ), .Z(n13177) );
  XOR \SUBBYTES[6].a/U4112  ( .A(n13179), .B(n13178), .Z(\SUBBYTES[6].a/w845 )
         );
  XOR \SUBBYTES[6].a/U4111  ( .A(\w1[6][97] ), .B(n13180), .Z(n13178) );
  XOR \SUBBYTES[6].a/U4110  ( .A(\SUBBYTES[6].a/w820 ), .B(
        \SUBBYTES[6].a/w822 ), .Z(n13179) );
  XOR \SUBBYTES[6].a/U4109  ( .A(\SUBBYTES[6].a/w804 ), .B(
        \SUBBYTES[6].a/w805 ), .Z(n13180) );
  XOR \SUBBYTES[6].a/U4108  ( .A(\w1[6][105] ), .B(n13181), .Z(n13475) );
  XOR \SUBBYTES[6].a/U4107  ( .A(\w1[6][107] ), .B(\w1[6][106] ), .Z(n13181)
         );
  XOR \SUBBYTES[6].a/U4106  ( .A(\w1[6][110] ), .B(n13475), .Z(
        \SUBBYTES[6].a/w687 ) );
  XOR \SUBBYTES[6].a/U4105  ( .A(\w1[6][104] ), .B(\SUBBYTES[6].a/w687 ), .Z(
        \SUBBYTES[6].a/w574 ) );
  XOR \SUBBYTES[6].a/U4104  ( .A(\w1[6][104] ), .B(n13182), .Z(
        \SUBBYTES[6].a/w575 ) );
  XOR \SUBBYTES[6].a/U4103  ( .A(\w1[6][110] ), .B(\w1[6][109] ), .Z(n13182)
         );
  XOR \SUBBYTES[6].a/U4102  ( .A(\w1[6][109] ), .B(n13475), .Z(
        \SUBBYTES[6].a/w705 ) );
  XOR \SUBBYTES[6].a/U4101  ( .A(n13184), .B(n13183), .Z(\SUBBYTES[6].a/w698 )
         );
  XOR \SUBBYTES[6].a/U4100  ( .A(\w1[6][107] ), .B(\w1[6][105] ), .Z(n13183)
         );
  XOR \SUBBYTES[6].a/U4099  ( .A(\w1[6][111] ), .B(\w1[6][108] ), .Z(n13184)
         );
  XOR \SUBBYTES[6].a/U4098  ( .A(\w1[6][104] ), .B(\SUBBYTES[6].a/w698 ), .Z(
        \SUBBYTES[6].a/w577 ) );
  XOR \SUBBYTES[6].a/U4097  ( .A(n13186), .B(n13185), .Z(\SUBBYTES[6].a/w685 )
         );
  XOR \SUBBYTES[6].a/U4096  ( .A(\SUBBYTES[6].a/w646 ), .B(n1039), .Z(n13185)
         );
  XOR \SUBBYTES[6].a/U4095  ( .A(\SUBBYTES[6].a/w639 ), .B(
        \SUBBYTES[6].a/w642 ), .Z(n13186) );
  XOR \SUBBYTES[6].a/U4094  ( .A(n13188), .B(n13187), .Z(\SUBBYTES[6].a/w686 )
         );
  XOR \SUBBYTES[6].a/U4093  ( .A(\SUBBYTES[6].a/w646 ), .B(n12237), .Z(n13187)
         );
  XOR \SUBBYTES[6].a/U4092  ( .A(\SUBBYTES[6].a/w639 ), .B(n12236), .Z(n13188)
         );
  XOR \SUBBYTES[6].a/U4091  ( .A(\SUBBYTES[6].a/w698 ), .B(n13189), .Z(
        \SUBBYTES[6].a/w688 ) );
  XOR \SUBBYTES[6].a/U4090  ( .A(\w1[6][110] ), .B(\w1[6][109] ), .Z(n13189)
         );
  XOR \SUBBYTES[6].a/U4089  ( .A(n13191), .B(n13190), .Z(\SUBBYTES[6].a/w689 )
         );
  XOR \SUBBYTES[6].a/U4088  ( .A(n12237), .B(n1039), .Z(n13190) );
  XOR \SUBBYTES[6].a/U4087  ( .A(n12236), .B(\SUBBYTES[6].a/w642 ), .Z(n13191)
         );
  XOR \SUBBYTES[6].a/U4086  ( .A(\w1[6][111] ), .B(\w1[6][106] ), .Z(n13481)
         );
  XOR \SUBBYTES[6].a/U4085  ( .A(n13481), .B(n13192), .Z(\SUBBYTES[6].a/w690 )
         );
  XOR \SUBBYTES[6].a/U4084  ( .A(\w1[6][109] ), .B(\w1[6][108] ), .Z(n13192)
         );
  XOR \SUBBYTES[6].a/U4083  ( .A(\w1[6][111] ), .B(\SUBBYTES[6].a/w575 ), .Z(
        \SUBBYTES[6].a/w578 ) );
  XOR \SUBBYTES[6].a/U4082  ( .A(\w1[6][105] ), .B(\SUBBYTES[6].a/w575 ), .Z(
        \SUBBYTES[6].a/w579 ) );
  XOR \SUBBYTES[6].a/U4081  ( .A(\w1[6][108] ), .B(\SUBBYTES[6].a/w575 ), .Z(
        \SUBBYTES[6].a/w580 ) );
  XOR \SUBBYTES[6].a/U4080  ( .A(\SUBBYTES[6].a/w579 ), .B(n13481), .Z(
        \SUBBYTES[6].a/w581 ) );
  XOR \SUBBYTES[6].a/U4079  ( .A(n13481), .B(n13193), .Z(\SUBBYTES[6].a/w666 )
         );
  XOR \SUBBYTES[6].a/U4078  ( .A(\w1[6][108] ), .B(\w1[6][105] ), .Z(n13193)
         );
  XOR \SUBBYTES[6].a/U4077  ( .A(n13195), .B(n13194), .Z(n13478) );
  XOR \SUBBYTES[6].a/U4076  ( .A(\w1[6][108] ), .B(n13196), .Z(n13194) );
  XOR \SUBBYTES[6].a/U4075  ( .A(\SUBBYTES[6].a/w631 ), .B(\w1[6][110] ), .Z(
        n13195) );
  XOR \SUBBYTES[6].a/U4074  ( .A(\SUBBYTES[6].a/w605 ), .B(
        \SUBBYTES[6].a/w612 ), .Z(n13196) );
  XOR \SUBBYTES[6].a/U4073  ( .A(n13198), .B(n13197), .Z(n13476) );
  XOR \SUBBYTES[6].a/U4072  ( .A(\w1[6][105] ), .B(n13199), .Z(n13197) );
  XOR \SUBBYTES[6].a/U4071  ( .A(\SUBBYTES[6].a/w630 ), .B(\w1[6][109] ), .Z(
        n13198) );
  XOR \SUBBYTES[6].a/U4070  ( .A(\SUBBYTES[6].a/w606 ), .B(
        \SUBBYTES[6].a/w613 ), .Z(n13199) );
  XOR \SUBBYTES[6].a/U4069  ( .A(n13478), .B(n13476), .Z(\SUBBYTES[6].a/w636 )
         );
  XOR \SUBBYTES[6].a/U4068  ( .A(\w1[6][109] ), .B(n13200), .Z(n13479) );
  XOR \SUBBYTES[6].a/U4067  ( .A(\SUBBYTES[6].a/w598 ), .B(
        \SUBBYTES[6].a/w608 ), .Z(n13200) );
  XOR \SUBBYTES[6].a/U4066  ( .A(n13202), .B(n13201), .Z(\SUBBYTES[6].a/w623 )
         );
  XOR \SUBBYTES[6].a/U4065  ( .A(n13479), .B(n13203), .Z(n13201) );
  XOR \SUBBYTES[6].a/U4064  ( .A(\w1[6][108] ), .B(\SUBBYTES[6].a/w687 ), .Z(
        n13202) );
  XOR \SUBBYTES[6].a/U4063  ( .A(\SUBBYTES[6].a/w600 ), .B(
        \SUBBYTES[6].a/w605 ), .Z(n13203) );
  XOR \SUBBYTES[6].a/U4062  ( .A(n13205), .B(n13204), .Z(n13477) );
  XOR \SUBBYTES[6].a/U4061  ( .A(\SUBBYTES[6].a/w633 ), .B(\w1[6][111] ), .Z(
        n13204) );
  XOR \SUBBYTES[6].a/U4060  ( .A(\SUBBYTES[6].a/w608 ), .B(
        \SUBBYTES[6].a/w615 ), .Z(n13205) );
  XOR \SUBBYTES[6].a/U4059  ( .A(n13476), .B(n13477), .Z(\SUBBYTES[6].a/w635 )
         );
  XOR \SUBBYTES[6].a/U4058  ( .A(\w1[6][107] ), .B(n13206), .Z(n13480) );
  XOR \SUBBYTES[6].a/U4057  ( .A(\SUBBYTES[6].a/w597 ), .B(
        \SUBBYTES[6].a/w600 ), .Z(n13206) );
  XOR \SUBBYTES[6].a/U4056  ( .A(n13208), .B(n13207), .Z(\SUBBYTES[6].a/w624 )
         );
  XOR \SUBBYTES[6].a/U4055  ( .A(n13480), .B(n13209), .Z(n13207) );
  XOR \SUBBYTES[6].a/U4054  ( .A(\w1[6][110] ), .B(\SUBBYTES[6].a/w666 ), .Z(
        n13208) );
  XOR \SUBBYTES[6].a/U4053  ( .A(\SUBBYTES[6].a/w605 ), .B(
        \SUBBYTES[6].a/w606 ), .Z(n13209) );
  XOR \SUBBYTES[6].a/U4052  ( .A(n13478), .B(n13477), .Z(\SUBBYTES[6].a/w644 )
         );
  XOR \SUBBYTES[6].a/U4051  ( .A(n13211), .B(n13210), .Z(\SUBBYTES[6].a/w645 )
         );
  XOR \SUBBYTES[6].a/U4050  ( .A(\w1[6][111] ), .B(n13479), .Z(n13210) );
  XOR \SUBBYTES[6].a/U4049  ( .A(\SUBBYTES[6].a/w597 ), .B(
        \SUBBYTES[6].a/w606 ), .Z(n13211) );
  XOR \SUBBYTES[6].a/U4048  ( .A(n13213), .B(n13212), .Z(\SUBBYTES[6].a/w621 )
         );
  XOR \SUBBYTES[6].a/U4047  ( .A(n13215), .B(n13214), .Z(n13212) );
  XOR \SUBBYTES[6].a/U4046  ( .A(\w1[6][111] ), .B(\SUBBYTES[6].a/w705 ), .Z(
        n13213) );
  XOR \SUBBYTES[6].a/U4045  ( .A(\SUBBYTES[6].a/w612 ), .B(
        \SUBBYTES[6].a/w615 ), .Z(n13214) );
  XOR \SUBBYTES[6].a/U4044  ( .A(\SUBBYTES[6].a/w598 ), .B(
        \SUBBYTES[6].a/w600 ), .Z(n13215) );
  XOR \SUBBYTES[6].a/U4043  ( .A(n13217), .B(n13216), .Z(\SUBBYTES[6].a/w622 )
         );
  XOR \SUBBYTES[6].a/U4042  ( .A(n13480), .B(n13218), .Z(n13216) );
  XOR \SUBBYTES[6].a/U4041  ( .A(\w1[6][109] ), .B(n13481), .Z(n13217) );
  XOR \SUBBYTES[6].a/U4040  ( .A(\SUBBYTES[6].a/w612 ), .B(
        \SUBBYTES[6].a/w613 ), .Z(n13218) );
  XOR \SUBBYTES[6].a/U4039  ( .A(n13220), .B(n13219), .Z(\SUBBYTES[6].a/w638 )
         );
  XOR \SUBBYTES[6].a/U4038  ( .A(\w1[6][105] ), .B(n13221), .Z(n13219) );
  XOR \SUBBYTES[6].a/U4037  ( .A(\SUBBYTES[6].a/w613 ), .B(
        \SUBBYTES[6].a/w615 ), .Z(n13220) );
  XOR \SUBBYTES[6].a/U4036  ( .A(\SUBBYTES[6].a/w597 ), .B(
        \SUBBYTES[6].a/w598 ), .Z(n13221) );
  XOR \SUBBYTES[6].a/U4035  ( .A(\w1[6][113] ), .B(n13222), .Z(n13482) );
  XOR \SUBBYTES[6].a/U4034  ( .A(\w1[6][115] ), .B(\w1[6][114] ), .Z(n13222)
         );
  XOR \SUBBYTES[6].a/U4033  ( .A(\w1[6][118] ), .B(n13482), .Z(
        \SUBBYTES[6].a/w480 ) );
  XOR \SUBBYTES[6].a/U4032  ( .A(\w1[6][112] ), .B(\SUBBYTES[6].a/w480 ), .Z(
        \SUBBYTES[6].a/w367 ) );
  XOR \SUBBYTES[6].a/U4031  ( .A(\w1[6][112] ), .B(n13223), .Z(
        \SUBBYTES[6].a/w368 ) );
  XOR \SUBBYTES[6].a/U4030  ( .A(\w1[6][118] ), .B(\w1[6][117] ), .Z(n13223)
         );
  XOR \SUBBYTES[6].a/U4029  ( .A(\w1[6][117] ), .B(n13482), .Z(
        \SUBBYTES[6].a/w498 ) );
  XOR \SUBBYTES[6].a/U4028  ( .A(n13225), .B(n13224), .Z(\SUBBYTES[6].a/w491 )
         );
  XOR \SUBBYTES[6].a/U4027  ( .A(\w1[6][115] ), .B(\w1[6][113] ), .Z(n13224)
         );
  XOR \SUBBYTES[6].a/U4026  ( .A(\w1[6][119] ), .B(\w1[6][116] ), .Z(n13225)
         );
  XOR \SUBBYTES[6].a/U4025  ( .A(\w1[6][112] ), .B(\SUBBYTES[6].a/w491 ), .Z(
        \SUBBYTES[6].a/w370 ) );
  XOR \SUBBYTES[6].a/U4024  ( .A(n13227), .B(n13226), .Z(\SUBBYTES[6].a/w478 )
         );
  XOR \SUBBYTES[6].a/U4023  ( .A(\SUBBYTES[6].a/w439 ), .B(n1038), .Z(n13226)
         );
  XOR \SUBBYTES[6].a/U4022  ( .A(\SUBBYTES[6].a/w432 ), .B(
        \SUBBYTES[6].a/w435 ), .Z(n13227) );
  XOR \SUBBYTES[6].a/U4021  ( .A(n13229), .B(n13228), .Z(\SUBBYTES[6].a/w479 )
         );
  XOR \SUBBYTES[6].a/U4020  ( .A(\SUBBYTES[6].a/w439 ), .B(n12235), .Z(n13228)
         );
  XOR \SUBBYTES[6].a/U4019  ( .A(\SUBBYTES[6].a/w432 ), .B(n12234), .Z(n13229)
         );
  XOR \SUBBYTES[6].a/U4018  ( .A(\SUBBYTES[6].a/w491 ), .B(n13230), .Z(
        \SUBBYTES[6].a/w481 ) );
  XOR \SUBBYTES[6].a/U4017  ( .A(\w1[6][118] ), .B(\w1[6][117] ), .Z(n13230)
         );
  XOR \SUBBYTES[6].a/U4016  ( .A(n13232), .B(n13231), .Z(\SUBBYTES[6].a/w482 )
         );
  XOR \SUBBYTES[6].a/U4015  ( .A(n12235), .B(n1038), .Z(n13231) );
  XOR \SUBBYTES[6].a/U4014  ( .A(n12234), .B(\SUBBYTES[6].a/w435 ), .Z(n13232)
         );
  XOR \SUBBYTES[6].a/U4013  ( .A(\w1[6][119] ), .B(\w1[6][114] ), .Z(n13488)
         );
  XOR \SUBBYTES[6].a/U4012  ( .A(n13488), .B(n13233), .Z(\SUBBYTES[6].a/w483 )
         );
  XOR \SUBBYTES[6].a/U4011  ( .A(\w1[6][117] ), .B(\w1[6][116] ), .Z(n13233)
         );
  XOR \SUBBYTES[6].a/U4010  ( .A(\w1[6][119] ), .B(\SUBBYTES[6].a/w368 ), .Z(
        \SUBBYTES[6].a/w371 ) );
  XOR \SUBBYTES[6].a/U4009  ( .A(\w1[6][113] ), .B(\SUBBYTES[6].a/w368 ), .Z(
        \SUBBYTES[6].a/w372 ) );
  XOR \SUBBYTES[6].a/U4008  ( .A(\w1[6][116] ), .B(\SUBBYTES[6].a/w368 ), .Z(
        \SUBBYTES[6].a/w373 ) );
  XOR \SUBBYTES[6].a/U4007  ( .A(\SUBBYTES[6].a/w372 ), .B(n13488), .Z(
        \SUBBYTES[6].a/w374 ) );
  XOR \SUBBYTES[6].a/U4006  ( .A(n13488), .B(n13234), .Z(\SUBBYTES[6].a/w459 )
         );
  XOR \SUBBYTES[6].a/U4005  ( .A(\w1[6][116] ), .B(\w1[6][113] ), .Z(n13234)
         );
  XOR \SUBBYTES[6].a/U4004  ( .A(n13236), .B(n13235), .Z(n13485) );
  XOR \SUBBYTES[6].a/U4003  ( .A(\w1[6][116] ), .B(n13237), .Z(n13235) );
  XOR \SUBBYTES[6].a/U4002  ( .A(\SUBBYTES[6].a/w424 ), .B(\w1[6][118] ), .Z(
        n13236) );
  XOR \SUBBYTES[6].a/U4001  ( .A(\SUBBYTES[6].a/w398 ), .B(
        \SUBBYTES[6].a/w405 ), .Z(n13237) );
  XOR \SUBBYTES[6].a/U4000  ( .A(n13239), .B(n13238), .Z(n13483) );
  XOR \SUBBYTES[6].a/U3999  ( .A(\w1[6][113] ), .B(n13240), .Z(n13238) );
  XOR \SUBBYTES[6].a/U3998  ( .A(\SUBBYTES[6].a/w423 ), .B(\w1[6][117] ), .Z(
        n13239) );
  XOR \SUBBYTES[6].a/U3997  ( .A(\SUBBYTES[6].a/w399 ), .B(
        \SUBBYTES[6].a/w406 ), .Z(n13240) );
  XOR \SUBBYTES[6].a/U3996  ( .A(n13485), .B(n13483), .Z(\SUBBYTES[6].a/w429 )
         );
  XOR \SUBBYTES[6].a/U3995  ( .A(\w1[6][117] ), .B(n13241), .Z(n13486) );
  XOR \SUBBYTES[6].a/U3994  ( .A(\SUBBYTES[6].a/w391 ), .B(
        \SUBBYTES[6].a/w401 ), .Z(n13241) );
  XOR \SUBBYTES[6].a/U3993  ( .A(n13243), .B(n13242), .Z(\SUBBYTES[6].a/w416 )
         );
  XOR \SUBBYTES[6].a/U3992  ( .A(n13486), .B(n13244), .Z(n13242) );
  XOR \SUBBYTES[6].a/U3991  ( .A(\w1[6][116] ), .B(\SUBBYTES[6].a/w480 ), .Z(
        n13243) );
  XOR \SUBBYTES[6].a/U3990  ( .A(\SUBBYTES[6].a/w393 ), .B(
        \SUBBYTES[6].a/w398 ), .Z(n13244) );
  XOR \SUBBYTES[6].a/U3989  ( .A(n13246), .B(n13245), .Z(n13484) );
  XOR \SUBBYTES[6].a/U3988  ( .A(\SUBBYTES[6].a/w426 ), .B(\w1[6][119] ), .Z(
        n13245) );
  XOR \SUBBYTES[6].a/U3987  ( .A(\SUBBYTES[6].a/w401 ), .B(
        \SUBBYTES[6].a/w408 ), .Z(n13246) );
  XOR \SUBBYTES[6].a/U3986  ( .A(n13483), .B(n13484), .Z(\SUBBYTES[6].a/w428 )
         );
  XOR \SUBBYTES[6].a/U3985  ( .A(\w1[6][115] ), .B(n13247), .Z(n13487) );
  XOR \SUBBYTES[6].a/U3984  ( .A(\SUBBYTES[6].a/w390 ), .B(
        \SUBBYTES[6].a/w393 ), .Z(n13247) );
  XOR \SUBBYTES[6].a/U3983  ( .A(n13249), .B(n13248), .Z(\SUBBYTES[6].a/w417 )
         );
  XOR \SUBBYTES[6].a/U3982  ( .A(n13487), .B(n13250), .Z(n13248) );
  XOR \SUBBYTES[6].a/U3981  ( .A(\w1[6][118] ), .B(\SUBBYTES[6].a/w459 ), .Z(
        n13249) );
  XOR \SUBBYTES[6].a/U3980  ( .A(\SUBBYTES[6].a/w398 ), .B(
        \SUBBYTES[6].a/w399 ), .Z(n13250) );
  XOR \SUBBYTES[6].a/U3979  ( .A(n13485), .B(n13484), .Z(\SUBBYTES[6].a/w437 )
         );
  XOR \SUBBYTES[6].a/U3978  ( .A(n13252), .B(n13251), .Z(\SUBBYTES[6].a/w438 )
         );
  XOR \SUBBYTES[6].a/U3977  ( .A(\w1[6][119] ), .B(n13486), .Z(n13251) );
  XOR \SUBBYTES[6].a/U3976  ( .A(\SUBBYTES[6].a/w390 ), .B(
        \SUBBYTES[6].a/w399 ), .Z(n13252) );
  XOR \SUBBYTES[6].a/U3975  ( .A(n13254), .B(n13253), .Z(\SUBBYTES[6].a/w414 )
         );
  XOR \SUBBYTES[6].a/U3974  ( .A(n13256), .B(n13255), .Z(n13253) );
  XOR \SUBBYTES[6].a/U3973  ( .A(\w1[6][119] ), .B(\SUBBYTES[6].a/w498 ), .Z(
        n13254) );
  XOR \SUBBYTES[6].a/U3972  ( .A(\SUBBYTES[6].a/w405 ), .B(
        \SUBBYTES[6].a/w408 ), .Z(n13255) );
  XOR \SUBBYTES[6].a/U3971  ( .A(\SUBBYTES[6].a/w391 ), .B(
        \SUBBYTES[6].a/w393 ), .Z(n13256) );
  XOR \SUBBYTES[6].a/U3970  ( .A(n13258), .B(n13257), .Z(\SUBBYTES[6].a/w415 )
         );
  XOR \SUBBYTES[6].a/U3969  ( .A(n13487), .B(n13259), .Z(n13257) );
  XOR \SUBBYTES[6].a/U3968  ( .A(\w1[6][117] ), .B(n13488), .Z(n13258) );
  XOR \SUBBYTES[6].a/U3967  ( .A(\SUBBYTES[6].a/w405 ), .B(
        \SUBBYTES[6].a/w406 ), .Z(n13259) );
  XOR \SUBBYTES[6].a/U3966  ( .A(n13261), .B(n13260), .Z(\SUBBYTES[6].a/w431 )
         );
  XOR \SUBBYTES[6].a/U3965  ( .A(\w1[6][113] ), .B(n13262), .Z(n13260) );
  XOR \SUBBYTES[6].a/U3964  ( .A(\SUBBYTES[6].a/w406 ), .B(
        \SUBBYTES[6].a/w408 ), .Z(n13261) );
  XOR \SUBBYTES[6].a/U3963  ( .A(\SUBBYTES[6].a/w390 ), .B(
        \SUBBYTES[6].a/w391 ), .Z(n13262) );
  XOR \SUBBYTES[6].a/U3962  ( .A(\w1[6][121] ), .B(n13263), .Z(n13489) );
  XOR \SUBBYTES[6].a/U3961  ( .A(\w1[6][123] ), .B(\w1[6][122] ), .Z(n13263)
         );
  XOR \SUBBYTES[6].a/U3960  ( .A(\w1[6][126] ), .B(n13489), .Z(
        \SUBBYTES[6].a/w273 ) );
  XOR \SUBBYTES[6].a/U3959  ( .A(\w1[6][120] ), .B(\SUBBYTES[6].a/w273 ), .Z(
        \SUBBYTES[6].a/w160 ) );
  XOR \SUBBYTES[6].a/U3958  ( .A(\w1[6][120] ), .B(n13264), .Z(
        \SUBBYTES[6].a/w161 ) );
  XOR \SUBBYTES[6].a/U3957  ( .A(\w1[6][126] ), .B(\w1[6][125] ), .Z(n13264)
         );
  XOR \SUBBYTES[6].a/U3956  ( .A(\w1[6][125] ), .B(n13489), .Z(
        \SUBBYTES[6].a/w291 ) );
  XOR \SUBBYTES[6].a/U3955  ( .A(n13266), .B(n13265), .Z(\SUBBYTES[6].a/w284 )
         );
  XOR \SUBBYTES[6].a/U3954  ( .A(\w1[6][123] ), .B(\w1[6][121] ), .Z(n13265)
         );
  XOR \SUBBYTES[6].a/U3953  ( .A(\w1[6][127] ), .B(\w1[6][124] ), .Z(n13266)
         );
  XOR \SUBBYTES[6].a/U3952  ( .A(\w1[6][120] ), .B(\SUBBYTES[6].a/w284 ), .Z(
        \SUBBYTES[6].a/w163 ) );
  XOR \SUBBYTES[6].a/U3951  ( .A(n13268), .B(n13267), .Z(\SUBBYTES[6].a/w271 )
         );
  XOR \SUBBYTES[6].a/U3950  ( .A(\SUBBYTES[6].a/w232 ), .B(n1037), .Z(n13267)
         );
  XOR \SUBBYTES[6].a/U3949  ( .A(\SUBBYTES[6].a/w225 ), .B(
        \SUBBYTES[6].a/w228 ), .Z(n13268) );
  XOR \SUBBYTES[6].a/U3948  ( .A(n13270), .B(n13269), .Z(\SUBBYTES[6].a/w272 )
         );
  XOR \SUBBYTES[6].a/U3947  ( .A(\SUBBYTES[6].a/w232 ), .B(n12233), .Z(n13269)
         );
  XOR \SUBBYTES[6].a/U3946  ( .A(\SUBBYTES[6].a/w225 ), .B(n12232), .Z(n13270)
         );
  XOR \SUBBYTES[6].a/U3945  ( .A(\SUBBYTES[6].a/w284 ), .B(n13271), .Z(
        \SUBBYTES[6].a/w274 ) );
  XOR \SUBBYTES[6].a/U3944  ( .A(\w1[6][126] ), .B(\w1[6][125] ), .Z(n13271)
         );
  XOR \SUBBYTES[6].a/U3943  ( .A(n13273), .B(n13272), .Z(\SUBBYTES[6].a/w275 )
         );
  XOR \SUBBYTES[6].a/U3942  ( .A(n12233), .B(n1037), .Z(n13272) );
  XOR \SUBBYTES[6].a/U3941  ( .A(n12232), .B(\SUBBYTES[6].a/w228 ), .Z(n13273)
         );
  XOR \SUBBYTES[6].a/U3940  ( .A(\w1[6][127] ), .B(\w1[6][122] ), .Z(n13495)
         );
  XOR \SUBBYTES[6].a/U3939  ( .A(n13495), .B(n13274), .Z(\SUBBYTES[6].a/w276 )
         );
  XOR \SUBBYTES[6].a/U3938  ( .A(\w1[6][125] ), .B(\w1[6][124] ), .Z(n13274)
         );
  XOR \SUBBYTES[6].a/U3937  ( .A(\w1[6][127] ), .B(\SUBBYTES[6].a/w161 ), .Z(
        \SUBBYTES[6].a/w164 ) );
  XOR \SUBBYTES[6].a/U3936  ( .A(\w1[6][121] ), .B(\SUBBYTES[6].a/w161 ), .Z(
        \SUBBYTES[6].a/w165 ) );
  XOR \SUBBYTES[6].a/U3935  ( .A(\w1[6][124] ), .B(\SUBBYTES[6].a/w161 ), .Z(
        \SUBBYTES[6].a/w166 ) );
  XOR \SUBBYTES[6].a/U3934  ( .A(\SUBBYTES[6].a/w165 ), .B(n13495), .Z(
        \SUBBYTES[6].a/w167 ) );
  XOR \SUBBYTES[6].a/U3933  ( .A(n13495), .B(n13275), .Z(\SUBBYTES[6].a/w252 )
         );
  XOR \SUBBYTES[6].a/U3932  ( .A(\w1[6][124] ), .B(\w1[6][121] ), .Z(n13275)
         );
  XOR \SUBBYTES[6].a/U3931  ( .A(n13277), .B(n13276), .Z(n13492) );
  XOR \SUBBYTES[6].a/U3930  ( .A(\w1[6][124] ), .B(n13278), .Z(n13276) );
  XOR \SUBBYTES[6].a/U3929  ( .A(\SUBBYTES[6].a/w217 ), .B(\w1[6][126] ), .Z(
        n13277) );
  XOR \SUBBYTES[6].a/U3928  ( .A(\SUBBYTES[6].a/w191 ), .B(
        \SUBBYTES[6].a/w198 ), .Z(n13278) );
  XOR \SUBBYTES[6].a/U3927  ( .A(n13280), .B(n13279), .Z(n13490) );
  XOR \SUBBYTES[6].a/U3926  ( .A(\w1[6][121] ), .B(n13281), .Z(n13279) );
  XOR \SUBBYTES[6].a/U3925  ( .A(\SUBBYTES[6].a/w216 ), .B(\w1[6][125] ), .Z(
        n13280) );
  XOR \SUBBYTES[6].a/U3924  ( .A(\SUBBYTES[6].a/w192 ), .B(
        \SUBBYTES[6].a/w199 ), .Z(n13281) );
  XOR \SUBBYTES[6].a/U3923  ( .A(n13492), .B(n13490), .Z(\SUBBYTES[6].a/w222 )
         );
  XOR \SUBBYTES[6].a/U3922  ( .A(\w1[6][125] ), .B(n13282), .Z(n13493) );
  XOR \SUBBYTES[6].a/U3921  ( .A(\SUBBYTES[6].a/w184 ), .B(
        \SUBBYTES[6].a/w194 ), .Z(n13282) );
  XOR \SUBBYTES[6].a/U3920  ( .A(n13284), .B(n13283), .Z(\SUBBYTES[6].a/w209 )
         );
  XOR \SUBBYTES[6].a/U3919  ( .A(n13493), .B(n13285), .Z(n13283) );
  XOR \SUBBYTES[6].a/U3918  ( .A(\w1[6][124] ), .B(\SUBBYTES[6].a/w273 ), .Z(
        n13284) );
  XOR \SUBBYTES[6].a/U3917  ( .A(\SUBBYTES[6].a/w186 ), .B(
        \SUBBYTES[6].a/w191 ), .Z(n13285) );
  XOR \SUBBYTES[6].a/U3916  ( .A(n13287), .B(n13286), .Z(n13491) );
  XOR \SUBBYTES[6].a/U3915  ( .A(\SUBBYTES[6].a/w219 ), .B(\w1[6][127] ), .Z(
        n13286) );
  XOR \SUBBYTES[6].a/U3914  ( .A(\SUBBYTES[6].a/w194 ), .B(
        \SUBBYTES[6].a/w201 ), .Z(n13287) );
  XOR \SUBBYTES[6].a/U3913  ( .A(n13490), .B(n13491), .Z(\SUBBYTES[6].a/w221 )
         );
  XOR \SUBBYTES[6].a/U3912  ( .A(\w1[6][123] ), .B(n13288), .Z(n13494) );
  XOR \SUBBYTES[6].a/U3911  ( .A(\SUBBYTES[6].a/w183 ), .B(
        \SUBBYTES[6].a/w186 ), .Z(n13288) );
  XOR \SUBBYTES[6].a/U3910  ( .A(n13290), .B(n13289), .Z(\SUBBYTES[6].a/w210 )
         );
  XOR \SUBBYTES[6].a/U3909  ( .A(n13494), .B(n13291), .Z(n13289) );
  XOR \SUBBYTES[6].a/U3908  ( .A(\w1[6][126] ), .B(\SUBBYTES[6].a/w252 ), .Z(
        n13290) );
  XOR \SUBBYTES[6].a/U3907  ( .A(\SUBBYTES[6].a/w191 ), .B(
        \SUBBYTES[6].a/w192 ), .Z(n13291) );
  XOR \SUBBYTES[6].a/U3906  ( .A(n13492), .B(n13491), .Z(\SUBBYTES[6].a/w230 )
         );
  XOR \SUBBYTES[6].a/U3905  ( .A(n13293), .B(n13292), .Z(\SUBBYTES[6].a/w231 )
         );
  XOR \SUBBYTES[6].a/U3904  ( .A(\w1[6][127] ), .B(n13493), .Z(n13292) );
  XOR \SUBBYTES[6].a/U3903  ( .A(\SUBBYTES[6].a/w183 ), .B(
        \SUBBYTES[6].a/w192 ), .Z(n13293) );
  XOR \SUBBYTES[6].a/U3902  ( .A(n13295), .B(n13294), .Z(\SUBBYTES[6].a/w207 )
         );
  XOR \SUBBYTES[6].a/U3901  ( .A(n13297), .B(n13296), .Z(n13294) );
  XOR \SUBBYTES[6].a/U3900  ( .A(\w1[6][127] ), .B(\SUBBYTES[6].a/w291 ), .Z(
        n13295) );
  XOR \SUBBYTES[6].a/U3899  ( .A(\SUBBYTES[6].a/w198 ), .B(
        \SUBBYTES[6].a/w201 ), .Z(n13296) );
  XOR \SUBBYTES[6].a/U3898  ( .A(\SUBBYTES[6].a/w184 ), .B(
        \SUBBYTES[6].a/w186 ), .Z(n13297) );
  XOR \SUBBYTES[6].a/U3897  ( .A(n13299), .B(n13298), .Z(\SUBBYTES[6].a/w208 )
         );
  XOR \SUBBYTES[6].a/U3896  ( .A(n13494), .B(n13300), .Z(n13298) );
  XOR \SUBBYTES[6].a/U3895  ( .A(\w1[6][125] ), .B(n13495), .Z(n13299) );
  XOR \SUBBYTES[6].a/U3894  ( .A(\SUBBYTES[6].a/w198 ), .B(
        \SUBBYTES[6].a/w199 ), .Z(n13300) );
  XOR \SUBBYTES[6].a/U3893  ( .A(n13302), .B(n13301), .Z(\SUBBYTES[6].a/w224 )
         );
  XOR \SUBBYTES[6].a/U3892  ( .A(\w1[6][121] ), .B(n13303), .Z(n13301) );
  XOR \SUBBYTES[6].a/U3891  ( .A(\SUBBYTES[6].a/w199 ), .B(
        \SUBBYTES[6].a/w201 ), .Z(n13302) );
  XOR \SUBBYTES[6].a/U3890  ( .A(\SUBBYTES[6].a/w183 ), .B(
        \SUBBYTES[6].a/w184 ), .Z(n13303) );
  XOR \SUBBYTES[5].a/U5649  ( .A(\SUBBYTES[5].a/w3390 ), .B(
        \SUBBYTES[5].a/w3391 ), .Z(n12025) );
  XOR \SUBBYTES[5].a/U5648  ( .A(n12025), .B(n10984), .Z(n12024) );
  XOR \SUBBYTES[5].a/U5647  ( .A(\SUBBYTES[5].a/w3383 ), .B(
        \SUBBYTES[5].a/w3400 ), .Z(n10984) );
  XOR \SUBBYTES[5].a/U5645  ( .A(\SUBBYTES[5].a/w3382 ), .B(
        \SUBBYTES[5].a/w3397 ), .Z(n10985) );
  XOR \SUBBYTES[5].a/U5644  ( .A(n12025), .B(n10986), .Z(n12216) );
  XOR \SUBBYTES[5].a/U5643  ( .A(\SUBBYTES[5].a/w3397 ), .B(
        \SUBBYTES[5].a/w3398 ), .Z(n10986) );
  XOR \SUBBYTES[5].a/U5642  ( .A(\SUBBYTES[5].a/w3359 ), .B(n10987), .Z(n12027) );
  XOR \SUBBYTES[5].a/U5641  ( .A(\SUBBYTES[5].a/w3350 ), .B(
        \SUBBYTES[5].a/w3351 ), .Z(n10987) );
  XOR \SUBBYTES[5].a/U5639  ( .A(\SUBBYTES[5].a/w3361 ), .B(n12216), .Z(n10988) );
  XOR \SUBBYTES[5].a/U5638  ( .A(n10990), .B(n10989), .Z(n12028) );
  XOR \SUBBYTES[5].a/U5637  ( .A(n10992), .B(n10991), .Z(n10989) );
  XOR \SUBBYTES[5].a/U5636  ( .A(\SUBBYTES[5].a/w3397 ), .B(
        \SUBBYTES[5].a/w3398 ), .Z(n10990) );
  XOR \SUBBYTES[5].a/U5635  ( .A(\SUBBYTES[5].a/w3361 ), .B(
        \SUBBYTES[5].a/w3385 ), .Z(n10991) );
  XOR \SUBBYTES[5].a/U5634  ( .A(\SUBBYTES[5].a/w3350 ), .B(
        \SUBBYTES[5].a/w3359 ), .Z(n10992) );
  XOR \SUBBYTES[5].a/U5633  ( .A(\SUBBYTES[5].a/w3382 ), .B(n10993), .Z(n12026) );
  XOR \SUBBYTES[5].a/U5632  ( .A(\SUBBYTES[5].a/w3365 ), .B(
        \SUBBYTES[5].a/w3368 ), .Z(n10993) );
  XOR \SUBBYTES[5].a/U5630  ( .A(\SUBBYTES[5].a/w3353 ), .B(n12028), .Z(n10994) );
  XOR \SUBBYTES[5].a/U5628  ( .A(\SUBBYTES[5].a/w3385 ), .B(
        \SUBBYTES[5].a/w3398 ), .Z(n10995) );
  XOR \SUBBYTES[5].a/U5626  ( .A(n10999), .B(n10998), .Z(n10996) );
  XOR \SUBBYTES[5].a/U5625  ( .A(n11001), .B(n11000), .Z(n10997) );
  XOR \SUBBYTES[5].a/U5624  ( .A(\SUBBYTES[5].a/w3397 ), .B(
        \SUBBYTES[5].a/w3400 ), .Z(n10998) );
  XOR \SUBBYTES[5].a/U5623  ( .A(\SUBBYTES[5].a/w3390 ), .B(
        \SUBBYTES[5].a/w3393 ), .Z(n10999) );
  XOR \SUBBYTES[5].a/U5622  ( .A(\SUBBYTES[5].a/w3365 ), .B(
        \SUBBYTES[5].a/w3366 ), .Z(n11000) );
  XOR \SUBBYTES[5].a/U5621  ( .A(\SUBBYTES[5].a/w3350 ), .B(
        \SUBBYTES[5].a/w3353 ), .Z(n11001) );
  XOR \SUBBYTES[5].a/U5619  ( .A(n12025), .B(n11004), .Z(n11002) );
  XOR \SUBBYTES[5].a/U5618  ( .A(n12027), .B(n12026), .Z(n11003) );
  XOR \SUBBYTES[5].a/U5617  ( .A(\SUBBYTES[5].a/w3358 ), .B(
        \SUBBYTES[5].a/w3385 ), .Z(n11004) );
  XOR \SUBBYTES[5].a/U5615  ( .A(n12028), .B(n11007), .Z(n11005) );
  XOR \SUBBYTES[5].a/U5614  ( .A(\SUBBYTES[5].a/w3391 ), .B(
        \SUBBYTES[5].a/w3393 ), .Z(n11006) );
  XOR \SUBBYTES[5].a/U5613  ( .A(\SUBBYTES[5].a/w3351 ), .B(
        \SUBBYTES[5].a/w3383 ), .Z(n11007) );
  XOR \SUBBYTES[5].a/U5612  ( .A(\SUBBYTES[5].a/w3183 ), .B(
        \SUBBYTES[5].a/w3184 ), .Z(n12030) );
  XOR \SUBBYTES[5].a/U5611  ( .A(n12030), .B(n11008), .Z(n12029) );
  XOR \SUBBYTES[5].a/U5610  ( .A(\SUBBYTES[5].a/w3176 ), .B(
        \SUBBYTES[5].a/w3193 ), .Z(n11008) );
  XOR \SUBBYTES[5].a/U5608  ( .A(\SUBBYTES[5].a/w3175 ), .B(
        \SUBBYTES[5].a/w3190 ), .Z(n11009) );
  XOR \SUBBYTES[5].a/U5607  ( .A(n12030), .B(n11010), .Z(n12217) );
  XOR \SUBBYTES[5].a/U5606  ( .A(\SUBBYTES[5].a/w3190 ), .B(
        \SUBBYTES[5].a/w3191 ), .Z(n11010) );
  XOR \SUBBYTES[5].a/U5605  ( .A(\SUBBYTES[5].a/w3152 ), .B(n11011), .Z(n12032) );
  XOR \SUBBYTES[5].a/U5604  ( .A(\SUBBYTES[5].a/w3143 ), .B(
        \SUBBYTES[5].a/w3144 ), .Z(n11011) );
  XOR \SUBBYTES[5].a/U5602  ( .A(\SUBBYTES[5].a/w3154 ), .B(n12217), .Z(n11012) );
  XOR \SUBBYTES[5].a/U5601  ( .A(n11014), .B(n11013), .Z(n12033) );
  XOR \SUBBYTES[5].a/U5600  ( .A(n11016), .B(n11015), .Z(n11013) );
  XOR \SUBBYTES[5].a/U5599  ( .A(\SUBBYTES[5].a/w3190 ), .B(
        \SUBBYTES[5].a/w3191 ), .Z(n11014) );
  XOR \SUBBYTES[5].a/U5598  ( .A(\SUBBYTES[5].a/w3154 ), .B(
        \SUBBYTES[5].a/w3178 ), .Z(n11015) );
  XOR \SUBBYTES[5].a/U5597  ( .A(\SUBBYTES[5].a/w3143 ), .B(
        \SUBBYTES[5].a/w3152 ), .Z(n11016) );
  XOR \SUBBYTES[5].a/U5596  ( .A(\SUBBYTES[5].a/w3175 ), .B(n11017), .Z(n12031) );
  XOR \SUBBYTES[5].a/U5595  ( .A(\SUBBYTES[5].a/w3158 ), .B(
        \SUBBYTES[5].a/w3161 ), .Z(n11017) );
  XOR \SUBBYTES[5].a/U5593  ( .A(\SUBBYTES[5].a/w3146 ), .B(n12033), .Z(n11018) );
  XOR \SUBBYTES[5].a/U5591  ( .A(\SUBBYTES[5].a/w3178 ), .B(
        \SUBBYTES[5].a/w3191 ), .Z(n11019) );
  XOR \SUBBYTES[5].a/U5589  ( .A(n11023), .B(n11022), .Z(n11020) );
  XOR \SUBBYTES[5].a/U5588  ( .A(n11025), .B(n11024), .Z(n11021) );
  XOR \SUBBYTES[5].a/U5587  ( .A(\SUBBYTES[5].a/w3190 ), .B(
        \SUBBYTES[5].a/w3193 ), .Z(n11022) );
  XOR \SUBBYTES[5].a/U5586  ( .A(\SUBBYTES[5].a/w3183 ), .B(
        \SUBBYTES[5].a/w3186 ), .Z(n11023) );
  XOR \SUBBYTES[5].a/U5585  ( .A(\SUBBYTES[5].a/w3158 ), .B(
        \SUBBYTES[5].a/w3159 ), .Z(n11024) );
  XOR \SUBBYTES[5].a/U5584  ( .A(\SUBBYTES[5].a/w3143 ), .B(
        \SUBBYTES[5].a/w3146 ), .Z(n11025) );
  XOR \SUBBYTES[5].a/U5582  ( .A(n12030), .B(n11028), .Z(n11026) );
  XOR \SUBBYTES[5].a/U5581  ( .A(n12032), .B(n12031), .Z(n11027) );
  XOR \SUBBYTES[5].a/U5580  ( .A(\SUBBYTES[5].a/w3151 ), .B(
        \SUBBYTES[5].a/w3178 ), .Z(n11028) );
  XOR \SUBBYTES[5].a/U5578  ( .A(n12033), .B(n11031), .Z(n11029) );
  XOR \SUBBYTES[5].a/U5577  ( .A(\SUBBYTES[5].a/w3184 ), .B(
        \SUBBYTES[5].a/w3186 ), .Z(n11030) );
  XOR \SUBBYTES[5].a/U5576  ( .A(\SUBBYTES[5].a/w3144 ), .B(
        \SUBBYTES[5].a/w3176 ), .Z(n11031) );
  XOR \SUBBYTES[5].a/U5575  ( .A(\SUBBYTES[5].a/w2976 ), .B(
        \SUBBYTES[5].a/w2977 ), .Z(n12035) );
  XOR \SUBBYTES[5].a/U5574  ( .A(n12035), .B(n11032), .Z(n12034) );
  XOR \SUBBYTES[5].a/U5573  ( .A(\SUBBYTES[5].a/w2969 ), .B(
        \SUBBYTES[5].a/w2986 ), .Z(n11032) );
  XOR \SUBBYTES[5].a/U5571  ( .A(\SUBBYTES[5].a/w2968 ), .B(
        \SUBBYTES[5].a/w2983 ), .Z(n11033) );
  XOR \SUBBYTES[5].a/U5570  ( .A(n12035), .B(n11034), .Z(n12218) );
  XOR \SUBBYTES[5].a/U5569  ( .A(\SUBBYTES[5].a/w2983 ), .B(
        \SUBBYTES[5].a/w2984 ), .Z(n11034) );
  XOR \SUBBYTES[5].a/U5568  ( .A(\SUBBYTES[5].a/w2945 ), .B(n11035), .Z(n12037) );
  XOR \SUBBYTES[5].a/U5567  ( .A(\SUBBYTES[5].a/w2936 ), .B(
        \SUBBYTES[5].a/w2937 ), .Z(n11035) );
  XOR \SUBBYTES[5].a/U5565  ( .A(\SUBBYTES[5].a/w2947 ), .B(n12218), .Z(n11036) );
  XOR \SUBBYTES[5].a/U5564  ( .A(n11038), .B(n11037), .Z(n12038) );
  XOR \SUBBYTES[5].a/U5563  ( .A(n11040), .B(n11039), .Z(n11037) );
  XOR \SUBBYTES[5].a/U5562  ( .A(\SUBBYTES[5].a/w2983 ), .B(
        \SUBBYTES[5].a/w2984 ), .Z(n11038) );
  XOR \SUBBYTES[5].a/U5561  ( .A(\SUBBYTES[5].a/w2947 ), .B(
        \SUBBYTES[5].a/w2971 ), .Z(n11039) );
  XOR \SUBBYTES[5].a/U5560  ( .A(\SUBBYTES[5].a/w2936 ), .B(
        \SUBBYTES[5].a/w2945 ), .Z(n11040) );
  XOR \SUBBYTES[5].a/U5559  ( .A(\SUBBYTES[5].a/w2968 ), .B(n11041), .Z(n12036) );
  XOR \SUBBYTES[5].a/U5558  ( .A(\SUBBYTES[5].a/w2951 ), .B(
        \SUBBYTES[5].a/w2954 ), .Z(n11041) );
  XOR \SUBBYTES[5].a/U5556  ( .A(\SUBBYTES[5].a/w2939 ), .B(n12038), .Z(n11042) );
  XOR \SUBBYTES[5].a/U5554  ( .A(\SUBBYTES[5].a/w2971 ), .B(
        \SUBBYTES[5].a/w2984 ), .Z(n11043) );
  XOR \SUBBYTES[5].a/U5552  ( .A(n11047), .B(n11046), .Z(n11044) );
  XOR \SUBBYTES[5].a/U5551  ( .A(n11049), .B(n11048), .Z(n11045) );
  XOR \SUBBYTES[5].a/U5550  ( .A(\SUBBYTES[5].a/w2983 ), .B(
        \SUBBYTES[5].a/w2986 ), .Z(n11046) );
  XOR \SUBBYTES[5].a/U5549  ( .A(\SUBBYTES[5].a/w2976 ), .B(
        \SUBBYTES[5].a/w2979 ), .Z(n11047) );
  XOR \SUBBYTES[5].a/U5548  ( .A(\SUBBYTES[5].a/w2951 ), .B(
        \SUBBYTES[5].a/w2952 ), .Z(n11048) );
  XOR \SUBBYTES[5].a/U5547  ( .A(\SUBBYTES[5].a/w2936 ), .B(
        \SUBBYTES[5].a/w2939 ), .Z(n11049) );
  XOR \SUBBYTES[5].a/U5545  ( .A(n12035), .B(n11052), .Z(n11050) );
  XOR \SUBBYTES[5].a/U5544  ( .A(n12037), .B(n12036), .Z(n11051) );
  XOR \SUBBYTES[5].a/U5543  ( .A(\SUBBYTES[5].a/w2944 ), .B(
        \SUBBYTES[5].a/w2971 ), .Z(n11052) );
  XOR \SUBBYTES[5].a/U5541  ( .A(n12038), .B(n11055), .Z(n11053) );
  XOR \SUBBYTES[5].a/U5540  ( .A(\SUBBYTES[5].a/w2977 ), .B(
        \SUBBYTES[5].a/w2979 ), .Z(n11054) );
  XOR \SUBBYTES[5].a/U5539  ( .A(\SUBBYTES[5].a/w2937 ), .B(
        \SUBBYTES[5].a/w2969 ), .Z(n11055) );
  XOR \SUBBYTES[5].a/U5538  ( .A(\SUBBYTES[5].a/w2769 ), .B(
        \SUBBYTES[5].a/w2770 ), .Z(n12040) );
  XOR \SUBBYTES[5].a/U5537  ( .A(n12040), .B(n11056), .Z(n12039) );
  XOR \SUBBYTES[5].a/U5536  ( .A(\SUBBYTES[5].a/w2762 ), .B(
        \SUBBYTES[5].a/w2779 ), .Z(n11056) );
  XOR \SUBBYTES[5].a/U5534  ( .A(\SUBBYTES[5].a/w2761 ), .B(
        \SUBBYTES[5].a/w2776 ), .Z(n11057) );
  XOR \SUBBYTES[5].a/U5533  ( .A(n12040), .B(n11058), .Z(n12219) );
  XOR \SUBBYTES[5].a/U5532  ( .A(\SUBBYTES[5].a/w2776 ), .B(
        \SUBBYTES[5].a/w2777 ), .Z(n11058) );
  XOR \SUBBYTES[5].a/U5531  ( .A(\SUBBYTES[5].a/w2738 ), .B(n11059), .Z(n12042) );
  XOR \SUBBYTES[5].a/U5530  ( .A(\SUBBYTES[5].a/w2729 ), .B(
        \SUBBYTES[5].a/w2730 ), .Z(n11059) );
  XOR \SUBBYTES[5].a/U5528  ( .A(\SUBBYTES[5].a/w2740 ), .B(n12219), .Z(n11060) );
  XOR \SUBBYTES[5].a/U5527  ( .A(n11062), .B(n11061), .Z(n12043) );
  XOR \SUBBYTES[5].a/U5526  ( .A(n11064), .B(n11063), .Z(n11061) );
  XOR \SUBBYTES[5].a/U5525  ( .A(\SUBBYTES[5].a/w2776 ), .B(
        \SUBBYTES[5].a/w2777 ), .Z(n11062) );
  XOR \SUBBYTES[5].a/U5524  ( .A(\SUBBYTES[5].a/w2740 ), .B(
        \SUBBYTES[5].a/w2764 ), .Z(n11063) );
  XOR \SUBBYTES[5].a/U5523  ( .A(\SUBBYTES[5].a/w2729 ), .B(
        \SUBBYTES[5].a/w2738 ), .Z(n11064) );
  XOR \SUBBYTES[5].a/U5522  ( .A(\SUBBYTES[5].a/w2761 ), .B(n11065), .Z(n12041) );
  XOR \SUBBYTES[5].a/U5521  ( .A(\SUBBYTES[5].a/w2744 ), .B(
        \SUBBYTES[5].a/w2747 ), .Z(n11065) );
  XOR \SUBBYTES[5].a/U5519  ( .A(\SUBBYTES[5].a/w2732 ), .B(n12043), .Z(n11066) );
  XOR \SUBBYTES[5].a/U5517  ( .A(\SUBBYTES[5].a/w2764 ), .B(
        \SUBBYTES[5].a/w2777 ), .Z(n11067) );
  XOR \SUBBYTES[5].a/U5515  ( .A(n11071), .B(n11070), .Z(n11068) );
  XOR \SUBBYTES[5].a/U5514  ( .A(n11073), .B(n11072), .Z(n11069) );
  XOR \SUBBYTES[5].a/U5513  ( .A(\SUBBYTES[5].a/w2776 ), .B(
        \SUBBYTES[5].a/w2779 ), .Z(n11070) );
  XOR \SUBBYTES[5].a/U5512  ( .A(\SUBBYTES[5].a/w2769 ), .B(
        \SUBBYTES[5].a/w2772 ), .Z(n11071) );
  XOR \SUBBYTES[5].a/U5511  ( .A(\SUBBYTES[5].a/w2744 ), .B(
        \SUBBYTES[5].a/w2745 ), .Z(n11072) );
  XOR \SUBBYTES[5].a/U5510  ( .A(\SUBBYTES[5].a/w2729 ), .B(
        \SUBBYTES[5].a/w2732 ), .Z(n11073) );
  XOR \SUBBYTES[5].a/U5508  ( .A(n12040), .B(n11076), .Z(n11074) );
  XOR \SUBBYTES[5].a/U5507  ( .A(n12042), .B(n12041), .Z(n11075) );
  XOR \SUBBYTES[5].a/U5506  ( .A(\SUBBYTES[5].a/w2737 ), .B(
        \SUBBYTES[5].a/w2764 ), .Z(n11076) );
  XOR \SUBBYTES[5].a/U5504  ( .A(n12043), .B(n11079), .Z(n11077) );
  XOR \SUBBYTES[5].a/U5503  ( .A(\SUBBYTES[5].a/w2770 ), .B(
        \SUBBYTES[5].a/w2772 ), .Z(n11078) );
  XOR \SUBBYTES[5].a/U5502  ( .A(\SUBBYTES[5].a/w2730 ), .B(
        \SUBBYTES[5].a/w2762 ), .Z(n11079) );
  XOR \SUBBYTES[5].a/U5501  ( .A(\SUBBYTES[5].a/w2562 ), .B(
        \SUBBYTES[5].a/w2563 ), .Z(n12045) );
  XOR \SUBBYTES[5].a/U5500  ( .A(n12045), .B(n11080), .Z(n12044) );
  XOR \SUBBYTES[5].a/U5499  ( .A(\SUBBYTES[5].a/w2555 ), .B(
        \SUBBYTES[5].a/w2572 ), .Z(n11080) );
  XOR \SUBBYTES[5].a/U5497  ( .A(\SUBBYTES[5].a/w2554 ), .B(
        \SUBBYTES[5].a/w2569 ), .Z(n11081) );
  XOR \SUBBYTES[5].a/U5496  ( .A(n12045), .B(n11082), .Z(n12220) );
  XOR \SUBBYTES[5].a/U5495  ( .A(\SUBBYTES[5].a/w2569 ), .B(
        \SUBBYTES[5].a/w2570 ), .Z(n11082) );
  XOR \SUBBYTES[5].a/U5494  ( .A(\SUBBYTES[5].a/w2531 ), .B(n11083), .Z(n12047) );
  XOR \SUBBYTES[5].a/U5493  ( .A(\SUBBYTES[5].a/w2522 ), .B(
        \SUBBYTES[5].a/w2523 ), .Z(n11083) );
  XOR \SUBBYTES[5].a/U5491  ( .A(\SUBBYTES[5].a/w2533 ), .B(n12220), .Z(n11084) );
  XOR \SUBBYTES[5].a/U5490  ( .A(n11086), .B(n11085), .Z(n12048) );
  XOR \SUBBYTES[5].a/U5489  ( .A(n11088), .B(n11087), .Z(n11085) );
  XOR \SUBBYTES[5].a/U5488  ( .A(\SUBBYTES[5].a/w2569 ), .B(
        \SUBBYTES[5].a/w2570 ), .Z(n11086) );
  XOR \SUBBYTES[5].a/U5487  ( .A(\SUBBYTES[5].a/w2533 ), .B(
        \SUBBYTES[5].a/w2557 ), .Z(n11087) );
  XOR \SUBBYTES[5].a/U5486  ( .A(\SUBBYTES[5].a/w2522 ), .B(
        \SUBBYTES[5].a/w2531 ), .Z(n11088) );
  XOR \SUBBYTES[5].a/U5485  ( .A(\SUBBYTES[5].a/w2554 ), .B(n11089), .Z(n12046) );
  XOR \SUBBYTES[5].a/U5484  ( .A(\SUBBYTES[5].a/w2537 ), .B(
        \SUBBYTES[5].a/w2540 ), .Z(n11089) );
  XOR \SUBBYTES[5].a/U5482  ( .A(\SUBBYTES[5].a/w2525 ), .B(n12048), .Z(n11090) );
  XOR \SUBBYTES[5].a/U5480  ( .A(\SUBBYTES[5].a/w2557 ), .B(
        \SUBBYTES[5].a/w2570 ), .Z(n11091) );
  XOR \SUBBYTES[5].a/U5478  ( .A(n11095), .B(n11094), .Z(n11092) );
  XOR \SUBBYTES[5].a/U5477  ( .A(n11097), .B(n11096), .Z(n11093) );
  XOR \SUBBYTES[5].a/U5476  ( .A(\SUBBYTES[5].a/w2569 ), .B(
        \SUBBYTES[5].a/w2572 ), .Z(n11094) );
  XOR \SUBBYTES[5].a/U5475  ( .A(\SUBBYTES[5].a/w2562 ), .B(
        \SUBBYTES[5].a/w2565 ), .Z(n11095) );
  XOR \SUBBYTES[5].a/U5474  ( .A(\SUBBYTES[5].a/w2537 ), .B(
        \SUBBYTES[5].a/w2538 ), .Z(n11096) );
  XOR \SUBBYTES[5].a/U5473  ( .A(\SUBBYTES[5].a/w2522 ), .B(
        \SUBBYTES[5].a/w2525 ), .Z(n11097) );
  XOR \SUBBYTES[5].a/U5471  ( .A(n12045), .B(n11100), .Z(n11098) );
  XOR \SUBBYTES[5].a/U5470  ( .A(n12047), .B(n12046), .Z(n11099) );
  XOR \SUBBYTES[5].a/U5469  ( .A(\SUBBYTES[5].a/w2530 ), .B(
        \SUBBYTES[5].a/w2557 ), .Z(n11100) );
  XOR \SUBBYTES[5].a/U5467  ( .A(n12048), .B(n11103), .Z(n11101) );
  XOR \SUBBYTES[5].a/U5466  ( .A(\SUBBYTES[5].a/w2563 ), .B(
        \SUBBYTES[5].a/w2565 ), .Z(n11102) );
  XOR \SUBBYTES[5].a/U5465  ( .A(\SUBBYTES[5].a/w2523 ), .B(
        \SUBBYTES[5].a/w2555 ), .Z(n11103) );
  XOR \SUBBYTES[5].a/U5464  ( .A(\SUBBYTES[5].a/w2355 ), .B(
        \SUBBYTES[5].a/w2356 ), .Z(n12050) );
  XOR \SUBBYTES[5].a/U5463  ( .A(n12050), .B(n11104), .Z(n12049) );
  XOR \SUBBYTES[5].a/U5462  ( .A(\SUBBYTES[5].a/w2348 ), .B(
        \SUBBYTES[5].a/w2365 ), .Z(n11104) );
  XOR \SUBBYTES[5].a/U5460  ( .A(\SUBBYTES[5].a/w2347 ), .B(
        \SUBBYTES[5].a/w2362 ), .Z(n11105) );
  XOR \SUBBYTES[5].a/U5459  ( .A(n12050), .B(n11106), .Z(n12221) );
  XOR \SUBBYTES[5].a/U5458  ( .A(\SUBBYTES[5].a/w2362 ), .B(
        \SUBBYTES[5].a/w2363 ), .Z(n11106) );
  XOR \SUBBYTES[5].a/U5457  ( .A(\SUBBYTES[5].a/w2324 ), .B(n11107), .Z(n12052) );
  XOR \SUBBYTES[5].a/U5456  ( .A(\SUBBYTES[5].a/w2315 ), .B(
        \SUBBYTES[5].a/w2316 ), .Z(n11107) );
  XOR \SUBBYTES[5].a/U5454  ( .A(\SUBBYTES[5].a/w2326 ), .B(n12221), .Z(n11108) );
  XOR \SUBBYTES[5].a/U5453  ( .A(n11110), .B(n11109), .Z(n12053) );
  XOR \SUBBYTES[5].a/U5452  ( .A(n11112), .B(n11111), .Z(n11109) );
  XOR \SUBBYTES[5].a/U5451  ( .A(\SUBBYTES[5].a/w2362 ), .B(
        \SUBBYTES[5].a/w2363 ), .Z(n11110) );
  XOR \SUBBYTES[5].a/U5450  ( .A(\SUBBYTES[5].a/w2326 ), .B(
        \SUBBYTES[5].a/w2350 ), .Z(n11111) );
  XOR \SUBBYTES[5].a/U5449  ( .A(\SUBBYTES[5].a/w2315 ), .B(
        \SUBBYTES[5].a/w2324 ), .Z(n11112) );
  XOR \SUBBYTES[5].a/U5448  ( .A(\SUBBYTES[5].a/w2347 ), .B(n11113), .Z(n12051) );
  XOR \SUBBYTES[5].a/U5447  ( .A(\SUBBYTES[5].a/w2330 ), .B(
        \SUBBYTES[5].a/w2333 ), .Z(n11113) );
  XOR \SUBBYTES[5].a/U5445  ( .A(\SUBBYTES[5].a/w2318 ), .B(n12053), .Z(n11114) );
  XOR \SUBBYTES[5].a/U5443  ( .A(\SUBBYTES[5].a/w2350 ), .B(
        \SUBBYTES[5].a/w2363 ), .Z(n11115) );
  XOR \SUBBYTES[5].a/U5441  ( .A(n11119), .B(n11118), .Z(n11116) );
  XOR \SUBBYTES[5].a/U5440  ( .A(n11121), .B(n11120), .Z(n11117) );
  XOR \SUBBYTES[5].a/U5439  ( .A(\SUBBYTES[5].a/w2362 ), .B(
        \SUBBYTES[5].a/w2365 ), .Z(n11118) );
  XOR \SUBBYTES[5].a/U5438  ( .A(\SUBBYTES[5].a/w2355 ), .B(
        \SUBBYTES[5].a/w2358 ), .Z(n11119) );
  XOR \SUBBYTES[5].a/U5437  ( .A(\SUBBYTES[5].a/w2330 ), .B(
        \SUBBYTES[5].a/w2331 ), .Z(n11120) );
  XOR \SUBBYTES[5].a/U5436  ( .A(\SUBBYTES[5].a/w2315 ), .B(
        \SUBBYTES[5].a/w2318 ), .Z(n11121) );
  XOR \SUBBYTES[5].a/U5434  ( .A(n12050), .B(n11124), .Z(n11122) );
  XOR \SUBBYTES[5].a/U5433  ( .A(n12052), .B(n12051), .Z(n11123) );
  XOR \SUBBYTES[5].a/U5432  ( .A(\SUBBYTES[5].a/w2323 ), .B(
        \SUBBYTES[5].a/w2350 ), .Z(n11124) );
  XOR \SUBBYTES[5].a/U5430  ( .A(n12053), .B(n11127), .Z(n11125) );
  XOR \SUBBYTES[5].a/U5429  ( .A(\SUBBYTES[5].a/w2356 ), .B(
        \SUBBYTES[5].a/w2358 ), .Z(n11126) );
  XOR \SUBBYTES[5].a/U5428  ( .A(\SUBBYTES[5].a/w2316 ), .B(
        \SUBBYTES[5].a/w2348 ), .Z(n11127) );
  XOR \SUBBYTES[5].a/U5427  ( .A(\SUBBYTES[5].a/w2148 ), .B(
        \SUBBYTES[5].a/w2149 ), .Z(n12055) );
  XOR \SUBBYTES[5].a/U5426  ( .A(n12055), .B(n11128), .Z(n12054) );
  XOR \SUBBYTES[5].a/U5425  ( .A(\SUBBYTES[5].a/w2141 ), .B(
        \SUBBYTES[5].a/w2158 ), .Z(n11128) );
  XOR \SUBBYTES[5].a/U5423  ( .A(\SUBBYTES[5].a/w2140 ), .B(
        \SUBBYTES[5].a/w2155 ), .Z(n11129) );
  XOR \SUBBYTES[5].a/U5422  ( .A(n12055), .B(n11130), .Z(n12222) );
  XOR \SUBBYTES[5].a/U5421  ( .A(\SUBBYTES[5].a/w2155 ), .B(
        \SUBBYTES[5].a/w2156 ), .Z(n11130) );
  XOR \SUBBYTES[5].a/U5420  ( .A(\SUBBYTES[5].a/w2117 ), .B(n11131), .Z(n12057) );
  XOR \SUBBYTES[5].a/U5419  ( .A(\SUBBYTES[5].a/w2108 ), .B(
        \SUBBYTES[5].a/w2109 ), .Z(n11131) );
  XOR \SUBBYTES[5].a/U5417  ( .A(\SUBBYTES[5].a/w2119 ), .B(n12222), .Z(n11132) );
  XOR \SUBBYTES[5].a/U5416  ( .A(n11134), .B(n11133), .Z(n12058) );
  XOR \SUBBYTES[5].a/U5415  ( .A(n11136), .B(n11135), .Z(n11133) );
  XOR \SUBBYTES[5].a/U5414  ( .A(\SUBBYTES[5].a/w2155 ), .B(
        \SUBBYTES[5].a/w2156 ), .Z(n11134) );
  XOR \SUBBYTES[5].a/U5413  ( .A(\SUBBYTES[5].a/w2119 ), .B(
        \SUBBYTES[5].a/w2143 ), .Z(n11135) );
  XOR \SUBBYTES[5].a/U5412  ( .A(\SUBBYTES[5].a/w2108 ), .B(
        \SUBBYTES[5].a/w2117 ), .Z(n11136) );
  XOR \SUBBYTES[5].a/U5411  ( .A(\SUBBYTES[5].a/w2140 ), .B(n11137), .Z(n12056) );
  XOR \SUBBYTES[5].a/U5410  ( .A(\SUBBYTES[5].a/w2123 ), .B(
        \SUBBYTES[5].a/w2126 ), .Z(n11137) );
  XOR \SUBBYTES[5].a/U5408  ( .A(\SUBBYTES[5].a/w2111 ), .B(n12058), .Z(n11138) );
  XOR \SUBBYTES[5].a/U5406  ( .A(\SUBBYTES[5].a/w2143 ), .B(
        \SUBBYTES[5].a/w2156 ), .Z(n11139) );
  XOR \SUBBYTES[5].a/U5404  ( .A(n11143), .B(n11142), .Z(n11140) );
  XOR \SUBBYTES[5].a/U5403  ( .A(n11145), .B(n11144), .Z(n11141) );
  XOR \SUBBYTES[5].a/U5402  ( .A(\SUBBYTES[5].a/w2155 ), .B(
        \SUBBYTES[5].a/w2158 ), .Z(n11142) );
  XOR \SUBBYTES[5].a/U5401  ( .A(\SUBBYTES[5].a/w2148 ), .B(
        \SUBBYTES[5].a/w2151 ), .Z(n11143) );
  XOR \SUBBYTES[5].a/U5400  ( .A(\SUBBYTES[5].a/w2123 ), .B(
        \SUBBYTES[5].a/w2124 ), .Z(n11144) );
  XOR \SUBBYTES[5].a/U5399  ( .A(\SUBBYTES[5].a/w2108 ), .B(
        \SUBBYTES[5].a/w2111 ), .Z(n11145) );
  XOR \SUBBYTES[5].a/U5397  ( .A(n12055), .B(n11148), .Z(n11146) );
  XOR \SUBBYTES[5].a/U5396  ( .A(n12057), .B(n12056), .Z(n11147) );
  XOR \SUBBYTES[5].a/U5395  ( .A(\SUBBYTES[5].a/w2116 ), .B(
        \SUBBYTES[5].a/w2143 ), .Z(n11148) );
  XOR \SUBBYTES[5].a/U5393  ( .A(n12058), .B(n11151), .Z(n11149) );
  XOR \SUBBYTES[5].a/U5392  ( .A(\SUBBYTES[5].a/w2149 ), .B(
        \SUBBYTES[5].a/w2151 ), .Z(n11150) );
  XOR \SUBBYTES[5].a/U5391  ( .A(\SUBBYTES[5].a/w2109 ), .B(
        \SUBBYTES[5].a/w2141 ), .Z(n11151) );
  XOR \SUBBYTES[5].a/U5390  ( .A(\SUBBYTES[5].a/w1941 ), .B(
        \SUBBYTES[5].a/w1942 ), .Z(n12060) );
  XOR \SUBBYTES[5].a/U5389  ( .A(n12060), .B(n11152), .Z(n12059) );
  XOR \SUBBYTES[5].a/U5388  ( .A(\SUBBYTES[5].a/w1934 ), .B(
        \SUBBYTES[5].a/w1951 ), .Z(n11152) );
  XOR \SUBBYTES[5].a/U5386  ( .A(\SUBBYTES[5].a/w1933 ), .B(
        \SUBBYTES[5].a/w1948 ), .Z(n11153) );
  XOR \SUBBYTES[5].a/U5385  ( .A(n12060), .B(n11154), .Z(n12223) );
  XOR \SUBBYTES[5].a/U5384  ( .A(\SUBBYTES[5].a/w1948 ), .B(
        \SUBBYTES[5].a/w1949 ), .Z(n11154) );
  XOR \SUBBYTES[5].a/U5383  ( .A(\SUBBYTES[5].a/w1910 ), .B(n11155), .Z(n12062) );
  XOR \SUBBYTES[5].a/U5382  ( .A(\SUBBYTES[5].a/w1901 ), .B(
        \SUBBYTES[5].a/w1902 ), .Z(n11155) );
  XOR \SUBBYTES[5].a/U5380  ( .A(\SUBBYTES[5].a/w1912 ), .B(n12223), .Z(n11156) );
  XOR \SUBBYTES[5].a/U5379  ( .A(n11158), .B(n11157), .Z(n12063) );
  XOR \SUBBYTES[5].a/U5378  ( .A(n11160), .B(n11159), .Z(n11157) );
  XOR \SUBBYTES[5].a/U5377  ( .A(\SUBBYTES[5].a/w1948 ), .B(
        \SUBBYTES[5].a/w1949 ), .Z(n11158) );
  XOR \SUBBYTES[5].a/U5376  ( .A(\SUBBYTES[5].a/w1912 ), .B(
        \SUBBYTES[5].a/w1936 ), .Z(n11159) );
  XOR \SUBBYTES[5].a/U5375  ( .A(\SUBBYTES[5].a/w1901 ), .B(
        \SUBBYTES[5].a/w1910 ), .Z(n11160) );
  XOR \SUBBYTES[5].a/U5374  ( .A(\SUBBYTES[5].a/w1933 ), .B(n11161), .Z(n12061) );
  XOR \SUBBYTES[5].a/U5373  ( .A(\SUBBYTES[5].a/w1916 ), .B(
        \SUBBYTES[5].a/w1919 ), .Z(n11161) );
  XOR \SUBBYTES[5].a/U5371  ( .A(\SUBBYTES[5].a/w1904 ), .B(n12063), .Z(n11162) );
  XOR \SUBBYTES[5].a/U5369  ( .A(\SUBBYTES[5].a/w1936 ), .B(
        \SUBBYTES[5].a/w1949 ), .Z(n11163) );
  XOR \SUBBYTES[5].a/U5367  ( .A(n11167), .B(n11166), .Z(n11164) );
  XOR \SUBBYTES[5].a/U5366  ( .A(n11169), .B(n11168), .Z(n11165) );
  XOR \SUBBYTES[5].a/U5365  ( .A(\SUBBYTES[5].a/w1948 ), .B(
        \SUBBYTES[5].a/w1951 ), .Z(n11166) );
  XOR \SUBBYTES[5].a/U5364  ( .A(\SUBBYTES[5].a/w1941 ), .B(
        \SUBBYTES[5].a/w1944 ), .Z(n11167) );
  XOR \SUBBYTES[5].a/U5363  ( .A(\SUBBYTES[5].a/w1916 ), .B(
        \SUBBYTES[5].a/w1917 ), .Z(n11168) );
  XOR \SUBBYTES[5].a/U5362  ( .A(\SUBBYTES[5].a/w1901 ), .B(
        \SUBBYTES[5].a/w1904 ), .Z(n11169) );
  XOR \SUBBYTES[5].a/U5360  ( .A(n12060), .B(n11172), .Z(n11170) );
  XOR \SUBBYTES[5].a/U5359  ( .A(n12062), .B(n12061), .Z(n11171) );
  XOR \SUBBYTES[5].a/U5358  ( .A(\SUBBYTES[5].a/w1909 ), .B(
        \SUBBYTES[5].a/w1936 ), .Z(n11172) );
  XOR \SUBBYTES[5].a/U5356  ( .A(n12063), .B(n11175), .Z(n11173) );
  XOR \SUBBYTES[5].a/U5355  ( .A(\SUBBYTES[5].a/w1942 ), .B(
        \SUBBYTES[5].a/w1944 ), .Z(n11174) );
  XOR \SUBBYTES[5].a/U5354  ( .A(\SUBBYTES[5].a/w1902 ), .B(
        \SUBBYTES[5].a/w1934 ), .Z(n11175) );
  XOR \SUBBYTES[5].a/U5353  ( .A(\SUBBYTES[5].a/w1734 ), .B(
        \SUBBYTES[5].a/w1735 ), .Z(n12065) );
  XOR \SUBBYTES[5].a/U5352  ( .A(n12065), .B(n11176), .Z(n12064) );
  XOR \SUBBYTES[5].a/U5351  ( .A(\SUBBYTES[5].a/w1727 ), .B(
        \SUBBYTES[5].a/w1744 ), .Z(n11176) );
  XOR \SUBBYTES[5].a/U5349  ( .A(\SUBBYTES[5].a/w1726 ), .B(
        \SUBBYTES[5].a/w1741 ), .Z(n11177) );
  XOR \SUBBYTES[5].a/U5348  ( .A(n12065), .B(n11178), .Z(n12224) );
  XOR \SUBBYTES[5].a/U5347  ( .A(\SUBBYTES[5].a/w1741 ), .B(
        \SUBBYTES[5].a/w1742 ), .Z(n11178) );
  XOR \SUBBYTES[5].a/U5346  ( .A(\SUBBYTES[5].a/w1703 ), .B(n11179), .Z(n12067) );
  XOR \SUBBYTES[5].a/U5345  ( .A(\SUBBYTES[5].a/w1694 ), .B(
        \SUBBYTES[5].a/w1695 ), .Z(n11179) );
  XOR \SUBBYTES[5].a/U5343  ( .A(\SUBBYTES[5].a/w1705 ), .B(n12224), .Z(n11180) );
  XOR \SUBBYTES[5].a/U5342  ( .A(n11182), .B(n11181), .Z(n12068) );
  XOR \SUBBYTES[5].a/U5341  ( .A(n11184), .B(n11183), .Z(n11181) );
  XOR \SUBBYTES[5].a/U5340  ( .A(\SUBBYTES[5].a/w1741 ), .B(
        \SUBBYTES[5].a/w1742 ), .Z(n11182) );
  XOR \SUBBYTES[5].a/U5339  ( .A(\SUBBYTES[5].a/w1705 ), .B(
        \SUBBYTES[5].a/w1729 ), .Z(n11183) );
  XOR \SUBBYTES[5].a/U5338  ( .A(\SUBBYTES[5].a/w1694 ), .B(
        \SUBBYTES[5].a/w1703 ), .Z(n11184) );
  XOR \SUBBYTES[5].a/U5337  ( .A(\SUBBYTES[5].a/w1726 ), .B(n11185), .Z(n12066) );
  XOR \SUBBYTES[5].a/U5336  ( .A(\SUBBYTES[5].a/w1709 ), .B(
        \SUBBYTES[5].a/w1712 ), .Z(n11185) );
  XOR \SUBBYTES[5].a/U5334  ( .A(\SUBBYTES[5].a/w1697 ), .B(n12068), .Z(n11186) );
  XOR \SUBBYTES[5].a/U5332  ( .A(\SUBBYTES[5].a/w1729 ), .B(
        \SUBBYTES[5].a/w1742 ), .Z(n11187) );
  XOR \SUBBYTES[5].a/U5330  ( .A(n11191), .B(n11190), .Z(n11188) );
  XOR \SUBBYTES[5].a/U5329  ( .A(n11193), .B(n11192), .Z(n11189) );
  XOR \SUBBYTES[5].a/U5328  ( .A(\SUBBYTES[5].a/w1741 ), .B(
        \SUBBYTES[5].a/w1744 ), .Z(n11190) );
  XOR \SUBBYTES[5].a/U5327  ( .A(\SUBBYTES[5].a/w1734 ), .B(
        \SUBBYTES[5].a/w1737 ), .Z(n11191) );
  XOR \SUBBYTES[5].a/U5326  ( .A(\SUBBYTES[5].a/w1709 ), .B(
        \SUBBYTES[5].a/w1710 ), .Z(n11192) );
  XOR \SUBBYTES[5].a/U5325  ( .A(\SUBBYTES[5].a/w1694 ), .B(
        \SUBBYTES[5].a/w1697 ), .Z(n11193) );
  XOR \SUBBYTES[5].a/U5323  ( .A(n12065), .B(n11196), .Z(n11194) );
  XOR \SUBBYTES[5].a/U5322  ( .A(n12067), .B(n12066), .Z(n11195) );
  XOR \SUBBYTES[5].a/U5321  ( .A(\SUBBYTES[5].a/w1702 ), .B(
        \SUBBYTES[5].a/w1729 ), .Z(n11196) );
  XOR \SUBBYTES[5].a/U5319  ( .A(n12068), .B(n11199), .Z(n11197) );
  XOR \SUBBYTES[5].a/U5318  ( .A(\SUBBYTES[5].a/w1735 ), .B(
        \SUBBYTES[5].a/w1737 ), .Z(n11198) );
  XOR \SUBBYTES[5].a/U5317  ( .A(\SUBBYTES[5].a/w1695 ), .B(
        \SUBBYTES[5].a/w1727 ), .Z(n11199) );
  XOR \SUBBYTES[5].a/U5316  ( .A(\SUBBYTES[5].a/w1527 ), .B(
        \SUBBYTES[5].a/w1528 ), .Z(n12070) );
  XOR \SUBBYTES[5].a/U5315  ( .A(n12070), .B(n11200), .Z(n12069) );
  XOR \SUBBYTES[5].a/U5314  ( .A(\SUBBYTES[5].a/w1520 ), .B(
        \SUBBYTES[5].a/w1537 ), .Z(n11200) );
  XOR \SUBBYTES[5].a/U5312  ( .A(\SUBBYTES[5].a/w1519 ), .B(
        \SUBBYTES[5].a/w1534 ), .Z(n11201) );
  XOR \SUBBYTES[5].a/U5311  ( .A(n12070), .B(n11202), .Z(n12225) );
  XOR \SUBBYTES[5].a/U5310  ( .A(\SUBBYTES[5].a/w1534 ), .B(
        \SUBBYTES[5].a/w1535 ), .Z(n11202) );
  XOR \SUBBYTES[5].a/U5309  ( .A(\SUBBYTES[5].a/w1496 ), .B(n11203), .Z(n12072) );
  XOR \SUBBYTES[5].a/U5308  ( .A(\SUBBYTES[5].a/w1487 ), .B(
        \SUBBYTES[5].a/w1488 ), .Z(n11203) );
  XOR \SUBBYTES[5].a/U5306  ( .A(\SUBBYTES[5].a/w1498 ), .B(n12225), .Z(n11204) );
  XOR \SUBBYTES[5].a/U5305  ( .A(n11206), .B(n11205), .Z(n12073) );
  XOR \SUBBYTES[5].a/U5304  ( .A(n11208), .B(n11207), .Z(n11205) );
  XOR \SUBBYTES[5].a/U5303  ( .A(\SUBBYTES[5].a/w1534 ), .B(
        \SUBBYTES[5].a/w1535 ), .Z(n11206) );
  XOR \SUBBYTES[5].a/U5302  ( .A(\SUBBYTES[5].a/w1498 ), .B(
        \SUBBYTES[5].a/w1522 ), .Z(n11207) );
  XOR \SUBBYTES[5].a/U5301  ( .A(\SUBBYTES[5].a/w1487 ), .B(
        \SUBBYTES[5].a/w1496 ), .Z(n11208) );
  XOR \SUBBYTES[5].a/U5300  ( .A(\SUBBYTES[5].a/w1519 ), .B(n11209), .Z(n12071) );
  XOR \SUBBYTES[5].a/U5299  ( .A(\SUBBYTES[5].a/w1502 ), .B(
        \SUBBYTES[5].a/w1505 ), .Z(n11209) );
  XOR \SUBBYTES[5].a/U5297  ( .A(\SUBBYTES[5].a/w1490 ), .B(n12073), .Z(n11210) );
  XOR \SUBBYTES[5].a/U5295  ( .A(\SUBBYTES[5].a/w1522 ), .B(
        \SUBBYTES[5].a/w1535 ), .Z(n11211) );
  XOR \SUBBYTES[5].a/U5293  ( .A(n11215), .B(n11214), .Z(n11212) );
  XOR \SUBBYTES[5].a/U5292  ( .A(n11217), .B(n11216), .Z(n11213) );
  XOR \SUBBYTES[5].a/U5291  ( .A(\SUBBYTES[5].a/w1534 ), .B(
        \SUBBYTES[5].a/w1537 ), .Z(n11214) );
  XOR \SUBBYTES[5].a/U5290  ( .A(\SUBBYTES[5].a/w1527 ), .B(
        \SUBBYTES[5].a/w1530 ), .Z(n11215) );
  XOR \SUBBYTES[5].a/U5289  ( .A(\SUBBYTES[5].a/w1502 ), .B(
        \SUBBYTES[5].a/w1503 ), .Z(n11216) );
  XOR \SUBBYTES[5].a/U5288  ( .A(\SUBBYTES[5].a/w1487 ), .B(
        \SUBBYTES[5].a/w1490 ), .Z(n11217) );
  XOR \SUBBYTES[5].a/U5286  ( .A(n12070), .B(n11220), .Z(n11218) );
  XOR \SUBBYTES[5].a/U5285  ( .A(n12072), .B(n12071), .Z(n11219) );
  XOR \SUBBYTES[5].a/U5284  ( .A(\SUBBYTES[5].a/w1495 ), .B(
        \SUBBYTES[5].a/w1522 ), .Z(n11220) );
  XOR \SUBBYTES[5].a/U5282  ( .A(n12073), .B(n11223), .Z(n11221) );
  XOR \SUBBYTES[5].a/U5281  ( .A(\SUBBYTES[5].a/w1528 ), .B(
        \SUBBYTES[5].a/w1530 ), .Z(n11222) );
  XOR \SUBBYTES[5].a/U5280  ( .A(\SUBBYTES[5].a/w1488 ), .B(
        \SUBBYTES[5].a/w1520 ), .Z(n11223) );
  XOR \SUBBYTES[5].a/U5279  ( .A(\SUBBYTES[5].a/w1320 ), .B(
        \SUBBYTES[5].a/w1321 ), .Z(n12075) );
  XOR \SUBBYTES[5].a/U5278  ( .A(n12075), .B(n11224), .Z(n12074) );
  XOR \SUBBYTES[5].a/U5277  ( .A(\SUBBYTES[5].a/w1313 ), .B(
        \SUBBYTES[5].a/w1330 ), .Z(n11224) );
  XOR \SUBBYTES[5].a/U5275  ( .A(\SUBBYTES[5].a/w1312 ), .B(
        \SUBBYTES[5].a/w1327 ), .Z(n11225) );
  XOR \SUBBYTES[5].a/U5274  ( .A(n12075), .B(n11226), .Z(n12226) );
  XOR \SUBBYTES[5].a/U5273  ( .A(\SUBBYTES[5].a/w1327 ), .B(
        \SUBBYTES[5].a/w1328 ), .Z(n11226) );
  XOR \SUBBYTES[5].a/U5272  ( .A(\SUBBYTES[5].a/w1289 ), .B(n11227), .Z(n12077) );
  XOR \SUBBYTES[5].a/U5271  ( .A(\SUBBYTES[5].a/w1280 ), .B(
        \SUBBYTES[5].a/w1281 ), .Z(n11227) );
  XOR \SUBBYTES[5].a/U5269  ( .A(\SUBBYTES[5].a/w1291 ), .B(n12226), .Z(n11228) );
  XOR \SUBBYTES[5].a/U5268  ( .A(n11230), .B(n11229), .Z(n12078) );
  XOR \SUBBYTES[5].a/U5267  ( .A(n11232), .B(n11231), .Z(n11229) );
  XOR \SUBBYTES[5].a/U5266  ( .A(\SUBBYTES[5].a/w1327 ), .B(
        \SUBBYTES[5].a/w1328 ), .Z(n11230) );
  XOR \SUBBYTES[5].a/U5265  ( .A(\SUBBYTES[5].a/w1291 ), .B(
        \SUBBYTES[5].a/w1315 ), .Z(n11231) );
  XOR \SUBBYTES[5].a/U5264  ( .A(\SUBBYTES[5].a/w1280 ), .B(
        \SUBBYTES[5].a/w1289 ), .Z(n11232) );
  XOR \SUBBYTES[5].a/U5263  ( .A(\SUBBYTES[5].a/w1312 ), .B(n11233), .Z(n12076) );
  XOR \SUBBYTES[5].a/U5262  ( .A(\SUBBYTES[5].a/w1295 ), .B(
        \SUBBYTES[5].a/w1298 ), .Z(n11233) );
  XOR \SUBBYTES[5].a/U5260  ( .A(\SUBBYTES[5].a/w1283 ), .B(n12078), .Z(n11234) );
  XOR \SUBBYTES[5].a/U5258  ( .A(\SUBBYTES[5].a/w1315 ), .B(
        \SUBBYTES[5].a/w1328 ), .Z(n11235) );
  XOR \SUBBYTES[5].a/U5256  ( .A(n11239), .B(n11238), .Z(n11236) );
  XOR \SUBBYTES[5].a/U5255  ( .A(n11241), .B(n11240), .Z(n11237) );
  XOR \SUBBYTES[5].a/U5254  ( .A(\SUBBYTES[5].a/w1327 ), .B(
        \SUBBYTES[5].a/w1330 ), .Z(n11238) );
  XOR \SUBBYTES[5].a/U5253  ( .A(\SUBBYTES[5].a/w1320 ), .B(
        \SUBBYTES[5].a/w1323 ), .Z(n11239) );
  XOR \SUBBYTES[5].a/U5252  ( .A(\SUBBYTES[5].a/w1295 ), .B(
        \SUBBYTES[5].a/w1296 ), .Z(n11240) );
  XOR \SUBBYTES[5].a/U5251  ( .A(\SUBBYTES[5].a/w1280 ), .B(
        \SUBBYTES[5].a/w1283 ), .Z(n11241) );
  XOR \SUBBYTES[5].a/U5249  ( .A(n12075), .B(n11244), .Z(n11242) );
  XOR \SUBBYTES[5].a/U5248  ( .A(n12077), .B(n12076), .Z(n11243) );
  XOR \SUBBYTES[5].a/U5247  ( .A(\SUBBYTES[5].a/w1288 ), .B(
        \SUBBYTES[5].a/w1315 ), .Z(n11244) );
  XOR \SUBBYTES[5].a/U5245  ( .A(n12078), .B(n11247), .Z(n11245) );
  XOR \SUBBYTES[5].a/U5244  ( .A(\SUBBYTES[5].a/w1321 ), .B(
        \SUBBYTES[5].a/w1323 ), .Z(n11246) );
  XOR \SUBBYTES[5].a/U5243  ( .A(\SUBBYTES[5].a/w1281 ), .B(
        \SUBBYTES[5].a/w1313 ), .Z(n11247) );
  XOR \SUBBYTES[5].a/U5242  ( .A(\SUBBYTES[5].a/w1113 ), .B(
        \SUBBYTES[5].a/w1114 ), .Z(n12080) );
  XOR \SUBBYTES[5].a/U5241  ( .A(n12080), .B(n11248), .Z(n12079) );
  XOR \SUBBYTES[5].a/U5240  ( .A(\SUBBYTES[5].a/w1106 ), .B(
        \SUBBYTES[5].a/w1123 ), .Z(n11248) );
  XOR \SUBBYTES[5].a/U5238  ( .A(\SUBBYTES[5].a/w1105 ), .B(
        \SUBBYTES[5].a/w1120 ), .Z(n11249) );
  XOR \SUBBYTES[5].a/U5237  ( .A(n12080), .B(n11250), .Z(n12227) );
  XOR \SUBBYTES[5].a/U5236  ( .A(\SUBBYTES[5].a/w1120 ), .B(
        \SUBBYTES[5].a/w1121 ), .Z(n11250) );
  XOR \SUBBYTES[5].a/U5235  ( .A(\SUBBYTES[5].a/w1082 ), .B(n11251), .Z(n12082) );
  XOR \SUBBYTES[5].a/U5234  ( .A(\SUBBYTES[5].a/w1073 ), .B(
        \SUBBYTES[5].a/w1074 ), .Z(n11251) );
  XOR \SUBBYTES[5].a/U5232  ( .A(\SUBBYTES[5].a/w1084 ), .B(n12227), .Z(n11252) );
  XOR \SUBBYTES[5].a/U5231  ( .A(n11254), .B(n11253), .Z(n12083) );
  XOR \SUBBYTES[5].a/U5230  ( .A(n11256), .B(n11255), .Z(n11253) );
  XOR \SUBBYTES[5].a/U5229  ( .A(\SUBBYTES[5].a/w1120 ), .B(
        \SUBBYTES[5].a/w1121 ), .Z(n11254) );
  XOR \SUBBYTES[5].a/U5228  ( .A(\SUBBYTES[5].a/w1084 ), .B(
        \SUBBYTES[5].a/w1108 ), .Z(n11255) );
  XOR \SUBBYTES[5].a/U5227  ( .A(\SUBBYTES[5].a/w1073 ), .B(
        \SUBBYTES[5].a/w1082 ), .Z(n11256) );
  XOR \SUBBYTES[5].a/U5226  ( .A(\SUBBYTES[5].a/w1105 ), .B(n11257), .Z(n12081) );
  XOR \SUBBYTES[5].a/U5225  ( .A(\SUBBYTES[5].a/w1088 ), .B(
        \SUBBYTES[5].a/w1091 ), .Z(n11257) );
  XOR \SUBBYTES[5].a/U5223  ( .A(\SUBBYTES[5].a/w1076 ), .B(n12083), .Z(n11258) );
  XOR \SUBBYTES[5].a/U5221  ( .A(\SUBBYTES[5].a/w1108 ), .B(
        \SUBBYTES[5].a/w1121 ), .Z(n11259) );
  XOR \SUBBYTES[5].a/U5219  ( .A(n11263), .B(n11262), .Z(n11260) );
  XOR \SUBBYTES[5].a/U5218  ( .A(n11265), .B(n11264), .Z(n11261) );
  XOR \SUBBYTES[5].a/U5217  ( .A(\SUBBYTES[5].a/w1120 ), .B(
        \SUBBYTES[5].a/w1123 ), .Z(n11262) );
  XOR \SUBBYTES[5].a/U5216  ( .A(\SUBBYTES[5].a/w1113 ), .B(
        \SUBBYTES[5].a/w1116 ), .Z(n11263) );
  XOR \SUBBYTES[5].a/U5215  ( .A(\SUBBYTES[5].a/w1088 ), .B(
        \SUBBYTES[5].a/w1089 ), .Z(n11264) );
  XOR \SUBBYTES[5].a/U5214  ( .A(\SUBBYTES[5].a/w1073 ), .B(
        \SUBBYTES[5].a/w1076 ), .Z(n11265) );
  XOR \SUBBYTES[5].a/U5212  ( .A(n12080), .B(n11268), .Z(n11266) );
  XOR \SUBBYTES[5].a/U5211  ( .A(n12082), .B(n12081), .Z(n11267) );
  XOR \SUBBYTES[5].a/U5210  ( .A(\SUBBYTES[5].a/w1081 ), .B(
        \SUBBYTES[5].a/w1108 ), .Z(n11268) );
  XOR \SUBBYTES[5].a/U5208  ( .A(n12083), .B(n11271), .Z(n11269) );
  XOR \SUBBYTES[5].a/U5207  ( .A(\SUBBYTES[5].a/w1114 ), .B(
        \SUBBYTES[5].a/w1116 ), .Z(n11270) );
  XOR \SUBBYTES[5].a/U5206  ( .A(\SUBBYTES[5].a/w1074 ), .B(
        \SUBBYTES[5].a/w1106 ), .Z(n11271) );
  XOR \SUBBYTES[5].a/U5205  ( .A(\SUBBYTES[5].a/w906 ), .B(
        \SUBBYTES[5].a/w907 ), .Z(n12085) );
  XOR \SUBBYTES[5].a/U5204  ( .A(n12085), .B(n11272), .Z(n12084) );
  XOR \SUBBYTES[5].a/U5203  ( .A(\SUBBYTES[5].a/w899 ), .B(
        \SUBBYTES[5].a/w916 ), .Z(n11272) );
  XOR \SUBBYTES[5].a/U5201  ( .A(\SUBBYTES[5].a/w898 ), .B(
        \SUBBYTES[5].a/w913 ), .Z(n11273) );
  XOR \SUBBYTES[5].a/U5200  ( .A(n12085), .B(n11274), .Z(n12228) );
  XOR \SUBBYTES[5].a/U5199  ( .A(\SUBBYTES[5].a/w913 ), .B(
        \SUBBYTES[5].a/w914 ), .Z(n11274) );
  XOR \SUBBYTES[5].a/U5198  ( .A(\SUBBYTES[5].a/w875 ), .B(n11275), .Z(n12087)
         );
  XOR \SUBBYTES[5].a/U5197  ( .A(\SUBBYTES[5].a/w866 ), .B(
        \SUBBYTES[5].a/w867 ), .Z(n11275) );
  XOR \SUBBYTES[5].a/U5195  ( .A(\SUBBYTES[5].a/w877 ), .B(n12228), .Z(n11276)
         );
  XOR \SUBBYTES[5].a/U5194  ( .A(n11278), .B(n11277), .Z(n12088) );
  XOR \SUBBYTES[5].a/U5193  ( .A(n11280), .B(n11279), .Z(n11277) );
  XOR \SUBBYTES[5].a/U5192  ( .A(\SUBBYTES[5].a/w913 ), .B(
        \SUBBYTES[5].a/w914 ), .Z(n11278) );
  XOR \SUBBYTES[5].a/U5191  ( .A(\SUBBYTES[5].a/w877 ), .B(
        \SUBBYTES[5].a/w901 ), .Z(n11279) );
  XOR \SUBBYTES[5].a/U5190  ( .A(\SUBBYTES[5].a/w866 ), .B(
        \SUBBYTES[5].a/w875 ), .Z(n11280) );
  XOR \SUBBYTES[5].a/U5189  ( .A(\SUBBYTES[5].a/w898 ), .B(n11281), .Z(n12086)
         );
  XOR \SUBBYTES[5].a/U5188  ( .A(\SUBBYTES[5].a/w881 ), .B(
        \SUBBYTES[5].a/w884 ), .Z(n11281) );
  XOR \SUBBYTES[5].a/U5186  ( .A(\SUBBYTES[5].a/w869 ), .B(n12088), .Z(n11282)
         );
  XOR \SUBBYTES[5].a/U5184  ( .A(\SUBBYTES[5].a/w901 ), .B(
        \SUBBYTES[5].a/w914 ), .Z(n11283) );
  XOR \SUBBYTES[5].a/U5182  ( .A(n11287), .B(n11286), .Z(n11284) );
  XOR \SUBBYTES[5].a/U5181  ( .A(n11289), .B(n11288), .Z(n11285) );
  XOR \SUBBYTES[5].a/U5180  ( .A(\SUBBYTES[5].a/w913 ), .B(
        \SUBBYTES[5].a/w916 ), .Z(n11286) );
  XOR \SUBBYTES[5].a/U5179  ( .A(\SUBBYTES[5].a/w906 ), .B(
        \SUBBYTES[5].a/w909 ), .Z(n11287) );
  XOR \SUBBYTES[5].a/U5178  ( .A(\SUBBYTES[5].a/w881 ), .B(
        \SUBBYTES[5].a/w882 ), .Z(n11288) );
  XOR \SUBBYTES[5].a/U5177  ( .A(\SUBBYTES[5].a/w866 ), .B(
        \SUBBYTES[5].a/w869 ), .Z(n11289) );
  XOR \SUBBYTES[5].a/U5175  ( .A(n12085), .B(n11292), .Z(n11290) );
  XOR \SUBBYTES[5].a/U5174  ( .A(n12087), .B(n12086), .Z(n11291) );
  XOR \SUBBYTES[5].a/U5173  ( .A(\SUBBYTES[5].a/w874 ), .B(
        \SUBBYTES[5].a/w901 ), .Z(n11292) );
  XOR \SUBBYTES[5].a/U5171  ( .A(n12088), .B(n11295), .Z(n11293) );
  XOR \SUBBYTES[5].a/U5170  ( .A(\SUBBYTES[5].a/w907 ), .B(
        \SUBBYTES[5].a/w909 ), .Z(n11294) );
  XOR \SUBBYTES[5].a/U5169  ( .A(\SUBBYTES[5].a/w867 ), .B(
        \SUBBYTES[5].a/w899 ), .Z(n11295) );
  XOR \SUBBYTES[5].a/U5168  ( .A(\SUBBYTES[5].a/w699 ), .B(
        \SUBBYTES[5].a/w700 ), .Z(n12090) );
  XOR \SUBBYTES[5].a/U5167  ( .A(n12090), .B(n11296), .Z(n12089) );
  XOR \SUBBYTES[5].a/U5166  ( .A(\SUBBYTES[5].a/w692 ), .B(
        \SUBBYTES[5].a/w709 ), .Z(n11296) );
  XOR \SUBBYTES[5].a/U5164  ( .A(\SUBBYTES[5].a/w691 ), .B(
        \SUBBYTES[5].a/w706 ), .Z(n11297) );
  XOR \SUBBYTES[5].a/U5163  ( .A(n12090), .B(n11298), .Z(n12229) );
  XOR \SUBBYTES[5].a/U5162  ( .A(\SUBBYTES[5].a/w706 ), .B(
        \SUBBYTES[5].a/w707 ), .Z(n11298) );
  XOR \SUBBYTES[5].a/U5161  ( .A(\SUBBYTES[5].a/w668 ), .B(n11299), .Z(n12092)
         );
  XOR \SUBBYTES[5].a/U5160  ( .A(\SUBBYTES[5].a/w659 ), .B(
        \SUBBYTES[5].a/w660 ), .Z(n11299) );
  XOR \SUBBYTES[5].a/U5158  ( .A(\SUBBYTES[5].a/w670 ), .B(n12229), .Z(n11300)
         );
  XOR \SUBBYTES[5].a/U5157  ( .A(n11302), .B(n11301), .Z(n12093) );
  XOR \SUBBYTES[5].a/U5156  ( .A(n11304), .B(n11303), .Z(n11301) );
  XOR \SUBBYTES[5].a/U5155  ( .A(\SUBBYTES[5].a/w706 ), .B(
        \SUBBYTES[5].a/w707 ), .Z(n11302) );
  XOR \SUBBYTES[5].a/U5154  ( .A(\SUBBYTES[5].a/w670 ), .B(
        \SUBBYTES[5].a/w694 ), .Z(n11303) );
  XOR \SUBBYTES[5].a/U5153  ( .A(\SUBBYTES[5].a/w659 ), .B(
        \SUBBYTES[5].a/w668 ), .Z(n11304) );
  XOR \SUBBYTES[5].a/U5152  ( .A(\SUBBYTES[5].a/w691 ), .B(n11305), .Z(n12091)
         );
  XOR \SUBBYTES[5].a/U5151  ( .A(\SUBBYTES[5].a/w674 ), .B(
        \SUBBYTES[5].a/w677 ), .Z(n11305) );
  XOR \SUBBYTES[5].a/U5149  ( .A(\SUBBYTES[5].a/w662 ), .B(n12093), .Z(n11306)
         );
  XOR \SUBBYTES[5].a/U5147  ( .A(\SUBBYTES[5].a/w694 ), .B(
        \SUBBYTES[5].a/w707 ), .Z(n11307) );
  XOR \SUBBYTES[5].a/U5145  ( .A(n11311), .B(n11310), .Z(n11308) );
  XOR \SUBBYTES[5].a/U5144  ( .A(n11313), .B(n11312), .Z(n11309) );
  XOR \SUBBYTES[5].a/U5143  ( .A(\SUBBYTES[5].a/w706 ), .B(
        \SUBBYTES[5].a/w709 ), .Z(n11310) );
  XOR \SUBBYTES[5].a/U5142  ( .A(\SUBBYTES[5].a/w699 ), .B(
        \SUBBYTES[5].a/w702 ), .Z(n11311) );
  XOR \SUBBYTES[5].a/U5141  ( .A(\SUBBYTES[5].a/w674 ), .B(
        \SUBBYTES[5].a/w675 ), .Z(n11312) );
  XOR \SUBBYTES[5].a/U5140  ( .A(\SUBBYTES[5].a/w659 ), .B(
        \SUBBYTES[5].a/w662 ), .Z(n11313) );
  XOR \SUBBYTES[5].a/U5138  ( .A(n12090), .B(n11316), .Z(n11314) );
  XOR \SUBBYTES[5].a/U5137  ( .A(n12092), .B(n12091), .Z(n11315) );
  XOR \SUBBYTES[5].a/U5136  ( .A(\SUBBYTES[5].a/w667 ), .B(
        \SUBBYTES[5].a/w694 ), .Z(n11316) );
  XOR \SUBBYTES[5].a/U5134  ( .A(n12093), .B(n11319), .Z(n11317) );
  XOR \SUBBYTES[5].a/U5133  ( .A(\SUBBYTES[5].a/w700 ), .B(
        \SUBBYTES[5].a/w702 ), .Z(n11318) );
  XOR \SUBBYTES[5].a/U5132  ( .A(\SUBBYTES[5].a/w660 ), .B(
        \SUBBYTES[5].a/w692 ), .Z(n11319) );
  XOR \SUBBYTES[5].a/U5131  ( .A(\SUBBYTES[5].a/w492 ), .B(
        \SUBBYTES[5].a/w493 ), .Z(n12095) );
  XOR \SUBBYTES[5].a/U5130  ( .A(n12095), .B(n11320), .Z(n12094) );
  XOR \SUBBYTES[5].a/U5129  ( .A(\SUBBYTES[5].a/w485 ), .B(
        \SUBBYTES[5].a/w502 ), .Z(n11320) );
  XOR \SUBBYTES[5].a/U5127  ( .A(\SUBBYTES[5].a/w484 ), .B(
        \SUBBYTES[5].a/w499 ), .Z(n11321) );
  XOR \SUBBYTES[5].a/U5126  ( .A(n12095), .B(n11322), .Z(n12230) );
  XOR \SUBBYTES[5].a/U5125  ( .A(\SUBBYTES[5].a/w499 ), .B(
        \SUBBYTES[5].a/w500 ), .Z(n11322) );
  XOR \SUBBYTES[5].a/U5124  ( .A(\SUBBYTES[5].a/w461 ), .B(n11323), .Z(n12097)
         );
  XOR \SUBBYTES[5].a/U5123  ( .A(\SUBBYTES[5].a/w452 ), .B(
        \SUBBYTES[5].a/w453 ), .Z(n11323) );
  XOR \SUBBYTES[5].a/U5121  ( .A(\SUBBYTES[5].a/w463 ), .B(n12230), .Z(n11324)
         );
  XOR \SUBBYTES[5].a/U5120  ( .A(n11326), .B(n11325), .Z(n12098) );
  XOR \SUBBYTES[5].a/U5119  ( .A(n11328), .B(n11327), .Z(n11325) );
  XOR \SUBBYTES[5].a/U5118  ( .A(\SUBBYTES[5].a/w499 ), .B(
        \SUBBYTES[5].a/w500 ), .Z(n11326) );
  XOR \SUBBYTES[5].a/U5117  ( .A(\SUBBYTES[5].a/w463 ), .B(
        \SUBBYTES[5].a/w487 ), .Z(n11327) );
  XOR \SUBBYTES[5].a/U5116  ( .A(\SUBBYTES[5].a/w452 ), .B(
        \SUBBYTES[5].a/w461 ), .Z(n11328) );
  XOR \SUBBYTES[5].a/U5115  ( .A(\SUBBYTES[5].a/w484 ), .B(n11329), .Z(n12096)
         );
  XOR \SUBBYTES[5].a/U5114  ( .A(\SUBBYTES[5].a/w467 ), .B(
        \SUBBYTES[5].a/w470 ), .Z(n11329) );
  XOR \SUBBYTES[5].a/U5112  ( .A(\SUBBYTES[5].a/w455 ), .B(n12098), .Z(n11330)
         );
  XOR \SUBBYTES[5].a/U5110  ( .A(\SUBBYTES[5].a/w487 ), .B(
        \SUBBYTES[5].a/w500 ), .Z(n11331) );
  XOR \SUBBYTES[5].a/U5108  ( .A(n11335), .B(n11334), .Z(n11332) );
  XOR \SUBBYTES[5].a/U5107  ( .A(n11337), .B(n11336), .Z(n11333) );
  XOR \SUBBYTES[5].a/U5106  ( .A(\SUBBYTES[5].a/w499 ), .B(
        \SUBBYTES[5].a/w502 ), .Z(n11334) );
  XOR \SUBBYTES[5].a/U5105  ( .A(\SUBBYTES[5].a/w492 ), .B(
        \SUBBYTES[5].a/w495 ), .Z(n11335) );
  XOR \SUBBYTES[5].a/U5104  ( .A(\SUBBYTES[5].a/w467 ), .B(
        \SUBBYTES[5].a/w468 ), .Z(n11336) );
  XOR \SUBBYTES[5].a/U5103  ( .A(\SUBBYTES[5].a/w452 ), .B(
        \SUBBYTES[5].a/w455 ), .Z(n11337) );
  XOR \SUBBYTES[5].a/U5101  ( .A(n12095), .B(n11340), .Z(n11338) );
  XOR \SUBBYTES[5].a/U5100  ( .A(n12097), .B(n12096), .Z(n11339) );
  XOR \SUBBYTES[5].a/U5099  ( .A(\SUBBYTES[5].a/w460 ), .B(
        \SUBBYTES[5].a/w487 ), .Z(n11340) );
  XOR \SUBBYTES[5].a/U5097  ( .A(n12098), .B(n11343), .Z(n11341) );
  XOR \SUBBYTES[5].a/U5096  ( .A(\SUBBYTES[5].a/w493 ), .B(
        \SUBBYTES[5].a/w495 ), .Z(n11342) );
  XOR \SUBBYTES[5].a/U5095  ( .A(\SUBBYTES[5].a/w453 ), .B(
        \SUBBYTES[5].a/w485 ), .Z(n11343) );
  XOR \SUBBYTES[5].a/U5094  ( .A(\SUBBYTES[5].a/w285 ), .B(
        \SUBBYTES[5].a/w286 ), .Z(n12100) );
  XOR \SUBBYTES[5].a/U5093  ( .A(n12100), .B(n11344), .Z(n12099) );
  XOR \SUBBYTES[5].a/U5092  ( .A(\SUBBYTES[5].a/w278 ), .B(
        \SUBBYTES[5].a/w295 ), .Z(n11344) );
  XOR \SUBBYTES[5].a/U5090  ( .A(\SUBBYTES[5].a/w277 ), .B(
        \SUBBYTES[5].a/w292 ), .Z(n11345) );
  XOR \SUBBYTES[5].a/U5089  ( .A(n12100), .B(n11346), .Z(n12231) );
  XOR \SUBBYTES[5].a/U5088  ( .A(\SUBBYTES[5].a/w292 ), .B(
        \SUBBYTES[5].a/w293 ), .Z(n11346) );
  XOR \SUBBYTES[5].a/U5087  ( .A(\SUBBYTES[5].a/w254 ), .B(n11347), .Z(n12102)
         );
  XOR \SUBBYTES[5].a/U5086  ( .A(\SUBBYTES[5].a/w245 ), .B(
        \SUBBYTES[5].a/w246 ), .Z(n11347) );
  XOR \SUBBYTES[5].a/U5084  ( .A(\SUBBYTES[5].a/w256 ), .B(n12231), .Z(n11348)
         );
  XOR \SUBBYTES[5].a/U5083  ( .A(n11350), .B(n11349), .Z(n12103) );
  XOR \SUBBYTES[5].a/U5082  ( .A(n11352), .B(n11351), .Z(n11349) );
  XOR \SUBBYTES[5].a/U5081  ( .A(\SUBBYTES[5].a/w292 ), .B(
        \SUBBYTES[5].a/w293 ), .Z(n11350) );
  XOR \SUBBYTES[5].a/U5080  ( .A(\SUBBYTES[5].a/w256 ), .B(
        \SUBBYTES[5].a/w280 ), .Z(n11351) );
  XOR \SUBBYTES[5].a/U5079  ( .A(\SUBBYTES[5].a/w245 ), .B(
        \SUBBYTES[5].a/w254 ), .Z(n11352) );
  XOR \SUBBYTES[5].a/U5078  ( .A(\SUBBYTES[5].a/w277 ), .B(n11353), .Z(n12101)
         );
  XOR \SUBBYTES[5].a/U5077  ( .A(\SUBBYTES[5].a/w260 ), .B(
        \SUBBYTES[5].a/w263 ), .Z(n11353) );
  XOR \SUBBYTES[5].a/U5075  ( .A(\SUBBYTES[5].a/w248 ), .B(n12103), .Z(n11354)
         );
  XOR \SUBBYTES[5].a/U5073  ( .A(\SUBBYTES[5].a/w280 ), .B(
        \SUBBYTES[5].a/w293 ), .Z(n11355) );
  XOR \SUBBYTES[5].a/U5071  ( .A(n11359), .B(n11358), .Z(n11356) );
  XOR \SUBBYTES[5].a/U5070  ( .A(n11361), .B(n11360), .Z(n11357) );
  XOR \SUBBYTES[5].a/U5069  ( .A(\SUBBYTES[5].a/w292 ), .B(
        \SUBBYTES[5].a/w295 ), .Z(n11358) );
  XOR \SUBBYTES[5].a/U5068  ( .A(\SUBBYTES[5].a/w285 ), .B(
        \SUBBYTES[5].a/w288 ), .Z(n11359) );
  XOR \SUBBYTES[5].a/U5067  ( .A(\SUBBYTES[5].a/w260 ), .B(
        \SUBBYTES[5].a/w261 ), .Z(n11360) );
  XOR \SUBBYTES[5].a/U5066  ( .A(\SUBBYTES[5].a/w245 ), .B(
        \SUBBYTES[5].a/w248 ), .Z(n11361) );
  XOR \SUBBYTES[5].a/U5064  ( .A(n12100), .B(n11364), .Z(n11362) );
  XOR \SUBBYTES[5].a/U5063  ( .A(n12102), .B(n12101), .Z(n11363) );
  XOR \SUBBYTES[5].a/U5062  ( .A(\SUBBYTES[5].a/w253 ), .B(
        \SUBBYTES[5].a/w280 ), .Z(n11364) );
  XOR \SUBBYTES[5].a/U5060  ( .A(n12103), .B(n11367), .Z(n11365) );
  XOR \SUBBYTES[5].a/U5059  ( .A(\SUBBYTES[5].a/w286 ), .B(
        \SUBBYTES[5].a/w288 ), .Z(n11366) );
  XOR \SUBBYTES[5].a/U5058  ( .A(\SUBBYTES[5].a/w246 ), .B(
        \SUBBYTES[5].a/w278 ), .Z(n11367) );
  XOR \SUBBYTES[5].a/U5057  ( .A(\w1[5][1] ), .B(n11368), .Z(n12104) );
  XOR \SUBBYTES[5].a/U5056  ( .A(\w1[5][3] ), .B(\w1[5][2] ), .Z(n11368) );
  XOR \SUBBYTES[5].a/U5055  ( .A(\w1[5][6] ), .B(n12104), .Z(
        \SUBBYTES[5].a/w3378 ) );
  XOR \SUBBYTES[5].a/U5054  ( .A(\w1[5][0] ), .B(\SUBBYTES[5].a/w3378 ), .Z(
        \SUBBYTES[5].a/w3265 ) );
  XOR \SUBBYTES[5].a/U5053  ( .A(\w1[5][0] ), .B(n11369), .Z(
        \SUBBYTES[5].a/w3266 ) );
  XOR \SUBBYTES[5].a/U5052  ( .A(\w1[5][6] ), .B(\w1[5][5] ), .Z(n11369) );
  XOR \SUBBYTES[5].a/U5051  ( .A(\w1[5][5] ), .B(n12104), .Z(
        \SUBBYTES[5].a/w3396 ) );
  XOR \SUBBYTES[5].a/U5050  ( .A(n11371), .B(n11370), .Z(\SUBBYTES[5].a/w3389 ) );
  XOR \SUBBYTES[5].a/U5049  ( .A(\w1[5][3] ), .B(\w1[5][1] ), .Z(n11370) );
  XOR \SUBBYTES[5].a/U5048  ( .A(\w1[5][7] ), .B(\w1[5][4] ), .Z(n11371) );
  XOR \SUBBYTES[5].a/U5047  ( .A(\w1[5][0] ), .B(\SUBBYTES[5].a/w3389 ), .Z(
        \SUBBYTES[5].a/w3268 ) );
  XOR \SUBBYTES[5].a/U5046  ( .A(n11373), .B(n11372), .Z(\SUBBYTES[5].a/w3376 ) );
  XOR \SUBBYTES[5].a/U5045  ( .A(\SUBBYTES[5].a/w3337 ), .B(n1036), .Z(n11372)
         );
  XOR \SUBBYTES[5].a/U5044  ( .A(\SUBBYTES[5].a/w3330 ), .B(
        \SUBBYTES[5].a/w3333 ), .Z(n11373) );
  XOR \SUBBYTES[5].a/U5043  ( .A(n11375), .B(n11374), .Z(\SUBBYTES[5].a/w3377 ) );
  XOR \SUBBYTES[5].a/U5042  ( .A(\SUBBYTES[5].a/w3337 ), .B(n10983), .Z(n11374) );
  XOR \SUBBYTES[5].a/U5041  ( .A(\SUBBYTES[5].a/w3330 ), .B(n10982), .Z(n11375) );
  XOR \SUBBYTES[5].a/U5040  ( .A(\SUBBYTES[5].a/w3389 ), .B(n11376), .Z(
        \SUBBYTES[5].a/w3379 ) );
  XOR \SUBBYTES[5].a/U5039  ( .A(\w1[5][6] ), .B(\w1[5][5] ), .Z(n11376) );
  XOR \SUBBYTES[5].a/U5038  ( .A(n11378), .B(n11377), .Z(\SUBBYTES[5].a/w3380 ) );
  XOR \SUBBYTES[5].a/U5037  ( .A(n10983), .B(n1036), .Z(n11377) );
  XOR \SUBBYTES[5].a/U5036  ( .A(n10982), .B(\SUBBYTES[5].a/w3333 ), .Z(n11378) );
  XOR \SUBBYTES[5].a/U5035  ( .A(\w1[5][7] ), .B(\w1[5][2] ), .Z(n12110) );
  XOR \SUBBYTES[5].a/U5034  ( .A(n12110), .B(n11379), .Z(\SUBBYTES[5].a/w3381 ) );
  XOR \SUBBYTES[5].a/U5033  ( .A(\w1[5][5] ), .B(\w1[5][4] ), .Z(n11379) );
  XOR \SUBBYTES[5].a/U5032  ( .A(\w1[5][7] ), .B(\SUBBYTES[5].a/w3266 ), .Z(
        \SUBBYTES[5].a/w3269 ) );
  XOR \SUBBYTES[5].a/U5031  ( .A(\w1[5][1] ), .B(\SUBBYTES[5].a/w3266 ), .Z(
        \SUBBYTES[5].a/w3270 ) );
  XOR \SUBBYTES[5].a/U5030  ( .A(\w1[5][4] ), .B(\SUBBYTES[5].a/w3266 ), .Z(
        \SUBBYTES[5].a/w3271 ) );
  XOR \SUBBYTES[5].a/U5029  ( .A(\SUBBYTES[5].a/w3270 ), .B(n12110), .Z(
        \SUBBYTES[5].a/w3272 ) );
  XOR \SUBBYTES[5].a/U5028  ( .A(n12110), .B(n11380), .Z(\SUBBYTES[5].a/w3357 ) );
  XOR \SUBBYTES[5].a/U5027  ( .A(\w1[5][4] ), .B(\w1[5][1] ), .Z(n11380) );
  XOR \SUBBYTES[5].a/U5026  ( .A(n11382), .B(n11381), .Z(n12107) );
  XOR \SUBBYTES[5].a/U5025  ( .A(\w1[5][4] ), .B(n11383), .Z(n11381) );
  XOR \SUBBYTES[5].a/U5024  ( .A(\SUBBYTES[5].a/w3322 ), .B(\w1[5][6] ), .Z(
        n11382) );
  XOR \SUBBYTES[5].a/U5023  ( .A(\SUBBYTES[5].a/w3296 ), .B(
        \SUBBYTES[5].a/w3303 ), .Z(n11383) );
  XOR \SUBBYTES[5].a/U5022  ( .A(n11385), .B(n11384), .Z(n12105) );
  XOR \SUBBYTES[5].a/U5021  ( .A(\w1[5][1] ), .B(n11386), .Z(n11384) );
  XOR \SUBBYTES[5].a/U5020  ( .A(\SUBBYTES[5].a/w3321 ), .B(\w1[5][5] ), .Z(
        n11385) );
  XOR \SUBBYTES[5].a/U5019  ( .A(\SUBBYTES[5].a/w3297 ), .B(
        \SUBBYTES[5].a/w3304 ), .Z(n11386) );
  XOR \SUBBYTES[5].a/U5018  ( .A(n12107), .B(n12105), .Z(\SUBBYTES[5].a/w3327 ) );
  XOR \SUBBYTES[5].a/U5017  ( .A(\w1[5][5] ), .B(n11387), .Z(n12108) );
  XOR \SUBBYTES[5].a/U5016  ( .A(\SUBBYTES[5].a/w3289 ), .B(
        \SUBBYTES[5].a/w3299 ), .Z(n11387) );
  XOR \SUBBYTES[5].a/U5015  ( .A(n11389), .B(n11388), .Z(\SUBBYTES[5].a/w3314 ) );
  XOR \SUBBYTES[5].a/U5014  ( .A(n12108), .B(n11390), .Z(n11388) );
  XOR \SUBBYTES[5].a/U5013  ( .A(\w1[5][4] ), .B(\SUBBYTES[5].a/w3378 ), .Z(
        n11389) );
  XOR \SUBBYTES[5].a/U5012  ( .A(\SUBBYTES[5].a/w3291 ), .B(
        \SUBBYTES[5].a/w3296 ), .Z(n11390) );
  XOR \SUBBYTES[5].a/U5011  ( .A(n11392), .B(n11391), .Z(n12106) );
  XOR \SUBBYTES[5].a/U5010  ( .A(\SUBBYTES[5].a/w3324 ), .B(\w1[5][7] ), .Z(
        n11391) );
  XOR \SUBBYTES[5].a/U5009  ( .A(\SUBBYTES[5].a/w3299 ), .B(
        \SUBBYTES[5].a/w3306 ), .Z(n11392) );
  XOR \SUBBYTES[5].a/U5008  ( .A(n12105), .B(n12106), .Z(\SUBBYTES[5].a/w3326 ) );
  XOR \SUBBYTES[5].a/U5007  ( .A(\w1[5][3] ), .B(n11393), .Z(n12109) );
  XOR \SUBBYTES[5].a/U5006  ( .A(\SUBBYTES[5].a/w3288 ), .B(
        \SUBBYTES[5].a/w3291 ), .Z(n11393) );
  XOR \SUBBYTES[5].a/U5005  ( .A(n11395), .B(n11394), .Z(\SUBBYTES[5].a/w3315 ) );
  XOR \SUBBYTES[5].a/U5004  ( .A(n12109), .B(n11396), .Z(n11394) );
  XOR \SUBBYTES[5].a/U5003  ( .A(\w1[5][6] ), .B(\SUBBYTES[5].a/w3357 ), .Z(
        n11395) );
  XOR \SUBBYTES[5].a/U5002  ( .A(\SUBBYTES[5].a/w3296 ), .B(
        \SUBBYTES[5].a/w3297 ), .Z(n11396) );
  XOR \SUBBYTES[5].a/U5001  ( .A(n12107), .B(n12106), .Z(\SUBBYTES[5].a/w3335 ) );
  XOR \SUBBYTES[5].a/U5000  ( .A(n11398), .B(n11397), .Z(\SUBBYTES[5].a/w3336 ) );
  XOR \SUBBYTES[5].a/U4999  ( .A(\w1[5][7] ), .B(n12108), .Z(n11397) );
  XOR \SUBBYTES[5].a/U4998  ( .A(\SUBBYTES[5].a/w3288 ), .B(
        \SUBBYTES[5].a/w3297 ), .Z(n11398) );
  XOR \SUBBYTES[5].a/U4997  ( .A(n11400), .B(n11399), .Z(\SUBBYTES[5].a/w3312 ) );
  XOR \SUBBYTES[5].a/U4996  ( .A(n11402), .B(n11401), .Z(n11399) );
  XOR \SUBBYTES[5].a/U4995  ( .A(\w1[5][7] ), .B(\SUBBYTES[5].a/w3396 ), .Z(
        n11400) );
  XOR \SUBBYTES[5].a/U4994  ( .A(\SUBBYTES[5].a/w3303 ), .B(
        \SUBBYTES[5].a/w3306 ), .Z(n11401) );
  XOR \SUBBYTES[5].a/U4993  ( .A(\SUBBYTES[5].a/w3289 ), .B(
        \SUBBYTES[5].a/w3291 ), .Z(n11402) );
  XOR \SUBBYTES[5].a/U4992  ( .A(n11404), .B(n11403), .Z(\SUBBYTES[5].a/w3313 ) );
  XOR \SUBBYTES[5].a/U4991  ( .A(n12109), .B(n11405), .Z(n11403) );
  XOR \SUBBYTES[5].a/U4990  ( .A(\w1[5][5] ), .B(n12110), .Z(n11404) );
  XOR \SUBBYTES[5].a/U4989  ( .A(\SUBBYTES[5].a/w3303 ), .B(
        \SUBBYTES[5].a/w3304 ), .Z(n11405) );
  XOR \SUBBYTES[5].a/U4988  ( .A(n11407), .B(n11406), .Z(\SUBBYTES[5].a/w3329 ) );
  XOR \SUBBYTES[5].a/U4987  ( .A(\w1[5][1] ), .B(n11408), .Z(n11406) );
  XOR \SUBBYTES[5].a/U4986  ( .A(\SUBBYTES[5].a/w3304 ), .B(
        \SUBBYTES[5].a/w3306 ), .Z(n11407) );
  XOR \SUBBYTES[5].a/U4985  ( .A(\SUBBYTES[5].a/w3288 ), .B(
        \SUBBYTES[5].a/w3289 ), .Z(n11408) );
  XOR \SUBBYTES[5].a/U4984  ( .A(\w1[5][9] ), .B(n11409), .Z(n12111) );
  XOR \SUBBYTES[5].a/U4983  ( .A(\w1[5][11] ), .B(\w1[5][10] ), .Z(n11409) );
  XOR \SUBBYTES[5].a/U4982  ( .A(\w1[5][14] ), .B(n12111), .Z(
        \SUBBYTES[5].a/w3171 ) );
  XOR \SUBBYTES[5].a/U4981  ( .A(\w1[5][8] ), .B(\SUBBYTES[5].a/w3171 ), .Z(
        \SUBBYTES[5].a/w3058 ) );
  XOR \SUBBYTES[5].a/U4980  ( .A(\w1[5][8] ), .B(n11410), .Z(
        \SUBBYTES[5].a/w3059 ) );
  XOR \SUBBYTES[5].a/U4979  ( .A(\w1[5][14] ), .B(\w1[5][13] ), .Z(n11410) );
  XOR \SUBBYTES[5].a/U4978  ( .A(\w1[5][13] ), .B(n12111), .Z(
        \SUBBYTES[5].a/w3189 ) );
  XOR \SUBBYTES[5].a/U4977  ( .A(n11412), .B(n11411), .Z(\SUBBYTES[5].a/w3182 ) );
  XOR \SUBBYTES[5].a/U4976  ( .A(\w1[5][11] ), .B(\w1[5][9] ), .Z(n11411) );
  XOR \SUBBYTES[5].a/U4975  ( .A(\w1[5][15] ), .B(\w1[5][12] ), .Z(n11412) );
  XOR \SUBBYTES[5].a/U4974  ( .A(\w1[5][8] ), .B(\SUBBYTES[5].a/w3182 ), .Z(
        \SUBBYTES[5].a/w3061 ) );
  XOR \SUBBYTES[5].a/U4973  ( .A(n11414), .B(n11413), .Z(\SUBBYTES[5].a/w3169 ) );
  XOR \SUBBYTES[5].a/U4972  ( .A(\SUBBYTES[5].a/w3130 ), .B(n1035), .Z(n11413)
         );
  XOR \SUBBYTES[5].a/U4971  ( .A(\SUBBYTES[5].a/w3123 ), .B(
        \SUBBYTES[5].a/w3126 ), .Z(n11414) );
  XOR \SUBBYTES[5].a/U4970  ( .A(n11416), .B(n11415), .Z(\SUBBYTES[5].a/w3170 ) );
  XOR \SUBBYTES[5].a/U4969  ( .A(\SUBBYTES[5].a/w3130 ), .B(n10981), .Z(n11415) );
  XOR \SUBBYTES[5].a/U4968  ( .A(\SUBBYTES[5].a/w3123 ), .B(n10980), .Z(n11416) );
  XOR \SUBBYTES[5].a/U4967  ( .A(\SUBBYTES[5].a/w3182 ), .B(n11417), .Z(
        \SUBBYTES[5].a/w3172 ) );
  XOR \SUBBYTES[5].a/U4966  ( .A(\w1[5][14] ), .B(\w1[5][13] ), .Z(n11417) );
  XOR \SUBBYTES[5].a/U4965  ( .A(n11419), .B(n11418), .Z(\SUBBYTES[5].a/w3173 ) );
  XOR \SUBBYTES[5].a/U4964  ( .A(n10981), .B(n1035), .Z(n11418) );
  XOR \SUBBYTES[5].a/U4963  ( .A(n10980), .B(\SUBBYTES[5].a/w3126 ), .Z(n11419) );
  XOR \SUBBYTES[5].a/U4962  ( .A(\w1[5][15] ), .B(\w1[5][10] ), .Z(n12117) );
  XOR \SUBBYTES[5].a/U4961  ( .A(n12117), .B(n11420), .Z(\SUBBYTES[5].a/w3174 ) );
  XOR \SUBBYTES[5].a/U4960  ( .A(\w1[5][13] ), .B(\w1[5][12] ), .Z(n11420) );
  XOR \SUBBYTES[5].a/U4959  ( .A(\w1[5][15] ), .B(\SUBBYTES[5].a/w3059 ), .Z(
        \SUBBYTES[5].a/w3062 ) );
  XOR \SUBBYTES[5].a/U4958  ( .A(\w1[5][9] ), .B(\SUBBYTES[5].a/w3059 ), .Z(
        \SUBBYTES[5].a/w3063 ) );
  XOR \SUBBYTES[5].a/U4957  ( .A(\w1[5][12] ), .B(\SUBBYTES[5].a/w3059 ), .Z(
        \SUBBYTES[5].a/w3064 ) );
  XOR \SUBBYTES[5].a/U4956  ( .A(\SUBBYTES[5].a/w3063 ), .B(n12117), .Z(
        \SUBBYTES[5].a/w3065 ) );
  XOR \SUBBYTES[5].a/U4955  ( .A(n12117), .B(n11421), .Z(\SUBBYTES[5].a/w3150 ) );
  XOR \SUBBYTES[5].a/U4954  ( .A(\w1[5][12] ), .B(\w1[5][9] ), .Z(n11421) );
  XOR \SUBBYTES[5].a/U4953  ( .A(n11423), .B(n11422), .Z(n12114) );
  XOR \SUBBYTES[5].a/U4952  ( .A(\w1[5][12] ), .B(n11424), .Z(n11422) );
  XOR \SUBBYTES[5].a/U4951  ( .A(\SUBBYTES[5].a/w3115 ), .B(\w1[5][14] ), .Z(
        n11423) );
  XOR \SUBBYTES[5].a/U4950  ( .A(\SUBBYTES[5].a/w3089 ), .B(
        \SUBBYTES[5].a/w3096 ), .Z(n11424) );
  XOR \SUBBYTES[5].a/U4949  ( .A(n11426), .B(n11425), .Z(n12112) );
  XOR \SUBBYTES[5].a/U4948  ( .A(\w1[5][9] ), .B(n11427), .Z(n11425) );
  XOR \SUBBYTES[5].a/U4947  ( .A(\SUBBYTES[5].a/w3114 ), .B(\w1[5][13] ), .Z(
        n11426) );
  XOR \SUBBYTES[5].a/U4946  ( .A(\SUBBYTES[5].a/w3090 ), .B(
        \SUBBYTES[5].a/w3097 ), .Z(n11427) );
  XOR \SUBBYTES[5].a/U4945  ( .A(n12114), .B(n12112), .Z(\SUBBYTES[5].a/w3120 ) );
  XOR \SUBBYTES[5].a/U4944  ( .A(\w1[5][13] ), .B(n11428), .Z(n12115) );
  XOR \SUBBYTES[5].a/U4943  ( .A(\SUBBYTES[5].a/w3082 ), .B(
        \SUBBYTES[5].a/w3092 ), .Z(n11428) );
  XOR \SUBBYTES[5].a/U4942  ( .A(n11430), .B(n11429), .Z(\SUBBYTES[5].a/w3107 ) );
  XOR \SUBBYTES[5].a/U4941  ( .A(n12115), .B(n11431), .Z(n11429) );
  XOR \SUBBYTES[5].a/U4940  ( .A(\w1[5][12] ), .B(\SUBBYTES[5].a/w3171 ), .Z(
        n11430) );
  XOR \SUBBYTES[5].a/U4939  ( .A(\SUBBYTES[5].a/w3084 ), .B(
        \SUBBYTES[5].a/w3089 ), .Z(n11431) );
  XOR \SUBBYTES[5].a/U4938  ( .A(n11433), .B(n11432), .Z(n12113) );
  XOR \SUBBYTES[5].a/U4937  ( .A(\SUBBYTES[5].a/w3117 ), .B(\w1[5][15] ), .Z(
        n11432) );
  XOR \SUBBYTES[5].a/U4936  ( .A(\SUBBYTES[5].a/w3092 ), .B(
        \SUBBYTES[5].a/w3099 ), .Z(n11433) );
  XOR \SUBBYTES[5].a/U4935  ( .A(n12112), .B(n12113), .Z(\SUBBYTES[5].a/w3119 ) );
  XOR \SUBBYTES[5].a/U4934  ( .A(\w1[5][11] ), .B(n11434), .Z(n12116) );
  XOR \SUBBYTES[5].a/U4933  ( .A(\SUBBYTES[5].a/w3081 ), .B(
        \SUBBYTES[5].a/w3084 ), .Z(n11434) );
  XOR \SUBBYTES[5].a/U4932  ( .A(n11436), .B(n11435), .Z(\SUBBYTES[5].a/w3108 ) );
  XOR \SUBBYTES[5].a/U4931  ( .A(n12116), .B(n11437), .Z(n11435) );
  XOR \SUBBYTES[5].a/U4930  ( .A(\w1[5][14] ), .B(\SUBBYTES[5].a/w3150 ), .Z(
        n11436) );
  XOR \SUBBYTES[5].a/U4929  ( .A(\SUBBYTES[5].a/w3089 ), .B(
        \SUBBYTES[5].a/w3090 ), .Z(n11437) );
  XOR \SUBBYTES[5].a/U4928  ( .A(n12114), .B(n12113), .Z(\SUBBYTES[5].a/w3128 ) );
  XOR \SUBBYTES[5].a/U4927  ( .A(n11439), .B(n11438), .Z(\SUBBYTES[5].a/w3129 ) );
  XOR \SUBBYTES[5].a/U4926  ( .A(\w1[5][15] ), .B(n12115), .Z(n11438) );
  XOR \SUBBYTES[5].a/U4925  ( .A(\SUBBYTES[5].a/w3081 ), .B(
        \SUBBYTES[5].a/w3090 ), .Z(n11439) );
  XOR \SUBBYTES[5].a/U4924  ( .A(n11441), .B(n11440), .Z(\SUBBYTES[5].a/w3105 ) );
  XOR \SUBBYTES[5].a/U4923  ( .A(n11443), .B(n11442), .Z(n11440) );
  XOR \SUBBYTES[5].a/U4922  ( .A(\w1[5][15] ), .B(\SUBBYTES[5].a/w3189 ), .Z(
        n11441) );
  XOR \SUBBYTES[5].a/U4921  ( .A(\SUBBYTES[5].a/w3096 ), .B(
        \SUBBYTES[5].a/w3099 ), .Z(n11442) );
  XOR \SUBBYTES[5].a/U4920  ( .A(\SUBBYTES[5].a/w3082 ), .B(
        \SUBBYTES[5].a/w3084 ), .Z(n11443) );
  XOR \SUBBYTES[5].a/U4919  ( .A(n11445), .B(n11444), .Z(\SUBBYTES[5].a/w3106 ) );
  XOR \SUBBYTES[5].a/U4918  ( .A(n12116), .B(n11446), .Z(n11444) );
  XOR \SUBBYTES[5].a/U4917  ( .A(\w1[5][13] ), .B(n12117), .Z(n11445) );
  XOR \SUBBYTES[5].a/U4916  ( .A(\SUBBYTES[5].a/w3096 ), .B(
        \SUBBYTES[5].a/w3097 ), .Z(n11446) );
  XOR \SUBBYTES[5].a/U4915  ( .A(n11448), .B(n11447), .Z(\SUBBYTES[5].a/w3122 ) );
  XOR \SUBBYTES[5].a/U4914  ( .A(\w1[5][9] ), .B(n11449), .Z(n11447) );
  XOR \SUBBYTES[5].a/U4913  ( .A(\SUBBYTES[5].a/w3097 ), .B(
        \SUBBYTES[5].a/w3099 ), .Z(n11448) );
  XOR \SUBBYTES[5].a/U4912  ( .A(\SUBBYTES[5].a/w3081 ), .B(
        \SUBBYTES[5].a/w3082 ), .Z(n11449) );
  XOR \SUBBYTES[5].a/U4911  ( .A(\w1[5][17] ), .B(n11450), .Z(n12118) );
  XOR \SUBBYTES[5].a/U4910  ( .A(\w1[5][19] ), .B(\w1[5][18] ), .Z(n11450) );
  XOR \SUBBYTES[5].a/U4909  ( .A(\w1[5][22] ), .B(n12118), .Z(
        \SUBBYTES[5].a/w2964 ) );
  XOR \SUBBYTES[5].a/U4908  ( .A(\w1[5][16] ), .B(\SUBBYTES[5].a/w2964 ), .Z(
        \SUBBYTES[5].a/w2851 ) );
  XOR \SUBBYTES[5].a/U4907  ( .A(\w1[5][16] ), .B(n11451), .Z(
        \SUBBYTES[5].a/w2852 ) );
  XOR \SUBBYTES[5].a/U4906  ( .A(\w1[5][22] ), .B(\w1[5][21] ), .Z(n11451) );
  XOR \SUBBYTES[5].a/U4905  ( .A(\w1[5][21] ), .B(n12118), .Z(
        \SUBBYTES[5].a/w2982 ) );
  XOR \SUBBYTES[5].a/U4904  ( .A(n11453), .B(n11452), .Z(\SUBBYTES[5].a/w2975 ) );
  XOR \SUBBYTES[5].a/U4903  ( .A(\w1[5][19] ), .B(\w1[5][17] ), .Z(n11452) );
  XOR \SUBBYTES[5].a/U4902  ( .A(\w1[5][23] ), .B(\w1[5][20] ), .Z(n11453) );
  XOR \SUBBYTES[5].a/U4901  ( .A(\w1[5][16] ), .B(\SUBBYTES[5].a/w2975 ), .Z(
        \SUBBYTES[5].a/w2854 ) );
  XOR \SUBBYTES[5].a/U4900  ( .A(n11455), .B(n11454), .Z(\SUBBYTES[5].a/w2962 ) );
  XOR \SUBBYTES[5].a/U4899  ( .A(\SUBBYTES[5].a/w2923 ), .B(n1034), .Z(n11454)
         );
  XOR \SUBBYTES[5].a/U4898  ( .A(\SUBBYTES[5].a/w2916 ), .B(
        \SUBBYTES[5].a/w2919 ), .Z(n11455) );
  XOR \SUBBYTES[5].a/U4897  ( .A(n11457), .B(n11456), .Z(\SUBBYTES[5].a/w2963 ) );
  XOR \SUBBYTES[5].a/U4896  ( .A(\SUBBYTES[5].a/w2923 ), .B(n10979), .Z(n11456) );
  XOR \SUBBYTES[5].a/U4895  ( .A(\SUBBYTES[5].a/w2916 ), .B(n10978), .Z(n11457) );
  XOR \SUBBYTES[5].a/U4894  ( .A(\SUBBYTES[5].a/w2975 ), .B(n11458), .Z(
        \SUBBYTES[5].a/w2965 ) );
  XOR \SUBBYTES[5].a/U4893  ( .A(\w1[5][22] ), .B(\w1[5][21] ), .Z(n11458) );
  XOR \SUBBYTES[5].a/U4892  ( .A(n11460), .B(n11459), .Z(\SUBBYTES[5].a/w2966 ) );
  XOR \SUBBYTES[5].a/U4891  ( .A(n10979), .B(n1034), .Z(n11459) );
  XOR \SUBBYTES[5].a/U4890  ( .A(n10978), .B(\SUBBYTES[5].a/w2919 ), .Z(n11460) );
  XOR \SUBBYTES[5].a/U4889  ( .A(\w1[5][23] ), .B(\w1[5][18] ), .Z(n12124) );
  XOR \SUBBYTES[5].a/U4888  ( .A(n12124), .B(n11461), .Z(\SUBBYTES[5].a/w2967 ) );
  XOR \SUBBYTES[5].a/U4887  ( .A(\w1[5][21] ), .B(\w1[5][20] ), .Z(n11461) );
  XOR \SUBBYTES[5].a/U4886  ( .A(\w1[5][23] ), .B(\SUBBYTES[5].a/w2852 ), .Z(
        \SUBBYTES[5].a/w2855 ) );
  XOR \SUBBYTES[5].a/U4885  ( .A(\w1[5][17] ), .B(\SUBBYTES[5].a/w2852 ), .Z(
        \SUBBYTES[5].a/w2856 ) );
  XOR \SUBBYTES[5].a/U4884  ( .A(\w1[5][20] ), .B(\SUBBYTES[5].a/w2852 ), .Z(
        \SUBBYTES[5].a/w2857 ) );
  XOR \SUBBYTES[5].a/U4883  ( .A(\SUBBYTES[5].a/w2856 ), .B(n12124), .Z(
        \SUBBYTES[5].a/w2858 ) );
  XOR \SUBBYTES[5].a/U4882  ( .A(n12124), .B(n11462), .Z(\SUBBYTES[5].a/w2943 ) );
  XOR \SUBBYTES[5].a/U4881  ( .A(\w1[5][20] ), .B(\w1[5][17] ), .Z(n11462) );
  XOR \SUBBYTES[5].a/U4880  ( .A(n11464), .B(n11463), .Z(n12121) );
  XOR \SUBBYTES[5].a/U4879  ( .A(\w1[5][20] ), .B(n11465), .Z(n11463) );
  XOR \SUBBYTES[5].a/U4878  ( .A(\SUBBYTES[5].a/w2908 ), .B(\w1[5][22] ), .Z(
        n11464) );
  XOR \SUBBYTES[5].a/U4877  ( .A(\SUBBYTES[5].a/w2882 ), .B(
        \SUBBYTES[5].a/w2889 ), .Z(n11465) );
  XOR \SUBBYTES[5].a/U4876  ( .A(n11467), .B(n11466), .Z(n12119) );
  XOR \SUBBYTES[5].a/U4875  ( .A(\w1[5][17] ), .B(n11468), .Z(n11466) );
  XOR \SUBBYTES[5].a/U4874  ( .A(\SUBBYTES[5].a/w2907 ), .B(\w1[5][21] ), .Z(
        n11467) );
  XOR \SUBBYTES[5].a/U4873  ( .A(\SUBBYTES[5].a/w2883 ), .B(
        \SUBBYTES[5].a/w2890 ), .Z(n11468) );
  XOR \SUBBYTES[5].a/U4872  ( .A(n12121), .B(n12119), .Z(\SUBBYTES[5].a/w2913 ) );
  XOR \SUBBYTES[5].a/U4871  ( .A(\w1[5][21] ), .B(n11469), .Z(n12122) );
  XOR \SUBBYTES[5].a/U4870  ( .A(\SUBBYTES[5].a/w2875 ), .B(
        \SUBBYTES[5].a/w2885 ), .Z(n11469) );
  XOR \SUBBYTES[5].a/U4869  ( .A(n11471), .B(n11470), .Z(\SUBBYTES[5].a/w2900 ) );
  XOR \SUBBYTES[5].a/U4868  ( .A(n12122), .B(n11472), .Z(n11470) );
  XOR \SUBBYTES[5].a/U4867  ( .A(\w1[5][20] ), .B(\SUBBYTES[5].a/w2964 ), .Z(
        n11471) );
  XOR \SUBBYTES[5].a/U4866  ( .A(\SUBBYTES[5].a/w2877 ), .B(
        \SUBBYTES[5].a/w2882 ), .Z(n11472) );
  XOR \SUBBYTES[5].a/U4865  ( .A(n11474), .B(n11473), .Z(n12120) );
  XOR \SUBBYTES[5].a/U4864  ( .A(\SUBBYTES[5].a/w2910 ), .B(\w1[5][23] ), .Z(
        n11473) );
  XOR \SUBBYTES[5].a/U4863  ( .A(\SUBBYTES[5].a/w2885 ), .B(
        \SUBBYTES[5].a/w2892 ), .Z(n11474) );
  XOR \SUBBYTES[5].a/U4862  ( .A(n12119), .B(n12120), .Z(\SUBBYTES[5].a/w2912 ) );
  XOR \SUBBYTES[5].a/U4861  ( .A(\w1[5][19] ), .B(n11475), .Z(n12123) );
  XOR \SUBBYTES[5].a/U4860  ( .A(\SUBBYTES[5].a/w2874 ), .B(
        \SUBBYTES[5].a/w2877 ), .Z(n11475) );
  XOR \SUBBYTES[5].a/U4859  ( .A(n11477), .B(n11476), .Z(\SUBBYTES[5].a/w2901 ) );
  XOR \SUBBYTES[5].a/U4858  ( .A(n12123), .B(n11478), .Z(n11476) );
  XOR \SUBBYTES[5].a/U4857  ( .A(\w1[5][22] ), .B(\SUBBYTES[5].a/w2943 ), .Z(
        n11477) );
  XOR \SUBBYTES[5].a/U4856  ( .A(\SUBBYTES[5].a/w2882 ), .B(
        \SUBBYTES[5].a/w2883 ), .Z(n11478) );
  XOR \SUBBYTES[5].a/U4855  ( .A(n12121), .B(n12120), .Z(\SUBBYTES[5].a/w2921 ) );
  XOR \SUBBYTES[5].a/U4854  ( .A(n11480), .B(n11479), .Z(\SUBBYTES[5].a/w2922 ) );
  XOR \SUBBYTES[5].a/U4853  ( .A(\w1[5][23] ), .B(n12122), .Z(n11479) );
  XOR \SUBBYTES[5].a/U4852  ( .A(\SUBBYTES[5].a/w2874 ), .B(
        \SUBBYTES[5].a/w2883 ), .Z(n11480) );
  XOR \SUBBYTES[5].a/U4851  ( .A(n11482), .B(n11481), .Z(\SUBBYTES[5].a/w2898 ) );
  XOR \SUBBYTES[5].a/U4850  ( .A(n11484), .B(n11483), .Z(n11481) );
  XOR \SUBBYTES[5].a/U4849  ( .A(\w1[5][23] ), .B(\SUBBYTES[5].a/w2982 ), .Z(
        n11482) );
  XOR \SUBBYTES[5].a/U4848  ( .A(\SUBBYTES[5].a/w2889 ), .B(
        \SUBBYTES[5].a/w2892 ), .Z(n11483) );
  XOR \SUBBYTES[5].a/U4847  ( .A(\SUBBYTES[5].a/w2875 ), .B(
        \SUBBYTES[5].a/w2877 ), .Z(n11484) );
  XOR \SUBBYTES[5].a/U4846  ( .A(n11486), .B(n11485), .Z(\SUBBYTES[5].a/w2899 ) );
  XOR \SUBBYTES[5].a/U4845  ( .A(n12123), .B(n11487), .Z(n11485) );
  XOR \SUBBYTES[5].a/U4844  ( .A(\w1[5][21] ), .B(n12124), .Z(n11486) );
  XOR \SUBBYTES[5].a/U4843  ( .A(\SUBBYTES[5].a/w2889 ), .B(
        \SUBBYTES[5].a/w2890 ), .Z(n11487) );
  XOR \SUBBYTES[5].a/U4842  ( .A(n11489), .B(n11488), .Z(\SUBBYTES[5].a/w2915 ) );
  XOR \SUBBYTES[5].a/U4841  ( .A(\w1[5][17] ), .B(n11490), .Z(n11488) );
  XOR \SUBBYTES[5].a/U4840  ( .A(\SUBBYTES[5].a/w2890 ), .B(
        \SUBBYTES[5].a/w2892 ), .Z(n11489) );
  XOR \SUBBYTES[5].a/U4839  ( .A(\SUBBYTES[5].a/w2874 ), .B(
        \SUBBYTES[5].a/w2875 ), .Z(n11490) );
  XOR \SUBBYTES[5].a/U4838  ( .A(\w1[5][25] ), .B(n11491), .Z(n12125) );
  XOR \SUBBYTES[5].a/U4837  ( .A(\w1[5][27] ), .B(\w1[5][26] ), .Z(n11491) );
  XOR \SUBBYTES[5].a/U4836  ( .A(\w1[5][30] ), .B(n12125), .Z(
        \SUBBYTES[5].a/w2757 ) );
  XOR \SUBBYTES[5].a/U4835  ( .A(\w1[5][24] ), .B(\SUBBYTES[5].a/w2757 ), .Z(
        \SUBBYTES[5].a/w2644 ) );
  XOR \SUBBYTES[5].a/U4834  ( .A(\w1[5][24] ), .B(n11492), .Z(
        \SUBBYTES[5].a/w2645 ) );
  XOR \SUBBYTES[5].a/U4833  ( .A(\w1[5][30] ), .B(\w1[5][29] ), .Z(n11492) );
  XOR \SUBBYTES[5].a/U4832  ( .A(\w1[5][29] ), .B(n12125), .Z(
        \SUBBYTES[5].a/w2775 ) );
  XOR \SUBBYTES[5].a/U4831  ( .A(n11494), .B(n11493), .Z(\SUBBYTES[5].a/w2768 ) );
  XOR \SUBBYTES[5].a/U4830  ( .A(\w1[5][27] ), .B(\w1[5][25] ), .Z(n11493) );
  XOR \SUBBYTES[5].a/U4829  ( .A(\w1[5][31] ), .B(\w1[5][28] ), .Z(n11494) );
  XOR \SUBBYTES[5].a/U4828  ( .A(\w1[5][24] ), .B(\SUBBYTES[5].a/w2768 ), .Z(
        \SUBBYTES[5].a/w2647 ) );
  XOR \SUBBYTES[5].a/U4827  ( .A(n11496), .B(n11495), .Z(\SUBBYTES[5].a/w2755 ) );
  XOR \SUBBYTES[5].a/U4826  ( .A(\SUBBYTES[5].a/w2716 ), .B(n1033), .Z(n11495)
         );
  XOR \SUBBYTES[5].a/U4825  ( .A(\SUBBYTES[5].a/w2709 ), .B(
        \SUBBYTES[5].a/w2712 ), .Z(n11496) );
  XOR \SUBBYTES[5].a/U4824  ( .A(n11498), .B(n11497), .Z(\SUBBYTES[5].a/w2756 ) );
  XOR \SUBBYTES[5].a/U4823  ( .A(\SUBBYTES[5].a/w2716 ), .B(n10977), .Z(n11497) );
  XOR \SUBBYTES[5].a/U4822  ( .A(\SUBBYTES[5].a/w2709 ), .B(n10976), .Z(n11498) );
  XOR \SUBBYTES[5].a/U4821  ( .A(\SUBBYTES[5].a/w2768 ), .B(n11499), .Z(
        \SUBBYTES[5].a/w2758 ) );
  XOR \SUBBYTES[5].a/U4820  ( .A(\w1[5][30] ), .B(\w1[5][29] ), .Z(n11499) );
  XOR \SUBBYTES[5].a/U4819  ( .A(n11501), .B(n11500), .Z(\SUBBYTES[5].a/w2759 ) );
  XOR \SUBBYTES[5].a/U4818  ( .A(n10977), .B(n1033), .Z(n11500) );
  XOR \SUBBYTES[5].a/U4817  ( .A(n10976), .B(\SUBBYTES[5].a/w2712 ), .Z(n11501) );
  XOR \SUBBYTES[5].a/U4816  ( .A(\w1[5][31] ), .B(\w1[5][26] ), .Z(n12131) );
  XOR \SUBBYTES[5].a/U4815  ( .A(n12131), .B(n11502), .Z(\SUBBYTES[5].a/w2760 ) );
  XOR \SUBBYTES[5].a/U4814  ( .A(\w1[5][29] ), .B(\w1[5][28] ), .Z(n11502) );
  XOR \SUBBYTES[5].a/U4813  ( .A(\w1[5][31] ), .B(\SUBBYTES[5].a/w2645 ), .Z(
        \SUBBYTES[5].a/w2648 ) );
  XOR \SUBBYTES[5].a/U4812  ( .A(\w1[5][25] ), .B(\SUBBYTES[5].a/w2645 ), .Z(
        \SUBBYTES[5].a/w2649 ) );
  XOR \SUBBYTES[5].a/U4811  ( .A(\w1[5][28] ), .B(\SUBBYTES[5].a/w2645 ), .Z(
        \SUBBYTES[5].a/w2650 ) );
  XOR \SUBBYTES[5].a/U4810  ( .A(\SUBBYTES[5].a/w2649 ), .B(n12131), .Z(
        \SUBBYTES[5].a/w2651 ) );
  XOR \SUBBYTES[5].a/U4809  ( .A(n12131), .B(n11503), .Z(\SUBBYTES[5].a/w2736 ) );
  XOR \SUBBYTES[5].a/U4808  ( .A(\w1[5][28] ), .B(\w1[5][25] ), .Z(n11503) );
  XOR \SUBBYTES[5].a/U4807  ( .A(n11505), .B(n11504), .Z(n12128) );
  XOR \SUBBYTES[5].a/U4806  ( .A(\w1[5][28] ), .B(n11506), .Z(n11504) );
  XOR \SUBBYTES[5].a/U4805  ( .A(\SUBBYTES[5].a/w2701 ), .B(\w1[5][30] ), .Z(
        n11505) );
  XOR \SUBBYTES[5].a/U4804  ( .A(\SUBBYTES[5].a/w2675 ), .B(
        \SUBBYTES[5].a/w2682 ), .Z(n11506) );
  XOR \SUBBYTES[5].a/U4803  ( .A(n11508), .B(n11507), .Z(n12126) );
  XOR \SUBBYTES[5].a/U4802  ( .A(\w1[5][25] ), .B(n11509), .Z(n11507) );
  XOR \SUBBYTES[5].a/U4801  ( .A(\SUBBYTES[5].a/w2700 ), .B(\w1[5][29] ), .Z(
        n11508) );
  XOR \SUBBYTES[5].a/U4800  ( .A(\SUBBYTES[5].a/w2676 ), .B(
        \SUBBYTES[5].a/w2683 ), .Z(n11509) );
  XOR \SUBBYTES[5].a/U4799  ( .A(n12128), .B(n12126), .Z(\SUBBYTES[5].a/w2706 ) );
  XOR \SUBBYTES[5].a/U4798  ( .A(\w1[5][29] ), .B(n11510), .Z(n12129) );
  XOR \SUBBYTES[5].a/U4797  ( .A(\SUBBYTES[5].a/w2668 ), .B(
        \SUBBYTES[5].a/w2678 ), .Z(n11510) );
  XOR \SUBBYTES[5].a/U4796  ( .A(n11512), .B(n11511), .Z(\SUBBYTES[5].a/w2693 ) );
  XOR \SUBBYTES[5].a/U4795  ( .A(n12129), .B(n11513), .Z(n11511) );
  XOR \SUBBYTES[5].a/U4794  ( .A(\w1[5][28] ), .B(\SUBBYTES[5].a/w2757 ), .Z(
        n11512) );
  XOR \SUBBYTES[5].a/U4793  ( .A(\SUBBYTES[5].a/w2670 ), .B(
        \SUBBYTES[5].a/w2675 ), .Z(n11513) );
  XOR \SUBBYTES[5].a/U4792  ( .A(n11515), .B(n11514), .Z(n12127) );
  XOR \SUBBYTES[5].a/U4791  ( .A(\SUBBYTES[5].a/w2703 ), .B(\w1[5][31] ), .Z(
        n11514) );
  XOR \SUBBYTES[5].a/U4790  ( .A(\SUBBYTES[5].a/w2678 ), .B(
        \SUBBYTES[5].a/w2685 ), .Z(n11515) );
  XOR \SUBBYTES[5].a/U4789  ( .A(n12126), .B(n12127), .Z(\SUBBYTES[5].a/w2705 ) );
  XOR \SUBBYTES[5].a/U4788  ( .A(\w1[5][27] ), .B(n11516), .Z(n12130) );
  XOR \SUBBYTES[5].a/U4787  ( .A(\SUBBYTES[5].a/w2667 ), .B(
        \SUBBYTES[5].a/w2670 ), .Z(n11516) );
  XOR \SUBBYTES[5].a/U4786  ( .A(n11518), .B(n11517), .Z(\SUBBYTES[5].a/w2694 ) );
  XOR \SUBBYTES[5].a/U4785  ( .A(n12130), .B(n11519), .Z(n11517) );
  XOR \SUBBYTES[5].a/U4784  ( .A(\w1[5][30] ), .B(\SUBBYTES[5].a/w2736 ), .Z(
        n11518) );
  XOR \SUBBYTES[5].a/U4783  ( .A(\SUBBYTES[5].a/w2675 ), .B(
        \SUBBYTES[5].a/w2676 ), .Z(n11519) );
  XOR \SUBBYTES[5].a/U4782  ( .A(n12128), .B(n12127), .Z(\SUBBYTES[5].a/w2714 ) );
  XOR \SUBBYTES[5].a/U4781  ( .A(n11521), .B(n11520), .Z(\SUBBYTES[5].a/w2715 ) );
  XOR \SUBBYTES[5].a/U4780  ( .A(\w1[5][31] ), .B(n12129), .Z(n11520) );
  XOR \SUBBYTES[5].a/U4779  ( .A(\SUBBYTES[5].a/w2667 ), .B(
        \SUBBYTES[5].a/w2676 ), .Z(n11521) );
  XOR \SUBBYTES[5].a/U4778  ( .A(n11523), .B(n11522), .Z(\SUBBYTES[5].a/w2691 ) );
  XOR \SUBBYTES[5].a/U4777  ( .A(n11525), .B(n11524), .Z(n11522) );
  XOR \SUBBYTES[5].a/U4776  ( .A(\w1[5][31] ), .B(\SUBBYTES[5].a/w2775 ), .Z(
        n11523) );
  XOR \SUBBYTES[5].a/U4775  ( .A(\SUBBYTES[5].a/w2682 ), .B(
        \SUBBYTES[5].a/w2685 ), .Z(n11524) );
  XOR \SUBBYTES[5].a/U4774  ( .A(\SUBBYTES[5].a/w2668 ), .B(
        \SUBBYTES[5].a/w2670 ), .Z(n11525) );
  XOR \SUBBYTES[5].a/U4773  ( .A(n11527), .B(n11526), .Z(\SUBBYTES[5].a/w2692 ) );
  XOR \SUBBYTES[5].a/U4772  ( .A(n12130), .B(n11528), .Z(n11526) );
  XOR \SUBBYTES[5].a/U4771  ( .A(\w1[5][29] ), .B(n12131), .Z(n11527) );
  XOR \SUBBYTES[5].a/U4770  ( .A(\SUBBYTES[5].a/w2682 ), .B(
        \SUBBYTES[5].a/w2683 ), .Z(n11528) );
  XOR \SUBBYTES[5].a/U4769  ( .A(n11530), .B(n11529), .Z(\SUBBYTES[5].a/w2708 ) );
  XOR \SUBBYTES[5].a/U4768  ( .A(\w1[5][25] ), .B(n11531), .Z(n11529) );
  XOR \SUBBYTES[5].a/U4767  ( .A(\SUBBYTES[5].a/w2683 ), .B(
        \SUBBYTES[5].a/w2685 ), .Z(n11530) );
  XOR \SUBBYTES[5].a/U4766  ( .A(\SUBBYTES[5].a/w2667 ), .B(
        \SUBBYTES[5].a/w2668 ), .Z(n11531) );
  XOR \SUBBYTES[5].a/U4765  ( .A(\w1[5][33] ), .B(n11532), .Z(n12132) );
  XOR \SUBBYTES[5].a/U4764  ( .A(\w1[5][35] ), .B(\w1[5][34] ), .Z(n11532) );
  XOR \SUBBYTES[5].a/U4763  ( .A(\w1[5][38] ), .B(n12132), .Z(
        \SUBBYTES[5].a/w2550 ) );
  XOR \SUBBYTES[5].a/U4762  ( .A(\w1[5][32] ), .B(\SUBBYTES[5].a/w2550 ), .Z(
        \SUBBYTES[5].a/w2437 ) );
  XOR \SUBBYTES[5].a/U4761  ( .A(\w1[5][32] ), .B(n11533), .Z(
        \SUBBYTES[5].a/w2438 ) );
  XOR \SUBBYTES[5].a/U4760  ( .A(\w1[5][38] ), .B(\w1[5][37] ), .Z(n11533) );
  XOR \SUBBYTES[5].a/U4759  ( .A(\w1[5][37] ), .B(n12132), .Z(
        \SUBBYTES[5].a/w2568 ) );
  XOR \SUBBYTES[5].a/U4758  ( .A(n11535), .B(n11534), .Z(\SUBBYTES[5].a/w2561 ) );
  XOR \SUBBYTES[5].a/U4757  ( .A(\w1[5][35] ), .B(\w1[5][33] ), .Z(n11534) );
  XOR \SUBBYTES[5].a/U4756  ( .A(\w1[5][39] ), .B(\w1[5][36] ), .Z(n11535) );
  XOR \SUBBYTES[5].a/U4755  ( .A(\w1[5][32] ), .B(\SUBBYTES[5].a/w2561 ), .Z(
        \SUBBYTES[5].a/w2440 ) );
  XOR \SUBBYTES[5].a/U4754  ( .A(n11537), .B(n11536), .Z(\SUBBYTES[5].a/w2548 ) );
  XOR \SUBBYTES[5].a/U4753  ( .A(\SUBBYTES[5].a/w2509 ), .B(n1032), .Z(n11536)
         );
  XOR \SUBBYTES[5].a/U4752  ( .A(\SUBBYTES[5].a/w2502 ), .B(
        \SUBBYTES[5].a/w2505 ), .Z(n11537) );
  XOR \SUBBYTES[5].a/U4751  ( .A(n11539), .B(n11538), .Z(\SUBBYTES[5].a/w2549 ) );
  XOR \SUBBYTES[5].a/U4750  ( .A(\SUBBYTES[5].a/w2509 ), .B(n10975), .Z(n11538) );
  XOR \SUBBYTES[5].a/U4749  ( .A(\SUBBYTES[5].a/w2502 ), .B(n10974), .Z(n11539) );
  XOR \SUBBYTES[5].a/U4748  ( .A(\SUBBYTES[5].a/w2561 ), .B(n11540), .Z(
        \SUBBYTES[5].a/w2551 ) );
  XOR \SUBBYTES[5].a/U4747  ( .A(\w1[5][38] ), .B(\w1[5][37] ), .Z(n11540) );
  XOR \SUBBYTES[5].a/U4746  ( .A(n11542), .B(n11541), .Z(\SUBBYTES[5].a/w2552 ) );
  XOR \SUBBYTES[5].a/U4745  ( .A(n10975), .B(n1032), .Z(n11541) );
  XOR \SUBBYTES[5].a/U4744  ( .A(n10974), .B(\SUBBYTES[5].a/w2505 ), .Z(n11542) );
  XOR \SUBBYTES[5].a/U4743  ( .A(\w1[5][39] ), .B(\w1[5][34] ), .Z(n12138) );
  XOR \SUBBYTES[5].a/U4742  ( .A(n12138), .B(n11543), .Z(\SUBBYTES[5].a/w2553 ) );
  XOR \SUBBYTES[5].a/U4741  ( .A(\w1[5][37] ), .B(\w1[5][36] ), .Z(n11543) );
  XOR \SUBBYTES[5].a/U4740  ( .A(\w1[5][39] ), .B(\SUBBYTES[5].a/w2438 ), .Z(
        \SUBBYTES[5].a/w2441 ) );
  XOR \SUBBYTES[5].a/U4739  ( .A(\w1[5][33] ), .B(\SUBBYTES[5].a/w2438 ), .Z(
        \SUBBYTES[5].a/w2442 ) );
  XOR \SUBBYTES[5].a/U4738  ( .A(\w1[5][36] ), .B(\SUBBYTES[5].a/w2438 ), .Z(
        \SUBBYTES[5].a/w2443 ) );
  XOR \SUBBYTES[5].a/U4737  ( .A(\SUBBYTES[5].a/w2442 ), .B(n12138), .Z(
        \SUBBYTES[5].a/w2444 ) );
  XOR \SUBBYTES[5].a/U4736  ( .A(n12138), .B(n11544), .Z(\SUBBYTES[5].a/w2529 ) );
  XOR \SUBBYTES[5].a/U4735  ( .A(\w1[5][36] ), .B(\w1[5][33] ), .Z(n11544) );
  XOR \SUBBYTES[5].a/U4734  ( .A(n11546), .B(n11545), .Z(n12135) );
  XOR \SUBBYTES[5].a/U4733  ( .A(\w1[5][36] ), .B(n11547), .Z(n11545) );
  XOR \SUBBYTES[5].a/U4732  ( .A(\SUBBYTES[5].a/w2494 ), .B(\w1[5][38] ), .Z(
        n11546) );
  XOR \SUBBYTES[5].a/U4731  ( .A(\SUBBYTES[5].a/w2468 ), .B(
        \SUBBYTES[5].a/w2475 ), .Z(n11547) );
  XOR \SUBBYTES[5].a/U4730  ( .A(n11549), .B(n11548), .Z(n12133) );
  XOR \SUBBYTES[5].a/U4729  ( .A(\w1[5][33] ), .B(n11550), .Z(n11548) );
  XOR \SUBBYTES[5].a/U4728  ( .A(\SUBBYTES[5].a/w2493 ), .B(\w1[5][37] ), .Z(
        n11549) );
  XOR \SUBBYTES[5].a/U4727  ( .A(\SUBBYTES[5].a/w2469 ), .B(
        \SUBBYTES[5].a/w2476 ), .Z(n11550) );
  XOR \SUBBYTES[5].a/U4726  ( .A(n12135), .B(n12133), .Z(\SUBBYTES[5].a/w2499 ) );
  XOR \SUBBYTES[5].a/U4725  ( .A(\w1[5][37] ), .B(n11551), .Z(n12136) );
  XOR \SUBBYTES[5].a/U4724  ( .A(\SUBBYTES[5].a/w2461 ), .B(
        \SUBBYTES[5].a/w2471 ), .Z(n11551) );
  XOR \SUBBYTES[5].a/U4723  ( .A(n11553), .B(n11552), .Z(\SUBBYTES[5].a/w2486 ) );
  XOR \SUBBYTES[5].a/U4722  ( .A(n12136), .B(n11554), .Z(n11552) );
  XOR \SUBBYTES[5].a/U4721  ( .A(\w1[5][36] ), .B(\SUBBYTES[5].a/w2550 ), .Z(
        n11553) );
  XOR \SUBBYTES[5].a/U4720  ( .A(\SUBBYTES[5].a/w2463 ), .B(
        \SUBBYTES[5].a/w2468 ), .Z(n11554) );
  XOR \SUBBYTES[5].a/U4719  ( .A(n11556), .B(n11555), .Z(n12134) );
  XOR \SUBBYTES[5].a/U4718  ( .A(\SUBBYTES[5].a/w2496 ), .B(\w1[5][39] ), .Z(
        n11555) );
  XOR \SUBBYTES[5].a/U4717  ( .A(\SUBBYTES[5].a/w2471 ), .B(
        \SUBBYTES[5].a/w2478 ), .Z(n11556) );
  XOR \SUBBYTES[5].a/U4716  ( .A(n12133), .B(n12134), .Z(\SUBBYTES[5].a/w2498 ) );
  XOR \SUBBYTES[5].a/U4715  ( .A(\w1[5][35] ), .B(n11557), .Z(n12137) );
  XOR \SUBBYTES[5].a/U4714  ( .A(\SUBBYTES[5].a/w2460 ), .B(
        \SUBBYTES[5].a/w2463 ), .Z(n11557) );
  XOR \SUBBYTES[5].a/U4713  ( .A(n11559), .B(n11558), .Z(\SUBBYTES[5].a/w2487 ) );
  XOR \SUBBYTES[5].a/U4712  ( .A(n12137), .B(n11560), .Z(n11558) );
  XOR \SUBBYTES[5].a/U4711  ( .A(\w1[5][38] ), .B(\SUBBYTES[5].a/w2529 ), .Z(
        n11559) );
  XOR \SUBBYTES[5].a/U4710  ( .A(\SUBBYTES[5].a/w2468 ), .B(
        \SUBBYTES[5].a/w2469 ), .Z(n11560) );
  XOR \SUBBYTES[5].a/U4709  ( .A(n12135), .B(n12134), .Z(\SUBBYTES[5].a/w2507 ) );
  XOR \SUBBYTES[5].a/U4708  ( .A(n11562), .B(n11561), .Z(\SUBBYTES[5].a/w2508 ) );
  XOR \SUBBYTES[5].a/U4707  ( .A(\w1[5][39] ), .B(n12136), .Z(n11561) );
  XOR \SUBBYTES[5].a/U4706  ( .A(\SUBBYTES[5].a/w2460 ), .B(
        \SUBBYTES[5].a/w2469 ), .Z(n11562) );
  XOR \SUBBYTES[5].a/U4705  ( .A(n11564), .B(n11563), .Z(\SUBBYTES[5].a/w2484 ) );
  XOR \SUBBYTES[5].a/U4704  ( .A(n11566), .B(n11565), .Z(n11563) );
  XOR \SUBBYTES[5].a/U4703  ( .A(\w1[5][39] ), .B(\SUBBYTES[5].a/w2568 ), .Z(
        n11564) );
  XOR \SUBBYTES[5].a/U4702  ( .A(\SUBBYTES[5].a/w2475 ), .B(
        \SUBBYTES[5].a/w2478 ), .Z(n11565) );
  XOR \SUBBYTES[5].a/U4701  ( .A(\SUBBYTES[5].a/w2461 ), .B(
        \SUBBYTES[5].a/w2463 ), .Z(n11566) );
  XOR \SUBBYTES[5].a/U4700  ( .A(n11568), .B(n11567), .Z(\SUBBYTES[5].a/w2485 ) );
  XOR \SUBBYTES[5].a/U4699  ( .A(n12137), .B(n11569), .Z(n11567) );
  XOR \SUBBYTES[5].a/U4698  ( .A(\w1[5][37] ), .B(n12138), .Z(n11568) );
  XOR \SUBBYTES[5].a/U4697  ( .A(\SUBBYTES[5].a/w2475 ), .B(
        \SUBBYTES[5].a/w2476 ), .Z(n11569) );
  XOR \SUBBYTES[5].a/U4696  ( .A(n11571), .B(n11570), .Z(\SUBBYTES[5].a/w2501 ) );
  XOR \SUBBYTES[5].a/U4695  ( .A(\w1[5][33] ), .B(n11572), .Z(n11570) );
  XOR \SUBBYTES[5].a/U4694  ( .A(\SUBBYTES[5].a/w2476 ), .B(
        \SUBBYTES[5].a/w2478 ), .Z(n11571) );
  XOR \SUBBYTES[5].a/U4693  ( .A(\SUBBYTES[5].a/w2460 ), .B(
        \SUBBYTES[5].a/w2461 ), .Z(n11572) );
  XOR \SUBBYTES[5].a/U4692  ( .A(\w1[5][41] ), .B(n11573), .Z(n12139) );
  XOR \SUBBYTES[5].a/U4691  ( .A(\w1[5][43] ), .B(\w1[5][42] ), .Z(n11573) );
  XOR \SUBBYTES[5].a/U4690  ( .A(\w1[5][46] ), .B(n12139), .Z(
        \SUBBYTES[5].a/w2343 ) );
  XOR \SUBBYTES[5].a/U4689  ( .A(\w1[5][40] ), .B(\SUBBYTES[5].a/w2343 ), .Z(
        \SUBBYTES[5].a/w2230 ) );
  XOR \SUBBYTES[5].a/U4688  ( .A(\w1[5][40] ), .B(n11574), .Z(
        \SUBBYTES[5].a/w2231 ) );
  XOR \SUBBYTES[5].a/U4687  ( .A(\w1[5][46] ), .B(\w1[5][45] ), .Z(n11574) );
  XOR \SUBBYTES[5].a/U4686  ( .A(\w1[5][45] ), .B(n12139), .Z(
        \SUBBYTES[5].a/w2361 ) );
  XOR \SUBBYTES[5].a/U4685  ( .A(n11576), .B(n11575), .Z(\SUBBYTES[5].a/w2354 ) );
  XOR \SUBBYTES[5].a/U4684  ( .A(\w1[5][43] ), .B(\w1[5][41] ), .Z(n11575) );
  XOR \SUBBYTES[5].a/U4683  ( .A(\w1[5][47] ), .B(\w1[5][44] ), .Z(n11576) );
  XOR \SUBBYTES[5].a/U4682  ( .A(\w1[5][40] ), .B(\SUBBYTES[5].a/w2354 ), .Z(
        \SUBBYTES[5].a/w2233 ) );
  XOR \SUBBYTES[5].a/U4681  ( .A(n11578), .B(n11577), .Z(\SUBBYTES[5].a/w2341 ) );
  XOR \SUBBYTES[5].a/U4680  ( .A(\SUBBYTES[5].a/w2302 ), .B(n1031), .Z(n11577)
         );
  XOR \SUBBYTES[5].a/U4679  ( .A(\SUBBYTES[5].a/w2295 ), .B(
        \SUBBYTES[5].a/w2298 ), .Z(n11578) );
  XOR \SUBBYTES[5].a/U4678  ( .A(n11580), .B(n11579), .Z(\SUBBYTES[5].a/w2342 ) );
  XOR \SUBBYTES[5].a/U4677  ( .A(\SUBBYTES[5].a/w2302 ), .B(n10973), .Z(n11579) );
  XOR \SUBBYTES[5].a/U4676  ( .A(\SUBBYTES[5].a/w2295 ), .B(n10972), .Z(n11580) );
  XOR \SUBBYTES[5].a/U4675  ( .A(\SUBBYTES[5].a/w2354 ), .B(n11581), .Z(
        \SUBBYTES[5].a/w2344 ) );
  XOR \SUBBYTES[5].a/U4674  ( .A(\w1[5][46] ), .B(\w1[5][45] ), .Z(n11581) );
  XOR \SUBBYTES[5].a/U4673  ( .A(n11583), .B(n11582), .Z(\SUBBYTES[5].a/w2345 ) );
  XOR \SUBBYTES[5].a/U4672  ( .A(n10973), .B(n1031), .Z(n11582) );
  XOR \SUBBYTES[5].a/U4671  ( .A(n10972), .B(\SUBBYTES[5].a/w2298 ), .Z(n11583) );
  XOR \SUBBYTES[5].a/U4670  ( .A(\w1[5][47] ), .B(\w1[5][42] ), .Z(n12145) );
  XOR \SUBBYTES[5].a/U4669  ( .A(n12145), .B(n11584), .Z(\SUBBYTES[5].a/w2346 ) );
  XOR \SUBBYTES[5].a/U4668  ( .A(\w1[5][45] ), .B(\w1[5][44] ), .Z(n11584) );
  XOR \SUBBYTES[5].a/U4667  ( .A(\w1[5][47] ), .B(\SUBBYTES[5].a/w2231 ), .Z(
        \SUBBYTES[5].a/w2234 ) );
  XOR \SUBBYTES[5].a/U4666  ( .A(\w1[5][41] ), .B(\SUBBYTES[5].a/w2231 ), .Z(
        \SUBBYTES[5].a/w2235 ) );
  XOR \SUBBYTES[5].a/U4665  ( .A(\w1[5][44] ), .B(\SUBBYTES[5].a/w2231 ), .Z(
        \SUBBYTES[5].a/w2236 ) );
  XOR \SUBBYTES[5].a/U4664  ( .A(\SUBBYTES[5].a/w2235 ), .B(n12145), .Z(
        \SUBBYTES[5].a/w2237 ) );
  XOR \SUBBYTES[5].a/U4663  ( .A(n12145), .B(n11585), .Z(\SUBBYTES[5].a/w2322 ) );
  XOR \SUBBYTES[5].a/U4662  ( .A(\w1[5][44] ), .B(\w1[5][41] ), .Z(n11585) );
  XOR \SUBBYTES[5].a/U4661  ( .A(n11587), .B(n11586), .Z(n12142) );
  XOR \SUBBYTES[5].a/U4660  ( .A(\w1[5][44] ), .B(n11588), .Z(n11586) );
  XOR \SUBBYTES[5].a/U4659  ( .A(\SUBBYTES[5].a/w2287 ), .B(\w1[5][46] ), .Z(
        n11587) );
  XOR \SUBBYTES[5].a/U4658  ( .A(\SUBBYTES[5].a/w2261 ), .B(
        \SUBBYTES[5].a/w2268 ), .Z(n11588) );
  XOR \SUBBYTES[5].a/U4657  ( .A(n11590), .B(n11589), .Z(n12140) );
  XOR \SUBBYTES[5].a/U4656  ( .A(\w1[5][41] ), .B(n11591), .Z(n11589) );
  XOR \SUBBYTES[5].a/U4655  ( .A(\SUBBYTES[5].a/w2286 ), .B(\w1[5][45] ), .Z(
        n11590) );
  XOR \SUBBYTES[5].a/U4654  ( .A(\SUBBYTES[5].a/w2262 ), .B(
        \SUBBYTES[5].a/w2269 ), .Z(n11591) );
  XOR \SUBBYTES[5].a/U4653  ( .A(n12142), .B(n12140), .Z(\SUBBYTES[5].a/w2292 ) );
  XOR \SUBBYTES[5].a/U4652  ( .A(\w1[5][45] ), .B(n11592), .Z(n12143) );
  XOR \SUBBYTES[5].a/U4651  ( .A(\SUBBYTES[5].a/w2254 ), .B(
        \SUBBYTES[5].a/w2264 ), .Z(n11592) );
  XOR \SUBBYTES[5].a/U4650  ( .A(n11594), .B(n11593), .Z(\SUBBYTES[5].a/w2279 ) );
  XOR \SUBBYTES[5].a/U4649  ( .A(n12143), .B(n11595), .Z(n11593) );
  XOR \SUBBYTES[5].a/U4648  ( .A(\w1[5][44] ), .B(\SUBBYTES[5].a/w2343 ), .Z(
        n11594) );
  XOR \SUBBYTES[5].a/U4647  ( .A(\SUBBYTES[5].a/w2256 ), .B(
        \SUBBYTES[5].a/w2261 ), .Z(n11595) );
  XOR \SUBBYTES[5].a/U4646  ( .A(n11597), .B(n11596), .Z(n12141) );
  XOR \SUBBYTES[5].a/U4645  ( .A(\SUBBYTES[5].a/w2289 ), .B(\w1[5][47] ), .Z(
        n11596) );
  XOR \SUBBYTES[5].a/U4644  ( .A(\SUBBYTES[5].a/w2264 ), .B(
        \SUBBYTES[5].a/w2271 ), .Z(n11597) );
  XOR \SUBBYTES[5].a/U4643  ( .A(n12140), .B(n12141), .Z(\SUBBYTES[5].a/w2291 ) );
  XOR \SUBBYTES[5].a/U4642  ( .A(\w1[5][43] ), .B(n11598), .Z(n12144) );
  XOR \SUBBYTES[5].a/U4641  ( .A(\SUBBYTES[5].a/w2253 ), .B(
        \SUBBYTES[5].a/w2256 ), .Z(n11598) );
  XOR \SUBBYTES[5].a/U4640  ( .A(n11600), .B(n11599), .Z(\SUBBYTES[5].a/w2280 ) );
  XOR \SUBBYTES[5].a/U4639  ( .A(n12144), .B(n11601), .Z(n11599) );
  XOR \SUBBYTES[5].a/U4638  ( .A(\w1[5][46] ), .B(\SUBBYTES[5].a/w2322 ), .Z(
        n11600) );
  XOR \SUBBYTES[5].a/U4637  ( .A(\SUBBYTES[5].a/w2261 ), .B(
        \SUBBYTES[5].a/w2262 ), .Z(n11601) );
  XOR \SUBBYTES[5].a/U4636  ( .A(n12142), .B(n12141), .Z(\SUBBYTES[5].a/w2300 ) );
  XOR \SUBBYTES[5].a/U4635  ( .A(n11603), .B(n11602), .Z(\SUBBYTES[5].a/w2301 ) );
  XOR \SUBBYTES[5].a/U4634  ( .A(\w1[5][47] ), .B(n12143), .Z(n11602) );
  XOR \SUBBYTES[5].a/U4633  ( .A(\SUBBYTES[5].a/w2253 ), .B(
        \SUBBYTES[5].a/w2262 ), .Z(n11603) );
  XOR \SUBBYTES[5].a/U4632  ( .A(n11605), .B(n11604), .Z(\SUBBYTES[5].a/w2277 ) );
  XOR \SUBBYTES[5].a/U4631  ( .A(n11607), .B(n11606), .Z(n11604) );
  XOR \SUBBYTES[5].a/U4630  ( .A(\w1[5][47] ), .B(\SUBBYTES[5].a/w2361 ), .Z(
        n11605) );
  XOR \SUBBYTES[5].a/U4629  ( .A(\SUBBYTES[5].a/w2268 ), .B(
        \SUBBYTES[5].a/w2271 ), .Z(n11606) );
  XOR \SUBBYTES[5].a/U4628  ( .A(\SUBBYTES[5].a/w2254 ), .B(
        \SUBBYTES[5].a/w2256 ), .Z(n11607) );
  XOR \SUBBYTES[5].a/U4627  ( .A(n11609), .B(n11608), .Z(\SUBBYTES[5].a/w2278 ) );
  XOR \SUBBYTES[5].a/U4626  ( .A(n12144), .B(n11610), .Z(n11608) );
  XOR \SUBBYTES[5].a/U4625  ( .A(\w1[5][45] ), .B(n12145), .Z(n11609) );
  XOR \SUBBYTES[5].a/U4624  ( .A(\SUBBYTES[5].a/w2268 ), .B(
        \SUBBYTES[5].a/w2269 ), .Z(n11610) );
  XOR \SUBBYTES[5].a/U4623  ( .A(n11612), .B(n11611), .Z(\SUBBYTES[5].a/w2294 ) );
  XOR \SUBBYTES[5].a/U4622  ( .A(\w1[5][41] ), .B(n11613), .Z(n11611) );
  XOR \SUBBYTES[5].a/U4621  ( .A(\SUBBYTES[5].a/w2269 ), .B(
        \SUBBYTES[5].a/w2271 ), .Z(n11612) );
  XOR \SUBBYTES[5].a/U4620  ( .A(\SUBBYTES[5].a/w2253 ), .B(
        \SUBBYTES[5].a/w2254 ), .Z(n11613) );
  XOR \SUBBYTES[5].a/U4619  ( .A(\w1[5][49] ), .B(n11614), .Z(n12146) );
  XOR \SUBBYTES[5].a/U4618  ( .A(\w1[5][51] ), .B(\w1[5][50] ), .Z(n11614) );
  XOR \SUBBYTES[5].a/U4617  ( .A(\w1[5][54] ), .B(n12146), .Z(
        \SUBBYTES[5].a/w2136 ) );
  XOR \SUBBYTES[5].a/U4616  ( .A(\w1[5][48] ), .B(\SUBBYTES[5].a/w2136 ), .Z(
        \SUBBYTES[5].a/w2023 ) );
  XOR \SUBBYTES[5].a/U4615  ( .A(\w1[5][48] ), .B(n11615), .Z(
        \SUBBYTES[5].a/w2024 ) );
  XOR \SUBBYTES[5].a/U4614  ( .A(\w1[5][54] ), .B(\w1[5][53] ), .Z(n11615) );
  XOR \SUBBYTES[5].a/U4613  ( .A(\w1[5][53] ), .B(n12146), .Z(
        \SUBBYTES[5].a/w2154 ) );
  XOR \SUBBYTES[5].a/U4612  ( .A(n11617), .B(n11616), .Z(\SUBBYTES[5].a/w2147 ) );
  XOR \SUBBYTES[5].a/U4611  ( .A(\w1[5][51] ), .B(\w1[5][49] ), .Z(n11616) );
  XOR \SUBBYTES[5].a/U4610  ( .A(\w1[5][55] ), .B(\w1[5][52] ), .Z(n11617) );
  XOR \SUBBYTES[5].a/U4609  ( .A(\w1[5][48] ), .B(\SUBBYTES[5].a/w2147 ), .Z(
        \SUBBYTES[5].a/w2026 ) );
  XOR \SUBBYTES[5].a/U4608  ( .A(n11619), .B(n11618), .Z(\SUBBYTES[5].a/w2134 ) );
  XOR \SUBBYTES[5].a/U4607  ( .A(\SUBBYTES[5].a/w2095 ), .B(n1030), .Z(n11618)
         );
  XOR \SUBBYTES[5].a/U4606  ( .A(\SUBBYTES[5].a/w2088 ), .B(
        \SUBBYTES[5].a/w2091 ), .Z(n11619) );
  XOR \SUBBYTES[5].a/U4605  ( .A(n11621), .B(n11620), .Z(\SUBBYTES[5].a/w2135 ) );
  XOR \SUBBYTES[5].a/U4604  ( .A(\SUBBYTES[5].a/w2095 ), .B(n10971), .Z(n11620) );
  XOR \SUBBYTES[5].a/U4603  ( .A(\SUBBYTES[5].a/w2088 ), .B(n10970), .Z(n11621) );
  XOR \SUBBYTES[5].a/U4602  ( .A(\SUBBYTES[5].a/w2147 ), .B(n11622), .Z(
        \SUBBYTES[5].a/w2137 ) );
  XOR \SUBBYTES[5].a/U4601  ( .A(\w1[5][54] ), .B(\w1[5][53] ), .Z(n11622) );
  XOR \SUBBYTES[5].a/U4600  ( .A(n11624), .B(n11623), .Z(\SUBBYTES[5].a/w2138 ) );
  XOR \SUBBYTES[5].a/U4599  ( .A(n10971), .B(n1030), .Z(n11623) );
  XOR \SUBBYTES[5].a/U4598  ( .A(n10970), .B(\SUBBYTES[5].a/w2091 ), .Z(n11624) );
  XOR \SUBBYTES[5].a/U4597  ( .A(\w1[5][55] ), .B(\w1[5][50] ), .Z(n12152) );
  XOR \SUBBYTES[5].a/U4596  ( .A(n12152), .B(n11625), .Z(\SUBBYTES[5].a/w2139 ) );
  XOR \SUBBYTES[5].a/U4595  ( .A(\w1[5][53] ), .B(\w1[5][52] ), .Z(n11625) );
  XOR \SUBBYTES[5].a/U4594  ( .A(\w1[5][55] ), .B(\SUBBYTES[5].a/w2024 ), .Z(
        \SUBBYTES[5].a/w2027 ) );
  XOR \SUBBYTES[5].a/U4593  ( .A(\w1[5][49] ), .B(\SUBBYTES[5].a/w2024 ), .Z(
        \SUBBYTES[5].a/w2028 ) );
  XOR \SUBBYTES[5].a/U4592  ( .A(\w1[5][52] ), .B(\SUBBYTES[5].a/w2024 ), .Z(
        \SUBBYTES[5].a/w2029 ) );
  XOR \SUBBYTES[5].a/U4591  ( .A(\SUBBYTES[5].a/w2028 ), .B(n12152), .Z(
        \SUBBYTES[5].a/w2030 ) );
  XOR \SUBBYTES[5].a/U4590  ( .A(n12152), .B(n11626), .Z(\SUBBYTES[5].a/w2115 ) );
  XOR \SUBBYTES[5].a/U4589  ( .A(\w1[5][52] ), .B(\w1[5][49] ), .Z(n11626) );
  XOR \SUBBYTES[5].a/U4588  ( .A(n11628), .B(n11627), .Z(n12149) );
  XOR \SUBBYTES[5].a/U4587  ( .A(\w1[5][52] ), .B(n11629), .Z(n11627) );
  XOR \SUBBYTES[5].a/U4586  ( .A(\SUBBYTES[5].a/w2080 ), .B(\w1[5][54] ), .Z(
        n11628) );
  XOR \SUBBYTES[5].a/U4585  ( .A(\SUBBYTES[5].a/w2054 ), .B(
        \SUBBYTES[5].a/w2061 ), .Z(n11629) );
  XOR \SUBBYTES[5].a/U4584  ( .A(n11631), .B(n11630), .Z(n12147) );
  XOR \SUBBYTES[5].a/U4583  ( .A(\w1[5][49] ), .B(n11632), .Z(n11630) );
  XOR \SUBBYTES[5].a/U4582  ( .A(\SUBBYTES[5].a/w2079 ), .B(\w1[5][53] ), .Z(
        n11631) );
  XOR \SUBBYTES[5].a/U4581  ( .A(\SUBBYTES[5].a/w2055 ), .B(
        \SUBBYTES[5].a/w2062 ), .Z(n11632) );
  XOR \SUBBYTES[5].a/U4580  ( .A(n12149), .B(n12147), .Z(\SUBBYTES[5].a/w2085 ) );
  XOR \SUBBYTES[5].a/U4579  ( .A(\w1[5][53] ), .B(n11633), .Z(n12150) );
  XOR \SUBBYTES[5].a/U4578  ( .A(\SUBBYTES[5].a/w2047 ), .B(
        \SUBBYTES[5].a/w2057 ), .Z(n11633) );
  XOR \SUBBYTES[5].a/U4577  ( .A(n11635), .B(n11634), .Z(\SUBBYTES[5].a/w2072 ) );
  XOR \SUBBYTES[5].a/U4576  ( .A(n12150), .B(n11636), .Z(n11634) );
  XOR \SUBBYTES[5].a/U4575  ( .A(\w1[5][52] ), .B(\SUBBYTES[5].a/w2136 ), .Z(
        n11635) );
  XOR \SUBBYTES[5].a/U4574  ( .A(\SUBBYTES[5].a/w2049 ), .B(
        \SUBBYTES[5].a/w2054 ), .Z(n11636) );
  XOR \SUBBYTES[5].a/U4573  ( .A(n11638), .B(n11637), .Z(n12148) );
  XOR \SUBBYTES[5].a/U4572  ( .A(\SUBBYTES[5].a/w2082 ), .B(\w1[5][55] ), .Z(
        n11637) );
  XOR \SUBBYTES[5].a/U4571  ( .A(\SUBBYTES[5].a/w2057 ), .B(
        \SUBBYTES[5].a/w2064 ), .Z(n11638) );
  XOR \SUBBYTES[5].a/U4570  ( .A(n12147), .B(n12148), .Z(\SUBBYTES[5].a/w2084 ) );
  XOR \SUBBYTES[5].a/U4569  ( .A(\w1[5][51] ), .B(n11639), .Z(n12151) );
  XOR \SUBBYTES[5].a/U4568  ( .A(\SUBBYTES[5].a/w2046 ), .B(
        \SUBBYTES[5].a/w2049 ), .Z(n11639) );
  XOR \SUBBYTES[5].a/U4567  ( .A(n11641), .B(n11640), .Z(\SUBBYTES[5].a/w2073 ) );
  XOR \SUBBYTES[5].a/U4566  ( .A(n12151), .B(n11642), .Z(n11640) );
  XOR \SUBBYTES[5].a/U4565  ( .A(\w1[5][54] ), .B(\SUBBYTES[5].a/w2115 ), .Z(
        n11641) );
  XOR \SUBBYTES[5].a/U4564  ( .A(\SUBBYTES[5].a/w2054 ), .B(
        \SUBBYTES[5].a/w2055 ), .Z(n11642) );
  XOR \SUBBYTES[5].a/U4563  ( .A(n12149), .B(n12148), .Z(\SUBBYTES[5].a/w2093 ) );
  XOR \SUBBYTES[5].a/U4562  ( .A(n11644), .B(n11643), .Z(\SUBBYTES[5].a/w2094 ) );
  XOR \SUBBYTES[5].a/U4561  ( .A(\w1[5][55] ), .B(n12150), .Z(n11643) );
  XOR \SUBBYTES[5].a/U4560  ( .A(\SUBBYTES[5].a/w2046 ), .B(
        \SUBBYTES[5].a/w2055 ), .Z(n11644) );
  XOR \SUBBYTES[5].a/U4559  ( .A(n11646), .B(n11645), .Z(\SUBBYTES[5].a/w2070 ) );
  XOR \SUBBYTES[5].a/U4558  ( .A(n11648), .B(n11647), .Z(n11645) );
  XOR \SUBBYTES[5].a/U4557  ( .A(\w1[5][55] ), .B(\SUBBYTES[5].a/w2154 ), .Z(
        n11646) );
  XOR \SUBBYTES[5].a/U4556  ( .A(\SUBBYTES[5].a/w2061 ), .B(
        \SUBBYTES[5].a/w2064 ), .Z(n11647) );
  XOR \SUBBYTES[5].a/U4555  ( .A(\SUBBYTES[5].a/w2047 ), .B(
        \SUBBYTES[5].a/w2049 ), .Z(n11648) );
  XOR \SUBBYTES[5].a/U4554  ( .A(n11650), .B(n11649), .Z(\SUBBYTES[5].a/w2071 ) );
  XOR \SUBBYTES[5].a/U4553  ( .A(n12151), .B(n11651), .Z(n11649) );
  XOR \SUBBYTES[5].a/U4552  ( .A(\w1[5][53] ), .B(n12152), .Z(n11650) );
  XOR \SUBBYTES[5].a/U4551  ( .A(\SUBBYTES[5].a/w2061 ), .B(
        \SUBBYTES[5].a/w2062 ), .Z(n11651) );
  XOR \SUBBYTES[5].a/U4550  ( .A(n11653), .B(n11652), .Z(\SUBBYTES[5].a/w2087 ) );
  XOR \SUBBYTES[5].a/U4549  ( .A(\w1[5][49] ), .B(n11654), .Z(n11652) );
  XOR \SUBBYTES[5].a/U4548  ( .A(\SUBBYTES[5].a/w2062 ), .B(
        \SUBBYTES[5].a/w2064 ), .Z(n11653) );
  XOR \SUBBYTES[5].a/U4547  ( .A(\SUBBYTES[5].a/w2046 ), .B(
        \SUBBYTES[5].a/w2047 ), .Z(n11654) );
  XOR \SUBBYTES[5].a/U4546  ( .A(\w1[5][57] ), .B(n11655), .Z(n12153) );
  XOR \SUBBYTES[5].a/U4545  ( .A(\w1[5][59] ), .B(\w1[5][58] ), .Z(n11655) );
  XOR \SUBBYTES[5].a/U4544  ( .A(\w1[5][62] ), .B(n12153), .Z(
        \SUBBYTES[5].a/w1929 ) );
  XOR \SUBBYTES[5].a/U4543  ( .A(\w1[5][56] ), .B(\SUBBYTES[5].a/w1929 ), .Z(
        \SUBBYTES[5].a/w1816 ) );
  XOR \SUBBYTES[5].a/U4542  ( .A(\w1[5][56] ), .B(n11656), .Z(
        \SUBBYTES[5].a/w1817 ) );
  XOR \SUBBYTES[5].a/U4541  ( .A(\w1[5][62] ), .B(\w1[5][61] ), .Z(n11656) );
  XOR \SUBBYTES[5].a/U4540  ( .A(\w1[5][61] ), .B(n12153), .Z(
        \SUBBYTES[5].a/w1947 ) );
  XOR \SUBBYTES[5].a/U4539  ( .A(n11658), .B(n11657), .Z(\SUBBYTES[5].a/w1940 ) );
  XOR \SUBBYTES[5].a/U4538  ( .A(\w1[5][59] ), .B(\w1[5][57] ), .Z(n11657) );
  XOR \SUBBYTES[5].a/U4537  ( .A(\w1[5][63] ), .B(\w1[5][60] ), .Z(n11658) );
  XOR \SUBBYTES[5].a/U4536  ( .A(\w1[5][56] ), .B(\SUBBYTES[5].a/w1940 ), .Z(
        \SUBBYTES[5].a/w1819 ) );
  XOR \SUBBYTES[5].a/U4535  ( .A(n11660), .B(n11659), .Z(\SUBBYTES[5].a/w1927 ) );
  XOR \SUBBYTES[5].a/U4534  ( .A(\SUBBYTES[5].a/w1888 ), .B(n1029), .Z(n11659)
         );
  XOR \SUBBYTES[5].a/U4533  ( .A(\SUBBYTES[5].a/w1881 ), .B(
        \SUBBYTES[5].a/w1884 ), .Z(n11660) );
  XOR \SUBBYTES[5].a/U4532  ( .A(n11662), .B(n11661), .Z(\SUBBYTES[5].a/w1928 ) );
  XOR \SUBBYTES[5].a/U4531  ( .A(\SUBBYTES[5].a/w1888 ), .B(n10969), .Z(n11661) );
  XOR \SUBBYTES[5].a/U4530  ( .A(\SUBBYTES[5].a/w1881 ), .B(n10968), .Z(n11662) );
  XOR \SUBBYTES[5].a/U4529  ( .A(\SUBBYTES[5].a/w1940 ), .B(n11663), .Z(
        \SUBBYTES[5].a/w1930 ) );
  XOR \SUBBYTES[5].a/U4528  ( .A(\w1[5][62] ), .B(\w1[5][61] ), .Z(n11663) );
  XOR \SUBBYTES[5].a/U4527  ( .A(n11665), .B(n11664), .Z(\SUBBYTES[5].a/w1931 ) );
  XOR \SUBBYTES[5].a/U4526  ( .A(n10969), .B(n1029), .Z(n11664) );
  XOR \SUBBYTES[5].a/U4525  ( .A(n10968), .B(\SUBBYTES[5].a/w1884 ), .Z(n11665) );
  XOR \SUBBYTES[5].a/U4524  ( .A(\w1[5][63] ), .B(\w1[5][58] ), .Z(n12159) );
  XOR \SUBBYTES[5].a/U4523  ( .A(n12159), .B(n11666), .Z(\SUBBYTES[5].a/w1932 ) );
  XOR \SUBBYTES[5].a/U4522  ( .A(\w1[5][61] ), .B(\w1[5][60] ), .Z(n11666) );
  XOR \SUBBYTES[5].a/U4521  ( .A(\w1[5][63] ), .B(\SUBBYTES[5].a/w1817 ), .Z(
        \SUBBYTES[5].a/w1820 ) );
  XOR \SUBBYTES[5].a/U4520  ( .A(\w1[5][57] ), .B(\SUBBYTES[5].a/w1817 ), .Z(
        \SUBBYTES[5].a/w1821 ) );
  XOR \SUBBYTES[5].a/U4519  ( .A(\w1[5][60] ), .B(\SUBBYTES[5].a/w1817 ), .Z(
        \SUBBYTES[5].a/w1822 ) );
  XOR \SUBBYTES[5].a/U4518  ( .A(\SUBBYTES[5].a/w1821 ), .B(n12159), .Z(
        \SUBBYTES[5].a/w1823 ) );
  XOR \SUBBYTES[5].a/U4517  ( .A(n12159), .B(n11667), .Z(\SUBBYTES[5].a/w1908 ) );
  XOR \SUBBYTES[5].a/U4516  ( .A(\w1[5][60] ), .B(\w1[5][57] ), .Z(n11667) );
  XOR \SUBBYTES[5].a/U4515  ( .A(n11669), .B(n11668), .Z(n12156) );
  XOR \SUBBYTES[5].a/U4514  ( .A(\w1[5][60] ), .B(n11670), .Z(n11668) );
  XOR \SUBBYTES[5].a/U4513  ( .A(\SUBBYTES[5].a/w1873 ), .B(\w1[5][62] ), .Z(
        n11669) );
  XOR \SUBBYTES[5].a/U4512  ( .A(\SUBBYTES[5].a/w1847 ), .B(
        \SUBBYTES[5].a/w1854 ), .Z(n11670) );
  XOR \SUBBYTES[5].a/U4511  ( .A(n11672), .B(n11671), .Z(n12154) );
  XOR \SUBBYTES[5].a/U4510  ( .A(\w1[5][57] ), .B(n11673), .Z(n11671) );
  XOR \SUBBYTES[5].a/U4509  ( .A(\SUBBYTES[5].a/w1872 ), .B(\w1[5][61] ), .Z(
        n11672) );
  XOR \SUBBYTES[5].a/U4508  ( .A(\SUBBYTES[5].a/w1848 ), .B(
        \SUBBYTES[5].a/w1855 ), .Z(n11673) );
  XOR \SUBBYTES[5].a/U4507  ( .A(n12156), .B(n12154), .Z(\SUBBYTES[5].a/w1878 ) );
  XOR \SUBBYTES[5].a/U4506  ( .A(\w1[5][61] ), .B(n11674), .Z(n12157) );
  XOR \SUBBYTES[5].a/U4505  ( .A(\SUBBYTES[5].a/w1840 ), .B(
        \SUBBYTES[5].a/w1850 ), .Z(n11674) );
  XOR \SUBBYTES[5].a/U4504  ( .A(n11676), .B(n11675), .Z(\SUBBYTES[5].a/w1865 ) );
  XOR \SUBBYTES[5].a/U4503  ( .A(n12157), .B(n11677), .Z(n11675) );
  XOR \SUBBYTES[5].a/U4502  ( .A(\w1[5][60] ), .B(\SUBBYTES[5].a/w1929 ), .Z(
        n11676) );
  XOR \SUBBYTES[5].a/U4501  ( .A(\SUBBYTES[5].a/w1842 ), .B(
        \SUBBYTES[5].a/w1847 ), .Z(n11677) );
  XOR \SUBBYTES[5].a/U4500  ( .A(n11679), .B(n11678), .Z(n12155) );
  XOR \SUBBYTES[5].a/U4499  ( .A(\SUBBYTES[5].a/w1875 ), .B(\w1[5][63] ), .Z(
        n11678) );
  XOR \SUBBYTES[5].a/U4498  ( .A(\SUBBYTES[5].a/w1850 ), .B(
        \SUBBYTES[5].a/w1857 ), .Z(n11679) );
  XOR \SUBBYTES[5].a/U4497  ( .A(n12154), .B(n12155), .Z(\SUBBYTES[5].a/w1877 ) );
  XOR \SUBBYTES[5].a/U4496  ( .A(\w1[5][59] ), .B(n11680), .Z(n12158) );
  XOR \SUBBYTES[5].a/U4495  ( .A(\SUBBYTES[5].a/w1839 ), .B(
        \SUBBYTES[5].a/w1842 ), .Z(n11680) );
  XOR \SUBBYTES[5].a/U4494  ( .A(n11682), .B(n11681), .Z(\SUBBYTES[5].a/w1866 ) );
  XOR \SUBBYTES[5].a/U4493  ( .A(n12158), .B(n11683), .Z(n11681) );
  XOR \SUBBYTES[5].a/U4492  ( .A(\w1[5][62] ), .B(\SUBBYTES[5].a/w1908 ), .Z(
        n11682) );
  XOR \SUBBYTES[5].a/U4491  ( .A(\SUBBYTES[5].a/w1847 ), .B(
        \SUBBYTES[5].a/w1848 ), .Z(n11683) );
  XOR \SUBBYTES[5].a/U4490  ( .A(n12156), .B(n12155), .Z(\SUBBYTES[5].a/w1886 ) );
  XOR \SUBBYTES[5].a/U4489  ( .A(n11685), .B(n11684), .Z(\SUBBYTES[5].a/w1887 ) );
  XOR \SUBBYTES[5].a/U4488  ( .A(\w1[5][63] ), .B(n12157), .Z(n11684) );
  XOR \SUBBYTES[5].a/U4487  ( .A(\SUBBYTES[5].a/w1839 ), .B(
        \SUBBYTES[5].a/w1848 ), .Z(n11685) );
  XOR \SUBBYTES[5].a/U4486  ( .A(n11687), .B(n11686), .Z(\SUBBYTES[5].a/w1863 ) );
  XOR \SUBBYTES[5].a/U4485  ( .A(n11689), .B(n11688), .Z(n11686) );
  XOR \SUBBYTES[5].a/U4484  ( .A(\w1[5][63] ), .B(\SUBBYTES[5].a/w1947 ), .Z(
        n11687) );
  XOR \SUBBYTES[5].a/U4483  ( .A(\SUBBYTES[5].a/w1854 ), .B(
        \SUBBYTES[5].a/w1857 ), .Z(n11688) );
  XOR \SUBBYTES[5].a/U4482  ( .A(\SUBBYTES[5].a/w1840 ), .B(
        \SUBBYTES[5].a/w1842 ), .Z(n11689) );
  XOR \SUBBYTES[5].a/U4481  ( .A(n11691), .B(n11690), .Z(\SUBBYTES[5].a/w1864 ) );
  XOR \SUBBYTES[5].a/U4480  ( .A(n12158), .B(n11692), .Z(n11690) );
  XOR \SUBBYTES[5].a/U4479  ( .A(\w1[5][61] ), .B(n12159), .Z(n11691) );
  XOR \SUBBYTES[5].a/U4478  ( .A(\SUBBYTES[5].a/w1854 ), .B(
        \SUBBYTES[5].a/w1855 ), .Z(n11692) );
  XOR \SUBBYTES[5].a/U4477  ( .A(n11694), .B(n11693), .Z(\SUBBYTES[5].a/w1880 ) );
  XOR \SUBBYTES[5].a/U4476  ( .A(\w1[5][57] ), .B(n11695), .Z(n11693) );
  XOR \SUBBYTES[5].a/U4475  ( .A(\SUBBYTES[5].a/w1855 ), .B(
        \SUBBYTES[5].a/w1857 ), .Z(n11694) );
  XOR \SUBBYTES[5].a/U4474  ( .A(\SUBBYTES[5].a/w1839 ), .B(
        \SUBBYTES[5].a/w1840 ), .Z(n11695) );
  XOR \SUBBYTES[5].a/U4473  ( .A(\w1[5][65] ), .B(n11696), .Z(n12160) );
  XOR \SUBBYTES[5].a/U4472  ( .A(\w1[5][67] ), .B(\w1[5][66] ), .Z(n11696) );
  XOR \SUBBYTES[5].a/U4471  ( .A(\w1[5][70] ), .B(n12160), .Z(
        \SUBBYTES[5].a/w1722 ) );
  XOR \SUBBYTES[5].a/U4470  ( .A(\w1[5][64] ), .B(\SUBBYTES[5].a/w1722 ), .Z(
        \SUBBYTES[5].a/w1609 ) );
  XOR \SUBBYTES[5].a/U4469  ( .A(\w1[5][64] ), .B(n11697), .Z(
        \SUBBYTES[5].a/w1610 ) );
  XOR \SUBBYTES[5].a/U4468  ( .A(\w1[5][70] ), .B(\w1[5][69] ), .Z(n11697) );
  XOR \SUBBYTES[5].a/U4467  ( .A(\w1[5][69] ), .B(n12160), .Z(
        \SUBBYTES[5].a/w1740 ) );
  XOR \SUBBYTES[5].a/U4466  ( .A(n11699), .B(n11698), .Z(\SUBBYTES[5].a/w1733 ) );
  XOR \SUBBYTES[5].a/U4465  ( .A(\w1[5][67] ), .B(\w1[5][65] ), .Z(n11698) );
  XOR \SUBBYTES[5].a/U4464  ( .A(\w1[5][71] ), .B(\w1[5][68] ), .Z(n11699) );
  XOR \SUBBYTES[5].a/U4463  ( .A(\w1[5][64] ), .B(\SUBBYTES[5].a/w1733 ), .Z(
        \SUBBYTES[5].a/w1612 ) );
  XOR \SUBBYTES[5].a/U4462  ( .A(n11701), .B(n11700), .Z(\SUBBYTES[5].a/w1720 ) );
  XOR \SUBBYTES[5].a/U4461  ( .A(\SUBBYTES[5].a/w1681 ), .B(n1028), .Z(n11700)
         );
  XOR \SUBBYTES[5].a/U4460  ( .A(\SUBBYTES[5].a/w1674 ), .B(
        \SUBBYTES[5].a/w1677 ), .Z(n11701) );
  XOR \SUBBYTES[5].a/U4459  ( .A(n11703), .B(n11702), .Z(\SUBBYTES[5].a/w1721 ) );
  XOR \SUBBYTES[5].a/U4458  ( .A(\SUBBYTES[5].a/w1681 ), .B(n10967), .Z(n11702) );
  XOR \SUBBYTES[5].a/U4457  ( .A(\SUBBYTES[5].a/w1674 ), .B(n10966), .Z(n11703) );
  XOR \SUBBYTES[5].a/U4456  ( .A(\SUBBYTES[5].a/w1733 ), .B(n11704), .Z(
        \SUBBYTES[5].a/w1723 ) );
  XOR \SUBBYTES[5].a/U4455  ( .A(\w1[5][70] ), .B(\w1[5][69] ), .Z(n11704) );
  XOR \SUBBYTES[5].a/U4454  ( .A(n11706), .B(n11705), .Z(\SUBBYTES[5].a/w1724 ) );
  XOR \SUBBYTES[5].a/U4453  ( .A(n10967), .B(n1028), .Z(n11705) );
  XOR \SUBBYTES[5].a/U4452  ( .A(n10966), .B(\SUBBYTES[5].a/w1677 ), .Z(n11706) );
  XOR \SUBBYTES[5].a/U4451  ( .A(\w1[5][71] ), .B(\w1[5][66] ), .Z(n12166) );
  XOR \SUBBYTES[5].a/U4450  ( .A(n12166), .B(n11707), .Z(\SUBBYTES[5].a/w1725 ) );
  XOR \SUBBYTES[5].a/U4449  ( .A(\w1[5][69] ), .B(\w1[5][68] ), .Z(n11707) );
  XOR \SUBBYTES[5].a/U4448  ( .A(\w1[5][71] ), .B(\SUBBYTES[5].a/w1610 ), .Z(
        \SUBBYTES[5].a/w1613 ) );
  XOR \SUBBYTES[5].a/U4447  ( .A(\w1[5][65] ), .B(\SUBBYTES[5].a/w1610 ), .Z(
        \SUBBYTES[5].a/w1614 ) );
  XOR \SUBBYTES[5].a/U4446  ( .A(\w1[5][68] ), .B(\SUBBYTES[5].a/w1610 ), .Z(
        \SUBBYTES[5].a/w1615 ) );
  XOR \SUBBYTES[5].a/U4445  ( .A(\SUBBYTES[5].a/w1614 ), .B(n12166), .Z(
        \SUBBYTES[5].a/w1616 ) );
  XOR \SUBBYTES[5].a/U4444  ( .A(n12166), .B(n11708), .Z(\SUBBYTES[5].a/w1701 ) );
  XOR \SUBBYTES[5].a/U4443  ( .A(\w1[5][68] ), .B(\w1[5][65] ), .Z(n11708) );
  XOR \SUBBYTES[5].a/U4442  ( .A(n11710), .B(n11709), .Z(n12163) );
  XOR \SUBBYTES[5].a/U4441  ( .A(\w1[5][68] ), .B(n11711), .Z(n11709) );
  XOR \SUBBYTES[5].a/U4440  ( .A(\SUBBYTES[5].a/w1666 ), .B(\w1[5][70] ), .Z(
        n11710) );
  XOR \SUBBYTES[5].a/U4439  ( .A(\SUBBYTES[5].a/w1640 ), .B(
        \SUBBYTES[5].a/w1647 ), .Z(n11711) );
  XOR \SUBBYTES[5].a/U4438  ( .A(n11713), .B(n11712), .Z(n12161) );
  XOR \SUBBYTES[5].a/U4437  ( .A(\w1[5][65] ), .B(n11714), .Z(n11712) );
  XOR \SUBBYTES[5].a/U4436  ( .A(\SUBBYTES[5].a/w1665 ), .B(\w1[5][69] ), .Z(
        n11713) );
  XOR \SUBBYTES[5].a/U4435  ( .A(\SUBBYTES[5].a/w1641 ), .B(
        \SUBBYTES[5].a/w1648 ), .Z(n11714) );
  XOR \SUBBYTES[5].a/U4434  ( .A(n12163), .B(n12161), .Z(\SUBBYTES[5].a/w1671 ) );
  XOR \SUBBYTES[5].a/U4433  ( .A(\w1[5][69] ), .B(n11715), .Z(n12164) );
  XOR \SUBBYTES[5].a/U4432  ( .A(\SUBBYTES[5].a/w1633 ), .B(
        \SUBBYTES[5].a/w1643 ), .Z(n11715) );
  XOR \SUBBYTES[5].a/U4431  ( .A(n11717), .B(n11716), .Z(\SUBBYTES[5].a/w1658 ) );
  XOR \SUBBYTES[5].a/U4430  ( .A(n12164), .B(n11718), .Z(n11716) );
  XOR \SUBBYTES[5].a/U4429  ( .A(\w1[5][68] ), .B(\SUBBYTES[5].a/w1722 ), .Z(
        n11717) );
  XOR \SUBBYTES[5].a/U4428  ( .A(\SUBBYTES[5].a/w1635 ), .B(
        \SUBBYTES[5].a/w1640 ), .Z(n11718) );
  XOR \SUBBYTES[5].a/U4427  ( .A(n11720), .B(n11719), .Z(n12162) );
  XOR \SUBBYTES[5].a/U4426  ( .A(\SUBBYTES[5].a/w1668 ), .B(\w1[5][71] ), .Z(
        n11719) );
  XOR \SUBBYTES[5].a/U4425  ( .A(\SUBBYTES[5].a/w1643 ), .B(
        \SUBBYTES[5].a/w1650 ), .Z(n11720) );
  XOR \SUBBYTES[5].a/U4424  ( .A(n12161), .B(n12162), .Z(\SUBBYTES[5].a/w1670 ) );
  XOR \SUBBYTES[5].a/U4423  ( .A(\w1[5][67] ), .B(n11721), .Z(n12165) );
  XOR \SUBBYTES[5].a/U4422  ( .A(\SUBBYTES[5].a/w1632 ), .B(
        \SUBBYTES[5].a/w1635 ), .Z(n11721) );
  XOR \SUBBYTES[5].a/U4421  ( .A(n11723), .B(n11722), .Z(\SUBBYTES[5].a/w1659 ) );
  XOR \SUBBYTES[5].a/U4420  ( .A(n12165), .B(n11724), .Z(n11722) );
  XOR \SUBBYTES[5].a/U4419  ( .A(\w1[5][70] ), .B(\SUBBYTES[5].a/w1701 ), .Z(
        n11723) );
  XOR \SUBBYTES[5].a/U4418  ( .A(\SUBBYTES[5].a/w1640 ), .B(
        \SUBBYTES[5].a/w1641 ), .Z(n11724) );
  XOR \SUBBYTES[5].a/U4417  ( .A(n12163), .B(n12162), .Z(\SUBBYTES[5].a/w1679 ) );
  XOR \SUBBYTES[5].a/U4416  ( .A(n11726), .B(n11725), .Z(\SUBBYTES[5].a/w1680 ) );
  XOR \SUBBYTES[5].a/U4415  ( .A(\w1[5][71] ), .B(n12164), .Z(n11725) );
  XOR \SUBBYTES[5].a/U4414  ( .A(\SUBBYTES[5].a/w1632 ), .B(
        \SUBBYTES[5].a/w1641 ), .Z(n11726) );
  XOR \SUBBYTES[5].a/U4413  ( .A(n11728), .B(n11727), .Z(\SUBBYTES[5].a/w1656 ) );
  XOR \SUBBYTES[5].a/U4412  ( .A(n11730), .B(n11729), .Z(n11727) );
  XOR \SUBBYTES[5].a/U4411  ( .A(\w1[5][71] ), .B(\SUBBYTES[5].a/w1740 ), .Z(
        n11728) );
  XOR \SUBBYTES[5].a/U4410  ( .A(\SUBBYTES[5].a/w1647 ), .B(
        \SUBBYTES[5].a/w1650 ), .Z(n11729) );
  XOR \SUBBYTES[5].a/U4409  ( .A(\SUBBYTES[5].a/w1633 ), .B(
        \SUBBYTES[5].a/w1635 ), .Z(n11730) );
  XOR \SUBBYTES[5].a/U4408  ( .A(n11732), .B(n11731), .Z(\SUBBYTES[5].a/w1657 ) );
  XOR \SUBBYTES[5].a/U4407  ( .A(n12165), .B(n11733), .Z(n11731) );
  XOR \SUBBYTES[5].a/U4406  ( .A(\w1[5][69] ), .B(n12166), .Z(n11732) );
  XOR \SUBBYTES[5].a/U4405  ( .A(\SUBBYTES[5].a/w1647 ), .B(
        \SUBBYTES[5].a/w1648 ), .Z(n11733) );
  XOR \SUBBYTES[5].a/U4404  ( .A(n11735), .B(n11734), .Z(\SUBBYTES[5].a/w1673 ) );
  XOR \SUBBYTES[5].a/U4403  ( .A(\w1[5][65] ), .B(n11736), .Z(n11734) );
  XOR \SUBBYTES[5].a/U4402  ( .A(\SUBBYTES[5].a/w1648 ), .B(
        \SUBBYTES[5].a/w1650 ), .Z(n11735) );
  XOR \SUBBYTES[5].a/U4401  ( .A(\SUBBYTES[5].a/w1632 ), .B(
        \SUBBYTES[5].a/w1633 ), .Z(n11736) );
  XOR \SUBBYTES[5].a/U4400  ( .A(\w1[5][73] ), .B(n11737), .Z(n12167) );
  XOR \SUBBYTES[5].a/U4399  ( .A(\w1[5][75] ), .B(\w1[5][74] ), .Z(n11737) );
  XOR \SUBBYTES[5].a/U4398  ( .A(\w1[5][78] ), .B(n12167), .Z(
        \SUBBYTES[5].a/w1515 ) );
  XOR \SUBBYTES[5].a/U4397  ( .A(\w1[5][72] ), .B(\SUBBYTES[5].a/w1515 ), .Z(
        \SUBBYTES[5].a/w1402 ) );
  XOR \SUBBYTES[5].a/U4396  ( .A(\w1[5][72] ), .B(n11738), .Z(
        \SUBBYTES[5].a/w1403 ) );
  XOR \SUBBYTES[5].a/U4395  ( .A(\w1[5][78] ), .B(\w1[5][77] ), .Z(n11738) );
  XOR \SUBBYTES[5].a/U4394  ( .A(\w1[5][77] ), .B(n12167), .Z(
        \SUBBYTES[5].a/w1533 ) );
  XOR \SUBBYTES[5].a/U4393  ( .A(n11740), .B(n11739), .Z(\SUBBYTES[5].a/w1526 ) );
  XOR \SUBBYTES[5].a/U4392  ( .A(\w1[5][75] ), .B(\w1[5][73] ), .Z(n11739) );
  XOR \SUBBYTES[5].a/U4391  ( .A(\w1[5][79] ), .B(\w1[5][76] ), .Z(n11740) );
  XOR \SUBBYTES[5].a/U4390  ( .A(\w1[5][72] ), .B(\SUBBYTES[5].a/w1526 ), .Z(
        \SUBBYTES[5].a/w1405 ) );
  XOR \SUBBYTES[5].a/U4389  ( .A(n11742), .B(n11741), .Z(\SUBBYTES[5].a/w1513 ) );
  XOR \SUBBYTES[5].a/U4388  ( .A(\SUBBYTES[5].a/w1474 ), .B(n1027), .Z(n11741)
         );
  XOR \SUBBYTES[5].a/U4387  ( .A(\SUBBYTES[5].a/w1467 ), .B(
        \SUBBYTES[5].a/w1470 ), .Z(n11742) );
  XOR \SUBBYTES[5].a/U4386  ( .A(n11744), .B(n11743), .Z(\SUBBYTES[5].a/w1514 ) );
  XOR \SUBBYTES[5].a/U4385  ( .A(\SUBBYTES[5].a/w1474 ), .B(n10965), .Z(n11743) );
  XOR \SUBBYTES[5].a/U4384  ( .A(\SUBBYTES[5].a/w1467 ), .B(n10964), .Z(n11744) );
  XOR \SUBBYTES[5].a/U4383  ( .A(\SUBBYTES[5].a/w1526 ), .B(n11745), .Z(
        \SUBBYTES[5].a/w1516 ) );
  XOR \SUBBYTES[5].a/U4382  ( .A(\w1[5][78] ), .B(\w1[5][77] ), .Z(n11745) );
  XOR \SUBBYTES[5].a/U4381  ( .A(n11747), .B(n11746), .Z(\SUBBYTES[5].a/w1517 ) );
  XOR \SUBBYTES[5].a/U4380  ( .A(n10965), .B(n1027), .Z(n11746) );
  XOR \SUBBYTES[5].a/U4379  ( .A(n10964), .B(\SUBBYTES[5].a/w1470 ), .Z(n11747) );
  XOR \SUBBYTES[5].a/U4378  ( .A(\w1[5][79] ), .B(\w1[5][74] ), .Z(n12173) );
  XOR \SUBBYTES[5].a/U4377  ( .A(n12173), .B(n11748), .Z(\SUBBYTES[5].a/w1518 ) );
  XOR \SUBBYTES[5].a/U4376  ( .A(\w1[5][77] ), .B(\w1[5][76] ), .Z(n11748) );
  XOR \SUBBYTES[5].a/U4375  ( .A(\w1[5][79] ), .B(\SUBBYTES[5].a/w1403 ), .Z(
        \SUBBYTES[5].a/w1406 ) );
  XOR \SUBBYTES[5].a/U4374  ( .A(\w1[5][73] ), .B(\SUBBYTES[5].a/w1403 ), .Z(
        \SUBBYTES[5].a/w1407 ) );
  XOR \SUBBYTES[5].a/U4373  ( .A(\w1[5][76] ), .B(\SUBBYTES[5].a/w1403 ), .Z(
        \SUBBYTES[5].a/w1408 ) );
  XOR \SUBBYTES[5].a/U4372  ( .A(\SUBBYTES[5].a/w1407 ), .B(n12173), .Z(
        \SUBBYTES[5].a/w1409 ) );
  XOR \SUBBYTES[5].a/U4371  ( .A(n12173), .B(n11749), .Z(\SUBBYTES[5].a/w1494 ) );
  XOR \SUBBYTES[5].a/U4370  ( .A(\w1[5][76] ), .B(\w1[5][73] ), .Z(n11749) );
  XOR \SUBBYTES[5].a/U4369  ( .A(n11751), .B(n11750), .Z(n12170) );
  XOR \SUBBYTES[5].a/U4368  ( .A(\w1[5][76] ), .B(n11752), .Z(n11750) );
  XOR \SUBBYTES[5].a/U4367  ( .A(\SUBBYTES[5].a/w1459 ), .B(\w1[5][78] ), .Z(
        n11751) );
  XOR \SUBBYTES[5].a/U4366  ( .A(\SUBBYTES[5].a/w1433 ), .B(
        \SUBBYTES[5].a/w1440 ), .Z(n11752) );
  XOR \SUBBYTES[5].a/U4365  ( .A(n11754), .B(n11753), .Z(n12168) );
  XOR \SUBBYTES[5].a/U4364  ( .A(\w1[5][73] ), .B(n11755), .Z(n11753) );
  XOR \SUBBYTES[5].a/U4363  ( .A(\SUBBYTES[5].a/w1458 ), .B(\w1[5][77] ), .Z(
        n11754) );
  XOR \SUBBYTES[5].a/U4362  ( .A(\SUBBYTES[5].a/w1434 ), .B(
        \SUBBYTES[5].a/w1441 ), .Z(n11755) );
  XOR \SUBBYTES[5].a/U4361  ( .A(n12170), .B(n12168), .Z(\SUBBYTES[5].a/w1464 ) );
  XOR \SUBBYTES[5].a/U4360  ( .A(\w1[5][77] ), .B(n11756), .Z(n12171) );
  XOR \SUBBYTES[5].a/U4359  ( .A(\SUBBYTES[5].a/w1426 ), .B(
        \SUBBYTES[5].a/w1436 ), .Z(n11756) );
  XOR \SUBBYTES[5].a/U4358  ( .A(n11758), .B(n11757), .Z(\SUBBYTES[5].a/w1451 ) );
  XOR \SUBBYTES[5].a/U4357  ( .A(n12171), .B(n11759), .Z(n11757) );
  XOR \SUBBYTES[5].a/U4356  ( .A(\w1[5][76] ), .B(\SUBBYTES[5].a/w1515 ), .Z(
        n11758) );
  XOR \SUBBYTES[5].a/U4355  ( .A(\SUBBYTES[5].a/w1428 ), .B(
        \SUBBYTES[5].a/w1433 ), .Z(n11759) );
  XOR \SUBBYTES[5].a/U4354  ( .A(n11761), .B(n11760), .Z(n12169) );
  XOR \SUBBYTES[5].a/U4353  ( .A(\SUBBYTES[5].a/w1461 ), .B(\w1[5][79] ), .Z(
        n11760) );
  XOR \SUBBYTES[5].a/U4352  ( .A(\SUBBYTES[5].a/w1436 ), .B(
        \SUBBYTES[5].a/w1443 ), .Z(n11761) );
  XOR \SUBBYTES[5].a/U4351  ( .A(n12168), .B(n12169), .Z(\SUBBYTES[5].a/w1463 ) );
  XOR \SUBBYTES[5].a/U4350  ( .A(\w1[5][75] ), .B(n11762), .Z(n12172) );
  XOR \SUBBYTES[5].a/U4349  ( .A(\SUBBYTES[5].a/w1425 ), .B(
        \SUBBYTES[5].a/w1428 ), .Z(n11762) );
  XOR \SUBBYTES[5].a/U4348  ( .A(n11764), .B(n11763), .Z(\SUBBYTES[5].a/w1452 ) );
  XOR \SUBBYTES[5].a/U4347  ( .A(n12172), .B(n11765), .Z(n11763) );
  XOR \SUBBYTES[5].a/U4346  ( .A(\w1[5][78] ), .B(\SUBBYTES[5].a/w1494 ), .Z(
        n11764) );
  XOR \SUBBYTES[5].a/U4345  ( .A(\SUBBYTES[5].a/w1433 ), .B(
        \SUBBYTES[5].a/w1434 ), .Z(n11765) );
  XOR \SUBBYTES[5].a/U4344  ( .A(n12170), .B(n12169), .Z(\SUBBYTES[5].a/w1472 ) );
  XOR \SUBBYTES[5].a/U4343  ( .A(n11767), .B(n11766), .Z(\SUBBYTES[5].a/w1473 ) );
  XOR \SUBBYTES[5].a/U4342  ( .A(\w1[5][79] ), .B(n12171), .Z(n11766) );
  XOR \SUBBYTES[5].a/U4341  ( .A(\SUBBYTES[5].a/w1425 ), .B(
        \SUBBYTES[5].a/w1434 ), .Z(n11767) );
  XOR \SUBBYTES[5].a/U4340  ( .A(n11769), .B(n11768), .Z(\SUBBYTES[5].a/w1449 ) );
  XOR \SUBBYTES[5].a/U4339  ( .A(n11771), .B(n11770), .Z(n11768) );
  XOR \SUBBYTES[5].a/U4338  ( .A(\w1[5][79] ), .B(\SUBBYTES[5].a/w1533 ), .Z(
        n11769) );
  XOR \SUBBYTES[5].a/U4337  ( .A(\SUBBYTES[5].a/w1440 ), .B(
        \SUBBYTES[5].a/w1443 ), .Z(n11770) );
  XOR \SUBBYTES[5].a/U4336  ( .A(\SUBBYTES[5].a/w1426 ), .B(
        \SUBBYTES[5].a/w1428 ), .Z(n11771) );
  XOR \SUBBYTES[5].a/U4335  ( .A(n11773), .B(n11772), .Z(\SUBBYTES[5].a/w1450 ) );
  XOR \SUBBYTES[5].a/U4334  ( .A(n12172), .B(n11774), .Z(n11772) );
  XOR \SUBBYTES[5].a/U4333  ( .A(\w1[5][77] ), .B(n12173), .Z(n11773) );
  XOR \SUBBYTES[5].a/U4332  ( .A(\SUBBYTES[5].a/w1440 ), .B(
        \SUBBYTES[5].a/w1441 ), .Z(n11774) );
  XOR \SUBBYTES[5].a/U4331  ( .A(n11776), .B(n11775), .Z(\SUBBYTES[5].a/w1466 ) );
  XOR \SUBBYTES[5].a/U4330  ( .A(\w1[5][73] ), .B(n11777), .Z(n11775) );
  XOR \SUBBYTES[5].a/U4329  ( .A(\SUBBYTES[5].a/w1441 ), .B(
        \SUBBYTES[5].a/w1443 ), .Z(n11776) );
  XOR \SUBBYTES[5].a/U4328  ( .A(\SUBBYTES[5].a/w1425 ), .B(
        \SUBBYTES[5].a/w1426 ), .Z(n11777) );
  XOR \SUBBYTES[5].a/U4327  ( .A(\w1[5][81] ), .B(n11778), .Z(n12174) );
  XOR \SUBBYTES[5].a/U4326  ( .A(\w1[5][83] ), .B(\w1[5][82] ), .Z(n11778) );
  XOR \SUBBYTES[5].a/U4325  ( .A(\w1[5][86] ), .B(n12174), .Z(
        \SUBBYTES[5].a/w1308 ) );
  XOR \SUBBYTES[5].a/U4324  ( .A(\w1[5][80] ), .B(\SUBBYTES[5].a/w1308 ), .Z(
        \SUBBYTES[5].a/w1195 ) );
  XOR \SUBBYTES[5].a/U4323  ( .A(\w1[5][80] ), .B(n11779), .Z(
        \SUBBYTES[5].a/w1196 ) );
  XOR \SUBBYTES[5].a/U4322  ( .A(\w1[5][86] ), .B(\w1[5][85] ), .Z(n11779) );
  XOR \SUBBYTES[5].a/U4321  ( .A(\w1[5][85] ), .B(n12174), .Z(
        \SUBBYTES[5].a/w1326 ) );
  XOR \SUBBYTES[5].a/U4320  ( .A(n11781), .B(n11780), .Z(\SUBBYTES[5].a/w1319 ) );
  XOR \SUBBYTES[5].a/U4319  ( .A(\w1[5][83] ), .B(\w1[5][81] ), .Z(n11780) );
  XOR \SUBBYTES[5].a/U4318  ( .A(\w1[5][87] ), .B(\w1[5][84] ), .Z(n11781) );
  XOR \SUBBYTES[5].a/U4317  ( .A(\w1[5][80] ), .B(\SUBBYTES[5].a/w1319 ), .Z(
        \SUBBYTES[5].a/w1198 ) );
  XOR \SUBBYTES[5].a/U4316  ( .A(n11783), .B(n11782), .Z(\SUBBYTES[5].a/w1306 ) );
  XOR \SUBBYTES[5].a/U4315  ( .A(\SUBBYTES[5].a/w1267 ), .B(n1026), .Z(n11782)
         );
  XOR \SUBBYTES[5].a/U4314  ( .A(\SUBBYTES[5].a/w1260 ), .B(
        \SUBBYTES[5].a/w1263 ), .Z(n11783) );
  XOR \SUBBYTES[5].a/U4313  ( .A(n11785), .B(n11784), .Z(\SUBBYTES[5].a/w1307 ) );
  XOR \SUBBYTES[5].a/U4312  ( .A(\SUBBYTES[5].a/w1267 ), .B(n10963), .Z(n11784) );
  XOR \SUBBYTES[5].a/U4311  ( .A(\SUBBYTES[5].a/w1260 ), .B(n10962), .Z(n11785) );
  XOR \SUBBYTES[5].a/U4310  ( .A(\SUBBYTES[5].a/w1319 ), .B(n11786), .Z(
        \SUBBYTES[5].a/w1309 ) );
  XOR \SUBBYTES[5].a/U4309  ( .A(\w1[5][86] ), .B(\w1[5][85] ), .Z(n11786) );
  XOR \SUBBYTES[5].a/U4308  ( .A(n11788), .B(n11787), .Z(\SUBBYTES[5].a/w1310 ) );
  XOR \SUBBYTES[5].a/U4307  ( .A(n10963), .B(n1026), .Z(n11787) );
  XOR \SUBBYTES[5].a/U4306  ( .A(n10962), .B(\SUBBYTES[5].a/w1263 ), .Z(n11788) );
  XOR \SUBBYTES[5].a/U4305  ( .A(\w1[5][87] ), .B(\w1[5][82] ), .Z(n12180) );
  XOR \SUBBYTES[5].a/U4304  ( .A(n12180), .B(n11789), .Z(\SUBBYTES[5].a/w1311 ) );
  XOR \SUBBYTES[5].a/U4303  ( .A(\w1[5][85] ), .B(\w1[5][84] ), .Z(n11789) );
  XOR \SUBBYTES[5].a/U4302  ( .A(\w1[5][87] ), .B(\SUBBYTES[5].a/w1196 ), .Z(
        \SUBBYTES[5].a/w1199 ) );
  XOR \SUBBYTES[5].a/U4301  ( .A(\w1[5][81] ), .B(\SUBBYTES[5].a/w1196 ), .Z(
        \SUBBYTES[5].a/w1200 ) );
  XOR \SUBBYTES[5].a/U4300  ( .A(\w1[5][84] ), .B(\SUBBYTES[5].a/w1196 ), .Z(
        \SUBBYTES[5].a/w1201 ) );
  XOR \SUBBYTES[5].a/U4299  ( .A(\SUBBYTES[5].a/w1200 ), .B(n12180), .Z(
        \SUBBYTES[5].a/w1202 ) );
  XOR \SUBBYTES[5].a/U4298  ( .A(n12180), .B(n11790), .Z(\SUBBYTES[5].a/w1287 ) );
  XOR \SUBBYTES[5].a/U4297  ( .A(\w1[5][84] ), .B(\w1[5][81] ), .Z(n11790) );
  XOR \SUBBYTES[5].a/U4296  ( .A(n11792), .B(n11791), .Z(n12177) );
  XOR \SUBBYTES[5].a/U4295  ( .A(\w1[5][84] ), .B(n11793), .Z(n11791) );
  XOR \SUBBYTES[5].a/U4294  ( .A(\SUBBYTES[5].a/w1252 ), .B(\w1[5][86] ), .Z(
        n11792) );
  XOR \SUBBYTES[5].a/U4293  ( .A(\SUBBYTES[5].a/w1226 ), .B(
        \SUBBYTES[5].a/w1233 ), .Z(n11793) );
  XOR \SUBBYTES[5].a/U4292  ( .A(n11795), .B(n11794), .Z(n12175) );
  XOR \SUBBYTES[5].a/U4291  ( .A(\w1[5][81] ), .B(n11796), .Z(n11794) );
  XOR \SUBBYTES[5].a/U4290  ( .A(\SUBBYTES[5].a/w1251 ), .B(\w1[5][85] ), .Z(
        n11795) );
  XOR \SUBBYTES[5].a/U4289  ( .A(\SUBBYTES[5].a/w1227 ), .B(
        \SUBBYTES[5].a/w1234 ), .Z(n11796) );
  XOR \SUBBYTES[5].a/U4288  ( .A(n12177), .B(n12175), .Z(\SUBBYTES[5].a/w1257 ) );
  XOR \SUBBYTES[5].a/U4287  ( .A(\w1[5][85] ), .B(n11797), .Z(n12178) );
  XOR \SUBBYTES[5].a/U4286  ( .A(\SUBBYTES[5].a/w1219 ), .B(
        \SUBBYTES[5].a/w1229 ), .Z(n11797) );
  XOR \SUBBYTES[5].a/U4285  ( .A(n11799), .B(n11798), .Z(\SUBBYTES[5].a/w1244 ) );
  XOR \SUBBYTES[5].a/U4284  ( .A(n12178), .B(n11800), .Z(n11798) );
  XOR \SUBBYTES[5].a/U4283  ( .A(\w1[5][84] ), .B(\SUBBYTES[5].a/w1308 ), .Z(
        n11799) );
  XOR \SUBBYTES[5].a/U4282  ( .A(\SUBBYTES[5].a/w1221 ), .B(
        \SUBBYTES[5].a/w1226 ), .Z(n11800) );
  XOR \SUBBYTES[5].a/U4281  ( .A(n11802), .B(n11801), .Z(n12176) );
  XOR \SUBBYTES[5].a/U4280  ( .A(\SUBBYTES[5].a/w1254 ), .B(\w1[5][87] ), .Z(
        n11801) );
  XOR \SUBBYTES[5].a/U4279  ( .A(\SUBBYTES[5].a/w1229 ), .B(
        \SUBBYTES[5].a/w1236 ), .Z(n11802) );
  XOR \SUBBYTES[5].a/U4278  ( .A(n12175), .B(n12176), .Z(\SUBBYTES[5].a/w1256 ) );
  XOR \SUBBYTES[5].a/U4277  ( .A(\w1[5][83] ), .B(n11803), .Z(n12179) );
  XOR \SUBBYTES[5].a/U4276  ( .A(\SUBBYTES[5].a/w1218 ), .B(
        \SUBBYTES[5].a/w1221 ), .Z(n11803) );
  XOR \SUBBYTES[5].a/U4275  ( .A(n11805), .B(n11804), .Z(\SUBBYTES[5].a/w1245 ) );
  XOR \SUBBYTES[5].a/U4274  ( .A(n12179), .B(n11806), .Z(n11804) );
  XOR \SUBBYTES[5].a/U4273  ( .A(\w1[5][86] ), .B(\SUBBYTES[5].a/w1287 ), .Z(
        n11805) );
  XOR \SUBBYTES[5].a/U4272  ( .A(\SUBBYTES[5].a/w1226 ), .B(
        \SUBBYTES[5].a/w1227 ), .Z(n11806) );
  XOR \SUBBYTES[5].a/U4271  ( .A(n12177), .B(n12176), .Z(\SUBBYTES[5].a/w1265 ) );
  XOR \SUBBYTES[5].a/U4270  ( .A(n11808), .B(n11807), .Z(\SUBBYTES[5].a/w1266 ) );
  XOR \SUBBYTES[5].a/U4269  ( .A(\w1[5][87] ), .B(n12178), .Z(n11807) );
  XOR \SUBBYTES[5].a/U4268  ( .A(\SUBBYTES[5].a/w1218 ), .B(
        \SUBBYTES[5].a/w1227 ), .Z(n11808) );
  XOR \SUBBYTES[5].a/U4267  ( .A(n11810), .B(n11809), .Z(\SUBBYTES[5].a/w1242 ) );
  XOR \SUBBYTES[5].a/U4266  ( .A(n11812), .B(n11811), .Z(n11809) );
  XOR \SUBBYTES[5].a/U4265  ( .A(\w1[5][87] ), .B(\SUBBYTES[5].a/w1326 ), .Z(
        n11810) );
  XOR \SUBBYTES[5].a/U4264  ( .A(\SUBBYTES[5].a/w1233 ), .B(
        \SUBBYTES[5].a/w1236 ), .Z(n11811) );
  XOR \SUBBYTES[5].a/U4263  ( .A(\SUBBYTES[5].a/w1219 ), .B(
        \SUBBYTES[5].a/w1221 ), .Z(n11812) );
  XOR \SUBBYTES[5].a/U4262  ( .A(n11814), .B(n11813), .Z(\SUBBYTES[5].a/w1243 ) );
  XOR \SUBBYTES[5].a/U4261  ( .A(n12179), .B(n11815), .Z(n11813) );
  XOR \SUBBYTES[5].a/U4260  ( .A(\w1[5][85] ), .B(n12180), .Z(n11814) );
  XOR \SUBBYTES[5].a/U4259  ( .A(\SUBBYTES[5].a/w1233 ), .B(
        \SUBBYTES[5].a/w1234 ), .Z(n11815) );
  XOR \SUBBYTES[5].a/U4258  ( .A(n11817), .B(n11816), .Z(\SUBBYTES[5].a/w1259 ) );
  XOR \SUBBYTES[5].a/U4257  ( .A(\w1[5][81] ), .B(n11818), .Z(n11816) );
  XOR \SUBBYTES[5].a/U4256  ( .A(\SUBBYTES[5].a/w1234 ), .B(
        \SUBBYTES[5].a/w1236 ), .Z(n11817) );
  XOR \SUBBYTES[5].a/U4255  ( .A(\SUBBYTES[5].a/w1218 ), .B(
        \SUBBYTES[5].a/w1219 ), .Z(n11818) );
  XOR \SUBBYTES[5].a/U4254  ( .A(\w1[5][89] ), .B(n11819), .Z(n12181) );
  XOR \SUBBYTES[5].a/U4253  ( .A(\w1[5][91] ), .B(\w1[5][90] ), .Z(n11819) );
  XOR \SUBBYTES[5].a/U4252  ( .A(\w1[5][94] ), .B(n12181), .Z(
        \SUBBYTES[5].a/w1101 ) );
  XOR \SUBBYTES[5].a/U4251  ( .A(\w1[5][88] ), .B(\SUBBYTES[5].a/w1101 ), .Z(
        \SUBBYTES[5].a/w988 ) );
  XOR \SUBBYTES[5].a/U4250  ( .A(\w1[5][88] ), .B(n11820), .Z(
        \SUBBYTES[5].a/w989 ) );
  XOR \SUBBYTES[5].a/U4249  ( .A(\w1[5][94] ), .B(\w1[5][93] ), .Z(n11820) );
  XOR \SUBBYTES[5].a/U4248  ( .A(\w1[5][93] ), .B(n12181), .Z(
        \SUBBYTES[5].a/w1119 ) );
  XOR \SUBBYTES[5].a/U4247  ( .A(n11822), .B(n11821), .Z(\SUBBYTES[5].a/w1112 ) );
  XOR \SUBBYTES[5].a/U4246  ( .A(\w1[5][91] ), .B(\w1[5][89] ), .Z(n11821) );
  XOR \SUBBYTES[5].a/U4245  ( .A(\w1[5][95] ), .B(\w1[5][92] ), .Z(n11822) );
  XOR \SUBBYTES[5].a/U4244  ( .A(\w1[5][88] ), .B(\SUBBYTES[5].a/w1112 ), .Z(
        \SUBBYTES[5].a/w991 ) );
  XOR \SUBBYTES[5].a/U4243  ( .A(n11824), .B(n11823), .Z(\SUBBYTES[5].a/w1099 ) );
  XOR \SUBBYTES[5].a/U4242  ( .A(\SUBBYTES[5].a/w1060 ), .B(n1025), .Z(n11823)
         );
  XOR \SUBBYTES[5].a/U4241  ( .A(\SUBBYTES[5].a/w1053 ), .B(
        \SUBBYTES[5].a/w1056 ), .Z(n11824) );
  XOR \SUBBYTES[5].a/U4240  ( .A(n11826), .B(n11825), .Z(\SUBBYTES[5].a/w1100 ) );
  XOR \SUBBYTES[5].a/U4239  ( .A(\SUBBYTES[5].a/w1060 ), .B(n10961), .Z(n11825) );
  XOR \SUBBYTES[5].a/U4238  ( .A(\SUBBYTES[5].a/w1053 ), .B(n10960), .Z(n11826) );
  XOR \SUBBYTES[5].a/U4237  ( .A(\SUBBYTES[5].a/w1112 ), .B(n11827), .Z(
        \SUBBYTES[5].a/w1102 ) );
  XOR \SUBBYTES[5].a/U4236  ( .A(\w1[5][94] ), .B(\w1[5][93] ), .Z(n11827) );
  XOR \SUBBYTES[5].a/U4235  ( .A(n11829), .B(n11828), .Z(\SUBBYTES[5].a/w1103 ) );
  XOR \SUBBYTES[5].a/U4234  ( .A(n10961), .B(n1025), .Z(n11828) );
  XOR \SUBBYTES[5].a/U4233  ( .A(n10960), .B(\SUBBYTES[5].a/w1056 ), .Z(n11829) );
  XOR \SUBBYTES[5].a/U4232  ( .A(\w1[5][95] ), .B(\w1[5][90] ), .Z(n12187) );
  XOR \SUBBYTES[5].a/U4231  ( .A(n12187), .B(n11830), .Z(\SUBBYTES[5].a/w1104 ) );
  XOR \SUBBYTES[5].a/U4230  ( .A(\w1[5][93] ), .B(\w1[5][92] ), .Z(n11830) );
  XOR \SUBBYTES[5].a/U4229  ( .A(\w1[5][95] ), .B(\SUBBYTES[5].a/w989 ), .Z(
        \SUBBYTES[5].a/w992 ) );
  XOR \SUBBYTES[5].a/U4228  ( .A(\w1[5][89] ), .B(\SUBBYTES[5].a/w989 ), .Z(
        \SUBBYTES[5].a/w993 ) );
  XOR \SUBBYTES[5].a/U4227  ( .A(\w1[5][92] ), .B(\SUBBYTES[5].a/w989 ), .Z(
        \SUBBYTES[5].a/w994 ) );
  XOR \SUBBYTES[5].a/U4226  ( .A(\SUBBYTES[5].a/w993 ), .B(n12187), .Z(
        \SUBBYTES[5].a/w995 ) );
  XOR \SUBBYTES[5].a/U4225  ( .A(n12187), .B(n11831), .Z(\SUBBYTES[5].a/w1080 ) );
  XOR \SUBBYTES[5].a/U4224  ( .A(\w1[5][92] ), .B(\w1[5][89] ), .Z(n11831) );
  XOR \SUBBYTES[5].a/U4223  ( .A(n11833), .B(n11832), .Z(n12184) );
  XOR \SUBBYTES[5].a/U4222  ( .A(\w1[5][92] ), .B(n11834), .Z(n11832) );
  XOR \SUBBYTES[5].a/U4221  ( .A(\SUBBYTES[5].a/w1045 ), .B(\w1[5][94] ), .Z(
        n11833) );
  XOR \SUBBYTES[5].a/U4220  ( .A(\SUBBYTES[5].a/w1019 ), .B(
        \SUBBYTES[5].a/w1026 ), .Z(n11834) );
  XOR \SUBBYTES[5].a/U4219  ( .A(n11836), .B(n11835), .Z(n12182) );
  XOR \SUBBYTES[5].a/U4218  ( .A(\w1[5][89] ), .B(n11837), .Z(n11835) );
  XOR \SUBBYTES[5].a/U4217  ( .A(\SUBBYTES[5].a/w1044 ), .B(\w1[5][93] ), .Z(
        n11836) );
  XOR \SUBBYTES[5].a/U4216  ( .A(\SUBBYTES[5].a/w1020 ), .B(
        \SUBBYTES[5].a/w1027 ), .Z(n11837) );
  XOR \SUBBYTES[5].a/U4215  ( .A(n12184), .B(n12182), .Z(\SUBBYTES[5].a/w1050 ) );
  XOR \SUBBYTES[5].a/U4214  ( .A(\w1[5][93] ), .B(n11838), .Z(n12185) );
  XOR \SUBBYTES[5].a/U4213  ( .A(\SUBBYTES[5].a/w1012 ), .B(
        \SUBBYTES[5].a/w1022 ), .Z(n11838) );
  XOR \SUBBYTES[5].a/U4212  ( .A(n11840), .B(n11839), .Z(\SUBBYTES[5].a/w1037 ) );
  XOR \SUBBYTES[5].a/U4211  ( .A(n12185), .B(n11841), .Z(n11839) );
  XOR \SUBBYTES[5].a/U4210  ( .A(\w1[5][92] ), .B(\SUBBYTES[5].a/w1101 ), .Z(
        n11840) );
  XOR \SUBBYTES[5].a/U4209  ( .A(\SUBBYTES[5].a/w1014 ), .B(
        \SUBBYTES[5].a/w1019 ), .Z(n11841) );
  XOR \SUBBYTES[5].a/U4208  ( .A(n11843), .B(n11842), .Z(n12183) );
  XOR \SUBBYTES[5].a/U4207  ( .A(\SUBBYTES[5].a/w1047 ), .B(\w1[5][95] ), .Z(
        n11842) );
  XOR \SUBBYTES[5].a/U4206  ( .A(\SUBBYTES[5].a/w1022 ), .B(
        \SUBBYTES[5].a/w1029 ), .Z(n11843) );
  XOR \SUBBYTES[5].a/U4205  ( .A(n12182), .B(n12183), .Z(\SUBBYTES[5].a/w1049 ) );
  XOR \SUBBYTES[5].a/U4204  ( .A(\w1[5][91] ), .B(n11844), .Z(n12186) );
  XOR \SUBBYTES[5].a/U4203  ( .A(\SUBBYTES[5].a/w1011 ), .B(
        \SUBBYTES[5].a/w1014 ), .Z(n11844) );
  XOR \SUBBYTES[5].a/U4202  ( .A(n11846), .B(n11845), .Z(\SUBBYTES[5].a/w1038 ) );
  XOR \SUBBYTES[5].a/U4201  ( .A(n12186), .B(n11847), .Z(n11845) );
  XOR \SUBBYTES[5].a/U4200  ( .A(\w1[5][94] ), .B(\SUBBYTES[5].a/w1080 ), .Z(
        n11846) );
  XOR \SUBBYTES[5].a/U4199  ( .A(\SUBBYTES[5].a/w1019 ), .B(
        \SUBBYTES[5].a/w1020 ), .Z(n11847) );
  XOR \SUBBYTES[5].a/U4198  ( .A(n12184), .B(n12183), .Z(\SUBBYTES[5].a/w1058 ) );
  XOR \SUBBYTES[5].a/U4197  ( .A(n11849), .B(n11848), .Z(\SUBBYTES[5].a/w1059 ) );
  XOR \SUBBYTES[5].a/U4196  ( .A(\w1[5][95] ), .B(n12185), .Z(n11848) );
  XOR \SUBBYTES[5].a/U4195  ( .A(\SUBBYTES[5].a/w1011 ), .B(
        \SUBBYTES[5].a/w1020 ), .Z(n11849) );
  XOR \SUBBYTES[5].a/U4194  ( .A(n11851), .B(n11850), .Z(\SUBBYTES[5].a/w1035 ) );
  XOR \SUBBYTES[5].a/U4193  ( .A(n11853), .B(n11852), .Z(n11850) );
  XOR \SUBBYTES[5].a/U4192  ( .A(\w1[5][95] ), .B(\SUBBYTES[5].a/w1119 ), .Z(
        n11851) );
  XOR \SUBBYTES[5].a/U4191  ( .A(\SUBBYTES[5].a/w1026 ), .B(
        \SUBBYTES[5].a/w1029 ), .Z(n11852) );
  XOR \SUBBYTES[5].a/U4190  ( .A(\SUBBYTES[5].a/w1012 ), .B(
        \SUBBYTES[5].a/w1014 ), .Z(n11853) );
  XOR \SUBBYTES[5].a/U4189  ( .A(n11855), .B(n11854), .Z(\SUBBYTES[5].a/w1036 ) );
  XOR \SUBBYTES[5].a/U4188  ( .A(n12186), .B(n11856), .Z(n11854) );
  XOR \SUBBYTES[5].a/U4187  ( .A(\w1[5][93] ), .B(n12187), .Z(n11855) );
  XOR \SUBBYTES[5].a/U4186  ( .A(\SUBBYTES[5].a/w1026 ), .B(
        \SUBBYTES[5].a/w1027 ), .Z(n11856) );
  XOR \SUBBYTES[5].a/U4185  ( .A(n11858), .B(n11857), .Z(\SUBBYTES[5].a/w1052 ) );
  XOR \SUBBYTES[5].a/U4184  ( .A(\w1[5][89] ), .B(n11859), .Z(n11857) );
  XOR \SUBBYTES[5].a/U4183  ( .A(\SUBBYTES[5].a/w1027 ), .B(
        \SUBBYTES[5].a/w1029 ), .Z(n11858) );
  XOR \SUBBYTES[5].a/U4182  ( .A(\SUBBYTES[5].a/w1011 ), .B(
        \SUBBYTES[5].a/w1012 ), .Z(n11859) );
  XOR \SUBBYTES[5].a/U4181  ( .A(\w1[5][97] ), .B(n11860), .Z(n12188) );
  XOR \SUBBYTES[5].a/U4180  ( .A(\w1[5][99] ), .B(\w1[5][98] ), .Z(n11860) );
  XOR \SUBBYTES[5].a/U4179  ( .A(\w1[5][102] ), .B(n12188), .Z(
        \SUBBYTES[5].a/w894 ) );
  XOR \SUBBYTES[5].a/U4178  ( .A(\w1[5][96] ), .B(\SUBBYTES[5].a/w894 ), .Z(
        \SUBBYTES[5].a/w781 ) );
  XOR \SUBBYTES[5].a/U4177  ( .A(\w1[5][96] ), .B(n11861), .Z(
        \SUBBYTES[5].a/w782 ) );
  XOR \SUBBYTES[5].a/U4176  ( .A(\w1[5][102] ), .B(\w1[5][101] ), .Z(n11861)
         );
  XOR \SUBBYTES[5].a/U4175  ( .A(\w1[5][101] ), .B(n12188), .Z(
        \SUBBYTES[5].a/w912 ) );
  XOR \SUBBYTES[5].a/U4174  ( .A(n11863), .B(n11862), .Z(\SUBBYTES[5].a/w905 )
         );
  XOR \SUBBYTES[5].a/U4173  ( .A(\w1[5][99] ), .B(\w1[5][97] ), .Z(n11862) );
  XOR \SUBBYTES[5].a/U4172  ( .A(\w1[5][103] ), .B(\w1[5][100] ), .Z(n11863)
         );
  XOR \SUBBYTES[5].a/U4171  ( .A(\w1[5][96] ), .B(\SUBBYTES[5].a/w905 ), .Z(
        \SUBBYTES[5].a/w784 ) );
  XOR \SUBBYTES[5].a/U4170  ( .A(n11865), .B(n11864), .Z(\SUBBYTES[5].a/w892 )
         );
  XOR \SUBBYTES[5].a/U4169  ( .A(\SUBBYTES[5].a/w853 ), .B(n1024), .Z(n11864)
         );
  XOR \SUBBYTES[5].a/U4168  ( .A(\SUBBYTES[5].a/w846 ), .B(
        \SUBBYTES[5].a/w849 ), .Z(n11865) );
  XOR \SUBBYTES[5].a/U4167  ( .A(n11867), .B(n11866), .Z(\SUBBYTES[5].a/w893 )
         );
  XOR \SUBBYTES[5].a/U4166  ( .A(\SUBBYTES[5].a/w853 ), .B(n10959), .Z(n11866)
         );
  XOR \SUBBYTES[5].a/U4165  ( .A(\SUBBYTES[5].a/w846 ), .B(n10958), .Z(n11867)
         );
  XOR \SUBBYTES[5].a/U4164  ( .A(\SUBBYTES[5].a/w905 ), .B(n11868), .Z(
        \SUBBYTES[5].a/w895 ) );
  XOR \SUBBYTES[5].a/U4163  ( .A(\w1[5][102] ), .B(\w1[5][101] ), .Z(n11868)
         );
  XOR \SUBBYTES[5].a/U4162  ( .A(n11870), .B(n11869), .Z(\SUBBYTES[5].a/w896 )
         );
  XOR \SUBBYTES[5].a/U4161  ( .A(n10959), .B(n1024), .Z(n11869) );
  XOR \SUBBYTES[5].a/U4160  ( .A(n10958), .B(\SUBBYTES[5].a/w849 ), .Z(n11870)
         );
  XOR \SUBBYTES[5].a/U4159  ( .A(\w1[5][103] ), .B(\w1[5][98] ), .Z(n12194) );
  XOR \SUBBYTES[5].a/U4158  ( .A(n12194), .B(n11871), .Z(\SUBBYTES[5].a/w897 )
         );
  XOR \SUBBYTES[5].a/U4157  ( .A(\w1[5][101] ), .B(\w1[5][100] ), .Z(n11871)
         );
  XOR \SUBBYTES[5].a/U4156  ( .A(\w1[5][103] ), .B(\SUBBYTES[5].a/w782 ), .Z(
        \SUBBYTES[5].a/w785 ) );
  XOR \SUBBYTES[5].a/U4155  ( .A(\w1[5][97] ), .B(\SUBBYTES[5].a/w782 ), .Z(
        \SUBBYTES[5].a/w786 ) );
  XOR \SUBBYTES[5].a/U4154  ( .A(\w1[5][100] ), .B(\SUBBYTES[5].a/w782 ), .Z(
        \SUBBYTES[5].a/w787 ) );
  XOR \SUBBYTES[5].a/U4153  ( .A(\SUBBYTES[5].a/w786 ), .B(n12194), .Z(
        \SUBBYTES[5].a/w788 ) );
  XOR \SUBBYTES[5].a/U4152  ( .A(n12194), .B(n11872), .Z(\SUBBYTES[5].a/w873 )
         );
  XOR \SUBBYTES[5].a/U4151  ( .A(\w1[5][100] ), .B(\w1[5][97] ), .Z(n11872) );
  XOR \SUBBYTES[5].a/U4150  ( .A(n11874), .B(n11873), .Z(n12191) );
  XOR \SUBBYTES[5].a/U4149  ( .A(\w1[5][100] ), .B(n11875), .Z(n11873) );
  XOR \SUBBYTES[5].a/U4148  ( .A(\SUBBYTES[5].a/w838 ), .B(\w1[5][102] ), .Z(
        n11874) );
  XOR \SUBBYTES[5].a/U4147  ( .A(\SUBBYTES[5].a/w812 ), .B(
        \SUBBYTES[5].a/w819 ), .Z(n11875) );
  XOR \SUBBYTES[5].a/U4146  ( .A(n11877), .B(n11876), .Z(n12189) );
  XOR \SUBBYTES[5].a/U4145  ( .A(\w1[5][97] ), .B(n11878), .Z(n11876) );
  XOR \SUBBYTES[5].a/U4144  ( .A(\SUBBYTES[5].a/w837 ), .B(\w1[5][101] ), .Z(
        n11877) );
  XOR \SUBBYTES[5].a/U4143  ( .A(\SUBBYTES[5].a/w813 ), .B(
        \SUBBYTES[5].a/w820 ), .Z(n11878) );
  XOR \SUBBYTES[5].a/U4142  ( .A(n12191), .B(n12189), .Z(\SUBBYTES[5].a/w843 )
         );
  XOR \SUBBYTES[5].a/U4141  ( .A(\w1[5][101] ), .B(n11879), .Z(n12192) );
  XOR \SUBBYTES[5].a/U4140  ( .A(\SUBBYTES[5].a/w805 ), .B(
        \SUBBYTES[5].a/w815 ), .Z(n11879) );
  XOR \SUBBYTES[5].a/U4139  ( .A(n11881), .B(n11880), .Z(\SUBBYTES[5].a/w830 )
         );
  XOR \SUBBYTES[5].a/U4138  ( .A(n12192), .B(n11882), .Z(n11880) );
  XOR \SUBBYTES[5].a/U4137  ( .A(\w1[5][100] ), .B(\SUBBYTES[5].a/w894 ), .Z(
        n11881) );
  XOR \SUBBYTES[5].a/U4136  ( .A(\SUBBYTES[5].a/w807 ), .B(
        \SUBBYTES[5].a/w812 ), .Z(n11882) );
  XOR \SUBBYTES[5].a/U4135  ( .A(n11884), .B(n11883), .Z(n12190) );
  XOR \SUBBYTES[5].a/U4134  ( .A(\SUBBYTES[5].a/w840 ), .B(\w1[5][103] ), .Z(
        n11883) );
  XOR \SUBBYTES[5].a/U4133  ( .A(\SUBBYTES[5].a/w815 ), .B(
        \SUBBYTES[5].a/w822 ), .Z(n11884) );
  XOR \SUBBYTES[5].a/U4132  ( .A(n12189), .B(n12190), .Z(\SUBBYTES[5].a/w842 )
         );
  XOR \SUBBYTES[5].a/U4131  ( .A(\w1[5][99] ), .B(n11885), .Z(n12193) );
  XOR \SUBBYTES[5].a/U4130  ( .A(\SUBBYTES[5].a/w804 ), .B(
        \SUBBYTES[5].a/w807 ), .Z(n11885) );
  XOR \SUBBYTES[5].a/U4129  ( .A(n11887), .B(n11886), .Z(\SUBBYTES[5].a/w831 )
         );
  XOR \SUBBYTES[5].a/U4128  ( .A(n12193), .B(n11888), .Z(n11886) );
  XOR \SUBBYTES[5].a/U4127  ( .A(\w1[5][102] ), .B(\SUBBYTES[5].a/w873 ), .Z(
        n11887) );
  XOR \SUBBYTES[5].a/U4126  ( .A(\SUBBYTES[5].a/w812 ), .B(
        \SUBBYTES[5].a/w813 ), .Z(n11888) );
  XOR \SUBBYTES[5].a/U4125  ( .A(n12191), .B(n12190), .Z(\SUBBYTES[5].a/w851 )
         );
  XOR \SUBBYTES[5].a/U4124  ( .A(n11890), .B(n11889), .Z(\SUBBYTES[5].a/w852 )
         );
  XOR \SUBBYTES[5].a/U4123  ( .A(\w1[5][103] ), .B(n12192), .Z(n11889) );
  XOR \SUBBYTES[5].a/U4122  ( .A(\SUBBYTES[5].a/w804 ), .B(
        \SUBBYTES[5].a/w813 ), .Z(n11890) );
  XOR \SUBBYTES[5].a/U4121  ( .A(n11892), .B(n11891), .Z(\SUBBYTES[5].a/w828 )
         );
  XOR \SUBBYTES[5].a/U4120  ( .A(n11894), .B(n11893), .Z(n11891) );
  XOR \SUBBYTES[5].a/U4119  ( .A(\w1[5][103] ), .B(\SUBBYTES[5].a/w912 ), .Z(
        n11892) );
  XOR \SUBBYTES[5].a/U4118  ( .A(\SUBBYTES[5].a/w819 ), .B(
        \SUBBYTES[5].a/w822 ), .Z(n11893) );
  XOR \SUBBYTES[5].a/U4117  ( .A(\SUBBYTES[5].a/w805 ), .B(
        \SUBBYTES[5].a/w807 ), .Z(n11894) );
  XOR \SUBBYTES[5].a/U4116  ( .A(n11896), .B(n11895), .Z(\SUBBYTES[5].a/w829 )
         );
  XOR \SUBBYTES[5].a/U4115  ( .A(n12193), .B(n11897), .Z(n11895) );
  XOR \SUBBYTES[5].a/U4114  ( .A(\w1[5][101] ), .B(n12194), .Z(n11896) );
  XOR \SUBBYTES[5].a/U4113  ( .A(\SUBBYTES[5].a/w819 ), .B(
        \SUBBYTES[5].a/w820 ), .Z(n11897) );
  XOR \SUBBYTES[5].a/U4112  ( .A(n11899), .B(n11898), .Z(\SUBBYTES[5].a/w845 )
         );
  XOR \SUBBYTES[5].a/U4111  ( .A(\w1[5][97] ), .B(n11900), .Z(n11898) );
  XOR \SUBBYTES[5].a/U4110  ( .A(\SUBBYTES[5].a/w820 ), .B(
        \SUBBYTES[5].a/w822 ), .Z(n11899) );
  XOR \SUBBYTES[5].a/U4109  ( .A(\SUBBYTES[5].a/w804 ), .B(
        \SUBBYTES[5].a/w805 ), .Z(n11900) );
  XOR \SUBBYTES[5].a/U4108  ( .A(\w1[5][105] ), .B(n11901), .Z(n12195) );
  XOR \SUBBYTES[5].a/U4107  ( .A(\w1[5][107] ), .B(\w1[5][106] ), .Z(n11901)
         );
  XOR \SUBBYTES[5].a/U4106  ( .A(\w1[5][110] ), .B(n12195), .Z(
        \SUBBYTES[5].a/w687 ) );
  XOR \SUBBYTES[5].a/U4105  ( .A(\w1[5][104] ), .B(\SUBBYTES[5].a/w687 ), .Z(
        \SUBBYTES[5].a/w574 ) );
  XOR \SUBBYTES[5].a/U4104  ( .A(\w1[5][104] ), .B(n11902), .Z(
        \SUBBYTES[5].a/w575 ) );
  XOR \SUBBYTES[5].a/U4103  ( .A(\w1[5][110] ), .B(\w1[5][109] ), .Z(n11902)
         );
  XOR \SUBBYTES[5].a/U4102  ( .A(\w1[5][109] ), .B(n12195), .Z(
        \SUBBYTES[5].a/w705 ) );
  XOR \SUBBYTES[5].a/U4101  ( .A(n11904), .B(n11903), .Z(\SUBBYTES[5].a/w698 )
         );
  XOR \SUBBYTES[5].a/U4100  ( .A(\w1[5][107] ), .B(\w1[5][105] ), .Z(n11903)
         );
  XOR \SUBBYTES[5].a/U4099  ( .A(\w1[5][111] ), .B(\w1[5][108] ), .Z(n11904)
         );
  XOR \SUBBYTES[5].a/U4098  ( .A(\w1[5][104] ), .B(\SUBBYTES[5].a/w698 ), .Z(
        \SUBBYTES[5].a/w577 ) );
  XOR \SUBBYTES[5].a/U4097  ( .A(n11906), .B(n11905), .Z(\SUBBYTES[5].a/w685 )
         );
  XOR \SUBBYTES[5].a/U4096  ( .A(\SUBBYTES[5].a/w646 ), .B(n1023), .Z(n11905)
         );
  XOR \SUBBYTES[5].a/U4095  ( .A(\SUBBYTES[5].a/w639 ), .B(
        \SUBBYTES[5].a/w642 ), .Z(n11906) );
  XOR \SUBBYTES[5].a/U4094  ( .A(n11908), .B(n11907), .Z(\SUBBYTES[5].a/w686 )
         );
  XOR \SUBBYTES[5].a/U4093  ( .A(\SUBBYTES[5].a/w646 ), .B(n10957), .Z(n11907)
         );
  XOR \SUBBYTES[5].a/U4092  ( .A(\SUBBYTES[5].a/w639 ), .B(n10956), .Z(n11908)
         );
  XOR \SUBBYTES[5].a/U4091  ( .A(\SUBBYTES[5].a/w698 ), .B(n11909), .Z(
        \SUBBYTES[5].a/w688 ) );
  XOR \SUBBYTES[5].a/U4090  ( .A(\w1[5][110] ), .B(\w1[5][109] ), .Z(n11909)
         );
  XOR \SUBBYTES[5].a/U4089  ( .A(n11911), .B(n11910), .Z(\SUBBYTES[5].a/w689 )
         );
  XOR \SUBBYTES[5].a/U4088  ( .A(n10957), .B(n1023), .Z(n11910) );
  XOR \SUBBYTES[5].a/U4087  ( .A(n10956), .B(\SUBBYTES[5].a/w642 ), .Z(n11911)
         );
  XOR \SUBBYTES[5].a/U4086  ( .A(\w1[5][111] ), .B(\w1[5][106] ), .Z(n12201)
         );
  XOR \SUBBYTES[5].a/U4085  ( .A(n12201), .B(n11912), .Z(\SUBBYTES[5].a/w690 )
         );
  XOR \SUBBYTES[5].a/U4084  ( .A(\w1[5][109] ), .B(\w1[5][108] ), .Z(n11912)
         );
  XOR \SUBBYTES[5].a/U4083  ( .A(\w1[5][111] ), .B(\SUBBYTES[5].a/w575 ), .Z(
        \SUBBYTES[5].a/w578 ) );
  XOR \SUBBYTES[5].a/U4082  ( .A(\w1[5][105] ), .B(\SUBBYTES[5].a/w575 ), .Z(
        \SUBBYTES[5].a/w579 ) );
  XOR \SUBBYTES[5].a/U4081  ( .A(\w1[5][108] ), .B(\SUBBYTES[5].a/w575 ), .Z(
        \SUBBYTES[5].a/w580 ) );
  XOR \SUBBYTES[5].a/U4080  ( .A(\SUBBYTES[5].a/w579 ), .B(n12201), .Z(
        \SUBBYTES[5].a/w581 ) );
  XOR \SUBBYTES[5].a/U4079  ( .A(n12201), .B(n11913), .Z(\SUBBYTES[5].a/w666 )
         );
  XOR \SUBBYTES[5].a/U4078  ( .A(\w1[5][108] ), .B(\w1[5][105] ), .Z(n11913)
         );
  XOR \SUBBYTES[5].a/U4077  ( .A(n11915), .B(n11914), .Z(n12198) );
  XOR \SUBBYTES[5].a/U4076  ( .A(\w1[5][108] ), .B(n11916), .Z(n11914) );
  XOR \SUBBYTES[5].a/U4075  ( .A(\SUBBYTES[5].a/w631 ), .B(\w1[5][110] ), .Z(
        n11915) );
  XOR \SUBBYTES[5].a/U4074  ( .A(\SUBBYTES[5].a/w605 ), .B(
        \SUBBYTES[5].a/w612 ), .Z(n11916) );
  XOR \SUBBYTES[5].a/U4073  ( .A(n11918), .B(n11917), .Z(n12196) );
  XOR \SUBBYTES[5].a/U4072  ( .A(\w1[5][105] ), .B(n11919), .Z(n11917) );
  XOR \SUBBYTES[5].a/U4071  ( .A(\SUBBYTES[5].a/w630 ), .B(\w1[5][109] ), .Z(
        n11918) );
  XOR \SUBBYTES[5].a/U4070  ( .A(\SUBBYTES[5].a/w606 ), .B(
        \SUBBYTES[5].a/w613 ), .Z(n11919) );
  XOR \SUBBYTES[5].a/U4069  ( .A(n12198), .B(n12196), .Z(\SUBBYTES[5].a/w636 )
         );
  XOR \SUBBYTES[5].a/U4068  ( .A(\w1[5][109] ), .B(n11920), .Z(n12199) );
  XOR \SUBBYTES[5].a/U4067  ( .A(\SUBBYTES[5].a/w598 ), .B(
        \SUBBYTES[5].a/w608 ), .Z(n11920) );
  XOR \SUBBYTES[5].a/U4066  ( .A(n11922), .B(n11921), .Z(\SUBBYTES[5].a/w623 )
         );
  XOR \SUBBYTES[5].a/U4065  ( .A(n12199), .B(n11923), .Z(n11921) );
  XOR \SUBBYTES[5].a/U4064  ( .A(\w1[5][108] ), .B(\SUBBYTES[5].a/w687 ), .Z(
        n11922) );
  XOR \SUBBYTES[5].a/U4063  ( .A(\SUBBYTES[5].a/w600 ), .B(
        \SUBBYTES[5].a/w605 ), .Z(n11923) );
  XOR \SUBBYTES[5].a/U4062  ( .A(n11925), .B(n11924), .Z(n12197) );
  XOR \SUBBYTES[5].a/U4061  ( .A(\SUBBYTES[5].a/w633 ), .B(\w1[5][111] ), .Z(
        n11924) );
  XOR \SUBBYTES[5].a/U4060  ( .A(\SUBBYTES[5].a/w608 ), .B(
        \SUBBYTES[5].a/w615 ), .Z(n11925) );
  XOR \SUBBYTES[5].a/U4059  ( .A(n12196), .B(n12197), .Z(\SUBBYTES[5].a/w635 )
         );
  XOR \SUBBYTES[5].a/U4058  ( .A(\w1[5][107] ), .B(n11926), .Z(n12200) );
  XOR \SUBBYTES[5].a/U4057  ( .A(\SUBBYTES[5].a/w597 ), .B(
        \SUBBYTES[5].a/w600 ), .Z(n11926) );
  XOR \SUBBYTES[5].a/U4056  ( .A(n11928), .B(n11927), .Z(\SUBBYTES[5].a/w624 )
         );
  XOR \SUBBYTES[5].a/U4055  ( .A(n12200), .B(n11929), .Z(n11927) );
  XOR \SUBBYTES[5].a/U4054  ( .A(\w1[5][110] ), .B(\SUBBYTES[5].a/w666 ), .Z(
        n11928) );
  XOR \SUBBYTES[5].a/U4053  ( .A(\SUBBYTES[5].a/w605 ), .B(
        \SUBBYTES[5].a/w606 ), .Z(n11929) );
  XOR \SUBBYTES[5].a/U4052  ( .A(n12198), .B(n12197), .Z(\SUBBYTES[5].a/w644 )
         );
  XOR \SUBBYTES[5].a/U4051  ( .A(n11931), .B(n11930), .Z(\SUBBYTES[5].a/w645 )
         );
  XOR \SUBBYTES[5].a/U4050  ( .A(\w1[5][111] ), .B(n12199), .Z(n11930) );
  XOR \SUBBYTES[5].a/U4049  ( .A(\SUBBYTES[5].a/w597 ), .B(
        \SUBBYTES[5].a/w606 ), .Z(n11931) );
  XOR \SUBBYTES[5].a/U4048  ( .A(n11933), .B(n11932), .Z(\SUBBYTES[5].a/w621 )
         );
  XOR \SUBBYTES[5].a/U4047  ( .A(n11935), .B(n11934), .Z(n11932) );
  XOR \SUBBYTES[5].a/U4046  ( .A(\w1[5][111] ), .B(\SUBBYTES[5].a/w705 ), .Z(
        n11933) );
  XOR \SUBBYTES[5].a/U4045  ( .A(\SUBBYTES[5].a/w612 ), .B(
        \SUBBYTES[5].a/w615 ), .Z(n11934) );
  XOR \SUBBYTES[5].a/U4044  ( .A(\SUBBYTES[5].a/w598 ), .B(
        \SUBBYTES[5].a/w600 ), .Z(n11935) );
  XOR \SUBBYTES[5].a/U4043  ( .A(n11937), .B(n11936), .Z(\SUBBYTES[5].a/w622 )
         );
  XOR \SUBBYTES[5].a/U4042  ( .A(n12200), .B(n11938), .Z(n11936) );
  XOR \SUBBYTES[5].a/U4041  ( .A(\w1[5][109] ), .B(n12201), .Z(n11937) );
  XOR \SUBBYTES[5].a/U4040  ( .A(\SUBBYTES[5].a/w612 ), .B(
        \SUBBYTES[5].a/w613 ), .Z(n11938) );
  XOR \SUBBYTES[5].a/U4039  ( .A(n11940), .B(n11939), .Z(\SUBBYTES[5].a/w638 )
         );
  XOR \SUBBYTES[5].a/U4038  ( .A(\w1[5][105] ), .B(n11941), .Z(n11939) );
  XOR \SUBBYTES[5].a/U4037  ( .A(\SUBBYTES[5].a/w613 ), .B(
        \SUBBYTES[5].a/w615 ), .Z(n11940) );
  XOR \SUBBYTES[5].a/U4036  ( .A(\SUBBYTES[5].a/w597 ), .B(
        \SUBBYTES[5].a/w598 ), .Z(n11941) );
  XOR \SUBBYTES[5].a/U4035  ( .A(\w1[5][113] ), .B(n11942), .Z(n12202) );
  XOR \SUBBYTES[5].a/U4034  ( .A(\w1[5][115] ), .B(\w1[5][114] ), .Z(n11942)
         );
  XOR \SUBBYTES[5].a/U4033  ( .A(\w1[5][118] ), .B(n12202), .Z(
        \SUBBYTES[5].a/w480 ) );
  XOR \SUBBYTES[5].a/U4032  ( .A(\w1[5][112] ), .B(\SUBBYTES[5].a/w480 ), .Z(
        \SUBBYTES[5].a/w367 ) );
  XOR \SUBBYTES[5].a/U4031  ( .A(\w1[5][112] ), .B(n11943), .Z(
        \SUBBYTES[5].a/w368 ) );
  XOR \SUBBYTES[5].a/U4030  ( .A(\w1[5][118] ), .B(\w1[5][117] ), .Z(n11943)
         );
  XOR \SUBBYTES[5].a/U4029  ( .A(\w1[5][117] ), .B(n12202), .Z(
        \SUBBYTES[5].a/w498 ) );
  XOR \SUBBYTES[5].a/U4028  ( .A(n11945), .B(n11944), .Z(\SUBBYTES[5].a/w491 )
         );
  XOR \SUBBYTES[5].a/U4027  ( .A(\w1[5][115] ), .B(\w1[5][113] ), .Z(n11944)
         );
  XOR \SUBBYTES[5].a/U4026  ( .A(\w1[5][119] ), .B(\w1[5][116] ), .Z(n11945)
         );
  XOR \SUBBYTES[5].a/U4025  ( .A(\w1[5][112] ), .B(\SUBBYTES[5].a/w491 ), .Z(
        \SUBBYTES[5].a/w370 ) );
  XOR \SUBBYTES[5].a/U4024  ( .A(n11947), .B(n11946), .Z(\SUBBYTES[5].a/w478 )
         );
  XOR \SUBBYTES[5].a/U4023  ( .A(\SUBBYTES[5].a/w439 ), .B(n1022), .Z(n11946)
         );
  XOR \SUBBYTES[5].a/U4022  ( .A(\SUBBYTES[5].a/w432 ), .B(
        \SUBBYTES[5].a/w435 ), .Z(n11947) );
  XOR \SUBBYTES[5].a/U4021  ( .A(n11949), .B(n11948), .Z(\SUBBYTES[5].a/w479 )
         );
  XOR \SUBBYTES[5].a/U4020  ( .A(\SUBBYTES[5].a/w439 ), .B(n10955), .Z(n11948)
         );
  XOR \SUBBYTES[5].a/U4019  ( .A(\SUBBYTES[5].a/w432 ), .B(n10954), .Z(n11949)
         );
  XOR \SUBBYTES[5].a/U4018  ( .A(\SUBBYTES[5].a/w491 ), .B(n11950), .Z(
        \SUBBYTES[5].a/w481 ) );
  XOR \SUBBYTES[5].a/U4017  ( .A(\w1[5][118] ), .B(\w1[5][117] ), .Z(n11950)
         );
  XOR \SUBBYTES[5].a/U4016  ( .A(n11952), .B(n11951), .Z(\SUBBYTES[5].a/w482 )
         );
  XOR \SUBBYTES[5].a/U4015  ( .A(n10955), .B(n1022), .Z(n11951) );
  XOR \SUBBYTES[5].a/U4014  ( .A(n10954), .B(\SUBBYTES[5].a/w435 ), .Z(n11952)
         );
  XOR \SUBBYTES[5].a/U4013  ( .A(\w1[5][119] ), .B(\w1[5][114] ), .Z(n12208)
         );
  XOR \SUBBYTES[5].a/U4012  ( .A(n12208), .B(n11953), .Z(\SUBBYTES[5].a/w483 )
         );
  XOR \SUBBYTES[5].a/U4011  ( .A(\w1[5][117] ), .B(\w1[5][116] ), .Z(n11953)
         );
  XOR \SUBBYTES[5].a/U4010  ( .A(\w1[5][119] ), .B(\SUBBYTES[5].a/w368 ), .Z(
        \SUBBYTES[5].a/w371 ) );
  XOR \SUBBYTES[5].a/U4009  ( .A(\w1[5][113] ), .B(\SUBBYTES[5].a/w368 ), .Z(
        \SUBBYTES[5].a/w372 ) );
  XOR \SUBBYTES[5].a/U4008  ( .A(\w1[5][116] ), .B(\SUBBYTES[5].a/w368 ), .Z(
        \SUBBYTES[5].a/w373 ) );
  XOR \SUBBYTES[5].a/U4007  ( .A(\SUBBYTES[5].a/w372 ), .B(n12208), .Z(
        \SUBBYTES[5].a/w374 ) );
  XOR \SUBBYTES[5].a/U4006  ( .A(n12208), .B(n11954), .Z(\SUBBYTES[5].a/w459 )
         );
  XOR \SUBBYTES[5].a/U4005  ( .A(\w1[5][116] ), .B(\w1[5][113] ), .Z(n11954)
         );
  XOR \SUBBYTES[5].a/U4004  ( .A(n11956), .B(n11955), .Z(n12205) );
  XOR \SUBBYTES[5].a/U4003  ( .A(\w1[5][116] ), .B(n11957), .Z(n11955) );
  XOR \SUBBYTES[5].a/U4002  ( .A(\SUBBYTES[5].a/w424 ), .B(\w1[5][118] ), .Z(
        n11956) );
  XOR \SUBBYTES[5].a/U4001  ( .A(\SUBBYTES[5].a/w398 ), .B(
        \SUBBYTES[5].a/w405 ), .Z(n11957) );
  XOR \SUBBYTES[5].a/U4000  ( .A(n11959), .B(n11958), .Z(n12203) );
  XOR \SUBBYTES[5].a/U3999  ( .A(\w1[5][113] ), .B(n11960), .Z(n11958) );
  XOR \SUBBYTES[5].a/U3998  ( .A(\SUBBYTES[5].a/w423 ), .B(\w1[5][117] ), .Z(
        n11959) );
  XOR \SUBBYTES[5].a/U3997  ( .A(\SUBBYTES[5].a/w399 ), .B(
        \SUBBYTES[5].a/w406 ), .Z(n11960) );
  XOR \SUBBYTES[5].a/U3996  ( .A(n12205), .B(n12203), .Z(\SUBBYTES[5].a/w429 )
         );
  XOR \SUBBYTES[5].a/U3995  ( .A(\w1[5][117] ), .B(n11961), .Z(n12206) );
  XOR \SUBBYTES[5].a/U3994  ( .A(\SUBBYTES[5].a/w391 ), .B(
        \SUBBYTES[5].a/w401 ), .Z(n11961) );
  XOR \SUBBYTES[5].a/U3993  ( .A(n11963), .B(n11962), .Z(\SUBBYTES[5].a/w416 )
         );
  XOR \SUBBYTES[5].a/U3992  ( .A(n12206), .B(n11964), .Z(n11962) );
  XOR \SUBBYTES[5].a/U3991  ( .A(\w1[5][116] ), .B(\SUBBYTES[5].a/w480 ), .Z(
        n11963) );
  XOR \SUBBYTES[5].a/U3990  ( .A(\SUBBYTES[5].a/w393 ), .B(
        \SUBBYTES[5].a/w398 ), .Z(n11964) );
  XOR \SUBBYTES[5].a/U3989  ( .A(n11966), .B(n11965), .Z(n12204) );
  XOR \SUBBYTES[5].a/U3988  ( .A(\SUBBYTES[5].a/w426 ), .B(\w1[5][119] ), .Z(
        n11965) );
  XOR \SUBBYTES[5].a/U3987  ( .A(\SUBBYTES[5].a/w401 ), .B(
        \SUBBYTES[5].a/w408 ), .Z(n11966) );
  XOR \SUBBYTES[5].a/U3986  ( .A(n12203), .B(n12204), .Z(\SUBBYTES[5].a/w428 )
         );
  XOR \SUBBYTES[5].a/U3985  ( .A(\w1[5][115] ), .B(n11967), .Z(n12207) );
  XOR \SUBBYTES[5].a/U3984  ( .A(\SUBBYTES[5].a/w390 ), .B(
        \SUBBYTES[5].a/w393 ), .Z(n11967) );
  XOR \SUBBYTES[5].a/U3983  ( .A(n11969), .B(n11968), .Z(\SUBBYTES[5].a/w417 )
         );
  XOR \SUBBYTES[5].a/U3982  ( .A(n12207), .B(n11970), .Z(n11968) );
  XOR \SUBBYTES[5].a/U3981  ( .A(\w1[5][118] ), .B(\SUBBYTES[5].a/w459 ), .Z(
        n11969) );
  XOR \SUBBYTES[5].a/U3980  ( .A(\SUBBYTES[5].a/w398 ), .B(
        \SUBBYTES[5].a/w399 ), .Z(n11970) );
  XOR \SUBBYTES[5].a/U3979  ( .A(n12205), .B(n12204), .Z(\SUBBYTES[5].a/w437 )
         );
  XOR \SUBBYTES[5].a/U3978  ( .A(n11972), .B(n11971), .Z(\SUBBYTES[5].a/w438 )
         );
  XOR \SUBBYTES[5].a/U3977  ( .A(\w1[5][119] ), .B(n12206), .Z(n11971) );
  XOR \SUBBYTES[5].a/U3976  ( .A(\SUBBYTES[5].a/w390 ), .B(
        \SUBBYTES[5].a/w399 ), .Z(n11972) );
  XOR \SUBBYTES[5].a/U3975  ( .A(n11974), .B(n11973), .Z(\SUBBYTES[5].a/w414 )
         );
  XOR \SUBBYTES[5].a/U3974  ( .A(n11976), .B(n11975), .Z(n11973) );
  XOR \SUBBYTES[5].a/U3973  ( .A(\w1[5][119] ), .B(\SUBBYTES[5].a/w498 ), .Z(
        n11974) );
  XOR \SUBBYTES[5].a/U3972  ( .A(\SUBBYTES[5].a/w405 ), .B(
        \SUBBYTES[5].a/w408 ), .Z(n11975) );
  XOR \SUBBYTES[5].a/U3971  ( .A(\SUBBYTES[5].a/w391 ), .B(
        \SUBBYTES[5].a/w393 ), .Z(n11976) );
  XOR \SUBBYTES[5].a/U3970  ( .A(n11978), .B(n11977), .Z(\SUBBYTES[5].a/w415 )
         );
  XOR \SUBBYTES[5].a/U3969  ( .A(n12207), .B(n11979), .Z(n11977) );
  XOR \SUBBYTES[5].a/U3968  ( .A(\w1[5][117] ), .B(n12208), .Z(n11978) );
  XOR \SUBBYTES[5].a/U3967  ( .A(\SUBBYTES[5].a/w405 ), .B(
        \SUBBYTES[5].a/w406 ), .Z(n11979) );
  XOR \SUBBYTES[5].a/U3966  ( .A(n11981), .B(n11980), .Z(\SUBBYTES[5].a/w431 )
         );
  XOR \SUBBYTES[5].a/U3965  ( .A(\w1[5][113] ), .B(n11982), .Z(n11980) );
  XOR \SUBBYTES[5].a/U3964  ( .A(\SUBBYTES[5].a/w406 ), .B(
        \SUBBYTES[5].a/w408 ), .Z(n11981) );
  XOR \SUBBYTES[5].a/U3963  ( .A(\SUBBYTES[5].a/w390 ), .B(
        \SUBBYTES[5].a/w391 ), .Z(n11982) );
  XOR \SUBBYTES[5].a/U3962  ( .A(\w1[5][121] ), .B(n11983), .Z(n12209) );
  XOR \SUBBYTES[5].a/U3961  ( .A(\w1[5][123] ), .B(\w1[5][122] ), .Z(n11983)
         );
  XOR \SUBBYTES[5].a/U3960  ( .A(\w1[5][126] ), .B(n12209), .Z(
        \SUBBYTES[5].a/w273 ) );
  XOR \SUBBYTES[5].a/U3959  ( .A(\w1[5][120] ), .B(\SUBBYTES[5].a/w273 ), .Z(
        \SUBBYTES[5].a/w160 ) );
  XOR \SUBBYTES[5].a/U3958  ( .A(\w1[5][120] ), .B(n11984), .Z(
        \SUBBYTES[5].a/w161 ) );
  XOR \SUBBYTES[5].a/U3957  ( .A(\w1[5][126] ), .B(\w1[5][125] ), .Z(n11984)
         );
  XOR \SUBBYTES[5].a/U3956  ( .A(\w1[5][125] ), .B(n12209), .Z(
        \SUBBYTES[5].a/w291 ) );
  XOR \SUBBYTES[5].a/U3955  ( .A(n11986), .B(n11985), .Z(\SUBBYTES[5].a/w284 )
         );
  XOR \SUBBYTES[5].a/U3954  ( .A(\w1[5][123] ), .B(\w1[5][121] ), .Z(n11985)
         );
  XOR \SUBBYTES[5].a/U3953  ( .A(\w1[5][127] ), .B(\w1[5][124] ), .Z(n11986)
         );
  XOR \SUBBYTES[5].a/U3952  ( .A(\w1[5][120] ), .B(\SUBBYTES[5].a/w284 ), .Z(
        \SUBBYTES[5].a/w163 ) );
  XOR \SUBBYTES[5].a/U3951  ( .A(n11988), .B(n11987), .Z(\SUBBYTES[5].a/w271 )
         );
  XOR \SUBBYTES[5].a/U3950  ( .A(\SUBBYTES[5].a/w232 ), .B(n1021), .Z(n11987)
         );
  XOR \SUBBYTES[5].a/U3949  ( .A(\SUBBYTES[5].a/w225 ), .B(
        \SUBBYTES[5].a/w228 ), .Z(n11988) );
  XOR \SUBBYTES[5].a/U3948  ( .A(n11990), .B(n11989), .Z(\SUBBYTES[5].a/w272 )
         );
  XOR \SUBBYTES[5].a/U3947  ( .A(\SUBBYTES[5].a/w232 ), .B(n10953), .Z(n11989)
         );
  XOR \SUBBYTES[5].a/U3946  ( .A(\SUBBYTES[5].a/w225 ), .B(n10952), .Z(n11990)
         );
  XOR \SUBBYTES[5].a/U3945  ( .A(\SUBBYTES[5].a/w284 ), .B(n11991), .Z(
        \SUBBYTES[5].a/w274 ) );
  XOR \SUBBYTES[5].a/U3944  ( .A(\w1[5][126] ), .B(\w1[5][125] ), .Z(n11991)
         );
  XOR \SUBBYTES[5].a/U3943  ( .A(n11993), .B(n11992), .Z(\SUBBYTES[5].a/w275 )
         );
  XOR \SUBBYTES[5].a/U3942  ( .A(n10953), .B(n1021), .Z(n11992) );
  XOR \SUBBYTES[5].a/U3941  ( .A(n10952), .B(\SUBBYTES[5].a/w228 ), .Z(n11993)
         );
  XOR \SUBBYTES[5].a/U3940  ( .A(\w1[5][127] ), .B(\w1[5][122] ), .Z(n12215)
         );
  XOR \SUBBYTES[5].a/U3939  ( .A(n12215), .B(n11994), .Z(\SUBBYTES[5].a/w276 )
         );
  XOR \SUBBYTES[5].a/U3938  ( .A(\w1[5][125] ), .B(\w1[5][124] ), .Z(n11994)
         );
  XOR \SUBBYTES[5].a/U3937  ( .A(\w1[5][127] ), .B(\SUBBYTES[5].a/w161 ), .Z(
        \SUBBYTES[5].a/w164 ) );
  XOR \SUBBYTES[5].a/U3936  ( .A(\w1[5][121] ), .B(\SUBBYTES[5].a/w161 ), .Z(
        \SUBBYTES[5].a/w165 ) );
  XOR \SUBBYTES[5].a/U3935  ( .A(\w1[5][124] ), .B(\SUBBYTES[5].a/w161 ), .Z(
        \SUBBYTES[5].a/w166 ) );
  XOR \SUBBYTES[5].a/U3934  ( .A(\SUBBYTES[5].a/w165 ), .B(n12215), .Z(
        \SUBBYTES[5].a/w167 ) );
  XOR \SUBBYTES[5].a/U3933  ( .A(n12215), .B(n11995), .Z(\SUBBYTES[5].a/w252 )
         );
  XOR \SUBBYTES[5].a/U3932  ( .A(\w1[5][124] ), .B(\w1[5][121] ), .Z(n11995)
         );
  XOR \SUBBYTES[5].a/U3931  ( .A(n11997), .B(n11996), .Z(n12212) );
  XOR \SUBBYTES[5].a/U3930  ( .A(\w1[5][124] ), .B(n11998), .Z(n11996) );
  XOR \SUBBYTES[5].a/U3929  ( .A(\SUBBYTES[5].a/w217 ), .B(\w1[5][126] ), .Z(
        n11997) );
  XOR \SUBBYTES[5].a/U3928  ( .A(\SUBBYTES[5].a/w191 ), .B(
        \SUBBYTES[5].a/w198 ), .Z(n11998) );
  XOR \SUBBYTES[5].a/U3927  ( .A(n12000), .B(n11999), .Z(n12210) );
  XOR \SUBBYTES[5].a/U3926  ( .A(\w1[5][121] ), .B(n12001), .Z(n11999) );
  XOR \SUBBYTES[5].a/U3925  ( .A(\SUBBYTES[5].a/w216 ), .B(\w1[5][125] ), .Z(
        n12000) );
  XOR \SUBBYTES[5].a/U3924  ( .A(\SUBBYTES[5].a/w192 ), .B(
        \SUBBYTES[5].a/w199 ), .Z(n12001) );
  XOR \SUBBYTES[5].a/U3923  ( .A(n12212), .B(n12210), .Z(\SUBBYTES[5].a/w222 )
         );
  XOR \SUBBYTES[5].a/U3922  ( .A(\w1[5][125] ), .B(n12002), .Z(n12213) );
  XOR \SUBBYTES[5].a/U3921  ( .A(\SUBBYTES[5].a/w184 ), .B(
        \SUBBYTES[5].a/w194 ), .Z(n12002) );
  XOR \SUBBYTES[5].a/U3920  ( .A(n12004), .B(n12003), .Z(\SUBBYTES[5].a/w209 )
         );
  XOR \SUBBYTES[5].a/U3919  ( .A(n12213), .B(n12005), .Z(n12003) );
  XOR \SUBBYTES[5].a/U3918  ( .A(\w1[5][124] ), .B(\SUBBYTES[5].a/w273 ), .Z(
        n12004) );
  XOR \SUBBYTES[5].a/U3917  ( .A(\SUBBYTES[5].a/w186 ), .B(
        \SUBBYTES[5].a/w191 ), .Z(n12005) );
  XOR \SUBBYTES[5].a/U3916  ( .A(n12007), .B(n12006), .Z(n12211) );
  XOR \SUBBYTES[5].a/U3915  ( .A(\SUBBYTES[5].a/w219 ), .B(\w1[5][127] ), .Z(
        n12006) );
  XOR \SUBBYTES[5].a/U3914  ( .A(\SUBBYTES[5].a/w194 ), .B(
        \SUBBYTES[5].a/w201 ), .Z(n12007) );
  XOR \SUBBYTES[5].a/U3913  ( .A(n12210), .B(n12211), .Z(\SUBBYTES[5].a/w221 )
         );
  XOR \SUBBYTES[5].a/U3912  ( .A(\w1[5][123] ), .B(n12008), .Z(n12214) );
  XOR \SUBBYTES[5].a/U3911  ( .A(\SUBBYTES[5].a/w183 ), .B(
        \SUBBYTES[5].a/w186 ), .Z(n12008) );
  XOR \SUBBYTES[5].a/U3910  ( .A(n12010), .B(n12009), .Z(\SUBBYTES[5].a/w210 )
         );
  XOR \SUBBYTES[5].a/U3909  ( .A(n12214), .B(n12011), .Z(n12009) );
  XOR \SUBBYTES[5].a/U3908  ( .A(\w1[5][126] ), .B(\SUBBYTES[5].a/w252 ), .Z(
        n12010) );
  XOR \SUBBYTES[5].a/U3907  ( .A(\SUBBYTES[5].a/w191 ), .B(
        \SUBBYTES[5].a/w192 ), .Z(n12011) );
  XOR \SUBBYTES[5].a/U3906  ( .A(n12212), .B(n12211), .Z(\SUBBYTES[5].a/w230 )
         );
  XOR \SUBBYTES[5].a/U3905  ( .A(n12013), .B(n12012), .Z(\SUBBYTES[5].a/w231 )
         );
  XOR \SUBBYTES[5].a/U3904  ( .A(\w1[5][127] ), .B(n12213), .Z(n12012) );
  XOR \SUBBYTES[5].a/U3903  ( .A(\SUBBYTES[5].a/w183 ), .B(
        \SUBBYTES[5].a/w192 ), .Z(n12013) );
  XOR \SUBBYTES[5].a/U3902  ( .A(n12015), .B(n12014), .Z(\SUBBYTES[5].a/w207 )
         );
  XOR \SUBBYTES[5].a/U3901  ( .A(n12017), .B(n12016), .Z(n12014) );
  XOR \SUBBYTES[5].a/U3900  ( .A(\w1[5][127] ), .B(\SUBBYTES[5].a/w291 ), .Z(
        n12015) );
  XOR \SUBBYTES[5].a/U3899  ( .A(\SUBBYTES[5].a/w198 ), .B(
        \SUBBYTES[5].a/w201 ), .Z(n12016) );
  XOR \SUBBYTES[5].a/U3898  ( .A(\SUBBYTES[5].a/w184 ), .B(
        \SUBBYTES[5].a/w186 ), .Z(n12017) );
  XOR \SUBBYTES[5].a/U3897  ( .A(n12019), .B(n12018), .Z(\SUBBYTES[5].a/w208 )
         );
  XOR \SUBBYTES[5].a/U3896  ( .A(n12214), .B(n12020), .Z(n12018) );
  XOR \SUBBYTES[5].a/U3895  ( .A(\w1[5][125] ), .B(n12215), .Z(n12019) );
  XOR \SUBBYTES[5].a/U3894  ( .A(\SUBBYTES[5].a/w198 ), .B(
        \SUBBYTES[5].a/w199 ), .Z(n12020) );
  XOR \SUBBYTES[5].a/U3893  ( .A(n12022), .B(n12021), .Z(\SUBBYTES[5].a/w224 )
         );
  XOR \SUBBYTES[5].a/U3892  ( .A(\w1[5][121] ), .B(n12023), .Z(n12021) );
  XOR \SUBBYTES[5].a/U3891  ( .A(\SUBBYTES[5].a/w199 ), .B(
        \SUBBYTES[5].a/w201 ), .Z(n12022) );
  XOR \SUBBYTES[5].a/U3890  ( .A(\SUBBYTES[5].a/w183 ), .B(
        \SUBBYTES[5].a/w184 ), .Z(n12023) );
  XOR \SUBBYTES[4].a/U5649  ( .A(\SUBBYTES[4].a/w3390 ), .B(
        \SUBBYTES[4].a/w3391 ), .Z(n10745) );
  XOR \SUBBYTES[4].a/U5648  ( .A(n10745), .B(n9704), .Z(n10744) );
  XOR \SUBBYTES[4].a/U5647  ( .A(\SUBBYTES[4].a/w3383 ), .B(
        \SUBBYTES[4].a/w3400 ), .Z(n9704) );
  XOR \SUBBYTES[4].a/U5645  ( .A(\SUBBYTES[4].a/w3382 ), .B(
        \SUBBYTES[4].a/w3397 ), .Z(n9705) );
  XOR \SUBBYTES[4].a/U5644  ( .A(n10745), .B(n9706), .Z(n10936) );
  XOR \SUBBYTES[4].a/U5643  ( .A(\SUBBYTES[4].a/w3397 ), .B(
        \SUBBYTES[4].a/w3398 ), .Z(n9706) );
  XOR \SUBBYTES[4].a/U5642  ( .A(\SUBBYTES[4].a/w3359 ), .B(n9707), .Z(n10747)
         );
  XOR \SUBBYTES[4].a/U5641  ( .A(\SUBBYTES[4].a/w3350 ), .B(
        \SUBBYTES[4].a/w3351 ), .Z(n9707) );
  XOR \SUBBYTES[4].a/U5639  ( .A(\SUBBYTES[4].a/w3361 ), .B(n10936), .Z(n9708)
         );
  XOR \SUBBYTES[4].a/U5638  ( .A(n9710), .B(n9709), .Z(n10748) );
  XOR \SUBBYTES[4].a/U5637  ( .A(n9712), .B(n9711), .Z(n9709) );
  XOR \SUBBYTES[4].a/U5636  ( .A(\SUBBYTES[4].a/w3397 ), .B(
        \SUBBYTES[4].a/w3398 ), .Z(n9710) );
  XOR \SUBBYTES[4].a/U5635  ( .A(\SUBBYTES[4].a/w3361 ), .B(
        \SUBBYTES[4].a/w3385 ), .Z(n9711) );
  XOR \SUBBYTES[4].a/U5634  ( .A(\SUBBYTES[4].a/w3350 ), .B(
        \SUBBYTES[4].a/w3359 ), .Z(n9712) );
  XOR \SUBBYTES[4].a/U5633  ( .A(\SUBBYTES[4].a/w3382 ), .B(n9713), .Z(n10746)
         );
  XOR \SUBBYTES[4].a/U5632  ( .A(\SUBBYTES[4].a/w3365 ), .B(
        \SUBBYTES[4].a/w3368 ), .Z(n9713) );
  XOR \SUBBYTES[4].a/U5630  ( .A(\SUBBYTES[4].a/w3353 ), .B(n10748), .Z(n9714)
         );
  XOR \SUBBYTES[4].a/U5628  ( .A(\SUBBYTES[4].a/w3385 ), .B(
        \SUBBYTES[4].a/w3398 ), .Z(n9715) );
  XOR \SUBBYTES[4].a/U5626  ( .A(n9719), .B(n9718), .Z(n9716) );
  XOR \SUBBYTES[4].a/U5625  ( .A(n9721), .B(n9720), .Z(n9717) );
  XOR \SUBBYTES[4].a/U5624  ( .A(\SUBBYTES[4].a/w3397 ), .B(
        \SUBBYTES[4].a/w3400 ), .Z(n9718) );
  XOR \SUBBYTES[4].a/U5623  ( .A(\SUBBYTES[4].a/w3390 ), .B(
        \SUBBYTES[4].a/w3393 ), .Z(n9719) );
  XOR \SUBBYTES[4].a/U5622  ( .A(\SUBBYTES[4].a/w3365 ), .B(
        \SUBBYTES[4].a/w3366 ), .Z(n9720) );
  XOR \SUBBYTES[4].a/U5621  ( .A(\SUBBYTES[4].a/w3350 ), .B(
        \SUBBYTES[4].a/w3353 ), .Z(n9721) );
  XOR \SUBBYTES[4].a/U5619  ( .A(n10745), .B(n9724), .Z(n9722) );
  XOR \SUBBYTES[4].a/U5618  ( .A(n10747), .B(n10746), .Z(n9723) );
  XOR \SUBBYTES[4].a/U5617  ( .A(\SUBBYTES[4].a/w3358 ), .B(
        \SUBBYTES[4].a/w3385 ), .Z(n9724) );
  XOR \SUBBYTES[4].a/U5615  ( .A(n10748), .B(n9727), .Z(n9725) );
  XOR \SUBBYTES[4].a/U5614  ( .A(\SUBBYTES[4].a/w3391 ), .B(
        \SUBBYTES[4].a/w3393 ), .Z(n9726) );
  XOR \SUBBYTES[4].a/U5613  ( .A(\SUBBYTES[4].a/w3351 ), .B(
        \SUBBYTES[4].a/w3383 ), .Z(n9727) );
  XOR \SUBBYTES[4].a/U5612  ( .A(\SUBBYTES[4].a/w3183 ), .B(
        \SUBBYTES[4].a/w3184 ), .Z(n10750) );
  XOR \SUBBYTES[4].a/U5611  ( .A(n10750), .B(n9728), .Z(n10749) );
  XOR \SUBBYTES[4].a/U5610  ( .A(\SUBBYTES[4].a/w3176 ), .B(
        \SUBBYTES[4].a/w3193 ), .Z(n9728) );
  XOR \SUBBYTES[4].a/U5608  ( .A(\SUBBYTES[4].a/w3175 ), .B(
        \SUBBYTES[4].a/w3190 ), .Z(n9729) );
  XOR \SUBBYTES[4].a/U5607  ( .A(n10750), .B(n9730), .Z(n10937) );
  XOR \SUBBYTES[4].a/U5606  ( .A(\SUBBYTES[4].a/w3190 ), .B(
        \SUBBYTES[4].a/w3191 ), .Z(n9730) );
  XOR \SUBBYTES[4].a/U5605  ( .A(\SUBBYTES[4].a/w3152 ), .B(n9731), .Z(n10752)
         );
  XOR \SUBBYTES[4].a/U5604  ( .A(\SUBBYTES[4].a/w3143 ), .B(
        \SUBBYTES[4].a/w3144 ), .Z(n9731) );
  XOR \SUBBYTES[4].a/U5602  ( .A(\SUBBYTES[4].a/w3154 ), .B(n10937), .Z(n9732)
         );
  XOR \SUBBYTES[4].a/U5601  ( .A(n9734), .B(n9733), .Z(n10753) );
  XOR \SUBBYTES[4].a/U5600  ( .A(n9736), .B(n9735), .Z(n9733) );
  XOR \SUBBYTES[4].a/U5599  ( .A(\SUBBYTES[4].a/w3190 ), .B(
        \SUBBYTES[4].a/w3191 ), .Z(n9734) );
  XOR \SUBBYTES[4].a/U5598  ( .A(\SUBBYTES[4].a/w3154 ), .B(
        \SUBBYTES[4].a/w3178 ), .Z(n9735) );
  XOR \SUBBYTES[4].a/U5597  ( .A(\SUBBYTES[4].a/w3143 ), .B(
        \SUBBYTES[4].a/w3152 ), .Z(n9736) );
  XOR \SUBBYTES[4].a/U5596  ( .A(\SUBBYTES[4].a/w3175 ), .B(n9737), .Z(n10751)
         );
  XOR \SUBBYTES[4].a/U5595  ( .A(\SUBBYTES[4].a/w3158 ), .B(
        \SUBBYTES[4].a/w3161 ), .Z(n9737) );
  XOR \SUBBYTES[4].a/U5593  ( .A(\SUBBYTES[4].a/w3146 ), .B(n10753), .Z(n9738)
         );
  XOR \SUBBYTES[4].a/U5591  ( .A(\SUBBYTES[4].a/w3178 ), .B(
        \SUBBYTES[4].a/w3191 ), .Z(n9739) );
  XOR \SUBBYTES[4].a/U5589  ( .A(n9743), .B(n9742), .Z(n9740) );
  XOR \SUBBYTES[4].a/U5588  ( .A(n9745), .B(n9744), .Z(n9741) );
  XOR \SUBBYTES[4].a/U5587  ( .A(\SUBBYTES[4].a/w3190 ), .B(
        \SUBBYTES[4].a/w3193 ), .Z(n9742) );
  XOR \SUBBYTES[4].a/U5586  ( .A(\SUBBYTES[4].a/w3183 ), .B(
        \SUBBYTES[4].a/w3186 ), .Z(n9743) );
  XOR \SUBBYTES[4].a/U5585  ( .A(\SUBBYTES[4].a/w3158 ), .B(
        \SUBBYTES[4].a/w3159 ), .Z(n9744) );
  XOR \SUBBYTES[4].a/U5584  ( .A(\SUBBYTES[4].a/w3143 ), .B(
        \SUBBYTES[4].a/w3146 ), .Z(n9745) );
  XOR \SUBBYTES[4].a/U5582  ( .A(n10750), .B(n9748), .Z(n9746) );
  XOR \SUBBYTES[4].a/U5581  ( .A(n10752), .B(n10751), .Z(n9747) );
  XOR \SUBBYTES[4].a/U5580  ( .A(\SUBBYTES[4].a/w3151 ), .B(
        \SUBBYTES[4].a/w3178 ), .Z(n9748) );
  XOR \SUBBYTES[4].a/U5578  ( .A(n10753), .B(n9751), .Z(n9749) );
  XOR \SUBBYTES[4].a/U5577  ( .A(\SUBBYTES[4].a/w3184 ), .B(
        \SUBBYTES[4].a/w3186 ), .Z(n9750) );
  XOR \SUBBYTES[4].a/U5576  ( .A(\SUBBYTES[4].a/w3144 ), .B(
        \SUBBYTES[4].a/w3176 ), .Z(n9751) );
  XOR \SUBBYTES[4].a/U5575  ( .A(\SUBBYTES[4].a/w2976 ), .B(
        \SUBBYTES[4].a/w2977 ), .Z(n10755) );
  XOR \SUBBYTES[4].a/U5574  ( .A(n10755), .B(n9752), .Z(n10754) );
  XOR \SUBBYTES[4].a/U5573  ( .A(\SUBBYTES[4].a/w2969 ), .B(
        \SUBBYTES[4].a/w2986 ), .Z(n9752) );
  XOR \SUBBYTES[4].a/U5571  ( .A(\SUBBYTES[4].a/w2968 ), .B(
        \SUBBYTES[4].a/w2983 ), .Z(n9753) );
  XOR \SUBBYTES[4].a/U5570  ( .A(n10755), .B(n9754), .Z(n10938) );
  XOR \SUBBYTES[4].a/U5569  ( .A(\SUBBYTES[4].a/w2983 ), .B(
        \SUBBYTES[4].a/w2984 ), .Z(n9754) );
  XOR \SUBBYTES[4].a/U5568  ( .A(\SUBBYTES[4].a/w2945 ), .B(n9755), .Z(n10757)
         );
  XOR \SUBBYTES[4].a/U5567  ( .A(\SUBBYTES[4].a/w2936 ), .B(
        \SUBBYTES[4].a/w2937 ), .Z(n9755) );
  XOR \SUBBYTES[4].a/U5565  ( .A(\SUBBYTES[4].a/w2947 ), .B(n10938), .Z(n9756)
         );
  XOR \SUBBYTES[4].a/U5564  ( .A(n9758), .B(n9757), .Z(n10758) );
  XOR \SUBBYTES[4].a/U5563  ( .A(n9760), .B(n9759), .Z(n9757) );
  XOR \SUBBYTES[4].a/U5562  ( .A(\SUBBYTES[4].a/w2983 ), .B(
        \SUBBYTES[4].a/w2984 ), .Z(n9758) );
  XOR \SUBBYTES[4].a/U5561  ( .A(\SUBBYTES[4].a/w2947 ), .B(
        \SUBBYTES[4].a/w2971 ), .Z(n9759) );
  XOR \SUBBYTES[4].a/U5560  ( .A(\SUBBYTES[4].a/w2936 ), .B(
        \SUBBYTES[4].a/w2945 ), .Z(n9760) );
  XOR \SUBBYTES[4].a/U5559  ( .A(\SUBBYTES[4].a/w2968 ), .B(n9761), .Z(n10756)
         );
  XOR \SUBBYTES[4].a/U5558  ( .A(\SUBBYTES[4].a/w2951 ), .B(
        \SUBBYTES[4].a/w2954 ), .Z(n9761) );
  XOR \SUBBYTES[4].a/U5556  ( .A(\SUBBYTES[4].a/w2939 ), .B(n10758), .Z(n9762)
         );
  XOR \SUBBYTES[4].a/U5554  ( .A(\SUBBYTES[4].a/w2971 ), .B(
        \SUBBYTES[4].a/w2984 ), .Z(n9763) );
  XOR \SUBBYTES[4].a/U5552  ( .A(n9767), .B(n9766), .Z(n9764) );
  XOR \SUBBYTES[4].a/U5551  ( .A(n9769), .B(n9768), .Z(n9765) );
  XOR \SUBBYTES[4].a/U5550  ( .A(\SUBBYTES[4].a/w2983 ), .B(
        \SUBBYTES[4].a/w2986 ), .Z(n9766) );
  XOR \SUBBYTES[4].a/U5549  ( .A(\SUBBYTES[4].a/w2976 ), .B(
        \SUBBYTES[4].a/w2979 ), .Z(n9767) );
  XOR \SUBBYTES[4].a/U5548  ( .A(\SUBBYTES[4].a/w2951 ), .B(
        \SUBBYTES[4].a/w2952 ), .Z(n9768) );
  XOR \SUBBYTES[4].a/U5547  ( .A(\SUBBYTES[4].a/w2936 ), .B(
        \SUBBYTES[4].a/w2939 ), .Z(n9769) );
  XOR \SUBBYTES[4].a/U5545  ( .A(n10755), .B(n9772), .Z(n9770) );
  XOR \SUBBYTES[4].a/U5544  ( .A(n10757), .B(n10756), .Z(n9771) );
  XOR \SUBBYTES[4].a/U5543  ( .A(\SUBBYTES[4].a/w2944 ), .B(
        \SUBBYTES[4].a/w2971 ), .Z(n9772) );
  XOR \SUBBYTES[4].a/U5541  ( .A(n10758), .B(n9775), .Z(n9773) );
  XOR \SUBBYTES[4].a/U5540  ( .A(\SUBBYTES[4].a/w2977 ), .B(
        \SUBBYTES[4].a/w2979 ), .Z(n9774) );
  XOR \SUBBYTES[4].a/U5539  ( .A(\SUBBYTES[4].a/w2937 ), .B(
        \SUBBYTES[4].a/w2969 ), .Z(n9775) );
  XOR \SUBBYTES[4].a/U5538  ( .A(\SUBBYTES[4].a/w2769 ), .B(
        \SUBBYTES[4].a/w2770 ), .Z(n10760) );
  XOR \SUBBYTES[4].a/U5537  ( .A(n10760), .B(n9776), .Z(n10759) );
  XOR \SUBBYTES[4].a/U5536  ( .A(\SUBBYTES[4].a/w2762 ), .B(
        \SUBBYTES[4].a/w2779 ), .Z(n9776) );
  XOR \SUBBYTES[4].a/U5534  ( .A(\SUBBYTES[4].a/w2761 ), .B(
        \SUBBYTES[4].a/w2776 ), .Z(n9777) );
  XOR \SUBBYTES[4].a/U5533  ( .A(n10760), .B(n9778), .Z(n10939) );
  XOR \SUBBYTES[4].a/U5532  ( .A(\SUBBYTES[4].a/w2776 ), .B(
        \SUBBYTES[4].a/w2777 ), .Z(n9778) );
  XOR \SUBBYTES[4].a/U5531  ( .A(\SUBBYTES[4].a/w2738 ), .B(n9779), .Z(n10762)
         );
  XOR \SUBBYTES[4].a/U5530  ( .A(\SUBBYTES[4].a/w2729 ), .B(
        \SUBBYTES[4].a/w2730 ), .Z(n9779) );
  XOR \SUBBYTES[4].a/U5528  ( .A(\SUBBYTES[4].a/w2740 ), .B(n10939), .Z(n9780)
         );
  XOR \SUBBYTES[4].a/U5527  ( .A(n9782), .B(n9781), .Z(n10763) );
  XOR \SUBBYTES[4].a/U5526  ( .A(n9784), .B(n9783), .Z(n9781) );
  XOR \SUBBYTES[4].a/U5525  ( .A(\SUBBYTES[4].a/w2776 ), .B(
        \SUBBYTES[4].a/w2777 ), .Z(n9782) );
  XOR \SUBBYTES[4].a/U5524  ( .A(\SUBBYTES[4].a/w2740 ), .B(
        \SUBBYTES[4].a/w2764 ), .Z(n9783) );
  XOR \SUBBYTES[4].a/U5523  ( .A(\SUBBYTES[4].a/w2729 ), .B(
        \SUBBYTES[4].a/w2738 ), .Z(n9784) );
  XOR \SUBBYTES[4].a/U5522  ( .A(\SUBBYTES[4].a/w2761 ), .B(n9785), .Z(n10761)
         );
  XOR \SUBBYTES[4].a/U5521  ( .A(\SUBBYTES[4].a/w2744 ), .B(
        \SUBBYTES[4].a/w2747 ), .Z(n9785) );
  XOR \SUBBYTES[4].a/U5519  ( .A(\SUBBYTES[4].a/w2732 ), .B(n10763), .Z(n9786)
         );
  XOR \SUBBYTES[4].a/U5517  ( .A(\SUBBYTES[4].a/w2764 ), .B(
        \SUBBYTES[4].a/w2777 ), .Z(n9787) );
  XOR \SUBBYTES[4].a/U5515  ( .A(n9791), .B(n9790), .Z(n9788) );
  XOR \SUBBYTES[4].a/U5514  ( .A(n9793), .B(n9792), .Z(n9789) );
  XOR \SUBBYTES[4].a/U5513  ( .A(\SUBBYTES[4].a/w2776 ), .B(
        \SUBBYTES[4].a/w2779 ), .Z(n9790) );
  XOR \SUBBYTES[4].a/U5512  ( .A(\SUBBYTES[4].a/w2769 ), .B(
        \SUBBYTES[4].a/w2772 ), .Z(n9791) );
  XOR \SUBBYTES[4].a/U5511  ( .A(\SUBBYTES[4].a/w2744 ), .B(
        \SUBBYTES[4].a/w2745 ), .Z(n9792) );
  XOR \SUBBYTES[4].a/U5510  ( .A(\SUBBYTES[4].a/w2729 ), .B(
        \SUBBYTES[4].a/w2732 ), .Z(n9793) );
  XOR \SUBBYTES[4].a/U5508  ( .A(n10760), .B(n9796), .Z(n9794) );
  XOR \SUBBYTES[4].a/U5507  ( .A(n10762), .B(n10761), .Z(n9795) );
  XOR \SUBBYTES[4].a/U5506  ( .A(\SUBBYTES[4].a/w2737 ), .B(
        \SUBBYTES[4].a/w2764 ), .Z(n9796) );
  XOR \SUBBYTES[4].a/U5504  ( .A(n10763), .B(n9799), .Z(n9797) );
  XOR \SUBBYTES[4].a/U5503  ( .A(\SUBBYTES[4].a/w2770 ), .B(
        \SUBBYTES[4].a/w2772 ), .Z(n9798) );
  XOR \SUBBYTES[4].a/U5502  ( .A(\SUBBYTES[4].a/w2730 ), .B(
        \SUBBYTES[4].a/w2762 ), .Z(n9799) );
  XOR \SUBBYTES[4].a/U5501  ( .A(\SUBBYTES[4].a/w2562 ), .B(
        \SUBBYTES[4].a/w2563 ), .Z(n10765) );
  XOR \SUBBYTES[4].a/U5500  ( .A(n10765), .B(n9800), .Z(n10764) );
  XOR \SUBBYTES[4].a/U5499  ( .A(\SUBBYTES[4].a/w2555 ), .B(
        \SUBBYTES[4].a/w2572 ), .Z(n9800) );
  XOR \SUBBYTES[4].a/U5497  ( .A(\SUBBYTES[4].a/w2554 ), .B(
        \SUBBYTES[4].a/w2569 ), .Z(n9801) );
  XOR \SUBBYTES[4].a/U5496  ( .A(n10765), .B(n9802), .Z(n10940) );
  XOR \SUBBYTES[4].a/U5495  ( .A(\SUBBYTES[4].a/w2569 ), .B(
        \SUBBYTES[4].a/w2570 ), .Z(n9802) );
  XOR \SUBBYTES[4].a/U5494  ( .A(\SUBBYTES[4].a/w2531 ), .B(n9803), .Z(n10767)
         );
  XOR \SUBBYTES[4].a/U5493  ( .A(\SUBBYTES[4].a/w2522 ), .B(
        \SUBBYTES[4].a/w2523 ), .Z(n9803) );
  XOR \SUBBYTES[4].a/U5491  ( .A(\SUBBYTES[4].a/w2533 ), .B(n10940), .Z(n9804)
         );
  XOR \SUBBYTES[4].a/U5490  ( .A(n9806), .B(n9805), .Z(n10768) );
  XOR \SUBBYTES[4].a/U5489  ( .A(n9808), .B(n9807), .Z(n9805) );
  XOR \SUBBYTES[4].a/U5488  ( .A(\SUBBYTES[4].a/w2569 ), .B(
        \SUBBYTES[4].a/w2570 ), .Z(n9806) );
  XOR \SUBBYTES[4].a/U5487  ( .A(\SUBBYTES[4].a/w2533 ), .B(
        \SUBBYTES[4].a/w2557 ), .Z(n9807) );
  XOR \SUBBYTES[4].a/U5486  ( .A(\SUBBYTES[4].a/w2522 ), .B(
        \SUBBYTES[4].a/w2531 ), .Z(n9808) );
  XOR \SUBBYTES[4].a/U5485  ( .A(\SUBBYTES[4].a/w2554 ), .B(n9809), .Z(n10766)
         );
  XOR \SUBBYTES[4].a/U5484  ( .A(\SUBBYTES[4].a/w2537 ), .B(
        \SUBBYTES[4].a/w2540 ), .Z(n9809) );
  XOR \SUBBYTES[4].a/U5482  ( .A(\SUBBYTES[4].a/w2525 ), .B(n10768), .Z(n9810)
         );
  XOR \SUBBYTES[4].a/U5480  ( .A(\SUBBYTES[4].a/w2557 ), .B(
        \SUBBYTES[4].a/w2570 ), .Z(n9811) );
  XOR \SUBBYTES[4].a/U5478  ( .A(n9815), .B(n9814), .Z(n9812) );
  XOR \SUBBYTES[4].a/U5477  ( .A(n9817), .B(n9816), .Z(n9813) );
  XOR \SUBBYTES[4].a/U5476  ( .A(\SUBBYTES[4].a/w2569 ), .B(
        \SUBBYTES[4].a/w2572 ), .Z(n9814) );
  XOR \SUBBYTES[4].a/U5475  ( .A(\SUBBYTES[4].a/w2562 ), .B(
        \SUBBYTES[4].a/w2565 ), .Z(n9815) );
  XOR \SUBBYTES[4].a/U5474  ( .A(\SUBBYTES[4].a/w2537 ), .B(
        \SUBBYTES[4].a/w2538 ), .Z(n9816) );
  XOR \SUBBYTES[4].a/U5473  ( .A(\SUBBYTES[4].a/w2522 ), .B(
        \SUBBYTES[4].a/w2525 ), .Z(n9817) );
  XOR \SUBBYTES[4].a/U5471  ( .A(n10765), .B(n9820), .Z(n9818) );
  XOR \SUBBYTES[4].a/U5470  ( .A(n10767), .B(n10766), .Z(n9819) );
  XOR \SUBBYTES[4].a/U5469  ( .A(\SUBBYTES[4].a/w2530 ), .B(
        \SUBBYTES[4].a/w2557 ), .Z(n9820) );
  XOR \SUBBYTES[4].a/U5467  ( .A(n10768), .B(n9823), .Z(n9821) );
  XOR \SUBBYTES[4].a/U5466  ( .A(\SUBBYTES[4].a/w2563 ), .B(
        \SUBBYTES[4].a/w2565 ), .Z(n9822) );
  XOR \SUBBYTES[4].a/U5465  ( .A(\SUBBYTES[4].a/w2523 ), .B(
        \SUBBYTES[4].a/w2555 ), .Z(n9823) );
  XOR \SUBBYTES[4].a/U5464  ( .A(\SUBBYTES[4].a/w2355 ), .B(
        \SUBBYTES[4].a/w2356 ), .Z(n10770) );
  XOR \SUBBYTES[4].a/U5463  ( .A(n10770), .B(n9824), .Z(n10769) );
  XOR \SUBBYTES[4].a/U5462  ( .A(\SUBBYTES[4].a/w2348 ), .B(
        \SUBBYTES[4].a/w2365 ), .Z(n9824) );
  XOR \SUBBYTES[4].a/U5460  ( .A(\SUBBYTES[4].a/w2347 ), .B(
        \SUBBYTES[4].a/w2362 ), .Z(n9825) );
  XOR \SUBBYTES[4].a/U5459  ( .A(n10770), .B(n9826), .Z(n10941) );
  XOR \SUBBYTES[4].a/U5458  ( .A(\SUBBYTES[4].a/w2362 ), .B(
        \SUBBYTES[4].a/w2363 ), .Z(n9826) );
  XOR \SUBBYTES[4].a/U5457  ( .A(\SUBBYTES[4].a/w2324 ), .B(n9827), .Z(n10772)
         );
  XOR \SUBBYTES[4].a/U5456  ( .A(\SUBBYTES[4].a/w2315 ), .B(
        \SUBBYTES[4].a/w2316 ), .Z(n9827) );
  XOR \SUBBYTES[4].a/U5454  ( .A(\SUBBYTES[4].a/w2326 ), .B(n10941), .Z(n9828)
         );
  XOR \SUBBYTES[4].a/U5453  ( .A(n9830), .B(n9829), .Z(n10773) );
  XOR \SUBBYTES[4].a/U5452  ( .A(n9832), .B(n9831), .Z(n9829) );
  XOR \SUBBYTES[4].a/U5451  ( .A(\SUBBYTES[4].a/w2362 ), .B(
        \SUBBYTES[4].a/w2363 ), .Z(n9830) );
  XOR \SUBBYTES[4].a/U5450  ( .A(\SUBBYTES[4].a/w2326 ), .B(
        \SUBBYTES[4].a/w2350 ), .Z(n9831) );
  XOR \SUBBYTES[4].a/U5449  ( .A(\SUBBYTES[4].a/w2315 ), .B(
        \SUBBYTES[4].a/w2324 ), .Z(n9832) );
  XOR \SUBBYTES[4].a/U5448  ( .A(\SUBBYTES[4].a/w2347 ), .B(n9833), .Z(n10771)
         );
  XOR \SUBBYTES[4].a/U5447  ( .A(\SUBBYTES[4].a/w2330 ), .B(
        \SUBBYTES[4].a/w2333 ), .Z(n9833) );
  XOR \SUBBYTES[4].a/U5445  ( .A(\SUBBYTES[4].a/w2318 ), .B(n10773), .Z(n9834)
         );
  XOR \SUBBYTES[4].a/U5443  ( .A(\SUBBYTES[4].a/w2350 ), .B(
        \SUBBYTES[4].a/w2363 ), .Z(n9835) );
  XOR \SUBBYTES[4].a/U5441  ( .A(n9839), .B(n9838), .Z(n9836) );
  XOR \SUBBYTES[4].a/U5440  ( .A(n9841), .B(n9840), .Z(n9837) );
  XOR \SUBBYTES[4].a/U5439  ( .A(\SUBBYTES[4].a/w2362 ), .B(
        \SUBBYTES[4].a/w2365 ), .Z(n9838) );
  XOR \SUBBYTES[4].a/U5438  ( .A(\SUBBYTES[4].a/w2355 ), .B(
        \SUBBYTES[4].a/w2358 ), .Z(n9839) );
  XOR \SUBBYTES[4].a/U5437  ( .A(\SUBBYTES[4].a/w2330 ), .B(
        \SUBBYTES[4].a/w2331 ), .Z(n9840) );
  XOR \SUBBYTES[4].a/U5436  ( .A(\SUBBYTES[4].a/w2315 ), .B(
        \SUBBYTES[4].a/w2318 ), .Z(n9841) );
  XOR \SUBBYTES[4].a/U5434  ( .A(n10770), .B(n9844), .Z(n9842) );
  XOR \SUBBYTES[4].a/U5433  ( .A(n10772), .B(n10771), .Z(n9843) );
  XOR \SUBBYTES[4].a/U5432  ( .A(\SUBBYTES[4].a/w2323 ), .B(
        \SUBBYTES[4].a/w2350 ), .Z(n9844) );
  XOR \SUBBYTES[4].a/U5430  ( .A(n10773), .B(n9847), .Z(n9845) );
  XOR \SUBBYTES[4].a/U5429  ( .A(\SUBBYTES[4].a/w2356 ), .B(
        \SUBBYTES[4].a/w2358 ), .Z(n9846) );
  XOR \SUBBYTES[4].a/U5428  ( .A(\SUBBYTES[4].a/w2316 ), .B(
        \SUBBYTES[4].a/w2348 ), .Z(n9847) );
  XOR \SUBBYTES[4].a/U5427  ( .A(\SUBBYTES[4].a/w2148 ), .B(
        \SUBBYTES[4].a/w2149 ), .Z(n10775) );
  XOR \SUBBYTES[4].a/U5426  ( .A(n10775), .B(n9848), .Z(n10774) );
  XOR \SUBBYTES[4].a/U5425  ( .A(\SUBBYTES[4].a/w2141 ), .B(
        \SUBBYTES[4].a/w2158 ), .Z(n9848) );
  XOR \SUBBYTES[4].a/U5423  ( .A(\SUBBYTES[4].a/w2140 ), .B(
        \SUBBYTES[4].a/w2155 ), .Z(n9849) );
  XOR \SUBBYTES[4].a/U5422  ( .A(n10775), .B(n9850), .Z(n10942) );
  XOR \SUBBYTES[4].a/U5421  ( .A(\SUBBYTES[4].a/w2155 ), .B(
        \SUBBYTES[4].a/w2156 ), .Z(n9850) );
  XOR \SUBBYTES[4].a/U5420  ( .A(\SUBBYTES[4].a/w2117 ), .B(n9851), .Z(n10777)
         );
  XOR \SUBBYTES[4].a/U5419  ( .A(\SUBBYTES[4].a/w2108 ), .B(
        \SUBBYTES[4].a/w2109 ), .Z(n9851) );
  XOR \SUBBYTES[4].a/U5417  ( .A(\SUBBYTES[4].a/w2119 ), .B(n10942), .Z(n9852)
         );
  XOR \SUBBYTES[4].a/U5416  ( .A(n9854), .B(n9853), .Z(n10778) );
  XOR \SUBBYTES[4].a/U5415  ( .A(n9856), .B(n9855), .Z(n9853) );
  XOR \SUBBYTES[4].a/U5414  ( .A(\SUBBYTES[4].a/w2155 ), .B(
        \SUBBYTES[4].a/w2156 ), .Z(n9854) );
  XOR \SUBBYTES[4].a/U5413  ( .A(\SUBBYTES[4].a/w2119 ), .B(
        \SUBBYTES[4].a/w2143 ), .Z(n9855) );
  XOR \SUBBYTES[4].a/U5412  ( .A(\SUBBYTES[4].a/w2108 ), .B(
        \SUBBYTES[4].a/w2117 ), .Z(n9856) );
  XOR \SUBBYTES[4].a/U5411  ( .A(\SUBBYTES[4].a/w2140 ), .B(n9857), .Z(n10776)
         );
  XOR \SUBBYTES[4].a/U5410  ( .A(\SUBBYTES[4].a/w2123 ), .B(
        \SUBBYTES[4].a/w2126 ), .Z(n9857) );
  XOR \SUBBYTES[4].a/U5408  ( .A(\SUBBYTES[4].a/w2111 ), .B(n10778), .Z(n9858)
         );
  XOR \SUBBYTES[4].a/U5406  ( .A(\SUBBYTES[4].a/w2143 ), .B(
        \SUBBYTES[4].a/w2156 ), .Z(n9859) );
  XOR \SUBBYTES[4].a/U5404  ( .A(n9863), .B(n9862), .Z(n9860) );
  XOR \SUBBYTES[4].a/U5403  ( .A(n9865), .B(n9864), .Z(n9861) );
  XOR \SUBBYTES[4].a/U5402  ( .A(\SUBBYTES[4].a/w2155 ), .B(
        \SUBBYTES[4].a/w2158 ), .Z(n9862) );
  XOR \SUBBYTES[4].a/U5401  ( .A(\SUBBYTES[4].a/w2148 ), .B(
        \SUBBYTES[4].a/w2151 ), .Z(n9863) );
  XOR \SUBBYTES[4].a/U5400  ( .A(\SUBBYTES[4].a/w2123 ), .B(
        \SUBBYTES[4].a/w2124 ), .Z(n9864) );
  XOR \SUBBYTES[4].a/U5399  ( .A(\SUBBYTES[4].a/w2108 ), .B(
        \SUBBYTES[4].a/w2111 ), .Z(n9865) );
  XOR \SUBBYTES[4].a/U5397  ( .A(n10775), .B(n9868), .Z(n9866) );
  XOR \SUBBYTES[4].a/U5396  ( .A(n10777), .B(n10776), .Z(n9867) );
  XOR \SUBBYTES[4].a/U5395  ( .A(\SUBBYTES[4].a/w2116 ), .B(
        \SUBBYTES[4].a/w2143 ), .Z(n9868) );
  XOR \SUBBYTES[4].a/U5393  ( .A(n10778), .B(n9871), .Z(n9869) );
  XOR \SUBBYTES[4].a/U5392  ( .A(\SUBBYTES[4].a/w2149 ), .B(
        \SUBBYTES[4].a/w2151 ), .Z(n9870) );
  XOR \SUBBYTES[4].a/U5391  ( .A(\SUBBYTES[4].a/w2109 ), .B(
        \SUBBYTES[4].a/w2141 ), .Z(n9871) );
  XOR \SUBBYTES[4].a/U5390  ( .A(\SUBBYTES[4].a/w1941 ), .B(
        \SUBBYTES[4].a/w1942 ), .Z(n10780) );
  XOR \SUBBYTES[4].a/U5389  ( .A(n10780), .B(n9872), .Z(n10779) );
  XOR \SUBBYTES[4].a/U5388  ( .A(\SUBBYTES[4].a/w1934 ), .B(
        \SUBBYTES[4].a/w1951 ), .Z(n9872) );
  XOR \SUBBYTES[4].a/U5386  ( .A(\SUBBYTES[4].a/w1933 ), .B(
        \SUBBYTES[4].a/w1948 ), .Z(n9873) );
  XOR \SUBBYTES[4].a/U5385  ( .A(n10780), .B(n9874), .Z(n10943) );
  XOR \SUBBYTES[4].a/U5384  ( .A(\SUBBYTES[4].a/w1948 ), .B(
        \SUBBYTES[4].a/w1949 ), .Z(n9874) );
  XOR \SUBBYTES[4].a/U5383  ( .A(\SUBBYTES[4].a/w1910 ), .B(n9875), .Z(n10782)
         );
  XOR \SUBBYTES[4].a/U5382  ( .A(\SUBBYTES[4].a/w1901 ), .B(
        \SUBBYTES[4].a/w1902 ), .Z(n9875) );
  XOR \SUBBYTES[4].a/U5380  ( .A(\SUBBYTES[4].a/w1912 ), .B(n10943), .Z(n9876)
         );
  XOR \SUBBYTES[4].a/U5379  ( .A(n9878), .B(n9877), .Z(n10783) );
  XOR \SUBBYTES[4].a/U5378  ( .A(n9880), .B(n9879), .Z(n9877) );
  XOR \SUBBYTES[4].a/U5377  ( .A(\SUBBYTES[4].a/w1948 ), .B(
        \SUBBYTES[4].a/w1949 ), .Z(n9878) );
  XOR \SUBBYTES[4].a/U5376  ( .A(\SUBBYTES[4].a/w1912 ), .B(
        \SUBBYTES[4].a/w1936 ), .Z(n9879) );
  XOR \SUBBYTES[4].a/U5375  ( .A(\SUBBYTES[4].a/w1901 ), .B(
        \SUBBYTES[4].a/w1910 ), .Z(n9880) );
  XOR \SUBBYTES[4].a/U5374  ( .A(\SUBBYTES[4].a/w1933 ), .B(n9881), .Z(n10781)
         );
  XOR \SUBBYTES[4].a/U5373  ( .A(\SUBBYTES[4].a/w1916 ), .B(
        \SUBBYTES[4].a/w1919 ), .Z(n9881) );
  XOR \SUBBYTES[4].a/U5371  ( .A(\SUBBYTES[4].a/w1904 ), .B(n10783), .Z(n9882)
         );
  XOR \SUBBYTES[4].a/U5369  ( .A(\SUBBYTES[4].a/w1936 ), .B(
        \SUBBYTES[4].a/w1949 ), .Z(n9883) );
  XOR \SUBBYTES[4].a/U5367  ( .A(n9887), .B(n9886), .Z(n9884) );
  XOR \SUBBYTES[4].a/U5366  ( .A(n9889), .B(n9888), .Z(n9885) );
  XOR \SUBBYTES[4].a/U5365  ( .A(\SUBBYTES[4].a/w1948 ), .B(
        \SUBBYTES[4].a/w1951 ), .Z(n9886) );
  XOR \SUBBYTES[4].a/U5364  ( .A(\SUBBYTES[4].a/w1941 ), .B(
        \SUBBYTES[4].a/w1944 ), .Z(n9887) );
  XOR \SUBBYTES[4].a/U5363  ( .A(\SUBBYTES[4].a/w1916 ), .B(
        \SUBBYTES[4].a/w1917 ), .Z(n9888) );
  XOR \SUBBYTES[4].a/U5362  ( .A(\SUBBYTES[4].a/w1901 ), .B(
        \SUBBYTES[4].a/w1904 ), .Z(n9889) );
  XOR \SUBBYTES[4].a/U5360  ( .A(n10780), .B(n9892), .Z(n9890) );
  XOR \SUBBYTES[4].a/U5359  ( .A(n10782), .B(n10781), .Z(n9891) );
  XOR \SUBBYTES[4].a/U5358  ( .A(\SUBBYTES[4].a/w1909 ), .B(
        \SUBBYTES[4].a/w1936 ), .Z(n9892) );
  XOR \SUBBYTES[4].a/U5356  ( .A(n10783), .B(n9895), .Z(n9893) );
  XOR \SUBBYTES[4].a/U5355  ( .A(\SUBBYTES[4].a/w1942 ), .B(
        \SUBBYTES[4].a/w1944 ), .Z(n9894) );
  XOR \SUBBYTES[4].a/U5354  ( .A(\SUBBYTES[4].a/w1902 ), .B(
        \SUBBYTES[4].a/w1934 ), .Z(n9895) );
  XOR \SUBBYTES[4].a/U5353  ( .A(\SUBBYTES[4].a/w1734 ), .B(
        \SUBBYTES[4].a/w1735 ), .Z(n10785) );
  XOR \SUBBYTES[4].a/U5352  ( .A(n10785), .B(n9896), .Z(n10784) );
  XOR \SUBBYTES[4].a/U5351  ( .A(\SUBBYTES[4].a/w1727 ), .B(
        \SUBBYTES[4].a/w1744 ), .Z(n9896) );
  XOR \SUBBYTES[4].a/U5349  ( .A(\SUBBYTES[4].a/w1726 ), .B(
        \SUBBYTES[4].a/w1741 ), .Z(n9897) );
  XOR \SUBBYTES[4].a/U5348  ( .A(n10785), .B(n9898), .Z(n10944) );
  XOR \SUBBYTES[4].a/U5347  ( .A(\SUBBYTES[4].a/w1741 ), .B(
        \SUBBYTES[4].a/w1742 ), .Z(n9898) );
  XOR \SUBBYTES[4].a/U5346  ( .A(\SUBBYTES[4].a/w1703 ), .B(n9899), .Z(n10787)
         );
  XOR \SUBBYTES[4].a/U5345  ( .A(\SUBBYTES[4].a/w1694 ), .B(
        \SUBBYTES[4].a/w1695 ), .Z(n9899) );
  XOR \SUBBYTES[4].a/U5343  ( .A(\SUBBYTES[4].a/w1705 ), .B(n10944), .Z(n9900)
         );
  XOR \SUBBYTES[4].a/U5342  ( .A(n9902), .B(n9901), .Z(n10788) );
  XOR \SUBBYTES[4].a/U5341  ( .A(n9904), .B(n9903), .Z(n9901) );
  XOR \SUBBYTES[4].a/U5340  ( .A(\SUBBYTES[4].a/w1741 ), .B(
        \SUBBYTES[4].a/w1742 ), .Z(n9902) );
  XOR \SUBBYTES[4].a/U5339  ( .A(\SUBBYTES[4].a/w1705 ), .B(
        \SUBBYTES[4].a/w1729 ), .Z(n9903) );
  XOR \SUBBYTES[4].a/U5338  ( .A(\SUBBYTES[4].a/w1694 ), .B(
        \SUBBYTES[4].a/w1703 ), .Z(n9904) );
  XOR \SUBBYTES[4].a/U5337  ( .A(\SUBBYTES[4].a/w1726 ), .B(n9905), .Z(n10786)
         );
  XOR \SUBBYTES[4].a/U5336  ( .A(\SUBBYTES[4].a/w1709 ), .B(
        \SUBBYTES[4].a/w1712 ), .Z(n9905) );
  XOR \SUBBYTES[4].a/U5334  ( .A(\SUBBYTES[4].a/w1697 ), .B(n10788), .Z(n9906)
         );
  XOR \SUBBYTES[4].a/U5332  ( .A(\SUBBYTES[4].a/w1729 ), .B(
        \SUBBYTES[4].a/w1742 ), .Z(n9907) );
  XOR \SUBBYTES[4].a/U5330  ( .A(n9911), .B(n9910), .Z(n9908) );
  XOR \SUBBYTES[4].a/U5329  ( .A(n9913), .B(n9912), .Z(n9909) );
  XOR \SUBBYTES[4].a/U5328  ( .A(\SUBBYTES[4].a/w1741 ), .B(
        \SUBBYTES[4].a/w1744 ), .Z(n9910) );
  XOR \SUBBYTES[4].a/U5327  ( .A(\SUBBYTES[4].a/w1734 ), .B(
        \SUBBYTES[4].a/w1737 ), .Z(n9911) );
  XOR \SUBBYTES[4].a/U5326  ( .A(\SUBBYTES[4].a/w1709 ), .B(
        \SUBBYTES[4].a/w1710 ), .Z(n9912) );
  XOR \SUBBYTES[4].a/U5325  ( .A(\SUBBYTES[4].a/w1694 ), .B(
        \SUBBYTES[4].a/w1697 ), .Z(n9913) );
  XOR \SUBBYTES[4].a/U5323  ( .A(n10785), .B(n9916), .Z(n9914) );
  XOR \SUBBYTES[4].a/U5322  ( .A(n10787), .B(n10786), .Z(n9915) );
  XOR \SUBBYTES[4].a/U5321  ( .A(\SUBBYTES[4].a/w1702 ), .B(
        \SUBBYTES[4].a/w1729 ), .Z(n9916) );
  XOR \SUBBYTES[4].a/U5319  ( .A(n10788), .B(n9919), .Z(n9917) );
  XOR \SUBBYTES[4].a/U5318  ( .A(\SUBBYTES[4].a/w1735 ), .B(
        \SUBBYTES[4].a/w1737 ), .Z(n9918) );
  XOR \SUBBYTES[4].a/U5317  ( .A(\SUBBYTES[4].a/w1695 ), .B(
        \SUBBYTES[4].a/w1727 ), .Z(n9919) );
  XOR \SUBBYTES[4].a/U5316  ( .A(\SUBBYTES[4].a/w1527 ), .B(
        \SUBBYTES[4].a/w1528 ), .Z(n10790) );
  XOR \SUBBYTES[4].a/U5315  ( .A(n10790), .B(n9920), .Z(n10789) );
  XOR \SUBBYTES[4].a/U5314  ( .A(\SUBBYTES[4].a/w1520 ), .B(
        \SUBBYTES[4].a/w1537 ), .Z(n9920) );
  XOR \SUBBYTES[4].a/U5312  ( .A(\SUBBYTES[4].a/w1519 ), .B(
        \SUBBYTES[4].a/w1534 ), .Z(n9921) );
  XOR \SUBBYTES[4].a/U5311  ( .A(n10790), .B(n9922), .Z(n10945) );
  XOR \SUBBYTES[4].a/U5310  ( .A(\SUBBYTES[4].a/w1534 ), .B(
        \SUBBYTES[4].a/w1535 ), .Z(n9922) );
  XOR \SUBBYTES[4].a/U5309  ( .A(\SUBBYTES[4].a/w1496 ), .B(n9923), .Z(n10792)
         );
  XOR \SUBBYTES[4].a/U5308  ( .A(\SUBBYTES[4].a/w1487 ), .B(
        \SUBBYTES[4].a/w1488 ), .Z(n9923) );
  XOR \SUBBYTES[4].a/U5306  ( .A(\SUBBYTES[4].a/w1498 ), .B(n10945), .Z(n9924)
         );
  XOR \SUBBYTES[4].a/U5305  ( .A(n9926), .B(n9925), .Z(n10793) );
  XOR \SUBBYTES[4].a/U5304  ( .A(n9928), .B(n9927), .Z(n9925) );
  XOR \SUBBYTES[4].a/U5303  ( .A(\SUBBYTES[4].a/w1534 ), .B(
        \SUBBYTES[4].a/w1535 ), .Z(n9926) );
  XOR \SUBBYTES[4].a/U5302  ( .A(\SUBBYTES[4].a/w1498 ), .B(
        \SUBBYTES[4].a/w1522 ), .Z(n9927) );
  XOR \SUBBYTES[4].a/U5301  ( .A(\SUBBYTES[4].a/w1487 ), .B(
        \SUBBYTES[4].a/w1496 ), .Z(n9928) );
  XOR \SUBBYTES[4].a/U5300  ( .A(\SUBBYTES[4].a/w1519 ), .B(n9929), .Z(n10791)
         );
  XOR \SUBBYTES[4].a/U5299  ( .A(\SUBBYTES[4].a/w1502 ), .B(
        \SUBBYTES[4].a/w1505 ), .Z(n9929) );
  XOR \SUBBYTES[4].a/U5297  ( .A(\SUBBYTES[4].a/w1490 ), .B(n10793), .Z(n9930)
         );
  XOR \SUBBYTES[4].a/U5295  ( .A(\SUBBYTES[4].a/w1522 ), .B(
        \SUBBYTES[4].a/w1535 ), .Z(n9931) );
  XOR \SUBBYTES[4].a/U5293  ( .A(n9935), .B(n9934), .Z(n9932) );
  XOR \SUBBYTES[4].a/U5292  ( .A(n9937), .B(n9936), .Z(n9933) );
  XOR \SUBBYTES[4].a/U5291  ( .A(\SUBBYTES[4].a/w1534 ), .B(
        \SUBBYTES[4].a/w1537 ), .Z(n9934) );
  XOR \SUBBYTES[4].a/U5290  ( .A(\SUBBYTES[4].a/w1527 ), .B(
        \SUBBYTES[4].a/w1530 ), .Z(n9935) );
  XOR \SUBBYTES[4].a/U5289  ( .A(\SUBBYTES[4].a/w1502 ), .B(
        \SUBBYTES[4].a/w1503 ), .Z(n9936) );
  XOR \SUBBYTES[4].a/U5288  ( .A(\SUBBYTES[4].a/w1487 ), .B(
        \SUBBYTES[4].a/w1490 ), .Z(n9937) );
  XOR \SUBBYTES[4].a/U5286  ( .A(n10790), .B(n9940), .Z(n9938) );
  XOR \SUBBYTES[4].a/U5285  ( .A(n10792), .B(n10791), .Z(n9939) );
  XOR \SUBBYTES[4].a/U5284  ( .A(\SUBBYTES[4].a/w1495 ), .B(
        \SUBBYTES[4].a/w1522 ), .Z(n9940) );
  XOR \SUBBYTES[4].a/U5282  ( .A(n10793), .B(n9943), .Z(n9941) );
  XOR \SUBBYTES[4].a/U5281  ( .A(\SUBBYTES[4].a/w1528 ), .B(
        \SUBBYTES[4].a/w1530 ), .Z(n9942) );
  XOR \SUBBYTES[4].a/U5280  ( .A(\SUBBYTES[4].a/w1488 ), .B(
        \SUBBYTES[4].a/w1520 ), .Z(n9943) );
  XOR \SUBBYTES[4].a/U5279  ( .A(\SUBBYTES[4].a/w1320 ), .B(
        \SUBBYTES[4].a/w1321 ), .Z(n10795) );
  XOR \SUBBYTES[4].a/U5278  ( .A(n10795), .B(n9944), .Z(n10794) );
  XOR \SUBBYTES[4].a/U5277  ( .A(\SUBBYTES[4].a/w1313 ), .B(
        \SUBBYTES[4].a/w1330 ), .Z(n9944) );
  XOR \SUBBYTES[4].a/U5275  ( .A(\SUBBYTES[4].a/w1312 ), .B(
        \SUBBYTES[4].a/w1327 ), .Z(n9945) );
  XOR \SUBBYTES[4].a/U5274  ( .A(n10795), .B(n9946), .Z(n10946) );
  XOR \SUBBYTES[4].a/U5273  ( .A(\SUBBYTES[4].a/w1327 ), .B(
        \SUBBYTES[4].a/w1328 ), .Z(n9946) );
  XOR \SUBBYTES[4].a/U5272  ( .A(\SUBBYTES[4].a/w1289 ), .B(n9947), .Z(n10797)
         );
  XOR \SUBBYTES[4].a/U5271  ( .A(\SUBBYTES[4].a/w1280 ), .B(
        \SUBBYTES[4].a/w1281 ), .Z(n9947) );
  XOR \SUBBYTES[4].a/U5269  ( .A(\SUBBYTES[4].a/w1291 ), .B(n10946), .Z(n9948)
         );
  XOR \SUBBYTES[4].a/U5268  ( .A(n9950), .B(n9949), .Z(n10798) );
  XOR \SUBBYTES[4].a/U5267  ( .A(n9952), .B(n9951), .Z(n9949) );
  XOR \SUBBYTES[4].a/U5266  ( .A(\SUBBYTES[4].a/w1327 ), .B(
        \SUBBYTES[4].a/w1328 ), .Z(n9950) );
  XOR \SUBBYTES[4].a/U5265  ( .A(\SUBBYTES[4].a/w1291 ), .B(
        \SUBBYTES[4].a/w1315 ), .Z(n9951) );
  XOR \SUBBYTES[4].a/U5264  ( .A(\SUBBYTES[4].a/w1280 ), .B(
        \SUBBYTES[4].a/w1289 ), .Z(n9952) );
  XOR \SUBBYTES[4].a/U5263  ( .A(\SUBBYTES[4].a/w1312 ), .B(n9953), .Z(n10796)
         );
  XOR \SUBBYTES[4].a/U5262  ( .A(\SUBBYTES[4].a/w1295 ), .B(
        \SUBBYTES[4].a/w1298 ), .Z(n9953) );
  XOR \SUBBYTES[4].a/U5260  ( .A(\SUBBYTES[4].a/w1283 ), .B(n10798), .Z(n9954)
         );
  XOR \SUBBYTES[4].a/U5258  ( .A(\SUBBYTES[4].a/w1315 ), .B(
        \SUBBYTES[4].a/w1328 ), .Z(n9955) );
  XOR \SUBBYTES[4].a/U5256  ( .A(n9959), .B(n9958), .Z(n9956) );
  XOR \SUBBYTES[4].a/U5255  ( .A(n9961), .B(n9960), .Z(n9957) );
  XOR \SUBBYTES[4].a/U5254  ( .A(\SUBBYTES[4].a/w1327 ), .B(
        \SUBBYTES[4].a/w1330 ), .Z(n9958) );
  XOR \SUBBYTES[4].a/U5253  ( .A(\SUBBYTES[4].a/w1320 ), .B(
        \SUBBYTES[4].a/w1323 ), .Z(n9959) );
  XOR \SUBBYTES[4].a/U5252  ( .A(\SUBBYTES[4].a/w1295 ), .B(
        \SUBBYTES[4].a/w1296 ), .Z(n9960) );
  XOR \SUBBYTES[4].a/U5251  ( .A(\SUBBYTES[4].a/w1280 ), .B(
        \SUBBYTES[4].a/w1283 ), .Z(n9961) );
  XOR \SUBBYTES[4].a/U5249  ( .A(n10795), .B(n9964), .Z(n9962) );
  XOR \SUBBYTES[4].a/U5248  ( .A(n10797), .B(n10796), .Z(n9963) );
  XOR \SUBBYTES[4].a/U5247  ( .A(\SUBBYTES[4].a/w1288 ), .B(
        \SUBBYTES[4].a/w1315 ), .Z(n9964) );
  XOR \SUBBYTES[4].a/U5245  ( .A(n10798), .B(n9967), .Z(n9965) );
  XOR \SUBBYTES[4].a/U5244  ( .A(\SUBBYTES[4].a/w1321 ), .B(
        \SUBBYTES[4].a/w1323 ), .Z(n9966) );
  XOR \SUBBYTES[4].a/U5243  ( .A(\SUBBYTES[4].a/w1281 ), .B(
        \SUBBYTES[4].a/w1313 ), .Z(n9967) );
  XOR \SUBBYTES[4].a/U5242  ( .A(\SUBBYTES[4].a/w1113 ), .B(
        \SUBBYTES[4].a/w1114 ), .Z(n10800) );
  XOR \SUBBYTES[4].a/U5241  ( .A(n10800), .B(n9968), .Z(n10799) );
  XOR \SUBBYTES[4].a/U5240  ( .A(\SUBBYTES[4].a/w1106 ), .B(
        \SUBBYTES[4].a/w1123 ), .Z(n9968) );
  XOR \SUBBYTES[4].a/U5238  ( .A(\SUBBYTES[4].a/w1105 ), .B(
        \SUBBYTES[4].a/w1120 ), .Z(n9969) );
  XOR \SUBBYTES[4].a/U5237  ( .A(n10800), .B(n9970), .Z(n10947) );
  XOR \SUBBYTES[4].a/U5236  ( .A(\SUBBYTES[4].a/w1120 ), .B(
        \SUBBYTES[4].a/w1121 ), .Z(n9970) );
  XOR \SUBBYTES[4].a/U5235  ( .A(\SUBBYTES[4].a/w1082 ), .B(n9971), .Z(n10802)
         );
  XOR \SUBBYTES[4].a/U5234  ( .A(\SUBBYTES[4].a/w1073 ), .B(
        \SUBBYTES[4].a/w1074 ), .Z(n9971) );
  XOR \SUBBYTES[4].a/U5232  ( .A(\SUBBYTES[4].a/w1084 ), .B(n10947), .Z(n9972)
         );
  XOR \SUBBYTES[4].a/U5231  ( .A(n9974), .B(n9973), .Z(n10803) );
  XOR \SUBBYTES[4].a/U5230  ( .A(n9976), .B(n9975), .Z(n9973) );
  XOR \SUBBYTES[4].a/U5229  ( .A(\SUBBYTES[4].a/w1120 ), .B(
        \SUBBYTES[4].a/w1121 ), .Z(n9974) );
  XOR \SUBBYTES[4].a/U5228  ( .A(\SUBBYTES[4].a/w1084 ), .B(
        \SUBBYTES[4].a/w1108 ), .Z(n9975) );
  XOR \SUBBYTES[4].a/U5227  ( .A(\SUBBYTES[4].a/w1073 ), .B(
        \SUBBYTES[4].a/w1082 ), .Z(n9976) );
  XOR \SUBBYTES[4].a/U5226  ( .A(\SUBBYTES[4].a/w1105 ), .B(n9977), .Z(n10801)
         );
  XOR \SUBBYTES[4].a/U5225  ( .A(\SUBBYTES[4].a/w1088 ), .B(
        \SUBBYTES[4].a/w1091 ), .Z(n9977) );
  XOR \SUBBYTES[4].a/U5223  ( .A(\SUBBYTES[4].a/w1076 ), .B(n10803), .Z(n9978)
         );
  XOR \SUBBYTES[4].a/U5221  ( .A(\SUBBYTES[4].a/w1108 ), .B(
        \SUBBYTES[4].a/w1121 ), .Z(n9979) );
  XOR \SUBBYTES[4].a/U5219  ( .A(n9983), .B(n9982), .Z(n9980) );
  XOR \SUBBYTES[4].a/U5218  ( .A(n9985), .B(n9984), .Z(n9981) );
  XOR \SUBBYTES[4].a/U5217  ( .A(\SUBBYTES[4].a/w1120 ), .B(
        \SUBBYTES[4].a/w1123 ), .Z(n9982) );
  XOR \SUBBYTES[4].a/U5216  ( .A(\SUBBYTES[4].a/w1113 ), .B(
        \SUBBYTES[4].a/w1116 ), .Z(n9983) );
  XOR \SUBBYTES[4].a/U5215  ( .A(\SUBBYTES[4].a/w1088 ), .B(
        \SUBBYTES[4].a/w1089 ), .Z(n9984) );
  XOR \SUBBYTES[4].a/U5214  ( .A(\SUBBYTES[4].a/w1073 ), .B(
        \SUBBYTES[4].a/w1076 ), .Z(n9985) );
  XOR \SUBBYTES[4].a/U5212  ( .A(n10800), .B(n9988), .Z(n9986) );
  XOR \SUBBYTES[4].a/U5211  ( .A(n10802), .B(n10801), .Z(n9987) );
  XOR \SUBBYTES[4].a/U5210  ( .A(\SUBBYTES[4].a/w1081 ), .B(
        \SUBBYTES[4].a/w1108 ), .Z(n9988) );
  XOR \SUBBYTES[4].a/U5208  ( .A(n10803), .B(n9991), .Z(n9989) );
  XOR \SUBBYTES[4].a/U5207  ( .A(\SUBBYTES[4].a/w1114 ), .B(
        \SUBBYTES[4].a/w1116 ), .Z(n9990) );
  XOR \SUBBYTES[4].a/U5206  ( .A(\SUBBYTES[4].a/w1074 ), .B(
        \SUBBYTES[4].a/w1106 ), .Z(n9991) );
  XOR \SUBBYTES[4].a/U5205  ( .A(\SUBBYTES[4].a/w906 ), .B(
        \SUBBYTES[4].a/w907 ), .Z(n10805) );
  XOR \SUBBYTES[4].a/U5204  ( .A(n10805), .B(n9992), .Z(n10804) );
  XOR \SUBBYTES[4].a/U5203  ( .A(\SUBBYTES[4].a/w899 ), .B(
        \SUBBYTES[4].a/w916 ), .Z(n9992) );
  XOR \SUBBYTES[4].a/U5201  ( .A(\SUBBYTES[4].a/w898 ), .B(
        \SUBBYTES[4].a/w913 ), .Z(n9993) );
  XOR \SUBBYTES[4].a/U5200  ( .A(n10805), .B(n9994), .Z(n10948) );
  XOR \SUBBYTES[4].a/U5199  ( .A(\SUBBYTES[4].a/w913 ), .B(
        \SUBBYTES[4].a/w914 ), .Z(n9994) );
  XOR \SUBBYTES[4].a/U5198  ( .A(\SUBBYTES[4].a/w875 ), .B(n9995), .Z(n10807)
         );
  XOR \SUBBYTES[4].a/U5197  ( .A(\SUBBYTES[4].a/w866 ), .B(
        \SUBBYTES[4].a/w867 ), .Z(n9995) );
  XOR \SUBBYTES[4].a/U5195  ( .A(\SUBBYTES[4].a/w877 ), .B(n10948), .Z(n9996)
         );
  XOR \SUBBYTES[4].a/U5194  ( .A(n9998), .B(n9997), .Z(n10808) );
  XOR \SUBBYTES[4].a/U5193  ( .A(n10000), .B(n9999), .Z(n9997) );
  XOR \SUBBYTES[4].a/U5192  ( .A(\SUBBYTES[4].a/w913 ), .B(
        \SUBBYTES[4].a/w914 ), .Z(n9998) );
  XOR \SUBBYTES[4].a/U5191  ( .A(\SUBBYTES[4].a/w877 ), .B(
        \SUBBYTES[4].a/w901 ), .Z(n9999) );
  XOR \SUBBYTES[4].a/U5190  ( .A(\SUBBYTES[4].a/w866 ), .B(
        \SUBBYTES[4].a/w875 ), .Z(n10000) );
  XOR \SUBBYTES[4].a/U5189  ( .A(\SUBBYTES[4].a/w898 ), .B(n10001), .Z(n10806)
         );
  XOR \SUBBYTES[4].a/U5188  ( .A(\SUBBYTES[4].a/w881 ), .B(
        \SUBBYTES[4].a/w884 ), .Z(n10001) );
  XOR \SUBBYTES[4].a/U5186  ( .A(\SUBBYTES[4].a/w869 ), .B(n10808), .Z(n10002)
         );
  XOR \SUBBYTES[4].a/U5184  ( .A(\SUBBYTES[4].a/w901 ), .B(
        \SUBBYTES[4].a/w914 ), .Z(n10003) );
  XOR \SUBBYTES[4].a/U5182  ( .A(n10007), .B(n10006), .Z(n10004) );
  XOR \SUBBYTES[4].a/U5181  ( .A(n10009), .B(n10008), .Z(n10005) );
  XOR \SUBBYTES[4].a/U5180  ( .A(\SUBBYTES[4].a/w913 ), .B(
        \SUBBYTES[4].a/w916 ), .Z(n10006) );
  XOR \SUBBYTES[4].a/U5179  ( .A(\SUBBYTES[4].a/w906 ), .B(
        \SUBBYTES[4].a/w909 ), .Z(n10007) );
  XOR \SUBBYTES[4].a/U5178  ( .A(\SUBBYTES[4].a/w881 ), .B(
        \SUBBYTES[4].a/w882 ), .Z(n10008) );
  XOR \SUBBYTES[4].a/U5177  ( .A(\SUBBYTES[4].a/w866 ), .B(
        \SUBBYTES[4].a/w869 ), .Z(n10009) );
  XOR \SUBBYTES[4].a/U5175  ( .A(n10805), .B(n10012), .Z(n10010) );
  XOR \SUBBYTES[4].a/U5174  ( .A(n10807), .B(n10806), .Z(n10011) );
  XOR \SUBBYTES[4].a/U5173  ( .A(\SUBBYTES[4].a/w874 ), .B(
        \SUBBYTES[4].a/w901 ), .Z(n10012) );
  XOR \SUBBYTES[4].a/U5171  ( .A(n10808), .B(n10015), .Z(n10013) );
  XOR \SUBBYTES[4].a/U5170  ( .A(\SUBBYTES[4].a/w907 ), .B(
        \SUBBYTES[4].a/w909 ), .Z(n10014) );
  XOR \SUBBYTES[4].a/U5169  ( .A(\SUBBYTES[4].a/w867 ), .B(
        \SUBBYTES[4].a/w899 ), .Z(n10015) );
  XOR \SUBBYTES[4].a/U5168  ( .A(\SUBBYTES[4].a/w699 ), .B(
        \SUBBYTES[4].a/w700 ), .Z(n10810) );
  XOR \SUBBYTES[4].a/U5167  ( .A(n10810), .B(n10016), .Z(n10809) );
  XOR \SUBBYTES[4].a/U5166  ( .A(\SUBBYTES[4].a/w692 ), .B(
        \SUBBYTES[4].a/w709 ), .Z(n10016) );
  XOR \SUBBYTES[4].a/U5164  ( .A(\SUBBYTES[4].a/w691 ), .B(
        \SUBBYTES[4].a/w706 ), .Z(n10017) );
  XOR \SUBBYTES[4].a/U5163  ( .A(n10810), .B(n10018), .Z(n10949) );
  XOR \SUBBYTES[4].a/U5162  ( .A(\SUBBYTES[4].a/w706 ), .B(
        \SUBBYTES[4].a/w707 ), .Z(n10018) );
  XOR \SUBBYTES[4].a/U5161  ( .A(\SUBBYTES[4].a/w668 ), .B(n10019), .Z(n10812)
         );
  XOR \SUBBYTES[4].a/U5160  ( .A(\SUBBYTES[4].a/w659 ), .B(
        \SUBBYTES[4].a/w660 ), .Z(n10019) );
  XOR \SUBBYTES[4].a/U5158  ( .A(\SUBBYTES[4].a/w670 ), .B(n10949), .Z(n10020)
         );
  XOR \SUBBYTES[4].a/U5157  ( .A(n10022), .B(n10021), .Z(n10813) );
  XOR \SUBBYTES[4].a/U5156  ( .A(n10024), .B(n10023), .Z(n10021) );
  XOR \SUBBYTES[4].a/U5155  ( .A(\SUBBYTES[4].a/w706 ), .B(
        \SUBBYTES[4].a/w707 ), .Z(n10022) );
  XOR \SUBBYTES[4].a/U5154  ( .A(\SUBBYTES[4].a/w670 ), .B(
        \SUBBYTES[4].a/w694 ), .Z(n10023) );
  XOR \SUBBYTES[4].a/U5153  ( .A(\SUBBYTES[4].a/w659 ), .B(
        \SUBBYTES[4].a/w668 ), .Z(n10024) );
  XOR \SUBBYTES[4].a/U5152  ( .A(\SUBBYTES[4].a/w691 ), .B(n10025), .Z(n10811)
         );
  XOR \SUBBYTES[4].a/U5151  ( .A(\SUBBYTES[4].a/w674 ), .B(
        \SUBBYTES[4].a/w677 ), .Z(n10025) );
  XOR \SUBBYTES[4].a/U5149  ( .A(\SUBBYTES[4].a/w662 ), .B(n10813), .Z(n10026)
         );
  XOR \SUBBYTES[4].a/U5147  ( .A(\SUBBYTES[4].a/w694 ), .B(
        \SUBBYTES[4].a/w707 ), .Z(n10027) );
  XOR \SUBBYTES[4].a/U5145  ( .A(n10031), .B(n10030), .Z(n10028) );
  XOR \SUBBYTES[4].a/U5144  ( .A(n10033), .B(n10032), .Z(n10029) );
  XOR \SUBBYTES[4].a/U5143  ( .A(\SUBBYTES[4].a/w706 ), .B(
        \SUBBYTES[4].a/w709 ), .Z(n10030) );
  XOR \SUBBYTES[4].a/U5142  ( .A(\SUBBYTES[4].a/w699 ), .B(
        \SUBBYTES[4].a/w702 ), .Z(n10031) );
  XOR \SUBBYTES[4].a/U5141  ( .A(\SUBBYTES[4].a/w674 ), .B(
        \SUBBYTES[4].a/w675 ), .Z(n10032) );
  XOR \SUBBYTES[4].a/U5140  ( .A(\SUBBYTES[4].a/w659 ), .B(
        \SUBBYTES[4].a/w662 ), .Z(n10033) );
  XOR \SUBBYTES[4].a/U5138  ( .A(n10810), .B(n10036), .Z(n10034) );
  XOR \SUBBYTES[4].a/U5137  ( .A(n10812), .B(n10811), .Z(n10035) );
  XOR \SUBBYTES[4].a/U5136  ( .A(\SUBBYTES[4].a/w667 ), .B(
        \SUBBYTES[4].a/w694 ), .Z(n10036) );
  XOR \SUBBYTES[4].a/U5134  ( .A(n10813), .B(n10039), .Z(n10037) );
  XOR \SUBBYTES[4].a/U5133  ( .A(\SUBBYTES[4].a/w700 ), .B(
        \SUBBYTES[4].a/w702 ), .Z(n10038) );
  XOR \SUBBYTES[4].a/U5132  ( .A(\SUBBYTES[4].a/w660 ), .B(
        \SUBBYTES[4].a/w692 ), .Z(n10039) );
  XOR \SUBBYTES[4].a/U5131  ( .A(\SUBBYTES[4].a/w492 ), .B(
        \SUBBYTES[4].a/w493 ), .Z(n10815) );
  XOR \SUBBYTES[4].a/U5130  ( .A(n10815), .B(n10040), .Z(n10814) );
  XOR \SUBBYTES[4].a/U5129  ( .A(\SUBBYTES[4].a/w485 ), .B(
        \SUBBYTES[4].a/w502 ), .Z(n10040) );
  XOR \SUBBYTES[4].a/U5127  ( .A(\SUBBYTES[4].a/w484 ), .B(
        \SUBBYTES[4].a/w499 ), .Z(n10041) );
  XOR \SUBBYTES[4].a/U5126  ( .A(n10815), .B(n10042), .Z(n10950) );
  XOR \SUBBYTES[4].a/U5125  ( .A(\SUBBYTES[4].a/w499 ), .B(
        \SUBBYTES[4].a/w500 ), .Z(n10042) );
  XOR \SUBBYTES[4].a/U5124  ( .A(\SUBBYTES[4].a/w461 ), .B(n10043), .Z(n10817)
         );
  XOR \SUBBYTES[4].a/U5123  ( .A(\SUBBYTES[4].a/w452 ), .B(
        \SUBBYTES[4].a/w453 ), .Z(n10043) );
  XOR \SUBBYTES[4].a/U5121  ( .A(\SUBBYTES[4].a/w463 ), .B(n10950), .Z(n10044)
         );
  XOR \SUBBYTES[4].a/U5120  ( .A(n10046), .B(n10045), .Z(n10818) );
  XOR \SUBBYTES[4].a/U5119  ( .A(n10048), .B(n10047), .Z(n10045) );
  XOR \SUBBYTES[4].a/U5118  ( .A(\SUBBYTES[4].a/w499 ), .B(
        \SUBBYTES[4].a/w500 ), .Z(n10046) );
  XOR \SUBBYTES[4].a/U5117  ( .A(\SUBBYTES[4].a/w463 ), .B(
        \SUBBYTES[4].a/w487 ), .Z(n10047) );
  XOR \SUBBYTES[4].a/U5116  ( .A(\SUBBYTES[4].a/w452 ), .B(
        \SUBBYTES[4].a/w461 ), .Z(n10048) );
  XOR \SUBBYTES[4].a/U5115  ( .A(\SUBBYTES[4].a/w484 ), .B(n10049), .Z(n10816)
         );
  XOR \SUBBYTES[4].a/U5114  ( .A(\SUBBYTES[4].a/w467 ), .B(
        \SUBBYTES[4].a/w470 ), .Z(n10049) );
  XOR \SUBBYTES[4].a/U5112  ( .A(\SUBBYTES[4].a/w455 ), .B(n10818), .Z(n10050)
         );
  XOR \SUBBYTES[4].a/U5110  ( .A(\SUBBYTES[4].a/w487 ), .B(
        \SUBBYTES[4].a/w500 ), .Z(n10051) );
  XOR \SUBBYTES[4].a/U5108  ( .A(n10055), .B(n10054), .Z(n10052) );
  XOR \SUBBYTES[4].a/U5107  ( .A(n10057), .B(n10056), .Z(n10053) );
  XOR \SUBBYTES[4].a/U5106  ( .A(\SUBBYTES[4].a/w499 ), .B(
        \SUBBYTES[4].a/w502 ), .Z(n10054) );
  XOR \SUBBYTES[4].a/U5105  ( .A(\SUBBYTES[4].a/w492 ), .B(
        \SUBBYTES[4].a/w495 ), .Z(n10055) );
  XOR \SUBBYTES[4].a/U5104  ( .A(\SUBBYTES[4].a/w467 ), .B(
        \SUBBYTES[4].a/w468 ), .Z(n10056) );
  XOR \SUBBYTES[4].a/U5103  ( .A(\SUBBYTES[4].a/w452 ), .B(
        \SUBBYTES[4].a/w455 ), .Z(n10057) );
  XOR \SUBBYTES[4].a/U5101  ( .A(n10815), .B(n10060), .Z(n10058) );
  XOR \SUBBYTES[4].a/U5100  ( .A(n10817), .B(n10816), .Z(n10059) );
  XOR \SUBBYTES[4].a/U5099  ( .A(\SUBBYTES[4].a/w460 ), .B(
        \SUBBYTES[4].a/w487 ), .Z(n10060) );
  XOR \SUBBYTES[4].a/U5097  ( .A(n10818), .B(n10063), .Z(n10061) );
  XOR \SUBBYTES[4].a/U5096  ( .A(\SUBBYTES[4].a/w493 ), .B(
        \SUBBYTES[4].a/w495 ), .Z(n10062) );
  XOR \SUBBYTES[4].a/U5095  ( .A(\SUBBYTES[4].a/w453 ), .B(
        \SUBBYTES[4].a/w485 ), .Z(n10063) );
  XOR \SUBBYTES[4].a/U5094  ( .A(\SUBBYTES[4].a/w285 ), .B(
        \SUBBYTES[4].a/w286 ), .Z(n10820) );
  XOR \SUBBYTES[4].a/U5093  ( .A(n10820), .B(n10064), .Z(n10819) );
  XOR \SUBBYTES[4].a/U5092  ( .A(\SUBBYTES[4].a/w278 ), .B(
        \SUBBYTES[4].a/w295 ), .Z(n10064) );
  XOR \SUBBYTES[4].a/U5090  ( .A(\SUBBYTES[4].a/w277 ), .B(
        \SUBBYTES[4].a/w292 ), .Z(n10065) );
  XOR \SUBBYTES[4].a/U5089  ( .A(n10820), .B(n10066), .Z(n10951) );
  XOR \SUBBYTES[4].a/U5088  ( .A(\SUBBYTES[4].a/w292 ), .B(
        \SUBBYTES[4].a/w293 ), .Z(n10066) );
  XOR \SUBBYTES[4].a/U5087  ( .A(\SUBBYTES[4].a/w254 ), .B(n10067), .Z(n10822)
         );
  XOR \SUBBYTES[4].a/U5086  ( .A(\SUBBYTES[4].a/w245 ), .B(
        \SUBBYTES[4].a/w246 ), .Z(n10067) );
  XOR \SUBBYTES[4].a/U5084  ( .A(\SUBBYTES[4].a/w256 ), .B(n10951), .Z(n10068)
         );
  XOR \SUBBYTES[4].a/U5083  ( .A(n10070), .B(n10069), .Z(n10823) );
  XOR \SUBBYTES[4].a/U5082  ( .A(n10072), .B(n10071), .Z(n10069) );
  XOR \SUBBYTES[4].a/U5081  ( .A(\SUBBYTES[4].a/w292 ), .B(
        \SUBBYTES[4].a/w293 ), .Z(n10070) );
  XOR \SUBBYTES[4].a/U5080  ( .A(\SUBBYTES[4].a/w256 ), .B(
        \SUBBYTES[4].a/w280 ), .Z(n10071) );
  XOR \SUBBYTES[4].a/U5079  ( .A(\SUBBYTES[4].a/w245 ), .B(
        \SUBBYTES[4].a/w254 ), .Z(n10072) );
  XOR \SUBBYTES[4].a/U5078  ( .A(\SUBBYTES[4].a/w277 ), .B(n10073), .Z(n10821)
         );
  XOR \SUBBYTES[4].a/U5077  ( .A(\SUBBYTES[4].a/w260 ), .B(
        \SUBBYTES[4].a/w263 ), .Z(n10073) );
  XOR \SUBBYTES[4].a/U5075  ( .A(\SUBBYTES[4].a/w248 ), .B(n10823), .Z(n10074)
         );
  XOR \SUBBYTES[4].a/U5073  ( .A(\SUBBYTES[4].a/w280 ), .B(
        \SUBBYTES[4].a/w293 ), .Z(n10075) );
  XOR \SUBBYTES[4].a/U5071  ( .A(n10079), .B(n10078), .Z(n10076) );
  XOR \SUBBYTES[4].a/U5070  ( .A(n10081), .B(n10080), .Z(n10077) );
  XOR \SUBBYTES[4].a/U5069  ( .A(\SUBBYTES[4].a/w292 ), .B(
        \SUBBYTES[4].a/w295 ), .Z(n10078) );
  XOR \SUBBYTES[4].a/U5068  ( .A(\SUBBYTES[4].a/w285 ), .B(
        \SUBBYTES[4].a/w288 ), .Z(n10079) );
  XOR \SUBBYTES[4].a/U5067  ( .A(\SUBBYTES[4].a/w260 ), .B(
        \SUBBYTES[4].a/w261 ), .Z(n10080) );
  XOR \SUBBYTES[4].a/U5066  ( .A(\SUBBYTES[4].a/w245 ), .B(
        \SUBBYTES[4].a/w248 ), .Z(n10081) );
  XOR \SUBBYTES[4].a/U5064  ( .A(n10820), .B(n10084), .Z(n10082) );
  XOR \SUBBYTES[4].a/U5063  ( .A(n10822), .B(n10821), .Z(n10083) );
  XOR \SUBBYTES[4].a/U5062  ( .A(\SUBBYTES[4].a/w253 ), .B(
        \SUBBYTES[4].a/w280 ), .Z(n10084) );
  XOR \SUBBYTES[4].a/U5060  ( .A(n10823), .B(n10087), .Z(n10085) );
  XOR \SUBBYTES[4].a/U5059  ( .A(\SUBBYTES[4].a/w286 ), .B(
        \SUBBYTES[4].a/w288 ), .Z(n10086) );
  XOR \SUBBYTES[4].a/U5058  ( .A(\SUBBYTES[4].a/w246 ), .B(
        \SUBBYTES[4].a/w278 ), .Z(n10087) );
  XOR \SUBBYTES[4].a/U5057  ( .A(\w1[4][1] ), .B(n10088), .Z(n10824) );
  XOR \SUBBYTES[4].a/U5056  ( .A(\w1[4][3] ), .B(\w1[4][2] ), .Z(n10088) );
  XOR \SUBBYTES[4].a/U5055  ( .A(\w1[4][6] ), .B(n10824), .Z(
        \SUBBYTES[4].a/w3378 ) );
  XOR \SUBBYTES[4].a/U5054  ( .A(\w1[4][0] ), .B(\SUBBYTES[4].a/w3378 ), .Z(
        \SUBBYTES[4].a/w3265 ) );
  XOR \SUBBYTES[4].a/U5053  ( .A(\w1[4][0] ), .B(n10089), .Z(
        \SUBBYTES[4].a/w3266 ) );
  XOR \SUBBYTES[4].a/U5052  ( .A(\w1[4][6] ), .B(\w1[4][5] ), .Z(n10089) );
  XOR \SUBBYTES[4].a/U5051  ( .A(\w1[4][5] ), .B(n10824), .Z(
        \SUBBYTES[4].a/w3396 ) );
  XOR \SUBBYTES[4].a/U5050  ( .A(n10091), .B(n10090), .Z(\SUBBYTES[4].a/w3389 ) );
  XOR \SUBBYTES[4].a/U5049  ( .A(\w1[4][3] ), .B(\w1[4][1] ), .Z(n10090) );
  XOR \SUBBYTES[4].a/U5048  ( .A(\w1[4][7] ), .B(\w1[4][4] ), .Z(n10091) );
  XOR \SUBBYTES[4].a/U5047  ( .A(\w1[4][0] ), .B(\SUBBYTES[4].a/w3389 ), .Z(
        \SUBBYTES[4].a/w3268 ) );
  XOR \SUBBYTES[4].a/U5046  ( .A(n10093), .B(n10092), .Z(\SUBBYTES[4].a/w3376 ) );
  XOR \SUBBYTES[4].a/U5045  ( .A(\SUBBYTES[4].a/w3337 ), .B(n1020), .Z(n10092)
         );
  XOR \SUBBYTES[4].a/U5044  ( .A(\SUBBYTES[4].a/w3330 ), .B(
        \SUBBYTES[4].a/w3333 ), .Z(n10093) );
  XOR \SUBBYTES[4].a/U5043  ( .A(n10095), .B(n10094), .Z(\SUBBYTES[4].a/w3377 ) );
  XOR \SUBBYTES[4].a/U5042  ( .A(\SUBBYTES[4].a/w3337 ), .B(n9703), .Z(n10094)
         );
  XOR \SUBBYTES[4].a/U5041  ( .A(\SUBBYTES[4].a/w3330 ), .B(n9702), .Z(n10095)
         );
  XOR \SUBBYTES[4].a/U5040  ( .A(\SUBBYTES[4].a/w3389 ), .B(n10096), .Z(
        \SUBBYTES[4].a/w3379 ) );
  XOR \SUBBYTES[4].a/U5039  ( .A(\w1[4][6] ), .B(\w1[4][5] ), .Z(n10096) );
  XOR \SUBBYTES[4].a/U5038  ( .A(n10098), .B(n10097), .Z(\SUBBYTES[4].a/w3380 ) );
  XOR \SUBBYTES[4].a/U5037  ( .A(n9703), .B(n1020), .Z(n10097) );
  XOR \SUBBYTES[4].a/U5036  ( .A(n9702), .B(\SUBBYTES[4].a/w3333 ), .Z(n10098)
         );
  XOR \SUBBYTES[4].a/U5035  ( .A(\w1[4][7] ), .B(\w1[4][2] ), .Z(n10830) );
  XOR \SUBBYTES[4].a/U5034  ( .A(n10830), .B(n10099), .Z(\SUBBYTES[4].a/w3381 ) );
  XOR \SUBBYTES[4].a/U5033  ( .A(\w1[4][5] ), .B(\w1[4][4] ), .Z(n10099) );
  XOR \SUBBYTES[4].a/U5032  ( .A(\w1[4][7] ), .B(\SUBBYTES[4].a/w3266 ), .Z(
        \SUBBYTES[4].a/w3269 ) );
  XOR \SUBBYTES[4].a/U5031  ( .A(\w1[4][1] ), .B(\SUBBYTES[4].a/w3266 ), .Z(
        \SUBBYTES[4].a/w3270 ) );
  XOR \SUBBYTES[4].a/U5030  ( .A(\w1[4][4] ), .B(\SUBBYTES[4].a/w3266 ), .Z(
        \SUBBYTES[4].a/w3271 ) );
  XOR \SUBBYTES[4].a/U5029  ( .A(\SUBBYTES[4].a/w3270 ), .B(n10830), .Z(
        \SUBBYTES[4].a/w3272 ) );
  XOR \SUBBYTES[4].a/U5028  ( .A(n10830), .B(n10100), .Z(\SUBBYTES[4].a/w3357 ) );
  XOR \SUBBYTES[4].a/U5027  ( .A(\w1[4][4] ), .B(\w1[4][1] ), .Z(n10100) );
  XOR \SUBBYTES[4].a/U5026  ( .A(n10102), .B(n10101), .Z(n10827) );
  XOR \SUBBYTES[4].a/U5025  ( .A(\w1[4][4] ), .B(n10103), .Z(n10101) );
  XOR \SUBBYTES[4].a/U5024  ( .A(\SUBBYTES[4].a/w3322 ), .B(\w1[4][6] ), .Z(
        n10102) );
  XOR \SUBBYTES[4].a/U5023  ( .A(\SUBBYTES[4].a/w3296 ), .B(
        \SUBBYTES[4].a/w3303 ), .Z(n10103) );
  XOR \SUBBYTES[4].a/U5022  ( .A(n10105), .B(n10104), .Z(n10825) );
  XOR \SUBBYTES[4].a/U5021  ( .A(\w1[4][1] ), .B(n10106), .Z(n10104) );
  XOR \SUBBYTES[4].a/U5020  ( .A(\SUBBYTES[4].a/w3321 ), .B(\w1[4][5] ), .Z(
        n10105) );
  XOR \SUBBYTES[4].a/U5019  ( .A(\SUBBYTES[4].a/w3297 ), .B(
        \SUBBYTES[4].a/w3304 ), .Z(n10106) );
  XOR \SUBBYTES[4].a/U5018  ( .A(n10827), .B(n10825), .Z(\SUBBYTES[4].a/w3327 ) );
  XOR \SUBBYTES[4].a/U5017  ( .A(\w1[4][5] ), .B(n10107), .Z(n10828) );
  XOR \SUBBYTES[4].a/U5016  ( .A(\SUBBYTES[4].a/w3289 ), .B(
        \SUBBYTES[4].a/w3299 ), .Z(n10107) );
  XOR \SUBBYTES[4].a/U5015  ( .A(n10109), .B(n10108), .Z(\SUBBYTES[4].a/w3314 ) );
  XOR \SUBBYTES[4].a/U5014  ( .A(n10828), .B(n10110), .Z(n10108) );
  XOR \SUBBYTES[4].a/U5013  ( .A(\w1[4][4] ), .B(\SUBBYTES[4].a/w3378 ), .Z(
        n10109) );
  XOR \SUBBYTES[4].a/U5012  ( .A(\SUBBYTES[4].a/w3291 ), .B(
        \SUBBYTES[4].a/w3296 ), .Z(n10110) );
  XOR \SUBBYTES[4].a/U5011  ( .A(n10112), .B(n10111), .Z(n10826) );
  XOR \SUBBYTES[4].a/U5010  ( .A(\SUBBYTES[4].a/w3324 ), .B(\w1[4][7] ), .Z(
        n10111) );
  XOR \SUBBYTES[4].a/U5009  ( .A(\SUBBYTES[4].a/w3299 ), .B(
        \SUBBYTES[4].a/w3306 ), .Z(n10112) );
  XOR \SUBBYTES[4].a/U5008  ( .A(n10825), .B(n10826), .Z(\SUBBYTES[4].a/w3326 ) );
  XOR \SUBBYTES[4].a/U5007  ( .A(\w1[4][3] ), .B(n10113), .Z(n10829) );
  XOR \SUBBYTES[4].a/U5006  ( .A(\SUBBYTES[4].a/w3288 ), .B(
        \SUBBYTES[4].a/w3291 ), .Z(n10113) );
  XOR \SUBBYTES[4].a/U5005  ( .A(n10115), .B(n10114), .Z(\SUBBYTES[4].a/w3315 ) );
  XOR \SUBBYTES[4].a/U5004  ( .A(n10829), .B(n10116), .Z(n10114) );
  XOR \SUBBYTES[4].a/U5003  ( .A(\w1[4][6] ), .B(\SUBBYTES[4].a/w3357 ), .Z(
        n10115) );
  XOR \SUBBYTES[4].a/U5002  ( .A(\SUBBYTES[4].a/w3296 ), .B(
        \SUBBYTES[4].a/w3297 ), .Z(n10116) );
  XOR \SUBBYTES[4].a/U5001  ( .A(n10827), .B(n10826), .Z(\SUBBYTES[4].a/w3335 ) );
  XOR \SUBBYTES[4].a/U5000  ( .A(n10118), .B(n10117), .Z(\SUBBYTES[4].a/w3336 ) );
  XOR \SUBBYTES[4].a/U4999  ( .A(\w1[4][7] ), .B(n10828), .Z(n10117) );
  XOR \SUBBYTES[4].a/U4998  ( .A(\SUBBYTES[4].a/w3288 ), .B(
        \SUBBYTES[4].a/w3297 ), .Z(n10118) );
  XOR \SUBBYTES[4].a/U4997  ( .A(n10120), .B(n10119), .Z(\SUBBYTES[4].a/w3312 ) );
  XOR \SUBBYTES[4].a/U4996  ( .A(n10122), .B(n10121), .Z(n10119) );
  XOR \SUBBYTES[4].a/U4995  ( .A(\w1[4][7] ), .B(\SUBBYTES[4].a/w3396 ), .Z(
        n10120) );
  XOR \SUBBYTES[4].a/U4994  ( .A(\SUBBYTES[4].a/w3303 ), .B(
        \SUBBYTES[4].a/w3306 ), .Z(n10121) );
  XOR \SUBBYTES[4].a/U4993  ( .A(\SUBBYTES[4].a/w3289 ), .B(
        \SUBBYTES[4].a/w3291 ), .Z(n10122) );
  XOR \SUBBYTES[4].a/U4992  ( .A(n10124), .B(n10123), .Z(\SUBBYTES[4].a/w3313 ) );
  XOR \SUBBYTES[4].a/U4991  ( .A(n10829), .B(n10125), .Z(n10123) );
  XOR \SUBBYTES[4].a/U4990  ( .A(\w1[4][5] ), .B(n10830), .Z(n10124) );
  XOR \SUBBYTES[4].a/U4989  ( .A(\SUBBYTES[4].a/w3303 ), .B(
        \SUBBYTES[4].a/w3304 ), .Z(n10125) );
  XOR \SUBBYTES[4].a/U4988  ( .A(n10127), .B(n10126), .Z(\SUBBYTES[4].a/w3329 ) );
  XOR \SUBBYTES[4].a/U4987  ( .A(\w1[4][1] ), .B(n10128), .Z(n10126) );
  XOR \SUBBYTES[4].a/U4986  ( .A(\SUBBYTES[4].a/w3304 ), .B(
        \SUBBYTES[4].a/w3306 ), .Z(n10127) );
  XOR \SUBBYTES[4].a/U4985  ( .A(\SUBBYTES[4].a/w3288 ), .B(
        \SUBBYTES[4].a/w3289 ), .Z(n10128) );
  XOR \SUBBYTES[4].a/U4984  ( .A(\w1[4][9] ), .B(n10129), .Z(n10831) );
  XOR \SUBBYTES[4].a/U4983  ( .A(\w1[4][11] ), .B(\w1[4][10] ), .Z(n10129) );
  XOR \SUBBYTES[4].a/U4982  ( .A(\w1[4][14] ), .B(n10831), .Z(
        \SUBBYTES[4].a/w3171 ) );
  XOR \SUBBYTES[4].a/U4981  ( .A(\w1[4][8] ), .B(\SUBBYTES[4].a/w3171 ), .Z(
        \SUBBYTES[4].a/w3058 ) );
  XOR \SUBBYTES[4].a/U4980  ( .A(\w1[4][8] ), .B(n10130), .Z(
        \SUBBYTES[4].a/w3059 ) );
  XOR \SUBBYTES[4].a/U4979  ( .A(\w1[4][14] ), .B(\w1[4][13] ), .Z(n10130) );
  XOR \SUBBYTES[4].a/U4978  ( .A(\w1[4][13] ), .B(n10831), .Z(
        \SUBBYTES[4].a/w3189 ) );
  XOR \SUBBYTES[4].a/U4977  ( .A(n10132), .B(n10131), .Z(\SUBBYTES[4].a/w3182 ) );
  XOR \SUBBYTES[4].a/U4976  ( .A(\w1[4][11] ), .B(\w1[4][9] ), .Z(n10131) );
  XOR \SUBBYTES[4].a/U4975  ( .A(\w1[4][15] ), .B(\w1[4][12] ), .Z(n10132) );
  XOR \SUBBYTES[4].a/U4974  ( .A(\w1[4][8] ), .B(\SUBBYTES[4].a/w3182 ), .Z(
        \SUBBYTES[4].a/w3061 ) );
  XOR \SUBBYTES[4].a/U4973  ( .A(n10134), .B(n10133), .Z(\SUBBYTES[4].a/w3169 ) );
  XOR \SUBBYTES[4].a/U4972  ( .A(\SUBBYTES[4].a/w3130 ), .B(n1019), .Z(n10133)
         );
  XOR \SUBBYTES[4].a/U4971  ( .A(\SUBBYTES[4].a/w3123 ), .B(
        \SUBBYTES[4].a/w3126 ), .Z(n10134) );
  XOR \SUBBYTES[4].a/U4970  ( .A(n10136), .B(n10135), .Z(\SUBBYTES[4].a/w3170 ) );
  XOR \SUBBYTES[4].a/U4969  ( .A(\SUBBYTES[4].a/w3130 ), .B(n9701), .Z(n10135)
         );
  XOR \SUBBYTES[4].a/U4968  ( .A(\SUBBYTES[4].a/w3123 ), .B(n9700), .Z(n10136)
         );
  XOR \SUBBYTES[4].a/U4967  ( .A(\SUBBYTES[4].a/w3182 ), .B(n10137), .Z(
        \SUBBYTES[4].a/w3172 ) );
  XOR \SUBBYTES[4].a/U4966  ( .A(\w1[4][14] ), .B(\w1[4][13] ), .Z(n10137) );
  XOR \SUBBYTES[4].a/U4965  ( .A(n10139), .B(n10138), .Z(\SUBBYTES[4].a/w3173 ) );
  XOR \SUBBYTES[4].a/U4964  ( .A(n9701), .B(n1019), .Z(n10138) );
  XOR \SUBBYTES[4].a/U4963  ( .A(n9700), .B(\SUBBYTES[4].a/w3126 ), .Z(n10139)
         );
  XOR \SUBBYTES[4].a/U4962  ( .A(\w1[4][15] ), .B(\w1[4][10] ), .Z(n10837) );
  XOR \SUBBYTES[4].a/U4961  ( .A(n10837), .B(n10140), .Z(\SUBBYTES[4].a/w3174 ) );
  XOR \SUBBYTES[4].a/U4960  ( .A(\w1[4][13] ), .B(\w1[4][12] ), .Z(n10140) );
  XOR \SUBBYTES[4].a/U4959  ( .A(\w1[4][15] ), .B(\SUBBYTES[4].a/w3059 ), .Z(
        \SUBBYTES[4].a/w3062 ) );
  XOR \SUBBYTES[4].a/U4958  ( .A(\w1[4][9] ), .B(\SUBBYTES[4].a/w3059 ), .Z(
        \SUBBYTES[4].a/w3063 ) );
  XOR \SUBBYTES[4].a/U4957  ( .A(\w1[4][12] ), .B(\SUBBYTES[4].a/w3059 ), .Z(
        \SUBBYTES[4].a/w3064 ) );
  XOR \SUBBYTES[4].a/U4956  ( .A(\SUBBYTES[4].a/w3063 ), .B(n10837), .Z(
        \SUBBYTES[4].a/w3065 ) );
  XOR \SUBBYTES[4].a/U4955  ( .A(n10837), .B(n10141), .Z(\SUBBYTES[4].a/w3150 ) );
  XOR \SUBBYTES[4].a/U4954  ( .A(\w1[4][12] ), .B(\w1[4][9] ), .Z(n10141) );
  XOR \SUBBYTES[4].a/U4953  ( .A(n10143), .B(n10142), .Z(n10834) );
  XOR \SUBBYTES[4].a/U4952  ( .A(\w1[4][12] ), .B(n10144), .Z(n10142) );
  XOR \SUBBYTES[4].a/U4951  ( .A(\SUBBYTES[4].a/w3115 ), .B(\w1[4][14] ), .Z(
        n10143) );
  XOR \SUBBYTES[4].a/U4950  ( .A(\SUBBYTES[4].a/w3089 ), .B(
        \SUBBYTES[4].a/w3096 ), .Z(n10144) );
  XOR \SUBBYTES[4].a/U4949  ( .A(n10146), .B(n10145), .Z(n10832) );
  XOR \SUBBYTES[4].a/U4948  ( .A(\w1[4][9] ), .B(n10147), .Z(n10145) );
  XOR \SUBBYTES[4].a/U4947  ( .A(\SUBBYTES[4].a/w3114 ), .B(\w1[4][13] ), .Z(
        n10146) );
  XOR \SUBBYTES[4].a/U4946  ( .A(\SUBBYTES[4].a/w3090 ), .B(
        \SUBBYTES[4].a/w3097 ), .Z(n10147) );
  XOR \SUBBYTES[4].a/U4945  ( .A(n10834), .B(n10832), .Z(\SUBBYTES[4].a/w3120 ) );
  XOR \SUBBYTES[4].a/U4944  ( .A(\w1[4][13] ), .B(n10148), .Z(n10835) );
  XOR \SUBBYTES[4].a/U4943  ( .A(\SUBBYTES[4].a/w3082 ), .B(
        \SUBBYTES[4].a/w3092 ), .Z(n10148) );
  XOR \SUBBYTES[4].a/U4942  ( .A(n10150), .B(n10149), .Z(\SUBBYTES[4].a/w3107 ) );
  XOR \SUBBYTES[4].a/U4941  ( .A(n10835), .B(n10151), .Z(n10149) );
  XOR \SUBBYTES[4].a/U4940  ( .A(\w1[4][12] ), .B(\SUBBYTES[4].a/w3171 ), .Z(
        n10150) );
  XOR \SUBBYTES[4].a/U4939  ( .A(\SUBBYTES[4].a/w3084 ), .B(
        \SUBBYTES[4].a/w3089 ), .Z(n10151) );
  XOR \SUBBYTES[4].a/U4938  ( .A(n10153), .B(n10152), .Z(n10833) );
  XOR \SUBBYTES[4].a/U4937  ( .A(\SUBBYTES[4].a/w3117 ), .B(\w1[4][15] ), .Z(
        n10152) );
  XOR \SUBBYTES[4].a/U4936  ( .A(\SUBBYTES[4].a/w3092 ), .B(
        \SUBBYTES[4].a/w3099 ), .Z(n10153) );
  XOR \SUBBYTES[4].a/U4935  ( .A(n10832), .B(n10833), .Z(\SUBBYTES[4].a/w3119 ) );
  XOR \SUBBYTES[4].a/U4934  ( .A(\w1[4][11] ), .B(n10154), .Z(n10836) );
  XOR \SUBBYTES[4].a/U4933  ( .A(\SUBBYTES[4].a/w3081 ), .B(
        \SUBBYTES[4].a/w3084 ), .Z(n10154) );
  XOR \SUBBYTES[4].a/U4932  ( .A(n10156), .B(n10155), .Z(\SUBBYTES[4].a/w3108 ) );
  XOR \SUBBYTES[4].a/U4931  ( .A(n10836), .B(n10157), .Z(n10155) );
  XOR \SUBBYTES[4].a/U4930  ( .A(\w1[4][14] ), .B(\SUBBYTES[4].a/w3150 ), .Z(
        n10156) );
  XOR \SUBBYTES[4].a/U4929  ( .A(\SUBBYTES[4].a/w3089 ), .B(
        \SUBBYTES[4].a/w3090 ), .Z(n10157) );
  XOR \SUBBYTES[4].a/U4928  ( .A(n10834), .B(n10833), .Z(\SUBBYTES[4].a/w3128 ) );
  XOR \SUBBYTES[4].a/U4927  ( .A(n10159), .B(n10158), .Z(\SUBBYTES[4].a/w3129 ) );
  XOR \SUBBYTES[4].a/U4926  ( .A(\w1[4][15] ), .B(n10835), .Z(n10158) );
  XOR \SUBBYTES[4].a/U4925  ( .A(\SUBBYTES[4].a/w3081 ), .B(
        \SUBBYTES[4].a/w3090 ), .Z(n10159) );
  XOR \SUBBYTES[4].a/U4924  ( .A(n10161), .B(n10160), .Z(\SUBBYTES[4].a/w3105 ) );
  XOR \SUBBYTES[4].a/U4923  ( .A(n10163), .B(n10162), .Z(n10160) );
  XOR \SUBBYTES[4].a/U4922  ( .A(\w1[4][15] ), .B(\SUBBYTES[4].a/w3189 ), .Z(
        n10161) );
  XOR \SUBBYTES[4].a/U4921  ( .A(\SUBBYTES[4].a/w3096 ), .B(
        \SUBBYTES[4].a/w3099 ), .Z(n10162) );
  XOR \SUBBYTES[4].a/U4920  ( .A(\SUBBYTES[4].a/w3082 ), .B(
        \SUBBYTES[4].a/w3084 ), .Z(n10163) );
  XOR \SUBBYTES[4].a/U4919  ( .A(n10165), .B(n10164), .Z(\SUBBYTES[4].a/w3106 ) );
  XOR \SUBBYTES[4].a/U4918  ( .A(n10836), .B(n10166), .Z(n10164) );
  XOR \SUBBYTES[4].a/U4917  ( .A(\w1[4][13] ), .B(n10837), .Z(n10165) );
  XOR \SUBBYTES[4].a/U4916  ( .A(\SUBBYTES[4].a/w3096 ), .B(
        \SUBBYTES[4].a/w3097 ), .Z(n10166) );
  XOR \SUBBYTES[4].a/U4915  ( .A(n10168), .B(n10167), .Z(\SUBBYTES[4].a/w3122 ) );
  XOR \SUBBYTES[4].a/U4914  ( .A(\w1[4][9] ), .B(n10169), .Z(n10167) );
  XOR \SUBBYTES[4].a/U4913  ( .A(\SUBBYTES[4].a/w3097 ), .B(
        \SUBBYTES[4].a/w3099 ), .Z(n10168) );
  XOR \SUBBYTES[4].a/U4912  ( .A(\SUBBYTES[4].a/w3081 ), .B(
        \SUBBYTES[4].a/w3082 ), .Z(n10169) );
  XOR \SUBBYTES[4].a/U4911  ( .A(\w1[4][17] ), .B(n10170), .Z(n10838) );
  XOR \SUBBYTES[4].a/U4910  ( .A(\w1[4][19] ), .B(\w1[4][18] ), .Z(n10170) );
  XOR \SUBBYTES[4].a/U4909  ( .A(\w1[4][22] ), .B(n10838), .Z(
        \SUBBYTES[4].a/w2964 ) );
  XOR \SUBBYTES[4].a/U4908  ( .A(\w1[4][16] ), .B(\SUBBYTES[4].a/w2964 ), .Z(
        \SUBBYTES[4].a/w2851 ) );
  XOR \SUBBYTES[4].a/U4907  ( .A(\w1[4][16] ), .B(n10171), .Z(
        \SUBBYTES[4].a/w2852 ) );
  XOR \SUBBYTES[4].a/U4906  ( .A(\w1[4][22] ), .B(\w1[4][21] ), .Z(n10171) );
  XOR \SUBBYTES[4].a/U4905  ( .A(\w1[4][21] ), .B(n10838), .Z(
        \SUBBYTES[4].a/w2982 ) );
  XOR \SUBBYTES[4].a/U4904  ( .A(n10173), .B(n10172), .Z(\SUBBYTES[4].a/w2975 ) );
  XOR \SUBBYTES[4].a/U4903  ( .A(\w1[4][19] ), .B(\w1[4][17] ), .Z(n10172) );
  XOR \SUBBYTES[4].a/U4902  ( .A(\w1[4][23] ), .B(\w1[4][20] ), .Z(n10173) );
  XOR \SUBBYTES[4].a/U4901  ( .A(\w1[4][16] ), .B(\SUBBYTES[4].a/w2975 ), .Z(
        \SUBBYTES[4].a/w2854 ) );
  XOR \SUBBYTES[4].a/U4900  ( .A(n10175), .B(n10174), .Z(\SUBBYTES[4].a/w2962 ) );
  XOR \SUBBYTES[4].a/U4899  ( .A(\SUBBYTES[4].a/w2923 ), .B(n1018), .Z(n10174)
         );
  XOR \SUBBYTES[4].a/U4898  ( .A(\SUBBYTES[4].a/w2916 ), .B(
        \SUBBYTES[4].a/w2919 ), .Z(n10175) );
  XOR \SUBBYTES[4].a/U4897  ( .A(n10177), .B(n10176), .Z(\SUBBYTES[4].a/w2963 ) );
  XOR \SUBBYTES[4].a/U4896  ( .A(\SUBBYTES[4].a/w2923 ), .B(n9699), .Z(n10176)
         );
  XOR \SUBBYTES[4].a/U4895  ( .A(\SUBBYTES[4].a/w2916 ), .B(n9698), .Z(n10177)
         );
  XOR \SUBBYTES[4].a/U4894  ( .A(\SUBBYTES[4].a/w2975 ), .B(n10178), .Z(
        \SUBBYTES[4].a/w2965 ) );
  XOR \SUBBYTES[4].a/U4893  ( .A(\w1[4][22] ), .B(\w1[4][21] ), .Z(n10178) );
  XOR \SUBBYTES[4].a/U4892  ( .A(n10180), .B(n10179), .Z(\SUBBYTES[4].a/w2966 ) );
  XOR \SUBBYTES[4].a/U4891  ( .A(n9699), .B(n1018), .Z(n10179) );
  XOR \SUBBYTES[4].a/U4890  ( .A(n9698), .B(\SUBBYTES[4].a/w2919 ), .Z(n10180)
         );
  XOR \SUBBYTES[4].a/U4889  ( .A(\w1[4][23] ), .B(\w1[4][18] ), .Z(n10844) );
  XOR \SUBBYTES[4].a/U4888  ( .A(n10844), .B(n10181), .Z(\SUBBYTES[4].a/w2967 ) );
  XOR \SUBBYTES[4].a/U4887  ( .A(\w1[4][21] ), .B(\w1[4][20] ), .Z(n10181) );
  XOR \SUBBYTES[4].a/U4886  ( .A(\w1[4][23] ), .B(\SUBBYTES[4].a/w2852 ), .Z(
        \SUBBYTES[4].a/w2855 ) );
  XOR \SUBBYTES[4].a/U4885  ( .A(\w1[4][17] ), .B(\SUBBYTES[4].a/w2852 ), .Z(
        \SUBBYTES[4].a/w2856 ) );
  XOR \SUBBYTES[4].a/U4884  ( .A(\w1[4][20] ), .B(\SUBBYTES[4].a/w2852 ), .Z(
        \SUBBYTES[4].a/w2857 ) );
  XOR \SUBBYTES[4].a/U4883  ( .A(\SUBBYTES[4].a/w2856 ), .B(n10844), .Z(
        \SUBBYTES[4].a/w2858 ) );
  XOR \SUBBYTES[4].a/U4882  ( .A(n10844), .B(n10182), .Z(\SUBBYTES[4].a/w2943 ) );
  XOR \SUBBYTES[4].a/U4881  ( .A(\w1[4][20] ), .B(\w1[4][17] ), .Z(n10182) );
  XOR \SUBBYTES[4].a/U4880  ( .A(n10184), .B(n10183), .Z(n10841) );
  XOR \SUBBYTES[4].a/U4879  ( .A(\w1[4][20] ), .B(n10185), .Z(n10183) );
  XOR \SUBBYTES[4].a/U4878  ( .A(\SUBBYTES[4].a/w2908 ), .B(\w1[4][22] ), .Z(
        n10184) );
  XOR \SUBBYTES[4].a/U4877  ( .A(\SUBBYTES[4].a/w2882 ), .B(
        \SUBBYTES[4].a/w2889 ), .Z(n10185) );
  XOR \SUBBYTES[4].a/U4876  ( .A(n10187), .B(n10186), .Z(n10839) );
  XOR \SUBBYTES[4].a/U4875  ( .A(\w1[4][17] ), .B(n10188), .Z(n10186) );
  XOR \SUBBYTES[4].a/U4874  ( .A(\SUBBYTES[4].a/w2907 ), .B(\w1[4][21] ), .Z(
        n10187) );
  XOR \SUBBYTES[4].a/U4873  ( .A(\SUBBYTES[4].a/w2883 ), .B(
        \SUBBYTES[4].a/w2890 ), .Z(n10188) );
  XOR \SUBBYTES[4].a/U4872  ( .A(n10841), .B(n10839), .Z(\SUBBYTES[4].a/w2913 ) );
  XOR \SUBBYTES[4].a/U4871  ( .A(\w1[4][21] ), .B(n10189), .Z(n10842) );
  XOR \SUBBYTES[4].a/U4870  ( .A(\SUBBYTES[4].a/w2875 ), .B(
        \SUBBYTES[4].a/w2885 ), .Z(n10189) );
  XOR \SUBBYTES[4].a/U4869  ( .A(n10191), .B(n10190), .Z(\SUBBYTES[4].a/w2900 ) );
  XOR \SUBBYTES[4].a/U4868  ( .A(n10842), .B(n10192), .Z(n10190) );
  XOR \SUBBYTES[4].a/U4867  ( .A(\w1[4][20] ), .B(\SUBBYTES[4].a/w2964 ), .Z(
        n10191) );
  XOR \SUBBYTES[4].a/U4866  ( .A(\SUBBYTES[4].a/w2877 ), .B(
        \SUBBYTES[4].a/w2882 ), .Z(n10192) );
  XOR \SUBBYTES[4].a/U4865  ( .A(n10194), .B(n10193), .Z(n10840) );
  XOR \SUBBYTES[4].a/U4864  ( .A(\SUBBYTES[4].a/w2910 ), .B(\w1[4][23] ), .Z(
        n10193) );
  XOR \SUBBYTES[4].a/U4863  ( .A(\SUBBYTES[4].a/w2885 ), .B(
        \SUBBYTES[4].a/w2892 ), .Z(n10194) );
  XOR \SUBBYTES[4].a/U4862  ( .A(n10839), .B(n10840), .Z(\SUBBYTES[4].a/w2912 ) );
  XOR \SUBBYTES[4].a/U4861  ( .A(\w1[4][19] ), .B(n10195), .Z(n10843) );
  XOR \SUBBYTES[4].a/U4860  ( .A(\SUBBYTES[4].a/w2874 ), .B(
        \SUBBYTES[4].a/w2877 ), .Z(n10195) );
  XOR \SUBBYTES[4].a/U4859  ( .A(n10197), .B(n10196), .Z(\SUBBYTES[4].a/w2901 ) );
  XOR \SUBBYTES[4].a/U4858  ( .A(n10843), .B(n10198), .Z(n10196) );
  XOR \SUBBYTES[4].a/U4857  ( .A(\w1[4][22] ), .B(\SUBBYTES[4].a/w2943 ), .Z(
        n10197) );
  XOR \SUBBYTES[4].a/U4856  ( .A(\SUBBYTES[4].a/w2882 ), .B(
        \SUBBYTES[4].a/w2883 ), .Z(n10198) );
  XOR \SUBBYTES[4].a/U4855  ( .A(n10841), .B(n10840), .Z(\SUBBYTES[4].a/w2921 ) );
  XOR \SUBBYTES[4].a/U4854  ( .A(n10200), .B(n10199), .Z(\SUBBYTES[4].a/w2922 ) );
  XOR \SUBBYTES[4].a/U4853  ( .A(\w1[4][23] ), .B(n10842), .Z(n10199) );
  XOR \SUBBYTES[4].a/U4852  ( .A(\SUBBYTES[4].a/w2874 ), .B(
        \SUBBYTES[4].a/w2883 ), .Z(n10200) );
  XOR \SUBBYTES[4].a/U4851  ( .A(n10202), .B(n10201), .Z(\SUBBYTES[4].a/w2898 ) );
  XOR \SUBBYTES[4].a/U4850  ( .A(n10204), .B(n10203), .Z(n10201) );
  XOR \SUBBYTES[4].a/U4849  ( .A(\w1[4][23] ), .B(\SUBBYTES[4].a/w2982 ), .Z(
        n10202) );
  XOR \SUBBYTES[4].a/U4848  ( .A(\SUBBYTES[4].a/w2889 ), .B(
        \SUBBYTES[4].a/w2892 ), .Z(n10203) );
  XOR \SUBBYTES[4].a/U4847  ( .A(\SUBBYTES[4].a/w2875 ), .B(
        \SUBBYTES[4].a/w2877 ), .Z(n10204) );
  XOR \SUBBYTES[4].a/U4846  ( .A(n10206), .B(n10205), .Z(\SUBBYTES[4].a/w2899 ) );
  XOR \SUBBYTES[4].a/U4845  ( .A(n10843), .B(n10207), .Z(n10205) );
  XOR \SUBBYTES[4].a/U4844  ( .A(\w1[4][21] ), .B(n10844), .Z(n10206) );
  XOR \SUBBYTES[4].a/U4843  ( .A(\SUBBYTES[4].a/w2889 ), .B(
        \SUBBYTES[4].a/w2890 ), .Z(n10207) );
  XOR \SUBBYTES[4].a/U4842  ( .A(n10209), .B(n10208), .Z(\SUBBYTES[4].a/w2915 ) );
  XOR \SUBBYTES[4].a/U4841  ( .A(\w1[4][17] ), .B(n10210), .Z(n10208) );
  XOR \SUBBYTES[4].a/U4840  ( .A(\SUBBYTES[4].a/w2890 ), .B(
        \SUBBYTES[4].a/w2892 ), .Z(n10209) );
  XOR \SUBBYTES[4].a/U4839  ( .A(\SUBBYTES[4].a/w2874 ), .B(
        \SUBBYTES[4].a/w2875 ), .Z(n10210) );
  XOR \SUBBYTES[4].a/U4838  ( .A(\w1[4][25] ), .B(n10211), .Z(n10845) );
  XOR \SUBBYTES[4].a/U4837  ( .A(\w1[4][27] ), .B(\w1[4][26] ), .Z(n10211) );
  XOR \SUBBYTES[4].a/U4836  ( .A(\w1[4][30] ), .B(n10845), .Z(
        \SUBBYTES[4].a/w2757 ) );
  XOR \SUBBYTES[4].a/U4835  ( .A(\w1[4][24] ), .B(\SUBBYTES[4].a/w2757 ), .Z(
        \SUBBYTES[4].a/w2644 ) );
  XOR \SUBBYTES[4].a/U4834  ( .A(\w1[4][24] ), .B(n10212), .Z(
        \SUBBYTES[4].a/w2645 ) );
  XOR \SUBBYTES[4].a/U4833  ( .A(\w1[4][30] ), .B(\w1[4][29] ), .Z(n10212) );
  XOR \SUBBYTES[4].a/U4832  ( .A(\w1[4][29] ), .B(n10845), .Z(
        \SUBBYTES[4].a/w2775 ) );
  XOR \SUBBYTES[4].a/U4831  ( .A(n10214), .B(n10213), .Z(\SUBBYTES[4].a/w2768 ) );
  XOR \SUBBYTES[4].a/U4830  ( .A(\w1[4][27] ), .B(\w1[4][25] ), .Z(n10213) );
  XOR \SUBBYTES[4].a/U4829  ( .A(\w1[4][31] ), .B(\w1[4][28] ), .Z(n10214) );
  XOR \SUBBYTES[4].a/U4828  ( .A(\w1[4][24] ), .B(\SUBBYTES[4].a/w2768 ), .Z(
        \SUBBYTES[4].a/w2647 ) );
  XOR \SUBBYTES[4].a/U4827  ( .A(n10216), .B(n10215), .Z(\SUBBYTES[4].a/w2755 ) );
  XOR \SUBBYTES[4].a/U4826  ( .A(\SUBBYTES[4].a/w2716 ), .B(n1017), .Z(n10215)
         );
  XOR \SUBBYTES[4].a/U4825  ( .A(\SUBBYTES[4].a/w2709 ), .B(
        \SUBBYTES[4].a/w2712 ), .Z(n10216) );
  XOR \SUBBYTES[4].a/U4824  ( .A(n10218), .B(n10217), .Z(\SUBBYTES[4].a/w2756 ) );
  XOR \SUBBYTES[4].a/U4823  ( .A(\SUBBYTES[4].a/w2716 ), .B(n9697), .Z(n10217)
         );
  XOR \SUBBYTES[4].a/U4822  ( .A(\SUBBYTES[4].a/w2709 ), .B(n9696), .Z(n10218)
         );
  XOR \SUBBYTES[4].a/U4821  ( .A(\SUBBYTES[4].a/w2768 ), .B(n10219), .Z(
        \SUBBYTES[4].a/w2758 ) );
  XOR \SUBBYTES[4].a/U4820  ( .A(\w1[4][30] ), .B(\w1[4][29] ), .Z(n10219) );
  XOR \SUBBYTES[4].a/U4819  ( .A(n10221), .B(n10220), .Z(\SUBBYTES[4].a/w2759 ) );
  XOR \SUBBYTES[4].a/U4818  ( .A(n9697), .B(n1017), .Z(n10220) );
  XOR \SUBBYTES[4].a/U4817  ( .A(n9696), .B(\SUBBYTES[4].a/w2712 ), .Z(n10221)
         );
  XOR \SUBBYTES[4].a/U4816  ( .A(\w1[4][31] ), .B(\w1[4][26] ), .Z(n10851) );
  XOR \SUBBYTES[4].a/U4815  ( .A(n10851), .B(n10222), .Z(\SUBBYTES[4].a/w2760 ) );
  XOR \SUBBYTES[4].a/U4814  ( .A(\w1[4][29] ), .B(\w1[4][28] ), .Z(n10222) );
  XOR \SUBBYTES[4].a/U4813  ( .A(\w1[4][31] ), .B(\SUBBYTES[4].a/w2645 ), .Z(
        \SUBBYTES[4].a/w2648 ) );
  XOR \SUBBYTES[4].a/U4812  ( .A(\w1[4][25] ), .B(\SUBBYTES[4].a/w2645 ), .Z(
        \SUBBYTES[4].a/w2649 ) );
  XOR \SUBBYTES[4].a/U4811  ( .A(\w1[4][28] ), .B(\SUBBYTES[4].a/w2645 ), .Z(
        \SUBBYTES[4].a/w2650 ) );
  XOR \SUBBYTES[4].a/U4810  ( .A(\SUBBYTES[4].a/w2649 ), .B(n10851), .Z(
        \SUBBYTES[4].a/w2651 ) );
  XOR \SUBBYTES[4].a/U4809  ( .A(n10851), .B(n10223), .Z(\SUBBYTES[4].a/w2736 ) );
  XOR \SUBBYTES[4].a/U4808  ( .A(\w1[4][28] ), .B(\w1[4][25] ), .Z(n10223) );
  XOR \SUBBYTES[4].a/U4807  ( .A(n10225), .B(n10224), .Z(n10848) );
  XOR \SUBBYTES[4].a/U4806  ( .A(\w1[4][28] ), .B(n10226), .Z(n10224) );
  XOR \SUBBYTES[4].a/U4805  ( .A(\SUBBYTES[4].a/w2701 ), .B(\w1[4][30] ), .Z(
        n10225) );
  XOR \SUBBYTES[4].a/U4804  ( .A(\SUBBYTES[4].a/w2675 ), .B(
        \SUBBYTES[4].a/w2682 ), .Z(n10226) );
  XOR \SUBBYTES[4].a/U4803  ( .A(n10228), .B(n10227), .Z(n10846) );
  XOR \SUBBYTES[4].a/U4802  ( .A(\w1[4][25] ), .B(n10229), .Z(n10227) );
  XOR \SUBBYTES[4].a/U4801  ( .A(\SUBBYTES[4].a/w2700 ), .B(\w1[4][29] ), .Z(
        n10228) );
  XOR \SUBBYTES[4].a/U4800  ( .A(\SUBBYTES[4].a/w2676 ), .B(
        \SUBBYTES[4].a/w2683 ), .Z(n10229) );
  XOR \SUBBYTES[4].a/U4799  ( .A(n10848), .B(n10846), .Z(\SUBBYTES[4].a/w2706 ) );
  XOR \SUBBYTES[4].a/U4798  ( .A(\w1[4][29] ), .B(n10230), .Z(n10849) );
  XOR \SUBBYTES[4].a/U4797  ( .A(\SUBBYTES[4].a/w2668 ), .B(
        \SUBBYTES[4].a/w2678 ), .Z(n10230) );
  XOR \SUBBYTES[4].a/U4796  ( .A(n10232), .B(n10231), .Z(\SUBBYTES[4].a/w2693 ) );
  XOR \SUBBYTES[4].a/U4795  ( .A(n10849), .B(n10233), .Z(n10231) );
  XOR \SUBBYTES[4].a/U4794  ( .A(\w1[4][28] ), .B(\SUBBYTES[4].a/w2757 ), .Z(
        n10232) );
  XOR \SUBBYTES[4].a/U4793  ( .A(\SUBBYTES[4].a/w2670 ), .B(
        \SUBBYTES[4].a/w2675 ), .Z(n10233) );
  XOR \SUBBYTES[4].a/U4792  ( .A(n10235), .B(n10234), .Z(n10847) );
  XOR \SUBBYTES[4].a/U4791  ( .A(\SUBBYTES[4].a/w2703 ), .B(\w1[4][31] ), .Z(
        n10234) );
  XOR \SUBBYTES[4].a/U4790  ( .A(\SUBBYTES[4].a/w2678 ), .B(
        \SUBBYTES[4].a/w2685 ), .Z(n10235) );
  XOR \SUBBYTES[4].a/U4789  ( .A(n10846), .B(n10847), .Z(\SUBBYTES[4].a/w2705 ) );
  XOR \SUBBYTES[4].a/U4788  ( .A(\w1[4][27] ), .B(n10236), .Z(n10850) );
  XOR \SUBBYTES[4].a/U4787  ( .A(\SUBBYTES[4].a/w2667 ), .B(
        \SUBBYTES[4].a/w2670 ), .Z(n10236) );
  XOR \SUBBYTES[4].a/U4786  ( .A(n10238), .B(n10237), .Z(\SUBBYTES[4].a/w2694 ) );
  XOR \SUBBYTES[4].a/U4785  ( .A(n10850), .B(n10239), .Z(n10237) );
  XOR \SUBBYTES[4].a/U4784  ( .A(\w1[4][30] ), .B(\SUBBYTES[4].a/w2736 ), .Z(
        n10238) );
  XOR \SUBBYTES[4].a/U4783  ( .A(\SUBBYTES[4].a/w2675 ), .B(
        \SUBBYTES[4].a/w2676 ), .Z(n10239) );
  XOR \SUBBYTES[4].a/U4782  ( .A(n10848), .B(n10847), .Z(\SUBBYTES[4].a/w2714 ) );
  XOR \SUBBYTES[4].a/U4781  ( .A(n10241), .B(n10240), .Z(\SUBBYTES[4].a/w2715 ) );
  XOR \SUBBYTES[4].a/U4780  ( .A(\w1[4][31] ), .B(n10849), .Z(n10240) );
  XOR \SUBBYTES[4].a/U4779  ( .A(\SUBBYTES[4].a/w2667 ), .B(
        \SUBBYTES[4].a/w2676 ), .Z(n10241) );
  XOR \SUBBYTES[4].a/U4778  ( .A(n10243), .B(n10242), .Z(\SUBBYTES[4].a/w2691 ) );
  XOR \SUBBYTES[4].a/U4777  ( .A(n10245), .B(n10244), .Z(n10242) );
  XOR \SUBBYTES[4].a/U4776  ( .A(\w1[4][31] ), .B(\SUBBYTES[4].a/w2775 ), .Z(
        n10243) );
  XOR \SUBBYTES[4].a/U4775  ( .A(\SUBBYTES[4].a/w2682 ), .B(
        \SUBBYTES[4].a/w2685 ), .Z(n10244) );
  XOR \SUBBYTES[4].a/U4774  ( .A(\SUBBYTES[4].a/w2668 ), .B(
        \SUBBYTES[4].a/w2670 ), .Z(n10245) );
  XOR \SUBBYTES[4].a/U4773  ( .A(n10247), .B(n10246), .Z(\SUBBYTES[4].a/w2692 ) );
  XOR \SUBBYTES[4].a/U4772  ( .A(n10850), .B(n10248), .Z(n10246) );
  XOR \SUBBYTES[4].a/U4771  ( .A(\w1[4][29] ), .B(n10851), .Z(n10247) );
  XOR \SUBBYTES[4].a/U4770  ( .A(\SUBBYTES[4].a/w2682 ), .B(
        \SUBBYTES[4].a/w2683 ), .Z(n10248) );
  XOR \SUBBYTES[4].a/U4769  ( .A(n10250), .B(n10249), .Z(\SUBBYTES[4].a/w2708 ) );
  XOR \SUBBYTES[4].a/U4768  ( .A(\w1[4][25] ), .B(n10251), .Z(n10249) );
  XOR \SUBBYTES[4].a/U4767  ( .A(\SUBBYTES[4].a/w2683 ), .B(
        \SUBBYTES[4].a/w2685 ), .Z(n10250) );
  XOR \SUBBYTES[4].a/U4766  ( .A(\SUBBYTES[4].a/w2667 ), .B(
        \SUBBYTES[4].a/w2668 ), .Z(n10251) );
  XOR \SUBBYTES[4].a/U4765  ( .A(\w1[4][33] ), .B(n10252), .Z(n10852) );
  XOR \SUBBYTES[4].a/U4764  ( .A(\w1[4][35] ), .B(\w1[4][34] ), .Z(n10252) );
  XOR \SUBBYTES[4].a/U4763  ( .A(\w1[4][38] ), .B(n10852), .Z(
        \SUBBYTES[4].a/w2550 ) );
  XOR \SUBBYTES[4].a/U4762  ( .A(\w1[4][32] ), .B(\SUBBYTES[4].a/w2550 ), .Z(
        \SUBBYTES[4].a/w2437 ) );
  XOR \SUBBYTES[4].a/U4761  ( .A(\w1[4][32] ), .B(n10253), .Z(
        \SUBBYTES[4].a/w2438 ) );
  XOR \SUBBYTES[4].a/U4760  ( .A(\w1[4][38] ), .B(\w1[4][37] ), .Z(n10253) );
  XOR \SUBBYTES[4].a/U4759  ( .A(\w1[4][37] ), .B(n10852), .Z(
        \SUBBYTES[4].a/w2568 ) );
  XOR \SUBBYTES[4].a/U4758  ( .A(n10255), .B(n10254), .Z(\SUBBYTES[4].a/w2561 ) );
  XOR \SUBBYTES[4].a/U4757  ( .A(\w1[4][35] ), .B(\w1[4][33] ), .Z(n10254) );
  XOR \SUBBYTES[4].a/U4756  ( .A(\w1[4][39] ), .B(\w1[4][36] ), .Z(n10255) );
  XOR \SUBBYTES[4].a/U4755  ( .A(\w1[4][32] ), .B(\SUBBYTES[4].a/w2561 ), .Z(
        \SUBBYTES[4].a/w2440 ) );
  XOR \SUBBYTES[4].a/U4754  ( .A(n10257), .B(n10256), .Z(\SUBBYTES[4].a/w2548 ) );
  XOR \SUBBYTES[4].a/U4753  ( .A(\SUBBYTES[4].a/w2509 ), .B(n1016), .Z(n10256)
         );
  XOR \SUBBYTES[4].a/U4752  ( .A(\SUBBYTES[4].a/w2502 ), .B(
        \SUBBYTES[4].a/w2505 ), .Z(n10257) );
  XOR \SUBBYTES[4].a/U4751  ( .A(n10259), .B(n10258), .Z(\SUBBYTES[4].a/w2549 ) );
  XOR \SUBBYTES[4].a/U4750  ( .A(\SUBBYTES[4].a/w2509 ), .B(n9695), .Z(n10258)
         );
  XOR \SUBBYTES[4].a/U4749  ( .A(\SUBBYTES[4].a/w2502 ), .B(n9694), .Z(n10259)
         );
  XOR \SUBBYTES[4].a/U4748  ( .A(\SUBBYTES[4].a/w2561 ), .B(n10260), .Z(
        \SUBBYTES[4].a/w2551 ) );
  XOR \SUBBYTES[4].a/U4747  ( .A(\w1[4][38] ), .B(\w1[4][37] ), .Z(n10260) );
  XOR \SUBBYTES[4].a/U4746  ( .A(n10262), .B(n10261), .Z(\SUBBYTES[4].a/w2552 ) );
  XOR \SUBBYTES[4].a/U4745  ( .A(n9695), .B(n1016), .Z(n10261) );
  XOR \SUBBYTES[4].a/U4744  ( .A(n9694), .B(\SUBBYTES[4].a/w2505 ), .Z(n10262)
         );
  XOR \SUBBYTES[4].a/U4743  ( .A(\w1[4][39] ), .B(\w1[4][34] ), .Z(n10858) );
  XOR \SUBBYTES[4].a/U4742  ( .A(n10858), .B(n10263), .Z(\SUBBYTES[4].a/w2553 ) );
  XOR \SUBBYTES[4].a/U4741  ( .A(\w1[4][37] ), .B(\w1[4][36] ), .Z(n10263) );
  XOR \SUBBYTES[4].a/U4740  ( .A(\w1[4][39] ), .B(\SUBBYTES[4].a/w2438 ), .Z(
        \SUBBYTES[4].a/w2441 ) );
  XOR \SUBBYTES[4].a/U4739  ( .A(\w1[4][33] ), .B(\SUBBYTES[4].a/w2438 ), .Z(
        \SUBBYTES[4].a/w2442 ) );
  XOR \SUBBYTES[4].a/U4738  ( .A(\w1[4][36] ), .B(\SUBBYTES[4].a/w2438 ), .Z(
        \SUBBYTES[4].a/w2443 ) );
  XOR \SUBBYTES[4].a/U4737  ( .A(\SUBBYTES[4].a/w2442 ), .B(n10858), .Z(
        \SUBBYTES[4].a/w2444 ) );
  XOR \SUBBYTES[4].a/U4736  ( .A(n10858), .B(n10264), .Z(\SUBBYTES[4].a/w2529 ) );
  XOR \SUBBYTES[4].a/U4735  ( .A(\w1[4][36] ), .B(\w1[4][33] ), .Z(n10264) );
  XOR \SUBBYTES[4].a/U4734  ( .A(n10266), .B(n10265), .Z(n10855) );
  XOR \SUBBYTES[4].a/U4733  ( .A(\w1[4][36] ), .B(n10267), .Z(n10265) );
  XOR \SUBBYTES[4].a/U4732  ( .A(\SUBBYTES[4].a/w2494 ), .B(\w1[4][38] ), .Z(
        n10266) );
  XOR \SUBBYTES[4].a/U4731  ( .A(\SUBBYTES[4].a/w2468 ), .B(
        \SUBBYTES[4].a/w2475 ), .Z(n10267) );
  XOR \SUBBYTES[4].a/U4730  ( .A(n10269), .B(n10268), .Z(n10853) );
  XOR \SUBBYTES[4].a/U4729  ( .A(\w1[4][33] ), .B(n10270), .Z(n10268) );
  XOR \SUBBYTES[4].a/U4728  ( .A(\SUBBYTES[4].a/w2493 ), .B(\w1[4][37] ), .Z(
        n10269) );
  XOR \SUBBYTES[4].a/U4727  ( .A(\SUBBYTES[4].a/w2469 ), .B(
        \SUBBYTES[4].a/w2476 ), .Z(n10270) );
  XOR \SUBBYTES[4].a/U4726  ( .A(n10855), .B(n10853), .Z(\SUBBYTES[4].a/w2499 ) );
  XOR \SUBBYTES[4].a/U4725  ( .A(\w1[4][37] ), .B(n10271), .Z(n10856) );
  XOR \SUBBYTES[4].a/U4724  ( .A(\SUBBYTES[4].a/w2461 ), .B(
        \SUBBYTES[4].a/w2471 ), .Z(n10271) );
  XOR \SUBBYTES[4].a/U4723  ( .A(n10273), .B(n10272), .Z(\SUBBYTES[4].a/w2486 ) );
  XOR \SUBBYTES[4].a/U4722  ( .A(n10856), .B(n10274), .Z(n10272) );
  XOR \SUBBYTES[4].a/U4721  ( .A(\w1[4][36] ), .B(\SUBBYTES[4].a/w2550 ), .Z(
        n10273) );
  XOR \SUBBYTES[4].a/U4720  ( .A(\SUBBYTES[4].a/w2463 ), .B(
        \SUBBYTES[4].a/w2468 ), .Z(n10274) );
  XOR \SUBBYTES[4].a/U4719  ( .A(n10276), .B(n10275), .Z(n10854) );
  XOR \SUBBYTES[4].a/U4718  ( .A(\SUBBYTES[4].a/w2496 ), .B(\w1[4][39] ), .Z(
        n10275) );
  XOR \SUBBYTES[4].a/U4717  ( .A(\SUBBYTES[4].a/w2471 ), .B(
        \SUBBYTES[4].a/w2478 ), .Z(n10276) );
  XOR \SUBBYTES[4].a/U4716  ( .A(n10853), .B(n10854), .Z(\SUBBYTES[4].a/w2498 ) );
  XOR \SUBBYTES[4].a/U4715  ( .A(\w1[4][35] ), .B(n10277), .Z(n10857) );
  XOR \SUBBYTES[4].a/U4714  ( .A(\SUBBYTES[4].a/w2460 ), .B(
        \SUBBYTES[4].a/w2463 ), .Z(n10277) );
  XOR \SUBBYTES[4].a/U4713  ( .A(n10279), .B(n10278), .Z(\SUBBYTES[4].a/w2487 ) );
  XOR \SUBBYTES[4].a/U4712  ( .A(n10857), .B(n10280), .Z(n10278) );
  XOR \SUBBYTES[4].a/U4711  ( .A(\w1[4][38] ), .B(\SUBBYTES[4].a/w2529 ), .Z(
        n10279) );
  XOR \SUBBYTES[4].a/U4710  ( .A(\SUBBYTES[4].a/w2468 ), .B(
        \SUBBYTES[4].a/w2469 ), .Z(n10280) );
  XOR \SUBBYTES[4].a/U4709  ( .A(n10855), .B(n10854), .Z(\SUBBYTES[4].a/w2507 ) );
  XOR \SUBBYTES[4].a/U4708  ( .A(n10282), .B(n10281), .Z(\SUBBYTES[4].a/w2508 ) );
  XOR \SUBBYTES[4].a/U4707  ( .A(\w1[4][39] ), .B(n10856), .Z(n10281) );
  XOR \SUBBYTES[4].a/U4706  ( .A(\SUBBYTES[4].a/w2460 ), .B(
        \SUBBYTES[4].a/w2469 ), .Z(n10282) );
  XOR \SUBBYTES[4].a/U4705  ( .A(n10284), .B(n10283), .Z(\SUBBYTES[4].a/w2484 ) );
  XOR \SUBBYTES[4].a/U4704  ( .A(n10286), .B(n10285), .Z(n10283) );
  XOR \SUBBYTES[4].a/U4703  ( .A(\w1[4][39] ), .B(\SUBBYTES[4].a/w2568 ), .Z(
        n10284) );
  XOR \SUBBYTES[4].a/U4702  ( .A(\SUBBYTES[4].a/w2475 ), .B(
        \SUBBYTES[4].a/w2478 ), .Z(n10285) );
  XOR \SUBBYTES[4].a/U4701  ( .A(\SUBBYTES[4].a/w2461 ), .B(
        \SUBBYTES[4].a/w2463 ), .Z(n10286) );
  XOR \SUBBYTES[4].a/U4700  ( .A(n10288), .B(n10287), .Z(\SUBBYTES[4].a/w2485 ) );
  XOR \SUBBYTES[4].a/U4699  ( .A(n10857), .B(n10289), .Z(n10287) );
  XOR \SUBBYTES[4].a/U4698  ( .A(\w1[4][37] ), .B(n10858), .Z(n10288) );
  XOR \SUBBYTES[4].a/U4697  ( .A(\SUBBYTES[4].a/w2475 ), .B(
        \SUBBYTES[4].a/w2476 ), .Z(n10289) );
  XOR \SUBBYTES[4].a/U4696  ( .A(n10291), .B(n10290), .Z(\SUBBYTES[4].a/w2501 ) );
  XOR \SUBBYTES[4].a/U4695  ( .A(\w1[4][33] ), .B(n10292), .Z(n10290) );
  XOR \SUBBYTES[4].a/U4694  ( .A(\SUBBYTES[4].a/w2476 ), .B(
        \SUBBYTES[4].a/w2478 ), .Z(n10291) );
  XOR \SUBBYTES[4].a/U4693  ( .A(\SUBBYTES[4].a/w2460 ), .B(
        \SUBBYTES[4].a/w2461 ), .Z(n10292) );
  XOR \SUBBYTES[4].a/U4692  ( .A(\w1[4][41] ), .B(n10293), .Z(n10859) );
  XOR \SUBBYTES[4].a/U4691  ( .A(\w1[4][43] ), .B(\w1[4][42] ), .Z(n10293) );
  XOR \SUBBYTES[4].a/U4690  ( .A(\w1[4][46] ), .B(n10859), .Z(
        \SUBBYTES[4].a/w2343 ) );
  XOR \SUBBYTES[4].a/U4689  ( .A(\w1[4][40] ), .B(\SUBBYTES[4].a/w2343 ), .Z(
        \SUBBYTES[4].a/w2230 ) );
  XOR \SUBBYTES[4].a/U4688  ( .A(\w1[4][40] ), .B(n10294), .Z(
        \SUBBYTES[4].a/w2231 ) );
  XOR \SUBBYTES[4].a/U4687  ( .A(\w1[4][46] ), .B(\w1[4][45] ), .Z(n10294) );
  XOR \SUBBYTES[4].a/U4686  ( .A(\w1[4][45] ), .B(n10859), .Z(
        \SUBBYTES[4].a/w2361 ) );
  XOR \SUBBYTES[4].a/U4685  ( .A(n10296), .B(n10295), .Z(\SUBBYTES[4].a/w2354 ) );
  XOR \SUBBYTES[4].a/U4684  ( .A(\w1[4][43] ), .B(\w1[4][41] ), .Z(n10295) );
  XOR \SUBBYTES[4].a/U4683  ( .A(\w1[4][47] ), .B(\w1[4][44] ), .Z(n10296) );
  XOR \SUBBYTES[4].a/U4682  ( .A(\w1[4][40] ), .B(\SUBBYTES[4].a/w2354 ), .Z(
        \SUBBYTES[4].a/w2233 ) );
  XOR \SUBBYTES[4].a/U4681  ( .A(n10298), .B(n10297), .Z(\SUBBYTES[4].a/w2341 ) );
  XOR \SUBBYTES[4].a/U4680  ( .A(\SUBBYTES[4].a/w2302 ), .B(n1015), .Z(n10297)
         );
  XOR \SUBBYTES[4].a/U4679  ( .A(\SUBBYTES[4].a/w2295 ), .B(
        \SUBBYTES[4].a/w2298 ), .Z(n10298) );
  XOR \SUBBYTES[4].a/U4678  ( .A(n10300), .B(n10299), .Z(\SUBBYTES[4].a/w2342 ) );
  XOR \SUBBYTES[4].a/U4677  ( .A(\SUBBYTES[4].a/w2302 ), .B(n9693), .Z(n10299)
         );
  XOR \SUBBYTES[4].a/U4676  ( .A(\SUBBYTES[4].a/w2295 ), .B(n9692), .Z(n10300)
         );
  XOR \SUBBYTES[4].a/U4675  ( .A(\SUBBYTES[4].a/w2354 ), .B(n10301), .Z(
        \SUBBYTES[4].a/w2344 ) );
  XOR \SUBBYTES[4].a/U4674  ( .A(\w1[4][46] ), .B(\w1[4][45] ), .Z(n10301) );
  XOR \SUBBYTES[4].a/U4673  ( .A(n10303), .B(n10302), .Z(\SUBBYTES[4].a/w2345 ) );
  XOR \SUBBYTES[4].a/U4672  ( .A(n9693), .B(n1015), .Z(n10302) );
  XOR \SUBBYTES[4].a/U4671  ( .A(n9692), .B(\SUBBYTES[4].a/w2298 ), .Z(n10303)
         );
  XOR \SUBBYTES[4].a/U4670  ( .A(\w1[4][47] ), .B(\w1[4][42] ), .Z(n10865) );
  XOR \SUBBYTES[4].a/U4669  ( .A(n10865), .B(n10304), .Z(\SUBBYTES[4].a/w2346 ) );
  XOR \SUBBYTES[4].a/U4668  ( .A(\w1[4][45] ), .B(\w1[4][44] ), .Z(n10304) );
  XOR \SUBBYTES[4].a/U4667  ( .A(\w1[4][47] ), .B(\SUBBYTES[4].a/w2231 ), .Z(
        \SUBBYTES[4].a/w2234 ) );
  XOR \SUBBYTES[4].a/U4666  ( .A(\w1[4][41] ), .B(\SUBBYTES[4].a/w2231 ), .Z(
        \SUBBYTES[4].a/w2235 ) );
  XOR \SUBBYTES[4].a/U4665  ( .A(\w1[4][44] ), .B(\SUBBYTES[4].a/w2231 ), .Z(
        \SUBBYTES[4].a/w2236 ) );
  XOR \SUBBYTES[4].a/U4664  ( .A(\SUBBYTES[4].a/w2235 ), .B(n10865), .Z(
        \SUBBYTES[4].a/w2237 ) );
  XOR \SUBBYTES[4].a/U4663  ( .A(n10865), .B(n10305), .Z(\SUBBYTES[4].a/w2322 ) );
  XOR \SUBBYTES[4].a/U4662  ( .A(\w1[4][44] ), .B(\w1[4][41] ), .Z(n10305) );
  XOR \SUBBYTES[4].a/U4661  ( .A(n10307), .B(n10306), .Z(n10862) );
  XOR \SUBBYTES[4].a/U4660  ( .A(\w1[4][44] ), .B(n10308), .Z(n10306) );
  XOR \SUBBYTES[4].a/U4659  ( .A(\SUBBYTES[4].a/w2287 ), .B(\w1[4][46] ), .Z(
        n10307) );
  XOR \SUBBYTES[4].a/U4658  ( .A(\SUBBYTES[4].a/w2261 ), .B(
        \SUBBYTES[4].a/w2268 ), .Z(n10308) );
  XOR \SUBBYTES[4].a/U4657  ( .A(n10310), .B(n10309), .Z(n10860) );
  XOR \SUBBYTES[4].a/U4656  ( .A(\w1[4][41] ), .B(n10311), .Z(n10309) );
  XOR \SUBBYTES[4].a/U4655  ( .A(\SUBBYTES[4].a/w2286 ), .B(\w1[4][45] ), .Z(
        n10310) );
  XOR \SUBBYTES[4].a/U4654  ( .A(\SUBBYTES[4].a/w2262 ), .B(
        \SUBBYTES[4].a/w2269 ), .Z(n10311) );
  XOR \SUBBYTES[4].a/U4653  ( .A(n10862), .B(n10860), .Z(\SUBBYTES[4].a/w2292 ) );
  XOR \SUBBYTES[4].a/U4652  ( .A(\w1[4][45] ), .B(n10312), .Z(n10863) );
  XOR \SUBBYTES[4].a/U4651  ( .A(\SUBBYTES[4].a/w2254 ), .B(
        \SUBBYTES[4].a/w2264 ), .Z(n10312) );
  XOR \SUBBYTES[4].a/U4650  ( .A(n10314), .B(n10313), .Z(\SUBBYTES[4].a/w2279 ) );
  XOR \SUBBYTES[4].a/U4649  ( .A(n10863), .B(n10315), .Z(n10313) );
  XOR \SUBBYTES[4].a/U4648  ( .A(\w1[4][44] ), .B(\SUBBYTES[4].a/w2343 ), .Z(
        n10314) );
  XOR \SUBBYTES[4].a/U4647  ( .A(\SUBBYTES[4].a/w2256 ), .B(
        \SUBBYTES[4].a/w2261 ), .Z(n10315) );
  XOR \SUBBYTES[4].a/U4646  ( .A(n10317), .B(n10316), .Z(n10861) );
  XOR \SUBBYTES[4].a/U4645  ( .A(\SUBBYTES[4].a/w2289 ), .B(\w1[4][47] ), .Z(
        n10316) );
  XOR \SUBBYTES[4].a/U4644  ( .A(\SUBBYTES[4].a/w2264 ), .B(
        \SUBBYTES[4].a/w2271 ), .Z(n10317) );
  XOR \SUBBYTES[4].a/U4643  ( .A(n10860), .B(n10861), .Z(\SUBBYTES[4].a/w2291 ) );
  XOR \SUBBYTES[4].a/U4642  ( .A(\w1[4][43] ), .B(n10318), .Z(n10864) );
  XOR \SUBBYTES[4].a/U4641  ( .A(\SUBBYTES[4].a/w2253 ), .B(
        \SUBBYTES[4].a/w2256 ), .Z(n10318) );
  XOR \SUBBYTES[4].a/U4640  ( .A(n10320), .B(n10319), .Z(\SUBBYTES[4].a/w2280 ) );
  XOR \SUBBYTES[4].a/U4639  ( .A(n10864), .B(n10321), .Z(n10319) );
  XOR \SUBBYTES[4].a/U4638  ( .A(\w1[4][46] ), .B(\SUBBYTES[4].a/w2322 ), .Z(
        n10320) );
  XOR \SUBBYTES[4].a/U4637  ( .A(\SUBBYTES[4].a/w2261 ), .B(
        \SUBBYTES[4].a/w2262 ), .Z(n10321) );
  XOR \SUBBYTES[4].a/U4636  ( .A(n10862), .B(n10861), .Z(\SUBBYTES[4].a/w2300 ) );
  XOR \SUBBYTES[4].a/U4635  ( .A(n10323), .B(n10322), .Z(\SUBBYTES[4].a/w2301 ) );
  XOR \SUBBYTES[4].a/U4634  ( .A(\w1[4][47] ), .B(n10863), .Z(n10322) );
  XOR \SUBBYTES[4].a/U4633  ( .A(\SUBBYTES[4].a/w2253 ), .B(
        \SUBBYTES[4].a/w2262 ), .Z(n10323) );
  XOR \SUBBYTES[4].a/U4632  ( .A(n10325), .B(n10324), .Z(\SUBBYTES[4].a/w2277 ) );
  XOR \SUBBYTES[4].a/U4631  ( .A(n10327), .B(n10326), .Z(n10324) );
  XOR \SUBBYTES[4].a/U4630  ( .A(\w1[4][47] ), .B(\SUBBYTES[4].a/w2361 ), .Z(
        n10325) );
  XOR \SUBBYTES[4].a/U4629  ( .A(\SUBBYTES[4].a/w2268 ), .B(
        \SUBBYTES[4].a/w2271 ), .Z(n10326) );
  XOR \SUBBYTES[4].a/U4628  ( .A(\SUBBYTES[4].a/w2254 ), .B(
        \SUBBYTES[4].a/w2256 ), .Z(n10327) );
  XOR \SUBBYTES[4].a/U4627  ( .A(n10329), .B(n10328), .Z(\SUBBYTES[4].a/w2278 ) );
  XOR \SUBBYTES[4].a/U4626  ( .A(n10864), .B(n10330), .Z(n10328) );
  XOR \SUBBYTES[4].a/U4625  ( .A(\w1[4][45] ), .B(n10865), .Z(n10329) );
  XOR \SUBBYTES[4].a/U4624  ( .A(\SUBBYTES[4].a/w2268 ), .B(
        \SUBBYTES[4].a/w2269 ), .Z(n10330) );
  XOR \SUBBYTES[4].a/U4623  ( .A(n10332), .B(n10331), .Z(\SUBBYTES[4].a/w2294 ) );
  XOR \SUBBYTES[4].a/U4622  ( .A(\w1[4][41] ), .B(n10333), .Z(n10331) );
  XOR \SUBBYTES[4].a/U4621  ( .A(\SUBBYTES[4].a/w2269 ), .B(
        \SUBBYTES[4].a/w2271 ), .Z(n10332) );
  XOR \SUBBYTES[4].a/U4620  ( .A(\SUBBYTES[4].a/w2253 ), .B(
        \SUBBYTES[4].a/w2254 ), .Z(n10333) );
  XOR \SUBBYTES[4].a/U4619  ( .A(\w1[4][49] ), .B(n10334), .Z(n10866) );
  XOR \SUBBYTES[4].a/U4618  ( .A(\w1[4][51] ), .B(\w1[4][50] ), .Z(n10334) );
  XOR \SUBBYTES[4].a/U4617  ( .A(\w1[4][54] ), .B(n10866), .Z(
        \SUBBYTES[4].a/w2136 ) );
  XOR \SUBBYTES[4].a/U4616  ( .A(\w1[4][48] ), .B(\SUBBYTES[4].a/w2136 ), .Z(
        \SUBBYTES[4].a/w2023 ) );
  XOR \SUBBYTES[4].a/U4615  ( .A(\w1[4][48] ), .B(n10335), .Z(
        \SUBBYTES[4].a/w2024 ) );
  XOR \SUBBYTES[4].a/U4614  ( .A(\w1[4][54] ), .B(\w1[4][53] ), .Z(n10335) );
  XOR \SUBBYTES[4].a/U4613  ( .A(\w1[4][53] ), .B(n10866), .Z(
        \SUBBYTES[4].a/w2154 ) );
  XOR \SUBBYTES[4].a/U4612  ( .A(n10337), .B(n10336), .Z(\SUBBYTES[4].a/w2147 ) );
  XOR \SUBBYTES[4].a/U4611  ( .A(\w1[4][51] ), .B(\w1[4][49] ), .Z(n10336) );
  XOR \SUBBYTES[4].a/U4610  ( .A(\w1[4][55] ), .B(\w1[4][52] ), .Z(n10337) );
  XOR \SUBBYTES[4].a/U4609  ( .A(\w1[4][48] ), .B(\SUBBYTES[4].a/w2147 ), .Z(
        \SUBBYTES[4].a/w2026 ) );
  XOR \SUBBYTES[4].a/U4608  ( .A(n10339), .B(n10338), .Z(\SUBBYTES[4].a/w2134 ) );
  XOR \SUBBYTES[4].a/U4607  ( .A(\SUBBYTES[4].a/w2095 ), .B(n1014), .Z(n10338)
         );
  XOR \SUBBYTES[4].a/U4606  ( .A(\SUBBYTES[4].a/w2088 ), .B(
        \SUBBYTES[4].a/w2091 ), .Z(n10339) );
  XOR \SUBBYTES[4].a/U4605  ( .A(n10341), .B(n10340), .Z(\SUBBYTES[4].a/w2135 ) );
  XOR \SUBBYTES[4].a/U4604  ( .A(\SUBBYTES[4].a/w2095 ), .B(n9691), .Z(n10340)
         );
  XOR \SUBBYTES[4].a/U4603  ( .A(\SUBBYTES[4].a/w2088 ), .B(n9690), .Z(n10341)
         );
  XOR \SUBBYTES[4].a/U4602  ( .A(\SUBBYTES[4].a/w2147 ), .B(n10342), .Z(
        \SUBBYTES[4].a/w2137 ) );
  XOR \SUBBYTES[4].a/U4601  ( .A(\w1[4][54] ), .B(\w1[4][53] ), .Z(n10342) );
  XOR \SUBBYTES[4].a/U4600  ( .A(n10344), .B(n10343), .Z(\SUBBYTES[4].a/w2138 ) );
  XOR \SUBBYTES[4].a/U4599  ( .A(n9691), .B(n1014), .Z(n10343) );
  XOR \SUBBYTES[4].a/U4598  ( .A(n9690), .B(\SUBBYTES[4].a/w2091 ), .Z(n10344)
         );
  XOR \SUBBYTES[4].a/U4597  ( .A(\w1[4][55] ), .B(\w1[4][50] ), .Z(n10872) );
  XOR \SUBBYTES[4].a/U4596  ( .A(n10872), .B(n10345), .Z(\SUBBYTES[4].a/w2139 ) );
  XOR \SUBBYTES[4].a/U4595  ( .A(\w1[4][53] ), .B(\w1[4][52] ), .Z(n10345) );
  XOR \SUBBYTES[4].a/U4594  ( .A(\w1[4][55] ), .B(\SUBBYTES[4].a/w2024 ), .Z(
        \SUBBYTES[4].a/w2027 ) );
  XOR \SUBBYTES[4].a/U4593  ( .A(\w1[4][49] ), .B(\SUBBYTES[4].a/w2024 ), .Z(
        \SUBBYTES[4].a/w2028 ) );
  XOR \SUBBYTES[4].a/U4592  ( .A(\w1[4][52] ), .B(\SUBBYTES[4].a/w2024 ), .Z(
        \SUBBYTES[4].a/w2029 ) );
  XOR \SUBBYTES[4].a/U4591  ( .A(\SUBBYTES[4].a/w2028 ), .B(n10872), .Z(
        \SUBBYTES[4].a/w2030 ) );
  XOR \SUBBYTES[4].a/U4590  ( .A(n10872), .B(n10346), .Z(\SUBBYTES[4].a/w2115 ) );
  XOR \SUBBYTES[4].a/U4589  ( .A(\w1[4][52] ), .B(\w1[4][49] ), .Z(n10346) );
  XOR \SUBBYTES[4].a/U4588  ( .A(n10348), .B(n10347), .Z(n10869) );
  XOR \SUBBYTES[4].a/U4587  ( .A(\w1[4][52] ), .B(n10349), .Z(n10347) );
  XOR \SUBBYTES[4].a/U4586  ( .A(\SUBBYTES[4].a/w2080 ), .B(\w1[4][54] ), .Z(
        n10348) );
  XOR \SUBBYTES[4].a/U4585  ( .A(\SUBBYTES[4].a/w2054 ), .B(
        \SUBBYTES[4].a/w2061 ), .Z(n10349) );
  XOR \SUBBYTES[4].a/U4584  ( .A(n10351), .B(n10350), .Z(n10867) );
  XOR \SUBBYTES[4].a/U4583  ( .A(\w1[4][49] ), .B(n10352), .Z(n10350) );
  XOR \SUBBYTES[4].a/U4582  ( .A(\SUBBYTES[4].a/w2079 ), .B(\w1[4][53] ), .Z(
        n10351) );
  XOR \SUBBYTES[4].a/U4581  ( .A(\SUBBYTES[4].a/w2055 ), .B(
        \SUBBYTES[4].a/w2062 ), .Z(n10352) );
  XOR \SUBBYTES[4].a/U4580  ( .A(n10869), .B(n10867), .Z(\SUBBYTES[4].a/w2085 ) );
  XOR \SUBBYTES[4].a/U4579  ( .A(\w1[4][53] ), .B(n10353), .Z(n10870) );
  XOR \SUBBYTES[4].a/U4578  ( .A(\SUBBYTES[4].a/w2047 ), .B(
        \SUBBYTES[4].a/w2057 ), .Z(n10353) );
  XOR \SUBBYTES[4].a/U4577  ( .A(n10355), .B(n10354), .Z(\SUBBYTES[4].a/w2072 ) );
  XOR \SUBBYTES[4].a/U4576  ( .A(n10870), .B(n10356), .Z(n10354) );
  XOR \SUBBYTES[4].a/U4575  ( .A(\w1[4][52] ), .B(\SUBBYTES[4].a/w2136 ), .Z(
        n10355) );
  XOR \SUBBYTES[4].a/U4574  ( .A(\SUBBYTES[4].a/w2049 ), .B(
        \SUBBYTES[4].a/w2054 ), .Z(n10356) );
  XOR \SUBBYTES[4].a/U4573  ( .A(n10358), .B(n10357), .Z(n10868) );
  XOR \SUBBYTES[4].a/U4572  ( .A(\SUBBYTES[4].a/w2082 ), .B(\w1[4][55] ), .Z(
        n10357) );
  XOR \SUBBYTES[4].a/U4571  ( .A(\SUBBYTES[4].a/w2057 ), .B(
        \SUBBYTES[4].a/w2064 ), .Z(n10358) );
  XOR \SUBBYTES[4].a/U4570  ( .A(n10867), .B(n10868), .Z(\SUBBYTES[4].a/w2084 ) );
  XOR \SUBBYTES[4].a/U4569  ( .A(\w1[4][51] ), .B(n10359), .Z(n10871) );
  XOR \SUBBYTES[4].a/U4568  ( .A(\SUBBYTES[4].a/w2046 ), .B(
        \SUBBYTES[4].a/w2049 ), .Z(n10359) );
  XOR \SUBBYTES[4].a/U4567  ( .A(n10361), .B(n10360), .Z(\SUBBYTES[4].a/w2073 ) );
  XOR \SUBBYTES[4].a/U4566  ( .A(n10871), .B(n10362), .Z(n10360) );
  XOR \SUBBYTES[4].a/U4565  ( .A(\w1[4][54] ), .B(\SUBBYTES[4].a/w2115 ), .Z(
        n10361) );
  XOR \SUBBYTES[4].a/U4564  ( .A(\SUBBYTES[4].a/w2054 ), .B(
        \SUBBYTES[4].a/w2055 ), .Z(n10362) );
  XOR \SUBBYTES[4].a/U4563  ( .A(n10869), .B(n10868), .Z(\SUBBYTES[4].a/w2093 ) );
  XOR \SUBBYTES[4].a/U4562  ( .A(n10364), .B(n10363), .Z(\SUBBYTES[4].a/w2094 ) );
  XOR \SUBBYTES[4].a/U4561  ( .A(\w1[4][55] ), .B(n10870), .Z(n10363) );
  XOR \SUBBYTES[4].a/U4560  ( .A(\SUBBYTES[4].a/w2046 ), .B(
        \SUBBYTES[4].a/w2055 ), .Z(n10364) );
  XOR \SUBBYTES[4].a/U4559  ( .A(n10366), .B(n10365), .Z(\SUBBYTES[4].a/w2070 ) );
  XOR \SUBBYTES[4].a/U4558  ( .A(n10368), .B(n10367), .Z(n10365) );
  XOR \SUBBYTES[4].a/U4557  ( .A(\w1[4][55] ), .B(\SUBBYTES[4].a/w2154 ), .Z(
        n10366) );
  XOR \SUBBYTES[4].a/U4556  ( .A(\SUBBYTES[4].a/w2061 ), .B(
        \SUBBYTES[4].a/w2064 ), .Z(n10367) );
  XOR \SUBBYTES[4].a/U4555  ( .A(\SUBBYTES[4].a/w2047 ), .B(
        \SUBBYTES[4].a/w2049 ), .Z(n10368) );
  XOR \SUBBYTES[4].a/U4554  ( .A(n10370), .B(n10369), .Z(\SUBBYTES[4].a/w2071 ) );
  XOR \SUBBYTES[4].a/U4553  ( .A(n10871), .B(n10371), .Z(n10369) );
  XOR \SUBBYTES[4].a/U4552  ( .A(\w1[4][53] ), .B(n10872), .Z(n10370) );
  XOR \SUBBYTES[4].a/U4551  ( .A(\SUBBYTES[4].a/w2061 ), .B(
        \SUBBYTES[4].a/w2062 ), .Z(n10371) );
  XOR \SUBBYTES[4].a/U4550  ( .A(n10373), .B(n10372), .Z(\SUBBYTES[4].a/w2087 ) );
  XOR \SUBBYTES[4].a/U4549  ( .A(\w1[4][49] ), .B(n10374), .Z(n10372) );
  XOR \SUBBYTES[4].a/U4548  ( .A(\SUBBYTES[4].a/w2062 ), .B(
        \SUBBYTES[4].a/w2064 ), .Z(n10373) );
  XOR \SUBBYTES[4].a/U4547  ( .A(\SUBBYTES[4].a/w2046 ), .B(
        \SUBBYTES[4].a/w2047 ), .Z(n10374) );
  XOR \SUBBYTES[4].a/U4546  ( .A(\w1[4][57] ), .B(n10375), .Z(n10873) );
  XOR \SUBBYTES[4].a/U4545  ( .A(\w1[4][59] ), .B(\w1[4][58] ), .Z(n10375) );
  XOR \SUBBYTES[4].a/U4544  ( .A(\w1[4][62] ), .B(n10873), .Z(
        \SUBBYTES[4].a/w1929 ) );
  XOR \SUBBYTES[4].a/U4543  ( .A(\w1[4][56] ), .B(\SUBBYTES[4].a/w1929 ), .Z(
        \SUBBYTES[4].a/w1816 ) );
  XOR \SUBBYTES[4].a/U4542  ( .A(\w1[4][56] ), .B(n10376), .Z(
        \SUBBYTES[4].a/w1817 ) );
  XOR \SUBBYTES[4].a/U4541  ( .A(\w1[4][62] ), .B(\w1[4][61] ), .Z(n10376) );
  XOR \SUBBYTES[4].a/U4540  ( .A(\w1[4][61] ), .B(n10873), .Z(
        \SUBBYTES[4].a/w1947 ) );
  XOR \SUBBYTES[4].a/U4539  ( .A(n10378), .B(n10377), .Z(\SUBBYTES[4].a/w1940 ) );
  XOR \SUBBYTES[4].a/U4538  ( .A(\w1[4][59] ), .B(\w1[4][57] ), .Z(n10377) );
  XOR \SUBBYTES[4].a/U4537  ( .A(\w1[4][63] ), .B(\w1[4][60] ), .Z(n10378) );
  XOR \SUBBYTES[4].a/U4536  ( .A(\w1[4][56] ), .B(\SUBBYTES[4].a/w1940 ), .Z(
        \SUBBYTES[4].a/w1819 ) );
  XOR \SUBBYTES[4].a/U4535  ( .A(n10380), .B(n10379), .Z(\SUBBYTES[4].a/w1927 ) );
  XOR \SUBBYTES[4].a/U4534  ( .A(\SUBBYTES[4].a/w1888 ), .B(n1013), .Z(n10379)
         );
  XOR \SUBBYTES[4].a/U4533  ( .A(\SUBBYTES[4].a/w1881 ), .B(
        \SUBBYTES[4].a/w1884 ), .Z(n10380) );
  XOR \SUBBYTES[4].a/U4532  ( .A(n10382), .B(n10381), .Z(\SUBBYTES[4].a/w1928 ) );
  XOR \SUBBYTES[4].a/U4531  ( .A(\SUBBYTES[4].a/w1888 ), .B(n9689), .Z(n10381)
         );
  XOR \SUBBYTES[4].a/U4530  ( .A(\SUBBYTES[4].a/w1881 ), .B(n9688), .Z(n10382)
         );
  XOR \SUBBYTES[4].a/U4529  ( .A(\SUBBYTES[4].a/w1940 ), .B(n10383), .Z(
        \SUBBYTES[4].a/w1930 ) );
  XOR \SUBBYTES[4].a/U4528  ( .A(\w1[4][62] ), .B(\w1[4][61] ), .Z(n10383) );
  XOR \SUBBYTES[4].a/U4527  ( .A(n10385), .B(n10384), .Z(\SUBBYTES[4].a/w1931 ) );
  XOR \SUBBYTES[4].a/U4526  ( .A(n9689), .B(n1013), .Z(n10384) );
  XOR \SUBBYTES[4].a/U4525  ( .A(n9688), .B(\SUBBYTES[4].a/w1884 ), .Z(n10385)
         );
  XOR \SUBBYTES[4].a/U4524  ( .A(\w1[4][63] ), .B(\w1[4][58] ), .Z(n10879) );
  XOR \SUBBYTES[4].a/U4523  ( .A(n10879), .B(n10386), .Z(\SUBBYTES[4].a/w1932 ) );
  XOR \SUBBYTES[4].a/U4522  ( .A(\w1[4][61] ), .B(\w1[4][60] ), .Z(n10386) );
  XOR \SUBBYTES[4].a/U4521  ( .A(\w1[4][63] ), .B(\SUBBYTES[4].a/w1817 ), .Z(
        \SUBBYTES[4].a/w1820 ) );
  XOR \SUBBYTES[4].a/U4520  ( .A(\w1[4][57] ), .B(\SUBBYTES[4].a/w1817 ), .Z(
        \SUBBYTES[4].a/w1821 ) );
  XOR \SUBBYTES[4].a/U4519  ( .A(\w1[4][60] ), .B(\SUBBYTES[4].a/w1817 ), .Z(
        \SUBBYTES[4].a/w1822 ) );
  XOR \SUBBYTES[4].a/U4518  ( .A(\SUBBYTES[4].a/w1821 ), .B(n10879), .Z(
        \SUBBYTES[4].a/w1823 ) );
  XOR \SUBBYTES[4].a/U4517  ( .A(n10879), .B(n10387), .Z(\SUBBYTES[4].a/w1908 ) );
  XOR \SUBBYTES[4].a/U4516  ( .A(\w1[4][60] ), .B(\w1[4][57] ), .Z(n10387) );
  XOR \SUBBYTES[4].a/U4515  ( .A(n10389), .B(n10388), .Z(n10876) );
  XOR \SUBBYTES[4].a/U4514  ( .A(\w1[4][60] ), .B(n10390), .Z(n10388) );
  XOR \SUBBYTES[4].a/U4513  ( .A(\SUBBYTES[4].a/w1873 ), .B(\w1[4][62] ), .Z(
        n10389) );
  XOR \SUBBYTES[4].a/U4512  ( .A(\SUBBYTES[4].a/w1847 ), .B(
        \SUBBYTES[4].a/w1854 ), .Z(n10390) );
  XOR \SUBBYTES[4].a/U4511  ( .A(n10392), .B(n10391), .Z(n10874) );
  XOR \SUBBYTES[4].a/U4510  ( .A(\w1[4][57] ), .B(n10393), .Z(n10391) );
  XOR \SUBBYTES[4].a/U4509  ( .A(\SUBBYTES[4].a/w1872 ), .B(\w1[4][61] ), .Z(
        n10392) );
  XOR \SUBBYTES[4].a/U4508  ( .A(\SUBBYTES[4].a/w1848 ), .B(
        \SUBBYTES[4].a/w1855 ), .Z(n10393) );
  XOR \SUBBYTES[4].a/U4507  ( .A(n10876), .B(n10874), .Z(\SUBBYTES[4].a/w1878 ) );
  XOR \SUBBYTES[4].a/U4506  ( .A(\w1[4][61] ), .B(n10394), .Z(n10877) );
  XOR \SUBBYTES[4].a/U4505  ( .A(\SUBBYTES[4].a/w1840 ), .B(
        \SUBBYTES[4].a/w1850 ), .Z(n10394) );
  XOR \SUBBYTES[4].a/U4504  ( .A(n10396), .B(n10395), .Z(\SUBBYTES[4].a/w1865 ) );
  XOR \SUBBYTES[4].a/U4503  ( .A(n10877), .B(n10397), .Z(n10395) );
  XOR \SUBBYTES[4].a/U4502  ( .A(\w1[4][60] ), .B(\SUBBYTES[4].a/w1929 ), .Z(
        n10396) );
  XOR \SUBBYTES[4].a/U4501  ( .A(\SUBBYTES[4].a/w1842 ), .B(
        \SUBBYTES[4].a/w1847 ), .Z(n10397) );
  XOR \SUBBYTES[4].a/U4500  ( .A(n10399), .B(n10398), .Z(n10875) );
  XOR \SUBBYTES[4].a/U4499  ( .A(\SUBBYTES[4].a/w1875 ), .B(\w1[4][63] ), .Z(
        n10398) );
  XOR \SUBBYTES[4].a/U4498  ( .A(\SUBBYTES[4].a/w1850 ), .B(
        \SUBBYTES[4].a/w1857 ), .Z(n10399) );
  XOR \SUBBYTES[4].a/U4497  ( .A(n10874), .B(n10875), .Z(\SUBBYTES[4].a/w1877 ) );
  XOR \SUBBYTES[4].a/U4496  ( .A(\w1[4][59] ), .B(n10400), .Z(n10878) );
  XOR \SUBBYTES[4].a/U4495  ( .A(\SUBBYTES[4].a/w1839 ), .B(
        \SUBBYTES[4].a/w1842 ), .Z(n10400) );
  XOR \SUBBYTES[4].a/U4494  ( .A(n10402), .B(n10401), .Z(\SUBBYTES[4].a/w1866 ) );
  XOR \SUBBYTES[4].a/U4493  ( .A(n10878), .B(n10403), .Z(n10401) );
  XOR \SUBBYTES[4].a/U4492  ( .A(\w1[4][62] ), .B(\SUBBYTES[4].a/w1908 ), .Z(
        n10402) );
  XOR \SUBBYTES[4].a/U4491  ( .A(\SUBBYTES[4].a/w1847 ), .B(
        \SUBBYTES[4].a/w1848 ), .Z(n10403) );
  XOR \SUBBYTES[4].a/U4490  ( .A(n10876), .B(n10875), .Z(\SUBBYTES[4].a/w1886 ) );
  XOR \SUBBYTES[4].a/U4489  ( .A(n10405), .B(n10404), .Z(\SUBBYTES[4].a/w1887 ) );
  XOR \SUBBYTES[4].a/U4488  ( .A(\w1[4][63] ), .B(n10877), .Z(n10404) );
  XOR \SUBBYTES[4].a/U4487  ( .A(\SUBBYTES[4].a/w1839 ), .B(
        \SUBBYTES[4].a/w1848 ), .Z(n10405) );
  XOR \SUBBYTES[4].a/U4486  ( .A(n10407), .B(n10406), .Z(\SUBBYTES[4].a/w1863 ) );
  XOR \SUBBYTES[4].a/U4485  ( .A(n10409), .B(n10408), .Z(n10406) );
  XOR \SUBBYTES[4].a/U4484  ( .A(\w1[4][63] ), .B(\SUBBYTES[4].a/w1947 ), .Z(
        n10407) );
  XOR \SUBBYTES[4].a/U4483  ( .A(\SUBBYTES[4].a/w1854 ), .B(
        \SUBBYTES[4].a/w1857 ), .Z(n10408) );
  XOR \SUBBYTES[4].a/U4482  ( .A(\SUBBYTES[4].a/w1840 ), .B(
        \SUBBYTES[4].a/w1842 ), .Z(n10409) );
  XOR \SUBBYTES[4].a/U4481  ( .A(n10411), .B(n10410), .Z(\SUBBYTES[4].a/w1864 ) );
  XOR \SUBBYTES[4].a/U4480  ( .A(n10878), .B(n10412), .Z(n10410) );
  XOR \SUBBYTES[4].a/U4479  ( .A(\w1[4][61] ), .B(n10879), .Z(n10411) );
  XOR \SUBBYTES[4].a/U4478  ( .A(\SUBBYTES[4].a/w1854 ), .B(
        \SUBBYTES[4].a/w1855 ), .Z(n10412) );
  XOR \SUBBYTES[4].a/U4477  ( .A(n10414), .B(n10413), .Z(\SUBBYTES[4].a/w1880 ) );
  XOR \SUBBYTES[4].a/U4476  ( .A(\w1[4][57] ), .B(n10415), .Z(n10413) );
  XOR \SUBBYTES[4].a/U4475  ( .A(\SUBBYTES[4].a/w1855 ), .B(
        \SUBBYTES[4].a/w1857 ), .Z(n10414) );
  XOR \SUBBYTES[4].a/U4474  ( .A(\SUBBYTES[4].a/w1839 ), .B(
        \SUBBYTES[4].a/w1840 ), .Z(n10415) );
  XOR \SUBBYTES[4].a/U4473  ( .A(\w1[4][65] ), .B(n10416), .Z(n10880) );
  XOR \SUBBYTES[4].a/U4472  ( .A(\w1[4][67] ), .B(\w1[4][66] ), .Z(n10416) );
  XOR \SUBBYTES[4].a/U4471  ( .A(\w1[4][70] ), .B(n10880), .Z(
        \SUBBYTES[4].a/w1722 ) );
  XOR \SUBBYTES[4].a/U4470  ( .A(\w1[4][64] ), .B(\SUBBYTES[4].a/w1722 ), .Z(
        \SUBBYTES[4].a/w1609 ) );
  XOR \SUBBYTES[4].a/U4469  ( .A(\w1[4][64] ), .B(n10417), .Z(
        \SUBBYTES[4].a/w1610 ) );
  XOR \SUBBYTES[4].a/U4468  ( .A(\w1[4][70] ), .B(\w1[4][69] ), .Z(n10417) );
  XOR \SUBBYTES[4].a/U4467  ( .A(\w1[4][69] ), .B(n10880), .Z(
        \SUBBYTES[4].a/w1740 ) );
  XOR \SUBBYTES[4].a/U4466  ( .A(n10419), .B(n10418), .Z(\SUBBYTES[4].a/w1733 ) );
  XOR \SUBBYTES[4].a/U4465  ( .A(\w1[4][67] ), .B(\w1[4][65] ), .Z(n10418) );
  XOR \SUBBYTES[4].a/U4464  ( .A(\w1[4][71] ), .B(\w1[4][68] ), .Z(n10419) );
  XOR \SUBBYTES[4].a/U4463  ( .A(\w1[4][64] ), .B(\SUBBYTES[4].a/w1733 ), .Z(
        \SUBBYTES[4].a/w1612 ) );
  XOR \SUBBYTES[4].a/U4462  ( .A(n10421), .B(n10420), .Z(\SUBBYTES[4].a/w1720 ) );
  XOR \SUBBYTES[4].a/U4461  ( .A(\SUBBYTES[4].a/w1681 ), .B(n1012), .Z(n10420)
         );
  XOR \SUBBYTES[4].a/U4460  ( .A(\SUBBYTES[4].a/w1674 ), .B(
        \SUBBYTES[4].a/w1677 ), .Z(n10421) );
  XOR \SUBBYTES[4].a/U4459  ( .A(n10423), .B(n10422), .Z(\SUBBYTES[4].a/w1721 ) );
  XOR \SUBBYTES[4].a/U4458  ( .A(\SUBBYTES[4].a/w1681 ), .B(n9687), .Z(n10422)
         );
  XOR \SUBBYTES[4].a/U4457  ( .A(\SUBBYTES[4].a/w1674 ), .B(n9686), .Z(n10423)
         );
  XOR \SUBBYTES[4].a/U4456  ( .A(\SUBBYTES[4].a/w1733 ), .B(n10424), .Z(
        \SUBBYTES[4].a/w1723 ) );
  XOR \SUBBYTES[4].a/U4455  ( .A(\w1[4][70] ), .B(\w1[4][69] ), .Z(n10424) );
  XOR \SUBBYTES[4].a/U4454  ( .A(n10426), .B(n10425), .Z(\SUBBYTES[4].a/w1724 ) );
  XOR \SUBBYTES[4].a/U4453  ( .A(n9687), .B(n1012), .Z(n10425) );
  XOR \SUBBYTES[4].a/U4452  ( .A(n9686), .B(\SUBBYTES[4].a/w1677 ), .Z(n10426)
         );
  XOR \SUBBYTES[4].a/U4451  ( .A(\w1[4][71] ), .B(\w1[4][66] ), .Z(n10886) );
  XOR \SUBBYTES[4].a/U4450  ( .A(n10886), .B(n10427), .Z(\SUBBYTES[4].a/w1725 ) );
  XOR \SUBBYTES[4].a/U4449  ( .A(\w1[4][69] ), .B(\w1[4][68] ), .Z(n10427) );
  XOR \SUBBYTES[4].a/U4448  ( .A(\w1[4][71] ), .B(\SUBBYTES[4].a/w1610 ), .Z(
        \SUBBYTES[4].a/w1613 ) );
  XOR \SUBBYTES[4].a/U4447  ( .A(\w1[4][65] ), .B(\SUBBYTES[4].a/w1610 ), .Z(
        \SUBBYTES[4].a/w1614 ) );
  XOR \SUBBYTES[4].a/U4446  ( .A(\w1[4][68] ), .B(\SUBBYTES[4].a/w1610 ), .Z(
        \SUBBYTES[4].a/w1615 ) );
  XOR \SUBBYTES[4].a/U4445  ( .A(\SUBBYTES[4].a/w1614 ), .B(n10886), .Z(
        \SUBBYTES[4].a/w1616 ) );
  XOR \SUBBYTES[4].a/U4444  ( .A(n10886), .B(n10428), .Z(\SUBBYTES[4].a/w1701 ) );
  XOR \SUBBYTES[4].a/U4443  ( .A(\w1[4][68] ), .B(\w1[4][65] ), .Z(n10428) );
  XOR \SUBBYTES[4].a/U4442  ( .A(n10430), .B(n10429), .Z(n10883) );
  XOR \SUBBYTES[4].a/U4441  ( .A(\w1[4][68] ), .B(n10431), .Z(n10429) );
  XOR \SUBBYTES[4].a/U4440  ( .A(\SUBBYTES[4].a/w1666 ), .B(\w1[4][70] ), .Z(
        n10430) );
  XOR \SUBBYTES[4].a/U4439  ( .A(\SUBBYTES[4].a/w1640 ), .B(
        \SUBBYTES[4].a/w1647 ), .Z(n10431) );
  XOR \SUBBYTES[4].a/U4438  ( .A(n10433), .B(n10432), .Z(n10881) );
  XOR \SUBBYTES[4].a/U4437  ( .A(\w1[4][65] ), .B(n10434), .Z(n10432) );
  XOR \SUBBYTES[4].a/U4436  ( .A(\SUBBYTES[4].a/w1665 ), .B(\w1[4][69] ), .Z(
        n10433) );
  XOR \SUBBYTES[4].a/U4435  ( .A(\SUBBYTES[4].a/w1641 ), .B(
        \SUBBYTES[4].a/w1648 ), .Z(n10434) );
  XOR \SUBBYTES[4].a/U4434  ( .A(n10883), .B(n10881), .Z(\SUBBYTES[4].a/w1671 ) );
  XOR \SUBBYTES[4].a/U4433  ( .A(\w1[4][69] ), .B(n10435), .Z(n10884) );
  XOR \SUBBYTES[4].a/U4432  ( .A(\SUBBYTES[4].a/w1633 ), .B(
        \SUBBYTES[4].a/w1643 ), .Z(n10435) );
  XOR \SUBBYTES[4].a/U4431  ( .A(n10437), .B(n10436), .Z(\SUBBYTES[4].a/w1658 ) );
  XOR \SUBBYTES[4].a/U4430  ( .A(n10884), .B(n10438), .Z(n10436) );
  XOR \SUBBYTES[4].a/U4429  ( .A(\w1[4][68] ), .B(\SUBBYTES[4].a/w1722 ), .Z(
        n10437) );
  XOR \SUBBYTES[4].a/U4428  ( .A(\SUBBYTES[4].a/w1635 ), .B(
        \SUBBYTES[4].a/w1640 ), .Z(n10438) );
  XOR \SUBBYTES[4].a/U4427  ( .A(n10440), .B(n10439), .Z(n10882) );
  XOR \SUBBYTES[4].a/U4426  ( .A(\SUBBYTES[4].a/w1668 ), .B(\w1[4][71] ), .Z(
        n10439) );
  XOR \SUBBYTES[4].a/U4425  ( .A(\SUBBYTES[4].a/w1643 ), .B(
        \SUBBYTES[4].a/w1650 ), .Z(n10440) );
  XOR \SUBBYTES[4].a/U4424  ( .A(n10881), .B(n10882), .Z(\SUBBYTES[4].a/w1670 ) );
  XOR \SUBBYTES[4].a/U4423  ( .A(\w1[4][67] ), .B(n10441), .Z(n10885) );
  XOR \SUBBYTES[4].a/U4422  ( .A(\SUBBYTES[4].a/w1632 ), .B(
        \SUBBYTES[4].a/w1635 ), .Z(n10441) );
  XOR \SUBBYTES[4].a/U4421  ( .A(n10443), .B(n10442), .Z(\SUBBYTES[4].a/w1659 ) );
  XOR \SUBBYTES[4].a/U4420  ( .A(n10885), .B(n10444), .Z(n10442) );
  XOR \SUBBYTES[4].a/U4419  ( .A(\w1[4][70] ), .B(\SUBBYTES[4].a/w1701 ), .Z(
        n10443) );
  XOR \SUBBYTES[4].a/U4418  ( .A(\SUBBYTES[4].a/w1640 ), .B(
        \SUBBYTES[4].a/w1641 ), .Z(n10444) );
  XOR \SUBBYTES[4].a/U4417  ( .A(n10883), .B(n10882), .Z(\SUBBYTES[4].a/w1679 ) );
  XOR \SUBBYTES[4].a/U4416  ( .A(n10446), .B(n10445), .Z(\SUBBYTES[4].a/w1680 ) );
  XOR \SUBBYTES[4].a/U4415  ( .A(\w1[4][71] ), .B(n10884), .Z(n10445) );
  XOR \SUBBYTES[4].a/U4414  ( .A(\SUBBYTES[4].a/w1632 ), .B(
        \SUBBYTES[4].a/w1641 ), .Z(n10446) );
  XOR \SUBBYTES[4].a/U4413  ( .A(n10448), .B(n10447), .Z(\SUBBYTES[4].a/w1656 ) );
  XOR \SUBBYTES[4].a/U4412  ( .A(n10450), .B(n10449), .Z(n10447) );
  XOR \SUBBYTES[4].a/U4411  ( .A(\w1[4][71] ), .B(\SUBBYTES[4].a/w1740 ), .Z(
        n10448) );
  XOR \SUBBYTES[4].a/U4410  ( .A(\SUBBYTES[4].a/w1647 ), .B(
        \SUBBYTES[4].a/w1650 ), .Z(n10449) );
  XOR \SUBBYTES[4].a/U4409  ( .A(\SUBBYTES[4].a/w1633 ), .B(
        \SUBBYTES[4].a/w1635 ), .Z(n10450) );
  XOR \SUBBYTES[4].a/U4408  ( .A(n10452), .B(n10451), .Z(\SUBBYTES[4].a/w1657 ) );
  XOR \SUBBYTES[4].a/U4407  ( .A(n10885), .B(n10453), .Z(n10451) );
  XOR \SUBBYTES[4].a/U4406  ( .A(\w1[4][69] ), .B(n10886), .Z(n10452) );
  XOR \SUBBYTES[4].a/U4405  ( .A(\SUBBYTES[4].a/w1647 ), .B(
        \SUBBYTES[4].a/w1648 ), .Z(n10453) );
  XOR \SUBBYTES[4].a/U4404  ( .A(n10455), .B(n10454), .Z(\SUBBYTES[4].a/w1673 ) );
  XOR \SUBBYTES[4].a/U4403  ( .A(\w1[4][65] ), .B(n10456), .Z(n10454) );
  XOR \SUBBYTES[4].a/U4402  ( .A(\SUBBYTES[4].a/w1648 ), .B(
        \SUBBYTES[4].a/w1650 ), .Z(n10455) );
  XOR \SUBBYTES[4].a/U4401  ( .A(\SUBBYTES[4].a/w1632 ), .B(
        \SUBBYTES[4].a/w1633 ), .Z(n10456) );
  XOR \SUBBYTES[4].a/U4400  ( .A(\w1[4][73] ), .B(n10457), .Z(n10887) );
  XOR \SUBBYTES[4].a/U4399  ( .A(\w1[4][75] ), .B(\w1[4][74] ), .Z(n10457) );
  XOR \SUBBYTES[4].a/U4398  ( .A(\w1[4][78] ), .B(n10887), .Z(
        \SUBBYTES[4].a/w1515 ) );
  XOR \SUBBYTES[4].a/U4397  ( .A(\w1[4][72] ), .B(\SUBBYTES[4].a/w1515 ), .Z(
        \SUBBYTES[4].a/w1402 ) );
  XOR \SUBBYTES[4].a/U4396  ( .A(\w1[4][72] ), .B(n10458), .Z(
        \SUBBYTES[4].a/w1403 ) );
  XOR \SUBBYTES[4].a/U4395  ( .A(\w1[4][78] ), .B(\w1[4][77] ), .Z(n10458) );
  XOR \SUBBYTES[4].a/U4394  ( .A(\w1[4][77] ), .B(n10887), .Z(
        \SUBBYTES[4].a/w1533 ) );
  XOR \SUBBYTES[4].a/U4393  ( .A(n10460), .B(n10459), .Z(\SUBBYTES[4].a/w1526 ) );
  XOR \SUBBYTES[4].a/U4392  ( .A(\w1[4][75] ), .B(\w1[4][73] ), .Z(n10459) );
  XOR \SUBBYTES[4].a/U4391  ( .A(\w1[4][79] ), .B(\w1[4][76] ), .Z(n10460) );
  XOR \SUBBYTES[4].a/U4390  ( .A(\w1[4][72] ), .B(\SUBBYTES[4].a/w1526 ), .Z(
        \SUBBYTES[4].a/w1405 ) );
  XOR \SUBBYTES[4].a/U4389  ( .A(n10462), .B(n10461), .Z(\SUBBYTES[4].a/w1513 ) );
  XOR \SUBBYTES[4].a/U4388  ( .A(\SUBBYTES[4].a/w1474 ), .B(n1011), .Z(n10461)
         );
  XOR \SUBBYTES[4].a/U4387  ( .A(\SUBBYTES[4].a/w1467 ), .B(
        \SUBBYTES[4].a/w1470 ), .Z(n10462) );
  XOR \SUBBYTES[4].a/U4386  ( .A(n10464), .B(n10463), .Z(\SUBBYTES[4].a/w1514 ) );
  XOR \SUBBYTES[4].a/U4385  ( .A(\SUBBYTES[4].a/w1474 ), .B(n9685), .Z(n10463)
         );
  XOR \SUBBYTES[4].a/U4384  ( .A(\SUBBYTES[4].a/w1467 ), .B(n9684), .Z(n10464)
         );
  XOR \SUBBYTES[4].a/U4383  ( .A(\SUBBYTES[4].a/w1526 ), .B(n10465), .Z(
        \SUBBYTES[4].a/w1516 ) );
  XOR \SUBBYTES[4].a/U4382  ( .A(\w1[4][78] ), .B(\w1[4][77] ), .Z(n10465) );
  XOR \SUBBYTES[4].a/U4381  ( .A(n10467), .B(n10466), .Z(\SUBBYTES[4].a/w1517 ) );
  XOR \SUBBYTES[4].a/U4380  ( .A(n9685), .B(n1011), .Z(n10466) );
  XOR \SUBBYTES[4].a/U4379  ( .A(n9684), .B(\SUBBYTES[4].a/w1470 ), .Z(n10467)
         );
  XOR \SUBBYTES[4].a/U4378  ( .A(\w1[4][79] ), .B(\w1[4][74] ), .Z(n10893) );
  XOR \SUBBYTES[4].a/U4377  ( .A(n10893), .B(n10468), .Z(\SUBBYTES[4].a/w1518 ) );
  XOR \SUBBYTES[4].a/U4376  ( .A(\w1[4][77] ), .B(\w1[4][76] ), .Z(n10468) );
  XOR \SUBBYTES[4].a/U4375  ( .A(\w1[4][79] ), .B(\SUBBYTES[4].a/w1403 ), .Z(
        \SUBBYTES[4].a/w1406 ) );
  XOR \SUBBYTES[4].a/U4374  ( .A(\w1[4][73] ), .B(\SUBBYTES[4].a/w1403 ), .Z(
        \SUBBYTES[4].a/w1407 ) );
  XOR \SUBBYTES[4].a/U4373  ( .A(\w1[4][76] ), .B(\SUBBYTES[4].a/w1403 ), .Z(
        \SUBBYTES[4].a/w1408 ) );
  XOR \SUBBYTES[4].a/U4372  ( .A(\SUBBYTES[4].a/w1407 ), .B(n10893), .Z(
        \SUBBYTES[4].a/w1409 ) );
  XOR \SUBBYTES[4].a/U4371  ( .A(n10893), .B(n10469), .Z(\SUBBYTES[4].a/w1494 ) );
  XOR \SUBBYTES[4].a/U4370  ( .A(\w1[4][76] ), .B(\w1[4][73] ), .Z(n10469) );
  XOR \SUBBYTES[4].a/U4369  ( .A(n10471), .B(n10470), .Z(n10890) );
  XOR \SUBBYTES[4].a/U4368  ( .A(\w1[4][76] ), .B(n10472), .Z(n10470) );
  XOR \SUBBYTES[4].a/U4367  ( .A(\SUBBYTES[4].a/w1459 ), .B(\w1[4][78] ), .Z(
        n10471) );
  XOR \SUBBYTES[4].a/U4366  ( .A(\SUBBYTES[4].a/w1433 ), .B(
        \SUBBYTES[4].a/w1440 ), .Z(n10472) );
  XOR \SUBBYTES[4].a/U4365  ( .A(n10474), .B(n10473), .Z(n10888) );
  XOR \SUBBYTES[4].a/U4364  ( .A(\w1[4][73] ), .B(n10475), .Z(n10473) );
  XOR \SUBBYTES[4].a/U4363  ( .A(\SUBBYTES[4].a/w1458 ), .B(\w1[4][77] ), .Z(
        n10474) );
  XOR \SUBBYTES[4].a/U4362  ( .A(\SUBBYTES[4].a/w1434 ), .B(
        \SUBBYTES[4].a/w1441 ), .Z(n10475) );
  XOR \SUBBYTES[4].a/U4361  ( .A(n10890), .B(n10888), .Z(\SUBBYTES[4].a/w1464 ) );
  XOR \SUBBYTES[4].a/U4360  ( .A(\w1[4][77] ), .B(n10476), .Z(n10891) );
  XOR \SUBBYTES[4].a/U4359  ( .A(\SUBBYTES[4].a/w1426 ), .B(
        \SUBBYTES[4].a/w1436 ), .Z(n10476) );
  XOR \SUBBYTES[4].a/U4358  ( .A(n10478), .B(n10477), .Z(\SUBBYTES[4].a/w1451 ) );
  XOR \SUBBYTES[4].a/U4357  ( .A(n10891), .B(n10479), .Z(n10477) );
  XOR \SUBBYTES[4].a/U4356  ( .A(\w1[4][76] ), .B(\SUBBYTES[4].a/w1515 ), .Z(
        n10478) );
  XOR \SUBBYTES[4].a/U4355  ( .A(\SUBBYTES[4].a/w1428 ), .B(
        \SUBBYTES[4].a/w1433 ), .Z(n10479) );
  XOR \SUBBYTES[4].a/U4354  ( .A(n10481), .B(n10480), .Z(n10889) );
  XOR \SUBBYTES[4].a/U4353  ( .A(\SUBBYTES[4].a/w1461 ), .B(\w1[4][79] ), .Z(
        n10480) );
  XOR \SUBBYTES[4].a/U4352  ( .A(\SUBBYTES[4].a/w1436 ), .B(
        \SUBBYTES[4].a/w1443 ), .Z(n10481) );
  XOR \SUBBYTES[4].a/U4351  ( .A(n10888), .B(n10889), .Z(\SUBBYTES[4].a/w1463 ) );
  XOR \SUBBYTES[4].a/U4350  ( .A(\w1[4][75] ), .B(n10482), .Z(n10892) );
  XOR \SUBBYTES[4].a/U4349  ( .A(\SUBBYTES[4].a/w1425 ), .B(
        \SUBBYTES[4].a/w1428 ), .Z(n10482) );
  XOR \SUBBYTES[4].a/U4348  ( .A(n10484), .B(n10483), .Z(\SUBBYTES[4].a/w1452 ) );
  XOR \SUBBYTES[4].a/U4347  ( .A(n10892), .B(n10485), .Z(n10483) );
  XOR \SUBBYTES[4].a/U4346  ( .A(\w1[4][78] ), .B(\SUBBYTES[4].a/w1494 ), .Z(
        n10484) );
  XOR \SUBBYTES[4].a/U4345  ( .A(\SUBBYTES[4].a/w1433 ), .B(
        \SUBBYTES[4].a/w1434 ), .Z(n10485) );
  XOR \SUBBYTES[4].a/U4344  ( .A(n10890), .B(n10889), .Z(\SUBBYTES[4].a/w1472 ) );
  XOR \SUBBYTES[4].a/U4343  ( .A(n10487), .B(n10486), .Z(\SUBBYTES[4].a/w1473 ) );
  XOR \SUBBYTES[4].a/U4342  ( .A(\w1[4][79] ), .B(n10891), .Z(n10486) );
  XOR \SUBBYTES[4].a/U4341  ( .A(\SUBBYTES[4].a/w1425 ), .B(
        \SUBBYTES[4].a/w1434 ), .Z(n10487) );
  XOR \SUBBYTES[4].a/U4340  ( .A(n10489), .B(n10488), .Z(\SUBBYTES[4].a/w1449 ) );
  XOR \SUBBYTES[4].a/U4339  ( .A(n10491), .B(n10490), .Z(n10488) );
  XOR \SUBBYTES[4].a/U4338  ( .A(\w1[4][79] ), .B(\SUBBYTES[4].a/w1533 ), .Z(
        n10489) );
  XOR \SUBBYTES[4].a/U4337  ( .A(\SUBBYTES[4].a/w1440 ), .B(
        \SUBBYTES[4].a/w1443 ), .Z(n10490) );
  XOR \SUBBYTES[4].a/U4336  ( .A(\SUBBYTES[4].a/w1426 ), .B(
        \SUBBYTES[4].a/w1428 ), .Z(n10491) );
  XOR \SUBBYTES[4].a/U4335  ( .A(n10493), .B(n10492), .Z(\SUBBYTES[4].a/w1450 ) );
  XOR \SUBBYTES[4].a/U4334  ( .A(n10892), .B(n10494), .Z(n10492) );
  XOR \SUBBYTES[4].a/U4333  ( .A(\w1[4][77] ), .B(n10893), .Z(n10493) );
  XOR \SUBBYTES[4].a/U4332  ( .A(\SUBBYTES[4].a/w1440 ), .B(
        \SUBBYTES[4].a/w1441 ), .Z(n10494) );
  XOR \SUBBYTES[4].a/U4331  ( .A(n10496), .B(n10495), .Z(\SUBBYTES[4].a/w1466 ) );
  XOR \SUBBYTES[4].a/U4330  ( .A(\w1[4][73] ), .B(n10497), .Z(n10495) );
  XOR \SUBBYTES[4].a/U4329  ( .A(\SUBBYTES[4].a/w1441 ), .B(
        \SUBBYTES[4].a/w1443 ), .Z(n10496) );
  XOR \SUBBYTES[4].a/U4328  ( .A(\SUBBYTES[4].a/w1425 ), .B(
        \SUBBYTES[4].a/w1426 ), .Z(n10497) );
  XOR \SUBBYTES[4].a/U4327  ( .A(\w1[4][81] ), .B(n10498), .Z(n10894) );
  XOR \SUBBYTES[4].a/U4326  ( .A(\w1[4][83] ), .B(\w1[4][82] ), .Z(n10498) );
  XOR \SUBBYTES[4].a/U4325  ( .A(\w1[4][86] ), .B(n10894), .Z(
        \SUBBYTES[4].a/w1308 ) );
  XOR \SUBBYTES[4].a/U4324  ( .A(\w1[4][80] ), .B(\SUBBYTES[4].a/w1308 ), .Z(
        \SUBBYTES[4].a/w1195 ) );
  XOR \SUBBYTES[4].a/U4323  ( .A(\w1[4][80] ), .B(n10499), .Z(
        \SUBBYTES[4].a/w1196 ) );
  XOR \SUBBYTES[4].a/U4322  ( .A(\w1[4][86] ), .B(\w1[4][85] ), .Z(n10499) );
  XOR \SUBBYTES[4].a/U4321  ( .A(\w1[4][85] ), .B(n10894), .Z(
        \SUBBYTES[4].a/w1326 ) );
  XOR \SUBBYTES[4].a/U4320  ( .A(n10501), .B(n10500), .Z(\SUBBYTES[4].a/w1319 ) );
  XOR \SUBBYTES[4].a/U4319  ( .A(\w1[4][83] ), .B(\w1[4][81] ), .Z(n10500) );
  XOR \SUBBYTES[4].a/U4318  ( .A(\w1[4][87] ), .B(\w1[4][84] ), .Z(n10501) );
  XOR \SUBBYTES[4].a/U4317  ( .A(\w1[4][80] ), .B(\SUBBYTES[4].a/w1319 ), .Z(
        \SUBBYTES[4].a/w1198 ) );
  XOR \SUBBYTES[4].a/U4316  ( .A(n10503), .B(n10502), .Z(\SUBBYTES[4].a/w1306 ) );
  XOR \SUBBYTES[4].a/U4315  ( .A(\SUBBYTES[4].a/w1267 ), .B(n1010), .Z(n10502)
         );
  XOR \SUBBYTES[4].a/U4314  ( .A(\SUBBYTES[4].a/w1260 ), .B(
        \SUBBYTES[4].a/w1263 ), .Z(n10503) );
  XOR \SUBBYTES[4].a/U4313  ( .A(n10505), .B(n10504), .Z(\SUBBYTES[4].a/w1307 ) );
  XOR \SUBBYTES[4].a/U4312  ( .A(\SUBBYTES[4].a/w1267 ), .B(n9683), .Z(n10504)
         );
  XOR \SUBBYTES[4].a/U4311  ( .A(\SUBBYTES[4].a/w1260 ), .B(n9682), .Z(n10505)
         );
  XOR \SUBBYTES[4].a/U4310  ( .A(\SUBBYTES[4].a/w1319 ), .B(n10506), .Z(
        \SUBBYTES[4].a/w1309 ) );
  XOR \SUBBYTES[4].a/U4309  ( .A(\w1[4][86] ), .B(\w1[4][85] ), .Z(n10506) );
  XOR \SUBBYTES[4].a/U4308  ( .A(n10508), .B(n10507), .Z(\SUBBYTES[4].a/w1310 ) );
  XOR \SUBBYTES[4].a/U4307  ( .A(n9683), .B(n1010), .Z(n10507) );
  XOR \SUBBYTES[4].a/U4306  ( .A(n9682), .B(\SUBBYTES[4].a/w1263 ), .Z(n10508)
         );
  XOR \SUBBYTES[4].a/U4305  ( .A(\w1[4][87] ), .B(\w1[4][82] ), .Z(n10900) );
  XOR \SUBBYTES[4].a/U4304  ( .A(n10900), .B(n10509), .Z(\SUBBYTES[4].a/w1311 ) );
  XOR \SUBBYTES[4].a/U4303  ( .A(\w1[4][85] ), .B(\w1[4][84] ), .Z(n10509) );
  XOR \SUBBYTES[4].a/U4302  ( .A(\w1[4][87] ), .B(\SUBBYTES[4].a/w1196 ), .Z(
        \SUBBYTES[4].a/w1199 ) );
  XOR \SUBBYTES[4].a/U4301  ( .A(\w1[4][81] ), .B(\SUBBYTES[4].a/w1196 ), .Z(
        \SUBBYTES[4].a/w1200 ) );
  XOR \SUBBYTES[4].a/U4300  ( .A(\w1[4][84] ), .B(\SUBBYTES[4].a/w1196 ), .Z(
        \SUBBYTES[4].a/w1201 ) );
  XOR \SUBBYTES[4].a/U4299  ( .A(\SUBBYTES[4].a/w1200 ), .B(n10900), .Z(
        \SUBBYTES[4].a/w1202 ) );
  XOR \SUBBYTES[4].a/U4298  ( .A(n10900), .B(n10510), .Z(\SUBBYTES[4].a/w1287 ) );
  XOR \SUBBYTES[4].a/U4297  ( .A(\w1[4][84] ), .B(\w1[4][81] ), .Z(n10510) );
  XOR \SUBBYTES[4].a/U4296  ( .A(n10512), .B(n10511), .Z(n10897) );
  XOR \SUBBYTES[4].a/U4295  ( .A(\w1[4][84] ), .B(n10513), .Z(n10511) );
  XOR \SUBBYTES[4].a/U4294  ( .A(\SUBBYTES[4].a/w1252 ), .B(\w1[4][86] ), .Z(
        n10512) );
  XOR \SUBBYTES[4].a/U4293  ( .A(\SUBBYTES[4].a/w1226 ), .B(
        \SUBBYTES[4].a/w1233 ), .Z(n10513) );
  XOR \SUBBYTES[4].a/U4292  ( .A(n10515), .B(n10514), .Z(n10895) );
  XOR \SUBBYTES[4].a/U4291  ( .A(\w1[4][81] ), .B(n10516), .Z(n10514) );
  XOR \SUBBYTES[4].a/U4290  ( .A(\SUBBYTES[4].a/w1251 ), .B(\w1[4][85] ), .Z(
        n10515) );
  XOR \SUBBYTES[4].a/U4289  ( .A(\SUBBYTES[4].a/w1227 ), .B(
        \SUBBYTES[4].a/w1234 ), .Z(n10516) );
  XOR \SUBBYTES[4].a/U4288  ( .A(n10897), .B(n10895), .Z(\SUBBYTES[4].a/w1257 ) );
  XOR \SUBBYTES[4].a/U4287  ( .A(\w1[4][85] ), .B(n10517), .Z(n10898) );
  XOR \SUBBYTES[4].a/U4286  ( .A(\SUBBYTES[4].a/w1219 ), .B(
        \SUBBYTES[4].a/w1229 ), .Z(n10517) );
  XOR \SUBBYTES[4].a/U4285  ( .A(n10519), .B(n10518), .Z(\SUBBYTES[4].a/w1244 ) );
  XOR \SUBBYTES[4].a/U4284  ( .A(n10898), .B(n10520), .Z(n10518) );
  XOR \SUBBYTES[4].a/U4283  ( .A(\w1[4][84] ), .B(\SUBBYTES[4].a/w1308 ), .Z(
        n10519) );
  XOR \SUBBYTES[4].a/U4282  ( .A(\SUBBYTES[4].a/w1221 ), .B(
        \SUBBYTES[4].a/w1226 ), .Z(n10520) );
  XOR \SUBBYTES[4].a/U4281  ( .A(n10522), .B(n10521), .Z(n10896) );
  XOR \SUBBYTES[4].a/U4280  ( .A(\SUBBYTES[4].a/w1254 ), .B(\w1[4][87] ), .Z(
        n10521) );
  XOR \SUBBYTES[4].a/U4279  ( .A(\SUBBYTES[4].a/w1229 ), .B(
        \SUBBYTES[4].a/w1236 ), .Z(n10522) );
  XOR \SUBBYTES[4].a/U4278  ( .A(n10895), .B(n10896), .Z(\SUBBYTES[4].a/w1256 ) );
  XOR \SUBBYTES[4].a/U4277  ( .A(\w1[4][83] ), .B(n10523), .Z(n10899) );
  XOR \SUBBYTES[4].a/U4276  ( .A(\SUBBYTES[4].a/w1218 ), .B(
        \SUBBYTES[4].a/w1221 ), .Z(n10523) );
  XOR \SUBBYTES[4].a/U4275  ( .A(n10525), .B(n10524), .Z(\SUBBYTES[4].a/w1245 ) );
  XOR \SUBBYTES[4].a/U4274  ( .A(n10899), .B(n10526), .Z(n10524) );
  XOR \SUBBYTES[4].a/U4273  ( .A(\w1[4][86] ), .B(\SUBBYTES[4].a/w1287 ), .Z(
        n10525) );
  XOR \SUBBYTES[4].a/U4272  ( .A(\SUBBYTES[4].a/w1226 ), .B(
        \SUBBYTES[4].a/w1227 ), .Z(n10526) );
  XOR \SUBBYTES[4].a/U4271  ( .A(n10897), .B(n10896), .Z(\SUBBYTES[4].a/w1265 ) );
  XOR \SUBBYTES[4].a/U4270  ( .A(n10528), .B(n10527), .Z(\SUBBYTES[4].a/w1266 ) );
  XOR \SUBBYTES[4].a/U4269  ( .A(\w1[4][87] ), .B(n10898), .Z(n10527) );
  XOR \SUBBYTES[4].a/U4268  ( .A(\SUBBYTES[4].a/w1218 ), .B(
        \SUBBYTES[4].a/w1227 ), .Z(n10528) );
  XOR \SUBBYTES[4].a/U4267  ( .A(n10530), .B(n10529), .Z(\SUBBYTES[4].a/w1242 ) );
  XOR \SUBBYTES[4].a/U4266  ( .A(n10532), .B(n10531), .Z(n10529) );
  XOR \SUBBYTES[4].a/U4265  ( .A(\w1[4][87] ), .B(\SUBBYTES[4].a/w1326 ), .Z(
        n10530) );
  XOR \SUBBYTES[4].a/U4264  ( .A(\SUBBYTES[4].a/w1233 ), .B(
        \SUBBYTES[4].a/w1236 ), .Z(n10531) );
  XOR \SUBBYTES[4].a/U4263  ( .A(\SUBBYTES[4].a/w1219 ), .B(
        \SUBBYTES[4].a/w1221 ), .Z(n10532) );
  XOR \SUBBYTES[4].a/U4262  ( .A(n10534), .B(n10533), .Z(\SUBBYTES[4].a/w1243 ) );
  XOR \SUBBYTES[4].a/U4261  ( .A(n10899), .B(n10535), .Z(n10533) );
  XOR \SUBBYTES[4].a/U4260  ( .A(\w1[4][85] ), .B(n10900), .Z(n10534) );
  XOR \SUBBYTES[4].a/U4259  ( .A(\SUBBYTES[4].a/w1233 ), .B(
        \SUBBYTES[4].a/w1234 ), .Z(n10535) );
  XOR \SUBBYTES[4].a/U4258  ( .A(n10537), .B(n10536), .Z(\SUBBYTES[4].a/w1259 ) );
  XOR \SUBBYTES[4].a/U4257  ( .A(\w1[4][81] ), .B(n10538), .Z(n10536) );
  XOR \SUBBYTES[4].a/U4256  ( .A(\SUBBYTES[4].a/w1234 ), .B(
        \SUBBYTES[4].a/w1236 ), .Z(n10537) );
  XOR \SUBBYTES[4].a/U4255  ( .A(\SUBBYTES[4].a/w1218 ), .B(
        \SUBBYTES[4].a/w1219 ), .Z(n10538) );
  XOR \SUBBYTES[4].a/U4254  ( .A(\w1[4][89] ), .B(n10539), .Z(n10901) );
  XOR \SUBBYTES[4].a/U4253  ( .A(\w1[4][91] ), .B(\w1[4][90] ), .Z(n10539) );
  XOR \SUBBYTES[4].a/U4252  ( .A(\w1[4][94] ), .B(n10901), .Z(
        \SUBBYTES[4].a/w1101 ) );
  XOR \SUBBYTES[4].a/U4251  ( .A(\w1[4][88] ), .B(\SUBBYTES[4].a/w1101 ), .Z(
        \SUBBYTES[4].a/w988 ) );
  XOR \SUBBYTES[4].a/U4250  ( .A(\w1[4][88] ), .B(n10540), .Z(
        \SUBBYTES[4].a/w989 ) );
  XOR \SUBBYTES[4].a/U4249  ( .A(\w1[4][94] ), .B(\w1[4][93] ), .Z(n10540) );
  XOR \SUBBYTES[4].a/U4248  ( .A(\w1[4][93] ), .B(n10901), .Z(
        \SUBBYTES[4].a/w1119 ) );
  XOR \SUBBYTES[4].a/U4247  ( .A(n10542), .B(n10541), .Z(\SUBBYTES[4].a/w1112 ) );
  XOR \SUBBYTES[4].a/U4246  ( .A(\w1[4][91] ), .B(\w1[4][89] ), .Z(n10541) );
  XOR \SUBBYTES[4].a/U4245  ( .A(\w1[4][95] ), .B(\w1[4][92] ), .Z(n10542) );
  XOR \SUBBYTES[4].a/U4244  ( .A(\w1[4][88] ), .B(\SUBBYTES[4].a/w1112 ), .Z(
        \SUBBYTES[4].a/w991 ) );
  XOR \SUBBYTES[4].a/U4243  ( .A(n10544), .B(n10543), .Z(\SUBBYTES[4].a/w1099 ) );
  XOR \SUBBYTES[4].a/U4242  ( .A(\SUBBYTES[4].a/w1060 ), .B(n1009), .Z(n10543)
         );
  XOR \SUBBYTES[4].a/U4241  ( .A(\SUBBYTES[4].a/w1053 ), .B(
        \SUBBYTES[4].a/w1056 ), .Z(n10544) );
  XOR \SUBBYTES[4].a/U4240  ( .A(n10546), .B(n10545), .Z(\SUBBYTES[4].a/w1100 ) );
  XOR \SUBBYTES[4].a/U4239  ( .A(\SUBBYTES[4].a/w1060 ), .B(n9681), .Z(n10545)
         );
  XOR \SUBBYTES[4].a/U4238  ( .A(\SUBBYTES[4].a/w1053 ), .B(n9680), .Z(n10546)
         );
  XOR \SUBBYTES[4].a/U4237  ( .A(\SUBBYTES[4].a/w1112 ), .B(n10547), .Z(
        \SUBBYTES[4].a/w1102 ) );
  XOR \SUBBYTES[4].a/U4236  ( .A(\w1[4][94] ), .B(\w1[4][93] ), .Z(n10547) );
  XOR \SUBBYTES[4].a/U4235  ( .A(n10549), .B(n10548), .Z(\SUBBYTES[4].a/w1103 ) );
  XOR \SUBBYTES[4].a/U4234  ( .A(n9681), .B(n1009), .Z(n10548) );
  XOR \SUBBYTES[4].a/U4233  ( .A(n9680), .B(\SUBBYTES[4].a/w1056 ), .Z(n10549)
         );
  XOR \SUBBYTES[4].a/U4232  ( .A(\w1[4][95] ), .B(\w1[4][90] ), .Z(n10907) );
  XOR \SUBBYTES[4].a/U4231  ( .A(n10907), .B(n10550), .Z(\SUBBYTES[4].a/w1104 ) );
  XOR \SUBBYTES[4].a/U4230  ( .A(\w1[4][93] ), .B(\w1[4][92] ), .Z(n10550) );
  XOR \SUBBYTES[4].a/U4229  ( .A(\w1[4][95] ), .B(\SUBBYTES[4].a/w989 ), .Z(
        \SUBBYTES[4].a/w992 ) );
  XOR \SUBBYTES[4].a/U4228  ( .A(\w1[4][89] ), .B(\SUBBYTES[4].a/w989 ), .Z(
        \SUBBYTES[4].a/w993 ) );
  XOR \SUBBYTES[4].a/U4227  ( .A(\w1[4][92] ), .B(\SUBBYTES[4].a/w989 ), .Z(
        \SUBBYTES[4].a/w994 ) );
  XOR \SUBBYTES[4].a/U4226  ( .A(\SUBBYTES[4].a/w993 ), .B(n10907), .Z(
        \SUBBYTES[4].a/w995 ) );
  XOR \SUBBYTES[4].a/U4225  ( .A(n10907), .B(n10551), .Z(\SUBBYTES[4].a/w1080 ) );
  XOR \SUBBYTES[4].a/U4224  ( .A(\w1[4][92] ), .B(\w1[4][89] ), .Z(n10551) );
  XOR \SUBBYTES[4].a/U4223  ( .A(n10553), .B(n10552), .Z(n10904) );
  XOR \SUBBYTES[4].a/U4222  ( .A(\w1[4][92] ), .B(n10554), .Z(n10552) );
  XOR \SUBBYTES[4].a/U4221  ( .A(\SUBBYTES[4].a/w1045 ), .B(\w1[4][94] ), .Z(
        n10553) );
  XOR \SUBBYTES[4].a/U4220  ( .A(\SUBBYTES[4].a/w1019 ), .B(
        \SUBBYTES[4].a/w1026 ), .Z(n10554) );
  XOR \SUBBYTES[4].a/U4219  ( .A(n10556), .B(n10555), .Z(n10902) );
  XOR \SUBBYTES[4].a/U4218  ( .A(\w1[4][89] ), .B(n10557), .Z(n10555) );
  XOR \SUBBYTES[4].a/U4217  ( .A(\SUBBYTES[4].a/w1044 ), .B(\w1[4][93] ), .Z(
        n10556) );
  XOR \SUBBYTES[4].a/U4216  ( .A(\SUBBYTES[4].a/w1020 ), .B(
        \SUBBYTES[4].a/w1027 ), .Z(n10557) );
  XOR \SUBBYTES[4].a/U4215  ( .A(n10904), .B(n10902), .Z(\SUBBYTES[4].a/w1050 ) );
  XOR \SUBBYTES[4].a/U4214  ( .A(\w1[4][93] ), .B(n10558), .Z(n10905) );
  XOR \SUBBYTES[4].a/U4213  ( .A(\SUBBYTES[4].a/w1012 ), .B(
        \SUBBYTES[4].a/w1022 ), .Z(n10558) );
  XOR \SUBBYTES[4].a/U4212  ( .A(n10560), .B(n10559), .Z(\SUBBYTES[4].a/w1037 ) );
  XOR \SUBBYTES[4].a/U4211  ( .A(n10905), .B(n10561), .Z(n10559) );
  XOR \SUBBYTES[4].a/U4210  ( .A(\w1[4][92] ), .B(\SUBBYTES[4].a/w1101 ), .Z(
        n10560) );
  XOR \SUBBYTES[4].a/U4209  ( .A(\SUBBYTES[4].a/w1014 ), .B(
        \SUBBYTES[4].a/w1019 ), .Z(n10561) );
  XOR \SUBBYTES[4].a/U4208  ( .A(n10563), .B(n10562), .Z(n10903) );
  XOR \SUBBYTES[4].a/U4207  ( .A(\SUBBYTES[4].a/w1047 ), .B(\w1[4][95] ), .Z(
        n10562) );
  XOR \SUBBYTES[4].a/U4206  ( .A(\SUBBYTES[4].a/w1022 ), .B(
        \SUBBYTES[4].a/w1029 ), .Z(n10563) );
  XOR \SUBBYTES[4].a/U4205  ( .A(n10902), .B(n10903), .Z(\SUBBYTES[4].a/w1049 ) );
  XOR \SUBBYTES[4].a/U4204  ( .A(\w1[4][91] ), .B(n10564), .Z(n10906) );
  XOR \SUBBYTES[4].a/U4203  ( .A(\SUBBYTES[4].a/w1011 ), .B(
        \SUBBYTES[4].a/w1014 ), .Z(n10564) );
  XOR \SUBBYTES[4].a/U4202  ( .A(n10566), .B(n10565), .Z(\SUBBYTES[4].a/w1038 ) );
  XOR \SUBBYTES[4].a/U4201  ( .A(n10906), .B(n10567), .Z(n10565) );
  XOR \SUBBYTES[4].a/U4200  ( .A(\w1[4][94] ), .B(\SUBBYTES[4].a/w1080 ), .Z(
        n10566) );
  XOR \SUBBYTES[4].a/U4199  ( .A(\SUBBYTES[4].a/w1019 ), .B(
        \SUBBYTES[4].a/w1020 ), .Z(n10567) );
  XOR \SUBBYTES[4].a/U4198  ( .A(n10904), .B(n10903), .Z(\SUBBYTES[4].a/w1058 ) );
  XOR \SUBBYTES[4].a/U4197  ( .A(n10569), .B(n10568), .Z(\SUBBYTES[4].a/w1059 ) );
  XOR \SUBBYTES[4].a/U4196  ( .A(\w1[4][95] ), .B(n10905), .Z(n10568) );
  XOR \SUBBYTES[4].a/U4195  ( .A(\SUBBYTES[4].a/w1011 ), .B(
        \SUBBYTES[4].a/w1020 ), .Z(n10569) );
  XOR \SUBBYTES[4].a/U4194  ( .A(n10571), .B(n10570), .Z(\SUBBYTES[4].a/w1035 ) );
  XOR \SUBBYTES[4].a/U4193  ( .A(n10573), .B(n10572), .Z(n10570) );
  XOR \SUBBYTES[4].a/U4192  ( .A(\w1[4][95] ), .B(\SUBBYTES[4].a/w1119 ), .Z(
        n10571) );
  XOR \SUBBYTES[4].a/U4191  ( .A(\SUBBYTES[4].a/w1026 ), .B(
        \SUBBYTES[4].a/w1029 ), .Z(n10572) );
  XOR \SUBBYTES[4].a/U4190  ( .A(\SUBBYTES[4].a/w1012 ), .B(
        \SUBBYTES[4].a/w1014 ), .Z(n10573) );
  XOR \SUBBYTES[4].a/U4189  ( .A(n10575), .B(n10574), .Z(\SUBBYTES[4].a/w1036 ) );
  XOR \SUBBYTES[4].a/U4188  ( .A(n10906), .B(n10576), .Z(n10574) );
  XOR \SUBBYTES[4].a/U4187  ( .A(\w1[4][93] ), .B(n10907), .Z(n10575) );
  XOR \SUBBYTES[4].a/U4186  ( .A(\SUBBYTES[4].a/w1026 ), .B(
        \SUBBYTES[4].a/w1027 ), .Z(n10576) );
  XOR \SUBBYTES[4].a/U4185  ( .A(n10578), .B(n10577), .Z(\SUBBYTES[4].a/w1052 ) );
  XOR \SUBBYTES[4].a/U4184  ( .A(\w1[4][89] ), .B(n10579), .Z(n10577) );
  XOR \SUBBYTES[4].a/U4183  ( .A(\SUBBYTES[4].a/w1027 ), .B(
        \SUBBYTES[4].a/w1029 ), .Z(n10578) );
  XOR \SUBBYTES[4].a/U4182  ( .A(\SUBBYTES[4].a/w1011 ), .B(
        \SUBBYTES[4].a/w1012 ), .Z(n10579) );
  XOR \SUBBYTES[4].a/U4181  ( .A(\w1[4][97] ), .B(n10580), .Z(n10908) );
  XOR \SUBBYTES[4].a/U4180  ( .A(\w1[4][99] ), .B(\w1[4][98] ), .Z(n10580) );
  XOR \SUBBYTES[4].a/U4179  ( .A(\w1[4][102] ), .B(n10908), .Z(
        \SUBBYTES[4].a/w894 ) );
  XOR \SUBBYTES[4].a/U4178  ( .A(\w1[4][96] ), .B(\SUBBYTES[4].a/w894 ), .Z(
        \SUBBYTES[4].a/w781 ) );
  XOR \SUBBYTES[4].a/U4177  ( .A(\w1[4][96] ), .B(n10581), .Z(
        \SUBBYTES[4].a/w782 ) );
  XOR \SUBBYTES[4].a/U4176  ( .A(\w1[4][102] ), .B(\w1[4][101] ), .Z(n10581)
         );
  XOR \SUBBYTES[4].a/U4175  ( .A(\w1[4][101] ), .B(n10908), .Z(
        \SUBBYTES[4].a/w912 ) );
  XOR \SUBBYTES[4].a/U4174  ( .A(n10583), .B(n10582), .Z(\SUBBYTES[4].a/w905 )
         );
  XOR \SUBBYTES[4].a/U4173  ( .A(\w1[4][99] ), .B(\w1[4][97] ), .Z(n10582) );
  XOR \SUBBYTES[4].a/U4172  ( .A(\w1[4][103] ), .B(\w1[4][100] ), .Z(n10583)
         );
  XOR \SUBBYTES[4].a/U4171  ( .A(\w1[4][96] ), .B(\SUBBYTES[4].a/w905 ), .Z(
        \SUBBYTES[4].a/w784 ) );
  XOR \SUBBYTES[4].a/U4170  ( .A(n10585), .B(n10584), .Z(\SUBBYTES[4].a/w892 )
         );
  XOR \SUBBYTES[4].a/U4169  ( .A(\SUBBYTES[4].a/w853 ), .B(n1008), .Z(n10584)
         );
  XOR \SUBBYTES[4].a/U4168  ( .A(\SUBBYTES[4].a/w846 ), .B(
        \SUBBYTES[4].a/w849 ), .Z(n10585) );
  XOR \SUBBYTES[4].a/U4167  ( .A(n10587), .B(n10586), .Z(\SUBBYTES[4].a/w893 )
         );
  XOR \SUBBYTES[4].a/U4166  ( .A(\SUBBYTES[4].a/w853 ), .B(n9679), .Z(n10586)
         );
  XOR \SUBBYTES[4].a/U4165  ( .A(\SUBBYTES[4].a/w846 ), .B(n9678), .Z(n10587)
         );
  XOR \SUBBYTES[4].a/U4164  ( .A(\SUBBYTES[4].a/w905 ), .B(n10588), .Z(
        \SUBBYTES[4].a/w895 ) );
  XOR \SUBBYTES[4].a/U4163  ( .A(\w1[4][102] ), .B(\w1[4][101] ), .Z(n10588)
         );
  XOR \SUBBYTES[4].a/U4162  ( .A(n10590), .B(n10589), .Z(\SUBBYTES[4].a/w896 )
         );
  XOR \SUBBYTES[4].a/U4161  ( .A(n9679), .B(n1008), .Z(n10589) );
  XOR \SUBBYTES[4].a/U4160  ( .A(n9678), .B(\SUBBYTES[4].a/w849 ), .Z(n10590)
         );
  XOR \SUBBYTES[4].a/U4159  ( .A(\w1[4][103] ), .B(\w1[4][98] ), .Z(n10914) );
  XOR \SUBBYTES[4].a/U4158  ( .A(n10914), .B(n10591), .Z(\SUBBYTES[4].a/w897 )
         );
  XOR \SUBBYTES[4].a/U4157  ( .A(\w1[4][101] ), .B(\w1[4][100] ), .Z(n10591)
         );
  XOR \SUBBYTES[4].a/U4156  ( .A(\w1[4][103] ), .B(\SUBBYTES[4].a/w782 ), .Z(
        \SUBBYTES[4].a/w785 ) );
  XOR \SUBBYTES[4].a/U4155  ( .A(\w1[4][97] ), .B(\SUBBYTES[4].a/w782 ), .Z(
        \SUBBYTES[4].a/w786 ) );
  XOR \SUBBYTES[4].a/U4154  ( .A(\w1[4][100] ), .B(\SUBBYTES[4].a/w782 ), .Z(
        \SUBBYTES[4].a/w787 ) );
  XOR \SUBBYTES[4].a/U4153  ( .A(\SUBBYTES[4].a/w786 ), .B(n10914), .Z(
        \SUBBYTES[4].a/w788 ) );
  XOR \SUBBYTES[4].a/U4152  ( .A(n10914), .B(n10592), .Z(\SUBBYTES[4].a/w873 )
         );
  XOR \SUBBYTES[4].a/U4151  ( .A(\w1[4][100] ), .B(\w1[4][97] ), .Z(n10592) );
  XOR \SUBBYTES[4].a/U4150  ( .A(n10594), .B(n10593), .Z(n10911) );
  XOR \SUBBYTES[4].a/U4149  ( .A(\w1[4][100] ), .B(n10595), .Z(n10593) );
  XOR \SUBBYTES[4].a/U4148  ( .A(\SUBBYTES[4].a/w838 ), .B(\w1[4][102] ), .Z(
        n10594) );
  XOR \SUBBYTES[4].a/U4147  ( .A(\SUBBYTES[4].a/w812 ), .B(
        \SUBBYTES[4].a/w819 ), .Z(n10595) );
  XOR \SUBBYTES[4].a/U4146  ( .A(n10597), .B(n10596), .Z(n10909) );
  XOR \SUBBYTES[4].a/U4145  ( .A(\w1[4][97] ), .B(n10598), .Z(n10596) );
  XOR \SUBBYTES[4].a/U4144  ( .A(\SUBBYTES[4].a/w837 ), .B(\w1[4][101] ), .Z(
        n10597) );
  XOR \SUBBYTES[4].a/U4143  ( .A(\SUBBYTES[4].a/w813 ), .B(
        \SUBBYTES[4].a/w820 ), .Z(n10598) );
  XOR \SUBBYTES[4].a/U4142  ( .A(n10911), .B(n10909), .Z(\SUBBYTES[4].a/w843 )
         );
  XOR \SUBBYTES[4].a/U4141  ( .A(\w1[4][101] ), .B(n10599), .Z(n10912) );
  XOR \SUBBYTES[4].a/U4140  ( .A(\SUBBYTES[4].a/w805 ), .B(
        \SUBBYTES[4].a/w815 ), .Z(n10599) );
  XOR \SUBBYTES[4].a/U4139  ( .A(n10601), .B(n10600), .Z(\SUBBYTES[4].a/w830 )
         );
  XOR \SUBBYTES[4].a/U4138  ( .A(n10912), .B(n10602), .Z(n10600) );
  XOR \SUBBYTES[4].a/U4137  ( .A(\w1[4][100] ), .B(\SUBBYTES[4].a/w894 ), .Z(
        n10601) );
  XOR \SUBBYTES[4].a/U4136  ( .A(\SUBBYTES[4].a/w807 ), .B(
        \SUBBYTES[4].a/w812 ), .Z(n10602) );
  XOR \SUBBYTES[4].a/U4135  ( .A(n10604), .B(n10603), .Z(n10910) );
  XOR \SUBBYTES[4].a/U4134  ( .A(\SUBBYTES[4].a/w840 ), .B(\w1[4][103] ), .Z(
        n10603) );
  XOR \SUBBYTES[4].a/U4133  ( .A(\SUBBYTES[4].a/w815 ), .B(
        \SUBBYTES[4].a/w822 ), .Z(n10604) );
  XOR \SUBBYTES[4].a/U4132  ( .A(n10909), .B(n10910), .Z(\SUBBYTES[4].a/w842 )
         );
  XOR \SUBBYTES[4].a/U4131  ( .A(\w1[4][99] ), .B(n10605), .Z(n10913) );
  XOR \SUBBYTES[4].a/U4130  ( .A(\SUBBYTES[4].a/w804 ), .B(
        \SUBBYTES[4].a/w807 ), .Z(n10605) );
  XOR \SUBBYTES[4].a/U4129  ( .A(n10607), .B(n10606), .Z(\SUBBYTES[4].a/w831 )
         );
  XOR \SUBBYTES[4].a/U4128  ( .A(n10913), .B(n10608), .Z(n10606) );
  XOR \SUBBYTES[4].a/U4127  ( .A(\w1[4][102] ), .B(\SUBBYTES[4].a/w873 ), .Z(
        n10607) );
  XOR \SUBBYTES[4].a/U4126  ( .A(\SUBBYTES[4].a/w812 ), .B(
        \SUBBYTES[4].a/w813 ), .Z(n10608) );
  XOR \SUBBYTES[4].a/U4125  ( .A(n10911), .B(n10910), .Z(\SUBBYTES[4].a/w851 )
         );
  XOR \SUBBYTES[4].a/U4124  ( .A(n10610), .B(n10609), .Z(\SUBBYTES[4].a/w852 )
         );
  XOR \SUBBYTES[4].a/U4123  ( .A(\w1[4][103] ), .B(n10912), .Z(n10609) );
  XOR \SUBBYTES[4].a/U4122  ( .A(\SUBBYTES[4].a/w804 ), .B(
        \SUBBYTES[4].a/w813 ), .Z(n10610) );
  XOR \SUBBYTES[4].a/U4121  ( .A(n10612), .B(n10611), .Z(\SUBBYTES[4].a/w828 )
         );
  XOR \SUBBYTES[4].a/U4120  ( .A(n10614), .B(n10613), .Z(n10611) );
  XOR \SUBBYTES[4].a/U4119  ( .A(\w1[4][103] ), .B(\SUBBYTES[4].a/w912 ), .Z(
        n10612) );
  XOR \SUBBYTES[4].a/U4118  ( .A(\SUBBYTES[4].a/w819 ), .B(
        \SUBBYTES[4].a/w822 ), .Z(n10613) );
  XOR \SUBBYTES[4].a/U4117  ( .A(\SUBBYTES[4].a/w805 ), .B(
        \SUBBYTES[4].a/w807 ), .Z(n10614) );
  XOR \SUBBYTES[4].a/U4116  ( .A(n10616), .B(n10615), .Z(\SUBBYTES[4].a/w829 )
         );
  XOR \SUBBYTES[4].a/U4115  ( .A(n10913), .B(n10617), .Z(n10615) );
  XOR \SUBBYTES[4].a/U4114  ( .A(\w1[4][101] ), .B(n10914), .Z(n10616) );
  XOR \SUBBYTES[4].a/U4113  ( .A(\SUBBYTES[4].a/w819 ), .B(
        \SUBBYTES[4].a/w820 ), .Z(n10617) );
  XOR \SUBBYTES[4].a/U4112  ( .A(n10619), .B(n10618), .Z(\SUBBYTES[4].a/w845 )
         );
  XOR \SUBBYTES[4].a/U4111  ( .A(\w1[4][97] ), .B(n10620), .Z(n10618) );
  XOR \SUBBYTES[4].a/U4110  ( .A(\SUBBYTES[4].a/w820 ), .B(
        \SUBBYTES[4].a/w822 ), .Z(n10619) );
  XOR \SUBBYTES[4].a/U4109  ( .A(\SUBBYTES[4].a/w804 ), .B(
        \SUBBYTES[4].a/w805 ), .Z(n10620) );
  XOR \SUBBYTES[4].a/U4108  ( .A(\w1[4][105] ), .B(n10621), .Z(n10915) );
  XOR \SUBBYTES[4].a/U4107  ( .A(\w1[4][107] ), .B(\w1[4][106] ), .Z(n10621)
         );
  XOR \SUBBYTES[4].a/U4106  ( .A(\w1[4][110] ), .B(n10915), .Z(
        \SUBBYTES[4].a/w687 ) );
  XOR \SUBBYTES[4].a/U4105  ( .A(\w1[4][104] ), .B(\SUBBYTES[4].a/w687 ), .Z(
        \SUBBYTES[4].a/w574 ) );
  XOR \SUBBYTES[4].a/U4104  ( .A(\w1[4][104] ), .B(n10622), .Z(
        \SUBBYTES[4].a/w575 ) );
  XOR \SUBBYTES[4].a/U4103  ( .A(\w1[4][110] ), .B(\w1[4][109] ), .Z(n10622)
         );
  XOR \SUBBYTES[4].a/U4102  ( .A(\w1[4][109] ), .B(n10915), .Z(
        \SUBBYTES[4].a/w705 ) );
  XOR \SUBBYTES[4].a/U4101  ( .A(n10624), .B(n10623), .Z(\SUBBYTES[4].a/w698 )
         );
  XOR \SUBBYTES[4].a/U4100  ( .A(\w1[4][107] ), .B(\w1[4][105] ), .Z(n10623)
         );
  XOR \SUBBYTES[4].a/U4099  ( .A(\w1[4][111] ), .B(\w1[4][108] ), .Z(n10624)
         );
  XOR \SUBBYTES[4].a/U4098  ( .A(\w1[4][104] ), .B(\SUBBYTES[4].a/w698 ), .Z(
        \SUBBYTES[4].a/w577 ) );
  XOR \SUBBYTES[4].a/U4097  ( .A(n10626), .B(n10625), .Z(\SUBBYTES[4].a/w685 )
         );
  XOR \SUBBYTES[4].a/U4096  ( .A(\SUBBYTES[4].a/w646 ), .B(n1007), .Z(n10625)
         );
  XOR \SUBBYTES[4].a/U4095  ( .A(\SUBBYTES[4].a/w639 ), .B(
        \SUBBYTES[4].a/w642 ), .Z(n10626) );
  XOR \SUBBYTES[4].a/U4094  ( .A(n10628), .B(n10627), .Z(\SUBBYTES[4].a/w686 )
         );
  XOR \SUBBYTES[4].a/U4093  ( .A(\SUBBYTES[4].a/w646 ), .B(n9677), .Z(n10627)
         );
  XOR \SUBBYTES[4].a/U4092  ( .A(\SUBBYTES[4].a/w639 ), .B(n9676), .Z(n10628)
         );
  XOR \SUBBYTES[4].a/U4091  ( .A(\SUBBYTES[4].a/w698 ), .B(n10629), .Z(
        \SUBBYTES[4].a/w688 ) );
  XOR \SUBBYTES[4].a/U4090  ( .A(\w1[4][110] ), .B(\w1[4][109] ), .Z(n10629)
         );
  XOR \SUBBYTES[4].a/U4089  ( .A(n10631), .B(n10630), .Z(\SUBBYTES[4].a/w689 )
         );
  XOR \SUBBYTES[4].a/U4088  ( .A(n9677), .B(n1007), .Z(n10630) );
  XOR \SUBBYTES[4].a/U4087  ( .A(n9676), .B(\SUBBYTES[4].a/w642 ), .Z(n10631)
         );
  XOR \SUBBYTES[4].a/U4086  ( .A(\w1[4][111] ), .B(\w1[4][106] ), .Z(n10921)
         );
  XOR \SUBBYTES[4].a/U4085  ( .A(n10921), .B(n10632), .Z(\SUBBYTES[4].a/w690 )
         );
  XOR \SUBBYTES[4].a/U4084  ( .A(\w1[4][109] ), .B(\w1[4][108] ), .Z(n10632)
         );
  XOR \SUBBYTES[4].a/U4083  ( .A(\w1[4][111] ), .B(\SUBBYTES[4].a/w575 ), .Z(
        \SUBBYTES[4].a/w578 ) );
  XOR \SUBBYTES[4].a/U4082  ( .A(\w1[4][105] ), .B(\SUBBYTES[4].a/w575 ), .Z(
        \SUBBYTES[4].a/w579 ) );
  XOR \SUBBYTES[4].a/U4081  ( .A(\w1[4][108] ), .B(\SUBBYTES[4].a/w575 ), .Z(
        \SUBBYTES[4].a/w580 ) );
  XOR \SUBBYTES[4].a/U4080  ( .A(\SUBBYTES[4].a/w579 ), .B(n10921), .Z(
        \SUBBYTES[4].a/w581 ) );
  XOR \SUBBYTES[4].a/U4079  ( .A(n10921), .B(n10633), .Z(\SUBBYTES[4].a/w666 )
         );
  XOR \SUBBYTES[4].a/U4078  ( .A(\w1[4][108] ), .B(\w1[4][105] ), .Z(n10633)
         );
  XOR \SUBBYTES[4].a/U4077  ( .A(n10635), .B(n10634), .Z(n10918) );
  XOR \SUBBYTES[4].a/U4076  ( .A(\w1[4][108] ), .B(n10636), .Z(n10634) );
  XOR \SUBBYTES[4].a/U4075  ( .A(\SUBBYTES[4].a/w631 ), .B(\w1[4][110] ), .Z(
        n10635) );
  XOR \SUBBYTES[4].a/U4074  ( .A(\SUBBYTES[4].a/w605 ), .B(
        \SUBBYTES[4].a/w612 ), .Z(n10636) );
  XOR \SUBBYTES[4].a/U4073  ( .A(n10638), .B(n10637), .Z(n10916) );
  XOR \SUBBYTES[4].a/U4072  ( .A(\w1[4][105] ), .B(n10639), .Z(n10637) );
  XOR \SUBBYTES[4].a/U4071  ( .A(\SUBBYTES[4].a/w630 ), .B(\w1[4][109] ), .Z(
        n10638) );
  XOR \SUBBYTES[4].a/U4070  ( .A(\SUBBYTES[4].a/w606 ), .B(
        \SUBBYTES[4].a/w613 ), .Z(n10639) );
  XOR \SUBBYTES[4].a/U4069  ( .A(n10918), .B(n10916), .Z(\SUBBYTES[4].a/w636 )
         );
  XOR \SUBBYTES[4].a/U4068  ( .A(\w1[4][109] ), .B(n10640), .Z(n10919) );
  XOR \SUBBYTES[4].a/U4067  ( .A(\SUBBYTES[4].a/w598 ), .B(
        \SUBBYTES[4].a/w608 ), .Z(n10640) );
  XOR \SUBBYTES[4].a/U4066  ( .A(n10642), .B(n10641), .Z(\SUBBYTES[4].a/w623 )
         );
  XOR \SUBBYTES[4].a/U4065  ( .A(n10919), .B(n10643), .Z(n10641) );
  XOR \SUBBYTES[4].a/U4064  ( .A(\w1[4][108] ), .B(\SUBBYTES[4].a/w687 ), .Z(
        n10642) );
  XOR \SUBBYTES[4].a/U4063  ( .A(\SUBBYTES[4].a/w600 ), .B(
        \SUBBYTES[4].a/w605 ), .Z(n10643) );
  XOR \SUBBYTES[4].a/U4062  ( .A(n10645), .B(n10644), .Z(n10917) );
  XOR \SUBBYTES[4].a/U4061  ( .A(\SUBBYTES[4].a/w633 ), .B(\w1[4][111] ), .Z(
        n10644) );
  XOR \SUBBYTES[4].a/U4060  ( .A(\SUBBYTES[4].a/w608 ), .B(
        \SUBBYTES[4].a/w615 ), .Z(n10645) );
  XOR \SUBBYTES[4].a/U4059  ( .A(n10916), .B(n10917), .Z(\SUBBYTES[4].a/w635 )
         );
  XOR \SUBBYTES[4].a/U4058  ( .A(\w1[4][107] ), .B(n10646), .Z(n10920) );
  XOR \SUBBYTES[4].a/U4057  ( .A(\SUBBYTES[4].a/w597 ), .B(
        \SUBBYTES[4].a/w600 ), .Z(n10646) );
  XOR \SUBBYTES[4].a/U4056  ( .A(n10648), .B(n10647), .Z(\SUBBYTES[4].a/w624 )
         );
  XOR \SUBBYTES[4].a/U4055  ( .A(n10920), .B(n10649), .Z(n10647) );
  XOR \SUBBYTES[4].a/U4054  ( .A(\w1[4][110] ), .B(\SUBBYTES[4].a/w666 ), .Z(
        n10648) );
  XOR \SUBBYTES[4].a/U4053  ( .A(\SUBBYTES[4].a/w605 ), .B(
        \SUBBYTES[4].a/w606 ), .Z(n10649) );
  XOR \SUBBYTES[4].a/U4052  ( .A(n10918), .B(n10917), .Z(\SUBBYTES[4].a/w644 )
         );
  XOR \SUBBYTES[4].a/U4051  ( .A(n10651), .B(n10650), .Z(\SUBBYTES[4].a/w645 )
         );
  XOR \SUBBYTES[4].a/U4050  ( .A(\w1[4][111] ), .B(n10919), .Z(n10650) );
  XOR \SUBBYTES[4].a/U4049  ( .A(\SUBBYTES[4].a/w597 ), .B(
        \SUBBYTES[4].a/w606 ), .Z(n10651) );
  XOR \SUBBYTES[4].a/U4048  ( .A(n10653), .B(n10652), .Z(\SUBBYTES[4].a/w621 )
         );
  XOR \SUBBYTES[4].a/U4047  ( .A(n10655), .B(n10654), .Z(n10652) );
  XOR \SUBBYTES[4].a/U4046  ( .A(\w1[4][111] ), .B(\SUBBYTES[4].a/w705 ), .Z(
        n10653) );
  XOR \SUBBYTES[4].a/U4045  ( .A(\SUBBYTES[4].a/w612 ), .B(
        \SUBBYTES[4].a/w615 ), .Z(n10654) );
  XOR \SUBBYTES[4].a/U4044  ( .A(\SUBBYTES[4].a/w598 ), .B(
        \SUBBYTES[4].a/w600 ), .Z(n10655) );
  XOR \SUBBYTES[4].a/U4043  ( .A(n10657), .B(n10656), .Z(\SUBBYTES[4].a/w622 )
         );
  XOR \SUBBYTES[4].a/U4042  ( .A(n10920), .B(n10658), .Z(n10656) );
  XOR \SUBBYTES[4].a/U4041  ( .A(\w1[4][109] ), .B(n10921), .Z(n10657) );
  XOR \SUBBYTES[4].a/U4040  ( .A(\SUBBYTES[4].a/w612 ), .B(
        \SUBBYTES[4].a/w613 ), .Z(n10658) );
  XOR \SUBBYTES[4].a/U4039  ( .A(n10660), .B(n10659), .Z(\SUBBYTES[4].a/w638 )
         );
  XOR \SUBBYTES[4].a/U4038  ( .A(\w1[4][105] ), .B(n10661), .Z(n10659) );
  XOR \SUBBYTES[4].a/U4037  ( .A(\SUBBYTES[4].a/w613 ), .B(
        \SUBBYTES[4].a/w615 ), .Z(n10660) );
  XOR \SUBBYTES[4].a/U4036  ( .A(\SUBBYTES[4].a/w597 ), .B(
        \SUBBYTES[4].a/w598 ), .Z(n10661) );
  XOR \SUBBYTES[4].a/U4035  ( .A(\w1[4][113] ), .B(n10662), .Z(n10922) );
  XOR \SUBBYTES[4].a/U4034  ( .A(\w1[4][115] ), .B(\w1[4][114] ), .Z(n10662)
         );
  XOR \SUBBYTES[4].a/U4033  ( .A(\w1[4][118] ), .B(n10922), .Z(
        \SUBBYTES[4].a/w480 ) );
  XOR \SUBBYTES[4].a/U4032  ( .A(\w1[4][112] ), .B(\SUBBYTES[4].a/w480 ), .Z(
        \SUBBYTES[4].a/w367 ) );
  XOR \SUBBYTES[4].a/U4031  ( .A(\w1[4][112] ), .B(n10663), .Z(
        \SUBBYTES[4].a/w368 ) );
  XOR \SUBBYTES[4].a/U4030  ( .A(\w1[4][118] ), .B(\w1[4][117] ), .Z(n10663)
         );
  XOR \SUBBYTES[4].a/U4029  ( .A(\w1[4][117] ), .B(n10922), .Z(
        \SUBBYTES[4].a/w498 ) );
  XOR \SUBBYTES[4].a/U4028  ( .A(n10665), .B(n10664), .Z(\SUBBYTES[4].a/w491 )
         );
  XOR \SUBBYTES[4].a/U4027  ( .A(\w1[4][115] ), .B(\w1[4][113] ), .Z(n10664)
         );
  XOR \SUBBYTES[4].a/U4026  ( .A(\w1[4][119] ), .B(\w1[4][116] ), .Z(n10665)
         );
  XOR \SUBBYTES[4].a/U4025  ( .A(\w1[4][112] ), .B(\SUBBYTES[4].a/w491 ), .Z(
        \SUBBYTES[4].a/w370 ) );
  XOR \SUBBYTES[4].a/U4024  ( .A(n10667), .B(n10666), .Z(\SUBBYTES[4].a/w478 )
         );
  XOR \SUBBYTES[4].a/U4023  ( .A(\SUBBYTES[4].a/w439 ), .B(n1006), .Z(n10666)
         );
  XOR \SUBBYTES[4].a/U4022  ( .A(\SUBBYTES[4].a/w432 ), .B(
        \SUBBYTES[4].a/w435 ), .Z(n10667) );
  XOR \SUBBYTES[4].a/U4021  ( .A(n10669), .B(n10668), .Z(\SUBBYTES[4].a/w479 )
         );
  XOR \SUBBYTES[4].a/U4020  ( .A(\SUBBYTES[4].a/w439 ), .B(n9675), .Z(n10668)
         );
  XOR \SUBBYTES[4].a/U4019  ( .A(\SUBBYTES[4].a/w432 ), .B(n9674), .Z(n10669)
         );
  XOR \SUBBYTES[4].a/U4018  ( .A(\SUBBYTES[4].a/w491 ), .B(n10670), .Z(
        \SUBBYTES[4].a/w481 ) );
  XOR \SUBBYTES[4].a/U4017  ( .A(\w1[4][118] ), .B(\w1[4][117] ), .Z(n10670)
         );
  XOR \SUBBYTES[4].a/U4016  ( .A(n10672), .B(n10671), .Z(\SUBBYTES[4].a/w482 )
         );
  XOR \SUBBYTES[4].a/U4015  ( .A(n9675), .B(n1006), .Z(n10671) );
  XOR \SUBBYTES[4].a/U4014  ( .A(n9674), .B(\SUBBYTES[4].a/w435 ), .Z(n10672)
         );
  XOR \SUBBYTES[4].a/U4013  ( .A(\w1[4][119] ), .B(\w1[4][114] ), .Z(n10928)
         );
  XOR \SUBBYTES[4].a/U4012  ( .A(n10928), .B(n10673), .Z(\SUBBYTES[4].a/w483 )
         );
  XOR \SUBBYTES[4].a/U4011  ( .A(\w1[4][117] ), .B(\w1[4][116] ), .Z(n10673)
         );
  XOR \SUBBYTES[4].a/U4010  ( .A(\w1[4][119] ), .B(\SUBBYTES[4].a/w368 ), .Z(
        \SUBBYTES[4].a/w371 ) );
  XOR \SUBBYTES[4].a/U4009  ( .A(\w1[4][113] ), .B(\SUBBYTES[4].a/w368 ), .Z(
        \SUBBYTES[4].a/w372 ) );
  XOR \SUBBYTES[4].a/U4008  ( .A(\w1[4][116] ), .B(\SUBBYTES[4].a/w368 ), .Z(
        \SUBBYTES[4].a/w373 ) );
  XOR \SUBBYTES[4].a/U4007  ( .A(\SUBBYTES[4].a/w372 ), .B(n10928), .Z(
        \SUBBYTES[4].a/w374 ) );
  XOR \SUBBYTES[4].a/U4006  ( .A(n10928), .B(n10674), .Z(\SUBBYTES[4].a/w459 )
         );
  XOR \SUBBYTES[4].a/U4005  ( .A(\w1[4][116] ), .B(\w1[4][113] ), .Z(n10674)
         );
  XOR \SUBBYTES[4].a/U4004  ( .A(n10676), .B(n10675), .Z(n10925) );
  XOR \SUBBYTES[4].a/U4003  ( .A(\w1[4][116] ), .B(n10677), .Z(n10675) );
  XOR \SUBBYTES[4].a/U4002  ( .A(\SUBBYTES[4].a/w424 ), .B(\w1[4][118] ), .Z(
        n10676) );
  XOR \SUBBYTES[4].a/U4001  ( .A(\SUBBYTES[4].a/w398 ), .B(
        \SUBBYTES[4].a/w405 ), .Z(n10677) );
  XOR \SUBBYTES[4].a/U4000  ( .A(n10679), .B(n10678), .Z(n10923) );
  XOR \SUBBYTES[4].a/U3999  ( .A(\w1[4][113] ), .B(n10680), .Z(n10678) );
  XOR \SUBBYTES[4].a/U3998  ( .A(\SUBBYTES[4].a/w423 ), .B(\w1[4][117] ), .Z(
        n10679) );
  XOR \SUBBYTES[4].a/U3997  ( .A(\SUBBYTES[4].a/w399 ), .B(
        \SUBBYTES[4].a/w406 ), .Z(n10680) );
  XOR \SUBBYTES[4].a/U3996  ( .A(n10925), .B(n10923), .Z(\SUBBYTES[4].a/w429 )
         );
  XOR \SUBBYTES[4].a/U3995  ( .A(\w1[4][117] ), .B(n10681), .Z(n10926) );
  XOR \SUBBYTES[4].a/U3994  ( .A(\SUBBYTES[4].a/w391 ), .B(
        \SUBBYTES[4].a/w401 ), .Z(n10681) );
  XOR \SUBBYTES[4].a/U3993  ( .A(n10683), .B(n10682), .Z(\SUBBYTES[4].a/w416 )
         );
  XOR \SUBBYTES[4].a/U3992  ( .A(n10926), .B(n10684), .Z(n10682) );
  XOR \SUBBYTES[4].a/U3991  ( .A(\w1[4][116] ), .B(\SUBBYTES[4].a/w480 ), .Z(
        n10683) );
  XOR \SUBBYTES[4].a/U3990  ( .A(\SUBBYTES[4].a/w393 ), .B(
        \SUBBYTES[4].a/w398 ), .Z(n10684) );
  XOR \SUBBYTES[4].a/U3989  ( .A(n10686), .B(n10685), .Z(n10924) );
  XOR \SUBBYTES[4].a/U3988  ( .A(\SUBBYTES[4].a/w426 ), .B(\w1[4][119] ), .Z(
        n10685) );
  XOR \SUBBYTES[4].a/U3987  ( .A(\SUBBYTES[4].a/w401 ), .B(
        \SUBBYTES[4].a/w408 ), .Z(n10686) );
  XOR \SUBBYTES[4].a/U3986  ( .A(n10923), .B(n10924), .Z(\SUBBYTES[4].a/w428 )
         );
  XOR \SUBBYTES[4].a/U3985  ( .A(\w1[4][115] ), .B(n10687), .Z(n10927) );
  XOR \SUBBYTES[4].a/U3984  ( .A(\SUBBYTES[4].a/w390 ), .B(
        \SUBBYTES[4].a/w393 ), .Z(n10687) );
  XOR \SUBBYTES[4].a/U3983  ( .A(n10689), .B(n10688), .Z(\SUBBYTES[4].a/w417 )
         );
  XOR \SUBBYTES[4].a/U3982  ( .A(n10927), .B(n10690), .Z(n10688) );
  XOR \SUBBYTES[4].a/U3981  ( .A(\w1[4][118] ), .B(\SUBBYTES[4].a/w459 ), .Z(
        n10689) );
  XOR \SUBBYTES[4].a/U3980  ( .A(\SUBBYTES[4].a/w398 ), .B(
        \SUBBYTES[4].a/w399 ), .Z(n10690) );
  XOR \SUBBYTES[4].a/U3979  ( .A(n10925), .B(n10924), .Z(\SUBBYTES[4].a/w437 )
         );
  XOR \SUBBYTES[4].a/U3978  ( .A(n10692), .B(n10691), .Z(\SUBBYTES[4].a/w438 )
         );
  XOR \SUBBYTES[4].a/U3977  ( .A(\w1[4][119] ), .B(n10926), .Z(n10691) );
  XOR \SUBBYTES[4].a/U3976  ( .A(\SUBBYTES[4].a/w390 ), .B(
        \SUBBYTES[4].a/w399 ), .Z(n10692) );
  XOR \SUBBYTES[4].a/U3975  ( .A(n10694), .B(n10693), .Z(\SUBBYTES[4].a/w414 )
         );
  XOR \SUBBYTES[4].a/U3974  ( .A(n10696), .B(n10695), .Z(n10693) );
  XOR \SUBBYTES[4].a/U3973  ( .A(\w1[4][119] ), .B(\SUBBYTES[4].a/w498 ), .Z(
        n10694) );
  XOR \SUBBYTES[4].a/U3972  ( .A(\SUBBYTES[4].a/w405 ), .B(
        \SUBBYTES[4].a/w408 ), .Z(n10695) );
  XOR \SUBBYTES[4].a/U3971  ( .A(\SUBBYTES[4].a/w391 ), .B(
        \SUBBYTES[4].a/w393 ), .Z(n10696) );
  XOR \SUBBYTES[4].a/U3970  ( .A(n10698), .B(n10697), .Z(\SUBBYTES[4].a/w415 )
         );
  XOR \SUBBYTES[4].a/U3969  ( .A(n10927), .B(n10699), .Z(n10697) );
  XOR \SUBBYTES[4].a/U3968  ( .A(\w1[4][117] ), .B(n10928), .Z(n10698) );
  XOR \SUBBYTES[4].a/U3967  ( .A(\SUBBYTES[4].a/w405 ), .B(
        \SUBBYTES[4].a/w406 ), .Z(n10699) );
  XOR \SUBBYTES[4].a/U3966  ( .A(n10701), .B(n10700), .Z(\SUBBYTES[4].a/w431 )
         );
  XOR \SUBBYTES[4].a/U3965  ( .A(\w1[4][113] ), .B(n10702), .Z(n10700) );
  XOR \SUBBYTES[4].a/U3964  ( .A(\SUBBYTES[4].a/w406 ), .B(
        \SUBBYTES[4].a/w408 ), .Z(n10701) );
  XOR \SUBBYTES[4].a/U3963  ( .A(\SUBBYTES[4].a/w390 ), .B(
        \SUBBYTES[4].a/w391 ), .Z(n10702) );
  XOR \SUBBYTES[4].a/U3962  ( .A(\w1[4][121] ), .B(n10703), .Z(n10929) );
  XOR \SUBBYTES[4].a/U3961  ( .A(\w1[4][123] ), .B(\w1[4][122] ), .Z(n10703)
         );
  XOR \SUBBYTES[4].a/U3960  ( .A(\w1[4][126] ), .B(n10929), .Z(
        \SUBBYTES[4].a/w273 ) );
  XOR \SUBBYTES[4].a/U3959  ( .A(\w1[4][120] ), .B(\SUBBYTES[4].a/w273 ), .Z(
        \SUBBYTES[4].a/w160 ) );
  XOR \SUBBYTES[4].a/U3958  ( .A(\w1[4][120] ), .B(n10704), .Z(
        \SUBBYTES[4].a/w161 ) );
  XOR \SUBBYTES[4].a/U3957  ( .A(\w1[4][126] ), .B(\w1[4][125] ), .Z(n10704)
         );
  XOR \SUBBYTES[4].a/U3956  ( .A(\w1[4][125] ), .B(n10929), .Z(
        \SUBBYTES[4].a/w291 ) );
  XOR \SUBBYTES[4].a/U3955  ( .A(n10706), .B(n10705), .Z(\SUBBYTES[4].a/w284 )
         );
  XOR \SUBBYTES[4].a/U3954  ( .A(\w1[4][123] ), .B(\w1[4][121] ), .Z(n10705)
         );
  XOR \SUBBYTES[4].a/U3953  ( .A(\w1[4][127] ), .B(\w1[4][124] ), .Z(n10706)
         );
  XOR \SUBBYTES[4].a/U3952  ( .A(\w1[4][120] ), .B(\SUBBYTES[4].a/w284 ), .Z(
        \SUBBYTES[4].a/w163 ) );
  XOR \SUBBYTES[4].a/U3951  ( .A(n10708), .B(n10707), .Z(\SUBBYTES[4].a/w271 )
         );
  XOR \SUBBYTES[4].a/U3950  ( .A(\SUBBYTES[4].a/w232 ), .B(n1005), .Z(n10707)
         );
  XOR \SUBBYTES[4].a/U3949  ( .A(\SUBBYTES[4].a/w225 ), .B(
        \SUBBYTES[4].a/w228 ), .Z(n10708) );
  XOR \SUBBYTES[4].a/U3948  ( .A(n10710), .B(n10709), .Z(\SUBBYTES[4].a/w272 )
         );
  XOR \SUBBYTES[4].a/U3947  ( .A(\SUBBYTES[4].a/w232 ), .B(n9673), .Z(n10709)
         );
  XOR \SUBBYTES[4].a/U3946  ( .A(\SUBBYTES[4].a/w225 ), .B(n9672), .Z(n10710)
         );
  XOR \SUBBYTES[4].a/U3945  ( .A(\SUBBYTES[4].a/w284 ), .B(n10711), .Z(
        \SUBBYTES[4].a/w274 ) );
  XOR \SUBBYTES[4].a/U3944  ( .A(\w1[4][126] ), .B(\w1[4][125] ), .Z(n10711)
         );
  XOR \SUBBYTES[4].a/U3943  ( .A(n10713), .B(n10712), .Z(\SUBBYTES[4].a/w275 )
         );
  XOR \SUBBYTES[4].a/U3942  ( .A(n9673), .B(n1005), .Z(n10712) );
  XOR \SUBBYTES[4].a/U3941  ( .A(n9672), .B(\SUBBYTES[4].a/w228 ), .Z(n10713)
         );
  XOR \SUBBYTES[4].a/U3940  ( .A(\w1[4][127] ), .B(\w1[4][122] ), .Z(n10935)
         );
  XOR \SUBBYTES[4].a/U3939  ( .A(n10935), .B(n10714), .Z(\SUBBYTES[4].a/w276 )
         );
  XOR \SUBBYTES[4].a/U3938  ( .A(\w1[4][125] ), .B(\w1[4][124] ), .Z(n10714)
         );
  XOR \SUBBYTES[4].a/U3937  ( .A(\w1[4][127] ), .B(\SUBBYTES[4].a/w161 ), .Z(
        \SUBBYTES[4].a/w164 ) );
  XOR \SUBBYTES[4].a/U3936  ( .A(\w1[4][121] ), .B(\SUBBYTES[4].a/w161 ), .Z(
        \SUBBYTES[4].a/w165 ) );
  XOR \SUBBYTES[4].a/U3935  ( .A(\w1[4][124] ), .B(\SUBBYTES[4].a/w161 ), .Z(
        \SUBBYTES[4].a/w166 ) );
  XOR \SUBBYTES[4].a/U3934  ( .A(\SUBBYTES[4].a/w165 ), .B(n10935), .Z(
        \SUBBYTES[4].a/w167 ) );
  XOR \SUBBYTES[4].a/U3933  ( .A(n10935), .B(n10715), .Z(\SUBBYTES[4].a/w252 )
         );
  XOR \SUBBYTES[4].a/U3932  ( .A(\w1[4][124] ), .B(\w1[4][121] ), .Z(n10715)
         );
  XOR \SUBBYTES[4].a/U3931  ( .A(n10717), .B(n10716), .Z(n10932) );
  XOR \SUBBYTES[4].a/U3930  ( .A(\w1[4][124] ), .B(n10718), .Z(n10716) );
  XOR \SUBBYTES[4].a/U3929  ( .A(\SUBBYTES[4].a/w217 ), .B(\w1[4][126] ), .Z(
        n10717) );
  XOR \SUBBYTES[4].a/U3928  ( .A(\SUBBYTES[4].a/w191 ), .B(
        \SUBBYTES[4].a/w198 ), .Z(n10718) );
  XOR \SUBBYTES[4].a/U3927  ( .A(n10720), .B(n10719), .Z(n10930) );
  XOR \SUBBYTES[4].a/U3926  ( .A(\w1[4][121] ), .B(n10721), .Z(n10719) );
  XOR \SUBBYTES[4].a/U3925  ( .A(\SUBBYTES[4].a/w216 ), .B(\w1[4][125] ), .Z(
        n10720) );
  XOR \SUBBYTES[4].a/U3924  ( .A(\SUBBYTES[4].a/w192 ), .B(
        \SUBBYTES[4].a/w199 ), .Z(n10721) );
  XOR \SUBBYTES[4].a/U3923  ( .A(n10932), .B(n10930), .Z(\SUBBYTES[4].a/w222 )
         );
  XOR \SUBBYTES[4].a/U3922  ( .A(\w1[4][125] ), .B(n10722), .Z(n10933) );
  XOR \SUBBYTES[4].a/U3921  ( .A(\SUBBYTES[4].a/w184 ), .B(
        \SUBBYTES[4].a/w194 ), .Z(n10722) );
  XOR \SUBBYTES[4].a/U3920  ( .A(n10724), .B(n10723), .Z(\SUBBYTES[4].a/w209 )
         );
  XOR \SUBBYTES[4].a/U3919  ( .A(n10933), .B(n10725), .Z(n10723) );
  XOR \SUBBYTES[4].a/U3918  ( .A(\w1[4][124] ), .B(\SUBBYTES[4].a/w273 ), .Z(
        n10724) );
  XOR \SUBBYTES[4].a/U3917  ( .A(\SUBBYTES[4].a/w186 ), .B(
        \SUBBYTES[4].a/w191 ), .Z(n10725) );
  XOR \SUBBYTES[4].a/U3916  ( .A(n10727), .B(n10726), .Z(n10931) );
  XOR \SUBBYTES[4].a/U3915  ( .A(\SUBBYTES[4].a/w219 ), .B(\w1[4][127] ), .Z(
        n10726) );
  XOR \SUBBYTES[4].a/U3914  ( .A(\SUBBYTES[4].a/w194 ), .B(
        \SUBBYTES[4].a/w201 ), .Z(n10727) );
  XOR \SUBBYTES[4].a/U3913  ( .A(n10930), .B(n10931), .Z(\SUBBYTES[4].a/w221 )
         );
  XOR \SUBBYTES[4].a/U3912  ( .A(\w1[4][123] ), .B(n10728), .Z(n10934) );
  XOR \SUBBYTES[4].a/U3911  ( .A(\SUBBYTES[4].a/w183 ), .B(
        \SUBBYTES[4].a/w186 ), .Z(n10728) );
  XOR \SUBBYTES[4].a/U3910  ( .A(n10730), .B(n10729), .Z(\SUBBYTES[4].a/w210 )
         );
  XOR \SUBBYTES[4].a/U3909  ( .A(n10934), .B(n10731), .Z(n10729) );
  XOR \SUBBYTES[4].a/U3908  ( .A(\w1[4][126] ), .B(\SUBBYTES[4].a/w252 ), .Z(
        n10730) );
  XOR \SUBBYTES[4].a/U3907  ( .A(\SUBBYTES[4].a/w191 ), .B(
        \SUBBYTES[4].a/w192 ), .Z(n10731) );
  XOR \SUBBYTES[4].a/U3906  ( .A(n10932), .B(n10931), .Z(\SUBBYTES[4].a/w230 )
         );
  XOR \SUBBYTES[4].a/U3905  ( .A(n10733), .B(n10732), .Z(\SUBBYTES[4].a/w231 )
         );
  XOR \SUBBYTES[4].a/U3904  ( .A(\w1[4][127] ), .B(n10933), .Z(n10732) );
  XOR \SUBBYTES[4].a/U3903  ( .A(\SUBBYTES[4].a/w183 ), .B(
        \SUBBYTES[4].a/w192 ), .Z(n10733) );
  XOR \SUBBYTES[4].a/U3902  ( .A(n10735), .B(n10734), .Z(\SUBBYTES[4].a/w207 )
         );
  XOR \SUBBYTES[4].a/U3901  ( .A(n10737), .B(n10736), .Z(n10734) );
  XOR \SUBBYTES[4].a/U3900  ( .A(\w1[4][127] ), .B(\SUBBYTES[4].a/w291 ), .Z(
        n10735) );
  XOR \SUBBYTES[4].a/U3899  ( .A(\SUBBYTES[4].a/w198 ), .B(
        \SUBBYTES[4].a/w201 ), .Z(n10736) );
  XOR \SUBBYTES[4].a/U3898  ( .A(\SUBBYTES[4].a/w184 ), .B(
        \SUBBYTES[4].a/w186 ), .Z(n10737) );
  XOR \SUBBYTES[4].a/U3897  ( .A(n10739), .B(n10738), .Z(\SUBBYTES[4].a/w208 )
         );
  XOR \SUBBYTES[4].a/U3896  ( .A(n10934), .B(n10740), .Z(n10738) );
  XOR \SUBBYTES[4].a/U3895  ( .A(\w1[4][125] ), .B(n10935), .Z(n10739) );
  XOR \SUBBYTES[4].a/U3894  ( .A(\SUBBYTES[4].a/w198 ), .B(
        \SUBBYTES[4].a/w199 ), .Z(n10740) );
  XOR \SUBBYTES[4].a/U3893  ( .A(n10742), .B(n10741), .Z(\SUBBYTES[4].a/w224 )
         );
  XOR \SUBBYTES[4].a/U3892  ( .A(\w1[4][121] ), .B(n10743), .Z(n10741) );
  XOR \SUBBYTES[4].a/U3891  ( .A(\SUBBYTES[4].a/w199 ), .B(
        \SUBBYTES[4].a/w201 ), .Z(n10742) );
  XOR \SUBBYTES[4].a/U3890  ( .A(\SUBBYTES[4].a/w183 ), .B(
        \SUBBYTES[4].a/w184 ), .Z(n10743) );
  XOR \SUBBYTES[3].a/U5649  ( .A(\SUBBYTES[3].a/w3390 ), .B(
        \SUBBYTES[3].a/w3391 ), .Z(n9465) );
  XOR \SUBBYTES[3].a/U5648  ( .A(n9465), .B(n8424), .Z(n9464) );
  XOR \SUBBYTES[3].a/U5647  ( .A(\SUBBYTES[3].a/w3383 ), .B(
        \SUBBYTES[3].a/w3400 ), .Z(n8424) );
  XOR \SUBBYTES[3].a/U5645  ( .A(\SUBBYTES[3].a/w3382 ), .B(
        \SUBBYTES[3].a/w3397 ), .Z(n8425) );
  XOR \SUBBYTES[3].a/U5644  ( .A(n9465), .B(n8426), .Z(n9656) );
  XOR \SUBBYTES[3].a/U5643  ( .A(\SUBBYTES[3].a/w3397 ), .B(
        \SUBBYTES[3].a/w3398 ), .Z(n8426) );
  XOR \SUBBYTES[3].a/U5642  ( .A(\SUBBYTES[3].a/w3359 ), .B(n8427), .Z(n9467)
         );
  XOR \SUBBYTES[3].a/U5641  ( .A(\SUBBYTES[3].a/w3350 ), .B(
        \SUBBYTES[3].a/w3351 ), .Z(n8427) );
  XOR \SUBBYTES[3].a/U5639  ( .A(\SUBBYTES[3].a/w3361 ), .B(n9656), .Z(n8428)
         );
  XOR \SUBBYTES[3].a/U5638  ( .A(n8430), .B(n8429), .Z(n9468) );
  XOR \SUBBYTES[3].a/U5637  ( .A(n8432), .B(n8431), .Z(n8429) );
  XOR \SUBBYTES[3].a/U5636  ( .A(\SUBBYTES[3].a/w3397 ), .B(
        \SUBBYTES[3].a/w3398 ), .Z(n8430) );
  XOR \SUBBYTES[3].a/U5635  ( .A(\SUBBYTES[3].a/w3361 ), .B(
        \SUBBYTES[3].a/w3385 ), .Z(n8431) );
  XOR \SUBBYTES[3].a/U5634  ( .A(\SUBBYTES[3].a/w3350 ), .B(
        \SUBBYTES[3].a/w3359 ), .Z(n8432) );
  XOR \SUBBYTES[3].a/U5633  ( .A(\SUBBYTES[3].a/w3382 ), .B(n8433), .Z(n9466)
         );
  XOR \SUBBYTES[3].a/U5632  ( .A(\SUBBYTES[3].a/w3365 ), .B(
        \SUBBYTES[3].a/w3368 ), .Z(n8433) );
  XOR \SUBBYTES[3].a/U5630  ( .A(\SUBBYTES[3].a/w3353 ), .B(n9468), .Z(n8434)
         );
  XOR \SUBBYTES[3].a/U5628  ( .A(\SUBBYTES[3].a/w3385 ), .B(
        \SUBBYTES[3].a/w3398 ), .Z(n8435) );
  XOR \SUBBYTES[3].a/U5626  ( .A(n8439), .B(n8438), .Z(n8436) );
  XOR \SUBBYTES[3].a/U5625  ( .A(n8441), .B(n8440), .Z(n8437) );
  XOR \SUBBYTES[3].a/U5624  ( .A(\SUBBYTES[3].a/w3397 ), .B(
        \SUBBYTES[3].a/w3400 ), .Z(n8438) );
  XOR \SUBBYTES[3].a/U5623  ( .A(\SUBBYTES[3].a/w3390 ), .B(
        \SUBBYTES[3].a/w3393 ), .Z(n8439) );
  XOR \SUBBYTES[3].a/U5622  ( .A(\SUBBYTES[3].a/w3365 ), .B(
        \SUBBYTES[3].a/w3366 ), .Z(n8440) );
  XOR \SUBBYTES[3].a/U5621  ( .A(\SUBBYTES[3].a/w3350 ), .B(
        \SUBBYTES[3].a/w3353 ), .Z(n8441) );
  XOR \SUBBYTES[3].a/U5619  ( .A(n9465), .B(n8444), .Z(n8442) );
  XOR \SUBBYTES[3].a/U5618  ( .A(n9467), .B(n9466), .Z(n8443) );
  XOR \SUBBYTES[3].a/U5617  ( .A(\SUBBYTES[3].a/w3358 ), .B(
        \SUBBYTES[3].a/w3385 ), .Z(n8444) );
  XOR \SUBBYTES[3].a/U5615  ( .A(n9468), .B(n8447), .Z(n8445) );
  XOR \SUBBYTES[3].a/U5614  ( .A(\SUBBYTES[3].a/w3391 ), .B(
        \SUBBYTES[3].a/w3393 ), .Z(n8446) );
  XOR \SUBBYTES[3].a/U5613  ( .A(\SUBBYTES[3].a/w3351 ), .B(
        \SUBBYTES[3].a/w3383 ), .Z(n8447) );
  XOR \SUBBYTES[3].a/U5612  ( .A(\SUBBYTES[3].a/w3183 ), .B(
        \SUBBYTES[3].a/w3184 ), .Z(n9470) );
  XOR \SUBBYTES[3].a/U5611  ( .A(n9470), .B(n8448), .Z(n9469) );
  XOR \SUBBYTES[3].a/U5610  ( .A(\SUBBYTES[3].a/w3176 ), .B(
        \SUBBYTES[3].a/w3193 ), .Z(n8448) );
  XOR \SUBBYTES[3].a/U5608  ( .A(\SUBBYTES[3].a/w3175 ), .B(
        \SUBBYTES[3].a/w3190 ), .Z(n8449) );
  XOR \SUBBYTES[3].a/U5607  ( .A(n9470), .B(n8450), .Z(n9657) );
  XOR \SUBBYTES[3].a/U5606  ( .A(\SUBBYTES[3].a/w3190 ), .B(
        \SUBBYTES[3].a/w3191 ), .Z(n8450) );
  XOR \SUBBYTES[3].a/U5605  ( .A(\SUBBYTES[3].a/w3152 ), .B(n8451), .Z(n9472)
         );
  XOR \SUBBYTES[3].a/U5604  ( .A(\SUBBYTES[3].a/w3143 ), .B(
        \SUBBYTES[3].a/w3144 ), .Z(n8451) );
  XOR \SUBBYTES[3].a/U5602  ( .A(\SUBBYTES[3].a/w3154 ), .B(n9657), .Z(n8452)
         );
  XOR \SUBBYTES[3].a/U5601  ( .A(n8454), .B(n8453), .Z(n9473) );
  XOR \SUBBYTES[3].a/U5600  ( .A(n8456), .B(n8455), .Z(n8453) );
  XOR \SUBBYTES[3].a/U5599  ( .A(\SUBBYTES[3].a/w3190 ), .B(
        \SUBBYTES[3].a/w3191 ), .Z(n8454) );
  XOR \SUBBYTES[3].a/U5598  ( .A(\SUBBYTES[3].a/w3154 ), .B(
        \SUBBYTES[3].a/w3178 ), .Z(n8455) );
  XOR \SUBBYTES[3].a/U5597  ( .A(\SUBBYTES[3].a/w3143 ), .B(
        \SUBBYTES[3].a/w3152 ), .Z(n8456) );
  XOR \SUBBYTES[3].a/U5596  ( .A(\SUBBYTES[3].a/w3175 ), .B(n8457), .Z(n9471)
         );
  XOR \SUBBYTES[3].a/U5595  ( .A(\SUBBYTES[3].a/w3158 ), .B(
        \SUBBYTES[3].a/w3161 ), .Z(n8457) );
  XOR \SUBBYTES[3].a/U5593  ( .A(\SUBBYTES[3].a/w3146 ), .B(n9473), .Z(n8458)
         );
  XOR \SUBBYTES[3].a/U5591  ( .A(\SUBBYTES[3].a/w3178 ), .B(
        \SUBBYTES[3].a/w3191 ), .Z(n8459) );
  XOR \SUBBYTES[3].a/U5589  ( .A(n8463), .B(n8462), .Z(n8460) );
  XOR \SUBBYTES[3].a/U5588  ( .A(n8465), .B(n8464), .Z(n8461) );
  XOR \SUBBYTES[3].a/U5587  ( .A(\SUBBYTES[3].a/w3190 ), .B(
        \SUBBYTES[3].a/w3193 ), .Z(n8462) );
  XOR \SUBBYTES[3].a/U5586  ( .A(\SUBBYTES[3].a/w3183 ), .B(
        \SUBBYTES[3].a/w3186 ), .Z(n8463) );
  XOR \SUBBYTES[3].a/U5585  ( .A(\SUBBYTES[3].a/w3158 ), .B(
        \SUBBYTES[3].a/w3159 ), .Z(n8464) );
  XOR \SUBBYTES[3].a/U5584  ( .A(\SUBBYTES[3].a/w3143 ), .B(
        \SUBBYTES[3].a/w3146 ), .Z(n8465) );
  XOR \SUBBYTES[3].a/U5582  ( .A(n9470), .B(n8468), .Z(n8466) );
  XOR \SUBBYTES[3].a/U5581  ( .A(n9472), .B(n9471), .Z(n8467) );
  XOR \SUBBYTES[3].a/U5580  ( .A(\SUBBYTES[3].a/w3151 ), .B(
        \SUBBYTES[3].a/w3178 ), .Z(n8468) );
  XOR \SUBBYTES[3].a/U5578  ( .A(n9473), .B(n8471), .Z(n8469) );
  XOR \SUBBYTES[3].a/U5577  ( .A(\SUBBYTES[3].a/w3184 ), .B(
        \SUBBYTES[3].a/w3186 ), .Z(n8470) );
  XOR \SUBBYTES[3].a/U5576  ( .A(\SUBBYTES[3].a/w3144 ), .B(
        \SUBBYTES[3].a/w3176 ), .Z(n8471) );
  XOR \SUBBYTES[3].a/U5575  ( .A(\SUBBYTES[3].a/w2976 ), .B(
        \SUBBYTES[3].a/w2977 ), .Z(n9475) );
  XOR \SUBBYTES[3].a/U5574  ( .A(n9475), .B(n8472), .Z(n9474) );
  XOR \SUBBYTES[3].a/U5573  ( .A(\SUBBYTES[3].a/w2969 ), .B(
        \SUBBYTES[3].a/w2986 ), .Z(n8472) );
  XOR \SUBBYTES[3].a/U5571  ( .A(\SUBBYTES[3].a/w2968 ), .B(
        \SUBBYTES[3].a/w2983 ), .Z(n8473) );
  XOR \SUBBYTES[3].a/U5570  ( .A(n9475), .B(n8474), .Z(n9658) );
  XOR \SUBBYTES[3].a/U5569  ( .A(\SUBBYTES[3].a/w2983 ), .B(
        \SUBBYTES[3].a/w2984 ), .Z(n8474) );
  XOR \SUBBYTES[3].a/U5568  ( .A(\SUBBYTES[3].a/w2945 ), .B(n8475), .Z(n9477)
         );
  XOR \SUBBYTES[3].a/U5567  ( .A(\SUBBYTES[3].a/w2936 ), .B(
        \SUBBYTES[3].a/w2937 ), .Z(n8475) );
  XOR \SUBBYTES[3].a/U5565  ( .A(\SUBBYTES[3].a/w2947 ), .B(n9658), .Z(n8476)
         );
  XOR \SUBBYTES[3].a/U5564  ( .A(n8478), .B(n8477), .Z(n9478) );
  XOR \SUBBYTES[3].a/U5563  ( .A(n8480), .B(n8479), .Z(n8477) );
  XOR \SUBBYTES[3].a/U5562  ( .A(\SUBBYTES[3].a/w2983 ), .B(
        \SUBBYTES[3].a/w2984 ), .Z(n8478) );
  XOR \SUBBYTES[3].a/U5561  ( .A(\SUBBYTES[3].a/w2947 ), .B(
        \SUBBYTES[3].a/w2971 ), .Z(n8479) );
  XOR \SUBBYTES[3].a/U5560  ( .A(\SUBBYTES[3].a/w2936 ), .B(
        \SUBBYTES[3].a/w2945 ), .Z(n8480) );
  XOR \SUBBYTES[3].a/U5559  ( .A(\SUBBYTES[3].a/w2968 ), .B(n8481), .Z(n9476)
         );
  XOR \SUBBYTES[3].a/U5558  ( .A(\SUBBYTES[3].a/w2951 ), .B(
        \SUBBYTES[3].a/w2954 ), .Z(n8481) );
  XOR \SUBBYTES[3].a/U5556  ( .A(\SUBBYTES[3].a/w2939 ), .B(n9478), .Z(n8482)
         );
  XOR \SUBBYTES[3].a/U5554  ( .A(\SUBBYTES[3].a/w2971 ), .B(
        \SUBBYTES[3].a/w2984 ), .Z(n8483) );
  XOR \SUBBYTES[3].a/U5552  ( .A(n8487), .B(n8486), .Z(n8484) );
  XOR \SUBBYTES[3].a/U5551  ( .A(n8489), .B(n8488), .Z(n8485) );
  XOR \SUBBYTES[3].a/U5550  ( .A(\SUBBYTES[3].a/w2983 ), .B(
        \SUBBYTES[3].a/w2986 ), .Z(n8486) );
  XOR \SUBBYTES[3].a/U5549  ( .A(\SUBBYTES[3].a/w2976 ), .B(
        \SUBBYTES[3].a/w2979 ), .Z(n8487) );
  XOR \SUBBYTES[3].a/U5548  ( .A(\SUBBYTES[3].a/w2951 ), .B(
        \SUBBYTES[3].a/w2952 ), .Z(n8488) );
  XOR \SUBBYTES[3].a/U5547  ( .A(\SUBBYTES[3].a/w2936 ), .B(
        \SUBBYTES[3].a/w2939 ), .Z(n8489) );
  XOR \SUBBYTES[3].a/U5545  ( .A(n9475), .B(n8492), .Z(n8490) );
  XOR \SUBBYTES[3].a/U5544  ( .A(n9477), .B(n9476), .Z(n8491) );
  XOR \SUBBYTES[3].a/U5543  ( .A(\SUBBYTES[3].a/w2944 ), .B(
        \SUBBYTES[3].a/w2971 ), .Z(n8492) );
  XOR \SUBBYTES[3].a/U5541  ( .A(n9478), .B(n8495), .Z(n8493) );
  XOR \SUBBYTES[3].a/U5540  ( .A(\SUBBYTES[3].a/w2977 ), .B(
        \SUBBYTES[3].a/w2979 ), .Z(n8494) );
  XOR \SUBBYTES[3].a/U5539  ( .A(\SUBBYTES[3].a/w2937 ), .B(
        \SUBBYTES[3].a/w2969 ), .Z(n8495) );
  XOR \SUBBYTES[3].a/U5538  ( .A(\SUBBYTES[3].a/w2769 ), .B(
        \SUBBYTES[3].a/w2770 ), .Z(n9480) );
  XOR \SUBBYTES[3].a/U5537  ( .A(n9480), .B(n8496), .Z(n9479) );
  XOR \SUBBYTES[3].a/U5536  ( .A(\SUBBYTES[3].a/w2762 ), .B(
        \SUBBYTES[3].a/w2779 ), .Z(n8496) );
  XOR \SUBBYTES[3].a/U5534  ( .A(\SUBBYTES[3].a/w2761 ), .B(
        \SUBBYTES[3].a/w2776 ), .Z(n8497) );
  XOR \SUBBYTES[3].a/U5533  ( .A(n9480), .B(n8498), .Z(n9659) );
  XOR \SUBBYTES[3].a/U5532  ( .A(\SUBBYTES[3].a/w2776 ), .B(
        \SUBBYTES[3].a/w2777 ), .Z(n8498) );
  XOR \SUBBYTES[3].a/U5531  ( .A(\SUBBYTES[3].a/w2738 ), .B(n8499), .Z(n9482)
         );
  XOR \SUBBYTES[3].a/U5530  ( .A(\SUBBYTES[3].a/w2729 ), .B(
        \SUBBYTES[3].a/w2730 ), .Z(n8499) );
  XOR \SUBBYTES[3].a/U5528  ( .A(\SUBBYTES[3].a/w2740 ), .B(n9659), .Z(n8500)
         );
  XOR \SUBBYTES[3].a/U5527  ( .A(n8502), .B(n8501), .Z(n9483) );
  XOR \SUBBYTES[3].a/U5526  ( .A(n8504), .B(n8503), .Z(n8501) );
  XOR \SUBBYTES[3].a/U5525  ( .A(\SUBBYTES[3].a/w2776 ), .B(
        \SUBBYTES[3].a/w2777 ), .Z(n8502) );
  XOR \SUBBYTES[3].a/U5524  ( .A(\SUBBYTES[3].a/w2740 ), .B(
        \SUBBYTES[3].a/w2764 ), .Z(n8503) );
  XOR \SUBBYTES[3].a/U5523  ( .A(\SUBBYTES[3].a/w2729 ), .B(
        \SUBBYTES[3].a/w2738 ), .Z(n8504) );
  XOR \SUBBYTES[3].a/U5522  ( .A(\SUBBYTES[3].a/w2761 ), .B(n8505), .Z(n9481)
         );
  XOR \SUBBYTES[3].a/U5521  ( .A(\SUBBYTES[3].a/w2744 ), .B(
        \SUBBYTES[3].a/w2747 ), .Z(n8505) );
  XOR \SUBBYTES[3].a/U5519  ( .A(\SUBBYTES[3].a/w2732 ), .B(n9483), .Z(n8506)
         );
  XOR \SUBBYTES[3].a/U5517  ( .A(\SUBBYTES[3].a/w2764 ), .B(
        \SUBBYTES[3].a/w2777 ), .Z(n8507) );
  XOR \SUBBYTES[3].a/U5515  ( .A(n8511), .B(n8510), .Z(n8508) );
  XOR \SUBBYTES[3].a/U5514  ( .A(n8513), .B(n8512), .Z(n8509) );
  XOR \SUBBYTES[3].a/U5513  ( .A(\SUBBYTES[3].a/w2776 ), .B(
        \SUBBYTES[3].a/w2779 ), .Z(n8510) );
  XOR \SUBBYTES[3].a/U5512  ( .A(\SUBBYTES[3].a/w2769 ), .B(
        \SUBBYTES[3].a/w2772 ), .Z(n8511) );
  XOR \SUBBYTES[3].a/U5511  ( .A(\SUBBYTES[3].a/w2744 ), .B(
        \SUBBYTES[3].a/w2745 ), .Z(n8512) );
  XOR \SUBBYTES[3].a/U5510  ( .A(\SUBBYTES[3].a/w2729 ), .B(
        \SUBBYTES[3].a/w2732 ), .Z(n8513) );
  XOR \SUBBYTES[3].a/U5508  ( .A(n9480), .B(n8516), .Z(n8514) );
  XOR \SUBBYTES[3].a/U5507  ( .A(n9482), .B(n9481), .Z(n8515) );
  XOR \SUBBYTES[3].a/U5506  ( .A(\SUBBYTES[3].a/w2737 ), .B(
        \SUBBYTES[3].a/w2764 ), .Z(n8516) );
  XOR \SUBBYTES[3].a/U5504  ( .A(n9483), .B(n8519), .Z(n8517) );
  XOR \SUBBYTES[3].a/U5503  ( .A(\SUBBYTES[3].a/w2770 ), .B(
        \SUBBYTES[3].a/w2772 ), .Z(n8518) );
  XOR \SUBBYTES[3].a/U5502  ( .A(\SUBBYTES[3].a/w2730 ), .B(
        \SUBBYTES[3].a/w2762 ), .Z(n8519) );
  XOR \SUBBYTES[3].a/U5501  ( .A(\SUBBYTES[3].a/w2562 ), .B(
        \SUBBYTES[3].a/w2563 ), .Z(n9485) );
  XOR \SUBBYTES[3].a/U5500  ( .A(n9485), .B(n8520), .Z(n9484) );
  XOR \SUBBYTES[3].a/U5499  ( .A(\SUBBYTES[3].a/w2555 ), .B(
        \SUBBYTES[3].a/w2572 ), .Z(n8520) );
  XOR \SUBBYTES[3].a/U5497  ( .A(\SUBBYTES[3].a/w2554 ), .B(
        \SUBBYTES[3].a/w2569 ), .Z(n8521) );
  XOR \SUBBYTES[3].a/U5496  ( .A(n9485), .B(n8522), .Z(n9660) );
  XOR \SUBBYTES[3].a/U5495  ( .A(\SUBBYTES[3].a/w2569 ), .B(
        \SUBBYTES[3].a/w2570 ), .Z(n8522) );
  XOR \SUBBYTES[3].a/U5494  ( .A(\SUBBYTES[3].a/w2531 ), .B(n8523), .Z(n9487)
         );
  XOR \SUBBYTES[3].a/U5493  ( .A(\SUBBYTES[3].a/w2522 ), .B(
        \SUBBYTES[3].a/w2523 ), .Z(n8523) );
  XOR \SUBBYTES[3].a/U5491  ( .A(\SUBBYTES[3].a/w2533 ), .B(n9660), .Z(n8524)
         );
  XOR \SUBBYTES[3].a/U5490  ( .A(n8526), .B(n8525), .Z(n9488) );
  XOR \SUBBYTES[3].a/U5489  ( .A(n8528), .B(n8527), .Z(n8525) );
  XOR \SUBBYTES[3].a/U5488  ( .A(\SUBBYTES[3].a/w2569 ), .B(
        \SUBBYTES[3].a/w2570 ), .Z(n8526) );
  XOR \SUBBYTES[3].a/U5487  ( .A(\SUBBYTES[3].a/w2533 ), .B(
        \SUBBYTES[3].a/w2557 ), .Z(n8527) );
  XOR \SUBBYTES[3].a/U5486  ( .A(\SUBBYTES[3].a/w2522 ), .B(
        \SUBBYTES[3].a/w2531 ), .Z(n8528) );
  XOR \SUBBYTES[3].a/U5485  ( .A(\SUBBYTES[3].a/w2554 ), .B(n8529), .Z(n9486)
         );
  XOR \SUBBYTES[3].a/U5484  ( .A(\SUBBYTES[3].a/w2537 ), .B(
        \SUBBYTES[3].a/w2540 ), .Z(n8529) );
  XOR \SUBBYTES[3].a/U5482  ( .A(\SUBBYTES[3].a/w2525 ), .B(n9488), .Z(n8530)
         );
  XOR \SUBBYTES[3].a/U5480  ( .A(\SUBBYTES[3].a/w2557 ), .B(
        \SUBBYTES[3].a/w2570 ), .Z(n8531) );
  XOR \SUBBYTES[3].a/U5478  ( .A(n8535), .B(n8534), .Z(n8532) );
  XOR \SUBBYTES[3].a/U5477  ( .A(n8537), .B(n8536), .Z(n8533) );
  XOR \SUBBYTES[3].a/U5476  ( .A(\SUBBYTES[3].a/w2569 ), .B(
        \SUBBYTES[3].a/w2572 ), .Z(n8534) );
  XOR \SUBBYTES[3].a/U5475  ( .A(\SUBBYTES[3].a/w2562 ), .B(
        \SUBBYTES[3].a/w2565 ), .Z(n8535) );
  XOR \SUBBYTES[3].a/U5474  ( .A(\SUBBYTES[3].a/w2537 ), .B(
        \SUBBYTES[3].a/w2538 ), .Z(n8536) );
  XOR \SUBBYTES[3].a/U5473  ( .A(\SUBBYTES[3].a/w2522 ), .B(
        \SUBBYTES[3].a/w2525 ), .Z(n8537) );
  XOR \SUBBYTES[3].a/U5471  ( .A(n9485), .B(n8540), .Z(n8538) );
  XOR \SUBBYTES[3].a/U5470  ( .A(n9487), .B(n9486), .Z(n8539) );
  XOR \SUBBYTES[3].a/U5469  ( .A(\SUBBYTES[3].a/w2530 ), .B(
        \SUBBYTES[3].a/w2557 ), .Z(n8540) );
  XOR \SUBBYTES[3].a/U5467  ( .A(n9488), .B(n8543), .Z(n8541) );
  XOR \SUBBYTES[3].a/U5466  ( .A(\SUBBYTES[3].a/w2563 ), .B(
        \SUBBYTES[3].a/w2565 ), .Z(n8542) );
  XOR \SUBBYTES[3].a/U5465  ( .A(\SUBBYTES[3].a/w2523 ), .B(
        \SUBBYTES[3].a/w2555 ), .Z(n8543) );
  XOR \SUBBYTES[3].a/U5464  ( .A(\SUBBYTES[3].a/w2355 ), .B(
        \SUBBYTES[3].a/w2356 ), .Z(n9490) );
  XOR \SUBBYTES[3].a/U5463  ( .A(n9490), .B(n8544), .Z(n9489) );
  XOR \SUBBYTES[3].a/U5462  ( .A(\SUBBYTES[3].a/w2348 ), .B(
        \SUBBYTES[3].a/w2365 ), .Z(n8544) );
  XOR \SUBBYTES[3].a/U5460  ( .A(\SUBBYTES[3].a/w2347 ), .B(
        \SUBBYTES[3].a/w2362 ), .Z(n8545) );
  XOR \SUBBYTES[3].a/U5459  ( .A(n9490), .B(n8546), .Z(n9661) );
  XOR \SUBBYTES[3].a/U5458  ( .A(\SUBBYTES[3].a/w2362 ), .B(
        \SUBBYTES[3].a/w2363 ), .Z(n8546) );
  XOR \SUBBYTES[3].a/U5457  ( .A(\SUBBYTES[3].a/w2324 ), .B(n8547), .Z(n9492)
         );
  XOR \SUBBYTES[3].a/U5456  ( .A(\SUBBYTES[3].a/w2315 ), .B(
        \SUBBYTES[3].a/w2316 ), .Z(n8547) );
  XOR \SUBBYTES[3].a/U5454  ( .A(\SUBBYTES[3].a/w2326 ), .B(n9661), .Z(n8548)
         );
  XOR \SUBBYTES[3].a/U5453  ( .A(n8550), .B(n8549), .Z(n9493) );
  XOR \SUBBYTES[3].a/U5452  ( .A(n8552), .B(n8551), .Z(n8549) );
  XOR \SUBBYTES[3].a/U5451  ( .A(\SUBBYTES[3].a/w2362 ), .B(
        \SUBBYTES[3].a/w2363 ), .Z(n8550) );
  XOR \SUBBYTES[3].a/U5450  ( .A(\SUBBYTES[3].a/w2326 ), .B(
        \SUBBYTES[3].a/w2350 ), .Z(n8551) );
  XOR \SUBBYTES[3].a/U5449  ( .A(\SUBBYTES[3].a/w2315 ), .B(
        \SUBBYTES[3].a/w2324 ), .Z(n8552) );
  XOR \SUBBYTES[3].a/U5448  ( .A(\SUBBYTES[3].a/w2347 ), .B(n8553), .Z(n9491)
         );
  XOR \SUBBYTES[3].a/U5447  ( .A(\SUBBYTES[3].a/w2330 ), .B(
        \SUBBYTES[3].a/w2333 ), .Z(n8553) );
  XOR \SUBBYTES[3].a/U5445  ( .A(\SUBBYTES[3].a/w2318 ), .B(n9493), .Z(n8554)
         );
  XOR \SUBBYTES[3].a/U5443  ( .A(\SUBBYTES[3].a/w2350 ), .B(
        \SUBBYTES[3].a/w2363 ), .Z(n8555) );
  XOR \SUBBYTES[3].a/U5441  ( .A(n8559), .B(n8558), .Z(n8556) );
  XOR \SUBBYTES[3].a/U5440  ( .A(n8561), .B(n8560), .Z(n8557) );
  XOR \SUBBYTES[3].a/U5439  ( .A(\SUBBYTES[3].a/w2362 ), .B(
        \SUBBYTES[3].a/w2365 ), .Z(n8558) );
  XOR \SUBBYTES[3].a/U5438  ( .A(\SUBBYTES[3].a/w2355 ), .B(
        \SUBBYTES[3].a/w2358 ), .Z(n8559) );
  XOR \SUBBYTES[3].a/U5437  ( .A(\SUBBYTES[3].a/w2330 ), .B(
        \SUBBYTES[3].a/w2331 ), .Z(n8560) );
  XOR \SUBBYTES[3].a/U5436  ( .A(\SUBBYTES[3].a/w2315 ), .B(
        \SUBBYTES[3].a/w2318 ), .Z(n8561) );
  XOR \SUBBYTES[3].a/U5434  ( .A(n9490), .B(n8564), .Z(n8562) );
  XOR \SUBBYTES[3].a/U5433  ( .A(n9492), .B(n9491), .Z(n8563) );
  XOR \SUBBYTES[3].a/U5432  ( .A(\SUBBYTES[3].a/w2323 ), .B(
        \SUBBYTES[3].a/w2350 ), .Z(n8564) );
  XOR \SUBBYTES[3].a/U5430  ( .A(n9493), .B(n8567), .Z(n8565) );
  XOR \SUBBYTES[3].a/U5429  ( .A(\SUBBYTES[3].a/w2356 ), .B(
        \SUBBYTES[3].a/w2358 ), .Z(n8566) );
  XOR \SUBBYTES[3].a/U5428  ( .A(\SUBBYTES[3].a/w2316 ), .B(
        \SUBBYTES[3].a/w2348 ), .Z(n8567) );
  XOR \SUBBYTES[3].a/U5427  ( .A(\SUBBYTES[3].a/w2148 ), .B(
        \SUBBYTES[3].a/w2149 ), .Z(n9495) );
  XOR \SUBBYTES[3].a/U5426  ( .A(n9495), .B(n8568), .Z(n9494) );
  XOR \SUBBYTES[3].a/U5425  ( .A(\SUBBYTES[3].a/w2141 ), .B(
        \SUBBYTES[3].a/w2158 ), .Z(n8568) );
  XOR \SUBBYTES[3].a/U5423  ( .A(\SUBBYTES[3].a/w2140 ), .B(
        \SUBBYTES[3].a/w2155 ), .Z(n8569) );
  XOR \SUBBYTES[3].a/U5422  ( .A(n9495), .B(n8570), .Z(n9662) );
  XOR \SUBBYTES[3].a/U5421  ( .A(\SUBBYTES[3].a/w2155 ), .B(
        \SUBBYTES[3].a/w2156 ), .Z(n8570) );
  XOR \SUBBYTES[3].a/U5420  ( .A(\SUBBYTES[3].a/w2117 ), .B(n8571), .Z(n9497)
         );
  XOR \SUBBYTES[3].a/U5419  ( .A(\SUBBYTES[3].a/w2108 ), .B(
        \SUBBYTES[3].a/w2109 ), .Z(n8571) );
  XOR \SUBBYTES[3].a/U5417  ( .A(\SUBBYTES[3].a/w2119 ), .B(n9662), .Z(n8572)
         );
  XOR \SUBBYTES[3].a/U5416  ( .A(n8574), .B(n8573), .Z(n9498) );
  XOR \SUBBYTES[3].a/U5415  ( .A(n8576), .B(n8575), .Z(n8573) );
  XOR \SUBBYTES[3].a/U5414  ( .A(\SUBBYTES[3].a/w2155 ), .B(
        \SUBBYTES[3].a/w2156 ), .Z(n8574) );
  XOR \SUBBYTES[3].a/U5413  ( .A(\SUBBYTES[3].a/w2119 ), .B(
        \SUBBYTES[3].a/w2143 ), .Z(n8575) );
  XOR \SUBBYTES[3].a/U5412  ( .A(\SUBBYTES[3].a/w2108 ), .B(
        \SUBBYTES[3].a/w2117 ), .Z(n8576) );
  XOR \SUBBYTES[3].a/U5411  ( .A(\SUBBYTES[3].a/w2140 ), .B(n8577), .Z(n9496)
         );
  XOR \SUBBYTES[3].a/U5410  ( .A(\SUBBYTES[3].a/w2123 ), .B(
        \SUBBYTES[3].a/w2126 ), .Z(n8577) );
  XOR \SUBBYTES[3].a/U5408  ( .A(\SUBBYTES[3].a/w2111 ), .B(n9498), .Z(n8578)
         );
  XOR \SUBBYTES[3].a/U5406  ( .A(\SUBBYTES[3].a/w2143 ), .B(
        \SUBBYTES[3].a/w2156 ), .Z(n8579) );
  XOR \SUBBYTES[3].a/U5404  ( .A(n8583), .B(n8582), .Z(n8580) );
  XOR \SUBBYTES[3].a/U5403  ( .A(n8585), .B(n8584), .Z(n8581) );
  XOR \SUBBYTES[3].a/U5402  ( .A(\SUBBYTES[3].a/w2155 ), .B(
        \SUBBYTES[3].a/w2158 ), .Z(n8582) );
  XOR \SUBBYTES[3].a/U5401  ( .A(\SUBBYTES[3].a/w2148 ), .B(
        \SUBBYTES[3].a/w2151 ), .Z(n8583) );
  XOR \SUBBYTES[3].a/U5400  ( .A(\SUBBYTES[3].a/w2123 ), .B(
        \SUBBYTES[3].a/w2124 ), .Z(n8584) );
  XOR \SUBBYTES[3].a/U5399  ( .A(\SUBBYTES[3].a/w2108 ), .B(
        \SUBBYTES[3].a/w2111 ), .Z(n8585) );
  XOR \SUBBYTES[3].a/U5397  ( .A(n9495), .B(n8588), .Z(n8586) );
  XOR \SUBBYTES[3].a/U5396  ( .A(n9497), .B(n9496), .Z(n8587) );
  XOR \SUBBYTES[3].a/U5395  ( .A(\SUBBYTES[3].a/w2116 ), .B(
        \SUBBYTES[3].a/w2143 ), .Z(n8588) );
  XOR \SUBBYTES[3].a/U5393  ( .A(n9498), .B(n8591), .Z(n8589) );
  XOR \SUBBYTES[3].a/U5392  ( .A(\SUBBYTES[3].a/w2149 ), .B(
        \SUBBYTES[3].a/w2151 ), .Z(n8590) );
  XOR \SUBBYTES[3].a/U5391  ( .A(\SUBBYTES[3].a/w2109 ), .B(
        \SUBBYTES[3].a/w2141 ), .Z(n8591) );
  XOR \SUBBYTES[3].a/U5390  ( .A(\SUBBYTES[3].a/w1941 ), .B(
        \SUBBYTES[3].a/w1942 ), .Z(n9500) );
  XOR \SUBBYTES[3].a/U5389  ( .A(n9500), .B(n8592), .Z(n9499) );
  XOR \SUBBYTES[3].a/U5388  ( .A(\SUBBYTES[3].a/w1934 ), .B(
        \SUBBYTES[3].a/w1951 ), .Z(n8592) );
  XOR \SUBBYTES[3].a/U5386  ( .A(\SUBBYTES[3].a/w1933 ), .B(
        \SUBBYTES[3].a/w1948 ), .Z(n8593) );
  XOR \SUBBYTES[3].a/U5385  ( .A(n9500), .B(n8594), .Z(n9663) );
  XOR \SUBBYTES[3].a/U5384  ( .A(\SUBBYTES[3].a/w1948 ), .B(
        \SUBBYTES[3].a/w1949 ), .Z(n8594) );
  XOR \SUBBYTES[3].a/U5383  ( .A(\SUBBYTES[3].a/w1910 ), .B(n8595), .Z(n9502)
         );
  XOR \SUBBYTES[3].a/U5382  ( .A(\SUBBYTES[3].a/w1901 ), .B(
        \SUBBYTES[3].a/w1902 ), .Z(n8595) );
  XOR \SUBBYTES[3].a/U5380  ( .A(\SUBBYTES[3].a/w1912 ), .B(n9663), .Z(n8596)
         );
  XOR \SUBBYTES[3].a/U5379  ( .A(n8598), .B(n8597), .Z(n9503) );
  XOR \SUBBYTES[3].a/U5378  ( .A(n8600), .B(n8599), .Z(n8597) );
  XOR \SUBBYTES[3].a/U5377  ( .A(\SUBBYTES[3].a/w1948 ), .B(
        \SUBBYTES[3].a/w1949 ), .Z(n8598) );
  XOR \SUBBYTES[3].a/U5376  ( .A(\SUBBYTES[3].a/w1912 ), .B(
        \SUBBYTES[3].a/w1936 ), .Z(n8599) );
  XOR \SUBBYTES[3].a/U5375  ( .A(\SUBBYTES[3].a/w1901 ), .B(
        \SUBBYTES[3].a/w1910 ), .Z(n8600) );
  XOR \SUBBYTES[3].a/U5374  ( .A(\SUBBYTES[3].a/w1933 ), .B(n8601), .Z(n9501)
         );
  XOR \SUBBYTES[3].a/U5373  ( .A(\SUBBYTES[3].a/w1916 ), .B(
        \SUBBYTES[3].a/w1919 ), .Z(n8601) );
  XOR \SUBBYTES[3].a/U5371  ( .A(\SUBBYTES[3].a/w1904 ), .B(n9503), .Z(n8602)
         );
  XOR \SUBBYTES[3].a/U5369  ( .A(\SUBBYTES[3].a/w1936 ), .B(
        \SUBBYTES[3].a/w1949 ), .Z(n8603) );
  XOR \SUBBYTES[3].a/U5367  ( .A(n8607), .B(n8606), .Z(n8604) );
  XOR \SUBBYTES[3].a/U5366  ( .A(n8609), .B(n8608), .Z(n8605) );
  XOR \SUBBYTES[3].a/U5365  ( .A(\SUBBYTES[3].a/w1948 ), .B(
        \SUBBYTES[3].a/w1951 ), .Z(n8606) );
  XOR \SUBBYTES[3].a/U5364  ( .A(\SUBBYTES[3].a/w1941 ), .B(
        \SUBBYTES[3].a/w1944 ), .Z(n8607) );
  XOR \SUBBYTES[3].a/U5363  ( .A(\SUBBYTES[3].a/w1916 ), .B(
        \SUBBYTES[3].a/w1917 ), .Z(n8608) );
  XOR \SUBBYTES[3].a/U5362  ( .A(\SUBBYTES[3].a/w1901 ), .B(
        \SUBBYTES[3].a/w1904 ), .Z(n8609) );
  XOR \SUBBYTES[3].a/U5360  ( .A(n9500), .B(n8612), .Z(n8610) );
  XOR \SUBBYTES[3].a/U5359  ( .A(n9502), .B(n9501), .Z(n8611) );
  XOR \SUBBYTES[3].a/U5358  ( .A(\SUBBYTES[3].a/w1909 ), .B(
        \SUBBYTES[3].a/w1936 ), .Z(n8612) );
  XOR \SUBBYTES[3].a/U5356  ( .A(n9503), .B(n8615), .Z(n8613) );
  XOR \SUBBYTES[3].a/U5355  ( .A(\SUBBYTES[3].a/w1942 ), .B(
        \SUBBYTES[3].a/w1944 ), .Z(n8614) );
  XOR \SUBBYTES[3].a/U5354  ( .A(\SUBBYTES[3].a/w1902 ), .B(
        \SUBBYTES[3].a/w1934 ), .Z(n8615) );
  XOR \SUBBYTES[3].a/U5353  ( .A(\SUBBYTES[3].a/w1734 ), .B(
        \SUBBYTES[3].a/w1735 ), .Z(n9505) );
  XOR \SUBBYTES[3].a/U5352  ( .A(n9505), .B(n8616), .Z(n9504) );
  XOR \SUBBYTES[3].a/U5351  ( .A(\SUBBYTES[3].a/w1727 ), .B(
        \SUBBYTES[3].a/w1744 ), .Z(n8616) );
  XOR \SUBBYTES[3].a/U5349  ( .A(\SUBBYTES[3].a/w1726 ), .B(
        \SUBBYTES[3].a/w1741 ), .Z(n8617) );
  XOR \SUBBYTES[3].a/U5348  ( .A(n9505), .B(n8618), .Z(n9664) );
  XOR \SUBBYTES[3].a/U5347  ( .A(\SUBBYTES[3].a/w1741 ), .B(
        \SUBBYTES[3].a/w1742 ), .Z(n8618) );
  XOR \SUBBYTES[3].a/U5346  ( .A(\SUBBYTES[3].a/w1703 ), .B(n8619), .Z(n9507)
         );
  XOR \SUBBYTES[3].a/U5345  ( .A(\SUBBYTES[3].a/w1694 ), .B(
        \SUBBYTES[3].a/w1695 ), .Z(n8619) );
  XOR \SUBBYTES[3].a/U5343  ( .A(\SUBBYTES[3].a/w1705 ), .B(n9664), .Z(n8620)
         );
  XOR \SUBBYTES[3].a/U5342  ( .A(n8622), .B(n8621), .Z(n9508) );
  XOR \SUBBYTES[3].a/U5341  ( .A(n8624), .B(n8623), .Z(n8621) );
  XOR \SUBBYTES[3].a/U5340  ( .A(\SUBBYTES[3].a/w1741 ), .B(
        \SUBBYTES[3].a/w1742 ), .Z(n8622) );
  XOR \SUBBYTES[3].a/U5339  ( .A(\SUBBYTES[3].a/w1705 ), .B(
        \SUBBYTES[3].a/w1729 ), .Z(n8623) );
  XOR \SUBBYTES[3].a/U5338  ( .A(\SUBBYTES[3].a/w1694 ), .B(
        \SUBBYTES[3].a/w1703 ), .Z(n8624) );
  XOR \SUBBYTES[3].a/U5337  ( .A(\SUBBYTES[3].a/w1726 ), .B(n8625), .Z(n9506)
         );
  XOR \SUBBYTES[3].a/U5336  ( .A(\SUBBYTES[3].a/w1709 ), .B(
        \SUBBYTES[3].a/w1712 ), .Z(n8625) );
  XOR \SUBBYTES[3].a/U5334  ( .A(\SUBBYTES[3].a/w1697 ), .B(n9508), .Z(n8626)
         );
  XOR \SUBBYTES[3].a/U5332  ( .A(\SUBBYTES[3].a/w1729 ), .B(
        \SUBBYTES[3].a/w1742 ), .Z(n8627) );
  XOR \SUBBYTES[3].a/U5330  ( .A(n8631), .B(n8630), .Z(n8628) );
  XOR \SUBBYTES[3].a/U5329  ( .A(n8633), .B(n8632), .Z(n8629) );
  XOR \SUBBYTES[3].a/U5328  ( .A(\SUBBYTES[3].a/w1741 ), .B(
        \SUBBYTES[3].a/w1744 ), .Z(n8630) );
  XOR \SUBBYTES[3].a/U5327  ( .A(\SUBBYTES[3].a/w1734 ), .B(
        \SUBBYTES[3].a/w1737 ), .Z(n8631) );
  XOR \SUBBYTES[3].a/U5326  ( .A(\SUBBYTES[3].a/w1709 ), .B(
        \SUBBYTES[3].a/w1710 ), .Z(n8632) );
  XOR \SUBBYTES[3].a/U5325  ( .A(\SUBBYTES[3].a/w1694 ), .B(
        \SUBBYTES[3].a/w1697 ), .Z(n8633) );
  XOR \SUBBYTES[3].a/U5323  ( .A(n9505), .B(n8636), .Z(n8634) );
  XOR \SUBBYTES[3].a/U5322  ( .A(n9507), .B(n9506), .Z(n8635) );
  XOR \SUBBYTES[3].a/U5321  ( .A(\SUBBYTES[3].a/w1702 ), .B(
        \SUBBYTES[3].a/w1729 ), .Z(n8636) );
  XOR \SUBBYTES[3].a/U5319  ( .A(n9508), .B(n8639), .Z(n8637) );
  XOR \SUBBYTES[3].a/U5318  ( .A(\SUBBYTES[3].a/w1735 ), .B(
        \SUBBYTES[3].a/w1737 ), .Z(n8638) );
  XOR \SUBBYTES[3].a/U5317  ( .A(\SUBBYTES[3].a/w1695 ), .B(
        \SUBBYTES[3].a/w1727 ), .Z(n8639) );
  XOR \SUBBYTES[3].a/U5316  ( .A(\SUBBYTES[3].a/w1527 ), .B(
        \SUBBYTES[3].a/w1528 ), .Z(n9510) );
  XOR \SUBBYTES[3].a/U5315  ( .A(n9510), .B(n8640), .Z(n9509) );
  XOR \SUBBYTES[3].a/U5314  ( .A(\SUBBYTES[3].a/w1520 ), .B(
        \SUBBYTES[3].a/w1537 ), .Z(n8640) );
  XOR \SUBBYTES[3].a/U5312  ( .A(\SUBBYTES[3].a/w1519 ), .B(
        \SUBBYTES[3].a/w1534 ), .Z(n8641) );
  XOR \SUBBYTES[3].a/U5311  ( .A(n9510), .B(n8642), .Z(n9665) );
  XOR \SUBBYTES[3].a/U5310  ( .A(\SUBBYTES[3].a/w1534 ), .B(
        \SUBBYTES[3].a/w1535 ), .Z(n8642) );
  XOR \SUBBYTES[3].a/U5309  ( .A(\SUBBYTES[3].a/w1496 ), .B(n8643), .Z(n9512)
         );
  XOR \SUBBYTES[3].a/U5308  ( .A(\SUBBYTES[3].a/w1487 ), .B(
        \SUBBYTES[3].a/w1488 ), .Z(n8643) );
  XOR \SUBBYTES[3].a/U5306  ( .A(\SUBBYTES[3].a/w1498 ), .B(n9665), .Z(n8644)
         );
  XOR \SUBBYTES[3].a/U5305  ( .A(n8646), .B(n8645), .Z(n9513) );
  XOR \SUBBYTES[3].a/U5304  ( .A(n8648), .B(n8647), .Z(n8645) );
  XOR \SUBBYTES[3].a/U5303  ( .A(\SUBBYTES[3].a/w1534 ), .B(
        \SUBBYTES[3].a/w1535 ), .Z(n8646) );
  XOR \SUBBYTES[3].a/U5302  ( .A(\SUBBYTES[3].a/w1498 ), .B(
        \SUBBYTES[3].a/w1522 ), .Z(n8647) );
  XOR \SUBBYTES[3].a/U5301  ( .A(\SUBBYTES[3].a/w1487 ), .B(
        \SUBBYTES[3].a/w1496 ), .Z(n8648) );
  XOR \SUBBYTES[3].a/U5300  ( .A(\SUBBYTES[3].a/w1519 ), .B(n8649), .Z(n9511)
         );
  XOR \SUBBYTES[3].a/U5299  ( .A(\SUBBYTES[3].a/w1502 ), .B(
        \SUBBYTES[3].a/w1505 ), .Z(n8649) );
  XOR \SUBBYTES[3].a/U5297  ( .A(\SUBBYTES[3].a/w1490 ), .B(n9513), .Z(n8650)
         );
  XOR \SUBBYTES[3].a/U5295  ( .A(\SUBBYTES[3].a/w1522 ), .B(
        \SUBBYTES[3].a/w1535 ), .Z(n8651) );
  XOR \SUBBYTES[3].a/U5293  ( .A(n8655), .B(n8654), .Z(n8652) );
  XOR \SUBBYTES[3].a/U5292  ( .A(n8657), .B(n8656), .Z(n8653) );
  XOR \SUBBYTES[3].a/U5291  ( .A(\SUBBYTES[3].a/w1534 ), .B(
        \SUBBYTES[3].a/w1537 ), .Z(n8654) );
  XOR \SUBBYTES[3].a/U5290  ( .A(\SUBBYTES[3].a/w1527 ), .B(
        \SUBBYTES[3].a/w1530 ), .Z(n8655) );
  XOR \SUBBYTES[3].a/U5289  ( .A(\SUBBYTES[3].a/w1502 ), .B(
        \SUBBYTES[3].a/w1503 ), .Z(n8656) );
  XOR \SUBBYTES[3].a/U5288  ( .A(\SUBBYTES[3].a/w1487 ), .B(
        \SUBBYTES[3].a/w1490 ), .Z(n8657) );
  XOR \SUBBYTES[3].a/U5286  ( .A(n9510), .B(n8660), .Z(n8658) );
  XOR \SUBBYTES[3].a/U5285  ( .A(n9512), .B(n9511), .Z(n8659) );
  XOR \SUBBYTES[3].a/U5284  ( .A(\SUBBYTES[3].a/w1495 ), .B(
        \SUBBYTES[3].a/w1522 ), .Z(n8660) );
  XOR \SUBBYTES[3].a/U5282  ( .A(n9513), .B(n8663), .Z(n8661) );
  XOR \SUBBYTES[3].a/U5281  ( .A(\SUBBYTES[3].a/w1528 ), .B(
        \SUBBYTES[3].a/w1530 ), .Z(n8662) );
  XOR \SUBBYTES[3].a/U5280  ( .A(\SUBBYTES[3].a/w1488 ), .B(
        \SUBBYTES[3].a/w1520 ), .Z(n8663) );
  XOR \SUBBYTES[3].a/U5279  ( .A(\SUBBYTES[3].a/w1320 ), .B(
        \SUBBYTES[3].a/w1321 ), .Z(n9515) );
  XOR \SUBBYTES[3].a/U5278  ( .A(n9515), .B(n8664), .Z(n9514) );
  XOR \SUBBYTES[3].a/U5277  ( .A(\SUBBYTES[3].a/w1313 ), .B(
        \SUBBYTES[3].a/w1330 ), .Z(n8664) );
  XOR \SUBBYTES[3].a/U5275  ( .A(\SUBBYTES[3].a/w1312 ), .B(
        \SUBBYTES[3].a/w1327 ), .Z(n8665) );
  XOR \SUBBYTES[3].a/U5274  ( .A(n9515), .B(n8666), .Z(n9666) );
  XOR \SUBBYTES[3].a/U5273  ( .A(\SUBBYTES[3].a/w1327 ), .B(
        \SUBBYTES[3].a/w1328 ), .Z(n8666) );
  XOR \SUBBYTES[3].a/U5272  ( .A(\SUBBYTES[3].a/w1289 ), .B(n8667), .Z(n9517)
         );
  XOR \SUBBYTES[3].a/U5271  ( .A(\SUBBYTES[3].a/w1280 ), .B(
        \SUBBYTES[3].a/w1281 ), .Z(n8667) );
  XOR \SUBBYTES[3].a/U5269  ( .A(\SUBBYTES[3].a/w1291 ), .B(n9666), .Z(n8668)
         );
  XOR \SUBBYTES[3].a/U5268  ( .A(n8670), .B(n8669), .Z(n9518) );
  XOR \SUBBYTES[3].a/U5267  ( .A(n8672), .B(n8671), .Z(n8669) );
  XOR \SUBBYTES[3].a/U5266  ( .A(\SUBBYTES[3].a/w1327 ), .B(
        \SUBBYTES[3].a/w1328 ), .Z(n8670) );
  XOR \SUBBYTES[3].a/U5265  ( .A(\SUBBYTES[3].a/w1291 ), .B(
        \SUBBYTES[3].a/w1315 ), .Z(n8671) );
  XOR \SUBBYTES[3].a/U5264  ( .A(\SUBBYTES[3].a/w1280 ), .B(
        \SUBBYTES[3].a/w1289 ), .Z(n8672) );
  XOR \SUBBYTES[3].a/U5263  ( .A(\SUBBYTES[3].a/w1312 ), .B(n8673), .Z(n9516)
         );
  XOR \SUBBYTES[3].a/U5262  ( .A(\SUBBYTES[3].a/w1295 ), .B(
        \SUBBYTES[3].a/w1298 ), .Z(n8673) );
  XOR \SUBBYTES[3].a/U5260  ( .A(\SUBBYTES[3].a/w1283 ), .B(n9518), .Z(n8674)
         );
  XOR \SUBBYTES[3].a/U5258  ( .A(\SUBBYTES[3].a/w1315 ), .B(
        \SUBBYTES[3].a/w1328 ), .Z(n8675) );
  XOR \SUBBYTES[3].a/U5256  ( .A(n8679), .B(n8678), .Z(n8676) );
  XOR \SUBBYTES[3].a/U5255  ( .A(n8681), .B(n8680), .Z(n8677) );
  XOR \SUBBYTES[3].a/U5254  ( .A(\SUBBYTES[3].a/w1327 ), .B(
        \SUBBYTES[3].a/w1330 ), .Z(n8678) );
  XOR \SUBBYTES[3].a/U5253  ( .A(\SUBBYTES[3].a/w1320 ), .B(
        \SUBBYTES[3].a/w1323 ), .Z(n8679) );
  XOR \SUBBYTES[3].a/U5252  ( .A(\SUBBYTES[3].a/w1295 ), .B(
        \SUBBYTES[3].a/w1296 ), .Z(n8680) );
  XOR \SUBBYTES[3].a/U5251  ( .A(\SUBBYTES[3].a/w1280 ), .B(
        \SUBBYTES[3].a/w1283 ), .Z(n8681) );
  XOR \SUBBYTES[3].a/U5249  ( .A(n9515), .B(n8684), .Z(n8682) );
  XOR \SUBBYTES[3].a/U5248  ( .A(n9517), .B(n9516), .Z(n8683) );
  XOR \SUBBYTES[3].a/U5247  ( .A(\SUBBYTES[3].a/w1288 ), .B(
        \SUBBYTES[3].a/w1315 ), .Z(n8684) );
  XOR \SUBBYTES[3].a/U5245  ( .A(n9518), .B(n8687), .Z(n8685) );
  XOR \SUBBYTES[3].a/U5244  ( .A(\SUBBYTES[3].a/w1321 ), .B(
        \SUBBYTES[3].a/w1323 ), .Z(n8686) );
  XOR \SUBBYTES[3].a/U5243  ( .A(\SUBBYTES[3].a/w1281 ), .B(
        \SUBBYTES[3].a/w1313 ), .Z(n8687) );
  XOR \SUBBYTES[3].a/U5242  ( .A(\SUBBYTES[3].a/w1113 ), .B(
        \SUBBYTES[3].a/w1114 ), .Z(n9520) );
  XOR \SUBBYTES[3].a/U5241  ( .A(n9520), .B(n8688), .Z(n9519) );
  XOR \SUBBYTES[3].a/U5240  ( .A(\SUBBYTES[3].a/w1106 ), .B(
        \SUBBYTES[3].a/w1123 ), .Z(n8688) );
  XOR \SUBBYTES[3].a/U5238  ( .A(\SUBBYTES[3].a/w1105 ), .B(
        \SUBBYTES[3].a/w1120 ), .Z(n8689) );
  XOR \SUBBYTES[3].a/U5237  ( .A(n9520), .B(n8690), .Z(n9667) );
  XOR \SUBBYTES[3].a/U5236  ( .A(\SUBBYTES[3].a/w1120 ), .B(
        \SUBBYTES[3].a/w1121 ), .Z(n8690) );
  XOR \SUBBYTES[3].a/U5235  ( .A(\SUBBYTES[3].a/w1082 ), .B(n8691), .Z(n9522)
         );
  XOR \SUBBYTES[3].a/U5234  ( .A(\SUBBYTES[3].a/w1073 ), .B(
        \SUBBYTES[3].a/w1074 ), .Z(n8691) );
  XOR \SUBBYTES[3].a/U5232  ( .A(\SUBBYTES[3].a/w1084 ), .B(n9667), .Z(n8692)
         );
  XOR \SUBBYTES[3].a/U5231  ( .A(n8694), .B(n8693), .Z(n9523) );
  XOR \SUBBYTES[3].a/U5230  ( .A(n8696), .B(n8695), .Z(n8693) );
  XOR \SUBBYTES[3].a/U5229  ( .A(\SUBBYTES[3].a/w1120 ), .B(
        \SUBBYTES[3].a/w1121 ), .Z(n8694) );
  XOR \SUBBYTES[3].a/U5228  ( .A(\SUBBYTES[3].a/w1084 ), .B(
        \SUBBYTES[3].a/w1108 ), .Z(n8695) );
  XOR \SUBBYTES[3].a/U5227  ( .A(\SUBBYTES[3].a/w1073 ), .B(
        \SUBBYTES[3].a/w1082 ), .Z(n8696) );
  XOR \SUBBYTES[3].a/U5226  ( .A(\SUBBYTES[3].a/w1105 ), .B(n8697), .Z(n9521)
         );
  XOR \SUBBYTES[3].a/U5225  ( .A(\SUBBYTES[3].a/w1088 ), .B(
        \SUBBYTES[3].a/w1091 ), .Z(n8697) );
  XOR \SUBBYTES[3].a/U5223  ( .A(\SUBBYTES[3].a/w1076 ), .B(n9523), .Z(n8698)
         );
  XOR \SUBBYTES[3].a/U5221  ( .A(\SUBBYTES[3].a/w1108 ), .B(
        \SUBBYTES[3].a/w1121 ), .Z(n8699) );
  XOR \SUBBYTES[3].a/U5219  ( .A(n8703), .B(n8702), .Z(n8700) );
  XOR \SUBBYTES[3].a/U5218  ( .A(n8705), .B(n8704), .Z(n8701) );
  XOR \SUBBYTES[3].a/U5217  ( .A(\SUBBYTES[3].a/w1120 ), .B(
        \SUBBYTES[3].a/w1123 ), .Z(n8702) );
  XOR \SUBBYTES[3].a/U5216  ( .A(\SUBBYTES[3].a/w1113 ), .B(
        \SUBBYTES[3].a/w1116 ), .Z(n8703) );
  XOR \SUBBYTES[3].a/U5215  ( .A(\SUBBYTES[3].a/w1088 ), .B(
        \SUBBYTES[3].a/w1089 ), .Z(n8704) );
  XOR \SUBBYTES[3].a/U5214  ( .A(\SUBBYTES[3].a/w1073 ), .B(
        \SUBBYTES[3].a/w1076 ), .Z(n8705) );
  XOR \SUBBYTES[3].a/U5212  ( .A(n9520), .B(n8708), .Z(n8706) );
  XOR \SUBBYTES[3].a/U5211  ( .A(n9522), .B(n9521), .Z(n8707) );
  XOR \SUBBYTES[3].a/U5210  ( .A(\SUBBYTES[3].a/w1081 ), .B(
        \SUBBYTES[3].a/w1108 ), .Z(n8708) );
  XOR \SUBBYTES[3].a/U5208  ( .A(n9523), .B(n8711), .Z(n8709) );
  XOR \SUBBYTES[3].a/U5207  ( .A(\SUBBYTES[3].a/w1114 ), .B(
        \SUBBYTES[3].a/w1116 ), .Z(n8710) );
  XOR \SUBBYTES[3].a/U5206  ( .A(\SUBBYTES[3].a/w1074 ), .B(
        \SUBBYTES[3].a/w1106 ), .Z(n8711) );
  XOR \SUBBYTES[3].a/U5205  ( .A(\SUBBYTES[3].a/w906 ), .B(
        \SUBBYTES[3].a/w907 ), .Z(n9525) );
  XOR \SUBBYTES[3].a/U5204  ( .A(n9525), .B(n8712), .Z(n9524) );
  XOR \SUBBYTES[3].a/U5203  ( .A(\SUBBYTES[3].a/w899 ), .B(
        \SUBBYTES[3].a/w916 ), .Z(n8712) );
  XOR \SUBBYTES[3].a/U5201  ( .A(\SUBBYTES[3].a/w898 ), .B(
        \SUBBYTES[3].a/w913 ), .Z(n8713) );
  XOR \SUBBYTES[3].a/U5200  ( .A(n9525), .B(n8714), .Z(n9668) );
  XOR \SUBBYTES[3].a/U5199  ( .A(\SUBBYTES[3].a/w913 ), .B(
        \SUBBYTES[3].a/w914 ), .Z(n8714) );
  XOR \SUBBYTES[3].a/U5198  ( .A(\SUBBYTES[3].a/w875 ), .B(n8715), .Z(n9527)
         );
  XOR \SUBBYTES[3].a/U5197  ( .A(\SUBBYTES[3].a/w866 ), .B(
        \SUBBYTES[3].a/w867 ), .Z(n8715) );
  XOR \SUBBYTES[3].a/U5195  ( .A(\SUBBYTES[3].a/w877 ), .B(n9668), .Z(n8716)
         );
  XOR \SUBBYTES[3].a/U5194  ( .A(n8718), .B(n8717), .Z(n9528) );
  XOR \SUBBYTES[3].a/U5193  ( .A(n8720), .B(n8719), .Z(n8717) );
  XOR \SUBBYTES[3].a/U5192  ( .A(\SUBBYTES[3].a/w913 ), .B(
        \SUBBYTES[3].a/w914 ), .Z(n8718) );
  XOR \SUBBYTES[3].a/U5191  ( .A(\SUBBYTES[3].a/w877 ), .B(
        \SUBBYTES[3].a/w901 ), .Z(n8719) );
  XOR \SUBBYTES[3].a/U5190  ( .A(\SUBBYTES[3].a/w866 ), .B(
        \SUBBYTES[3].a/w875 ), .Z(n8720) );
  XOR \SUBBYTES[3].a/U5189  ( .A(\SUBBYTES[3].a/w898 ), .B(n8721), .Z(n9526)
         );
  XOR \SUBBYTES[3].a/U5188  ( .A(\SUBBYTES[3].a/w881 ), .B(
        \SUBBYTES[3].a/w884 ), .Z(n8721) );
  XOR \SUBBYTES[3].a/U5186  ( .A(\SUBBYTES[3].a/w869 ), .B(n9528), .Z(n8722)
         );
  XOR \SUBBYTES[3].a/U5184  ( .A(\SUBBYTES[3].a/w901 ), .B(
        \SUBBYTES[3].a/w914 ), .Z(n8723) );
  XOR \SUBBYTES[3].a/U5182  ( .A(n8727), .B(n8726), .Z(n8724) );
  XOR \SUBBYTES[3].a/U5181  ( .A(n8729), .B(n8728), .Z(n8725) );
  XOR \SUBBYTES[3].a/U5180  ( .A(\SUBBYTES[3].a/w913 ), .B(
        \SUBBYTES[3].a/w916 ), .Z(n8726) );
  XOR \SUBBYTES[3].a/U5179  ( .A(\SUBBYTES[3].a/w906 ), .B(
        \SUBBYTES[3].a/w909 ), .Z(n8727) );
  XOR \SUBBYTES[3].a/U5178  ( .A(\SUBBYTES[3].a/w881 ), .B(
        \SUBBYTES[3].a/w882 ), .Z(n8728) );
  XOR \SUBBYTES[3].a/U5177  ( .A(\SUBBYTES[3].a/w866 ), .B(
        \SUBBYTES[3].a/w869 ), .Z(n8729) );
  XOR \SUBBYTES[3].a/U5175  ( .A(n9525), .B(n8732), .Z(n8730) );
  XOR \SUBBYTES[3].a/U5174  ( .A(n9527), .B(n9526), .Z(n8731) );
  XOR \SUBBYTES[3].a/U5173  ( .A(\SUBBYTES[3].a/w874 ), .B(
        \SUBBYTES[3].a/w901 ), .Z(n8732) );
  XOR \SUBBYTES[3].a/U5171  ( .A(n9528), .B(n8735), .Z(n8733) );
  XOR \SUBBYTES[3].a/U5170  ( .A(\SUBBYTES[3].a/w907 ), .B(
        \SUBBYTES[3].a/w909 ), .Z(n8734) );
  XOR \SUBBYTES[3].a/U5169  ( .A(\SUBBYTES[3].a/w867 ), .B(
        \SUBBYTES[3].a/w899 ), .Z(n8735) );
  XOR \SUBBYTES[3].a/U5168  ( .A(\SUBBYTES[3].a/w699 ), .B(
        \SUBBYTES[3].a/w700 ), .Z(n9530) );
  XOR \SUBBYTES[3].a/U5167  ( .A(n9530), .B(n8736), .Z(n9529) );
  XOR \SUBBYTES[3].a/U5166  ( .A(\SUBBYTES[3].a/w692 ), .B(
        \SUBBYTES[3].a/w709 ), .Z(n8736) );
  XOR \SUBBYTES[3].a/U5164  ( .A(\SUBBYTES[3].a/w691 ), .B(
        \SUBBYTES[3].a/w706 ), .Z(n8737) );
  XOR \SUBBYTES[3].a/U5163  ( .A(n9530), .B(n8738), .Z(n9669) );
  XOR \SUBBYTES[3].a/U5162  ( .A(\SUBBYTES[3].a/w706 ), .B(
        \SUBBYTES[3].a/w707 ), .Z(n8738) );
  XOR \SUBBYTES[3].a/U5161  ( .A(\SUBBYTES[3].a/w668 ), .B(n8739), .Z(n9532)
         );
  XOR \SUBBYTES[3].a/U5160  ( .A(\SUBBYTES[3].a/w659 ), .B(
        \SUBBYTES[3].a/w660 ), .Z(n8739) );
  XOR \SUBBYTES[3].a/U5158  ( .A(\SUBBYTES[3].a/w670 ), .B(n9669), .Z(n8740)
         );
  XOR \SUBBYTES[3].a/U5157  ( .A(n8742), .B(n8741), .Z(n9533) );
  XOR \SUBBYTES[3].a/U5156  ( .A(n8744), .B(n8743), .Z(n8741) );
  XOR \SUBBYTES[3].a/U5155  ( .A(\SUBBYTES[3].a/w706 ), .B(
        \SUBBYTES[3].a/w707 ), .Z(n8742) );
  XOR \SUBBYTES[3].a/U5154  ( .A(\SUBBYTES[3].a/w670 ), .B(
        \SUBBYTES[3].a/w694 ), .Z(n8743) );
  XOR \SUBBYTES[3].a/U5153  ( .A(\SUBBYTES[3].a/w659 ), .B(
        \SUBBYTES[3].a/w668 ), .Z(n8744) );
  XOR \SUBBYTES[3].a/U5152  ( .A(\SUBBYTES[3].a/w691 ), .B(n8745), .Z(n9531)
         );
  XOR \SUBBYTES[3].a/U5151  ( .A(\SUBBYTES[3].a/w674 ), .B(
        \SUBBYTES[3].a/w677 ), .Z(n8745) );
  XOR \SUBBYTES[3].a/U5149  ( .A(\SUBBYTES[3].a/w662 ), .B(n9533), .Z(n8746)
         );
  XOR \SUBBYTES[3].a/U5147  ( .A(\SUBBYTES[3].a/w694 ), .B(
        \SUBBYTES[3].a/w707 ), .Z(n8747) );
  XOR \SUBBYTES[3].a/U5145  ( .A(n8751), .B(n8750), .Z(n8748) );
  XOR \SUBBYTES[3].a/U5144  ( .A(n8753), .B(n8752), .Z(n8749) );
  XOR \SUBBYTES[3].a/U5143  ( .A(\SUBBYTES[3].a/w706 ), .B(
        \SUBBYTES[3].a/w709 ), .Z(n8750) );
  XOR \SUBBYTES[3].a/U5142  ( .A(\SUBBYTES[3].a/w699 ), .B(
        \SUBBYTES[3].a/w702 ), .Z(n8751) );
  XOR \SUBBYTES[3].a/U5141  ( .A(\SUBBYTES[3].a/w674 ), .B(
        \SUBBYTES[3].a/w675 ), .Z(n8752) );
  XOR \SUBBYTES[3].a/U5140  ( .A(\SUBBYTES[3].a/w659 ), .B(
        \SUBBYTES[3].a/w662 ), .Z(n8753) );
  XOR \SUBBYTES[3].a/U5138  ( .A(n9530), .B(n8756), .Z(n8754) );
  XOR \SUBBYTES[3].a/U5137  ( .A(n9532), .B(n9531), .Z(n8755) );
  XOR \SUBBYTES[3].a/U5136  ( .A(\SUBBYTES[3].a/w667 ), .B(
        \SUBBYTES[3].a/w694 ), .Z(n8756) );
  XOR \SUBBYTES[3].a/U5134  ( .A(n9533), .B(n8759), .Z(n8757) );
  XOR \SUBBYTES[3].a/U5133  ( .A(\SUBBYTES[3].a/w700 ), .B(
        \SUBBYTES[3].a/w702 ), .Z(n8758) );
  XOR \SUBBYTES[3].a/U5132  ( .A(\SUBBYTES[3].a/w660 ), .B(
        \SUBBYTES[3].a/w692 ), .Z(n8759) );
  XOR \SUBBYTES[3].a/U5131  ( .A(\SUBBYTES[3].a/w492 ), .B(
        \SUBBYTES[3].a/w493 ), .Z(n9535) );
  XOR \SUBBYTES[3].a/U5130  ( .A(n9535), .B(n8760), .Z(n9534) );
  XOR \SUBBYTES[3].a/U5129  ( .A(\SUBBYTES[3].a/w485 ), .B(
        \SUBBYTES[3].a/w502 ), .Z(n8760) );
  XOR \SUBBYTES[3].a/U5127  ( .A(\SUBBYTES[3].a/w484 ), .B(
        \SUBBYTES[3].a/w499 ), .Z(n8761) );
  XOR \SUBBYTES[3].a/U5126  ( .A(n9535), .B(n8762), .Z(n9670) );
  XOR \SUBBYTES[3].a/U5125  ( .A(\SUBBYTES[3].a/w499 ), .B(
        \SUBBYTES[3].a/w500 ), .Z(n8762) );
  XOR \SUBBYTES[3].a/U5124  ( .A(\SUBBYTES[3].a/w461 ), .B(n8763), .Z(n9537)
         );
  XOR \SUBBYTES[3].a/U5123  ( .A(\SUBBYTES[3].a/w452 ), .B(
        \SUBBYTES[3].a/w453 ), .Z(n8763) );
  XOR \SUBBYTES[3].a/U5121  ( .A(\SUBBYTES[3].a/w463 ), .B(n9670), .Z(n8764)
         );
  XOR \SUBBYTES[3].a/U5120  ( .A(n8766), .B(n8765), .Z(n9538) );
  XOR \SUBBYTES[3].a/U5119  ( .A(n8768), .B(n8767), .Z(n8765) );
  XOR \SUBBYTES[3].a/U5118  ( .A(\SUBBYTES[3].a/w499 ), .B(
        \SUBBYTES[3].a/w500 ), .Z(n8766) );
  XOR \SUBBYTES[3].a/U5117  ( .A(\SUBBYTES[3].a/w463 ), .B(
        \SUBBYTES[3].a/w487 ), .Z(n8767) );
  XOR \SUBBYTES[3].a/U5116  ( .A(\SUBBYTES[3].a/w452 ), .B(
        \SUBBYTES[3].a/w461 ), .Z(n8768) );
  XOR \SUBBYTES[3].a/U5115  ( .A(\SUBBYTES[3].a/w484 ), .B(n8769), .Z(n9536)
         );
  XOR \SUBBYTES[3].a/U5114  ( .A(\SUBBYTES[3].a/w467 ), .B(
        \SUBBYTES[3].a/w470 ), .Z(n8769) );
  XOR \SUBBYTES[3].a/U5112  ( .A(\SUBBYTES[3].a/w455 ), .B(n9538), .Z(n8770)
         );
  XOR \SUBBYTES[3].a/U5110  ( .A(\SUBBYTES[3].a/w487 ), .B(
        \SUBBYTES[3].a/w500 ), .Z(n8771) );
  XOR \SUBBYTES[3].a/U5108  ( .A(n8775), .B(n8774), .Z(n8772) );
  XOR \SUBBYTES[3].a/U5107  ( .A(n8777), .B(n8776), .Z(n8773) );
  XOR \SUBBYTES[3].a/U5106  ( .A(\SUBBYTES[3].a/w499 ), .B(
        \SUBBYTES[3].a/w502 ), .Z(n8774) );
  XOR \SUBBYTES[3].a/U5105  ( .A(\SUBBYTES[3].a/w492 ), .B(
        \SUBBYTES[3].a/w495 ), .Z(n8775) );
  XOR \SUBBYTES[3].a/U5104  ( .A(\SUBBYTES[3].a/w467 ), .B(
        \SUBBYTES[3].a/w468 ), .Z(n8776) );
  XOR \SUBBYTES[3].a/U5103  ( .A(\SUBBYTES[3].a/w452 ), .B(
        \SUBBYTES[3].a/w455 ), .Z(n8777) );
  XOR \SUBBYTES[3].a/U5101  ( .A(n9535), .B(n8780), .Z(n8778) );
  XOR \SUBBYTES[3].a/U5100  ( .A(n9537), .B(n9536), .Z(n8779) );
  XOR \SUBBYTES[3].a/U5099  ( .A(\SUBBYTES[3].a/w460 ), .B(
        \SUBBYTES[3].a/w487 ), .Z(n8780) );
  XOR \SUBBYTES[3].a/U5097  ( .A(n9538), .B(n8783), .Z(n8781) );
  XOR \SUBBYTES[3].a/U5096  ( .A(\SUBBYTES[3].a/w493 ), .B(
        \SUBBYTES[3].a/w495 ), .Z(n8782) );
  XOR \SUBBYTES[3].a/U5095  ( .A(\SUBBYTES[3].a/w453 ), .B(
        \SUBBYTES[3].a/w485 ), .Z(n8783) );
  XOR \SUBBYTES[3].a/U5094  ( .A(\SUBBYTES[3].a/w285 ), .B(
        \SUBBYTES[3].a/w286 ), .Z(n9540) );
  XOR \SUBBYTES[3].a/U5093  ( .A(n9540), .B(n8784), .Z(n9539) );
  XOR \SUBBYTES[3].a/U5092  ( .A(\SUBBYTES[3].a/w278 ), .B(
        \SUBBYTES[3].a/w295 ), .Z(n8784) );
  XOR \SUBBYTES[3].a/U5090  ( .A(\SUBBYTES[3].a/w277 ), .B(
        \SUBBYTES[3].a/w292 ), .Z(n8785) );
  XOR \SUBBYTES[3].a/U5089  ( .A(n9540), .B(n8786), .Z(n9671) );
  XOR \SUBBYTES[3].a/U5088  ( .A(\SUBBYTES[3].a/w292 ), .B(
        \SUBBYTES[3].a/w293 ), .Z(n8786) );
  XOR \SUBBYTES[3].a/U5087  ( .A(\SUBBYTES[3].a/w254 ), .B(n8787), .Z(n9542)
         );
  XOR \SUBBYTES[3].a/U5086  ( .A(\SUBBYTES[3].a/w245 ), .B(
        \SUBBYTES[3].a/w246 ), .Z(n8787) );
  XOR \SUBBYTES[3].a/U5084  ( .A(\SUBBYTES[3].a/w256 ), .B(n9671), .Z(n8788)
         );
  XOR \SUBBYTES[3].a/U5083  ( .A(n8790), .B(n8789), .Z(n9543) );
  XOR \SUBBYTES[3].a/U5082  ( .A(n8792), .B(n8791), .Z(n8789) );
  XOR \SUBBYTES[3].a/U5081  ( .A(\SUBBYTES[3].a/w292 ), .B(
        \SUBBYTES[3].a/w293 ), .Z(n8790) );
  XOR \SUBBYTES[3].a/U5080  ( .A(\SUBBYTES[3].a/w256 ), .B(
        \SUBBYTES[3].a/w280 ), .Z(n8791) );
  XOR \SUBBYTES[3].a/U5079  ( .A(\SUBBYTES[3].a/w245 ), .B(
        \SUBBYTES[3].a/w254 ), .Z(n8792) );
  XOR \SUBBYTES[3].a/U5078  ( .A(\SUBBYTES[3].a/w277 ), .B(n8793), .Z(n9541)
         );
  XOR \SUBBYTES[3].a/U5077  ( .A(\SUBBYTES[3].a/w260 ), .B(
        \SUBBYTES[3].a/w263 ), .Z(n8793) );
  XOR \SUBBYTES[3].a/U5075  ( .A(\SUBBYTES[3].a/w248 ), .B(n9543), .Z(n8794)
         );
  XOR \SUBBYTES[3].a/U5073  ( .A(\SUBBYTES[3].a/w280 ), .B(
        \SUBBYTES[3].a/w293 ), .Z(n8795) );
  XOR \SUBBYTES[3].a/U5071  ( .A(n8799), .B(n8798), .Z(n8796) );
  XOR \SUBBYTES[3].a/U5070  ( .A(n8801), .B(n8800), .Z(n8797) );
  XOR \SUBBYTES[3].a/U5069  ( .A(\SUBBYTES[3].a/w292 ), .B(
        \SUBBYTES[3].a/w295 ), .Z(n8798) );
  XOR \SUBBYTES[3].a/U5068  ( .A(\SUBBYTES[3].a/w285 ), .B(
        \SUBBYTES[3].a/w288 ), .Z(n8799) );
  XOR \SUBBYTES[3].a/U5067  ( .A(\SUBBYTES[3].a/w260 ), .B(
        \SUBBYTES[3].a/w261 ), .Z(n8800) );
  XOR \SUBBYTES[3].a/U5066  ( .A(\SUBBYTES[3].a/w245 ), .B(
        \SUBBYTES[3].a/w248 ), .Z(n8801) );
  XOR \SUBBYTES[3].a/U5064  ( .A(n9540), .B(n8804), .Z(n8802) );
  XOR \SUBBYTES[3].a/U5063  ( .A(n9542), .B(n9541), .Z(n8803) );
  XOR \SUBBYTES[3].a/U5062  ( .A(\SUBBYTES[3].a/w253 ), .B(
        \SUBBYTES[3].a/w280 ), .Z(n8804) );
  XOR \SUBBYTES[3].a/U5060  ( .A(n9543), .B(n8807), .Z(n8805) );
  XOR \SUBBYTES[3].a/U5059  ( .A(\SUBBYTES[3].a/w286 ), .B(
        \SUBBYTES[3].a/w288 ), .Z(n8806) );
  XOR \SUBBYTES[3].a/U5058  ( .A(\SUBBYTES[3].a/w246 ), .B(
        \SUBBYTES[3].a/w278 ), .Z(n8807) );
  XOR \SUBBYTES[3].a/U5057  ( .A(\w1[3][1] ), .B(n8808), .Z(n9544) );
  XOR \SUBBYTES[3].a/U5056  ( .A(\w1[3][3] ), .B(\w1[3][2] ), .Z(n8808) );
  XOR \SUBBYTES[3].a/U5055  ( .A(\w1[3][6] ), .B(n9544), .Z(
        \SUBBYTES[3].a/w3378 ) );
  XOR \SUBBYTES[3].a/U5054  ( .A(\w1[3][0] ), .B(\SUBBYTES[3].a/w3378 ), .Z(
        \SUBBYTES[3].a/w3265 ) );
  XOR \SUBBYTES[3].a/U5053  ( .A(\w1[3][0] ), .B(n8809), .Z(
        \SUBBYTES[3].a/w3266 ) );
  XOR \SUBBYTES[3].a/U5052  ( .A(\w1[3][6] ), .B(\w1[3][5] ), .Z(n8809) );
  XOR \SUBBYTES[3].a/U5051  ( .A(\w1[3][5] ), .B(n9544), .Z(
        \SUBBYTES[3].a/w3396 ) );
  XOR \SUBBYTES[3].a/U5050  ( .A(n8811), .B(n8810), .Z(\SUBBYTES[3].a/w3389 )
         );
  XOR \SUBBYTES[3].a/U5049  ( .A(\w1[3][3] ), .B(\w1[3][1] ), .Z(n8810) );
  XOR \SUBBYTES[3].a/U5048  ( .A(\w1[3][7] ), .B(\w1[3][4] ), .Z(n8811) );
  XOR \SUBBYTES[3].a/U5047  ( .A(\w1[3][0] ), .B(\SUBBYTES[3].a/w3389 ), .Z(
        \SUBBYTES[3].a/w3268 ) );
  XOR \SUBBYTES[3].a/U5046  ( .A(n8813), .B(n8812), .Z(\SUBBYTES[3].a/w3376 )
         );
  XOR \SUBBYTES[3].a/U5045  ( .A(\SUBBYTES[3].a/w3337 ), .B(n1004), .Z(n8812)
         );
  XOR \SUBBYTES[3].a/U5044  ( .A(\SUBBYTES[3].a/w3330 ), .B(
        \SUBBYTES[3].a/w3333 ), .Z(n8813) );
  XOR \SUBBYTES[3].a/U5043  ( .A(n8815), .B(n8814), .Z(\SUBBYTES[3].a/w3377 )
         );
  XOR \SUBBYTES[3].a/U5042  ( .A(\SUBBYTES[3].a/w3337 ), .B(n8423), .Z(n8814)
         );
  XOR \SUBBYTES[3].a/U5041  ( .A(\SUBBYTES[3].a/w3330 ), .B(n8422), .Z(n8815)
         );
  XOR \SUBBYTES[3].a/U5040  ( .A(\SUBBYTES[3].a/w3389 ), .B(n8816), .Z(
        \SUBBYTES[3].a/w3379 ) );
  XOR \SUBBYTES[3].a/U5039  ( .A(\w1[3][6] ), .B(\w1[3][5] ), .Z(n8816) );
  XOR \SUBBYTES[3].a/U5038  ( .A(n8818), .B(n8817), .Z(\SUBBYTES[3].a/w3380 )
         );
  XOR \SUBBYTES[3].a/U5037  ( .A(n8423), .B(n1004), .Z(n8817) );
  XOR \SUBBYTES[3].a/U5036  ( .A(n8422), .B(\SUBBYTES[3].a/w3333 ), .Z(n8818)
         );
  XOR \SUBBYTES[3].a/U5035  ( .A(\w1[3][7] ), .B(\w1[3][2] ), .Z(n9550) );
  XOR \SUBBYTES[3].a/U5034  ( .A(n9550), .B(n8819), .Z(\SUBBYTES[3].a/w3381 )
         );
  XOR \SUBBYTES[3].a/U5033  ( .A(\w1[3][5] ), .B(\w1[3][4] ), .Z(n8819) );
  XOR \SUBBYTES[3].a/U5032  ( .A(\w1[3][7] ), .B(\SUBBYTES[3].a/w3266 ), .Z(
        \SUBBYTES[3].a/w3269 ) );
  XOR \SUBBYTES[3].a/U5031  ( .A(\w1[3][1] ), .B(\SUBBYTES[3].a/w3266 ), .Z(
        \SUBBYTES[3].a/w3270 ) );
  XOR \SUBBYTES[3].a/U5030  ( .A(\w1[3][4] ), .B(\SUBBYTES[3].a/w3266 ), .Z(
        \SUBBYTES[3].a/w3271 ) );
  XOR \SUBBYTES[3].a/U5029  ( .A(\SUBBYTES[3].a/w3270 ), .B(n9550), .Z(
        \SUBBYTES[3].a/w3272 ) );
  XOR \SUBBYTES[3].a/U5028  ( .A(n9550), .B(n8820), .Z(\SUBBYTES[3].a/w3357 )
         );
  XOR \SUBBYTES[3].a/U5027  ( .A(\w1[3][4] ), .B(\w1[3][1] ), .Z(n8820) );
  XOR \SUBBYTES[3].a/U5026  ( .A(n8822), .B(n8821), .Z(n9547) );
  XOR \SUBBYTES[3].a/U5025  ( .A(\w1[3][4] ), .B(n8823), .Z(n8821) );
  XOR \SUBBYTES[3].a/U5024  ( .A(\SUBBYTES[3].a/w3322 ), .B(\w1[3][6] ), .Z(
        n8822) );
  XOR \SUBBYTES[3].a/U5023  ( .A(\SUBBYTES[3].a/w3296 ), .B(
        \SUBBYTES[3].a/w3303 ), .Z(n8823) );
  XOR \SUBBYTES[3].a/U5022  ( .A(n8825), .B(n8824), .Z(n9545) );
  XOR \SUBBYTES[3].a/U5021  ( .A(\w1[3][1] ), .B(n8826), .Z(n8824) );
  XOR \SUBBYTES[3].a/U5020  ( .A(\SUBBYTES[3].a/w3321 ), .B(\w1[3][5] ), .Z(
        n8825) );
  XOR \SUBBYTES[3].a/U5019  ( .A(\SUBBYTES[3].a/w3297 ), .B(
        \SUBBYTES[3].a/w3304 ), .Z(n8826) );
  XOR \SUBBYTES[3].a/U5018  ( .A(n9547), .B(n9545), .Z(\SUBBYTES[3].a/w3327 )
         );
  XOR \SUBBYTES[3].a/U5017  ( .A(\w1[3][5] ), .B(n8827), .Z(n9548) );
  XOR \SUBBYTES[3].a/U5016  ( .A(\SUBBYTES[3].a/w3289 ), .B(
        \SUBBYTES[3].a/w3299 ), .Z(n8827) );
  XOR \SUBBYTES[3].a/U5015  ( .A(n8829), .B(n8828), .Z(\SUBBYTES[3].a/w3314 )
         );
  XOR \SUBBYTES[3].a/U5014  ( .A(n9548), .B(n8830), .Z(n8828) );
  XOR \SUBBYTES[3].a/U5013  ( .A(\w1[3][4] ), .B(\SUBBYTES[3].a/w3378 ), .Z(
        n8829) );
  XOR \SUBBYTES[3].a/U5012  ( .A(\SUBBYTES[3].a/w3291 ), .B(
        \SUBBYTES[3].a/w3296 ), .Z(n8830) );
  XOR \SUBBYTES[3].a/U5011  ( .A(n8832), .B(n8831), .Z(n9546) );
  XOR \SUBBYTES[3].a/U5010  ( .A(\SUBBYTES[3].a/w3324 ), .B(\w1[3][7] ), .Z(
        n8831) );
  XOR \SUBBYTES[3].a/U5009  ( .A(\SUBBYTES[3].a/w3299 ), .B(
        \SUBBYTES[3].a/w3306 ), .Z(n8832) );
  XOR \SUBBYTES[3].a/U5008  ( .A(n9545), .B(n9546), .Z(\SUBBYTES[3].a/w3326 )
         );
  XOR \SUBBYTES[3].a/U5007  ( .A(\w1[3][3] ), .B(n8833), .Z(n9549) );
  XOR \SUBBYTES[3].a/U5006  ( .A(\SUBBYTES[3].a/w3288 ), .B(
        \SUBBYTES[3].a/w3291 ), .Z(n8833) );
  XOR \SUBBYTES[3].a/U5005  ( .A(n8835), .B(n8834), .Z(\SUBBYTES[3].a/w3315 )
         );
  XOR \SUBBYTES[3].a/U5004  ( .A(n9549), .B(n8836), .Z(n8834) );
  XOR \SUBBYTES[3].a/U5003  ( .A(\w1[3][6] ), .B(\SUBBYTES[3].a/w3357 ), .Z(
        n8835) );
  XOR \SUBBYTES[3].a/U5002  ( .A(\SUBBYTES[3].a/w3296 ), .B(
        \SUBBYTES[3].a/w3297 ), .Z(n8836) );
  XOR \SUBBYTES[3].a/U5001  ( .A(n9547), .B(n9546), .Z(\SUBBYTES[3].a/w3335 )
         );
  XOR \SUBBYTES[3].a/U5000  ( .A(n8838), .B(n8837), .Z(\SUBBYTES[3].a/w3336 )
         );
  XOR \SUBBYTES[3].a/U4999  ( .A(\w1[3][7] ), .B(n9548), .Z(n8837) );
  XOR \SUBBYTES[3].a/U4998  ( .A(\SUBBYTES[3].a/w3288 ), .B(
        \SUBBYTES[3].a/w3297 ), .Z(n8838) );
  XOR \SUBBYTES[3].a/U4997  ( .A(n8840), .B(n8839), .Z(\SUBBYTES[3].a/w3312 )
         );
  XOR \SUBBYTES[3].a/U4996  ( .A(n8842), .B(n8841), .Z(n8839) );
  XOR \SUBBYTES[3].a/U4995  ( .A(\w1[3][7] ), .B(\SUBBYTES[3].a/w3396 ), .Z(
        n8840) );
  XOR \SUBBYTES[3].a/U4994  ( .A(\SUBBYTES[3].a/w3303 ), .B(
        \SUBBYTES[3].a/w3306 ), .Z(n8841) );
  XOR \SUBBYTES[3].a/U4993  ( .A(\SUBBYTES[3].a/w3289 ), .B(
        \SUBBYTES[3].a/w3291 ), .Z(n8842) );
  XOR \SUBBYTES[3].a/U4992  ( .A(n8844), .B(n8843), .Z(\SUBBYTES[3].a/w3313 )
         );
  XOR \SUBBYTES[3].a/U4991  ( .A(n9549), .B(n8845), .Z(n8843) );
  XOR \SUBBYTES[3].a/U4990  ( .A(\w1[3][5] ), .B(n9550), .Z(n8844) );
  XOR \SUBBYTES[3].a/U4989  ( .A(\SUBBYTES[3].a/w3303 ), .B(
        \SUBBYTES[3].a/w3304 ), .Z(n8845) );
  XOR \SUBBYTES[3].a/U4988  ( .A(n8847), .B(n8846), .Z(\SUBBYTES[3].a/w3329 )
         );
  XOR \SUBBYTES[3].a/U4987  ( .A(\w1[3][1] ), .B(n8848), .Z(n8846) );
  XOR \SUBBYTES[3].a/U4986  ( .A(\SUBBYTES[3].a/w3304 ), .B(
        \SUBBYTES[3].a/w3306 ), .Z(n8847) );
  XOR \SUBBYTES[3].a/U4985  ( .A(\SUBBYTES[3].a/w3288 ), .B(
        \SUBBYTES[3].a/w3289 ), .Z(n8848) );
  XOR \SUBBYTES[3].a/U4984  ( .A(\w1[3][9] ), .B(n8849), .Z(n9551) );
  XOR \SUBBYTES[3].a/U4983  ( .A(\w1[3][11] ), .B(\w1[3][10] ), .Z(n8849) );
  XOR \SUBBYTES[3].a/U4982  ( .A(\w1[3][14] ), .B(n9551), .Z(
        \SUBBYTES[3].a/w3171 ) );
  XOR \SUBBYTES[3].a/U4981  ( .A(\w1[3][8] ), .B(\SUBBYTES[3].a/w3171 ), .Z(
        \SUBBYTES[3].a/w3058 ) );
  XOR \SUBBYTES[3].a/U4980  ( .A(\w1[3][8] ), .B(n8850), .Z(
        \SUBBYTES[3].a/w3059 ) );
  XOR \SUBBYTES[3].a/U4979  ( .A(\w1[3][14] ), .B(\w1[3][13] ), .Z(n8850) );
  XOR \SUBBYTES[3].a/U4978  ( .A(\w1[3][13] ), .B(n9551), .Z(
        \SUBBYTES[3].a/w3189 ) );
  XOR \SUBBYTES[3].a/U4977  ( .A(n8852), .B(n8851), .Z(\SUBBYTES[3].a/w3182 )
         );
  XOR \SUBBYTES[3].a/U4976  ( .A(\w1[3][11] ), .B(\w1[3][9] ), .Z(n8851) );
  XOR \SUBBYTES[3].a/U4975  ( .A(\w1[3][15] ), .B(\w1[3][12] ), .Z(n8852) );
  XOR \SUBBYTES[3].a/U4974  ( .A(\w1[3][8] ), .B(\SUBBYTES[3].a/w3182 ), .Z(
        \SUBBYTES[3].a/w3061 ) );
  XOR \SUBBYTES[3].a/U4973  ( .A(n8854), .B(n8853), .Z(\SUBBYTES[3].a/w3169 )
         );
  XOR \SUBBYTES[3].a/U4972  ( .A(\SUBBYTES[3].a/w3130 ), .B(n1003), .Z(n8853)
         );
  XOR \SUBBYTES[3].a/U4971  ( .A(\SUBBYTES[3].a/w3123 ), .B(
        \SUBBYTES[3].a/w3126 ), .Z(n8854) );
  XOR \SUBBYTES[3].a/U4970  ( .A(n8856), .B(n8855), .Z(\SUBBYTES[3].a/w3170 )
         );
  XOR \SUBBYTES[3].a/U4969  ( .A(\SUBBYTES[3].a/w3130 ), .B(n8421), .Z(n8855)
         );
  XOR \SUBBYTES[3].a/U4968  ( .A(\SUBBYTES[3].a/w3123 ), .B(n8420), .Z(n8856)
         );
  XOR \SUBBYTES[3].a/U4967  ( .A(\SUBBYTES[3].a/w3182 ), .B(n8857), .Z(
        \SUBBYTES[3].a/w3172 ) );
  XOR \SUBBYTES[3].a/U4966  ( .A(\w1[3][14] ), .B(\w1[3][13] ), .Z(n8857) );
  XOR \SUBBYTES[3].a/U4965  ( .A(n8859), .B(n8858), .Z(\SUBBYTES[3].a/w3173 )
         );
  XOR \SUBBYTES[3].a/U4964  ( .A(n8421), .B(n1003), .Z(n8858) );
  XOR \SUBBYTES[3].a/U4963  ( .A(n8420), .B(\SUBBYTES[3].a/w3126 ), .Z(n8859)
         );
  XOR \SUBBYTES[3].a/U4962  ( .A(\w1[3][15] ), .B(\w1[3][10] ), .Z(n9557) );
  XOR \SUBBYTES[3].a/U4961  ( .A(n9557), .B(n8860), .Z(\SUBBYTES[3].a/w3174 )
         );
  XOR \SUBBYTES[3].a/U4960  ( .A(\w1[3][13] ), .B(\w1[3][12] ), .Z(n8860) );
  XOR \SUBBYTES[3].a/U4959  ( .A(\w1[3][15] ), .B(\SUBBYTES[3].a/w3059 ), .Z(
        \SUBBYTES[3].a/w3062 ) );
  XOR \SUBBYTES[3].a/U4958  ( .A(\w1[3][9] ), .B(\SUBBYTES[3].a/w3059 ), .Z(
        \SUBBYTES[3].a/w3063 ) );
  XOR \SUBBYTES[3].a/U4957  ( .A(\w1[3][12] ), .B(\SUBBYTES[3].a/w3059 ), .Z(
        \SUBBYTES[3].a/w3064 ) );
  XOR \SUBBYTES[3].a/U4956  ( .A(\SUBBYTES[3].a/w3063 ), .B(n9557), .Z(
        \SUBBYTES[3].a/w3065 ) );
  XOR \SUBBYTES[3].a/U4955  ( .A(n9557), .B(n8861), .Z(\SUBBYTES[3].a/w3150 )
         );
  XOR \SUBBYTES[3].a/U4954  ( .A(\w1[3][12] ), .B(\w1[3][9] ), .Z(n8861) );
  XOR \SUBBYTES[3].a/U4953  ( .A(n8863), .B(n8862), .Z(n9554) );
  XOR \SUBBYTES[3].a/U4952  ( .A(\w1[3][12] ), .B(n8864), .Z(n8862) );
  XOR \SUBBYTES[3].a/U4951  ( .A(\SUBBYTES[3].a/w3115 ), .B(\w1[3][14] ), .Z(
        n8863) );
  XOR \SUBBYTES[3].a/U4950  ( .A(\SUBBYTES[3].a/w3089 ), .B(
        \SUBBYTES[3].a/w3096 ), .Z(n8864) );
  XOR \SUBBYTES[3].a/U4949  ( .A(n8866), .B(n8865), .Z(n9552) );
  XOR \SUBBYTES[3].a/U4948  ( .A(\w1[3][9] ), .B(n8867), .Z(n8865) );
  XOR \SUBBYTES[3].a/U4947  ( .A(\SUBBYTES[3].a/w3114 ), .B(\w1[3][13] ), .Z(
        n8866) );
  XOR \SUBBYTES[3].a/U4946  ( .A(\SUBBYTES[3].a/w3090 ), .B(
        \SUBBYTES[3].a/w3097 ), .Z(n8867) );
  XOR \SUBBYTES[3].a/U4945  ( .A(n9554), .B(n9552), .Z(\SUBBYTES[3].a/w3120 )
         );
  XOR \SUBBYTES[3].a/U4944  ( .A(\w1[3][13] ), .B(n8868), .Z(n9555) );
  XOR \SUBBYTES[3].a/U4943  ( .A(\SUBBYTES[3].a/w3082 ), .B(
        \SUBBYTES[3].a/w3092 ), .Z(n8868) );
  XOR \SUBBYTES[3].a/U4942  ( .A(n8870), .B(n8869), .Z(\SUBBYTES[3].a/w3107 )
         );
  XOR \SUBBYTES[3].a/U4941  ( .A(n9555), .B(n8871), .Z(n8869) );
  XOR \SUBBYTES[3].a/U4940  ( .A(\w1[3][12] ), .B(\SUBBYTES[3].a/w3171 ), .Z(
        n8870) );
  XOR \SUBBYTES[3].a/U4939  ( .A(\SUBBYTES[3].a/w3084 ), .B(
        \SUBBYTES[3].a/w3089 ), .Z(n8871) );
  XOR \SUBBYTES[3].a/U4938  ( .A(n8873), .B(n8872), .Z(n9553) );
  XOR \SUBBYTES[3].a/U4937  ( .A(\SUBBYTES[3].a/w3117 ), .B(\w1[3][15] ), .Z(
        n8872) );
  XOR \SUBBYTES[3].a/U4936  ( .A(\SUBBYTES[3].a/w3092 ), .B(
        \SUBBYTES[3].a/w3099 ), .Z(n8873) );
  XOR \SUBBYTES[3].a/U4935  ( .A(n9552), .B(n9553), .Z(\SUBBYTES[3].a/w3119 )
         );
  XOR \SUBBYTES[3].a/U4934  ( .A(\w1[3][11] ), .B(n8874), .Z(n9556) );
  XOR \SUBBYTES[3].a/U4933  ( .A(\SUBBYTES[3].a/w3081 ), .B(
        \SUBBYTES[3].a/w3084 ), .Z(n8874) );
  XOR \SUBBYTES[3].a/U4932  ( .A(n8876), .B(n8875), .Z(\SUBBYTES[3].a/w3108 )
         );
  XOR \SUBBYTES[3].a/U4931  ( .A(n9556), .B(n8877), .Z(n8875) );
  XOR \SUBBYTES[3].a/U4930  ( .A(\w1[3][14] ), .B(\SUBBYTES[3].a/w3150 ), .Z(
        n8876) );
  XOR \SUBBYTES[3].a/U4929  ( .A(\SUBBYTES[3].a/w3089 ), .B(
        \SUBBYTES[3].a/w3090 ), .Z(n8877) );
  XOR \SUBBYTES[3].a/U4928  ( .A(n9554), .B(n9553), .Z(\SUBBYTES[3].a/w3128 )
         );
  XOR \SUBBYTES[3].a/U4927  ( .A(n8879), .B(n8878), .Z(\SUBBYTES[3].a/w3129 )
         );
  XOR \SUBBYTES[3].a/U4926  ( .A(\w1[3][15] ), .B(n9555), .Z(n8878) );
  XOR \SUBBYTES[3].a/U4925  ( .A(\SUBBYTES[3].a/w3081 ), .B(
        \SUBBYTES[3].a/w3090 ), .Z(n8879) );
  XOR \SUBBYTES[3].a/U4924  ( .A(n8881), .B(n8880), .Z(\SUBBYTES[3].a/w3105 )
         );
  XOR \SUBBYTES[3].a/U4923  ( .A(n8883), .B(n8882), .Z(n8880) );
  XOR \SUBBYTES[3].a/U4922  ( .A(\w1[3][15] ), .B(\SUBBYTES[3].a/w3189 ), .Z(
        n8881) );
  XOR \SUBBYTES[3].a/U4921  ( .A(\SUBBYTES[3].a/w3096 ), .B(
        \SUBBYTES[3].a/w3099 ), .Z(n8882) );
  XOR \SUBBYTES[3].a/U4920  ( .A(\SUBBYTES[3].a/w3082 ), .B(
        \SUBBYTES[3].a/w3084 ), .Z(n8883) );
  XOR \SUBBYTES[3].a/U4919  ( .A(n8885), .B(n8884), .Z(\SUBBYTES[3].a/w3106 )
         );
  XOR \SUBBYTES[3].a/U4918  ( .A(n9556), .B(n8886), .Z(n8884) );
  XOR \SUBBYTES[3].a/U4917  ( .A(\w1[3][13] ), .B(n9557), .Z(n8885) );
  XOR \SUBBYTES[3].a/U4916  ( .A(\SUBBYTES[3].a/w3096 ), .B(
        \SUBBYTES[3].a/w3097 ), .Z(n8886) );
  XOR \SUBBYTES[3].a/U4915  ( .A(n8888), .B(n8887), .Z(\SUBBYTES[3].a/w3122 )
         );
  XOR \SUBBYTES[3].a/U4914  ( .A(\w1[3][9] ), .B(n8889), .Z(n8887) );
  XOR \SUBBYTES[3].a/U4913  ( .A(\SUBBYTES[3].a/w3097 ), .B(
        \SUBBYTES[3].a/w3099 ), .Z(n8888) );
  XOR \SUBBYTES[3].a/U4912  ( .A(\SUBBYTES[3].a/w3081 ), .B(
        \SUBBYTES[3].a/w3082 ), .Z(n8889) );
  XOR \SUBBYTES[3].a/U4911  ( .A(\w1[3][17] ), .B(n8890), .Z(n9558) );
  XOR \SUBBYTES[3].a/U4910  ( .A(\w1[3][19] ), .B(\w1[3][18] ), .Z(n8890) );
  XOR \SUBBYTES[3].a/U4909  ( .A(\w1[3][22] ), .B(n9558), .Z(
        \SUBBYTES[3].a/w2964 ) );
  XOR \SUBBYTES[3].a/U4908  ( .A(\w1[3][16] ), .B(\SUBBYTES[3].a/w2964 ), .Z(
        \SUBBYTES[3].a/w2851 ) );
  XOR \SUBBYTES[3].a/U4907  ( .A(\w1[3][16] ), .B(n8891), .Z(
        \SUBBYTES[3].a/w2852 ) );
  XOR \SUBBYTES[3].a/U4906  ( .A(\w1[3][22] ), .B(\w1[3][21] ), .Z(n8891) );
  XOR \SUBBYTES[3].a/U4905  ( .A(\w1[3][21] ), .B(n9558), .Z(
        \SUBBYTES[3].a/w2982 ) );
  XOR \SUBBYTES[3].a/U4904  ( .A(n8893), .B(n8892), .Z(\SUBBYTES[3].a/w2975 )
         );
  XOR \SUBBYTES[3].a/U4903  ( .A(\w1[3][19] ), .B(\w1[3][17] ), .Z(n8892) );
  XOR \SUBBYTES[3].a/U4902  ( .A(\w1[3][23] ), .B(\w1[3][20] ), .Z(n8893) );
  XOR \SUBBYTES[3].a/U4901  ( .A(\w1[3][16] ), .B(\SUBBYTES[3].a/w2975 ), .Z(
        \SUBBYTES[3].a/w2854 ) );
  XOR \SUBBYTES[3].a/U4900  ( .A(n8895), .B(n8894), .Z(\SUBBYTES[3].a/w2962 )
         );
  XOR \SUBBYTES[3].a/U4899  ( .A(\SUBBYTES[3].a/w2923 ), .B(n1002), .Z(n8894)
         );
  XOR \SUBBYTES[3].a/U4898  ( .A(\SUBBYTES[3].a/w2916 ), .B(
        \SUBBYTES[3].a/w2919 ), .Z(n8895) );
  XOR \SUBBYTES[3].a/U4897  ( .A(n8897), .B(n8896), .Z(\SUBBYTES[3].a/w2963 )
         );
  XOR \SUBBYTES[3].a/U4896  ( .A(\SUBBYTES[3].a/w2923 ), .B(n8419), .Z(n8896)
         );
  XOR \SUBBYTES[3].a/U4895  ( .A(\SUBBYTES[3].a/w2916 ), .B(n8418), .Z(n8897)
         );
  XOR \SUBBYTES[3].a/U4894  ( .A(\SUBBYTES[3].a/w2975 ), .B(n8898), .Z(
        \SUBBYTES[3].a/w2965 ) );
  XOR \SUBBYTES[3].a/U4893  ( .A(\w1[3][22] ), .B(\w1[3][21] ), .Z(n8898) );
  XOR \SUBBYTES[3].a/U4892  ( .A(n8900), .B(n8899), .Z(\SUBBYTES[3].a/w2966 )
         );
  XOR \SUBBYTES[3].a/U4891  ( .A(n8419), .B(n1002), .Z(n8899) );
  XOR \SUBBYTES[3].a/U4890  ( .A(n8418), .B(\SUBBYTES[3].a/w2919 ), .Z(n8900)
         );
  XOR \SUBBYTES[3].a/U4889  ( .A(\w1[3][23] ), .B(\w1[3][18] ), .Z(n9564) );
  XOR \SUBBYTES[3].a/U4888  ( .A(n9564), .B(n8901), .Z(\SUBBYTES[3].a/w2967 )
         );
  XOR \SUBBYTES[3].a/U4887  ( .A(\w1[3][21] ), .B(\w1[3][20] ), .Z(n8901) );
  XOR \SUBBYTES[3].a/U4886  ( .A(\w1[3][23] ), .B(\SUBBYTES[3].a/w2852 ), .Z(
        \SUBBYTES[3].a/w2855 ) );
  XOR \SUBBYTES[3].a/U4885  ( .A(\w1[3][17] ), .B(\SUBBYTES[3].a/w2852 ), .Z(
        \SUBBYTES[3].a/w2856 ) );
  XOR \SUBBYTES[3].a/U4884  ( .A(\w1[3][20] ), .B(\SUBBYTES[3].a/w2852 ), .Z(
        \SUBBYTES[3].a/w2857 ) );
  XOR \SUBBYTES[3].a/U4883  ( .A(\SUBBYTES[3].a/w2856 ), .B(n9564), .Z(
        \SUBBYTES[3].a/w2858 ) );
  XOR \SUBBYTES[3].a/U4882  ( .A(n9564), .B(n8902), .Z(\SUBBYTES[3].a/w2943 )
         );
  XOR \SUBBYTES[3].a/U4881  ( .A(\w1[3][20] ), .B(\w1[3][17] ), .Z(n8902) );
  XOR \SUBBYTES[3].a/U4880  ( .A(n8904), .B(n8903), .Z(n9561) );
  XOR \SUBBYTES[3].a/U4879  ( .A(\w1[3][20] ), .B(n8905), .Z(n8903) );
  XOR \SUBBYTES[3].a/U4878  ( .A(\SUBBYTES[3].a/w2908 ), .B(\w1[3][22] ), .Z(
        n8904) );
  XOR \SUBBYTES[3].a/U4877  ( .A(\SUBBYTES[3].a/w2882 ), .B(
        \SUBBYTES[3].a/w2889 ), .Z(n8905) );
  XOR \SUBBYTES[3].a/U4876  ( .A(n8907), .B(n8906), .Z(n9559) );
  XOR \SUBBYTES[3].a/U4875  ( .A(\w1[3][17] ), .B(n8908), .Z(n8906) );
  XOR \SUBBYTES[3].a/U4874  ( .A(\SUBBYTES[3].a/w2907 ), .B(\w1[3][21] ), .Z(
        n8907) );
  XOR \SUBBYTES[3].a/U4873  ( .A(\SUBBYTES[3].a/w2883 ), .B(
        \SUBBYTES[3].a/w2890 ), .Z(n8908) );
  XOR \SUBBYTES[3].a/U4872  ( .A(n9561), .B(n9559), .Z(\SUBBYTES[3].a/w2913 )
         );
  XOR \SUBBYTES[3].a/U4871  ( .A(\w1[3][21] ), .B(n8909), .Z(n9562) );
  XOR \SUBBYTES[3].a/U4870  ( .A(\SUBBYTES[3].a/w2875 ), .B(
        \SUBBYTES[3].a/w2885 ), .Z(n8909) );
  XOR \SUBBYTES[3].a/U4869  ( .A(n8911), .B(n8910), .Z(\SUBBYTES[3].a/w2900 )
         );
  XOR \SUBBYTES[3].a/U4868  ( .A(n9562), .B(n8912), .Z(n8910) );
  XOR \SUBBYTES[3].a/U4867  ( .A(\w1[3][20] ), .B(\SUBBYTES[3].a/w2964 ), .Z(
        n8911) );
  XOR \SUBBYTES[3].a/U4866  ( .A(\SUBBYTES[3].a/w2877 ), .B(
        \SUBBYTES[3].a/w2882 ), .Z(n8912) );
  XOR \SUBBYTES[3].a/U4865  ( .A(n8914), .B(n8913), .Z(n9560) );
  XOR \SUBBYTES[3].a/U4864  ( .A(\SUBBYTES[3].a/w2910 ), .B(\w1[3][23] ), .Z(
        n8913) );
  XOR \SUBBYTES[3].a/U4863  ( .A(\SUBBYTES[3].a/w2885 ), .B(
        \SUBBYTES[3].a/w2892 ), .Z(n8914) );
  XOR \SUBBYTES[3].a/U4862  ( .A(n9559), .B(n9560), .Z(\SUBBYTES[3].a/w2912 )
         );
  XOR \SUBBYTES[3].a/U4861  ( .A(\w1[3][19] ), .B(n8915), .Z(n9563) );
  XOR \SUBBYTES[3].a/U4860  ( .A(\SUBBYTES[3].a/w2874 ), .B(
        \SUBBYTES[3].a/w2877 ), .Z(n8915) );
  XOR \SUBBYTES[3].a/U4859  ( .A(n8917), .B(n8916), .Z(\SUBBYTES[3].a/w2901 )
         );
  XOR \SUBBYTES[3].a/U4858  ( .A(n9563), .B(n8918), .Z(n8916) );
  XOR \SUBBYTES[3].a/U4857  ( .A(\w1[3][22] ), .B(\SUBBYTES[3].a/w2943 ), .Z(
        n8917) );
  XOR \SUBBYTES[3].a/U4856  ( .A(\SUBBYTES[3].a/w2882 ), .B(
        \SUBBYTES[3].a/w2883 ), .Z(n8918) );
  XOR \SUBBYTES[3].a/U4855  ( .A(n9561), .B(n9560), .Z(\SUBBYTES[3].a/w2921 )
         );
  XOR \SUBBYTES[3].a/U4854  ( .A(n8920), .B(n8919), .Z(\SUBBYTES[3].a/w2922 )
         );
  XOR \SUBBYTES[3].a/U4853  ( .A(\w1[3][23] ), .B(n9562), .Z(n8919) );
  XOR \SUBBYTES[3].a/U4852  ( .A(\SUBBYTES[3].a/w2874 ), .B(
        \SUBBYTES[3].a/w2883 ), .Z(n8920) );
  XOR \SUBBYTES[3].a/U4851  ( .A(n8922), .B(n8921), .Z(\SUBBYTES[3].a/w2898 )
         );
  XOR \SUBBYTES[3].a/U4850  ( .A(n8924), .B(n8923), .Z(n8921) );
  XOR \SUBBYTES[3].a/U4849  ( .A(\w1[3][23] ), .B(\SUBBYTES[3].a/w2982 ), .Z(
        n8922) );
  XOR \SUBBYTES[3].a/U4848  ( .A(\SUBBYTES[3].a/w2889 ), .B(
        \SUBBYTES[3].a/w2892 ), .Z(n8923) );
  XOR \SUBBYTES[3].a/U4847  ( .A(\SUBBYTES[3].a/w2875 ), .B(
        \SUBBYTES[3].a/w2877 ), .Z(n8924) );
  XOR \SUBBYTES[3].a/U4846  ( .A(n8926), .B(n8925), .Z(\SUBBYTES[3].a/w2899 )
         );
  XOR \SUBBYTES[3].a/U4845  ( .A(n9563), .B(n8927), .Z(n8925) );
  XOR \SUBBYTES[3].a/U4844  ( .A(\w1[3][21] ), .B(n9564), .Z(n8926) );
  XOR \SUBBYTES[3].a/U4843  ( .A(\SUBBYTES[3].a/w2889 ), .B(
        \SUBBYTES[3].a/w2890 ), .Z(n8927) );
  XOR \SUBBYTES[3].a/U4842  ( .A(n8929), .B(n8928), .Z(\SUBBYTES[3].a/w2915 )
         );
  XOR \SUBBYTES[3].a/U4841  ( .A(\w1[3][17] ), .B(n8930), .Z(n8928) );
  XOR \SUBBYTES[3].a/U4840  ( .A(\SUBBYTES[3].a/w2890 ), .B(
        \SUBBYTES[3].a/w2892 ), .Z(n8929) );
  XOR \SUBBYTES[3].a/U4839  ( .A(\SUBBYTES[3].a/w2874 ), .B(
        \SUBBYTES[3].a/w2875 ), .Z(n8930) );
  XOR \SUBBYTES[3].a/U4838  ( .A(\w1[3][25] ), .B(n8931), .Z(n9565) );
  XOR \SUBBYTES[3].a/U4837  ( .A(\w1[3][27] ), .B(\w1[3][26] ), .Z(n8931) );
  XOR \SUBBYTES[3].a/U4836  ( .A(\w1[3][30] ), .B(n9565), .Z(
        \SUBBYTES[3].a/w2757 ) );
  XOR \SUBBYTES[3].a/U4835  ( .A(\w1[3][24] ), .B(\SUBBYTES[3].a/w2757 ), .Z(
        \SUBBYTES[3].a/w2644 ) );
  XOR \SUBBYTES[3].a/U4834  ( .A(\w1[3][24] ), .B(n8932), .Z(
        \SUBBYTES[3].a/w2645 ) );
  XOR \SUBBYTES[3].a/U4833  ( .A(\w1[3][30] ), .B(\w1[3][29] ), .Z(n8932) );
  XOR \SUBBYTES[3].a/U4832  ( .A(\w1[3][29] ), .B(n9565), .Z(
        \SUBBYTES[3].a/w2775 ) );
  XOR \SUBBYTES[3].a/U4831  ( .A(n8934), .B(n8933), .Z(\SUBBYTES[3].a/w2768 )
         );
  XOR \SUBBYTES[3].a/U4830  ( .A(\w1[3][27] ), .B(\w1[3][25] ), .Z(n8933) );
  XOR \SUBBYTES[3].a/U4829  ( .A(\w1[3][31] ), .B(\w1[3][28] ), .Z(n8934) );
  XOR \SUBBYTES[3].a/U4828  ( .A(\w1[3][24] ), .B(\SUBBYTES[3].a/w2768 ), .Z(
        \SUBBYTES[3].a/w2647 ) );
  XOR \SUBBYTES[3].a/U4827  ( .A(n8936), .B(n8935), .Z(\SUBBYTES[3].a/w2755 )
         );
  XOR \SUBBYTES[3].a/U4826  ( .A(\SUBBYTES[3].a/w2716 ), .B(n1001), .Z(n8935)
         );
  XOR \SUBBYTES[3].a/U4825  ( .A(\SUBBYTES[3].a/w2709 ), .B(
        \SUBBYTES[3].a/w2712 ), .Z(n8936) );
  XOR \SUBBYTES[3].a/U4824  ( .A(n8938), .B(n8937), .Z(\SUBBYTES[3].a/w2756 )
         );
  XOR \SUBBYTES[3].a/U4823  ( .A(\SUBBYTES[3].a/w2716 ), .B(n8417), .Z(n8937)
         );
  XOR \SUBBYTES[3].a/U4822  ( .A(\SUBBYTES[3].a/w2709 ), .B(n8416), .Z(n8938)
         );
  XOR \SUBBYTES[3].a/U4821  ( .A(\SUBBYTES[3].a/w2768 ), .B(n8939), .Z(
        \SUBBYTES[3].a/w2758 ) );
  XOR \SUBBYTES[3].a/U4820  ( .A(\w1[3][30] ), .B(\w1[3][29] ), .Z(n8939) );
  XOR \SUBBYTES[3].a/U4819  ( .A(n8941), .B(n8940), .Z(\SUBBYTES[3].a/w2759 )
         );
  XOR \SUBBYTES[3].a/U4818  ( .A(n8417), .B(n1001), .Z(n8940) );
  XOR \SUBBYTES[3].a/U4817  ( .A(n8416), .B(\SUBBYTES[3].a/w2712 ), .Z(n8941)
         );
  XOR \SUBBYTES[3].a/U4816  ( .A(\w1[3][31] ), .B(\w1[3][26] ), .Z(n9571) );
  XOR \SUBBYTES[3].a/U4815  ( .A(n9571), .B(n8942), .Z(\SUBBYTES[3].a/w2760 )
         );
  XOR \SUBBYTES[3].a/U4814  ( .A(\w1[3][29] ), .B(\w1[3][28] ), .Z(n8942) );
  XOR \SUBBYTES[3].a/U4813  ( .A(\w1[3][31] ), .B(\SUBBYTES[3].a/w2645 ), .Z(
        \SUBBYTES[3].a/w2648 ) );
  XOR \SUBBYTES[3].a/U4812  ( .A(\w1[3][25] ), .B(\SUBBYTES[3].a/w2645 ), .Z(
        \SUBBYTES[3].a/w2649 ) );
  XOR \SUBBYTES[3].a/U4811  ( .A(\w1[3][28] ), .B(\SUBBYTES[3].a/w2645 ), .Z(
        \SUBBYTES[3].a/w2650 ) );
  XOR \SUBBYTES[3].a/U4810  ( .A(\SUBBYTES[3].a/w2649 ), .B(n9571), .Z(
        \SUBBYTES[3].a/w2651 ) );
  XOR \SUBBYTES[3].a/U4809  ( .A(n9571), .B(n8943), .Z(\SUBBYTES[3].a/w2736 )
         );
  XOR \SUBBYTES[3].a/U4808  ( .A(\w1[3][28] ), .B(\w1[3][25] ), .Z(n8943) );
  XOR \SUBBYTES[3].a/U4807  ( .A(n8945), .B(n8944), .Z(n9568) );
  XOR \SUBBYTES[3].a/U4806  ( .A(\w1[3][28] ), .B(n8946), .Z(n8944) );
  XOR \SUBBYTES[3].a/U4805  ( .A(\SUBBYTES[3].a/w2701 ), .B(\w1[3][30] ), .Z(
        n8945) );
  XOR \SUBBYTES[3].a/U4804  ( .A(\SUBBYTES[3].a/w2675 ), .B(
        \SUBBYTES[3].a/w2682 ), .Z(n8946) );
  XOR \SUBBYTES[3].a/U4803  ( .A(n8948), .B(n8947), .Z(n9566) );
  XOR \SUBBYTES[3].a/U4802  ( .A(\w1[3][25] ), .B(n8949), .Z(n8947) );
  XOR \SUBBYTES[3].a/U4801  ( .A(\SUBBYTES[3].a/w2700 ), .B(\w1[3][29] ), .Z(
        n8948) );
  XOR \SUBBYTES[3].a/U4800  ( .A(\SUBBYTES[3].a/w2676 ), .B(
        \SUBBYTES[3].a/w2683 ), .Z(n8949) );
  XOR \SUBBYTES[3].a/U4799  ( .A(n9568), .B(n9566), .Z(\SUBBYTES[3].a/w2706 )
         );
  XOR \SUBBYTES[3].a/U4798  ( .A(\w1[3][29] ), .B(n8950), .Z(n9569) );
  XOR \SUBBYTES[3].a/U4797  ( .A(\SUBBYTES[3].a/w2668 ), .B(
        \SUBBYTES[3].a/w2678 ), .Z(n8950) );
  XOR \SUBBYTES[3].a/U4796  ( .A(n8952), .B(n8951), .Z(\SUBBYTES[3].a/w2693 )
         );
  XOR \SUBBYTES[3].a/U4795  ( .A(n9569), .B(n8953), .Z(n8951) );
  XOR \SUBBYTES[3].a/U4794  ( .A(\w1[3][28] ), .B(\SUBBYTES[3].a/w2757 ), .Z(
        n8952) );
  XOR \SUBBYTES[3].a/U4793  ( .A(\SUBBYTES[3].a/w2670 ), .B(
        \SUBBYTES[3].a/w2675 ), .Z(n8953) );
  XOR \SUBBYTES[3].a/U4792  ( .A(n8955), .B(n8954), .Z(n9567) );
  XOR \SUBBYTES[3].a/U4791  ( .A(\SUBBYTES[3].a/w2703 ), .B(\w1[3][31] ), .Z(
        n8954) );
  XOR \SUBBYTES[3].a/U4790  ( .A(\SUBBYTES[3].a/w2678 ), .B(
        \SUBBYTES[3].a/w2685 ), .Z(n8955) );
  XOR \SUBBYTES[3].a/U4789  ( .A(n9566), .B(n9567), .Z(\SUBBYTES[3].a/w2705 )
         );
  XOR \SUBBYTES[3].a/U4788  ( .A(\w1[3][27] ), .B(n8956), .Z(n9570) );
  XOR \SUBBYTES[3].a/U4787  ( .A(\SUBBYTES[3].a/w2667 ), .B(
        \SUBBYTES[3].a/w2670 ), .Z(n8956) );
  XOR \SUBBYTES[3].a/U4786  ( .A(n8958), .B(n8957), .Z(\SUBBYTES[3].a/w2694 )
         );
  XOR \SUBBYTES[3].a/U4785  ( .A(n9570), .B(n8959), .Z(n8957) );
  XOR \SUBBYTES[3].a/U4784  ( .A(\w1[3][30] ), .B(\SUBBYTES[3].a/w2736 ), .Z(
        n8958) );
  XOR \SUBBYTES[3].a/U4783  ( .A(\SUBBYTES[3].a/w2675 ), .B(
        \SUBBYTES[3].a/w2676 ), .Z(n8959) );
  XOR \SUBBYTES[3].a/U4782  ( .A(n9568), .B(n9567), .Z(\SUBBYTES[3].a/w2714 )
         );
  XOR \SUBBYTES[3].a/U4781  ( .A(n8961), .B(n8960), .Z(\SUBBYTES[3].a/w2715 )
         );
  XOR \SUBBYTES[3].a/U4780  ( .A(\w1[3][31] ), .B(n9569), .Z(n8960) );
  XOR \SUBBYTES[3].a/U4779  ( .A(\SUBBYTES[3].a/w2667 ), .B(
        \SUBBYTES[3].a/w2676 ), .Z(n8961) );
  XOR \SUBBYTES[3].a/U4778  ( .A(n8963), .B(n8962), .Z(\SUBBYTES[3].a/w2691 )
         );
  XOR \SUBBYTES[3].a/U4777  ( .A(n8965), .B(n8964), .Z(n8962) );
  XOR \SUBBYTES[3].a/U4776  ( .A(\w1[3][31] ), .B(\SUBBYTES[3].a/w2775 ), .Z(
        n8963) );
  XOR \SUBBYTES[3].a/U4775  ( .A(\SUBBYTES[3].a/w2682 ), .B(
        \SUBBYTES[3].a/w2685 ), .Z(n8964) );
  XOR \SUBBYTES[3].a/U4774  ( .A(\SUBBYTES[3].a/w2668 ), .B(
        \SUBBYTES[3].a/w2670 ), .Z(n8965) );
  XOR \SUBBYTES[3].a/U4773  ( .A(n8967), .B(n8966), .Z(\SUBBYTES[3].a/w2692 )
         );
  XOR \SUBBYTES[3].a/U4772  ( .A(n9570), .B(n8968), .Z(n8966) );
  XOR \SUBBYTES[3].a/U4771  ( .A(\w1[3][29] ), .B(n9571), .Z(n8967) );
  XOR \SUBBYTES[3].a/U4770  ( .A(\SUBBYTES[3].a/w2682 ), .B(
        \SUBBYTES[3].a/w2683 ), .Z(n8968) );
  XOR \SUBBYTES[3].a/U4769  ( .A(n8970), .B(n8969), .Z(\SUBBYTES[3].a/w2708 )
         );
  XOR \SUBBYTES[3].a/U4768  ( .A(\w1[3][25] ), .B(n8971), .Z(n8969) );
  XOR \SUBBYTES[3].a/U4767  ( .A(\SUBBYTES[3].a/w2683 ), .B(
        \SUBBYTES[3].a/w2685 ), .Z(n8970) );
  XOR \SUBBYTES[3].a/U4766  ( .A(\SUBBYTES[3].a/w2667 ), .B(
        \SUBBYTES[3].a/w2668 ), .Z(n8971) );
  XOR \SUBBYTES[3].a/U4765  ( .A(\w1[3][33] ), .B(n8972), .Z(n9572) );
  XOR \SUBBYTES[3].a/U4764  ( .A(\w1[3][35] ), .B(\w1[3][34] ), .Z(n8972) );
  XOR \SUBBYTES[3].a/U4763  ( .A(\w1[3][38] ), .B(n9572), .Z(
        \SUBBYTES[3].a/w2550 ) );
  XOR \SUBBYTES[3].a/U4762  ( .A(\w1[3][32] ), .B(\SUBBYTES[3].a/w2550 ), .Z(
        \SUBBYTES[3].a/w2437 ) );
  XOR \SUBBYTES[3].a/U4761  ( .A(\w1[3][32] ), .B(n8973), .Z(
        \SUBBYTES[3].a/w2438 ) );
  XOR \SUBBYTES[3].a/U4760  ( .A(\w1[3][38] ), .B(\w1[3][37] ), .Z(n8973) );
  XOR \SUBBYTES[3].a/U4759  ( .A(\w1[3][37] ), .B(n9572), .Z(
        \SUBBYTES[3].a/w2568 ) );
  XOR \SUBBYTES[3].a/U4758  ( .A(n8975), .B(n8974), .Z(\SUBBYTES[3].a/w2561 )
         );
  XOR \SUBBYTES[3].a/U4757  ( .A(\w1[3][35] ), .B(\w1[3][33] ), .Z(n8974) );
  XOR \SUBBYTES[3].a/U4756  ( .A(\w1[3][39] ), .B(\w1[3][36] ), .Z(n8975) );
  XOR \SUBBYTES[3].a/U4755  ( .A(\w1[3][32] ), .B(\SUBBYTES[3].a/w2561 ), .Z(
        \SUBBYTES[3].a/w2440 ) );
  XOR \SUBBYTES[3].a/U4754  ( .A(n8977), .B(n8976), .Z(\SUBBYTES[3].a/w2548 )
         );
  XOR \SUBBYTES[3].a/U4753  ( .A(\SUBBYTES[3].a/w2509 ), .B(n1000), .Z(n8976)
         );
  XOR \SUBBYTES[3].a/U4752  ( .A(\SUBBYTES[3].a/w2502 ), .B(
        \SUBBYTES[3].a/w2505 ), .Z(n8977) );
  XOR \SUBBYTES[3].a/U4751  ( .A(n8979), .B(n8978), .Z(\SUBBYTES[3].a/w2549 )
         );
  XOR \SUBBYTES[3].a/U4750  ( .A(\SUBBYTES[3].a/w2509 ), .B(n8415), .Z(n8978)
         );
  XOR \SUBBYTES[3].a/U4749  ( .A(\SUBBYTES[3].a/w2502 ), .B(n8414), .Z(n8979)
         );
  XOR \SUBBYTES[3].a/U4748  ( .A(\SUBBYTES[3].a/w2561 ), .B(n8980), .Z(
        \SUBBYTES[3].a/w2551 ) );
  XOR \SUBBYTES[3].a/U4747  ( .A(\w1[3][38] ), .B(\w1[3][37] ), .Z(n8980) );
  XOR \SUBBYTES[3].a/U4746  ( .A(n8982), .B(n8981), .Z(\SUBBYTES[3].a/w2552 )
         );
  XOR \SUBBYTES[3].a/U4745  ( .A(n8415), .B(n1000), .Z(n8981) );
  XOR \SUBBYTES[3].a/U4744  ( .A(n8414), .B(\SUBBYTES[3].a/w2505 ), .Z(n8982)
         );
  XOR \SUBBYTES[3].a/U4743  ( .A(\w1[3][39] ), .B(\w1[3][34] ), .Z(n9578) );
  XOR \SUBBYTES[3].a/U4742  ( .A(n9578), .B(n8983), .Z(\SUBBYTES[3].a/w2553 )
         );
  XOR \SUBBYTES[3].a/U4741  ( .A(\w1[3][37] ), .B(\w1[3][36] ), .Z(n8983) );
  XOR \SUBBYTES[3].a/U4740  ( .A(\w1[3][39] ), .B(\SUBBYTES[3].a/w2438 ), .Z(
        \SUBBYTES[3].a/w2441 ) );
  XOR \SUBBYTES[3].a/U4739  ( .A(\w1[3][33] ), .B(\SUBBYTES[3].a/w2438 ), .Z(
        \SUBBYTES[3].a/w2442 ) );
  XOR \SUBBYTES[3].a/U4738  ( .A(\w1[3][36] ), .B(\SUBBYTES[3].a/w2438 ), .Z(
        \SUBBYTES[3].a/w2443 ) );
  XOR \SUBBYTES[3].a/U4737  ( .A(\SUBBYTES[3].a/w2442 ), .B(n9578), .Z(
        \SUBBYTES[3].a/w2444 ) );
  XOR \SUBBYTES[3].a/U4736  ( .A(n9578), .B(n8984), .Z(\SUBBYTES[3].a/w2529 )
         );
  XOR \SUBBYTES[3].a/U4735  ( .A(\w1[3][36] ), .B(\w1[3][33] ), .Z(n8984) );
  XOR \SUBBYTES[3].a/U4734  ( .A(n8986), .B(n8985), .Z(n9575) );
  XOR \SUBBYTES[3].a/U4733  ( .A(\w1[3][36] ), .B(n8987), .Z(n8985) );
  XOR \SUBBYTES[3].a/U4732  ( .A(\SUBBYTES[3].a/w2494 ), .B(\w1[3][38] ), .Z(
        n8986) );
  XOR \SUBBYTES[3].a/U4731  ( .A(\SUBBYTES[3].a/w2468 ), .B(
        \SUBBYTES[3].a/w2475 ), .Z(n8987) );
  XOR \SUBBYTES[3].a/U4730  ( .A(n8989), .B(n8988), .Z(n9573) );
  XOR \SUBBYTES[3].a/U4729  ( .A(\w1[3][33] ), .B(n8990), .Z(n8988) );
  XOR \SUBBYTES[3].a/U4728  ( .A(\SUBBYTES[3].a/w2493 ), .B(\w1[3][37] ), .Z(
        n8989) );
  XOR \SUBBYTES[3].a/U4727  ( .A(\SUBBYTES[3].a/w2469 ), .B(
        \SUBBYTES[3].a/w2476 ), .Z(n8990) );
  XOR \SUBBYTES[3].a/U4726  ( .A(n9575), .B(n9573), .Z(\SUBBYTES[3].a/w2499 )
         );
  XOR \SUBBYTES[3].a/U4725  ( .A(\w1[3][37] ), .B(n8991), .Z(n9576) );
  XOR \SUBBYTES[3].a/U4724  ( .A(\SUBBYTES[3].a/w2461 ), .B(
        \SUBBYTES[3].a/w2471 ), .Z(n8991) );
  XOR \SUBBYTES[3].a/U4723  ( .A(n8993), .B(n8992), .Z(\SUBBYTES[3].a/w2486 )
         );
  XOR \SUBBYTES[3].a/U4722  ( .A(n9576), .B(n8994), .Z(n8992) );
  XOR \SUBBYTES[3].a/U4721  ( .A(\w1[3][36] ), .B(\SUBBYTES[3].a/w2550 ), .Z(
        n8993) );
  XOR \SUBBYTES[3].a/U4720  ( .A(\SUBBYTES[3].a/w2463 ), .B(
        \SUBBYTES[3].a/w2468 ), .Z(n8994) );
  XOR \SUBBYTES[3].a/U4719  ( .A(n8996), .B(n8995), .Z(n9574) );
  XOR \SUBBYTES[3].a/U4718  ( .A(\SUBBYTES[3].a/w2496 ), .B(\w1[3][39] ), .Z(
        n8995) );
  XOR \SUBBYTES[3].a/U4717  ( .A(\SUBBYTES[3].a/w2471 ), .B(
        \SUBBYTES[3].a/w2478 ), .Z(n8996) );
  XOR \SUBBYTES[3].a/U4716  ( .A(n9573), .B(n9574), .Z(\SUBBYTES[3].a/w2498 )
         );
  XOR \SUBBYTES[3].a/U4715  ( .A(\w1[3][35] ), .B(n8997), .Z(n9577) );
  XOR \SUBBYTES[3].a/U4714  ( .A(\SUBBYTES[3].a/w2460 ), .B(
        \SUBBYTES[3].a/w2463 ), .Z(n8997) );
  XOR \SUBBYTES[3].a/U4713  ( .A(n8999), .B(n8998), .Z(\SUBBYTES[3].a/w2487 )
         );
  XOR \SUBBYTES[3].a/U4712  ( .A(n9577), .B(n9000), .Z(n8998) );
  XOR \SUBBYTES[3].a/U4711  ( .A(\w1[3][38] ), .B(\SUBBYTES[3].a/w2529 ), .Z(
        n8999) );
  XOR \SUBBYTES[3].a/U4710  ( .A(\SUBBYTES[3].a/w2468 ), .B(
        \SUBBYTES[3].a/w2469 ), .Z(n9000) );
  XOR \SUBBYTES[3].a/U4709  ( .A(n9575), .B(n9574), .Z(\SUBBYTES[3].a/w2507 )
         );
  XOR \SUBBYTES[3].a/U4708  ( .A(n9002), .B(n9001), .Z(\SUBBYTES[3].a/w2508 )
         );
  XOR \SUBBYTES[3].a/U4707  ( .A(\w1[3][39] ), .B(n9576), .Z(n9001) );
  XOR \SUBBYTES[3].a/U4706  ( .A(\SUBBYTES[3].a/w2460 ), .B(
        \SUBBYTES[3].a/w2469 ), .Z(n9002) );
  XOR \SUBBYTES[3].a/U4705  ( .A(n9004), .B(n9003), .Z(\SUBBYTES[3].a/w2484 )
         );
  XOR \SUBBYTES[3].a/U4704  ( .A(n9006), .B(n9005), .Z(n9003) );
  XOR \SUBBYTES[3].a/U4703  ( .A(\w1[3][39] ), .B(\SUBBYTES[3].a/w2568 ), .Z(
        n9004) );
  XOR \SUBBYTES[3].a/U4702  ( .A(\SUBBYTES[3].a/w2475 ), .B(
        \SUBBYTES[3].a/w2478 ), .Z(n9005) );
  XOR \SUBBYTES[3].a/U4701  ( .A(\SUBBYTES[3].a/w2461 ), .B(
        \SUBBYTES[3].a/w2463 ), .Z(n9006) );
  XOR \SUBBYTES[3].a/U4700  ( .A(n9008), .B(n9007), .Z(\SUBBYTES[3].a/w2485 )
         );
  XOR \SUBBYTES[3].a/U4699  ( .A(n9577), .B(n9009), .Z(n9007) );
  XOR \SUBBYTES[3].a/U4698  ( .A(\w1[3][37] ), .B(n9578), .Z(n9008) );
  XOR \SUBBYTES[3].a/U4697  ( .A(\SUBBYTES[3].a/w2475 ), .B(
        \SUBBYTES[3].a/w2476 ), .Z(n9009) );
  XOR \SUBBYTES[3].a/U4696  ( .A(n9011), .B(n9010), .Z(\SUBBYTES[3].a/w2501 )
         );
  XOR \SUBBYTES[3].a/U4695  ( .A(\w1[3][33] ), .B(n9012), .Z(n9010) );
  XOR \SUBBYTES[3].a/U4694  ( .A(\SUBBYTES[3].a/w2476 ), .B(
        \SUBBYTES[3].a/w2478 ), .Z(n9011) );
  XOR \SUBBYTES[3].a/U4693  ( .A(\SUBBYTES[3].a/w2460 ), .B(
        \SUBBYTES[3].a/w2461 ), .Z(n9012) );
  XOR \SUBBYTES[3].a/U4692  ( .A(\w1[3][41] ), .B(n9013), .Z(n9579) );
  XOR \SUBBYTES[3].a/U4691  ( .A(\w1[3][43] ), .B(\w1[3][42] ), .Z(n9013) );
  XOR \SUBBYTES[3].a/U4690  ( .A(\w1[3][46] ), .B(n9579), .Z(
        \SUBBYTES[3].a/w2343 ) );
  XOR \SUBBYTES[3].a/U4689  ( .A(\w1[3][40] ), .B(\SUBBYTES[3].a/w2343 ), .Z(
        \SUBBYTES[3].a/w2230 ) );
  XOR \SUBBYTES[3].a/U4688  ( .A(\w1[3][40] ), .B(n9014), .Z(
        \SUBBYTES[3].a/w2231 ) );
  XOR \SUBBYTES[3].a/U4687  ( .A(\w1[3][46] ), .B(\w1[3][45] ), .Z(n9014) );
  XOR \SUBBYTES[3].a/U4686  ( .A(\w1[3][45] ), .B(n9579), .Z(
        \SUBBYTES[3].a/w2361 ) );
  XOR \SUBBYTES[3].a/U4685  ( .A(n9016), .B(n9015), .Z(\SUBBYTES[3].a/w2354 )
         );
  XOR \SUBBYTES[3].a/U4684  ( .A(\w1[3][43] ), .B(\w1[3][41] ), .Z(n9015) );
  XOR \SUBBYTES[3].a/U4683  ( .A(\w1[3][47] ), .B(\w1[3][44] ), .Z(n9016) );
  XOR \SUBBYTES[3].a/U4682  ( .A(\w1[3][40] ), .B(\SUBBYTES[3].a/w2354 ), .Z(
        \SUBBYTES[3].a/w2233 ) );
  XOR \SUBBYTES[3].a/U4681  ( .A(n9018), .B(n9017), .Z(\SUBBYTES[3].a/w2341 )
         );
  XOR \SUBBYTES[3].a/U4680  ( .A(\SUBBYTES[3].a/w2302 ), .B(n999), .Z(n9017)
         );
  XOR \SUBBYTES[3].a/U4679  ( .A(\SUBBYTES[3].a/w2295 ), .B(
        \SUBBYTES[3].a/w2298 ), .Z(n9018) );
  XOR \SUBBYTES[3].a/U4678  ( .A(n9020), .B(n9019), .Z(\SUBBYTES[3].a/w2342 )
         );
  XOR \SUBBYTES[3].a/U4677  ( .A(\SUBBYTES[3].a/w2302 ), .B(n8413), .Z(n9019)
         );
  XOR \SUBBYTES[3].a/U4676  ( .A(\SUBBYTES[3].a/w2295 ), .B(n8412), .Z(n9020)
         );
  XOR \SUBBYTES[3].a/U4675  ( .A(\SUBBYTES[3].a/w2354 ), .B(n9021), .Z(
        \SUBBYTES[3].a/w2344 ) );
  XOR \SUBBYTES[3].a/U4674  ( .A(\w1[3][46] ), .B(\w1[3][45] ), .Z(n9021) );
  XOR \SUBBYTES[3].a/U4673  ( .A(n9023), .B(n9022), .Z(\SUBBYTES[3].a/w2345 )
         );
  XOR \SUBBYTES[3].a/U4672  ( .A(n8413), .B(n999), .Z(n9022) );
  XOR \SUBBYTES[3].a/U4671  ( .A(n8412), .B(\SUBBYTES[3].a/w2298 ), .Z(n9023)
         );
  XOR \SUBBYTES[3].a/U4670  ( .A(\w1[3][47] ), .B(\w1[3][42] ), .Z(n9585) );
  XOR \SUBBYTES[3].a/U4669  ( .A(n9585), .B(n9024), .Z(\SUBBYTES[3].a/w2346 )
         );
  XOR \SUBBYTES[3].a/U4668  ( .A(\w1[3][45] ), .B(\w1[3][44] ), .Z(n9024) );
  XOR \SUBBYTES[3].a/U4667  ( .A(\w1[3][47] ), .B(\SUBBYTES[3].a/w2231 ), .Z(
        \SUBBYTES[3].a/w2234 ) );
  XOR \SUBBYTES[3].a/U4666  ( .A(\w1[3][41] ), .B(\SUBBYTES[3].a/w2231 ), .Z(
        \SUBBYTES[3].a/w2235 ) );
  XOR \SUBBYTES[3].a/U4665  ( .A(\w1[3][44] ), .B(\SUBBYTES[3].a/w2231 ), .Z(
        \SUBBYTES[3].a/w2236 ) );
  XOR \SUBBYTES[3].a/U4664  ( .A(\SUBBYTES[3].a/w2235 ), .B(n9585), .Z(
        \SUBBYTES[3].a/w2237 ) );
  XOR \SUBBYTES[3].a/U4663  ( .A(n9585), .B(n9025), .Z(\SUBBYTES[3].a/w2322 )
         );
  XOR \SUBBYTES[3].a/U4662  ( .A(\w1[3][44] ), .B(\w1[3][41] ), .Z(n9025) );
  XOR \SUBBYTES[3].a/U4661  ( .A(n9027), .B(n9026), .Z(n9582) );
  XOR \SUBBYTES[3].a/U4660  ( .A(\w1[3][44] ), .B(n9028), .Z(n9026) );
  XOR \SUBBYTES[3].a/U4659  ( .A(\SUBBYTES[3].a/w2287 ), .B(\w1[3][46] ), .Z(
        n9027) );
  XOR \SUBBYTES[3].a/U4658  ( .A(\SUBBYTES[3].a/w2261 ), .B(
        \SUBBYTES[3].a/w2268 ), .Z(n9028) );
  XOR \SUBBYTES[3].a/U4657  ( .A(n9030), .B(n9029), .Z(n9580) );
  XOR \SUBBYTES[3].a/U4656  ( .A(\w1[3][41] ), .B(n9031), .Z(n9029) );
  XOR \SUBBYTES[3].a/U4655  ( .A(\SUBBYTES[3].a/w2286 ), .B(\w1[3][45] ), .Z(
        n9030) );
  XOR \SUBBYTES[3].a/U4654  ( .A(\SUBBYTES[3].a/w2262 ), .B(
        \SUBBYTES[3].a/w2269 ), .Z(n9031) );
  XOR \SUBBYTES[3].a/U4653  ( .A(n9582), .B(n9580), .Z(\SUBBYTES[3].a/w2292 )
         );
  XOR \SUBBYTES[3].a/U4652  ( .A(\w1[3][45] ), .B(n9032), .Z(n9583) );
  XOR \SUBBYTES[3].a/U4651  ( .A(\SUBBYTES[3].a/w2254 ), .B(
        \SUBBYTES[3].a/w2264 ), .Z(n9032) );
  XOR \SUBBYTES[3].a/U4650  ( .A(n9034), .B(n9033), .Z(\SUBBYTES[3].a/w2279 )
         );
  XOR \SUBBYTES[3].a/U4649  ( .A(n9583), .B(n9035), .Z(n9033) );
  XOR \SUBBYTES[3].a/U4648  ( .A(\w1[3][44] ), .B(\SUBBYTES[3].a/w2343 ), .Z(
        n9034) );
  XOR \SUBBYTES[3].a/U4647  ( .A(\SUBBYTES[3].a/w2256 ), .B(
        \SUBBYTES[3].a/w2261 ), .Z(n9035) );
  XOR \SUBBYTES[3].a/U4646  ( .A(n9037), .B(n9036), .Z(n9581) );
  XOR \SUBBYTES[3].a/U4645  ( .A(\SUBBYTES[3].a/w2289 ), .B(\w1[3][47] ), .Z(
        n9036) );
  XOR \SUBBYTES[3].a/U4644  ( .A(\SUBBYTES[3].a/w2264 ), .B(
        \SUBBYTES[3].a/w2271 ), .Z(n9037) );
  XOR \SUBBYTES[3].a/U4643  ( .A(n9580), .B(n9581), .Z(\SUBBYTES[3].a/w2291 )
         );
  XOR \SUBBYTES[3].a/U4642  ( .A(\w1[3][43] ), .B(n9038), .Z(n9584) );
  XOR \SUBBYTES[3].a/U4641  ( .A(\SUBBYTES[3].a/w2253 ), .B(
        \SUBBYTES[3].a/w2256 ), .Z(n9038) );
  XOR \SUBBYTES[3].a/U4640  ( .A(n9040), .B(n9039), .Z(\SUBBYTES[3].a/w2280 )
         );
  XOR \SUBBYTES[3].a/U4639  ( .A(n9584), .B(n9041), .Z(n9039) );
  XOR \SUBBYTES[3].a/U4638  ( .A(\w1[3][46] ), .B(\SUBBYTES[3].a/w2322 ), .Z(
        n9040) );
  XOR \SUBBYTES[3].a/U4637  ( .A(\SUBBYTES[3].a/w2261 ), .B(
        \SUBBYTES[3].a/w2262 ), .Z(n9041) );
  XOR \SUBBYTES[3].a/U4636  ( .A(n9582), .B(n9581), .Z(\SUBBYTES[3].a/w2300 )
         );
  XOR \SUBBYTES[3].a/U4635  ( .A(n9043), .B(n9042), .Z(\SUBBYTES[3].a/w2301 )
         );
  XOR \SUBBYTES[3].a/U4634  ( .A(\w1[3][47] ), .B(n9583), .Z(n9042) );
  XOR \SUBBYTES[3].a/U4633  ( .A(\SUBBYTES[3].a/w2253 ), .B(
        \SUBBYTES[3].a/w2262 ), .Z(n9043) );
  XOR \SUBBYTES[3].a/U4632  ( .A(n9045), .B(n9044), .Z(\SUBBYTES[3].a/w2277 )
         );
  XOR \SUBBYTES[3].a/U4631  ( .A(n9047), .B(n9046), .Z(n9044) );
  XOR \SUBBYTES[3].a/U4630  ( .A(\w1[3][47] ), .B(\SUBBYTES[3].a/w2361 ), .Z(
        n9045) );
  XOR \SUBBYTES[3].a/U4629  ( .A(\SUBBYTES[3].a/w2268 ), .B(
        \SUBBYTES[3].a/w2271 ), .Z(n9046) );
  XOR \SUBBYTES[3].a/U4628  ( .A(\SUBBYTES[3].a/w2254 ), .B(
        \SUBBYTES[3].a/w2256 ), .Z(n9047) );
  XOR \SUBBYTES[3].a/U4627  ( .A(n9049), .B(n9048), .Z(\SUBBYTES[3].a/w2278 )
         );
  XOR \SUBBYTES[3].a/U4626  ( .A(n9584), .B(n9050), .Z(n9048) );
  XOR \SUBBYTES[3].a/U4625  ( .A(\w1[3][45] ), .B(n9585), .Z(n9049) );
  XOR \SUBBYTES[3].a/U4624  ( .A(\SUBBYTES[3].a/w2268 ), .B(
        \SUBBYTES[3].a/w2269 ), .Z(n9050) );
  XOR \SUBBYTES[3].a/U4623  ( .A(n9052), .B(n9051), .Z(\SUBBYTES[3].a/w2294 )
         );
  XOR \SUBBYTES[3].a/U4622  ( .A(\w1[3][41] ), .B(n9053), .Z(n9051) );
  XOR \SUBBYTES[3].a/U4621  ( .A(\SUBBYTES[3].a/w2269 ), .B(
        \SUBBYTES[3].a/w2271 ), .Z(n9052) );
  XOR \SUBBYTES[3].a/U4620  ( .A(\SUBBYTES[3].a/w2253 ), .B(
        \SUBBYTES[3].a/w2254 ), .Z(n9053) );
  XOR \SUBBYTES[3].a/U4619  ( .A(\w1[3][49] ), .B(n9054), .Z(n9586) );
  XOR \SUBBYTES[3].a/U4618  ( .A(\w1[3][51] ), .B(\w1[3][50] ), .Z(n9054) );
  XOR \SUBBYTES[3].a/U4617  ( .A(\w1[3][54] ), .B(n9586), .Z(
        \SUBBYTES[3].a/w2136 ) );
  XOR \SUBBYTES[3].a/U4616  ( .A(\w1[3][48] ), .B(\SUBBYTES[3].a/w2136 ), .Z(
        \SUBBYTES[3].a/w2023 ) );
  XOR \SUBBYTES[3].a/U4615  ( .A(\w1[3][48] ), .B(n9055), .Z(
        \SUBBYTES[3].a/w2024 ) );
  XOR \SUBBYTES[3].a/U4614  ( .A(\w1[3][54] ), .B(\w1[3][53] ), .Z(n9055) );
  XOR \SUBBYTES[3].a/U4613  ( .A(\w1[3][53] ), .B(n9586), .Z(
        \SUBBYTES[3].a/w2154 ) );
  XOR \SUBBYTES[3].a/U4612  ( .A(n9057), .B(n9056), .Z(\SUBBYTES[3].a/w2147 )
         );
  XOR \SUBBYTES[3].a/U4611  ( .A(\w1[3][51] ), .B(\w1[3][49] ), .Z(n9056) );
  XOR \SUBBYTES[3].a/U4610  ( .A(\w1[3][55] ), .B(\w1[3][52] ), .Z(n9057) );
  XOR \SUBBYTES[3].a/U4609  ( .A(\w1[3][48] ), .B(\SUBBYTES[3].a/w2147 ), .Z(
        \SUBBYTES[3].a/w2026 ) );
  XOR \SUBBYTES[3].a/U4608  ( .A(n9059), .B(n9058), .Z(\SUBBYTES[3].a/w2134 )
         );
  XOR \SUBBYTES[3].a/U4607  ( .A(\SUBBYTES[3].a/w2095 ), .B(n998), .Z(n9058)
         );
  XOR \SUBBYTES[3].a/U4606  ( .A(\SUBBYTES[3].a/w2088 ), .B(
        \SUBBYTES[3].a/w2091 ), .Z(n9059) );
  XOR \SUBBYTES[3].a/U4605  ( .A(n9061), .B(n9060), .Z(\SUBBYTES[3].a/w2135 )
         );
  XOR \SUBBYTES[3].a/U4604  ( .A(\SUBBYTES[3].a/w2095 ), .B(n8411), .Z(n9060)
         );
  XOR \SUBBYTES[3].a/U4603  ( .A(\SUBBYTES[3].a/w2088 ), .B(n8410), .Z(n9061)
         );
  XOR \SUBBYTES[3].a/U4602  ( .A(\SUBBYTES[3].a/w2147 ), .B(n9062), .Z(
        \SUBBYTES[3].a/w2137 ) );
  XOR \SUBBYTES[3].a/U4601  ( .A(\w1[3][54] ), .B(\w1[3][53] ), .Z(n9062) );
  XOR \SUBBYTES[3].a/U4600  ( .A(n9064), .B(n9063), .Z(\SUBBYTES[3].a/w2138 )
         );
  XOR \SUBBYTES[3].a/U4599  ( .A(n8411), .B(n998), .Z(n9063) );
  XOR \SUBBYTES[3].a/U4598  ( .A(n8410), .B(\SUBBYTES[3].a/w2091 ), .Z(n9064)
         );
  XOR \SUBBYTES[3].a/U4597  ( .A(\w1[3][55] ), .B(\w1[3][50] ), .Z(n9592) );
  XOR \SUBBYTES[3].a/U4596  ( .A(n9592), .B(n9065), .Z(\SUBBYTES[3].a/w2139 )
         );
  XOR \SUBBYTES[3].a/U4595  ( .A(\w1[3][53] ), .B(\w1[3][52] ), .Z(n9065) );
  XOR \SUBBYTES[3].a/U4594  ( .A(\w1[3][55] ), .B(\SUBBYTES[3].a/w2024 ), .Z(
        \SUBBYTES[3].a/w2027 ) );
  XOR \SUBBYTES[3].a/U4593  ( .A(\w1[3][49] ), .B(\SUBBYTES[3].a/w2024 ), .Z(
        \SUBBYTES[3].a/w2028 ) );
  XOR \SUBBYTES[3].a/U4592  ( .A(\w1[3][52] ), .B(\SUBBYTES[3].a/w2024 ), .Z(
        \SUBBYTES[3].a/w2029 ) );
  XOR \SUBBYTES[3].a/U4591  ( .A(\SUBBYTES[3].a/w2028 ), .B(n9592), .Z(
        \SUBBYTES[3].a/w2030 ) );
  XOR \SUBBYTES[3].a/U4590  ( .A(n9592), .B(n9066), .Z(\SUBBYTES[3].a/w2115 )
         );
  XOR \SUBBYTES[3].a/U4589  ( .A(\w1[3][52] ), .B(\w1[3][49] ), .Z(n9066) );
  XOR \SUBBYTES[3].a/U4588  ( .A(n9068), .B(n9067), .Z(n9589) );
  XOR \SUBBYTES[3].a/U4587  ( .A(\w1[3][52] ), .B(n9069), .Z(n9067) );
  XOR \SUBBYTES[3].a/U4586  ( .A(\SUBBYTES[3].a/w2080 ), .B(\w1[3][54] ), .Z(
        n9068) );
  XOR \SUBBYTES[3].a/U4585  ( .A(\SUBBYTES[3].a/w2054 ), .B(
        \SUBBYTES[3].a/w2061 ), .Z(n9069) );
  XOR \SUBBYTES[3].a/U4584  ( .A(n9071), .B(n9070), .Z(n9587) );
  XOR \SUBBYTES[3].a/U4583  ( .A(\w1[3][49] ), .B(n9072), .Z(n9070) );
  XOR \SUBBYTES[3].a/U4582  ( .A(\SUBBYTES[3].a/w2079 ), .B(\w1[3][53] ), .Z(
        n9071) );
  XOR \SUBBYTES[3].a/U4581  ( .A(\SUBBYTES[3].a/w2055 ), .B(
        \SUBBYTES[3].a/w2062 ), .Z(n9072) );
  XOR \SUBBYTES[3].a/U4580  ( .A(n9589), .B(n9587), .Z(\SUBBYTES[3].a/w2085 )
         );
  XOR \SUBBYTES[3].a/U4579  ( .A(\w1[3][53] ), .B(n9073), .Z(n9590) );
  XOR \SUBBYTES[3].a/U4578  ( .A(\SUBBYTES[3].a/w2047 ), .B(
        \SUBBYTES[3].a/w2057 ), .Z(n9073) );
  XOR \SUBBYTES[3].a/U4577  ( .A(n9075), .B(n9074), .Z(\SUBBYTES[3].a/w2072 )
         );
  XOR \SUBBYTES[3].a/U4576  ( .A(n9590), .B(n9076), .Z(n9074) );
  XOR \SUBBYTES[3].a/U4575  ( .A(\w1[3][52] ), .B(\SUBBYTES[3].a/w2136 ), .Z(
        n9075) );
  XOR \SUBBYTES[3].a/U4574  ( .A(\SUBBYTES[3].a/w2049 ), .B(
        \SUBBYTES[3].a/w2054 ), .Z(n9076) );
  XOR \SUBBYTES[3].a/U4573  ( .A(n9078), .B(n9077), .Z(n9588) );
  XOR \SUBBYTES[3].a/U4572  ( .A(\SUBBYTES[3].a/w2082 ), .B(\w1[3][55] ), .Z(
        n9077) );
  XOR \SUBBYTES[3].a/U4571  ( .A(\SUBBYTES[3].a/w2057 ), .B(
        \SUBBYTES[3].a/w2064 ), .Z(n9078) );
  XOR \SUBBYTES[3].a/U4570  ( .A(n9587), .B(n9588), .Z(\SUBBYTES[3].a/w2084 )
         );
  XOR \SUBBYTES[3].a/U4569  ( .A(\w1[3][51] ), .B(n9079), .Z(n9591) );
  XOR \SUBBYTES[3].a/U4568  ( .A(\SUBBYTES[3].a/w2046 ), .B(
        \SUBBYTES[3].a/w2049 ), .Z(n9079) );
  XOR \SUBBYTES[3].a/U4567  ( .A(n9081), .B(n9080), .Z(\SUBBYTES[3].a/w2073 )
         );
  XOR \SUBBYTES[3].a/U4566  ( .A(n9591), .B(n9082), .Z(n9080) );
  XOR \SUBBYTES[3].a/U4565  ( .A(\w1[3][54] ), .B(\SUBBYTES[3].a/w2115 ), .Z(
        n9081) );
  XOR \SUBBYTES[3].a/U4564  ( .A(\SUBBYTES[3].a/w2054 ), .B(
        \SUBBYTES[3].a/w2055 ), .Z(n9082) );
  XOR \SUBBYTES[3].a/U4563  ( .A(n9589), .B(n9588), .Z(\SUBBYTES[3].a/w2093 )
         );
  XOR \SUBBYTES[3].a/U4562  ( .A(n9084), .B(n9083), .Z(\SUBBYTES[3].a/w2094 )
         );
  XOR \SUBBYTES[3].a/U4561  ( .A(\w1[3][55] ), .B(n9590), .Z(n9083) );
  XOR \SUBBYTES[3].a/U4560  ( .A(\SUBBYTES[3].a/w2046 ), .B(
        \SUBBYTES[3].a/w2055 ), .Z(n9084) );
  XOR \SUBBYTES[3].a/U4559  ( .A(n9086), .B(n9085), .Z(\SUBBYTES[3].a/w2070 )
         );
  XOR \SUBBYTES[3].a/U4558  ( .A(n9088), .B(n9087), .Z(n9085) );
  XOR \SUBBYTES[3].a/U4557  ( .A(\w1[3][55] ), .B(\SUBBYTES[3].a/w2154 ), .Z(
        n9086) );
  XOR \SUBBYTES[3].a/U4556  ( .A(\SUBBYTES[3].a/w2061 ), .B(
        \SUBBYTES[3].a/w2064 ), .Z(n9087) );
  XOR \SUBBYTES[3].a/U4555  ( .A(\SUBBYTES[3].a/w2047 ), .B(
        \SUBBYTES[3].a/w2049 ), .Z(n9088) );
  XOR \SUBBYTES[3].a/U4554  ( .A(n9090), .B(n9089), .Z(\SUBBYTES[3].a/w2071 )
         );
  XOR \SUBBYTES[3].a/U4553  ( .A(n9591), .B(n9091), .Z(n9089) );
  XOR \SUBBYTES[3].a/U4552  ( .A(\w1[3][53] ), .B(n9592), .Z(n9090) );
  XOR \SUBBYTES[3].a/U4551  ( .A(\SUBBYTES[3].a/w2061 ), .B(
        \SUBBYTES[3].a/w2062 ), .Z(n9091) );
  XOR \SUBBYTES[3].a/U4550  ( .A(n9093), .B(n9092), .Z(\SUBBYTES[3].a/w2087 )
         );
  XOR \SUBBYTES[3].a/U4549  ( .A(\w1[3][49] ), .B(n9094), .Z(n9092) );
  XOR \SUBBYTES[3].a/U4548  ( .A(\SUBBYTES[3].a/w2062 ), .B(
        \SUBBYTES[3].a/w2064 ), .Z(n9093) );
  XOR \SUBBYTES[3].a/U4547  ( .A(\SUBBYTES[3].a/w2046 ), .B(
        \SUBBYTES[3].a/w2047 ), .Z(n9094) );
  XOR \SUBBYTES[3].a/U4546  ( .A(\w1[3][57] ), .B(n9095), .Z(n9593) );
  XOR \SUBBYTES[3].a/U4545  ( .A(\w1[3][59] ), .B(\w1[3][58] ), .Z(n9095) );
  XOR \SUBBYTES[3].a/U4544  ( .A(\w1[3][62] ), .B(n9593), .Z(
        \SUBBYTES[3].a/w1929 ) );
  XOR \SUBBYTES[3].a/U4543  ( .A(\w1[3][56] ), .B(\SUBBYTES[3].a/w1929 ), .Z(
        \SUBBYTES[3].a/w1816 ) );
  XOR \SUBBYTES[3].a/U4542  ( .A(\w1[3][56] ), .B(n9096), .Z(
        \SUBBYTES[3].a/w1817 ) );
  XOR \SUBBYTES[3].a/U4541  ( .A(\w1[3][62] ), .B(\w1[3][61] ), .Z(n9096) );
  XOR \SUBBYTES[3].a/U4540  ( .A(\w1[3][61] ), .B(n9593), .Z(
        \SUBBYTES[3].a/w1947 ) );
  XOR \SUBBYTES[3].a/U4539  ( .A(n9098), .B(n9097), .Z(\SUBBYTES[3].a/w1940 )
         );
  XOR \SUBBYTES[3].a/U4538  ( .A(\w1[3][59] ), .B(\w1[3][57] ), .Z(n9097) );
  XOR \SUBBYTES[3].a/U4537  ( .A(\w1[3][63] ), .B(\w1[3][60] ), .Z(n9098) );
  XOR \SUBBYTES[3].a/U4536  ( .A(\w1[3][56] ), .B(\SUBBYTES[3].a/w1940 ), .Z(
        \SUBBYTES[3].a/w1819 ) );
  XOR \SUBBYTES[3].a/U4535  ( .A(n9100), .B(n9099), .Z(\SUBBYTES[3].a/w1927 )
         );
  XOR \SUBBYTES[3].a/U4534  ( .A(\SUBBYTES[3].a/w1888 ), .B(n997), .Z(n9099)
         );
  XOR \SUBBYTES[3].a/U4533  ( .A(\SUBBYTES[3].a/w1881 ), .B(
        \SUBBYTES[3].a/w1884 ), .Z(n9100) );
  XOR \SUBBYTES[3].a/U4532  ( .A(n9102), .B(n9101), .Z(\SUBBYTES[3].a/w1928 )
         );
  XOR \SUBBYTES[3].a/U4531  ( .A(\SUBBYTES[3].a/w1888 ), .B(n8409), .Z(n9101)
         );
  XOR \SUBBYTES[3].a/U4530  ( .A(\SUBBYTES[3].a/w1881 ), .B(n8408), .Z(n9102)
         );
  XOR \SUBBYTES[3].a/U4529  ( .A(\SUBBYTES[3].a/w1940 ), .B(n9103), .Z(
        \SUBBYTES[3].a/w1930 ) );
  XOR \SUBBYTES[3].a/U4528  ( .A(\w1[3][62] ), .B(\w1[3][61] ), .Z(n9103) );
  XOR \SUBBYTES[3].a/U4527  ( .A(n9105), .B(n9104), .Z(\SUBBYTES[3].a/w1931 )
         );
  XOR \SUBBYTES[3].a/U4526  ( .A(n8409), .B(n997), .Z(n9104) );
  XOR \SUBBYTES[3].a/U4525  ( .A(n8408), .B(\SUBBYTES[3].a/w1884 ), .Z(n9105)
         );
  XOR \SUBBYTES[3].a/U4524  ( .A(\w1[3][63] ), .B(\w1[3][58] ), .Z(n9599) );
  XOR \SUBBYTES[3].a/U4523  ( .A(n9599), .B(n9106), .Z(\SUBBYTES[3].a/w1932 )
         );
  XOR \SUBBYTES[3].a/U4522  ( .A(\w1[3][61] ), .B(\w1[3][60] ), .Z(n9106) );
  XOR \SUBBYTES[3].a/U4521  ( .A(\w1[3][63] ), .B(\SUBBYTES[3].a/w1817 ), .Z(
        \SUBBYTES[3].a/w1820 ) );
  XOR \SUBBYTES[3].a/U4520  ( .A(\w1[3][57] ), .B(\SUBBYTES[3].a/w1817 ), .Z(
        \SUBBYTES[3].a/w1821 ) );
  XOR \SUBBYTES[3].a/U4519  ( .A(\w1[3][60] ), .B(\SUBBYTES[3].a/w1817 ), .Z(
        \SUBBYTES[3].a/w1822 ) );
  XOR \SUBBYTES[3].a/U4518  ( .A(\SUBBYTES[3].a/w1821 ), .B(n9599), .Z(
        \SUBBYTES[3].a/w1823 ) );
  XOR \SUBBYTES[3].a/U4517  ( .A(n9599), .B(n9107), .Z(\SUBBYTES[3].a/w1908 )
         );
  XOR \SUBBYTES[3].a/U4516  ( .A(\w1[3][60] ), .B(\w1[3][57] ), .Z(n9107) );
  XOR \SUBBYTES[3].a/U4515  ( .A(n9109), .B(n9108), .Z(n9596) );
  XOR \SUBBYTES[3].a/U4514  ( .A(\w1[3][60] ), .B(n9110), .Z(n9108) );
  XOR \SUBBYTES[3].a/U4513  ( .A(\SUBBYTES[3].a/w1873 ), .B(\w1[3][62] ), .Z(
        n9109) );
  XOR \SUBBYTES[3].a/U4512  ( .A(\SUBBYTES[3].a/w1847 ), .B(
        \SUBBYTES[3].a/w1854 ), .Z(n9110) );
  XOR \SUBBYTES[3].a/U4511  ( .A(n9112), .B(n9111), .Z(n9594) );
  XOR \SUBBYTES[3].a/U4510  ( .A(\w1[3][57] ), .B(n9113), .Z(n9111) );
  XOR \SUBBYTES[3].a/U4509  ( .A(\SUBBYTES[3].a/w1872 ), .B(\w1[3][61] ), .Z(
        n9112) );
  XOR \SUBBYTES[3].a/U4508  ( .A(\SUBBYTES[3].a/w1848 ), .B(
        \SUBBYTES[3].a/w1855 ), .Z(n9113) );
  XOR \SUBBYTES[3].a/U4507  ( .A(n9596), .B(n9594), .Z(\SUBBYTES[3].a/w1878 )
         );
  XOR \SUBBYTES[3].a/U4506  ( .A(\w1[3][61] ), .B(n9114), .Z(n9597) );
  XOR \SUBBYTES[3].a/U4505  ( .A(\SUBBYTES[3].a/w1840 ), .B(
        \SUBBYTES[3].a/w1850 ), .Z(n9114) );
  XOR \SUBBYTES[3].a/U4504  ( .A(n9116), .B(n9115), .Z(\SUBBYTES[3].a/w1865 )
         );
  XOR \SUBBYTES[3].a/U4503  ( .A(n9597), .B(n9117), .Z(n9115) );
  XOR \SUBBYTES[3].a/U4502  ( .A(\w1[3][60] ), .B(\SUBBYTES[3].a/w1929 ), .Z(
        n9116) );
  XOR \SUBBYTES[3].a/U4501  ( .A(\SUBBYTES[3].a/w1842 ), .B(
        \SUBBYTES[3].a/w1847 ), .Z(n9117) );
  XOR \SUBBYTES[3].a/U4500  ( .A(n9119), .B(n9118), .Z(n9595) );
  XOR \SUBBYTES[3].a/U4499  ( .A(\SUBBYTES[3].a/w1875 ), .B(\w1[3][63] ), .Z(
        n9118) );
  XOR \SUBBYTES[3].a/U4498  ( .A(\SUBBYTES[3].a/w1850 ), .B(
        \SUBBYTES[3].a/w1857 ), .Z(n9119) );
  XOR \SUBBYTES[3].a/U4497  ( .A(n9594), .B(n9595), .Z(\SUBBYTES[3].a/w1877 )
         );
  XOR \SUBBYTES[3].a/U4496  ( .A(\w1[3][59] ), .B(n9120), .Z(n9598) );
  XOR \SUBBYTES[3].a/U4495  ( .A(\SUBBYTES[3].a/w1839 ), .B(
        \SUBBYTES[3].a/w1842 ), .Z(n9120) );
  XOR \SUBBYTES[3].a/U4494  ( .A(n9122), .B(n9121), .Z(\SUBBYTES[3].a/w1866 )
         );
  XOR \SUBBYTES[3].a/U4493  ( .A(n9598), .B(n9123), .Z(n9121) );
  XOR \SUBBYTES[3].a/U4492  ( .A(\w1[3][62] ), .B(\SUBBYTES[3].a/w1908 ), .Z(
        n9122) );
  XOR \SUBBYTES[3].a/U4491  ( .A(\SUBBYTES[3].a/w1847 ), .B(
        \SUBBYTES[3].a/w1848 ), .Z(n9123) );
  XOR \SUBBYTES[3].a/U4490  ( .A(n9596), .B(n9595), .Z(\SUBBYTES[3].a/w1886 )
         );
  XOR \SUBBYTES[3].a/U4489  ( .A(n9125), .B(n9124), .Z(\SUBBYTES[3].a/w1887 )
         );
  XOR \SUBBYTES[3].a/U4488  ( .A(\w1[3][63] ), .B(n9597), .Z(n9124) );
  XOR \SUBBYTES[3].a/U4487  ( .A(\SUBBYTES[3].a/w1839 ), .B(
        \SUBBYTES[3].a/w1848 ), .Z(n9125) );
  XOR \SUBBYTES[3].a/U4486  ( .A(n9127), .B(n9126), .Z(\SUBBYTES[3].a/w1863 )
         );
  XOR \SUBBYTES[3].a/U4485  ( .A(n9129), .B(n9128), .Z(n9126) );
  XOR \SUBBYTES[3].a/U4484  ( .A(\w1[3][63] ), .B(\SUBBYTES[3].a/w1947 ), .Z(
        n9127) );
  XOR \SUBBYTES[3].a/U4483  ( .A(\SUBBYTES[3].a/w1854 ), .B(
        \SUBBYTES[3].a/w1857 ), .Z(n9128) );
  XOR \SUBBYTES[3].a/U4482  ( .A(\SUBBYTES[3].a/w1840 ), .B(
        \SUBBYTES[3].a/w1842 ), .Z(n9129) );
  XOR \SUBBYTES[3].a/U4481  ( .A(n9131), .B(n9130), .Z(\SUBBYTES[3].a/w1864 )
         );
  XOR \SUBBYTES[3].a/U4480  ( .A(n9598), .B(n9132), .Z(n9130) );
  XOR \SUBBYTES[3].a/U4479  ( .A(\w1[3][61] ), .B(n9599), .Z(n9131) );
  XOR \SUBBYTES[3].a/U4478  ( .A(\SUBBYTES[3].a/w1854 ), .B(
        \SUBBYTES[3].a/w1855 ), .Z(n9132) );
  XOR \SUBBYTES[3].a/U4477  ( .A(n9134), .B(n9133), .Z(\SUBBYTES[3].a/w1880 )
         );
  XOR \SUBBYTES[3].a/U4476  ( .A(\w1[3][57] ), .B(n9135), .Z(n9133) );
  XOR \SUBBYTES[3].a/U4475  ( .A(\SUBBYTES[3].a/w1855 ), .B(
        \SUBBYTES[3].a/w1857 ), .Z(n9134) );
  XOR \SUBBYTES[3].a/U4474  ( .A(\SUBBYTES[3].a/w1839 ), .B(
        \SUBBYTES[3].a/w1840 ), .Z(n9135) );
  XOR \SUBBYTES[3].a/U4473  ( .A(\w1[3][65] ), .B(n9136), .Z(n9600) );
  XOR \SUBBYTES[3].a/U4472  ( .A(\w1[3][67] ), .B(\w1[3][66] ), .Z(n9136) );
  XOR \SUBBYTES[3].a/U4471  ( .A(\w1[3][70] ), .B(n9600), .Z(
        \SUBBYTES[3].a/w1722 ) );
  XOR \SUBBYTES[3].a/U4470  ( .A(\w1[3][64] ), .B(\SUBBYTES[3].a/w1722 ), .Z(
        \SUBBYTES[3].a/w1609 ) );
  XOR \SUBBYTES[3].a/U4469  ( .A(\w1[3][64] ), .B(n9137), .Z(
        \SUBBYTES[3].a/w1610 ) );
  XOR \SUBBYTES[3].a/U4468  ( .A(\w1[3][70] ), .B(\w1[3][69] ), .Z(n9137) );
  XOR \SUBBYTES[3].a/U4467  ( .A(\w1[3][69] ), .B(n9600), .Z(
        \SUBBYTES[3].a/w1740 ) );
  XOR \SUBBYTES[3].a/U4466  ( .A(n9139), .B(n9138), .Z(\SUBBYTES[3].a/w1733 )
         );
  XOR \SUBBYTES[3].a/U4465  ( .A(\w1[3][67] ), .B(\w1[3][65] ), .Z(n9138) );
  XOR \SUBBYTES[3].a/U4464  ( .A(\w1[3][71] ), .B(\w1[3][68] ), .Z(n9139) );
  XOR \SUBBYTES[3].a/U4463  ( .A(\w1[3][64] ), .B(\SUBBYTES[3].a/w1733 ), .Z(
        \SUBBYTES[3].a/w1612 ) );
  XOR \SUBBYTES[3].a/U4462  ( .A(n9141), .B(n9140), .Z(\SUBBYTES[3].a/w1720 )
         );
  XOR \SUBBYTES[3].a/U4461  ( .A(\SUBBYTES[3].a/w1681 ), .B(n996), .Z(n9140)
         );
  XOR \SUBBYTES[3].a/U4460  ( .A(\SUBBYTES[3].a/w1674 ), .B(
        \SUBBYTES[3].a/w1677 ), .Z(n9141) );
  XOR \SUBBYTES[3].a/U4459  ( .A(n9143), .B(n9142), .Z(\SUBBYTES[3].a/w1721 )
         );
  XOR \SUBBYTES[3].a/U4458  ( .A(\SUBBYTES[3].a/w1681 ), .B(n8407), .Z(n9142)
         );
  XOR \SUBBYTES[3].a/U4457  ( .A(\SUBBYTES[3].a/w1674 ), .B(n8406), .Z(n9143)
         );
  XOR \SUBBYTES[3].a/U4456  ( .A(\SUBBYTES[3].a/w1733 ), .B(n9144), .Z(
        \SUBBYTES[3].a/w1723 ) );
  XOR \SUBBYTES[3].a/U4455  ( .A(\w1[3][70] ), .B(\w1[3][69] ), .Z(n9144) );
  XOR \SUBBYTES[3].a/U4454  ( .A(n9146), .B(n9145), .Z(\SUBBYTES[3].a/w1724 )
         );
  XOR \SUBBYTES[3].a/U4453  ( .A(n8407), .B(n996), .Z(n9145) );
  XOR \SUBBYTES[3].a/U4452  ( .A(n8406), .B(\SUBBYTES[3].a/w1677 ), .Z(n9146)
         );
  XOR \SUBBYTES[3].a/U4451  ( .A(\w1[3][71] ), .B(\w1[3][66] ), .Z(n9606) );
  XOR \SUBBYTES[3].a/U4450  ( .A(n9606), .B(n9147), .Z(\SUBBYTES[3].a/w1725 )
         );
  XOR \SUBBYTES[3].a/U4449  ( .A(\w1[3][69] ), .B(\w1[3][68] ), .Z(n9147) );
  XOR \SUBBYTES[3].a/U4448  ( .A(\w1[3][71] ), .B(\SUBBYTES[3].a/w1610 ), .Z(
        \SUBBYTES[3].a/w1613 ) );
  XOR \SUBBYTES[3].a/U4447  ( .A(\w1[3][65] ), .B(\SUBBYTES[3].a/w1610 ), .Z(
        \SUBBYTES[3].a/w1614 ) );
  XOR \SUBBYTES[3].a/U4446  ( .A(\w1[3][68] ), .B(\SUBBYTES[3].a/w1610 ), .Z(
        \SUBBYTES[3].a/w1615 ) );
  XOR \SUBBYTES[3].a/U4445  ( .A(\SUBBYTES[3].a/w1614 ), .B(n9606), .Z(
        \SUBBYTES[3].a/w1616 ) );
  XOR \SUBBYTES[3].a/U4444  ( .A(n9606), .B(n9148), .Z(\SUBBYTES[3].a/w1701 )
         );
  XOR \SUBBYTES[3].a/U4443  ( .A(\w1[3][68] ), .B(\w1[3][65] ), .Z(n9148) );
  XOR \SUBBYTES[3].a/U4442  ( .A(n9150), .B(n9149), .Z(n9603) );
  XOR \SUBBYTES[3].a/U4441  ( .A(\w1[3][68] ), .B(n9151), .Z(n9149) );
  XOR \SUBBYTES[3].a/U4440  ( .A(\SUBBYTES[3].a/w1666 ), .B(\w1[3][70] ), .Z(
        n9150) );
  XOR \SUBBYTES[3].a/U4439  ( .A(\SUBBYTES[3].a/w1640 ), .B(
        \SUBBYTES[3].a/w1647 ), .Z(n9151) );
  XOR \SUBBYTES[3].a/U4438  ( .A(n9153), .B(n9152), .Z(n9601) );
  XOR \SUBBYTES[3].a/U4437  ( .A(\w1[3][65] ), .B(n9154), .Z(n9152) );
  XOR \SUBBYTES[3].a/U4436  ( .A(\SUBBYTES[3].a/w1665 ), .B(\w1[3][69] ), .Z(
        n9153) );
  XOR \SUBBYTES[3].a/U4435  ( .A(\SUBBYTES[3].a/w1641 ), .B(
        \SUBBYTES[3].a/w1648 ), .Z(n9154) );
  XOR \SUBBYTES[3].a/U4434  ( .A(n9603), .B(n9601), .Z(\SUBBYTES[3].a/w1671 )
         );
  XOR \SUBBYTES[3].a/U4433  ( .A(\w1[3][69] ), .B(n9155), .Z(n9604) );
  XOR \SUBBYTES[3].a/U4432  ( .A(\SUBBYTES[3].a/w1633 ), .B(
        \SUBBYTES[3].a/w1643 ), .Z(n9155) );
  XOR \SUBBYTES[3].a/U4431  ( .A(n9157), .B(n9156), .Z(\SUBBYTES[3].a/w1658 )
         );
  XOR \SUBBYTES[3].a/U4430  ( .A(n9604), .B(n9158), .Z(n9156) );
  XOR \SUBBYTES[3].a/U4429  ( .A(\w1[3][68] ), .B(\SUBBYTES[3].a/w1722 ), .Z(
        n9157) );
  XOR \SUBBYTES[3].a/U4428  ( .A(\SUBBYTES[3].a/w1635 ), .B(
        \SUBBYTES[3].a/w1640 ), .Z(n9158) );
  XOR \SUBBYTES[3].a/U4427  ( .A(n9160), .B(n9159), .Z(n9602) );
  XOR \SUBBYTES[3].a/U4426  ( .A(\SUBBYTES[3].a/w1668 ), .B(\w1[3][71] ), .Z(
        n9159) );
  XOR \SUBBYTES[3].a/U4425  ( .A(\SUBBYTES[3].a/w1643 ), .B(
        \SUBBYTES[3].a/w1650 ), .Z(n9160) );
  XOR \SUBBYTES[3].a/U4424  ( .A(n9601), .B(n9602), .Z(\SUBBYTES[3].a/w1670 )
         );
  XOR \SUBBYTES[3].a/U4423  ( .A(\w1[3][67] ), .B(n9161), .Z(n9605) );
  XOR \SUBBYTES[3].a/U4422  ( .A(\SUBBYTES[3].a/w1632 ), .B(
        \SUBBYTES[3].a/w1635 ), .Z(n9161) );
  XOR \SUBBYTES[3].a/U4421  ( .A(n9163), .B(n9162), .Z(\SUBBYTES[3].a/w1659 )
         );
  XOR \SUBBYTES[3].a/U4420  ( .A(n9605), .B(n9164), .Z(n9162) );
  XOR \SUBBYTES[3].a/U4419  ( .A(\w1[3][70] ), .B(\SUBBYTES[3].a/w1701 ), .Z(
        n9163) );
  XOR \SUBBYTES[3].a/U4418  ( .A(\SUBBYTES[3].a/w1640 ), .B(
        \SUBBYTES[3].a/w1641 ), .Z(n9164) );
  XOR \SUBBYTES[3].a/U4417  ( .A(n9603), .B(n9602), .Z(\SUBBYTES[3].a/w1679 )
         );
  XOR \SUBBYTES[3].a/U4416  ( .A(n9166), .B(n9165), .Z(\SUBBYTES[3].a/w1680 )
         );
  XOR \SUBBYTES[3].a/U4415  ( .A(\w1[3][71] ), .B(n9604), .Z(n9165) );
  XOR \SUBBYTES[3].a/U4414  ( .A(\SUBBYTES[3].a/w1632 ), .B(
        \SUBBYTES[3].a/w1641 ), .Z(n9166) );
  XOR \SUBBYTES[3].a/U4413  ( .A(n9168), .B(n9167), .Z(\SUBBYTES[3].a/w1656 )
         );
  XOR \SUBBYTES[3].a/U4412  ( .A(n9170), .B(n9169), .Z(n9167) );
  XOR \SUBBYTES[3].a/U4411  ( .A(\w1[3][71] ), .B(\SUBBYTES[3].a/w1740 ), .Z(
        n9168) );
  XOR \SUBBYTES[3].a/U4410  ( .A(\SUBBYTES[3].a/w1647 ), .B(
        \SUBBYTES[3].a/w1650 ), .Z(n9169) );
  XOR \SUBBYTES[3].a/U4409  ( .A(\SUBBYTES[3].a/w1633 ), .B(
        \SUBBYTES[3].a/w1635 ), .Z(n9170) );
  XOR \SUBBYTES[3].a/U4408  ( .A(n9172), .B(n9171), .Z(\SUBBYTES[3].a/w1657 )
         );
  XOR \SUBBYTES[3].a/U4407  ( .A(n9605), .B(n9173), .Z(n9171) );
  XOR \SUBBYTES[3].a/U4406  ( .A(\w1[3][69] ), .B(n9606), .Z(n9172) );
  XOR \SUBBYTES[3].a/U4405  ( .A(\SUBBYTES[3].a/w1647 ), .B(
        \SUBBYTES[3].a/w1648 ), .Z(n9173) );
  XOR \SUBBYTES[3].a/U4404  ( .A(n9175), .B(n9174), .Z(\SUBBYTES[3].a/w1673 )
         );
  XOR \SUBBYTES[3].a/U4403  ( .A(\w1[3][65] ), .B(n9176), .Z(n9174) );
  XOR \SUBBYTES[3].a/U4402  ( .A(\SUBBYTES[3].a/w1648 ), .B(
        \SUBBYTES[3].a/w1650 ), .Z(n9175) );
  XOR \SUBBYTES[3].a/U4401  ( .A(\SUBBYTES[3].a/w1632 ), .B(
        \SUBBYTES[3].a/w1633 ), .Z(n9176) );
  XOR \SUBBYTES[3].a/U4400  ( .A(\w1[3][73] ), .B(n9177), .Z(n9607) );
  XOR \SUBBYTES[3].a/U4399  ( .A(\w1[3][75] ), .B(\w1[3][74] ), .Z(n9177) );
  XOR \SUBBYTES[3].a/U4398  ( .A(\w1[3][78] ), .B(n9607), .Z(
        \SUBBYTES[3].a/w1515 ) );
  XOR \SUBBYTES[3].a/U4397  ( .A(\w1[3][72] ), .B(\SUBBYTES[3].a/w1515 ), .Z(
        \SUBBYTES[3].a/w1402 ) );
  XOR \SUBBYTES[3].a/U4396  ( .A(\w1[3][72] ), .B(n9178), .Z(
        \SUBBYTES[3].a/w1403 ) );
  XOR \SUBBYTES[3].a/U4395  ( .A(\w1[3][78] ), .B(\w1[3][77] ), .Z(n9178) );
  XOR \SUBBYTES[3].a/U4394  ( .A(\w1[3][77] ), .B(n9607), .Z(
        \SUBBYTES[3].a/w1533 ) );
  XOR \SUBBYTES[3].a/U4393  ( .A(n9180), .B(n9179), .Z(\SUBBYTES[3].a/w1526 )
         );
  XOR \SUBBYTES[3].a/U4392  ( .A(\w1[3][75] ), .B(\w1[3][73] ), .Z(n9179) );
  XOR \SUBBYTES[3].a/U4391  ( .A(\w1[3][79] ), .B(\w1[3][76] ), .Z(n9180) );
  XOR \SUBBYTES[3].a/U4390  ( .A(\w1[3][72] ), .B(\SUBBYTES[3].a/w1526 ), .Z(
        \SUBBYTES[3].a/w1405 ) );
  XOR \SUBBYTES[3].a/U4389  ( .A(n9182), .B(n9181), .Z(\SUBBYTES[3].a/w1513 )
         );
  XOR \SUBBYTES[3].a/U4388  ( .A(\SUBBYTES[3].a/w1474 ), .B(n995), .Z(n9181)
         );
  XOR \SUBBYTES[3].a/U4387  ( .A(\SUBBYTES[3].a/w1467 ), .B(
        \SUBBYTES[3].a/w1470 ), .Z(n9182) );
  XOR \SUBBYTES[3].a/U4386  ( .A(n9184), .B(n9183), .Z(\SUBBYTES[3].a/w1514 )
         );
  XOR \SUBBYTES[3].a/U4385  ( .A(\SUBBYTES[3].a/w1474 ), .B(n8405), .Z(n9183)
         );
  XOR \SUBBYTES[3].a/U4384  ( .A(\SUBBYTES[3].a/w1467 ), .B(n8404), .Z(n9184)
         );
  XOR \SUBBYTES[3].a/U4383  ( .A(\SUBBYTES[3].a/w1526 ), .B(n9185), .Z(
        \SUBBYTES[3].a/w1516 ) );
  XOR \SUBBYTES[3].a/U4382  ( .A(\w1[3][78] ), .B(\w1[3][77] ), .Z(n9185) );
  XOR \SUBBYTES[3].a/U4381  ( .A(n9187), .B(n9186), .Z(\SUBBYTES[3].a/w1517 )
         );
  XOR \SUBBYTES[3].a/U4380  ( .A(n8405), .B(n995), .Z(n9186) );
  XOR \SUBBYTES[3].a/U4379  ( .A(n8404), .B(\SUBBYTES[3].a/w1470 ), .Z(n9187)
         );
  XOR \SUBBYTES[3].a/U4378  ( .A(\w1[3][79] ), .B(\w1[3][74] ), .Z(n9613) );
  XOR \SUBBYTES[3].a/U4377  ( .A(n9613), .B(n9188), .Z(\SUBBYTES[3].a/w1518 )
         );
  XOR \SUBBYTES[3].a/U4376  ( .A(\w1[3][77] ), .B(\w1[3][76] ), .Z(n9188) );
  XOR \SUBBYTES[3].a/U4375  ( .A(\w1[3][79] ), .B(\SUBBYTES[3].a/w1403 ), .Z(
        \SUBBYTES[3].a/w1406 ) );
  XOR \SUBBYTES[3].a/U4374  ( .A(\w1[3][73] ), .B(\SUBBYTES[3].a/w1403 ), .Z(
        \SUBBYTES[3].a/w1407 ) );
  XOR \SUBBYTES[3].a/U4373  ( .A(\w1[3][76] ), .B(\SUBBYTES[3].a/w1403 ), .Z(
        \SUBBYTES[3].a/w1408 ) );
  XOR \SUBBYTES[3].a/U4372  ( .A(\SUBBYTES[3].a/w1407 ), .B(n9613), .Z(
        \SUBBYTES[3].a/w1409 ) );
  XOR \SUBBYTES[3].a/U4371  ( .A(n9613), .B(n9189), .Z(\SUBBYTES[3].a/w1494 )
         );
  XOR \SUBBYTES[3].a/U4370  ( .A(\w1[3][76] ), .B(\w1[3][73] ), .Z(n9189) );
  XOR \SUBBYTES[3].a/U4369  ( .A(n9191), .B(n9190), .Z(n9610) );
  XOR \SUBBYTES[3].a/U4368  ( .A(\w1[3][76] ), .B(n9192), .Z(n9190) );
  XOR \SUBBYTES[3].a/U4367  ( .A(\SUBBYTES[3].a/w1459 ), .B(\w1[3][78] ), .Z(
        n9191) );
  XOR \SUBBYTES[3].a/U4366  ( .A(\SUBBYTES[3].a/w1433 ), .B(
        \SUBBYTES[3].a/w1440 ), .Z(n9192) );
  XOR \SUBBYTES[3].a/U4365  ( .A(n9194), .B(n9193), .Z(n9608) );
  XOR \SUBBYTES[3].a/U4364  ( .A(\w1[3][73] ), .B(n9195), .Z(n9193) );
  XOR \SUBBYTES[3].a/U4363  ( .A(\SUBBYTES[3].a/w1458 ), .B(\w1[3][77] ), .Z(
        n9194) );
  XOR \SUBBYTES[3].a/U4362  ( .A(\SUBBYTES[3].a/w1434 ), .B(
        \SUBBYTES[3].a/w1441 ), .Z(n9195) );
  XOR \SUBBYTES[3].a/U4361  ( .A(n9610), .B(n9608), .Z(\SUBBYTES[3].a/w1464 )
         );
  XOR \SUBBYTES[3].a/U4360  ( .A(\w1[3][77] ), .B(n9196), .Z(n9611) );
  XOR \SUBBYTES[3].a/U4359  ( .A(\SUBBYTES[3].a/w1426 ), .B(
        \SUBBYTES[3].a/w1436 ), .Z(n9196) );
  XOR \SUBBYTES[3].a/U4358  ( .A(n9198), .B(n9197), .Z(\SUBBYTES[3].a/w1451 )
         );
  XOR \SUBBYTES[3].a/U4357  ( .A(n9611), .B(n9199), .Z(n9197) );
  XOR \SUBBYTES[3].a/U4356  ( .A(\w1[3][76] ), .B(\SUBBYTES[3].a/w1515 ), .Z(
        n9198) );
  XOR \SUBBYTES[3].a/U4355  ( .A(\SUBBYTES[3].a/w1428 ), .B(
        \SUBBYTES[3].a/w1433 ), .Z(n9199) );
  XOR \SUBBYTES[3].a/U4354  ( .A(n9201), .B(n9200), .Z(n9609) );
  XOR \SUBBYTES[3].a/U4353  ( .A(\SUBBYTES[3].a/w1461 ), .B(\w1[3][79] ), .Z(
        n9200) );
  XOR \SUBBYTES[3].a/U4352  ( .A(\SUBBYTES[3].a/w1436 ), .B(
        \SUBBYTES[3].a/w1443 ), .Z(n9201) );
  XOR \SUBBYTES[3].a/U4351  ( .A(n9608), .B(n9609), .Z(\SUBBYTES[3].a/w1463 )
         );
  XOR \SUBBYTES[3].a/U4350  ( .A(\w1[3][75] ), .B(n9202), .Z(n9612) );
  XOR \SUBBYTES[3].a/U4349  ( .A(\SUBBYTES[3].a/w1425 ), .B(
        \SUBBYTES[3].a/w1428 ), .Z(n9202) );
  XOR \SUBBYTES[3].a/U4348  ( .A(n9204), .B(n9203), .Z(\SUBBYTES[3].a/w1452 )
         );
  XOR \SUBBYTES[3].a/U4347  ( .A(n9612), .B(n9205), .Z(n9203) );
  XOR \SUBBYTES[3].a/U4346  ( .A(\w1[3][78] ), .B(\SUBBYTES[3].a/w1494 ), .Z(
        n9204) );
  XOR \SUBBYTES[3].a/U4345  ( .A(\SUBBYTES[3].a/w1433 ), .B(
        \SUBBYTES[3].a/w1434 ), .Z(n9205) );
  XOR \SUBBYTES[3].a/U4344  ( .A(n9610), .B(n9609), .Z(\SUBBYTES[3].a/w1472 )
         );
  XOR \SUBBYTES[3].a/U4343  ( .A(n9207), .B(n9206), .Z(\SUBBYTES[3].a/w1473 )
         );
  XOR \SUBBYTES[3].a/U4342  ( .A(\w1[3][79] ), .B(n9611), .Z(n9206) );
  XOR \SUBBYTES[3].a/U4341  ( .A(\SUBBYTES[3].a/w1425 ), .B(
        \SUBBYTES[3].a/w1434 ), .Z(n9207) );
  XOR \SUBBYTES[3].a/U4340  ( .A(n9209), .B(n9208), .Z(\SUBBYTES[3].a/w1449 )
         );
  XOR \SUBBYTES[3].a/U4339  ( .A(n9211), .B(n9210), .Z(n9208) );
  XOR \SUBBYTES[3].a/U4338  ( .A(\w1[3][79] ), .B(\SUBBYTES[3].a/w1533 ), .Z(
        n9209) );
  XOR \SUBBYTES[3].a/U4337  ( .A(\SUBBYTES[3].a/w1440 ), .B(
        \SUBBYTES[3].a/w1443 ), .Z(n9210) );
  XOR \SUBBYTES[3].a/U4336  ( .A(\SUBBYTES[3].a/w1426 ), .B(
        \SUBBYTES[3].a/w1428 ), .Z(n9211) );
  XOR \SUBBYTES[3].a/U4335  ( .A(n9213), .B(n9212), .Z(\SUBBYTES[3].a/w1450 )
         );
  XOR \SUBBYTES[3].a/U4334  ( .A(n9612), .B(n9214), .Z(n9212) );
  XOR \SUBBYTES[3].a/U4333  ( .A(\w1[3][77] ), .B(n9613), .Z(n9213) );
  XOR \SUBBYTES[3].a/U4332  ( .A(\SUBBYTES[3].a/w1440 ), .B(
        \SUBBYTES[3].a/w1441 ), .Z(n9214) );
  XOR \SUBBYTES[3].a/U4331  ( .A(n9216), .B(n9215), .Z(\SUBBYTES[3].a/w1466 )
         );
  XOR \SUBBYTES[3].a/U4330  ( .A(\w1[3][73] ), .B(n9217), .Z(n9215) );
  XOR \SUBBYTES[3].a/U4329  ( .A(\SUBBYTES[3].a/w1441 ), .B(
        \SUBBYTES[3].a/w1443 ), .Z(n9216) );
  XOR \SUBBYTES[3].a/U4328  ( .A(\SUBBYTES[3].a/w1425 ), .B(
        \SUBBYTES[3].a/w1426 ), .Z(n9217) );
  XOR \SUBBYTES[3].a/U4327  ( .A(\w1[3][81] ), .B(n9218), .Z(n9614) );
  XOR \SUBBYTES[3].a/U4326  ( .A(\w1[3][83] ), .B(\w1[3][82] ), .Z(n9218) );
  XOR \SUBBYTES[3].a/U4325  ( .A(\w1[3][86] ), .B(n9614), .Z(
        \SUBBYTES[3].a/w1308 ) );
  XOR \SUBBYTES[3].a/U4324  ( .A(\w1[3][80] ), .B(\SUBBYTES[3].a/w1308 ), .Z(
        \SUBBYTES[3].a/w1195 ) );
  XOR \SUBBYTES[3].a/U4323  ( .A(\w1[3][80] ), .B(n9219), .Z(
        \SUBBYTES[3].a/w1196 ) );
  XOR \SUBBYTES[3].a/U4322  ( .A(\w1[3][86] ), .B(\w1[3][85] ), .Z(n9219) );
  XOR \SUBBYTES[3].a/U4321  ( .A(\w1[3][85] ), .B(n9614), .Z(
        \SUBBYTES[3].a/w1326 ) );
  XOR \SUBBYTES[3].a/U4320  ( .A(n9221), .B(n9220), .Z(\SUBBYTES[3].a/w1319 )
         );
  XOR \SUBBYTES[3].a/U4319  ( .A(\w1[3][83] ), .B(\w1[3][81] ), .Z(n9220) );
  XOR \SUBBYTES[3].a/U4318  ( .A(\w1[3][87] ), .B(\w1[3][84] ), .Z(n9221) );
  XOR \SUBBYTES[3].a/U4317  ( .A(\w1[3][80] ), .B(\SUBBYTES[3].a/w1319 ), .Z(
        \SUBBYTES[3].a/w1198 ) );
  XOR \SUBBYTES[3].a/U4316  ( .A(n9223), .B(n9222), .Z(\SUBBYTES[3].a/w1306 )
         );
  XOR \SUBBYTES[3].a/U4315  ( .A(\SUBBYTES[3].a/w1267 ), .B(n994), .Z(n9222)
         );
  XOR \SUBBYTES[3].a/U4314  ( .A(\SUBBYTES[3].a/w1260 ), .B(
        \SUBBYTES[3].a/w1263 ), .Z(n9223) );
  XOR \SUBBYTES[3].a/U4313  ( .A(n9225), .B(n9224), .Z(\SUBBYTES[3].a/w1307 )
         );
  XOR \SUBBYTES[3].a/U4312  ( .A(\SUBBYTES[3].a/w1267 ), .B(n8403), .Z(n9224)
         );
  XOR \SUBBYTES[3].a/U4311  ( .A(\SUBBYTES[3].a/w1260 ), .B(n8402), .Z(n9225)
         );
  XOR \SUBBYTES[3].a/U4310  ( .A(\SUBBYTES[3].a/w1319 ), .B(n9226), .Z(
        \SUBBYTES[3].a/w1309 ) );
  XOR \SUBBYTES[3].a/U4309  ( .A(\w1[3][86] ), .B(\w1[3][85] ), .Z(n9226) );
  XOR \SUBBYTES[3].a/U4308  ( .A(n9228), .B(n9227), .Z(\SUBBYTES[3].a/w1310 )
         );
  XOR \SUBBYTES[3].a/U4307  ( .A(n8403), .B(n994), .Z(n9227) );
  XOR \SUBBYTES[3].a/U4306  ( .A(n8402), .B(\SUBBYTES[3].a/w1263 ), .Z(n9228)
         );
  XOR \SUBBYTES[3].a/U4305  ( .A(\w1[3][87] ), .B(\w1[3][82] ), .Z(n9620) );
  XOR \SUBBYTES[3].a/U4304  ( .A(n9620), .B(n9229), .Z(\SUBBYTES[3].a/w1311 )
         );
  XOR \SUBBYTES[3].a/U4303  ( .A(\w1[3][85] ), .B(\w1[3][84] ), .Z(n9229) );
  XOR \SUBBYTES[3].a/U4302  ( .A(\w1[3][87] ), .B(\SUBBYTES[3].a/w1196 ), .Z(
        \SUBBYTES[3].a/w1199 ) );
  XOR \SUBBYTES[3].a/U4301  ( .A(\w1[3][81] ), .B(\SUBBYTES[3].a/w1196 ), .Z(
        \SUBBYTES[3].a/w1200 ) );
  XOR \SUBBYTES[3].a/U4300  ( .A(\w1[3][84] ), .B(\SUBBYTES[3].a/w1196 ), .Z(
        \SUBBYTES[3].a/w1201 ) );
  XOR \SUBBYTES[3].a/U4299  ( .A(\SUBBYTES[3].a/w1200 ), .B(n9620), .Z(
        \SUBBYTES[3].a/w1202 ) );
  XOR \SUBBYTES[3].a/U4298  ( .A(n9620), .B(n9230), .Z(\SUBBYTES[3].a/w1287 )
         );
  XOR \SUBBYTES[3].a/U4297  ( .A(\w1[3][84] ), .B(\w1[3][81] ), .Z(n9230) );
  XOR \SUBBYTES[3].a/U4296  ( .A(n9232), .B(n9231), .Z(n9617) );
  XOR \SUBBYTES[3].a/U4295  ( .A(\w1[3][84] ), .B(n9233), .Z(n9231) );
  XOR \SUBBYTES[3].a/U4294  ( .A(\SUBBYTES[3].a/w1252 ), .B(\w1[3][86] ), .Z(
        n9232) );
  XOR \SUBBYTES[3].a/U4293  ( .A(\SUBBYTES[3].a/w1226 ), .B(
        \SUBBYTES[3].a/w1233 ), .Z(n9233) );
  XOR \SUBBYTES[3].a/U4292  ( .A(n9235), .B(n9234), .Z(n9615) );
  XOR \SUBBYTES[3].a/U4291  ( .A(\w1[3][81] ), .B(n9236), .Z(n9234) );
  XOR \SUBBYTES[3].a/U4290  ( .A(\SUBBYTES[3].a/w1251 ), .B(\w1[3][85] ), .Z(
        n9235) );
  XOR \SUBBYTES[3].a/U4289  ( .A(\SUBBYTES[3].a/w1227 ), .B(
        \SUBBYTES[3].a/w1234 ), .Z(n9236) );
  XOR \SUBBYTES[3].a/U4288  ( .A(n9617), .B(n9615), .Z(\SUBBYTES[3].a/w1257 )
         );
  XOR \SUBBYTES[3].a/U4287  ( .A(\w1[3][85] ), .B(n9237), .Z(n9618) );
  XOR \SUBBYTES[3].a/U4286  ( .A(\SUBBYTES[3].a/w1219 ), .B(
        \SUBBYTES[3].a/w1229 ), .Z(n9237) );
  XOR \SUBBYTES[3].a/U4285  ( .A(n9239), .B(n9238), .Z(\SUBBYTES[3].a/w1244 )
         );
  XOR \SUBBYTES[3].a/U4284  ( .A(n9618), .B(n9240), .Z(n9238) );
  XOR \SUBBYTES[3].a/U4283  ( .A(\w1[3][84] ), .B(\SUBBYTES[3].a/w1308 ), .Z(
        n9239) );
  XOR \SUBBYTES[3].a/U4282  ( .A(\SUBBYTES[3].a/w1221 ), .B(
        \SUBBYTES[3].a/w1226 ), .Z(n9240) );
  XOR \SUBBYTES[3].a/U4281  ( .A(n9242), .B(n9241), .Z(n9616) );
  XOR \SUBBYTES[3].a/U4280  ( .A(\SUBBYTES[3].a/w1254 ), .B(\w1[3][87] ), .Z(
        n9241) );
  XOR \SUBBYTES[3].a/U4279  ( .A(\SUBBYTES[3].a/w1229 ), .B(
        \SUBBYTES[3].a/w1236 ), .Z(n9242) );
  XOR \SUBBYTES[3].a/U4278  ( .A(n9615), .B(n9616), .Z(\SUBBYTES[3].a/w1256 )
         );
  XOR \SUBBYTES[3].a/U4277  ( .A(\w1[3][83] ), .B(n9243), .Z(n9619) );
  XOR \SUBBYTES[3].a/U4276  ( .A(\SUBBYTES[3].a/w1218 ), .B(
        \SUBBYTES[3].a/w1221 ), .Z(n9243) );
  XOR \SUBBYTES[3].a/U4275  ( .A(n9245), .B(n9244), .Z(\SUBBYTES[3].a/w1245 )
         );
  XOR \SUBBYTES[3].a/U4274  ( .A(n9619), .B(n9246), .Z(n9244) );
  XOR \SUBBYTES[3].a/U4273  ( .A(\w1[3][86] ), .B(\SUBBYTES[3].a/w1287 ), .Z(
        n9245) );
  XOR \SUBBYTES[3].a/U4272  ( .A(\SUBBYTES[3].a/w1226 ), .B(
        \SUBBYTES[3].a/w1227 ), .Z(n9246) );
  XOR \SUBBYTES[3].a/U4271  ( .A(n9617), .B(n9616), .Z(\SUBBYTES[3].a/w1265 )
         );
  XOR \SUBBYTES[3].a/U4270  ( .A(n9248), .B(n9247), .Z(\SUBBYTES[3].a/w1266 )
         );
  XOR \SUBBYTES[3].a/U4269  ( .A(\w1[3][87] ), .B(n9618), .Z(n9247) );
  XOR \SUBBYTES[3].a/U4268  ( .A(\SUBBYTES[3].a/w1218 ), .B(
        \SUBBYTES[3].a/w1227 ), .Z(n9248) );
  XOR \SUBBYTES[3].a/U4267  ( .A(n9250), .B(n9249), .Z(\SUBBYTES[3].a/w1242 )
         );
  XOR \SUBBYTES[3].a/U4266  ( .A(n9252), .B(n9251), .Z(n9249) );
  XOR \SUBBYTES[3].a/U4265  ( .A(\w1[3][87] ), .B(\SUBBYTES[3].a/w1326 ), .Z(
        n9250) );
  XOR \SUBBYTES[3].a/U4264  ( .A(\SUBBYTES[3].a/w1233 ), .B(
        \SUBBYTES[3].a/w1236 ), .Z(n9251) );
  XOR \SUBBYTES[3].a/U4263  ( .A(\SUBBYTES[3].a/w1219 ), .B(
        \SUBBYTES[3].a/w1221 ), .Z(n9252) );
  XOR \SUBBYTES[3].a/U4262  ( .A(n9254), .B(n9253), .Z(\SUBBYTES[3].a/w1243 )
         );
  XOR \SUBBYTES[3].a/U4261  ( .A(n9619), .B(n9255), .Z(n9253) );
  XOR \SUBBYTES[3].a/U4260  ( .A(\w1[3][85] ), .B(n9620), .Z(n9254) );
  XOR \SUBBYTES[3].a/U4259  ( .A(\SUBBYTES[3].a/w1233 ), .B(
        \SUBBYTES[3].a/w1234 ), .Z(n9255) );
  XOR \SUBBYTES[3].a/U4258  ( .A(n9257), .B(n9256), .Z(\SUBBYTES[3].a/w1259 )
         );
  XOR \SUBBYTES[3].a/U4257  ( .A(\w1[3][81] ), .B(n9258), .Z(n9256) );
  XOR \SUBBYTES[3].a/U4256  ( .A(\SUBBYTES[3].a/w1234 ), .B(
        \SUBBYTES[3].a/w1236 ), .Z(n9257) );
  XOR \SUBBYTES[3].a/U4255  ( .A(\SUBBYTES[3].a/w1218 ), .B(
        \SUBBYTES[3].a/w1219 ), .Z(n9258) );
  XOR \SUBBYTES[3].a/U4254  ( .A(\w1[3][89] ), .B(n9259), .Z(n9621) );
  XOR \SUBBYTES[3].a/U4253  ( .A(\w1[3][91] ), .B(\w1[3][90] ), .Z(n9259) );
  XOR \SUBBYTES[3].a/U4252  ( .A(\w1[3][94] ), .B(n9621), .Z(
        \SUBBYTES[3].a/w1101 ) );
  XOR \SUBBYTES[3].a/U4251  ( .A(\w1[3][88] ), .B(\SUBBYTES[3].a/w1101 ), .Z(
        \SUBBYTES[3].a/w988 ) );
  XOR \SUBBYTES[3].a/U4250  ( .A(\w1[3][88] ), .B(n9260), .Z(
        \SUBBYTES[3].a/w989 ) );
  XOR \SUBBYTES[3].a/U4249  ( .A(\w1[3][94] ), .B(\w1[3][93] ), .Z(n9260) );
  XOR \SUBBYTES[3].a/U4248  ( .A(\w1[3][93] ), .B(n9621), .Z(
        \SUBBYTES[3].a/w1119 ) );
  XOR \SUBBYTES[3].a/U4247  ( .A(n9262), .B(n9261), .Z(\SUBBYTES[3].a/w1112 )
         );
  XOR \SUBBYTES[3].a/U4246  ( .A(\w1[3][91] ), .B(\w1[3][89] ), .Z(n9261) );
  XOR \SUBBYTES[3].a/U4245  ( .A(\w1[3][95] ), .B(\w1[3][92] ), .Z(n9262) );
  XOR \SUBBYTES[3].a/U4244  ( .A(\w1[3][88] ), .B(\SUBBYTES[3].a/w1112 ), .Z(
        \SUBBYTES[3].a/w991 ) );
  XOR \SUBBYTES[3].a/U4243  ( .A(n9264), .B(n9263), .Z(\SUBBYTES[3].a/w1099 )
         );
  XOR \SUBBYTES[3].a/U4242  ( .A(\SUBBYTES[3].a/w1060 ), .B(n993), .Z(n9263)
         );
  XOR \SUBBYTES[3].a/U4241  ( .A(\SUBBYTES[3].a/w1053 ), .B(
        \SUBBYTES[3].a/w1056 ), .Z(n9264) );
  XOR \SUBBYTES[3].a/U4240  ( .A(n9266), .B(n9265), .Z(\SUBBYTES[3].a/w1100 )
         );
  XOR \SUBBYTES[3].a/U4239  ( .A(\SUBBYTES[3].a/w1060 ), .B(n8401), .Z(n9265)
         );
  XOR \SUBBYTES[3].a/U4238  ( .A(\SUBBYTES[3].a/w1053 ), .B(n8400), .Z(n9266)
         );
  XOR \SUBBYTES[3].a/U4237  ( .A(\SUBBYTES[3].a/w1112 ), .B(n9267), .Z(
        \SUBBYTES[3].a/w1102 ) );
  XOR \SUBBYTES[3].a/U4236  ( .A(\w1[3][94] ), .B(\w1[3][93] ), .Z(n9267) );
  XOR \SUBBYTES[3].a/U4235  ( .A(n9269), .B(n9268), .Z(\SUBBYTES[3].a/w1103 )
         );
  XOR \SUBBYTES[3].a/U4234  ( .A(n8401), .B(n993), .Z(n9268) );
  XOR \SUBBYTES[3].a/U4233  ( .A(n8400), .B(\SUBBYTES[3].a/w1056 ), .Z(n9269)
         );
  XOR \SUBBYTES[3].a/U4232  ( .A(\w1[3][95] ), .B(\w1[3][90] ), .Z(n9627) );
  XOR \SUBBYTES[3].a/U4231  ( .A(n9627), .B(n9270), .Z(\SUBBYTES[3].a/w1104 )
         );
  XOR \SUBBYTES[3].a/U4230  ( .A(\w1[3][93] ), .B(\w1[3][92] ), .Z(n9270) );
  XOR \SUBBYTES[3].a/U4229  ( .A(\w1[3][95] ), .B(\SUBBYTES[3].a/w989 ), .Z(
        \SUBBYTES[3].a/w992 ) );
  XOR \SUBBYTES[3].a/U4228  ( .A(\w1[3][89] ), .B(\SUBBYTES[3].a/w989 ), .Z(
        \SUBBYTES[3].a/w993 ) );
  XOR \SUBBYTES[3].a/U4227  ( .A(\w1[3][92] ), .B(\SUBBYTES[3].a/w989 ), .Z(
        \SUBBYTES[3].a/w994 ) );
  XOR \SUBBYTES[3].a/U4226  ( .A(\SUBBYTES[3].a/w993 ), .B(n9627), .Z(
        \SUBBYTES[3].a/w995 ) );
  XOR \SUBBYTES[3].a/U4225  ( .A(n9627), .B(n9271), .Z(\SUBBYTES[3].a/w1080 )
         );
  XOR \SUBBYTES[3].a/U4224  ( .A(\w1[3][92] ), .B(\w1[3][89] ), .Z(n9271) );
  XOR \SUBBYTES[3].a/U4223  ( .A(n9273), .B(n9272), .Z(n9624) );
  XOR \SUBBYTES[3].a/U4222  ( .A(\w1[3][92] ), .B(n9274), .Z(n9272) );
  XOR \SUBBYTES[3].a/U4221  ( .A(\SUBBYTES[3].a/w1045 ), .B(\w1[3][94] ), .Z(
        n9273) );
  XOR \SUBBYTES[3].a/U4220  ( .A(\SUBBYTES[3].a/w1019 ), .B(
        \SUBBYTES[3].a/w1026 ), .Z(n9274) );
  XOR \SUBBYTES[3].a/U4219  ( .A(n9276), .B(n9275), .Z(n9622) );
  XOR \SUBBYTES[3].a/U4218  ( .A(\w1[3][89] ), .B(n9277), .Z(n9275) );
  XOR \SUBBYTES[3].a/U4217  ( .A(\SUBBYTES[3].a/w1044 ), .B(\w1[3][93] ), .Z(
        n9276) );
  XOR \SUBBYTES[3].a/U4216  ( .A(\SUBBYTES[3].a/w1020 ), .B(
        \SUBBYTES[3].a/w1027 ), .Z(n9277) );
  XOR \SUBBYTES[3].a/U4215  ( .A(n9624), .B(n9622), .Z(\SUBBYTES[3].a/w1050 )
         );
  XOR \SUBBYTES[3].a/U4214  ( .A(\w1[3][93] ), .B(n9278), .Z(n9625) );
  XOR \SUBBYTES[3].a/U4213  ( .A(\SUBBYTES[3].a/w1012 ), .B(
        \SUBBYTES[3].a/w1022 ), .Z(n9278) );
  XOR \SUBBYTES[3].a/U4212  ( .A(n9280), .B(n9279), .Z(\SUBBYTES[3].a/w1037 )
         );
  XOR \SUBBYTES[3].a/U4211  ( .A(n9625), .B(n9281), .Z(n9279) );
  XOR \SUBBYTES[3].a/U4210  ( .A(\w1[3][92] ), .B(\SUBBYTES[3].a/w1101 ), .Z(
        n9280) );
  XOR \SUBBYTES[3].a/U4209  ( .A(\SUBBYTES[3].a/w1014 ), .B(
        \SUBBYTES[3].a/w1019 ), .Z(n9281) );
  XOR \SUBBYTES[3].a/U4208  ( .A(n9283), .B(n9282), .Z(n9623) );
  XOR \SUBBYTES[3].a/U4207  ( .A(\SUBBYTES[3].a/w1047 ), .B(\w1[3][95] ), .Z(
        n9282) );
  XOR \SUBBYTES[3].a/U4206  ( .A(\SUBBYTES[3].a/w1022 ), .B(
        \SUBBYTES[3].a/w1029 ), .Z(n9283) );
  XOR \SUBBYTES[3].a/U4205  ( .A(n9622), .B(n9623), .Z(\SUBBYTES[3].a/w1049 )
         );
  XOR \SUBBYTES[3].a/U4204  ( .A(\w1[3][91] ), .B(n9284), .Z(n9626) );
  XOR \SUBBYTES[3].a/U4203  ( .A(\SUBBYTES[3].a/w1011 ), .B(
        \SUBBYTES[3].a/w1014 ), .Z(n9284) );
  XOR \SUBBYTES[3].a/U4202  ( .A(n9286), .B(n9285), .Z(\SUBBYTES[3].a/w1038 )
         );
  XOR \SUBBYTES[3].a/U4201  ( .A(n9626), .B(n9287), .Z(n9285) );
  XOR \SUBBYTES[3].a/U4200  ( .A(\w1[3][94] ), .B(\SUBBYTES[3].a/w1080 ), .Z(
        n9286) );
  XOR \SUBBYTES[3].a/U4199  ( .A(\SUBBYTES[3].a/w1019 ), .B(
        \SUBBYTES[3].a/w1020 ), .Z(n9287) );
  XOR \SUBBYTES[3].a/U4198  ( .A(n9624), .B(n9623), .Z(\SUBBYTES[3].a/w1058 )
         );
  XOR \SUBBYTES[3].a/U4197  ( .A(n9289), .B(n9288), .Z(\SUBBYTES[3].a/w1059 )
         );
  XOR \SUBBYTES[3].a/U4196  ( .A(\w1[3][95] ), .B(n9625), .Z(n9288) );
  XOR \SUBBYTES[3].a/U4195  ( .A(\SUBBYTES[3].a/w1011 ), .B(
        \SUBBYTES[3].a/w1020 ), .Z(n9289) );
  XOR \SUBBYTES[3].a/U4194  ( .A(n9291), .B(n9290), .Z(\SUBBYTES[3].a/w1035 )
         );
  XOR \SUBBYTES[3].a/U4193  ( .A(n9293), .B(n9292), .Z(n9290) );
  XOR \SUBBYTES[3].a/U4192  ( .A(\w1[3][95] ), .B(\SUBBYTES[3].a/w1119 ), .Z(
        n9291) );
  XOR \SUBBYTES[3].a/U4191  ( .A(\SUBBYTES[3].a/w1026 ), .B(
        \SUBBYTES[3].a/w1029 ), .Z(n9292) );
  XOR \SUBBYTES[3].a/U4190  ( .A(\SUBBYTES[3].a/w1012 ), .B(
        \SUBBYTES[3].a/w1014 ), .Z(n9293) );
  XOR \SUBBYTES[3].a/U4189  ( .A(n9295), .B(n9294), .Z(\SUBBYTES[3].a/w1036 )
         );
  XOR \SUBBYTES[3].a/U4188  ( .A(n9626), .B(n9296), .Z(n9294) );
  XOR \SUBBYTES[3].a/U4187  ( .A(\w1[3][93] ), .B(n9627), .Z(n9295) );
  XOR \SUBBYTES[3].a/U4186  ( .A(\SUBBYTES[3].a/w1026 ), .B(
        \SUBBYTES[3].a/w1027 ), .Z(n9296) );
  XOR \SUBBYTES[3].a/U4185  ( .A(n9298), .B(n9297), .Z(\SUBBYTES[3].a/w1052 )
         );
  XOR \SUBBYTES[3].a/U4184  ( .A(\w1[3][89] ), .B(n9299), .Z(n9297) );
  XOR \SUBBYTES[3].a/U4183  ( .A(\SUBBYTES[3].a/w1027 ), .B(
        \SUBBYTES[3].a/w1029 ), .Z(n9298) );
  XOR \SUBBYTES[3].a/U4182  ( .A(\SUBBYTES[3].a/w1011 ), .B(
        \SUBBYTES[3].a/w1012 ), .Z(n9299) );
  XOR \SUBBYTES[3].a/U4181  ( .A(\w1[3][97] ), .B(n9300), .Z(n9628) );
  XOR \SUBBYTES[3].a/U4180  ( .A(\w1[3][99] ), .B(\w1[3][98] ), .Z(n9300) );
  XOR \SUBBYTES[3].a/U4179  ( .A(\w1[3][102] ), .B(n9628), .Z(
        \SUBBYTES[3].a/w894 ) );
  XOR \SUBBYTES[3].a/U4178  ( .A(\w1[3][96] ), .B(\SUBBYTES[3].a/w894 ), .Z(
        \SUBBYTES[3].a/w781 ) );
  XOR \SUBBYTES[3].a/U4177  ( .A(\w1[3][96] ), .B(n9301), .Z(
        \SUBBYTES[3].a/w782 ) );
  XOR \SUBBYTES[3].a/U4176  ( .A(\w1[3][102] ), .B(\w1[3][101] ), .Z(n9301) );
  XOR \SUBBYTES[3].a/U4175  ( .A(\w1[3][101] ), .B(n9628), .Z(
        \SUBBYTES[3].a/w912 ) );
  XOR \SUBBYTES[3].a/U4174  ( .A(n9303), .B(n9302), .Z(\SUBBYTES[3].a/w905 )
         );
  XOR \SUBBYTES[3].a/U4173  ( .A(\w1[3][99] ), .B(\w1[3][97] ), .Z(n9302) );
  XOR \SUBBYTES[3].a/U4172  ( .A(\w1[3][103] ), .B(\w1[3][100] ), .Z(n9303) );
  XOR \SUBBYTES[3].a/U4171  ( .A(\w1[3][96] ), .B(\SUBBYTES[3].a/w905 ), .Z(
        \SUBBYTES[3].a/w784 ) );
  XOR \SUBBYTES[3].a/U4170  ( .A(n9305), .B(n9304), .Z(\SUBBYTES[3].a/w892 )
         );
  XOR \SUBBYTES[3].a/U4169  ( .A(\SUBBYTES[3].a/w853 ), .B(n992), .Z(n9304) );
  XOR \SUBBYTES[3].a/U4168  ( .A(\SUBBYTES[3].a/w846 ), .B(
        \SUBBYTES[3].a/w849 ), .Z(n9305) );
  XOR \SUBBYTES[3].a/U4167  ( .A(n9307), .B(n9306), .Z(\SUBBYTES[3].a/w893 )
         );
  XOR \SUBBYTES[3].a/U4166  ( .A(\SUBBYTES[3].a/w853 ), .B(n8399), .Z(n9306)
         );
  XOR \SUBBYTES[3].a/U4165  ( .A(\SUBBYTES[3].a/w846 ), .B(n8398), .Z(n9307)
         );
  XOR \SUBBYTES[3].a/U4164  ( .A(\SUBBYTES[3].a/w905 ), .B(n9308), .Z(
        \SUBBYTES[3].a/w895 ) );
  XOR \SUBBYTES[3].a/U4163  ( .A(\w1[3][102] ), .B(\w1[3][101] ), .Z(n9308) );
  XOR \SUBBYTES[3].a/U4162  ( .A(n9310), .B(n9309), .Z(\SUBBYTES[3].a/w896 )
         );
  XOR \SUBBYTES[3].a/U4161  ( .A(n8399), .B(n992), .Z(n9309) );
  XOR \SUBBYTES[3].a/U4160  ( .A(n8398), .B(\SUBBYTES[3].a/w849 ), .Z(n9310)
         );
  XOR \SUBBYTES[3].a/U4159  ( .A(\w1[3][103] ), .B(\w1[3][98] ), .Z(n9634) );
  XOR \SUBBYTES[3].a/U4158  ( .A(n9634), .B(n9311), .Z(\SUBBYTES[3].a/w897 )
         );
  XOR \SUBBYTES[3].a/U4157  ( .A(\w1[3][101] ), .B(\w1[3][100] ), .Z(n9311) );
  XOR \SUBBYTES[3].a/U4156  ( .A(\w1[3][103] ), .B(\SUBBYTES[3].a/w782 ), .Z(
        \SUBBYTES[3].a/w785 ) );
  XOR \SUBBYTES[3].a/U4155  ( .A(\w1[3][97] ), .B(\SUBBYTES[3].a/w782 ), .Z(
        \SUBBYTES[3].a/w786 ) );
  XOR \SUBBYTES[3].a/U4154  ( .A(\w1[3][100] ), .B(\SUBBYTES[3].a/w782 ), .Z(
        \SUBBYTES[3].a/w787 ) );
  XOR \SUBBYTES[3].a/U4153  ( .A(\SUBBYTES[3].a/w786 ), .B(n9634), .Z(
        \SUBBYTES[3].a/w788 ) );
  XOR \SUBBYTES[3].a/U4152  ( .A(n9634), .B(n9312), .Z(\SUBBYTES[3].a/w873 )
         );
  XOR \SUBBYTES[3].a/U4151  ( .A(\w1[3][100] ), .B(\w1[3][97] ), .Z(n9312) );
  XOR \SUBBYTES[3].a/U4150  ( .A(n9314), .B(n9313), .Z(n9631) );
  XOR \SUBBYTES[3].a/U4149  ( .A(\w1[3][100] ), .B(n9315), .Z(n9313) );
  XOR \SUBBYTES[3].a/U4148  ( .A(\SUBBYTES[3].a/w838 ), .B(\w1[3][102] ), .Z(
        n9314) );
  XOR \SUBBYTES[3].a/U4147  ( .A(\SUBBYTES[3].a/w812 ), .B(
        \SUBBYTES[3].a/w819 ), .Z(n9315) );
  XOR \SUBBYTES[3].a/U4146  ( .A(n9317), .B(n9316), .Z(n9629) );
  XOR \SUBBYTES[3].a/U4145  ( .A(\w1[3][97] ), .B(n9318), .Z(n9316) );
  XOR \SUBBYTES[3].a/U4144  ( .A(\SUBBYTES[3].a/w837 ), .B(\w1[3][101] ), .Z(
        n9317) );
  XOR \SUBBYTES[3].a/U4143  ( .A(\SUBBYTES[3].a/w813 ), .B(
        \SUBBYTES[3].a/w820 ), .Z(n9318) );
  XOR \SUBBYTES[3].a/U4142  ( .A(n9631), .B(n9629), .Z(\SUBBYTES[3].a/w843 )
         );
  XOR \SUBBYTES[3].a/U4141  ( .A(\w1[3][101] ), .B(n9319), .Z(n9632) );
  XOR \SUBBYTES[3].a/U4140  ( .A(\SUBBYTES[3].a/w805 ), .B(
        \SUBBYTES[3].a/w815 ), .Z(n9319) );
  XOR \SUBBYTES[3].a/U4139  ( .A(n9321), .B(n9320), .Z(\SUBBYTES[3].a/w830 )
         );
  XOR \SUBBYTES[3].a/U4138  ( .A(n9632), .B(n9322), .Z(n9320) );
  XOR \SUBBYTES[3].a/U4137  ( .A(\w1[3][100] ), .B(\SUBBYTES[3].a/w894 ), .Z(
        n9321) );
  XOR \SUBBYTES[3].a/U4136  ( .A(\SUBBYTES[3].a/w807 ), .B(
        \SUBBYTES[3].a/w812 ), .Z(n9322) );
  XOR \SUBBYTES[3].a/U4135  ( .A(n9324), .B(n9323), .Z(n9630) );
  XOR \SUBBYTES[3].a/U4134  ( .A(\SUBBYTES[3].a/w840 ), .B(\w1[3][103] ), .Z(
        n9323) );
  XOR \SUBBYTES[3].a/U4133  ( .A(\SUBBYTES[3].a/w815 ), .B(
        \SUBBYTES[3].a/w822 ), .Z(n9324) );
  XOR \SUBBYTES[3].a/U4132  ( .A(n9629), .B(n9630), .Z(\SUBBYTES[3].a/w842 )
         );
  XOR \SUBBYTES[3].a/U4131  ( .A(\w1[3][99] ), .B(n9325), .Z(n9633) );
  XOR \SUBBYTES[3].a/U4130  ( .A(\SUBBYTES[3].a/w804 ), .B(
        \SUBBYTES[3].a/w807 ), .Z(n9325) );
  XOR \SUBBYTES[3].a/U4129  ( .A(n9327), .B(n9326), .Z(\SUBBYTES[3].a/w831 )
         );
  XOR \SUBBYTES[3].a/U4128  ( .A(n9633), .B(n9328), .Z(n9326) );
  XOR \SUBBYTES[3].a/U4127  ( .A(\w1[3][102] ), .B(\SUBBYTES[3].a/w873 ), .Z(
        n9327) );
  XOR \SUBBYTES[3].a/U4126  ( .A(\SUBBYTES[3].a/w812 ), .B(
        \SUBBYTES[3].a/w813 ), .Z(n9328) );
  XOR \SUBBYTES[3].a/U4125  ( .A(n9631), .B(n9630), .Z(\SUBBYTES[3].a/w851 )
         );
  XOR \SUBBYTES[3].a/U4124  ( .A(n9330), .B(n9329), .Z(\SUBBYTES[3].a/w852 )
         );
  XOR \SUBBYTES[3].a/U4123  ( .A(\w1[3][103] ), .B(n9632), .Z(n9329) );
  XOR \SUBBYTES[3].a/U4122  ( .A(\SUBBYTES[3].a/w804 ), .B(
        \SUBBYTES[3].a/w813 ), .Z(n9330) );
  XOR \SUBBYTES[3].a/U4121  ( .A(n9332), .B(n9331), .Z(\SUBBYTES[3].a/w828 )
         );
  XOR \SUBBYTES[3].a/U4120  ( .A(n9334), .B(n9333), .Z(n9331) );
  XOR \SUBBYTES[3].a/U4119  ( .A(\w1[3][103] ), .B(\SUBBYTES[3].a/w912 ), .Z(
        n9332) );
  XOR \SUBBYTES[3].a/U4118  ( .A(\SUBBYTES[3].a/w819 ), .B(
        \SUBBYTES[3].a/w822 ), .Z(n9333) );
  XOR \SUBBYTES[3].a/U4117  ( .A(\SUBBYTES[3].a/w805 ), .B(
        \SUBBYTES[3].a/w807 ), .Z(n9334) );
  XOR \SUBBYTES[3].a/U4116  ( .A(n9336), .B(n9335), .Z(\SUBBYTES[3].a/w829 )
         );
  XOR \SUBBYTES[3].a/U4115  ( .A(n9633), .B(n9337), .Z(n9335) );
  XOR \SUBBYTES[3].a/U4114  ( .A(\w1[3][101] ), .B(n9634), .Z(n9336) );
  XOR \SUBBYTES[3].a/U4113  ( .A(\SUBBYTES[3].a/w819 ), .B(
        \SUBBYTES[3].a/w820 ), .Z(n9337) );
  XOR \SUBBYTES[3].a/U4112  ( .A(n9339), .B(n9338), .Z(\SUBBYTES[3].a/w845 )
         );
  XOR \SUBBYTES[3].a/U4111  ( .A(\w1[3][97] ), .B(n9340), .Z(n9338) );
  XOR \SUBBYTES[3].a/U4110  ( .A(\SUBBYTES[3].a/w820 ), .B(
        \SUBBYTES[3].a/w822 ), .Z(n9339) );
  XOR \SUBBYTES[3].a/U4109  ( .A(\SUBBYTES[3].a/w804 ), .B(
        \SUBBYTES[3].a/w805 ), .Z(n9340) );
  XOR \SUBBYTES[3].a/U4108  ( .A(\w1[3][105] ), .B(n9341), .Z(n9635) );
  XOR \SUBBYTES[3].a/U4107  ( .A(\w1[3][107] ), .B(\w1[3][106] ), .Z(n9341) );
  XOR \SUBBYTES[3].a/U4106  ( .A(\w1[3][110] ), .B(n9635), .Z(
        \SUBBYTES[3].a/w687 ) );
  XOR \SUBBYTES[3].a/U4105  ( .A(\w1[3][104] ), .B(\SUBBYTES[3].a/w687 ), .Z(
        \SUBBYTES[3].a/w574 ) );
  XOR \SUBBYTES[3].a/U4104  ( .A(\w1[3][104] ), .B(n9342), .Z(
        \SUBBYTES[3].a/w575 ) );
  XOR \SUBBYTES[3].a/U4103  ( .A(\w1[3][110] ), .B(\w1[3][109] ), .Z(n9342) );
  XOR \SUBBYTES[3].a/U4102  ( .A(\w1[3][109] ), .B(n9635), .Z(
        \SUBBYTES[3].a/w705 ) );
  XOR \SUBBYTES[3].a/U4101  ( .A(n9344), .B(n9343), .Z(\SUBBYTES[3].a/w698 )
         );
  XOR \SUBBYTES[3].a/U4100  ( .A(\w1[3][107] ), .B(\w1[3][105] ), .Z(n9343) );
  XOR \SUBBYTES[3].a/U4099  ( .A(\w1[3][111] ), .B(\w1[3][108] ), .Z(n9344) );
  XOR \SUBBYTES[3].a/U4098  ( .A(\w1[3][104] ), .B(\SUBBYTES[3].a/w698 ), .Z(
        \SUBBYTES[3].a/w577 ) );
  XOR \SUBBYTES[3].a/U4097  ( .A(n9346), .B(n9345), .Z(\SUBBYTES[3].a/w685 )
         );
  XOR \SUBBYTES[3].a/U4096  ( .A(\SUBBYTES[3].a/w646 ), .B(n991), .Z(n9345) );
  XOR \SUBBYTES[3].a/U4095  ( .A(\SUBBYTES[3].a/w639 ), .B(
        \SUBBYTES[3].a/w642 ), .Z(n9346) );
  XOR \SUBBYTES[3].a/U4094  ( .A(n9348), .B(n9347), .Z(\SUBBYTES[3].a/w686 )
         );
  XOR \SUBBYTES[3].a/U4093  ( .A(\SUBBYTES[3].a/w646 ), .B(n8397), .Z(n9347)
         );
  XOR \SUBBYTES[3].a/U4092  ( .A(\SUBBYTES[3].a/w639 ), .B(n8396), .Z(n9348)
         );
  XOR \SUBBYTES[3].a/U4091  ( .A(\SUBBYTES[3].a/w698 ), .B(n9349), .Z(
        \SUBBYTES[3].a/w688 ) );
  XOR \SUBBYTES[3].a/U4090  ( .A(\w1[3][110] ), .B(\w1[3][109] ), .Z(n9349) );
  XOR \SUBBYTES[3].a/U4089  ( .A(n9351), .B(n9350), .Z(\SUBBYTES[3].a/w689 )
         );
  XOR \SUBBYTES[3].a/U4088  ( .A(n8397), .B(n991), .Z(n9350) );
  XOR \SUBBYTES[3].a/U4087  ( .A(n8396), .B(\SUBBYTES[3].a/w642 ), .Z(n9351)
         );
  XOR \SUBBYTES[3].a/U4086  ( .A(\w1[3][111] ), .B(\w1[3][106] ), .Z(n9641) );
  XOR \SUBBYTES[3].a/U4085  ( .A(n9641), .B(n9352), .Z(\SUBBYTES[3].a/w690 )
         );
  XOR \SUBBYTES[3].a/U4084  ( .A(\w1[3][109] ), .B(\w1[3][108] ), .Z(n9352) );
  XOR \SUBBYTES[3].a/U4083  ( .A(\w1[3][111] ), .B(\SUBBYTES[3].a/w575 ), .Z(
        \SUBBYTES[3].a/w578 ) );
  XOR \SUBBYTES[3].a/U4082  ( .A(\w1[3][105] ), .B(\SUBBYTES[3].a/w575 ), .Z(
        \SUBBYTES[3].a/w579 ) );
  XOR \SUBBYTES[3].a/U4081  ( .A(\w1[3][108] ), .B(\SUBBYTES[3].a/w575 ), .Z(
        \SUBBYTES[3].a/w580 ) );
  XOR \SUBBYTES[3].a/U4080  ( .A(\SUBBYTES[3].a/w579 ), .B(n9641), .Z(
        \SUBBYTES[3].a/w581 ) );
  XOR \SUBBYTES[3].a/U4079  ( .A(n9641), .B(n9353), .Z(\SUBBYTES[3].a/w666 )
         );
  XOR \SUBBYTES[3].a/U4078  ( .A(\w1[3][108] ), .B(\w1[3][105] ), .Z(n9353) );
  XOR \SUBBYTES[3].a/U4077  ( .A(n9355), .B(n9354), .Z(n9638) );
  XOR \SUBBYTES[3].a/U4076  ( .A(\w1[3][108] ), .B(n9356), .Z(n9354) );
  XOR \SUBBYTES[3].a/U4075  ( .A(\SUBBYTES[3].a/w631 ), .B(\w1[3][110] ), .Z(
        n9355) );
  XOR \SUBBYTES[3].a/U4074  ( .A(\SUBBYTES[3].a/w605 ), .B(
        \SUBBYTES[3].a/w612 ), .Z(n9356) );
  XOR \SUBBYTES[3].a/U4073  ( .A(n9358), .B(n9357), .Z(n9636) );
  XOR \SUBBYTES[3].a/U4072  ( .A(\w1[3][105] ), .B(n9359), .Z(n9357) );
  XOR \SUBBYTES[3].a/U4071  ( .A(\SUBBYTES[3].a/w630 ), .B(\w1[3][109] ), .Z(
        n9358) );
  XOR \SUBBYTES[3].a/U4070  ( .A(\SUBBYTES[3].a/w606 ), .B(
        \SUBBYTES[3].a/w613 ), .Z(n9359) );
  XOR \SUBBYTES[3].a/U4069  ( .A(n9638), .B(n9636), .Z(\SUBBYTES[3].a/w636 )
         );
  XOR \SUBBYTES[3].a/U4068  ( .A(\w1[3][109] ), .B(n9360), .Z(n9639) );
  XOR \SUBBYTES[3].a/U4067  ( .A(\SUBBYTES[3].a/w598 ), .B(
        \SUBBYTES[3].a/w608 ), .Z(n9360) );
  XOR \SUBBYTES[3].a/U4066  ( .A(n9362), .B(n9361), .Z(\SUBBYTES[3].a/w623 )
         );
  XOR \SUBBYTES[3].a/U4065  ( .A(n9639), .B(n9363), .Z(n9361) );
  XOR \SUBBYTES[3].a/U4064  ( .A(\w1[3][108] ), .B(\SUBBYTES[3].a/w687 ), .Z(
        n9362) );
  XOR \SUBBYTES[3].a/U4063  ( .A(\SUBBYTES[3].a/w600 ), .B(
        \SUBBYTES[3].a/w605 ), .Z(n9363) );
  XOR \SUBBYTES[3].a/U4062  ( .A(n9365), .B(n9364), .Z(n9637) );
  XOR \SUBBYTES[3].a/U4061  ( .A(\SUBBYTES[3].a/w633 ), .B(\w1[3][111] ), .Z(
        n9364) );
  XOR \SUBBYTES[3].a/U4060  ( .A(\SUBBYTES[3].a/w608 ), .B(
        \SUBBYTES[3].a/w615 ), .Z(n9365) );
  XOR \SUBBYTES[3].a/U4059  ( .A(n9636), .B(n9637), .Z(\SUBBYTES[3].a/w635 )
         );
  XOR \SUBBYTES[3].a/U4058  ( .A(\w1[3][107] ), .B(n9366), .Z(n9640) );
  XOR \SUBBYTES[3].a/U4057  ( .A(\SUBBYTES[3].a/w597 ), .B(
        \SUBBYTES[3].a/w600 ), .Z(n9366) );
  XOR \SUBBYTES[3].a/U4056  ( .A(n9368), .B(n9367), .Z(\SUBBYTES[3].a/w624 )
         );
  XOR \SUBBYTES[3].a/U4055  ( .A(n9640), .B(n9369), .Z(n9367) );
  XOR \SUBBYTES[3].a/U4054  ( .A(\w1[3][110] ), .B(\SUBBYTES[3].a/w666 ), .Z(
        n9368) );
  XOR \SUBBYTES[3].a/U4053  ( .A(\SUBBYTES[3].a/w605 ), .B(
        \SUBBYTES[3].a/w606 ), .Z(n9369) );
  XOR \SUBBYTES[3].a/U4052  ( .A(n9638), .B(n9637), .Z(\SUBBYTES[3].a/w644 )
         );
  XOR \SUBBYTES[3].a/U4051  ( .A(n9371), .B(n9370), .Z(\SUBBYTES[3].a/w645 )
         );
  XOR \SUBBYTES[3].a/U4050  ( .A(\w1[3][111] ), .B(n9639), .Z(n9370) );
  XOR \SUBBYTES[3].a/U4049  ( .A(\SUBBYTES[3].a/w597 ), .B(
        \SUBBYTES[3].a/w606 ), .Z(n9371) );
  XOR \SUBBYTES[3].a/U4048  ( .A(n9373), .B(n9372), .Z(\SUBBYTES[3].a/w621 )
         );
  XOR \SUBBYTES[3].a/U4047  ( .A(n9375), .B(n9374), .Z(n9372) );
  XOR \SUBBYTES[3].a/U4046  ( .A(\w1[3][111] ), .B(\SUBBYTES[3].a/w705 ), .Z(
        n9373) );
  XOR \SUBBYTES[3].a/U4045  ( .A(\SUBBYTES[3].a/w612 ), .B(
        \SUBBYTES[3].a/w615 ), .Z(n9374) );
  XOR \SUBBYTES[3].a/U4044  ( .A(\SUBBYTES[3].a/w598 ), .B(
        \SUBBYTES[3].a/w600 ), .Z(n9375) );
  XOR \SUBBYTES[3].a/U4043  ( .A(n9377), .B(n9376), .Z(\SUBBYTES[3].a/w622 )
         );
  XOR \SUBBYTES[3].a/U4042  ( .A(n9640), .B(n9378), .Z(n9376) );
  XOR \SUBBYTES[3].a/U4041  ( .A(\w1[3][109] ), .B(n9641), .Z(n9377) );
  XOR \SUBBYTES[3].a/U4040  ( .A(\SUBBYTES[3].a/w612 ), .B(
        \SUBBYTES[3].a/w613 ), .Z(n9378) );
  XOR \SUBBYTES[3].a/U4039  ( .A(n9380), .B(n9379), .Z(\SUBBYTES[3].a/w638 )
         );
  XOR \SUBBYTES[3].a/U4038  ( .A(\w1[3][105] ), .B(n9381), .Z(n9379) );
  XOR \SUBBYTES[3].a/U4037  ( .A(\SUBBYTES[3].a/w613 ), .B(
        \SUBBYTES[3].a/w615 ), .Z(n9380) );
  XOR \SUBBYTES[3].a/U4036  ( .A(\SUBBYTES[3].a/w597 ), .B(
        \SUBBYTES[3].a/w598 ), .Z(n9381) );
  XOR \SUBBYTES[3].a/U4035  ( .A(\w1[3][113] ), .B(n9382), .Z(n9642) );
  XOR \SUBBYTES[3].a/U4034  ( .A(\w1[3][115] ), .B(\w1[3][114] ), .Z(n9382) );
  XOR \SUBBYTES[3].a/U4033  ( .A(\w1[3][118] ), .B(n9642), .Z(
        \SUBBYTES[3].a/w480 ) );
  XOR \SUBBYTES[3].a/U4032  ( .A(\w1[3][112] ), .B(\SUBBYTES[3].a/w480 ), .Z(
        \SUBBYTES[3].a/w367 ) );
  XOR \SUBBYTES[3].a/U4031  ( .A(\w1[3][112] ), .B(n9383), .Z(
        \SUBBYTES[3].a/w368 ) );
  XOR \SUBBYTES[3].a/U4030  ( .A(\w1[3][118] ), .B(\w1[3][117] ), .Z(n9383) );
  XOR \SUBBYTES[3].a/U4029  ( .A(\w1[3][117] ), .B(n9642), .Z(
        \SUBBYTES[3].a/w498 ) );
  XOR \SUBBYTES[3].a/U4028  ( .A(n9385), .B(n9384), .Z(\SUBBYTES[3].a/w491 )
         );
  XOR \SUBBYTES[3].a/U4027  ( .A(\w1[3][115] ), .B(\w1[3][113] ), .Z(n9384) );
  XOR \SUBBYTES[3].a/U4026  ( .A(\w1[3][119] ), .B(\w1[3][116] ), .Z(n9385) );
  XOR \SUBBYTES[3].a/U4025  ( .A(\w1[3][112] ), .B(\SUBBYTES[3].a/w491 ), .Z(
        \SUBBYTES[3].a/w370 ) );
  XOR \SUBBYTES[3].a/U4024  ( .A(n9387), .B(n9386), .Z(\SUBBYTES[3].a/w478 )
         );
  XOR \SUBBYTES[3].a/U4023  ( .A(\SUBBYTES[3].a/w439 ), .B(n990), .Z(n9386) );
  XOR \SUBBYTES[3].a/U4022  ( .A(\SUBBYTES[3].a/w432 ), .B(
        \SUBBYTES[3].a/w435 ), .Z(n9387) );
  XOR \SUBBYTES[3].a/U4021  ( .A(n9389), .B(n9388), .Z(\SUBBYTES[3].a/w479 )
         );
  XOR \SUBBYTES[3].a/U4020  ( .A(\SUBBYTES[3].a/w439 ), .B(n8395), .Z(n9388)
         );
  XOR \SUBBYTES[3].a/U4019  ( .A(\SUBBYTES[3].a/w432 ), .B(n8394), .Z(n9389)
         );
  XOR \SUBBYTES[3].a/U4018  ( .A(\SUBBYTES[3].a/w491 ), .B(n9390), .Z(
        \SUBBYTES[3].a/w481 ) );
  XOR \SUBBYTES[3].a/U4017  ( .A(\w1[3][118] ), .B(\w1[3][117] ), .Z(n9390) );
  XOR \SUBBYTES[3].a/U4016  ( .A(n9392), .B(n9391), .Z(\SUBBYTES[3].a/w482 )
         );
  XOR \SUBBYTES[3].a/U4015  ( .A(n8395), .B(n990), .Z(n9391) );
  XOR \SUBBYTES[3].a/U4014  ( .A(n8394), .B(\SUBBYTES[3].a/w435 ), .Z(n9392)
         );
  XOR \SUBBYTES[3].a/U4013  ( .A(\w1[3][119] ), .B(\w1[3][114] ), .Z(n9648) );
  XOR \SUBBYTES[3].a/U4012  ( .A(n9648), .B(n9393), .Z(\SUBBYTES[3].a/w483 )
         );
  XOR \SUBBYTES[3].a/U4011  ( .A(\w1[3][117] ), .B(\w1[3][116] ), .Z(n9393) );
  XOR \SUBBYTES[3].a/U4010  ( .A(\w1[3][119] ), .B(\SUBBYTES[3].a/w368 ), .Z(
        \SUBBYTES[3].a/w371 ) );
  XOR \SUBBYTES[3].a/U4009  ( .A(\w1[3][113] ), .B(\SUBBYTES[3].a/w368 ), .Z(
        \SUBBYTES[3].a/w372 ) );
  XOR \SUBBYTES[3].a/U4008  ( .A(\w1[3][116] ), .B(\SUBBYTES[3].a/w368 ), .Z(
        \SUBBYTES[3].a/w373 ) );
  XOR \SUBBYTES[3].a/U4007  ( .A(\SUBBYTES[3].a/w372 ), .B(n9648), .Z(
        \SUBBYTES[3].a/w374 ) );
  XOR \SUBBYTES[3].a/U4006  ( .A(n9648), .B(n9394), .Z(\SUBBYTES[3].a/w459 )
         );
  XOR \SUBBYTES[3].a/U4005  ( .A(\w1[3][116] ), .B(\w1[3][113] ), .Z(n9394) );
  XOR \SUBBYTES[3].a/U4004  ( .A(n9396), .B(n9395), .Z(n9645) );
  XOR \SUBBYTES[3].a/U4003  ( .A(\w1[3][116] ), .B(n9397), .Z(n9395) );
  XOR \SUBBYTES[3].a/U4002  ( .A(\SUBBYTES[3].a/w424 ), .B(\w1[3][118] ), .Z(
        n9396) );
  XOR \SUBBYTES[3].a/U4001  ( .A(\SUBBYTES[3].a/w398 ), .B(
        \SUBBYTES[3].a/w405 ), .Z(n9397) );
  XOR \SUBBYTES[3].a/U4000  ( .A(n9399), .B(n9398), .Z(n9643) );
  XOR \SUBBYTES[3].a/U3999  ( .A(\w1[3][113] ), .B(n9400), .Z(n9398) );
  XOR \SUBBYTES[3].a/U3998  ( .A(\SUBBYTES[3].a/w423 ), .B(\w1[3][117] ), .Z(
        n9399) );
  XOR \SUBBYTES[3].a/U3997  ( .A(\SUBBYTES[3].a/w399 ), .B(
        \SUBBYTES[3].a/w406 ), .Z(n9400) );
  XOR \SUBBYTES[3].a/U3996  ( .A(n9645), .B(n9643), .Z(\SUBBYTES[3].a/w429 )
         );
  XOR \SUBBYTES[3].a/U3995  ( .A(\w1[3][117] ), .B(n9401), .Z(n9646) );
  XOR \SUBBYTES[3].a/U3994  ( .A(\SUBBYTES[3].a/w391 ), .B(
        \SUBBYTES[3].a/w401 ), .Z(n9401) );
  XOR \SUBBYTES[3].a/U3993  ( .A(n9403), .B(n9402), .Z(\SUBBYTES[3].a/w416 )
         );
  XOR \SUBBYTES[3].a/U3992  ( .A(n9646), .B(n9404), .Z(n9402) );
  XOR \SUBBYTES[3].a/U3991  ( .A(\w1[3][116] ), .B(\SUBBYTES[3].a/w480 ), .Z(
        n9403) );
  XOR \SUBBYTES[3].a/U3990  ( .A(\SUBBYTES[3].a/w393 ), .B(
        \SUBBYTES[3].a/w398 ), .Z(n9404) );
  XOR \SUBBYTES[3].a/U3989  ( .A(n9406), .B(n9405), .Z(n9644) );
  XOR \SUBBYTES[3].a/U3988  ( .A(\SUBBYTES[3].a/w426 ), .B(\w1[3][119] ), .Z(
        n9405) );
  XOR \SUBBYTES[3].a/U3987  ( .A(\SUBBYTES[3].a/w401 ), .B(
        \SUBBYTES[3].a/w408 ), .Z(n9406) );
  XOR \SUBBYTES[3].a/U3986  ( .A(n9643), .B(n9644), .Z(\SUBBYTES[3].a/w428 )
         );
  XOR \SUBBYTES[3].a/U3985  ( .A(\w1[3][115] ), .B(n9407), .Z(n9647) );
  XOR \SUBBYTES[3].a/U3984  ( .A(\SUBBYTES[3].a/w390 ), .B(
        \SUBBYTES[3].a/w393 ), .Z(n9407) );
  XOR \SUBBYTES[3].a/U3983  ( .A(n9409), .B(n9408), .Z(\SUBBYTES[3].a/w417 )
         );
  XOR \SUBBYTES[3].a/U3982  ( .A(n9647), .B(n9410), .Z(n9408) );
  XOR \SUBBYTES[3].a/U3981  ( .A(\w1[3][118] ), .B(\SUBBYTES[3].a/w459 ), .Z(
        n9409) );
  XOR \SUBBYTES[3].a/U3980  ( .A(\SUBBYTES[3].a/w398 ), .B(
        \SUBBYTES[3].a/w399 ), .Z(n9410) );
  XOR \SUBBYTES[3].a/U3979  ( .A(n9645), .B(n9644), .Z(\SUBBYTES[3].a/w437 )
         );
  XOR \SUBBYTES[3].a/U3978  ( .A(n9412), .B(n9411), .Z(\SUBBYTES[3].a/w438 )
         );
  XOR \SUBBYTES[3].a/U3977  ( .A(\w1[3][119] ), .B(n9646), .Z(n9411) );
  XOR \SUBBYTES[3].a/U3976  ( .A(\SUBBYTES[3].a/w390 ), .B(
        \SUBBYTES[3].a/w399 ), .Z(n9412) );
  XOR \SUBBYTES[3].a/U3975  ( .A(n9414), .B(n9413), .Z(\SUBBYTES[3].a/w414 )
         );
  XOR \SUBBYTES[3].a/U3974  ( .A(n9416), .B(n9415), .Z(n9413) );
  XOR \SUBBYTES[3].a/U3973  ( .A(\w1[3][119] ), .B(\SUBBYTES[3].a/w498 ), .Z(
        n9414) );
  XOR \SUBBYTES[3].a/U3972  ( .A(\SUBBYTES[3].a/w405 ), .B(
        \SUBBYTES[3].a/w408 ), .Z(n9415) );
  XOR \SUBBYTES[3].a/U3971  ( .A(\SUBBYTES[3].a/w391 ), .B(
        \SUBBYTES[3].a/w393 ), .Z(n9416) );
  XOR \SUBBYTES[3].a/U3970  ( .A(n9418), .B(n9417), .Z(\SUBBYTES[3].a/w415 )
         );
  XOR \SUBBYTES[3].a/U3969  ( .A(n9647), .B(n9419), .Z(n9417) );
  XOR \SUBBYTES[3].a/U3968  ( .A(\w1[3][117] ), .B(n9648), .Z(n9418) );
  XOR \SUBBYTES[3].a/U3967  ( .A(\SUBBYTES[3].a/w405 ), .B(
        \SUBBYTES[3].a/w406 ), .Z(n9419) );
  XOR \SUBBYTES[3].a/U3966  ( .A(n9421), .B(n9420), .Z(\SUBBYTES[3].a/w431 )
         );
  XOR \SUBBYTES[3].a/U3965  ( .A(\w1[3][113] ), .B(n9422), .Z(n9420) );
  XOR \SUBBYTES[3].a/U3964  ( .A(\SUBBYTES[3].a/w406 ), .B(
        \SUBBYTES[3].a/w408 ), .Z(n9421) );
  XOR \SUBBYTES[3].a/U3963  ( .A(\SUBBYTES[3].a/w390 ), .B(
        \SUBBYTES[3].a/w391 ), .Z(n9422) );
  XOR \SUBBYTES[3].a/U3962  ( .A(\w1[3][121] ), .B(n9423), .Z(n9649) );
  XOR \SUBBYTES[3].a/U3961  ( .A(\w1[3][123] ), .B(\w1[3][122] ), .Z(n9423) );
  XOR \SUBBYTES[3].a/U3960  ( .A(\w1[3][126] ), .B(n9649), .Z(
        \SUBBYTES[3].a/w273 ) );
  XOR \SUBBYTES[3].a/U3959  ( .A(\w1[3][120] ), .B(\SUBBYTES[3].a/w273 ), .Z(
        \SUBBYTES[3].a/w160 ) );
  XOR \SUBBYTES[3].a/U3958  ( .A(\w1[3][120] ), .B(n9424), .Z(
        \SUBBYTES[3].a/w161 ) );
  XOR \SUBBYTES[3].a/U3957  ( .A(\w1[3][126] ), .B(\w1[3][125] ), .Z(n9424) );
  XOR \SUBBYTES[3].a/U3956  ( .A(\w1[3][125] ), .B(n9649), .Z(
        \SUBBYTES[3].a/w291 ) );
  XOR \SUBBYTES[3].a/U3955  ( .A(n9426), .B(n9425), .Z(\SUBBYTES[3].a/w284 )
         );
  XOR \SUBBYTES[3].a/U3954  ( .A(\w1[3][123] ), .B(\w1[3][121] ), .Z(n9425) );
  XOR \SUBBYTES[3].a/U3953  ( .A(\w1[3][127] ), .B(\w1[3][124] ), .Z(n9426) );
  XOR \SUBBYTES[3].a/U3952  ( .A(\w1[3][120] ), .B(\SUBBYTES[3].a/w284 ), .Z(
        \SUBBYTES[3].a/w163 ) );
  XOR \SUBBYTES[3].a/U3951  ( .A(n9428), .B(n9427), .Z(\SUBBYTES[3].a/w271 )
         );
  XOR \SUBBYTES[3].a/U3950  ( .A(\SUBBYTES[3].a/w232 ), .B(n989), .Z(n9427) );
  XOR \SUBBYTES[3].a/U3949  ( .A(\SUBBYTES[3].a/w225 ), .B(
        \SUBBYTES[3].a/w228 ), .Z(n9428) );
  XOR \SUBBYTES[3].a/U3948  ( .A(n9430), .B(n9429), .Z(\SUBBYTES[3].a/w272 )
         );
  XOR \SUBBYTES[3].a/U3947  ( .A(\SUBBYTES[3].a/w232 ), .B(n8393), .Z(n9429)
         );
  XOR \SUBBYTES[3].a/U3946  ( .A(\SUBBYTES[3].a/w225 ), .B(n8392), .Z(n9430)
         );
  XOR \SUBBYTES[3].a/U3945  ( .A(\SUBBYTES[3].a/w284 ), .B(n9431), .Z(
        \SUBBYTES[3].a/w274 ) );
  XOR \SUBBYTES[3].a/U3944  ( .A(\w1[3][126] ), .B(\w1[3][125] ), .Z(n9431) );
  XOR \SUBBYTES[3].a/U3943  ( .A(n9433), .B(n9432), .Z(\SUBBYTES[3].a/w275 )
         );
  XOR \SUBBYTES[3].a/U3942  ( .A(n8393), .B(n989), .Z(n9432) );
  XOR \SUBBYTES[3].a/U3941  ( .A(n8392), .B(\SUBBYTES[3].a/w228 ), .Z(n9433)
         );
  XOR \SUBBYTES[3].a/U3940  ( .A(\w1[3][127] ), .B(\w1[3][122] ), .Z(n9655) );
  XOR \SUBBYTES[3].a/U3939  ( .A(n9655), .B(n9434), .Z(\SUBBYTES[3].a/w276 )
         );
  XOR \SUBBYTES[3].a/U3938  ( .A(\w1[3][125] ), .B(\w1[3][124] ), .Z(n9434) );
  XOR \SUBBYTES[3].a/U3937  ( .A(\w1[3][127] ), .B(\SUBBYTES[3].a/w161 ), .Z(
        \SUBBYTES[3].a/w164 ) );
  XOR \SUBBYTES[3].a/U3936  ( .A(\w1[3][121] ), .B(\SUBBYTES[3].a/w161 ), .Z(
        \SUBBYTES[3].a/w165 ) );
  XOR \SUBBYTES[3].a/U3935  ( .A(\w1[3][124] ), .B(\SUBBYTES[3].a/w161 ), .Z(
        \SUBBYTES[3].a/w166 ) );
  XOR \SUBBYTES[3].a/U3934  ( .A(\SUBBYTES[3].a/w165 ), .B(n9655), .Z(
        \SUBBYTES[3].a/w167 ) );
  XOR \SUBBYTES[3].a/U3933  ( .A(n9655), .B(n9435), .Z(\SUBBYTES[3].a/w252 )
         );
  XOR \SUBBYTES[3].a/U3932  ( .A(\w1[3][124] ), .B(\w1[3][121] ), .Z(n9435) );
  XOR \SUBBYTES[3].a/U3931  ( .A(n9437), .B(n9436), .Z(n9652) );
  XOR \SUBBYTES[3].a/U3930  ( .A(\w1[3][124] ), .B(n9438), .Z(n9436) );
  XOR \SUBBYTES[3].a/U3929  ( .A(\SUBBYTES[3].a/w217 ), .B(\w1[3][126] ), .Z(
        n9437) );
  XOR \SUBBYTES[3].a/U3928  ( .A(\SUBBYTES[3].a/w191 ), .B(
        \SUBBYTES[3].a/w198 ), .Z(n9438) );
  XOR \SUBBYTES[3].a/U3927  ( .A(n9440), .B(n9439), .Z(n9650) );
  XOR \SUBBYTES[3].a/U3926  ( .A(\w1[3][121] ), .B(n9441), .Z(n9439) );
  XOR \SUBBYTES[3].a/U3925  ( .A(\SUBBYTES[3].a/w216 ), .B(\w1[3][125] ), .Z(
        n9440) );
  XOR \SUBBYTES[3].a/U3924  ( .A(\SUBBYTES[3].a/w192 ), .B(
        \SUBBYTES[3].a/w199 ), .Z(n9441) );
  XOR \SUBBYTES[3].a/U3923  ( .A(n9652), .B(n9650), .Z(\SUBBYTES[3].a/w222 )
         );
  XOR \SUBBYTES[3].a/U3922  ( .A(\w1[3][125] ), .B(n9442), .Z(n9653) );
  XOR \SUBBYTES[3].a/U3921  ( .A(\SUBBYTES[3].a/w184 ), .B(
        \SUBBYTES[3].a/w194 ), .Z(n9442) );
  XOR \SUBBYTES[3].a/U3920  ( .A(n9444), .B(n9443), .Z(\SUBBYTES[3].a/w209 )
         );
  XOR \SUBBYTES[3].a/U3919  ( .A(n9653), .B(n9445), .Z(n9443) );
  XOR \SUBBYTES[3].a/U3918  ( .A(\w1[3][124] ), .B(\SUBBYTES[3].a/w273 ), .Z(
        n9444) );
  XOR \SUBBYTES[3].a/U3917  ( .A(\SUBBYTES[3].a/w186 ), .B(
        \SUBBYTES[3].a/w191 ), .Z(n9445) );
  XOR \SUBBYTES[3].a/U3916  ( .A(n9447), .B(n9446), .Z(n9651) );
  XOR \SUBBYTES[3].a/U3915  ( .A(\SUBBYTES[3].a/w219 ), .B(\w1[3][127] ), .Z(
        n9446) );
  XOR \SUBBYTES[3].a/U3914  ( .A(\SUBBYTES[3].a/w194 ), .B(
        \SUBBYTES[3].a/w201 ), .Z(n9447) );
  XOR \SUBBYTES[3].a/U3913  ( .A(n9650), .B(n9651), .Z(\SUBBYTES[3].a/w221 )
         );
  XOR \SUBBYTES[3].a/U3912  ( .A(\w1[3][123] ), .B(n9448), .Z(n9654) );
  XOR \SUBBYTES[3].a/U3911  ( .A(\SUBBYTES[3].a/w183 ), .B(
        \SUBBYTES[3].a/w186 ), .Z(n9448) );
  XOR \SUBBYTES[3].a/U3910  ( .A(n9450), .B(n9449), .Z(\SUBBYTES[3].a/w210 )
         );
  XOR \SUBBYTES[3].a/U3909  ( .A(n9654), .B(n9451), .Z(n9449) );
  XOR \SUBBYTES[3].a/U3908  ( .A(\w1[3][126] ), .B(\SUBBYTES[3].a/w252 ), .Z(
        n9450) );
  XOR \SUBBYTES[3].a/U3907  ( .A(\SUBBYTES[3].a/w191 ), .B(
        \SUBBYTES[3].a/w192 ), .Z(n9451) );
  XOR \SUBBYTES[3].a/U3906  ( .A(n9652), .B(n9651), .Z(\SUBBYTES[3].a/w230 )
         );
  XOR \SUBBYTES[3].a/U3905  ( .A(n9453), .B(n9452), .Z(\SUBBYTES[3].a/w231 )
         );
  XOR \SUBBYTES[3].a/U3904  ( .A(\w1[3][127] ), .B(n9653), .Z(n9452) );
  XOR \SUBBYTES[3].a/U3903  ( .A(\SUBBYTES[3].a/w183 ), .B(
        \SUBBYTES[3].a/w192 ), .Z(n9453) );
  XOR \SUBBYTES[3].a/U3902  ( .A(n9455), .B(n9454), .Z(\SUBBYTES[3].a/w207 )
         );
  XOR \SUBBYTES[3].a/U3901  ( .A(n9457), .B(n9456), .Z(n9454) );
  XOR \SUBBYTES[3].a/U3900  ( .A(\w1[3][127] ), .B(\SUBBYTES[3].a/w291 ), .Z(
        n9455) );
  XOR \SUBBYTES[3].a/U3899  ( .A(\SUBBYTES[3].a/w198 ), .B(
        \SUBBYTES[3].a/w201 ), .Z(n9456) );
  XOR \SUBBYTES[3].a/U3898  ( .A(\SUBBYTES[3].a/w184 ), .B(
        \SUBBYTES[3].a/w186 ), .Z(n9457) );
  XOR \SUBBYTES[3].a/U3897  ( .A(n9459), .B(n9458), .Z(\SUBBYTES[3].a/w208 )
         );
  XOR \SUBBYTES[3].a/U3896  ( .A(n9654), .B(n9460), .Z(n9458) );
  XOR \SUBBYTES[3].a/U3895  ( .A(\w1[3][125] ), .B(n9655), .Z(n9459) );
  XOR \SUBBYTES[3].a/U3894  ( .A(\SUBBYTES[3].a/w198 ), .B(
        \SUBBYTES[3].a/w199 ), .Z(n9460) );
  XOR \SUBBYTES[3].a/U3893  ( .A(n9462), .B(n9461), .Z(\SUBBYTES[3].a/w224 )
         );
  XOR \SUBBYTES[3].a/U3892  ( .A(\w1[3][121] ), .B(n9463), .Z(n9461) );
  XOR \SUBBYTES[3].a/U3891  ( .A(\SUBBYTES[3].a/w199 ), .B(
        \SUBBYTES[3].a/w201 ), .Z(n9462) );
  XOR \SUBBYTES[3].a/U3890  ( .A(\SUBBYTES[3].a/w183 ), .B(
        \SUBBYTES[3].a/w184 ), .Z(n9463) );
  XOR \SUBBYTES[2].a/U5649  ( .A(\SUBBYTES[2].a/w3390 ), .B(
        \SUBBYTES[2].a/w3391 ), .Z(n8185) );
  XOR \SUBBYTES[2].a/U5648  ( .A(n8185), .B(n7144), .Z(n8184) );
  XOR \SUBBYTES[2].a/U5647  ( .A(\SUBBYTES[2].a/w3383 ), .B(
        \SUBBYTES[2].a/w3400 ), .Z(n7144) );
  XOR \SUBBYTES[2].a/U5645  ( .A(\SUBBYTES[2].a/w3382 ), .B(
        \SUBBYTES[2].a/w3397 ), .Z(n7145) );
  XOR \SUBBYTES[2].a/U5644  ( .A(n8185), .B(n7146), .Z(n8376) );
  XOR \SUBBYTES[2].a/U5643  ( .A(\SUBBYTES[2].a/w3397 ), .B(
        \SUBBYTES[2].a/w3398 ), .Z(n7146) );
  XOR \SUBBYTES[2].a/U5642  ( .A(\SUBBYTES[2].a/w3359 ), .B(n7147), .Z(n8187)
         );
  XOR \SUBBYTES[2].a/U5641  ( .A(\SUBBYTES[2].a/w3350 ), .B(
        \SUBBYTES[2].a/w3351 ), .Z(n7147) );
  XOR \SUBBYTES[2].a/U5639  ( .A(\SUBBYTES[2].a/w3361 ), .B(n8376), .Z(n7148)
         );
  XOR \SUBBYTES[2].a/U5638  ( .A(n7150), .B(n7149), .Z(n8188) );
  XOR \SUBBYTES[2].a/U5637  ( .A(n7152), .B(n7151), .Z(n7149) );
  XOR \SUBBYTES[2].a/U5636  ( .A(\SUBBYTES[2].a/w3397 ), .B(
        \SUBBYTES[2].a/w3398 ), .Z(n7150) );
  XOR \SUBBYTES[2].a/U5635  ( .A(\SUBBYTES[2].a/w3361 ), .B(
        \SUBBYTES[2].a/w3385 ), .Z(n7151) );
  XOR \SUBBYTES[2].a/U5634  ( .A(\SUBBYTES[2].a/w3350 ), .B(
        \SUBBYTES[2].a/w3359 ), .Z(n7152) );
  XOR \SUBBYTES[2].a/U5633  ( .A(\SUBBYTES[2].a/w3382 ), .B(n7153), .Z(n8186)
         );
  XOR \SUBBYTES[2].a/U5632  ( .A(\SUBBYTES[2].a/w3365 ), .B(
        \SUBBYTES[2].a/w3368 ), .Z(n7153) );
  XOR \SUBBYTES[2].a/U5630  ( .A(\SUBBYTES[2].a/w3353 ), .B(n8188), .Z(n7154)
         );
  XOR \SUBBYTES[2].a/U5628  ( .A(\SUBBYTES[2].a/w3385 ), .B(
        \SUBBYTES[2].a/w3398 ), .Z(n7155) );
  XOR \SUBBYTES[2].a/U5626  ( .A(n7159), .B(n7158), .Z(n7156) );
  XOR \SUBBYTES[2].a/U5625  ( .A(n7161), .B(n7160), .Z(n7157) );
  XOR \SUBBYTES[2].a/U5624  ( .A(\SUBBYTES[2].a/w3397 ), .B(
        \SUBBYTES[2].a/w3400 ), .Z(n7158) );
  XOR \SUBBYTES[2].a/U5623  ( .A(\SUBBYTES[2].a/w3390 ), .B(
        \SUBBYTES[2].a/w3393 ), .Z(n7159) );
  XOR \SUBBYTES[2].a/U5622  ( .A(\SUBBYTES[2].a/w3365 ), .B(
        \SUBBYTES[2].a/w3366 ), .Z(n7160) );
  XOR \SUBBYTES[2].a/U5621  ( .A(\SUBBYTES[2].a/w3350 ), .B(
        \SUBBYTES[2].a/w3353 ), .Z(n7161) );
  XOR \SUBBYTES[2].a/U5619  ( .A(n8185), .B(n7164), .Z(n7162) );
  XOR \SUBBYTES[2].a/U5618  ( .A(n8187), .B(n8186), .Z(n7163) );
  XOR \SUBBYTES[2].a/U5617  ( .A(\SUBBYTES[2].a/w3358 ), .B(
        \SUBBYTES[2].a/w3385 ), .Z(n7164) );
  XOR \SUBBYTES[2].a/U5615  ( .A(n8188), .B(n7167), .Z(n7165) );
  XOR \SUBBYTES[2].a/U5614  ( .A(\SUBBYTES[2].a/w3391 ), .B(
        \SUBBYTES[2].a/w3393 ), .Z(n7166) );
  XOR \SUBBYTES[2].a/U5613  ( .A(\SUBBYTES[2].a/w3351 ), .B(
        \SUBBYTES[2].a/w3383 ), .Z(n7167) );
  XOR \SUBBYTES[2].a/U5612  ( .A(\SUBBYTES[2].a/w3183 ), .B(
        \SUBBYTES[2].a/w3184 ), .Z(n8190) );
  XOR \SUBBYTES[2].a/U5611  ( .A(n8190), .B(n7168), .Z(n8189) );
  XOR \SUBBYTES[2].a/U5610  ( .A(\SUBBYTES[2].a/w3176 ), .B(
        \SUBBYTES[2].a/w3193 ), .Z(n7168) );
  XOR \SUBBYTES[2].a/U5608  ( .A(\SUBBYTES[2].a/w3175 ), .B(
        \SUBBYTES[2].a/w3190 ), .Z(n7169) );
  XOR \SUBBYTES[2].a/U5607  ( .A(n8190), .B(n7170), .Z(n8377) );
  XOR \SUBBYTES[2].a/U5606  ( .A(\SUBBYTES[2].a/w3190 ), .B(
        \SUBBYTES[2].a/w3191 ), .Z(n7170) );
  XOR \SUBBYTES[2].a/U5605  ( .A(\SUBBYTES[2].a/w3152 ), .B(n7171), .Z(n8192)
         );
  XOR \SUBBYTES[2].a/U5604  ( .A(\SUBBYTES[2].a/w3143 ), .B(
        \SUBBYTES[2].a/w3144 ), .Z(n7171) );
  XOR \SUBBYTES[2].a/U5602  ( .A(\SUBBYTES[2].a/w3154 ), .B(n8377), .Z(n7172)
         );
  XOR \SUBBYTES[2].a/U5601  ( .A(n7174), .B(n7173), .Z(n8193) );
  XOR \SUBBYTES[2].a/U5600  ( .A(n7176), .B(n7175), .Z(n7173) );
  XOR \SUBBYTES[2].a/U5599  ( .A(\SUBBYTES[2].a/w3190 ), .B(
        \SUBBYTES[2].a/w3191 ), .Z(n7174) );
  XOR \SUBBYTES[2].a/U5598  ( .A(\SUBBYTES[2].a/w3154 ), .B(
        \SUBBYTES[2].a/w3178 ), .Z(n7175) );
  XOR \SUBBYTES[2].a/U5597  ( .A(\SUBBYTES[2].a/w3143 ), .B(
        \SUBBYTES[2].a/w3152 ), .Z(n7176) );
  XOR \SUBBYTES[2].a/U5596  ( .A(\SUBBYTES[2].a/w3175 ), .B(n7177), .Z(n8191)
         );
  XOR \SUBBYTES[2].a/U5595  ( .A(\SUBBYTES[2].a/w3158 ), .B(
        \SUBBYTES[2].a/w3161 ), .Z(n7177) );
  XOR \SUBBYTES[2].a/U5593  ( .A(\SUBBYTES[2].a/w3146 ), .B(n8193), .Z(n7178)
         );
  XOR \SUBBYTES[2].a/U5591  ( .A(\SUBBYTES[2].a/w3178 ), .B(
        \SUBBYTES[2].a/w3191 ), .Z(n7179) );
  XOR \SUBBYTES[2].a/U5589  ( .A(n7183), .B(n7182), .Z(n7180) );
  XOR \SUBBYTES[2].a/U5588  ( .A(n7185), .B(n7184), .Z(n7181) );
  XOR \SUBBYTES[2].a/U5587  ( .A(\SUBBYTES[2].a/w3190 ), .B(
        \SUBBYTES[2].a/w3193 ), .Z(n7182) );
  XOR \SUBBYTES[2].a/U5586  ( .A(\SUBBYTES[2].a/w3183 ), .B(
        \SUBBYTES[2].a/w3186 ), .Z(n7183) );
  XOR \SUBBYTES[2].a/U5585  ( .A(\SUBBYTES[2].a/w3158 ), .B(
        \SUBBYTES[2].a/w3159 ), .Z(n7184) );
  XOR \SUBBYTES[2].a/U5584  ( .A(\SUBBYTES[2].a/w3143 ), .B(
        \SUBBYTES[2].a/w3146 ), .Z(n7185) );
  XOR \SUBBYTES[2].a/U5582  ( .A(n8190), .B(n7188), .Z(n7186) );
  XOR \SUBBYTES[2].a/U5581  ( .A(n8192), .B(n8191), .Z(n7187) );
  XOR \SUBBYTES[2].a/U5580  ( .A(\SUBBYTES[2].a/w3151 ), .B(
        \SUBBYTES[2].a/w3178 ), .Z(n7188) );
  XOR \SUBBYTES[2].a/U5578  ( .A(n8193), .B(n7191), .Z(n7189) );
  XOR \SUBBYTES[2].a/U5577  ( .A(\SUBBYTES[2].a/w3184 ), .B(
        \SUBBYTES[2].a/w3186 ), .Z(n7190) );
  XOR \SUBBYTES[2].a/U5576  ( .A(\SUBBYTES[2].a/w3144 ), .B(
        \SUBBYTES[2].a/w3176 ), .Z(n7191) );
  XOR \SUBBYTES[2].a/U5575  ( .A(\SUBBYTES[2].a/w2976 ), .B(
        \SUBBYTES[2].a/w2977 ), .Z(n8195) );
  XOR \SUBBYTES[2].a/U5574  ( .A(n8195), .B(n7192), .Z(n8194) );
  XOR \SUBBYTES[2].a/U5573  ( .A(\SUBBYTES[2].a/w2969 ), .B(
        \SUBBYTES[2].a/w2986 ), .Z(n7192) );
  XOR \SUBBYTES[2].a/U5571  ( .A(\SUBBYTES[2].a/w2968 ), .B(
        \SUBBYTES[2].a/w2983 ), .Z(n7193) );
  XOR \SUBBYTES[2].a/U5570  ( .A(n8195), .B(n7194), .Z(n8378) );
  XOR \SUBBYTES[2].a/U5569  ( .A(\SUBBYTES[2].a/w2983 ), .B(
        \SUBBYTES[2].a/w2984 ), .Z(n7194) );
  XOR \SUBBYTES[2].a/U5568  ( .A(\SUBBYTES[2].a/w2945 ), .B(n7195), .Z(n8197)
         );
  XOR \SUBBYTES[2].a/U5567  ( .A(\SUBBYTES[2].a/w2936 ), .B(
        \SUBBYTES[2].a/w2937 ), .Z(n7195) );
  XOR \SUBBYTES[2].a/U5565  ( .A(\SUBBYTES[2].a/w2947 ), .B(n8378), .Z(n7196)
         );
  XOR \SUBBYTES[2].a/U5564  ( .A(n7198), .B(n7197), .Z(n8198) );
  XOR \SUBBYTES[2].a/U5563  ( .A(n7200), .B(n7199), .Z(n7197) );
  XOR \SUBBYTES[2].a/U5562  ( .A(\SUBBYTES[2].a/w2983 ), .B(
        \SUBBYTES[2].a/w2984 ), .Z(n7198) );
  XOR \SUBBYTES[2].a/U5561  ( .A(\SUBBYTES[2].a/w2947 ), .B(
        \SUBBYTES[2].a/w2971 ), .Z(n7199) );
  XOR \SUBBYTES[2].a/U5560  ( .A(\SUBBYTES[2].a/w2936 ), .B(
        \SUBBYTES[2].a/w2945 ), .Z(n7200) );
  XOR \SUBBYTES[2].a/U5559  ( .A(\SUBBYTES[2].a/w2968 ), .B(n7201), .Z(n8196)
         );
  XOR \SUBBYTES[2].a/U5558  ( .A(\SUBBYTES[2].a/w2951 ), .B(
        \SUBBYTES[2].a/w2954 ), .Z(n7201) );
  XOR \SUBBYTES[2].a/U5556  ( .A(\SUBBYTES[2].a/w2939 ), .B(n8198), .Z(n7202)
         );
  XOR \SUBBYTES[2].a/U5554  ( .A(\SUBBYTES[2].a/w2971 ), .B(
        \SUBBYTES[2].a/w2984 ), .Z(n7203) );
  XOR \SUBBYTES[2].a/U5552  ( .A(n7207), .B(n7206), .Z(n7204) );
  XOR \SUBBYTES[2].a/U5551  ( .A(n7209), .B(n7208), .Z(n7205) );
  XOR \SUBBYTES[2].a/U5550  ( .A(\SUBBYTES[2].a/w2983 ), .B(
        \SUBBYTES[2].a/w2986 ), .Z(n7206) );
  XOR \SUBBYTES[2].a/U5549  ( .A(\SUBBYTES[2].a/w2976 ), .B(
        \SUBBYTES[2].a/w2979 ), .Z(n7207) );
  XOR \SUBBYTES[2].a/U5548  ( .A(\SUBBYTES[2].a/w2951 ), .B(
        \SUBBYTES[2].a/w2952 ), .Z(n7208) );
  XOR \SUBBYTES[2].a/U5547  ( .A(\SUBBYTES[2].a/w2936 ), .B(
        \SUBBYTES[2].a/w2939 ), .Z(n7209) );
  XOR \SUBBYTES[2].a/U5545  ( .A(n8195), .B(n7212), .Z(n7210) );
  XOR \SUBBYTES[2].a/U5544  ( .A(n8197), .B(n8196), .Z(n7211) );
  XOR \SUBBYTES[2].a/U5543  ( .A(\SUBBYTES[2].a/w2944 ), .B(
        \SUBBYTES[2].a/w2971 ), .Z(n7212) );
  XOR \SUBBYTES[2].a/U5541  ( .A(n8198), .B(n7215), .Z(n7213) );
  XOR \SUBBYTES[2].a/U5540  ( .A(\SUBBYTES[2].a/w2977 ), .B(
        \SUBBYTES[2].a/w2979 ), .Z(n7214) );
  XOR \SUBBYTES[2].a/U5539  ( .A(\SUBBYTES[2].a/w2937 ), .B(
        \SUBBYTES[2].a/w2969 ), .Z(n7215) );
  XOR \SUBBYTES[2].a/U5538  ( .A(\SUBBYTES[2].a/w2769 ), .B(
        \SUBBYTES[2].a/w2770 ), .Z(n8200) );
  XOR \SUBBYTES[2].a/U5537  ( .A(n8200), .B(n7216), .Z(n8199) );
  XOR \SUBBYTES[2].a/U5536  ( .A(\SUBBYTES[2].a/w2762 ), .B(
        \SUBBYTES[2].a/w2779 ), .Z(n7216) );
  XOR \SUBBYTES[2].a/U5534  ( .A(\SUBBYTES[2].a/w2761 ), .B(
        \SUBBYTES[2].a/w2776 ), .Z(n7217) );
  XOR \SUBBYTES[2].a/U5533  ( .A(n8200), .B(n7218), .Z(n8379) );
  XOR \SUBBYTES[2].a/U5532  ( .A(\SUBBYTES[2].a/w2776 ), .B(
        \SUBBYTES[2].a/w2777 ), .Z(n7218) );
  XOR \SUBBYTES[2].a/U5531  ( .A(\SUBBYTES[2].a/w2738 ), .B(n7219), .Z(n8202)
         );
  XOR \SUBBYTES[2].a/U5530  ( .A(\SUBBYTES[2].a/w2729 ), .B(
        \SUBBYTES[2].a/w2730 ), .Z(n7219) );
  XOR \SUBBYTES[2].a/U5528  ( .A(\SUBBYTES[2].a/w2740 ), .B(n8379), .Z(n7220)
         );
  XOR \SUBBYTES[2].a/U5527  ( .A(n7222), .B(n7221), .Z(n8203) );
  XOR \SUBBYTES[2].a/U5526  ( .A(n7224), .B(n7223), .Z(n7221) );
  XOR \SUBBYTES[2].a/U5525  ( .A(\SUBBYTES[2].a/w2776 ), .B(
        \SUBBYTES[2].a/w2777 ), .Z(n7222) );
  XOR \SUBBYTES[2].a/U5524  ( .A(\SUBBYTES[2].a/w2740 ), .B(
        \SUBBYTES[2].a/w2764 ), .Z(n7223) );
  XOR \SUBBYTES[2].a/U5523  ( .A(\SUBBYTES[2].a/w2729 ), .B(
        \SUBBYTES[2].a/w2738 ), .Z(n7224) );
  XOR \SUBBYTES[2].a/U5522  ( .A(\SUBBYTES[2].a/w2761 ), .B(n7225), .Z(n8201)
         );
  XOR \SUBBYTES[2].a/U5521  ( .A(\SUBBYTES[2].a/w2744 ), .B(
        \SUBBYTES[2].a/w2747 ), .Z(n7225) );
  XOR \SUBBYTES[2].a/U5519  ( .A(\SUBBYTES[2].a/w2732 ), .B(n8203), .Z(n7226)
         );
  XOR \SUBBYTES[2].a/U5517  ( .A(\SUBBYTES[2].a/w2764 ), .B(
        \SUBBYTES[2].a/w2777 ), .Z(n7227) );
  XOR \SUBBYTES[2].a/U5515  ( .A(n7231), .B(n7230), .Z(n7228) );
  XOR \SUBBYTES[2].a/U5514  ( .A(n7233), .B(n7232), .Z(n7229) );
  XOR \SUBBYTES[2].a/U5513  ( .A(\SUBBYTES[2].a/w2776 ), .B(
        \SUBBYTES[2].a/w2779 ), .Z(n7230) );
  XOR \SUBBYTES[2].a/U5512  ( .A(\SUBBYTES[2].a/w2769 ), .B(
        \SUBBYTES[2].a/w2772 ), .Z(n7231) );
  XOR \SUBBYTES[2].a/U5511  ( .A(\SUBBYTES[2].a/w2744 ), .B(
        \SUBBYTES[2].a/w2745 ), .Z(n7232) );
  XOR \SUBBYTES[2].a/U5510  ( .A(\SUBBYTES[2].a/w2729 ), .B(
        \SUBBYTES[2].a/w2732 ), .Z(n7233) );
  XOR \SUBBYTES[2].a/U5508  ( .A(n8200), .B(n7236), .Z(n7234) );
  XOR \SUBBYTES[2].a/U5507  ( .A(n8202), .B(n8201), .Z(n7235) );
  XOR \SUBBYTES[2].a/U5506  ( .A(\SUBBYTES[2].a/w2737 ), .B(
        \SUBBYTES[2].a/w2764 ), .Z(n7236) );
  XOR \SUBBYTES[2].a/U5504  ( .A(n8203), .B(n7239), .Z(n7237) );
  XOR \SUBBYTES[2].a/U5503  ( .A(\SUBBYTES[2].a/w2770 ), .B(
        \SUBBYTES[2].a/w2772 ), .Z(n7238) );
  XOR \SUBBYTES[2].a/U5502  ( .A(\SUBBYTES[2].a/w2730 ), .B(
        \SUBBYTES[2].a/w2762 ), .Z(n7239) );
  XOR \SUBBYTES[2].a/U5501  ( .A(\SUBBYTES[2].a/w2562 ), .B(
        \SUBBYTES[2].a/w2563 ), .Z(n8205) );
  XOR \SUBBYTES[2].a/U5500  ( .A(n8205), .B(n7240), .Z(n8204) );
  XOR \SUBBYTES[2].a/U5499  ( .A(\SUBBYTES[2].a/w2555 ), .B(
        \SUBBYTES[2].a/w2572 ), .Z(n7240) );
  XOR \SUBBYTES[2].a/U5497  ( .A(\SUBBYTES[2].a/w2554 ), .B(
        \SUBBYTES[2].a/w2569 ), .Z(n7241) );
  XOR \SUBBYTES[2].a/U5496  ( .A(n8205), .B(n7242), .Z(n8380) );
  XOR \SUBBYTES[2].a/U5495  ( .A(\SUBBYTES[2].a/w2569 ), .B(
        \SUBBYTES[2].a/w2570 ), .Z(n7242) );
  XOR \SUBBYTES[2].a/U5494  ( .A(\SUBBYTES[2].a/w2531 ), .B(n7243), .Z(n8207)
         );
  XOR \SUBBYTES[2].a/U5493  ( .A(\SUBBYTES[2].a/w2522 ), .B(
        \SUBBYTES[2].a/w2523 ), .Z(n7243) );
  XOR \SUBBYTES[2].a/U5491  ( .A(\SUBBYTES[2].a/w2533 ), .B(n8380), .Z(n7244)
         );
  XOR \SUBBYTES[2].a/U5490  ( .A(n7246), .B(n7245), .Z(n8208) );
  XOR \SUBBYTES[2].a/U5489  ( .A(n7248), .B(n7247), .Z(n7245) );
  XOR \SUBBYTES[2].a/U5488  ( .A(\SUBBYTES[2].a/w2569 ), .B(
        \SUBBYTES[2].a/w2570 ), .Z(n7246) );
  XOR \SUBBYTES[2].a/U5487  ( .A(\SUBBYTES[2].a/w2533 ), .B(
        \SUBBYTES[2].a/w2557 ), .Z(n7247) );
  XOR \SUBBYTES[2].a/U5486  ( .A(\SUBBYTES[2].a/w2522 ), .B(
        \SUBBYTES[2].a/w2531 ), .Z(n7248) );
  XOR \SUBBYTES[2].a/U5485  ( .A(\SUBBYTES[2].a/w2554 ), .B(n7249), .Z(n8206)
         );
  XOR \SUBBYTES[2].a/U5484  ( .A(\SUBBYTES[2].a/w2537 ), .B(
        \SUBBYTES[2].a/w2540 ), .Z(n7249) );
  XOR \SUBBYTES[2].a/U5482  ( .A(\SUBBYTES[2].a/w2525 ), .B(n8208), .Z(n7250)
         );
  XOR \SUBBYTES[2].a/U5480  ( .A(\SUBBYTES[2].a/w2557 ), .B(
        \SUBBYTES[2].a/w2570 ), .Z(n7251) );
  XOR \SUBBYTES[2].a/U5478  ( .A(n7255), .B(n7254), .Z(n7252) );
  XOR \SUBBYTES[2].a/U5477  ( .A(n7257), .B(n7256), .Z(n7253) );
  XOR \SUBBYTES[2].a/U5476  ( .A(\SUBBYTES[2].a/w2569 ), .B(
        \SUBBYTES[2].a/w2572 ), .Z(n7254) );
  XOR \SUBBYTES[2].a/U5475  ( .A(\SUBBYTES[2].a/w2562 ), .B(
        \SUBBYTES[2].a/w2565 ), .Z(n7255) );
  XOR \SUBBYTES[2].a/U5474  ( .A(\SUBBYTES[2].a/w2537 ), .B(
        \SUBBYTES[2].a/w2538 ), .Z(n7256) );
  XOR \SUBBYTES[2].a/U5473  ( .A(\SUBBYTES[2].a/w2522 ), .B(
        \SUBBYTES[2].a/w2525 ), .Z(n7257) );
  XOR \SUBBYTES[2].a/U5471  ( .A(n8205), .B(n7260), .Z(n7258) );
  XOR \SUBBYTES[2].a/U5470  ( .A(n8207), .B(n8206), .Z(n7259) );
  XOR \SUBBYTES[2].a/U5469  ( .A(\SUBBYTES[2].a/w2530 ), .B(
        \SUBBYTES[2].a/w2557 ), .Z(n7260) );
  XOR \SUBBYTES[2].a/U5467  ( .A(n8208), .B(n7263), .Z(n7261) );
  XOR \SUBBYTES[2].a/U5466  ( .A(\SUBBYTES[2].a/w2563 ), .B(
        \SUBBYTES[2].a/w2565 ), .Z(n7262) );
  XOR \SUBBYTES[2].a/U5465  ( .A(\SUBBYTES[2].a/w2523 ), .B(
        \SUBBYTES[2].a/w2555 ), .Z(n7263) );
  XOR \SUBBYTES[2].a/U5464  ( .A(\SUBBYTES[2].a/w2355 ), .B(
        \SUBBYTES[2].a/w2356 ), .Z(n8210) );
  XOR \SUBBYTES[2].a/U5463  ( .A(n8210), .B(n7264), .Z(n8209) );
  XOR \SUBBYTES[2].a/U5462  ( .A(\SUBBYTES[2].a/w2348 ), .B(
        \SUBBYTES[2].a/w2365 ), .Z(n7264) );
  XOR \SUBBYTES[2].a/U5460  ( .A(\SUBBYTES[2].a/w2347 ), .B(
        \SUBBYTES[2].a/w2362 ), .Z(n7265) );
  XOR \SUBBYTES[2].a/U5459  ( .A(n8210), .B(n7266), .Z(n8381) );
  XOR \SUBBYTES[2].a/U5458  ( .A(\SUBBYTES[2].a/w2362 ), .B(
        \SUBBYTES[2].a/w2363 ), .Z(n7266) );
  XOR \SUBBYTES[2].a/U5457  ( .A(\SUBBYTES[2].a/w2324 ), .B(n7267), .Z(n8212)
         );
  XOR \SUBBYTES[2].a/U5456  ( .A(\SUBBYTES[2].a/w2315 ), .B(
        \SUBBYTES[2].a/w2316 ), .Z(n7267) );
  XOR \SUBBYTES[2].a/U5454  ( .A(\SUBBYTES[2].a/w2326 ), .B(n8381), .Z(n7268)
         );
  XOR \SUBBYTES[2].a/U5453  ( .A(n7270), .B(n7269), .Z(n8213) );
  XOR \SUBBYTES[2].a/U5452  ( .A(n7272), .B(n7271), .Z(n7269) );
  XOR \SUBBYTES[2].a/U5451  ( .A(\SUBBYTES[2].a/w2362 ), .B(
        \SUBBYTES[2].a/w2363 ), .Z(n7270) );
  XOR \SUBBYTES[2].a/U5450  ( .A(\SUBBYTES[2].a/w2326 ), .B(
        \SUBBYTES[2].a/w2350 ), .Z(n7271) );
  XOR \SUBBYTES[2].a/U5449  ( .A(\SUBBYTES[2].a/w2315 ), .B(
        \SUBBYTES[2].a/w2324 ), .Z(n7272) );
  XOR \SUBBYTES[2].a/U5448  ( .A(\SUBBYTES[2].a/w2347 ), .B(n7273), .Z(n8211)
         );
  XOR \SUBBYTES[2].a/U5447  ( .A(\SUBBYTES[2].a/w2330 ), .B(
        \SUBBYTES[2].a/w2333 ), .Z(n7273) );
  XOR \SUBBYTES[2].a/U5445  ( .A(\SUBBYTES[2].a/w2318 ), .B(n8213), .Z(n7274)
         );
  XOR \SUBBYTES[2].a/U5443  ( .A(\SUBBYTES[2].a/w2350 ), .B(
        \SUBBYTES[2].a/w2363 ), .Z(n7275) );
  XOR \SUBBYTES[2].a/U5441  ( .A(n7279), .B(n7278), .Z(n7276) );
  XOR \SUBBYTES[2].a/U5440  ( .A(n7281), .B(n7280), .Z(n7277) );
  XOR \SUBBYTES[2].a/U5439  ( .A(\SUBBYTES[2].a/w2362 ), .B(
        \SUBBYTES[2].a/w2365 ), .Z(n7278) );
  XOR \SUBBYTES[2].a/U5438  ( .A(\SUBBYTES[2].a/w2355 ), .B(
        \SUBBYTES[2].a/w2358 ), .Z(n7279) );
  XOR \SUBBYTES[2].a/U5437  ( .A(\SUBBYTES[2].a/w2330 ), .B(
        \SUBBYTES[2].a/w2331 ), .Z(n7280) );
  XOR \SUBBYTES[2].a/U5436  ( .A(\SUBBYTES[2].a/w2315 ), .B(
        \SUBBYTES[2].a/w2318 ), .Z(n7281) );
  XOR \SUBBYTES[2].a/U5434  ( .A(n8210), .B(n7284), .Z(n7282) );
  XOR \SUBBYTES[2].a/U5433  ( .A(n8212), .B(n8211), .Z(n7283) );
  XOR \SUBBYTES[2].a/U5432  ( .A(\SUBBYTES[2].a/w2323 ), .B(
        \SUBBYTES[2].a/w2350 ), .Z(n7284) );
  XOR \SUBBYTES[2].a/U5430  ( .A(n8213), .B(n7287), .Z(n7285) );
  XOR \SUBBYTES[2].a/U5429  ( .A(\SUBBYTES[2].a/w2356 ), .B(
        \SUBBYTES[2].a/w2358 ), .Z(n7286) );
  XOR \SUBBYTES[2].a/U5428  ( .A(\SUBBYTES[2].a/w2316 ), .B(
        \SUBBYTES[2].a/w2348 ), .Z(n7287) );
  XOR \SUBBYTES[2].a/U5427  ( .A(\SUBBYTES[2].a/w2148 ), .B(
        \SUBBYTES[2].a/w2149 ), .Z(n8215) );
  XOR \SUBBYTES[2].a/U5426  ( .A(n8215), .B(n7288), .Z(n8214) );
  XOR \SUBBYTES[2].a/U5425  ( .A(\SUBBYTES[2].a/w2141 ), .B(
        \SUBBYTES[2].a/w2158 ), .Z(n7288) );
  XOR \SUBBYTES[2].a/U5423  ( .A(\SUBBYTES[2].a/w2140 ), .B(
        \SUBBYTES[2].a/w2155 ), .Z(n7289) );
  XOR \SUBBYTES[2].a/U5422  ( .A(n8215), .B(n7290), .Z(n8382) );
  XOR \SUBBYTES[2].a/U5421  ( .A(\SUBBYTES[2].a/w2155 ), .B(
        \SUBBYTES[2].a/w2156 ), .Z(n7290) );
  XOR \SUBBYTES[2].a/U5420  ( .A(\SUBBYTES[2].a/w2117 ), .B(n7291), .Z(n8217)
         );
  XOR \SUBBYTES[2].a/U5419  ( .A(\SUBBYTES[2].a/w2108 ), .B(
        \SUBBYTES[2].a/w2109 ), .Z(n7291) );
  XOR \SUBBYTES[2].a/U5417  ( .A(\SUBBYTES[2].a/w2119 ), .B(n8382), .Z(n7292)
         );
  XOR \SUBBYTES[2].a/U5416  ( .A(n7294), .B(n7293), .Z(n8218) );
  XOR \SUBBYTES[2].a/U5415  ( .A(n7296), .B(n7295), .Z(n7293) );
  XOR \SUBBYTES[2].a/U5414  ( .A(\SUBBYTES[2].a/w2155 ), .B(
        \SUBBYTES[2].a/w2156 ), .Z(n7294) );
  XOR \SUBBYTES[2].a/U5413  ( .A(\SUBBYTES[2].a/w2119 ), .B(
        \SUBBYTES[2].a/w2143 ), .Z(n7295) );
  XOR \SUBBYTES[2].a/U5412  ( .A(\SUBBYTES[2].a/w2108 ), .B(
        \SUBBYTES[2].a/w2117 ), .Z(n7296) );
  XOR \SUBBYTES[2].a/U5411  ( .A(\SUBBYTES[2].a/w2140 ), .B(n7297), .Z(n8216)
         );
  XOR \SUBBYTES[2].a/U5410  ( .A(\SUBBYTES[2].a/w2123 ), .B(
        \SUBBYTES[2].a/w2126 ), .Z(n7297) );
  XOR \SUBBYTES[2].a/U5408  ( .A(\SUBBYTES[2].a/w2111 ), .B(n8218), .Z(n7298)
         );
  XOR \SUBBYTES[2].a/U5406  ( .A(\SUBBYTES[2].a/w2143 ), .B(
        \SUBBYTES[2].a/w2156 ), .Z(n7299) );
  XOR \SUBBYTES[2].a/U5404  ( .A(n7303), .B(n7302), .Z(n7300) );
  XOR \SUBBYTES[2].a/U5403  ( .A(n7305), .B(n7304), .Z(n7301) );
  XOR \SUBBYTES[2].a/U5402  ( .A(\SUBBYTES[2].a/w2155 ), .B(
        \SUBBYTES[2].a/w2158 ), .Z(n7302) );
  XOR \SUBBYTES[2].a/U5401  ( .A(\SUBBYTES[2].a/w2148 ), .B(
        \SUBBYTES[2].a/w2151 ), .Z(n7303) );
  XOR \SUBBYTES[2].a/U5400  ( .A(\SUBBYTES[2].a/w2123 ), .B(
        \SUBBYTES[2].a/w2124 ), .Z(n7304) );
  XOR \SUBBYTES[2].a/U5399  ( .A(\SUBBYTES[2].a/w2108 ), .B(
        \SUBBYTES[2].a/w2111 ), .Z(n7305) );
  XOR \SUBBYTES[2].a/U5397  ( .A(n8215), .B(n7308), .Z(n7306) );
  XOR \SUBBYTES[2].a/U5396  ( .A(n8217), .B(n8216), .Z(n7307) );
  XOR \SUBBYTES[2].a/U5395  ( .A(\SUBBYTES[2].a/w2116 ), .B(
        \SUBBYTES[2].a/w2143 ), .Z(n7308) );
  XOR \SUBBYTES[2].a/U5393  ( .A(n8218), .B(n7311), .Z(n7309) );
  XOR \SUBBYTES[2].a/U5392  ( .A(\SUBBYTES[2].a/w2149 ), .B(
        \SUBBYTES[2].a/w2151 ), .Z(n7310) );
  XOR \SUBBYTES[2].a/U5391  ( .A(\SUBBYTES[2].a/w2109 ), .B(
        \SUBBYTES[2].a/w2141 ), .Z(n7311) );
  XOR \SUBBYTES[2].a/U5390  ( .A(\SUBBYTES[2].a/w1941 ), .B(
        \SUBBYTES[2].a/w1942 ), .Z(n8220) );
  XOR \SUBBYTES[2].a/U5389  ( .A(n8220), .B(n7312), .Z(n8219) );
  XOR \SUBBYTES[2].a/U5388  ( .A(\SUBBYTES[2].a/w1934 ), .B(
        \SUBBYTES[2].a/w1951 ), .Z(n7312) );
  XOR \SUBBYTES[2].a/U5386  ( .A(\SUBBYTES[2].a/w1933 ), .B(
        \SUBBYTES[2].a/w1948 ), .Z(n7313) );
  XOR \SUBBYTES[2].a/U5385  ( .A(n8220), .B(n7314), .Z(n8383) );
  XOR \SUBBYTES[2].a/U5384  ( .A(\SUBBYTES[2].a/w1948 ), .B(
        \SUBBYTES[2].a/w1949 ), .Z(n7314) );
  XOR \SUBBYTES[2].a/U5383  ( .A(\SUBBYTES[2].a/w1910 ), .B(n7315), .Z(n8222)
         );
  XOR \SUBBYTES[2].a/U5382  ( .A(\SUBBYTES[2].a/w1901 ), .B(
        \SUBBYTES[2].a/w1902 ), .Z(n7315) );
  XOR \SUBBYTES[2].a/U5380  ( .A(\SUBBYTES[2].a/w1912 ), .B(n8383), .Z(n7316)
         );
  XOR \SUBBYTES[2].a/U5379  ( .A(n7318), .B(n7317), .Z(n8223) );
  XOR \SUBBYTES[2].a/U5378  ( .A(n7320), .B(n7319), .Z(n7317) );
  XOR \SUBBYTES[2].a/U5377  ( .A(\SUBBYTES[2].a/w1948 ), .B(
        \SUBBYTES[2].a/w1949 ), .Z(n7318) );
  XOR \SUBBYTES[2].a/U5376  ( .A(\SUBBYTES[2].a/w1912 ), .B(
        \SUBBYTES[2].a/w1936 ), .Z(n7319) );
  XOR \SUBBYTES[2].a/U5375  ( .A(\SUBBYTES[2].a/w1901 ), .B(
        \SUBBYTES[2].a/w1910 ), .Z(n7320) );
  XOR \SUBBYTES[2].a/U5374  ( .A(\SUBBYTES[2].a/w1933 ), .B(n7321), .Z(n8221)
         );
  XOR \SUBBYTES[2].a/U5373  ( .A(\SUBBYTES[2].a/w1916 ), .B(
        \SUBBYTES[2].a/w1919 ), .Z(n7321) );
  XOR \SUBBYTES[2].a/U5371  ( .A(\SUBBYTES[2].a/w1904 ), .B(n8223), .Z(n7322)
         );
  XOR \SUBBYTES[2].a/U5369  ( .A(\SUBBYTES[2].a/w1936 ), .B(
        \SUBBYTES[2].a/w1949 ), .Z(n7323) );
  XOR \SUBBYTES[2].a/U5367  ( .A(n7327), .B(n7326), .Z(n7324) );
  XOR \SUBBYTES[2].a/U5366  ( .A(n7329), .B(n7328), .Z(n7325) );
  XOR \SUBBYTES[2].a/U5365  ( .A(\SUBBYTES[2].a/w1948 ), .B(
        \SUBBYTES[2].a/w1951 ), .Z(n7326) );
  XOR \SUBBYTES[2].a/U5364  ( .A(\SUBBYTES[2].a/w1941 ), .B(
        \SUBBYTES[2].a/w1944 ), .Z(n7327) );
  XOR \SUBBYTES[2].a/U5363  ( .A(\SUBBYTES[2].a/w1916 ), .B(
        \SUBBYTES[2].a/w1917 ), .Z(n7328) );
  XOR \SUBBYTES[2].a/U5362  ( .A(\SUBBYTES[2].a/w1901 ), .B(
        \SUBBYTES[2].a/w1904 ), .Z(n7329) );
  XOR \SUBBYTES[2].a/U5360  ( .A(n8220), .B(n7332), .Z(n7330) );
  XOR \SUBBYTES[2].a/U5359  ( .A(n8222), .B(n8221), .Z(n7331) );
  XOR \SUBBYTES[2].a/U5358  ( .A(\SUBBYTES[2].a/w1909 ), .B(
        \SUBBYTES[2].a/w1936 ), .Z(n7332) );
  XOR \SUBBYTES[2].a/U5356  ( .A(n8223), .B(n7335), .Z(n7333) );
  XOR \SUBBYTES[2].a/U5355  ( .A(\SUBBYTES[2].a/w1942 ), .B(
        \SUBBYTES[2].a/w1944 ), .Z(n7334) );
  XOR \SUBBYTES[2].a/U5354  ( .A(\SUBBYTES[2].a/w1902 ), .B(
        \SUBBYTES[2].a/w1934 ), .Z(n7335) );
  XOR \SUBBYTES[2].a/U5353  ( .A(\SUBBYTES[2].a/w1734 ), .B(
        \SUBBYTES[2].a/w1735 ), .Z(n8225) );
  XOR \SUBBYTES[2].a/U5352  ( .A(n8225), .B(n7336), .Z(n8224) );
  XOR \SUBBYTES[2].a/U5351  ( .A(\SUBBYTES[2].a/w1727 ), .B(
        \SUBBYTES[2].a/w1744 ), .Z(n7336) );
  XOR \SUBBYTES[2].a/U5349  ( .A(\SUBBYTES[2].a/w1726 ), .B(
        \SUBBYTES[2].a/w1741 ), .Z(n7337) );
  XOR \SUBBYTES[2].a/U5348  ( .A(n8225), .B(n7338), .Z(n8384) );
  XOR \SUBBYTES[2].a/U5347  ( .A(\SUBBYTES[2].a/w1741 ), .B(
        \SUBBYTES[2].a/w1742 ), .Z(n7338) );
  XOR \SUBBYTES[2].a/U5346  ( .A(\SUBBYTES[2].a/w1703 ), .B(n7339), .Z(n8227)
         );
  XOR \SUBBYTES[2].a/U5345  ( .A(\SUBBYTES[2].a/w1694 ), .B(
        \SUBBYTES[2].a/w1695 ), .Z(n7339) );
  XOR \SUBBYTES[2].a/U5343  ( .A(\SUBBYTES[2].a/w1705 ), .B(n8384), .Z(n7340)
         );
  XOR \SUBBYTES[2].a/U5342  ( .A(n7342), .B(n7341), .Z(n8228) );
  XOR \SUBBYTES[2].a/U5341  ( .A(n7344), .B(n7343), .Z(n7341) );
  XOR \SUBBYTES[2].a/U5340  ( .A(\SUBBYTES[2].a/w1741 ), .B(
        \SUBBYTES[2].a/w1742 ), .Z(n7342) );
  XOR \SUBBYTES[2].a/U5339  ( .A(\SUBBYTES[2].a/w1705 ), .B(
        \SUBBYTES[2].a/w1729 ), .Z(n7343) );
  XOR \SUBBYTES[2].a/U5338  ( .A(\SUBBYTES[2].a/w1694 ), .B(
        \SUBBYTES[2].a/w1703 ), .Z(n7344) );
  XOR \SUBBYTES[2].a/U5337  ( .A(\SUBBYTES[2].a/w1726 ), .B(n7345), .Z(n8226)
         );
  XOR \SUBBYTES[2].a/U5336  ( .A(\SUBBYTES[2].a/w1709 ), .B(
        \SUBBYTES[2].a/w1712 ), .Z(n7345) );
  XOR \SUBBYTES[2].a/U5334  ( .A(\SUBBYTES[2].a/w1697 ), .B(n8228), .Z(n7346)
         );
  XOR \SUBBYTES[2].a/U5332  ( .A(\SUBBYTES[2].a/w1729 ), .B(
        \SUBBYTES[2].a/w1742 ), .Z(n7347) );
  XOR \SUBBYTES[2].a/U5330  ( .A(n7351), .B(n7350), .Z(n7348) );
  XOR \SUBBYTES[2].a/U5329  ( .A(n7353), .B(n7352), .Z(n7349) );
  XOR \SUBBYTES[2].a/U5328  ( .A(\SUBBYTES[2].a/w1741 ), .B(
        \SUBBYTES[2].a/w1744 ), .Z(n7350) );
  XOR \SUBBYTES[2].a/U5327  ( .A(\SUBBYTES[2].a/w1734 ), .B(
        \SUBBYTES[2].a/w1737 ), .Z(n7351) );
  XOR \SUBBYTES[2].a/U5326  ( .A(\SUBBYTES[2].a/w1709 ), .B(
        \SUBBYTES[2].a/w1710 ), .Z(n7352) );
  XOR \SUBBYTES[2].a/U5325  ( .A(\SUBBYTES[2].a/w1694 ), .B(
        \SUBBYTES[2].a/w1697 ), .Z(n7353) );
  XOR \SUBBYTES[2].a/U5323  ( .A(n8225), .B(n7356), .Z(n7354) );
  XOR \SUBBYTES[2].a/U5322  ( .A(n8227), .B(n8226), .Z(n7355) );
  XOR \SUBBYTES[2].a/U5321  ( .A(\SUBBYTES[2].a/w1702 ), .B(
        \SUBBYTES[2].a/w1729 ), .Z(n7356) );
  XOR \SUBBYTES[2].a/U5319  ( .A(n8228), .B(n7359), .Z(n7357) );
  XOR \SUBBYTES[2].a/U5318  ( .A(\SUBBYTES[2].a/w1735 ), .B(
        \SUBBYTES[2].a/w1737 ), .Z(n7358) );
  XOR \SUBBYTES[2].a/U5317  ( .A(\SUBBYTES[2].a/w1695 ), .B(
        \SUBBYTES[2].a/w1727 ), .Z(n7359) );
  XOR \SUBBYTES[2].a/U5316  ( .A(\SUBBYTES[2].a/w1527 ), .B(
        \SUBBYTES[2].a/w1528 ), .Z(n8230) );
  XOR \SUBBYTES[2].a/U5315  ( .A(n8230), .B(n7360), .Z(n8229) );
  XOR \SUBBYTES[2].a/U5314  ( .A(\SUBBYTES[2].a/w1520 ), .B(
        \SUBBYTES[2].a/w1537 ), .Z(n7360) );
  XOR \SUBBYTES[2].a/U5312  ( .A(\SUBBYTES[2].a/w1519 ), .B(
        \SUBBYTES[2].a/w1534 ), .Z(n7361) );
  XOR \SUBBYTES[2].a/U5311  ( .A(n8230), .B(n7362), .Z(n8385) );
  XOR \SUBBYTES[2].a/U5310  ( .A(\SUBBYTES[2].a/w1534 ), .B(
        \SUBBYTES[2].a/w1535 ), .Z(n7362) );
  XOR \SUBBYTES[2].a/U5309  ( .A(\SUBBYTES[2].a/w1496 ), .B(n7363), .Z(n8232)
         );
  XOR \SUBBYTES[2].a/U5308  ( .A(\SUBBYTES[2].a/w1487 ), .B(
        \SUBBYTES[2].a/w1488 ), .Z(n7363) );
  XOR \SUBBYTES[2].a/U5306  ( .A(\SUBBYTES[2].a/w1498 ), .B(n8385), .Z(n7364)
         );
  XOR \SUBBYTES[2].a/U5305  ( .A(n7366), .B(n7365), .Z(n8233) );
  XOR \SUBBYTES[2].a/U5304  ( .A(n7368), .B(n7367), .Z(n7365) );
  XOR \SUBBYTES[2].a/U5303  ( .A(\SUBBYTES[2].a/w1534 ), .B(
        \SUBBYTES[2].a/w1535 ), .Z(n7366) );
  XOR \SUBBYTES[2].a/U5302  ( .A(\SUBBYTES[2].a/w1498 ), .B(
        \SUBBYTES[2].a/w1522 ), .Z(n7367) );
  XOR \SUBBYTES[2].a/U5301  ( .A(\SUBBYTES[2].a/w1487 ), .B(
        \SUBBYTES[2].a/w1496 ), .Z(n7368) );
  XOR \SUBBYTES[2].a/U5300  ( .A(\SUBBYTES[2].a/w1519 ), .B(n7369), .Z(n8231)
         );
  XOR \SUBBYTES[2].a/U5299  ( .A(\SUBBYTES[2].a/w1502 ), .B(
        \SUBBYTES[2].a/w1505 ), .Z(n7369) );
  XOR \SUBBYTES[2].a/U5297  ( .A(\SUBBYTES[2].a/w1490 ), .B(n8233), .Z(n7370)
         );
  XOR \SUBBYTES[2].a/U5295  ( .A(\SUBBYTES[2].a/w1522 ), .B(
        \SUBBYTES[2].a/w1535 ), .Z(n7371) );
  XOR \SUBBYTES[2].a/U5293  ( .A(n7375), .B(n7374), .Z(n7372) );
  XOR \SUBBYTES[2].a/U5292  ( .A(n7377), .B(n7376), .Z(n7373) );
  XOR \SUBBYTES[2].a/U5291  ( .A(\SUBBYTES[2].a/w1534 ), .B(
        \SUBBYTES[2].a/w1537 ), .Z(n7374) );
  XOR \SUBBYTES[2].a/U5290  ( .A(\SUBBYTES[2].a/w1527 ), .B(
        \SUBBYTES[2].a/w1530 ), .Z(n7375) );
  XOR \SUBBYTES[2].a/U5289  ( .A(\SUBBYTES[2].a/w1502 ), .B(
        \SUBBYTES[2].a/w1503 ), .Z(n7376) );
  XOR \SUBBYTES[2].a/U5288  ( .A(\SUBBYTES[2].a/w1487 ), .B(
        \SUBBYTES[2].a/w1490 ), .Z(n7377) );
  XOR \SUBBYTES[2].a/U5286  ( .A(n8230), .B(n7380), .Z(n7378) );
  XOR \SUBBYTES[2].a/U5285  ( .A(n8232), .B(n8231), .Z(n7379) );
  XOR \SUBBYTES[2].a/U5284  ( .A(\SUBBYTES[2].a/w1495 ), .B(
        \SUBBYTES[2].a/w1522 ), .Z(n7380) );
  XOR \SUBBYTES[2].a/U5282  ( .A(n8233), .B(n7383), .Z(n7381) );
  XOR \SUBBYTES[2].a/U5281  ( .A(\SUBBYTES[2].a/w1528 ), .B(
        \SUBBYTES[2].a/w1530 ), .Z(n7382) );
  XOR \SUBBYTES[2].a/U5280  ( .A(\SUBBYTES[2].a/w1488 ), .B(
        \SUBBYTES[2].a/w1520 ), .Z(n7383) );
  XOR \SUBBYTES[2].a/U5279  ( .A(\SUBBYTES[2].a/w1320 ), .B(
        \SUBBYTES[2].a/w1321 ), .Z(n8235) );
  XOR \SUBBYTES[2].a/U5278  ( .A(n8235), .B(n7384), .Z(n8234) );
  XOR \SUBBYTES[2].a/U5277  ( .A(\SUBBYTES[2].a/w1313 ), .B(
        \SUBBYTES[2].a/w1330 ), .Z(n7384) );
  XOR \SUBBYTES[2].a/U5275  ( .A(\SUBBYTES[2].a/w1312 ), .B(
        \SUBBYTES[2].a/w1327 ), .Z(n7385) );
  XOR \SUBBYTES[2].a/U5274  ( .A(n8235), .B(n7386), .Z(n8386) );
  XOR \SUBBYTES[2].a/U5273  ( .A(\SUBBYTES[2].a/w1327 ), .B(
        \SUBBYTES[2].a/w1328 ), .Z(n7386) );
  XOR \SUBBYTES[2].a/U5272  ( .A(\SUBBYTES[2].a/w1289 ), .B(n7387), .Z(n8237)
         );
  XOR \SUBBYTES[2].a/U5271  ( .A(\SUBBYTES[2].a/w1280 ), .B(
        \SUBBYTES[2].a/w1281 ), .Z(n7387) );
  XOR \SUBBYTES[2].a/U5269  ( .A(\SUBBYTES[2].a/w1291 ), .B(n8386), .Z(n7388)
         );
  XOR \SUBBYTES[2].a/U5268  ( .A(n7390), .B(n7389), .Z(n8238) );
  XOR \SUBBYTES[2].a/U5267  ( .A(n7392), .B(n7391), .Z(n7389) );
  XOR \SUBBYTES[2].a/U5266  ( .A(\SUBBYTES[2].a/w1327 ), .B(
        \SUBBYTES[2].a/w1328 ), .Z(n7390) );
  XOR \SUBBYTES[2].a/U5265  ( .A(\SUBBYTES[2].a/w1291 ), .B(
        \SUBBYTES[2].a/w1315 ), .Z(n7391) );
  XOR \SUBBYTES[2].a/U5264  ( .A(\SUBBYTES[2].a/w1280 ), .B(
        \SUBBYTES[2].a/w1289 ), .Z(n7392) );
  XOR \SUBBYTES[2].a/U5263  ( .A(\SUBBYTES[2].a/w1312 ), .B(n7393), .Z(n8236)
         );
  XOR \SUBBYTES[2].a/U5262  ( .A(\SUBBYTES[2].a/w1295 ), .B(
        \SUBBYTES[2].a/w1298 ), .Z(n7393) );
  XOR \SUBBYTES[2].a/U5260  ( .A(\SUBBYTES[2].a/w1283 ), .B(n8238), .Z(n7394)
         );
  XOR \SUBBYTES[2].a/U5258  ( .A(\SUBBYTES[2].a/w1315 ), .B(
        \SUBBYTES[2].a/w1328 ), .Z(n7395) );
  XOR \SUBBYTES[2].a/U5256  ( .A(n7399), .B(n7398), .Z(n7396) );
  XOR \SUBBYTES[2].a/U5255  ( .A(n7401), .B(n7400), .Z(n7397) );
  XOR \SUBBYTES[2].a/U5254  ( .A(\SUBBYTES[2].a/w1327 ), .B(
        \SUBBYTES[2].a/w1330 ), .Z(n7398) );
  XOR \SUBBYTES[2].a/U5253  ( .A(\SUBBYTES[2].a/w1320 ), .B(
        \SUBBYTES[2].a/w1323 ), .Z(n7399) );
  XOR \SUBBYTES[2].a/U5252  ( .A(\SUBBYTES[2].a/w1295 ), .B(
        \SUBBYTES[2].a/w1296 ), .Z(n7400) );
  XOR \SUBBYTES[2].a/U5251  ( .A(\SUBBYTES[2].a/w1280 ), .B(
        \SUBBYTES[2].a/w1283 ), .Z(n7401) );
  XOR \SUBBYTES[2].a/U5249  ( .A(n8235), .B(n7404), .Z(n7402) );
  XOR \SUBBYTES[2].a/U5248  ( .A(n8237), .B(n8236), .Z(n7403) );
  XOR \SUBBYTES[2].a/U5247  ( .A(\SUBBYTES[2].a/w1288 ), .B(
        \SUBBYTES[2].a/w1315 ), .Z(n7404) );
  XOR \SUBBYTES[2].a/U5245  ( .A(n8238), .B(n7407), .Z(n7405) );
  XOR \SUBBYTES[2].a/U5244  ( .A(\SUBBYTES[2].a/w1321 ), .B(
        \SUBBYTES[2].a/w1323 ), .Z(n7406) );
  XOR \SUBBYTES[2].a/U5243  ( .A(\SUBBYTES[2].a/w1281 ), .B(
        \SUBBYTES[2].a/w1313 ), .Z(n7407) );
  XOR \SUBBYTES[2].a/U5242  ( .A(\SUBBYTES[2].a/w1113 ), .B(
        \SUBBYTES[2].a/w1114 ), .Z(n8240) );
  XOR \SUBBYTES[2].a/U5241  ( .A(n8240), .B(n7408), .Z(n8239) );
  XOR \SUBBYTES[2].a/U5240  ( .A(\SUBBYTES[2].a/w1106 ), .B(
        \SUBBYTES[2].a/w1123 ), .Z(n7408) );
  XOR \SUBBYTES[2].a/U5238  ( .A(\SUBBYTES[2].a/w1105 ), .B(
        \SUBBYTES[2].a/w1120 ), .Z(n7409) );
  XOR \SUBBYTES[2].a/U5237  ( .A(n8240), .B(n7410), .Z(n8387) );
  XOR \SUBBYTES[2].a/U5236  ( .A(\SUBBYTES[2].a/w1120 ), .B(
        \SUBBYTES[2].a/w1121 ), .Z(n7410) );
  XOR \SUBBYTES[2].a/U5235  ( .A(\SUBBYTES[2].a/w1082 ), .B(n7411), .Z(n8242)
         );
  XOR \SUBBYTES[2].a/U5234  ( .A(\SUBBYTES[2].a/w1073 ), .B(
        \SUBBYTES[2].a/w1074 ), .Z(n7411) );
  XOR \SUBBYTES[2].a/U5232  ( .A(\SUBBYTES[2].a/w1084 ), .B(n8387), .Z(n7412)
         );
  XOR \SUBBYTES[2].a/U5231  ( .A(n7414), .B(n7413), .Z(n8243) );
  XOR \SUBBYTES[2].a/U5230  ( .A(n7416), .B(n7415), .Z(n7413) );
  XOR \SUBBYTES[2].a/U5229  ( .A(\SUBBYTES[2].a/w1120 ), .B(
        \SUBBYTES[2].a/w1121 ), .Z(n7414) );
  XOR \SUBBYTES[2].a/U5228  ( .A(\SUBBYTES[2].a/w1084 ), .B(
        \SUBBYTES[2].a/w1108 ), .Z(n7415) );
  XOR \SUBBYTES[2].a/U5227  ( .A(\SUBBYTES[2].a/w1073 ), .B(
        \SUBBYTES[2].a/w1082 ), .Z(n7416) );
  XOR \SUBBYTES[2].a/U5226  ( .A(\SUBBYTES[2].a/w1105 ), .B(n7417), .Z(n8241)
         );
  XOR \SUBBYTES[2].a/U5225  ( .A(\SUBBYTES[2].a/w1088 ), .B(
        \SUBBYTES[2].a/w1091 ), .Z(n7417) );
  XOR \SUBBYTES[2].a/U5223  ( .A(\SUBBYTES[2].a/w1076 ), .B(n8243), .Z(n7418)
         );
  XOR \SUBBYTES[2].a/U5221  ( .A(\SUBBYTES[2].a/w1108 ), .B(
        \SUBBYTES[2].a/w1121 ), .Z(n7419) );
  XOR \SUBBYTES[2].a/U5219  ( .A(n7423), .B(n7422), .Z(n7420) );
  XOR \SUBBYTES[2].a/U5218  ( .A(n7425), .B(n7424), .Z(n7421) );
  XOR \SUBBYTES[2].a/U5217  ( .A(\SUBBYTES[2].a/w1120 ), .B(
        \SUBBYTES[2].a/w1123 ), .Z(n7422) );
  XOR \SUBBYTES[2].a/U5216  ( .A(\SUBBYTES[2].a/w1113 ), .B(
        \SUBBYTES[2].a/w1116 ), .Z(n7423) );
  XOR \SUBBYTES[2].a/U5215  ( .A(\SUBBYTES[2].a/w1088 ), .B(
        \SUBBYTES[2].a/w1089 ), .Z(n7424) );
  XOR \SUBBYTES[2].a/U5214  ( .A(\SUBBYTES[2].a/w1073 ), .B(
        \SUBBYTES[2].a/w1076 ), .Z(n7425) );
  XOR \SUBBYTES[2].a/U5212  ( .A(n8240), .B(n7428), .Z(n7426) );
  XOR \SUBBYTES[2].a/U5211  ( .A(n8242), .B(n8241), .Z(n7427) );
  XOR \SUBBYTES[2].a/U5210  ( .A(\SUBBYTES[2].a/w1081 ), .B(
        \SUBBYTES[2].a/w1108 ), .Z(n7428) );
  XOR \SUBBYTES[2].a/U5208  ( .A(n8243), .B(n7431), .Z(n7429) );
  XOR \SUBBYTES[2].a/U5207  ( .A(\SUBBYTES[2].a/w1114 ), .B(
        \SUBBYTES[2].a/w1116 ), .Z(n7430) );
  XOR \SUBBYTES[2].a/U5206  ( .A(\SUBBYTES[2].a/w1074 ), .B(
        \SUBBYTES[2].a/w1106 ), .Z(n7431) );
  XOR \SUBBYTES[2].a/U5205  ( .A(\SUBBYTES[2].a/w906 ), .B(
        \SUBBYTES[2].a/w907 ), .Z(n8245) );
  XOR \SUBBYTES[2].a/U5204  ( .A(n8245), .B(n7432), .Z(n8244) );
  XOR \SUBBYTES[2].a/U5203  ( .A(\SUBBYTES[2].a/w899 ), .B(
        \SUBBYTES[2].a/w916 ), .Z(n7432) );
  XOR \SUBBYTES[2].a/U5201  ( .A(\SUBBYTES[2].a/w898 ), .B(
        \SUBBYTES[2].a/w913 ), .Z(n7433) );
  XOR \SUBBYTES[2].a/U5200  ( .A(n8245), .B(n7434), .Z(n8388) );
  XOR \SUBBYTES[2].a/U5199  ( .A(\SUBBYTES[2].a/w913 ), .B(
        \SUBBYTES[2].a/w914 ), .Z(n7434) );
  XOR \SUBBYTES[2].a/U5198  ( .A(\SUBBYTES[2].a/w875 ), .B(n7435), .Z(n8247)
         );
  XOR \SUBBYTES[2].a/U5197  ( .A(\SUBBYTES[2].a/w866 ), .B(
        \SUBBYTES[2].a/w867 ), .Z(n7435) );
  XOR \SUBBYTES[2].a/U5195  ( .A(\SUBBYTES[2].a/w877 ), .B(n8388), .Z(n7436)
         );
  XOR \SUBBYTES[2].a/U5194  ( .A(n7438), .B(n7437), .Z(n8248) );
  XOR \SUBBYTES[2].a/U5193  ( .A(n7440), .B(n7439), .Z(n7437) );
  XOR \SUBBYTES[2].a/U5192  ( .A(\SUBBYTES[2].a/w913 ), .B(
        \SUBBYTES[2].a/w914 ), .Z(n7438) );
  XOR \SUBBYTES[2].a/U5191  ( .A(\SUBBYTES[2].a/w877 ), .B(
        \SUBBYTES[2].a/w901 ), .Z(n7439) );
  XOR \SUBBYTES[2].a/U5190  ( .A(\SUBBYTES[2].a/w866 ), .B(
        \SUBBYTES[2].a/w875 ), .Z(n7440) );
  XOR \SUBBYTES[2].a/U5189  ( .A(\SUBBYTES[2].a/w898 ), .B(n7441), .Z(n8246)
         );
  XOR \SUBBYTES[2].a/U5188  ( .A(\SUBBYTES[2].a/w881 ), .B(
        \SUBBYTES[2].a/w884 ), .Z(n7441) );
  XOR \SUBBYTES[2].a/U5186  ( .A(\SUBBYTES[2].a/w869 ), .B(n8248), .Z(n7442)
         );
  XOR \SUBBYTES[2].a/U5184  ( .A(\SUBBYTES[2].a/w901 ), .B(
        \SUBBYTES[2].a/w914 ), .Z(n7443) );
  XOR \SUBBYTES[2].a/U5182  ( .A(n7447), .B(n7446), .Z(n7444) );
  XOR \SUBBYTES[2].a/U5181  ( .A(n7449), .B(n7448), .Z(n7445) );
  XOR \SUBBYTES[2].a/U5180  ( .A(\SUBBYTES[2].a/w913 ), .B(
        \SUBBYTES[2].a/w916 ), .Z(n7446) );
  XOR \SUBBYTES[2].a/U5179  ( .A(\SUBBYTES[2].a/w906 ), .B(
        \SUBBYTES[2].a/w909 ), .Z(n7447) );
  XOR \SUBBYTES[2].a/U5178  ( .A(\SUBBYTES[2].a/w881 ), .B(
        \SUBBYTES[2].a/w882 ), .Z(n7448) );
  XOR \SUBBYTES[2].a/U5177  ( .A(\SUBBYTES[2].a/w866 ), .B(
        \SUBBYTES[2].a/w869 ), .Z(n7449) );
  XOR \SUBBYTES[2].a/U5175  ( .A(n8245), .B(n7452), .Z(n7450) );
  XOR \SUBBYTES[2].a/U5174  ( .A(n8247), .B(n8246), .Z(n7451) );
  XOR \SUBBYTES[2].a/U5173  ( .A(\SUBBYTES[2].a/w874 ), .B(
        \SUBBYTES[2].a/w901 ), .Z(n7452) );
  XOR \SUBBYTES[2].a/U5171  ( .A(n8248), .B(n7455), .Z(n7453) );
  XOR \SUBBYTES[2].a/U5170  ( .A(\SUBBYTES[2].a/w907 ), .B(
        \SUBBYTES[2].a/w909 ), .Z(n7454) );
  XOR \SUBBYTES[2].a/U5169  ( .A(\SUBBYTES[2].a/w867 ), .B(
        \SUBBYTES[2].a/w899 ), .Z(n7455) );
  XOR \SUBBYTES[2].a/U5168  ( .A(\SUBBYTES[2].a/w699 ), .B(
        \SUBBYTES[2].a/w700 ), .Z(n8250) );
  XOR \SUBBYTES[2].a/U5167  ( .A(n8250), .B(n7456), .Z(n8249) );
  XOR \SUBBYTES[2].a/U5166  ( .A(\SUBBYTES[2].a/w692 ), .B(
        \SUBBYTES[2].a/w709 ), .Z(n7456) );
  XOR \SUBBYTES[2].a/U5164  ( .A(\SUBBYTES[2].a/w691 ), .B(
        \SUBBYTES[2].a/w706 ), .Z(n7457) );
  XOR \SUBBYTES[2].a/U5163  ( .A(n8250), .B(n7458), .Z(n8389) );
  XOR \SUBBYTES[2].a/U5162  ( .A(\SUBBYTES[2].a/w706 ), .B(
        \SUBBYTES[2].a/w707 ), .Z(n7458) );
  XOR \SUBBYTES[2].a/U5161  ( .A(\SUBBYTES[2].a/w668 ), .B(n7459), .Z(n8252)
         );
  XOR \SUBBYTES[2].a/U5160  ( .A(\SUBBYTES[2].a/w659 ), .B(
        \SUBBYTES[2].a/w660 ), .Z(n7459) );
  XOR \SUBBYTES[2].a/U5158  ( .A(\SUBBYTES[2].a/w670 ), .B(n8389), .Z(n7460)
         );
  XOR \SUBBYTES[2].a/U5157  ( .A(n7462), .B(n7461), .Z(n8253) );
  XOR \SUBBYTES[2].a/U5156  ( .A(n7464), .B(n7463), .Z(n7461) );
  XOR \SUBBYTES[2].a/U5155  ( .A(\SUBBYTES[2].a/w706 ), .B(
        \SUBBYTES[2].a/w707 ), .Z(n7462) );
  XOR \SUBBYTES[2].a/U5154  ( .A(\SUBBYTES[2].a/w670 ), .B(
        \SUBBYTES[2].a/w694 ), .Z(n7463) );
  XOR \SUBBYTES[2].a/U5153  ( .A(\SUBBYTES[2].a/w659 ), .B(
        \SUBBYTES[2].a/w668 ), .Z(n7464) );
  XOR \SUBBYTES[2].a/U5152  ( .A(\SUBBYTES[2].a/w691 ), .B(n7465), .Z(n8251)
         );
  XOR \SUBBYTES[2].a/U5151  ( .A(\SUBBYTES[2].a/w674 ), .B(
        \SUBBYTES[2].a/w677 ), .Z(n7465) );
  XOR \SUBBYTES[2].a/U5149  ( .A(\SUBBYTES[2].a/w662 ), .B(n8253), .Z(n7466)
         );
  XOR \SUBBYTES[2].a/U5147  ( .A(\SUBBYTES[2].a/w694 ), .B(
        \SUBBYTES[2].a/w707 ), .Z(n7467) );
  XOR \SUBBYTES[2].a/U5145  ( .A(n7471), .B(n7470), .Z(n7468) );
  XOR \SUBBYTES[2].a/U5144  ( .A(n7473), .B(n7472), .Z(n7469) );
  XOR \SUBBYTES[2].a/U5143  ( .A(\SUBBYTES[2].a/w706 ), .B(
        \SUBBYTES[2].a/w709 ), .Z(n7470) );
  XOR \SUBBYTES[2].a/U5142  ( .A(\SUBBYTES[2].a/w699 ), .B(
        \SUBBYTES[2].a/w702 ), .Z(n7471) );
  XOR \SUBBYTES[2].a/U5141  ( .A(\SUBBYTES[2].a/w674 ), .B(
        \SUBBYTES[2].a/w675 ), .Z(n7472) );
  XOR \SUBBYTES[2].a/U5140  ( .A(\SUBBYTES[2].a/w659 ), .B(
        \SUBBYTES[2].a/w662 ), .Z(n7473) );
  XOR \SUBBYTES[2].a/U5138  ( .A(n8250), .B(n7476), .Z(n7474) );
  XOR \SUBBYTES[2].a/U5137  ( .A(n8252), .B(n8251), .Z(n7475) );
  XOR \SUBBYTES[2].a/U5136  ( .A(\SUBBYTES[2].a/w667 ), .B(
        \SUBBYTES[2].a/w694 ), .Z(n7476) );
  XOR \SUBBYTES[2].a/U5134  ( .A(n8253), .B(n7479), .Z(n7477) );
  XOR \SUBBYTES[2].a/U5133  ( .A(\SUBBYTES[2].a/w700 ), .B(
        \SUBBYTES[2].a/w702 ), .Z(n7478) );
  XOR \SUBBYTES[2].a/U5132  ( .A(\SUBBYTES[2].a/w660 ), .B(
        \SUBBYTES[2].a/w692 ), .Z(n7479) );
  XOR \SUBBYTES[2].a/U5131  ( .A(\SUBBYTES[2].a/w492 ), .B(
        \SUBBYTES[2].a/w493 ), .Z(n8255) );
  XOR \SUBBYTES[2].a/U5130  ( .A(n8255), .B(n7480), .Z(n8254) );
  XOR \SUBBYTES[2].a/U5129  ( .A(\SUBBYTES[2].a/w485 ), .B(
        \SUBBYTES[2].a/w502 ), .Z(n7480) );
  XOR \SUBBYTES[2].a/U5127  ( .A(\SUBBYTES[2].a/w484 ), .B(
        \SUBBYTES[2].a/w499 ), .Z(n7481) );
  XOR \SUBBYTES[2].a/U5126  ( .A(n8255), .B(n7482), .Z(n8390) );
  XOR \SUBBYTES[2].a/U5125  ( .A(\SUBBYTES[2].a/w499 ), .B(
        \SUBBYTES[2].a/w500 ), .Z(n7482) );
  XOR \SUBBYTES[2].a/U5124  ( .A(\SUBBYTES[2].a/w461 ), .B(n7483), .Z(n8257)
         );
  XOR \SUBBYTES[2].a/U5123  ( .A(\SUBBYTES[2].a/w452 ), .B(
        \SUBBYTES[2].a/w453 ), .Z(n7483) );
  XOR \SUBBYTES[2].a/U5121  ( .A(\SUBBYTES[2].a/w463 ), .B(n8390), .Z(n7484)
         );
  XOR \SUBBYTES[2].a/U5120  ( .A(n7486), .B(n7485), .Z(n8258) );
  XOR \SUBBYTES[2].a/U5119  ( .A(n7488), .B(n7487), .Z(n7485) );
  XOR \SUBBYTES[2].a/U5118  ( .A(\SUBBYTES[2].a/w499 ), .B(
        \SUBBYTES[2].a/w500 ), .Z(n7486) );
  XOR \SUBBYTES[2].a/U5117  ( .A(\SUBBYTES[2].a/w463 ), .B(
        \SUBBYTES[2].a/w487 ), .Z(n7487) );
  XOR \SUBBYTES[2].a/U5116  ( .A(\SUBBYTES[2].a/w452 ), .B(
        \SUBBYTES[2].a/w461 ), .Z(n7488) );
  XOR \SUBBYTES[2].a/U5115  ( .A(\SUBBYTES[2].a/w484 ), .B(n7489), .Z(n8256)
         );
  XOR \SUBBYTES[2].a/U5114  ( .A(\SUBBYTES[2].a/w467 ), .B(
        \SUBBYTES[2].a/w470 ), .Z(n7489) );
  XOR \SUBBYTES[2].a/U5112  ( .A(\SUBBYTES[2].a/w455 ), .B(n8258), .Z(n7490)
         );
  XOR \SUBBYTES[2].a/U5110  ( .A(\SUBBYTES[2].a/w487 ), .B(
        \SUBBYTES[2].a/w500 ), .Z(n7491) );
  XOR \SUBBYTES[2].a/U5108  ( .A(n7495), .B(n7494), .Z(n7492) );
  XOR \SUBBYTES[2].a/U5107  ( .A(n7497), .B(n7496), .Z(n7493) );
  XOR \SUBBYTES[2].a/U5106  ( .A(\SUBBYTES[2].a/w499 ), .B(
        \SUBBYTES[2].a/w502 ), .Z(n7494) );
  XOR \SUBBYTES[2].a/U5105  ( .A(\SUBBYTES[2].a/w492 ), .B(
        \SUBBYTES[2].a/w495 ), .Z(n7495) );
  XOR \SUBBYTES[2].a/U5104  ( .A(\SUBBYTES[2].a/w467 ), .B(
        \SUBBYTES[2].a/w468 ), .Z(n7496) );
  XOR \SUBBYTES[2].a/U5103  ( .A(\SUBBYTES[2].a/w452 ), .B(
        \SUBBYTES[2].a/w455 ), .Z(n7497) );
  XOR \SUBBYTES[2].a/U5101  ( .A(n8255), .B(n7500), .Z(n7498) );
  XOR \SUBBYTES[2].a/U5100  ( .A(n8257), .B(n8256), .Z(n7499) );
  XOR \SUBBYTES[2].a/U5099  ( .A(\SUBBYTES[2].a/w460 ), .B(
        \SUBBYTES[2].a/w487 ), .Z(n7500) );
  XOR \SUBBYTES[2].a/U5097  ( .A(n8258), .B(n7503), .Z(n7501) );
  XOR \SUBBYTES[2].a/U5096  ( .A(\SUBBYTES[2].a/w493 ), .B(
        \SUBBYTES[2].a/w495 ), .Z(n7502) );
  XOR \SUBBYTES[2].a/U5095  ( .A(\SUBBYTES[2].a/w453 ), .B(
        \SUBBYTES[2].a/w485 ), .Z(n7503) );
  XOR \SUBBYTES[2].a/U5094  ( .A(\SUBBYTES[2].a/w285 ), .B(
        \SUBBYTES[2].a/w286 ), .Z(n8260) );
  XOR \SUBBYTES[2].a/U5093  ( .A(n8260), .B(n7504), .Z(n8259) );
  XOR \SUBBYTES[2].a/U5092  ( .A(\SUBBYTES[2].a/w278 ), .B(
        \SUBBYTES[2].a/w295 ), .Z(n7504) );
  XOR \SUBBYTES[2].a/U5090  ( .A(\SUBBYTES[2].a/w277 ), .B(
        \SUBBYTES[2].a/w292 ), .Z(n7505) );
  XOR \SUBBYTES[2].a/U5089  ( .A(n8260), .B(n7506), .Z(n8391) );
  XOR \SUBBYTES[2].a/U5088  ( .A(\SUBBYTES[2].a/w292 ), .B(
        \SUBBYTES[2].a/w293 ), .Z(n7506) );
  XOR \SUBBYTES[2].a/U5087  ( .A(\SUBBYTES[2].a/w254 ), .B(n7507), .Z(n8262)
         );
  XOR \SUBBYTES[2].a/U5086  ( .A(\SUBBYTES[2].a/w245 ), .B(
        \SUBBYTES[2].a/w246 ), .Z(n7507) );
  XOR \SUBBYTES[2].a/U5084  ( .A(\SUBBYTES[2].a/w256 ), .B(n8391), .Z(n7508)
         );
  XOR \SUBBYTES[2].a/U5083  ( .A(n7510), .B(n7509), .Z(n8263) );
  XOR \SUBBYTES[2].a/U5082  ( .A(n7512), .B(n7511), .Z(n7509) );
  XOR \SUBBYTES[2].a/U5081  ( .A(\SUBBYTES[2].a/w292 ), .B(
        \SUBBYTES[2].a/w293 ), .Z(n7510) );
  XOR \SUBBYTES[2].a/U5080  ( .A(\SUBBYTES[2].a/w256 ), .B(
        \SUBBYTES[2].a/w280 ), .Z(n7511) );
  XOR \SUBBYTES[2].a/U5079  ( .A(\SUBBYTES[2].a/w245 ), .B(
        \SUBBYTES[2].a/w254 ), .Z(n7512) );
  XOR \SUBBYTES[2].a/U5078  ( .A(\SUBBYTES[2].a/w277 ), .B(n7513), .Z(n8261)
         );
  XOR \SUBBYTES[2].a/U5077  ( .A(\SUBBYTES[2].a/w260 ), .B(
        \SUBBYTES[2].a/w263 ), .Z(n7513) );
  XOR \SUBBYTES[2].a/U5075  ( .A(\SUBBYTES[2].a/w248 ), .B(n8263), .Z(n7514)
         );
  XOR \SUBBYTES[2].a/U5073  ( .A(\SUBBYTES[2].a/w280 ), .B(
        \SUBBYTES[2].a/w293 ), .Z(n7515) );
  XOR \SUBBYTES[2].a/U5071  ( .A(n7519), .B(n7518), .Z(n7516) );
  XOR \SUBBYTES[2].a/U5070  ( .A(n7521), .B(n7520), .Z(n7517) );
  XOR \SUBBYTES[2].a/U5069  ( .A(\SUBBYTES[2].a/w292 ), .B(
        \SUBBYTES[2].a/w295 ), .Z(n7518) );
  XOR \SUBBYTES[2].a/U5068  ( .A(\SUBBYTES[2].a/w285 ), .B(
        \SUBBYTES[2].a/w288 ), .Z(n7519) );
  XOR \SUBBYTES[2].a/U5067  ( .A(\SUBBYTES[2].a/w260 ), .B(
        \SUBBYTES[2].a/w261 ), .Z(n7520) );
  XOR \SUBBYTES[2].a/U5066  ( .A(\SUBBYTES[2].a/w245 ), .B(
        \SUBBYTES[2].a/w248 ), .Z(n7521) );
  XOR \SUBBYTES[2].a/U5064  ( .A(n8260), .B(n7524), .Z(n7522) );
  XOR \SUBBYTES[2].a/U5063  ( .A(n8262), .B(n8261), .Z(n7523) );
  XOR \SUBBYTES[2].a/U5062  ( .A(\SUBBYTES[2].a/w253 ), .B(
        \SUBBYTES[2].a/w280 ), .Z(n7524) );
  XOR \SUBBYTES[2].a/U5060  ( .A(n8263), .B(n7527), .Z(n7525) );
  XOR \SUBBYTES[2].a/U5059  ( .A(\SUBBYTES[2].a/w286 ), .B(
        \SUBBYTES[2].a/w288 ), .Z(n7526) );
  XOR \SUBBYTES[2].a/U5058  ( .A(\SUBBYTES[2].a/w246 ), .B(
        \SUBBYTES[2].a/w278 ), .Z(n7527) );
  XOR \SUBBYTES[2].a/U5057  ( .A(\w1[2][1] ), .B(n7528), .Z(n8264) );
  XOR \SUBBYTES[2].a/U5056  ( .A(\w1[2][3] ), .B(\w1[2][2] ), .Z(n7528) );
  XOR \SUBBYTES[2].a/U5055  ( .A(\w1[2][6] ), .B(n8264), .Z(
        \SUBBYTES[2].a/w3378 ) );
  XOR \SUBBYTES[2].a/U5054  ( .A(\w1[2][0] ), .B(\SUBBYTES[2].a/w3378 ), .Z(
        \SUBBYTES[2].a/w3265 ) );
  XOR \SUBBYTES[2].a/U5053  ( .A(\w1[2][0] ), .B(n7529), .Z(
        \SUBBYTES[2].a/w3266 ) );
  XOR \SUBBYTES[2].a/U5052  ( .A(\w1[2][6] ), .B(\w1[2][5] ), .Z(n7529) );
  XOR \SUBBYTES[2].a/U5051  ( .A(\w1[2][5] ), .B(n8264), .Z(
        \SUBBYTES[2].a/w3396 ) );
  XOR \SUBBYTES[2].a/U5050  ( .A(n7531), .B(n7530), .Z(\SUBBYTES[2].a/w3389 )
         );
  XOR \SUBBYTES[2].a/U5049  ( .A(\w1[2][3] ), .B(\w1[2][1] ), .Z(n7530) );
  XOR \SUBBYTES[2].a/U5048  ( .A(\w1[2][7] ), .B(\w1[2][4] ), .Z(n7531) );
  XOR \SUBBYTES[2].a/U5047  ( .A(\w1[2][0] ), .B(\SUBBYTES[2].a/w3389 ), .Z(
        \SUBBYTES[2].a/w3268 ) );
  XOR \SUBBYTES[2].a/U5046  ( .A(n7533), .B(n7532), .Z(\SUBBYTES[2].a/w3376 )
         );
  XOR \SUBBYTES[2].a/U5045  ( .A(\SUBBYTES[2].a/w3337 ), .B(n988), .Z(n7532)
         );
  XOR \SUBBYTES[2].a/U5044  ( .A(\SUBBYTES[2].a/w3330 ), .B(
        \SUBBYTES[2].a/w3333 ), .Z(n7533) );
  XOR \SUBBYTES[2].a/U5043  ( .A(n7535), .B(n7534), .Z(\SUBBYTES[2].a/w3377 )
         );
  XOR \SUBBYTES[2].a/U5042  ( .A(\SUBBYTES[2].a/w3337 ), .B(n7143), .Z(n7534)
         );
  XOR \SUBBYTES[2].a/U5041  ( .A(\SUBBYTES[2].a/w3330 ), .B(n7142), .Z(n7535)
         );
  XOR \SUBBYTES[2].a/U5040  ( .A(\SUBBYTES[2].a/w3389 ), .B(n7536), .Z(
        \SUBBYTES[2].a/w3379 ) );
  XOR \SUBBYTES[2].a/U5039  ( .A(\w1[2][6] ), .B(\w1[2][5] ), .Z(n7536) );
  XOR \SUBBYTES[2].a/U5038  ( .A(n7538), .B(n7537), .Z(\SUBBYTES[2].a/w3380 )
         );
  XOR \SUBBYTES[2].a/U5037  ( .A(n7143), .B(n988), .Z(n7537) );
  XOR \SUBBYTES[2].a/U5036  ( .A(n7142), .B(\SUBBYTES[2].a/w3333 ), .Z(n7538)
         );
  XOR \SUBBYTES[2].a/U5035  ( .A(\w1[2][7] ), .B(\w1[2][2] ), .Z(n8270) );
  XOR \SUBBYTES[2].a/U5034  ( .A(n8270), .B(n7539), .Z(\SUBBYTES[2].a/w3381 )
         );
  XOR \SUBBYTES[2].a/U5033  ( .A(\w1[2][5] ), .B(\w1[2][4] ), .Z(n7539) );
  XOR \SUBBYTES[2].a/U5032  ( .A(\w1[2][7] ), .B(\SUBBYTES[2].a/w3266 ), .Z(
        \SUBBYTES[2].a/w3269 ) );
  XOR \SUBBYTES[2].a/U5031  ( .A(\w1[2][1] ), .B(\SUBBYTES[2].a/w3266 ), .Z(
        \SUBBYTES[2].a/w3270 ) );
  XOR \SUBBYTES[2].a/U5030  ( .A(\w1[2][4] ), .B(\SUBBYTES[2].a/w3266 ), .Z(
        \SUBBYTES[2].a/w3271 ) );
  XOR \SUBBYTES[2].a/U5029  ( .A(\SUBBYTES[2].a/w3270 ), .B(n8270), .Z(
        \SUBBYTES[2].a/w3272 ) );
  XOR \SUBBYTES[2].a/U5028  ( .A(n8270), .B(n7540), .Z(\SUBBYTES[2].a/w3357 )
         );
  XOR \SUBBYTES[2].a/U5027  ( .A(\w1[2][4] ), .B(\w1[2][1] ), .Z(n7540) );
  XOR \SUBBYTES[2].a/U5026  ( .A(n7542), .B(n7541), .Z(n8267) );
  XOR \SUBBYTES[2].a/U5025  ( .A(\w1[2][4] ), .B(n7543), .Z(n7541) );
  XOR \SUBBYTES[2].a/U5024  ( .A(\SUBBYTES[2].a/w3322 ), .B(\w1[2][6] ), .Z(
        n7542) );
  XOR \SUBBYTES[2].a/U5023  ( .A(\SUBBYTES[2].a/w3296 ), .B(
        \SUBBYTES[2].a/w3303 ), .Z(n7543) );
  XOR \SUBBYTES[2].a/U5022  ( .A(n7545), .B(n7544), .Z(n8265) );
  XOR \SUBBYTES[2].a/U5021  ( .A(\w1[2][1] ), .B(n7546), .Z(n7544) );
  XOR \SUBBYTES[2].a/U5020  ( .A(\SUBBYTES[2].a/w3321 ), .B(\w1[2][5] ), .Z(
        n7545) );
  XOR \SUBBYTES[2].a/U5019  ( .A(\SUBBYTES[2].a/w3297 ), .B(
        \SUBBYTES[2].a/w3304 ), .Z(n7546) );
  XOR \SUBBYTES[2].a/U5018  ( .A(n8267), .B(n8265), .Z(\SUBBYTES[2].a/w3327 )
         );
  XOR \SUBBYTES[2].a/U5017  ( .A(\w1[2][5] ), .B(n7547), .Z(n8268) );
  XOR \SUBBYTES[2].a/U5016  ( .A(\SUBBYTES[2].a/w3289 ), .B(
        \SUBBYTES[2].a/w3299 ), .Z(n7547) );
  XOR \SUBBYTES[2].a/U5015  ( .A(n7549), .B(n7548), .Z(\SUBBYTES[2].a/w3314 )
         );
  XOR \SUBBYTES[2].a/U5014  ( .A(n8268), .B(n7550), .Z(n7548) );
  XOR \SUBBYTES[2].a/U5013  ( .A(\w1[2][4] ), .B(\SUBBYTES[2].a/w3378 ), .Z(
        n7549) );
  XOR \SUBBYTES[2].a/U5012  ( .A(\SUBBYTES[2].a/w3291 ), .B(
        \SUBBYTES[2].a/w3296 ), .Z(n7550) );
  XOR \SUBBYTES[2].a/U5011  ( .A(n7552), .B(n7551), .Z(n8266) );
  XOR \SUBBYTES[2].a/U5010  ( .A(\SUBBYTES[2].a/w3324 ), .B(\w1[2][7] ), .Z(
        n7551) );
  XOR \SUBBYTES[2].a/U5009  ( .A(\SUBBYTES[2].a/w3299 ), .B(
        \SUBBYTES[2].a/w3306 ), .Z(n7552) );
  XOR \SUBBYTES[2].a/U5008  ( .A(n8265), .B(n8266), .Z(\SUBBYTES[2].a/w3326 )
         );
  XOR \SUBBYTES[2].a/U5007  ( .A(\w1[2][3] ), .B(n7553), .Z(n8269) );
  XOR \SUBBYTES[2].a/U5006  ( .A(\SUBBYTES[2].a/w3288 ), .B(
        \SUBBYTES[2].a/w3291 ), .Z(n7553) );
  XOR \SUBBYTES[2].a/U5005  ( .A(n7555), .B(n7554), .Z(\SUBBYTES[2].a/w3315 )
         );
  XOR \SUBBYTES[2].a/U5004  ( .A(n8269), .B(n7556), .Z(n7554) );
  XOR \SUBBYTES[2].a/U5003  ( .A(\w1[2][6] ), .B(\SUBBYTES[2].a/w3357 ), .Z(
        n7555) );
  XOR \SUBBYTES[2].a/U5002  ( .A(\SUBBYTES[2].a/w3296 ), .B(
        \SUBBYTES[2].a/w3297 ), .Z(n7556) );
  XOR \SUBBYTES[2].a/U5001  ( .A(n8267), .B(n8266), .Z(\SUBBYTES[2].a/w3335 )
         );
  XOR \SUBBYTES[2].a/U5000  ( .A(n7558), .B(n7557), .Z(\SUBBYTES[2].a/w3336 )
         );
  XOR \SUBBYTES[2].a/U4999  ( .A(\w1[2][7] ), .B(n8268), .Z(n7557) );
  XOR \SUBBYTES[2].a/U4998  ( .A(\SUBBYTES[2].a/w3288 ), .B(
        \SUBBYTES[2].a/w3297 ), .Z(n7558) );
  XOR \SUBBYTES[2].a/U4997  ( .A(n7560), .B(n7559), .Z(\SUBBYTES[2].a/w3312 )
         );
  XOR \SUBBYTES[2].a/U4996  ( .A(n7562), .B(n7561), .Z(n7559) );
  XOR \SUBBYTES[2].a/U4995  ( .A(\w1[2][7] ), .B(\SUBBYTES[2].a/w3396 ), .Z(
        n7560) );
  XOR \SUBBYTES[2].a/U4994  ( .A(\SUBBYTES[2].a/w3303 ), .B(
        \SUBBYTES[2].a/w3306 ), .Z(n7561) );
  XOR \SUBBYTES[2].a/U4993  ( .A(\SUBBYTES[2].a/w3289 ), .B(
        \SUBBYTES[2].a/w3291 ), .Z(n7562) );
  XOR \SUBBYTES[2].a/U4992  ( .A(n7564), .B(n7563), .Z(\SUBBYTES[2].a/w3313 )
         );
  XOR \SUBBYTES[2].a/U4991  ( .A(n8269), .B(n7565), .Z(n7563) );
  XOR \SUBBYTES[2].a/U4990  ( .A(\w1[2][5] ), .B(n8270), .Z(n7564) );
  XOR \SUBBYTES[2].a/U4989  ( .A(\SUBBYTES[2].a/w3303 ), .B(
        \SUBBYTES[2].a/w3304 ), .Z(n7565) );
  XOR \SUBBYTES[2].a/U4988  ( .A(n7567), .B(n7566), .Z(\SUBBYTES[2].a/w3329 )
         );
  XOR \SUBBYTES[2].a/U4987  ( .A(\w1[2][1] ), .B(n7568), .Z(n7566) );
  XOR \SUBBYTES[2].a/U4986  ( .A(\SUBBYTES[2].a/w3304 ), .B(
        \SUBBYTES[2].a/w3306 ), .Z(n7567) );
  XOR \SUBBYTES[2].a/U4985  ( .A(\SUBBYTES[2].a/w3288 ), .B(
        \SUBBYTES[2].a/w3289 ), .Z(n7568) );
  XOR \SUBBYTES[2].a/U4984  ( .A(\w1[2][9] ), .B(n7569), .Z(n8271) );
  XOR \SUBBYTES[2].a/U4983  ( .A(\w1[2][11] ), .B(\w1[2][10] ), .Z(n7569) );
  XOR \SUBBYTES[2].a/U4982  ( .A(\w1[2][14] ), .B(n8271), .Z(
        \SUBBYTES[2].a/w3171 ) );
  XOR \SUBBYTES[2].a/U4981  ( .A(\w1[2][8] ), .B(\SUBBYTES[2].a/w3171 ), .Z(
        \SUBBYTES[2].a/w3058 ) );
  XOR \SUBBYTES[2].a/U4980  ( .A(\w1[2][8] ), .B(n7570), .Z(
        \SUBBYTES[2].a/w3059 ) );
  XOR \SUBBYTES[2].a/U4979  ( .A(\w1[2][14] ), .B(\w1[2][13] ), .Z(n7570) );
  XOR \SUBBYTES[2].a/U4978  ( .A(\w1[2][13] ), .B(n8271), .Z(
        \SUBBYTES[2].a/w3189 ) );
  XOR \SUBBYTES[2].a/U4977  ( .A(n7572), .B(n7571), .Z(\SUBBYTES[2].a/w3182 )
         );
  XOR \SUBBYTES[2].a/U4976  ( .A(\w1[2][11] ), .B(\w1[2][9] ), .Z(n7571) );
  XOR \SUBBYTES[2].a/U4975  ( .A(\w1[2][15] ), .B(\w1[2][12] ), .Z(n7572) );
  XOR \SUBBYTES[2].a/U4974  ( .A(\w1[2][8] ), .B(\SUBBYTES[2].a/w3182 ), .Z(
        \SUBBYTES[2].a/w3061 ) );
  XOR \SUBBYTES[2].a/U4973  ( .A(n7574), .B(n7573), .Z(\SUBBYTES[2].a/w3169 )
         );
  XOR \SUBBYTES[2].a/U4972  ( .A(\SUBBYTES[2].a/w3130 ), .B(n987), .Z(n7573)
         );
  XOR \SUBBYTES[2].a/U4971  ( .A(\SUBBYTES[2].a/w3123 ), .B(
        \SUBBYTES[2].a/w3126 ), .Z(n7574) );
  XOR \SUBBYTES[2].a/U4970  ( .A(n7576), .B(n7575), .Z(\SUBBYTES[2].a/w3170 )
         );
  XOR \SUBBYTES[2].a/U4969  ( .A(\SUBBYTES[2].a/w3130 ), .B(n7141), .Z(n7575)
         );
  XOR \SUBBYTES[2].a/U4968  ( .A(\SUBBYTES[2].a/w3123 ), .B(n7140), .Z(n7576)
         );
  XOR \SUBBYTES[2].a/U4967  ( .A(\SUBBYTES[2].a/w3182 ), .B(n7577), .Z(
        \SUBBYTES[2].a/w3172 ) );
  XOR \SUBBYTES[2].a/U4966  ( .A(\w1[2][14] ), .B(\w1[2][13] ), .Z(n7577) );
  XOR \SUBBYTES[2].a/U4965  ( .A(n7579), .B(n7578), .Z(\SUBBYTES[2].a/w3173 )
         );
  XOR \SUBBYTES[2].a/U4964  ( .A(n7141), .B(n987), .Z(n7578) );
  XOR \SUBBYTES[2].a/U4963  ( .A(n7140), .B(\SUBBYTES[2].a/w3126 ), .Z(n7579)
         );
  XOR \SUBBYTES[2].a/U4962  ( .A(\w1[2][15] ), .B(\w1[2][10] ), .Z(n8277) );
  XOR \SUBBYTES[2].a/U4961  ( .A(n8277), .B(n7580), .Z(\SUBBYTES[2].a/w3174 )
         );
  XOR \SUBBYTES[2].a/U4960  ( .A(\w1[2][13] ), .B(\w1[2][12] ), .Z(n7580) );
  XOR \SUBBYTES[2].a/U4959  ( .A(\w1[2][15] ), .B(\SUBBYTES[2].a/w3059 ), .Z(
        \SUBBYTES[2].a/w3062 ) );
  XOR \SUBBYTES[2].a/U4958  ( .A(\w1[2][9] ), .B(\SUBBYTES[2].a/w3059 ), .Z(
        \SUBBYTES[2].a/w3063 ) );
  XOR \SUBBYTES[2].a/U4957  ( .A(\w1[2][12] ), .B(\SUBBYTES[2].a/w3059 ), .Z(
        \SUBBYTES[2].a/w3064 ) );
  XOR \SUBBYTES[2].a/U4956  ( .A(\SUBBYTES[2].a/w3063 ), .B(n8277), .Z(
        \SUBBYTES[2].a/w3065 ) );
  XOR \SUBBYTES[2].a/U4955  ( .A(n8277), .B(n7581), .Z(\SUBBYTES[2].a/w3150 )
         );
  XOR \SUBBYTES[2].a/U4954  ( .A(\w1[2][12] ), .B(\w1[2][9] ), .Z(n7581) );
  XOR \SUBBYTES[2].a/U4953  ( .A(n7583), .B(n7582), .Z(n8274) );
  XOR \SUBBYTES[2].a/U4952  ( .A(\w1[2][12] ), .B(n7584), .Z(n7582) );
  XOR \SUBBYTES[2].a/U4951  ( .A(\SUBBYTES[2].a/w3115 ), .B(\w1[2][14] ), .Z(
        n7583) );
  XOR \SUBBYTES[2].a/U4950  ( .A(\SUBBYTES[2].a/w3089 ), .B(
        \SUBBYTES[2].a/w3096 ), .Z(n7584) );
  XOR \SUBBYTES[2].a/U4949  ( .A(n7586), .B(n7585), .Z(n8272) );
  XOR \SUBBYTES[2].a/U4948  ( .A(\w1[2][9] ), .B(n7587), .Z(n7585) );
  XOR \SUBBYTES[2].a/U4947  ( .A(\SUBBYTES[2].a/w3114 ), .B(\w1[2][13] ), .Z(
        n7586) );
  XOR \SUBBYTES[2].a/U4946  ( .A(\SUBBYTES[2].a/w3090 ), .B(
        \SUBBYTES[2].a/w3097 ), .Z(n7587) );
  XOR \SUBBYTES[2].a/U4945  ( .A(n8274), .B(n8272), .Z(\SUBBYTES[2].a/w3120 )
         );
  XOR \SUBBYTES[2].a/U4944  ( .A(\w1[2][13] ), .B(n7588), .Z(n8275) );
  XOR \SUBBYTES[2].a/U4943  ( .A(\SUBBYTES[2].a/w3082 ), .B(
        \SUBBYTES[2].a/w3092 ), .Z(n7588) );
  XOR \SUBBYTES[2].a/U4942  ( .A(n7590), .B(n7589), .Z(\SUBBYTES[2].a/w3107 )
         );
  XOR \SUBBYTES[2].a/U4941  ( .A(n8275), .B(n7591), .Z(n7589) );
  XOR \SUBBYTES[2].a/U4940  ( .A(\w1[2][12] ), .B(\SUBBYTES[2].a/w3171 ), .Z(
        n7590) );
  XOR \SUBBYTES[2].a/U4939  ( .A(\SUBBYTES[2].a/w3084 ), .B(
        \SUBBYTES[2].a/w3089 ), .Z(n7591) );
  XOR \SUBBYTES[2].a/U4938  ( .A(n7593), .B(n7592), .Z(n8273) );
  XOR \SUBBYTES[2].a/U4937  ( .A(\SUBBYTES[2].a/w3117 ), .B(\w1[2][15] ), .Z(
        n7592) );
  XOR \SUBBYTES[2].a/U4936  ( .A(\SUBBYTES[2].a/w3092 ), .B(
        \SUBBYTES[2].a/w3099 ), .Z(n7593) );
  XOR \SUBBYTES[2].a/U4935  ( .A(n8272), .B(n8273), .Z(\SUBBYTES[2].a/w3119 )
         );
  XOR \SUBBYTES[2].a/U4934  ( .A(\w1[2][11] ), .B(n7594), .Z(n8276) );
  XOR \SUBBYTES[2].a/U4933  ( .A(\SUBBYTES[2].a/w3081 ), .B(
        \SUBBYTES[2].a/w3084 ), .Z(n7594) );
  XOR \SUBBYTES[2].a/U4932  ( .A(n7596), .B(n7595), .Z(\SUBBYTES[2].a/w3108 )
         );
  XOR \SUBBYTES[2].a/U4931  ( .A(n8276), .B(n7597), .Z(n7595) );
  XOR \SUBBYTES[2].a/U4930  ( .A(\w1[2][14] ), .B(\SUBBYTES[2].a/w3150 ), .Z(
        n7596) );
  XOR \SUBBYTES[2].a/U4929  ( .A(\SUBBYTES[2].a/w3089 ), .B(
        \SUBBYTES[2].a/w3090 ), .Z(n7597) );
  XOR \SUBBYTES[2].a/U4928  ( .A(n8274), .B(n8273), .Z(\SUBBYTES[2].a/w3128 )
         );
  XOR \SUBBYTES[2].a/U4927  ( .A(n7599), .B(n7598), .Z(\SUBBYTES[2].a/w3129 )
         );
  XOR \SUBBYTES[2].a/U4926  ( .A(\w1[2][15] ), .B(n8275), .Z(n7598) );
  XOR \SUBBYTES[2].a/U4925  ( .A(\SUBBYTES[2].a/w3081 ), .B(
        \SUBBYTES[2].a/w3090 ), .Z(n7599) );
  XOR \SUBBYTES[2].a/U4924  ( .A(n7601), .B(n7600), .Z(\SUBBYTES[2].a/w3105 )
         );
  XOR \SUBBYTES[2].a/U4923  ( .A(n7603), .B(n7602), .Z(n7600) );
  XOR \SUBBYTES[2].a/U4922  ( .A(\w1[2][15] ), .B(\SUBBYTES[2].a/w3189 ), .Z(
        n7601) );
  XOR \SUBBYTES[2].a/U4921  ( .A(\SUBBYTES[2].a/w3096 ), .B(
        \SUBBYTES[2].a/w3099 ), .Z(n7602) );
  XOR \SUBBYTES[2].a/U4920  ( .A(\SUBBYTES[2].a/w3082 ), .B(
        \SUBBYTES[2].a/w3084 ), .Z(n7603) );
  XOR \SUBBYTES[2].a/U4919  ( .A(n7605), .B(n7604), .Z(\SUBBYTES[2].a/w3106 )
         );
  XOR \SUBBYTES[2].a/U4918  ( .A(n8276), .B(n7606), .Z(n7604) );
  XOR \SUBBYTES[2].a/U4917  ( .A(\w1[2][13] ), .B(n8277), .Z(n7605) );
  XOR \SUBBYTES[2].a/U4916  ( .A(\SUBBYTES[2].a/w3096 ), .B(
        \SUBBYTES[2].a/w3097 ), .Z(n7606) );
  XOR \SUBBYTES[2].a/U4915  ( .A(n7608), .B(n7607), .Z(\SUBBYTES[2].a/w3122 )
         );
  XOR \SUBBYTES[2].a/U4914  ( .A(\w1[2][9] ), .B(n7609), .Z(n7607) );
  XOR \SUBBYTES[2].a/U4913  ( .A(\SUBBYTES[2].a/w3097 ), .B(
        \SUBBYTES[2].a/w3099 ), .Z(n7608) );
  XOR \SUBBYTES[2].a/U4912  ( .A(\SUBBYTES[2].a/w3081 ), .B(
        \SUBBYTES[2].a/w3082 ), .Z(n7609) );
  XOR \SUBBYTES[2].a/U4911  ( .A(\w1[2][17] ), .B(n7610), .Z(n8278) );
  XOR \SUBBYTES[2].a/U4910  ( .A(\w1[2][19] ), .B(\w1[2][18] ), .Z(n7610) );
  XOR \SUBBYTES[2].a/U4909  ( .A(\w1[2][22] ), .B(n8278), .Z(
        \SUBBYTES[2].a/w2964 ) );
  XOR \SUBBYTES[2].a/U4908  ( .A(\w1[2][16] ), .B(\SUBBYTES[2].a/w2964 ), .Z(
        \SUBBYTES[2].a/w2851 ) );
  XOR \SUBBYTES[2].a/U4907  ( .A(\w1[2][16] ), .B(n7611), .Z(
        \SUBBYTES[2].a/w2852 ) );
  XOR \SUBBYTES[2].a/U4906  ( .A(\w1[2][22] ), .B(\w1[2][21] ), .Z(n7611) );
  XOR \SUBBYTES[2].a/U4905  ( .A(\w1[2][21] ), .B(n8278), .Z(
        \SUBBYTES[2].a/w2982 ) );
  XOR \SUBBYTES[2].a/U4904  ( .A(n7613), .B(n7612), .Z(\SUBBYTES[2].a/w2975 )
         );
  XOR \SUBBYTES[2].a/U4903  ( .A(\w1[2][19] ), .B(\w1[2][17] ), .Z(n7612) );
  XOR \SUBBYTES[2].a/U4902  ( .A(\w1[2][23] ), .B(\w1[2][20] ), .Z(n7613) );
  XOR \SUBBYTES[2].a/U4901  ( .A(\w1[2][16] ), .B(\SUBBYTES[2].a/w2975 ), .Z(
        \SUBBYTES[2].a/w2854 ) );
  XOR \SUBBYTES[2].a/U4900  ( .A(n7615), .B(n7614), .Z(\SUBBYTES[2].a/w2962 )
         );
  XOR \SUBBYTES[2].a/U4899  ( .A(\SUBBYTES[2].a/w2923 ), .B(n986), .Z(n7614)
         );
  XOR \SUBBYTES[2].a/U4898  ( .A(\SUBBYTES[2].a/w2916 ), .B(
        \SUBBYTES[2].a/w2919 ), .Z(n7615) );
  XOR \SUBBYTES[2].a/U4897  ( .A(n7617), .B(n7616), .Z(\SUBBYTES[2].a/w2963 )
         );
  XOR \SUBBYTES[2].a/U4896  ( .A(\SUBBYTES[2].a/w2923 ), .B(n7139), .Z(n7616)
         );
  XOR \SUBBYTES[2].a/U4895  ( .A(\SUBBYTES[2].a/w2916 ), .B(n7138), .Z(n7617)
         );
  XOR \SUBBYTES[2].a/U4894  ( .A(\SUBBYTES[2].a/w2975 ), .B(n7618), .Z(
        \SUBBYTES[2].a/w2965 ) );
  XOR \SUBBYTES[2].a/U4893  ( .A(\w1[2][22] ), .B(\w1[2][21] ), .Z(n7618) );
  XOR \SUBBYTES[2].a/U4892  ( .A(n7620), .B(n7619), .Z(\SUBBYTES[2].a/w2966 )
         );
  XOR \SUBBYTES[2].a/U4891  ( .A(n7139), .B(n986), .Z(n7619) );
  XOR \SUBBYTES[2].a/U4890  ( .A(n7138), .B(\SUBBYTES[2].a/w2919 ), .Z(n7620)
         );
  XOR \SUBBYTES[2].a/U4889  ( .A(\w1[2][23] ), .B(\w1[2][18] ), .Z(n8284) );
  XOR \SUBBYTES[2].a/U4888  ( .A(n8284), .B(n7621), .Z(\SUBBYTES[2].a/w2967 )
         );
  XOR \SUBBYTES[2].a/U4887  ( .A(\w1[2][21] ), .B(\w1[2][20] ), .Z(n7621) );
  XOR \SUBBYTES[2].a/U4886  ( .A(\w1[2][23] ), .B(\SUBBYTES[2].a/w2852 ), .Z(
        \SUBBYTES[2].a/w2855 ) );
  XOR \SUBBYTES[2].a/U4885  ( .A(\w1[2][17] ), .B(\SUBBYTES[2].a/w2852 ), .Z(
        \SUBBYTES[2].a/w2856 ) );
  XOR \SUBBYTES[2].a/U4884  ( .A(\w1[2][20] ), .B(\SUBBYTES[2].a/w2852 ), .Z(
        \SUBBYTES[2].a/w2857 ) );
  XOR \SUBBYTES[2].a/U4883  ( .A(\SUBBYTES[2].a/w2856 ), .B(n8284), .Z(
        \SUBBYTES[2].a/w2858 ) );
  XOR \SUBBYTES[2].a/U4882  ( .A(n8284), .B(n7622), .Z(\SUBBYTES[2].a/w2943 )
         );
  XOR \SUBBYTES[2].a/U4881  ( .A(\w1[2][20] ), .B(\w1[2][17] ), .Z(n7622) );
  XOR \SUBBYTES[2].a/U4880  ( .A(n7624), .B(n7623), .Z(n8281) );
  XOR \SUBBYTES[2].a/U4879  ( .A(\w1[2][20] ), .B(n7625), .Z(n7623) );
  XOR \SUBBYTES[2].a/U4878  ( .A(\SUBBYTES[2].a/w2908 ), .B(\w1[2][22] ), .Z(
        n7624) );
  XOR \SUBBYTES[2].a/U4877  ( .A(\SUBBYTES[2].a/w2882 ), .B(
        \SUBBYTES[2].a/w2889 ), .Z(n7625) );
  XOR \SUBBYTES[2].a/U4876  ( .A(n7627), .B(n7626), .Z(n8279) );
  XOR \SUBBYTES[2].a/U4875  ( .A(\w1[2][17] ), .B(n7628), .Z(n7626) );
  XOR \SUBBYTES[2].a/U4874  ( .A(\SUBBYTES[2].a/w2907 ), .B(\w1[2][21] ), .Z(
        n7627) );
  XOR \SUBBYTES[2].a/U4873  ( .A(\SUBBYTES[2].a/w2883 ), .B(
        \SUBBYTES[2].a/w2890 ), .Z(n7628) );
  XOR \SUBBYTES[2].a/U4872  ( .A(n8281), .B(n8279), .Z(\SUBBYTES[2].a/w2913 )
         );
  XOR \SUBBYTES[2].a/U4871  ( .A(\w1[2][21] ), .B(n7629), .Z(n8282) );
  XOR \SUBBYTES[2].a/U4870  ( .A(\SUBBYTES[2].a/w2875 ), .B(
        \SUBBYTES[2].a/w2885 ), .Z(n7629) );
  XOR \SUBBYTES[2].a/U4869  ( .A(n7631), .B(n7630), .Z(\SUBBYTES[2].a/w2900 )
         );
  XOR \SUBBYTES[2].a/U4868  ( .A(n8282), .B(n7632), .Z(n7630) );
  XOR \SUBBYTES[2].a/U4867  ( .A(\w1[2][20] ), .B(\SUBBYTES[2].a/w2964 ), .Z(
        n7631) );
  XOR \SUBBYTES[2].a/U4866  ( .A(\SUBBYTES[2].a/w2877 ), .B(
        \SUBBYTES[2].a/w2882 ), .Z(n7632) );
  XOR \SUBBYTES[2].a/U4865  ( .A(n7634), .B(n7633), .Z(n8280) );
  XOR \SUBBYTES[2].a/U4864  ( .A(\SUBBYTES[2].a/w2910 ), .B(\w1[2][23] ), .Z(
        n7633) );
  XOR \SUBBYTES[2].a/U4863  ( .A(\SUBBYTES[2].a/w2885 ), .B(
        \SUBBYTES[2].a/w2892 ), .Z(n7634) );
  XOR \SUBBYTES[2].a/U4862  ( .A(n8279), .B(n8280), .Z(\SUBBYTES[2].a/w2912 )
         );
  XOR \SUBBYTES[2].a/U4861  ( .A(\w1[2][19] ), .B(n7635), .Z(n8283) );
  XOR \SUBBYTES[2].a/U4860  ( .A(\SUBBYTES[2].a/w2874 ), .B(
        \SUBBYTES[2].a/w2877 ), .Z(n7635) );
  XOR \SUBBYTES[2].a/U4859  ( .A(n7637), .B(n7636), .Z(\SUBBYTES[2].a/w2901 )
         );
  XOR \SUBBYTES[2].a/U4858  ( .A(n8283), .B(n7638), .Z(n7636) );
  XOR \SUBBYTES[2].a/U4857  ( .A(\w1[2][22] ), .B(\SUBBYTES[2].a/w2943 ), .Z(
        n7637) );
  XOR \SUBBYTES[2].a/U4856  ( .A(\SUBBYTES[2].a/w2882 ), .B(
        \SUBBYTES[2].a/w2883 ), .Z(n7638) );
  XOR \SUBBYTES[2].a/U4855  ( .A(n8281), .B(n8280), .Z(\SUBBYTES[2].a/w2921 )
         );
  XOR \SUBBYTES[2].a/U4854  ( .A(n7640), .B(n7639), .Z(\SUBBYTES[2].a/w2922 )
         );
  XOR \SUBBYTES[2].a/U4853  ( .A(\w1[2][23] ), .B(n8282), .Z(n7639) );
  XOR \SUBBYTES[2].a/U4852  ( .A(\SUBBYTES[2].a/w2874 ), .B(
        \SUBBYTES[2].a/w2883 ), .Z(n7640) );
  XOR \SUBBYTES[2].a/U4851  ( .A(n7642), .B(n7641), .Z(\SUBBYTES[2].a/w2898 )
         );
  XOR \SUBBYTES[2].a/U4850  ( .A(n7644), .B(n7643), .Z(n7641) );
  XOR \SUBBYTES[2].a/U4849  ( .A(\w1[2][23] ), .B(\SUBBYTES[2].a/w2982 ), .Z(
        n7642) );
  XOR \SUBBYTES[2].a/U4848  ( .A(\SUBBYTES[2].a/w2889 ), .B(
        \SUBBYTES[2].a/w2892 ), .Z(n7643) );
  XOR \SUBBYTES[2].a/U4847  ( .A(\SUBBYTES[2].a/w2875 ), .B(
        \SUBBYTES[2].a/w2877 ), .Z(n7644) );
  XOR \SUBBYTES[2].a/U4846  ( .A(n7646), .B(n7645), .Z(\SUBBYTES[2].a/w2899 )
         );
  XOR \SUBBYTES[2].a/U4845  ( .A(n8283), .B(n7647), .Z(n7645) );
  XOR \SUBBYTES[2].a/U4844  ( .A(\w1[2][21] ), .B(n8284), .Z(n7646) );
  XOR \SUBBYTES[2].a/U4843  ( .A(\SUBBYTES[2].a/w2889 ), .B(
        \SUBBYTES[2].a/w2890 ), .Z(n7647) );
  XOR \SUBBYTES[2].a/U4842  ( .A(n7649), .B(n7648), .Z(\SUBBYTES[2].a/w2915 )
         );
  XOR \SUBBYTES[2].a/U4841  ( .A(\w1[2][17] ), .B(n7650), .Z(n7648) );
  XOR \SUBBYTES[2].a/U4840  ( .A(\SUBBYTES[2].a/w2890 ), .B(
        \SUBBYTES[2].a/w2892 ), .Z(n7649) );
  XOR \SUBBYTES[2].a/U4839  ( .A(\SUBBYTES[2].a/w2874 ), .B(
        \SUBBYTES[2].a/w2875 ), .Z(n7650) );
  XOR \SUBBYTES[2].a/U4838  ( .A(\w1[2][25] ), .B(n7651), .Z(n8285) );
  XOR \SUBBYTES[2].a/U4837  ( .A(\w1[2][27] ), .B(\w1[2][26] ), .Z(n7651) );
  XOR \SUBBYTES[2].a/U4836  ( .A(\w1[2][30] ), .B(n8285), .Z(
        \SUBBYTES[2].a/w2757 ) );
  XOR \SUBBYTES[2].a/U4835  ( .A(\w1[2][24] ), .B(\SUBBYTES[2].a/w2757 ), .Z(
        \SUBBYTES[2].a/w2644 ) );
  XOR \SUBBYTES[2].a/U4834  ( .A(\w1[2][24] ), .B(n7652), .Z(
        \SUBBYTES[2].a/w2645 ) );
  XOR \SUBBYTES[2].a/U4833  ( .A(\w1[2][30] ), .B(\w1[2][29] ), .Z(n7652) );
  XOR \SUBBYTES[2].a/U4832  ( .A(\w1[2][29] ), .B(n8285), .Z(
        \SUBBYTES[2].a/w2775 ) );
  XOR \SUBBYTES[2].a/U4831  ( .A(n7654), .B(n7653), .Z(\SUBBYTES[2].a/w2768 )
         );
  XOR \SUBBYTES[2].a/U4830  ( .A(\w1[2][27] ), .B(\w1[2][25] ), .Z(n7653) );
  XOR \SUBBYTES[2].a/U4829  ( .A(\w1[2][31] ), .B(\w1[2][28] ), .Z(n7654) );
  XOR \SUBBYTES[2].a/U4828  ( .A(\w1[2][24] ), .B(\SUBBYTES[2].a/w2768 ), .Z(
        \SUBBYTES[2].a/w2647 ) );
  XOR \SUBBYTES[2].a/U4827  ( .A(n7656), .B(n7655), .Z(\SUBBYTES[2].a/w2755 )
         );
  XOR \SUBBYTES[2].a/U4826  ( .A(\SUBBYTES[2].a/w2716 ), .B(n985), .Z(n7655)
         );
  XOR \SUBBYTES[2].a/U4825  ( .A(\SUBBYTES[2].a/w2709 ), .B(
        \SUBBYTES[2].a/w2712 ), .Z(n7656) );
  XOR \SUBBYTES[2].a/U4824  ( .A(n7658), .B(n7657), .Z(\SUBBYTES[2].a/w2756 )
         );
  XOR \SUBBYTES[2].a/U4823  ( .A(\SUBBYTES[2].a/w2716 ), .B(n7137), .Z(n7657)
         );
  XOR \SUBBYTES[2].a/U4822  ( .A(\SUBBYTES[2].a/w2709 ), .B(n7136), .Z(n7658)
         );
  XOR \SUBBYTES[2].a/U4821  ( .A(\SUBBYTES[2].a/w2768 ), .B(n7659), .Z(
        \SUBBYTES[2].a/w2758 ) );
  XOR \SUBBYTES[2].a/U4820  ( .A(\w1[2][30] ), .B(\w1[2][29] ), .Z(n7659) );
  XOR \SUBBYTES[2].a/U4819  ( .A(n7661), .B(n7660), .Z(\SUBBYTES[2].a/w2759 )
         );
  XOR \SUBBYTES[2].a/U4818  ( .A(n7137), .B(n985), .Z(n7660) );
  XOR \SUBBYTES[2].a/U4817  ( .A(n7136), .B(\SUBBYTES[2].a/w2712 ), .Z(n7661)
         );
  XOR \SUBBYTES[2].a/U4816  ( .A(\w1[2][31] ), .B(\w1[2][26] ), .Z(n8291) );
  XOR \SUBBYTES[2].a/U4815  ( .A(n8291), .B(n7662), .Z(\SUBBYTES[2].a/w2760 )
         );
  XOR \SUBBYTES[2].a/U4814  ( .A(\w1[2][29] ), .B(\w1[2][28] ), .Z(n7662) );
  XOR \SUBBYTES[2].a/U4813  ( .A(\w1[2][31] ), .B(\SUBBYTES[2].a/w2645 ), .Z(
        \SUBBYTES[2].a/w2648 ) );
  XOR \SUBBYTES[2].a/U4812  ( .A(\w1[2][25] ), .B(\SUBBYTES[2].a/w2645 ), .Z(
        \SUBBYTES[2].a/w2649 ) );
  XOR \SUBBYTES[2].a/U4811  ( .A(\w1[2][28] ), .B(\SUBBYTES[2].a/w2645 ), .Z(
        \SUBBYTES[2].a/w2650 ) );
  XOR \SUBBYTES[2].a/U4810  ( .A(\SUBBYTES[2].a/w2649 ), .B(n8291), .Z(
        \SUBBYTES[2].a/w2651 ) );
  XOR \SUBBYTES[2].a/U4809  ( .A(n8291), .B(n7663), .Z(\SUBBYTES[2].a/w2736 )
         );
  XOR \SUBBYTES[2].a/U4808  ( .A(\w1[2][28] ), .B(\w1[2][25] ), .Z(n7663) );
  XOR \SUBBYTES[2].a/U4807  ( .A(n7665), .B(n7664), .Z(n8288) );
  XOR \SUBBYTES[2].a/U4806  ( .A(\w1[2][28] ), .B(n7666), .Z(n7664) );
  XOR \SUBBYTES[2].a/U4805  ( .A(\SUBBYTES[2].a/w2701 ), .B(\w1[2][30] ), .Z(
        n7665) );
  XOR \SUBBYTES[2].a/U4804  ( .A(\SUBBYTES[2].a/w2675 ), .B(
        \SUBBYTES[2].a/w2682 ), .Z(n7666) );
  XOR \SUBBYTES[2].a/U4803  ( .A(n7668), .B(n7667), .Z(n8286) );
  XOR \SUBBYTES[2].a/U4802  ( .A(\w1[2][25] ), .B(n7669), .Z(n7667) );
  XOR \SUBBYTES[2].a/U4801  ( .A(\SUBBYTES[2].a/w2700 ), .B(\w1[2][29] ), .Z(
        n7668) );
  XOR \SUBBYTES[2].a/U4800  ( .A(\SUBBYTES[2].a/w2676 ), .B(
        \SUBBYTES[2].a/w2683 ), .Z(n7669) );
  XOR \SUBBYTES[2].a/U4799  ( .A(n8288), .B(n8286), .Z(\SUBBYTES[2].a/w2706 )
         );
  XOR \SUBBYTES[2].a/U4798  ( .A(\w1[2][29] ), .B(n7670), .Z(n8289) );
  XOR \SUBBYTES[2].a/U4797  ( .A(\SUBBYTES[2].a/w2668 ), .B(
        \SUBBYTES[2].a/w2678 ), .Z(n7670) );
  XOR \SUBBYTES[2].a/U4796  ( .A(n7672), .B(n7671), .Z(\SUBBYTES[2].a/w2693 )
         );
  XOR \SUBBYTES[2].a/U4795  ( .A(n8289), .B(n7673), .Z(n7671) );
  XOR \SUBBYTES[2].a/U4794  ( .A(\w1[2][28] ), .B(\SUBBYTES[2].a/w2757 ), .Z(
        n7672) );
  XOR \SUBBYTES[2].a/U4793  ( .A(\SUBBYTES[2].a/w2670 ), .B(
        \SUBBYTES[2].a/w2675 ), .Z(n7673) );
  XOR \SUBBYTES[2].a/U4792  ( .A(n7675), .B(n7674), .Z(n8287) );
  XOR \SUBBYTES[2].a/U4791  ( .A(\SUBBYTES[2].a/w2703 ), .B(\w1[2][31] ), .Z(
        n7674) );
  XOR \SUBBYTES[2].a/U4790  ( .A(\SUBBYTES[2].a/w2678 ), .B(
        \SUBBYTES[2].a/w2685 ), .Z(n7675) );
  XOR \SUBBYTES[2].a/U4789  ( .A(n8286), .B(n8287), .Z(\SUBBYTES[2].a/w2705 )
         );
  XOR \SUBBYTES[2].a/U4788  ( .A(\w1[2][27] ), .B(n7676), .Z(n8290) );
  XOR \SUBBYTES[2].a/U4787  ( .A(\SUBBYTES[2].a/w2667 ), .B(
        \SUBBYTES[2].a/w2670 ), .Z(n7676) );
  XOR \SUBBYTES[2].a/U4786  ( .A(n7678), .B(n7677), .Z(\SUBBYTES[2].a/w2694 )
         );
  XOR \SUBBYTES[2].a/U4785  ( .A(n8290), .B(n7679), .Z(n7677) );
  XOR \SUBBYTES[2].a/U4784  ( .A(\w1[2][30] ), .B(\SUBBYTES[2].a/w2736 ), .Z(
        n7678) );
  XOR \SUBBYTES[2].a/U4783  ( .A(\SUBBYTES[2].a/w2675 ), .B(
        \SUBBYTES[2].a/w2676 ), .Z(n7679) );
  XOR \SUBBYTES[2].a/U4782  ( .A(n8288), .B(n8287), .Z(\SUBBYTES[2].a/w2714 )
         );
  XOR \SUBBYTES[2].a/U4781  ( .A(n7681), .B(n7680), .Z(\SUBBYTES[2].a/w2715 )
         );
  XOR \SUBBYTES[2].a/U4780  ( .A(\w1[2][31] ), .B(n8289), .Z(n7680) );
  XOR \SUBBYTES[2].a/U4779  ( .A(\SUBBYTES[2].a/w2667 ), .B(
        \SUBBYTES[2].a/w2676 ), .Z(n7681) );
  XOR \SUBBYTES[2].a/U4778  ( .A(n7683), .B(n7682), .Z(\SUBBYTES[2].a/w2691 )
         );
  XOR \SUBBYTES[2].a/U4777  ( .A(n7685), .B(n7684), .Z(n7682) );
  XOR \SUBBYTES[2].a/U4776  ( .A(\w1[2][31] ), .B(\SUBBYTES[2].a/w2775 ), .Z(
        n7683) );
  XOR \SUBBYTES[2].a/U4775  ( .A(\SUBBYTES[2].a/w2682 ), .B(
        \SUBBYTES[2].a/w2685 ), .Z(n7684) );
  XOR \SUBBYTES[2].a/U4774  ( .A(\SUBBYTES[2].a/w2668 ), .B(
        \SUBBYTES[2].a/w2670 ), .Z(n7685) );
  XOR \SUBBYTES[2].a/U4773  ( .A(n7687), .B(n7686), .Z(\SUBBYTES[2].a/w2692 )
         );
  XOR \SUBBYTES[2].a/U4772  ( .A(n8290), .B(n7688), .Z(n7686) );
  XOR \SUBBYTES[2].a/U4771  ( .A(\w1[2][29] ), .B(n8291), .Z(n7687) );
  XOR \SUBBYTES[2].a/U4770  ( .A(\SUBBYTES[2].a/w2682 ), .B(
        \SUBBYTES[2].a/w2683 ), .Z(n7688) );
  XOR \SUBBYTES[2].a/U4769  ( .A(n7690), .B(n7689), .Z(\SUBBYTES[2].a/w2708 )
         );
  XOR \SUBBYTES[2].a/U4768  ( .A(\w1[2][25] ), .B(n7691), .Z(n7689) );
  XOR \SUBBYTES[2].a/U4767  ( .A(\SUBBYTES[2].a/w2683 ), .B(
        \SUBBYTES[2].a/w2685 ), .Z(n7690) );
  XOR \SUBBYTES[2].a/U4766  ( .A(\SUBBYTES[2].a/w2667 ), .B(
        \SUBBYTES[2].a/w2668 ), .Z(n7691) );
  XOR \SUBBYTES[2].a/U4765  ( .A(\w1[2][33] ), .B(n7692), .Z(n8292) );
  XOR \SUBBYTES[2].a/U4764  ( .A(\w1[2][35] ), .B(\w1[2][34] ), .Z(n7692) );
  XOR \SUBBYTES[2].a/U4763  ( .A(\w1[2][38] ), .B(n8292), .Z(
        \SUBBYTES[2].a/w2550 ) );
  XOR \SUBBYTES[2].a/U4762  ( .A(\w1[2][32] ), .B(\SUBBYTES[2].a/w2550 ), .Z(
        \SUBBYTES[2].a/w2437 ) );
  XOR \SUBBYTES[2].a/U4761  ( .A(\w1[2][32] ), .B(n7693), .Z(
        \SUBBYTES[2].a/w2438 ) );
  XOR \SUBBYTES[2].a/U4760  ( .A(\w1[2][38] ), .B(\w1[2][37] ), .Z(n7693) );
  XOR \SUBBYTES[2].a/U4759  ( .A(\w1[2][37] ), .B(n8292), .Z(
        \SUBBYTES[2].a/w2568 ) );
  XOR \SUBBYTES[2].a/U4758  ( .A(n7695), .B(n7694), .Z(\SUBBYTES[2].a/w2561 )
         );
  XOR \SUBBYTES[2].a/U4757  ( .A(\w1[2][35] ), .B(\w1[2][33] ), .Z(n7694) );
  XOR \SUBBYTES[2].a/U4756  ( .A(\w1[2][39] ), .B(\w1[2][36] ), .Z(n7695) );
  XOR \SUBBYTES[2].a/U4755  ( .A(\w1[2][32] ), .B(\SUBBYTES[2].a/w2561 ), .Z(
        \SUBBYTES[2].a/w2440 ) );
  XOR \SUBBYTES[2].a/U4754  ( .A(n7697), .B(n7696), .Z(\SUBBYTES[2].a/w2548 )
         );
  XOR \SUBBYTES[2].a/U4753  ( .A(\SUBBYTES[2].a/w2509 ), .B(n984), .Z(n7696)
         );
  XOR \SUBBYTES[2].a/U4752  ( .A(\SUBBYTES[2].a/w2502 ), .B(
        \SUBBYTES[2].a/w2505 ), .Z(n7697) );
  XOR \SUBBYTES[2].a/U4751  ( .A(n7699), .B(n7698), .Z(\SUBBYTES[2].a/w2549 )
         );
  XOR \SUBBYTES[2].a/U4750  ( .A(\SUBBYTES[2].a/w2509 ), .B(n7135), .Z(n7698)
         );
  XOR \SUBBYTES[2].a/U4749  ( .A(\SUBBYTES[2].a/w2502 ), .B(n7134), .Z(n7699)
         );
  XOR \SUBBYTES[2].a/U4748  ( .A(\SUBBYTES[2].a/w2561 ), .B(n7700), .Z(
        \SUBBYTES[2].a/w2551 ) );
  XOR \SUBBYTES[2].a/U4747  ( .A(\w1[2][38] ), .B(\w1[2][37] ), .Z(n7700) );
  XOR \SUBBYTES[2].a/U4746  ( .A(n7702), .B(n7701), .Z(\SUBBYTES[2].a/w2552 )
         );
  XOR \SUBBYTES[2].a/U4745  ( .A(n7135), .B(n984), .Z(n7701) );
  XOR \SUBBYTES[2].a/U4744  ( .A(n7134), .B(\SUBBYTES[2].a/w2505 ), .Z(n7702)
         );
  XOR \SUBBYTES[2].a/U4743  ( .A(\w1[2][39] ), .B(\w1[2][34] ), .Z(n8298) );
  XOR \SUBBYTES[2].a/U4742  ( .A(n8298), .B(n7703), .Z(\SUBBYTES[2].a/w2553 )
         );
  XOR \SUBBYTES[2].a/U4741  ( .A(\w1[2][37] ), .B(\w1[2][36] ), .Z(n7703) );
  XOR \SUBBYTES[2].a/U4740  ( .A(\w1[2][39] ), .B(\SUBBYTES[2].a/w2438 ), .Z(
        \SUBBYTES[2].a/w2441 ) );
  XOR \SUBBYTES[2].a/U4739  ( .A(\w1[2][33] ), .B(\SUBBYTES[2].a/w2438 ), .Z(
        \SUBBYTES[2].a/w2442 ) );
  XOR \SUBBYTES[2].a/U4738  ( .A(\w1[2][36] ), .B(\SUBBYTES[2].a/w2438 ), .Z(
        \SUBBYTES[2].a/w2443 ) );
  XOR \SUBBYTES[2].a/U4737  ( .A(\SUBBYTES[2].a/w2442 ), .B(n8298), .Z(
        \SUBBYTES[2].a/w2444 ) );
  XOR \SUBBYTES[2].a/U4736  ( .A(n8298), .B(n7704), .Z(\SUBBYTES[2].a/w2529 )
         );
  XOR \SUBBYTES[2].a/U4735  ( .A(\w1[2][36] ), .B(\w1[2][33] ), .Z(n7704) );
  XOR \SUBBYTES[2].a/U4734  ( .A(n7706), .B(n7705), .Z(n8295) );
  XOR \SUBBYTES[2].a/U4733  ( .A(\w1[2][36] ), .B(n7707), .Z(n7705) );
  XOR \SUBBYTES[2].a/U4732  ( .A(\SUBBYTES[2].a/w2494 ), .B(\w1[2][38] ), .Z(
        n7706) );
  XOR \SUBBYTES[2].a/U4731  ( .A(\SUBBYTES[2].a/w2468 ), .B(
        \SUBBYTES[2].a/w2475 ), .Z(n7707) );
  XOR \SUBBYTES[2].a/U4730  ( .A(n7709), .B(n7708), .Z(n8293) );
  XOR \SUBBYTES[2].a/U4729  ( .A(\w1[2][33] ), .B(n7710), .Z(n7708) );
  XOR \SUBBYTES[2].a/U4728  ( .A(\SUBBYTES[2].a/w2493 ), .B(\w1[2][37] ), .Z(
        n7709) );
  XOR \SUBBYTES[2].a/U4727  ( .A(\SUBBYTES[2].a/w2469 ), .B(
        \SUBBYTES[2].a/w2476 ), .Z(n7710) );
  XOR \SUBBYTES[2].a/U4726  ( .A(n8295), .B(n8293), .Z(\SUBBYTES[2].a/w2499 )
         );
  XOR \SUBBYTES[2].a/U4725  ( .A(\w1[2][37] ), .B(n7711), .Z(n8296) );
  XOR \SUBBYTES[2].a/U4724  ( .A(\SUBBYTES[2].a/w2461 ), .B(
        \SUBBYTES[2].a/w2471 ), .Z(n7711) );
  XOR \SUBBYTES[2].a/U4723  ( .A(n7713), .B(n7712), .Z(\SUBBYTES[2].a/w2486 )
         );
  XOR \SUBBYTES[2].a/U4722  ( .A(n8296), .B(n7714), .Z(n7712) );
  XOR \SUBBYTES[2].a/U4721  ( .A(\w1[2][36] ), .B(\SUBBYTES[2].a/w2550 ), .Z(
        n7713) );
  XOR \SUBBYTES[2].a/U4720  ( .A(\SUBBYTES[2].a/w2463 ), .B(
        \SUBBYTES[2].a/w2468 ), .Z(n7714) );
  XOR \SUBBYTES[2].a/U4719  ( .A(n7716), .B(n7715), .Z(n8294) );
  XOR \SUBBYTES[2].a/U4718  ( .A(\SUBBYTES[2].a/w2496 ), .B(\w1[2][39] ), .Z(
        n7715) );
  XOR \SUBBYTES[2].a/U4717  ( .A(\SUBBYTES[2].a/w2471 ), .B(
        \SUBBYTES[2].a/w2478 ), .Z(n7716) );
  XOR \SUBBYTES[2].a/U4716  ( .A(n8293), .B(n8294), .Z(\SUBBYTES[2].a/w2498 )
         );
  XOR \SUBBYTES[2].a/U4715  ( .A(\w1[2][35] ), .B(n7717), .Z(n8297) );
  XOR \SUBBYTES[2].a/U4714  ( .A(\SUBBYTES[2].a/w2460 ), .B(
        \SUBBYTES[2].a/w2463 ), .Z(n7717) );
  XOR \SUBBYTES[2].a/U4713  ( .A(n7719), .B(n7718), .Z(\SUBBYTES[2].a/w2487 )
         );
  XOR \SUBBYTES[2].a/U4712  ( .A(n8297), .B(n7720), .Z(n7718) );
  XOR \SUBBYTES[2].a/U4711  ( .A(\w1[2][38] ), .B(\SUBBYTES[2].a/w2529 ), .Z(
        n7719) );
  XOR \SUBBYTES[2].a/U4710  ( .A(\SUBBYTES[2].a/w2468 ), .B(
        \SUBBYTES[2].a/w2469 ), .Z(n7720) );
  XOR \SUBBYTES[2].a/U4709  ( .A(n8295), .B(n8294), .Z(\SUBBYTES[2].a/w2507 )
         );
  XOR \SUBBYTES[2].a/U4708  ( .A(n7722), .B(n7721), .Z(\SUBBYTES[2].a/w2508 )
         );
  XOR \SUBBYTES[2].a/U4707  ( .A(\w1[2][39] ), .B(n8296), .Z(n7721) );
  XOR \SUBBYTES[2].a/U4706  ( .A(\SUBBYTES[2].a/w2460 ), .B(
        \SUBBYTES[2].a/w2469 ), .Z(n7722) );
  XOR \SUBBYTES[2].a/U4705  ( .A(n7724), .B(n7723), .Z(\SUBBYTES[2].a/w2484 )
         );
  XOR \SUBBYTES[2].a/U4704  ( .A(n7726), .B(n7725), .Z(n7723) );
  XOR \SUBBYTES[2].a/U4703  ( .A(\w1[2][39] ), .B(\SUBBYTES[2].a/w2568 ), .Z(
        n7724) );
  XOR \SUBBYTES[2].a/U4702  ( .A(\SUBBYTES[2].a/w2475 ), .B(
        \SUBBYTES[2].a/w2478 ), .Z(n7725) );
  XOR \SUBBYTES[2].a/U4701  ( .A(\SUBBYTES[2].a/w2461 ), .B(
        \SUBBYTES[2].a/w2463 ), .Z(n7726) );
  XOR \SUBBYTES[2].a/U4700  ( .A(n7728), .B(n7727), .Z(\SUBBYTES[2].a/w2485 )
         );
  XOR \SUBBYTES[2].a/U4699  ( .A(n8297), .B(n7729), .Z(n7727) );
  XOR \SUBBYTES[2].a/U4698  ( .A(\w1[2][37] ), .B(n8298), .Z(n7728) );
  XOR \SUBBYTES[2].a/U4697  ( .A(\SUBBYTES[2].a/w2475 ), .B(
        \SUBBYTES[2].a/w2476 ), .Z(n7729) );
  XOR \SUBBYTES[2].a/U4696  ( .A(n7731), .B(n7730), .Z(\SUBBYTES[2].a/w2501 )
         );
  XOR \SUBBYTES[2].a/U4695  ( .A(\w1[2][33] ), .B(n7732), .Z(n7730) );
  XOR \SUBBYTES[2].a/U4694  ( .A(\SUBBYTES[2].a/w2476 ), .B(
        \SUBBYTES[2].a/w2478 ), .Z(n7731) );
  XOR \SUBBYTES[2].a/U4693  ( .A(\SUBBYTES[2].a/w2460 ), .B(
        \SUBBYTES[2].a/w2461 ), .Z(n7732) );
  XOR \SUBBYTES[2].a/U4692  ( .A(\w1[2][41] ), .B(n7733), .Z(n8299) );
  XOR \SUBBYTES[2].a/U4691  ( .A(\w1[2][43] ), .B(\w1[2][42] ), .Z(n7733) );
  XOR \SUBBYTES[2].a/U4690  ( .A(\w1[2][46] ), .B(n8299), .Z(
        \SUBBYTES[2].a/w2343 ) );
  XOR \SUBBYTES[2].a/U4689  ( .A(\w1[2][40] ), .B(\SUBBYTES[2].a/w2343 ), .Z(
        \SUBBYTES[2].a/w2230 ) );
  XOR \SUBBYTES[2].a/U4688  ( .A(\w1[2][40] ), .B(n7734), .Z(
        \SUBBYTES[2].a/w2231 ) );
  XOR \SUBBYTES[2].a/U4687  ( .A(\w1[2][46] ), .B(\w1[2][45] ), .Z(n7734) );
  XOR \SUBBYTES[2].a/U4686  ( .A(\w1[2][45] ), .B(n8299), .Z(
        \SUBBYTES[2].a/w2361 ) );
  XOR \SUBBYTES[2].a/U4685  ( .A(n7736), .B(n7735), .Z(\SUBBYTES[2].a/w2354 )
         );
  XOR \SUBBYTES[2].a/U4684  ( .A(\w1[2][43] ), .B(\w1[2][41] ), .Z(n7735) );
  XOR \SUBBYTES[2].a/U4683  ( .A(\w1[2][47] ), .B(\w1[2][44] ), .Z(n7736) );
  XOR \SUBBYTES[2].a/U4682  ( .A(\w1[2][40] ), .B(\SUBBYTES[2].a/w2354 ), .Z(
        \SUBBYTES[2].a/w2233 ) );
  XOR \SUBBYTES[2].a/U4681  ( .A(n7738), .B(n7737), .Z(\SUBBYTES[2].a/w2341 )
         );
  XOR \SUBBYTES[2].a/U4680  ( .A(\SUBBYTES[2].a/w2302 ), .B(n983), .Z(n7737)
         );
  XOR \SUBBYTES[2].a/U4679  ( .A(\SUBBYTES[2].a/w2295 ), .B(
        \SUBBYTES[2].a/w2298 ), .Z(n7738) );
  XOR \SUBBYTES[2].a/U4678  ( .A(n7740), .B(n7739), .Z(\SUBBYTES[2].a/w2342 )
         );
  XOR \SUBBYTES[2].a/U4677  ( .A(\SUBBYTES[2].a/w2302 ), .B(n7133), .Z(n7739)
         );
  XOR \SUBBYTES[2].a/U4676  ( .A(\SUBBYTES[2].a/w2295 ), .B(n7132), .Z(n7740)
         );
  XOR \SUBBYTES[2].a/U4675  ( .A(\SUBBYTES[2].a/w2354 ), .B(n7741), .Z(
        \SUBBYTES[2].a/w2344 ) );
  XOR \SUBBYTES[2].a/U4674  ( .A(\w1[2][46] ), .B(\w1[2][45] ), .Z(n7741) );
  XOR \SUBBYTES[2].a/U4673  ( .A(n7743), .B(n7742), .Z(\SUBBYTES[2].a/w2345 )
         );
  XOR \SUBBYTES[2].a/U4672  ( .A(n7133), .B(n983), .Z(n7742) );
  XOR \SUBBYTES[2].a/U4671  ( .A(n7132), .B(\SUBBYTES[2].a/w2298 ), .Z(n7743)
         );
  XOR \SUBBYTES[2].a/U4670  ( .A(\w1[2][47] ), .B(\w1[2][42] ), .Z(n8305) );
  XOR \SUBBYTES[2].a/U4669  ( .A(n8305), .B(n7744), .Z(\SUBBYTES[2].a/w2346 )
         );
  XOR \SUBBYTES[2].a/U4668  ( .A(\w1[2][45] ), .B(\w1[2][44] ), .Z(n7744) );
  XOR \SUBBYTES[2].a/U4667  ( .A(\w1[2][47] ), .B(\SUBBYTES[2].a/w2231 ), .Z(
        \SUBBYTES[2].a/w2234 ) );
  XOR \SUBBYTES[2].a/U4666  ( .A(\w1[2][41] ), .B(\SUBBYTES[2].a/w2231 ), .Z(
        \SUBBYTES[2].a/w2235 ) );
  XOR \SUBBYTES[2].a/U4665  ( .A(\w1[2][44] ), .B(\SUBBYTES[2].a/w2231 ), .Z(
        \SUBBYTES[2].a/w2236 ) );
  XOR \SUBBYTES[2].a/U4664  ( .A(\SUBBYTES[2].a/w2235 ), .B(n8305), .Z(
        \SUBBYTES[2].a/w2237 ) );
  XOR \SUBBYTES[2].a/U4663  ( .A(n8305), .B(n7745), .Z(\SUBBYTES[2].a/w2322 )
         );
  XOR \SUBBYTES[2].a/U4662  ( .A(\w1[2][44] ), .B(\w1[2][41] ), .Z(n7745) );
  XOR \SUBBYTES[2].a/U4661  ( .A(n7747), .B(n7746), .Z(n8302) );
  XOR \SUBBYTES[2].a/U4660  ( .A(\w1[2][44] ), .B(n7748), .Z(n7746) );
  XOR \SUBBYTES[2].a/U4659  ( .A(\SUBBYTES[2].a/w2287 ), .B(\w1[2][46] ), .Z(
        n7747) );
  XOR \SUBBYTES[2].a/U4658  ( .A(\SUBBYTES[2].a/w2261 ), .B(
        \SUBBYTES[2].a/w2268 ), .Z(n7748) );
  XOR \SUBBYTES[2].a/U4657  ( .A(n7750), .B(n7749), .Z(n8300) );
  XOR \SUBBYTES[2].a/U4656  ( .A(\w1[2][41] ), .B(n7751), .Z(n7749) );
  XOR \SUBBYTES[2].a/U4655  ( .A(\SUBBYTES[2].a/w2286 ), .B(\w1[2][45] ), .Z(
        n7750) );
  XOR \SUBBYTES[2].a/U4654  ( .A(\SUBBYTES[2].a/w2262 ), .B(
        \SUBBYTES[2].a/w2269 ), .Z(n7751) );
  XOR \SUBBYTES[2].a/U4653  ( .A(n8302), .B(n8300), .Z(\SUBBYTES[2].a/w2292 )
         );
  XOR \SUBBYTES[2].a/U4652  ( .A(\w1[2][45] ), .B(n7752), .Z(n8303) );
  XOR \SUBBYTES[2].a/U4651  ( .A(\SUBBYTES[2].a/w2254 ), .B(
        \SUBBYTES[2].a/w2264 ), .Z(n7752) );
  XOR \SUBBYTES[2].a/U4650  ( .A(n7754), .B(n7753), .Z(\SUBBYTES[2].a/w2279 )
         );
  XOR \SUBBYTES[2].a/U4649  ( .A(n8303), .B(n7755), .Z(n7753) );
  XOR \SUBBYTES[2].a/U4648  ( .A(\w1[2][44] ), .B(\SUBBYTES[2].a/w2343 ), .Z(
        n7754) );
  XOR \SUBBYTES[2].a/U4647  ( .A(\SUBBYTES[2].a/w2256 ), .B(
        \SUBBYTES[2].a/w2261 ), .Z(n7755) );
  XOR \SUBBYTES[2].a/U4646  ( .A(n7757), .B(n7756), .Z(n8301) );
  XOR \SUBBYTES[2].a/U4645  ( .A(\SUBBYTES[2].a/w2289 ), .B(\w1[2][47] ), .Z(
        n7756) );
  XOR \SUBBYTES[2].a/U4644  ( .A(\SUBBYTES[2].a/w2264 ), .B(
        \SUBBYTES[2].a/w2271 ), .Z(n7757) );
  XOR \SUBBYTES[2].a/U4643  ( .A(n8300), .B(n8301), .Z(\SUBBYTES[2].a/w2291 )
         );
  XOR \SUBBYTES[2].a/U4642  ( .A(\w1[2][43] ), .B(n7758), .Z(n8304) );
  XOR \SUBBYTES[2].a/U4641  ( .A(\SUBBYTES[2].a/w2253 ), .B(
        \SUBBYTES[2].a/w2256 ), .Z(n7758) );
  XOR \SUBBYTES[2].a/U4640  ( .A(n7760), .B(n7759), .Z(\SUBBYTES[2].a/w2280 )
         );
  XOR \SUBBYTES[2].a/U4639  ( .A(n8304), .B(n7761), .Z(n7759) );
  XOR \SUBBYTES[2].a/U4638  ( .A(\w1[2][46] ), .B(\SUBBYTES[2].a/w2322 ), .Z(
        n7760) );
  XOR \SUBBYTES[2].a/U4637  ( .A(\SUBBYTES[2].a/w2261 ), .B(
        \SUBBYTES[2].a/w2262 ), .Z(n7761) );
  XOR \SUBBYTES[2].a/U4636  ( .A(n8302), .B(n8301), .Z(\SUBBYTES[2].a/w2300 )
         );
  XOR \SUBBYTES[2].a/U4635  ( .A(n7763), .B(n7762), .Z(\SUBBYTES[2].a/w2301 )
         );
  XOR \SUBBYTES[2].a/U4634  ( .A(\w1[2][47] ), .B(n8303), .Z(n7762) );
  XOR \SUBBYTES[2].a/U4633  ( .A(\SUBBYTES[2].a/w2253 ), .B(
        \SUBBYTES[2].a/w2262 ), .Z(n7763) );
  XOR \SUBBYTES[2].a/U4632  ( .A(n7765), .B(n7764), .Z(\SUBBYTES[2].a/w2277 )
         );
  XOR \SUBBYTES[2].a/U4631  ( .A(n7767), .B(n7766), .Z(n7764) );
  XOR \SUBBYTES[2].a/U4630  ( .A(\w1[2][47] ), .B(\SUBBYTES[2].a/w2361 ), .Z(
        n7765) );
  XOR \SUBBYTES[2].a/U4629  ( .A(\SUBBYTES[2].a/w2268 ), .B(
        \SUBBYTES[2].a/w2271 ), .Z(n7766) );
  XOR \SUBBYTES[2].a/U4628  ( .A(\SUBBYTES[2].a/w2254 ), .B(
        \SUBBYTES[2].a/w2256 ), .Z(n7767) );
  XOR \SUBBYTES[2].a/U4627  ( .A(n7769), .B(n7768), .Z(\SUBBYTES[2].a/w2278 )
         );
  XOR \SUBBYTES[2].a/U4626  ( .A(n8304), .B(n7770), .Z(n7768) );
  XOR \SUBBYTES[2].a/U4625  ( .A(\w1[2][45] ), .B(n8305), .Z(n7769) );
  XOR \SUBBYTES[2].a/U4624  ( .A(\SUBBYTES[2].a/w2268 ), .B(
        \SUBBYTES[2].a/w2269 ), .Z(n7770) );
  XOR \SUBBYTES[2].a/U4623  ( .A(n7772), .B(n7771), .Z(\SUBBYTES[2].a/w2294 )
         );
  XOR \SUBBYTES[2].a/U4622  ( .A(\w1[2][41] ), .B(n7773), .Z(n7771) );
  XOR \SUBBYTES[2].a/U4621  ( .A(\SUBBYTES[2].a/w2269 ), .B(
        \SUBBYTES[2].a/w2271 ), .Z(n7772) );
  XOR \SUBBYTES[2].a/U4620  ( .A(\SUBBYTES[2].a/w2253 ), .B(
        \SUBBYTES[2].a/w2254 ), .Z(n7773) );
  XOR \SUBBYTES[2].a/U4619  ( .A(\w1[2][49] ), .B(n7774), .Z(n8306) );
  XOR \SUBBYTES[2].a/U4618  ( .A(\w1[2][51] ), .B(\w1[2][50] ), .Z(n7774) );
  XOR \SUBBYTES[2].a/U4617  ( .A(\w1[2][54] ), .B(n8306), .Z(
        \SUBBYTES[2].a/w2136 ) );
  XOR \SUBBYTES[2].a/U4616  ( .A(\w1[2][48] ), .B(\SUBBYTES[2].a/w2136 ), .Z(
        \SUBBYTES[2].a/w2023 ) );
  XOR \SUBBYTES[2].a/U4615  ( .A(\w1[2][48] ), .B(n7775), .Z(
        \SUBBYTES[2].a/w2024 ) );
  XOR \SUBBYTES[2].a/U4614  ( .A(\w1[2][54] ), .B(\w1[2][53] ), .Z(n7775) );
  XOR \SUBBYTES[2].a/U4613  ( .A(\w1[2][53] ), .B(n8306), .Z(
        \SUBBYTES[2].a/w2154 ) );
  XOR \SUBBYTES[2].a/U4612  ( .A(n7777), .B(n7776), .Z(\SUBBYTES[2].a/w2147 )
         );
  XOR \SUBBYTES[2].a/U4611  ( .A(\w1[2][51] ), .B(\w1[2][49] ), .Z(n7776) );
  XOR \SUBBYTES[2].a/U4610  ( .A(\w1[2][55] ), .B(\w1[2][52] ), .Z(n7777) );
  XOR \SUBBYTES[2].a/U4609  ( .A(\w1[2][48] ), .B(\SUBBYTES[2].a/w2147 ), .Z(
        \SUBBYTES[2].a/w2026 ) );
  XOR \SUBBYTES[2].a/U4608  ( .A(n7779), .B(n7778), .Z(\SUBBYTES[2].a/w2134 )
         );
  XOR \SUBBYTES[2].a/U4607  ( .A(\SUBBYTES[2].a/w2095 ), .B(n982), .Z(n7778)
         );
  XOR \SUBBYTES[2].a/U4606  ( .A(\SUBBYTES[2].a/w2088 ), .B(
        \SUBBYTES[2].a/w2091 ), .Z(n7779) );
  XOR \SUBBYTES[2].a/U4605  ( .A(n7781), .B(n7780), .Z(\SUBBYTES[2].a/w2135 )
         );
  XOR \SUBBYTES[2].a/U4604  ( .A(\SUBBYTES[2].a/w2095 ), .B(n7131), .Z(n7780)
         );
  XOR \SUBBYTES[2].a/U4603  ( .A(\SUBBYTES[2].a/w2088 ), .B(n7130), .Z(n7781)
         );
  XOR \SUBBYTES[2].a/U4602  ( .A(\SUBBYTES[2].a/w2147 ), .B(n7782), .Z(
        \SUBBYTES[2].a/w2137 ) );
  XOR \SUBBYTES[2].a/U4601  ( .A(\w1[2][54] ), .B(\w1[2][53] ), .Z(n7782) );
  XOR \SUBBYTES[2].a/U4600  ( .A(n7784), .B(n7783), .Z(\SUBBYTES[2].a/w2138 )
         );
  XOR \SUBBYTES[2].a/U4599  ( .A(n7131), .B(n982), .Z(n7783) );
  XOR \SUBBYTES[2].a/U4598  ( .A(n7130), .B(\SUBBYTES[2].a/w2091 ), .Z(n7784)
         );
  XOR \SUBBYTES[2].a/U4597  ( .A(\w1[2][55] ), .B(\w1[2][50] ), .Z(n8312) );
  XOR \SUBBYTES[2].a/U4596  ( .A(n8312), .B(n7785), .Z(\SUBBYTES[2].a/w2139 )
         );
  XOR \SUBBYTES[2].a/U4595  ( .A(\w1[2][53] ), .B(\w1[2][52] ), .Z(n7785) );
  XOR \SUBBYTES[2].a/U4594  ( .A(\w1[2][55] ), .B(\SUBBYTES[2].a/w2024 ), .Z(
        \SUBBYTES[2].a/w2027 ) );
  XOR \SUBBYTES[2].a/U4593  ( .A(\w1[2][49] ), .B(\SUBBYTES[2].a/w2024 ), .Z(
        \SUBBYTES[2].a/w2028 ) );
  XOR \SUBBYTES[2].a/U4592  ( .A(\w1[2][52] ), .B(\SUBBYTES[2].a/w2024 ), .Z(
        \SUBBYTES[2].a/w2029 ) );
  XOR \SUBBYTES[2].a/U4591  ( .A(\SUBBYTES[2].a/w2028 ), .B(n8312), .Z(
        \SUBBYTES[2].a/w2030 ) );
  XOR \SUBBYTES[2].a/U4590  ( .A(n8312), .B(n7786), .Z(\SUBBYTES[2].a/w2115 )
         );
  XOR \SUBBYTES[2].a/U4589  ( .A(\w1[2][52] ), .B(\w1[2][49] ), .Z(n7786) );
  XOR \SUBBYTES[2].a/U4588  ( .A(n7788), .B(n7787), .Z(n8309) );
  XOR \SUBBYTES[2].a/U4587  ( .A(\w1[2][52] ), .B(n7789), .Z(n7787) );
  XOR \SUBBYTES[2].a/U4586  ( .A(\SUBBYTES[2].a/w2080 ), .B(\w1[2][54] ), .Z(
        n7788) );
  XOR \SUBBYTES[2].a/U4585  ( .A(\SUBBYTES[2].a/w2054 ), .B(
        \SUBBYTES[2].a/w2061 ), .Z(n7789) );
  XOR \SUBBYTES[2].a/U4584  ( .A(n7791), .B(n7790), .Z(n8307) );
  XOR \SUBBYTES[2].a/U4583  ( .A(\w1[2][49] ), .B(n7792), .Z(n7790) );
  XOR \SUBBYTES[2].a/U4582  ( .A(\SUBBYTES[2].a/w2079 ), .B(\w1[2][53] ), .Z(
        n7791) );
  XOR \SUBBYTES[2].a/U4581  ( .A(\SUBBYTES[2].a/w2055 ), .B(
        \SUBBYTES[2].a/w2062 ), .Z(n7792) );
  XOR \SUBBYTES[2].a/U4580  ( .A(n8309), .B(n8307), .Z(\SUBBYTES[2].a/w2085 )
         );
  XOR \SUBBYTES[2].a/U4579  ( .A(\w1[2][53] ), .B(n7793), .Z(n8310) );
  XOR \SUBBYTES[2].a/U4578  ( .A(\SUBBYTES[2].a/w2047 ), .B(
        \SUBBYTES[2].a/w2057 ), .Z(n7793) );
  XOR \SUBBYTES[2].a/U4577  ( .A(n7795), .B(n7794), .Z(\SUBBYTES[2].a/w2072 )
         );
  XOR \SUBBYTES[2].a/U4576  ( .A(n8310), .B(n7796), .Z(n7794) );
  XOR \SUBBYTES[2].a/U4575  ( .A(\w1[2][52] ), .B(\SUBBYTES[2].a/w2136 ), .Z(
        n7795) );
  XOR \SUBBYTES[2].a/U4574  ( .A(\SUBBYTES[2].a/w2049 ), .B(
        \SUBBYTES[2].a/w2054 ), .Z(n7796) );
  XOR \SUBBYTES[2].a/U4573  ( .A(n7798), .B(n7797), .Z(n8308) );
  XOR \SUBBYTES[2].a/U4572  ( .A(\SUBBYTES[2].a/w2082 ), .B(\w1[2][55] ), .Z(
        n7797) );
  XOR \SUBBYTES[2].a/U4571  ( .A(\SUBBYTES[2].a/w2057 ), .B(
        \SUBBYTES[2].a/w2064 ), .Z(n7798) );
  XOR \SUBBYTES[2].a/U4570  ( .A(n8307), .B(n8308), .Z(\SUBBYTES[2].a/w2084 )
         );
  XOR \SUBBYTES[2].a/U4569  ( .A(\w1[2][51] ), .B(n7799), .Z(n8311) );
  XOR \SUBBYTES[2].a/U4568  ( .A(\SUBBYTES[2].a/w2046 ), .B(
        \SUBBYTES[2].a/w2049 ), .Z(n7799) );
  XOR \SUBBYTES[2].a/U4567  ( .A(n7801), .B(n7800), .Z(\SUBBYTES[2].a/w2073 )
         );
  XOR \SUBBYTES[2].a/U4566  ( .A(n8311), .B(n7802), .Z(n7800) );
  XOR \SUBBYTES[2].a/U4565  ( .A(\w1[2][54] ), .B(\SUBBYTES[2].a/w2115 ), .Z(
        n7801) );
  XOR \SUBBYTES[2].a/U4564  ( .A(\SUBBYTES[2].a/w2054 ), .B(
        \SUBBYTES[2].a/w2055 ), .Z(n7802) );
  XOR \SUBBYTES[2].a/U4563  ( .A(n8309), .B(n8308), .Z(\SUBBYTES[2].a/w2093 )
         );
  XOR \SUBBYTES[2].a/U4562  ( .A(n7804), .B(n7803), .Z(\SUBBYTES[2].a/w2094 )
         );
  XOR \SUBBYTES[2].a/U4561  ( .A(\w1[2][55] ), .B(n8310), .Z(n7803) );
  XOR \SUBBYTES[2].a/U4560  ( .A(\SUBBYTES[2].a/w2046 ), .B(
        \SUBBYTES[2].a/w2055 ), .Z(n7804) );
  XOR \SUBBYTES[2].a/U4559  ( .A(n7806), .B(n7805), .Z(\SUBBYTES[2].a/w2070 )
         );
  XOR \SUBBYTES[2].a/U4558  ( .A(n7808), .B(n7807), .Z(n7805) );
  XOR \SUBBYTES[2].a/U4557  ( .A(\w1[2][55] ), .B(\SUBBYTES[2].a/w2154 ), .Z(
        n7806) );
  XOR \SUBBYTES[2].a/U4556  ( .A(\SUBBYTES[2].a/w2061 ), .B(
        \SUBBYTES[2].a/w2064 ), .Z(n7807) );
  XOR \SUBBYTES[2].a/U4555  ( .A(\SUBBYTES[2].a/w2047 ), .B(
        \SUBBYTES[2].a/w2049 ), .Z(n7808) );
  XOR \SUBBYTES[2].a/U4554  ( .A(n7810), .B(n7809), .Z(\SUBBYTES[2].a/w2071 )
         );
  XOR \SUBBYTES[2].a/U4553  ( .A(n8311), .B(n7811), .Z(n7809) );
  XOR \SUBBYTES[2].a/U4552  ( .A(\w1[2][53] ), .B(n8312), .Z(n7810) );
  XOR \SUBBYTES[2].a/U4551  ( .A(\SUBBYTES[2].a/w2061 ), .B(
        \SUBBYTES[2].a/w2062 ), .Z(n7811) );
  XOR \SUBBYTES[2].a/U4550  ( .A(n7813), .B(n7812), .Z(\SUBBYTES[2].a/w2087 )
         );
  XOR \SUBBYTES[2].a/U4549  ( .A(\w1[2][49] ), .B(n7814), .Z(n7812) );
  XOR \SUBBYTES[2].a/U4548  ( .A(\SUBBYTES[2].a/w2062 ), .B(
        \SUBBYTES[2].a/w2064 ), .Z(n7813) );
  XOR \SUBBYTES[2].a/U4547  ( .A(\SUBBYTES[2].a/w2046 ), .B(
        \SUBBYTES[2].a/w2047 ), .Z(n7814) );
  XOR \SUBBYTES[2].a/U4546  ( .A(\w1[2][57] ), .B(n7815), .Z(n8313) );
  XOR \SUBBYTES[2].a/U4545  ( .A(\w1[2][59] ), .B(\w1[2][58] ), .Z(n7815) );
  XOR \SUBBYTES[2].a/U4544  ( .A(\w1[2][62] ), .B(n8313), .Z(
        \SUBBYTES[2].a/w1929 ) );
  XOR \SUBBYTES[2].a/U4543  ( .A(\w1[2][56] ), .B(\SUBBYTES[2].a/w1929 ), .Z(
        \SUBBYTES[2].a/w1816 ) );
  XOR \SUBBYTES[2].a/U4542  ( .A(\w1[2][56] ), .B(n7816), .Z(
        \SUBBYTES[2].a/w1817 ) );
  XOR \SUBBYTES[2].a/U4541  ( .A(\w1[2][62] ), .B(\w1[2][61] ), .Z(n7816) );
  XOR \SUBBYTES[2].a/U4540  ( .A(\w1[2][61] ), .B(n8313), .Z(
        \SUBBYTES[2].a/w1947 ) );
  XOR \SUBBYTES[2].a/U4539  ( .A(n7818), .B(n7817), .Z(\SUBBYTES[2].a/w1940 )
         );
  XOR \SUBBYTES[2].a/U4538  ( .A(\w1[2][59] ), .B(\w1[2][57] ), .Z(n7817) );
  XOR \SUBBYTES[2].a/U4537  ( .A(\w1[2][63] ), .B(\w1[2][60] ), .Z(n7818) );
  XOR \SUBBYTES[2].a/U4536  ( .A(\w1[2][56] ), .B(\SUBBYTES[2].a/w1940 ), .Z(
        \SUBBYTES[2].a/w1819 ) );
  XOR \SUBBYTES[2].a/U4535  ( .A(n7820), .B(n7819), .Z(\SUBBYTES[2].a/w1927 )
         );
  XOR \SUBBYTES[2].a/U4534  ( .A(\SUBBYTES[2].a/w1888 ), .B(n981), .Z(n7819)
         );
  XOR \SUBBYTES[2].a/U4533  ( .A(\SUBBYTES[2].a/w1881 ), .B(
        \SUBBYTES[2].a/w1884 ), .Z(n7820) );
  XOR \SUBBYTES[2].a/U4532  ( .A(n7822), .B(n7821), .Z(\SUBBYTES[2].a/w1928 )
         );
  XOR \SUBBYTES[2].a/U4531  ( .A(\SUBBYTES[2].a/w1888 ), .B(n7129), .Z(n7821)
         );
  XOR \SUBBYTES[2].a/U4530  ( .A(\SUBBYTES[2].a/w1881 ), .B(n7128), .Z(n7822)
         );
  XOR \SUBBYTES[2].a/U4529  ( .A(\SUBBYTES[2].a/w1940 ), .B(n7823), .Z(
        \SUBBYTES[2].a/w1930 ) );
  XOR \SUBBYTES[2].a/U4528  ( .A(\w1[2][62] ), .B(\w1[2][61] ), .Z(n7823) );
  XOR \SUBBYTES[2].a/U4527  ( .A(n7825), .B(n7824), .Z(\SUBBYTES[2].a/w1931 )
         );
  XOR \SUBBYTES[2].a/U4526  ( .A(n7129), .B(n981), .Z(n7824) );
  XOR \SUBBYTES[2].a/U4525  ( .A(n7128), .B(\SUBBYTES[2].a/w1884 ), .Z(n7825)
         );
  XOR \SUBBYTES[2].a/U4524  ( .A(\w1[2][63] ), .B(\w1[2][58] ), .Z(n8319) );
  XOR \SUBBYTES[2].a/U4523  ( .A(n8319), .B(n7826), .Z(\SUBBYTES[2].a/w1932 )
         );
  XOR \SUBBYTES[2].a/U4522  ( .A(\w1[2][61] ), .B(\w1[2][60] ), .Z(n7826) );
  XOR \SUBBYTES[2].a/U4521  ( .A(\w1[2][63] ), .B(\SUBBYTES[2].a/w1817 ), .Z(
        \SUBBYTES[2].a/w1820 ) );
  XOR \SUBBYTES[2].a/U4520  ( .A(\w1[2][57] ), .B(\SUBBYTES[2].a/w1817 ), .Z(
        \SUBBYTES[2].a/w1821 ) );
  XOR \SUBBYTES[2].a/U4519  ( .A(\w1[2][60] ), .B(\SUBBYTES[2].a/w1817 ), .Z(
        \SUBBYTES[2].a/w1822 ) );
  XOR \SUBBYTES[2].a/U4518  ( .A(\SUBBYTES[2].a/w1821 ), .B(n8319), .Z(
        \SUBBYTES[2].a/w1823 ) );
  XOR \SUBBYTES[2].a/U4517  ( .A(n8319), .B(n7827), .Z(\SUBBYTES[2].a/w1908 )
         );
  XOR \SUBBYTES[2].a/U4516  ( .A(\w1[2][60] ), .B(\w1[2][57] ), .Z(n7827) );
  XOR \SUBBYTES[2].a/U4515  ( .A(n7829), .B(n7828), .Z(n8316) );
  XOR \SUBBYTES[2].a/U4514  ( .A(\w1[2][60] ), .B(n7830), .Z(n7828) );
  XOR \SUBBYTES[2].a/U4513  ( .A(\SUBBYTES[2].a/w1873 ), .B(\w1[2][62] ), .Z(
        n7829) );
  XOR \SUBBYTES[2].a/U4512  ( .A(\SUBBYTES[2].a/w1847 ), .B(
        \SUBBYTES[2].a/w1854 ), .Z(n7830) );
  XOR \SUBBYTES[2].a/U4511  ( .A(n7832), .B(n7831), .Z(n8314) );
  XOR \SUBBYTES[2].a/U4510  ( .A(\w1[2][57] ), .B(n7833), .Z(n7831) );
  XOR \SUBBYTES[2].a/U4509  ( .A(\SUBBYTES[2].a/w1872 ), .B(\w1[2][61] ), .Z(
        n7832) );
  XOR \SUBBYTES[2].a/U4508  ( .A(\SUBBYTES[2].a/w1848 ), .B(
        \SUBBYTES[2].a/w1855 ), .Z(n7833) );
  XOR \SUBBYTES[2].a/U4507  ( .A(n8316), .B(n8314), .Z(\SUBBYTES[2].a/w1878 )
         );
  XOR \SUBBYTES[2].a/U4506  ( .A(\w1[2][61] ), .B(n7834), .Z(n8317) );
  XOR \SUBBYTES[2].a/U4505  ( .A(\SUBBYTES[2].a/w1840 ), .B(
        \SUBBYTES[2].a/w1850 ), .Z(n7834) );
  XOR \SUBBYTES[2].a/U4504  ( .A(n7836), .B(n7835), .Z(\SUBBYTES[2].a/w1865 )
         );
  XOR \SUBBYTES[2].a/U4503  ( .A(n8317), .B(n7837), .Z(n7835) );
  XOR \SUBBYTES[2].a/U4502  ( .A(\w1[2][60] ), .B(\SUBBYTES[2].a/w1929 ), .Z(
        n7836) );
  XOR \SUBBYTES[2].a/U4501  ( .A(\SUBBYTES[2].a/w1842 ), .B(
        \SUBBYTES[2].a/w1847 ), .Z(n7837) );
  XOR \SUBBYTES[2].a/U4500  ( .A(n7839), .B(n7838), .Z(n8315) );
  XOR \SUBBYTES[2].a/U4499  ( .A(\SUBBYTES[2].a/w1875 ), .B(\w1[2][63] ), .Z(
        n7838) );
  XOR \SUBBYTES[2].a/U4498  ( .A(\SUBBYTES[2].a/w1850 ), .B(
        \SUBBYTES[2].a/w1857 ), .Z(n7839) );
  XOR \SUBBYTES[2].a/U4497  ( .A(n8314), .B(n8315), .Z(\SUBBYTES[2].a/w1877 )
         );
  XOR \SUBBYTES[2].a/U4496  ( .A(\w1[2][59] ), .B(n7840), .Z(n8318) );
  XOR \SUBBYTES[2].a/U4495  ( .A(\SUBBYTES[2].a/w1839 ), .B(
        \SUBBYTES[2].a/w1842 ), .Z(n7840) );
  XOR \SUBBYTES[2].a/U4494  ( .A(n7842), .B(n7841), .Z(\SUBBYTES[2].a/w1866 )
         );
  XOR \SUBBYTES[2].a/U4493  ( .A(n8318), .B(n7843), .Z(n7841) );
  XOR \SUBBYTES[2].a/U4492  ( .A(\w1[2][62] ), .B(\SUBBYTES[2].a/w1908 ), .Z(
        n7842) );
  XOR \SUBBYTES[2].a/U4491  ( .A(\SUBBYTES[2].a/w1847 ), .B(
        \SUBBYTES[2].a/w1848 ), .Z(n7843) );
  XOR \SUBBYTES[2].a/U4490  ( .A(n8316), .B(n8315), .Z(\SUBBYTES[2].a/w1886 )
         );
  XOR \SUBBYTES[2].a/U4489  ( .A(n7845), .B(n7844), .Z(\SUBBYTES[2].a/w1887 )
         );
  XOR \SUBBYTES[2].a/U4488  ( .A(\w1[2][63] ), .B(n8317), .Z(n7844) );
  XOR \SUBBYTES[2].a/U4487  ( .A(\SUBBYTES[2].a/w1839 ), .B(
        \SUBBYTES[2].a/w1848 ), .Z(n7845) );
  XOR \SUBBYTES[2].a/U4486  ( .A(n7847), .B(n7846), .Z(\SUBBYTES[2].a/w1863 )
         );
  XOR \SUBBYTES[2].a/U4485  ( .A(n7849), .B(n7848), .Z(n7846) );
  XOR \SUBBYTES[2].a/U4484  ( .A(\w1[2][63] ), .B(\SUBBYTES[2].a/w1947 ), .Z(
        n7847) );
  XOR \SUBBYTES[2].a/U4483  ( .A(\SUBBYTES[2].a/w1854 ), .B(
        \SUBBYTES[2].a/w1857 ), .Z(n7848) );
  XOR \SUBBYTES[2].a/U4482  ( .A(\SUBBYTES[2].a/w1840 ), .B(
        \SUBBYTES[2].a/w1842 ), .Z(n7849) );
  XOR \SUBBYTES[2].a/U4481  ( .A(n7851), .B(n7850), .Z(\SUBBYTES[2].a/w1864 )
         );
  XOR \SUBBYTES[2].a/U4480  ( .A(n8318), .B(n7852), .Z(n7850) );
  XOR \SUBBYTES[2].a/U4479  ( .A(\w1[2][61] ), .B(n8319), .Z(n7851) );
  XOR \SUBBYTES[2].a/U4478  ( .A(\SUBBYTES[2].a/w1854 ), .B(
        \SUBBYTES[2].a/w1855 ), .Z(n7852) );
  XOR \SUBBYTES[2].a/U4477  ( .A(n7854), .B(n7853), .Z(\SUBBYTES[2].a/w1880 )
         );
  XOR \SUBBYTES[2].a/U4476  ( .A(\w1[2][57] ), .B(n7855), .Z(n7853) );
  XOR \SUBBYTES[2].a/U4475  ( .A(\SUBBYTES[2].a/w1855 ), .B(
        \SUBBYTES[2].a/w1857 ), .Z(n7854) );
  XOR \SUBBYTES[2].a/U4474  ( .A(\SUBBYTES[2].a/w1839 ), .B(
        \SUBBYTES[2].a/w1840 ), .Z(n7855) );
  XOR \SUBBYTES[2].a/U4473  ( .A(\w1[2][65] ), .B(n7856), .Z(n8320) );
  XOR \SUBBYTES[2].a/U4472  ( .A(\w1[2][67] ), .B(\w1[2][66] ), .Z(n7856) );
  XOR \SUBBYTES[2].a/U4471  ( .A(\w1[2][70] ), .B(n8320), .Z(
        \SUBBYTES[2].a/w1722 ) );
  XOR \SUBBYTES[2].a/U4470  ( .A(\w1[2][64] ), .B(\SUBBYTES[2].a/w1722 ), .Z(
        \SUBBYTES[2].a/w1609 ) );
  XOR \SUBBYTES[2].a/U4469  ( .A(\w1[2][64] ), .B(n7857), .Z(
        \SUBBYTES[2].a/w1610 ) );
  XOR \SUBBYTES[2].a/U4468  ( .A(\w1[2][70] ), .B(\w1[2][69] ), .Z(n7857) );
  XOR \SUBBYTES[2].a/U4467  ( .A(\w1[2][69] ), .B(n8320), .Z(
        \SUBBYTES[2].a/w1740 ) );
  XOR \SUBBYTES[2].a/U4466  ( .A(n7859), .B(n7858), .Z(\SUBBYTES[2].a/w1733 )
         );
  XOR \SUBBYTES[2].a/U4465  ( .A(\w1[2][67] ), .B(\w1[2][65] ), .Z(n7858) );
  XOR \SUBBYTES[2].a/U4464  ( .A(\w1[2][71] ), .B(\w1[2][68] ), .Z(n7859) );
  XOR \SUBBYTES[2].a/U4463  ( .A(\w1[2][64] ), .B(\SUBBYTES[2].a/w1733 ), .Z(
        \SUBBYTES[2].a/w1612 ) );
  XOR \SUBBYTES[2].a/U4462  ( .A(n7861), .B(n7860), .Z(\SUBBYTES[2].a/w1720 )
         );
  XOR \SUBBYTES[2].a/U4461  ( .A(\SUBBYTES[2].a/w1681 ), .B(n980), .Z(n7860)
         );
  XOR \SUBBYTES[2].a/U4460  ( .A(\SUBBYTES[2].a/w1674 ), .B(
        \SUBBYTES[2].a/w1677 ), .Z(n7861) );
  XOR \SUBBYTES[2].a/U4459  ( .A(n7863), .B(n7862), .Z(\SUBBYTES[2].a/w1721 )
         );
  XOR \SUBBYTES[2].a/U4458  ( .A(\SUBBYTES[2].a/w1681 ), .B(n7127), .Z(n7862)
         );
  XOR \SUBBYTES[2].a/U4457  ( .A(\SUBBYTES[2].a/w1674 ), .B(n7126), .Z(n7863)
         );
  XOR \SUBBYTES[2].a/U4456  ( .A(\SUBBYTES[2].a/w1733 ), .B(n7864), .Z(
        \SUBBYTES[2].a/w1723 ) );
  XOR \SUBBYTES[2].a/U4455  ( .A(\w1[2][70] ), .B(\w1[2][69] ), .Z(n7864) );
  XOR \SUBBYTES[2].a/U4454  ( .A(n7866), .B(n7865), .Z(\SUBBYTES[2].a/w1724 )
         );
  XOR \SUBBYTES[2].a/U4453  ( .A(n7127), .B(n980), .Z(n7865) );
  XOR \SUBBYTES[2].a/U4452  ( .A(n7126), .B(\SUBBYTES[2].a/w1677 ), .Z(n7866)
         );
  XOR \SUBBYTES[2].a/U4451  ( .A(\w1[2][71] ), .B(\w1[2][66] ), .Z(n8326) );
  XOR \SUBBYTES[2].a/U4450  ( .A(n8326), .B(n7867), .Z(\SUBBYTES[2].a/w1725 )
         );
  XOR \SUBBYTES[2].a/U4449  ( .A(\w1[2][69] ), .B(\w1[2][68] ), .Z(n7867) );
  XOR \SUBBYTES[2].a/U4448  ( .A(\w1[2][71] ), .B(\SUBBYTES[2].a/w1610 ), .Z(
        \SUBBYTES[2].a/w1613 ) );
  XOR \SUBBYTES[2].a/U4447  ( .A(\w1[2][65] ), .B(\SUBBYTES[2].a/w1610 ), .Z(
        \SUBBYTES[2].a/w1614 ) );
  XOR \SUBBYTES[2].a/U4446  ( .A(\w1[2][68] ), .B(\SUBBYTES[2].a/w1610 ), .Z(
        \SUBBYTES[2].a/w1615 ) );
  XOR \SUBBYTES[2].a/U4445  ( .A(\SUBBYTES[2].a/w1614 ), .B(n8326), .Z(
        \SUBBYTES[2].a/w1616 ) );
  XOR \SUBBYTES[2].a/U4444  ( .A(n8326), .B(n7868), .Z(\SUBBYTES[2].a/w1701 )
         );
  XOR \SUBBYTES[2].a/U4443  ( .A(\w1[2][68] ), .B(\w1[2][65] ), .Z(n7868) );
  XOR \SUBBYTES[2].a/U4442  ( .A(n7870), .B(n7869), .Z(n8323) );
  XOR \SUBBYTES[2].a/U4441  ( .A(\w1[2][68] ), .B(n7871), .Z(n7869) );
  XOR \SUBBYTES[2].a/U4440  ( .A(\SUBBYTES[2].a/w1666 ), .B(\w1[2][70] ), .Z(
        n7870) );
  XOR \SUBBYTES[2].a/U4439  ( .A(\SUBBYTES[2].a/w1640 ), .B(
        \SUBBYTES[2].a/w1647 ), .Z(n7871) );
  XOR \SUBBYTES[2].a/U4438  ( .A(n7873), .B(n7872), .Z(n8321) );
  XOR \SUBBYTES[2].a/U4437  ( .A(\w1[2][65] ), .B(n7874), .Z(n7872) );
  XOR \SUBBYTES[2].a/U4436  ( .A(\SUBBYTES[2].a/w1665 ), .B(\w1[2][69] ), .Z(
        n7873) );
  XOR \SUBBYTES[2].a/U4435  ( .A(\SUBBYTES[2].a/w1641 ), .B(
        \SUBBYTES[2].a/w1648 ), .Z(n7874) );
  XOR \SUBBYTES[2].a/U4434  ( .A(n8323), .B(n8321), .Z(\SUBBYTES[2].a/w1671 )
         );
  XOR \SUBBYTES[2].a/U4433  ( .A(\w1[2][69] ), .B(n7875), .Z(n8324) );
  XOR \SUBBYTES[2].a/U4432  ( .A(\SUBBYTES[2].a/w1633 ), .B(
        \SUBBYTES[2].a/w1643 ), .Z(n7875) );
  XOR \SUBBYTES[2].a/U4431  ( .A(n7877), .B(n7876), .Z(\SUBBYTES[2].a/w1658 )
         );
  XOR \SUBBYTES[2].a/U4430  ( .A(n8324), .B(n7878), .Z(n7876) );
  XOR \SUBBYTES[2].a/U4429  ( .A(\w1[2][68] ), .B(\SUBBYTES[2].a/w1722 ), .Z(
        n7877) );
  XOR \SUBBYTES[2].a/U4428  ( .A(\SUBBYTES[2].a/w1635 ), .B(
        \SUBBYTES[2].a/w1640 ), .Z(n7878) );
  XOR \SUBBYTES[2].a/U4427  ( .A(n7880), .B(n7879), .Z(n8322) );
  XOR \SUBBYTES[2].a/U4426  ( .A(\SUBBYTES[2].a/w1668 ), .B(\w1[2][71] ), .Z(
        n7879) );
  XOR \SUBBYTES[2].a/U4425  ( .A(\SUBBYTES[2].a/w1643 ), .B(
        \SUBBYTES[2].a/w1650 ), .Z(n7880) );
  XOR \SUBBYTES[2].a/U4424  ( .A(n8321), .B(n8322), .Z(\SUBBYTES[2].a/w1670 )
         );
  XOR \SUBBYTES[2].a/U4423  ( .A(\w1[2][67] ), .B(n7881), .Z(n8325) );
  XOR \SUBBYTES[2].a/U4422  ( .A(\SUBBYTES[2].a/w1632 ), .B(
        \SUBBYTES[2].a/w1635 ), .Z(n7881) );
  XOR \SUBBYTES[2].a/U4421  ( .A(n7883), .B(n7882), .Z(\SUBBYTES[2].a/w1659 )
         );
  XOR \SUBBYTES[2].a/U4420  ( .A(n8325), .B(n7884), .Z(n7882) );
  XOR \SUBBYTES[2].a/U4419  ( .A(\w1[2][70] ), .B(\SUBBYTES[2].a/w1701 ), .Z(
        n7883) );
  XOR \SUBBYTES[2].a/U4418  ( .A(\SUBBYTES[2].a/w1640 ), .B(
        \SUBBYTES[2].a/w1641 ), .Z(n7884) );
  XOR \SUBBYTES[2].a/U4417  ( .A(n8323), .B(n8322), .Z(\SUBBYTES[2].a/w1679 )
         );
  XOR \SUBBYTES[2].a/U4416  ( .A(n7886), .B(n7885), .Z(\SUBBYTES[2].a/w1680 )
         );
  XOR \SUBBYTES[2].a/U4415  ( .A(\w1[2][71] ), .B(n8324), .Z(n7885) );
  XOR \SUBBYTES[2].a/U4414  ( .A(\SUBBYTES[2].a/w1632 ), .B(
        \SUBBYTES[2].a/w1641 ), .Z(n7886) );
  XOR \SUBBYTES[2].a/U4413  ( .A(n7888), .B(n7887), .Z(\SUBBYTES[2].a/w1656 )
         );
  XOR \SUBBYTES[2].a/U4412  ( .A(n7890), .B(n7889), .Z(n7887) );
  XOR \SUBBYTES[2].a/U4411  ( .A(\w1[2][71] ), .B(\SUBBYTES[2].a/w1740 ), .Z(
        n7888) );
  XOR \SUBBYTES[2].a/U4410  ( .A(\SUBBYTES[2].a/w1647 ), .B(
        \SUBBYTES[2].a/w1650 ), .Z(n7889) );
  XOR \SUBBYTES[2].a/U4409  ( .A(\SUBBYTES[2].a/w1633 ), .B(
        \SUBBYTES[2].a/w1635 ), .Z(n7890) );
  XOR \SUBBYTES[2].a/U4408  ( .A(n7892), .B(n7891), .Z(\SUBBYTES[2].a/w1657 )
         );
  XOR \SUBBYTES[2].a/U4407  ( .A(n8325), .B(n7893), .Z(n7891) );
  XOR \SUBBYTES[2].a/U4406  ( .A(\w1[2][69] ), .B(n8326), .Z(n7892) );
  XOR \SUBBYTES[2].a/U4405  ( .A(\SUBBYTES[2].a/w1647 ), .B(
        \SUBBYTES[2].a/w1648 ), .Z(n7893) );
  XOR \SUBBYTES[2].a/U4404  ( .A(n7895), .B(n7894), .Z(\SUBBYTES[2].a/w1673 )
         );
  XOR \SUBBYTES[2].a/U4403  ( .A(\w1[2][65] ), .B(n7896), .Z(n7894) );
  XOR \SUBBYTES[2].a/U4402  ( .A(\SUBBYTES[2].a/w1648 ), .B(
        \SUBBYTES[2].a/w1650 ), .Z(n7895) );
  XOR \SUBBYTES[2].a/U4401  ( .A(\SUBBYTES[2].a/w1632 ), .B(
        \SUBBYTES[2].a/w1633 ), .Z(n7896) );
  XOR \SUBBYTES[2].a/U4400  ( .A(\w1[2][73] ), .B(n7897), .Z(n8327) );
  XOR \SUBBYTES[2].a/U4399  ( .A(\w1[2][75] ), .B(\w1[2][74] ), .Z(n7897) );
  XOR \SUBBYTES[2].a/U4398  ( .A(\w1[2][78] ), .B(n8327), .Z(
        \SUBBYTES[2].a/w1515 ) );
  XOR \SUBBYTES[2].a/U4397  ( .A(\w1[2][72] ), .B(\SUBBYTES[2].a/w1515 ), .Z(
        \SUBBYTES[2].a/w1402 ) );
  XOR \SUBBYTES[2].a/U4396  ( .A(\w1[2][72] ), .B(n7898), .Z(
        \SUBBYTES[2].a/w1403 ) );
  XOR \SUBBYTES[2].a/U4395  ( .A(\w1[2][78] ), .B(\w1[2][77] ), .Z(n7898) );
  XOR \SUBBYTES[2].a/U4394  ( .A(\w1[2][77] ), .B(n8327), .Z(
        \SUBBYTES[2].a/w1533 ) );
  XOR \SUBBYTES[2].a/U4393  ( .A(n7900), .B(n7899), .Z(\SUBBYTES[2].a/w1526 )
         );
  XOR \SUBBYTES[2].a/U4392  ( .A(\w1[2][75] ), .B(\w1[2][73] ), .Z(n7899) );
  XOR \SUBBYTES[2].a/U4391  ( .A(\w1[2][79] ), .B(\w1[2][76] ), .Z(n7900) );
  XOR \SUBBYTES[2].a/U4390  ( .A(\w1[2][72] ), .B(\SUBBYTES[2].a/w1526 ), .Z(
        \SUBBYTES[2].a/w1405 ) );
  XOR \SUBBYTES[2].a/U4389  ( .A(n7902), .B(n7901), .Z(\SUBBYTES[2].a/w1513 )
         );
  XOR \SUBBYTES[2].a/U4388  ( .A(\SUBBYTES[2].a/w1474 ), .B(n979), .Z(n7901)
         );
  XOR \SUBBYTES[2].a/U4387  ( .A(\SUBBYTES[2].a/w1467 ), .B(
        \SUBBYTES[2].a/w1470 ), .Z(n7902) );
  XOR \SUBBYTES[2].a/U4386  ( .A(n7904), .B(n7903), .Z(\SUBBYTES[2].a/w1514 )
         );
  XOR \SUBBYTES[2].a/U4385  ( .A(\SUBBYTES[2].a/w1474 ), .B(n7125), .Z(n7903)
         );
  XOR \SUBBYTES[2].a/U4384  ( .A(\SUBBYTES[2].a/w1467 ), .B(n7124), .Z(n7904)
         );
  XOR \SUBBYTES[2].a/U4383  ( .A(\SUBBYTES[2].a/w1526 ), .B(n7905), .Z(
        \SUBBYTES[2].a/w1516 ) );
  XOR \SUBBYTES[2].a/U4382  ( .A(\w1[2][78] ), .B(\w1[2][77] ), .Z(n7905) );
  XOR \SUBBYTES[2].a/U4381  ( .A(n7907), .B(n7906), .Z(\SUBBYTES[2].a/w1517 )
         );
  XOR \SUBBYTES[2].a/U4380  ( .A(n7125), .B(n979), .Z(n7906) );
  XOR \SUBBYTES[2].a/U4379  ( .A(n7124), .B(\SUBBYTES[2].a/w1470 ), .Z(n7907)
         );
  XOR \SUBBYTES[2].a/U4378  ( .A(\w1[2][79] ), .B(\w1[2][74] ), .Z(n8333) );
  XOR \SUBBYTES[2].a/U4377  ( .A(n8333), .B(n7908), .Z(\SUBBYTES[2].a/w1518 )
         );
  XOR \SUBBYTES[2].a/U4376  ( .A(\w1[2][77] ), .B(\w1[2][76] ), .Z(n7908) );
  XOR \SUBBYTES[2].a/U4375  ( .A(\w1[2][79] ), .B(\SUBBYTES[2].a/w1403 ), .Z(
        \SUBBYTES[2].a/w1406 ) );
  XOR \SUBBYTES[2].a/U4374  ( .A(\w1[2][73] ), .B(\SUBBYTES[2].a/w1403 ), .Z(
        \SUBBYTES[2].a/w1407 ) );
  XOR \SUBBYTES[2].a/U4373  ( .A(\w1[2][76] ), .B(\SUBBYTES[2].a/w1403 ), .Z(
        \SUBBYTES[2].a/w1408 ) );
  XOR \SUBBYTES[2].a/U4372  ( .A(\SUBBYTES[2].a/w1407 ), .B(n8333), .Z(
        \SUBBYTES[2].a/w1409 ) );
  XOR \SUBBYTES[2].a/U4371  ( .A(n8333), .B(n7909), .Z(\SUBBYTES[2].a/w1494 )
         );
  XOR \SUBBYTES[2].a/U4370  ( .A(\w1[2][76] ), .B(\w1[2][73] ), .Z(n7909) );
  XOR \SUBBYTES[2].a/U4369  ( .A(n7911), .B(n7910), .Z(n8330) );
  XOR \SUBBYTES[2].a/U4368  ( .A(\w1[2][76] ), .B(n7912), .Z(n7910) );
  XOR \SUBBYTES[2].a/U4367  ( .A(\SUBBYTES[2].a/w1459 ), .B(\w1[2][78] ), .Z(
        n7911) );
  XOR \SUBBYTES[2].a/U4366  ( .A(\SUBBYTES[2].a/w1433 ), .B(
        \SUBBYTES[2].a/w1440 ), .Z(n7912) );
  XOR \SUBBYTES[2].a/U4365  ( .A(n7914), .B(n7913), .Z(n8328) );
  XOR \SUBBYTES[2].a/U4364  ( .A(\w1[2][73] ), .B(n7915), .Z(n7913) );
  XOR \SUBBYTES[2].a/U4363  ( .A(\SUBBYTES[2].a/w1458 ), .B(\w1[2][77] ), .Z(
        n7914) );
  XOR \SUBBYTES[2].a/U4362  ( .A(\SUBBYTES[2].a/w1434 ), .B(
        \SUBBYTES[2].a/w1441 ), .Z(n7915) );
  XOR \SUBBYTES[2].a/U4361  ( .A(n8330), .B(n8328), .Z(\SUBBYTES[2].a/w1464 )
         );
  XOR \SUBBYTES[2].a/U4360  ( .A(\w1[2][77] ), .B(n7916), .Z(n8331) );
  XOR \SUBBYTES[2].a/U4359  ( .A(\SUBBYTES[2].a/w1426 ), .B(
        \SUBBYTES[2].a/w1436 ), .Z(n7916) );
  XOR \SUBBYTES[2].a/U4358  ( .A(n7918), .B(n7917), .Z(\SUBBYTES[2].a/w1451 )
         );
  XOR \SUBBYTES[2].a/U4357  ( .A(n8331), .B(n7919), .Z(n7917) );
  XOR \SUBBYTES[2].a/U4356  ( .A(\w1[2][76] ), .B(\SUBBYTES[2].a/w1515 ), .Z(
        n7918) );
  XOR \SUBBYTES[2].a/U4355  ( .A(\SUBBYTES[2].a/w1428 ), .B(
        \SUBBYTES[2].a/w1433 ), .Z(n7919) );
  XOR \SUBBYTES[2].a/U4354  ( .A(n7921), .B(n7920), .Z(n8329) );
  XOR \SUBBYTES[2].a/U4353  ( .A(\SUBBYTES[2].a/w1461 ), .B(\w1[2][79] ), .Z(
        n7920) );
  XOR \SUBBYTES[2].a/U4352  ( .A(\SUBBYTES[2].a/w1436 ), .B(
        \SUBBYTES[2].a/w1443 ), .Z(n7921) );
  XOR \SUBBYTES[2].a/U4351  ( .A(n8328), .B(n8329), .Z(\SUBBYTES[2].a/w1463 )
         );
  XOR \SUBBYTES[2].a/U4350  ( .A(\w1[2][75] ), .B(n7922), .Z(n8332) );
  XOR \SUBBYTES[2].a/U4349  ( .A(\SUBBYTES[2].a/w1425 ), .B(
        \SUBBYTES[2].a/w1428 ), .Z(n7922) );
  XOR \SUBBYTES[2].a/U4348  ( .A(n7924), .B(n7923), .Z(\SUBBYTES[2].a/w1452 )
         );
  XOR \SUBBYTES[2].a/U4347  ( .A(n8332), .B(n7925), .Z(n7923) );
  XOR \SUBBYTES[2].a/U4346  ( .A(\w1[2][78] ), .B(\SUBBYTES[2].a/w1494 ), .Z(
        n7924) );
  XOR \SUBBYTES[2].a/U4345  ( .A(\SUBBYTES[2].a/w1433 ), .B(
        \SUBBYTES[2].a/w1434 ), .Z(n7925) );
  XOR \SUBBYTES[2].a/U4344  ( .A(n8330), .B(n8329), .Z(\SUBBYTES[2].a/w1472 )
         );
  XOR \SUBBYTES[2].a/U4343  ( .A(n7927), .B(n7926), .Z(\SUBBYTES[2].a/w1473 )
         );
  XOR \SUBBYTES[2].a/U4342  ( .A(\w1[2][79] ), .B(n8331), .Z(n7926) );
  XOR \SUBBYTES[2].a/U4341  ( .A(\SUBBYTES[2].a/w1425 ), .B(
        \SUBBYTES[2].a/w1434 ), .Z(n7927) );
  XOR \SUBBYTES[2].a/U4340  ( .A(n7929), .B(n7928), .Z(\SUBBYTES[2].a/w1449 )
         );
  XOR \SUBBYTES[2].a/U4339  ( .A(n7931), .B(n7930), .Z(n7928) );
  XOR \SUBBYTES[2].a/U4338  ( .A(\w1[2][79] ), .B(\SUBBYTES[2].a/w1533 ), .Z(
        n7929) );
  XOR \SUBBYTES[2].a/U4337  ( .A(\SUBBYTES[2].a/w1440 ), .B(
        \SUBBYTES[2].a/w1443 ), .Z(n7930) );
  XOR \SUBBYTES[2].a/U4336  ( .A(\SUBBYTES[2].a/w1426 ), .B(
        \SUBBYTES[2].a/w1428 ), .Z(n7931) );
  XOR \SUBBYTES[2].a/U4335  ( .A(n7933), .B(n7932), .Z(\SUBBYTES[2].a/w1450 )
         );
  XOR \SUBBYTES[2].a/U4334  ( .A(n8332), .B(n7934), .Z(n7932) );
  XOR \SUBBYTES[2].a/U4333  ( .A(\w1[2][77] ), .B(n8333), .Z(n7933) );
  XOR \SUBBYTES[2].a/U4332  ( .A(\SUBBYTES[2].a/w1440 ), .B(
        \SUBBYTES[2].a/w1441 ), .Z(n7934) );
  XOR \SUBBYTES[2].a/U4331  ( .A(n7936), .B(n7935), .Z(\SUBBYTES[2].a/w1466 )
         );
  XOR \SUBBYTES[2].a/U4330  ( .A(\w1[2][73] ), .B(n7937), .Z(n7935) );
  XOR \SUBBYTES[2].a/U4329  ( .A(\SUBBYTES[2].a/w1441 ), .B(
        \SUBBYTES[2].a/w1443 ), .Z(n7936) );
  XOR \SUBBYTES[2].a/U4328  ( .A(\SUBBYTES[2].a/w1425 ), .B(
        \SUBBYTES[2].a/w1426 ), .Z(n7937) );
  XOR \SUBBYTES[2].a/U4327  ( .A(\w1[2][81] ), .B(n7938), .Z(n8334) );
  XOR \SUBBYTES[2].a/U4326  ( .A(\w1[2][83] ), .B(\w1[2][82] ), .Z(n7938) );
  XOR \SUBBYTES[2].a/U4325  ( .A(\w1[2][86] ), .B(n8334), .Z(
        \SUBBYTES[2].a/w1308 ) );
  XOR \SUBBYTES[2].a/U4324  ( .A(\w1[2][80] ), .B(\SUBBYTES[2].a/w1308 ), .Z(
        \SUBBYTES[2].a/w1195 ) );
  XOR \SUBBYTES[2].a/U4323  ( .A(\w1[2][80] ), .B(n7939), .Z(
        \SUBBYTES[2].a/w1196 ) );
  XOR \SUBBYTES[2].a/U4322  ( .A(\w1[2][86] ), .B(\w1[2][85] ), .Z(n7939) );
  XOR \SUBBYTES[2].a/U4321  ( .A(\w1[2][85] ), .B(n8334), .Z(
        \SUBBYTES[2].a/w1326 ) );
  XOR \SUBBYTES[2].a/U4320  ( .A(n7941), .B(n7940), .Z(\SUBBYTES[2].a/w1319 )
         );
  XOR \SUBBYTES[2].a/U4319  ( .A(\w1[2][83] ), .B(\w1[2][81] ), .Z(n7940) );
  XOR \SUBBYTES[2].a/U4318  ( .A(\w1[2][87] ), .B(\w1[2][84] ), .Z(n7941) );
  XOR \SUBBYTES[2].a/U4317  ( .A(\w1[2][80] ), .B(\SUBBYTES[2].a/w1319 ), .Z(
        \SUBBYTES[2].a/w1198 ) );
  XOR \SUBBYTES[2].a/U4316  ( .A(n7943), .B(n7942), .Z(\SUBBYTES[2].a/w1306 )
         );
  XOR \SUBBYTES[2].a/U4315  ( .A(\SUBBYTES[2].a/w1267 ), .B(n978), .Z(n7942)
         );
  XOR \SUBBYTES[2].a/U4314  ( .A(\SUBBYTES[2].a/w1260 ), .B(
        \SUBBYTES[2].a/w1263 ), .Z(n7943) );
  XOR \SUBBYTES[2].a/U4313  ( .A(n7945), .B(n7944), .Z(\SUBBYTES[2].a/w1307 )
         );
  XOR \SUBBYTES[2].a/U4312  ( .A(\SUBBYTES[2].a/w1267 ), .B(n7123), .Z(n7944)
         );
  XOR \SUBBYTES[2].a/U4311  ( .A(\SUBBYTES[2].a/w1260 ), .B(n7122), .Z(n7945)
         );
  XOR \SUBBYTES[2].a/U4310  ( .A(\SUBBYTES[2].a/w1319 ), .B(n7946), .Z(
        \SUBBYTES[2].a/w1309 ) );
  XOR \SUBBYTES[2].a/U4309  ( .A(\w1[2][86] ), .B(\w1[2][85] ), .Z(n7946) );
  XOR \SUBBYTES[2].a/U4308  ( .A(n7948), .B(n7947), .Z(\SUBBYTES[2].a/w1310 )
         );
  XOR \SUBBYTES[2].a/U4307  ( .A(n7123), .B(n978), .Z(n7947) );
  XOR \SUBBYTES[2].a/U4306  ( .A(n7122), .B(\SUBBYTES[2].a/w1263 ), .Z(n7948)
         );
  XOR \SUBBYTES[2].a/U4305  ( .A(\w1[2][87] ), .B(\w1[2][82] ), .Z(n8340) );
  XOR \SUBBYTES[2].a/U4304  ( .A(n8340), .B(n7949), .Z(\SUBBYTES[2].a/w1311 )
         );
  XOR \SUBBYTES[2].a/U4303  ( .A(\w1[2][85] ), .B(\w1[2][84] ), .Z(n7949) );
  XOR \SUBBYTES[2].a/U4302  ( .A(\w1[2][87] ), .B(\SUBBYTES[2].a/w1196 ), .Z(
        \SUBBYTES[2].a/w1199 ) );
  XOR \SUBBYTES[2].a/U4301  ( .A(\w1[2][81] ), .B(\SUBBYTES[2].a/w1196 ), .Z(
        \SUBBYTES[2].a/w1200 ) );
  XOR \SUBBYTES[2].a/U4300  ( .A(\w1[2][84] ), .B(\SUBBYTES[2].a/w1196 ), .Z(
        \SUBBYTES[2].a/w1201 ) );
  XOR \SUBBYTES[2].a/U4299  ( .A(\SUBBYTES[2].a/w1200 ), .B(n8340), .Z(
        \SUBBYTES[2].a/w1202 ) );
  XOR \SUBBYTES[2].a/U4298  ( .A(n8340), .B(n7950), .Z(\SUBBYTES[2].a/w1287 )
         );
  XOR \SUBBYTES[2].a/U4297  ( .A(\w1[2][84] ), .B(\w1[2][81] ), .Z(n7950) );
  XOR \SUBBYTES[2].a/U4296  ( .A(n7952), .B(n7951), .Z(n8337) );
  XOR \SUBBYTES[2].a/U4295  ( .A(\w1[2][84] ), .B(n7953), .Z(n7951) );
  XOR \SUBBYTES[2].a/U4294  ( .A(\SUBBYTES[2].a/w1252 ), .B(\w1[2][86] ), .Z(
        n7952) );
  XOR \SUBBYTES[2].a/U4293  ( .A(\SUBBYTES[2].a/w1226 ), .B(
        \SUBBYTES[2].a/w1233 ), .Z(n7953) );
  XOR \SUBBYTES[2].a/U4292  ( .A(n7955), .B(n7954), .Z(n8335) );
  XOR \SUBBYTES[2].a/U4291  ( .A(\w1[2][81] ), .B(n7956), .Z(n7954) );
  XOR \SUBBYTES[2].a/U4290  ( .A(\SUBBYTES[2].a/w1251 ), .B(\w1[2][85] ), .Z(
        n7955) );
  XOR \SUBBYTES[2].a/U4289  ( .A(\SUBBYTES[2].a/w1227 ), .B(
        \SUBBYTES[2].a/w1234 ), .Z(n7956) );
  XOR \SUBBYTES[2].a/U4288  ( .A(n8337), .B(n8335), .Z(\SUBBYTES[2].a/w1257 )
         );
  XOR \SUBBYTES[2].a/U4287  ( .A(\w1[2][85] ), .B(n7957), .Z(n8338) );
  XOR \SUBBYTES[2].a/U4286  ( .A(\SUBBYTES[2].a/w1219 ), .B(
        \SUBBYTES[2].a/w1229 ), .Z(n7957) );
  XOR \SUBBYTES[2].a/U4285  ( .A(n7959), .B(n7958), .Z(\SUBBYTES[2].a/w1244 )
         );
  XOR \SUBBYTES[2].a/U4284  ( .A(n8338), .B(n7960), .Z(n7958) );
  XOR \SUBBYTES[2].a/U4283  ( .A(\w1[2][84] ), .B(\SUBBYTES[2].a/w1308 ), .Z(
        n7959) );
  XOR \SUBBYTES[2].a/U4282  ( .A(\SUBBYTES[2].a/w1221 ), .B(
        \SUBBYTES[2].a/w1226 ), .Z(n7960) );
  XOR \SUBBYTES[2].a/U4281  ( .A(n7962), .B(n7961), .Z(n8336) );
  XOR \SUBBYTES[2].a/U4280  ( .A(\SUBBYTES[2].a/w1254 ), .B(\w1[2][87] ), .Z(
        n7961) );
  XOR \SUBBYTES[2].a/U4279  ( .A(\SUBBYTES[2].a/w1229 ), .B(
        \SUBBYTES[2].a/w1236 ), .Z(n7962) );
  XOR \SUBBYTES[2].a/U4278  ( .A(n8335), .B(n8336), .Z(\SUBBYTES[2].a/w1256 )
         );
  XOR \SUBBYTES[2].a/U4277  ( .A(\w1[2][83] ), .B(n7963), .Z(n8339) );
  XOR \SUBBYTES[2].a/U4276  ( .A(\SUBBYTES[2].a/w1218 ), .B(
        \SUBBYTES[2].a/w1221 ), .Z(n7963) );
  XOR \SUBBYTES[2].a/U4275  ( .A(n7965), .B(n7964), .Z(\SUBBYTES[2].a/w1245 )
         );
  XOR \SUBBYTES[2].a/U4274  ( .A(n8339), .B(n7966), .Z(n7964) );
  XOR \SUBBYTES[2].a/U4273  ( .A(\w1[2][86] ), .B(\SUBBYTES[2].a/w1287 ), .Z(
        n7965) );
  XOR \SUBBYTES[2].a/U4272  ( .A(\SUBBYTES[2].a/w1226 ), .B(
        \SUBBYTES[2].a/w1227 ), .Z(n7966) );
  XOR \SUBBYTES[2].a/U4271  ( .A(n8337), .B(n8336), .Z(\SUBBYTES[2].a/w1265 )
         );
  XOR \SUBBYTES[2].a/U4270  ( .A(n7968), .B(n7967), .Z(\SUBBYTES[2].a/w1266 )
         );
  XOR \SUBBYTES[2].a/U4269  ( .A(\w1[2][87] ), .B(n8338), .Z(n7967) );
  XOR \SUBBYTES[2].a/U4268  ( .A(\SUBBYTES[2].a/w1218 ), .B(
        \SUBBYTES[2].a/w1227 ), .Z(n7968) );
  XOR \SUBBYTES[2].a/U4267  ( .A(n7970), .B(n7969), .Z(\SUBBYTES[2].a/w1242 )
         );
  XOR \SUBBYTES[2].a/U4266  ( .A(n7972), .B(n7971), .Z(n7969) );
  XOR \SUBBYTES[2].a/U4265  ( .A(\w1[2][87] ), .B(\SUBBYTES[2].a/w1326 ), .Z(
        n7970) );
  XOR \SUBBYTES[2].a/U4264  ( .A(\SUBBYTES[2].a/w1233 ), .B(
        \SUBBYTES[2].a/w1236 ), .Z(n7971) );
  XOR \SUBBYTES[2].a/U4263  ( .A(\SUBBYTES[2].a/w1219 ), .B(
        \SUBBYTES[2].a/w1221 ), .Z(n7972) );
  XOR \SUBBYTES[2].a/U4262  ( .A(n7974), .B(n7973), .Z(\SUBBYTES[2].a/w1243 )
         );
  XOR \SUBBYTES[2].a/U4261  ( .A(n8339), .B(n7975), .Z(n7973) );
  XOR \SUBBYTES[2].a/U4260  ( .A(\w1[2][85] ), .B(n8340), .Z(n7974) );
  XOR \SUBBYTES[2].a/U4259  ( .A(\SUBBYTES[2].a/w1233 ), .B(
        \SUBBYTES[2].a/w1234 ), .Z(n7975) );
  XOR \SUBBYTES[2].a/U4258  ( .A(n7977), .B(n7976), .Z(\SUBBYTES[2].a/w1259 )
         );
  XOR \SUBBYTES[2].a/U4257  ( .A(\w1[2][81] ), .B(n7978), .Z(n7976) );
  XOR \SUBBYTES[2].a/U4256  ( .A(\SUBBYTES[2].a/w1234 ), .B(
        \SUBBYTES[2].a/w1236 ), .Z(n7977) );
  XOR \SUBBYTES[2].a/U4255  ( .A(\SUBBYTES[2].a/w1218 ), .B(
        \SUBBYTES[2].a/w1219 ), .Z(n7978) );
  XOR \SUBBYTES[2].a/U4254  ( .A(\w1[2][89] ), .B(n7979), .Z(n8341) );
  XOR \SUBBYTES[2].a/U4253  ( .A(\w1[2][91] ), .B(\w1[2][90] ), .Z(n7979) );
  XOR \SUBBYTES[2].a/U4252  ( .A(\w1[2][94] ), .B(n8341), .Z(
        \SUBBYTES[2].a/w1101 ) );
  XOR \SUBBYTES[2].a/U4251  ( .A(\w1[2][88] ), .B(\SUBBYTES[2].a/w1101 ), .Z(
        \SUBBYTES[2].a/w988 ) );
  XOR \SUBBYTES[2].a/U4250  ( .A(\w1[2][88] ), .B(n7980), .Z(
        \SUBBYTES[2].a/w989 ) );
  XOR \SUBBYTES[2].a/U4249  ( .A(\w1[2][94] ), .B(\w1[2][93] ), .Z(n7980) );
  XOR \SUBBYTES[2].a/U4248  ( .A(\w1[2][93] ), .B(n8341), .Z(
        \SUBBYTES[2].a/w1119 ) );
  XOR \SUBBYTES[2].a/U4247  ( .A(n7982), .B(n7981), .Z(\SUBBYTES[2].a/w1112 )
         );
  XOR \SUBBYTES[2].a/U4246  ( .A(\w1[2][91] ), .B(\w1[2][89] ), .Z(n7981) );
  XOR \SUBBYTES[2].a/U4245  ( .A(\w1[2][95] ), .B(\w1[2][92] ), .Z(n7982) );
  XOR \SUBBYTES[2].a/U4244  ( .A(\w1[2][88] ), .B(\SUBBYTES[2].a/w1112 ), .Z(
        \SUBBYTES[2].a/w991 ) );
  XOR \SUBBYTES[2].a/U4243  ( .A(n7984), .B(n7983), .Z(\SUBBYTES[2].a/w1099 )
         );
  XOR \SUBBYTES[2].a/U4242  ( .A(\SUBBYTES[2].a/w1060 ), .B(n977), .Z(n7983)
         );
  XOR \SUBBYTES[2].a/U4241  ( .A(\SUBBYTES[2].a/w1053 ), .B(
        \SUBBYTES[2].a/w1056 ), .Z(n7984) );
  XOR \SUBBYTES[2].a/U4240  ( .A(n7986), .B(n7985), .Z(\SUBBYTES[2].a/w1100 )
         );
  XOR \SUBBYTES[2].a/U4239  ( .A(\SUBBYTES[2].a/w1060 ), .B(n7121), .Z(n7985)
         );
  XOR \SUBBYTES[2].a/U4238  ( .A(\SUBBYTES[2].a/w1053 ), .B(n7120), .Z(n7986)
         );
  XOR \SUBBYTES[2].a/U4237  ( .A(\SUBBYTES[2].a/w1112 ), .B(n7987), .Z(
        \SUBBYTES[2].a/w1102 ) );
  XOR \SUBBYTES[2].a/U4236  ( .A(\w1[2][94] ), .B(\w1[2][93] ), .Z(n7987) );
  XOR \SUBBYTES[2].a/U4235  ( .A(n7989), .B(n7988), .Z(\SUBBYTES[2].a/w1103 )
         );
  XOR \SUBBYTES[2].a/U4234  ( .A(n7121), .B(n977), .Z(n7988) );
  XOR \SUBBYTES[2].a/U4233  ( .A(n7120), .B(\SUBBYTES[2].a/w1056 ), .Z(n7989)
         );
  XOR \SUBBYTES[2].a/U4232  ( .A(\w1[2][95] ), .B(\w1[2][90] ), .Z(n8347) );
  XOR \SUBBYTES[2].a/U4231  ( .A(n8347), .B(n7990), .Z(\SUBBYTES[2].a/w1104 )
         );
  XOR \SUBBYTES[2].a/U4230  ( .A(\w1[2][93] ), .B(\w1[2][92] ), .Z(n7990) );
  XOR \SUBBYTES[2].a/U4229  ( .A(\w1[2][95] ), .B(\SUBBYTES[2].a/w989 ), .Z(
        \SUBBYTES[2].a/w992 ) );
  XOR \SUBBYTES[2].a/U4228  ( .A(\w1[2][89] ), .B(\SUBBYTES[2].a/w989 ), .Z(
        \SUBBYTES[2].a/w993 ) );
  XOR \SUBBYTES[2].a/U4227  ( .A(\w1[2][92] ), .B(\SUBBYTES[2].a/w989 ), .Z(
        \SUBBYTES[2].a/w994 ) );
  XOR \SUBBYTES[2].a/U4226  ( .A(\SUBBYTES[2].a/w993 ), .B(n8347), .Z(
        \SUBBYTES[2].a/w995 ) );
  XOR \SUBBYTES[2].a/U4225  ( .A(n8347), .B(n7991), .Z(\SUBBYTES[2].a/w1080 )
         );
  XOR \SUBBYTES[2].a/U4224  ( .A(\w1[2][92] ), .B(\w1[2][89] ), .Z(n7991) );
  XOR \SUBBYTES[2].a/U4223  ( .A(n7993), .B(n7992), .Z(n8344) );
  XOR \SUBBYTES[2].a/U4222  ( .A(\w1[2][92] ), .B(n7994), .Z(n7992) );
  XOR \SUBBYTES[2].a/U4221  ( .A(\SUBBYTES[2].a/w1045 ), .B(\w1[2][94] ), .Z(
        n7993) );
  XOR \SUBBYTES[2].a/U4220  ( .A(\SUBBYTES[2].a/w1019 ), .B(
        \SUBBYTES[2].a/w1026 ), .Z(n7994) );
  XOR \SUBBYTES[2].a/U4219  ( .A(n7996), .B(n7995), .Z(n8342) );
  XOR \SUBBYTES[2].a/U4218  ( .A(\w1[2][89] ), .B(n7997), .Z(n7995) );
  XOR \SUBBYTES[2].a/U4217  ( .A(\SUBBYTES[2].a/w1044 ), .B(\w1[2][93] ), .Z(
        n7996) );
  XOR \SUBBYTES[2].a/U4216  ( .A(\SUBBYTES[2].a/w1020 ), .B(
        \SUBBYTES[2].a/w1027 ), .Z(n7997) );
  XOR \SUBBYTES[2].a/U4215  ( .A(n8344), .B(n8342), .Z(\SUBBYTES[2].a/w1050 )
         );
  XOR \SUBBYTES[2].a/U4214  ( .A(\w1[2][93] ), .B(n7998), .Z(n8345) );
  XOR \SUBBYTES[2].a/U4213  ( .A(\SUBBYTES[2].a/w1012 ), .B(
        \SUBBYTES[2].a/w1022 ), .Z(n7998) );
  XOR \SUBBYTES[2].a/U4212  ( .A(n8000), .B(n7999), .Z(\SUBBYTES[2].a/w1037 )
         );
  XOR \SUBBYTES[2].a/U4211  ( .A(n8345), .B(n8001), .Z(n7999) );
  XOR \SUBBYTES[2].a/U4210  ( .A(\w1[2][92] ), .B(\SUBBYTES[2].a/w1101 ), .Z(
        n8000) );
  XOR \SUBBYTES[2].a/U4209  ( .A(\SUBBYTES[2].a/w1014 ), .B(
        \SUBBYTES[2].a/w1019 ), .Z(n8001) );
  XOR \SUBBYTES[2].a/U4208  ( .A(n8003), .B(n8002), .Z(n8343) );
  XOR \SUBBYTES[2].a/U4207  ( .A(\SUBBYTES[2].a/w1047 ), .B(\w1[2][95] ), .Z(
        n8002) );
  XOR \SUBBYTES[2].a/U4206  ( .A(\SUBBYTES[2].a/w1022 ), .B(
        \SUBBYTES[2].a/w1029 ), .Z(n8003) );
  XOR \SUBBYTES[2].a/U4205  ( .A(n8342), .B(n8343), .Z(\SUBBYTES[2].a/w1049 )
         );
  XOR \SUBBYTES[2].a/U4204  ( .A(\w1[2][91] ), .B(n8004), .Z(n8346) );
  XOR \SUBBYTES[2].a/U4203  ( .A(\SUBBYTES[2].a/w1011 ), .B(
        \SUBBYTES[2].a/w1014 ), .Z(n8004) );
  XOR \SUBBYTES[2].a/U4202  ( .A(n8006), .B(n8005), .Z(\SUBBYTES[2].a/w1038 )
         );
  XOR \SUBBYTES[2].a/U4201  ( .A(n8346), .B(n8007), .Z(n8005) );
  XOR \SUBBYTES[2].a/U4200  ( .A(\w1[2][94] ), .B(\SUBBYTES[2].a/w1080 ), .Z(
        n8006) );
  XOR \SUBBYTES[2].a/U4199  ( .A(\SUBBYTES[2].a/w1019 ), .B(
        \SUBBYTES[2].a/w1020 ), .Z(n8007) );
  XOR \SUBBYTES[2].a/U4198  ( .A(n8344), .B(n8343), .Z(\SUBBYTES[2].a/w1058 )
         );
  XOR \SUBBYTES[2].a/U4197  ( .A(n8009), .B(n8008), .Z(\SUBBYTES[2].a/w1059 )
         );
  XOR \SUBBYTES[2].a/U4196  ( .A(\w1[2][95] ), .B(n8345), .Z(n8008) );
  XOR \SUBBYTES[2].a/U4195  ( .A(\SUBBYTES[2].a/w1011 ), .B(
        \SUBBYTES[2].a/w1020 ), .Z(n8009) );
  XOR \SUBBYTES[2].a/U4194  ( .A(n8011), .B(n8010), .Z(\SUBBYTES[2].a/w1035 )
         );
  XOR \SUBBYTES[2].a/U4193  ( .A(n8013), .B(n8012), .Z(n8010) );
  XOR \SUBBYTES[2].a/U4192  ( .A(\w1[2][95] ), .B(\SUBBYTES[2].a/w1119 ), .Z(
        n8011) );
  XOR \SUBBYTES[2].a/U4191  ( .A(\SUBBYTES[2].a/w1026 ), .B(
        \SUBBYTES[2].a/w1029 ), .Z(n8012) );
  XOR \SUBBYTES[2].a/U4190  ( .A(\SUBBYTES[2].a/w1012 ), .B(
        \SUBBYTES[2].a/w1014 ), .Z(n8013) );
  XOR \SUBBYTES[2].a/U4189  ( .A(n8015), .B(n8014), .Z(\SUBBYTES[2].a/w1036 )
         );
  XOR \SUBBYTES[2].a/U4188  ( .A(n8346), .B(n8016), .Z(n8014) );
  XOR \SUBBYTES[2].a/U4187  ( .A(\w1[2][93] ), .B(n8347), .Z(n8015) );
  XOR \SUBBYTES[2].a/U4186  ( .A(\SUBBYTES[2].a/w1026 ), .B(
        \SUBBYTES[2].a/w1027 ), .Z(n8016) );
  XOR \SUBBYTES[2].a/U4185  ( .A(n8018), .B(n8017), .Z(\SUBBYTES[2].a/w1052 )
         );
  XOR \SUBBYTES[2].a/U4184  ( .A(\w1[2][89] ), .B(n8019), .Z(n8017) );
  XOR \SUBBYTES[2].a/U4183  ( .A(\SUBBYTES[2].a/w1027 ), .B(
        \SUBBYTES[2].a/w1029 ), .Z(n8018) );
  XOR \SUBBYTES[2].a/U4182  ( .A(\SUBBYTES[2].a/w1011 ), .B(
        \SUBBYTES[2].a/w1012 ), .Z(n8019) );
  XOR \SUBBYTES[2].a/U4181  ( .A(\w1[2][97] ), .B(n8020), .Z(n8348) );
  XOR \SUBBYTES[2].a/U4180  ( .A(\w1[2][99] ), .B(\w1[2][98] ), .Z(n8020) );
  XOR \SUBBYTES[2].a/U4179  ( .A(\w1[2][102] ), .B(n8348), .Z(
        \SUBBYTES[2].a/w894 ) );
  XOR \SUBBYTES[2].a/U4178  ( .A(\w1[2][96] ), .B(\SUBBYTES[2].a/w894 ), .Z(
        \SUBBYTES[2].a/w781 ) );
  XOR \SUBBYTES[2].a/U4177  ( .A(\w1[2][96] ), .B(n8021), .Z(
        \SUBBYTES[2].a/w782 ) );
  XOR \SUBBYTES[2].a/U4176  ( .A(\w1[2][102] ), .B(\w1[2][101] ), .Z(n8021) );
  XOR \SUBBYTES[2].a/U4175  ( .A(\w1[2][101] ), .B(n8348), .Z(
        \SUBBYTES[2].a/w912 ) );
  XOR \SUBBYTES[2].a/U4174  ( .A(n8023), .B(n8022), .Z(\SUBBYTES[2].a/w905 )
         );
  XOR \SUBBYTES[2].a/U4173  ( .A(\w1[2][99] ), .B(\w1[2][97] ), .Z(n8022) );
  XOR \SUBBYTES[2].a/U4172  ( .A(\w1[2][103] ), .B(\w1[2][100] ), .Z(n8023) );
  XOR \SUBBYTES[2].a/U4171  ( .A(\w1[2][96] ), .B(\SUBBYTES[2].a/w905 ), .Z(
        \SUBBYTES[2].a/w784 ) );
  XOR \SUBBYTES[2].a/U4170  ( .A(n8025), .B(n8024), .Z(\SUBBYTES[2].a/w892 )
         );
  XOR \SUBBYTES[2].a/U4169  ( .A(\SUBBYTES[2].a/w853 ), .B(n976), .Z(n8024) );
  XOR \SUBBYTES[2].a/U4168  ( .A(\SUBBYTES[2].a/w846 ), .B(
        \SUBBYTES[2].a/w849 ), .Z(n8025) );
  XOR \SUBBYTES[2].a/U4167  ( .A(n8027), .B(n8026), .Z(\SUBBYTES[2].a/w893 )
         );
  XOR \SUBBYTES[2].a/U4166  ( .A(\SUBBYTES[2].a/w853 ), .B(n7119), .Z(n8026)
         );
  XOR \SUBBYTES[2].a/U4165  ( .A(\SUBBYTES[2].a/w846 ), .B(n7118), .Z(n8027)
         );
  XOR \SUBBYTES[2].a/U4164  ( .A(\SUBBYTES[2].a/w905 ), .B(n8028), .Z(
        \SUBBYTES[2].a/w895 ) );
  XOR \SUBBYTES[2].a/U4163  ( .A(\w1[2][102] ), .B(\w1[2][101] ), .Z(n8028) );
  XOR \SUBBYTES[2].a/U4162  ( .A(n8030), .B(n8029), .Z(\SUBBYTES[2].a/w896 )
         );
  XOR \SUBBYTES[2].a/U4161  ( .A(n7119), .B(n976), .Z(n8029) );
  XOR \SUBBYTES[2].a/U4160  ( .A(n7118), .B(\SUBBYTES[2].a/w849 ), .Z(n8030)
         );
  XOR \SUBBYTES[2].a/U4159  ( .A(\w1[2][103] ), .B(\w1[2][98] ), .Z(n8354) );
  XOR \SUBBYTES[2].a/U4158  ( .A(n8354), .B(n8031), .Z(\SUBBYTES[2].a/w897 )
         );
  XOR \SUBBYTES[2].a/U4157  ( .A(\w1[2][101] ), .B(\w1[2][100] ), .Z(n8031) );
  XOR \SUBBYTES[2].a/U4156  ( .A(\w1[2][103] ), .B(\SUBBYTES[2].a/w782 ), .Z(
        \SUBBYTES[2].a/w785 ) );
  XOR \SUBBYTES[2].a/U4155  ( .A(\w1[2][97] ), .B(\SUBBYTES[2].a/w782 ), .Z(
        \SUBBYTES[2].a/w786 ) );
  XOR \SUBBYTES[2].a/U4154  ( .A(\w1[2][100] ), .B(\SUBBYTES[2].a/w782 ), .Z(
        \SUBBYTES[2].a/w787 ) );
  XOR \SUBBYTES[2].a/U4153  ( .A(\SUBBYTES[2].a/w786 ), .B(n8354), .Z(
        \SUBBYTES[2].a/w788 ) );
  XOR \SUBBYTES[2].a/U4152  ( .A(n8354), .B(n8032), .Z(\SUBBYTES[2].a/w873 )
         );
  XOR \SUBBYTES[2].a/U4151  ( .A(\w1[2][100] ), .B(\w1[2][97] ), .Z(n8032) );
  XOR \SUBBYTES[2].a/U4150  ( .A(n8034), .B(n8033), .Z(n8351) );
  XOR \SUBBYTES[2].a/U4149  ( .A(\w1[2][100] ), .B(n8035), .Z(n8033) );
  XOR \SUBBYTES[2].a/U4148  ( .A(\SUBBYTES[2].a/w838 ), .B(\w1[2][102] ), .Z(
        n8034) );
  XOR \SUBBYTES[2].a/U4147  ( .A(\SUBBYTES[2].a/w812 ), .B(
        \SUBBYTES[2].a/w819 ), .Z(n8035) );
  XOR \SUBBYTES[2].a/U4146  ( .A(n8037), .B(n8036), .Z(n8349) );
  XOR \SUBBYTES[2].a/U4145  ( .A(\w1[2][97] ), .B(n8038), .Z(n8036) );
  XOR \SUBBYTES[2].a/U4144  ( .A(\SUBBYTES[2].a/w837 ), .B(\w1[2][101] ), .Z(
        n8037) );
  XOR \SUBBYTES[2].a/U4143  ( .A(\SUBBYTES[2].a/w813 ), .B(
        \SUBBYTES[2].a/w820 ), .Z(n8038) );
  XOR \SUBBYTES[2].a/U4142  ( .A(n8351), .B(n8349), .Z(\SUBBYTES[2].a/w843 )
         );
  XOR \SUBBYTES[2].a/U4141  ( .A(\w1[2][101] ), .B(n8039), .Z(n8352) );
  XOR \SUBBYTES[2].a/U4140  ( .A(\SUBBYTES[2].a/w805 ), .B(
        \SUBBYTES[2].a/w815 ), .Z(n8039) );
  XOR \SUBBYTES[2].a/U4139  ( .A(n8041), .B(n8040), .Z(\SUBBYTES[2].a/w830 )
         );
  XOR \SUBBYTES[2].a/U4138  ( .A(n8352), .B(n8042), .Z(n8040) );
  XOR \SUBBYTES[2].a/U4137  ( .A(\w1[2][100] ), .B(\SUBBYTES[2].a/w894 ), .Z(
        n8041) );
  XOR \SUBBYTES[2].a/U4136  ( .A(\SUBBYTES[2].a/w807 ), .B(
        \SUBBYTES[2].a/w812 ), .Z(n8042) );
  XOR \SUBBYTES[2].a/U4135  ( .A(n8044), .B(n8043), .Z(n8350) );
  XOR \SUBBYTES[2].a/U4134  ( .A(\SUBBYTES[2].a/w840 ), .B(\w1[2][103] ), .Z(
        n8043) );
  XOR \SUBBYTES[2].a/U4133  ( .A(\SUBBYTES[2].a/w815 ), .B(
        \SUBBYTES[2].a/w822 ), .Z(n8044) );
  XOR \SUBBYTES[2].a/U4132  ( .A(n8349), .B(n8350), .Z(\SUBBYTES[2].a/w842 )
         );
  XOR \SUBBYTES[2].a/U4131  ( .A(\w1[2][99] ), .B(n8045), .Z(n8353) );
  XOR \SUBBYTES[2].a/U4130  ( .A(\SUBBYTES[2].a/w804 ), .B(
        \SUBBYTES[2].a/w807 ), .Z(n8045) );
  XOR \SUBBYTES[2].a/U4129  ( .A(n8047), .B(n8046), .Z(\SUBBYTES[2].a/w831 )
         );
  XOR \SUBBYTES[2].a/U4128  ( .A(n8353), .B(n8048), .Z(n8046) );
  XOR \SUBBYTES[2].a/U4127  ( .A(\w1[2][102] ), .B(\SUBBYTES[2].a/w873 ), .Z(
        n8047) );
  XOR \SUBBYTES[2].a/U4126  ( .A(\SUBBYTES[2].a/w812 ), .B(
        \SUBBYTES[2].a/w813 ), .Z(n8048) );
  XOR \SUBBYTES[2].a/U4125  ( .A(n8351), .B(n8350), .Z(\SUBBYTES[2].a/w851 )
         );
  XOR \SUBBYTES[2].a/U4124  ( .A(n8050), .B(n8049), .Z(\SUBBYTES[2].a/w852 )
         );
  XOR \SUBBYTES[2].a/U4123  ( .A(\w1[2][103] ), .B(n8352), .Z(n8049) );
  XOR \SUBBYTES[2].a/U4122  ( .A(\SUBBYTES[2].a/w804 ), .B(
        \SUBBYTES[2].a/w813 ), .Z(n8050) );
  XOR \SUBBYTES[2].a/U4121  ( .A(n8052), .B(n8051), .Z(\SUBBYTES[2].a/w828 )
         );
  XOR \SUBBYTES[2].a/U4120  ( .A(n8054), .B(n8053), .Z(n8051) );
  XOR \SUBBYTES[2].a/U4119  ( .A(\w1[2][103] ), .B(\SUBBYTES[2].a/w912 ), .Z(
        n8052) );
  XOR \SUBBYTES[2].a/U4118  ( .A(\SUBBYTES[2].a/w819 ), .B(
        \SUBBYTES[2].a/w822 ), .Z(n8053) );
  XOR \SUBBYTES[2].a/U4117  ( .A(\SUBBYTES[2].a/w805 ), .B(
        \SUBBYTES[2].a/w807 ), .Z(n8054) );
  XOR \SUBBYTES[2].a/U4116  ( .A(n8056), .B(n8055), .Z(\SUBBYTES[2].a/w829 )
         );
  XOR \SUBBYTES[2].a/U4115  ( .A(n8353), .B(n8057), .Z(n8055) );
  XOR \SUBBYTES[2].a/U4114  ( .A(\w1[2][101] ), .B(n8354), .Z(n8056) );
  XOR \SUBBYTES[2].a/U4113  ( .A(\SUBBYTES[2].a/w819 ), .B(
        \SUBBYTES[2].a/w820 ), .Z(n8057) );
  XOR \SUBBYTES[2].a/U4112  ( .A(n8059), .B(n8058), .Z(\SUBBYTES[2].a/w845 )
         );
  XOR \SUBBYTES[2].a/U4111  ( .A(\w1[2][97] ), .B(n8060), .Z(n8058) );
  XOR \SUBBYTES[2].a/U4110  ( .A(\SUBBYTES[2].a/w820 ), .B(
        \SUBBYTES[2].a/w822 ), .Z(n8059) );
  XOR \SUBBYTES[2].a/U4109  ( .A(\SUBBYTES[2].a/w804 ), .B(
        \SUBBYTES[2].a/w805 ), .Z(n8060) );
  XOR \SUBBYTES[2].a/U4108  ( .A(\w1[2][105] ), .B(n8061), .Z(n8355) );
  XOR \SUBBYTES[2].a/U4107  ( .A(\w1[2][107] ), .B(\w1[2][106] ), .Z(n8061) );
  XOR \SUBBYTES[2].a/U4106  ( .A(\w1[2][110] ), .B(n8355), .Z(
        \SUBBYTES[2].a/w687 ) );
  XOR \SUBBYTES[2].a/U4105  ( .A(\w1[2][104] ), .B(\SUBBYTES[2].a/w687 ), .Z(
        \SUBBYTES[2].a/w574 ) );
  XOR \SUBBYTES[2].a/U4104  ( .A(\w1[2][104] ), .B(n8062), .Z(
        \SUBBYTES[2].a/w575 ) );
  XOR \SUBBYTES[2].a/U4103  ( .A(\w1[2][110] ), .B(\w1[2][109] ), .Z(n8062) );
  XOR \SUBBYTES[2].a/U4102  ( .A(\w1[2][109] ), .B(n8355), .Z(
        \SUBBYTES[2].a/w705 ) );
  XOR \SUBBYTES[2].a/U4101  ( .A(n8064), .B(n8063), .Z(\SUBBYTES[2].a/w698 )
         );
  XOR \SUBBYTES[2].a/U4100  ( .A(\w1[2][107] ), .B(\w1[2][105] ), .Z(n8063) );
  XOR \SUBBYTES[2].a/U4099  ( .A(\w1[2][111] ), .B(\w1[2][108] ), .Z(n8064) );
  XOR \SUBBYTES[2].a/U4098  ( .A(\w1[2][104] ), .B(\SUBBYTES[2].a/w698 ), .Z(
        \SUBBYTES[2].a/w577 ) );
  XOR \SUBBYTES[2].a/U4097  ( .A(n8066), .B(n8065), .Z(\SUBBYTES[2].a/w685 )
         );
  XOR \SUBBYTES[2].a/U4096  ( .A(\SUBBYTES[2].a/w646 ), .B(n975), .Z(n8065) );
  XOR \SUBBYTES[2].a/U4095  ( .A(\SUBBYTES[2].a/w639 ), .B(
        \SUBBYTES[2].a/w642 ), .Z(n8066) );
  XOR \SUBBYTES[2].a/U4094  ( .A(n8068), .B(n8067), .Z(\SUBBYTES[2].a/w686 )
         );
  XOR \SUBBYTES[2].a/U4093  ( .A(\SUBBYTES[2].a/w646 ), .B(n7117), .Z(n8067)
         );
  XOR \SUBBYTES[2].a/U4092  ( .A(\SUBBYTES[2].a/w639 ), .B(n7116), .Z(n8068)
         );
  XOR \SUBBYTES[2].a/U4091  ( .A(\SUBBYTES[2].a/w698 ), .B(n8069), .Z(
        \SUBBYTES[2].a/w688 ) );
  XOR \SUBBYTES[2].a/U4090  ( .A(\w1[2][110] ), .B(\w1[2][109] ), .Z(n8069) );
  XOR \SUBBYTES[2].a/U4089  ( .A(n8071), .B(n8070), .Z(\SUBBYTES[2].a/w689 )
         );
  XOR \SUBBYTES[2].a/U4088  ( .A(n7117), .B(n975), .Z(n8070) );
  XOR \SUBBYTES[2].a/U4087  ( .A(n7116), .B(\SUBBYTES[2].a/w642 ), .Z(n8071)
         );
  XOR \SUBBYTES[2].a/U4086  ( .A(\w1[2][111] ), .B(\w1[2][106] ), .Z(n8361) );
  XOR \SUBBYTES[2].a/U4085  ( .A(n8361), .B(n8072), .Z(\SUBBYTES[2].a/w690 )
         );
  XOR \SUBBYTES[2].a/U4084  ( .A(\w1[2][109] ), .B(\w1[2][108] ), .Z(n8072) );
  XOR \SUBBYTES[2].a/U4083  ( .A(\w1[2][111] ), .B(\SUBBYTES[2].a/w575 ), .Z(
        \SUBBYTES[2].a/w578 ) );
  XOR \SUBBYTES[2].a/U4082  ( .A(\w1[2][105] ), .B(\SUBBYTES[2].a/w575 ), .Z(
        \SUBBYTES[2].a/w579 ) );
  XOR \SUBBYTES[2].a/U4081  ( .A(\w1[2][108] ), .B(\SUBBYTES[2].a/w575 ), .Z(
        \SUBBYTES[2].a/w580 ) );
  XOR \SUBBYTES[2].a/U4080  ( .A(\SUBBYTES[2].a/w579 ), .B(n8361), .Z(
        \SUBBYTES[2].a/w581 ) );
  XOR \SUBBYTES[2].a/U4079  ( .A(n8361), .B(n8073), .Z(\SUBBYTES[2].a/w666 )
         );
  XOR \SUBBYTES[2].a/U4078  ( .A(\w1[2][108] ), .B(\w1[2][105] ), .Z(n8073) );
  XOR \SUBBYTES[2].a/U4077  ( .A(n8075), .B(n8074), .Z(n8358) );
  XOR \SUBBYTES[2].a/U4076  ( .A(\w1[2][108] ), .B(n8076), .Z(n8074) );
  XOR \SUBBYTES[2].a/U4075  ( .A(\SUBBYTES[2].a/w631 ), .B(\w1[2][110] ), .Z(
        n8075) );
  XOR \SUBBYTES[2].a/U4074  ( .A(\SUBBYTES[2].a/w605 ), .B(
        \SUBBYTES[2].a/w612 ), .Z(n8076) );
  XOR \SUBBYTES[2].a/U4073  ( .A(n8078), .B(n8077), .Z(n8356) );
  XOR \SUBBYTES[2].a/U4072  ( .A(\w1[2][105] ), .B(n8079), .Z(n8077) );
  XOR \SUBBYTES[2].a/U4071  ( .A(\SUBBYTES[2].a/w630 ), .B(\w1[2][109] ), .Z(
        n8078) );
  XOR \SUBBYTES[2].a/U4070  ( .A(\SUBBYTES[2].a/w606 ), .B(
        \SUBBYTES[2].a/w613 ), .Z(n8079) );
  XOR \SUBBYTES[2].a/U4069  ( .A(n8358), .B(n8356), .Z(\SUBBYTES[2].a/w636 )
         );
  XOR \SUBBYTES[2].a/U4068  ( .A(\w1[2][109] ), .B(n8080), .Z(n8359) );
  XOR \SUBBYTES[2].a/U4067  ( .A(\SUBBYTES[2].a/w598 ), .B(
        \SUBBYTES[2].a/w608 ), .Z(n8080) );
  XOR \SUBBYTES[2].a/U4066  ( .A(n8082), .B(n8081), .Z(\SUBBYTES[2].a/w623 )
         );
  XOR \SUBBYTES[2].a/U4065  ( .A(n8359), .B(n8083), .Z(n8081) );
  XOR \SUBBYTES[2].a/U4064  ( .A(\w1[2][108] ), .B(\SUBBYTES[2].a/w687 ), .Z(
        n8082) );
  XOR \SUBBYTES[2].a/U4063  ( .A(\SUBBYTES[2].a/w600 ), .B(
        \SUBBYTES[2].a/w605 ), .Z(n8083) );
  XOR \SUBBYTES[2].a/U4062  ( .A(n8085), .B(n8084), .Z(n8357) );
  XOR \SUBBYTES[2].a/U4061  ( .A(\SUBBYTES[2].a/w633 ), .B(\w1[2][111] ), .Z(
        n8084) );
  XOR \SUBBYTES[2].a/U4060  ( .A(\SUBBYTES[2].a/w608 ), .B(
        \SUBBYTES[2].a/w615 ), .Z(n8085) );
  XOR \SUBBYTES[2].a/U4059  ( .A(n8356), .B(n8357), .Z(\SUBBYTES[2].a/w635 )
         );
  XOR \SUBBYTES[2].a/U4058  ( .A(\w1[2][107] ), .B(n8086), .Z(n8360) );
  XOR \SUBBYTES[2].a/U4057  ( .A(\SUBBYTES[2].a/w597 ), .B(
        \SUBBYTES[2].a/w600 ), .Z(n8086) );
  XOR \SUBBYTES[2].a/U4056  ( .A(n8088), .B(n8087), .Z(\SUBBYTES[2].a/w624 )
         );
  XOR \SUBBYTES[2].a/U4055  ( .A(n8360), .B(n8089), .Z(n8087) );
  XOR \SUBBYTES[2].a/U4054  ( .A(\w1[2][110] ), .B(\SUBBYTES[2].a/w666 ), .Z(
        n8088) );
  XOR \SUBBYTES[2].a/U4053  ( .A(\SUBBYTES[2].a/w605 ), .B(
        \SUBBYTES[2].a/w606 ), .Z(n8089) );
  XOR \SUBBYTES[2].a/U4052  ( .A(n8358), .B(n8357), .Z(\SUBBYTES[2].a/w644 )
         );
  XOR \SUBBYTES[2].a/U4051  ( .A(n8091), .B(n8090), .Z(\SUBBYTES[2].a/w645 )
         );
  XOR \SUBBYTES[2].a/U4050  ( .A(\w1[2][111] ), .B(n8359), .Z(n8090) );
  XOR \SUBBYTES[2].a/U4049  ( .A(\SUBBYTES[2].a/w597 ), .B(
        \SUBBYTES[2].a/w606 ), .Z(n8091) );
  XOR \SUBBYTES[2].a/U4048  ( .A(n8093), .B(n8092), .Z(\SUBBYTES[2].a/w621 )
         );
  XOR \SUBBYTES[2].a/U4047  ( .A(n8095), .B(n8094), .Z(n8092) );
  XOR \SUBBYTES[2].a/U4046  ( .A(\w1[2][111] ), .B(\SUBBYTES[2].a/w705 ), .Z(
        n8093) );
  XOR \SUBBYTES[2].a/U4045  ( .A(\SUBBYTES[2].a/w612 ), .B(
        \SUBBYTES[2].a/w615 ), .Z(n8094) );
  XOR \SUBBYTES[2].a/U4044  ( .A(\SUBBYTES[2].a/w598 ), .B(
        \SUBBYTES[2].a/w600 ), .Z(n8095) );
  XOR \SUBBYTES[2].a/U4043  ( .A(n8097), .B(n8096), .Z(\SUBBYTES[2].a/w622 )
         );
  XOR \SUBBYTES[2].a/U4042  ( .A(n8360), .B(n8098), .Z(n8096) );
  XOR \SUBBYTES[2].a/U4041  ( .A(\w1[2][109] ), .B(n8361), .Z(n8097) );
  XOR \SUBBYTES[2].a/U4040  ( .A(\SUBBYTES[2].a/w612 ), .B(
        \SUBBYTES[2].a/w613 ), .Z(n8098) );
  XOR \SUBBYTES[2].a/U4039  ( .A(n8100), .B(n8099), .Z(\SUBBYTES[2].a/w638 )
         );
  XOR \SUBBYTES[2].a/U4038  ( .A(\w1[2][105] ), .B(n8101), .Z(n8099) );
  XOR \SUBBYTES[2].a/U4037  ( .A(\SUBBYTES[2].a/w613 ), .B(
        \SUBBYTES[2].a/w615 ), .Z(n8100) );
  XOR \SUBBYTES[2].a/U4036  ( .A(\SUBBYTES[2].a/w597 ), .B(
        \SUBBYTES[2].a/w598 ), .Z(n8101) );
  XOR \SUBBYTES[2].a/U4035  ( .A(\w1[2][113] ), .B(n8102), .Z(n8362) );
  XOR \SUBBYTES[2].a/U4034  ( .A(\w1[2][115] ), .B(\w1[2][114] ), .Z(n8102) );
  XOR \SUBBYTES[2].a/U4033  ( .A(\w1[2][118] ), .B(n8362), .Z(
        \SUBBYTES[2].a/w480 ) );
  XOR \SUBBYTES[2].a/U4032  ( .A(\w1[2][112] ), .B(\SUBBYTES[2].a/w480 ), .Z(
        \SUBBYTES[2].a/w367 ) );
  XOR \SUBBYTES[2].a/U4031  ( .A(\w1[2][112] ), .B(n8103), .Z(
        \SUBBYTES[2].a/w368 ) );
  XOR \SUBBYTES[2].a/U4030  ( .A(\w1[2][118] ), .B(\w1[2][117] ), .Z(n8103) );
  XOR \SUBBYTES[2].a/U4029  ( .A(\w1[2][117] ), .B(n8362), .Z(
        \SUBBYTES[2].a/w498 ) );
  XOR \SUBBYTES[2].a/U4028  ( .A(n8105), .B(n8104), .Z(\SUBBYTES[2].a/w491 )
         );
  XOR \SUBBYTES[2].a/U4027  ( .A(\w1[2][115] ), .B(\w1[2][113] ), .Z(n8104) );
  XOR \SUBBYTES[2].a/U4026  ( .A(\w1[2][119] ), .B(\w1[2][116] ), .Z(n8105) );
  XOR \SUBBYTES[2].a/U4025  ( .A(\w1[2][112] ), .B(\SUBBYTES[2].a/w491 ), .Z(
        \SUBBYTES[2].a/w370 ) );
  XOR \SUBBYTES[2].a/U4024  ( .A(n8107), .B(n8106), .Z(\SUBBYTES[2].a/w478 )
         );
  XOR \SUBBYTES[2].a/U4023  ( .A(\SUBBYTES[2].a/w439 ), .B(n974), .Z(n8106) );
  XOR \SUBBYTES[2].a/U4022  ( .A(\SUBBYTES[2].a/w432 ), .B(
        \SUBBYTES[2].a/w435 ), .Z(n8107) );
  XOR \SUBBYTES[2].a/U4021  ( .A(n8109), .B(n8108), .Z(\SUBBYTES[2].a/w479 )
         );
  XOR \SUBBYTES[2].a/U4020  ( .A(\SUBBYTES[2].a/w439 ), .B(n7115), .Z(n8108)
         );
  XOR \SUBBYTES[2].a/U4019  ( .A(\SUBBYTES[2].a/w432 ), .B(n7114), .Z(n8109)
         );
  XOR \SUBBYTES[2].a/U4018  ( .A(\SUBBYTES[2].a/w491 ), .B(n8110), .Z(
        \SUBBYTES[2].a/w481 ) );
  XOR \SUBBYTES[2].a/U4017  ( .A(\w1[2][118] ), .B(\w1[2][117] ), .Z(n8110) );
  XOR \SUBBYTES[2].a/U4016  ( .A(n8112), .B(n8111), .Z(\SUBBYTES[2].a/w482 )
         );
  XOR \SUBBYTES[2].a/U4015  ( .A(n7115), .B(n974), .Z(n8111) );
  XOR \SUBBYTES[2].a/U4014  ( .A(n7114), .B(\SUBBYTES[2].a/w435 ), .Z(n8112)
         );
  XOR \SUBBYTES[2].a/U4013  ( .A(\w1[2][119] ), .B(\w1[2][114] ), .Z(n8368) );
  XOR \SUBBYTES[2].a/U4012  ( .A(n8368), .B(n8113), .Z(\SUBBYTES[2].a/w483 )
         );
  XOR \SUBBYTES[2].a/U4011  ( .A(\w1[2][117] ), .B(\w1[2][116] ), .Z(n8113) );
  XOR \SUBBYTES[2].a/U4010  ( .A(\w1[2][119] ), .B(\SUBBYTES[2].a/w368 ), .Z(
        \SUBBYTES[2].a/w371 ) );
  XOR \SUBBYTES[2].a/U4009  ( .A(\w1[2][113] ), .B(\SUBBYTES[2].a/w368 ), .Z(
        \SUBBYTES[2].a/w372 ) );
  XOR \SUBBYTES[2].a/U4008  ( .A(\w1[2][116] ), .B(\SUBBYTES[2].a/w368 ), .Z(
        \SUBBYTES[2].a/w373 ) );
  XOR \SUBBYTES[2].a/U4007  ( .A(\SUBBYTES[2].a/w372 ), .B(n8368), .Z(
        \SUBBYTES[2].a/w374 ) );
  XOR \SUBBYTES[2].a/U4006  ( .A(n8368), .B(n8114), .Z(\SUBBYTES[2].a/w459 )
         );
  XOR \SUBBYTES[2].a/U4005  ( .A(\w1[2][116] ), .B(\w1[2][113] ), .Z(n8114) );
  XOR \SUBBYTES[2].a/U4004  ( .A(n8116), .B(n8115), .Z(n8365) );
  XOR \SUBBYTES[2].a/U4003  ( .A(\w1[2][116] ), .B(n8117), .Z(n8115) );
  XOR \SUBBYTES[2].a/U4002  ( .A(\SUBBYTES[2].a/w424 ), .B(\w1[2][118] ), .Z(
        n8116) );
  XOR \SUBBYTES[2].a/U4001  ( .A(\SUBBYTES[2].a/w398 ), .B(
        \SUBBYTES[2].a/w405 ), .Z(n8117) );
  XOR \SUBBYTES[2].a/U4000  ( .A(n8119), .B(n8118), .Z(n8363) );
  XOR \SUBBYTES[2].a/U3999  ( .A(\w1[2][113] ), .B(n8120), .Z(n8118) );
  XOR \SUBBYTES[2].a/U3998  ( .A(\SUBBYTES[2].a/w423 ), .B(\w1[2][117] ), .Z(
        n8119) );
  XOR \SUBBYTES[2].a/U3997  ( .A(\SUBBYTES[2].a/w399 ), .B(
        \SUBBYTES[2].a/w406 ), .Z(n8120) );
  XOR \SUBBYTES[2].a/U3996  ( .A(n8365), .B(n8363), .Z(\SUBBYTES[2].a/w429 )
         );
  XOR \SUBBYTES[2].a/U3995  ( .A(\w1[2][117] ), .B(n8121), .Z(n8366) );
  XOR \SUBBYTES[2].a/U3994  ( .A(\SUBBYTES[2].a/w391 ), .B(
        \SUBBYTES[2].a/w401 ), .Z(n8121) );
  XOR \SUBBYTES[2].a/U3993  ( .A(n8123), .B(n8122), .Z(\SUBBYTES[2].a/w416 )
         );
  XOR \SUBBYTES[2].a/U3992  ( .A(n8366), .B(n8124), .Z(n8122) );
  XOR \SUBBYTES[2].a/U3991  ( .A(\w1[2][116] ), .B(\SUBBYTES[2].a/w480 ), .Z(
        n8123) );
  XOR \SUBBYTES[2].a/U3990  ( .A(\SUBBYTES[2].a/w393 ), .B(
        \SUBBYTES[2].a/w398 ), .Z(n8124) );
  XOR \SUBBYTES[2].a/U3989  ( .A(n8126), .B(n8125), .Z(n8364) );
  XOR \SUBBYTES[2].a/U3988  ( .A(\SUBBYTES[2].a/w426 ), .B(\w1[2][119] ), .Z(
        n8125) );
  XOR \SUBBYTES[2].a/U3987  ( .A(\SUBBYTES[2].a/w401 ), .B(
        \SUBBYTES[2].a/w408 ), .Z(n8126) );
  XOR \SUBBYTES[2].a/U3986  ( .A(n8363), .B(n8364), .Z(\SUBBYTES[2].a/w428 )
         );
  XOR \SUBBYTES[2].a/U3985  ( .A(\w1[2][115] ), .B(n8127), .Z(n8367) );
  XOR \SUBBYTES[2].a/U3984  ( .A(\SUBBYTES[2].a/w390 ), .B(
        \SUBBYTES[2].a/w393 ), .Z(n8127) );
  XOR \SUBBYTES[2].a/U3983  ( .A(n8129), .B(n8128), .Z(\SUBBYTES[2].a/w417 )
         );
  XOR \SUBBYTES[2].a/U3982  ( .A(n8367), .B(n8130), .Z(n8128) );
  XOR \SUBBYTES[2].a/U3981  ( .A(\w1[2][118] ), .B(\SUBBYTES[2].a/w459 ), .Z(
        n8129) );
  XOR \SUBBYTES[2].a/U3980  ( .A(\SUBBYTES[2].a/w398 ), .B(
        \SUBBYTES[2].a/w399 ), .Z(n8130) );
  XOR \SUBBYTES[2].a/U3979  ( .A(n8365), .B(n8364), .Z(\SUBBYTES[2].a/w437 )
         );
  XOR \SUBBYTES[2].a/U3978  ( .A(n8132), .B(n8131), .Z(\SUBBYTES[2].a/w438 )
         );
  XOR \SUBBYTES[2].a/U3977  ( .A(\w1[2][119] ), .B(n8366), .Z(n8131) );
  XOR \SUBBYTES[2].a/U3976  ( .A(\SUBBYTES[2].a/w390 ), .B(
        \SUBBYTES[2].a/w399 ), .Z(n8132) );
  XOR \SUBBYTES[2].a/U3975  ( .A(n8134), .B(n8133), .Z(\SUBBYTES[2].a/w414 )
         );
  XOR \SUBBYTES[2].a/U3974  ( .A(n8136), .B(n8135), .Z(n8133) );
  XOR \SUBBYTES[2].a/U3973  ( .A(\w1[2][119] ), .B(\SUBBYTES[2].a/w498 ), .Z(
        n8134) );
  XOR \SUBBYTES[2].a/U3972  ( .A(\SUBBYTES[2].a/w405 ), .B(
        \SUBBYTES[2].a/w408 ), .Z(n8135) );
  XOR \SUBBYTES[2].a/U3971  ( .A(\SUBBYTES[2].a/w391 ), .B(
        \SUBBYTES[2].a/w393 ), .Z(n8136) );
  XOR \SUBBYTES[2].a/U3970  ( .A(n8138), .B(n8137), .Z(\SUBBYTES[2].a/w415 )
         );
  XOR \SUBBYTES[2].a/U3969  ( .A(n8367), .B(n8139), .Z(n8137) );
  XOR \SUBBYTES[2].a/U3968  ( .A(\w1[2][117] ), .B(n8368), .Z(n8138) );
  XOR \SUBBYTES[2].a/U3967  ( .A(\SUBBYTES[2].a/w405 ), .B(
        \SUBBYTES[2].a/w406 ), .Z(n8139) );
  XOR \SUBBYTES[2].a/U3966  ( .A(n8141), .B(n8140), .Z(\SUBBYTES[2].a/w431 )
         );
  XOR \SUBBYTES[2].a/U3965  ( .A(\w1[2][113] ), .B(n8142), .Z(n8140) );
  XOR \SUBBYTES[2].a/U3964  ( .A(\SUBBYTES[2].a/w406 ), .B(
        \SUBBYTES[2].a/w408 ), .Z(n8141) );
  XOR \SUBBYTES[2].a/U3963  ( .A(\SUBBYTES[2].a/w390 ), .B(
        \SUBBYTES[2].a/w391 ), .Z(n8142) );
  XOR \SUBBYTES[2].a/U3962  ( .A(\w1[2][121] ), .B(n8143), .Z(n8369) );
  XOR \SUBBYTES[2].a/U3961  ( .A(\w1[2][123] ), .B(\w1[2][122] ), .Z(n8143) );
  XOR \SUBBYTES[2].a/U3960  ( .A(\w1[2][126] ), .B(n8369), .Z(
        \SUBBYTES[2].a/w273 ) );
  XOR \SUBBYTES[2].a/U3959  ( .A(\w1[2][120] ), .B(\SUBBYTES[2].a/w273 ), .Z(
        \SUBBYTES[2].a/w160 ) );
  XOR \SUBBYTES[2].a/U3958  ( .A(\w1[2][120] ), .B(n8144), .Z(
        \SUBBYTES[2].a/w161 ) );
  XOR \SUBBYTES[2].a/U3957  ( .A(\w1[2][126] ), .B(\w1[2][125] ), .Z(n8144) );
  XOR \SUBBYTES[2].a/U3956  ( .A(\w1[2][125] ), .B(n8369), .Z(
        \SUBBYTES[2].a/w291 ) );
  XOR \SUBBYTES[2].a/U3955  ( .A(n8146), .B(n8145), .Z(\SUBBYTES[2].a/w284 )
         );
  XOR \SUBBYTES[2].a/U3954  ( .A(\w1[2][123] ), .B(\w1[2][121] ), .Z(n8145) );
  XOR \SUBBYTES[2].a/U3953  ( .A(\w1[2][127] ), .B(\w1[2][124] ), .Z(n8146) );
  XOR \SUBBYTES[2].a/U3952  ( .A(\w1[2][120] ), .B(\SUBBYTES[2].a/w284 ), .Z(
        \SUBBYTES[2].a/w163 ) );
  XOR \SUBBYTES[2].a/U3951  ( .A(n8148), .B(n8147), .Z(\SUBBYTES[2].a/w271 )
         );
  XOR \SUBBYTES[2].a/U3950  ( .A(\SUBBYTES[2].a/w232 ), .B(n973), .Z(n8147) );
  XOR \SUBBYTES[2].a/U3949  ( .A(\SUBBYTES[2].a/w225 ), .B(
        \SUBBYTES[2].a/w228 ), .Z(n8148) );
  XOR \SUBBYTES[2].a/U3948  ( .A(n8150), .B(n8149), .Z(\SUBBYTES[2].a/w272 )
         );
  XOR \SUBBYTES[2].a/U3947  ( .A(\SUBBYTES[2].a/w232 ), .B(n7113), .Z(n8149)
         );
  XOR \SUBBYTES[2].a/U3946  ( .A(\SUBBYTES[2].a/w225 ), .B(n7112), .Z(n8150)
         );
  XOR \SUBBYTES[2].a/U3945  ( .A(\SUBBYTES[2].a/w284 ), .B(n8151), .Z(
        \SUBBYTES[2].a/w274 ) );
  XOR \SUBBYTES[2].a/U3944  ( .A(\w1[2][126] ), .B(\w1[2][125] ), .Z(n8151) );
  XOR \SUBBYTES[2].a/U3943  ( .A(n8153), .B(n8152), .Z(\SUBBYTES[2].a/w275 )
         );
  XOR \SUBBYTES[2].a/U3942  ( .A(n7113), .B(n973), .Z(n8152) );
  XOR \SUBBYTES[2].a/U3941  ( .A(n7112), .B(\SUBBYTES[2].a/w228 ), .Z(n8153)
         );
  XOR \SUBBYTES[2].a/U3940  ( .A(\w1[2][127] ), .B(\w1[2][122] ), .Z(n8375) );
  XOR \SUBBYTES[2].a/U3939  ( .A(n8375), .B(n8154), .Z(\SUBBYTES[2].a/w276 )
         );
  XOR \SUBBYTES[2].a/U3938  ( .A(\w1[2][125] ), .B(\w1[2][124] ), .Z(n8154) );
  XOR \SUBBYTES[2].a/U3937  ( .A(\w1[2][127] ), .B(\SUBBYTES[2].a/w161 ), .Z(
        \SUBBYTES[2].a/w164 ) );
  XOR \SUBBYTES[2].a/U3936  ( .A(\w1[2][121] ), .B(\SUBBYTES[2].a/w161 ), .Z(
        \SUBBYTES[2].a/w165 ) );
  XOR \SUBBYTES[2].a/U3935  ( .A(\w1[2][124] ), .B(\SUBBYTES[2].a/w161 ), .Z(
        \SUBBYTES[2].a/w166 ) );
  XOR \SUBBYTES[2].a/U3934  ( .A(\SUBBYTES[2].a/w165 ), .B(n8375), .Z(
        \SUBBYTES[2].a/w167 ) );
  XOR \SUBBYTES[2].a/U3933  ( .A(n8375), .B(n8155), .Z(\SUBBYTES[2].a/w252 )
         );
  XOR \SUBBYTES[2].a/U3932  ( .A(\w1[2][124] ), .B(\w1[2][121] ), .Z(n8155) );
  XOR \SUBBYTES[2].a/U3931  ( .A(n8157), .B(n8156), .Z(n8372) );
  XOR \SUBBYTES[2].a/U3930  ( .A(\w1[2][124] ), .B(n8158), .Z(n8156) );
  XOR \SUBBYTES[2].a/U3929  ( .A(\SUBBYTES[2].a/w217 ), .B(\w1[2][126] ), .Z(
        n8157) );
  XOR \SUBBYTES[2].a/U3928  ( .A(\SUBBYTES[2].a/w191 ), .B(
        \SUBBYTES[2].a/w198 ), .Z(n8158) );
  XOR \SUBBYTES[2].a/U3927  ( .A(n8160), .B(n8159), .Z(n8370) );
  XOR \SUBBYTES[2].a/U3926  ( .A(\w1[2][121] ), .B(n8161), .Z(n8159) );
  XOR \SUBBYTES[2].a/U3925  ( .A(\SUBBYTES[2].a/w216 ), .B(\w1[2][125] ), .Z(
        n8160) );
  XOR \SUBBYTES[2].a/U3924  ( .A(\SUBBYTES[2].a/w192 ), .B(
        \SUBBYTES[2].a/w199 ), .Z(n8161) );
  XOR \SUBBYTES[2].a/U3923  ( .A(n8372), .B(n8370), .Z(\SUBBYTES[2].a/w222 )
         );
  XOR \SUBBYTES[2].a/U3922  ( .A(\w1[2][125] ), .B(n8162), .Z(n8373) );
  XOR \SUBBYTES[2].a/U3921  ( .A(\SUBBYTES[2].a/w184 ), .B(
        \SUBBYTES[2].a/w194 ), .Z(n8162) );
  XOR \SUBBYTES[2].a/U3920  ( .A(n8164), .B(n8163), .Z(\SUBBYTES[2].a/w209 )
         );
  XOR \SUBBYTES[2].a/U3919  ( .A(n8373), .B(n8165), .Z(n8163) );
  XOR \SUBBYTES[2].a/U3918  ( .A(\w1[2][124] ), .B(\SUBBYTES[2].a/w273 ), .Z(
        n8164) );
  XOR \SUBBYTES[2].a/U3917  ( .A(\SUBBYTES[2].a/w186 ), .B(
        \SUBBYTES[2].a/w191 ), .Z(n8165) );
  XOR \SUBBYTES[2].a/U3916  ( .A(n8167), .B(n8166), .Z(n8371) );
  XOR \SUBBYTES[2].a/U3915  ( .A(\SUBBYTES[2].a/w219 ), .B(\w1[2][127] ), .Z(
        n8166) );
  XOR \SUBBYTES[2].a/U3914  ( .A(\SUBBYTES[2].a/w194 ), .B(
        \SUBBYTES[2].a/w201 ), .Z(n8167) );
  XOR \SUBBYTES[2].a/U3913  ( .A(n8370), .B(n8371), .Z(\SUBBYTES[2].a/w221 )
         );
  XOR \SUBBYTES[2].a/U3912  ( .A(\w1[2][123] ), .B(n8168), .Z(n8374) );
  XOR \SUBBYTES[2].a/U3911  ( .A(\SUBBYTES[2].a/w183 ), .B(
        \SUBBYTES[2].a/w186 ), .Z(n8168) );
  XOR \SUBBYTES[2].a/U3910  ( .A(n8170), .B(n8169), .Z(\SUBBYTES[2].a/w210 )
         );
  XOR \SUBBYTES[2].a/U3909  ( .A(n8374), .B(n8171), .Z(n8169) );
  XOR \SUBBYTES[2].a/U3908  ( .A(\w1[2][126] ), .B(\SUBBYTES[2].a/w252 ), .Z(
        n8170) );
  XOR \SUBBYTES[2].a/U3907  ( .A(\SUBBYTES[2].a/w191 ), .B(
        \SUBBYTES[2].a/w192 ), .Z(n8171) );
  XOR \SUBBYTES[2].a/U3906  ( .A(n8372), .B(n8371), .Z(\SUBBYTES[2].a/w230 )
         );
  XOR \SUBBYTES[2].a/U3905  ( .A(n8173), .B(n8172), .Z(\SUBBYTES[2].a/w231 )
         );
  XOR \SUBBYTES[2].a/U3904  ( .A(\w1[2][127] ), .B(n8373), .Z(n8172) );
  XOR \SUBBYTES[2].a/U3903  ( .A(\SUBBYTES[2].a/w183 ), .B(
        \SUBBYTES[2].a/w192 ), .Z(n8173) );
  XOR \SUBBYTES[2].a/U3902  ( .A(n8175), .B(n8174), .Z(\SUBBYTES[2].a/w207 )
         );
  XOR \SUBBYTES[2].a/U3901  ( .A(n8177), .B(n8176), .Z(n8174) );
  XOR \SUBBYTES[2].a/U3900  ( .A(\w1[2][127] ), .B(\SUBBYTES[2].a/w291 ), .Z(
        n8175) );
  XOR \SUBBYTES[2].a/U3899  ( .A(\SUBBYTES[2].a/w198 ), .B(
        \SUBBYTES[2].a/w201 ), .Z(n8176) );
  XOR \SUBBYTES[2].a/U3898  ( .A(\SUBBYTES[2].a/w184 ), .B(
        \SUBBYTES[2].a/w186 ), .Z(n8177) );
  XOR \SUBBYTES[2].a/U3897  ( .A(n8179), .B(n8178), .Z(\SUBBYTES[2].a/w208 )
         );
  XOR \SUBBYTES[2].a/U3896  ( .A(n8374), .B(n8180), .Z(n8178) );
  XOR \SUBBYTES[2].a/U3895  ( .A(\w1[2][125] ), .B(n8375), .Z(n8179) );
  XOR \SUBBYTES[2].a/U3894  ( .A(\SUBBYTES[2].a/w198 ), .B(
        \SUBBYTES[2].a/w199 ), .Z(n8180) );
  XOR \SUBBYTES[2].a/U3893  ( .A(n8182), .B(n8181), .Z(\SUBBYTES[2].a/w224 )
         );
  XOR \SUBBYTES[2].a/U3892  ( .A(\w1[2][121] ), .B(n8183), .Z(n8181) );
  XOR \SUBBYTES[2].a/U3891  ( .A(\SUBBYTES[2].a/w199 ), .B(
        \SUBBYTES[2].a/w201 ), .Z(n8182) );
  XOR \SUBBYTES[2].a/U3890  ( .A(\SUBBYTES[2].a/w183 ), .B(
        \SUBBYTES[2].a/w184 ), .Z(n8183) );
  XOR \SUBBYTES[1].a/U5649  ( .A(\SUBBYTES[1].a/w3390 ), .B(
        \SUBBYTES[1].a/w3391 ), .Z(n6905) );
  XOR \SUBBYTES[1].a/U5648  ( .A(n6905), .B(n5864), .Z(n6904) );
  XOR \SUBBYTES[1].a/U5647  ( .A(\SUBBYTES[1].a/w3383 ), .B(
        \SUBBYTES[1].a/w3400 ), .Z(n5864) );
  XOR \SUBBYTES[1].a/U5645  ( .A(\SUBBYTES[1].a/w3382 ), .B(
        \SUBBYTES[1].a/w3397 ), .Z(n5865) );
  XOR \SUBBYTES[1].a/U5644  ( .A(n6905), .B(n5866), .Z(n7096) );
  XOR \SUBBYTES[1].a/U5643  ( .A(\SUBBYTES[1].a/w3397 ), .B(
        \SUBBYTES[1].a/w3398 ), .Z(n5866) );
  XOR \SUBBYTES[1].a/U5642  ( .A(\SUBBYTES[1].a/w3359 ), .B(n5867), .Z(n6907)
         );
  XOR \SUBBYTES[1].a/U5641  ( .A(\SUBBYTES[1].a/w3350 ), .B(
        \SUBBYTES[1].a/w3351 ), .Z(n5867) );
  XOR \SUBBYTES[1].a/U5639  ( .A(\SUBBYTES[1].a/w3361 ), .B(n7096), .Z(n5868)
         );
  XOR \SUBBYTES[1].a/U5638  ( .A(n5870), .B(n5869), .Z(n6908) );
  XOR \SUBBYTES[1].a/U5637  ( .A(n5872), .B(n5871), .Z(n5869) );
  XOR \SUBBYTES[1].a/U5636  ( .A(\SUBBYTES[1].a/w3397 ), .B(
        \SUBBYTES[1].a/w3398 ), .Z(n5870) );
  XOR \SUBBYTES[1].a/U5635  ( .A(\SUBBYTES[1].a/w3361 ), .B(
        \SUBBYTES[1].a/w3385 ), .Z(n5871) );
  XOR \SUBBYTES[1].a/U5634  ( .A(\SUBBYTES[1].a/w3350 ), .B(
        \SUBBYTES[1].a/w3359 ), .Z(n5872) );
  XOR \SUBBYTES[1].a/U5633  ( .A(\SUBBYTES[1].a/w3382 ), .B(n5873), .Z(n6906)
         );
  XOR \SUBBYTES[1].a/U5632  ( .A(\SUBBYTES[1].a/w3365 ), .B(
        \SUBBYTES[1].a/w3368 ), .Z(n5873) );
  XOR \SUBBYTES[1].a/U5630  ( .A(\SUBBYTES[1].a/w3353 ), .B(n6908), .Z(n5874)
         );
  XOR \SUBBYTES[1].a/U5628  ( .A(\SUBBYTES[1].a/w3385 ), .B(
        \SUBBYTES[1].a/w3398 ), .Z(n5875) );
  XOR \SUBBYTES[1].a/U5626  ( .A(n5879), .B(n5878), .Z(n5876) );
  XOR \SUBBYTES[1].a/U5625  ( .A(n5881), .B(n5880), .Z(n5877) );
  XOR \SUBBYTES[1].a/U5624  ( .A(\SUBBYTES[1].a/w3397 ), .B(
        \SUBBYTES[1].a/w3400 ), .Z(n5878) );
  XOR \SUBBYTES[1].a/U5623  ( .A(\SUBBYTES[1].a/w3390 ), .B(
        \SUBBYTES[1].a/w3393 ), .Z(n5879) );
  XOR \SUBBYTES[1].a/U5622  ( .A(\SUBBYTES[1].a/w3365 ), .B(
        \SUBBYTES[1].a/w3366 ), .Z(n5880) );
  XOR \SUBBYTES[1].a/U5621  ( .A(\SUBBYTES[1].a/w3350 ), .B(
        \SUBBYTES[1].a/w3353 ), .Z(n5881) );
  XOR \SUBBYTES[1].a/U5619  ( .A(n6905), .B(n5884), .Z(n5882) );
  XOR \SUBBYTES[1].a/U5618  ( .A(n6907), .B(n6906), .Z(n5883) );
  XOR \SUBBYTES[1].a/U5617  ( .A(\SUBBYTES[1].a/w3358 ), .B(
        \SUBBYTES[1].a/w3385 ), .Z(n5884) );
  XOR \SUBBYTES[1].a/U5615  ( .A(n6908), .B(n5887), .Z(n5885) );
  XOR \SUBBYTES[1].a/U5614  ( .A(\SUBBYTES[1].a/w3391 ), .B(
        \SUBBYTES[1].a/w3393 ), .Z(n5886) );
  XOR \SUBBYTES[1].a/U5613  ( .A(\SUBBYTES[1].a/w3351 ), .B(
        \SUBBYTES[1].a/w3383 ), .Z(n5887) );
  XOR \SUBBYTES[1].a/U5612  ( .A(\SUBBYTES[1].a/w3183 ), .B(
        \SUBBYTES[1].a/w3184 ), .Z(n6910) );
  XOR \SUBBYTES[1].a/U5611  ( .A(n6910), .B(n5888), .Z(n6909) );
  XOR \SUBBYTES[1].a/U5610  ( .A(\SUBBYTES[1].a/w3176 ), .B(
        \SUBBYTES[1].a/w3193 ), .Z(n5888) );
  XOR \SUBBYTES[1].a/U5608  ( .A(\SUBBYTES[1].a/w3175 ), .B(
        \SUBBYTES[1].a/w3190 ), .Z(n5889) );
  XOR \SUBBYTES[1].a/U5607  ( .A(n6910), .B(n5890), .Z(n7097) );
  XOR \SUBBYTES[1].a/U5606  ( .A(\SUBBYTES[1].a/w3190 ), .B(
        \SUBBYTES[1].a/w3191 ), .Z(n5890) );
  XOR \SUBBYTES[1].a/U5605  ( .A(\SUBBYTES[1].a/w3152 ), .B(n5891), .Z(n6912)
         );
  XOR \SUBBYTES[1].a/U5604  ( .A(\SUBBYTES[1].a/w3143 ), .B(
        \SUBBYTES[1].a/w3144 ), .Z(n5891) );
  XOR \SUBBYTES[1].a/U5602  ( .A(\SUBBYTES[1].a/w3154 ), .B(n7097), .Z(n5892)
         );
  XOR \SUBBYTES[1].a/U5601  ( .A(n5894), .B(n5893), .Z(n6913) );
  XOR \SUBBYTES[1].a/U5600  ( .A(n5896), .B(n5895), .Z(n5893) );
  XOR \SUBBYTES[1].a/U5599  ( .A(\SUBBYTES[1].a/w3190 ), .B(
        \SUBBYTES[1].a/w3191 ), .Z(n5894) );
  XOR \SUBBYTES[1].a/U5598  ( .A(\SUBBYTES[1].a/w3154 ), .B(
        \SUBBYTES[1].a/w3178 ), .Z(n5895) );
  XOR \SUBBYTES[1].a/U5597  ( .A(\SUBBYTES[1].a/w3143 ), .B(
        \SUBBYTES[1].a/w3152 ), .Z(n5896) );
  XOR \SUBBYTES[1].a/U5596  ( .A(\SUBBYTES[1].a/w3175 ), .B(n5897), .Z(n6911)
         );
  XOR \SUBBYTES[1].a/U5595  ( .A(\SUBBYTES[1].a/w3158 ), .B(
        \SUBBYTES[1].a/w3161 ), .Z(n5897) );
  XOR \SUBBYTES[1].a/U5593  ( .A(\SUBBYTES[1].a/w3146 ), .B(n6913), .Z(n5898)
         );
  XOR \SUBBYTES[1].a/U5591  ( .A(\SUBBYTES[1].a/w3178 ), .B(
        \SUBBYTES[1].a/w3191 ), .Z(n5899) );
  XOR \SUBBYTES[1].a/U5589  ( .A(n5903), .B(n5902), .Z(n5900) );
  XOR \SUBBYTES[1].a/U5588  ( .A(n5905), .B(n5904), .Z(n5901) );
  XOR \SUBBYTES[1].a/U5587  ( .A(\SUBBYTES[1].a/w3190 ), .B(
        \SUBBYTES[1].a/w3193 ), .Z(n5902) );
  XOR \SUBBYTES[1].a/U5586  ( .A(\SUBBYTES[1].a/w3183 ), .B(
        \SUBBYTES[1].a/w3186 ), .Z(n5903) );
  XOR \SUBBYTES[1].a/U5585  ( .A(\SUBBYTES[1].a/w3158 ), .B(
        \SUBBYTES[1].a/w3159 ), .Z(n5904) );
  XOR \SUBBYTES[1].a/U5584  ( .A(\SUBBYTES[1].a/w3143 ), .B(
        \SUBBYTES[1].a/w3146 ), .Z(n5905) );
  XOR \SUBBYTES[1].a/U5582  ( .A(n6910), .B(n5908), .Z(n5906) );
  XOR \SUBBYTES[1].a/U5581  ( .A(n6912), .B(n6911), .Z(n5907) );
  XOR \SUBBYTES[1].a/U5580  ( .A(\SUBBYTES[1].a/w3151 ), .B(
        \SUBBYTES[1].a/w3178 ), .Z(n5908) );
  XOR \SUBBYTES[1].a/U5578  ( .A(n6913), .B(n5911), .Z(n5909) );
  XOR \SUBBYTES[1].a/U5577  ( .A(\SUBBYTES[1].a/w3184 ), .B(
        \SUBBYTES[1].a/w3186 ), .Z(n5910) );
  XOR \SUBBYTES[1].a/U5576  ( .A(\SUBBYTES[1].a/w3144 ), .B(
        \SUBBYTES[1].a/w3176 ), .Z(n5911) );
  XOR \SUBBYTES[1].a/U5575  ( .A(\SUBBYTES[1].a/w2976 ), .B(
        \SUBBYTES[1].a/w2977 ), .Z(n6915) );
  XOR \SUBBYTES[1].a/U5574  ( .A(n6915), .B(n5912), .Z(n6914) );
  XOR \SUBBYTES[1].a/U5573  ( .A(\SUBBYTES[1].a/w2969 ), .B(
        \SUBBYTES[1].a/w2986 ), .Z(n5912) );
  XOR \SUBBYTES[1].a/U5571  ( .A(\SUBBYTES[1].a/w2968 ), .B(
        \SUBBYTES[1].a/w2983 ), .Z(n5913) );
  XOR \SUBBYTES[1].a/U5570  ( .A(n6915), .B(n5914), .Z(n7098) );
  XOR \SUBBYTES[1].a/U5569  ( .A(\SUBBYTES[1].a/w2983 ), .B(
        \SUBBYTES[1].a/w2984 ), .Z(n5914) );
  XOR \SUBBYTES[1].a/U5568  ( .A(\SUBBYTES[1].a/w2945 ), .B(n5915), .Z(n6917)
         );
  XOR \SUBBYTES[1].a/U5567  ( .A(\SUBBYTES[1].a/w2936 ), .B(
        \SUBBYTES[1].a/w2937 ), .Z(n5915) );
  XOR \SUBBYTES[1].a/U5565  ( .A(\SUBBYTES[1].a/w2947 ), .B(n7098), .Z(n5916)
         );
  XOR \SUBBYTES[1].a/U5564  ( .A(n5918), .B(n5917), .Z(n6918) );
  XOR \SUBBYTES[1].a/U5563  ( .A(n5920), .B(n5919), .Z(n5917) );
  XOR \SUBBYTES[1].a/U5562  ( .A(\SUBBYTES[1].a/w2983 ), .B(
        \SUBBYTES[1].a/w2984 ), .Z(n5918) );
  XOR \SUBBYTES[1].a/U5561  ( .A(\SUBBYTES[1].a/w2947 ), .B(
        \SUBBYTES[1].a/w2971 ), .Z(n5919) );
  XOR \SUBBYTES[1].a/U5560  ( .A(\SUBBYTES[1].a/w2936 ), .B(
        \SUBBYTES[1].a/w2945 ), .Z(n5920) );
  XOR \SUBBYTES[1].a/U5559  ( .A(\SUBBYTES[1].a/w2968 ), .B(n5921), .Z(n6916)
         );
  XOR \SUBBYTES[1].a/U5558  ( .A(\SUBBYTES[1].a/w2951 ), .B(
        \SUBBYTES[1].a/w2954 ), .Z(n5921) );
  XOR \SUBBYTES[1].a/U5556  ( .A(\SUBBYTES[1].a/w2939 ), .B(n6918), .Z(n5922)
         );
  XOR \SUBBYTES[1].a/U5554  ( .A(\SUBBYTES[1].a/w2971 ), .B(
        \SUBBYTES[1].a/w2984 ), .Z(n5923) );
  XOR \SUBBYTES[1].a/U5552  ( .A(n5927), .B(n5926), .Z(n5924) );
  XOR \SUBBYTES[1].a/U5551  ( .A(n5929), .B(n5928), .Z(n5925) );
  XOR \SUBBYTES[1].a/U5550  ( .A(\SUBBYTES[1].a/w2983 ), .B(
        \SUBBYTES[1].a/w2986 ), .Z(n5926) );
  XOR \SUBBYTES[1].a/U5549  ( .A(\SUBBYTES[1].a/w2976 ), .B(
        \SUBBYTES[1].a/w2979 ), .Z(n5927) );
  XOR \SUBBYTES[1].a/U5548  ( .A(\SUBBYTES[1].a/w2951 ), .B(
        \SUBBYTES[1].a/w2952 ), .Z(n5928) );
  XOR \SUBBYTES[1].a/U5547  ( .A(\SUBBYTES[1].a/w2936 ), .B(
        \SUBBYTES[1].a/w2939 ), .Z(n5929) );
  XOR \SUBBYTES[1].a/U5545  ( .A(n6915), .B(n5932), .Z(n5930) );
  XOR \SUBBYTES[1].a/U5544  ( .A(n6917), .B(n6916), .Z(n5931) );
  XOR \SUBBYTES[1].a/U5543  ( .A(\SUBBYTES[1].a/w2944 ), .B(
        \SUBBYTES[1].a/w2971 ), .Z(n5932) );
  XOR \SUBBYTES[1].a/U5541  ( .A(n6918), .B(n5935), .Z(n5933) );
  XOR \SUBBYTES[1].a/U5540  ( .A(\SUBBYTES[1].a/w2977 ), .B(
        \SUBBYTES[1].a/w2979 ), .Z(n5934) );
  XOR \SUBBYTES[1].a/U5539  ( .A(\SUBBYTES[1].a/w2937 ), .B(
        \SUBBYTES[1].a/w2969 ), .Z(n5935) );
  XOR \SUBBYTES[1].a/U5538  ( .A(\SUBBYTES[1].a/w2769 ), .B(
        \SUBBYTES[1].a/w2770 ), .Z(n6920) );
  XOR \SUBBYTES[1].a/U5537  ( .A(n6920), .B(n5936), .Z(n6919) );
  XOR \SUBBYTES[1].a/U5536  ( .A(\SUBBYTES[1].a/w2762 ), .B(
        \SUBBYTES[1].a/w2779 ), .Z(n5936) );
  XOR \SUBBYTES[1].a/U5534  ( .A(\SUBBYTES[1].a/w2761 ), .B(
        \SUBBYTES[1].a/w2776 ), .Z(n5937) );
  XOR \SUBBYTES[1].a/U5533  ( .A(n6920), .B(n5938), .Z(n7099) );
  XOR \SUBBYTES[1].a/U5532  ( .A(\SUBBYTES[1].a/w2776 ), .B(
        \SUBBYTES[1].a/w2777 ), .Z(n5938) );
  XOR \SUBBYTES[1].a/U5531  ( .A(\SUBBYTES[1].a/w2738 ), .B(n5939), .Z(n6922)
         );
  XOR \SUBBYTES[1].a/U5530  ( .A(\SUBBYTES[1].a/w2729 ), .B(
        \SUBBYTES[1].a/w2730 ), .Z(n5939) );
  XOR \SUBBYTES[1].a/U5528  ( .A(\SUBBYTES[1].a/w2740 ), .B(n7099), .Z(n5940)
         );
  XOR \SUBBYTES[1].a/U5527  ( .A(n5942), .B(n5941), .Z(n6923) );
  XOR \SUBBYTES[1].a/U5526  ( .A(n5944), .B(n5943), .Z(n5941) );
  XOR \SUBBYTES[1].a/U5525  ( .A(\SUBBYTES[1].a/w2776 ), .B(
        \SUBBYTES[1].a/w2777 ), .Z(n5942) );
  XOR \SUBBYTES[1].a/U5524  ( .A(\SUBBYTES[1].a/w2740 ), .B(
        \SUBBYTES[1].a/w2764 ), .Z(n5943) );
  XOR \SUBBYTES[1].a/U5523  ( .A(\SUBBYTES[1].a/w2729 ), .B(
        \SUBBYTES[1].a/w2738 ), .Z(n5944) );
  XOR \SUBBYTES[1].a/U5522  ( .A(\SUBBYTES[1].a/w2761 ), .B(n5945), .Z(n6921)
         );
  XOR \SUBBYTES[1].a/U5521  ( .A(\SUBBYTES[1].a/w2744 ), .B(
        \SUBBYTES[1].a/w2747 ), .Z(n5945) );
  XOR \SUBBYTES[1].a/U5519  ( .A(\SUBBYTES[1].a/w2732 ), .B(n6923), .Z(n5946)
         );
  XOR \SUBBYTES[1].a/U5517  ( .A(\SUBBYTES[1].a/w2764 ), .B(
        \SUBBYTES[1].a/w2777 ), .Z(n5947) );
  XOR \SUBBYTES[1].a/U5515  ( .A(n5951), .B(n5950), .Z(n5948) );
  XOR \SUBBYTES[1].a/U5514  ( .A(n5953), .B(n5952), .Z(n5949) );
  XOR \SUBBYTES[1].a/U5513  ( .A(\SUBBYTES[1].a/w2776 ), .B(
        \SUBBYTES[1].a/w2779 ), .Z(n5950) );
  XOR \SUBBYTES[1].a/U5512  ( .A(\SUBBYTES[1].a/w2769 ), .B(
        \SUBBYTES[1].a/w2772 ), .Z(n5951) );
  XOR \SUBBYTES[1].a/U5511  ( .A(\SUBBYTES[1].a/w2744 ), .B(
        \SUBBYTES[1].a/w2745 ), .Z(n5952) );
  XOR \SUBBYTES[1].a/U5510  ( .A(\SUBBYTES[1].a/w2729 ), .B(
        \SUBBYTES[1].a/w2732 ), .Z(n5953) );
  XOR \SUBBYTES[1].a/U5508  ( .A(n6920), .B(n5956), .Z(n5954) );
  XOR \SUBBYTES[1].a/U5507  ( .A(n6922), .B(n6921), .Z(n5955) );
  XOR \SUBBYTES[1].a/U5506  ( .A(\SUBBYTES[1].a/w2737 ), .B(
        \SUBBYTES[1].a/w2764 ), .Z(n5956) );
  XOR \SUBBYTES[1].a/U5504  ( .A(n6923), .B(n5959), .Z(n5957) );
  XOR \SUBBYTES[1].a/U5503  ( .A(\SUBBYTES[1].a/w2770 ), .B(
        \SUBBYTES[1].a/w2772 ), .Z(n5958) );
  XOR \SUBBYTES[1].a/U5502  ( .A(\SUBBYTES[1].a/w2730 ), .B(
        \SUBBYTES[1].a/w2762 ), .Z(n5959) );
  XOR \SUBBYTES[1].a/U5501  ( .A(\SUBBYTES[1].a/w2562 ), .B(
        \SUBBYTES[1].a/w2563 ), .Z(n6925) );
  XOR \SUBBYTES[1].a/U5500  ( .A(n6925), .B(n5960), .Z(n6924) );
  XOR \SUBBYTES[1].a/U5499  ( .A(\SUBBYTES[1].a/w2555 ), .B(
        \SUBBYTES[1].a/w2572 ), .Z(n5960) );
  XOR \SUBBYTES[1].a/U5497  ( .A(\SUBBYTES[1].a/w2554 ), .B(
        \SUBBYTES[1].a/w2569 ), .Z(n5961) );
  XOR \SUBBYTES[1].a/U5496  ( .A(n6925), .B(n5962), .Z(n7100) );
  XOR \SUBBYTES[1].a/U5495  ( .A(\SUBBYTES[1].a/w2569 ), .B(
        \SUBBYTES[1].a/w2570 ), .Z(n5962) );
  XOR \SUBBYTES[1].a/U5494  ( .A(\SUBBYTES[1].a/w2531 ), .B(n5963), .Z(n6927)
         );
  XOR \SUBBYTES[1].a/U5493  ( .A(\SUBBYTES[1].a/w2522 ), .B(
        \SUBBYTES[1].a/w2523 ), .Z(n5963) );
  XOR \SUBBYTES[1].a/U5491  ( .A(\SUBBYTES[1].a/w2533 ), .B(n7100), .Z(n5964)
         );
  XOR \SUBBYTES[1].a/U5490  ( .A(n5966), .B(n5965), .Z(n6928) );
  XOR \SUBBYTES[1].a/U5489  ( .A(n5968), .B(n5967), .Z(n5965) );
  XOR \SUBBYTES[1].a/U5488  ( .A(\SUBBYTES[1].a/w2569 ), .B(
        \SUBBYTES[1].a/w2570 ), .Z(n5966) );
  XOR \SUBBYTES[1].a/U5487  ( .A(\SUBBYTES[1].a/w2533 ), .B(
        \SUBBYTES[1].a/w2557 ), .Z(n5967) );
  XOR \SUBBYTES[1].a/U5486  ( .A(\SUBBYTES[1].a/w2522 ), .B(
        \SUBBYTES[1].a/w2531 ), .Z(n5968) );
  XOR \SUBBYTES[1].a/U5485  ( .A(\SUBBYTES[1].a/w2554 ), .B(n5969), .Z(n6926)
         );
  XOR \SUBBYTES[1].a/U5484  ( .A(\SUBBYTES[1].a/w2537 ), .B(
        \SUBBYTES[1].a/w2540 ), .Z(n5969) );
  XOR \SUBBYTES[1].a/U5482  ( .A(\SUBBYTES[1].a/w2525 ), .B(n6928), .Z(n5970)
         );
  XOR \SUBBYTES[1].a/U5480  ( .A(\SUBBYTES[1].a/w2557 ), .B(
        \SUBBYTES[1].a/w2570 ), .Z(n5971) );
  XOR \SUBBYTES[1].a/U5478  ( .A(n5975), .B(n5974), .Z(n5972) );
  XOR \SUBBYTES[1].a/U5477  ( .A(n5977), .B(n5976), .Z(n5973) );
  XOR \SUBBYTES[1].a/U5476  ( .A(\SUBBYTES[1].a/w2569 ), .B(
        \SUBBYTES[1].a/w2572 ), .Z(n5974) );
  XOR \SUBBYTES[1].a/U5475  ( .A(\SUBBYTES[1].a/w2562 ), .B(
        \SUBBYTES[1].a/w2565 ), .Z(n5975) );
  XOR \SUBBYTES[1].a/U5474  ( .A(\SUBBYTES[1].a/w2537 ), .B(
        \SUBBYTES[1].a/w2538 ), .Z(n5976) );
  XOR \SUBBYTES[1].a/U5473  ( .A(\SUBBYTES[1].a/w2522 ), .B(
        \SUBBYTES[1].a/w2525 ), .Z(n5977) );
  XOR \SUBBYTES[1].a/U5471  ( .A(n6925), .B(n5980), .Z(n5978) );
  XOR \SUBBYTES[1].a/U5470  ( .A(n6927), .B(n6926), .Z(n5979) );
  XOR \SUBBYTES[1].a/U5469  ( .A(\SUBBYTES[1].a/w2530 ), .B(
        \SUBBYTES[1].a/w2557 ), .Z(n5980) );
  XOR \SUBBYTES[1].a/U5467  ( .A(n6928), .B(n5983), .Z(n5981) );
  XOR \SUBBYTES[1].a/U5466  ( .A(\SUBBYTES[1].a/w2563 ), .B(
        \SUBBYTES[1].a/w2565 ), .Z(n5982) );
  XOR \SUBBYTES[1].a/U5465  ( .A(\SUBBYTES[1].a/w2523 ), .B(
        \SUBBYTES[1].a/w2555 ), .Z(n5983) );
  XOR \SUBBYTES[1].a/U5464  ( .A(\SUBBYTES[1].a/w2355 ), .B(
        \SUBBYTES[1].a/w2356 ), .Z(n6930) );
  XOR \SUBBYTES[1].a/U5463  ( .A(n6930), .B(n5984), .Z(n6929) );
  XOR \SUBBYTES[1].a/U5462  ( .A(\SUBBYTES[1].a/w2348 ), .B(
        \SUBBYTES[1].a/w2365 ), .Z(n5984) );
  XOR \SUBBYTES[1].a/U5460  ( .A(\SUBBYTES[1].a/w2347 ), .B(
        \SUBBYTES[1].a/w2362 ), .Z(n5985) );
  XOR \SUBBYTES[1].a/U5459  ( .A(n6930), .B(n5986), .Z(n7101) );
  XOR \SUBBYTES[1].a/U5458  ( .A(\SUBBYTES[1].a/w2362 ), .B(
        \SUBBYTES[1].a/w2363 ), .Z(n5986) );
  XOR \SUBBYTES[1].a/U5457  ( .A(\SUBBYTES[1].a/w2324 ), .B(n5987), .Z(n6932)
         );
  XOR \SUBBYTES[1].a/U5456  ( .A(\SUBBYTES[1].a/w2315 ), .B(
        \SUBBYTES[1].a/w2316 ), .Z(n5987) );
  XOR \SUBBYTES[1].a/U5454  ( .A(\SUBBYTES[1].a/w2326 ), .B(n7101), .Z(n5988)
         );
  XOR \SUBBYTES[1].a/U5453  ( .A(n5990), .B(n5989), .Z(n6933) );
  XOR \SUBBYTES[1].a/U5452  ( .A(n5992), .B(n5991), .Z(n5989) );
  XOR \SUBBYTES[1].a/U5451  ( .A(\SUBBYTES[1].a/w2362 ), .B(
        \SUBBYTES[1].a/w2363 ), .Z(n5990) );
  XOR \SUBBYTES[1].a/U5450  ( .A(\SUBBYTES[1].a/w2326 ), .B(
        \SUBBYTES[1].a/w2350 ), .Z(n5991) );
  XOR \SUBBYTES[1].a/U5449  ( .A(\SUBBYTES[1].a/w2315 ), .B(
        \SUBBYTES[1].a/w2324 ), .Z(n5992) );
  XOR \SUBBYTES[1].a/U5448  ( .A(\SUBBYTES[1].a/w2347 ), .B(n5993), .Z(n6931)
         );
  XOR \SUBBYTES[1].a/U5447  ( .A(\SUBBYTES[1].a/w2330 ), .B(
        \SUBBYTES[1].a/w2333 ), .Z(n5993) );
  XOR \SUBBYTES[1].a/U5445  ( .A(\SUBBYTES[1].a/w2318 ), .B(n6933), .Z(n5994)
         );
  XOR \SUBBYTES[1].a/U5443  ( .A(\SUBBYTES[1].a/w2350 ), .B(
        \SUBBYTES[1].a/w2363 ), .Z(n5995) );
  XOR \SUBBYTES[1].a/U5441  ( .A(n5999), .B(n5998), .Z(n5996) );
  XOR \SUBBYTES[1].a/U5440  ( .A(n6001), .B(n6000), .Z(n5997) );
  XOR \SUBBYTES[1].a/U5439  ( .A(\SUBBYTES[1].a/w2362 ), .B(
        \SUBBYTES[1].a/w2365 ), .Z(n5998) );
  XOR \SUBBYTES[1].a/U5438  ( .A(\SUBBYTES[1].a/w2355 ), .B(
        \SUBBYTES[1].a/w2358 ), .Z(n5999) );
  XOR \SUBBYTES[1].a/U5437  ( .A(\SUBBYTES[1].a/w2330 ), .B(
        \SUBBYTES[1].a/w2331 ), .Z(n6000) );
  XOR \SUBBYTES[1].a/U5436  ( .A(\SUBBYTES[1].a/w2315 ), .B(
        \SUBBYTES[1].a/w2318 ), .Z(n6001) );
  XOR \SUBBYTES[1].a/U5434  ( .A(n6930), .B(n6004), .Z(n6002) );
  XOR \SUBBYTES[1].a/U5433  ( .A(n6932), .B(n6931), .Z(n6003) );
  XOR \SUBBYTES[1].a/U5432  ( .A(\SUBBYTES[1].a/w2323 ), .B(
        \SUBBYTES[1].a/w2350 ), .Z(n6004) );
  XOR \SUBBYTES[1].a/U5430  ( .A(n6933), .B(n6007), .Z(n6005) );
  XOR \SUBBYTES[1].a/U5429  ( .A(\SUBBYTES[1].a/w2356 ), .B(
        \SUBBYTES[1].a/w2358 ), .Z(n6006) );
  XOR \SUBBYTES[1].a/U5428  ( .A(\SUBBYTES[1].a/w2316 ), .B(
        \SUBBYTES[1].a/w2348 ), .Z(n6007) );
  XOR \SUBBYTES[1].a/U5427  ( .A(\SUBBYTES[1].a/w2148 ), .B(
        \SUBBYTES[1].a/w2149 ), .Z(n6935) );
  XOR \SUBBYTES[1].a/U5426  ( .A(n6935), .B(n6008), .Z(n6934) );
  XOR \SUBBYTES[1].a/U5425  ( .A(\SUBBYTES[1].a/w2141 ), .B(
        \SUBBYTES[1].a/w2158 ), .Z(n6008) );
  XOR \SUBBYTES[1].a/U5423  ( .A(\SUBBYTES[1].a/w2140 ), .B(
        \SUBBYTES[1].a/w2155 ), .Z(n6009) );
  XOR \SUBBYTES[1].a/U5422  ( .A(n6935), .B(n6010), .Z(n7102) );
  XOR \SUBBYTES[1].a/U5421  ( .A(\SUBBYTES[1].a/w2155 ), .B(
        \SUBBYTES[1].a/w2156 ), .Z(n6010) );
  XOR \SUBBYTES[1].a/U5420  ( .A(\SUBBYTES[1].a/w2117 ), .B(n6011), .Z(n6937)
         );
  XOR \SUBBYTES[1].a/U5419  ( .A(\SUBBYTES[1].a/w2108 ), .B(
        \SUBBYTES[1].a/w2109 ), .Z(n6011) );
  XOR \SUBBYTES[1].a/U5417  ( .A(\SUBBYTES[1].a/w2119 ), .B(n7102), .Z(n6012)
         );
  XOR \SUBBYTES[1].a/U5416  ( .A(n6014), .B(n6013), .Z(n6938) );
  XOR \SUBBYTES[1].a/U5415  ( .A(n6016), .B(n6015), .Z(n6013) );
  XOR \SUBBYTES[1].a/U5414  ( .A(\SUBBYTES[1].a/w2155 ), .B(
        \SUBBYTES[1].a/w2156 ), .Z(n6014) );
  XOR \SUBBYTES[1].a/U5413  ( .A(\SUBBYTES[1].a/w2119 ), .B(
        \SUBBYTES[1].a/w2143 ), .Z(n6015) );
  XOR \SUBBYTES[1].a/U5412  ( .A(\SUBBYTES[1].a/w2108 ), .B(
        \SUBBYTES[1].a/w2117 ), .Z(n6016) );
  XOR \SUBBYTES[1].a/U5411  ( .A(\SUBBYTES[1].a/w2140 ), .B(n6017), .Z(n6936)
         );
  XOR \SUBBYTES[1].a/U5410  ( .A(\SUBBYTES[1].a/w2123 ), .B(
        \SUBBYTES[1].a/w2126 ), .Z(n6017) );
  XOR \SUBBYTES[1].a/U5408  ( .A(\SUBBYTES[1].a/w2111 ), .B(n6938), .Z(n6018)
         );
  XOR \SUBBYTES[1].a/U5406  ( .A(\SUBBYTES[1].a/w2143 ), .B(
        \SUBBYTES[1].a/w2156 ), .Z(n6019) );
  XOR \SUBBYTES[1].a/U5404  ( .A(n6023), .B(n6022), .Z(n6020) );
  XOR \SUBBYTES[1].a/U5403  ( .A(n6025), .B(n6024), .Z(n6021) );
  XOR \SUBBYTES[1].a/U5402  ( .A(\SUBBYTES[1].a/w2155 ), .B(
        \SUBBYTES[1].a/w2158 ), .Z(n6022) );
  XOR \SUBBYTES[1].a/U5401  ( .A(\SUBBYTES[1].a/w2148 ), .B(
        \SUBBYTES[1].a/w2151 ), .Z(n6023) );
  XOR \SUBBYTES[1].a/U5400  ( .A(\SUBBYTES[1].a/w2123 ), .B(
        \SUBBYTES[1].a/w2124 ), .Z(n6024) );
  XOR \SUBBYTES[1].a/U5399  ( .A(\SUBBYTES[1].a/w2108 ), .B(
        \SUBBYTES[1].a/w2111 ), .Z(n6025) );
  XOR \SUBBYTES[1].a/U5397  ( .A(n6935), .B(n6028), .Z(n6026) );
  XOR \SUBBYTES[1].a/U5396  ( .A(n6937), .B(n6936), .Z(n6027) );
  XOR \SUBBYTES[1].a/U5395  ( .A(\SUBBYTES[1].a/w2116 ), .B(
        \SUBBYTES[1].a/w2143 ), .Z(n6028) );
  XOR \SUBBYTES[1].a/U5393  ( .A(n6938), .B(n6031), .Z(n6029) );
  XOR \SUBBYTES[1].a/U5392  ( .A(\SUBBYTES[1].a/w2149 ), .B(
        \SUBBYTES[1].a/w2151 ), .Z(n6030) );
  XOR \SUBBYTES[1].a/U5391  ( .A(\SUBBYTES[1].a/w2109 ), .B(
        \SUBBYTES[1].a/w2141 ), .Z(n6031) );
  XOR \SUBBYTES[1].a/U5390  ( .A(\SUBBYTES[1].a/w1941 ), .B(
        \SUBBYTES[1].a/w1942 ), .Z(n6940) );
  XOR \SUBBYTES[1].a/U5389  ( .A(n6940), .B(n6032), .Z(n6939) );
  XOR \SUBBYTES[1].a/U5388  ( .A(\SUBBYTES[1].a/w1934 ), .B(
        \SUBBYTES[1].a/w1951 ), .Z(n6032) );
  XOR \SUBBYTES[1].a/U5386  ( .A(\SUBBYTES[1].a/w1933 ), .B(
        \SUBBYTES[1].a/w1948 ), .Z(n6033) );
  XOR \SUBBYTES[1].a/U5385  ( .A(n6940), .B(n6034), .Z(n7103) );
  XOR \SUBBYTES[1].a/U5384  ( .A(\SUBBYTES[1].a/w1948 ), .B(
        \SUBBYTES[1].a/w1949 ), .Z(n6034) );
  XOR \SUBBYTES[1].a/U5383  ( .A(\SUBBYTES[1].a/w1910 ), .B(n6035), .Z(n6942)
         );
  XOR \SUBBYTES[1].a/U5382  ( .A(\SUBBYTES[1].a/w1901 ), .B(
        \SUBBYTES[1].a/w1902 ), .Z(n6035) );
  XOR \SUBBYTES[1].a/U5380  ( .A(\SUBBYTES[1].a/w1912 ), .B(n7103), .Z(n6036)
         );
  XOR \SUBBYTES[1].a/U5379  ( .A(n6038), .B(n6037), .Z(n6943) );
  XOR \SUBBYTES[1].a/U5378  ( .A(n6040), .B(n6039), .Z(n6037) );
  XOR \SUBBYTES[1].a/U5377  ( .A(\SUBBYTES[1].a/w1948 ), .B(
        \SUBBYTES[1].a/w1949 ), .Z(n6038) );
  XOR \SUBBYTES[1].a/U5376  ( .A(\SUBBYTES[1].a/w1912 ), .B(
        \SUBBYTES[1].a/w1936 ), .Z(n6039) );
  XOR \SUBBYTES[1].a/U5375  ( .A(\SUBBYTES[1].a/w1901 ), .B(
        \SUBBYTES[1].a/w1910 ), .Z(n6040) );
  XOR \SUBBYTES[1].a/U5374  ( .A(\SUBBYTES[1].a/w1933 ), .B(n6041), .Z(n6941)
         );
  XOR \SUBBYTES[1].a/U5373  ( .A(\SUBBYTES[1].a/w1916 ), .B(
        \SUBBYTES[1].a/w1919 ), .Z(n6041) );
  XOR \SUBBYTES[1].a/U5371  ( .A(\SUBBYTES[1].a/w1904 ), .B(n6943), .Z(n6042)
         );
  XOR \SUBBYTES[1].a/U5369  ( .A(\SUBBYTES[1].a/w1936 ), .B(
        \SUBBYTES[1].a/w1949 ), .Z(n6043) );
  XOR \SUBBYTES[1].a/U5367  ( .A(n6047), .B(n6046), .Z(n6044) );
  XOR \SUBBYTES[1].a/U5366  ( .A(n6049), .B(n6048), .Z(n6045) );
  XOR \SUBBYTES[1].a/U5365  ( .A(\SUBBYTES[1].a/w1948 ), .B(
        \SUBBYTES[1].a/w1951 ), .Z(n6046) );
  XOR \SUBBYTES[1].a/U5364  ( .A(\SUBBYTES[1].a/w1941 ), .B(
        \SUBBYTES[1].a/w1944 ), .Z(n6047) );
  XOR \SUBBYTES[1].a/U5363  ( .A(\SUBBYTES[1].a/w1916 ), .B(
        \SUBBYTES[1].a/w1917 ), .Z(n6048) );
  XOR \SUBBYTES[1].a/U5362  ( .A(\SUBBYTES[1].a/w1901 ), .B(
        \SUBBYTES[1].a/w1904 ), .Z(n6049) );
  XOR \SUBBYTES[1].a/U5360  ( .A(n6940), .B(n6052), .Z(n6050) );
  XOR \SUBBYTES[1].a/U5359  ( .A(n6942), .B(n6941), .Z(n6051) );
  XOR \SUBBYTES[1].a/U5358  ( .A(\SUBBYTES[1].a/w1909 ), .B(
        \SUBBYTES[1].a/w1936 ), .Z(n6052) );
  XOR \SUBBYTES[1].a/U5356  ( .A(n6943), .B(n6055), .Z(n6053) );
  XOR \SUBBYTES[1].a/U5355  ( .A(\SUBBYTES[1].a/w1942 ), .B(
        \SUBBYTES[1].a/w1944 ), .Z(n6054) );
  XOR \SUBBYTES[1].a/U5354  ( .A(\SUBBYTES[1].a/w1902 ), .B(
        \SUBBYTES[1].a/w1934 ), .Z(n6055) );
  XOR \SUBBYTES[1].a/U5353  ( .A(\SUBBYTES[1].a/w1734 ), .B(
        \SUBBYTES[1].a/w1735 ), .Z(n6945) );
  XOR \SUBBYTES[1].a/U5352  ( .A(n6945), .B(n6056), .Z(n6944) );
  XOR \SUBBYTES[1].a/U5351  ( .A(\SUBBYTES[1].a/w1727 ), .B(
        \SUBBYTES[1].a/w1744 ), .Z(n6056) );
  XOR \SUBBYTES[1].a/U5349  ( .A(\SUBBYTES[1].a/w1726 ), .B(
        \SUBBYTES[1].a/w1741 ), .Z(n6057) );
  XOR \SUBBYTES[1].a/U5348  ( .A(n6945), .B(n6058), .Z(n7104) );
  XOR \SUBBYTES[1].a/U5347  ( .A(\SUBBYTES[1].a/w1741 ), .B(
        \SUBBYTES[1].a/w1742 ), .Z(n6058) );
  XOR \SUBBYTES[1].a/U5346  ( .A(\SUBBYTES[1].a/w1703 ), .B(n6059), .Z(n6947)
         );
  XOR \SUBBYTES[1].a/U5345  ( .A(\SUBBYTES[1].a/w1694 ), .B(
        \SUBBYTES[1].a/w1695 ), .Z(n6059) );
  XOR \SUBBYTES[1].a/U5343  ( .A(\SUBBYTES[1].a/w1705 ), .B(n7104), .Z(n6060)
         );
  XOR \SUBBYTES[1].a/U5342  ( .A(n6062), .B(n6061), .Z(n6948) );
  XOR \SUBBYTES[1].a/U5341  ( .A(n6064), .B(n6063), .Z(n6061) );
  XOR \SUBBYTES[1].a/U5340  ( .A(\SUBBYTES[1].a/w1741 ), .B(
        \SUBBYTES[1].a/w1742 ), .Z(n6062) );
  XOR \SUBBYTES[1].a/U5339  ( .A(\SUBBYTES[1].a/w1705 ), .B(
        \SUBBYTES[1].a/w1729 ), .Z(n6063) );
  XOR \SUBBYTES[1].a/U5338  ( .A(\SUBBYTES[1].a/w1694 ), .B(
        \SUBBYTES[1].a/w1703 ), .Z(n6064) );
  XOR \SUBBYTES[1].a/U5337  ( .A(\SUBBYTES[1].a/w1726 ), .B(n6065), .Z(n6946)
         );
  XOR \SUBBYTES[1].a/U5336  ( .A(\SUBBYTES[1].a/w1709 ), .B(
        \SUBBYTES[1].a/w1712 ), .Z(n6065) );
  XOR \SUBBYTES[1].a/U5334  ( .A(\SUBBYTES[1].a/w1697 ), .B(n6948), .Z(n6066)
         );
  XOR \SUBBYTES[1].a/U5332  ( .A(\SUBBYTES[1].a/w1729 ), .B(
        \SUBBYTES[1].a/w1742 ), .Z(n6067) );
  XOR \SUBBYTES[1].a/U5330  ( .A(n6071), .B(n6070), .Z(n6068) );
  XOR \SUBBYTES[1].a/U5329  ( .A(n6073), .B(n6072), .Z(n6069) );
  XOR \SUBBYTES[1].a/U5328  ( .A(\SUBBYTES[1].a/w1741 ), .B(
        \SUBBYTES[1].a/w1744 ), .Z(n6070) );
  XOR \SUBBYTES[1].a/U5327  ( .A(\SUBBYTES[1].a/w1734 ), .B(
        \SUBBYTES[1].a/w1737 ), .Z(n6071) );
  XOR \SUBBYTES[1].a/U5326  ( .A(\SUBBYTES[1].a/w1709 ), .B(
        \SUBBYTES[1].a/w1710 ), .Z(n6072) );
  XOR \SUBBYTES[1].a/U5325  ( .A(\SUBBYTES[1].a/w1694 ), .B(
        \SUBBYTES[1].a/w1697 ), .Z(n6073) );
  XOR \SUBBYTES[1].a/U5323  ( .A(n6945), .B(n6076), .Z(n6074) );
  XOR \SUBBYTES[1].a/U5322  ( .A(n6947), .B(n6946), .Z(n6075) );
  XOR \SUBBYTES[1].a/U5321  ( .A(\SUBBYTES[1].a/w1702 ), .B(
        \SUBBYTES[1].a/w1729 ), .Z(n6076) );
  XOR \SUBBYTES[1].a/U5319  ( .A(n6948), .B(n6079), .Z(n6077) );
  XOR \SUBBYTES[1].a/U5318  ( .A(\SUBBYTES[1].a/w1735 ), .B(
        \SUBBYTES[1].a/w1737 ), .Z(n6078) );
  XOR \SUBBYTES[1].a/U5317  ( .A(\SUBBYTES[1].a/w1695 ), .B(
        \SUBBYTES[1].a/w1727 ), .Z(n6079) );
  XOR \SUBBYTES[1].a/U5316  ( .A(\SUBBYTES[1].a/w1527 ), .B(
        \SUBBYTES[1].a/w1528 ), .Z(n6950) );
  XOR \SUBBYTES[1].a/U5315  ( .A(n6950), .B(n6080), .Z(n6949) );
  XOR \SUBBYTES[1].a/U5314  ( .A(\SUBBYTES[1].a/w1520 ), .B(
        \SUBBYTES[1].a/w1537 ), .Z(n6080) );
  XOR \SUBBYTES[1].a/U5312  ( .A(\SUBBYTES[1].a/w1519 ), .B(
        \SUBBYTES[1].a/w1534 ), .Z(n6081) );
  XOR \SUBBYTES[1].a/U5311  ( .A(n6950), .B(n6082), .Z(n7105) );
  XOR \SUBBYTES[1].a/U5310  ( .A(\SUBBYTES[1].a/w1534 ), .B(
        \SUBBYTES[1].a/w1535 ), .Z(n6082) );
  XOR \SUBBYTES[1].a/U5309  ( .A(\SUBBYTES[1].a/w1496 ), .B(n6083), .Z(n6952)
         );
  XOR \SUBBYTES[1].a/U5308  ( .A(\SUBBYTES[1].a/w1487 ), .B(
        \SUBBYTES[1].a/w1488 ), .Z(n6083) );
  XOR \SUBBYTES[1].a/U5306  ( .A(\SUBBYTES[1].a/w1498 ), .B(n7105), .Z(n6084)
         );
  XOR \SUBBYTES[1].a/U5305  ( .A(n6086), .B(n6085), .Z(n6953) );
  XOR \SUBBYTES[1].a/U5304  ( .A(n6088), .B(n6087), .Z(n6085) );
  XOR \SUBBYTES[1].a/U5303  ( .A(\SUBBYTES[1].a/w1534 ), .B(
        \SUBBYTES[1].a/w1535 ), .Z(n6086) );
  XOR \SUBBYTES[1].a/U5302  ( .A(\SUBBYTES[1].a/w1498 ), .B(
        \SUBBYTES[1].a/w1522 ), .Z(n6087) );
  XOR \SUBBYTES[1].a/U5301  ( .A(\SUBBYTES[1].a/w1487 ), .B(
        \SUBBYTES[1].a/w1496 ), .Z(n6088) );
  XOR \SUBBYTES[1].a/U5300  ( .A(\SUBBYTES[1].a/w1519 ), .B(n6089), .Z(n6951)
         );
  XOR \SUBBYTES[1].a/U5299  ( .A(\SUBBYTES[1].a/w1502 ), .B(
        \SUBBYTES[1].a/w1505 ), .Z(n6089) );
  XOR \SUBBYTES[1].a/U5297  ( .A(\SUBBYTES[1].a/w1490 ), .B(n6953), .Z(n6090)
         );
  XOR \SUBBYTES[1].a/U5295  ( .A(\SUBBYTES[1].a/w1522 ), .B(
        \SUBBYTES[1].a/w1535 ), .Z(n6091) );
  XOR \SUBBYTES[1].a/U5293  ( .A(n6095), .B(n6094), .Z(n6092) );
  XOR \SUBBYTES[1].a/U5292  ( .A(n6097), .B(n6096), .Z(n6093) );
  XOR \SUBBYTES[1].a/U5291  ( .A(\SUBBYTES[1].a/w1534 ), .B(
        \SUBBYTES[1].a/w1537 ), .Z(n6094) );
  XOR \SUBBYTES[1].a/U5290  ( .A(\SUBBYTES[1].a/w1527 ), .B(
        \SUBBYTES[1].a/w1530 ), .Z(n6095) );
  XOR \SUBBYTES[1].a/U5289  ( .A(\SUBBYTES[1].a/w1502 ), .B(
        \SUBBYTES[1].a/w1503 ), .Z(n6096) );
  XOR \SUBBYTES[1].a/U5288  ( .A(\SUBBYTES[1].a/w1487 ), .B(
        \SUBBYTES[1].a/w1490 ), .Z(n6097) );
  XOR \SUBBYTES[1].a/U5286  ( .A(n6950), .B(n6100), .Z(n6098) );
  XOR \SUBBYTES[1].a/U5285  ( .A(n6952), .B(n6951), .Z(n6099) );
  XOR \SUBBYTES[1].a/U5284  ( .A(\SUBBYTES[1].a/w1495 ), .B(
        \SUBBYTES[1].a/w1522 ), .Z(n6100) );
  XOR \SUBBYTES[1].a/U5282  ( .A(n6953), .B(n6103), .Z(n6101) );
  XOR \SUBBYTES[1].a/U5281  ( .A(\SUBBYTES[1].a/w1528 ), .B(
        \SUBBYTES[1].a/w1530 ), .Z(n6102) );
  XOR \SUBBYTES[1].a/U5280  ( .A(\SUBBYTES[1].a/w1488 ), .B(
        \SUBBYTES[1].a/w1520 ), .Z(n6103) );
  XOR \SUBBYTES[1].a/U5279  ( .A(\SUBBYTES[1].a/w1320 ), .B(
        \SUBBYTES[1].a/w1321 ), .Z(n6955) );
  XOR \SUBBYTES[1].a/U5278  ( .A(n6955), .B(n6104), .Z(n6954) );
  XOR \SUBBYTES[1].a/U5277  ( .A(\SUBBYTES[1].a/w1313 ), .B(
        \SUBBYTES[1].a/w1330 ), .Z(n6104) );
  XOR \SUBBYTES[1].a/U5275  ( .A(\SUBBYTES[1].a/w1312 ), .B(
        \SUBBYTES[1].a/w1327 ), .Z(n6105) );
  XOR \SUBBYTES[1].a/U5274  ( .A(n6955), .B(n6106), .Z(n7106) );
  XOR \SUBBYTES[1].a/U5273  ( .A(\SUBBYTES[1].a/w1327 ), .B(
        \SUBBYTES[1].a/w1328 ), .Z(n6106) );
  XOR \SUBBYTES[1].a/U5272  ( .A(\SUBBYTES[1].a/w1289 ), .B(n6107), .Z(n6957)
         );
  XOR \SUBBYTES[1].a/U5271  ( .A(\SUBBYTES[1].a/w1280 ), .B(
        \SUBBYTES[1].a/w1281 ), .Z(n6107) );
  XOR \SUBBYTES[1].a/U5269  ( .A(\SUBBYTES[1].a/w1291 ), .B(n7106), .Z(n6108)
         );
  XOR \SUBBYTES[1].a/U5268  ( .A(n6110), .B(n6109), .Z(n6958) );
  XOR \SUBBYTES[1].a/U5267  ( .A(n6112), .B(n6111), .Z(n6109) );
  XOR \SUBBYTES[1].a/U5266  ( .A(\SUBBYTES[1].a/w1327 ), .B(
        \SUBBYTES[1].a/w1328 ), .Z(n6110) );
  XOR \SUBBYTES[1].a/U5265  ( .A(\SUBBYTES[1].a/w1291 ), .B(
        \SUBBYTES[1].a/w1315 ), .Z(n6111) );
  XOR \SUBBYTES[1].a/U5264  ( .A(\SUBBYTES[1].a/w1280 ), .B(
        \SUBBYTES[1].a/w1289 ), .Z(n6112) );
  XOR \SUBBYTES[1].a/U5263  ( .A(\SUBBYTES[1].a/w1312 ), .B(n6113), .Z(n6956)
         );
  XOR \SUBBYTES[1].a/U5262  ( .A(\SUBBYTES[1].a/w1295 ), .B(
        \SUBBYTES[1].a/w1298 ), .Z(n6113) );
  XOR \SUBBYTES[1].a/U5260  ( .A(\SUBBYTES[1].a/w1283 ), .B(n6958), .Z(n6114)
         );
  XOR \SUBBYTES[1].a/U5258  ( .A(\SUBBYTES[1].a/w1315 ), .B(
        \SUBBYTES[1].a/w1328 ), .Z(n6115) );
  XOR \SUBBYTES[1].a/U5256  ( .A(n6119), .B(n6118), .Z(n6116) );
  XOR \SUBBYTES[1].a/U5255  ( .A(n6121), .B(n6120), .Z(n6117) );
  XOR \SUBBYTES[1].a/U5254  ( .A(\SUBBYTES[1].a/w1327 ), .B(
        \SUBBYTES[1].a/w1330 ), .Z(n6118) );
  XOR \SUBBYTES[1].a/U5253  ( .A(\SUBBYTES[1].a/w1320 ), .B(
        \SUBBYTES[1].a/w1323 ), .Z(n6119) );
  XOR \SUBBYTES[1].a/U5252  ( .A(\SUBBYTES[1].a/w1295 ), .B(
        \SUBBYTES[1].a/w1296 ), .Z(n6120) );
  XOR \SUBBYTES[1].a/U5251  ( .A(\SUBBYTES[1].a/w1280 ), .B(
        \SUBBYTES[1].a/w1283 ), .Z(n6121) );
  XOR \SUBBYTES[1].a/U5249  ( .A(n6955), .B(n6124), .Z(n6122) );
  XOR \SUBBYTES[1].a/U5248  ( .A(n6957), .B(n6956), .Z(n6123) );
  XOR \SUBBYTES[1].a/U5247  ( .A(\SUBBYTES[1].a/w1288 ), .B(
        \SUBBYTES[1].a/w1315 ), .Z(n6124) );
  XOR \SUBBYTES[1].a/U5245  ( .A(n6958), .B(n6127), .Z(n6125) );
  XOR \SUBBYTES[1].a/U5244  ( .A(\SUBBYTES[1].a/w1321 ), .B(
        \SUBBYTES[1].a/w1323 ), .Z(n6126) );
  XOR \SUBBYTES[1].a/U5243  ( .A(\SUBBYTES[1].a/w1281 ), .B(
        \SUBBYTES[1].a/w1313 ), .Z(n6127) );
  XOR \SUBBYTES[1].a/U5242  ( .A(\SUBBYTES[1].a/w1113 ), .B(
        \SUBBYTES[1].a/w1114 ), .Z(n6960) );
  XOR \SUBBYTES[1].a/U5241  ( .A(n6960), .B(n6128), .Z(n6959) );
  XOR \SUBBYTES[1].a/U5240  ( .A(\SUBBYTES[1].a/w1106 ), .B(
        \SUBBYTES[1].a/w1123 ), .Z(n6128) );
  XOR \SUBBYTES[1].a/U5238  ( .A(\SUBBYTES[1].a/w1105 ), .B(
        \SUBBYTES[1].a/w1120 ), .Z(n6129) );
  XOR \SUBBYTES[1].a/U5237  ( .A(n6960), .B(n6130), .Z(n7107) );
  XOR \SUBBYTES[1].a/U5236  ( .A(\SUBBYTES[1].a/w1120 ), .B(
        \SUBBYTES[1].a/w1121 ), .Z(n6130) );
  XOR \SUBBYTES[1].a/U5235  ( .A(\SUBBYTES[1].a/w1082 ), .B(n6131), .Z(n6962)
         );
  XOR \SUBBYTES[1].a/U5234  ( .A(\SUBBYTES[1].a/w1073 ), .B(
        \SUBBYTES[1].a/w1074 ), .Z(n6131) );
  XOR \SUBBYTES[1].a/U5232  ( .A(\SUBBYTES[1].a/w1084 ), .B(n7107), .Z(n6132)
         );
  XOR \SUBBYTES[1].a/U5231  ( .A(n6134), .B(n6133), .Z(n6963) );
  XOR \SUBBYTES[1].a/U5230  ( .A(n6136), .B(n6135), .Z(n6133) );
  XOR \SUBBYTES[1].a/U5229  ( .A(\SUBBYTES[1].a/w1120 ), .B(
        \SUBBYTES[1].a/w1121 ), .Z(n6134) );
  XOR \SUBBYTES[1].a/U5228  ( .A(\SUBBYTES[1].a/w1084 ), .B(
        \SUBBYTES[1].a/w1108 ), .Z(n6135) );
  XOR \SUBBYTES[1].a/U5227  ( .A(\SUBBYTES[1].a/w1073 ), .B(
        \SUBBYTES[1].a/w1082 ), .Z(n6136) );
  XOR \SUBBYTES[1].a/U5226  ( .A(\SUBBYTES[1].a/w1105 ), .B(n6137), .Z(n6961)
         );
  XOR \SUBBYTES[1].a/U5225  ( .A(\SUBBYTES[1].a/w1088 ), .B(
        \SUBBYTES[1].a/w1091 ), .Z(n6137) );
  XOR \SUBBYTES[1].a/U5223  ( .A(\SUBBYTES[1].a/w1076 ), .B(n6963), .Z(n6138)
         );
  XOR \SUBBYTES[1].a/U5221  ( .A(\SUBBYTES[1].a/w1108 ), .B(
        \SUBBYTES[1].a/w1121 ), .Z(n6139) );
  XOR \SUBBYTES[1].a/U5219  ( .A(n6143), .B(n6142), .Z(n6140) );
  XOR \SUBBYTES[1].a/U5218  ( .A(n6145), .B(n6144), .Z(n6141) );
  XOR \SUBBYTES[1].a/U5217  ( .A(\SUBBYTES[1].a/w1120 ), .B(
        \SUBBYTES[1].a/w1123 ), .Z(n6142) );
  XOR \SUBBYTES[1].a/U5216  ( .A(\SUBBYTES[1].a/w1113 ), .B(
        \SUBBYTES[1].a/w1116 ), .Z(n6143) );
  XOR \SUBBYTES[1].a/U5215  ( .A(\SUBBYTES[1].a/w1088 ), .B(
        \SUBBYTES[1].a/w1089 ), .Z(n6144) );
  XOR \SUBBYTES[1].a/U5214  ( .A(\SUBBYTES[1].a/w1073 ), .B(
        \SUBBYTES[1].a/w1076 ), .Z(n6145) );
  XOR \SUBBYTES[1].a/U5212  ( .A(n6960), .B(n6148), .Z(n6146) );
  XOR \SUBBYTES[1].a/U5211  ( .A(n6962), .B(n6961), .Z(n6147) );
  XOR \SUBBYTES[1].a/U5210  ( .A(\SUBBYTES[1].a/w1081 ), .B(
        \SUBBYTES[1].a/w1108 ), .Z(n6148) );
  XOR \SUBBYTES[1].a/U5208  ( .A(n6963), .B(n6151), .Z(n6149) );
  XOR \SUBBYTES[1].a/U5207  ( .A(\SUBBYTES[1].a/w1114 ), .B(
        \SUBBYTES[1].a/w1116 ), .Z(n6150) );
  XOR \SUBBYTES[1].a/U5206  ( .A(\SUBBYTES[1].a/w1074 ), .B(
        \SUBBYTES[1].a/w1106 ), .Z(n6151) );
  XOR \SUBBYTES[1].a/U5205  ( .A(\SUBBYTES[1].a/w906 ), .B(
        \SUBBYTES[1].a/w907 ), .Z(n6965) );
  XOR \SUBBYTES[1].a/U5204  ( .A(n6965), .B(n6152), .Z(n6964) );
  XOR \SUBBYTES[1].a/U5203  ( .A(\SUBBYTES[1].a/w899 ), .B(
        \SUBBYTES[1].a/w916 ), .Z(n6152) );
  XOR \SUBBYTES[1].a/U5201  ( .A(\SUBBYTES[1].a/w898 ), .B(
        \SUBBYTES[1].a/w913 ), .Z(n6153) );
  XOR \SUBBYTES[1].a/U5200  ( .A(n6965), .B(n6154), .Z(n7108) );
  XOR \SUBBYTES[1].a/U5199  ( .A(\SUBBYTES[1].a/w913 ), .B(
        \SUBBYTES[1].a/w914 ), .Z(n6154) );
  XOR \SUBBYTES[1].a/U5198  ( .A(\SUBBYTES[1].a/w875 ), .B(n6155), .Z(n6967)
         );
  XOR \SUBBYTES[1].a/U5197  ( .A(\SUBBYTES[1].a/w866 ), .B(
        \SUBBYTES[1].a/w867 ), .Z(n6155) );
  XOR \SUBBYTES[1].a/U5195  ( .A(\SUBBYTES[1].a/w877 ), .B(n7108), .Z(n6156)
         );
  XOR \SUBBYTES[1].a/U5194  ( .A(n6158), .B(n6157), .Z(n6968) );
  XOR \SUBBYTES[1].a/U5193  ( .A(n6160), .B(n6159), .Z(n6157) );
  XOR \SUBBYTES[1].a/U5192  ( .A(\SUBBYTES[1].a/w913 ), .B(
        \SUBBYTES[1].a/w914 ), .Z(n6158) );
  XOR \SUBBYTES[1].a/U5191  ( .A(\SUBBYTES[1].a/w877 ), .B(
        \SUBBYTES[1].a/w901 ), .Z(n6159) );
  XOR \SUBBYTES[1].a/U5190  ( .A(\SUBBYTES[1].a/w866 ), .B(
        \SUBBYTES[1].a/w875 ), .Z(n6160) );
  XOR \SUBBYTES[1].a/U5189  ( .A(\SUBBYTES[1].a/w898 ), .B(n6161), .Z(n6966)
         );
  XOR \SUBBYTES[1].a/U5188  ( .A(\SUBBYTES[1].a/w881 ), .B(
        \SUBBYTES[1].a/w884 ), .Z(n6161) );
  XOR \SUBBYTES[1].a/U5186  ( .A(\SUBBYTES[1].a/w869 ), .B(n6968), .Z(n6162)
         );
  XOR \SUBBYTES[1].a/U5184  ( .A(\SUBBYTES[1].a/w901 ), .B(
        \SUBBYTES[1].a/w914 ), .Z(n6163) );
  XOR \SUBBYTES[1].a/U5182  ( .A(n6167), .B(n6166), .Z(n6164) );
  XOR \SUBBYTES[1].a/U5181  ( .A(n6169), .B(n6168), .Z(n6165) );
  XOR \SUBBYTES[1].a/U5180  ( .A(\SUBBYTES[1].a/w913 ), .B(
        \SUBBYTES[1].a/w916 ), .Z(n6166) );
  XOR \SUBBYTES[1].a/U5179  ( .A(\SUBBYTES[1].a/w906 ), .B(
        \SUBBYTES[1].a/w909 ), .Z(n6167) );
  XOR \SUBBYTES[1].a/U5178  ( .A(\SUBBYTES[1].a/w881 ), .B(
        \SUBBYTES[1].a/w882 ), .Z(n6168) );
  XOR \SUBBYTES[1].a/U5177  ( .A(\SUBBYTES[1].a/w866 ), .B(
        \SUBBYTES[1].a/w869 ), .Z(n6169) );
  XOR \SUBBYTES[1].a/U5175  ( .A(n6965), .B(n6172), .Z(n6170) );
  XOR \SUBBYTES[1].a/U5174  ( .A(n6967), .B(n6966), .Z(n6171) );
  XOR \SUBBYTES[1].a/U5173  ( .A(\SUBBYTES[1].a/w874 ), .B(
        \SUBBYTES[1].a/w901 ), .Z(n6172) );
  XOR \SUBBYTES[1].a/U5171  ( .A(n6968), .B(n6175), .Z(n6173) );
  XOR \SUBBYTES[1].a/U5170  ( .A(\SUBBYTES[1].a/w907 ), .B(
        \SUBBYTES[1].a/w909 ), .Z(n6174) );
  XOR \SUBBYTES[1].a/U5169  ( .A(\SUBBYTES[1].a/w867 ), .B(
        \SUBBYTES[1].a/w899 ), .Z(n6175) );
  XOR \SUBBYTES[1].a/U5168  ( .A(\SUBBYTES[1].a/w699 ), .B(
        \SUBBYTES[1].a/w700 ), .Z(n6970) );
  XOR \SUBBYTES[1].a/U5167  ( .A(n6970), .B(n6176), .Z(n6969) );
  XOR \SUBBYTES[1].a/U5166  ( .A(\SUBBYTES[1].a/w692 ), .B(
        \SUBBYTES[1].a/w709 ), .Z(n6176) );
  XOR \SUBBYTES[1].a/U5164  ( .A(\SUBBYTES[1].a/w691 ), .B(
        \SUBBYTES[1].a/w706 ), .Z(n6177) );
  XOR \SUBBYTES[1].a/U5163  ( .A(n6970), .B(n6178), .Z(n7109) );
  XOR \SUBBYTES[1].a/U5162  ( .A(\SUBBYTES[1].a/w706 ), .B(
        \SUBBYTES[1].a/w707 ), .Z(n6178) );
  XOR \SUBBYTES[1].a/U5161  ( .A(\SUBBYTES[1].a/w668 ), .B(n6179), .Z(n6972)
         );
  XOR \SUBBYTES[1].a/U5160  ( .A(\SUBBYTES[1].a/w659 ), .B(
        \SUBBYTES[1].a/w660 ), .Z(n6179) );
  XOR \SUBBYTES[1].a/U5158  ( .A(\SUBBYTES[1].a/w670 ), .B(n7109), .Z(n6180)
         );
  XOR \SUBBYTES[1].a/U5157  ( .A(n6182), .B(n6181), .Z(n6973) );
  XOR \SUBBYTES[1].a/U5156  ( .A(n6184), .B(n6183), .Z(n6181) );
  XOR \SUBBYTES[1].a/U5155  ( .A(\SUBBYTES[1].a/w706 ), .B(
        \SUBBYTES[1].a/w707 ), .Z(n6182) );
  XOR \SUBBYTES[1].a/U5154  ( .A(\SUBBYTES[1].a/w670 ), .B(
        \SUBBYTES[1].a/w694 ), .Z(n6183) );
  XOR \SUBBYTES[1].a/U5153  ( .A(\SUBBYTES[1].a/w659 ), .B(
        \SUBBYTES[1].a/w668 ), .Z(n6184) );
  XOR \SUBBYTES[1].a/U5152  ( .A(\SUBBYTES[1].a/w691 ), .B(n6185), .Z(n6971)
         );
  XOR \SUBBYTES[1].a/U5151  ( .A(\SUBBYTES[1].a/w674 ), .B(
        \SUBBYTES[1].a/w677 ), .Z(n6185) );
  XOR \SUBBYTES[1].a/U5149  ( .A(\SUBBYTES[1].a/w662 ), .B(n6973), .Z(n6186)
         );
  XOR \SUBBYTES[1].a/U5147  ( .A(\SUBBYTES[1].a/w694 ), .B(
        \SUBBYTES[1].a/w707 ), .Z(n6187) );
  XOR \SUBBYTES[1].a/U5145  ( .A(n6191), .B(n6190), .Z(n6188) );
  XOR \SUBBYTES[1].a/U5144  ( .A(n6193), .B(n6192), .Z(n6189) );
  XOR \SUBBYTES[1].a/U5143  ( .A(\SUBBYTES[1].a/w706 ), .B(
        \SUBBYTES[1].a/w709 ), .Z(n6190) );
  XOR \SUBBYTES[1].a/U5142  ( .A(\SUBBYTES[1].a/w699 ), .B(
        \SUBBYTES[1].a/w702 ), .Z(n6191) );
  XOR \SUBBYTES[1].a/U5141  ( .A(\SUBBYTES[1].a/w674 ), .B(
        \SUBBYTES[1].a/w675 ), .Z(n6192) );
  XOR \SUBBYTES[1].a/U5140  ( .A(\SUBBYTES[1].a/w659 ), .B(
        \SUBBYTES[1].a/w662 ), .Z(n6193) );
  XOR \SUBBYTES[1].a/U5138  ( .A(n6970), .B(n6196), .Z(n6194) );
  XOR \SUBBYTES[1].a/U5137  ( .A(n6972), .B(n6971), .Z(n6195) );
  XOR \SUBBYTES[1].a/U5136  ( .A(\SUBBYTES[1].a/w667 ), .B(
        \SUBBYTES[1].a/w694 ), .Z(n6196) );
  XOR \SUBBYTES[1].a/U5134  ( .A(n6973), .B(n6199), .Z(n6197) );
  XOR \SUBBYTES[1].a/U5133  ( .A(\SUBBYTES[1].a/w700 ), .B(
        \SUBBYTES[1].a/w702 ), .Z(n6198) );
  XOR \SUBBYTES[1].a/U5132  ( .A(\SUBBYTES[1].a/w660 ), .B(
        \SUBBYTES[1].a/w692 ), .Z(n6199) );
  XOR \SUBBYTES[1].a/U5131  ( .A(\SUBBYTES[1].a/w492 ), .B(
        \SUBBYTES[1].a/w493 ), .Z(n6975) );
  XOR \SUBBYTES[1].a/U5130  ( .A(n6975), .B(n6200), .Z(n6974) );
  XOR \SUBBYTES[1].a/U5129  ( .A(\SUBBYTES[1].a/w485 ), .B(
        \SUBBYTES[1].a/w502 ), .Z(n6200) );
  XOR \SUBBYTES[1].a/U5127  ( .A(\SUBBYTES[1].a/w484 ), .B(
        \SUBBYTES[1].a/w499 ), .Z(n6201) );
  XOR \SUBBYTES[1].a/U5126  ( .A(n6975), .B(n6202), .Z(n7110) );
  XOR \SUBBYTES[1].a/U5125  ( .A(\SUBBYTES[1].a/w499 ), .B(
        \SUBBYTES[1].a/w500 ), .Z(n6202) );
  XOR \SUBBYTES[1].a/U5124  ( .A(\SUBBYTES[1].a/w461 ), .B(n6203), .Z(n6977)
         );
  XOR \SUBBYTES[1].a/U5123  ( .A(\SUBBYTES[1].a/w452 ), .B(
        \SUBBYTES[1].a/w453 ), .Z(n6203) );
  XOR \SUBBYTES[1].a/U5121  ( .A(\SUBBYTES[1].a/w463 ), .B(n7110), .Z(n6204)
         );
  XOR \SUBBYTES[1].a/U5120  ( .A(n6206), .B(n6205), .Z(n6978) );
  XOR \SUBBYTES[1].a/U5119  ( .A(n6208), .B(n6207), .Z(n6205) );
  XOR \SUBBYTES[1].a/U5118  ( .A(\SUBBYTES[1].a/w499 ), .B(
        \SUBBYTES[1].a/w500 ), .Z(n6206) );
  XOR \SUBBYTES[1].a/U5117  ( .A(\SUBBYTES[1].a/w463 ), .B(
        \SUBBYTES[1].a/w487 ), .Z(n6207) );
  XOR \SUBBYTES[1].a/U5116  ( .A(\SUBBYTES[1].a/w452 ), .B(
        \SUBBYTES[1].a/w461 ), .Z(n6208) );
  XOR \SUBBYTES[1].a/U5115  ( .A(\SUBBYTES[1].a/w484 ), .B(n6209), .Z(n6976)
         );
  XOR \SUBBYTES[1].a/U5114  ( .A(\SUBBYTES[1].a/w467 ), .B(
        \SUBBYTES[1].a/w470 ), .Z(n6209) );
  XOR \SUBBYTES[1].a/U5112  ( .A(\SUBBYTES[1].a/w455 ), .B(n6978), .Z(n6210)
         );
  XOR \SUBBYTES[1].a/U5110  ( .A(\SUBBYTES[1].a/w487 ), .B(
        \SUBBYTES[1].a/w500 ), .Z(n6211) );
  XOR \SUBBYTES[1].a/U5108  ( .A(n6215), .B(n6214), .Z(n6212) );
  XOR \SUBBYTES[1].a/U5107  ( .A(n6217), .B(n6216), .Z(n6213) );
  XOR \SUBBYTES[1].a/U5106  ( .A(\SUBBYTES[1].a/w499 ), .B(
        \SUBBYTES[1].a/w502 ), .Z(n6214) );
  XOR \SUBBYTES[1].a/U5105  ( .A(\SUBBYTES[1].a/w492 ), .B(
        \SUBBYTES[1].a/w495 ), .Z(n6215) );
  XOR \SUBBYTES[1].a/U5104  ( .A(\SUBBYTES[1].a/w467 ), .B(
        \SUBBYTES[1].a/w468 ), .Z(n6216) );
  XOR \SUBBYTES[1].a/U5103  ( .A(\SUBBYTES[1].a/w452 ), .B(
        \SUBBYTES[1].a/w455 ), .Z(n6217) );
  XOR \SUBBYTES[1].a/U5101  ( .A(n6975), .B(n6220), .Z(n6218) );
  XOR \SUBBYTES[1].a/U5100  ( .A(n6977), .B(n6976), .Z(n6219) );
  XOR \SUBBYTES[1].a/U5099  ( .A(\SUBBYTES[1].a/w460 ), .B(
        \SUBBYTES[1].a/w487 ), .Z(n6220) );
  XOR \SUBBYTES[1].a/U5097  ( .A(n6978), .B(n6223), .Z(n6221) );
  XOR \SUBBYTES[1].a/U5096  ( .A(\SUBBYTES[1].a/w493 ), .B(
        \SUBBYTES[1].a/w495 ), .Z(n6222) );
  XOR \SUBBYTES[1].a/U5095  ( .A(\SUBBYTES[1].a/w453 ), .B(
        \SUBBYTES[1].a/w485 ), .Z(n6223) );
  XOR \SUBBYTES[1].a/U5094  ( .A(\SUBBYTES[1].a/w285 ), .B(
        \SUBBYTES[1].a/w286 ), .Z(n6980) );
  XOR \SUBBYTES[1].a/U5093  ( .A(n6980), .B(n6224), .Z(n6979) );
  XOR \SUBBYTES[1].a/U5092  ( .A(\SUBBYTES[1].a/w278 ), .B(
        \SUBBYTES[1].a/w295 ), .Z(n6224) );
  XOR \SUBBYTES[1].a/U5090  ( .A(\SUBBYTES[1].a/w277 ), .B(
        \SUBBYTES[1].a/w292 ), .Z(n6225) );
  XOR \SUBBYTES[1].a/U5089  ( .A(n6980), .B(n6226), .Z(n7111) );
  XOR \SUBBYTES[1].a/U5088  ( .A(\SUBBYTES[1].a/w292 ), .B(
        \SUBBYTES[1].a/w293 ), .Z(n6226) );
  XOR \SUBBYTES[1].a/U5087  ( .A(\SUBBYTES[1].a/w254 ), .B(n6227), .Z(n6982)
         );
  XOR \SUBBYTES[1].a/U5086  ( .A(\SUBBYTES[1].a/w245 ), .B(
        \SUBBYTES[1].a/w246 ), .Z(n6227) );
  XOR \SUBBYTES[1].a/U5084  ( .A(\SUBBYTES[1].a/w256 ), .B(n7111), .Z(n6228)
         );
  XOR \SUBBYTES[1].a/U5083  ( .A(n6230), .B(n6229), .Z(n6983) );
  XOR \SUBBYTES[1].a/U5082  ( .A(n6232), .B(n6231), .Z(n6229) );
  XOR \SUBBYTES[1].a/U5081  ( .A(\SUBBYTES[1].a/w292 ), .B(
        \SUBBYTES[1].a/w293 ), .Z(n6230) );
  XOR \SUBBYTES[1].a/U5080  ( .A(\SUBBYTES[1].a/w256 ), .B(
        \SUBBYTES[1].a/w280 ), .Z(n6231) );
  XOR \SUBBYTES[1].a/U5079  ( .A(\SUBBYTES[1].a/w245 ), .B(
        \SUBBYTES[1].a/w254 ), .Z(n6232) );
  XOR \SUBBYTES[1].a/U5078  ( .A(\SUBBYTES[1].a/w277 ), .B(n6233), .Z(n6981)
         );
  XOR \SUBBYTES[1].a/U5077  ( .A(\SUBBYTES[1].a/w260 ), .B(
        \SUBBYTES[1].a/w263 ), .Z(n6233) );
  XOR \SUBBYTES[1].a/U5075  ( .A(\SUBBYTES[1].a/w248 ), .B(n6983), .Z(n6234)
         );
  XOR \SUBBYTES[1].a/U5073  ( .A(\SUBBYTES[1].a/w280 ), .B(
        \SUBBYTES[1].a/w293 ), .Z(n6235) );
  XOR \SUBBYTES[1].a/U5071  ( .A(n6239), .B(n6238), .Z(n6236) );
  XOR \SUBBYTES[1].a/U5070  ( .A(n6241), .B(n6240), .Z(n6237) );
  XOR \SUBBYTES[1].a/U5069  ( .A(\SUBBYTES[1].a/w292 ), .B(
        \SUBBYTES[1].a/w295 ), .Z(n6238) );
  XOR \SUBBYTES[1].a/U5068  ( .A(\SUBBYTES[1].a/w285 ), .B(
        \SUBBYTES[1].a/w288 ), .Z(n6239) );
  XOR \SUBBYTES[1].a/U5067  ( .A(\SUBBYTES[1].a/w260 ), .B(
        \SUBBYTES[1].a/w261 ), .Z(n6240) );
  XOR \SUBBYTES[1].a/U5066  ( .A(\SUBBYTES[1].a/w245 ), .B(
        \SUBBYTES[1].a/w248 ), .Z(n6241) );
  XOR \SUBBYTES[1].a/U5064  ( .A(n6980), .B(n6244), .Z(n6242) );
  XOR \SUBBYTES[1].a/U5063  ( .A(n6982), .B(n6981), .Z(n6243) );
  XOR \SUBBYTES[1].a/U5062  ( .A(\SUBBYTES[1].a/w253 ), .B(
        \SUBBYTES[1].a/w280 ), .Z(n6244) );
  XOR \SUBBYTES[1].a/U5060  ( .A(n6983), .B(n6247), .Z(n6245) );
  XOR \SUBBYTES[1].a/U5059  ( .A(\SUBBYTES[1].a/w286 ), .B(
        \SUBBYTES[1].a/w288 ), .Z(n6246) );
  XOR \SUBBYTES[1].a/U5058  ( .A(\SUBBYTES[1].a/w246 ), .B(
        \SUBBYTES[1].a/w278 ), .Z(n6247) );
  XOR \SUBBYTES[1].a/U5057  ( .A(\w1[1][1] ), .B(n6248), .Z(n6984) );
  XOR \SUBBYTES[1].a/U5056  ( .A(\w1[1][3] ), .B(\w1[1][2] ), .Z(n6248) );
  XOR \SUBBYTES[1].a/U5055  ( .A(\w1[1][6] ), .B(n6984), .Z(
        \SUBBYTES[1].a/w3378 ) );
  XOR \SUBBYTES[1].a/U5054  ( .A(\w1[1][0] ), .B(\SUBBYTES[1].a/w3378 ), .Z(
        \SUBBYTES[1].a/w3265 ) );
  XOR \SUBBYTES[1].a/U5053  ( .A(\w1[1][0] ), .B(n6249), .Z(
        \SUBBYTES[1].a/w3266 ) );
  XOR \SUBBYTES[1].a/U5052  ( .A(\w1[1][6] ), .B(\w1[1][5] ), .Z(n6249) );
  XOR \SUBBYTES[1].a/U5051  ( .A(\w1[1][5] ), .B(n6984), .Z(
        \SUBBYTES[1].a/w3396 ) );
  XOR \SUBBYTES[1].a/U5050  ( .A(n6251), .B(n6250), .Z(\SUBBYTES[1].a/w3389 )
         );
  XOR \SUBBYTES[1].a/U5049  ( .A(\w1[1][3] ), .B(\w1[1][1] ), .Z(n6250) );
  XOR \SUBBYTES[1].a/U5048  ( .A(\w1[1][7] ), .B(\w1[1][4] ), .Z(n6251) );
  XOR \SUBBYTES[1].a/U5047  ( .A(\w1[1][0] ), .B(\SUBBYTES[1].a/w3389 ), .Z(
        \SUBBYTES[1].a/w3268 ) );
  XOR \SUBBYTES[1].a/U5046  ( .A(n6253), .B(n6252), .Z(\SUBBYTES[1].a/w3376 )
         );
  XOR \SUBBYTES[1].a/U5045  ( .A(\SUBBYTES[1].a/w3337 ), .B(n972), .Z(n6252)
         );
  XOR \SUBBYTES[1].a/U5044  ( .A(\SUBBYTES[1].a/w3330 ), .B(
        \SUBBYTES[1].a/w3333 ), .Z(n6253) );
  XOR \SUBBYTES[1].a/U5043  ( .A(n6255), .B(n6254), .Z(\SUBBYTES[1].a/w3377 )
         );
  XOR \SUBBYTES[1].a/U5042  ( .A(\SUBBYTES[1].a/w3337 ), .B(n5863), .Z(n6254)
         );
  XOR \SUBBYTES[1].a/U5041  ( .A(\SUBBYTES[1].a/w3330 ), .B(n5862), .Z(n6255)
         );
  XOR \SUBBYTES[1].a/U5040  ( .A(\SUBBYTES[1].a/w3389 ), .B(n6256), .Z(
        \SUBBYTES[1].a/w3379 ) );
  XOR \SUBBYTES[1].a/U5039  ( .A(\w1[1][6] ), .B(\w1[1][5] ), .Z(n6256) );
  XOR \SUBBYTES[1].a/U5038  ( .A(n6258), .B(n6257), .Z(\SUBBYTES[1].a/w3380 )
         );
  XOR \SUBBYTES[1].a/U5037  ( .A(n5863), .B(n972), .Z(n6257) );
  XOR \SUBBYTES[1].a/U5036  ( .A(n5862), .B(\SUBBYTES[1].a/w3333 ), .Z(n6258)
         );
  XOR \SUBBYTES[1].a/U5035  ( .A(\w1[1][7] ), .B(\w1[1][2] ), .Z(n6990) );
  XOR \SUBBYTES[1].a/U5034  ( .A(n6990), .B(n6259), .Z(\SUBBYTES[1].a/w3381 )
         );
  XOR \SUBBYTES[1].a/U5033  ( .A(\w1[1][5] ), .B(\w1[1][4] ), .Z(n6259) );
  XOR \SUBBYTES[1].a/U5032  ( .A(\w1[1][7] ), .B(\SUBBYTES[1].a/w3266 ), .Z(
        \SUBBYTES[1].a/w3269 ) );
  XOR \SUBBYTES[1].a/U5031  ( .A(\w1[1][1] ), .B(\SUBBYTES[1].a/w3266 ), .Z(
        \SUBBYTES[1].a/w3270 ) );
  XOR \SUBBYTES[1].a/U5030  ( .A(\w1[1][4] ), .B(\SUBBYTES[1].a/w3266 ), .Z(
        \SUBBYTES[1].a/w3271 ) );
  XOR \SUBBYTES[1].a/U5029  ( .A(\SUBBYTES[1].a/w3270 ), .B(n6990), .Z(
        \SUBBYTES[1].a/w3272 ) );
  XOR \SUBBYTES[1].a/U5028  ( .A(n6990), .B(n6260), .Z(\SUBBYTES[1].a/w3357 )
         );
  XOR \SUBBYTES[1].a/U5027  ( .A(\w1[1][4] ), .B(\w1[1][1] ), .Z(n6260) );
  XOR \SUBBYTES[1].a/U5026  ( .A(n6262), .B(n6261), .Z(n6987) );
  XOR \SUBBYTES[1].a/U5025  ( .A(\w1[1][4] ), .B(n6263), .Z(n6261) );
  XOR \SUBBYTES[1].a/U5024  ( .A(\SUBBYTES[1].a/w3322 ), .B(\w1[1][6] ), .Z(
        n6262) );
  XOR \SUBBYTES[1].a/U5023  ( .A(\SUBBYTES[1].a/w3296 ), .B(
        \SUBBYTES[1].a/w3303 ), .Z(n6263) );
  XOR \SUBBYTES[1].a/U5022  ( .A(n6265), .B(n6264), .Z(n6985) );
  XOR \SUBBYTES[1].a/U5021  ( .A(\w1[1][1] ), .B(n6266), .Z(n6264) );
  XOR \SUBBYTES[1].a/U5020  ( .A(\SUBBYTES[1].a/w3321 ), .B(\w1[1][5] ), .Z(
        n6265) );
  XOR \SUBBYTES[1].a/U5019  ( .A(\SUBBYTES[1].a/w3297 ), .B(
        \SUBBYTES[1].a/w3304 ), .Z(n6266) );
  XOR \SUBBYTES[1].a/U5018  ( .A(n6987), .B(n6985), .Z(\SUBBYTES[1].a/w3327 )
         );
  XOR \SUBBYTES[1].a/U5017  ( .A(\w1[1][5] ), .B(n6267), .Z(n6988) );
  XOR \SUBBYTES[1].a/U5016  ( .A(\SUBBYTES[1].a/w3289 ), .B(
        \SUBBYTES[1].a/w3299 ), .Z(n6267) );
  XOR \SUBBYTES[1].a/U5015  ( .A(n6269), .B(n6268), .Z(\SUBBYTES[1].a/w3314 )
         );
  XOR \SUBBYTES[1].a/U5014  ( .A(n6988), .B(n6270), .Z(n6268) );
  XOR \SUBBYTES[1].a/U5013  ( .A(\w1[1][4] ), .B(\SUBBYTES[1].a/w3378 ), .Z(
        n6269) );
  XOR \SUBBYTES[1].a/U5012  ( .A(\SUBBYTES[1].a/w3291 ), .B(
        \SUBBYTES[1].a/w3296 ), .Z(n6270) );
  XOR \SUBBYTES[1].a/U5011  ( .A(n6272), .B(n6271), .Z(n6986) );
  XOR \SUBBYTES[1].a/U5010  ( .A(\SUBBYTES[1].a/w3324 ), .B(\w1[1][7] ), .Z(
        n6271) );
  XOR \SUBBYTES[1].a/U5009  ( .A(\SUBBYTES[1].a/w3299 ), .B(
        \SUBBYTES[1].a/w3306 ), .Z(n6272) );
  XOR \SUBBYTES[1].a/U5008  ( .A(n6985), .B(n6986), .Z(\SUBBYTES[1].a/w3326 )
         );
  XOR \SUBBYTES[1].a/U5007  ( .A(\w1[1][3] ), .B(n6273), .Z(n6989) );
  XOR \SUBBYTES[1].a/U5006  ( .A(\SUBBYTES[1].a/w3288 ), .B(
        \SUBBYTES[1].a/w3291 ), .Z(n6273) );
  XOR \SUBBYTES[1].a/U5005  ( .A(n6275), .B(n6274), .Z(\SUBBYTES[1].a/w3315 )
         );
  XOR \SUBBYTES[1].a/U5004  ( .A(n6989), .B(n6276), .Z(n6274) );
  XOR \SUBBYTES[1].a/U5003  ( .A(\w1[1][6] ), .B(\SUBBYTES[1].a/w3357 ), .Z(
        n6275) );
  XOR \SUBBYTES[1].a/U5002  ( .A(\SUBBYTES[1].a/w3296 ), .B(
        \SUBBYTES[1].a/w3297 ), .Z(n6276) );
  XOR \SUBBYTES[1].a/U5001  ( .A(n6987), .B(n6986), .Z(\SUBBYTES[1].a/w3335 )
         );
  XOR \SUBBYTES[1].a/U5000  ( .A(n6278), .B(n6277), .Z(\SUBBYTES[1].a/w3336 )
         );
  XOR \SUBBYTES[1].a/U4999  ( .A(\w1[1][7] ), .B(n6988), .Z(n6277) );
  XOR \SUBBYTES[1].a/U4998  ( .A(\SUBBYTES[1].a/w3288 ), .B(
        \SUBBYTES[1].a/w3297 ), .Z(n6278) );
  XOR \SUBBYTES[1].a/U4997  ( .A(n6280), .B(n6279), .Z(\SUBBYTES[1].a/w3312 )
         );
  XOR \SUBBYTES[1].a/U4996  ( .A(n6282), .B(n6281), .Z(n6279) );
  XOR \SUBBYTES[1].a/U4995  ( .A(\w1[1][7] ), .B(\SUBBYTES[1].a/w3396 ), .Z(
        n6280) );
  XOR \SUBBYTES[1].a/U4994  ( .A(\SUBBYTES[1].a/w3303 ), .B(
        \SUBBYTES[1].a/w3306 ), .Z(n6281) );
  XOR \SUBBYTES[1].a/U4993  ( .A(\SUBBYTES[1].a/w3289 ), .B(
        \SUBBYTES[1].a/w3291 ), .Z(n6282) );
  XOR \SUBBYTES[1].a/U4992  ( .A(n6284), .B(n6283), .Z(\SUBBYTES[1].a/w3313 )
         );
  XOR \SUBBYTES[1].a/U4991  ( .A(n6989), .B(n6285), .Z(n6283) );
  XOR \SUBBYTES[1].a/U4990  ( .A(\w1[1][5] ), .B(n6990), .Z(n6284) );
  XOR \SUBBYTES[1].a/U4989  ( .A(\SUBBYTES[1].a/w3303 ), .B(
        \SUBBYTES[1].a/w3304 ), .Z(n6285) );
  XOR \SUBBYTES[1].a/U4988  ( .A(n6287), .B(n6286), .Z(\SUBBYTES[1].a/w3329 )
         );
  XOR \SUBBYTES[1].a/U4987  ( .A(\w1[1][1] ), .B(n6288), .Z(n6286) );
  XOR \SUBBYTES[1].a/U4986  ( .A(\SUBBYTES[1].a/w3304 ), .B(
        \SUBBYTES[1].a/w3306 ), .Z(n6287) );
  XOR \SUBBYTES[1].a/U4985  ( .A(\SUBBYTES[1].a/w3288 ), .B(
        \SUBBYTES[1].a/w3289 ), .Z(n6288) );
  XOR \SUBBYTES[1].a/U4984  ( .A(\w1[1][9] ), .B(n6289), .Z(n6991) );
  XOR \SUBBYTES[1].a/U4983  ( .A(\w1[1][11] ), .B(\w1[1][10] ), .Z(n6289) );
  XOR \SUBBYTES[1].a/U4982  ( .A(\w1[1][14] ), .B(n6991), .Z(
        \SUBBYTES[1].a/w3171 ) );
  XOR \SUBBYTES[1].a/U4981  ( .A(\w1[1][8] ), .B(\SUBBYTES[1].a/w3171 ), .Z(
        \SUBBYTES[1].a/w3058 ) );
  XOR \SUBBYTES[1].a/U4980  ( .A(\w1[1][8] ), .B(n6290), .Z(
        \SUBBYTES[1].a/w3059 ) );
  XOR \SUBBYTES[1].a/U4979  ( .A(\w1[1][14] ), .B(\w1[1][13] ), .Z(n6290) );
  XOR \SUBBYTES[1].a/U4978  ( .A(\w1[1][13] ), .B(n6991), .Z(
        \SUBBYTES[1].a/w3189 ) );
  XOR \SUBBYTES[1].a/U4977  ( .A(n6292), .B(n6291), .Z(\SUBBYTES[1].a/w3182 )
         );
  XOR \SUBBYTES[1].a/U4976  ( .A(\w1[1][11] ), .B(\w1[1][9] ), .Z(n6291) );
  XOR \SUBBYTES[1].a/U4975  ( .A(\w1[1][15] ), .B(\w1[1][12] ), .Z(n6292) );
  XOR \SUBBYTES[1].a/U4974  ( .A(\w1[1][8] ), .B(\SUBBYTES[1].a/w3182 ), .Z(
        \SUBBYTES[1].a/w3061 ) );
  XOR \SUBBYTES[1].a/U4973  ( .A(n6294), .B(n6293), .Z(\SUBBYTES[1].a/w3169 )
         );
  XOR \SUBBYTES[1].a/U4972  ( .A(\SUBBYTES[1].a/w3130 ), .B(n971), .Z(n6293)
         );
  XOR \SUBBYTES[1].a/U4971  ( .A(\SUBBYTES[1].a/w3123 ), .B(
        \SUBBYTES[1].a/w3126 ), .Z(n6294) );
  XOR \SUBBYTES[1].a/U4970  ( .A(n6296), .B(n6295), .Z(\SUBBYTES[1].a/w3170 )
         );
  XOR \SUBBYTES[1].a/U4969  ( .A(\SUBBYTES[1].a/w3130 ), .B(n5861), .Z(n6295)
         );
  XOR \SUBBYTES[1].a/U4968  ( .A(\SUBBYTES[1].a/w3123 ), .B(n5860), .Z(n6296)
         );
  XOR \SUBBYTES[1].a/U4967  ( .A(\SUBBYTES[1].a/w3182 ), .B(n6297), .Z(
        \SUBBYTES[1].a/w3172 ) );
  XOR \SUBBYTES[1].a/U4966  ( .A(\w1[1][14] ), .B(\w1[1][13] ), .Z(n6297) );
  XOR \SUBBYTES[1].a/U4965  ( .A(n6299), .B(n6298), .Z(\SUBBYTES[1].a/w3173 )
         );
  XOR \SUBBYTES[1].a/U4964  ( .A(n5861), .B(n971), .Z(n6298) );
  XOR \SUBBYTES[1].a/U4963  ( .A(n5860), .B(\SUBBYTES[1].a/w3126 ), .Z(n6299)
         );
  XOR \SUBBYTES[1].a/U4962  ( .A(\w1[1][15] ), .B(\w1[1][10] ), .Z(n6997) );
  XOR \SUBBYTES[1].a/U4961  ( .A(n6997), .B(n6300), .Z(\SUBBYTES[1].a/w3174 )
         );
  XOR \SUBBYTES[1].a/U4960  ( .A(\w1[1][13] ), .B(\w1[1][12] ), .Z(n6300) );
  XOR \SUBBYTES[1].a/U4959  ( .A(\w1[1][15] ), .B(\SUBBYTES[1].a/w3059 ), .Z(
        \SUBBYTES[1].a/w3062 ) );
  XOR \SUBBYTES[1].a/U4958  ( .A(\w1[1][9] ), .B(\SUBBYTES[1].a/w3059 ), .Z(
        \SUBBYTES[1].a/w3063 ) );
  XOR \SUBBYTES[1].a/U4957  ( .A(\w1[1][12] ), .B(\SUBBYTES[1].a/w3059 ), .Z(
        \SUBBYTES[1].a/w3064 ) );
  XOR \SUBBYTES[1].a/U4956  ( .A(\SUBBYTES[1].a/w3063 ), .B(n6997), .Z(
        \SUBBYTES[1].a/w3065 ) );
  XOR \SUBBYTES[1].a/U4955  ( .A(n6997), .B(n6301), .Z(\SUBBYTES[1].a/w3150 )
         );
  XOR \SUBBYTES[1].a/U4954  ( .A(\w1[1][12] ), .B(\w1[1][9] ), .Z(n6301) );
  XOR \SUBBYTES[1].a/U4953  ( .A(n6303), .B(n6302), .Z(n6994) );
  XOR \SUBBYTES[1].a/U4952  ( .A(\w1[1][12] ), .B(n6304), .Z(n6302) );
  XOR \SUBBYTES[1].a/U4951  ( .A(\SUBBYTES[1].a/w3115 ), .B(\w1[1][14] ), .Z(
        n6303) );
  XOR \SUBBYTES[1].a/U4950  ( .A(\SUBBYTES[1].a/w3089 ), .B(
        \SUBBYTES[1].a/w3096 ), .Z(n6304) );
  XOR \SUBBYTES[1].a/U4949  ( .A(n6306), .B(n6305), .Z(n6992) );
  XOR \SUBBYTES[1].a/U4948  ( .A(\w1[1][9] ), .B(n6307), .Z(n6305) );
  XOR \SUBBYTES[1].a/U4947  ( .A(\SUBBYTES[1].a/w3114 ), .B(\w1[1][13] ), .Z(
        n6306) );
  XOR \SUBBYTES[1].a/U4946  ( .A(\SUBBYTES[1].a/w3090 ), .B(
        \SUBBYTES[1].a/w3097 ), .Z(n6307) );
  XOR \SUBBYTES[1].a/U4945  ( .A(n6994), .B(n6992), .Z(\SUBBYTES[1].a/w3120 )
         );
  XOR \SUBBYTES[1].a/U4944  ( .A(\w1[1][13] ), .B(n6308), .Z(n6995) );
  XOR \SUBBYTES[1].a/U4943  ( .A(\SUBBYTES[1].a/w3082 ), .B(
        \SUBBYTES[1].a/w3092 ), .Z(n6308) );
  XOR \SUBBYTES[1].a/U4942  ( .A(n6310), .B(n6309), .Z(\SUBBYTES[1].a/w3107 )
         );
  XOR \SUBBYTES[1].a/U4941  ( .A(n6995), .B(n6311), .Z(n6309) );
  XOR \SUBBYTES[1].a/U4940  ( .A(\w1[1][12] ), .B(\SUBBYTES[1].a/w3171 ), .Z(
        n6310) );
  XOR \SUBBYTES[1].a/U4939  ( .A(\SUBBYTES[1].a/w3084 ), .B(
        \SUBBYTES[1].a/w3089 ), .Z(n6311) );
  XOR \SUBBYTES[1].a/U4938  ( .A(n6313), .B(n6312), .Z(n6993) );
  XOR \SUBBYTES[1].a/U4937  ( .A(\SUBBYTES[1].a/w3117 ), .B(\w1[1][15] ), .Z(
        n6312) );
  XOR \SUBBYTES[1].a/U4936  ( .A(\SUBBYTES[1].a/w3092 ), .B(
        \SUBBYTES[1].a/w3099 ), .Z(n6313) );
  XOR \SUBBYTES[1].a/U4935  ( .A(n6992), .B(n6993), .Z(\SUBBYTES[1].a/w3119 )
         );
  XOR \SUBBYTES[1].a/U4934  ( .A(\w1[1][11] ), .B(n6314), .Z(n6996) );
  XOR \SUBBYTES[1].a/U4933  ( .A(\SUBBYTES[1].a/w3081 ), .B(
        \SUBBYTES[1].a/w3084 ), .Z(n6314) );
  XOR \SUBBYTES[1].a/U4932  ( .A(n6316), .B(n6315), .Z(\SUBBYTES[1].a/w3108 )
         );
  XOR \SUBBYTES[1].a/U4931  ( .A(n6996), .B(n6317), .Z(n6315) );
  XOR \SUBBYTES[1].a/U4930  ( .A(\w1[1][14] ), .B(\SUBBYTES[1].a/w3150 ), .Z(
        n6316) );
  XOR \SUBBYTES[1].a/U4929  ( .A(\SUBBYTES[1].a/w3089 ), .B(
        \SUBBYTES[1].a/w3090 ), .Z(n6317) );
  XOR \SUBBYTES[1].a/U4928  ( .A(n6994), .B(n6993), .Z(\SUBBYTES[1].a/w3128 )
         );
  XOR \SUBBYTES[1].a/U4927  ( .A(n6319), .B(n6318), .Z(\SUBBYTES[1].a/w3129 )
         );
  XOR \SUBBYTES[1].a/U4926  ( .A(\w1[1][15] ), .B(n6995), .Z(n6318) );
  XOR \SUBBYTES[1].a/U4925  ( .A(\SUBBYTES[1].a/w3081 ), .B(
        \SUBBYTES[1].a/w3090 ), .Z(n6319) );
  XOR \SUBBYTES[1].a/U4924  ( .A(n6321), .B(n6320), .Z(\SUBBYTES[1].a/w3105 )
         );
  XOR \SUBBYTES[1].a/U4923  ( .A(n6323), .B(n6322), .Z(n6320) );
  XOR \SUBBYTES[1].a/U4922  ( .A(\w1[1][15] ), .B(\SUBBYTES[1].a/w3189 ), .Z(
        n6321) );
  XOR \SUBBYTES[1].a/U4921  ( .A(\SUBBYTES[1].a/w3096 ), .B(
        \SUBBYTES[1].a/w3099 ), .Z(n6322) );
  XOR \SUBBYTES[1].a/U4920  ( .A(\SUBBYTES[1].a/w3082 ), .B(
        \SUBBYTES[1].a/w3084 ), .Z(n6323) );
  XOR \SUBBYTES[1].a/U4919  ( .A(n6325), .B(n6324), .Z(\SUBBYTES[1].a/w3106 )
         );
  XOR \SUBBYTES[1].a/U4918  ( .A(n6996), .B(n6326), .Z(n6324) );
  XOR \SUBBYTES[1].a/U4917  ( .A(\w1[1][13] ), .B(n6997), .Z(n6325) );
  XOR \SUBBYTES[1].a/U4916  ( .A(\SUBBYTES[1].a/w3096 ), .B(
        \SUBBYTES[1].a/w3097 ), .Z(n6326) );
  XOR \SUBBYTES[1].a/U4915  ( .A(n6328), .B(n6327), .Z(\SUBBYTES[1].a/w3122 )
         );
  XOR \SUBBYTES[1].a/U4914  ( .A(\w1[1][9] ), .B(n6329), .Z(n6327) );
  XOR \SUBBYTES[1].a/U4913  ( .A(\SUBBYTES[1].a/w3097 ), .B(
        \SUBBYTES[1].a/w3099 ), .Z(n6328) );
  XOR \SUBBYTES[1].a/U4912  ( .A(\SUBBYTES[1].a/w3081 ), .B(
        \SUBBYTES[1].a/w3082 ), .Z(n6329) );
  XOR \SUBBYTES[1].a/U4911  ( .A(\w1[1][17] ), .B(n6330), .Z(n6998) );
  XOR \SUBBYTES[1].a/U4910  ( .A(\w1[1][19] ), .B(\w1[1][18] ), .Z(n6330) );
  XOR \SUBBYTES[1].a/U4909  ( .A(\w1[1][22] ), .B(n6998), .Z(
        \SUBBYTES[1].a/w2964 ) );
  XOR \SUBBYTES[1].a/U4908  ( .A(\w1[1][16] ), .B(\SUBBYTES[1].a/w2964 ), .Z(
        \SUBBYTES[1].a/w2851 ) );
  XOR \SUBBYTES[1].a/U4907  ( .A(\w1[1][16] ), .B(n6331), .Z(
        \SUBBYTES[1].a/w2852 ) );
  XOR \SUBBYTES[1].a/U4906  ( .A(\w1[1][22] ), .B(\w1[1][21] ), .Z(n6331) );
  XOR \SUBBYTES[1].a/U4905  ( .A(\w1[1][21] ), .B(n6998), .Z(
        \SUBBYTES[1].a/w2982 ) );
  XOR \SUBBYTES[1].a/U4904  ( .A(n6333), .B(n6332), .Z(\SUBBYTES[1].a/w2975 )
         );
  XOR \SUBBYTES[1].a/U4903  ( .A(\w1[1][19] ), .B(\w1[1][17] ), .Z(n6332) );
  XOR \SUBBYTES[1].a/U4902  ( .A(\w1[1][23] ), .B(\w1[1][20] ), .Z(n6333) );
  XOR \SUBBYTES[1].a/U4901  ( .A(\w1[1][16] ), .B(\SUBBYTES[1].a/w2975 ), .Z(
        \SUBBYTES[1].a/w2854 ) );
  XOR \SUBBYTES[1].a/U4900  ( .A(n6335), .B(n6334), .Z(\SUBBYTES[1].a/w2962 )
         );
  XOR \SUBBYTES[1].a/U4899  ( .A(\SUBBYTES[1].a/w2923 ), .B(n970), .Z(n6334)
         );
  XOR \SUBBYTES[1].a/U4898  ( .A(\SUBBYTES[1].a/w2916 ), .B(
        \SUBBYTES[1].a/w2919 ), .Z(n6335) );
  XOR \SUBBYTES[1].a/U4897  ( .A(n6337), .B(n6336), .Z(\SUBBYTES[1].a/w2963 )
         );
  XOR \SUBBYTES[1].a/U4896  ( .A(\SUBBYTES[1].a/w2923 ), .B(n5859), .Z(n6336)
         );
  XOR \SUBBYTES[1].a/U4895  ( .A(\SUBBYTES[1].a/w2916 ), .B(n5858), .Z(n6337)
         );
  XOR \SUBBYTES[1].a/U4894  ( .A(\SUBBYTES[1].a/w2975 ), .B(n6338), .Z(
        \SUBBYTES[1].a/w2965 ) );
  XOR \SUBBYTES[1].a/U4893  ( .A(\w1[1][22] ), .B(\w1[1][21] ), .Z(n6338) );
  XOR \SUBBYTES[1].a/U4892  ( .A(n6340), .B(n6339), .Z(\SUBBYTES[1].a/w2966 )
         );
  XOR \SUBBYTES[1].a/U4891  ( .A(n5859), .B(n970), .Z(n6339) );
  XOR \SUBBYTES[1].a/U4890  ( .A(n5858), .B(\SUBBYTES[1].a/w2919 ), .Z(n6340)
         );
  XOR \SUBBYTES[1].a/U4889  ( .A(\w1[1][23] ), .B(\w1[1][18] ), .Z(n7004) );
  XOR \SUBBYTES[1].a/U4888  ( .A(n7004), .B(n6341), .Z(\SUBBYTES[1].a/w2967 )
         );
  XOR \SUBBYTES[1].a/U4887  ( .A(\w1[1][21] ), .B(\w1[1][20] ), .Z(n6341) );
  XOR \SUBBYTES[1].a/U4886  ( .A(\w1[1][23] ), .B(\SUBBYTES[1].a/w2852 ), .Z(
        \SUBBYTES[1].a/w2855 ) );
  XOR \SUBBYTES[1].a/U4885  ( .A(\w1[1][17] ), .B(\SUBBYTES[1].a/w2852 ), .Z(
        \SUBBYTES[1].a/w2856 ) );
  XOR \SUBBYTES[1].a/U4884  ( .A(\w1[1][20] ), .B(\SUBBYTES[1].a/w2852 ), .Z(
        \SUBBYTES[1].a/w2857 ) );
  XOR \SUBBYTES[1].a/U4883  ( .A(\SUBBYTES[1].a/w2856 ), .B(n7004), .Z(
        \SUBBYTES[1].a/w2858 ) );
  XOR \SUBBYTES[1].a/U4882  ( .A(n7004), .B(n6342), .Z(\SUBBYTES[1].a/w2943 )
         );
  XOR \SUBBYTES[1].a/U4881  ( .A(\w1[1][20] ), .B(\w1[1][17] ), .Z(n6342) );
  XOR \SUBBYTES[1].a/U4880  ( .A(n6344), .B(n6343), .Z(n7001) );
  XOR \SUBBYTES[1].a/U4879  ( .A(\w1[1][20] ), .B(n6345), .Z(n6343) );
  XOR \SUBBYTES[1].a/U4878  ( .A(\SUBBYTES[1].a/w2908 ), .B(\w1[1][22] ), .Z(
        n6344) );
  XOR \SUBBYTES[1].a/U4877  ( .A(\SUBBYTES[1].a/w2882 ), .B(
        \SUBBYTES[1].a/w2889 ), .Z(n6345) );
  XOR \SUBBYTES[1].a/U4876  ( .A(n6347), .B(n6346), .Z(n6999) );
  XOR \SUBBYTES[1].a/U4875  ( .A(\w1[1][17] ), .B(n6348), .Z(n6346) );
  XOR \SUBBYTES[1].a/U4874  ( .A(\SUBBYTES[1].a/w2907 ), .B(\w1[1][21] ), .Z(
        n6347) );
  XOR \SUBBYTES[1].a/U4873  ( .A(\SUBBYTES[1].a/w2883 ), .B(
        \SUBBYTES[1].a/w2890 ), .Z(n6348) );
  XOR \SUBBYTES[1].a/U4872  ( .A(n7001), .B(n6999), .Z(\SUBBYTES[1].a/w2913 )
         );
  XOR \SUBBYTES[1].a/U4871  ( .A(\w1[1][21] ), .B(n6349), .Z(n7002) );
  XOR \SUBBYTES[1].a/U4870  ( .A(\SUBBYTES[1].a/w2875 ), .B(
        \SUBBYTES[1].a/w2885 ), .Z(n6349) );
  XOR \SUBBYTES[1].a/U4869  ( .A(n6351), .B(n6350), .Z(\SUBBYTES[1].a/w2900 )
         );
  XOR \SUBBYTES[1].a/U4868  ( .A(n7002), .B(n6352), .Z(n6350) );
  XOR \SUBBYTES[1].a/U4867  ( .A(\w1[1][20] ), .B(\SUBBYTES[1].a/w2964 ), .Z(
        n6351) );
  XOR \SUBBYTES[1].a/U4866  ( .A(\SUBBYTES[1].a/w2877 ), .B(
        \SUBBYTES[1].a/w2882 ), .Z(n6352) );
  XOR \SUBBYTES[1].a/U4865  ( .A(n6354), .B(n6353), .Z(n7000) );
  XOR \SUBBYTES[1].a/U4864  ( .A(\SUBBYTES[1].a/w2910 ), .B(\w1[1][23] ), .Z(
        n6353) );
  XOR \SUBBYTES[1].a/U4863  ( .A(\SUBBYTES[1].a/w2885 ), .B(
        \SUBBYTES[1].a/w2892 ), .Z(n6354) );
  XOR \SUBBYTES[1].a/U4862  ( .A(n6999), .B(n7000), .Z(\SUBBYTES[1].a/w2912 )
         );
  XOR \SUBBYTES[1].a/U4861  ( .A(\w1[1][19] ), .B(n6355), .Z(n7003) );
  XOR \SUBBYTES[1].a/U4860  ( .A(\SUBBYTES[1].a/w2874 ), .B(
        \SUBBYTES[1].a/w2877 ), .Z(n6355) );
  XOR \SUBBYTES[1].a/U4859  ( .A(n6357), .B(n6356), .Z(\SUBBYTES[1].a/w2901 )
         );
  XOR \SUBBYTES[1].a/U4858  ( .A(n7003), .B(n6358), .Z(n6356) );
  XOR \SUBBYTES[1].a/U4857  ( .A(\w1[1][22] ), .B(\SUBBYTES[1].a/w2943 ), .Z(
        n6357) );
  XOR \SUBBYTES[1].a/U4856  ( .A(\SUBBYTES[1].a/w2882 ), .B(
        \SUBBYTES[1].a/w2883 ), .Z(n6358) );
  XOR \SUBBYTES[1].a/U4855  ( .A(n7001), .B(n7000), .Z(\SUBBYTES[1].a/w2921 )
         );
  XOR \SUBBYTES[1].a/U4854  ( .A(n6360), .B(n6359), .Z(\SUBBYTES[1].a/w2922 )
         );
  XOR \SUBBYTES[1].a/U4853  ( .A(\w1[1][23] ), .B(n7002), .Z(n6359) );
  XOR \SUBBYTES[1].a/U4852  ( .A(\SUBBYTES[1].a/w2874 ), .B(
        \SUBBYTES[1].a/w2883 ), .Z(n6360) );
  XOR \SUBBYTES[1].a/U4851  ( .A(n6362), .B(n6361), .Z(\SUBBYTES[1].a/w2898 )
         );
  XOR \SUBBYTES[1].a/U4850  ( .A(n6364), .B(n6363), .Z(n6361) );
  XOR \SUBBYTES[1].a/U4849  ( .A(\w1[1][23] ), .B(\SUBBYTES[1].a/w2982 ), .Z(
        n6362) );
  XOR \SUBBYTES[1].a/U4848  ( .A(\SUBBYTES[1].a/w2889 ), .B(
        \SUBBYTES[1].a/w2892 ), .Z(n6363) );
  XOR \SUBBYTES[1].a/U4847  ( .A(\SUBBYTES[1].a/w2875 ), .B(
        \SUBBYTES[1].a/w2877 ), .Z(n6364) );
  XOR \SUBBYTES[1].a/U4846  ( .A(n6366), .B(n6365), .Z(\SUBBYTES[1].a/w2899 )
         );
  XOR \SUBBYTES[1].a/U4845  ( .A(n7003), .B(n6367), .Z(n6365) );
  XOR \SUBBYTES[1].a/U4844  ( .A(\w1[1][21] ), .B(n7004), .Z(n6366) );
  XOR \SUBBYTES[1].a/U4843  ( .A(\SUBBYTES[1].a/w2889 ), .B(
        \SUBBYTES[1].a/w2890 ), .Z(n6367) );
  XOR \SUBBYTES[1].a/U4842  ( .A(n6369), .B(n6368), .Z(\SUBBYTES[1].a/w2915 )
         );
  XOR \SUBBYTES[1].a/U4841  ( .A(\w1[1][17] ), .B(n6370), .Z(n6368) );
  XOR \SUBBYTES[1].a/U4840  ( .A(\SUBBYTES[1].a/w2890 ), .B(
        \SUBBYTES[1].a/w2892 ), .Z(n6369) );
  XOR \SUBBYTES[1].a/U4839  ( .A(\SUBBYTES[1].a/w2874 ), .B(
        \SUBBYTES[1].a/w2875 ), .Z(n6370) );
  XOR \SUBBYTES[1].a/U4838  ( .A(\w1[1][25] ), .B(n6371), .Z(n7005) );
  XOR \SUBBYTES[1].a/U4837  ( .A(\w1[1][27] ), .B(\w1[1][26] ), .Z(n6371) );
  XOR \SUBBYTES[1].a/U4836  ( .A(\w1[1][30] ), .B(n7005), .Z(
        \SUBBYTES[1].a/w2757 ) );
  XOR \SUBBYTES[1].a/U4835  ( .A(\w1[1][24] ), .B(\SUBBYTES[1].a/w2757 ), .Z(
        \SUBBYTES[1].a/w2644 ) );
  XOR \SUBBYTES[1].a/U4834  ( .A(\w1[1][24] ), .B(n6372), .Z(
        \SUBBYTES[1].a/w2645 ) );
  XOR \SUBBYTES[1].a/U4833  ( .A(\w1[1][30] ), .B(\w1[1][29] ), .Z(n6372) );
  XOR \SUBBYTES[1].a/U4832  ( .A(\w1[1][29] ), .B(n7005), .Z(
        \SUBBYTES[1].a/w2775 ) );
  XOR \SUBBYTES[1].a/U4831  ( .A(n6374), .B(n6373), .Z(\SUBBYTES[1].a/w2768 )
         );
  XOR \SUBBYTES[1].a/U4830  ( .A(\w1[1][27] ), .B(\w1[1][25] ), .Z(n6373) );
  XOR \SUBBYTES[1].a/U4829  ( .A(\w1[1][31] ), .B(\w1[1][28] ), .Z(n6374) );
  XOR \SUBBYTES[1].a/U4828  ( .A(\w1[1][24] ), .B(\SUBBYTES[1].a/w2768 ), .Z(
        \SUBBYTES[1].a/w2647 ) );
  XOR \SUBBYTES[1].a/U4827  ( .A(n6376), .B(n6375), .Z(\SUBBYTES[1].a/w2755 )
         );
  XOR \SUBBYTES[1].a/U4826  ( .A(\SUBBYTES[1].a/w2716 ), .B(n969), .Z(n6375)
         );
  XOR \SUBBYTES[1].a/U4825  ( .A(\SUBBYTES[1].a/w2709 ), .B(
        \SUBBYTES[1].a/w2712 ), .Z(n6376) );
  XOR \SUBBYTES[1].a/U4824  ( .A(n6378), .B(n6377), .Z(\SUBBYTES[1].a/w2756 )
         );
  XOR \SUBBYTES[1].a/U4823  ( .A(\SUBBYTES[1].a/w2716 ), .B(n5857), .Z(n6377)
         );
  XOR \SUBBYTES[1].a/U4822  ( .A(\SUBBYTES[1].a/w2709 ), .B(n5856), .Z(n6378)
         );
  XOR \SUBBYTES[1].a/U4821  ( .A(\SUBBYTES[1].a/w2768 ), .B(n6379), .Z(
        \SUBBYTES[1].a/w2758 ) );
  XOR \SUBBYTES[1].a/U4820  ( .A(\w1[1][30] ), .B(\w1[1][29] ), .Z(n6379) );
  XOR \SUBBYTES[1].a/U4819  ( .A(n6381), .B(n6380), .Z(\SUBBYTES[1].a/w2759 )
         );
  XOR \SUBBYTES[1].a/U4818  ( .A(n5857), .B(n969), .Z(n6380) );
  XOR \SUBBYTES[1].a/U4817  ( .A(n5856), .B(\SUBBYTES[1].a/w2712 ), .Z(n6381)
         );
  XOR \SUBBYTES[1].a/U4816  ( .A(\w1[1][31] ), .B(\w1[1][26] ), .Z(n7011) );
  XOR \SUBBYTES[1].a/U4815  ( .A(n7011), .B(n6382), .Z(\SUBBYTES[1].a/w2760 )
         );
  XOR \SUBBYTES[1].a/U4814  ( .A(\w1[1][29] ), .B(\w1[1][28] ), .Z(n6382) );
  XOR \SUBBYTES[1].a/U4813  ( .A(\w1[1][31] ), .B(\SUBBYTES[1].a/w2645 ), .Z(
        \SUBBYTES[1].a/w2648 ) );
  XOR \SUBBYTES[1].a/U4812  ( .A(\w1[1][25] ), .B(\SUBBYTES[1].a/w2645 ), .Z(
        \SUBBYTES[1].a/w2649 ) );
  XOR \SUBBYTES[1].a/U4811  ( .A(\w1[1][28] ), .B(\SUBBYTES[1].a/w2645 ), .Z(
        \SUBBYTES[1].a/w2650 ) );
  XOR \SUBBYTES[1].a/U4810  ( .A(\SUBBYTES[1].a/w2649 ), .B(n7011), .Z(
        \SUBBYTES[1].a/w2651 ) );
  XOR \SUBBYTES[1].a/U4809  ( .A(n7011), .B(n6383), .Z(\SUBBYTES[1].a/w2736 )
         );
  XOR \SUBBYTES[1].a/U4808  ( .A(\w1[1][28] ), .B(\w1[1][25] ), .Z(n6383) );
  XOR \SUBBYTES[1].a/U4807  ( .A(n6385), .B(n6384), .Z(n7008) );
  XOR \SUBBYTES[1].a/U4806  ( .A(\w1[1][28] ), .B(n6386), .Z(n6384) );
  XOR \SUBBYTES[1].a/U4805  ( .A(\SUBBYTES[1].a/w2701 ), .B(\w1[1][30] ), .Z(
        n6385) );
  XOR \SUBBYTES[1].a/U4804  ( .A(\SUBBYTES[1].a/w2675 ), .B(
        \SUBBYTES[1].a/w2682 ), .Z(n6386) );
  XOR \SUBBYTES[1].a/U4803  ( .A(n6388), .B(n6387), .Z(n7006) );
  XOR \SUBBYTES[1].a/U4802  ( .A(\w1[1][25] ), .B(n6389), .Z(n6387) );
  XOR \SUBBYTES[1].a/U4801  ( .A(\SUBBYTES[1].a/w2700 ), .B(\w1[1][29] ), .Z(
        n6388) );
  XOR \SUBBYTES[1].a/U4800  ( .A(\SUBBYTES[1].a/w2676 ), .B(
        \SUBBYTES[1].a/w2683 ), .Z(n6389) );
  XOR \SUBBYTES[1].a/U4799  ( .A(n7008), .B(n7006), .Z(\SUBBYTES[1].a/w2706 )
         );
  XOR \SUBBYTES[1].a/U4798  ( .A(\w1[1][29] ), .B(n6390), .Z(n7009) );
  XOR \SUBBYTES[1].a/U4797  ( .A(\SUBBYTES[1].a/w2668 ), .B(
        \SUBBYTES[1].a/w2678 ), .Z(n6390) );
  XOR \SUBBYTES[1].a/U4796  ( .A(n6392), .B(n6391), .Z(\SUBBYTES[1].a/w2693 )
         );
  XOR \SUBBYTES[1].a/U4795  ( .A(n7009), .B(n6393), .Z(n6391) );
  XOR \SUBBYTES[1].a/U4794  ( .A(\w1[1][28] ), .B(\SUBBYTES[1].a/w2757 ), .Z(
        n6392) );
  XOR \SUBBYTES[1].a/U4793  ( .A(\SUBBYTES[1].a/w2670 ), .B(
        \SUBBYTES[1].a/w2675 ), .Z(n6393) );
  XOR \SUBBYTES[1].a/U4792  ( .A(n6395), .B(n6394), .Z(n7007) );
  XOR \SUBBYTES[1].a/U4791  ( .A(\SUBBYTES[1].a/w2703 ), .B(\w1[1][31] ), .Z(
        n6394) );
  XOR \SUBBYTES[1].a/U4790  ( .A(\SUBBYTES[1].a/w2678 ), .B(
        \SUBBYTES[1].a/w2685 ), .Z(n6395) );
  XOR \SUBBYTES[1].a/U4789  ( .A(n7006), .B(n7007), .Z(\SUBBYTES[1].a/w2705 )
         );
  XOR \SUBBYTES[1].a/U4788  ( .A(\w1[1][27] ), .B(n6396), .Z(n7010) );
  XOR \SUBBYTES[1].a/U4787  ( .A(\SUBBYTES[1].a/w2667 ), .B(
        \SUBBYTES[1].a/w2670 ), .Z(n6396) );
  XOR \SUBBYTES[1].a/U4786  ( .A(n6398), .B(n6397), .Z(\SUBBYTES[1].a/w2694 )
         );
  XOR \SUBBYTES[1].a/U4785  ( .A(n7010), .B(n6399), .Z(n6397) );
  XOR \SUBBYTES[1].a/U4784  ( .A(\w1[1][30] ), .B(\SUBBYTES[1].a/w2736 ), .Z(
        n6398) );
  XOR \SUBBYTES[1].a/U4783  ( .A(\SUBBYTES[1].a/w2675 ), .B(
        \SUBBYTES[1].a/w2676 ), .Z(n6399) );
  XOR \SUBBYTES[1].a/U4782  ( .A(n7008), .B(n7007), .Z(\SUBBYTES[1].a/w2714 )
         );
  XOR \SUBBYTES[1].a/U4781  ( .A(n6401), .B(n6400), .Z(\SUBBYTES[1].a/w2715 )
         );
  XOR \SUBBYTES[1].a/U4780  ( .A(\w1[1][31] ), .B(n7009), .Z(n6400) );
  XOR \SUBBYTES[1].a/U4779  ( .A(\SUBBYTES[1].a/w2667 ), .B(
        \SUBBYTES[1].a/w2676 ), .Z(n6401) );
  XOR \SUBBYTES[1].a/U4778  ( .A(n6403), .B(n6402), .Z(\SUBBYTES[1].a/w2691 )
         );
  XOR \SUBBYTES[1].a/U4777  ( .A(n6405), .B(n6404), .Z(n6402) );
  XOR \SUBBYTES[1].a/U4776  ( .A(\w1[1][31] ), .B(\SUBBYTES[1].a/w2775 ), .Z(
        n6403) );
  XOR \SUBBYTES[1].a/U4775  ( .A(\SUBBYTES[1].a/w2682 ), .B(
        \SUBBYTES[1].a/w2685 ), .Z(n6404) );
  XOR \SUBBYTES[1].a/U4774  ( .A(\SUBBYTES[1].a/w2668 ), .B(
        \SUBBYTES[1].a/w2670 ), .Z(n6405) );
  XOR \SUBBYTES[1].a/U4773  ( .A(n6407), .B(n6406), .Z(\SUBBYTES[1].a/w2692 )
         );
  XOR \SUBBYTES[1].a/U4772  ( .A(n7010), .B(n6408), .Z(n6406) );
  XOR \SUBBYTES[1].a/U4771  ( .A(\w1[1][29] ), .B(n7011), .Z(n6407) );
  XOR \SUBBYTES[1].a/U4770  ( .A(\SUBBYTES[1].a/w2682 ), .B(
        \SUBBYTES[1].a/w2683 ), .Z(n6408) );
  XOR \SUBBYTES[1].a/U4769  ( .A(n6410), .B(n6409), .Z(\SUBBYTES[1].a/w2708 )
         );
  XOR \SUBBYTES[1].a/U4768  ( .A(\w1[1][25] ), .B(n6411), .Z(n6409) );
  XOR \SUBBYTES[1].a/U4767  ( .A(\SUBBYTES[1].a/w2683 ), .B(
        \SUBBYTES[1].a/w2685 ), .Z(n6410) );
  XOR \SUBBYTES[1].a/U4766  ( .A(\SUBBYTES[1].a/w2667 ), .B(
        \SUBBYTES[1].a/w2668 ), .Z(n6411) );
  XOR \SUBBYTES[1].a/U4765  ( .A(\w1[1][33] ), .B(n6412), .Z(n7012) );
  XOR \SUBBYTES[1].a/U4764  ( .A(\w1[1][35] ), .B(\w1[1][34] ), .Z(n6412) );
  XOR \SUBBYTES[1].a/U4763  ( .A(\w1[1][38] ), .B(n7012), .Z(
        \SUBBYTES[1].a/w2550 ) );
  XOR \SUBBYTES[1].a/U4762  ( .A(\w1[1][32] ), .B(\SUBBYTES[1].a/w2550 ), .Z(
        \SUBBYTES[1].a/w2437 ) );
  XOR \SUBBYTES[1].a/U4761  ( .A(\w1[1][32] ), .B(n6413), .Z(
        \SUBBYTES[1].a/w2438 ) );
  XOR \SUBBYTES[1].a/U4760  ( .A(\w1[1][38] ), .B(\w1[1][37] ), .Z(n6413) );
  XOR \SUBBYTES[1].a/U4759  ( .A(\w1[1][37] ), .B(n7012), .Z(
        \SUBBYTES[1].a/w2568 ) );
  XOR \SUBBYTES[1].a/U4758  ( .A(n6415), .B(n6414), .Z(\SUBBYTES[1].a/w2561 )
         );
  XOR \SUBBYTES[1].a/U4757  ( .A(\w1[1][35] ), .B(\w1[1][33] ), .Z(n6414) );
  XOR \SUBBYTES[1].a/U4756  ( .A(\w1[1][39] ), .B(\w1[1][36] ), .Z(n6415) );
  XOR \SUBBYTES[1].a/U4755  ( .A(\w1[1][32] ), .B(\SUBBYTES[1].a/w2561 ), .Z(
        \SUBBYTES[1].a/w2440 ) );
  XOR \SUBBYTES[1].a/U4754  ( .A(n6417), .B(n6416), .Z(\SUBBYTES[1].a/w2548 )
         );
  XOR \SUBBYTES[1].a/U4753  ( .A(\SUBBYTES[1].a/w2509 ), .B(n968), .Z(n6416)
         );
  XOR \SUBBYTES[1].a/U4752  ( .A(\SUBBYTES[1].a/w2502 ), .B(
        \SUBBYTES[1].a/w2505 ), .Z(n6417) );
  XOR \SUBBYTES[1].a/U4751  ( .A(n6419), .B(n6418), .Z(\SUBBYTES[1].a/w2549 )
         );
  XOR \SUBBYTES[1].a/U4750  ( .A(\SUBBYTES[1].a/w2509 ), .B(n5855), .Z(n6418)
         );
  XOR \SUBBYTES[1].a/U4749  ( .A(\SUBBYTES[1].a/w2502 ), .B(n5854), .Z(n6419)
         );
  XOR \SUBBYTES[1].a/U4748  ( .A(\SUBBYTES[1].a/w2561 ), .B(n6420), .Z(
        \SUBBYTES[1].a/w2551 ) );
  XOR \SUBBYTES[1].a/U4747  ( .A(\w1[1][38] ), .B(\w1[1][37] ), .Z(n6420) );
  XOR \SUBBYTES[1].a/U4746  ( .A(n6422), .B(n6421), .Z(\SUBBYTES[1].a/w2552 )
         );
  XOR \SUBBYTES[1].a/U4745  ( .A(n5855), .B(n968), .Z(n6421) );
  XOR \SUBBYTES[1].a/U4744  ( .A(n5854), .B(\SUBBYTES[1].a/w2505 ), .Z(n6422)
         );
  XOR \SUBBYTES[1].a/U4743  ( .A(\w1[1][39] ), .B(\w1[1][34] ), .Z(n7018) );
  XOR \SUBBYTES[1].a/U4742  ( .A(n7018), .B(n6423), .Z(\SUBBYTES[1].a/w2553 )
         );
  XOR \SUBBYTES[1].a/U4741  ( .A(\w1[1][37] ), .B(\w1[1][36] ), .Z(n6423) );
  XOR \SUBBYTES[1].a/U4740  ( .A(\w1[1][39] ), .B(\SUBBYTES[1].a/w2438 ), .Z(
        \SUBBYTES[1].a/w2441 ) );
  XOR \SUBBYTES[1].a/U4739  ( .A(\w1[1][33] ), .B(\SUBBYTES[1].a/w2438 ), .Z(
        \SUBBYTES[1].a/w2442 ) );
  XOR \SUBBYTES[1].a/U4738  ( .A(\w1[1][36] ), .B(\SUBBYTES[1].a/w2438 ), .Z(
        \SUBBYTES[1].a/w2443 ) );
  XOR \SUBBYTES[1].a/U4737  ( .A(\SUBBYTES[1].a/w2442 ), .B(n7018), .Z(
        \SUBBYTES[1].a/w2444 ) );
  XOR \SUBBYTES[1].a/U4736  ( .A(n7018), .B(n6424), .Z(\SUBBYTES[1].a/w2529 )
         );
  XOR \SUBBYTES[1].a/U4735  ( .A(\w1[1][36] ), .B(\w1[1][33] ), .Z(n6424) );
  XOR \SUBBYTES[1].a/U4734  ( .A(n6426), .B(n6425), .Z(n7015) );
  XOR \SUBBYTES[1].a/U4733  ( .A(\w1[1][36] ), .B(n6427), .Z(n6425) );
  XOR \SUBBYTES[1].a/U4732  ( .A(\SUBBYTES[1].a/w2494 ), .B(\w1[1][38] ), .Z(
        n6426) );
  XOR \SUBBYTES[1].a/U4731  ( .A(\SUBBYTES[1].a/w2468 ), .B(
        \SUBBYTES[1].a/w2475 ), .Z(n6427) );
  XOR \SUBBYTES[1].a/U4730  ( .A(n6429), .B(n6428), .Z(n7013) );
  XOR \SUBBYTES[1].a/U4729  ( .A(\w1[1][33] ), .B(n6430), .Z(n6428) );
  XOR \SUBBYTES[1].a/U4728  ( .A(\SUBBYTES[1].a/w2493 ), .B(\w1[1][37] ), .Z(
        n6429) );
  XOR \SUBBYTES[1].a/U4727  ( .A(\SUBBYTES[1].a/w2469 ), .B(
        \SUBBYTES[1].a/w2476 ), .Z(n6430) );
  XOR \SUBBYTES[1].a/U4726  ( .A(n7015), .B(n7013), .Z(\SUBBYTES[1].a/w2499 )
         );
  XOR \SUBBYTES[1].a/U4725  ( .A(\w1[1][37] ), .B(n6431), .Z(n7016) );
  XOR \SUBBYTES[1].a/U4724  ( .A(\SUBBYTES[1].a/w2461 ), .B(
        \SUBBYTES[1].a/w2471 ), .Z(n6431) );
  XOR \SUBBYTES[1].a/U4723  ( .A(n6433), .B(n6432), .Z(\SUBBYTES[1].a/w2486 )
         );
  XOR \SUBBYTES[1].a/U4722  ( .A(n7016), .B(n6434), .Z(n6432) );
  XOR \SUBBYTES[1].a/U4721  ( .A(\w1[1][36] ), .B(\SUBBYTES[1].a/w2550 ), .Z(
        n6433) );
  XOR \SUBBYTES[1].a/U4720  ( .A(\SUBBYTES[1].a/w2463 ), .B(
        \SUBBYTES[1].a/w2468 ), .Z(n6434) );
  XOR \SUBBYTES[1].a/U4719  ( .A(n6436), .B(n6435), .Z(n7014) );
  XOR \SUBBYTES[1].a/U4718  ( .A(\SUBBYTES[1].a/w2496 ), .B(\w1[1][39] ), .Z(
        n6435) );
  XOR \SUBBYTES[1].a/U4717  ( .A(\SUBBYTES[1].a/w2471 ), .B(
        \SUBBYTES[1].a/w2478 ), .Z(n6436) );
  XOR \SUBBYTES[1].a/U4716  ( .A(n7013), .B(n7014), .Z(\SUBBYTES[1].a/w2498 )
         );
  XOR \SUBBYTES[1].a/U4715  ( .A(\w1[1][35] ), .B(n6437), .Z(n7017) );
  XOR \SUBBYTES[1].a/U4714  ( .A(\SUBBYTES[1].a/w2460 ), .B(
        \SUBBYTES[1].a/w2463 ), .Z(n6437) );
  XOR \SUBBYTES[1].a/U4713  ( .A(n6439), .B(n6438), .Z(\SUBBYTES[1].a/w2487 )
         );
  XOR \SUBBYTES[1].a/U4712  ( .A(n7017), .B(n6440), .Z(n6438) );
  XOR \SUBBYTES[1].a/U4711  ( .A(\w1[1][38] ), .B(\SUBBYTES[1].a/w2529 ), .Z(
        n6439) );
  XOR \SUBBYTES[1].a/U4710  ( .A(\SUBBYTES[1].a/w2468 ), .B(
        \SUBBYTES[1].a/w2469 ), .Z(n6440) );
  XOR \SUBBYTES[1].a/U4709  ( .A(n7015), .B(n7014), .Z(\SUBBYTES[1].a/w2507 )
         );
  XOR \SUBBYTES[1].a/U4708  ( .A(n6442), .B(n6441), .Z(\SUBBYTES[1].a/w2508 )
         );
  XOR \SUBBYTES[1].a/U4707  ( .A(\w1[1][39] ), .B(n7016), .Z(n6441) );
  XOR \SUBBYTES[1].a/U4706  ( .A(\SUBBYTES[1].a/w2460 ), .B(
        \SUBBYTES[1].a/w2469 ), .Z(n6442) );
  XOR \SUBBYTES[1].a/U4705  ( .A(n6444), .B(n6443), .Z(\SUBBYTES[1].a/w2484 )
         );
  XOR \SUBBYTES[1].a/U4704  ( .A(n6446), .B(n6445), .Z(n6443) );
  XOR \SUBBYTES[1].a/U4703  ( .A(\w1[1][39] ), .B(\SUBBYTES[1].a/w2568 ), .Z(
        n6444) );
  XOR \SUBBYTES[1].a/U4702  ( .A(\SUBBYTES[1].a/w2475 ), .B(
        \SUBBYTES[1].a/w2478 ), .Z(n6445) );
  XOR \SUBBYTES[1].a/U4701  ( .A(\SUBBYTES[1].a/w2461 ), .B(
        \SUBBYTES[1].a/w2463 ), .Z(n6446) );
  XOR \SUBBYTES[1].a/U4700  ( .A(n6448), .B(n6447), .Z(\SUBBYTES[1].a/w2485 )
         );
  XOR \SUBBYTES[1].a/U4699  ( .A(n7017), .B(n6449), .Z(n6447) );
  XOR \SUBBYTES[1].a/U4698  ( .A(\w1[1][37] ), .B(n7018), .Z(n6448) );
  XOR \SUBBYTES[1].a/U4697  ( .A(\SUBBYTES[1].a/w2475 ), .B(
        \SUBBYTES[1].a/w2476 ), .Z(n6449) );
  XOR \SUBBYTES[1].a/U4696  ( .A(n6451), .B(n6450), .Z(\SUBBYTES[1].a/w2501 )
         );
  XOR \SUBBYTES[1].a/U4695  ( .A(\w1[1][33] ), .B(n6452), .Z(n6450) );
  XOR \SUBBYTES[1].a/U4694  ( .A(\SUBBYTES[1].a/w2476 ), .B(
        \SUBBYTES[1].a/w2478 ), .Z(n6451) );
  XOR \SUBBYTES[1].a/U4693  ( .A(\SUBBYTES[1].a/w2460 ), .B(
        \SUBBYTES[1].a/w2461 ), .Z(n6452) );
  XOR \SUBBYTES[1].a/U4692  ( .A(\w1[1][41] ), .B(n6453), .Z(n7019) );
  XOR \SUBBYTES[1].a/U4691  ( .A(\w1[1][43] ), .B(\w1[1][42] ), .Z(n6453) );
  XOR \SUBBYTES[1].a/U4690  ( .A(\w1[1][46] ), .B(n7019), .Z(
        \SUBBYTES[1].a/w2343 ) );
  XOR \SUBBYTES[1].a/U4689  ( .A(\w1[1][40] ), .B(\SUBBYTES[1].a/w2343 ), .Z(
        \SUBBYTES[1].a/w2230 ) );
  XOR \SUBBYTES[1].a/U4688  ( .A(\w1[1][40] ), .B(n6454), .Z(
        \SUBBYTES[1].a/w2231 ) );
  XOR \SUBBYTES[1].a/U4687  ( .A(\w1[1][46] ), .B(\w1[1][45] ), .Z(n6454) );
  XOR \SUBBYTES[1].a/U4686  ( .A(\w1[1][45] ), .B(n7019), .Z(
        \SUBBYTES[1].a/w2361 ) );
  XOR \SUBBYTES[1].a/U4685  ( .A(n6456), .B(n6455), .Z(\SUBBYTES[1].a/w2354 )
         );
  XOR \SUBBYTES[1].a/U4684  ( .A(\w1[1][43] ), .B(\w1[1][41] ), .Z(n6455) );
  XOR \SUBBYTES[1].a/U4683  ( .A(\w1[1][47] ), .B(\w1[1][44] ), .Z(n6456) );
  XOR \SUBBYTES[1].a/U4682  ( .A(\w1[1][40] ), .B(\SUBBYTES[1].a/w2354 ), .Z(
        \SUBBYTES[1].a/w2233 ) );
  XOR \SUBBYTES[1].a/U4681  ( .A(n6458), .B(n6457), .Z(\SUBBYTES[1].a/w2341 )
         );
  XOR \SUBBYTES[1].a/U4680  ( .A(\SUBBYTES[1].a/w2302 ), .B(n967), .Z(n6457)
         );
  XOR \SUBBYTES[1].a/U4679  ( .A(\SUBBYTES[1].a/w2295 ), .B(
        \SUBBYTES[1].a/w2298 ), .Z(n6458) );
  XOR \SUBBYTES[1].a/U4678  ( .A(n6460), .B(n6459), .Z(\SUBBYTES[1].a/w2342 )
         );
  XOR \SUBBYTES[1].a/U4677  ( .A(\SUBBYTES[1].a/w2302 ), .B(n5853), .Z(n6459)
         );
  XOR \SUBBYTES[1].a/U4676  ( .A(\SUBBYTES[1].a/w2295 ), .B(n5852), .Z(n6460)
         );
  XOR \SUBBYTES[1].a/U4675  ( .A(\SUBBYTES[1].a/w2354 ), .B(n6461), .Z(
        \SUBBYTES[1].a/w2344 ) );
  XOR \SUBBYTES[1].a/U4674  ( .A(\w1[1][46] ), .B(\w1[1][45] ), .Z(n6461) );
  XOR \SUBBYTES[1].a/U4673  ( .A(n6463), .B(n6462), .Z(\SUBBYTES[1].a/w2345 )
         );
  XOR \SUBBYTES[1].a/U4672  ( .A(n5853), .B(n967), .Z(n6462) );
  XOR \SUBBYTES[1].a/U4671  ( .A(n5852), .B(\SUBBYTES[1].a/w2298 ), .Z(n6463)
         );
  XOR \SUBBYTES[1].a/U4670  ( .A(\w1[1][47] ), .B(\w1[1][42] ), .Z(n7025) );
  XOR \SUBBYTES[1].a/U4669  ( .A(n7025), .B(n6464), .Z(\SUBBYTES[1].a/w2346 )
         );
  XOR \SUBBYTES[1].a/U4668  ( .A(\w1[1][45] ), .B(\w1[1][44] ), .Z(n6464) );
  XOR \SUBBYTES[1].a/U4667  ( .A(\w1[1][47] ), .B(\SUBBYTES[1].a/w2231 ), .Z(
        \SUBBYTES[1].a/w2234 ) );
  XOR \SUBBYTES[1].a/U4666  ( .A(\w1[1][41] ), .B(\SUBBYTES[1].a/w2231 ), .Z(
        \SUBBYTES[1].a/w2235 ) );
  XOR \SUBBYTES[1].a/U4665  ( .A(\w1[1][44] ), .B(\SUBBYTES[1].a/w2231 ), .Z(
        \SUBBYTES[1].a/w2236 ) );
  XOR \SUBBYTES[1].a/U4664  ( .A(\SUBBYTES[1].a/w2235 ), .B(n7025), .Z(
        \SUBBYTES[1].a/w2237 ) );
  XOR \SUBBYTES[1].a/U4663  ( .A(n7025), .B(n6465), .Z(\SUBBYTES[1].a/w2322 )
         );
  XOR \SUBBYTES[1].a/U4662  ( .A(\w1[1][44] ), .B(\w1[1][41] ), .Z(n6465) );
  XOR \SUBBYTES[1].a/U4661  ( .A(n6467), .B(n6466), .Z(n7022) );
  XOR \SUBBYTES[1].a/U4660  ( .A(\w1[1][44] ), .B(n6468), .Z(n6466) );
  XOR \SUBBYTES[1].a/U4659  ( .A(\SUBBYTES[1].a/w2287 ), .B(\w1[1][46] ), .Z(
        n6467) );
  XOR \SUBBYTES[1].a/U4658  ( .A(\SUBBYTES[1].a/w2261 ), .B(
        \SUBBYTES[1].a/w2268 ), .Z(n6468) );
  XOR \SUBBYTES[1].a/U4657  ( .A(n6470), .B(n6469), .Z(n7020) );
  XOR \SUBBYTES[1].a/U4656  ( .A(\w1[1][41] ), .B(n6471), .Z(n6469) );
  XOR \SUBBYTES[1].a/U4655  ( .A(\SUBBYTES[1].a/w2286 ), .B(\w1[1][45] ), .Z(
        n6470) );
  XOR \SUBBYTES[1].a/U4654  ( .A(\SUBBYTES[1].a/w2262 ), .B(
        \SUBBYTES[1].a/w2269 ), .Z(n6471) );
  XOR \SUBBYTES[1].a/U4653  ( .A(n7022), .B(n7020), .Z(\SUBBYTES[1].a/w2292 )
         );
  XOR \SUBBYTES[1].a/U4652  ( .A(\w1[1][45] ), .B(n6472), .Z(n7023) );
  XOR \SUBBYTES[1].a/U4651  ( .A(\SUBBYTES[1].a/w2254 ), .B(
        \SUBBYTES[1].a/w2264 ), .Z(n6472) );
  XOR \SUBBYTES[1].a/U4650  ( .A(n6474), .B(n6473), .Z(\SUBBYTES[1].a/w2279 )
         );
  XOR \SUBBYTES[1].a/U4649  ( .A(n7023), .B(n6475), .Z(n6473) );
  XOR \SUBBYTES[1].a/U4648  ( .A(\w1[1][44] ), .B(\SUBBYTES[1].a/w2343 ), .Z(
        n6474) );
  XOR \SUBBYTES[1].a/U4647  ( .A(\SUBBYTES[1].a/w2256 ), .B(
        \SUBBYTES[1].a/w2261 ), .Z(n6475) );
  XOR \SUBBYTES[1].a/U4646  ( .A(n6477), .B(n6476), .Z(n7021) );
  XOR \SUBBYTES[1].a/U4645  ( .A(\SUBBYTES[1].a/w2289 ), .B(\w1[1][47] ), .Z(
        n6476) );
  XOR \SUBBYTES[1].a/U4644  ( .A(\SUBBYTES[1].a/w2264 ), .B(
        \SUBBYTES[1].a/w2271 ), .Z(n6477) );
  XOR \SUBBYTES[1].a/U4643  ( .A(n7020), .B(n7021), .Z(\SUBBYTES[1].a/w2291 )
         );
  XOR \SUBBYTES[1].a/U4642  ( .A(\w1[1][43] ), .B(n6478), .Z(n7024) );
  XOR \SUBBYTES[1].a/U4641  ( .A(\SUBBYTES[1].a/w2253 ), .B(
        \SUBBYTES[1].a/w2256 ), .Z(n6478) );
  XOR \SUBBYTES[1].a/U4640  ( .A(n6480), .B(n6479), .Z(\SUBBYTES[1].a/w2280 )
         );
  XOR \SUBBYTES[1].a/U4639  ( .A(n7024), .B(n6481), .Z(n6479) );
  XOR \SUBBYTES[1].a/U4638  ( .A(\w1[1][46] ), .B(\SUBBYTES[1].a/w2322 ), .Z(
        n6480) );
  XOR \SUBBYTES[1].a/U4637  ( .A(\SUBBYTES[1].a/w2261 ), .B(
        \SUBBYTES[1].a/w2262 ), .Z(n6481) );
  XOR \SUBBYTES[1].a/U4636  ( .A(n7022), .B(n7021), .Z(\SUBBYTES[1].a/w2300 )
         );
  XOR \SUBBYTES[1].a/U4635  ( .A(n6483), .B(n6482), .Z(\SUBBYTES[1].a/w2301 )
         );
  XOR \SUBBYTES[1].a/U4634  ( .A(\w1[1][47] ), .B(n7023), .Z(n6482) );
  XOR \SUBBYTES[1].a/U4633  ( .A(\SUBBYTES[1].a/w2253 ), .B(
        \SUBBYTES[1].a/w2262 ), .Z(n6483) );
  XOR \SUBBYTES[1].a/U4632  ( .A(n6485), .B(n6484), .Z(\SUBBYTES[1].a/w2277 )
         );
  XOR \SUBBYTES[1].a/U4631  ( .A(n6487), .B(n6486), .Z(n6484) );
  XOR \SUBBYTES[1].a/U4630  ( .A(\w1[1][47] ), .B(\SUBBYTES[1].a/w2361 ), .Z(
        n6485) );
  XOR \SUBBYTES[1].a/U4629  ( .A(\SUBBYTES[1].a/w2268 ), .B(
        \SUBBYTES[1].a/w2271 ), .Z(n6486) );
  XOR \SUBBYTES[1].a/U4628  ( .A(\SUBBYTES[1].a/w2254 ), .B(
        \SUBBYTES[1].a/w2256 ), .Z(n6487) );
  XOR \SUBBYTES[1].a/U4627  ( .A(n6489), .B(n6488), .Z(\SUBBYTES[1].a/w2278 )
         );
  XOR \SUBBYTES[1].a/U4626  ( .A(n7024), .B(n6490), .Z(n6488) );
  XOR \SUBBYTES[1].a/U4625  ( .A(\w1[1][45] ), .B(n7025), .Z(n6489) );
  XOR \SUBBYTES[1].a/U4624  ( .A(\SUBBYTES[1].a/w2268 ), .B(
        \SUBBYTES[1].a/w2269 ), .Z(n6490) );
  XOR \SUBBYTES[1].a/U4623  ( .A(n6492), .B(n6491), .Z(\SUBBYTES[1].a/w2294 )
         );
  XOR \SUBBYTES[1].a/U4622  ( .A(\w1[1][41] ), .B(n6493), .Z(n6491) );
  XOR \SUBBYTES[1].a/U4621  ( .A(\SUBBYTES[1].a/w2269 ), .B(
        \SUBBYTES[1].a/w2271 ), .Z(n6492) );
  XOR \SUBBYTES[1].a/U4620  ( .A(\SUBBYTES[1].a/w2253 ), .B(
        \SUBBYTES[1].a/w2254 ), .Z(n6493) );
  XOR \SUBBYTES[1].a/U4619  ( .A(\w1[1][49] ), .B(n6494), .Z(n7026) );
  XOR \SUBBYTES[1].a/U4618  ( .A(\w1[1][51] ), .B(\w1[1][50] ), .Z(n6494) );
  XOR \SUBBYTES[1].a/U4617  ( .A(\w1[1][54] ), .B(n7026), .Z(
        \SUBBYTES[1].a/w2136 ) );
  XOR \SUBBYTES[1].a/U4616  ( .A(\w1[1][48] ), .B(\SUBBYTES[1].a/w2136 ), .Z(
        \SUBBYTES[1].a/w2023 ) );
  XOR \SUBBYTES[1].a/U4615  ( .A(\w1[1][48] ), .B(n6495), .Z(
        \SUBBYTES[1].a/w2024 ) );
  XOR \SUBBYTES[1].a/U4614  ( .A(\w1[1][54] ), .B(\w1[1][53] ), .Z(n6495) );
  XOR \SUBBYTES[1].a/U4613  ( .A(\w1[1][53] ), .B(n7026), .Z(
        \SUBBYTES[1].a/w2154 ) );
  XOR \SUBBYTES[1].a/U4612  ( .A(n6497), .B(n6496), .Z(\SUBBYTES[1].a/w2147 )
         );
  XOR \SUBBYTES[1].a/U4611  ( .A(\w1[1][51] ), .B(\w1[1][49] ), .Z(n6496) );
  XOR \SUBBYTES[1].a/U4610  ( .A(\w1[1][55] ), .B(\w1[1][52] ), .Z(n6497) );
  XOR \SUBBYTES[1].a/U4609  ( .A(\w1[1][48] ), .B(\SUBBYTES[1].a/w2147 ), .Z(
        \SUBBYTES[1].a/w2026 ) );
  XOR \SUBBYTES[1].a/U4608  ( .A(n6499), .B(n6498), .Z(\SUBBYTES[1].a/w2134 )
         );
  XOR \SUBBYTES[1].a/U4607  ( .A(\SUBBYTES[1].a/w2095 ), .B(n966), .Z(n6498)
         );
  XOR \SUBBYTES[1].a/U4606  ( .A(\SUBBYTES[1].a/w2088 ), .B(
        \SUBBYTES[1].a/w2091 ), .Z(n6499) );
  XOR \SUBBYTES[1].a/U4605  ( .A(n6501), .B(n6500), .Z(\SUBBYTES[1].a/w2135 )
         );
  XOR \SUBBYTES[1].a/U4604  ( .A(\SUBBYTES[1].a/w2095 ), .B(n5851), .Z(n6500)
         );
  XOR \SUBBYTES[1].a/U4603  ( .A(\SUBBYTES[1].a/w2088 ), .B(n5850), .Z(n6501)
         );
  XOR \SUBBYTES[1].a/U4602  ( .A(\SUBBYTES[1].a/w2147 ), .B(n6502), .Z(
        \SUBBYTES[1].a/w2137 ) );
  XOR \SUBBYTES[1].a/U4601  ( .A(\w1[1][54] ), .B(\w1[1][53] ), .Z(n6502) );
  XOR \SUBBYTES[1].a/U4600  ( .A(n6504), .B(n6503), .Z(\SUBBYTES[1].a/w2138 )
         );
  XOR \SUBBYTES[1].a/U4599  ( .A(n5851), .B(n966), .Z(n6503) );
  XOR \SUBBYTES[1].a/U4598  ( .A(n5850), .B(\SUBBYTES[1].a/w2091 ), .Z(n6504)
         );
  XOR \SUBBYTES[1].a/U4597  ( .A(\w1[1][55] ), .B(\w1[1][50] ), .Z(n7032) );
  XOR \SUBBYTES[1].a/U4596  ( .A(n7032), .B(n6505), .Z(\SUBBYTES[1].a/w2139 )
         );
  XOR \SUBBYTES[1].a/U4595  ( .A(\w1[1][53] ), .B(\w1[1][52] ), .Z(n6505) );
  XOR \SUBBYTES[1].a/U4594  ( .A(\w1[1][55] ), .B(\SUBBYTES[1].a/w2024 ), .Z(
        \SUBBYTES[1].a/w2027 ) );
  XOR \SUBBYTES[1].a/U4593  ( .A(\w1[1][49] ), .B(\SUBBYTES[1].a/w2024 ), .Z(
        \SUBBYTES[1].a/w2028 ) );
  XOR \SUBBYTES[1].a/U4592  ( .A(\w1[1][52] ), .B(\SUBBYTES[1].a/w2024 ), .Z(
        \SUBBYTES[1].a/w2029 ) );
  XOR \SUBBYTES[1].a/U4591  ( .A(\SUBBYTES[1].a/w2028 ), .B(n7032), .Z(
        \SUBBYTES[1].a/w2030 ) );
  XOR \SUBBYTES[1].a/U4590  ( .A(n7032), .B(n6506), .Z(\SUBBYTES[1].a/w2115 )
         );
  XOR \SUBBYTES[1].a/U4589  ( .A(\w1[1][52] ), .B(\w1[1][49] ), .Z(n6506) );
  XOR \SUBBYTES[1].a/U4588  ( .A(n6508), .B(n6507), .Z(n7029) );
  XOR \SUBBYTES[1].a/U4587  ( .A(\w1[1][52] ), .B(n6509), .Z(n6507) );
  XOR \SUBBYTES[1].a/U4586  ( .A(\SUBBYTES[1].a/w2080 ), .B(\w1[1][54] ), .Z(
        n6508) );
  XOR \SUBBYTES[1].a/U4585  ( .A(\SUBBYTES[1].a/w2054 ), .B(
        \SUBBYTES[1].a/w2061 ), .Z(n6509) );
  XOR \SUBBYTES[1].a/U4584  ( .A(n6511), .B(n6510), .Z(n7027) );
  XOR \SUBBYTES[1].a/U4583  ( .A(\w1[1][49] ), .B(n6512), .Z(n6510) );
  XOR \SUBBYTES[1].a/U4582  ( .A(\SUBBYTES[1].a/w2079 ), .B(\w1[1][53] ), .Z(
        n6511) );
  XOR \SUBBYTES[1].a/U4581  ( .A(\SUBBYTES[1].a/w2055 ), .B(
        \SUBBYTES[1].a/w2062 ), .Z(n6512) );
  XOR \SUBBYTES[1].a/U4580  ( .A(n7029), .B(n7027), .Z(\SUBBYTES[1].a/w2085 )
         );
  XOR \SUBBYTES[1].a/U4579  ( .A(\w1[1][53] ), .B(n6513), .Z(n7030) );
  XOR \SUBBYTES[1].a/U4578  ( .A(\SUBBYTES[1].a/w2047 ), .B(
        \SUBBYTES[1].a/w2057 ), .Z(n6513) );
  XOR \SUBBYTES[1].a/U4577  ( .A(n6515), .B(n6514), .Z(\SUBBYTES[1].a/w2072 )
         );
  XOR \SUBBYTES[1].a/U4576  ( .A(n7030), .B(n6516), .Z(n6514) );
  XOR \SUBBYTES[1].a/U4575  ( .A(\w1[1][52] ), .B(\SUBBYTES[1].a/w2136 ), .Z(
        n6515) );
  XOR \SUBBYTES[1].a/U4574  ( .A(\SUBBYTES[1].a/w2049 ), .B(
        \SUBBYTES[1].a/w2054 ), .Z(n6516) );
  XOR \SUBBYTES[1].a/U4573  ( .A(n6518), .B(n6517), .Z(n7028) );
  XOR \SUBBYTES[1].a/U4572  ( .A(\SUBBYTES[1].a/w2082 ), .B(\w1[1][55] ), .Z(
        n6517) );
  XOR \SUBBYTES[1].a/U4571  ( .A(\SUBBYTES[1].a/w2057 ), .B(
        \SUBBYTES[1].a/w2064 ), .Z(n6518) );
  XOR \SUBBYTES[1].a/U4570  ( .A(n7027), .B(n7028), .Z(\SUBBYTES[1].a/w2084 )
         );
  XOR \SUBBYTES[1].a/U4569  ( .A(\w1[1][51] ), .B(n6519), .Z(n7031) );
  XOR \SUBBYTES[1].a/U4568  ( .A(\SUBBYTES[1].a/w2046 ), .B(
        \SUBBYTES[1].a/w2049 ), .Z(n6519) );
  XOR \SUBBYTES[1].a/U4567  ( .A(n6521), .B(n6520), .Z(\SUBBYTES[1].a/w2073 )
         );
  XOR \SUBBYTES[1].a/U4566  ( .A(n7031), .B(n6522), .Z(n6520) );
  XOR \SUBBYTES[1].a/U4565  ( .A(\w1[1][54] ), .B(\SUBBYTES[1].a/w2115 ), .Z(
        n6521) );
  XOR \SUBBYTES[1].a/U4564  ( .A(\SUBBYTES[1].a/w2054 ), .B(
        \SUBBYTES[1].a/w2055 ), .Z(n6522) );
  XOR \SUBBYTES[1].a/U4563  ( .A(n7029), .B(n7028), .Z(\SUBBYTES[1].a/w2093 )
         );
  XOR \SUBBYTES[1].a/U4562  ( .A(n6524), .B(n6523), .Z(\SUBBYTES[1].a/w2094 )
         );
  XOR \SUBBYTES[1].a/U4561  ( .A(\w1[1][55] ), .B(n7030), .Z(n6523) );
  XOR \SUBBYTES[1].a/U4560  ( .A(\SUBBYTES[1].a/w2046 ), .B(
        \SUBBYTES[1].a/w2055 ), .Z(n6524) );
  XOR \SUBBYTES[1].a/U4559  ( .A(n6526), .B(n6525), .Z(\SUBBYTES[1].a/w2070 )
         );
  XOR \SUBBYTES[1].a/U4558  ( .A(n6528), .B(n6527), .Z(n6525) );
  XOR \SUBBYTES[1].a/U4557  ( .A(\w1[1][55] ), .B(\SUBBYTES[1].a/w2154 ), .Z(
        n6526) );
  XOR \SUBBYTES[1].a/U4556  ( .A(\SUBBYTES[1].a/w2061 ), .B(
        \SUBBYTES[1].a/w2064 ), .Z(n6527) );
  XOR \SUBBYTES[1].a/U4555  ( .A(\SUBBYTES[1].a/w2047 ), .B(
        \SUBBYTES[1].a/w2049 ), .Z(n6528) );
  XOR \SUBBYTES[1].a/U4554  ( .A(n6530), .B(n6529), .Z(\SUBBYTES[1].a/w2071 )
         );
  XOR \SUBBYTES[1].a/U4553  ( .A(n7031), .B(n6531), .Z(n6529) );
  XOR \SUBBYTES[1].a/U4552  ( .A(\w1[1][53] ), .B(n7032), .Z(n6530) );
  XOR \SUBBYTES[1].a/U4551  ( .A(\SUBBYTES[1].a/w2061 ), .B(
        \SUBBYTES[1].a/w2062 ), .Z(n6531) );
  XOR \SUBBYTES[1].a/U4550  ( .A(n6533), .B(n6532), .Z(\SUBBYTES[1].a/w2087 )
         );
  XOR \SUBBYTES[1].a/U4549  ( .A(\w1[1][49] ), .B(n6534), .Z(n6532) );
  XOR \SUBBYTES[1].a/U4548  ( .A(\SUBBYTES[1].a/w2062 ), .B(
        \SUBBYTES[1].a/w2064 ), .Z(n6533) );
  XOR \SUBBYTES[1].a/U4547  ( .A(\SUBBYTES[1].a/w2046 ), .B(
        \SUBBYTES[1].a/w2047 ), .Z(n6534) );
  XOR \SUBBYTES[1].a/U4546  ( .A(\w1[1][57] ), .B(n6535), .Z(n7033) );
  XOR \SUBBYTES[1].a/U4545  ( .A(\w1[1][59] ), .B(\w1[1][58] ), .Z(n6535) );
  XOR \SUBBYTES[1].a/U4544  ( .A(\w1[1][62] ), .B(n7033), .Z(
        \SUBBYTES[1].a/w1929 ) );
  XOR \SUBBYTES[1].a/U4543  ( .A(\w1[1][56] ), .B(\SUBBYTES[1].a/w1929 ), .Z(
        \SUBBYTES[1].a/w1816 ) );
  XOR \SUBBYTES[1].a/U4542  ( .A(\w1[1][56] ), .B(n6536), .Z(
        \SUBBYTES[1].a/w1817 ) );
  XOR \SUBBYTES[1].a/U4541  ( .A(\w1[1][62] ), .B(\w1[1][61] ), .Z(n6536) );
  XOR \SUBBYTES[1].a/U4540  ( .A(\w1[1][61] ), .B(n7033), .Z(
        \SUBBYTES[1].a/w1947 ) );
  XOR \SUBBYTES[1].a/U4539  ( .A(n6538), .B(n6537), .Z(\SUBBYTES[1].a/w1940 )
         );
  XOR \SUBBYTES[1].a/U4538  ( .A(\w1[1][59] ), .B(\w1[1][57] ), .Z(n6537) );
  XOR \SUBBYTES[1].a/U4537  ( .A(\w1[1][63] ), .B(\w1[1][60] ), .Z(n6538) );
  XOR \SUBBYTES[1].a/U4536  ( .A(\w1[1][56] ), .B(\SUBBYTES[1].a/w1940 ), .Z(
        \SUBBYTES[1].a/w1819 ) );
  XOR \SUBBYTES[1].a/U4535  ( .A(n6540), .B(n6539), .Z(\SUBBYTES[1].a/w1927 )
         );
  XOR \SUBBYTES[1].a/U4534  ( .A(\SUBBYTES[1].a/w1888 ), .B(n965), .Z(n6539)
         );
  XOR \SUBBYTES[1].a/U4533  ( .A(\SUBBYTES[1].a/w1881 ), .B(
        \SUBBYTES[1].a/w1884 ), .Z(n6540) );
  XOR \SUBBYTES[1].a/U4532  ( .A(n6542), .B(n6541), .Z(\SUBBYTES[1].a/w1928 )
         );
  XOR \SUBBYTES[1].a/U4531  ( .A(\SUBBYTES[1].a/w1888 ), .B(n5849), .Z(n6541)
         );
  XOR \SUBBYTES[1].a/U4530  ( .A(\SUBBYTES[1].a/w1881 ), .B(n5848), .Z(n6542)
         );
  XOR \SUBBYTES[1].a/U4529  ( .A(\SUBBYTES[1].a/w1940 ), .B(n6543), .Z(
        \SUBBYTES[1].a/w1930 ) );
  XOR \SUBBYTES[1].a/U4528  ( .A(\w1[1][62] ), .B(\w1[1][61] ), .Z(n6543) );
  XOR \SUBBYTES[1].a/U4527  ( .A(n6545), .B(n6544), .Z(\SUBBYTES[1].a/w1931 )
         );
  XOR \SUBBYTES[1].a/U4526  ( .A(n5849), .B(n965), .Z(n6544) );
  XOR \SUBBYTES[1].a/U4525  ( .A(n5848), .B(\SUBBYTES[1].a/w1884 ), .Z(n6545)
         );
  XOR \SUBBYTES[1].a/U4524  ( .A(\w1[1][63] ), .B(\w1[1][58] ), .Z(n7039) );
  XOR \SUBBYTES[1].a/U4523  ( .A(n7039), .B(n6546), .Z(\SUBBYTES[1].a/w1932 )
         );
  XOR \SUBBYTES[1].a/U4522  ( .A(\w1[1][61] ), .B(\w1[1][60] ), .Z(n6546) );
  XOR \SUBBYTES[1].a/U4521  ( .A(\w1[1][63] ), .B(\SUBBYTES[1].a/w1817 ), .Z(
        \SUBBYTES[1].a/w1820 ) );
  XOR \SUBBYTES[1].a/U4520  ( .A(\w1[1][57] ), .B(\SUBBYTES[1].a/w1817 ), .Z(
        \SUBBYTES[1].a/w1821 ) );
  XOR \SUBBYTES[1].a/U4519  ( .A(\w1[1][60] ), .B(\SUBBYTES[1].a/w1817 ), .Z(
        \SUBBYTES[1].a/w1822 ) );
  XOR \SUBBYTES[1].a/U4518  ( .A(\SUBBYTES[1].a/w1821 ), .B(n7039), .Z(
        \SUBBYTES[1].a/w1823 ) );
  XOR \SUBBYTES[1].a/U4517  ( .A(n7039), .B(n6547), .Z(\SUBBYTES[1].a/w1908 )
         );
  XOR \SUBBYTES[1].a/U4516  ( .A(\w1[1][60] ), .B(\w1[1][57] ), .Z(n6547) );
  XOR \SUBBYTES[1].a/U4515  ( .A(n6549), .B(n6548), .Z(n7036) );
  XOR \SUBBYTES[1].a/U4514  ( .A(\w1[1][60] ), .B(n6550), .Z(n6548) );
  XOR \SUBBYTES[1].a/U4513  ( .A(\SUBBYTES[1].a/w1873 ), .B(\w1[1][62] ), .Z(
        n6549) );
  XOR \SUBBYTES[1].a/U4512  ( .A(\SUBBYTES[1].a/w1847 ), .B(
        \SUBBYTES[1].a/w1854 ), .Z(n6550) );
  XOR \SUBBYTES[1].a/U4511  ( .A(n6552), .B(n6551), .Z(n7034) );
  XOR \SUBBYTES[1].a/U4510  ( .A(\w1[1][57] ), .B(n6553), .Z(n6551) );
  XOR \SUBBYTES[1].a/U4509  ( .A(\SUBBYTES[1].a/w1872 ), .B(\w1[1][61] ), .Z(
        n6552) );
  XOR \SUBBYTES[1].a/U4508  ( .A(\SUBBYTES[1].a/w1848 ), .B(
        \SUBBYTES[1].a/w1855 ), .Z(n6553) );
  XOR \SUBBYTES[1].a/U4507  ( .A(n7036), .B(n7034), .Z(\SUBBYTES[1].a/w1878 )
         );
  XOR \SUBBYTES[1].a/U4506  ( .A(\w1[1][61] ), .B(n6554), .Z(n7037) );
  XOR \SUBBYTES[1].a/U4505  ( .A(\SUBBYTES[1].a/w1840 ), .B(
        \SUBBYTES[1].a/w1850 ), .Z(n6554) );
  XOR \SUBBYTES[1].a/U4504  ( .A(n6556), .B(n6555), .Z(\SUBBYTES[1].a/w1865 )
         );
  XOR \SUBBYTES[1].a/U4503  ( .A(n7037), .B(n6557), .Z(n6555) );
  XOR \SUBBYTES[1].a/U4502  ( .A(\w1[1][60] ), .B(\SUBBYTES[1].a/w1929 ), .Z(
        n6556) );
  XOR \SUBBYTES[1].a/U4501  ( .A(\SUBBYTES[1].a/w1842 ), .B(
        \SUBBYTES[1].a/w1847 ), .Z(n6557) );
  XOR \SUBBYTES[1].a/U4500  ( .A(n6559), .B(n6558), .Z(n7035) );
  XOR \SUBBYTES[1].a/U4499  ( .A(\SUBBYTES[1].a/w1875 ), .B(\w1[1][63] ), .Z(
        n6558) );
  XOR \SUBBYTES[1].a/U4498  ( .A(\SUBBYTES[1].a/w1850 ), .B(
        \SUBBYTES[1].a/w1857 ), .Z(n6559) );
  XOR \SUBBYTES[1].a/U4497  ( .A(n7034), .B(n7035), .Z(\SUBBYTES[1].a/w1877 )
         );
  XOR \SUBBYTES[1].a/U4496  ( .A(\w1[1][59] ), .B(n6560), .Z(n7038) );
  XOR \SUBBYTES[1].a/U4495  ( .A(\SUBBYTES[1].a/w1839 ), .B(
        \SUBBYTES[1].a/w1842 ), .Z(n6560) );
  XOR \SUBBYTES[1].a/U4494  ( .A(n6562), .B(n6561), .Z(\SUBBYTES[1].a/w1866 )
         );
  XOR \SUBBYTES[1].a/U4493  ( .A(n7038), .B(n6563), .Z(n6561) );
  XOR \SUBBYTES[1].a/U4492  ( .A(\w1[1][62] ), .B(\SUBBYTES[1].a/w1908 ), .Z(
        n6562) );
  XOR \SUBBYTES[1].a/U4491  ( .A(\SUBBYTES[1].a/w1847 ), .B(
        \SUBBYTES[1].a/w1848 ), .Z(n6563) );
  XOR \SUBBYTES[1].a/U4490  ( .A(n7036), .B(n7035), .Z(\SUBBYTES[1].a/w1886 )
         );
  XOR \SUBBYTES[1].a/U4489  ( .A(n6565), .B(n6564), .Z(\SUBBYTES[1].a/w1887 )
         );
  XOR \SUBBYTES[1].a/U4488  ( .A(\w1[1][63] ), .B(n7037), .Z(n6564) );
  XOR \SUBBYTES[1].a/U4487  ( .A(\SUBBYTES[1].a/w1839 ), .B(
        \SUBBYTES[1].a/w1848 ), .Z(n6565) );
  XOR \SUBBYTES[1].a/U4486  ( .A(n6567), .B(n6566), .Z(\SUBBYTES[1].a/w1863 )
         );
  XOR \SUBBYTES[1].a/U4485  ( .A(n6569), .B(n6568), .Z(n6566) );
  XOR \SUBBYTES[1].a/U4484  ( .A(\w1[1][63] ), .B(\SUBBYTES[1].a/w1947 ), .Z(
        n6567) );
  XOR \SUBBYTES[1].a/U4483  ( .A(\SUBBYTES[1].a/w1854 ), .B(
        \SUBBYTES[1].a/w1857 ), .Z(n6568) );
  XOR \SUBBYTES[1].a/U4482  ( .A(\SUBBYTES[1].a/w1840 ), .B(
        \SUBBYTES[1].a/w1842 ), .Z(n6569) );
  XOR \SUBBYTES[1].a/U4481  ( .A(n6571), .B(n6570), .Z(\SUBBYTES[1].a/w1864 )
         );
  XOR \SUBBYTES[1].a/U4480  ( .A(n7038), .B(n6572), .Z(n6570) );
  XOR \SUBBYTES[1].a/U4479  ( .A(\w1[1][61] ), .B(n7039), .Z(n6571) );
  XOR \SUBBYTES[1].a/U4478  ( .A(\SUBBYTES[1].a/w1854 ), .B(
        \SUBBYTES[1].a/w1855 ), .Z(n6572) );
  XOR \SUBBYTES[1].a/U4477  ( .A(n6574), .B(n6573), .Z(\SUBBYTES[1].a/w1880 )
         );
  XOR \SUBBYTES[1].a/U4476  ( .A(\w1[1][57] ), .B(n6575), .Z(n6573) );
  XOR \SUBBYTES[1].a/U4475  ( .A(\SUBBYTES[1].a/w1855 ), .B(
        \SUBBYTES[1].a/w1857 ), .Z(n6574) );
  XOR \SUBBYTES[1].a/U4474  ( .A(\SUBBYTES[1].a/w1839 ), .B(
        \SUBBYTES[1].a/w1840 ), .Z(n6575) );
  XOR \SUBBYTES[1].a/U4473  ( .A(\w1[1][65] ), .B(n6576), .Z(n7040) );
  XOR \SUBBYTES[1].a/U4472  ( .A(\w1[1][67] ), .B(\w1[1][66] ), .Z(n6576) );
  XOR \SUBBYTES[1].a/U4471  ( .A(\w1[1][70] ), .B(n7040), .Z(
        \SUBBYTES[1].a/w1722 ) );
  XOR \SUBBYTES[1].a/U4470  ( .A(\w1[1][64] ), .B(\SUBBYTES[1].a/w1722 ), .Z(
        \SUBBYTES[1].a/w1609 ) );
  XOR \SUBBYTES[1].a/U4469  ( .A(\w1[1][64] ), .B(n6577), .Z(
        \SUBBYTES[1].a/w1610 ) );
  XOR \SUBBYTES[1].a/U4468  ( .A(\w1[1][70] ), .B(\w1[1][69] ), .Z(n6577) );
  XOR \SUBBYTES[1].a/U4467  ( .A(\w1[1][69] ), .B(n7040), .Z(
        \SUBBYTES[1].a/w1740 ) );
  XOR \SUBBYTES[1].a/U4466  ( .A(n6579), .B(n6578), .Z(\SUBBYTES[1].a/w1733 )
         );
  XOR \SUBBYTES[1].a/U4465  ( .A(\w1[1][67] ), .B(\w1[1][65] ), .Z(n6578) );
  XOR \SUBBYTES[1].a/U4464  ( .A(\w1[1][71] ), .B(\w1[1][68] ), .Z(n6579) );
  XOR \SUBBYTES[1].a/U4463  ( .A(\w1[1][64] ), .B(\SUBBYTES[1].a/w1733 ), .Z(
        \SUBBYTES[1].a/w1612 ) );
  XOR \SUBBYTES[1].a/U4462  ( .A(n6581), .B(n6580), .Z(\SUBBYTES[1].a/w1720 )
         );
  XOR \SUBBYTES[1].a/U4461  ( .A(\SUBBYTES[1].a/w1681 ), .B(n964), .Z(n6580)
         );
  XOR \SUBBYTES[1].a/U4460  ( .A(\SUBBYTES[1].a/w1674 ), .B(
        \SUBBYTES[1].a/w1677 ), .Z(n6581) );
  XOR \SUBBYTES[1].a/U4459  ( .A(n6583), .B(n6582), .Z(\SUBBYTES[1].a/w1721 )
         );
  XOR \SUBBYTES[1].a/U4458  ( .A(\SUBBYTES[1].a/w1681 ), .B(n5847), .Z(n6582)
         );
  XOR \SUBBYTES[1].a/U4457  ( .A(\SUBBYTES[1].a/w1674 ), .B(n5846), .Z(n6583)
         );
  XOR \SUBBYTES[1].a/U4456  ( .A(\SUBBYTES[1].a/w1733 ), .B(n6584), .Z(
        \SUBBYTES[1].a/w1723 ) );
  XOR \SUBBYTES[1].a/U4455  ( .A(\w1[1][70] ), .B(\w1[1][69] ), .Z(n6584) );
  XOR \SUBBYTES[1].a/U4454  ( .A(n6586), .B(n6585), .Z(\SUBBYTES[1].a/w1724 )
         );
  XOR \SUBBYTES[1].a/U4453  ( .A(n5847), .B(n964), .Z(n6585) );
  XOR \SUBBYTES[1].a/U4452  ( .A(n5846), .B(\SUBBYTES[1].a/w1677 ), .Z(n6586)
         );
  XOR \SUBBYTES[1].a/U4451  ( .A(\w1[1][71] ), .B(\w1[1][66] ), .Z(n7046) );
  XOR \SUBBYTES[1].a/U4450  ( .A(n7046), .B(n6587), .Z(\SUBBYTES[1].a/w1725 )
         );
  XOR \SUBBYTES[1].a/U4449  ( .A(\w1[1][69] ), .B(\w1[1][68] ), .Z(n6587) );
  XOR \SUBBYTES[1].a/U4448  ( .A(\w1[1][71] ), .B(\SUBBYTES[1].a/w1610 ), .Z(
        \SUBBYTES[1].a/w1613 ) );
  XOR \SUBBYTES[1].a/U4447  ( .A(\w1[1][65] ), .B(\SUBBYTES[1].a/w1610 ), .Z(
        \SUBBYTES[1].a/w1614 ) );
  XOR \SUBBYTES[1].a/U4446  ( .A(\w1[1][68] ), .B(\SUBBYTES[1].a/w1610 ), .Z(
        \SUBBYTES[1].a/w1615 ) );
  XOR \SUBBYTES[1].a/U4445  ( .A(\SUBBYTES[1].a/w1614 ), .B(n7046), .Z(
        \SUBBYTES[1].a/w1616 ) );
  XOR \SUBBYTES[1].a/U4444  ( .A(n7046), .B(n6588), .Z(\SUBBYTES[1].a/w1701 )
         );
  XOR \SUBBYTES[1].a/U4443  ( .A(\w1[1][68] ), .B(\w1[1][65] ), .Z(n6588) );
  XOR \SUBBYTES[1].a/U4442  ( .A(n6590), .B(n6589), .Z(n7043) );
  XOR \SUBBYTES[1].a/U4441  ( .A(\w1[1][68] ), .B(n6591), .Z(n6589) );
  XOR \SUBBYTES[1].a/U4440  ( .A(\SUBBYTES[1].a/w1666 ), .B(\w1[1][70] ), .Z(
        n6590) );
  XOR \SUBBYTES[1].a/U4439  ( .A(\SUBBYTES[1].a/w1640 ), .B(
        \SUBBYTES[1].a/w1647 ), .Z(n6591) );
  XOR \SUBBYTES[1].a/U4438  ( .A(n6593), .B(n6592), .Z(n7041) );
  XOR \SUBBYTES[1].a/U4437  ( .A(\w1[1][65] ), .B(n6594), .Z(n6592) );
  XOR \SUBBYTES[1].a/U4436  ( .A(\SUBBYTES[1].a/w1665 ), .B(\w1[1][69] ), .Z(
        n6593) );
  XOR \SUBBYTES[1].a/U4435  ( .A(\SUBBYTES[1].a/w1641 ), .B(
        \SUBBYTES[1].a/w1648 ), .Z(n6594) );
  XOR \SUBBYTES[1].a/U4434  ( .A(n7043), .B(n7041), .Z(\SUBBYTES[1].a/w1671 )
         );
  XOR \SUBBYTES[1].a/U4433  ( .A(\w1[1][69] ), .B(n6595), .Z(n7044) );
  XOR \SUBBYTES[1].a/U4432  ( .A(\SUBBYTES[1].a/w1633 ), .B(
        \SUBBYTES[1].a/w1643 ), .Z(n6595) );
  XOR \SUBBYTES[1].a/U4431  ( .A(n6597), .B(n6596), .Z(\SUBBYTES[1].a/w1658 )
         );
  XOR \SUBBYTES[1].a/U4430  ( .A(n7044), .B(n6598), .Z(n6596) );
  XOR \SUBBYTES[1].a/U4429  ( .A(\w1[1][68] ), .B(\SUBBYTES[1].a/w1722 ), .Z(
        n6597) );
  XOR \SUBBYTES[1].a/U4428  ( .A(\SUBBYTES[1].a/w1635 ), .B(
        \SUBBYTES[1].a/w1640 ), .Z(n6598) );
  XOR \SUBBYTES[1].a/U4427  ( .A(n6600), .B(n6599), .Z(n7042) );
  XOR \SUBBYTES[1].a/U4426  ( .A(\SUBBYTES[1].a/w1668 ), .B(\w1[1][71] ), .Z(
        n6599) );
  XOR \SUBBYTES[1].a/U4425  ( .A(\SUBBYTES[1].a/w1643 ), .B(
        \SUBBYTES[1].a/w1650 ), .Z(n6600) );
  XOR \SUBBYTES[1].a/U4424  ( .A(n7041), .B(n7042), .Z(\SUBBYTES[1].a/w1670 )
         );
  XOR \SUBBYTES[1].a/U4423  ( .A(\w1[1][67] ), .B(n6601), .Z(n7045) );
  XOR \SUBBYTES[1].a/U4422  ( .A(\SUBBYTES[1].a/w1632 ), .B(
        \SUBBYTES[1].a/w1635 ), .Z(n6601) );
  XOR \SUBBYTES[1].a/U4421  ( .A(n6603), .B(n6602), .Z(\SUBBYTES[1].a/w1659 )
         );
  XOR \SUBBYTES[1].a/U4420  ( .A(n7045), .B(n6604), .Z(n6602) );
  XOR \SUBBYTES[1].a/U4419  ( .A(\w1[1][70] ), .B(\SUBBYTES[1].a/w1701 ), .Z(
        n6603) );
  XOR \SUBBYTES[1].a/U4418  ( .A(\SUBBYTES[1].a/w1640 ), .B(
        \SUBBYTES[1].a/w1641 ), .Z(n6604) );
  XOR \SUBBYTES[1].a/U4417  ( .A(n7043), .B(n7042), .Z(\SUBBYTES[1].a/w1679 )
         );
  XOR \SUBBYTES[1].a/U4416  ( .A(n6606), .B(n6605), .Z(\SUBBYTES[1].a/w1680 )
         );
  XOR \SUBBYTES[1].a/U4415  ( .A(\w1[1][71] ), .B(n7044), .Z(n6605) );
  XOR \SUBBYTES[1].a/U4414  ( .A(\SUBBYTES[1].a/w1632 ), .B(
        \SUBBYTES[1].a/w1641 ), .Z(n6606) );
  XOR \SUBBYTES[1].a/U4413  ( .A(n6608), .B(n6607), .Z(\SUBBYTES[1].a/w1656 )
         );
  XOR \SUBBYTES[1].a/U4412  ( .A(n6610), .B(n6609), .Z(n6607) );
  XOR \SUBBYTES[1].a/U4411  ( .A(\w1[1][71] ), .B(\SUBBYTES[1].a/w1740 ), .Z(
        n6608) );
  XOR \SUBBYTES[1].a/U4410  ( .A(\SUBBYTES[1].a/w1647 ), .B(
        \SUBBYTES[1].a/w1650 ), .Z(n6609) );
  XOR \SUBBYTES[1].a/U4409  ( .A(\SUBBYTES[1].a/w1633 ), .B(
        \SUBBYTES[1].a/w1635 ), .Z(n6610) );
  XOR \SUBBYTES[1].a/U4408  ( .A(n6612), .B(n6611), .Z(\SUBBYTES[1].a/w1657 )
         );
  XOR \SUBBYTES[1].a/U4407  ( .A(n7045), .B(n6613), .Z(n6611) );
  XOR \SUBBYTES[1].a/U4406  ( .A(\w1[1][69] ), .B(n7046), .Z(n6612) );
  XOR \SUBBYTES[1].a/U4405  ( .A(\SUBBYTES[1].a/w1647 ), .B(
        \SUBBYTES[1].a/w1648 ), .Z(n6613) );
  XOR \SUBBYTES[1].a/U4404  ( .A(n6615), .B(n6614), .Z(\SUBBYTES[1].a/w1673 )
         );
  XOR \SUBBYTES[1].a/U4403  ( .A(\w1[1][65] ), .B(n6616), .Z(n6614) );
  XOR \SUBBYTES[1].a/U4402  ( .A(\SUBBYTES[1].a/w1648 ), .B(
        \SUBBYTES[1].a/w1650 ), .Z(n6615) );
  XOR \SUBBYTES[1].a/U4401  ( .A(\SUBBYTES[1].a/w1632 ), .B(
        \SUBBYTES[1].a/w1633 ), .Z(n6616) );
  XOR \SUBBYTES[1].a/U4400  ( .A(\w1[1][73] ), .B(n6617), .Z(n7047) );
  XOR \SUBBYTES[1].a/U4399  ( .A(\w1[1][75] ), .B(\w1[1][74] ), .Z(n6617) );
  XOR \SUBBYTES[1].a/U4398  ( .A(\w1[1][78] ), .B(n7047), .Z(
        \SUBBYTES[1].a/w1515 ) );
  XOR \SUBBYTES[1].a/U4397  ( .A(\w1[1][72] ), .B(\SUBBYTES[1].a/w1515 ), .Z(
        \SUBBYTES[1].a/w1402 ) );
  XOR \SUBBYTES[1].a/U4396  ( .A(\w1[1][72] ), .B(n6618), .Z(
        \SUBBYTES[1].a/w1403 ) );
  XOR \SUBBYTES[1].a/U4395  ( .A(\w1[1][78] ), .B(\w1[1][77] ), .Z(n6618) );
  XOR \SUBBYTES[1].a/U4394  ( .A(\w1[1][77] ), .B(n7047), .Z(
        \SUBBYTES[1].a/w1533 ) );
  XOR \SUBBYTES[1].a/U4393  ( .A(n6620), .B(n6619), .Z(\SUBBYTES[1].a/w1526 )
         );
  XOR \SUBBYTES[1].a/U4392  ( .A(\w1[1][75] ), .B(\w1[1][73] ), .Z(n6619) );
  XOR \SUBBYTES[1].a/U4391  ( .A(\w1[1][79] ), .B(\w1[1][76] ), .Z(n6620) );
  XOR \SUBBYTES[1].a/U4390  ( .A(\w1[1][72] ), .B(\SUBBYTES[1].a/w1526 ), .Z(
        \SUBBYTES[1].a/w1405 ) );
  XOR \SUBBYTES[1].a/U4389  ( .A(n6622), .B(n6621), .Z(\SUBBYTES[1].a/w1513 )
         );
  XOR \SUBBYTES[1].a/U4388  ( .A(\SUBBYTES[1].a/w1474 ), .B(n963), .Z(n6621)
         );
  XOR \SUBBYTES[1].a/U4387  ( .A(\SUBBYTES[1].a/w1467 ), .B(
        \SUBBYTES[1].a/w1470 ), .Z(n6622) );
  XOR \SUBBYTES[1].a/U4386  ( .A(n6624), .B(n6623), .Z(\SUBBYTES[1].a/w1514 )
         );
  XOR \SUBBYTES[1].a/U4385  ( .A(\SUBBYTES[1].a/w1474 ), .B(n5845), .Z(n6623)
         );
  XOR \SUBBYTES[1].a/U4384  ( .A(\SUBBYTES[1].a/w1467 ), .B(n5844), .Z(n6624)
         );
  XOR \SUBBYTES[1].a/U4383  ( .A(\SUBBYTES[1].a/w1526 ), .B(n6625), .Z(
        \SUBBYTES[1].a/w1516 ) );
  XOR \SUBBYTES[1].a/U4382  ( .A(\w1[1][78] ), .B(\w1[1][77] ), .Z(n6625) );
  XOR \SUBBYTES[1].a/U4381  ( .A(n6627), .B(n6626), .Z(\SUBBYTES[1].a/w1517 )
         );
  XOR \SUBBYTES[1].a/U4380  ( .A(n5845), .B(n963), .Z(n6626) );
  XOR \SUBBYTES[1].a/U4379  ( .A(n5844), .B(\SUBBYTES[1].a/w1470 ), .Z(n6627)
         );
  XOR \SUBBYTES[1].a/U4378  ( .A(\w1[1][79] ), .B(\w1[1][74] ), .Z(n7053) );
  XOR \SUBBYTES[1].a/U4377  ( .A(n7053), .B(n6628), .Z(\SUBBYTES[1].a/w1518 )
         );
  XOR \SUBBYTES[1].a/U4376  ( .A(\w1[1][77] ), .B(\w1[1][76] ), .Z(n6628) );
  XOR \SUBBYTES[1].a/U4375  ( .A(\w1[1][79] ), .B(\SUBBYTES[1].a/w1403 ), .Z(
        \SUBBYTES[1].a/w1406 ) );
  XOR \SUBBYTES[1].a/U4374  ( .A(\w1[1][73] ), .B(\SUBBYTES[1].a/w1403 ), .Z(
        \SUBBYTES[1].a/w1407 ) );
  XOR \SUBBYTES[1].a/U4373  ( .A(\w1[1][76] ), .B(\SUBBYTES[1].a/w1403 ), .Z(
        \SUBBYTES[1].a/w1408 ) );
  XOR \SUBBYTES[1].a/U4372  ( .A(\SUBBYTES[1].a/w1407 ), .B(n7053), .Z(
        \SUBBYTES[1].a/w1409 ) );
  XOR \SUBBYTES[1].a/U4371  ( .A(n7053), .B(n6629), .Z(\SUBBYTES[1].a/w1494 )
         );
  XOR \SUBBYTES[1].a/U4370  ( .A(\w1[1][76] ), .B(\w1[1][73] ), .Z(n6629) );
  XOR \SUBBYTES[1].a/U4369  ( .A(n6631), .B(n6630), .Z(n7050) );
  XOR \SUBBYTES[1].a/U4368  ( .A(\w1[1][76] ), .B(n6632), .Z(n6630) );
  XOR \SUBBYTES[1].a/U4367  ( .A(\SUBBYTES[1].a/w1459 ), .B(\w1[1][78] ), .Z(
        n6631) );
  XOR \SUBBYTES[1].a/U4366  ( .A(\SUBBYTES[1].a/w1433 ), .B(
        \SUBBYTES[1].a/w1440 ), .Z(n6632) );
  XOR \SUBBYTES[1].a/U4365  ( .A(n6634), .B(n6633), .Z(n7048) );
  XOR \SUBBYTES[1].a/U4364  ( .A(\w1[1][73] ), .B(n6635), .Z(n6633) );
  XOR \SUBBYTES[1].a/U4363  ( .A(\SUBBYTES[1].a/w1458 ), .B(\w1[1][77] ), .Z(
        n6634) );
  XOR \SUBBYTES[1].a/U4362  ( .A(\SUBBYTES[1].a/w1434 ), .B(
        \SUBBYTES[1].a/w1441 ), .Z(n6635) );
  XOR \SUBBYTES[1].a/U4361  ( .A(n7050), .B(n7048), .Z(\SUBBYTES[1].a/w1464 )
         );
  XOR \SUBBYTES[1].a/U4360  ( .A(\w1[1][77] ), .B(n6636), .Z(n7051) );
  XOR \SUBBYTES[1].a/U4359  ( .A(\SUBBYTES[1].a/w1426 ), .B(
        \SUBBYTES[1].a/w1436 ), .Z(n6636) );
  XOR \SUBBYTES[1].a/U4358  ( .A(n6638), .B(n6637), .Z(\SUBBYTES[1].a/w1451 )
         );
  XOR \SUBBYTES[1].a/U4357  ( .A(n7051), .B(n6639), .Z(n6637) );
  XOR \SUBBYTES[1].a/U4356  ( .A(\w1[1][76] ), .B(\SUBBYTES[1].a/w1515 ), .Z(
        n6638) );
  XOR \SUBBYTES[1].a/U4355  ( .A(\SUBBYTES[1].a/w1428 ), .B(
        \SUBBYTES[1].a/w1433 ), .Z(n6639) );
  XOR \SUBBYTES[1].a/U4354  ( .A(n6641), .B(n6640), .Z(n7049) );
  XOR \SUBBYTES[1].a/U4353  ( .A(\SUBBYTES[1].a/w1461 ), .B(\w1[1][79] ), .Z(
        n6640) );
  XOR \SUBBYTES[1].a/U4352  ( .A(\SUBBYTES[1].a/w1436 ), .B(
        \SUBBYTES[1].a/w1443 ), .Z(n6641) );
  XOR \SUBBYTES[1].a/U4351  ( .A(n7048), .B(n7049), .Z(\SUBBYTES[1].a/w1463 )
         );
  XOR \SUBBYTES[1].a/U4350  ( .A(\w1[1][75] ), .B(n6642), .Z(n7052) );
  XOR \SUBBYTES[1].a/U4349  ( .A(\SUBBYTES[1].a/w1425 ), .B(
        \SUBBYTES[1].a/w1428 ), .Z(n6642) );
  XOR \SUBBYTES[1].a/U4348  ( .A(n6644), .B(n6643), .Z(\SUBBYTES[1].a/w1452 )
         );
  XOR \SUBBYTES[1].a/U4347  ( .A(n7052), .B(n6645), .Z(n6643) );
  XOR \SUBBYTES[1].a/U4346  ( .A(\w1[1][78] ), .B(\SUBBYTES[1].a/w1494 ), .Z(
        n6644) );
  XOR \SUBBYTES[1].a/U4345  ( .A(\SUBBYTES[1].a/w1433 ), .B(
        \SUBBYTES[1].a/w1434 ), .Z(n6645) );
  XOR \SUBBYTES[1].a/U4344  ( .A(n7050), .B(n7049), .Z(\SUBBYTES[1].a/w1472 )
         );
  XOR \SUBBYTES[1].a/U4343  ( .A(n6647), .B(n6646), .Z(\SUBBYTES[1].a/w1473 )
         );
  XOR \SUBBYTES[1].a/U4342  ( .A(\w1[1][79] ), .B(n7051), .Z(n6646) );
  XOR \SUBBYTES[1].a/U4341  ( .A(\SUBBYTES[1].a/w1425 ), .B(
        \SUBBYTES[1].a/w1434 ), .Z(n6647) );
  XOR \SUBBYTES[1].a/U4340  ( .A(n6649), .B(n6648), .Z(\SUBBYTES[1].a/w1449 )
         );
  XOR \SUBBYTES[1].a/U4339  ( .A(n6651), .B(n6650), .Z(n6648) );
  XOR \SUBBYTES[1].a/U4338  ( .A(\w1[1][79] ), .B(\SUBBYTES[1].a/w1533 ), .Z(
        n6649) );
  XOR \SUBBYTES[1].a/U4337  ( .A(\SUBBYTES[1].a/w1440 ), .B(
        \SUBBYTES[1].a/w1443 ), .Z(n6650) );
  XOR \SUBBYTES[1].a/U4336  ( .A(\SUBBYTES[1].a/w1426 ), .B(
        \SUBBYTES[1].a/w1428 ), .Z(n6651) );
  XOR \SUBBYTES[1].a/U4335  ( .A(n6653), .B(n6652), .Z(\SUBBYTES[1].a/w1450 )
         );
  XOR \SUBBYTES[1].a/U4334  ( .A(n7052), .B(n6654), .Z(n6652) );
  XOR \SUBBYTES[1].a/U4333  ( .A(\w1[1][77] ), .B(n7053), .Z(n6653) );
  XOR \SUBBYTES[1].a/U4332  ( .A(\SUBBYTES[1].a/w1440 ), .B(
        \SUBBYTES[1].a/w1441 ), .Z(n6654) );
  XOR \SUBBYTES[1].a/U4331  ( .A(n6656), .B(n6655), .Z(\SUBBYTES[1].a/w1466 )
         );
  XOR \SUBBYTES[1].a/U4330  ( .A(\w1[1][73] ), .B(n6657), .Z(n6655) );
  XOR \SUBBYTES[1].a/U4329  ( .A(\SUBBYTES[1].a/w1441 ), .B(
        \SUBBYTES[1].a/w1443 ), .Z(n6656) );
  XOR \SUBBYTES[1].a/U4328  ( .A(\SUBBYTES[1].a/w1425 ), .B(
        \SUBBYTES[1].a/w1426 ), .Z(n6657) );
  XOR \SUBBYTES[1].a/U4327  ( .A(\w1[1][81] ), .B(n6658), .Z(n7054) );
  XOR \SUBBYTES[1].a/U4326  ( .A(\w1[1][83] ), .B(\w1[1][82] ), .Z(n6658) );
  XOR \SUBBYTES[1].a/U4325  ( .A(\w1[1][86] ), .B(n7054), .Z(
        \SUBBYTES[1].a/w1308 ) );
  XOR \SUBBYTES[1].a/U4324  ( .A(\w1[1][80] ), .B(\SUBBYTES[1].a/w1308 ), .Z(
        \SUBBYTES[1].a/w1195 ) );
  XOR \SUBBYTES[1].a/U4323  ( .A(\w1[1][80] ), .B(n6659), .Z(
        \SUBBYTES[1].a/w1196 ) );
  XOR \SUBBYTES[1].a/U4322  ( .A(\w1[1][86] ), .B(\w1[1][85] ), .Z(n6659) );
  XOR \SUBBYTES[1].a/U4321  ( .A(\w1[1][85] ), .B(n7054), .Z(
        \SUBBYTES[1].a/w1326 ) );
  XOR \SUBBYTES[1].a/U4320  ( .A(n6661), .B(n6660), .Z(\SUBBYTES[1].a/w1319 )
         );
  XOR \SUBBYTES[1].a/U4319  ( .A(\w1[1][83] ), .B(\w1[1][81] ), .Z(n6660) );
  XOR \SUBBYTES[1].a/U4318  ( .A(\w1[1][87] ), .B(\w1[1][84] ), .Z(n6661) );
  XOR \SUBBYTES[1].a/U4317  ( .A(\w1[1][80] ), .B(\SUBBYTES[1].a/w1319 ), .Z(
        \SUBBYTES[1].a/w1198 ) );
  XOR \SUBBYTES[1].a/U4316  ( .A(n6663), .B(n6662), .Z(\SUBBYTES[1].a/w1306 )
         );
  XOR \SUBBYTES[1].a/U4315  ( .A(\SUBBYTES[1].a/w1267 ), .B(n962), .Z(n6662)
         );
  XOR \SUBBYTES[1].a/U4314  ( .A(\SUBBYTES[1].a/w1260 ), .B(
        \SUBBYTES[1].a/w1263 ), .Z(n6663) );
  XOR \SUBBYTES[1].a/U4313  ( .A(n6665), .B(n6664), .Z(\SUBBYTES[1].a/w1307 )
         );
  XOR \SUBBYTES[1].a/U4312  ( .A(\SUBBYTES[1].a/w1267 ), .B(n5843), .Z(n6664)
         );
  XOR \SUBBYTES[1].a/U4311  ( .A(\SUBBYTES[1].a/w1260 ), .B(n5842), .Z(n6665)
         );
  XOR \SUBBYTES[1].a/U4310  ( .A(\SUBBYTES[1].a/w1319 ), .B(n6666), .Z(
        \SUBBYTES[1].a/w1309 ) );
  XOR \SUBBYTES[1].a/U4309  ( .A(\w1[1][86] ), .B(\w1[1][85] ), .Z(n6666) );
  XOR \SUBBYTES[1].a/U4308  ( .A(n6668), .B(n6667), .Z(\SUBBYTES[1].a/w1310 )
         );
  XOR \SUBBYTES[1].a/U4307  ( .A(n5843), .B(n962), .Z(n6667) );
  XOR \SUBBYTES[1].a/U4306  ( .A(n5842), .B(\SUBBYTES[1].a/w1263 ), .Z(n6668)
         );
  XOR \SUBBYTES[1].a/U4305  ( .A(\w1[1][87] ), .B(\w1[1][82] ), .Z(n7060) );
  XOR \SUBBYTES[1].a/U4304  ( .A(n7060), .B(n6669), .Z(\SUBBYTES[1].a/w1311 )
         );
  XOR \SUBBYTES[1].a/U4303  ( .A(\w1[1][85] ), .B(\w1[1][84] ), .Z(n6669) );
  XOR \SUBBYTES[1].a/U4302  ( .A(\w1[1][87] ), .B(\SUBBYTES[1].a/w1196 ), .Z(
        \SUBBYTES[1].a/w1199 ) );
  XOR \SUBBYTES[1].a/U4301  ( .A(\w1[1][81] ), .B(\SUBBYTES[1].a/w1196 ), .Z(
        \SUBBYTES[1].a/w1200 ) );
  XOR \SUBBYTES[1].a/U4300  ( .A(\w1[1][84] ), .B(\SUBBYTES[1].a/w1196 ), .Z(
        \SUBBYTES[1].a/w1201 ) );
  XOR \SUBBYTES[1].a/U4299  ( .A(\SUBBYTES[1].a/w1200 ), .B(n7060), .Z(
        \SUBBYTES[1].a/w1202 ) );
  XOR \SUBBYTES[1].a/U4298  ( .A(n7060), .B(n6670), .Z(\SUBBYTES[1].a/w1287 )
         );
  XOR \SUBBYTES[1].a/U4297  ( .A(\w1[1][84] ), .B(\w1[1][81] ), .Z(n6670) );
  XOR \SUBBYTES[1].a/U4296  ( .A(n6672), .B(n6671), .Z(n7057) );
  XOR \SUBBYTES[1].a/U4295  ( .A(\w1[1][84] ), .B(n6673), .Z(n6671) );
  XOR \SUBBYTES[1].a/U4294  ( .A(\SUBBYTES[1].a/w1252 ), .B(\w1[1][86] ), .Z(
        n6672) );
  XOR \SUBBYTES[1].a/U4293  ( .A(\SUBBYTES[1].a/w1226 ), .B(
        \SUBBYTES[1].a/w1233 ), .Z(n6673) );
  XOR \SUBBYTES[1].a/U4292  ( .A(n6675), .B(n6674), .Z(n7055) );
  XOR \SUBBYTES[1].a/U4291  ( .A(\w1[1][81] ), .B(n6676), .Z(n6674) );
  XOR \SUBBYTES[1].a/U4290  ( .A(\SUBBYTES[1].a/w1251 ), .B(\w1[1][85] ), .Z(
        n6675) );
  XOR \SUBBYTES[1].a/U4289  ( .A(\SUBBYTES[1].a/w1227 ), .B(
        \SUBBYTES[1].a/w1234 ), .Z(n6676) );
  XOR \SUBBYTES[1].a/U4288  ( .A(n7057), .B(n7055), .Z(\SUBBYTES[1].a/w1257 )
         );
  XOR \SUBBYTES[1].a/U4287  ( .A(\w1[1][85] ), .B(n6677), .Z(n7058) );
  XOR \SUBBYTES[1].a/U4286  ( .A(\SUBBYTES[1].a/w1219 ), .B(
        \SUBBYTES[1].a/w1229 ), .Z(n6677) );
  XOR \SUBBYTES[1].a/U4285  ( .A(n6679), .B(n6678), .Z(\SUBBYTES[1].a/w1244 )
         );
  XOR \SUBBYTES[1].a/U4284  ( .A(n7058), .B(n6680), .Z(n6678) );
  XOR \SUBBYTES[1].a/U4283  ( .A(\w1[1][84] ), .B(\SUBBYTES[1].a/w1308 ), .Z(
        n6679) );
  XOR \SUBBYTES[1].a/U4282  ( .A(\SUBBYTES[1].a/w1221 ), .B(
        \SUBBYTES[1].a/w1226 ), .Z(n6680) );
  XOR \SUBBYTES[1].a/U4281  ( .A(n6682), .B(n6681), .Z(n7056) );
  XOR \SUBBYTES[1].a/U4280  ( .A(\SUBBYTES[1].a/w1254 ), .B(\w1[1][87] ), .Z(
        n6681) );
  XOR \SUBBYTES[1].a/U4279  ( .A(\SUBBYTES[1].a/w1229 ), .B(
        \SUBBYTES[1].a/w1236 ), .Z(n6682) );
  XOR \SUBBYTES[1].a/U4278  ( .A(n7055), .B(n7056), .Z(\SUBBYTES[1].a/w1256 )
         );
  XOR \SUBBYTES[1].a/U4277  ( .A(\w1[1][83] ), .B(n6683), .Z(n7059) );
  XOR \SUBBYTES[1].a/U4276  ( .A(\SUBBYTES[1].a/w1218 ), .B(
        \SUBBYTES[1].a/w1221 ), .Z(n6683) );
  XOR \SUBBYTES[1].a/U4275  ( .A(n6685), .B(n6684), .Z(\SUBBYTES[1].a/w1245 )
         );
  XOR \SUBBYTES[1].a/U4274  ( .A(n7059), .B(n6686), .Z(n6684) );
  XOR \SUBBYTES[1].a/U4273  ( .A(\w1[1][86] ), .B(\SUBBYTES[1].a/w1287 ), .Z(
        n6685) );
  XOR \SUBBYTES[1].a/U4272  ( .A(\SUBBYTES[1].a/w1226 ), .B(
        \SUBBYTES[1].a/w1227 ), .Z(n6686) );
  XOR \SUBBYTES[1].a/U4271  ( .A(n7057), .B(n7056), .Z(\SUBBYTES[1].a/w1265 )
         );
  XOR \SUBBYTES[1].a/U4270  ( .A(n6688), .B(n6687), .Z(\SUBBYTES[1].a/w1266 )
         );
  XOR \SUBBYTES[1].a/U4269  ( .A(\w1[1][87] ), .B(n7058), .Z(n6687) );
  XOR \SUBBYTES[1].a/U4268  ( .A(\SUBBYTES[1].a/w1218 ), .B(
        \SUBBYTES[1].a/w1227 ), .Z(n6688) );
  XOR \SUBBYTES[1].a/U4267  ( .A(n6690), .B(n6689), .Z(\SUBBYTES[1].a/w1242 )
         );
  XOR \SUBBYTES[1].a/U4266  ( .A(n6692), .B(n6691), .Z(n6689) );
  XOR \SUBBYTES[1].a/U4265  ( .A(\w1[1][87] ), .B(\SUBBYTES[1].a/w1326 ), .Z(
        n6690) );
  XOR \SUBBYTES[1].a/U4264  ( .A(\SUBBYTES[1].a/w1233 ), .B(
        \SUBBYTES[1].a/w1236 ), .Z(n6691) );
  XOR \SUBBYTES[1].a/U4263  ( .A(\SUBBYTES[1].a/w1219 ), .B(
        \SUBBYTES[1].a/w1221 ), .Z(n6692) );
  XOR \SUBBYTES[1].a/U4262  ( .A(n6694), .B(n6693), .Z(\SUBBYTES[1].a/w1243 )
         );
  XOR \SUBBYTES[1].a/U4261  ( .A(n7059), .B(n6695), .Z(n6693) );
  XOR \SUBBYTES[1].a/U4260  ( .A(\w1[1][85] ), .B(n7060), .Z(n6694) );
  XOR \SUBBYTES[1].a/U4259  ( .A(\SUBBYTES[1].a/w1233 ), .B(
        \SUBBYTES[1].a/w1234 ), .Z(n6695) );
  XOR \SUBBYTES[1].a/U4258  ( .A(n6697), .B(n6696), .Z(\SUBBYTES[1].a/w1259 )
         );
  XOR \SUBBYTES[1].a/U4257  ( .A(\w1[1][81] ), .B(n6698), .Z(n6696) );
  XOR \SUBBYTES[1].a/U4256  ( .A(\SUBBYTES[1].a/w1234 ), .B(
        \SUBBYTES[1].a/w1236 ), .Z(n6697) );
  XOR \SUBBYTES[1].a/U4255  ( .A(\SUBBYTES[1].a/w1218 ), .B(
        \SUBBYTES[1].a/w1219 ), .Z(n6698) );
  XOR \SUBBYTES[1].a/U4254  ( .A(\w1[1][89] ), .B(n6699), .Z(n7061) );
  XOR \SUBBYTES[1].a/U4253  ( .A(\w1[1][91] ), .B(\w1[1][90] ), .Z(n6699) );
  XOR \SUBBYTES[1].a/U4252  ( .A(\w1[1][94] ), .B(n7061), .Z(
        \SUBBYTES[1].a/w1101 ) );
  XOR \SUBBYTES[1].a/U4251  ( .A(\w1[1][88] ), .B(\SUBBYTES[1].a/w1101 ), .Z(
        \SUBBYTES[1].a/w988 ) );
  XOR \SUBBYTES[1].a/U4250  ( .A(\w1[1][88] ), .B(n6700), .Z(
        \SUBBYTES[1].a/w989 ) );
  XOR \SUBBYTES[1].a/U4249  ( .A(\w1[1][94] ), .B(\w1[1][93] ), .Z(n6700) );
  XOR \SUBBYTES[1].a/U4248  ( .A(\w1[1][93] ), .B(n7061), .Z(
        \SUBBYTES[1].a/w1119 ) );
  XOR \SUBBYTES[1].a/U4247  ( .A(n6702), .B(n6701), .Z(\SUBBYTES[1].a/w1112 )
         );
  XOR \SUBBYTES[1].a/U4246  ( .A(\w1[1][91] ), .B(\w1[1][89] ), .Z(n6701) );
  XOR \SUBBYTES[1].a/U4245  ( .A(\w1[1][95] ), .B(\w1[1][92] ), .Z(n6702) );
  XOR \SUBBYTES[1].a/U4244  ( .A(\w1[1][88] ), .B(\SUBBYTES[1].a/w1112 ), .Z(
        \SUBBYTES[1].a/w991 ) );
  XOR \SUBBYTES[1].a/U4243  ( .A(n6704), .B(n6703), .Z(\SUBBYTES[1].a/w1099 )
         );
  XOR \SUBBYTES[1].a/U4242  ( .A(\SUBBYTES[1].a/w1060 ), .B(n961), .Z(n6703)
         );
  XOR \SUBBYTES[1].a/U4241  ( .A(\SUBBYTES[1].a/w1053 ), .B(
        \SUBBYTES[1].a/w1056 ), .Z(n6704) );
  XOR \SUBBYTES[1].a/U4240  ( .A(n6706), .B(n6705), .Z(\SUBBYTES[1].a/w1100 )
         );
  XOR \SUBBYTES[1].a/U4239  ( .A(\SUBBYTES[1].a/w1060 ), .B(n5841), .Z(n6705)
         );
  XOR \SUBBYTES[1].a/U4238  ( .A(\SUBBYTES[1].a/w1053 ), .B(n5840), .Z(n6706)
         );
  XOR \SUBBYTES[1].a/U4237  ( .A(\SUBBYTES[1].a/w1112 ), .B(n6707), .Z(
        \SUBBYTES[1].a/w1102 ) );
  XOR \SUBBYTES[1].a/U4236  ( .A(\w1[1][94] ), .B(\w1[1][93] ), .Z(n6707) );
  XOR \SUBBYTES[1].a/U4235  ( .A(n6709), .B(n6708), .Z(\SUBBYTES[1].a/w1103 )
         );
  XOR \SUBBYTES[1].a/U4234  ( .A(n5841), .B(n961), .Z(n6708) );
  XOR \SUBBYTES[1].a/U4233  ( .A(n5840), .B(\SUBBYTES[1].a/w1056 ), .Z(n6709)
         );
  XOR \SUBBYTES[1].a/U4232  ( .A(\w1[1][95] ), .B(\w1[1][90] ), .Z(n7067) );
  XOR \SUBBYTES[1].a/U4231  ( .A(n7067), .B(n6710), .Z(\SUBBYTES[1].a/w1104 )
         );
  XOR \SUBBYTES[1].a/U4230  ( .A(\w1[1][93] ), .B(\w1[1][92] ), .Z(n6710) );
  XOR \SUBBYTES[1].a/U4229  ( .A(\w1[1][95] ), .B(\SUBBYTES[1].a/w989 ), .Z(
        \SUBBYTES[1].a/w992 ) );
  XOR \SUBBYTES[1].a/U4228  ( .A(\w1[1][89] ), .B(\SUBBYTES[1].a/w989 ), .Z(
        \SUBBYTES[1].a/w993 ) );
  XOR \SUBBYTES[1].a/U4227  ( .A(\w1[1][92] ), .B(\SUBBYTES[1].a/w989 ), .Z(
        \SUBBYTES[1].a/w994 ) );
  XOR \SUBBYTES[1].a/U4226  ( .A(\SUBBYTES[1].a/w993 ), .B(n7067), .Z(
        \SUBBYTES[1].a/w995 ) );
  XOR \SUBBYTES[1].a/U4225  ( .A(n7067), .B(n6711), .Z(\SUBBYTES[1].a/w1080 )
         );
  XOR \SUBBYTES[1].a/U4224  ( .A(\w1[1][92] ), .B(\w1[1][89] ), .Z(n6711) );
  XOR \SUBBYTES[1].a/U4223  ( .A(n6713), .B(n6712), .Z(n7064) );
  XOR \SUBBYTES[1].a/U4222  ( .A(\w1[1][92] ), .B(n6714), .Z(n6712) );
  XOR \SUBBYTES[1].a/U4221  ( .A(\SUBBYTES[1].a/w1045 ), .B(\w1[1][94] ), .Z(
        n6713) );
  XOR \SUBBYTES[1].a/U4220  ( .A(\SUBBYTES[1].a/w1019 ), .B(
        \SUBBYTES[1].a/w1026 ), .Z(n6714) );
  XOR \SUBBYTES[1].a/U4219  ( .A(n6716), .B(n6715), .Z(n7062) );
  XOR \SUBBYTES[1].a/U4218  ( .A(\w1[1][89] ), .B(n6717), .Z(n6715) );
  XOR \SUBBYTES[1].a/U4217  ( .A(\SUBBYTES[1].a/w1044 ), .B(\w1[1][93] ), .Z(
        n6716) );
  XOR \SUBBYTES[1].a/U4216  ( .A(\SUBBYTES[1].a/w1020 ), .B(
        \SUBBYTES[1].a/w1027 ), .Z(n6717) );
  XOR \SUBBYTES[1].a/U4215  ( .A(n7064), .B(n7062), .Z(\SUBBYTES[1].a/w1050 )
         );
  XOR \SUBBYTES[1].a/U4214  ( .A(\w1[1][93] ), .B(n6718), .Z(n7065) );
  XOR \SUBBYTES[1].a/U4213  ( .A(\SUBBYTES[1].a/w1012 ), .B(
        \SUBBYTES[1].a/w1022 ), .Z(n6718) );
  XOR \SUBBYTES[1].a/U4212  ( .A(n6720), .B(n6719), .Z(\SUBBYTES[1].a/w1037 )
         );
  XOR \SUBBYTES[1].a/U4211  ( .A(n7065), .B(n6721), .Z(n6719) );
  XOR \SUBBYTES[1].a/U4210  ( .A(\w1[1][92] ), .B(\SUBBYTES[1].a/w1101 ), .Z(
        n6720) );
  XOR \SUBBYTES[1].a/U4209  ( .A(\SUBBYTES[1].a/w1014 ), .B(
        \SUBBYTES[1].a/w1019 ), .Z(n6721) );
  XOR \SUBBYTES[1].a/U4208  ( .A(n6723), .B(n6722), .Z(n7063) );
  XOR \SUBBYTES[1].a/U4207  ( .A(\SUBBYTES[1].a/w1047 ), .B(\w1[1][95] ), .Z(
        n6722) );
  XOR \SUBBYTES[1].a/U4206  ( .A(\SUBBYTES[1].a/w1022 ), .B(
        \SUBBYTES[1].a/w1029 ), .Z(n6723) );
  XOR \SUBBYTES[1].a/U4205  ( .A(n7062), .B(n7063), .Z(\SUBBYTES[1].a/w1049 )
         );
  XOR \SUBBYTES[1].a/U4204  ( .A(\w1[1][91] ), .B(n6724), .Z(n7066) );
  XOR \SUBBYTES[1].a/U4203  ( .A(\SUBBYTES[1].a/w1011 ), .B(
        \SUBBYTES[1].a/w1014 ), .Z(n6724) );
  XOR \SUBBYTES[1].a/U4202  ( .A(n6726), .B(n6725), .Z(\SUBBYTES[1].a/w1038 )
         );
  XOR \SUBBYTES[1].a/U4201  ( .A(n7066), .B(n6727), .Z(n6725) );
  XOR \SUBBYTES[1].a/U4200  ( .A(\w1[1][94] ), .B(\SUBBYTES[1].a/w1080 ), .Z(
        n6726) );
  XOR \SUBBYTES[1].a/U4199  ( .A(\SUBBYTES[1].a/w1019 ), .B(
        \SUBBYTES[1].a/w1020 ), .Z(n6727) );
  XOR \SUBBYTES[1].a/U4198  ( .A(n7064), .B(n7063), .Z(\SUBBYTES[1].a/w1058 )
         );
  XOR \SUBBYTES[1].a/U4197  ( .A(n6729), .B(n6728), .Z(\SUBBYTES[1].a/w1059 )
         );
  XOR \SUBBYTES[1].a/U4196  ( .A(\w1[1][95] ), .B(n7065), .Z(n6728) );
  XOR \SUBBYTES[1].a/U4195  ( .A(\SUBBYTES[1].a/w1011 ), .B(
        \SUBBYTES[1].a/w1020 ), .Z(n6729) );
  XOR \SUBBYTES[1].a/U4194  ( .A(n6731), .B(n6730), .Z(\SUBBYTES[1].a/w1035 )
         );
  XOR \SUBBYTES[1].a/U4193  ( .A(n6733), .B(n6732), .Z(n6730) );
  XOR \SUBBYTES[1].a/U4192  ( .A(\w1[1][95] ), .B(\SUBBYTES[1].a/w1119 ), .Z(
        n6731) );
  XOR \SUBBYTES[1].a/U4191  ( .A(\SUBBYTES[1].a/w1026 ), .B(
        \SUBBYTES[1].a/w1029 ), .Z(n6732) );
  XOR \SUBBYTES[1].a/U4190  ( .A(\SUBBYTES[1].a/w1012 ), .B(
        \SUBBYTES[1].a/w1014 ), .Z(n6733) );
  XOR \SUBBYTES[1].a/U4189  ( .A(n6735), .B(n6734), .Z(\SUBBYTES[1].a/w1036 )
         );
  XOR \SUBBYTES[1].a/U4188  ( .A(n7066), .B(n6736), .Z(n6734) );
  XOR \SUBBYTES[1].a/U4187  ( .A(\w1[1][93] ), .B(n7067), .Z(n6735) );
  XOR \SUBBYTES[1].a/U4186  ( .A(\SUBBYTES[1].a/w1026 ), .B(
        \SUBBYTES[1].a/w1027 ), .Z(n6736) );
  XOR \SUBBYTES[1].a/U4185  ( .A(n6738), .B(n6737), .Z(\SUBBYTES[1].a/w1052 )
         );
  XOR \SUBBYTES[1].a/U4184  ( .A(\w1[1][89] ), .B(n6739), .Z(n6737) );
  XOR \SUBBYTES[1].a/U4183  ( .A(\SUBBYTES[1].a/w1027 ), .B(
        \SUBBYTES[1].a/w1029 ), .Z(n6738) );
  XOR \SUBBYTES[1].a/U4182  ( .A(\SUBBYTES[1].a/w1011 ), .B(
        \SUBBYTES[1].a/w1012 ), .Z(n6739) );
  XOR \SUBBYTES[1].a/U4181  ( .A(\w1[1][97] ), .B(n6740), .Z(n7068) );
  XOR \SUBBYTES[1].a/U4180  ( .A(\w1[1][99] ), .B(\w1[1][98] ), .Z(n6740) );
  XOR \SUBBYTES[1].a/U4179  ( .A(\w1[1][102] ), .B(n7068), .Z(
        \SUBBYTES[1].a/w894 ) );
  XOR \SUBBYTES[1].a/U4178  ( .A(\w1[1][96] ), .B(\SUBBYTES[1].a/w894 ), .Z(
        \SUBBYTES[1].a/w781 ) );
  XOR \SUBBYTES[1].a/U4177  ( .A(\w1[1][96] ), .B(n6741), .Z(
        \SUBBYTES[1].a/w782 ) );
  XOR \SUBBYTES[1].a/U4176  ( .A(\w1[1][102] ), .B(\w1[1][101] ), .Z(n6741) );
  XOR \SUBBYTES[1].a/U4175  ( .A(\w1[1][101] ), .B(n7068), .Z(
        \SUBBYTES[1].a/w912 ) );
  XOR \SUBBYTES[1].a/U4174  ( .A(n6743), .B(n6742), .Z(\SUBBYTES[1].a/w905 )
         );
  XOR \SUBBYTES[1].a/U4173  ( .A(\w1[1][99] ), .B(\w1[1][97] ), .Z(n6742) );
  XOR \SUBBYTES[1].a/U4172  ( .A(\w1[1][103] ), .B(\w1[1][100] ), .Z(n6743) );
  XOR \SUBBYTES[1].a/U4171  ( .A(\w1[1][96] ), .B(\SUBBYTES[1].a/w905 ), .Z(
        \SUBBYTES[1].a/w784 ) );
  XOR \SUBBYTES[1].a/U4170  ( .A(n6745), .B(n6744), .Z(\SUBBYTES[1].a/w892 )
         );
  XOR \SUBBYTES[1].a/U4169  ( .A(\SUBBYTES[1].a/w853 ), .B(n960), .Z(n6744) );
  XOR \SUBBYTES[1].a/U4168  ( .A(\SUBBYTES[1].a/w846 ), .B(
        \SUBBYTES[1].a/w849 ), .Z(n6745) );
  XOR \SUBBYTES[1].a/U4167  ( .A(n6747), .B(n6746), .Z(\SUBBYTES[1].a/w893 )
         );
  XOR \SUBBYTES[1].a/U4166  ( .A(\SUBBYTES[1].a/w853 ), .B(n5839), .Z(n6746)
         );
  XOR \SUBBYTES[1].a/U4165  ( .A(\SUBBYTES[1].a/w846 ), .B(n5838), .Z(n6747)
         );
  XOR \SUBBYTES[1].a/U4164  ( .A(\SUBBYTES[1].a/w905 ), .B(n6748), .Z(
        \SUBBYTES[1].a/w895 ) );
  XOR \SUBBYTES[1].a/U4163  ( .A(\w1[1][102] ), .B(\w1[1][101] ), .Z(n6748) );
  XOR \SUBBYTES[1].a/U4162  ( .A(n6750), .B(n6749), .Z(\SUBBYTES[1].a/w896 )
         );
  XOR \SUBBYTES[1].a/U4161  ( .A(n5839), .B(n960), .Z(n6749) );
  XOR \SUBBYTES[1].a/U4160  ( .A(n5838), .B(\SUBBYTES[1].a/w849 ), .Z(n6750)
         );
  XOR \SUBBYTES[1].a/U4159  ( .A(\w1[1][103] ), .B(\w1[1][98] ), .Z(n7074) );
  XOR \SUBBYTES[1].a/U4158  ( .A(n7074), .B(n6751), .Z(\SUBBYTES[1].a/w897 )
         );
  XOR \SUBBYTES[1].a/U4157  ( .A(\w1[1][101] ), .B(\w1[1][100] ), .Z(n6751) );
  XOR \SUBBYTES[1].a/U4156  ( .A(\w1[1][103] ), .B(\SUBBYTES[1].a/w782 ), .Z(
        \SUBBYTES[1].a/w785 ) );
  XOR \SUBBYTES[1].a/U4155  ( .A(\w1[1][97] ), .B(\SUBBYTES[1].a/w782 ), .Z(
        \SUBBYTES[1].a/w786 ) );
  XOR \SUBBYTES[1].a/U4154  ( .A(\w1[1][100] ), .B(\SUBBYTES[1].a/w782 ), .Z(
        \SUBBYTES[1].a/w787 ) );
  XOR \SUBBYTES[1].a/U4153  ( .A(\SUBBYTES[1].a/w786 ), .B(n7074), .Z(
        \SUBBYTES[1].a/w788 ) );
  XOR \SUBBYTES[1].a/U4152  ( .A(n7074), .B(n6752), .Z(\SUBBYTES[1].a/w873 )
         );
  XOR \SUBBYTES[1].a/U4151  ( .A(\w1[1][100] ), .B(\w1[1][97] ), .Z(n6752) );
  XOR \SUBBYTES[1].a/U4150  ( .A(n6754), .B(n6753), .Z(n7071) );
  XOR \SUBBYTES[1].a/U4149  ( .A(\w1[1][100] ), .B(n6755), .Z(n6753) );
  XOR \SUBBYTES[1].a/U4148  ( .A(\SUBBYTES[1].a/w838 ), .B(\w1[1][102] ), .Z(
        n6754) );
  XOR \SUBBYTES[1].a/U4147  ( .A(\SUBBYTES[1].a/w812 ), .B(
        \SUBBYTES[1].a/w819 ), .Z(n6755) );
  XOR \SUBBYTES[1].a/U4146  ( .A(n6757), .B(n6756), .Z(n7069) );
  XOR \SUBBYTES[1].a/U4145  ( .A(\w1[1][97] ), .B(n6758), .Z(n6756) );
  XOR \SUBBYTES[1].a/U4144  ( .A(\SUBBYTES[1].a/w837 ), .B(\w1[1][101] ), .Z(
        n6757) );
  XOR \SUBBYTES[1].a/U4143  ( .A(\SUBBYTES[1].a/w813 ), .B(
        \SUBBYTES[1].a/w820 ), .Z(n6758) );
  XOR \SUBBYTES[1].a/U4142  ( .A(n7071), .B(n7069), .Z(\SUBBYTES[1].a/w843 )
         );
  XOR \SUBBYTES[1].a/U4141  ( .A(\w1[1][101] ), .B(n6759), .Z(n7072) );
  XOR \SUBBYTES[1].a/U4140  ( .A(\SUBBYTES[1].a/w805 ), .B(
        \SUBBYTES[1].a/w815 ), .Z(n6759) );
  XOR \SUBBYTES[1].a/U4139  ( .A(n6761), .B(n6760), .Z(\SUBBYTES[1].a/w830 )
         );
  XOR \SUBBYTES[1].a/U4138  ( .A(n7072), .B(n6762), .Z(n6760) );
  XOR \SUBBYTES[1].a/U4137  ( .A(\w1[1][100] ), .B(\SUBBYTES[1].a/w894 ), .Z(
        n6761) );
  XOR \SUBBYTES[1].a/U4136  ( .A(\SUBBYTES[1].a/w807 ), .B(
        \SUBBYTES[1].a/w812 ), .Z(n6762) );
  XOR \SUBBYTES[1].a/U4135  ( .A(n6764), .B(n6763), .Z(n7070) );
  XOR \SUBBYTES[1].a/U4134  ( .A(\SUBBYTES[1].a/w840 ), .B(\w1[1][103] ), .Z(
        n6763) );
  XOR \SUBBYTES[1].a/U4133  ( .A(\SUBBYTES[1].a/w815 ), .B(
        \SUBBYTES[1].a/w822 ), .Z(n6764) );
  XOR \SUBBYTES[1].a/U4132  ( .A(n7069), .B(n7070), .Z(\SUBBYTES[1].a/w842 )
         );
  XOR \SUBBYTES[1].a/U4131  ( .A(\w1[1][99] ), .B(n6765), .Z(n7073) );
  XOR \SUBBYTES[1].a/U4130  ( .A(\SUBBYTES[1].a/w804 ), .B(
        \SUBBYTES[1].a/w807 ), .Z(n6765) );
  XOR \SUBBYTES[1].a/U4129  ( .A(n6767), .B(n6766), .Z(\SUBBYTES[1].a/w831 )
         );
  XOR \SUBBYTES[1].a/U4128  ( .A(n7073), .B(n6768), .Z(n6766) );
  XOR \SUBBYTES[1].a/U4127  ( .A(\w1[1][102] ), .B(\SUBBYTES[1].a/w873 ), .Z(
        n6767) );
  XOR \SUBBYTES[1].a/U4126  ( .A(\SUBBYTES[1].a/w812 ), .B(
        \SUBBYTES[1].a/w813 ), .Z(n6768) );
  XOR \SUBBYTES[1].a/U4125  ( .A(n7071), .B(n7070), .Z(\SUBBYTES[1].a/w851 )
         );
  XOR \SUBBYTES[1].a/U4124  ( .A(n6770), .B(n6769), .Z(\SUBBYTES[1].a/w852 )
         );
  XOR \SUBBYTES[1].a/U4123  ( .A(\w1[1][103] ), .B(n7072), .Z(n6769) );
  XOR \SUBBYTES[1].a/U4122  ( .A(\SUBBYTES[1].a/w804 ), .B(
        \SUBBYTES[1].a/w813 ), .Z(n6770) );
  XOR \SUBBYTES[1].a/U4121  ( .A(n6772), .B(n6771), .Z(\SUBBYTES[1].a/w828 )
         );
  XOR \SUBBYTES[1].a/U4120  ( .A(n6774), .B(n6773), .Z(n6771) );
  XOR \SUBBYTES[1].a/U4119  ( .A(\w1[1][103] ), .B(\SUBBYTES[1].a/w912 ), .Z(
        n6772) );
  XOR \SUBBYTES[1].a/U4118  ( .A(\SUBBYTES[1].a/w819 ), .B(
        \SUBBYTES[1].a/w822 ), .Z(n6773) );
  XOR \SUBBYTES[1].a/U4117  ( .A(\SUBBYTES[1].a/w805 ), .B(
        \SUBBYTES[1].a/w807 ), .Z(n6774) );
  XOR \SUBBYTES[1].a/U4116  ( .A(n6776), .B(n6775), .Z(\SUBBYTES[1].a/w829 )
         );
  XOR \SUBBYTES[1].a/U4115  ( .A(n7073), .B(n6777), .Z(n6775) );
  XOR \SUBBYTES[1].a/U4114  ( .A(\w1[1][101] ), .B(n7074), .Z(n6776) );
  XOR \SUBBYTES[1].a/U4113  ( .A(\SUBBYTES[1].a/w819 ), .B(
        \SUBBYTES[1].a/w820 ), .Z(n6777) );
  XOR \SUBBYTES[1].a/U4112  ( .A(n6779), .B(n6778), .Z(\SUBBYTES[1].a/w845 )
         );
  XOR \SUBBYTES[1].a/U4111  ( .A(\w1[1][97] ), .B(n6780), .Z(n6778) );
  XOR \SUBBYTES[1].a/U4110  ( .A(\SUBBYTES[1].a/w820 ), .B(
        \SUBBYTES[1].a/w822 ), .Z(n6779) );
  XOR \SUBBYTES[1].a/U4109  ( .A(\SUBBYTES[1].a/w804 ), .B(
        \SUBBYTES[1].a/w805 ), .Z(n6780) );
  XOR \SUBBYTES[1].a/U4108  ( .A(\w1[1][105] ), .B(n6781), .Z(n7075) );
  XOR \SUBBYTES[1].a/U4107  ( .A(\w1[1][107] ), .B(\w1[1][106] ), .Z(n6781) );
  XOR \SUBBYTES[1].a/U4106  ( .A(\w1[1][110] ), .B(n7075), .Z(
        \SUBBYTES[1].a/w687 ) );
  XOR \SUBBYTES[1].a/U4105  ( .A(\w1[1][104] ), .B(\SUBBYTES[1].a/w687 ), .Z(
        \SUBBYTES[1].a/w574 ) );
  XOR \SUBBYTES[1].a/U4104  ( .A(\w1[1][104] ), .B(n6782), .Z(
        \SUBBYTES[1].a/w575 ) );
  XOR \SUBBYTES[1].a/U4103  ( .A(\w1[1][110] ), .B(\w1[1][109] ), .Z(n6782) );
  XOR \SUBBYTES[1].a/U4102  ( .A(\w1[1][109] ), .B(n7075), .Z(
        \SUBBYTES[1].a/w705 ) );
  XOR \SUBBYTES[1].a/U4101  ( .A(n6784), .B(n6783), .Z(\SUBBYTES[1].a/w698 )
         );
  XOR \SUBBYTES[1].a/U4100  ( .A(\w1[1][107] ), .B(\w1[1][105] ), .Z(n6783) );
  XOR \SUBBYTES[1].a/U4099  ( .A(\w1[1][111] ), .B(\w1[1][108] ), .Z(n6784) );
  XOR \SUBBYTES[1].a/U4098  ( .A(\w1[1][104] ), .B(\SUBBYTES[1].a/w698 ), .Z(
        \SUBBYTES[1].a/w577 ) );
  XOR \SUBBYTES[1].a/U4097  ( .A(n6786), .B(n6785), .Z(\SUBBYTES[1].a/w685 )
         );
  XOR \SUBBYTES[1].a/U4096  ( .A(\SUBBYTES[1].a/w646 ), .B(n959), .Z(n6785) );
  XOR \SUBBYTES[1].a/U4095  ( .A(\SUBBYTES[1].a/w639 ), .B(
        \SUBBYTES[1].a/w642 ), .Z(n6786) );
  XOR \SUBBYTES[1].a/U4094  ( .A(n6788), .B(n6787), .Z(\SUBBYTES[1].a/w686 )
         );
  XOR \SUBBYTES[1].a/U4093  ( .A(\SUBBYTES[1].a/w646 ), .B(n5837), .Z(n6787)
         );
  XOR \SUBBYTES[1].a/U4092  ( .A(\SUBBYTES[1].a/w639 ), .B(n5836), .Z(n6788)
         );
  XOR \SUBBYTES[1].a/U4091  ( .A(\SUBBYTES[1].a/w698 ), .B(n6789), .Z(
        \SUBBYTES[1].a/w688 ) );
  XOR \SUBBYTES[1].a/U4090  ( .A(\w1[1][110] ), .B(\w1[1][109] ), .Z(n6789) );
  XOR \SUBBYTES[1].a/U4089  ( .A(n6791), .B(n6790), .Z(\SUBBYTES[1].a/w689 )
         );
  XOR \SUBBYTES[1].a/U4088  ( .A(n5837), .B(n959), .Z(n6790) );
  XOR \SUBBYTES[1].a/U4087  ( .A(n5836), .B(\SUBBYTES[1].a/w642 ), .Z(n6791)
         );
  XOR \SUBBYTES[1].a/U4086  ( .A(\w1[1][111] ), .B(\w1[1][106] ), .Z(n7081) );
  XOR \SUBBYTES[1].a/U4085  ( .A(n7081), .B(n6792), .Z(\SUBBYTES[1].a/w690 )
         );
  XOR \SUBBYTES[1].a/U4084  ( .A(\w1[1][109] ), .B(\w1[1][108] ), .Z(n6792) );
  XOR \SUBBYTES[1].a/U4083  ( .A(\w1[1][111] ), .B(\SUBBYTES[1].a/w575 ), .Z(
        \SUBBYTES[1].a/w578 ) );
  XOR \SUBBYTES[1].a/U4082  ( .A(\w1[1][105] ), .B(\SUBBYTES[1].a/w575 ), .Z(
        \SUBBYTES[1].a/w579 ) );
  XOR \SUBBYTES[1].a/U4081  ( .A(\w1[1][108] ), .B(\SUBBYTES[1].a/w575 ), .Z(
        \SUBBYTES[1].a/w580 ) );
  XOR \SUBBYTES[1].a/U4080  ( .A(\SUBBYTES[1].a/w579 ), .B(n7081), .Z(
        \SUBBYTES[1].a/w581 ) );
  XOR \SUBBYTES[1].a/U4079  ( .A(n7081), .B(n6793), .Z(\SUBBYTES[1].a/w666 )
         );
  XOR \SUBBYTES[1].a/U4078  ( .A(\w1[1][108] ), .B(\w1[1][105] ), .Z(n6793) );
  XOR \SUBBYTES[1].a/U4077  ( .A(n6795), .B(n6794), .Z(n7078) );
  XOR \SUBBYTES[1].a/U4076  ( .A(\w1[1][108] ), .B(n6796), .Z(n6794) );
  XOR \SUBBYTES[1].a/U4075  ( .A(\SUBBYTES[1].a/w631 ), .B(\w1[1][110] ), .Z(
        n6795) );
  XOR \SUBBYTES[1].a/U4074  ( .A(\SUBBYTES[1].a/w605 ), .B(
        \SUBBYTES[1].a/w612 ), .Z(n6796) );
  XOR \SUBBYTES[1].a/U4073  ( .A(n6798), .B(n6797), .Z(n7076) );
  XOR \SUBBYTES[1].a/U4072  ( .A(\w1[1][105] ), .B(n6799), .Z(n6797) );
  XOR \SUBBYTES[1].a/U4071  ( .A(\SUBBYTES[1].a/w630 ), .B(\w1[1][109] ), .Z(
        n6798) );
  XOR \SUBBYTES[1].a/U4070  ( .A(\SUBBYTES[1].a/w606 ), .B(
        \SUBBYTES[1].a/w613 ), .Z(n6799) );
  XOR \SUBBYTES[1].a/U4069  ( .A(n7078), .B(n7076), .Z(\SUBBYTES[1].a/w636 )
         );
  XOR \SUBBYTES[1].a/U4068  ( .A(\w1[1][109] ), .B(n6800), .Z(n7079) );
  XOR \SUBBYTES[1].a/U4067  ( .A(\SUBBYTES[1].a/w598 ), .B(
        \SUBBYTES[1].a/w608 ), .Z(n6800) );
  XOR \SUBBYTES[1].a/U4066  ( .A(n6802), .B(n6801), .Z(\SUBBYTES[1].a/w623 )
         );
  XOR \SUBBYTES[1].a/U4065  ( .A(n7079), .B(n6803), .Z(n6801) );
  XOR \SUBBYTES[1].a/U4064  ( .A(\w1[1][108] ), .B(\SUBBYTES[1].a/w687 ), .Z(
        n6802) );
  XOR \SUBBYTES[1].a/U4063  ( .A(\SUBBYTES[1].a/w600 ), .B(
        \SUBBYTES[1].a/w605 ), .Z(n6803) );
  XOR \SUBBYTES[1].a/U4062  ( .A(n6805), .B(n6804), .Z(n7077) );
  XOR \SUBBYTES[1].a/U4061  ( .A(\SUBBYTES[1].a/w633 ), .B(\w1[1][111] ), .Z(
        n6804) );
  XOR \SUBBYTES[1].a/U4060  ( .A(\SUBBYTES[1].a/w608 ), .B(
        \SUBBYTES[1].a/w615 ), .Z(n6805) );
  XOR \SUBBYTES[1].a/U4059  ( .A(n7076), .B(n7077), .Z(\SUBBYTES[1].a/w635 )
         );
  XOR \SUBBYTES[1].a/U4058  ( .A(\w1[1][107] ), .B(n6806), .Z(n7080) );
  XOR \SUBBYTES[1].a/U4057  ( .A(\SUBBYTES[1].a/w597 ), .B(
        \SUBBYTES[1].a/w600 ), .Z(n6806) );
  XOR \SUBBYTES[1].a/U4056  ( .A(n6808), .B(n6807), .Z(\SUBBYTES[1].a/w624 )
         );
  XOR \SUBBYTES[1].a/U4055  ( .A(n7080), .B(n6809), .Z(n6807) );
  XOR \SUBBYTES[1].a/U4054  ( .A(\w1[1][110] ), .B(\SUBBYTES[1].a/w666 ), .Z(
        n6808) );
  XOR \SUBBYTES[1].a/U4053  ( .A(\SUBBYTES[1].a/w605 ), .B(
        \SUBBYTES[1].a/w606 ), .Z(n6809) );
  XOR \SUBBYTES[1].a/U4052  ( .A(n7078), .B(n7077), .Z(\SUBBYTES[1].a/w644 )
         );
  XOR \SUBBYTES[1].a/U4051  ( .A(n6811), .B(n6810), .Z(\SUBBYTES[1].a/w645 )
         );
  XOR \SUBBYTES[1].a/U4050  ( .A(\w1[1][111] ), .B(n7079), .Z(n6810) );
  XOR \SUBBYTES[1].a/U4049  ( .A(\SUBBYTES[1].a/w597 ), .B(
        \SUBBYTES[1].a/w606 ), .Z(n6811) );
  XOR \SUBBYTES[1].a/U4048  ( .A(n6813), .B(n6812), .Z(\SUBBYTES[1].a/w621 )
         );
  XOR \SUBBYTES[1].a/U4047  ( .A(n6815), .B(n6814), .Z(n6812) );
  XOR \SUBBYTES[1].a/U4046  ( .A(\w1[1][111] ), .B(\SUBBYTES[1].a/w705 ), .Z(
        n6813) );
  XOR \SUBBYTES[1].a/U4045  ( .A(\SUBBYTES[1].a/w612 ), .B(
        \SUBBYTES[1].a/w615 ), .Z(n6814) );
  XOR \SUBBYTES[1].a/U4044  ( .A(\SUBBYTES[1].a/w598 ), .B(
        \SUBBYTES[1].a/w600 ), .Z(n6815) );
  XOR \SUBBYTES[1].a/U4043  ( .A(n6817), .B(n6816), .Z(\SUBBYTES[1].a/w622 )
         );
  XOR \SUBBYTES[1].a/U4042  ( .A(n7080), .B(n6818), .Z(n6816) );
  XOR \SUBBYTES[1].a/U4041  ( .A(\w1[1][109] ), .B(n7081), .Z(n6817) );
  XOR \SUBBYTES[1].a/U4040  ( .A(\SUBBYTES[1].a/w612 ), .B(
        \SUBBYTES[1].a/w613 ), .Z(n6818) );
  XOR \SUBBYTES[1].a/U4039  ( .A(n6820), .B(n6819), .Z(\SUBBYTES[1].a/w638 )
         );
  XOR \SUBBYTES[1].a/U4038  ( .A(\w1[1][105] ), .B(n6821), .Z(n6819) );
  XOR \SUBBYTES[1].a/U4037  ( .A(\SUBBYTES[1].a/w613 ), .B(
        \SUBBYTES[1].a/w615 ), .Z(n6820) );
  XOR \SUBBYTES[1].a/U4036  ( .A(\SUBBYTES[1].a/w597 ), .B(
        \SUBBYTES[1].a/w598 ), .Z(n6821) );
  XOR \SUBBYTES[1].a/U4035  ( .A(\w1[1][113] ), .B(n6822), .Z(n7082) );
  XOR \SUBBYTES[1].a/U4034  ( .A(\w1[1][115] ), .B(\w1[1][114] ), .Z(n6822) );
  XOR \SUBBYTES[1].a/U4033  ( .A(\w1[1][118] ), .B(n7082), .Z(
        \SUBBYTES[1].a/w480 ) );
  XOR \SUBBYTES[1].a/U4032  ( .A(\w1[1][112] ), .B(\SUBBYTES[1].a/w480 ), .Z(
        \SUBBYTES[1].a/w367 ) );
  XOR \SUBBYTES[1].a/U4031  ( .A(\w1[1][112] ), .B(n6823), .Z(
        \SUBBYTES[1].a/w368 ) );
  XOR \SUBBYTES[1].a/U4030  ( .A(\w1[1][118] ), .B(\w1[1][117] ), .Z(n6823) );
  XOR \SUBBYTES[1].a/U4029  ( .A(\w1[1][117] ), .B(n7082), .Z(
        \SUBBYTES[1].a/w498 ) );
  XOR \SUBBYTES[1].a/U4028  ( .A(n6825), .B(n6824), .Z(\SUBBYTES[1].a/w491 )
         );
  XOR \SUBBYTES[1].a/U4027  ( .A(\w1[1][115] ), .B(\w1[1][113] ), .Z(n6824) );
  XOR \SUBBYTES[1].a/U4026  ( .A(\w1[1][119] ), .B(\w1[1][116] ), .Z(n6825) );
  XOR \SUBBYTES[1].a/U4025  ( .A(\w1[1][112] ), .B(\SUBBYTES[1].a/w491 ), .Z(
        \SUBBYTES[1].a/w370 ) );
  XOR \SUBBYTES[1].a/U4024  ( .A(n6827), .B(n6826), .Z(\SUBBYTES[1].a/w478 )
         );
  XOR \SUBBYTES[1].a/U4023  ( .A(\SUBBYTES[1].a/w439 ), .B(n958), .Z(n6826) );
  XOR \SUBBYTES[1].a/U4022  ( .A(\SUBBYTES[1].a/w432 ), .B(
        \SUBBYTES[1].a/w435 ), .Z(n6827) );
  XOR \SUBBYTES[1].a/U4021  ( .A(n6829), .B(n6828), .Z(\SUBBYTES[1].a/w479 )
         );
  XOR \SUBBYTES[1].a/U4020  ( .A(\SUBBYTES[1].a/w439 ), .B(n5835), .Z(n6828)
         );
  XOR \SUBBYTES[1].a/U4019  ( .A(\SUBBYTES[1].a/w432 ), .B(n5834), .Z(n6829)
         );
  XOR \SUBBYTES[1].a/U4018  ( .A(\SUBBYTES[1].a/w491 ), .B(n6830), .Z(
        \SUBBYTES[1].a/w481 ) );
  XOR \SUBBYTES[1].a/U4017  ( .A(\w1[1][118] ), .B(\w1[1][117] ), .Z(n6830) );
  XOR \SUBBYTES[1].a/U4016  ( .A(n6832), .B(n6831), .Z(\SUBBYTES[1].a/w482 )
         );
  XOR \SUBBYTES[1].a/U4015  ( .A(n5835), .B(n958), .Z(n6831) );
  XOR \SUBBYTES[1].a/U4014  ( .A(n5834), .B(\SUBBYTES[1].a/w435 ), .Z(n6832)
         );
  XOR \SUBBYTES[1].a/U4013  ( .A(\w1[1][119] ), .B(\w1[1][114] ), .Z(n7088) );
  XOR \SUBBYTES[1].a/U4012  ( .A(n7088), .B(n6833), .Z(\SUBBYTES[1].a/w483 )
         );
  XOR \SUBBYTES[1].a/U4011  ( .A(\w1[1][117] ), .B(\w1[1][116] ), .Z(n6833) );
  XOR \SUBBYTES[1].a/U4010  ( .A(\w1[1][119] ), .B(\SUBBYTES[1].a/w368 ), .Z(
        \SUBBYTES[1].a/w371 ) );
  XOR \SUBBYTES[1].a/U4009  ( .A(\w1[1][113] ), .B(\SUBBYTES[1].a/w368 ), .Z(
        \SUBBYTES[1].a/w372 ) );
  XOR \SUBBYTES[1].a/U4008  ( .A(\w1[1][116] ), .B(\SUBBYTES[1].a/w368 ), .Z(
        \SUBBYTES[1].a/w373 ) );
  XOR \SUBBYTES[1].a/U4007  ( .A(\SUBBYTES[1].a/w372 ), .B(n7088), .Z(
        \SUBBYTES[1].a/w374 ) );
  XOR \SUBBYTES[1].a/U4006  ( .A(n7088), .B(n6834), .Z(\SUBBYTES[1].a/w459 )
         );
  XOR \SUBBYTES[1].a/U4005  ( .A(\w1[1][116] ), .B(\w1[1][113] ), .Z(n6834) );
  XOR \SUBBYTES[1].a/U4004  ( .A(n6836), .B(n6835), .Z(n7085) );
  XOR \SUBBYTES[1].a/U4003  ( .A(\w1[1][116] ), .B(n6837), .Z(n6835) );
  XOR \SUBBYTES[1].a/U4002  ( .A(\SUBBYTES[1].a/w424 ), .B(\w1[1][118] ), .Z(
        n6836) );
  XOR \SUBBYTES[1].a/U4001  ( .A(\SUBBYTES[1].a/w398 ), .B(
        \SUBBYTES[1].a/w405 ), .Z(n6837) );
  XOR \SUBBYTES[1].a/U4000  ( .A(n6839), .B(n6838), .Z(n7083) );
  XOR \SUBBYTES[1].a/U3999  ( .A(\w1[1][113] ), .B(n6840), .Z(n6838) );
  XOR \SUBBYTES[1].a/U3998  ( .A(\SUBBYTES[1].a/w423 ), .B(\w1[1][117] ), .Z(
        n6839) );
  XOR \SUBBYTES[1].a/U3997  ( .A(\SUBBYTES[1].a/w399 ), .B(
        \SUBBYTES[1].a/w406 ), .Z(n6840) );
  XOR \SUBBYTES[1].a/U3996  ( .A(n7085), .B(n7083), .Z(\SUBBYTES[1].a/w429 )
         );
  XOR \SUBBYTES[1].a/U3995  ( .A(\w1[1][117] ), .B(n6841), .Z(n7086) );
  XOR \SUBBYTES[1].a/U3994  ( .A(\SUBBYTES[1].a/w391 ), .B(
        \SUBBYTES[1].a/w401 ), .Z(n6841) );
  XOR \SUBBYTES[1].a/U3993  ( .A(n6843), .B(n6842), .Z(\SUBBYTES[1].a/w416 )
         );
  XOR \SUBBYTES[1].a/U3992  ( .A(n7086), .B(n6844), .Z(n6842) );
  XOR \SUBBYTES[1].a/U3991  ( .A(\w1[1][116] ), .B(\SUBBYTES[1].a/w480 ), .Z(
        n6843) );
  XOR \SUBBYTES[1].a/U3990  ( .A(\SUBBYTES[1].a/w393 ), .B(
        \SUBBYTES[1].a/w398 ), .Z(n6844) );
  XOR \SUBBYTES[1].a/U3989  ( .A(n6846), .B(n6845), .Z(n7084) );
  XOR \SUBBYTES[1].a/U3988  ( .A(\SUBBYTES[1].a/w426 ), .B(\w1[1][119] ), .Z(
        n6845) );
  XOR \SUBBYTES[1].a/U3987  ( .A(\SUBBYTES[1].a/w401 ), .B(
        \SUBBYTES[1].a/w408 ), .Z(n6846) );
  XOR \SUBBYTES[1].a/U3986  ( .A(n7083), .B(n7084), .Z(\SUBBYTES[1].a/w428 )
         );
  XOR \SUBBYTES[1].a/U3985  ( .A(\w1[1][115] ), .B(n6847), .Z(n7087) );
  XOR \SUBBYTES[1].a/U3984  ( .A(\SUBBYTES[1].a/w390 ), .B(
        \SUBBYTES[1].a/w393 ), .Z(n6847) );
  XOR \SUBBYTES[1].a/U3983  ( .A(n6849), .B(n6848), .Z(\SUBBYTES[1].a/w417 )
         );
  XOR \SUBBYTES[1].a/U3982  ( .A(n7087), .B(n6850), .Z(n6848) );
  XOR \SUBBYTES[1].a/U3981  ( .A(\w1[1][118] ), .B(\SUBBYTES[1].a/w459 ), .Z(
        n6849) );
  XOR \SUBBYTES[1].a/U3980  ( .A(\SUBBYTES[1].a/w398 ), .B(
        \SUBBYTES[1].a/w399 ), .Z(n6850) );
  XOR \SUBBYTES[1].a/U3979  ( .A(n7085), .B(n7084), .Z(\SUBBYTES[1].a/w437 )
         );
  XOR \SUBBYTES[1].a/U3978  ( .A(n6852), .B(n6851), .Z(\SUBBYTES[1].a/w438 )
         );
  XOR \SUBBYTES[1].a/U3977  ( .A(\w1[1][119] ), .B(n7086), .Z(n6851) );
  XOR \SUBBYTES[1].a/U3976  ( .A(\SUBBYTES[1].a/w390 ), .B(
        \SUBBYTES[1].a/w399 ), .Z(n6852) );
  XOR \SUBBYTES[1].a/U3975  ( .A(n6854), .B(n6853), .Z(\SUBBYTES[1].a/w414 )
         );
  XOR \SUBBYTES[1].a/U3974  ( .A(n6856), .B(n6855), .Z(n6853) );
  XOR \SUBBYTES[1].a/U3973  ( .A(\w1[1][119] ), .B(\SUBBYTES[1].a/w498 ), .Z(
        n6854) );
  XOR \SUBBYTES[1].a/U3972  ( .A(\SUBBYTES[1].a/w405 ), .B(
        \SUBBYTES[1].a/w408 ), .Z(n6855) );
  XOR \SUBBYTES[1].a/U3971  ( .A(\SUBBYTES[1].a/w391 ), .B(
        \SUBBYTES[1].a/w393 ), .Z(n6856) );
  XOR \SUBBYTES[1].a/U3970  ( .A(n6858), .B(n6857), .Z(\SUBBYTES[1].a/w415 )
         );
  XOR \SUBBYTES[1].a/U3969  ( .A(n7087), .B(n6859), .Z(n6857) );
  XOR \SUBBYTES[1].a/U3968  ( .A(\w1[1][117] ), .B(n7088), .Z(n6858) );
  XOR \SUBBYTES[1].a/U3967  ( .A(\SUBBYTES[1].a/w405 ), .B(
        \SUBBYTES[1].a/w406 ), .Z(n6859) );
  XOR \SUBBYTES[1].a/U3966  ( .A(n6861), .B(n6860), .Z(\SUBBYTES[1].a/w431 )
         );
  XOR \SUBBYTES[1].a/U3965  ( .A(\w1[1][113] ), .B(n6862), .Z(n6860) );
  XOR \SUBBYTES[1].a/U3964  ( .A(\SUBBYTES[1].a/w406 ), .B(
        \SUBBYTES[1].a/w408 ), .Z(n6861) );
  XOR \SUBBYTES[1].a/U3963  ( .A(\SUBBYTES[1].a/w390 ), .B(
        \SUBBYTES[1].a/w391 ), .Z(n6862) );
  XOR \SUBBYTES[1].a/U3962  ( .A(\w1[1][121] ), .B(n6863), .Z(n7089) );
  XOR \SUBBYTES[1].a/U3961  ( .A(\w1[1][123] ), .B(\w1[1][122] ), .Z(n6863) );
  XOR \SUBBYTES[1].a/U3960  ( .A(\w1[1][126] ), .B(n7089), .Z(
        \SUBBYTES[1].a/w273 ) );
  XOR \SUBBYTES[1].a/U3959  ( .A(\w1[1][120] ), .B(\SUBBYTES[1].a/w273 ), .Z(
        \SUBBYTES[1].a/w160 ) );
  XOR \SUBBYTES[1].a/U3958  ( .A(\w1[1][120] ), .B(n6864), .Z(
        \SUBBYTES[1].a/w161 ) );
  XOR \SUBBYTES[1].a/U3957  ( .A(\w1[1][126] ), .B(\w1[1][125] ), .Z(n6864) );
  XOR \SUBBYTES[1].a/U3956  ( .A(\w1[1][125] ), .B(n7089), .Z(
        \SUBBYTES[1].a/w291 ) );
  XOR \SUBBYTES[1].a/U3955  ( .A(n6866), .B(n6865), .Z(\SUBBYTES[1].a/w284 )
         );
  XOR \SUBBYTES[1].a/U3954  ( .A(\w1[1][123] ), .B(\w1[1][121] ), .Z(n6865) );
  XOR \SUBBYTES[1].a/U3953  ( .A(\w1[1][127] ), .B(\w1[1][124] ), .Z(n6866) );
  XOR \SUBBYTES[1].a/U3952  ( .A(\w1[1][120] ), .B(\SUBBYTES[1].a/w284 ), .Z(
        \SUBBYTES[1].a/w163 ) );
  XOR \SUBBYTES[1].a/U3951  ( .A(n6868), .B(n6867), .Z(\SUBBYTES[1].a/w271 )
         );
  XOR \SUBBYTES[1].a/U3950  ( .A(\SUBBYTES[1].a/w232 ), .B(n957), .Z(n6867) );
  XOR \SUBBYTES[1].a/U3949  ( .A(\SUBBYTES[1].a/w225 ), .B(
        \SUBBYTES[1].a/w228 ), .Z(n6868) );
  XOR \SUBBYTES[1].a/U3948  ( .A(n6870), .B(n6869), .Z(\SUBBYTES[1].a/w272 )
         );
  XOR \SUBBYTES[1].a/U3947  ( .A(\SUBBYTES[1].a/w232 ), .B(n5833), .Z(n6869)
         );
  XOR \SUBBYTES[1].a/U3946  ( .A(\SUBBYTES[1].a/w225 ), .B(n5832), .Z(n6870)
         );
  XOR \SUBBYTES[1].a/U3945  ( .A(\SUBBYTES[1].a/w284 ), .B(n6871), .Z(
        \SUBBYTES[1].a/w274 ) );
  XOR \SUBBYTES[1].a/U3944  ( .A(\w1[1][126] ), .B(\w1[1][125] ), .Z(n6871) );
  XOR \SUBBYTES[1].a/U3943  ( .A(n6873), .B(n6872), .Z(\SUBBYTES[1].a/w275 )
         );
  XOR \SUBBYTES[1].a/U3942  ( .A(n5833), .B(n957), .Z(n6872) );
  XOR \SUBBYTES[1].a/U3941  ( .A(n5832), .B(\SUBBYTES[1].a/w228 ), .Z(n6873)
         );
  XOR \SUBBYTES[1].a/U3940  ( .A(\w1[1][127] ), .B(\w1[1][122] ), .Z(n7095) );
  XOR \SUBBYTES[1].a/U3939  ( .A(n7095), .B(n6874), .Z(\SUBBYTES[1].a/w276 )
         );
  XOR \SUBBYTES[1].a/U3938  ( .A(\w1[1][125] ), .B(\w1[1][124] ), .Z(n6874) );
  XOR \SUBBYTES[1].a/U3937  ( .A(\w1[1][127] ), .B(\SUBBYTES[1].a/w161 ), .Z(
        \SUBBYTES[1].a/w164 ) );
  XOR \SUBBYTES[1].a/U3936  ( .A(\w1[1][121] ), .B(\SUBBYTES[1].a/w161 ), .Z(
        \SUBBYTES[1].a/w165 ) );
  XOR \SUBBYTES[1].a/U3935  ( .A(\w1[1][124] ), .B(\SUBBYTES[1].a/w161 ), .Z(
        \SUBBYTES[1].a/w166 ) );
  XOR \SUBBYTES[1].a/U3934  ( .A(\SUBBYTES[1].a/w165 ), .B(n7095), .Z(
        \SUBBYTES[1].a/w167 ) );
  XOR \SUBBYTES[1].a/U3933  ( .A(n7095), .B(n6875), .Z(\SUBBYTES[1].a/w252 )
         );
  XOR \SUBBYTES[1].a/U3932  ( .A(\w1[1][124] ), .B(\w1[1][121] ), .Z(n6875) );
  XOR \SUBBYTES[1].a/U3931  ( .A(n6877), .B(n6876), .Z(n7092) );
  XOR \SUBBYTES[1].a/U3930  ( .A(\w1[1][124] ), .B(n6878), .Z(n6876) );
  XOR \SUBBYTES[1].a/U3929  ( .A(\SUBBYTES[1].a/w217 ), .B(\w1[1][126] ), .Z(
        n6877) );
  XOR \SUBBYTES[1].a/U3928  ( .A(\SUBBYTES[1].a/w191 ), .B(
        \SUBBYTES[1].a/w198 ), .Z(n6878) );
  XOR \SUBBYTES[1].a/U3927  ( .A(n6880), .B(n6879), .Z(n7090) );
  XOR \SUBBYTES[1].a/U3926  ( .A(\w1[1][121] ), .B(n6881), .Z(n6879) );
  XOR \SUBBYTES[1].a/U3925  ( .A(\SUBBYTES[1].a/w216 ), .B(\w1[1][125] ), .Z(
        n6880) );
  XOR \SUBBYTES[1].a/U3924  ( .A(\SUBBYTES[1].a/w192 ), .B(
        \SUBBYTES[1].a/w199 ), .Z(n6881) );
  XOR \SUBBYTES[1].a/U3923  ( .A(n7092), .B(n7090), .Z(\SUBBYTES[1].a/w222 )
         );
  XOR \SUBBYTES[1].a/U3922  ( .A(\w1[1][125] ), .B(n6882), .Z(n7093) );
  XOR \SUBBYTES[1].a/U3921  ( .A(\SUBBYTES[1].a/w184 ), .B(
        \SUBBYTES[1].a/w194 ), .Z(n6882) );
  XOR \SUBBYTES[1].a/U3920  ( .A(n6884), .B(n6883), .Z(\SUBBYTES[1].a/w209 )
         );
  XOR \SUBBYTES[1].a/U3919  ( .A(n7093), .B(n6885), .Z(n6883) );
  XOR \SUBBYTES[1].a/U3918  ( .A(\w1[1][124] ), .B(\SUBBYTES[1].a/w273 ), .Z(
        n6884) );
  XOR \SUBBYTES[1].a/U3917  ( .A(\SUBBYTES[1].a/w186 ), .B(
        \SUBBYTES[1].a/w191 ), .Z(n6885) );
  XOR \SUBBYTES[1].a/U3916  ( .A(n6887), .B(n6886), .Z(n7091) );
  XOR \SUBBYTES[1].a/U3915  ( .A(\SUBBYTES[1].a/w219 ), .B(\w1[1][127] ), .Z(
        n6886) );
  XOR \SUBBYTES[1].a/U3914  ( .A(\SUBBYTES[1].a/w194 ), .B(
        \SUBBYTES[1].a/w201 ), .Z(n6887) );
  XOR \SUBBYTES[1].a/U3913  ( .A(n7090), .B(n7091), .Z(\SUBBYTES[1].a/w221 )
         );
  XOR \SUBBYTES[1].a/U3912  ( .A(\w1[1][123] ), .B(n6888), .Z(n7094) );
  XOR \SUBBYTES[1].a/U3911  ( .A(\SUBBYTES[1].a/w183 ), .B(
        \SUBBYTES[1].a/w186 ), .Z(n6888) );
  XOR \SUBBYTES[1].a/U3910  ( .A(n6890), .B(n6889), .Z(\SUBBYTES[1].a/w210 )
         );
  XOR \SUBBYTES[1].a/U3909  ( .A(n7094), .B(n6891), .Z(n6889) );
  XOR \SUBBYTES[1].a/U3908  ( .A(\w1[1][126] ), .B(\SUBBYTES[1].a/w252 ), .Z(
        n6890) );
  XOR \SUBBYTES[1].a/U3907  ( .A(\SUBBYTES[1].a/w191 ), .B(
        \SUBBYTES[1].a/w192 ), .Z(n6891) );
  XOR \SUBBYTES[1].a/U3906  ( .A(n7092), .B(n7091), .Z(\SUBBYTES[1].a/w230 )
         );
  XOR \SUBBYTES[1].a/U3905  ( .A(n6893), .B(n6892), .Z(\SUBBYTES[1].a/w231 )
         );
  XOR \SUBBYTES[1].a/U3904  ( .A(\w1[1][127] ), .B(n7093), .Z(n6892) );
  XOR \SUBBYTES[1].a/U3903  ( .A(\SUBBYTES[1].a/w183 ), .B(
        \SUBBYTES[1].a/w192 ), .Z(n6893) );
  XOR \SUBBYTES[1].a/U3902  ( .A(n6895), .B(n6894), .Z(\SUBBYTES[1].a/w207 )
         );
  XOR \SUBBYTES[1].a/U3901  ( .A(n6897), .B(n6896), .Z(n6894) );
  XOR \SUBBYTES[1].a/U3900  ( .A(\w1[1][127] ), .B(\SUBBYTES[1].a/w291 ), .Z(
        n6895) );
  XOR \SUBBYTES[1].a/U3899  ( .A(\SUBBYTES[1].a/w198 ), .B(
        \SUBBYTES[1].a/w201 ), .Z(n6896) );
  XOR \SUBBYTES[1].a/U3898  ( .A(\SUBBYTES[1].a/w184 ), .B(
        \SUBBYTES[1].a/w186 ), .Z(n6897) );
  XOR \SUBBYTES[1].a/U3897  ( .A(n6899), .B(n6898), .Z(\SUBBYTES[1].a/w208 )
         );
  XOR \SUBBYTES[1].a/U3896  ( .A(n7094), .B(n6900), .Z(n6898) );
  XOR \SUBBYTES[1].a/U3895  ( .A(\w1[1][125] ), .B(n7095), .Z(n6899) );
  XOR \SUBBYTES[1].a/U3894  ( .A(\SUBBYTES[1].a/w198 ), .B(
        \SUBBYTES[1].a/w199 ), .Z(n6900) );
  XOR \SUBBYTES[1].a/U3893  ( .A(n6902), .B(n6901), .Z(\SUBBYTES[1].a/w224 )
         );
  XOR \SUBBYTES[1].a/U3892  ( .A(\w1[1][121] ), .B(n6903), .Z(n6901) );
  XOR \SUBBYTES[1].a/U3891  ( .A(\SUBBYTES[1].a/w199 ), .B(
        \SUBBYTES[1].a/w201 ), .Z(n6902) );
  XOR \SUBBYTES[1].a/U3890  ( .A(\SUBBYTES[1].a/w183 ), .B(
        \SUBBYTES[1].a/w184 ), .Z(n6903) );
  XOR \MIXCOLUMNS[8].d/U432  ( .A(n956), .B(n484), .Z(n5777) );
  XOR \MIXCOLUMNS[8].d/U431  ( .A(n5529), .B(n5528), .Z(\w0[9][0] ) );
  XOR \MIXCOLUMNS[8].d/U430  ( .A(n955), .B(n5777), .Z(n5528) );
  XOR \MIXCOLUMNS[8].d/U429  ( .A(n954), .B(n32), .Z(n5529) );
  XOR \MIXCOLUMNS[8].d/U428  ( .A(n954), .B(n483), .Z(n5762) );
  XOR \MIXCOLUMNS[8].d/U427  ( .A(n5531), .B(n5530), .Z(\w0[9][1] ) );
  XOR \MIXCOLUMNS[8].d/U426  ( .A(\w3[8][2] ), .B(n5762), .Z(n5530) );
  XOR \MIXCOLUMNS[8].d/U425  ( .A(\w3[8][26] ), .B(n482), .Z(n5531) );
  XOR \MIXCOLUMNS[8].d/U424  ( .A(\w3[8][26] ), .B(\w3[8][18] ), .Z(n5765) );
  XOR \MIXCOLUMNS[8].d/U423  ( .A(n5533), .B(n5532), .Z(\w0[9][2] ) );
  XOR \MIXCOLUMNS[8].d/U422  ( .A(n953), .B(n5765), .Z(n5532) );
  XOR \MIXCOLUMNS[8].d/U421  ( .A(n952), .B(\w3[8][10] ), .Z(n5533) );
  XOR \MIXCOLUMNS[8].d/U420  ( .A(n956), .B(n481), .Z(n5760) );
  XOR \MIXCOLUMNS[8].d/U419  ( .A(n952), .B(n480), .Z(n5767) );
  XOR \MIXCOLUMNS[8].d/U418  ( .A(n5535), .B(n5534), .Z(\w0[9][3] ) );
  XOR \MIXCOLUMNS[8].d/U417  ( .A(n5767), .B(n5536), .Z(n5534) );
  XOR \MIXCOLUMNS[8].d/U416  ( .A(n951), .B(n5760), .Z(n5535) );
  XOR \MIXCOLUMNS[8].d/U415  ( .A(n950), .B(n479), .Z(n5536) );
  XOR \MIXCOLUMNS[8].d/U414  ( .A(n950), .B(n478), .Z(n5769) );
  XOR \MIXCOLUMNS[8].d/U413  ( .A(n5538), .B(n5537), .Z(\w0[9][4] ) );
  XOR \MIXCOLUMNS[8].d/U412  ( .A(n5769), .B(n5539), .Z(n5537) );
  XOR \MIXCOLUMNS[8].d/U411  ( .A(n949), .B(n5760), .Z(n5538) );
  XOR \MIXCOLUMNS[8].d/U410  ( .A(n948), .B(n477), .Z(n5539) );
  XOR \MIXCOLUMNS[8].d/U409  ( .A(n948), .B(n476), .Z(n5771) );
  XOR \MIXCOLUMNS[8].d/U408  ( .A(n5541), .B(n5540), .Z(\w0[9][5] ) );
  XOR \MIXCOLUMNS[8].d/U407  ( .A(n947), .B(n5771), .Z(n5540) );
  XOR \MIXCOLUMNS[8].d/U406  ( .A(n946), .B(n475), .Z(n5541) );
  XOR \MIXCOLUMNS[8].d/U405  ( .A(n946), .B(n474), .Z(n5773) );
  XOR \MIXCOLUMNS[8].d/U404  ( .A(n5543), .B(n5542), .Z(\w0[9][6] ) );
  XOR \MIXCOLUMNS[8].d/U403  ( .A(n5773), .B(n5544), .Z(n5542) );
  XOR \MIXCOLUMNS[8].d/U402  ( .A(n945), .B(n5760), .Z(n5543) );
  XOR \MIXCOLUMNS[8].d/U401  ( .A(n944), .B(n473), .Z(n5544) );
  XOR \MIXCOLUMNS[8].d/U400  ( .A(n944), .B(n472), .Z(n5775) );
  XOR \MIXCOLUMNS[8].d/U399  ( .A(n5775), .B(n5545), .Z(\w0[9][7] ) );
  XOR \MIXCOLUMNS[8].d/U398  ( .A(n471), .B(n5760), .Z(n5545) );
  XOR \MIXCOLUMNS[8].d/U397  ( .A(n482), .B(n955), .Z(n5764) );
  XOR \MIXCOLUMNS[8].d/U396  ( .A(n5764), .B(n5546), .Z(\w0[9][8] ) );
  XOR \MIXCOLUMNS[8].d/U395  ( .A(n481), .B(n5777), .Z(n5546) );
  XOR \MIXCOLUMNS[8].d/U394  ( .A(\w3[8][10] ), .B(\w3[8][2] ), .Z(n5766) );
  XOR \MIXCOLUMNS[8].d/U393  ( .A(n5766), .B(n5547), .Z(\w0[9][9] ) );
  XOR \MIXCOLUMNS[8].d/U392  ( .A(n955), .B(n5762), .Z(n5547) );
  XOR \MIXCOLUMNS[8].d/U391  ( .A(n479), .B(n953), .Z(n5768) );
  XOR \MIXCOLUMNS[8].d/U390  ( .A(n5768), .B(n5548), .Z(\w0[9][10] ) );
  XOR \MIXCOLUMNS[8].d/U389  ( .A(\w3[8][2] ), .B(n5765), .Z(n5548) );
  XOR \MIXCOLUMNS[8].d/U388  ( .A(n32), .B(n481), .Z(n5763) );
  XOR \MIXCOLUMNS[8].d/U387  ( .A(n477), .B(n951), .Z(n5770) );
  XOR \MIXCOLUMNS[8].d/U386  ( .A(n5550), .B(n5549), .Z(\w0[9][11] ) );
  XOR \MIXCOLUMNS[8].d/U385  ( .A(n5767), .B(n5770), .Z(n5549) );
  XOR \MIXCOLUMNS[8].d/U384  ( .A(n953), .B(n5763), .Z(n5550) );
  XOR \MIXCOLUMNS[8].d/U383  ( .A(n475), .B(n949), .Z(n5772) );
  XOR \MIXCOLUMNS[8].d/U382  ( .A(n5552), .B(n5551), .Z(\w0[9][12] ) );
  XOR \MIXCOLUMNS[8].d/U381  ( .A(n5769), .B(n5772), .Z(n5551) );
  XOR \MIXCOLUMNS[8].d/U380  ( .A(n951), .B(n5763), .Z(n5552) );
  XOR \MIXCOLUMNS[8].d/U379  ( .A(n473), .B(n947), .Z(n5774) );
  XOR \MIXCOLUMNS[8].d/U378  ( .A(n5774), .B(n5553), .Z(\w0[9][13] ) );
  XOR \MIXCOLUMNS[8].d/U377  ( .A(n949), .B(n5771), .Z(n5553) );
  XOR \MIXCOLUMNS[8].d/U376  ( .A(n471), .B(n945), .Z(n5776) );
  XOR \MIXCOLUMNS[8].d/U375  ( .A(n5555), .B(n5554), .Z(\w0[9][14] ) );
  XOR \MIXCOLUMNS[8].d/U374  ( .A(n5773), .B(n5776), .Z(n5554) );
  XOR \MIXCOLUMNS[8].d/U373  ( .A(n947), .B(n5763), .Z(n5555) );
  XOR \MIXCOLUMNS[8].d/U372  ( .A(n5775), .B(n5556), .Z(\w0[9][15] ) );
  XOR \MIXCOLUMNS[8].d/U371  ( .A(n945), .B(n5763), .Z(n5556) );
  XOR \MIXCOLUMNS[8].d/U370  ( .A(n5558), .B(n5557), .Z(\w0[9][16] ) );
  XOR \MIXCOLUMNS[8].d/U369  ( .A(n482), .B(n5763), .Z(n5557) );
  XOR \MIXCOLUMNS[8].d/U368  ( .A(n956), .B(n483), .Z(n5558) );
  XOR \MIXCOLUMNS[8].d/U367  ( .A(n5560), .B(n5559), .Z(\w0[9][17] ) );
  XOR \MIXCOLUMNS[8].d/U366  ( .A(\w3[8][10] ), .B(n5764), .Z(n5559) );
  XOR \MIXCOLUMNS[8].d/U365  ( .A(n954), .B(\w3[8][18] ), .Z(n5560) );
  XOR \MIXCOLUMNS[8].d/U364  ( .A(n5562), .B(n5561), .Z(\w0[9][18] ) );
  XOR \MIXCOLUMNS[8].d/U363  ( .A(n479), .B(n5766), .Z(n5561) );
  XOR \MIXCOLUMNS[8].d/U362  ( .A(\w3[8][26] ), .B(n480), .Z(n5562) );
  XOR \MIXCOLUMNS[8].d/U361  ( .A(n484), .B(n32), .Z(n5761) );
  XOR \MIXCOLUMNS[8].d/U360  ( .A(n5564), .B(n5563), .Z(\w0[9][19] ) );
  XOR \MIXCOLUMNS[8].d/U359  ( .A(n5768), .B(n5565), .Z(n5563) );
  XOR \MIXCOLUMNS[8].d/U358  ( .A(n477), .B(n5761), .Z(n5564) );
  XOR \MIXCOLUMNS[8].d/U357  ( .A(n952), .B(n478), .Z(n5565) );
  XOR \MIXCOLUMNS[8].d/U356  ( .A(n5567), .B(n5566), .Z(\w0[9][20] ) );
  XOR \MIXCOLUMNS[8].d/U355  ( .A(n5770), .B(n5568), .Z(n5566) );
  XOR \MIXCOLUMNS[8].d/U354  ( .A(n475), .B(n5761), .Z(n5567) );
  XOR \MIXCOLUMNS[8].d/U353  ( .A(n950), .B(n476), .Z(n5568) );
  XOR \MIXCOLUMNS[8].d/U352  ( .A(n5570), .B(n5569), .Z(\w0[9][21] ) );
  XOR \MIXCOLUMNS[8].d/U351  ( .A(n473), .B(n5772), .Z(n5569) );
  XOR \MIXCOLUMNS[8].d/U350  ( .A(n948), .B(n474), .Z(n5570) );
  XOR \MIXCOLUMNS[8].d/U349  ( .A(n5572), .B(n5571), .Z(\w0[9][22] ) );
  XOR \MIXCOLUMNS[8].d/U348  ( .A(n5774), .B(n5573), .Z(n5571) );
  XOR \MIXCOLUMNS[8].d/U347  ( .A(n471), .B(n5761), .Z(n5572) );
  XOR \MIXCOLUMNS[8].d/U346  ( .A(n946), .B(n472), .Z(n5573) );
  XOR \MIXCOLUMNS[8].d/U345  ( .A(n5776), .B(n5574), .Z(\w0[9][23] ) );
  XOR \MIXCOLUMNS[8].d/U344  ( .A(n944), .B(n5761), .Z(n5574) );
  XOR \MIXCOLUMNS[8].d/U343  ( .A(n5762), .B(n5575), .Z(\w0[9][24] ) );
  XOR \MIXCOLUMNS[8].d/U342  ( .A(n484), .B(n5763), .Z(n5575) );
  XOR \MIXCOLUMNS[8].d/U341  ( .A(n5764), .B(n5576), .Z(\w0[9][25] ) );
  XOR \MIXCOLUMNS[8].d/U340  ( .A(n483), .B(n5765), .Z(n5576) );
  XOR \MIXCOLUMNS[8].d/U339  ( .A(n5766), .B(n5577), .Z(\w0[9][26] ) );
  XOR \MIXCOLUMNS[8].d/U338  ( .A(\w3[8][18] ), .B(n5767), .Z(n5577) );
  XOR \MIXCOLUMNS[8].d/U337  ( .A(n5579), .B(n5578), .Z(\w0[9][27] ) );
  XOR \MIXCOLUMNS[8].d/U336  ( .A(n5769), .B(n5768), .Z(n5578) );
  XOR \MIXCOLUMNS[8].d/U335  ( .A(n480), .B(n5777), .Z(n5579) );
  XOR \MIXCOLUMNS[8].d/U334  ( .A(n5581), .B(n5580), .Z(\w0[9][28] ) );
  XOR \MIXCOLUMNS[8].d/U333  ( .A(n5771), .B(n5770), .Z(n5580) );
  XOR \MIXCOLUMNS[8].d/U332  ( .A(n478), .B(n5777), .Z(n5581) );
  XOR \MIXCOLUMNS[8].d/U331  ( .A(n5772), .B(n5582), .Z(\w0[9][29] ) );
  XOR \MIXCOLUMNS[8].d/U330  ( .A(n476), .B(n5773), .Z(n5582) );
  XOR \MIXCOLUMNS[8].d/U329  ( .A(n5584), .B(n5583), .Z(\w0[9][30] ) );
  XOR \MIXCOLUMNS[8].d/U328  ( .A(n5775), .B(n5774), .Z(n5583) );
  XOR \MIXCOLUMNS[8].d/U327  ( .A(n474), .B(n5777), .Z(n5584) );
  XOR \MIXCOLUMNS[8].d/U326  ( .A(n5776), .B(n5585), .Z(\w0[9][31] ) );
  XOR \MIXCOLUMNS[8].d/U325  ( .A(n472), .B(n5777), .Z(n5585) );
  XOR \MIXCOLUMNS[8].d/U324  ( .A(n943), .B(n470), .Z(n5795) );
  XOR \MIXCOLUMNS[8].d/U323  ( .A(n5587), .B(n5586), .Z(\w0[9][32] ) );
  XOR \MIXCOLUMNS[8].d/U322  ( .A(n942), .B(n5795), .Z(n5586) );
  XOR \MIXCOLUMNS[8].d/U321  ( .A(n941), .B(n31), .Z(n5587) );
  XOR \MIXCOLUMNS[8].d/U320  ( .A(n941), .B(n469), .Z(n5780) );
  XOR \MIXCOLUMNS[8].d/U319  ( .A(n5589), .B(n5588), .Z(\w0[9][33] ) );
  XOR \MIXCOLUMNS[8].d/U318  ( .A(\w3[8][34] ), .B(n5780), .Z(n5588) );
  XOR \MIXCOLUMNS[8].d/U317  ( .A(\w3[8][58] ), .B(n468), .Z(n5589) );
  XOR \MIXCOLUMNS[8].d/U316  ( .A(\w3[8][58] ), .B(\w3[8][50] ), .Z(n5783) );
  XOR \MIXCOLUMNS[8].d/U315  ( .A(n5591), .B(n5590), .Z(\w0[9][34] ) );
  XOR \MIXCOLUMNS[8].d/U314  ( .A(n940), .B(n5783), .Z(n5590) );
  XOR \MIXCOLUMNS[8].d/U313  ( .A(n939), .B(\w3[8][42] ), .Z(n5591) );
  XOR \MIXCOLUMNS[8].d/U312  ( .A(n943), .B(n467), .Z(n5778) );
  XOR \MIXCOLUMNS[8].d/U311  ( .A(n939), .B(n466), .Z(n5785) );
  XOR \MIXCOLUMNS[8].d/U310  ( .A(n5593), .B(n5592), .Z(\w0[9][35] ) );
  XOR \MIXCOLUMNS[8].d/U309  ( .A(n5785), .B(n5594), .Z(n5592) );
  XOR \MIXCOLUMNS[8].d/U308  ( .A(n938), .B(n5778), .Z(n5593) );
  XOR \MIXCOLUMNS[8].d/U307  ( .A(n937), .B(n465), .Z(n5594) );
  XOR \MIXCOLUMNS[8].d/U306  ( .A(n937), .B(n464), .Z(n5787) );
  XOR \MIXCOLUMNS[8].d/U305  ( .A(n5596), .B(n5595), .Z(\w0[9][36] ) );
  XOR \MIXCOLUMNS[8].d/U304  ( .A(n5787), .B(n5597), .Z(n5595) );
  XOR \MIXCOLUMNS[8].d/U303  ( .A(n936), .B(n5778), .Z(n5596) );
  XOR \MIXCOLUMNS[8].d/U302  ( .A(n935), .B(n463), .Z(n5597) );
  XOR \MIXCOLUMNS[8].d/U301  ( .A(n935), .B(n462), .Z(n5789) );
  XOR \MIXCOLUMNS[8].d/U300  ( .A(n5599), .B(n5598), .Z(\w0[9][37] ) );
  XOR \MIXCOLUMNS[8].d/U299  ( .A(n934), .B(n5789), .Z(n5598) );
  XOR \MIXCOLUMNS[8].d/U298  ( .A(n933), .B(n461), .Z(n5599) );
  XOR \MIXCOLUMNS[8].d/U297  ( .A(n933), .B(n460), .Z(n5791) );
  XOR \MIXCOLUMNS[8].d/U296  ( .A(n5601), .B(n5600), .Z(\w0[9][38] ) );
  XOR \MIXCOLUMNS[8].d/U295  ( .A(n5791), .B(n5602), .Z(n5600) );
  XOR \MIXCOLUMNS[8].d/U294  ( .A(n932), .B(n5778), .Z(n5601) );
  XOR \MIXCOLUMNS[8].d/U293  ( .A(n931), .B(n459), .Z(n5602) );
  XOR \MIXCOLUMNS[8].d/U292  ( .A(n931), .B(n458), .Z(n5793) );
  XOR \MIXCOLUMNS[8].d/U291  ( .A(n5793), .B(n5603), .Z(\w0[9][39] ) );
  XOR \MIXCOLUMNS[8].d/U290  ( .A(n457), .B(n5778), .Z(n5603) );
  XOR \MIXCOLUMNS[8].d/U289  ( .A(n468), .B(n942), .Z(n5782) );
  XOR \MIXCOLUMNS[8].d/U288  ( .A(n5782), .B(n5604), .Z(\w0[9][40] ) );
  XOR \MIXCOLUMNS[8].d/U287  ( .A(n467), .B(n5795), .Z(n5604) );
  XOR \MIXCOLUMNS[8].d/U286  ( .A(\w3[8][42] ), .B(\w3[8][34] ), .Z(n5784) );
  XOR \MIXCOLUMNS[8].d/U285  ( .A(n5784), .B(n5605), .Z(\w0[9][41] ) );
  XOR \MIXCOLUMNS[8].d/U284  ( .A(n942), .B(n5780), .Z(n5605) );
  XOR \MIXCOLUMNS[8].d/U283  ( .A(n465), .B(n940), .Z(n5786) );
  XOR \MIXCOLUMNS[8].d/U282  ( .A(n5786), .B(n5606), .Z(\w0[9][42] ) );
  XOR \MIXCOLUMNS[8].d/U281  ( .A(\w3[8][34] ), .B(n5783), .Z(n5606) );
  XOR \MIXCOLUMNS[8].d/U280  ( .A(n31), .B(n467), .Z(n5781) );
  XOR \MIXCOLUMNS[8].d/U279  ( .A(n463), .B(n938), .Z(n5788) );
  XOR \MIXCOLUMNS[8].d/U278  ( .A(n5608), .B(n5607), .Z(\w0[9][43] ) );
  XOR \MIXCOLUMNS[8].d/U277  ( .A(n5785), .B(n5788), .Z(n5607) );
  XOR \MIXCOLUMNS[8].d/U276  ( .A(n940), .B(n5781), .Z(n5608) );
  XOR \MIXCOLUMNS[8].d/U275  ( .A(n461), .B(n936), .Z(n5790) );
  XOR \MIXCOLUMNS[8].d/U274  ( .A(n5610), .B(n5609), .Z(\w0[9][44] ) );
  XOR \MIXCOLUMNS[8].d/U273  ( .A(n5787), .B(n5790), .Z(n5609) );
  XOR \MIXCOLUMNS[8].d/U272  ( .A(n938), .B(n5781), .Z(n5610) );
  XOR \MIXCOLUMNS[8].d/U271  ( .A(n459), .B(n934), .Z(n5792) );
  XOR \MIXCOLUMNS[8].d/U270  ( .A(n5792), .B(n5611), .Z(\w0[9][45] ) );
  XOR \MIXCOLUMNS[8].d/U269  ( .A(n936), .B(n5789), .Z(n5611) );
  XOR \MIXCOLUMNS[8].d/U268  ( .A(n457), .B(n932), .Z(n5794) );
  XOR \MIXCOLUMNS[8].d/U267  ( .A(n5613), .B(n5612), .Z(\w0[9][46] ) );
  XOR \MIXCOLUMNS[8].d/U266  ( .A(n5791), .B(n5794), .Z(n5612) );
  XOR \MIXCOLUMNS[8].d/U265  ( .A(n934), .B(n5781), .Z(n5613) );
  XOR \MIXCOLUMNS[8].d/U264  ( .A(n5793), .B(n5614), .Z(\w0[9][47] ) );
  XOR \MIXCOLUMNS[8].d/U263  ( .A(n932), .B(n5781), .Z(n5614) );
  XOR \MIXCOLUMNS[8].d/U262  ( .A(n5616), .B(n5615), .Z(\w0[9][48] ) );
  XOR \MIXCOLUMNS[8].d/U261  ( .A(n468), .B(n5781), .Z(n5615) );
  XOR \MIXCOLUMNS[8].d/U260  ( .A(n943), .B(n469), .Z(n5616) );
  XOR \MIXCOLUMNS[8].d/U259  ( .A(n5618), .B(n5617), .Z(\w0[9][49] ) );
  XOR \MIXCOLUMNS[8].d/U258  ( .A(\w3[8][42] ), .B(n5782), .Z(n5617) );
  XOR \MIXCOLUMNS[8].d/U257  ( .A(n941), .B(\w3[8][50] ), .Z(n5618) );
  XOR \MIXCOLUMNS[8].d/U256  ( .A(n5620), .B(n5619), .Z(\w0[9][50] ) );
  XOR \MIXCOLUMNS[8].d/U255  ( .A(n465), .B(n5784), .Z(n5619) );
  XOR \MIXCOLUMNS[8].d/U254  ( .A(\w3[8][58] ), .B(n466), .Z(n5620) );
  XOR \MIXCOLUMNS[8].d/U253  ( .A(n470), .B(n31), .Z(n5779) );
  XOR \MIXCOLUMNS[8].d/U252  ( .A(n5622), .B(n5621), .Z(\w0[9][51] ) );
  XOR \MIXCOLUMNS[8].d/U251  ( .A(n5786), .B(n5623), .Z(n5621) );
  XOR \MIXCOLUMNS[8].d/U250  ( .A(n463), .B(n5779), .Z(n5622) );
  XOR \MIXCOLUMNS[8].d/U249  ( .A(n939), .B(n464), .Z(n5623) );
  XOR \MIXCOLUMNS[8].d/U248  ( .A(n5625), .B(n5624), .Z(\w0[9][52] ) );
  XOR \MIXCOLUMNS[8].d/U247  ( .A(n5788), .B(n5626), .Z(n5624) );
  XOR \MIXCOLUMNS[8].d/U246  ( .A(n461), .B(n5779), .Z(n5625) );
  XOR \MIXCOLUMNS[8].d/U245  ( .A(n937), .B(n462), .Z(n5626) );
  XOR \MIXCOLUMNS[8].d/U244  ( .A(n5628), .B(n5627), .Z(\w0[9][53] ) );
  XOR \MIXCOLUMNS[8].d/U243  ( .A(n459), .B(n5790), .Z(n5627) );
  XOR \MIXCOLUMNS[8].d/U242  ( .A(n935), .B(n460), .Z(n5628) );
  XOR \MIXCOLUMNS[8].d/U241  ( .A(n5630), .B(n5629), .Z(\w0[9][54] ) );
  XOR \MIXCOLUMNS[8].d/U240  ( .A(n5792), .B(n5631), .Z(n5629) );
  XOR \MIXCOLUMNS[8].d/U239  ( .A(n457), .B(n5779), .Z(n5630) );
  XOR \MIXCOLUMNS[8].d/U238  ( .A(n933), .B(n458), .Z(n5631) );
  XOR \MIXCOLUMNS[8].d/U237  ( .A(n5794), .B(n5632), .Z(\w0[9][55] ) );
  XOR \MIXCOLUMNS[8].d/U236  ( .A(n931), .B(n5779), .Z(n5632) );
  XOR \MIXCOLUMNS[8].d/U235  ( .A(n5780), .B(n5633), .Z(\w0[9][56] ) );
  XOR \MIXCOLUMNS[8].d/U234  ( .A(n470), .B(n5781), .Z(n5633) );
  XOR \MIXCOLUMNS[8].d/U233  ( .A(n5782), .B(n5634), .Z(\w0[9][57] ) );
  XOR \MIXCOLUMNS[8].d/U232  ( .A(n469), .B(n5783), .Z(n5634) );
  XOR \MIXCOLUMNS[8].d/U231  ( .A(n5784), .B(n5635), .Z(\w0[9][58] ) );
  XOR \MIXCOLUMNS[8].d/U230  ( .A(\w3[8][50] ), .B(n5785), .Z(n5635) );
  XOR \MIXCOLUMNS[8].d/U229  ( .A(n5637), .B(n5636), .Z(\w0[9][59] ) );
  XOR \MIXCOLUMNS[8].d/U228  ( .A(n5787), .B(n5786), .Z(n5636) );
  XOR \MIXCOLUMNS[8].d/U227  ( .A(n466), .B(n5795), .Z(n5637) );
  XOR \MIXCOLUMNS[8].d/U226  ( .A(n5639), .B(n5638), .Z(\w0[9][60] ) );
  XOR \MIXCOLUMNS[8].d/U225  ( .A(n5789), .B(n5788), .Z(n5638) );
  XOR \MIXCOLUMNS[8].d/U224  ( .A(n464), .B(n5795), .Z(n5639) );
  XOR \MIXCOLUMNS[8].d/U223  ( .A(n5790), .B(n5640), .Z(\w0[9][61] ) );
  XOR \MIXCOLUMNS[8].d/U222  ( .A(n462), .B(n5791), .Z(n5640) );
  XOR \MIXCOLUMNS[8].d/U221  ( .A(n5642), .B(n5641), .Z(\w0[9][62] ) );
  XOR \MIXCOLUMNS[8].d/U220  ( .A(n5793), .B(n5792), .Z(n5641) );
  XOR \MIXCOLUMNS[8].d/U219  ( .A(n460), .B(n5795), .Z(n5642) );
  XOR \MIXCOLUMNS[8].d/U218  ( .A(n5794), .B(n5643), .Z(\w0[9][63] ) );
  XOR \MIXCOLUMNS[8].d/U217  ( .A(n458), .B(n5795), .Z(n5643) );
  XOR \MIXCOLUMNS[8].d/U216  ( .A(n930), .B(n456), .Z(n5813) );
  XOR \MIXCOLUMNS[8].d/U215  ( .A(n5645), .B(n5644), .Z(\w0[9][64] ) );
  XOR \MIXCOLUMNS[8].d/U214  ( .A(n929), .B(n5813), .Z(n5644) );
  XOR \MIXCOLUMNS[8].d/U213  ( .A(n928), .B(n30), .Z(n5645) );
  XOR \MIXCOLUMNS[8].d/U212  ( .A(n928), .B(n455), .Z(n5798) );
  XOR \MIXCOLUMNS[8].d/U211  ( .A(n5647), .B(n5646), .Z(\w0[9][65] ) );
  XOR \MIXCOLUMNS[8].d/U210  ( .A(\w3[8][66] ), .B(n5798), .Z(n5646) );
  XOR \MIXCOLUMNS[8].d/U209  ( .A(\w3[8][90] ), .B(n454), .Z(n5647) );
  XOR \MIXCOLUMNS[8].d/U208  ( .A(\w3[8][90] ), .B(\w3[8][82] ), .Z(n5801) );
  XOR \MIXCOLUMNS[8].d/U207  ( .A(n5649), .B(n5648), .Z(\w0[9][66] ) );
  XOR \MIXCOLUMNS[8].d/U206  ( .A(n927), .B(n5801), .Z(n5648) );
  XOR \MIXCOLUMNS[8].d/U205  ( .A(n926), .B(\w3[8][74] ), .Z(n5649) );
  XOR \MIXCOLUMNS[8].d/U204  ( .A(n930), .B(n453), .Z(n5796) );
  XOR \MIXCOLUMNS[8].d/U203  ( .A(n926), .B(n452), .Z(n5803) );
  XOR \MIXCOLUMNS[8].d/U202  ( .A(n5651), .B(n5650), .Z(\w0[9][67] ) );
  XOR \MIXCOLUMNS[8].d/U201  ( .A(n5803), .B(n5652), .Z(n5650) );
  XOR \MIXCOLUMNS[8].d/U200  ( .A(n925), .B(n5796), .Z(n5651) );
  XOR \MIXCOLUMNS[8].d/U199  ( .A(n924), .B(n451), .Z(n5652) );
  XOR \MIXCOLUMNS[8].d/U198  ( .A(n924), .B(n450), .Z(n5805) );
  XOR \MIXCOLUMNS[8].d/U197  ( .A(n5654), .B(n5653), .Z(\w0[9][68] ) );
  XOR \MIXCOLUMNS[8].d/U196  ( .A(n5805), .B(n5655), .Z(n5653) );
  XOR \MIXCOLUMNS[8].d/U195  ( .A(n923), .B(n5796), .Z(n5654) );
  XOR \MIXCOLUMNS[8].d/U194  ( .A(n922), .B(n449), .Z(n5655) );
  XOR \MIXCOLUMNS[8].d/U193  ( .A(n922), .B(n448), .Z(n5807) );
  XOR \MIXCOLUMNS[8].d/U192  ( .A(n5657), .B(n5656), .Z(\w0[9][69] ) );
  XOR \MIXCOLUMNS[8].d/U191  ( .A(n921), .B(n5807), .Z(n5656) );
  XOR \MIXCOLUMNS[8].d/U190  ( .A(n920), .B(n447), .Z(n5657) );
  XOR \MIXCOLUMNS[8].d/U189  ( .A(n920), .B(n446), .Z(n5809) );
  XOR \MIXCOLUMNS[8].d/U188  ( .A(n5659), .B(n5658), .Z(\w0[9][70] ) );
  XOR \MIXCOLUMNS[8].d/U187  ( .A(n5809), .B(n5660), .Z(n5658) );
  XOR \MIXCOLUMNS[8].d/U186  ( .A(n919), .B(n5796), .Z(n5659) );
  XOR \MIXCOLUMNS[8].d/U185  ( .A(n918), .B(n445), .Z(n5660) );
  XOR \MIXCOLUMNS[8].d/U184  ( .A(n918), .B(n444), .Z(n5811) );
  XOR \MIXCOLUMNS[8].d/U183  ( .A(n5811), .B(n5661), .Z(\w0[9][71] ) );
  XOR \MIXCOLUMNS[8].d/U182  ( .A(n443), .B(n5796), .Z(n5661) );
  XOR \MIXCOLUMNS[8].d/U181  ( .A(n454), .B(n929), .Z(n5800) );
  XOR \MIXCOLUMNS[8].d/U180  ( .A(n5800), .B(n5662), .Z(\w0[9][72] ) );
  XOR \MIXCOLUMNS[8].d/U179  ( .A(n453), .B(n5813), .Z(n5662) );
  XOR \MIXCOLUMNS[8].d/U178  ( .A(\w3[8][74] ), .B(\w3[8][66] ), .Z(n5802) );
  XOR \MIXCOLUMNS[8].d/U177  ( .A(n5802), .B(n5663), .Z(\w0[9][73] ) );
  XOR \MIXCOLUMNS[8].d/U176  ( .A(n929), .B(n5798), .Z(n5663) );
  XOR \MIXCOLUMNS[8].d/U175  ( .A(n451), .B(n927), .Z(n5804) );
  XOR \MIXCOLUMNS[8].d/U174  ( .A(n5804), .B(n5664), .Z(\w0[9][74] ) );
  XOR \MIXCOLUMNS[8].d/U173  ( .A(\w3[8][66] ), .B(n5801), .Z(n5664) );
  XOR \MIXCOLUMNS[8].d/U172  ( .A(n30), .B(n453), .Z(n5799) );
  XOR \MIXCOLUMNS[8].d/U171  ( .A(n449), .B(n925), .Z(n5806) );
  XOR \MIXCOLUMNS[8].d/U170  ( .A(n5666), .B(n5665), .Z(\w0[9][75] ) );
  XOR \MIXCOLUMNS[8].d/U169  ( .A(n5803), .B(n5806), .Z(n5665) );
  XOR \MIXCOLUMNS[8].d/U168  ( .A(n927), .B(n5799), .Z(n5666) );
  XOR \MIXCOLUMNS[8].d/U167  ( .A(n447), .B(n923), .Z(n5808) );
  XOR \MIXCOLUMNS[8].d/U166  ( .A(n5668), .B(n5667), .Z(\w0[9][76] ) );
  XOR \MIXCOLUMNS[8].d/U165  ( .A(n5805), .B(n5808), .Z(n5667) );
  XOR \MIXCOLUMNS[8].d/U164  ( .A(n925), .B(n5799), .Z(n5668) );
  XOR \MIXCOLUMNS[8].d/U163  ( .A(n445), .B(n921), .Z(n5810) );
  XOR \MIXCOLUMNS[8].d/U162  ( .A(n5810), .B(n5669), .Z(\w0[9][77] ) );
  XOR \MIXCOLUMNS[8].d/U161  ( .A(n923), .B(n5807), .Z(n5669) );
  XOR \MIXCOLUMNS[8].d/U160  ( .A(n443), .B(n919), .Z(n5812) );
  XOR \MIXCOLUMNS[8].d/U159  ( .A(n5671), .B(n5670), .Z(\w0[9][78] ) );
  XOR \MIXCOLUMNS[8].d/U158  ( .A(n5809), .B(n5812), .Z(n5670) );
  XOR \MIXCOLUMNS[8].d/U157  ( .A(n921), .B(n5799), .Z(n5671) );
  XOR \MIXCOLUMNS[8].d/U156  ( .A(n5811), .B(n5672), .Z(\w0[9][79] ) );
  XOR \MIXCOLUMNS[8].d/U155  ( .A(n919), .B(n5799), .Z(n5672) );
  XOR \MIXCOLUMNS[8].d/U154  ( .A(n5674), .B(n5673), .Z(\w0[9][80] ) );
  XOR \MIXCOLUMNS[8].d/U153  ( .A(n454), .B(n5799), .Z(n5673) );
  XOR \MIXCOLUMNS[8].d/U152  ( .A(n930), .B(n455), .Z(n5674) );
  XOR \MIXCOLUMNS[8].d/U151  ( .A(n5676), .B(n5675), .Z(\w0[9][81] ) );
  XOR \MIXCOLUMNS[8].d/U150  ( .A(\w3[8][74] ), .B(n5800), .Z(n5675) );
  XOR \MIXCOLUMNS[8].d/U149  ( .A(n928), .B(\w3[8][82] ), .Z(n5676) );
  XOR \MIXCOLUMNS[8].d/U148  ( .A(n5678), .B(n5677), .Z(\w0[9][82] ) );
  XOR \MIXCOLUMNS[8].d/U147  ( .A(n451), .B(n5802), .Z(n5677) );
  XOR \MIXCOLUMNS[8].d/U146  ( .A(\w3[8][90] ), .B(n452), .Z(n5678) );
  XOR \MIXCOLUMNS[8].d/U145  ( .A(n456), .B(n30), .Z(n5797) );
  XOR \MIXCOLUMNS[8].d/U144  ( .A(n5680), .B(n5679), .Z(\w0[9][83] ) );
  XOR \MIXCOLUMNS[8].d/U143  ( .A(n5804), .B(n5681), .Z(n5679) );
  XOR \MIXCOLUMNS[8].d/U142  ( .A(n449), .B(n5797), .Z(n5680) );
  XOR \MIXCOLUMNS[8].d/U141  ( .A(n926), .B(n450), .Z(n5681) );
  XOR \MIXCOLUMNS[8].d/U140  ( .A(n5683), .B(n5682), .Z(\w0[9][84] ) );
  XOR \MIXCOLUMNS[8].d/U139  ( .A(n5806), .B(n5684), .Z(n5682) );
  XOR \MIXCOLUMNS[8].d/U138  ( .A(n447), .B(n5797), .Z(n5683) );
  XOR \MIXCOLUMNS[8].d/U137  ( .A(n924), .B(n448), .Z(n5684) );
  XOR \MIXCOLUMNS[8].d/U136  ( .A(n5686), .B(n5685), .Z(\w0[9][85] ) );
  XOR \MIXCOLUMNS[8].d/U135  ( .A(n445), .B(n5808), .Z(n5685) );
  XOR \MIXCOLUMNS[8].d/U134  ( .A(n922), .B(n446), .Z(n5686) );
  XOR \MIXCOLUMNS[8].d/U133  ( .A(n5688), .B(n5687), .Z(\w0[9][86] ) );
  XOR \MIXCOLUMNS[8].d/U132  ( .A(n5810), .B(n5689), .Z(n5687) );
  XOR \MIXCOLUMNS[8].d/U131  ( .A(n443), .B(n5797), .Z(n5688) );
  XOR \MIXCOLUMNS[8].d/U130  ( .A(n920), .B(n444), .Z(n5689) );
  XOR \MIXCOLUMNS[8].d/U129  ( .A(n5812), .B(n5690), .Z(\w0[9][87] ) );
  XOR \MIXCOLUMNS[8].d/U128  ( .A(n918), .B(n5797), .Z(n5690) );
  XOR \MIXCOLUMNS[8].d/U127  ( .A(n5798), .B(n5691), .Z(\w0[9][88] ) );
  XOR \MIXCOLUMNS[8].d/U126  ( .A(n456), .B(n5799), .Z(n5691) );
  XOR \MIXCOLUMNS[8].d/U125  ( .A(n5800), .B(n5692), .Z(\w0[9][89] ) );
  XOR \MIXCOLUMNS[8].d/U124  ( .A(n455), .B(n5801), .Z(n5692) );
  XOR \MIXCOLUMNS[8].d/U123  ( .A(n5802), .B(n5693), .Z(\w0[9][90] ) );
  XOR \MIXCOLUMNS[8].d/U122  ( .A(\w3[8][82] ), .B(n5803), .Z(n5693) );
  XOR \MIXCOLUMNS[8].d/U121  ( .A(n5695), .B(n5694), .Z(\w0[9][91] ) );
  XOR \MIXCOLUMNS[8].d/U120  ( .A(n5805), .B(n5804), .Z(n5694) );
  XOR \MIXCOLUMNS[8].d/U119  ( .A(n452), .B(n5813), .Z(n5695) );
  XOR \MIXCOLUMNS[8].d/U118  ( .A(n5697), .B(n5696), .Z(\w0[9][92] ) );
  XOR \MIXCOLUMNS[8].d/U117  ( .A(n5807), .B(n5806), .Z(n5696) );
  XOR \MIXCOLUMNS[8].d/U116  ( .A(n450), .B(n5813), .Z(n5697) );
  XOR \MIXCOLUMNS[8].d/U115  ( .A(n5808), .B(n5698), .Z(\w0[9][93] ) );
  XOR \MIXCOLUMNS[8].d/U114  ( .A(n448), .B(n5809), .Z(n5698) );
  XOR \MIXCOLUMNS[8].d/U113  ( .A(n5700), .B(n5699), .Z(\w0[9][94] ) );
  XOR \MIXCOLUMNS[8].d/U112  ( .A(n5811), .B(n5810), .Z(n5699) );
  XOR \MIXCOLUMNS[8].d/U111  ( .A(n446), .B(n5813), .Z(n5700) );
  XOR \MIXCOLUMNS[8].d/U110  ( .A(n5812), .B(n5701), .Z(\w0[9][95] ) );
  XOR \MIXCOLUMNS[8].d/U109  ( .A(n444), .B(n5813), .Z(n5701) );
  XOR \MIXCOLUMNS[8].d/U108  ( .A(n917), .B(n442), .Z(n5831) );
  XOR \MIXCOLUMNS[8].d/U107  ( .A(n5703), .B(n5702), .Z(\w0[9][96] ) );
  XOR \MIXCOLUMNS[8].d/U106  ( .A(n916), .B(n5831), .Z(n5702) );
  XOR \MIXCOLUMNS[8].d/U105  ( .A(n915), .B(n29), .Z(n5703) );
  XOR \MIXCOLUMNS[8].d/U104  ( .A(n915), .B(n441), .Z(n5816) );
  XOR \MIXCOLUMNS[8].d/U103  ( .A(n5705), .B(n5704), .Z(\w0[9][97] ) );
  XOR \MIXCOLUMNS[8].d/U102  ( .A(\w3[8][98] ), .B(n5816), .Z(n5704) );
  XOR \MIXCOLUMNS[8].d/U101  ( .A(\w3[8][122] ), .B(n440), .Z(n5705) );
  XOR \MIXCOLUMNS[8].d/U100  ( .A(\w3[8][122] ), .B(\w3[8][114] ), .Z(n5819)
         );
  XOR \MIXCOLUMNS[8].d/U99  ( .A(n5707), .B(n5706), .Z(\w0[9][98] ) );
  XOR \MIXCOLUMNS[8].d/U98  ( .A(n914), .B(n5819), .Z(n5706) );
  XOR \MIXCOLUMNS[8].d/U97  ( .A(n913), .B(\w3[8][106] ), .Z(n5707) );
  XOR \MIXCOLUMNS[8].d/U96  ( .A(n917), .B(n439), .Z(n5814) );
  XOR \MIXCOLUMNS[8].d/U95  ( .A(n913), .B(n438), .Z(n5821) );
  XOR \MIXCOLUMNS[8].d/U94  ( .A(n5709), .B(n5708), .Z(\w0[9][99] ) );
  XOR \MIXCOLUMNS[8].d/U93  ( .A(n5821), .B(n5710), .Z(n5708) );
  XOR \MIXCOLUMNS[8].d/U92  ( .A(n912), .B(n5814), .Z(n5709) );
  XOR \MIXCOLUMNS[8].d/U91  ( .A(n911), .B(n437), .Z(n5710) );
  XOR \MIXCOLUMNS[8].d/U90  ( .A(n911), .B(n436), .Z(n5823) );
  XOR \MIXCOLUMNS[8].d/U89  ( .A(n5712), .B(n5711), .Z(\w0[9][100] ) );
  XOR \MIXCOLUMNS[8].d/U88  ( .A(n5823), .B(n5713), .Z(n5711) );
  XOR \MIXCOLUMNS[8].d/U87  ( .A(n910), .B(n5814), .Z(n5712) );
  XOR \MIXCOLUMNS[8].d/U86  ( .A(n909), .B(n435), .Z(n5713) );
  XOR \MIXCOLUMNS[8].d/U85  ( .A(n909), .B(n434), .Z(n5825) );
  XOR \MIXCOLUMNS[8].d/U84  ( .A(n5715), .B(n5714), .Z(\w0[9][101] ) );
  XOR \MIXCOLUMNS[8].d/U83  ( .A(n908), .B(n5825), .Z(n5714) );
  XOR \MIXCOLUMNS[8].d/U82  ( .A(n907), .B(n433), .Z(n5715) );
  XOR \MIXCOLUMNS[8].d/U81  ( .A(n907), .B(n432), .Z(n5827) );
  XOR \MIXCOLUMNS[8].d/U80  ( .A(n5717), .B(n5716), .Z(\w0[9][102] ) );
  XOR \MIXCOLUMNS[8].d/U79  ( .A(n5827), .B(n5718), .Z(n5716) );
  XOR \MIXCOLUMNS[8].d/U78  ( .A(n906), .B(n5814), .Z(n5717) );
  XOR \MIXCOLUMNS[8].d/U77  ( .A(n905), .B(n431), .Z(n5718) );
  XOR \MIXCOLUMNS[8].d/U76  ( .A(n905), .B(n430), .Z(n5829) );
  XOR \MIXCOLUMNS[8].d/U75  ( .A(n5829), .B(n5719), .Z(\w0[9][103] ) );
  XOR \MIXCOLUMNS[8].d/U74  ( .A(n429), .B(n5814), .Z(n5719) );
  XOR \MIXCOLUMNS[8].d/U73  ( .A(n440), .B(n916), .Z(n5818) );
  XOR \MIXCOLUMNS[8].d/U72  ( .A(n5818), .B(n5720), .Z(\w0[9][104] ) );
  XOR \MIXCOLUMNS[8].d/U71  ( .A(n439), .B(n5831), .Z(n5720) );
  XOR \MIXCOLUMNS[8].d/U70  ( .A(\w3[8][106] ), .B(\w3[8][98] ), .Z(n5820) );
  XOR \MIXCOLUMNS[8].d/U69  ( .A(n5820), .B(n5721), .Z(\w0[9][105] ) );
  XOR \MIXCOLUMNS[8].d/U68  ( .A(n916), .B(n5816), .Z(n5721) );
  XOR \MIXCOLUMNS[8].d/U67  ( .A(n437), .B(n914), .Z(n5822) );
  XOR \MIXCOLUMNS[8].d/U66  ( .A(n5822), .B(n5722), .Z(\w0[9][106] ) );
  XOR \MIXCOLUMNS[8].d/U65  ( .A(\w3[8][98] ), .B(n5819), .Z(n5722) );
  XOR \MIXCOLUMNS[8].d/U64  ( .A(n29), .B(n439), .Z(n5817) );
  XOR \MIXCOLUMNS[8].d/U63  ( .A(n435), .B(n912), .Z(n5824) );
  XOR \MIXCOLUMNS[8].d/U62  ( .A(n5724), .B(n5723), .Z(\w0[9][107] ) );
  XOR \MIXCOLUMNS[8].d/U61  ( .A(n5821), .B(n5824), .Z(n5723) );
  XOR \MIXCOLUMNS[8].d/U60  ( .A(n914), .B(n5817), .Z(n5724) );
  XOR \MIXCOLUMNS[8].d/U59  ( .A(n433), .B(n910), .Z(n5826) );
  XOR \MIXCOLUMNS[8].d/U58  ( .A(n5726), .B(n5725), .Z(\w0[9][108] ) );
  XOR \MIXCOLUMNS[8].d/U57  ( .A(n5823), .B(n5826), .Z(n5725) );
  XOR \MIXCOLUMNS[8].d/U56  ( .A(n912), .B(n5817), .Z(n5726) );
  XOR \MIXCOLUMNS[8].d/U55  ( .A(n431), .B(n908), .Z(n5828) );
  XOR \MIXCOLUMNS[8].d/U54  ( .A(n5828), .B(n5727), .Z(\w0[9][109] ) );
  XOR \MIXCOLUMNS[8].d/U53  ( .A(n910), .B(n5825), .Z(n5727) );
  XOR \MIXCOLUMNS[8].d/U52  ( .A(n429), .B(n906), .Z(n5830) );
  XOR \MIXCOLUMNS[8].d/U51  ( .A(n5729), .B(n5728), .Z(\w0[9][110] ) );
  XOR \MIXCOLUMNS[8].d/U50  ( .A(n5827), .B(n5830), .Z(n5728) );
  XOR \MIXCOLUMNS[8].d/U49  ( .A(n908), .B(n5817), .Z(n5729) );
  XOR \MIXCOLUMNS[8].d/U48  ( .A(n5829), .B(n5730), .Z(\w0[9][111] ) );
  XOR \MIXCOLUMNS[8].d/U47  ( .A(n906), .B(n5817), .Z(n5730) );
  XOR \MIXCOLUMNS[8].d/U46  ( .A(n5732), .B(n5731), .Z(\w0[9][112] ) );
  XOR \MIXCOLUMNS[8].d/U45  ( .A(n440), .B(n5817), .Z(n5731) );
  XOR \MIXCOLUMNS[8].d/U44  ( .A(n917), .B(n441), .Z(n5732) );
  XOR \MIXCOLUMNS[8].d/U43  ( .A(n5734), .B(n5733), .Z(\w0[9][113] ) );
  XOR \MIXCOLUMNS[8].d/U42  ( .A(\w3[8][106] ), .B(n5818), .Z(n5733) );
  XOR \MIXCOLUMNS[8].d/U41  ( .A(n915), .B(\w3[8][114] ), .Z(n5734) );
  XOR \MIXCOLUMNS[8].d/U40  ( .A(n5736), .B(n5735), .Z(\w0[9][114] ) );
  XOR \MIXCOLUMNS[8].d/U39  ( .A(n437), .B(n5820), .Z(n5735) );
  XOR \MIXCOLUMNS[8].d/U38  ( .A(\w3[8][122] ), .B(n438), .Z(n5736) );
  XOR \MIXCOLUMNS[8].d/U37  ( .A(n442), .B(n29), .Z(n5815) );
  XOR \MIXCOLUMNS[8].d/U36  ( .A(n5738), .B(n5737), .Z(\w0[9][115] ) );
  XOR \MIXCOLUMNS[8].d/U35  ( .A(n5822), .B(n5739), .Z(n5737) );
  XOR \MIXCOLUMNS[8].d/U34  ( .A(n435), .B(n5815), .Z(n5738) );
  XOR \MIXCOLUMNS[8].d/U33  ( .A(n913), .B(n436), .Z(n5739) );
  XOR \MIXCOLUMNS[8].d/U32  ( .A(n5741), .B(n5740), .Z(\w0[9][116] ) );
  XOR \MIXCOLUMNS[8].d/U31  ( .A(n5824), .B(n5742), .Z(n5740) );
  XOR \MIXCOLUMNS[8].d/U30  ( .A(n433), .B(n5815), .Z(n5741) );
  XOR \MIXCOLUMNS[8].d/U29  ( .A(n911), .B(n434), .Z(n5742) );
  XOR \MIXCOLUMNS[8].d/U28  ( .A(n5744), .B(n5743), .Z(\w0[9][117] ) );
  XOR \MIXCOLUMNS[8].d/U27  ( .A(n431), .B(n5826), .Z(n5743) );
  XOR \MIXCOLUMNS[8].d/U26  ( .A(n909), .B(n432), .Z(n5744) );
  XOR \MIXCOLUMNS[8].d/U25  ( .A(n5746), .B(n5745), .Z(\w0[9][118] ) );
  XOR \MIXCOLUMNS[8].d/U24  ( .A(n5828), .B(n5747), .Z(n5745) );
  XOR \MIXCOLUMNS[8].d/U23  ( .A(n429), .B(n5815), .Z(n5746) );
  XOR \MIXCOLUMNS[8].d/U22  ( .A(n907), .B(n430), .Z(n5747) );
  XOR \MIXCOLUMNS[8].d/U21  ( .A(n5830), .B(n5748), .Z(\w0[9][119] ) );
  XOR \MIXCOLUMNS[8].d/U20  ( .A(n905), .B(n5815), .Z(n5748) );
  XOR \MIXCOLUMNS[8].d/U19  ( .A(n5816), .B(n5749), .Z(\w0[9][120] ) );
  XOR \MIXCOLUMNS[8].d/U18  ( .A(n442), .B(n5817), .Z(n5749) );
  XOR \MIXCOLUMNS[8].d/U17  ( .A(n5818), .B(n5750), .Z(\w0[9][121] ) );
  XOR \MIXCOLUMNS[8].d/U16  ( .A(n441), .B(n5819), .Z(n5750) );
  XOR \MIXCOLUMNS[8].d/U15  ( .A(n5820), .B(n5751), .Z(\w0[9][122] ) );
  XOR \MIXCOLUMNS[8].d/U14  ( .A(\w3[8][114] ), .B(n5821), .Z(n5751) );
  XOR \MIXCOLUMNS[8].d/U13  ( .A(n5753), .B(n5752), .Z(\w0[9][123] ) );
  XOR \MIXCOLUMNS[8].d/U12  ( .A(n5823), .B(n5822), .Z(n5752) );
  XOR \MIXCOLUMNS[8].d/U11  ( .A(n438), .B(n5831), .Z(n5753) );
  XOR \MIXCOLUMNS[8].d/U10  ( .A(n5755), .B(n5754), .Z(\w0[9][124] ) );
  XOR \MIXCOLUMNS[8].d/U9  ( .A(n5825), .B(n5824), .Z(n5754) );
  XOR \MIXCOLUMNS[8].d/U8  ( .A(n436), .B(n5831), .Z(n5755) );
  XOR \MIXCOLUMNS[8].d/U7  ( .A(n5826), .B(n5756), .Z(\w0[9][125] ) );
  XOR \MIXCOLUMNS[8].d/U6  ( .A(n434), .B(n5827), .Z(n5756) );
  XOR \MIXCOLUMNS[8].d/U5  ( .A(n5758), .B(n5757), .Z(\w0[9][126] ) );
  XOR \MIXCOLUMNS[8].d/U4  ( .A(n5829), .B(n5828), .Z(n5757) );
  XOR \MIXCOLUMNS[8].d/U3  ( .A(n432), .B(n5831), .Z(n5758) );
  XOR \MIXCOLUMNS[8].d/U2  ( .A(n5830), .B(n5759), .Z(\w0[9][127] ) );
  XOR \MIXCOLUMNS[8].d/U1  ( .A(n430), .B(n5831), .Z(n5759) );
  XOR \MIXCOLUMNS[7].d/U432  ( .A(n904), .B(n428), .Z(n5473) );
  XOR \MIXCOLUMNS[7].d/U431  ( .A(n5225), .B(n5224), .Z(\w0[8][0] ) );
  XOR \MIXCOLUMNS[7].d/U430  ( .A(n903), .B(n5473), .Z(n5224) );
  XOR \MIXCOLUMNS[7].d/U429  ( .A(n902), .B(n28), .Z(n5225) );
  XOR \MIXCOLUMNS[7].d/U428  ( .A(n902), .B(n427), .Z(n5458) );
  XOR \MIXCOLUMNS[7].d/U427  ( .A(n5227), .B(n5226), .Z(\w0[8][1] ) );
  XOR \MIXCOLUMNS[7].d/U426  ( .A(\w3[7][2] ), .B(n5458), .Z(n5226) );
  XOR \MIXCOLUMNS[7].d/U425  ( .A(\w3[7][26] ), .B(n426), .Z(n5227) );
  XOR \MIXCOLUMNS[7].d/U424  ( .A(\w3[7][26] ), .B(\w3[7][18] ), .Z(n5461) );
  XOR \MIXCOLUMNS[7].d/U423  ( .A(n5229), .B(n5228), .Z(\w0[8][2] ) );
  XOR \MIXCOLUMNS[7].d/U422  ( .A(n901), .B(n5461), .Z(n5228) );
  XOR \MIXCOLUMNS[7].d/U421  ( .A(n900), .B(\w3[7][10] ), .Z(n5229) );
  XOR \MIXCOLUMNS[7].d/U420  ( .A(n904), .B(n425), .Z(n5456) );
  XOR \MIXCOLUMNS[7].d/U419  ( .A(n900), .B(n424), .Z(n5463) );
  XOR \MIXCOLUMNS[7].d/U418  ( .A(n5231), .B(n5230), .Z(\w0[8][3] ) );
  XOR \MIXCOLUMNS[7].d/U417  ( .A(n5463), .B(n5232), .Z(n5230) );
  XOR \MIXCOLUMNS[7].d/U416  ( .A(n899), .B(n5456), .Z(n5231) );
  XOR \MIXCOLUMNS[7].d/U415  ( .A(n898), .B(n423), .Z(n5232) );
  XOR \MIXCOLUMNS[7].d/U414  ( .A(n898), .B(n422), .Z(n5465) );
  XOR \MIXCOLUMNS[7].d/U413  ( .A(n5234), .B(n5233), .Z(\w0[8][4] ) );
  XOR \MIXCOLUMNS[7].d/U412  ( .A(n5465), .B(n5235), .Z(n5233) );
  XOR \MIXCOLUMNS[7].d/U411  ( .A(n897), .B(n5456), .Z(n5234) );
  XOR \MIXCOLUMNS[7].d/U410  ( .A(n896), .B(n421), .Z(n5235) );
  XOR \MIXCOLUMNS[7].d/U409  ( .A(n896), .B(n420), .Z(n5467) );
  XOR \MIXCOLUMNS[7].d/U408  ( .A(n5237), .B(n5236), .Z(\w0[8][5] ) );
  XOR \MIXCOLUMNS[7].d/U407  ( .A(n895), .B(n5467), .Z(n5236) );
  XOR \MIXCOLUMNS[7].d/U406  ( .A(n894), .B(n419), .Z(n5237) );
  XOR \MIXCOLUMNS[7].d/U405  ( .A(n894), .B(n418), .Z(n5469) );
  XOR \MIXCOLUMNS[7].d/U404  ( .A(n5239), .B(n5238), .Z(\w0[8][6] ) );
  XOR \MIXCOLUMNS[7].d/U403  ( .A(n5469), .B(n5240), .Z(n5238) );
  XOR \MIXCOLUMNS[7].d/U402  ( .A(n893), .B(n5456), .Z(n5239) );
  XOR \MIXCOLUMNS[7].d/U401  ( .A(n892), .B(n417), .Z(n5240) );
  XOR \MIXCOLUMNS[7].d/U400  ( .A(n892), .B(n416), .Z(n5471) );
  XOR \MIXCOLUMNS[7].d/U399  ( .A(n5471), .B(n5241), .Z(\w0[8][7] ) );
  XOR \MIXCOLUMNS[7].d/U398  ( .A(n415), .B(n5456), .Z(n5241) );
  XOR \MIXCOLUMNS[7].d/U397  ( .A(n426), .B(n903), .Z(n5460) );
  XOR \MIXCOLUMNS[7].d/U396  ( .A(n5460), .B(n5242), .Z(\w0[8][8] ) );
  XOR \MIXCOLUMNS[7].d/U395  ( .A(n425), .B(n5473), .Z(n5242) );
  XOR \MIXCOLUMNS[7].d/U394  ( .A(\w3[7][10] ), .B(\w3[7][2] ), .Z(n5462) );
  XOR \MIXCOLUMNS[7].d/U393  ( .A(n5462), .B(n5243), .Z(\w0[8][9] ) );
  XOR \MIXCOLUMNS[7].d/U392  ( .A(n903), .B(n5458), .Z(n5243) );
  XOR \MIXCOLUMNS[7].d/U391  ( .A(n423), .B(n901), .Z(n5464) );
  XOR \MIXCOLUMNS[7].d/U390  ( .A(n5464), .B(n5244), .Z(\w0[8][10] ) );
  XOR \MIXCOLUMNS[7].d/U389  ( .A(\w3[7][2] ), .B(n5461), .Z(n5244) );
  XOR \MIXCOLUMNS[7].d/U388  ( .A(n28), .B(n425), .Z(n5459) );
  XOR \MIXCOLUMNS[7].d/U387  ( .A(n421), .B(n899), .Z(n5466) );
  XOR \MIXCOLUMNS[7].d/U386  ( .A(n5246), .B(n5245), .Z(\w0[8][11] ) );
  XOR \MIXCOLUMNS[7].d/U385  ( .A(n5463), .B(n5466), .Z(n5245) );
  XOR \MIXCOLUMNS[7].d/U384  ( .A(n901), .B(n5459), .Z(n5246) );
  XOR \MIXCOLUMNS[7].d/U383  ( .A(n419), .B(n897), .Z(n5468) );
  XOR \MIXCOLUMNS[7].d/U382  ( .A(n5248), .B(n5247), .Z(\w0[8][12] ) );
  XOR \MIXCOLUMNS[7].d/U381  ( .A(n5465), .B(n5468), .Z(n5247) );
  XOR \MIXCOLUMNS[7].d/U380  ( .A(n899), .B(n5459), .Z(n5248) );
  XOR \MIXCOLUMNS[7].d/U379  ( .A(n417), .B(n895), .Z(n5470) );
  XOR \MIXCOLUMNS[7].d/U378  ( .A(n5470), .B(n5249), .Z(\w0[8][13] ) );
  XOR \MIXCOLUMNS[7].d/U377  ( .A(n897), .B(n5467), .Z(n5249) );
  XOR \MIXCOLUMNS[7].d/U376  ( .A(n415), .B(n893), .Z(n5472) );
  XOR \MIXCOLUMNS[7].d/U375  ( .A(n5251), .B(n5250), .Z(\w0[8][14] ) );
  XOR \MIXCOLUMNS[7].d/U374  ( .A(n5469), .B(n5472), .Z(n5250) );
  XOR \MIXCOLUMNS[7].d/U373  ( .A(n895), .B(n5459), .Z(n5251) );
  XOR \MIXCOLUMNS[7].d/U372  ( .A(n5471), .B(n5252), .Z(\w0[8][15] ) );
  XOR \MIXCOLUMNS[7].d/U371  ( .A(n893), .B(n5459), .Z(n5252) );
  XOR \MIXCOLUMNS[7].d/U370  ( .A(n5254), .B(n5253), .Z(\w0[8][16] ) );
  XOR \MIXCOLUMNS[7].d/U369  ( .A(n426), .B(n5459), .Z(n5253) );
  XOR \MIXCOLUMNS[7].d/U368  ( .A(n904), .B(n427), .Z(n5254) );
  XOR \MIXCOLUMNS[7].d/U367  ( .A(n5256), .B(n5255), .Z(\w0[8][17] ) );
  XOR \MIXCOLUMNS[7].d/U366  ( .A(\w3[7][10] ), .B(n5460), .Z(n5255) );
  XOR \MIXCOLUMNS[7].d/U365  ( .A(n902), .B(\w3[7][18] ), .Z(n5256) );
  XOR \MIXCOLUMNS[7].d/U364  ( .A(n5258), .B(n5257), .Z(\w0[8][18] ) );
  XOR \MIXCOLUMNS[7].d/U363  ( .A(n423), .B(n5462), .Z(n5257) );
  XOR \MIXCOLUMNS[7].d/U362  ( .A(\w3[7][26] ), .B(n424), .Z(n5258) );
  XOR \MIXCOLUMNS[7].d/U361  ( .A(n428), .B(n28), .Z(n5457) );
  XOR \MIXCOLUMNS[7].d/U360  ( .A(n5260), .B(n5259), .Z(\w0[8][19] ) );
  XOR \MIXCOLUMNS[7].d/U359  ( .A(n5464), .B(n5261), .Z(n5259) );
  XOR \MIXCOLUMNS[7].d/U358  ( .A(n421), .B(n5457), .Z(n5260) );
  XOR \MIXCOLUMNS[7].d/U357  ( .A(n900), .B(n422), .Z(n5261) );
  XOR \MIXCOLUMNS[7].d/U356  ( .A(n5263), .B(n5262), .Z(\w0[8][20] ) );
  XOR \MIXCOLUMNS[7].d/U355  ( .A(n5466), .B(n5264), .Z(n5262) );
  XOR \MIXCOLUMNS[7].d/U354  ( .A(n419), .B(n5457), .Z(n5263) );
  XOR \MIXCOLUMNS[7].d/U353  ( .A(n898), .B(n420), .Z(n5264) );
  XOR \MIXCOLUMNS[7].d/U352  ( .A(n5266), .B(n5265), .Z(\w0[8][21] ) );
  XOR \MIXCOLUMNS[7].d/U351  ( .A(n417), .B(n5468), .Z(n5265) );
  XOR \MIXCOLUMNS[7].d/U350  ( .A(n896), .B(n418), .Z(n5266) );
  XOR \MIXCOLUMNS[7].d/U349  ( .A(n5268), .B(n5267), .Z(\w0[8][22] ) );
  XOR \MIXCOLUMNS[7].d/U348  ( .A(n5470), .B(n5269), .Z(n5267) );
  XOR \MIXCOLUMNS[7].d/U347  ( .A(n415), .B(n5457), .Z(n5268) );
  XOR \MIXCOLUMNS[7].d/U346  ( .A(n894), .B(n416), .Z(n5269) );
  XOR \MIXCOLUMNS[7].d/U345  ( .A(n5472), .B(n5270), .Z(\w0[8][23] ) );
  XOR \MIXCOLUMNS[7].d/U344  ( .A(n892), .B(n5457), .Z(n5270) );
  XOR \MIXCOLUMNS[7].d/U343  ( .A(n5458), .B(n5271), .Z(\w0[8][24] ) );
  XOR \MIXCOLUMNS[7].d/U342  ( .A(n428), .B(n5459), .Z(n5271) );
  XOR \MIXCOLUMNS[7].d/U341  ( .A(n5460), .B(n5272), .Z(\w0[8][25] ) );
  XOR \MIXCOLUMNS[7].d/U340  ( .A(n427), .B(n5461), .Z(n5272) );
  XOR \MIXCOLUMNS[7].d/U339  ( .A(n5462), .B(n5273), .Z(\w0[8][26] ) );
  XOR \MIXCOLUMNS[7].d/U338  ( .A(\w3[7][18] ), .B(n5463), .Z(n5273) );
  XOR \MIXCOLUMNS[7].d/U337  ( .A(n5275), .B(n5274), .Z(\w0[8][27] ) );
  XOR \MIXCOLUMNS[7].d/U336  ( .A(n5465), .B(n5464), .Z(n5274) );
  XOR \MIXCOLUMNS[7].d/U335  ( .A(n424), .B(n5473), .Z(n5275) );
  XOR \MIXCOLUMNS[7].d/U334  ( .A(n5277), .B(n5276), .Z(\w0[8][28] ) );
  XOR \MIXCOLUMNS[7].d/U333  ( .A(n5467), .B(n5466), .Z(n5276) );
  XOR \MIXCOLUMNS[7].d/U332  ( .A(n422), .B(n5473), .Z(n5277) );
  XOR \MIXCOLUMNS[7].d/U331  ( .A(n5468), .B(n5278), .Z(\w0[8][29] ) );
  XOR \MIXCOLUMNS[7].d/U330  ( .A(n420), .B(n5469), .Z(n5278) );
  XOR \MIXCOLUMNS[7].d/U329  ( .A(n5280), .B(n5279), .Z(\w0[8][30] ) );
  XOR \MIXCOLUMNS[7].d/U328  ( .A(n5471), .B(n5470), .Z(n5279) );
  XOR \MIXCOLUMNS[7].d/U327  ( .A(n418), .B(n5473), .Z(n5280) );
  XOR \MIXCOLUMNS[7].d/U326  ( .A(n5472), .B(n5281), .Z(\w0[8][31] ) );
  XOR \MIXCOLUMNS[7].d/U325  ( .A(n416), .B(n5473), .Z(n5281) );
  XOR \MIXCOLUMNS[7].d/U324  ( .A(n891), .B(n414), .Z(n5491) );
  XOR \MIXCOLUMNS[7].d/U323  ( .A(n5283), .B(n5282), .Z(\w0[8][32] ) );
  XOR \MIXCOLUMNS[7].d/U322  ( .A(n890), .B(n5491), .Z(n5282) );
  XOR \MIXCOLUMNS[7].d/U321  ( .A(n889), .B(n27), .Z(n5283) );
  XOR \MIXCOLUMNS[7].d/U320  ( .A(n889), .B(n413), .Z(n5476) );
  XOR \MIXCOLUMNS[7].d/U319  ( .A(n5285), .B(n5284), .Z(\w0[8][33] ) );
  XOR \MIXCOLUMNS[7].d/U318  ( .A(\w3[7][34] ), .B(n5476), .Z(n5284) );
  XOR \MIXCOLUMNS[7].d/U317  ( .A(\w3[7][58] ), .B(n412), .Z(n5285) );
  XOR \MIXCOLUMNS[7].d/U316  ( .A(\w3[7][58] ), .B(\w3[7][50] ), .Z(n5479) );
  XOR \MIXCOLUMNS[7].d/U315  ( .A(n5287), .B(n5286), .Z(\w0[8][34] ) );
  XOR \MIXCOLUMNS[7].d/U314  ( .A(n888), .B(n5479), .Z(n5286) );
  XOR \MIXCOLUMNS[7].d/U313  ( .A(n887), .B(\w3[7][42] ), .Z(n5287) );
  XOR \MIXCOLUMNS[7].d/U312  ( .A(n891), .B(n411), .Z(n5474) );
  XOR \MIXCOLUMNS[7].d/U311  ( .A(n887), .B(n410), .Z(n5481) );
  XOR \MIXCOLUMNS[7].d/U310  ( .A(n5289), .B(n5288), .Z(\w0[8][35] ) );
  XOR \MIXCOLUMNS[7].d/U309  ( .A(n5481), .B(n5290), .Z(n5288) );
  XOR \MIXCOLUMNS[7].d/U308  ( .A(n886), .B(n5474), .Z(n5289) );
  XOR \MIXCOLUMNS[7].d/U307  ( .A(n885), .B(n409), .Z(n5290) );
  XOR \MIXCOLUMNS[7].d/U306  ( .A(n885), .B(n408), .Z(n5483) );
  XOR \MIXCOLUMNS[7].d/U305  ( .A(n5292), .B(n5291), .Z(\w0[8][36] ) );
  XOR \MIXCOLUMNS[7].d/U304  ( .A(n5483), .B(n5293), .Z(n5291) );
  XOR \MIXCOLUMNS[7].d/U303  ( .A(n884), .B(n5474), .Z(n5292) );
  XOR \MIXCOLUMNS[7].d/U302  ( .A(n883), .B(n407), .Z(n5293) );
  XOR \MIXCOLUMNS[7].d/U301  ( .A(n883), .B(n406), .Z(n5485) );
  XOR \MIXCOLUMNS[7].d/U300  ( .A(n5295), .B(n5294), .Z(\w0[8][37] ) );
  XOR \MIXCOLUMNS[7].d/U299  ( .A(n882), .B(n5485), .Z(n5294) );
  XOR \MIXCOLUMNS[7].d/U298  ( .A(n881), .B(n405), .Z(n5295) );
  XOR \MIXCOLUMNS[7].d/U297  ( .A(n881), .B(n404), .Z(n5487) );
  XOR \MIXCOLUMNS[7].d/U296  ( .A(n5297), .B(n5296), .Z(\w0[8][38] ) );
  XOR \MIXCOLUMNS[7].d/U295  ( .A(n5487), .B(n5298), .Z(n5296) );
  XOR \MIXCOLUMNS[7].d/U294  ( .A(n880), .B(n5474), .Z(n5297) );
  XOR \MIXCOLUMNS[7].d/U293  ( .A(n879), .B(n403), .Z(n5298) );
  XOR \MIXCOLUMNS[7].d/U292  ( .A(n879), .B(n402), .Z(n5489) );
  XOR \MIXCOLUMNS[7].d/U291  ( .A(n5489), .B(n5299), .Z(\w0[8][39] ) );
  XOR \MIXCOLUMNS[7].d/U290  ( .A(n401), .B(n5474), .Z(n5299) );
  XOR \MIXCOLUMNS[7].d/U289  ( .A(n412), .B(n890), .Z(n5478) );
  XOR \MIXCOLUMNS[7].d/U288  ( .A(n5478), .B(n5300), .Z(\w0[8][40] ) );
  XOR \MIXCOLUMNS[7].d/U287  ( .A(n411), .B(n5491), .Z(n5300) );
  XOR \MIXCOLUMNS[7].d/U286  ( .A(\w3[7][42] ), .B(\w3[7][34] ), .Z(n5480) );
  XOR \MIXCOLUMNS[7].d/U285  ( .A(n5480), .B(n5301), .Z(\w0[8][41] ) );
  XOR \MIXCOLUMNS[7].d/U284  ( .A(n890), .B(n5476), .Z(n5301) );
  XOR \MIXCOLUMNS[7].d/U283  ( .A(n409), .B(n888), .Z(n5482) );
  XOR \MIXCOLUMNS[7].d/U282  ( .A(n5482), .B(n5302), .Z(\w0[8][42] ) );
  XOR \MIXCOLUMNS[7].d/U281  ( .A(\w3[7][34] ), .B(n5479), .Z(n5302) );
  XOR \MIXCOLUMNS[7].d/U280  ( .A(n27), .B(n411), .Z(n5477) );
  XOR \MIXCOLUMNS[7].d/U279  ( .A(n407), .B(n886), .Z(n5484) );
  XOR \MIXCOLUMNS[7].d/U278  ( .A(n5304), .B(n5303), .Z(\w0[8][43] ) );
  XOR \MIXCOLUMNS[7].d/U277  ( .A(n5481), .B(n5484), .Z(n5303) );
  XOR \MIXCOLUMNS[7].d/U276  ( .A(n888), .B(n5477), .Z(n5304) );
  XOR \MIXCOLUMNS[7].d/U275  ( .A(n405), .B(n884), .Z(n5486) );
  XOR \MIXCOLUMNS[7].d/U274  ( .A(n5306), .B(n5305), .Z(\w0[8][44] ) );
  XOR \MIXCOLUMNS[7].d/U273  ( .A(n5483), .B(n5486), .Z(n5305) );
  XOR \MIXCOLUMNS[7].d/U272  ( .A(n886), .B(n5477), .Z(n5306) );
  XOR \MIXCOLUMNS[7].d/U271  ( .A(n403), .B(n882), .Z(n5488) );
  XOR \MIXCOLUMNS[7].d/U270  ( .A(n5488), .B(n5307), .Z(\w0[8][45] ) );
  XOR \MIXCOLUMNS[7].d/U269  ( .A(n884), .B(n5485), .Z(n5307) );
  XOR \MIXCOLUMNS[7].d/U268  ( .A(n401), .B(n880), .Z(n5490) );
  XOR \MIXCOLUMNS[7].d/U267  ( .A(n5309), .B(n5308), .Z(\w0[8][46] ) );
  XOR \MIXCOLUMNS[7].d/U266  ( .A(n5487), .B(n5490), .Z(n5308) );
  XOR \MIXCOLUMNS[7].d/U265  ( .A(n882), .B(n5477), .Z(n5309) );
  XOR \MIXCOLUMNS[7].d/U264  ( .A(n5489), .B(n5310), .Z(\w0[8][47] ) );
  XOR \MIXCOLUMNS[7].d/U263  ( .A(n880), .B(n5477), .Z(n5310) );
  XOR \MIXCOLUMNS[7].d/U262  ( .A(n5312), .B(n5311), .Z(\w0[8][48] ) );
  XOR \MIXCOLUMNS[7].d/U261  ( .A(n412), .B(n5477), .Z(n5311) );
  XOR \MIXCOLUMNS[7].d/U260  ( .A(n891), .B(n413), .Z(n5312) );
  XOR \MIXCOLUMNS[7].d/U259  ( .A(n5314), .B(n5313), .Z(\w0[8][49] ) );
  XOR \MIXCOLUMNS[7].d/U258  ( .A(\w3[7][42] ), .B(n5478), .Z(n5313) );
  XOR \MIXCOLUMNS[7].d/U257  ( .A(n889), .B(\w3[7][50] ), .Z(n5314) );
  XOR \MIXCOLUMNS[7].d/U256  ( .A(n5316), .B(n5315), .Z(\w0[8][50] ) );
  XOR \MIXCOLUMNS[7].d/U255  ( .A(n409), .B(n5480), .Z(n5315) );
  XOR \MIXCOLUMNS[7].d/U254  ( .A(\w3[7][58] ), .B(n410), .Z(n5316) );
  XOR \MIXCOLUMNS[7].d/U253  ( .A(n414), .B(n27), .Z(n5475) );
  XOR \MIXCOLUMNS[7].d/U252  ( .A(n5318), .B(n5317), .Z(\w0[8][51] ) );
  XOR \MIXCOLUMNS[7].d/U251  ( .A(n5482), .B(n5319), .Z(n5317) );
  XOR \MIXCOLUMNS[7].d/U250  ( .A(n407), .B(n5475), .Z(n5318) );
  XOR \MIXCOLUMNS[7].d/U249  ( .A(n887), .B(n408), .Z(n5319) );
  XOR \MIXCOLUMNS[7].d/U248  ( .A(n5321), .B(n5320), .Z(\w0[8][52] ) );
  XOR \MIXCOLUMNS[7].d/U247  ( .A(n5484), .B(n5322), .Z(n5320) );
  XOR \MIXCOLUMNS[7].d/U246  ( .A(n405), .B(n5475), .Z(n5321) );
  XOR \MIXCOLUMNS[7].d/U245  ( .A(n885), .B(n406), .Z(n5322) );
  XOR \MIXCOLUMNS[7].d/U244  ( .A(n5324), .B(n5323), .Z(\w0[8][53] ) );
  XOR \MIXCOLUMNS[7].d/U243  ( .A(n403), .B(n5486), .Z(n5323) );
  XOR \MIXCOLUMNS[7].d/U242  ( .A(n883), .B(n404), .Z(n5324) );
  XOR \MIXCOLUMNS[7].d/U241  ( .A(n5326), .B(n5325), .Z(\w0[8][54] ) );
  XOR \MIXCOLUMNS[7].d/U240  ( .A(n5488), .B(n5327), .Z(n5325) );
  XOR \MIXCOLUMNS[7].d/U239  ( .A(n401), .B(n5475), .Z(n5326) );
  XOR \MIXCOLUMNS[7].d/U238  ( .A(n881), .B(n402), .Z(n5327) );
  XOR \MIXCOLUMNS[7].d/U237  ( .A(n5490), .B(n5328), .Z(\w0[8][55] ) );
  XOR \MIXCOLUMNS[7].d/U236  ( .A(n879), .B(n5475), .Z(n5328) );
  XOR \MIXCOLUMNS[7].d/U235  ( .A(n5476), .B(n5329), .Z(\w0[8][56] ) );
  XOR \MIXCOLUMNS[7].d/U234  ( .A(n414), .B(n5477), .Z(n5329) );
  XOR \MIXCOLUMNS[7].d/U233  ( .A(n5478), .B(n5330), .Z(\w0[8][57] ) );
  XOR \MIXCOLUMNS[7].d/U232  ( .A(n413), .B(n5479), .Z(n5330) );
  XOR \MIXCOLUMNS[7].d/U231  ( .A(n5480), .B(n5331), .Z(\w0[8][58] ) );
  XOR \MIXCOLUMNS[7].d/U230  ( .A(\w3[7][50] ), .B(n5481), .Z(n5331) );
  XOR \MIXCOLUMNS[7].d/U229  ( .A(n5333), .B(n5332), .Z(\w0[8][59] ) );
  XOR \MIXCOLUMNS[7].d/U228  ( .A(n5483), .B(n5482), .Z(n5332) );
  XOR \MIXCOLUMNS[7].d/U227  ( .A(n410), .B(n5491), .Z(n5333) );
  XOR \MIXCOLUMNS[7].d/U226  ( .A(n5335), .B(n5334), .Z(\w0[8][60] ) );
  XOR \MIXCOLUMNS[7].d/U225  ( .A(n5485), .B(n5484), .Z(n5334) );
  XOR \MIXCOLUMNS[7].d/U224  ( .A(n408), .B(n5491), .Z(n5335) );
  XOR \MIXCOLUMNS[7].d/U223  ( .A(n5486), .B(n5336), .Z(\w0[8][61] ) );
  XOR \MIXCOLUMNS[7].d/U222  ( .A(n406), .B(n5487), .Z(n5336) );
  XOR \MIXCOLUMNS[7].d/U221  ( .A(n5338), .B(n5337), .Z(\w0[8][62] ) );
  XOR \MIXCOLUMNS[7].d/U220  ( .A(n5489), .B(n5488), .Z(n5337) );
  XOR \MIXCOLUMNS[7].d/U219  ( .A(n404), .B(n5491), .Z(n5338) );
  XOR \MIXCOLUMNS[7].d/U218  ( .A(n5490), .B(n5339), .Z(\w0[8][63] ) );
  XOR \MIXCOLUMNS[7].d/U217  ( .A(n402), .B(n5491), .Z(n5339) );
  XOR \MIXCOLUMNS[7].d/U216  ( .A(n878), .B(n400), .Z(n5509) );
  XOR \MIXCOLUMNS[7].d/U215  ( .A(n5341), .B(n5340), .Z(\w0[8][64] ) );
  XOR \MIXCOLUMNS[7].d/U214  ( .A(n877), .B(n5509), .Z(n5340) );
  XOR \MIXCOLUMNS[7].d/U213  ( .A(n876), .B(n26), .Z(n5341) );
  XOR \MIXCOLUMNS[7].d/U212  ( .A(n876), .B(n399), .Z(n5494) );
  XOR \MIXCOLUMNS[7].d/U211  ( .A(n5343), .B(n5342), .Z(\w0[8][65] ) );
  XOR \MIXCOLUMNS[7].d/U210  ( .A(\w3[7][66] ), .B(n5494), .Z(n5342) );
  XOR \MIXCOLUMNS[7].d/U209  ( .A(\w3[7][90] ), .B(n398), .Z(n5343) );
  XOR \MIXCOLUMNS[7].d/U208  ( .A(\w3[7][90] ), .B(\w3[7][82] ), .Z(n5497) );
  XOR \MIXCOLUMNS[7].d/U207  ( .A(n5345), .B(n5344), .Z(\w0[8][66] ) );
  XOR \MIXCOLUMNS[7].d/U206  ( .A(n875), .B(n5497), .Z(n5344) );
  XOR \MIXCOLUMNS[7].d/U205  ( .A(n874), .B(\w3[7][74] ), .Z(n5345) );
  XOR \MIXCOLUMNS[7].d/U204  ( .A(n878), .B(n397), .Z(n5492) );
  XOR \MIXCOLUMNS[7].d/U203  ( .A(n874), .B(n396), .Z(n5499) );
  XOR \MIXCOLUMNS[7].d/U202  ( .A(n5347), .B(n5346), .Z(\w0[8][67] ) );
  XOR \MIXCOLUMNS[7].d/U201  ( .A(n5499), .B(n5348), .Z(n5346) );
  XOR \MIXCOLUMNS[7].d/U200  ( .A(n873), .B(n5492), .Z(n5347) );
  XOR \MIXCOLUMNS[7].d/U199  ( .A(n872), .B(n395), .Z(n5348) );
  XOR \MIXCOLUMNS[7].d/U198  ( .A(n872), .B(n394), .Z(n5501) );
  XOR \MIXCOLUMNS[7].d/U197  ( .A(n5350), .B(n5349), .Z(\w0[8][68] ) );
  XOR \MIXCOLUMNS[7].d/U196  ( .A(n5501), .B(n5351), .Z(n5349) );
  XOR \MIXCOLUMNS[7].d/U195  ( .A(n871), .B(n5492), .Z(n5350) );
  XOR \MIXCOLUMNS[7].d/U194  ( .A(n870), .B(n393), .Z(n5351) );
  XOR \MIXCOLUMNS[7].d/U193  ( .A(n870), .B(n392), .Z(n5503) );
  XOR \MIXCOLUMNS[7].d/U192  ( .A(n5353), .B(n5352), .Z(\w0[8][69] ) );
  XOR \MIXCOLUMNS[7].d/U191  ( .A(n869), .B(n5503), .Z(n5352) );
  XOR \MIXCOLUMNS[7].d/U190  ( .A(n868), .B(n391), .Z(n5353) );
  XOR \MIXCOLUMNS[7].d/U189  ( .A(n868), .B(n390), .Z(n5505) );
  XOR \MIXCOLUMNS[7].d/U188  ( .A(n5355), .B(n5354), .Z(\w0[8][70] ) );
  XOR \MIXCOLUMNS[7].d/U187  ( .A(n5505), .B(n5356), .Z(n5354) );
  XOR \MIXCOLUMNS[7].d/U186  ( .A(n867), .B(n5492), .Z(n5355) );
  XOR \MIXCOLUMNS[7].d/U185  ( .A(n866), .B(n389), .Z(n5356) );
  XOR \MIXCOLUMNS[7].d/U184  ( .A(n866), .B(n388), .Z(n5507) );
  XOR \MIXCOLUMNS[7].d/U183  ( .A(n5507), .B(n5357), .Z(\w0[8][71] ) );
  XOR \MIXCOLUMNS[7].d/U182  ( .A(n387), .B(n5492), .Z(n5357) );
  XOR \MIXCOLUMNS[7].d/U181  ( .A(n398), .B(n877), .Z(n5496) );
  XOR \MIXCOLUMNS[7].d/U180  ( .A(n5496), .B(n5358), .Z(\w0[8][72] ) );
  XOR \MIXCOLUMNS[7].d/U179  ( .A(n397), .B(n5509), .Z(n5358) );
  XOR \MIXCOLUMNS[7].d/U178  ( .A(\w3[7][74] ), .B(\w3[7][66] ), .Z(n5498) );
  XOR \MIXCOLUMNS[7].d/U177  ( .A(n5498), .B(n5359), .Z(\w0[8][73] ) );
  XOR \MIXCOLUMNS[7].d/U176  ( .A(n877), .B(n5494), .Z(n5359) );
  XOR \MIXCOLUMNS[7].d/U175  ( .A(n395), .B(n875), .Z(n5500) );
  XOR \MIXCOLUMNS[7].d/U174  ( .A(n5500), .B(n5360), .Z(\w0[8][74] ) );
  XOR \MIXCOLUMNS[7].d/U173  ( .A(\w3[7][66] ), .B(n5497), .Z(n5360) );
  XOR \MIXCOLUMNS[7].d/U172  ( .A(n26), .B(n397), .Z(n5495) );
  XOR \MIXCOLUMNS[7].d/U171  ( .A(n393), .B(n873), .Z(n5502) );
  XOR \MIXCOLUMNS[7].d/U170  ( .A(n5362), .B(n5361), .Z(\w0[8][75] ) );
  XOR \MIXCOLUMNS[7].d/U169  ( .A(n5499), .B(n5502), .Z(n5361) );
  XOR \MIXCOLUMNS[7].d/U168  ( .A(n875), .B(n5495), .Z(n5362) );
  XOR \MIXCOLUMNS[7].d/U167  ( .A(n391), .B(n871), .Z(n5504) );
  XOR \MIXCOLUMNS[7].d/U166  ( .A(n5364), .B(n5363), .Z(\w0[8][76] ) );
  XOR \MIXCOLUMNS[7].d/U165  ( .A(n5501), .B(n5504), .Z(n5363) );
  XOR \MIXCOLUMNS[7].d/U164  ( .A(n873), .B(n5495), .Z(n5364) );
  XOR \MIXCOLUMNS[7].d/U163  ( .A(n389), .B(n869), .Z(n5506) );
  XOR \MIXCOLUMNS[7].d/U162  ( .A(n5506), .B(n5365), .Z(\w0[8][77] ) );
  XOR \MIXCOLUMNS[7].d/U161  ( .A(n871), .B(n5503), .Z(n5365) );
  XOR \MIXCOLUMNS[7].d/U160  ( .A(n387), .B(n867), .Z(n5508) );
  XOR \MIXCOLUMNS[7].d/U159  ( .A(n5367), .B(n5366), .Z(\w0[8][78] ) );
  XOR \MIXCOLUMNS[7].d/U158  ( .A(n5505), .B(n5508), .Z(n5366) );
  XOR \MIXCOLUMNS[7].d/U157  ( .A(n869), .B(n5495), .Z(n5367) );
  XOR \MIXCOLUMNS[7].d/U156  ( .A(n5507), .B(n5368), .Z(\w0[8][79] ) );
  XOR \MIXCOLUMNS[7].d/U155  ( .A(n867), .B(n5495), .Z(n5368) );
  XOR \MIXCOLUMNS[7].d/U154  ( .A(n5370), .B(n5369), .Z(\w0[8][80] ) );
  XOR \MIXCOLUMNS[7].d/U153  ( .A(n398), .B(n5495), .Z(n5369) );
  XOR \MIXCOLUMNS[7].d/U152  ( .A(n878), .B(n399), .Z(n5370) );
  XOR \MIXCOLUMNS[7].d/U151  ( .A(n5372), .B(n5371), .Z(\w0[8][81] ) );
  XOR \MIXCOLUMNS[7].d/U150  ( .A(\w3[7][74] ), .B(n5496), .Z(n5371) );
  XOR \MIXCOLUMNS[7].d/U149  ( .A(n876), .B(\w3[7][82] ), .Z(n5372) );
  XOR \MIXCOLUMNS[7].d/U148  ( .A(n5374), .B(n5373), .Z(\w0[8][82] ) );
  XOR \MIXCOLUMNS[7].d/U147  ( .A(n395), .B(n5498), .Z(n5373) );
  XOR \MIXCOLUMNS[7].d/U146  ( .A(\w3[7][90] ), .B(n396), .Z(n5374) );
  XOR \MIXCOLUMNS[7].d/U145  ( .A(n400), .B(n26), .Z(n5493) );
  XOR \MIXCOLUMNS[7].d/U144  ( .A(n5376), .B(n5375), .Z(\w0[8][83] ) );
  XOR \MIXCOLUMNS[7].d/U143  ( .A(n5500), .B(n5377), .Z(n5375) );
  XOR \MIXCOLUMNS[7].d/U142  ( .A(n393), .B(n5493), .Z(n5376) );
  XOR \MIXCOLUMNS[7].d/U141  ( .A(n874), .B(n394), .Z(n5377) );
  XOR \MIXCOLUMNS[7].d/U140  ( .A(n5379), .B(n5378), .Z(\w0[8][84] ) );
  XOR \MIXCOLUMNS[7].d/U139  ( .A(n5502), .B(n5380), .Z(n5378) );
  XOR \MIXCOLUMNS[7].d/U138  ( .A(n391), .B(n5493), .Z(n5379) );
  XOR \MIXCOLUMNS[7].d/U137  ( .A(n872), .B(n392), .Z(n5380) );
  XOR \MIXCOLUMNS[7].d/U136  ( .A(n5382), .B(n5381), .Z(\w0[8][85] ) );
  XOR \MIXCOLUMNS[7].d/U135  ( .A(n389), .B(n5504), .Z(n5381) );
  XOR \MIXCOLUMNS[7].d/U134  ( .A(n870), .B(n390), .Z(n5382) );
  XOR \MIXCOLUMNS[7].d/U133  ( .A(n5384), .B(n5383), .Z(\w0[8][86] ) );
  XOR \MIXCOLUMNS[7].d/U132  ( .A(n5506), .B(n5385), .Z(n5383) );
  XOR \MIXCOLUMNS[7].d/U131  ( .A(n387), .B(n5493), .Z(n5384) );
  XOR \MIXCOLUMNS[7].d/U130  ( .A(n868), .B(n388), .Z(n5385) );
  XOR \MIXCOLUMNS[7].d/U129  ( .A(n5508), .B(n5386), .Z(\w0[8][87] ) );
  XOR \MIXCOLUMNS[7].d/U128  ( .A(n866), .B(n5493), .Z(n5386) );
  XOR \MIXCOLUMNS[7].d/U127  ( .A(n5494), .B(n5387), .Z(\w0[8][88] ) );
  XOR \MIXCOLUMNS[7].d/U126  ( .A(n400), .B(n5495), .Z(n5387) );
  XOR \MIXCOLUMNS[7].d/U125  ( .A(n5496), .B(n5388), .Z(\w0[8][89] ) );
  XOR \MIXCOLUMNS[7].d/U124  ( .A(n399), .B(n5497), .Z(n5388) );
  XOR \MIXCOLUMNS[7].d/U123  ( .A(n5498), .B(n5389), .Z(\w0[8][90] ) );
  XOR \MIXCOLUMNS[7].d/U122  ( .A(\w3[7][82] ), .B(n5499), .Z(n5389) );
  XOR \MIXCOLUMNS[7].d/U121  ( .A(n5391), .B(n5390), .Z(\w0[8][91] ) );
  XOR \MIXCOLUMNS[7].d/U120  ( .A(n5501), .B(n5500), .Z(n5390) );
  XOR \MIXCOLUMNS[7].d/U119  ( .A(n396), .B(n5509), .Z(n5391) );
  XOR \MIXCOLUMNS[7].d/U118  ( .A(n5393), .B(n5392), .Z(\w0[8][92] ) );
  XOR \MIXCOLUMNS[7].d/U117  ( .A(n5503), .B(n5502), .Z(n5392) );
  XOR \MIXCOLUMNS[7].d/U116  ( .A(n394), .B(n5509), .Z(n5393) );
  XOR \MIXCOLUMNS[7].d/U115  ( .A(n5504), .B(n5394), .Z(\w0[8][93] ) );
  XOR \MIXCOLUMNS[7].d/U114  ( .A(n392), .B(n5505), .Z(n5394) );
  XOR \MIXCOLUMNS[7].d/U113  ( .A(n5396), .B(n5395), .Z(\w0[8][94] ) );
  XOR \MIXCOLUMNS[7].d/U112  ( .A(n5507), .B(n5506), .Z(n5395) );
  XOR \MIXCOLUMNS[7].d/U111  ( .A(n390), .B(n5509), .Z(n5396) );
  XOR \MIXCOLUMNS[7].d/U110  ( .A(n5508), .B(n5397), .Z(\w0[8][95] ) );
  XOR \MIXCOLUMNS[7].d/U109  ( .A(n388), .B(n5509), .Z(n5397) );
  XOR \MIXCOLUMNS[7].d/U108  ( .A(n865), .B(n386), .Z(n5527) );
  XOR \MIXCOLUMNS[7].d/U107  ( .A(n5399), .B(n5398), .Z(\w0[8][96] ) );
  XOR \MIXCOLUMNS[7].d/U106  ( .A(n864), .B(n5527), .Z(n5398) );
  XOR \MIXCOLUMNS[7].d/U105  ( .A(n863), .B(n25), .Z(n5399) );
  XOR \MIXCOLUMNS[7].d/U104  ( .A(n863), .B(n385), .Z(n5512) );
  XOR \MIXCOLUMNS[7].d/U103  ( .A(n5401), .B(n5400), .Z(\w0[8][97] ) );
  XOR \MIXCOLUMNS[7].d/U102  ( .A(\w3[7][98] ), .B(n5512), .Z(n5400) );
  XOR \MIXCOLUMNS[7].d/U101  ( .A(\w3[7][122] ), .B(n384), .Z(n5401) );
  XOR \MIXCOLUMNS[7].d/U100  ( .A(\w3[7][122] ), .B(\w3[7][114] ), .Z(n5515)
         );
  XOR \MIXCOLUMNS[7].d/U99  ( .A(n5403), .B(n5402), .Z(\w0[8][98] ) );
  XOR \MIXCOLUMNS[7].d/U98  ( .A(n862), .B(n5515), .Z(n5402) );
  XOR \MIXCOLUMNS[7].d/U97  ( .A(n861), .B(\w3[7][106] ), .Z(n5403) );
  XOR \MIXCOLUMNS[7].d/U96  ( .A(n865), .B(n383), .Z(n5510) );
  XOR \MIXCOLUMNS[7].d/U95  ( .A(n861), .B(n382), .Z(n5517) );
  XOR \MIXCOLUMNS[7].d/U94  ( .A(n5405), .B(n5404), .Z(\w0[8][99] ) );
  XOR \MIXCOLUMNS[7].d/U93  ( .A(n5517), .B(n5406), .Z(n5404) );
  XOR \MIXCOLUMNS[7].d/U92  ( .A(n860), .B(n5510), .Z(n5405) );
  XOR \MIXCOLUMNS[7].d/U91  ( .A(n859), .B(n381), .Z(n5406) );
  XOR \MIXCOLUMNS[7].d/U90  ( .A(n859), .B(n380), .Z(n5519) );
  XOR \MIXCOLUMNS[7].d/U89  ( .A(n5408), .B(n5407), .Z(\w0[8][100] ) );
  XOR \MIXCOLUMNS[7].d/U88  ( .A(n5519), .B(n5409), .Z(n5407) );
  XOR \MIXCOLUMNS[7].d/U87  ( .A(n858), .B(n5510), .Z(n5408) );
  XOR \MIXCOLUMNS[7].d/U86  ( .A(n857), .B(n379), .Z(n5409) );
  XOR \MIXCOLUMNS[7].d/U85  ( .A(n857), .B(n378), .Z(n5521) );
  XOR \MIXCOLUMNS[7].d/U84  ( .A(n5411), .B(n5410), .Z(\w0[8][101] ) );
  XOR \MIXCOLUMNS[7].d/U83  ( .A(n856), .B(n5521), .Z(n5410) );
  XOR \MIXCOLUMNS[7].d/U82  ( .A(n855), .B(n377), .Z(n5411) );
  XOR \MIXCOLUMNS[7].d/U81  ( .A(n855), .B(n376), .Z(n5523) );
  XOR \MIXCOLUMNS[7].d/U80  ( .A(n5413), .B(n5412), .Z(\w0[8][102] ) );
  XOR \MIXCOLUMNS[7].d/U79  ( .A(n5523), .B(n5414), .Z(n5412) );
  XOR \MIXCOLUMNS[7].d/U78  ( .A(n854), .B(n5510), .Z(n5413) );
  XOR \MIXCOLUMNS[7].d/U77  ( .A(n853), .B(n375), .Z(n5414) );
  XOR \MIXCOLUMNS[7].d/U76  ( .A(n853), .B(n374), .Z(n5525) );
  XOR \MIXCOLUMNS[7].d/U75  ( .A(n5525), .B(n5415), .Z(\w0[8][103] ) );
  XOR \MIXCOLUMNS[7].d/U74  ( .A(n373), .B(n5510), .Z(n5415) );
  XOR \MIXCOLUMNS[7].d/U73  ( .A(n384), .B(n864), .Z(n5514) );
  XOR \MIXCOLUMNS[7].d/U72  ( .A(n5514), .B(n5416), .Z(\w0[8][104] ) );
  XOR \MIXCOLUMNS[7].d/U71  ( .A(n383), .B(n5527), .Z(n5416) );
  XOR \MIXCOLUMNS[7].d/U70  ( .A(\w3[7][106] ), .B(\w3[7][98] ), .Z(n5516) );
  XOR \MIXCOLUMNS[7].d/U69  ( .A(n5516), .B(n5417), .Z(\w0[8][105] ) );
  XOR \MIXCOLUMNS[7].d/U68  ( .A(n864), .B(n5512), .Z(n5417) );
  XOR \MIXCOLUMNS[7].d/U67  ( .A(n381), .B(n862), .Z(n5518) );
  XOR \MIXCOLUMNS[7].d/U66  ( .A(n5518), .B(n5418), .Z(\w0[8][106] ) );
  XOR \MIXCOLUMNS[7].d/U65  ( .A(\w3[7][98] ), .B(n5515), .Z(n5418) );
  XOR \MIXCOLUMNS[7].d/U64  ( .A(n25), .B(n383), .Z(n5513) );
  XOR \MIXCOLUMNS[7].d/U63  ( .A(n379), .B(n860), .Z(n5520) );
  XOR \MIXCOLUMNS[7].d/U62  ( .A(n5420), .B(n5419), .Z(\w0[8][107] ) );
  XOR \MIXCOLUMNS[7].d/U61  ( .A(n5517), .B(n5520), .Z(n5419) );
  XOR \MIXCOLUMNS[7].d/U60  ( .A(n862), .B(n5513), .Z(n5420) );
  XOR \MIXCOLUMNS[7].d/U59  ( .A(n377), .B(n858), .Z(n5522) );
  XOR \MIXCOLUMNS[7].d/U58  ( .A(n5422), .B(n5421), .Z(\w0[8][108] ) );
  XOR \MIXCOLUMNS[7].d/U57  ( .A(n5519), .B(n5522), .Z(n5421) );
  XOR \MIXCOLUMNS[7].d/U56  ( .A(n860), .B(n5513), .Z(n5422) );
  XOR \MIXCOLUMNS[7].d/U55  ( .A(n375), .B(n856), .Z(n5524) );
  XOR \MIXCOLUMNS[7].d/U54  ( .A(n5524), .B(n5423), .Z(\w0[8][109] ) );
  XOR \MIXCOLUMNS[7].d/U53  ( .A(n858), .B(n5521), .Z(n5423) );
  XOR \MIXCOLUMNS[7].d/U52  ( .A(n373), .B(n854), .Z(n5526) );
  XOR \MIXCOLUMNS[7].d/U51  ( .A(n5425), .B(n5424), .Z(\w0[8][110] ) );
  XOR \MIXCOLUMNS[7].d/U50  ( .A(n5523), .B(n5526), .Z(n5424) );
  XOR \MIXCOLUMNS[7].d/U49  ( .A(n856), .B(n5513), .Z(n5425) );
  XOR \MIXCOLUMNS[7].d/U48  ( .A(n5525), .B(n5426), .Z(\w0[8][111] ) );
  XOR \MIXCOLUMNS[7].d/U47  ( .A(n854), .B(n5513), .Z(n5426) );
  XOR \MIXCOLUMNS[7].d/U46  ( .A(n5428), .B(n5427), .Z(\w0[8][112] ) );
  XOR \MIXCOLUMNS[7].d/U45  ( .A(n384), .B(n5513), .Z(n5427) );
  XOR \MIXCOLUMNS[7].d/U44  ( .A(n865), .B(n385), .Z(n5428) );
  XOR \MIXCOLUMNS[7].d/U43  ( .A(n5430), .B(n5429), .Z(\w0[8][113] ) );
  XOR \MIXCOLUMNS[7].d/U42  ( .A(\w3[7][106] ), .B(n5514), .Z(n5429) );
  XOR \MIXCOLUMNS[7].d/U41  ( .A(n863), .B(\w3[7][114] ), .Z(n5430) );
  XOR \MIXCOLUMNS[7].d/U40  ( .A(n5432), .B(n5431), .Z(\w0[8][114] ) );
  XOR \MIXCOLUMNS[7].d/U39  ( .A(n381), .B(n5516), .Z(n5431) );
  XOR \MIXCOLUMNS[7].d/U38  ( .A(\w3[7][122] ), .B(n382), .Z(n5432) );
  XOR \MIXCOLUMNS[7].d/U37  ( .A(n386), .B(n25), .Z(n5511) );
  XOR \MIXCOLUMNS[7].d/U36  ( .A(n5434), .B(n5433), .Z(\w0[8][115] ) );
  XOR \MIXCOLUMNS[7].d/U35  ( .A(n5518), .B(n5435), .Z(n5433) );
  XOR \MIXCOLUMNS[7].d/U34  ( .A(n379), .B(n5511), .Z(n5434) );
  XOR \MIXCOLUMNS[7].d/U33  ( .A(n861), .B(n380), .Z(n5435) );
  XOR \MIXCOLUMNS[7].d/U32  ( .A(n5437), .B(n5436), .Z(\w0[8][116] ) );
  XOR \MIXCOLUMNS[7].d/U31  ( .A(n5520), .B(n5438), .Z(n5436) );
  XOR \MIXCOLUMNS[7].d/U30  ( .A(n377), .B(n5511), .Z(n5437) );
  XOR \MIXCOLUMNS[7].d/U29  ( .A(n859), .B(n378), .Z(n5438) );
  XOR \MIXCOLUMNS[7].d/U28  ( .A(n5440), .B(n5439), .Z(\w0[8][117] ) );
  XOR \MIXCOLUMNS[7].d/U27  ( .A(n375), .B(n5522), .Z(n5439) );
  XOR \MIXCOLUMNS[7].d/U26  ( .A(n857), .B(n376), .Z(n5440) );
  XOR \MIXCOLUMNS[7].d/U25  ( .A(n5442), .B(n5441), .Z(\w0[8][118] ) );
  XOR \MIXCOLUMNS[7].d/U24  ( .A(n5524), .B(n5443), .Z(n5441) );
  XOR \MIXCOLUMNS[7].d/U23  ( .A(n373), .B(n5511), .Z(n5442) );
  XOR \MIXCOLUMNS[7].d/U22  ( .A(n855), .B(n374), .Z(n5443) );
  XOR \MIXCOLUMNS[7].d/U21  ( .A(n5526), .B(n5444), .Z(\w0[8][119] ) );
  XOR \MIXCOLUMNS[7].d/U20  ( .A(n853), .B(n5511), .Z(n5444) );
  XOR \MIXCOLUMNS[7].d/U19  ( .A(n5512), .B(n5445), .Z(\w0[8][120] ) );
  XOR \MIXCOLUMNS[7].d/U18  ( .A(n386), .B(n5513), .Z(n5445) );
  XOR \MIXCOLUMNS[7].d/U17  ( .A(n5514), .B(n5446), .Z(\w0[8][121] ) );
  XOR \MIXCOLUMNS[7].d/U16  ( .A(n385), .B(n5515), .Z(n5446) );
  XOR \MIXCOLUMNS[7].d/U15  ( .A(n5516), .B(n5447), .Z(\w0[8][122] ) );
  XOR \MIXCOLUMNS[7].d/U14  ( .A(\w3[7][114] ), .B(n5517), .Z(n5447) );
  XOR \MIXCOLUMNS[7].d/U13  ( .A(n5449), .B(n5448), .Z(\w0[8][123] ) );
  XOR \MIXCOLUMNS[7].d/U12  ( .A(n5519), .B(n5518), .Z(n5448) );
  XOR \MIXCOLUMNS[7].d/U11  ( .A(n382), .B(n5527), .Z(n5449) );
  XOR \MIXCOLUMNS[7].d/U10  ( .A(n5451), .B(n5450), .Z(\w0[8][124] ) );
  XOR \MIXCOLUMNS[7].d/U9  ( .A(n5521), .B(n5520), .Z(n5450) );
  XOR \MIXCOLUMNS[7].d/U8  ( .A(n380), .B(n5527), .Z(n5451) );
  XOR \MIXCOLUMNS[7].d/U7  ( .A(n5522), .B(n5452), .Z(\w0[8][125] ) );
  XOR \MIXCOLUMNS[7].d/U6  ( .A(n378), .B(n5523), .Z(n5452) );
  XOR \MIXCOLUMNS[7].d/U5  ( .A(n5454), .B(n5453), .Z(\w0[8][126] ) );
  XOR \MIXCOLUMNS[7].d/U4  ( .A(n5525), .B(n5524), .Z(n5453) );
  XOR \MIXCOLUMNS[7].d/U3  ( .A(n376), .B(n5527), .Z(n5454) );
  XOR \MIXCOLUMNS[7].d/U2  ( .A(n5526), .B(n5455), .Z(\w0[8][127] ) );
  XOR \MIXCOLUMNS[7].d/U1  ( .A(n374), .B(n5527), .Z(n5455) );
  XOR \MIXCOLUMNS[6].d/U432  ( .A(n852), .B(n372), .Z(n5169) );
  XOR \MIXCOLUMNS[6].d/U431  ( .A(n4921), .B(n4920), .Z(\w0[7][0] ) );
  XOR \MIXCOLUMNS[6].d/U430  ( .A(n851), .B(n5169), .Z(n4920) );
  XOR \MIXCOLUMNS[6].d/U429  ( .A(n850), .B(n24), .Z(n4921) );
  XOR \MIXCOLUMNS[6].d/U428  ( .A(n850), .B(n371), .Z(n5154) );
  XOR \MIXCOLUMNS[6].d/U427  ( .A(n4923), .B(n4922), .Z(\w0[7][1] ) );
  XOR \MIXCOLUMNS[6].d/U426  ( .A(\w3[6][2] ), .B(n5154), .Z(n4922) );
  XOR \MIXCOLUMNS[6].d/U425  ( .A(\w3[6][26] ), .B(n370), .Z(n4923) );
  XOR \MIXCOLUMNS[6].d/U424  ( .A(\w3[6][26] ), .B(\w3[6][18] ), .Z(n5157) );
  XOR \MIXCOLUMNS[6].d/U423  ( .A(n4925), .B(n4924), .Z(\w0[7][2] ) );
  XOR \MIXCOLUMNS[6].d/U422  ( .A(n849), .B(n5157), .Z(n4924) );
  XOR \MIXCOLUMNS[6].d/U421  ( .A(n848), .B(\w3[6][10] ), .Z(n4925) );
  XOR \MIXCOLUMNS[6].d/U420  ( .A(n852), .B(n369), .Z(n5152) );
  XOR \MIXCOLUMNS[6].d/U419  ( .A(n848), .B(n368), .Z(n5159) );
  XOR \MIXCOLUMNS[6].d/U418  ( .A(n4927), .B(n4926), .Z(\w0[7][3] ) );
  XOR \MIXCOLUMNS[6].d/U417  ( .A(n5159), .B(n4928), .Z(n4926) );
  XOR \MIXCOLUMNS[6].d/U416  ( .A(n847), .B(n5152), .Z(n4927) );
  XOR \MIXCOLUMNS[6].d/U415  ( .A(n846), .B(n367), .Z(n4928) );
  XOR \MIXCOLUMNS[6].d/U414  ( .A(n846), .B(n366), .Z(n5161) );
  XOR \MIXCOLUMNS[6].d/U413  ( .A(n4930), .B(n4929), .Z(\w0[7][4] ) );
  XOR \MIXCOLUMNS[6].d/U412  ( .A(n5161), .B(n4931), .Z(n4929) );
  XOR \MIXCOLUMNS[6].d/U411  ( .A(n845), .B(n5152), .Z(n4930) );
  XOR \MIXCOLUMNS[6].d/U410  ( .A(n844), .B(n365), .Z(n4931) );
  XOR \MIXCOLUMNS[6].d/U409  ( .A(n844), .B(n364), .Z(n5163) );
  XOR \MIXCOLUMNS[6].d/U408  ( .A(n4933), .B(n4932), .Z(\w0[7][5] ) );
  XOR \MIXCOLUMNS[6].d/U407  ( .A(n843), .B(n5163), .Z(n4932) );
  XOR \MIXCOLUMNS[6].d/U406  ( .A(n842), .B(n363), .Z(n4933) );
  XOR \MIXCOLUMNS[6].d/U405  ( .A(n842), .B(n362), .Z(n5165) );
  XOR \MIXCOLUMNS[6].d/U404  ( .A(n4935), .B(n4934), .Z(\w0[7][6] ) );
  XOR \MIXCOLUMNS[6].d/U403  ( .A(n5165), .B(n4936), .Z(n4934) );
  XOR \MIXCOLUMNS[6].d/U402  ( .A(n841), .B(n5152), .Z(n4935) );
  XOR \MIXCOLUMNS[6].d/U401  ( .A(n840), .B(n361), .Z(n4936) );
  XOR \MIXCOLUMNS[6].d/U400  ( .A(n840), .B(n360), .Z(n5167) );
  XOR \MIXCOLUMNS[6].d/U399  ( .A(n5167), .B(n4937), .Z(\w0[7][7] ) );
  XOR \MIXCOLUMNS[6].d/U398  ( .A(n359), .B(n5152), .Z(n4937) );
  XOR \MIXCOLUMNS[6].d/U397  ( .A(n370), .B(n851), .Z(n5156) );
  XOR \MIXCOLUMNS[6].d/U396  ( .A(n5156), .B(n4938), .Z(\w0[7][8] ) );
  XOR \MIXCOLUMNS[6].d/U395  ( .A(n369), .B(n5169), .Z(n4938) );
  XOR \MIXCOLUMNS[6].d/U394  ( .A(\w3[6][10] ), .B(\w3[6][2] ), .Z(n5158) );
  XOR \MIXCOLUMNS[6].d/U393  ( .A(n5158), .B(n4939), .Z(\w0[7][9] ) );
  XOR \MIXCOLUMNS[6].d/U392  ( .A(n851), .B(n5154), .Z(n4939) );
  XOR \MIXCOLUMNS[6].d/U391  ( .A(n367), .B(n849), .Z(n5160) );
  XOR \MIXCOLUMNS[6].d/U390  ( .A(n5160), .B(n4940), .Z(\w0[7][10] ) );
  XOR \MIXCOLUMNS[6].d/U389  ( .A(\w3[6][2] ), .B(n5157), .Z(n4940) );
  XOR \MIXCOLUMNS[6].d/U388  ( .A(n24), .B(n369), .Z(n5155) );
  XOR \MIXCOLUMNS[6].d/U387  ( .A(n365), .B(n847), .Z(n5162) );
  XOR \MIXCOLUMNS[6].d/U386  ( .A(n4942), .B(n4941), .Z(\w0[7][11] ) );
  XOR \MIXCOLUMNS[6].d/U385  ( .A(n5159), .B(n5162), .Z(n4941) );
  XOR \MIXCOLUMNS[6].d/U384  ( .A(n849), .B(n5155), .Z(n4942) );
  XOR \MIXCOLUMNS[6].d/U383  ( .A(n363), .B(n845), .Z(n5164) );
  XOR \MIXCOLUMNS[6].d/U382  ( .A(n4944), .B(n4943), .Z(\w0[7][12] ) );
  XOR \MIXCOLUMNS[6].d/U381  ( .A(n5161), .B(n5164), .Z(n4943) );
  XOR \MIXCOLUMNS[6].d/U380  ( .A(n847), .B(n5155), .Z(n4944) );
  XOR \MIXCOLUMNS[6].d/U379  ( .A(n361), .B(n843), .Z(n5166) );
  XOR \MIXCOLUMNS[6].d/U378  ( .A(n5166), .B(n4945), .Z(\w0[7][13] ) );
  XOR \MIXCOLUMNS[6].d/U377  ( .A(n845), .B(n5163), .Z(n4945) );
  XOR \MIXCOLUMNS[6].d/U376  ( .A(n359), .B(n841), .Z(n5168) );
  XOR \MIXCOLUMNS[6].d/U375  ( .A(n4947), .B(n4946), .Z(\w0[7][14] ) );
  XOR \MIXCOLUMNS[6].d/U374  ( .A(n5165), .B(n5168), .Z(n4946) );
  XOR \MIXCOLUMNS[6].d/U373  ( .A(n843), .B(n5155), .Z(n4947) );
  XOR \MIXCOLUMNS[6].d/U372  ( .A(n5167), .B(n4948), .Z(\w0[7][15] ) );
  XOR \MIXCOLUMNS[6].d/U371  ( .A(n841), .B(n5155), .Z(n4948) );
  XOR \MIXCOLUMNS[6].d/U370  ( .A(n4950), .B(n4949), .Z(\w0[7][16] ) );
  XOR \MIXCOLUMNS[6].d/U369  ( .A(n370), .B(n5155), .Z(n4949) );
  XOR \MIXCOLUMNS[6].d/U368  ( .A(n852), .B(n371), .Z(n4950) );
  XOR \MIXCOLUMNS[6].d/U367  ( .A(n4952), .B(n4951), .Z(\w0[7][17] ) );
  XOR \MIXCOLUMNS[6].d/U366  ( .A(\w3[6][10] ), .B(n5156), .Z(n4951) );
  XOR \MIXCOLUMNS[6].d/U365  ( .A(n850), .B(\w3[6][18] ), .Z(n4952) );
  XOR \MIXCOLUMNS[6].d/U364  ( .A(n4954), .B(n4953), .Z(\w0[7][18] ) );
  XOR \MIXCOLUMNS[6].d/U363  ( .A(n367), .B(n5158), .Z(n4953) );
  XOR \MIXCOLUMNS[6].d/U362  ( .A(\w3[6][26] ), .B(n368), .Z(n4954) );
  XOR \MIXCOLUMNS[6].d/U361  ( .A(n372), .B(n24), .Z(n5153) );
  XOR \MIXCOLUMNS[6].d/U360  ( .A(n4956), .B(n4955), .Z(\w0[7][19] ) );
  XOR \MIXCOLUMNS[6].d/U359  ( .A(n5160), .B(n4957), .Z(n4955) );
  XOR \MIXCOLUMNS[6].d/U358  ( .A(n365), .B(n5153), .Z(n4956) );
  XOR \MIXCOLUMNS[6].d/U357  ( .A(n848), .B(n366), .Z(n4957) );
  XOR \MIXCOLUMNS[6].d/U356  ( .A(n4959), .B(n4958), .Z(\w0[7][20] ) );
  XOR \MIXCOLUMNS[6].d/U355  ( .A(n5162), .B(n4960), .Z(n4958) );
  XOR \MIXCOLUMNS[6].d/U354  ( .A(n363), .B(n5153), .Z(n4959) );
  XOR \MIXCOLUMNS[6].d/U353  ( .A(n846), .B(n364), .Z(n4960) );
  XOR \MIXCOLUMNS[6].d/U352  ( .A(n4962), .B(n4961), .Z(\w0[7][21] ) );
  XOR \MIXCOLUMNS[6].d/U351  ( .A(n361), .B(n5164), .Z(n4961) );
  XOR \MIXCOLUMNS[6].d/U350  ( .A(n844), .B(n362), .Z(n4962) );
  XOR \MIXCOLUMNS[6].d/U349  ( .A(n4964), .B(n4963), .Z(\w0[7][22] ) );
  XOR \MIXCOLUMNS[6].d/U348  ( .A(n5166), .B(n4965), .Z(n4963) );
  XOR \MIXCOLUMNS[6].d/U347  ( .A(n359), .B(n5153), .Z(n4964) );
  XOR \MIXCOLUMNS[6].d/U346  ( .A(n842), .B(n360), .Z(n4965) );
  XOR \MIXCOLUMNS[6].d/U345  ( .A(n5168), .B(n4966), .Z(\w0[7][23] ) );
  XOR \MIXCOLUMNS[6].d/U344  ( .A(n840), .B(n5153), .Z(n4966) );
  XOR \MIXCOLUMNS[6].d/U343  ( .A(n5154), .B(n4967), .Z(\w0[7][24] ) );
  XOR \MIXCOLUMNS[6].d/U342  ( .A(n372), .B(n5155), .Z(n4967) );
  XOR \MIXCOLUMNS[6].d/U341  ( .A(n5156), .B(n4968), .Z(\w0[7][25] ) );
  XOR \MIXCOLUMNS[6].d/U340  ( .A(n371), .B(n5157), .Z(n4968) );
  XOR \MIXCOLUMNS[6].d/U339  ( .A(n5158), .B(n4969), .Z(\w0[7][26] ) );
  XOR \MIXCOLUMNS[6].d/U338  ( .A(\w3[6][18] ), .B(n5159), .Z(n4969) );
  XOR \MIXCOLUMNS[6].d/U337  ( .A(n4971), .B(n4970), .Z(\w0[7][27] ) );
  XOR \MIXCOLUMNS[6].d/U336  ( .A(n5161), .B(n5160), .Z(n4970) );
  XOR \MIXCOLUMNS[6].d/U335  ( .A(n368), .B(n5169), .Z(n4971) );
  XOR \MIXCOLUMNS[6].d/U334  ( .A(n4973), .B(n4972), .Z(\w0[7][28] ) );
  XOR \MIXCOLUMNS[6].d/U333  ( .A(n5163), .B(n5162), .Z(n4972) );
  XOR \MIXCOLUMNS[6].d/U332  ( .A(n366), .B(n5169), .Z(n4973) );
  XOR \MIXCOLUMNS[6].d/U331  ( .A(n5164), .B(n4974), .Z(\w0[7][29] ) );
  XOR \MIXCOLUMNS[6].d/U330  ( .A(n364), .B(n5165), .Z(n4974) );
  XOR \MIXCOLUMNS[6].d/U329  ( .A(n4976), .B(n4975), .Z(\w0[7][30] ) );
  XOR \MIXCOLUMNS[6].d/U328  ( .A(n5167), .B(n5166), .Z(n4975) );
  XOR \MIXCOLUMNS[6].d/U327  ( .A(n362), .B(n5169), .Z(n4976) );
  XOR \MIXCOLUMNS[6].d/U326  ( .A(n5168), .B(n4977), .Z(\w0[7][31] ) );
  XOR \MIXCOLUMNS[6].d/U325  ( .A(n360), .B(n5169), .Z(n4977) );
  XOR \MIXCOLUMNS[6].d/U324  ( .A(n839), .B(n358), .Z(n5187) );
  XOR \MIXCOLUMNS[6].d/U323  ( .A(n4979), .B(n4978), .Z(\w0[7][32] ) );
  XOR \MIXCOLUMNS[6].d/U322  ( .A(n838), .B(n5187), .Z(n4978) );
  XOR \MIXCOLUMNS[6].d/U321  ( .A(n837), .B(n23), .Z(n4979) );
  XOR \MIXCOLUMNS[6].d/U320  ( .A(n837), .B(n357), .Z(n5172) );
  XOR \MIXCOLUMNS[6].d/U319  ( .A(n4981), .B(n4980), .Z(\w0[7][33] ) );
  XOR \MIXCOLUMNS[6].d/U318  ( .A(\w3[6][34] ), .B(n5172), .Z(n4980) );
  XOR \MIXCOLUMNS[6].d/U317  ( .A(\w3[6][58] ), .B(n356), .Z(n4981) );
  XOR \MIXCOLUMNS[6].d/U316  ( .A(\w3[6][58] ), .B(\w3[6][50] ), .Z(n5175) );
  XOR \MIXCOLUMNS[6].d/U315  ( .A(n4983), .B(n4982), .Z(\w0[7][34] ) );
  XOR \MIXCOLUMNS[6].d/U314  ( .A(n836), .B(n5175), .Z(n4982) );
  XOR \MIXCOLUMNS[6].d/U313  ( .A(n835), .B(\w3[6][42] ), .Z(n4983) );
  XOR \MIXCOLUMNS[6].d/U312  ( .A(n839), .B(n355), .Z(n5170) );
  XOR \MIXCOLUMNS[6].d/U311  ( .A(n835), .B(n354), .Z(n5177) );
  XOR \MIXCOLUMNS[6].d/U310  ( .A(n4985), .B(n4984), .Z(\w0[7][35] ) );
  XOR \MIXCOLUMNS[6].d/U309  ( .A(n5177), .B(n4986), .Z(n4984) );
  XOR \MIXCOLUMNS[6].d/U308  ( .A(n834), .B(n5170), .Z(n4985) );
  XOR \MIXCOLUMNS[6].d/U307  ( .A(n833), .B(n353), .Z(n4986) );
  XOR \MIXCOLUMNS[6].d/U306  ( .A(n833), .B(n352), .Z(n5179) );
  XOR \MIXCOLUMNS[6].d/U305  ( .A(n4988), .B(n4987), .Z(\w0[7][36] ) );
  XOR \MIXCOLUMNS[6].d/U304  ( .A(n5179), .B(n4989), .Z(n4987) );
  XOR \MIXCOLUMNS[6].d/U303  ( .A(n832), .B(n5170), .Z(n4988) );
  XOR \MIXCOLUMNS[6].d/U302  ( .A(n831), .B(n351), .Z(n4989) );
  XOR \MIXCOLUMNS[6].d/U301  ( .A(n831), .B(n350), .Z(n5181) );
  XOR \MIXCOLUMNS[6].d/U300  ( .A(n4991), .B(n4990), .Z(\w0[7][37] ) );
  XOR \MIXCOLUMNS[6].d/U299  ( .A(n830), .B(n5181), .Z(n4990) );
  XOR \MIXCOLUMNS[6].d/U298  ( .A(n829), .B(n349), .Z(n4991) );
  XOR \MIXCOLUMNS[6].d/U297  ( .A(n829), .B(n348), .Z(n5183) );
  XOR \MIXCOLUMNS[6].d/U296  ( .A(n4993), .B(n4992), .Z(\w0[7][38] ) );
  XOR \MIXCOLUMNS[6].d/U295  ( .A(n5183), .B(n4994), .Z(n4992) );
  XOR \MIXCOLUMNS[6].d/U294  ( .A(n828), .B(n5170), .Z(n4993) );
  XOR \MIXCOLUMNS[6].d/U293  ( .A(n827), .B(n347), .Z(n4994) );
  XOR \MIXCOLUMNS[6].d/U292  ( .A(n827), .B(n346), .Z(n5185) );
  XOR \MIXCOLUMNS[6].d/U291  ( .A(n5185), .B(n4995), .Z(\w0[7][39] ) );
  XOR \MIXCOLUMNS[6].d/U290  ( .A(n345), .B(n5170), .Z(n4995) );
  XOR \MIXCOLUMNS[6].d/U289  ( .A(n356), .B(n838), .Z(n5174) );
  XOR \MIXCOLUMNS[6].d/U288  ( .A(n5174), .B(n4996), .Z(\w0[7][40] ) );
  XOR \MIXCOLUMNS[6].d/U287  ( .A(n355), .B(n5187), .Z(n4996) );
  XOR \MIXCOLUMNS[6].d/U286  ( .A(\w3[6][42] ), .B(\w3[6][34] ), .Z(n5176) );
  XOR \MIXCOLUMNS[6].d/U285  ( .A(n5176), .B(n4997), .Z(\w0[7][41] ) );
  XOR \MIXCOLUMNS[6].d/U284  ( .A(n838), .B(n5172), .Z(n4997) );
  XOR \MIXCOLUMNS[6].d/U283  ( .A(n353), .B(n836), .Z(n5178) );
  XOR \MIXCOLUMNS[6].d/U282  ( .A(n5178), .B(n4998), .Z(\w0[7][42] ) );
  XOR \MIXCOLUMNS[6].d/U281  ( .A(\w3[6][34] ), .B(n5175), .Z(n4998) );
  XOR \MIXCOLUMNS[6].d/U280  ( .A(n23), .B(n355), .Z(n5173) );
  XOR \MIXCOLUMNS[6].d/U279  ( .A(n351), .B(n834), .Z(n5180) );
  XOR \MIXCOLUMNS[6].d/U278  ( .A(n5000), .B(n4999), .Z(\w0[7][43] ) );
  XOR \MIXCOLUMNS[6].d/U277  ( .A(n5177), .B(n5180), .Z(n4999) );
  XOR \MIXCOLUMNS[6].d/U276  ( .A(n836), .B(n5173), .Z(n5000) );
  XOR \MIXCOLUMNS[6].d/U275  ( .A(n349), .B(n832), .Z(n5182) );
  XOR \MIXCOLUMNS[6].d/U274  ( .A(n5002), .B(n5001), .Z(\w0[7][44] ) );
  XOR \MIXCOLUMNS[6].d/U273  ( .A(n5179), .B(n5182), .Z(n5001) );
  XOR \MIXCOLUMNS[6].d/U272  ( .A(n834), .B(n5173), .Z(n5002) );
  XOR \MIXCOLUMNS[6].d/U271  ( .A(n347), .B(n830), .Z(n5184) );
  XOR \MIXCOLUMNS[6].d/U270  ( .A(n5184), .B(n5003), .Z(\w0[7][45] ) );
  XOR \MIXCOLUMNS[6].d/U269  ( .A(n832), .B(n5181), .Z(n5003) );
  XOR \MIXCOLUMNS[6].d/U268  ( .A(n345), .B(n828), .Z(n5186) );
  XOR \MIXCOLUMNS[6].d/U267  ( .A(n5005), .B(n5004), .Z(\w0[7][46] ) );
  XOR \MIXCOLUMNS[6].d/U266  ( .A(n5183), .B(n5186), .Z(n5004) );
  XOR \MIXCOLUMNS[6].d/U265  ( .A(n830), .B(n5173), .Z(n5005) );
  XOR \MIXCOLUMNS[6].d/U264  ( .A(n5185), .B(n5006), .Z(\w0[7][47] ) );
  XOR \MIXCOLUMNS[6].d/U263  ( .A(n828), .B(n5173), .Z(n5006) );
  XOR \MIXCOLUMNS[6].d/U262  ( .A(n5008), .B(n5007), .Z(\w0[7][48] ) );
  XOR \MIXCOLUMNS[6].d/U261  ( .A(n356), .B(n5173), .Z(n5007) );
  XOR \MIXCOLUMNS[6].d/U260  ( .A(n839), .B(n357), .Z(n5008) );
  XOR \MIXCOLUMNS[6].d/U259  ( .A(n5010), .B(n5009), .Z(\w0[7][49] ) );
  XOR \MIXCOLUMNS[6].d/U258  ( .A(\w3[6][42] ), .B(n5174), .Z(n5009) );
  XOR \MIXCOLUMNS[6].d/U257  ( .A(n837), .B(\w3[6][50] ), .Z(n5010) );
  XOR \MIXCOLUMNS[6].d/U256  ( .A(n5012), .B(n5011), .Z(\w0[7][50] ) );
  XOR \MIXCOLUMNS[6].d/U255  ( .A(n353), .B(n5176), .Z(n5011) );
  XOR \MIXCOLUMNS[6].d/U254  ( .A(\w3[6][58] ), .B(n354), .Z(n5012) );
  XOR \MIXCOLUMNS[6].d/U253  ( .A(n358), .B(n23), .Z(n5171) );
  XOR \MIXCOLUMNS[6].d/U252  ( .A(n5014), .B(n5013), .Z(\w0[7][51] ) );
  XOR \MIXCOLUMNS[6].d/U251  ( .A(n5178), .B(n5015), .Z(n5013) );
  XOR \MIXCOLUMNS[6].d/U250  ( .A(n351), .B(n5171), .Z(n5014) );
  XOR \MIXCOLUMNS[6].d/U249  ( .A(n835), .B(n352), .Z(n5015) );
  XOR \MIXCOLUMNS[6].d/U248  ( .A(n5017), .B(n5016), .Z(\w0[7][52] ) );
  XOR \MIXCOLUMNS[6].d/U247  ( .A(n5180), .B(n5018), .Z(n5016) );
  XOR \MIXCOLUMNS[6].d/U246  ( .A(n349), .B(n5171), .Z(n5017) );
  XOR \MIXCOLUMNS[6].d/U245  ( .A(n833), .B(n350), .Z(n5018) );
  XOR \MIXCOLUMNS[6].d/U244  ( .A(n5020), .B(n5019), .Z(\w0[7][53] ) );
  XOR \MIXCOLUMNS[6].d/U243  ( .A(n347), .B(n5182), .Z(n5019) );
  XOR \MIXCOLUMNS[6].d/U242  ( .A(n831), .B(n348), .Z(n5020) );
  XOR \MIXCOLUMNS[6].d/U241  ( .A(n5022), .B(n5021), .Z(\w0[7][54] ) );
  XOR \MIXCOLUMNS[6].d/U240  ( .A(n5184), .B(n5023), .Z(n5021) );
  XOR \MIXCOLUMNS[6].d/U239  ( .A(n345), .B(n5171), .Z(n5022) );
  XOR \MIXCOLUMNS[6].d/U238  ( .A(n829), .B(n346), .Z(n5023) );
  XOR \MIXCOLUMNS[6].d/U237  ( .A(n5186), .B(n5024), .Z(\w0[7][55] ) );
  XOR \MIXCOLUMNS[6].d/U236  ( .A(n827), .B(n5171), .Z(n5024) );
  XOR \MIXCOLUMNS[6].d/U235  ( .A(n5172), .B(n5025), .Z(\w0[7][56] ) );
  XOR \MIXCOLUMNS[6].d/U234  ( .A(n358), .B(n5173), .Z(n5025) );
  XOR \MIXCOLUMNS[6].d/U233  ( .A(n5174), .B(n5026), .Z(\w0[7][57] ) );
  XOR \MIXCOLUMNS[6].d/U232  ( .A(n357), .B(n5175), .Z(n5026) );
  XOR \MIXCOLUMNS[6].d/U231  ( .A(n5176), .B(n5027), .Z(\w0[7][58] ) );
  XOR \MIXCOLUMNS[6].d/U230  ( .A(\w3[6][50] ), .B(n5177), .Z(n5027) );
  XOR \MIXCOLUMNS[6].d/U229  ( .A(n5029), .B(n5028), .Z(\w0[7][59] ) );
  XOR \MIXCOLUMNS[6].d/U228  ( .A(n5179), .B(n5178), .Z(n5028) );
  XOR \MIXCOLUMNS[6].d/U227  ( .A(n354), .B(n5187), .Z(n5029) );
  XOR \MIXCOLUMNS[6].d/U226  ( .A(n5031), .B(n5030), .Z(\w0[7][60] ) );
  XOR \MIXCOLUMNS[6].d/U225  ( .A(n5181), .B(n5180), .Z(n5030) );
  XOR \MIXCOLUMNS[6].d/U224  ( .A(n352), .B(n5187), .Z(n5031) );
  XOR \MIXCOLUMNS[6].d/U223  ( .A(n5182), .B(n5032), .Z(\w0[7][61] ) );
  XOR \MIXCOLUMNS[6].d/U222  ( .A(n350), .B(n5183), .Z(n5032) );
  XOR \MIXCOLUMNS[6].d/U221  ( .A(n5034), .B(n5033), .Z(\w0[7][62] ) );
  XOR \MIXCOLUMNS[6].d/U220  ( .A(n5185), .B(n5184), .Z(n5033) );
  XOR \MIXCOLUMNS[6].d/U219  ( .A(n348), .B(n5187), .Z(n5034) );
  XOR \MIXCOLUMNS[6].d/U218  ( .A(n5186), .B(n5035), .Z(\w0[7][63] ) );
  XOR \MIXCOLUMNS[6].d/U217  ( .A(n346), .B(n5187), .Z(n5035) );
  XOR \MIXCOLUMNS[6].d/U216  ( .A(n826), .B(n344), .Z(n5205) );
  XOR \MIXCOLUMNS[6].d/U215  ( .A(n5037), .B(n5036), .Z(\w0[7][64] ) );
  XOR \MIXCOLUMNS[6].d/U214  ( .A(n825), .B(n5205), .Z(n5036) );
  XOR \MIXCOLUMNS[6].d/U213  ( .A(n824), .B(n22), .Z(n5037) );
  XOR \MIXCOLUMNS[6].d/U212  ( .A(n824), .B(n343), .Z(n5190) );
  XOR \MIXCOLUMNS[6].d/U211  ( .A(n5039), .B(n5038), .Z(\w0[7][65] ) );
  XOR \MIXCOLUMNS[6].d/U210  ( .A(\w3[6][66] ), .B(n5190), .Z(n5038) );
  XOR \MIXCOLUMNS[6].d/U209  ( .A(\w3[6][90] ), .B(n342), .Z(n5039) );
  XOR \MIXCOLUMNS[6].d/U208  ( .A(\w3[6][90] ), .B(\w3[6][82] ), .Z(n5193) );
  XOR \MIXCOLUMNS[6].d/U207  ( .A(n5041), .B(n5040), .Z(\w0[7][66] ) );
  XOR \MIXCOLUMNS[6].d/U206  ( .A(n823), .B(n5193), .Z(n5040) );
  XOR \MIXCOLUMNS[6].d/U205  ( .A(n822), .B(\w3[6][74] ), .Z(n5041) );
  XOR \MIXCOLUMNS[6].d/U204  ( .A(n826), .B(n341), .Z(n5188) );
  XOR \MIXCOLUMNS[6].d/U203  ( .A(n822), .B(n340), .Z(n5195) );
  XOR \MIXCOLUMNS[6].d/U202  ( .A(n5043), .B(n5042), .Z(\w0[7][67] ) );
  XOR \MIXCOLUMNS[6].d/U201  ( .A(n5195), .B(n5044), .Z(n5042) );
  XOR \MIXCOLUMNS[6].d/U200  ( .A(n821), .B(n5188), .Z(n5043) );
  XOR \MIXCOLUMNS[6].d/U199  ( .A(n820), .B(n339), .Z(n5044) );
  XOR \MIXCOLUMNS[6].d/U198  ( .A(n820), .B(n338), .Z(n5197) );
  XOR \MIXCOLUMNS[6].d/U197  ( .A(n5046), .B(n5045), .Z(\w0[7][68] ) );
  XOR \MIXCOLUMNS[6].d/U196  ( .A(n5197), .B(n5047), .Z(n5045) );
  XOR \MIXCOLUMNS[6].d/U195  ( .A(n819), .B(n5188), .Z(n5046) );
  XOR \MIXCOLUMNS[6].d/U194  ( .A(n818), .B(n337), .Z(n5047) );
  XOR \MIXCOLUMNS[6].d/U193  ( .A(n818), .B(n336), .Z(n5199) );
  XOR \MIXCOLUMNS[6].d/U192  ( .A(n5049), .B(n5048), .Z(\w0[7][69] ) );
  XOR \MIXCOLUMNS[6].d/U191  ( .A(n817), .B(n5199), .Z(n5048) );
  XOR \MIXCOLUMNS[6].d/U190  ( .A(n816), .B(n335), .Z(n5049) );
  XOR \MIXCOLUMNS[6].d/U189  ( .A(n816), .B(n334), .Z(n5201) );
  XOR \MIXCOLUMNS[6].d/U188  ( .A(n5051), .B(n5050), .Z(\w0[7][70] ) );
  XOR \MIXCOLUMNS[6].d/U187  ( .A(n5201), .B(n5052), .Z(n5050) );
  XOR \MIXCOLUMNS[6].d/U186  ( .A(n815), .B(n5188), .Z(n5051) );
  XOR \MIXCOLUMNS[6].d/U185  ( .A(n814), .B(n333), .Z(n5052) );
  XOR \MIXCOLUMNS[6].d/U184  ( .A(n814), .B(n332), .Z(n5203) );
  XOR \MIXCOLUMNS[6].d/U183  ( .A(n5203), .B(n5053), .Z(\w0[7][71] ) );
  XOR \MIXCOLUMNS[6].d/U182  ( .A(n331), .B(n5188), .Z(n5053) );
  XOR \MIXCOLUMNS[6].d/U181  ( .A(n342), .B(n825), .Z(n5192) );
  XOR \MIXCOLUMNS[6].d/U180  ( .A(n5192), .B(n5054), .Z(\w0[7][72] ) );
  XOR \MIXCOLUMNS[6].d/U179  ( .A(n341), .B(n5205), .Z(n5054) );
  XOR \MIXCOLUMNS[6].d/U178  ( .A(\w3[6][74] ), .B(\w3[6][66] ), .Z(n5194) );
  XOR \MIXCOLUMNS[6].d/U177  ( .A(n5194), .B(n5055), .Z(\w0[7][73] ) );
  XOR \MIXCOLUMNS[6].d/U176  ( .A(n825), .B(n5190), .Z(n5055) );
  XOR \MIXCOLUMNS[6].d/U175  ( .A(n339), .B(n823), .Z(n5196) );
  XOR \MIXCOLUMNS[6].d/U174  ( .A(n5196), .B(n5056), .Z(\w0[7][74] ) );
  XOR \MIXCOLUMNS[6].d/U173  ( .A(\w3[6][66] ), .B(n5193), .Z(n5056) );
  XOR \MIXCOLUMNS[6].d/U172  ( .A(n22), .B(n341), .Z(n5191) );
  XOR \MIXCOLUMNS[6].d/U171  ( .A(n337), .B(n821), .Z(n5198) );
  XOR \MIXCOLUMNS[6].d/U170  ( .A(n5058), .B(n5057), .Z(\w0[7][75] ) );
  XOR \MIXCOLUMNS[6].d/U169  ( .A(n5195), .B(n5198), .Z(n5057) );
  XOR \MIXCOLUMNS[6].d/U168  ( .A(n823), .B(n5191), .Z(n5058) );
  XOR \MIXCOLUMNS[6].d/U167  ( .A(n335), .B(n819), .Z(n5200) );
  XOR \MIXCOLUMNS[6].d/U166  ( .A(n5060), .B(n5059), .Z(\w0[7][76] ) );
  XOR \MIXCOLUMNS[6].d/U165  ( .A(n5197), .B(n5200), .Z(n5059) );
  XOR \MIXCOLUMNS[6].d/U164  ( .A(n821), .B(n5191), .Z(n5060) );
  XOR \MIXCOLUMNS[6].d/U163  ( .A(n333), .B(n817), .Z(n5202) );
  XOR \MIXCOLUMNS[6].d/U162  ( .A(n5202), .B(n5061), .Z(\w0[7][77] ) );
  XOR \MIXCOLUMNS[6].d/U161  ( .A(n819), .B(n5199), .Z(n5061) );
  XOR \MIXCOLUMNS[6].d/U160  ( .A(n331), .B(n815), .Z(n5204) );
  XOR \MIXCOLUMNS[6].d/U159  ( .A(n5063), .B(n5062), .Z(\w0[7][78] ) );
  XOR \MIXCOLUMNS[6].d/U158  ( .A(n5201), .B(n5204), .Z(n5062) );
  XOR \MIXCOLUMNS[6].d/U157  ( .A(n817), .B(n5191), .Z(n5063) );
  XOR \MIXCOLUMNS[6].d/U156  ( .A(n5203), .B(n5064), .Z(\w0[7][79] ) );
  XOR \MIXCOLUMNS[6].d/U155  ( .A(n815), .B(n5191), .Z(n5064) );
  XOR \MIXCOLUMNS[6].d/U154  ( .A(n5066), .B(n5065), .Z(\w0[7][80] ) );
  XOR \MIXCOLUMNS[6].d/U153  ( .A(n342), .B(n5191), .Z(n5065) );
  XOR \MIXCOLUMNS[6].d/U152  ( .A(n826), .B(n343), .Z(n5066) );
  XOR \MIXCOLUMNS[6].d/U151  ( .A(n5068), .B(n5067), .Z(\w0[7][81] ) );
  XOR \MIXCOLUMNS[6].d/U150  ( .A(\w3[6][74] ), .B(n5192), .Z(n5067) );
  XOR \MIXCOLUMNS[6].d/U149  ( .A(n824), .B(\w3[6][82] ), .Z(n5068) );
  XOR \MIXCOLUMNS[6].d/U148  ( .A(n5070), .B(n5069), .Z(\w0[7][82] ) );
  XOR \MIXCOLUMNS[6].d/U147  ( .A(n339), .B(n5194), .Z(n5069) );
  XOR \MIXCOLUMNS[6].d/U146  ( .A(\w3[6][90] ), .B(n340), .Z(n5070) );
  XOR \MIXCOLUMNS[6].d/U145  ( .A(n344), .B(n22), .Z(n5189) );
  XOR \MIXCOLUMNS[6].d/U144  ( .A(n5072), .B(n5071), .Z(\w0[7][83] ) );
  XOR \MIXCOLUMNS[6].d/U143  ( .A(n5196), .B(n5073), .Z(n5071) );
  XOR \MIXCOLUMNS[6].d/U142  ( .A(n337), .B(n5189), .Z(n5072) );
  XOR \MIXCOLUMNS[6].d/U141  ( .A(n822), .B(n338), .Z(n5073) );
  XOR \MIXCOLUMNS[6].d/U140  ( .A(n5075), .B(n5074), .Z(\w0[7][84] ) );
  XOR \MIXCOLUMNS[6].d/U139  ( .A(n5198), .B(n5076), .Z(n5074) );
  XOR \MIXCOLUMNS[6].d/U138  ( .A(n335), .B(n5189), .Z(n5075) );
  XOR \MIXCOLUMNS[6].d/U137  ( .A(n820), .B(n336), .Z(n5076) );
  XOR \MIXCOLUMNS[6].d/U136  ( .A(n5078), .B(n5077), .Z(\w0[7][85] ) );
  XOR \MIXCOLUMNS[6].d/U135  ( .A(n333), .B(n5200), .Z(n5077) );
  XOR \MIXCOLUMNS[6].d/U134  ( .A(n818), .B(n334), .Z(n5078) );
  XOR \MIXCOLUMNS[6].d/U133  ( .A(n5080), .B(n5079), .Z(\w0[7][86] ) );
  XOR \MIXCOLUMNS[6].d/U132  ( .A(n5202), .B(n5081), .Z(n5079) );
  XOR \MIXCOLUMNS[6].d/U131  ( .A(n331), .B(n5189), .Z(n5080) );
  XOR \MIXCOLUMNS[6].d/U130  ( .A(n816), .B(n332), .Z(n5081) );
  XOR \MIXCOLUMNS[6].d/U129  ( .A(n5204), .B(n5082), .Z(\w0[7][87] ) );
  XOR \MIXCOLUMNS[6].d/U128  ( .A(n814), .B(n5189), .Z(n5082) );
  XOR \MIXCOLUMNS[6].d/U127  ( .A(n5190), .B(n5083), .Z(\w0[7][88] ) );
  XOR \MIXCOLUMNS[6].d/U126  ( .A(n344), .B(n5191), .Z(n5083) );
  XOR \MIXCOLUMNS[6].d/U125  ( .A(n5192), .B(n5084), .Z(\w0[7][89] ) );
  XOR \MIXCOLUMNS[6].d/U124  ( .A(n343), .B(n5193), .Z(n5084) );
  XOR \MIXCOLUMNS[6].d/U123  ( .A(n5194), .B(n5085), .Z(\w0[7][90] ) );
  XOR \MIXCOLUMNS[6].d/U122  ( .A(\w3[6][82] ), .B(n5195), .Z(n5085) );
  XOR \MIXCOLUMNS[6].d/U121  ( .A(n5087), .B(n5086), .Z(\w0[7][91] ) );
  XOR \MIXCOLUMNS[6].d/U120  ( .A(n5197), .B(n5196), .Z(n5086) );
  XOR \MIXCOLUMNS[6].d/U119  ( .A(n340), .B(n5205), .Z(n5087) );
  XOR \MIXCOLUMNS[6].d/U118  ( .A(n5089), .B(n5088), .Z(\w0[7][92] ) );
  XOR \MIXCOLUMNS[6].d/U117  ( .A(n5199), .B(n5198), .Z(n5088) );
  XOR \MIXCOLUMNS[6].d/U116  ( .A(n338), .B(n5205), .Z(n5089) );
  XOR \MIXCOLUMNS[6].d/U115  ( .A(n5200), .B(n5090), .Z(\w0[7][93] ) );
  XOR \MIXCOLUMNS[6].d/U114  ( .A(n336), .B(n5201), .Z(n5090) );
  XOR \MIXCOLUMNS[6].d/U113  ( .A(n5092), .B(n5091), .Z(\w0[7][94] ) );
  XOR \MIXCOLUMNS[6].d/U112  ( .A(n5203), .B(n5202), .Z(n5091) );
  XOR \MIXCOLUMNS[6].d/U111  ( .A(n334), .B(n5205), .Z(n5092) );
  XOR \MIXCOLUMNS[6].d/U110  ( .A(n5204), .B(n5093), .Z(\w0[7][95] ) );
  XOR \MIXCOLUMNS[6].d/U109  ( .A(n332), .B(n5205), .Z(n5093) );
  XOR \MIXCOLUMNS[6].d/U108  ( .A(n813), .B(n330), .Z(n5223) );
  XOR \MIXCOLUMNS[6].d/U107  ( .A(n5095), .B(n5094), .Z(\w0[7][96] ) );
  XOR \MIXCOLUMNS[6].d/U106  ( .A(n812), .B(n5223), .Z(n5094) );
  XOR \MIXCOLUMNS[6].d/U105  ( .A(n811), .B(n21), .Z(n5095) );
  XOR \MIXCOLUMNS[6].d/U104  ( .A(n811), .B(n329), .Z(n5208) );
  XOR \MIXCOLUMNS[6].d/U103  ( .A(n5097), .B(n5096), .Z(\w0[7][97] ) );
  XOR \MIXCOLUMNS[6].d/U102  ( .A(\w3[6][98] ), .B(n5208), .Z(n5096) );
  XOR \MIXCOLUMNS[6].d/U101  ( .A(\w3[6][122] ), .B(n328), .Z(n5097) );
  XOR \MIXCOLUMNS[6].d/U100  ( .A(\w3[6][122] ), .B(\w3[6][114] ), .Z(n5211)
         );
  XOR \MIXCOLUMNS[6].d/U99  ( .A(n5099), .B(n5098), .Z(\w0[7][98] ) );
  XOR \MIXCOLUMNS[6].d/U98  ( .A(n810), .B(n5211), .Z(n5098) );
  XOR \MIXCOLUMNS[6].d/U97  ( .A(n809), .B(\w3[6][106] ), .Z(n5099) );
  XOR \MIXCOLUMNS[6].d/U96  ( .A(n813), .B(n327), .Z(n5206) );
  XOR \MIXCOLUMNS[6].d/U95  ( .A(n809), .B(n326), .Z(n5213) );
  XOR \MIXCOLUMNS[6].d/U94  ( .A(n5101), .B(n5100), .Z(\w0[7][99] ) );
  XOR \MIXCOLUMNS[6].d/U93  ( .A(n5213), .B(n5102), .Z(n5100) );
  XOR \MIXCOLUMNS[6].d/U92  ( .A(n808), .B(n5206), .Z(n5101) );
  XOR \MIXCOLUMNS[6].d/U91  ( .A(n807), .B(n325), .Z(n5102) );
  XOR \MIXCOLUMNS[6].d/U90  ( .A(n807), .B(n324), .Z(n5215) );
  XOR \MIXCOLUMNS[6].d/U89  ( .A(n5104), .B(n5103), .Z(\w0[7][100] ) );
  XOR \MIXCOLUMNS[6].d/U88  ( .A(n5215), .B(n5105), .Z(n5103) );
  XOR \MIXCOLUMNS[6].d/U87  ( .A(n806), .B(n5206), .Z(n5104) );
  XOR \MIXCOLUMNS[6].d/U86  ( .A(n805), .B(n323), .Z(n5105) );
  XOR \MIXCOLUMNS[6].d/U85  ( .A(n805), .B(n322), .Z(n5217) );
  XOR \MIXCOLUMNS[6].d/U84  ( .A(n5107), .B(n5106), .Z(\w0[7][101] ) );
  XOR \MIXCOLUMNS[6].d/U83  ( .A(n804), .B(n5217), .Z(n5106) );
  XOR \MIXCOLUMNS[6].d/U82  ( .A(n803), .B(n321), .Z(n5107) );
  XOR \MIXCOLUMNS[6].d/U81  ( .A(n803), .B(n320), .Z(n5219) );
  XOR \MIXCOLUMNS[6].d/U80  ( .A(n5109), .B(n5108), .Z(\w0[7][102] ) );
  XOR \MIXCOLUMNS[6].d/U79  ( .A(n5219), .B(n5110), .Z(n5108) );
  XOR \MIXCOLUMNS[6].d/U78  ( .A(n802), .B(n5206), .Z(n5109) );
  XOR \MIXCOLUMNS[6].d/U77  ( .A(n801), .B(n319), .Z(n5110) );
  XOR \MIXCOLUMNS[6].d/U76  ( .A(n801), .B(n318), .Z(n5221) );
  XOR \MIXCOLUMNS[6].d/U75  ( .A(n5221), .B(n5111), .Z(\w0[7][103] ) );
  XOR \MIXCOLUMNS[6].d/U74  ( .A(n317), .B(n5206), .Z(n5111) );
  XOR \MIXCOLUMNS[6].d/U73  ( .A(n328), .B(n812), .Z(n5210) );
  XOR \MIXCOLUMNS[6].d/U72  ( .A(n5210), .B(n5112), .Z(\w0[7][104] ) );
  XOR \MIXCOLUMNS[6].d/U71  ( .A(n327), .B(n5223), .Z(n5112) );
  XOR \MIXCOLUMNS[6].d/U70  ( .A(\w3[6][106] ), .B(\w3[6][98] ), .Z(n5212) );
  XOR \MIXCOLUMNS[6].d/U69  ( .A(n5212), .B(n5113), .Z(\w0[7][105] ) );
  XOR \MIXCOLUMNS[6].d/U68  ( .A(n812), .B(n5208), .Z(n5113) );
  XOR \MIXCOLUMNS[6].d/U67  ( .A(n325), .B(n810), .Z(n5214) );
  XOR \MIXCOLUMNS[6].d/U66  ( .A(n5214), .B(n5114), .Z(\w0[7][106] ) );
  XOR \MIXCOLUMNS[6].d/U65  ( .A(\w3[6][98] ), .B(n5211), .Z(n5114) );
  XOR \MIXCOLUMNS[6].d/U64  ( .A(n21), .B(n327), .Z(n5209) );
  XOR \MIXCOLUMNS[6].d/U63  ( .A(n323), .B(n808), .Z(n5216) );
  XOR \MIXCOLUMNS[6].d/U62  ( .A(n5116), .B(n5115), .Z(\w0[7][107] ) );
  XOR \MIXCOLUMNS[6].d/U61  ( .A(n5213), .B(n5216), .Z(n5115) );
  XOR \MIXCOLUMNS[6].d/U60  ( .A(n810), .B(n5209), .Z(n5116) );
  XOR \MIXCOLUMNS[6].d/U59  ( .A(n321), .B(n806), .Z(n5218) );
  XOR \MIXCOLUMNS[6].d/U58  ( .A(n5118), .B(n5117), .Z(\w0[7][108] ) );
  XOR \MIXCOLUMNS[6].d/U57  ( .A(n5215), .B(n5218), .Z(n5117) );
  XOR \MIXCOLUMNS[6].d/U56  ( .A(n808), .B(n5209), .Z(n5118) );
  XOR \MIXCOLUMNS[6].d/U55  ( .A(n319), .B(n804), .Z(n5220) );
  XOR \MIXCOLUMNS[6].d/U54  ( .A(n5220), .B(n5119), .Z(\w0[7][109] ) );
  XOR \MIXCOLUMNS[6].d/U53  ( .A(n806), .B(n5217), .Z(n5119) );
  XOR \MIXCOLUMNS[6].d/U52  ( .A(n317), .B(n802), .Z(n5222) );
  XOR \MIXCOLUMNS[6].d/U51  ( .A(n5121), .B(n5120), .Z(\w0[7][110] ) );
  XOR \MIXCOLUMNS[6].d/U50  ( .A(n5219), .B(n5222), .Z(n5120) );
  XOR \MIXCOLUMNS[6].d/U49  ( .A(n804), .B(n5209), .Z(n5121) );
  XOR \MIXCOLUMNS[6].d/U48  ( .A(n5221), .B(n5122), .Z(\w0[7][111] ) );
  XOR \MIXCOLUMNS[6].d/U47  ( .A(n802), .B(n5209), .Z(n5122) );
  XOR \MIXCOLUMNS[6].d/U46  ( .A(n5124), .B(n5123), .Z(\w0[7][112] ) );
  XOR \MIXCOLUMNS[6].d/U45  ( .A(n328), .B(n5209), .Z(n5123) );
  XOR \MIXCOLUMNS[6].d/U44  ( .A(n813), .B(n329), .Z(n5124) );
  XOR \MIXCOLUMNS[6].d/U43  ( .A(n5126), .B(n5125), .Z(\w0[7][113] ) );
  XOR \MIXCOLUMNS[6].d/U42  ( .A(\w3[6][106] ), .B(n5210), .Z(n5125) );
  XOR \MIXCOLUMNS[6].d/U41  ( .A(n811), .B(\w3[6][114] ), .Z(n5126) );
  XOR \MIXCOLUMNS[6].d/U40  ( .A(n5128), .B(n5127), .Z(\w0[7][114] ) );
  XOR \MIXCOLUMNS[6].d/U39  ( .A(n325), .B(n5212), .Z(n5127) );
  XOR \MIXCOLUMNS[6].d/U38  ( .A(\w3[6][122] ), .B(n326), .Z(n5128) );
  XOR \MIXCOLUMNS[6].d/U37  ( .A(n330), .B(n21), .Z(n5207) );
  XOR \MIXCOLUMNS[6].d/U36  ( .A(n5130), .B(n5129), .Z(\w0[7][115] ) );
  XOR \MIXCOLUMNS[6].d/U35  ( .A(n5214), .B(n5131), .Z(n5129) );
  XOR \MIXCOLUMNS[6].d/U34  ( .A(n323), .B(n5207), .Z(n5130) );
  XOR \MIXCOLUMNS[6].d/U33  ( .A(n809), .B(n324), .Z(n5131) );
  XOR \MIXCOLUMNS[6].d/U32  ( .A(n5133), .B(n5132), .Z(\w0[7][116] ) );
  XOR \MIXCOLUMNS[6].d/U31  ( .A(n5216), .B(n5134), .Z(n5132) );
  XOR \MIXCOLUMNS[6].d/U30  ( .A(n321), .B(n5207), .Z(n5133) );
  XOR \MIXCOLUMNS[6].d/U29  ( .A(n807), .B(n322), .Z(n5134) );
  XOR \MIXCOLUMNS[6].d/U28  ( .A(n5136), .B(n5135), .Z(\w0[7][117] ) );
  XOR \MIXCOLUMNS[6].d/U27  ( .A(n319), .B(n5218), .Z(n5135) );
  XOR \MIXCOLUMNS[6].d/U26  ( .A(n805), .B(n320), .Z(n5136) );
  XOR \MIXCOLUMNS[6].d/U25  ( .A(n5138), .B(n5137), .Z(\w0[7][118] ) );
  XOR \MIXCOLUMNS[6].d/U24  ( .A(n5220), .B(n5139), .Z(n5137) );
  XOR \MIXCOLUMNS[6].d/U23  ( .A(n317), .B(n5207), .Z(n5138) );
  XOR \MIXCOLUMNS[6].d/U22  ( .A(n803), .B(n318), .Z(n5139) );
  XOR \MIXCOLUMNS[6].d/U21  ( .A(n5222), .B(n5140), .Z(\w0[7][119] ) );
  XOR \MIXCOLUMNS[6].d/U20  ( .A(n801), .B(n5207), .Z(n5140) );
  XOR \MIXCOLUMNS[6].d/U19  ( .A(n5208), .B(n5141), .Z(\w0[7][120] ) );
  XOR \MIXCOLUMNS[6].d/U18  ( .A(n330), .B(n5209), .Z(n5141) );
  XOR \MIXCOLUMNS[6].d/U17  ( .A(n5210), .B(n5142), .Z(\w0[7][121] ) );
  XOR \MIXCOLUMNS[6].d/U16  ( .A(n329), .B(n5211), .Z(n5142) );
  XOR \MIXCOLUMNS[6].d/U15  ( .A(n5212), .B(n5143), .Z(\w0[7][122] ) );
  XOR \MIXCOLUMNS[6].d/U14  ( .A(\w3[6][114] ), .B(n5213), .Z(n5143) );
  XOR \MIXCOLUMNS[6].d/U13  ( .A(n5145), .B(n5144), .Z(\w0[7][123] ) );
  XOR \MIXCOLUMNS[6].d/U12  ( .A(n5215), .B(n5214), .Z(n5144) );
  XOR \MIXCOLUMNS[6].d/U11  ( .A(n326), .B(n5223), .Z(n5145) );
  XOR \MIXCOLUMNS[6].d/U10  ( .A(n5147), .B(n5146), .Z(\w0[7][124] ) );
  XOR \MIXCOLUMNS[6].d/U9  ( .A(n5217), .B(n5216), .Z(n5146) );
  XOR \MIXCOLUMNS[6].d/U8  ( .A(n324), .B(n5223), .Z(n5147) );
  XOR \MIXCOLUMNS[6].d/U7  ( .A(n5218), .B(n5148), .Z(\w0[7][125] ) );
  XOR \MIXCOLUMNS[6].d/U6  ( .A(n322), .B(n5219), .Z(n5148) );
  XOR \MIXCOLUMNS[6].d/U5  ( .A(n5150), .B(n5149), .Z(\w0[7][126] ) );
  XOR \MIXCOLUMNS[6].d/U4  ( .A(n5221), .B(n5220), .Z(n5149) );
  XOR \MIXCOLUMNS[6].d/U3  ( .A(n320), .B(n5223), .Z(n5150) );
  XOR \MIXCOLUMNS[6].d/U2  ( .A(n5222), .B(n5151), .Z(\w0[7][127] ) );
  XOR \MIXCOLUMNS[6].d/U1  ( .A(n318), .B(n5223), .Z(n5151) );
  XOR \MIXCOLUMNS[5].d/U432  ( .A(n800), .B(n316), .Z(n4865) );
  XOR \MIXCOLUMNS[5].d/U431  ( .A(n4617), .B(n4616), .Z(\w0[6][0] ) );
  XOR \MIXCOLUMNS[5].d/U430  ( .A(n799), .B(n4865), .Z(n4616) );
  XOR \MIXCOLUMNS[5].d/U429  ( .A(n798), .B(n20), .Z(n4617) );
  XOR \MIXCOLUMNS[5].d/U428  ( .A(n798), .B(n315), .Z(n4850) );
  XOR \MIXCOLUMNS[5].d/U427  ( .A(n4619), .B(n4618), .Z(\w0[6][1] ) );
  XOR \MIXCOLUMNS[5].d/U426  ( .A(\w3[5][2] ), .B(n4850), .Z(n4618) );
  XOR \MIXCOLUMNS[5].d/U425  ( .A(\w3[5][26] ), .B(n314), .Z(n4619) );
  XOR \MIXCOLUMNS[5].d/U424  ( .A(\w3[5][26] ), .B(\w3[5][18] ), .Z(n4853) );
  XOR \MIXCOLUMNS[5].d/U423  ( .A(n4621), .B(n4620), .Z(\w0[6][2] ) );
  XOR \MIXCOLUMNS[5].d/U422  ( .A(n797), .B(n4853), .Z(n4620) );
  XOR \MIXCOLUMNS[5].d/U421  ( .A(n796), .B(\w3[5][10] ), .Z(n4621) );
  XOR \MIXCOLUMNS[5].d/U420  ( .A(n800), .B(n313), .Z(n4848) );
  XOR \MIXCOLUMNS[5].d/U419  ( .A(n796), .B(n312), .Z(n4855) );
  XOR \MIXCOLUMNS[5].d/U418  ( .A(n4623), .B(n4622), .Z(\w0[6][3] ) );
  XOR \MIXCOLUMNS[5].d/U417  ( .A(n4855), .B(n4624), .Z(n4622) );
  XOR \MIXCOLUMNS[5].d/U416  ( .A(n795), .B(n4848), .Z(n4623) );
  XOR \MIXCOLUMNS[5].d/U415  ( .A(n794), .B(n311), .Z(n4624) );
  XOR \MIXCOLUMNS[5].d/U414  ( .A(n794), .B(n310), .Z(n4857) );
  XOR \MIXCOLUMNS[5].d/U413  ( .A(n4626), .B(n4625), .Z(\w0[6][4] ) );
  XOR \MIXCOLUMNS[5].d/U412  ( .A(n4857), .B(n4627), .Z(n4625) );
  XOR \MIXCOLUMNS[5].d/U411  ( .A(n793), .B(n4848), .Z(n4626) );
  XOR \MIXCOLUMNS[5].d/U410  ( .A(n792), .B(n309), .Z(n4627) );
  XOR \MIXCOLUMNS[5].d/U409  ( .A(n792), .B(n308), .Z(n4859) );
  XOR \MIXCOLUMNS[5].d/U408  ( .A(n4629), .B(n4628), .Z(\w0[6][5] ) );
  XOR \MIXCOLUMNS[5].d/U407  ( .A(n791), .B(n4859), .Z(n4628) );
  XOR \MIXCOLUMNS[5].d/U406  ( .A(n790), .B(n307), .Z(n4629) );
  XOR \MIXCOLUMNS[5].d/U405  ( .A(n790), .B(n306), .Z(n4861) );
  XOR \MIXCOLUMNS[5].d/U404  ( .A(n4631), .B(n4630), .Z(\w0[6][6] ) );
  XOR \MIXCOLUMNS[5].d/U403  ( .A(n4861), .B(n4632), .Z(n4630) );
  XOR \MIXCOLUMNS[5].d/U402  ( .A(n789), .B(n4848), .Z(n4631) );
  XOR \MIXCOLUMNS[5].d/U401  ( .A(n788), .B(n305), .Z(n4632) );
  XOR \MIXCOLUMNS[5].d/U400  ( .A(n788), .B(n304), .Z(n4863) );
  XOR \MIXCOLUMNS[5].d/U399  ( .A(n4863), .B(n4633), .Z(\w0[6][7] ) );
  XOR \MIXCOLUMNS[5].d/U398  ( .A(n303), .B(n4848), .Z(n4633) );
  XOR \MIXCOLUMNS[5].d/U397  ( .A(n314), .B(n799), .Z(n4852) );
  XOR \MIXCOLUMNS[5].d/U396  ( .A(n4852), .B(n4634), .Z(\w0[6][8] ) );
  XOR \MIXCOLUMNS[5].d/U395  ( .A(n313), .B(n4865), .Z(n4634) );
  XOR \MIXCOLUMNS[5].d/U394  ( .A(\w3[5][10] ), .B(\w3[5][2] ), .Z(n4854) );
  XOR \MIXCOLUMNS[5].d/U393  ( .A(n4854), .B(n4635), .Z(\w0[6][9] ) );
  XOR \MIXCOLUMNS[5].d/U392  ( .A(n799), .B(n4850), .Z(n4635) );
  XOR \MIXCOLUMNS[5].d/U391  ( .A(n311), .B(n797), .Z(n4856) );
  XOR \MIXCOLUMNS[5].d/U390  ( .A(n4856), .B(n4636), .Z(\w0[6][10] ) );
  XOR \MIXCOLUMNS[5].d/U389  ( .A(\w3[5][2] ), .B(n4853), .Z(n4636) );
  XOR \MIXCOLUMNS[5].d/U388  ( .A(n20), .B(n313), .Z(n4851) );
  XOR \MIXCOLUMNS[5].d/U387  ( .A(n309), .B(n795), .Z(n4858) );
  XOR \MIXCOLUMNS[5].d/U386  ( .A(n4638), .B(n4637), .Z(\w0[6][11] ) );
  XOR \MIXCOLUMNS[5].d/U385  ( .A(n4855), .B(n4858), .Z(n4637) );
  XOR \MIXCOLUMNS[5].d/U384  ( .A(n797), .B(n4851), .Z(n4638) );
  XOR \MIXCOLUMNS[5].d/U383  ( .A(n307), .B(n793), .Z(n4860) );
  XOR \MIXCOLUMNS[5].d/U382  ( .A(n4640), .B(n4639), .Z(\w0[6][12] ) );
  XOR \MIXCOLUMNS[5].d/U381  ( .A(n4857), .B(n4860), .Z(n4639) );
  XOR \MIXCOLUMNS[5].d/U380  ( .A(n795), .B(n4851), .Z(n4640) );
  XOR \MIXCOLUMNS[5].d/U379  ( .A(n305), .B(n791), .Z(n4862) );
  XOR \MIXCOLUMNS[5].d/U378  ( .A(n4862), .B(n4641), .Z(\w0[6][13] ) );
  XOR \MIXCOLUMNS[5].d/U377  ( .A(n793), .B(n4859), .Z(n4641) );
  XOR \MIXCOLUMNS[5].d/U376  ( .A(n303), .B(n789), .Z(n4864) );
  XOR \MIXCOLUMNS[5].d/U375  ( .A(n4643), .B(n4642), .Z(\w0[6][14] ) );
  XOR \MIXCOLUMNS[5].d/U374  ( .A(n4861), .B(n4864), .Z(n4642) );
  XOR \MIXCOLUMNS[5].d/U373  ( .A(n791), .B(n4851), .Z(n4643) );
  XOR \MIXCOLUMNS[5].d/U372  ( .A(n4863), .B(n4644), .Z(\w0[6][15] ) );
  XOR \MIXCOLUMNS[5].d/U371  ( .A(n789), .B(n4851), .Z(n4644) );
  XOR \MIXCOLUMNS[5].d/U370  ( .A(n4646), .B(n4645), .Z(\w0[6][16] ) );
  XOR \MIXCOLUMNS[5].d/U369  ( .A(n314), .B(n4851), .Z(n4645) );
  XOR \MIXCOLUMNS[5].d/U368  ( .A(n800), .B(n315), .Z(n4646) );
  XOR \MIXCOLUMNS[5].d/U367  ( .A(n4648), .B(n4647), .Z(\w0[6][17] ) );
  XOR \MIXCOLUMNS[5].d/U366  ( .A(\w3[5][10] ), .B(n4852), .Z(n4647) );
  XOR \MIXCOLUMNS[5].d/U365  ( .A(n798), .B(\w3[5][18] ), .Z(n4648) );
  XOR \MIXCOLUMNS[5].d/U364  ( .A(n4650), .B(n4649), .Z(\w0[6][18] ) );
  XOR \MIXCOLUMNS[5].d/U363  ( .A(n311), .B(n4854), .Z(n4649) );
  XOR \MIXCOLUMNS[5].d/U362  ( .A(\w3[5][26] ), .B(n312), .Z(n4650) );
  XOR \MIXCOLUMNS[5].d/U361  ( .A(n316), .B(n20), .Z(n4849) );
  XOR \MIXCOLUMNS[5].d/U360  ( .A(n4652), .B(n4651), .Z(\w0[6][19] ) );
  XOR \MIXCOLUMNS[5].d/U359  ( .A(n4856), .B(n4653), .Z(n4651) );
  XOR \MIXCOLUMNS[5].d/U358  ( .A(n309), .B(n4849), .Z(n4652) );
  XOR \MIXCOLUMNS[5].d/U357  ( .A(n796), .B(n310), .Z(n4653) );
  XOR \MIXCOLUMNS[5].d/U356  ( .A(n4655), .B(n4654), .Z(\w0[6][20] ) );
  XOR \MIXCOLUMNS[5].d/U355  ( .A(n4858), .B(n4656), .Z(n4654) );
  XOR \MIXCOLUMNS[5].d/U354  ( .A(n307), .B(n4849), .Z(n4655) );
  XOR \MIXCOLUMNS[5].d/U353  ( .A(n794), .B(n308), .Z(n4656) );
  XOR \MIXCOLUMNS[5].d/U352  ( .A(n4658), .B(n4657), .Z(\w0[6][21] ) );
  XOR \MIXCOLUMNS[5].d/U351  ( .A(n305), .B(n4860), .Z(n4657) );
  XOR \MIXCOLUMNS[5].d/U350  ( .A(n792), .B(n306), .Z(n4658) );
  XOR \MIXCOLUMNS[5].d/U349  ( .A(n4660), .B(n4659), .Z(\w0[6][22] ) );
  XOR \MIXCOLUMNS[5].d/U348  ( .A(n4862), .B(n4661), .Z(n4659) );
  XOR \MIXCOLUMNS[5].d/U347  ( .A(n303), .B(n4849), .Z(n4660) );
  XOR \MIXCOLUMNS[5].d/U346  ( .A(n790), .B(n304), .Z(n4661) );
  XOR \MIXCOLUMNS[5].d/U345  ( .A(n4864), .B(n4662), .Z(\w0[6][23] ) );
  XOR \MIXCOLUMNS[5].d/U344  ( .A(n788), .B(n4849), .Z(n4662) );
  XOR \MIXCOLUMNS[5].d/U343  ( .A(n4850), .B(n4663), .Z(\w0[6][24] ) );
  XOR \MIXCOLUMNS[5].d/U342  ( .A(n316), .B(n4851), .Z(n4663) );
  XOR \MIXCOLUMNS[5].d/U341  ( .A(n4852), .B(n4664), .Z(\w0[6][25] ) );
  XOR \MIXCOLUMNS[5].d/U340  ( .A(n315), .B(n4853), .Z(n4664) );
  XOR \MIXCOLUMNS[5].d/U339  ( .A(n4854), .B(n4665), .Z(\w0[6][26] ) );
  XOR \MIXCOLUMNS[5].d/U338  ( .A(\w3[5][18] ), .B(n4855), .Z(n4665) );
  XOR \MIXCOLUMNS[5].d/U337  ( .A(n4667), .B(n4666), .Z(\w0[6][27] ) );
  XOR \MIXCOLUMNS[5].d/U336  ( .A(n4857), .B(n4856), .Z(n4666) );
  XOR \MIXCOLUMNS[5].d/U335  ( .A(n312), .B(n4865), .Z(n4667) );
  XOR \MIXCOLUMNS[5].d/U334  ( .A(n4669), .B(n4668), .Z(\w0[6][28] ) );
  XOR \MIXCOLUMNS[5].d/U333  ( .A(n4859), .B(n4858), .Z(n4668) );
  XOR \MIXCOLUMNS[5].d/U332  ( .A(n310), .B(n4865), .Z(n4669) );
  XOR \MIXCOLUMNS[5].d/U331  ( .A(n4860), .B(n4670), .Z(\w0[6][29] ) );
  XOR \MIXCOLUMNS[5].d/U330  ( .A(n308), .B(n4861), .Z(n4670) );
  XOR \MIXCOLUMNS[5].d/U329  ( .A(n4672), .B(n4671), .Z(\w0[6][30] ) );
  XOR \MIXCOLUMNS[5].d/U328  ( .A(n4863), .B(n4862), .Z(n4671) );
  XOR \MIXCOLUMNS[5].d/U327  ( .A(n306), .B(n4865), .Z(n4672) );
  XOR \MIXCOLUMNS[5].d/U326  ( .A(n4864), .B(n4673), .Z(\w0[6][31] ) );
  XOR \MIXCOLUMNS[5].d/U325  ( .A(n304), .B(n4865), .Z(n4673) );
  XOR \MIXCOLUMNS[5].d/U324  ( .A(n787), .B(n302), .Z(n4883) );
  XOR \MIXCOLUMNS[5].d/U323  ( .A(n4675), .B(n4674), .Z(\w0[6][32] ) );
  XOR \MIXCOLUMNS[5].d/U322  ( .A(n786), .B(n4883), .Z(n4674) );
  XOR \MIXCOLUMNS[5].d/U321  ( .A(n785), .B(n19), .Z(n4675) );
  XOR \MIXCOLUMNS[5].d/U320  ( .A(n785), .B(n301), .Z(n4868) );
  XOR \MIXCOLUMNS[5].d/U319  ( .A(n4677), .B(n4676), .Z(\w0[6][33] ) );
  XOR \MIXCOLUMNS[5].d/U318  ( .A(\w3[5][34] ), .B(n4868), .Z(n4676) );
  XOR \MIXCOLUMNS[5].d/U317  ( .A(\w3[5][58] ), .B(n300), .Z(n4677) );
  XOR \MIXCOLUMNS[5].d/U316  ( .A(\w3[5][58] ), .B(\w3[5][50] ), .Z(n4871) );
  XOR \MIXCOLUMNS[5].d/U315  ( .A(n4679), .B(n4678), .Z(\w0[6][34] ) );
  XOR \MIXCOLUMNS[5].d/U314  ( .A(n784), .B(n4871), .Z(n4678) );
  XOR \MIXCOLUMNS[5].d/U313  ( .A(n783), .B(\w3[5][42] ), .Z(n4679) );
  XOR \MIXCOLUMNS[5].d/U312  ( .A(n787), .B(n299), .Z(n4866) );
  XOR \MIXCOLUMNS[5].d/U311  ( .A(n783), .B(n298), .Z(n4873) );
  XOR \MIXCOLUMNS[5].d/U310  ( .A(n4681), .B(n4680), .Z(\w0[6][35] ) );
  XOR \MIXCOLUMNS[5].d/U309  ( .A(n4873), .B(n4682), .Z(n4680) );
  XOR \MIXCOLUMNS[5].d/U308  ( .A(n782), .B(n4866), .Z(n4681) );
  XOR \MIXCOLUMNS[5].d/U307  ( .A(n781), .B(n297), .Z(n4682) );
  XOR \MIXCOLUMNS[5].d/U306  ( .A(n781), .B(n296), .Z(n4875) );
  XOR \MIXCOLUMNS[5].d/U305  ( .A(n4684), .B(n4683), .Z(\w0[6][36] ) );
  XOR \MIXCOLUMNS[5].d/U304  ( .A(n4875), .B(n4685), .Z(n4683) );
  XOR \MIXCOLUMNS[5].d/U303  ( .A(n780), .B(n4866), .Z(n4684) );
  XOR \MIXCOLUMNS[5].d/U302  ( .A(n779), .B(n295), .Z(n4685) );
  XOR \MIXCOLUMNS[5].d/U301  ( .A(n779), .B(n294), .Z(n4877) );
  XOR \MIXCOLUMNS[5].d/U300  ( .A(n4687), .B(n4686), .Z(\w0[6][37] ) );
  XOR \MIXCOLUMNS[5].d/U299  ( .A(n778), .B(n4877), .Z(n4686) );
  XOR \MIXCOLUMNS[5].d/U298  ( .A(n777), .B(n293), .Z(n4687) );
  XOR \MIXCOLUMNS[5].d/U297  ( .A(n777), .B(n292), .Z(n4879) );
  XOR \MIXCOLUMNS[5].d/U296  ( .A(n4689), .B(n4688), .Z(\w0[6][38] ) );
  XOR \MIXCOLUMNS[5].d/U295  ( .A(n4879), .B(n4690), .Z(n4688) );
  XOR \MIXCOLUMNS[5].d/U294  ( .A(n776), .B(n4866), .Z(n4689) );
  XOR \MIXCOLUMNS[5].d/U293  ( .A(n775), .B(n291), .Z(n4690) );
  XOR \MIXCOLUMNS[5].d/U292  ( .A(n775), .B(n290), .Z(n4881) );
  XOR \MIXCOLUMNS[5].d/U291  ( .A(n4881), .B(n4691), .Z(\w0[6][39] ) );
  XOR \MIXCOLUMNS[5].d/U290  ( .A(n289), .B(n4866), .Z(n4691) );
  XOR \MIXCOLUMNS[5].d/U289  ( .A(n300), .B(n786), .Z(n4870) );
  XOR \MIXCOLUMNS[5].d/U288  ( .A(n4870), .B(n4692), .Z(\w0[6][40] ) );
  XOR \MIXCOLUMNS[5].d/U287  ( .A(n299), .B(n4883), .Z(n4692) );
  XOR \MIXCOLUMNS[5].d/U286  ( .A(\w3[5][42] ), .B(\w3[5][34] ), .Z(n4872) );
  XOR \MIXCOLUMNS[5].d/U285  ( .A(n4872), .B(n4693), .Z(\w0[6][41] ) );
  XOR \MIXCOLUMNS[5].d/U284  ( .A(n786), .B(n4868), .Z(n4693) );
  XOR \MIXCOLUMNS[5].d/U283  ( .A(n297), .B(n784), .Z(n4874) );
  XOR \MIXCOLUMNS[5].d/U282  ( .A(n4874), .B(n4694), .Z(\w0[6][42] ) );
  XOR \MIXCOLUMNS[5].d/U281  ( .A(\w3[5][34] ), .B(n4871), .Z(n4694) );
  XOR \MIXCOLUMNS[5].d/U280  ( .A(n19), .B(n299), .Z(n4869) );
  XOR \MIXCOLUMNS[5].d/U279  ( .A(n295), .B(n782), .Z(n4876) );
  XOR \MIXCOLUMNS[5].d/U278  ( .A(n4696), .B(n4695), .Z(\w0[6][43] ) );
  XOR \MIXCOLUMNS[5].d/U277  ( .A(n4873), .B(n4876), .Z(n4695) );
  XOR \MIXCOLUMNS[5].d/U276  ( .A(n784), .B(n4869), .Z(n4696) );
  XOR \MIXCOLUMNS[5].d/U275  ( .A(n293), .B(n780), .Z(n4878) );
  XOR \MIXCOLUMNS[5].d/U274  ( .A(n4698), .B(n4697), .Z(\w0[6][44] ) );
  XOR \MIXCOLUMNS[5].d/U273  ( .A(n4875), .B(n4878), .Z(n4697) );
  XOR \MIXCOLUMNS[5].d/U272  ( .A(n782), .B(n4869), .Z(n4698) );
  XOR \MIXCOLUMNS[5].d/U271  ( .A(n291), .B(n778), .Z(n4880) );
  XOR \MIXCOLUMNS[5].d/U270  ( .A(n4880), .B(n4699), .Z(\w0[6][45] ) );
  XOR \MIXCOLUMNS[5].d/U269  ( .A(n780), .B(n4877), .Z(n4699) );
  XOR \MIXCOLUMNS[5].d/U268  ( .A(n289), .B(n776), .Z(n4882) );
  XOR \MIXCOLUMNS[5].d/U267  ( .A(n4701), .B(n4700), .Z(\w0[6][46] ) );
  XOR \MIXCOLUMNS[5].d/U266  ( .A(n4879), .B(n4882), .Z(n4700) );
  XOR \MIXCOLUMNS[5].d/U265  ( .A(n778), .B(n4869), .Z(n4701) );
  XOR \MIXCOLUMNS[5].d/U264  ( .A(n4881), .B(n4702), .Z(\w0[6][47] ) );
  XOR \MIXCOLUMNS[5].d/U263  ( .A(n776), .B(n4869), .Z(n4702) );
  XOR \MIXCOLUMNS[5].d/U262  ( .A(n4704), .B(n4703), .Z(\w0[6][48] ) );
  XOR \MIXCOLUMNS[5].d/U261  ( .A(n300), .B(n4869), .Z(n4703) );
  XOR \MIXCOLUMNS[5].d/U260  ( .A(n787), .B(n301), .Z(n4704) );
  XOR \MIXCOLUMNS[5].d/U259  ( .A(n4706), .B(n4705), .Z(\w0[6][49] ) );
  XOR \MIXCOLUMNS[5].d/U258  ( .A(\w3[5][42] ), .B(n4870), .Z(n4705) );
  XOR \MIXCOLUMNS[5].d/U257  ( .A(n785), .B(\w3[5][50] ), .Z(n4706) );
  XOR \MIXCOLUMNS[5].d/U256  ( .A(n4708), .B(n4707), .Z(\w0[6][50] ) );
  XOR \MIXCOLUMNS[5].d/U255  ( .A(n297), .B(n4872), .Z(n4707) );
  XOR \MIXCOLUMNS[5].d/U254  ( .A(\w3[5][58] ), .B(n298), .Z(n4708) );
  XOR \MIXCOLUMNS[5].d/U253  ( .A(n302), .B(n19), .Z(n4867) );
  XOR \MIXCOLUMNS[5].d/U252  ( .A(n4710), .B(n4709), .Z(\w0[6][51] ) );
  XOR \MIXCOLUMNS[5].d/U251  ( .A(n4874), .B(n4711), .Z(n4709) );
  XOR \MIXCOLUMNS[5].d/U250  ( .A(n295), .B(n4867), .Z(n4710) );
  XOR \MIXCOLUMNS[5].d/U249  ( .A(n783), .B(n296), .Z(n4711) );
  XOR \MIXCOLUMNS[5].d/U248  ( .A(n4713), .B(n4712), .Z(\w0[6][52] ) );
  XOR \MIXCOLUMNS[5].d/U247  ( .A(n4876), .B(n4714), .Z(n4712) );
  XOR \MIXCOLUMNS[5].d/U246  ( .A(n293), .B(n4867), .Z(n4713) );
  XOR \MIXCOLUMNS[5].d/U245  ( .A(n781), .B(n294), .Z(n4714) );
  XOR \MIXCOLUMNS[5].d/U244  ( .A(n4716), .B(n4715), .Z(\w0[6][53] ) );
  XOR \MIXCOLUMNS[5].d/U243  ( .A(n291), .B(n4878), .Z(n4715) );
  XOR \MIXCOLUMNS[5].d/U242  ( .A(n779), .B(n292), .Z(n4716) );
  XOR \MIXCOLUMNS[5].d/U241  ( .A(n4718), .B(n4717), .Z(\w0[6][54] ) );
  XOR \MIXCOLUMNS[5].d/U240  ( .A(n4880), .B(n4719), .Z(n4717) );
  XOR \MIXCOLUMNS[5].d/U239  ( .A(n289), .B(n4867), .Z(n4718) );
  XOR \MIXCOLUMNS[5].d/U238  ( .A(n777), .B(n290), .Z(n4719) );
  XOR \MIXCOLUMNS[5].d/U237  ( .A(n4882), .B(n4720), .Z(\w0[6][55] ) );
  XOR \MIXCOLUMNS[5].d/U236  ( .A(n775), .B(n4867), .Z(n4720) );
  XOR \MIXCOLUMNS[5].d/U235  ( .A(n4868), .B(n4721), .Z(\w0[6][56] ) );
  XOR \MIXCOLUMNS[5].d/U234  ( .A(n302), .B(n4869), .Z(n4721) );
  XOR \MIXCOLUMNS[5].d/U233  ( .A(n4870), .B(n4722), .Z(\w0[6][57] ) );
  XOR \MIXCOLUMNS[5].d/U232  ( .A(n301), .B(n4871), .Z(n4722) );
  XOR \MIXCOLUMNS[5].d/U231  ( .A(n4872), .B(n4723), .Z(\w0[6][58] ) );
  XOR \MIXCOLUMNS[5].d/U230  ( .A(\w3[5][50] ), .B(n4873), .Z(n4723) );
  XOR \MIXCOLUMNS[5].d/U229  ( .A(n4725), .B(n4724), .Z(\w0[6][59] ) );
  XOR \MIXCOLUMNS[5].d/U228  ( .A(n4875), .B(n4874), .Z(n4724) );
  XOR \MIXCOLUMNS[5].d/U227  ( .A(n298), .B(n4883), .Z(n4725) );
  XOR \MIXCOLUMNS[5].d/U226  ( .A(n4727), .B(n4726), .Z(\w0[6][60] ) );
  XOR \MIXCOLUMNS[5].d/U225  ( .A(n4877), .B(n4876), .Z(n4726) );
  XOR \MIXCOLUMNS[5].d/U224  ( .A(n296), .B(n4883), .Z(n4727) );
  XOR \MIXCOLUMNS[5].d/U223  ( .A(n4878), .B(n4728), .Z(\w0[6][61] ) );
  XOR \MIXCOLUMNS[5].d/U222  ( .A(n294), .B(n4879), .Z(n4728) );
  XOR \MIXCOLUMNS[5].d/U221  ( .A(n4730), .B(n4729), .Z(\w0[6][62] ) );
  XOR \MIXCOLUMNS[5].d/U220  ( .A(n4881), .B(n4880), .Z(n4729) );
  XOR \MIXCOLUMNS[5].d/U219  ( .A(n292), .B(n4883), .Z(n4730) );
  XOR \MIXCOLUMNS[5].d/U218  ( .A(n4882), .B(n4731), .Z(\w0[6][63] ) );
  XOR \MIXCOLUMNS[5].d/U217  ( .A(n290), .B(n4883), .Z(n4731) );
  XOR \MIXCOLUMNS[5].d/U216  ( .A(n774), .B(n288), .Z(n4901) );
  XOR \MIXCOLUMNS[5].d/U215  ( .A(n4733), .B(n4732), .Z(\w0[6][64] ) );
  XOR \MIXCOLUMNS[5].d/U214  ( .A(n773), .B(n4901), .Z(n4732) );
  XOR \MIXCOLUMNS[5].d/U213  ( .A(n772), .B(n18), .Z(n4733) );
  XOR \MIXCOLUMNS[5].d/U212  ( .A(n772), .B(n287), .Z(n4886) );
  XOR \MIXCOLUMNS[5].d/U211  ( .A(n4735), .B(n4734), .Z(\w0[6][65] ) );
  XOR \MIXCOLUMNS[5].d/U210  ( .A(\w3[5][66] ), .B(n4886), .Z(n4734) );
  XOR \MIXCOLUMNS[5].d/U209  ( .A(\w3[5][90] ), .B(n286), .Z(n4735) );
  XOR \MIXCOLUMNS[5].d/U208  ( .A(\w3[5][90] ), .B(\w3[5][82] ), .Z(n4889) );
  XOR \MIXCOLUMNS[5].d/U207  ( .A(n4737), .B(n4736), .Z(\w0[6][66] ) );
  XOR \MIXCOLUMNS[5].d/U206  ( .A(n771), .B(n4889), .Z(n4736) );
  XOR \MIXCOLUMNS[5].d/U205  ( .A(n770), .B(\w3[5][74] ), .Z(n4737) );
  XOR \MIXCOLUMNS[5].d/U204  ( .A(n774), .B(n285), .Z(n4884) );
  XOR \MIXCOLUMNS[5].d/U203  ( .A(n770), .B(n284), .Z(n4891) );
  XOR \MIXCOLUMNS[5].d/U202  ( .A(n4739), .B(n4738), .Z(\w0[6][67] ) );
  XOR \MIXCOLUMNS[5].d/U201  ( .A(n4891), .B(n4740), .Z(n4738) );
  XOR \MIXCOLUMNS[5].d/U200  ( .A(n769), .B(n4884), .Z(n4739) );
  XOR \MIXCOLUMNS[5].d/U199  ( .A(n768), .B(n283), .Z(n4740) );
  XOR \MIXCOLUMNS[5].d/U198  ( .A(n768), .B(n282), .Z(n4893) );
  XOR \MIXCOLUMNS[5].d/U197  ( .A(n4742), .B(n4741), .Z(\w0[6][68] ) );
  XOR \MIXCOLUMNS[5].d/U196  ( .A(n4893), .B(n4743), .Z(n4741) );
  XOR \MIXCOLUMNS[5].d/U195  ( .A(n767), .B(n4884), .Z(n4742) );
  XOR \MIXCOLUMNS[5].d/U194  ( .A(n766), .B(n281), .Z(n4743) );
  XOR \MIXCOLUMNS[5].d/U193  ( .A(n766), .B(n280), .Z(n4895) );
  XOR \MIXCOLUMNS[5].d/U192  ( .A(n4745), .B(n4744), .Z(\w0[6][69] ) );
  XOR \MIXCOLUMNS[5].d/U191  ( .A(n765), .B(n4895), .Z(n4744) );
  XOR \MIXCOLUMNS[5].d/U190  ( .A(n764), .B(n279), .Z(n4745) );
  XOR \MIXCOLUMNS[5].d/U189  ( .A(n764), .B(n278), .Z(n4897) );
  XOR \MIXCOLUMNS[5].d/U188  ( .A(n4747), .B(n4746), .Z(\w0[6][70] ) );
  XOR \MIXCOLUMNS[5].d/U187  ( .A(n4897), .B(n4748), .Z(n4746) );
  XOR \MIXCOLUMNS[5].d/U186  ( .A(n763), .B(n4884), .Z(n4747) );
  XOR \MIXCOLUMNS[5].d/U185  ( .A(n762), .B(n277), .Z(n4748) );
  XOR \MIXCOLUMNS[5].d/U184  ( .A(n762), .B(n276), .Z(n4899) );
  XOR \MIXCOLUMNS[5].d/U183  ( .A(n4899), .B(n4749), .Z(\w0[6][71] ) );
  XOR \MIXCOLUMNS[5].d/U182  ( .A(n275), .B(n4884), .Z(n4749) );
  XOR \MIXCOLUMNS[5].d/U181  ( .A(n286), .B(n773), .Z(n4888) );
  XOR \MIXCOLUMNS[5].d/U180  ( .A(n4888), .B(n4750), .Z(\w0[6][72] ) );
  XOR \MIXCOLUMNS[5].d/U179  ( .A(n285), .B(n4901), .Z(n4750) );
  XOR \MIXCOLUMNS[5].d/U178  ( .A(\w3[5][74] ), .B(\w3[5][66] ), .Z(n4890) );
  XOR \MIXCOLUMNS[5].d/U177  ( .A(n4890), .B(n4751), .Z(\w0[6][73] ) );
  XOR \MIXCOLUMNS[5].d/U176  ( .A(n773), .B(n4886), .Z(n4751) );
  XOR \MIXCOLUMNS[5].d/U175  ( .A(n283), .B(n771), .Z(n4892) );
  XOR \MIXCOLUMNS[5].d/U174  ( .A(n4892), .B(n4752), .Z(\w0[6][74] ) );
  XOR \MIXCOLUMNS[5].d/U173  ( .A(\w3[5][66] ), .B(n4889), .Z(n4752) );
  XOR \MIXCOLUMNS[5].d/U172  ( .A(n18), .B(n285), .Z(n4887) );
  XOR \MIXCOLUMNS[5].d/U171  ( .A(n281), .B(n769), .Z(n4894) );
  XOR \MIXCOLUMNS[5].d/U170  ( .A(n4754), .B(n4753), .Z(\w0[6][75] ) );
  XOR \MIXCOLUMNS[5].d/U169  ( .A(n4891), .B(n4894), .Z(n4753) );
  XOR \MIXCOLUMNS[5].d/U168  ( .A(n771), .B(n4887), .Z(n4754) );
  XOR \MIXCOLUMNS[5].d/U167  ( .A(n279), .B(n767), .Z(n4896) );
  XOR \MIXCOLUMNS[5].d/U166  ( .A(n4756), .B(n4755), .Z(\w0[6][76] ) );
  XOR \MIXCOLUMNS[5].d/U165  ( .A(n4893), .B(n4896), .Z(n4755) );
  XOR \MIXCOLUMNS[5].d/U164  ( .A(n769), .B(n4887), .Z(n4756) );
  XOR \MIXCOLUMNS[5].d/U163  ( .A(n277), .B(n765), .Z(n4898) );
  XOR \MIXCOLUMNS[5].d/U162  ( .A(n4898), .B(n4757), .Z(\w0[6][77] ) );
  XOR \MIXCOLUMNS[5].d/U161  ( .A(n767), .B(n4895), .Z(n4757) );
  XOR \MIXCOLUMNS[5].d/U160  ( .A(n275), .B(n763), .Z(n4900) );
  XOR \MIXCOLUMNS[5].d/U159  ( .A(n4759), .B(n4758), .Z(\w0[6][78] ) );
  XOR \MIXCOLUMNS[5].d/U158  ( .A(n4897), .B(n4900), .Z(n4758) );
  XOR \MIXCOLUMNS[5].d/U157  ( .A(n765), .B(n4887), .Z(n4759) );
  XOR \MIXCOLUMNS[5].d/U156  ( .A(n4899), .B(n4760), .Z(\w0[6][79] ) );
  XOR \MIXCOLUMNS[5].d/U155  ( .A(n763), .B(n4887), .Z(n4760) );
  XOR \MIXCOLUMNS[5].d/U154  ( .A(n4762), .B(n4761), .Z(\w0[6][80] ) );
  XOR \MIXCOLUMNS[5].d/U153  ( .A(n286), .B(n4887), .Z(n4761) );
  XOR \MIXCOLUMNS[5].d/U152  ( .A(n774), .B(n287), .Z(n4762) );
  XOR \MIXCOLUMNS[5].d/U151  ( .A(n4764), .B(n4763), .Z(\w0[6][81] ) );
  XOR \MIXCOLUMNS[5].d/U150  ( .A(\w3[5][74] ), .B(n4888), .Z(n4763) );
  XOR \MIXCOLUMNS[5].d/U149  ( .A(n772), .B(\w3[5][82] ), .Z(n4764) );
  XOR \MIXCOLUMNS[5].d/U148  ( .A(n4766), .B(n4765), .Z(\w0[6][82] ) );
  XOR \MIXCOLUMNS[5].d/U147  ( .A(n283), .B(n4890), .Z(n4765) );
  XOR \MIXCOLUMNS[5].d/U146  ( .A(\w3[5][90] ), .B(n284), .Z(n4766) );
  XOR \MIXCOLUMNS[5].d/U145  ( .A(n288), .B(n18), .Z(n4885) );
  XOR \MIXCOLUMNS[5].d/U144  ( .A(n4768), .B(n4767), .Z(\w0[6][83] ) );
  XOR \MIXCOLUMNS[5].d/U143  ( .A(n4892), .B(n4769), .Z(n4767) );
  XOR \MIXCOLUMNS[5].d/U142  ( .A(n281), .B(n4885), .Z(n4768) );
  XOR \MIXCOLUMNS[5].d/U141  ( .A(n770), .B(n282), .Z(n4769) );
  XOR \MIXCOLUMNS[5].d/U140  ( .A(n4771), .B(n4770), .Z(\w0[6][84] ) );
  XOR \MIXCOLUMNS[5].d/U139  ( .A(n4894), .B(n4772), .Z(n4770) );
  XOR \MIXCOLUMNS[5].d/U138  ( .A(n279), .B(n4885), .Z(n4771) );
  XOR \MIXCOLUMNS[5].d/U137  ( .A(n768), .B(n280), .Z(n4772) );
  XOR \MIXCOLUMNS[5].d/U136  ( .A(n4774), .B(n4773), .Z(\w0[6][85] ) );
  XOR \MIXCOLUMNS[5].d/U135  ( .A(n277), .B(n4896), .Z(n4773) );
  XOR \MIXCOLUMNS[5].d/U134  ( .A(n766), .B(n278), .Z(n4774) );
  XOR \MIXCOLUMNS[5].d/U133  ( .A(n4776), .B(n4775), .Z(\w0[6][86] ) );
  XOR \MIXCOLUMNS[5].d/U132  ( .A(n4898), .B(n4777), .Z(n4775) );
  XOR \MIXCOLUMNS[5].d/U131  ( .A(n275), .B(n4885), .Z(n4776) );
  XOR \MIXCOLUMNS[5].d/U130  ( .A(n764), .B(n276), .Z(n4777) );
  XOR \MIXCOLUMNS[5].d/U129  ( .A(n4900), .B(n4778), .Z(\w0[6][87] ) );
  XOR \MIXCOLUMNS[5].d/U128  ( .A(n762), .B(n4885), .Z(n4778) );
  XOR \MIXCOLUMNS[5].d/U127  ( .A(n4886), .B(n4779), .Z(\w0[6][88] ) );
  XOR \MIXCOLUMNS[5].d/U126  ( .A(n288), .B(n4887), .Z(n4779) );
  XOR \MIXCOLUMNS[5].d/U125  ( .A(n4888), .B(n4780), .Z(\w0[6][89] ) );
  XOR \MIXCOLUMNS[5].d/U124  ( .A(n287), .B(n4889), .Z(n4780) );
  XOR \MIXCOLUMNS[5].d/U123  ( .A(n4890), .B(n4781), .Z(\w0[6][90] ) );
  XOR \MIXCOLUMNS[5].d/U122  ( .A(\w3[5][82] ), .B(n4891), .Z(n4781) );
  XOR \MIXCOLUMNS[5].d/U121  ( .A(n4783), .B(n4782), .Z(\w0[6][91] ) );
  XOR \MIXCOLUMNS[5].d/U120  ( .A(n4893), .B(n4892), .Z(n4782) );
  XOR \MIXCOLUMNS[5].d/U119  ( .A(n284), .B(n4901), .Z(n4783) );
  XOR \MIXCOLUMNS[5].d/U118  ( .A(n4785), .B(n4784), .Z(\w0[6][92] ) );
  XOR \MIXCOLUMNS[5].d/U117  ( .A(n4895), .B(n4894), .Z(n4784) );
  XOR \MIXCOLUMNS[5].d/U116  ( .A(n282), .B(n4901), .Z(n4785) );
  XOR \MIXCOLUMNS[5].d/U115  ( .A(n4896), .B(n4786), .Z(\w0[6][93] ) );
  XOR \MIXCOLUMNS[5].d/U114  ( .A(n280), .B(n4897), .Z(n4786) );
  XOR \MIXCOLUMNS[5].d/U113  ( .A(n4788), .B(n4787), .Z(\w0[6][94] ) );
  XOR \MIXCOLUMNS[5].d/U112  ( .A(n4899), .B(n4898), .Z(n4787) );
  XOR \MIXCOLUMNS[5].d/U111  ( .A(n278), .B(n4901), .Z(n4788) );
  XOR \MIXCOLUMNS[5].d/U110  ( .A(n4900), .B(n4789), .Z(\w0[6][95] ) );
  XOR \MIXCOLUMNS[5].d/U109  ( .A(n276), .B(n4901), .Z(n4789) );
  XOR \MIXCOLUMNS[5].d/U108  ( .A(n761), .B(n274), .Z(n4919) );
  XOR \MIXCOLUMNS[5].d/U107  ( .A(n4791), .B(n4790), .Z(\w0[6][96] ) );
  XOR \MIXCOLUMNS[5].d/U106  ( .A(n760), .B(n4919), .Z(n4790) );
  XOR \MIXCOLUMNS[5].d/U105  ( .A(n759), .B(n17), .Z(n4791) );
  XOR \MIXCOLUMNS[5].d/U104  ( .A(n759), .B(n273), .Z(n4904) );
  XOR \MIXCOLUMNS[5].d/U103  ( .A(n4793), .B(n4792), .Z(\w0[6][97] ) );
  XOR \MIXCOLUMNS[5].d/U102  ( .A(\w3[5][98] ), .B(n4904), .Z(n4792) );
  XOR \MIXCOLUMNS[5].d/U101  ( .A(\w3[5][122] ), .B(n272), .Z(n4793) );
  XOR \MIXCOLUMNS[5].d/U100  ( .A(\w3[5][122] ), .B(\w3[5][114] ), .Z(n4907)
         );
  XOR \MIXCOLUMNS[5].d/U99  ( .A(n4795), .B(n4794), .Z(\w0[6][98] ) );
  XOR \MIXCOLUMNS[5].d/U98  ( .A(n758), .B(n4907), .Z(n4794) );
  XOR \MIXCOLUMNS[5].d/U97  ( .A(n757), .B(\w3[5][106] ), .Z(n4795) );
  XOR \MIXCOLUMNS[5].d/U96  ( .A(n761), .B(n271), .Z(n4902) );
  XOR \MIXCOLUMNS[5].d/U95  ( .A(n757), .B(n270), .Z(n4909) );
  XOR \MIXCOLUMNS[5].d/U94  ( .A(n4797), .B(n4796), .Z(\w0[6][99] ) );
  XOR \MIXCOLUMNS[5].d/U93  ( .A(n4909), .B(n4798), .Z(n4796) );
  XOR \MIXCOLUMNS[5].d/U92  ( .A(n756), .B(n4902), .Z(n4797) );
  XOR \MIXCOLUMNS[5].d/U91  ( .A(n755), .B(n269), .Z(n4798) );
  XOR \MIXCOLUMNS[5].d/U90  ( .A(n755), .B(n268), .Z(n4911) );
  XOR \MIXCOLUMNS[5].d/U89  ( .A(n4800), .B(n4799), .Z(\w0[6][100] ) );
  XOR \MIXCOLUMNS[5].d/U88  ( .A(n4911), .B(n4801), .Z(n4799) );
  XOR \MIXCOLUMNS[5].d/U87  ( .A(n754), .B(n4902), .Z(n4800) );
  XOR \MIXCOLUMNS[5].d/U86  ( .A(n753), .B(n267), .Z(n4801) );
  XOR \MIXCOLUMNS[5].d/U85  ( .A(n753), .B(n266), .Z(n4913) );
  XOR \MIXCOLUMNS[5].d/U84  ( .A(n4803), .B(n4802), .Z(\w0[6][101] ) );
  XOR \MIXCOLUMNS[5].d/U83  ( .A(n752), .B(n4913), .Z(n4802) );
  XOR \MIXCOLUMNS[5].d/U82  ( .A(n751), .B(n265), .Z(n4803) );
  XOR \MIXCOLUMNS[5].d/U81  ( .A(n751), .B(n264), .Z(n4915) );
  XOR \MIXCOLUMNS[5].d/U80  ( .A(n4805), .B(n4804), .Z(\w0[6][102] ) );
  XOR \MIXCOLUMNS[5].d/U79  ( .A(n4915), .B(n4806), .Z(n4804) );
  XOR \MIXCOLUMNS[5].d/U78  ( .A(n750), .B(n4902), .Z(n4805) );
  XOR \MIXCOLUMNS[5].d/U77  ( .A(n749), .B(n263), .Z(n4806) );
  XOR \MIXCOLUMNS[5].d/U76  ( .A(n749), .B(n262), .Z(n4917) );
  XOR \MIXCOLUMNS[5].d/U75  ( .A(n4917), .B(n4807), .Z(\w0[6][103] ) );
  XOR \MIXCOLUMNS[5].d/U74  ( .A(n261), .B(n4902), .Z(n4807) );
  XOR \MIXCOLUMNS[5].d/U73  ( .A(n272), .B(n760), .Z(n4906) );
  XOR \MIXCOLUMNS[5].d/U72  ( .A(n4906), .B(n4808), .Z(\w0[6][104] ) );
  XOR \MIXCOLUMNS[5].d/U71  ( .A(n271), .B(n4919), .Z(n4808) );
  XOR \MIXCOLUMNS[5].d/U70  ( .A(\w3[5][106] ), .B(\w3[5][98] ), .Z(n4908) );
  XOR \MIXCOLUMNS[5].d/U69  ( .A(n4908), .B(n4809), .Z(\w0[6][105] ) );
  XOR \MIXCOLUMNS[5].d/U68  ( .A(n760), .B(n4904), .Z(n4809) );
  XOR \MIXCOLUMNS[5].d/U67  ( .A(n269), .B(n758), .Z(n4910) );
  XOR \MIXCOLUMNS[5].d/U66  ( .A(n4910), .B(n4810), .Z(\w0[6][106] ) );
  XOR \MIXCOLUMNS[5].d/U65  ( .A(\w3[5][98] ), .B(n4907), .Z(n4810) );
  XOR \MIXCOLUMNS[5].d/U64  ( .A(n17), .B(n271), .Z(n4905) );
  XOR \MIXCOLUMNS[5].d/U63  ( .A(n267), .B(n756), .Z(n4912) );
  XOR \MIXCOLUMNS[5].d/U62  ( .A(n4812), .B(n4811), .Z(\w0[6][107] ) );
  XOR \MIXCOLUMNS[5].d/U61  ( .A(n4909), .B(n4912), .Z(n4811) );
  XOR \MIXCOLUMNS[5].d/U60  ( .A(n758), .B(n4905), .Z(n4812) );
  XOR \MIXCOLUMNS[5].d/U59  ( .A(n265), .B(n754), .Z(n4914) );
  XOR \MIXCOLUMNS[5].d/U58  ( .A(n4814), .B(n4813), .Z(\w0[6][108] ) );
  XOR \MIXCOLUMNS[5].d/U57  ( .A(n4911), .B(n4914), .Z(n4813) );
  XOR \MIXCOLUMNS[5].d/U56  ( .A(n756), .B(n4905), .Z(n4814) );
  XOR \MIXCOLUMNS[5].d/U55  ( .A(n263), .B(n752), .Z(n4916) );
  XOR \MIXCOLUMNS[5].d/U54  ( .A(n4916), .B(n4815), .Z(\w0[6][109] ) );
  XOR \MIXCOLUMNS[5].d/U53  ( .A(n754), .B(n4913), .Z(n4815) );
  XOR \MIXCOLUMNS[5].d/U52  ( .A(n261), .B(n750), .Z(n4918) );
  XOR \MIXCOLUMNS[5].d/U51  ( .A(n4817), .B(n4816), .Z(\w0[6][110] ) );
  XOR \MIXCOLUMNS[5].d/U50  ( .A(n4915), .B(n4918), .Z(n4816) );
  XOR \MIXCOLUMNS[5].d/U49  ( .A(n752), .B(n4905), .Z(n4817) );
  XOR \MIXCOLUMNS[5].d/U48  ( .A(n4917), .B(n4818), .Z(\w0[6][111] ) );
  XOR \MIXCOLUMNS[5].d/U47  ( .A(n750), .B(n4905), .Z(n4818) );
  XOR \MIXCOLUMNS[5].d/U46  ( .A(n4820), .B(n4819), .Z(\w0[6][112] ) );
  XOR \MIXCOLUMNS[5].d/U45  ( .A(n272), .B(n4905), .Z(n4819) );
  XOR \MIXCOLUMNS[5].d/U44  ( .A(n761), .B(n273), .Z(n4820) );
  XOR \MIXCOLUMNS[5].d/U43  ( .A(n4822), .B(n4821), .Z(\w0[6][113] ) );
  XOR \MIXCOLUMNS[5].d/U42  ( .A(\w3[5][106] ), .B(n4906), .Z(n4821) );
  XOR \MIXCOLUMNS[5].d/U41  ( .A(n759), .B(\w3[5][114] ), .Z(n4822) );
  XOR \MIXCOLUMNS[5].d/U40  ( .A(n4824), .B(n4823), .Z(\w0[6][114] ) );
  XOR \MIXCOLUMNS[5].d/U39  ( .A(n269), .B(n4908), .Z(n4823) );
  XOR \MIXCOLUMNS[5].d/U38  ( .A(\w3[5][122] ), .B(n270), .Z(n4824) );
  XOR \MIXCOLUMNS[5].d/U37  ( .A(n274), .B(n17), .Z(n4903) );
  XOR \MIXCOLUMNS[5].d/U36  ( .A(n4826), .B(n4825), .Z(\w0[6][115] ) );
  XOR \MIXCOLUMNS[5].d/U35  ( .A(n4910), .B(n4827), .Z(n4825) );
  XOR \MIXCOLUMNS[5].d/U34  ( .A(n267), .B(n4903), .Z(n4826) );
  XOR \MIXCOLUMNS[5].d/U33  ( .A(n757), .B(n268), .Z(n4827) );
  XOR \MIXCOLUMNS[5].d/U32  ( .A(n4829), .B(n4828), .Z(\w0[6][116] ) );
  XOR \MIXCOLUMNS[5].d/U31  ( .A(n4912), .B(n4830), .Z(n4828) );
  XOR \MIXCOLUMNS[5].d/U30  ( .A(n265), .B(n4903), .Z(n4829) );
  XOR \MIXCOLUMNS[5].d/U29  ( .A(n755), .B(n266), .Z(n4830) );
  XOR \MIXCOLUMNS[5].d/U28  ( .A(n4832), .B(n4831), .Z(\w0[6][117] ) );
  XOR \MIXCOLUMNS[5].d/U27  ( .A(n263), .B(n4914), .Z(n4831) );
  XOR \MIXCOLUMNS[5].d/U26  ( .A(n753), .B(n264), .Z(n4832) );
  XOR \MIXCOLUMNS[5].d/U25  ( .A(n4834), .B(n4833), .Z(\w0[6][118] ) );
  XOR \MIXCOLUMNS[5].d/U24  ( .A(n4916), .B(n4835), .Z(n4833) );
  XOR \MIXCOLUMNS[5].d/U23  ( .A(n261), .B(n4903), .Z(n4834) );
  XOR \MIXCOLUMNS[5].d/U22  ( .A(n751), .B(n262), .Z(n4835) );
  XOR \MIXCOLUMNS[5].d/U21  ( .A(n4918), .B(n4836), .Z(\w0[6][119] ) );
  XOR \MIXCOLUMNS[5].d/U20  ( .A(n749), .B(n4903), .Z(n4836) );
  XOR \MIXCOLUMNS[5].d/U19  ( .A(n4904), .B(n4837), .Z(\w0[6][120] ) );
  XOR \MIXCOLUMNS[5].d/U18  ( .A(n274), .B(n4905), .Z(n4837) );
  XOR \MIXCOLUMNS[5].d/U17  ( .A(n4906), .B(n4838), .Z(\w0[6][121] ) );
  XOR \MIXCOLUMNS[5].d/U16  ( .A(n273), .B(n4907), .Z(n4838) );
  XOR \MIXCOLUMNS[5].d/U15  ( .A(n4908), .B(n4839), .Z(\w0[6][122] ) );
  XOR \MIXCOLUMNS[5].d/U14  ( .A(\w3[5][114] ), .B(n4909), .Z(n4839) );
  XOR \MIXCOLUMNS[5].d/U13  ( .A(n4841), .B(n4840), .Z(\w0[6][123] ) );
  XOR \MIXCOLUMNS[5].d/U12  ( .A(n4911), .B(n4910), .Z(n4840) );
  XOR \MIXCOLUMNS[5].d/U11  ( .A(n270), .B(n4919), .Z(n4841) );
  XOR \MIXCOLUMNS[5].d/U10  ( .A(n4843), .B(n4842), .Z(\w0[6][124] ) );
  XOR \MIXCOLUMNS[5].d/U9  ( .A(n4913), .B(n4912), .Z(n4842) );
  XOR \MIXCOLUMNS[5].d/U8  ( .A(n268), .B(n4919), .Z(n4843) );
  XOR \MIXCOLUMNS[5].d/U7  ( .A(n4914), .B(n4844), .Z(\w0[6][125] ) );
  XOR \MIXCOLUMNS[5].d/U6  ( .A(n266), .B(n4915), .Z(n4844) );
  XOR \MIXCOLUMNS[5].d/U5  ( .A(n4846), .B(n4845), .Z(\w0[6][126] ) );
  XOR \MIXCOLUMNS[5].d/U4  ( .A(n4917), .B(n4916), .Z(n4845) );
  XOR \MIXCOLUMNS[5].d/U3  ( .A(n264), .B(n4919), .Z(n4846) );
  XOR \MIXCOLUMNS[5].d/U2  ( .A(n4918), .B(n4847), .Z(\w0[6][127] ) );
  XOR \MIXCOLUMNS[5].d/U1  ( .A(n262), .B(n4919), .Z(n4847) );
  XOR \MIXCOLUMNS[4].d/U432  ( .A(n748), .B(n260), .Z(n4561) );
  XOR \MIXCOLUMNS[4].d/U431  ( .A(n4313), .B(n4312), .Z(\w0[5][0] ) );
  XOR \MIXCOLUMNS[4].d/U430  ( .A(n747), .B(n4561), .Z(n4312) );
  XOR \MIXCOLUMNS[4].d/U429  ( .A(n746), .B(n16), .Z(n4313) );
  XOR \MIXCOLUMNS[4].d/U428  ( .A(n746), .B(n259), .Z(n4546) );
  XOR \MIXCOLUMNS[4].d/U427  ( .A(n4315), .B(n4314), .Z(\w0[5][1] ) );
  XOR \MIXCOLUMNS[4].d/U426  ( .A(\w3[4][2] ), .B(n4546), .Z(n4314) );
  XOR \MIXCOLUMNS[4].d/U425  ( .A(\w3[4][26] ), .B(n258), .Z(n4315) );
  XOR \MIXCOLUMNS[4].d/U424  ( .A(\w3[4][26] ), .B(\w3[4][18] ), .Z(n4549) );
  XOR \MIXCOLUMNS[4].d/U423  ( .A(n4317), .B(n4316), .Z(\w0[5][2] ) );
  XOR \MIXCOLUMNS[4].d/U422  ( .A(n745), .B(n4549), .Z(n4316) );
  XOR \MIXCOLUMNS[4].d/U421  ( .A(n744), .B(\w3[4][10] ), .Z(n4317) );
  XOR \MIXCOLUMNS[4].d/U420  ( .A(n748), .B(n257), .Z(n4544) );
  XOR \MIXCOLUMNS[4].d/U419  ( .A(n744), .B(n256), .Z(n4551) );
  XOR \MIXCOLUMNS[4].d/U418  ( .A(n4319), .B(n4318), .Z(\w0[5][3] ) );
  XOR \MIXCOLUMNS[4].d/U417  ( .A(n4551), .B(n4320), .Z(n4318) );
  XOR \MIXCOLUMNS[4].d/U416  ( .A(n743), .B(n4544), .Z(n4319) );
  XOR \MIXCOLUMNS[4].d/U415  ( .A(n742), .B(n255), .Z(n4320) );
  XOR \MIXCOLUMNS[4].d/U414  ( .A(n742), .B(n254), .Z(n4553) );
  XOR \MIXCOLUMNS[4].d/U413  ( .A(n4322), .B(n4321), .Z(\w0[5][4] ) );
  XOR \MIXCOLUMNS[4].d/U412  ( .A(n4553), .B(n4323), .Z(n4321) );
  XOR \MIXCOLUMNS[4].d/U411  ( .A(n741), .B(n4544), .Z(n4322) );
  XOR \MIXCOLUMNS[4].d/U410  ( .A(n740), .B(n253), .Z(n4323) );
  XOR \MIXCOLUMNS[4].d/U409  ( .A(n740), .B(n252), .Z(n4555) );
  XOR \MIXCOLUMNS[4].d/U408  ( .A(n4325), .B(n4324), .Z(\w0[5][5] ) );
  XOR \MIXCOLUMNS[4].d/U407  ( .A(n739), .B(n4555), .Z(n4324) );
  XOR \MIXCOLUMNS[4].d/U406  ( .A(n738), .B(n251), .Z(n4325) );
  XOR \MIXCOLUMNS[4].d/U405  ( .A(n738), .B(n250), .Z(n4557) );
  XOR \MIXCOLUMNS[4].d/U404  ( .A(n4327), .B(n4326), .Z(\w0[5][6] ) );
  XOR \MIXCOLUMNS[4].d/U403  ( .A(n4557), .B(n4328), .Z(n4326) );
  XOR \MIXCOLUMNS[4].d/U402  ( .A(n737), .B(n4544), .Z(n4327) );
  XOR \MIXCOLUMNS[4].d/U401  ( .A(n736), .B(n249), .Z(n4328) );
  XOR \MIXCOLUMNS[4].d/U400  ( .A(n736), .B(n248), .Z(n4559) );
  XOR \MIXCOLUMNS[4].d/U399  ( .A(n4559), .B(n4329), .Z(\w0[5][7] ) );
  XOR \MIXCOLUMNS[4].d/U398  ( .A(n247), .B(n4544), .Z(n4329) );
  XOR \MIXCOLUMNS[4].d/U397  ( .A(n258), .B(n747), .Z(n4548) );
  XOR \MIXCOLUMNS[4].d/U396  ( .A(n4548), .B(n4330), .Z(\w0[5][8] ) );
  XOR \MIXCOLUMNS[4].d/U395  ( .A(n257), .B(n4561), .Z(n4330) );
  XOR \MIXCOLUMNS[4].d/U394  ( .A(\w3[4][10] ), .B(\w3[4][2] ), .Z(n4550) );
  XOR \MIXCOLUMNS[4].d/U393  ( .A(n4550), .B(n4331), .Z(\w0[5][9] ) );
  XOR \MIXCOLUMNS[4].d/U392  ( .A(n747), .B(n4546), .Z(n4331) );
  XOR \MIXCOLUMNS[4].d/U391  ( .A(n255), .B(n745), .Z(n4552) );
  XOR \MIXCOLUMNS[4].d/U390  ( .A(n4552), .B(n4332), .Z(\w0[5][10] ) );
  XOR \MIXCOLUMNS[4].d/U389  ( .A(\w3[4][2] ), .B(n4549), .Z(n4332) );
  XOR \MIXCOLUMNS[4].d/U388  ( .A(n16), .B(n257), .Z(n4547) );
  XOR \MIXCOLUMNS[4].d/U387  ( .A(n253), .B(n743), .Z(n4554) );
  XOR \MIXCOLUMNS[4].d/U386  ( .A(n4334), .B(n4333), .Z(\w0[5][11] ) );
  XOR \MIXCOLUMNS[4].d/U385  ( .A(n4551), .B(n4554), .Z(n4333) );
  XOR \MIXCOLUMNS[4].d/U384  ( .A(n745), .B(n4547), .Z(n4334) );
  XOR \MIXCOLUMNS[4].d/U383  ( .A(n251), .B(n741), .Z(n4556) );
  XOR \MIXCOLUMNS[4].d/U382  ( .A(n4336), .B(n4335), .Z(\w0[5][12] ) );
  XOR \MIXCOLUMNS[4].d/U381  ( .A(n4553), .B(n4556), .Z(n4335) );
  XOR \MIXCOLUMNS[4].d/U380  ( .A(n743), .B(n4547), .Z(n4336) );
  XOR \MIXCOLUMNS[4].d/U379  ( .A(n249), .B(n739), .Z(n4558) );
  XOR \MIXCOLUMNS[4].d/U378  ( .A(n4558), .B(n4337), .Z(\w0[5][13] ) );
  XOR \MIXCOLUMNS[4].d/U377  ( .A(n741), .B(n4555), .Z(n4337) );
  XOR \MIXCOLUMNS[4].d/U376  ( .A(n247), .B(n737), .Z(n4560) );
  XOR \MIXCOLUMNS[4].d/U375  ( .A(n4339), .B(n4338), .Z(\w0[5][14] ) );
  XOR \MIXCOLUMNS[4].d/U374  ( .A(n4557), .B(n4560), .Z(n4338) );
  XOR \MIXCOLUMNS[4].d/U373  ( .A(n739), .B(n4547), .Z(n4339) );
  XOR \MIXCOLUMNS[4].d/U372  ( .A(n4559), .B(n4340), .Z(\w0[5][15] ) );
  XOR \MIXCOLUMNS[4].d/U371  ( .A(n737), .B(n4547), .Z(n4340) );
  XOR \MIXCOLUMNS[4].d/U370  ( .A(n4342), .B(n4341), .Z(\w0[5][16] ) );
  XOR \MIXCOLUMNS[4].d/U369  ( .A(n258), .B(n4547), .Z(n4341) );
  XOR \MIXCOLUMNS[4].d/U368  ( .A(n748), .B(n259), .Z(n4342) );
  XOR \MIXCOLUMNS[4].d/U367  ( .A(n4344), .B(n4343), .Z(\w0[5][17] ) );
  XOR \MIXCOLUMNS[4].d/U366  ( .A(\w3[4][10] ), .B(n4548), .Z(n4343) );
  XOR \MIXCOLUMNS[4].d/U365  ( .A(n746), .B(\w3[4][18] ), .Z(n4344) );
  XOR \MIXCOLUMNS[4].d/U364  ( .A(n4346), .B(n4345), .Z(\w0[5][18] ) );
  XOR \MIXCOLUMNS[4].d/U363  ( .A(n255), .B(n4550), .Z(n4345) );
  XOR \MIXCOLUMNS[4].d/U362  ( .A(\w3[4][26] ), .B(n256), .Z(n4346) );
  XOR \MIXCOLUMNS[4].d/U361  ( .A(n260), .B(n16), .Z(n4545) );
  XOR \MIXCOLUMNS[4].d/U360  ( .A(n4348), .B(n4347), .Z(\w0[5][19] ) );
  XOR \MIXCOLUMNS[4].d/U359  ( .A(n4552), .B(n4349), .Z(n4347) );
  XOR \MIXCOLUMNS[4].d/U358  ( .A(n253), .B(n4545), .Z(n4348) );
  XOR \MIXCOLUMNS[4].d/U357  ( .A(n744), .B(n254), .Z(n4349) );
  XOR \MIXCOLUMNS[4].d/U356  ( .A(n4351), .B(n4350), .Z(\w0[5][20] ) );
  XOR \MIXCOLUMNS[4].d/U355  ( .A(n4554), .B(n4352), .Z(n4350) );
  XOR \MIXCOLUMNS[4].d/U354  ( .A(n251), .B(n4545), .Z(n4351) );
  XOR \MIXCOLUMNS[4].d/U353  ( .A(n742), .B(n252), .Z(n4352) );
  XOR \MIXCOLUMNS[4].d/U352  ( .A(n4354), .B(n4353), .Z(\w0[5][21] ) );
  XOR \MIXCOLUMNS[4].d/U351  ( .A(n249), .B(n4556), .Z(n4353) );
  XOR \MIXCOLUMNS[4].d/U350  ( .A(n740), .B(n250), .Z(n4354) );
  XOR \MIXCOLUMNS[4].d/U349  ( .A(n4356), .B(n4355), .Z(\w0[5][22] ) );
  XOR \MIXCOLUMNS[4].d/U348  ( .A(n4558), .B(n4357), .Z(n4355) );
  XOR \MIXCOLUMNS[4].d/U347  ( .A(n247), .B(n4545), .Z(n4356) );
  XOR \MIXCOLUMNS[4].d/U346  ( .A(n738), .B(n248), .Z(n4357) );
  XOR \MIXCOLUMNS[4].d/U345  ( .A(n4560), .B(n4358), .Z(\w0[5][23] ) );
  XOR \MIXCOLUMNS[4].d/U344  ( .A(n736), .B(n4545), .Z(n4358) );
  XOR \MIXCOLUMNS[4].d/U343  ( .A(n4546), .B(n4359), .Z(\w0[5][24] ) );
  XOR \MIXCOLUMNS[4].d/U342  ( .A(n260), .B(n4547), .Z(n4359) );
  XOR \MIXCOLUMNS[4].d/U341  ( .A(n4548), .B(n4360), .Z(\w0[5][25] ) );
  XOR \MIXCOLUMNS[4].d/U340  ( .A(n259), .B(n4549), .Z(n4360) );
  XOR \MIXCOLUMNS[4].d/U339  ( .A(n4550), .B(n4361), .Z(\w0[5][26] ) );
  XOR \MIXCOLUMNS[4].d/U338  ( .A(\w3[4][18] ), .B(n4551), .Z(n4361) );
  XOR \MIXCOLUMNS[4].d/U337  ( .A(n4363), .B(n4362), .Z(\w0[5][27] ) );
  XOR \MIXCOLUMNS[4].d/U336  ( .A(n4553), .B(n4552), .Z(n4362) );
  XOR \MIXCOLUMNS[4].d/U335  ( .A(n256), .B(n4561), .Z(n4363) );
  XOR \MIXCOLUMNS[4].d/U334  ( .A(n4365), .B(n4364), .Z(\w0[5][28] ) );
  XOR \MIXCOLUMNS[4].d/U333  ( .A(n4555), .B(n4554), .Z(n4364) );
  XOR \MIXCOLUMNS[4].d/U332  ( .A(n254), .B(n4561), .Z(n4365) );
  XOR \MIXCOLUMNS[4].d/U331  ( .A(n4556), .B(n4366), .Z(\w0[5][29] ) );
  XOR \MIXCOLUMNS[4].d/U330  ( .A(n252), .B(n4557), .Z(n4366) );
  XOR \MIXCOLUMNS[4].d/U329  ( .A(n4368), .B(n4367), .Z(\w0[5][30] ) );
  XOR \MIXCOLUMNS[4].d/U328  ( .A(n4559), .B(n4558), .Z(n4367) );
  XOR \MIXCOLUMNS[4].d/U327  ( .A(n250), .B(n4561), .Z(n4368) );
  XOR \MIXCOLUMNS[4].d/U326  ( .A(n4560), .B(n4369), .Z(\w0[5][31] ) );
  XOR \MIXCOLUMNS[4].d/U325  ( .A(n248), .B(n4561), .Z(n4369) );
  XOR \MIXCOLUMNS[4].d/U324  ( .A(n735), .B(n246), .Z(n4579) );
  XOR \MIXCOLUMNS[4].d/U323  ( .A(n4371), .B(n4370), .Z(\w0[5][32] ) );
  XOR \MIXCOLUMNS[4].d/U322  ( .A(n734), .B(n4579), .Z(n4370) );
  XOR \MIXCOLUMNS[4].d/U321  ( .A(n733), .B(n15), .Z(n4371) );
  XOR \MIXCOLUMNS[4].d/U320  ( .A(n733), .B(n245), .Z(n4564) );
  XOR \MIXCOLUMNS[4].d/U319  ( .A(n4373), .B(n4372), .Z(\w0[5][33] ) );
  XOR \MIXCOLUMNS[4].d/U318  ( .A(\w3[4][34] ), .B(n4564), .Z(n4372) );
  XOR \MIXCOLUMNS[4].d/U317  ( .A(\w3[4][58] ), .B(n244), .Z(n4373) );
  XOR \MIXCOLUMNS[4].d/U316  ( .A(\w3[4][58] ), .B(\w3[4][50] ), .Z(n4567) );
  XOR \MIXCOLUMNS[4].d/U315  ( .A(n4375), .B(n4374), .Z(\w0[5][34] ) );
  XOR \MIXCOLUMNS[4].d/U314  ( .A(n732), .B(n4567), .Z(n4374) );
  XOR \MIXCOLUMNS[4].d/U313  ( .A(n731), .B(\w3[4][42] ), .Z(n4375) );
  XOR \MIXCOLUMNS[4].d/U312  ( .A(n735), .B(n243), .Z(n4562) );
  XOR \MIXCOLUMNS[4].d/U311  ( .A(n731), .B(n242), .Z(n4569) );
  XOR \MIXCOLUMNS[4].d/U310  ( .A(n4377), .B(n4376), .Z(\w0[5][35] ) );
  XOR \MIXCOLUMNS[4].d/U309  ( .A(n4569), .B(n4378), .Z(n4376) );
  XOR \MIXCOLUMNS[4].d/U308  ( .A(n730), .B(n4562), .Z(n4377) );
  XOR \MIXCOLUMNS[4].d/U307  ( .A(n729), .B(n241), .Z(n4378) );
  XOR \MIXCOLUMNS[4].d/U306  ( .A(n729), .B(n240), .Z(n4571) );
  XOR \MIXCOLUMNS[4].d/U305  ( .A(n4380), .B(n4379), .Z(\w0[5][36] ) );
  XOR \MIXCOLUMNS[4].d/U304  ( .A(n4571), .B(n4381), .Z(n4379) );
  XOR \MIXCOLUMNS[4].d/U303  ( .A(n728), .B(n4562), .Z(n4380) );
  XOR \MIXCOLUMNS[4].d/U302  ( .A(n727), .B(n239), .Z(n4381) );
  XOR \MIXCOLUMNS[4].d/U301  ( .A(n727), .B(n238), .Z(n4573) );
  XOR \MIXCOLUMNS[4].d/U300  ( .A(n4383), .B(n4382), .Z(\w0[5][37] ) );
  XOR \MIXCOLUMNS[4].d/U299  ( .A(n726), .B(n4573), .Z(n4382) );
  XOR \MIXCOLUMNS[4].d/U298  ( .A(n725), .B(n237), .Z(n4383) );
  XOR \MIXCOLUMNS[4].d/U297  ( .A(n725), .B(n236), .Z(n4575) );
  XOR \MIXCOLUMNS[4].d/U296  ( .A(n4385), .B(n4384), .Z(\w0[5][38] ) );
  XOR \MIXCOLUMNS[4].d/U295  ( .A(n4575), .B(n4386), .Z(n4384) );
  XOR \MIXCOLUMNS[4].d/U294  ( .A(n724), .B(n4562), .Z(n4385) );
  XOR \MIXCOLUMNS[4].d/U293  ( .A(n723), .B(n235), .Z(n4386) );
  XOR \MIXCOLUMNS[4].d/U292  ( .A(n723), .B(n234), .Z(n4577) );
  XOR \MIXCOLUMNS[4].d/U291  ( .A(n4577), .B(n4387), .Z(\w0[5][39] ) );
  XOR \MIXCOLUMNS[4].d/U290  ( .A(n233), .B(n4562), .Z(n4387) );
  XOR \MIXCOLUMNS[4].d/U289  ( .A(n244), .B(n734), .Z(n4566) );
  XOR \MIXCOLUMNS[4].d/U288  ( .A(n4566), .B(n4388), .Z(\w0[5][40] ) );
  XOR \MIXCOLUMNS[4].d/U287  ( .A(n243), .B(n4579), .Z(n4388) );
  XOR \MIXCOLUMNS[4].d/U286  ( .A(\w3[4][42] ), .B(\w3[4][34] ), .Z(n4568) );
  XOR \MIXCOLUMNS[4].d/U285  ( .A(n4568), .B(n4389), .Z(\w0[5][41] ) );
  XOR \MIXCOLUMNS[4].d/U284  ( .A(n734), .B(n4564), .Z(n4389) );
  XOR \MIXCOLUMNS[4].d/U283  ( .A(n241), .B(n732), .Z(n4570) );
  XOR \MIXCOLUMNS[4].d/U282  ( .A(n4570), .B(n4390), .Z(\w0[5][42] ) );
  XOR \MIXCOLUMNS[4].d/U281  ( .A(\w3[4][34] ), .B(n4567), .Z(n4390) );
  XOR \MIXCOLUMNS[4].d/U280  ( .A(n15), .B(n243), .Z(n4565) );
  XOR \MIXCOLUMNS[4].d/U279  ( .A(n239), .B(n730), .Z(n4572) );
  XOR \MIXCOLUMNS[4].d/U278  ( .A(n4392), .B(n4391), .Z(\w0[5][43] ) );
  XOR \MIXCOLUMNS[4].d/U277  ( .A(n4569), .B(n4572), .Z(n4391) );
  XOR \MIXCOLUMNS[4].d/U276  ( .A(n732), .B(n4565), .Z(n4392) );
  XOR \MIXCOLUMNS[4].d/U275  ( .A(n237), .B(n728), .Z(n4574) );
  XOR \MIXCOLUMNS[4].d/U274  ( .A(n4394), .B(n4393), .Z(\w0[5][44] ) );
  XOR \MIXCOLUMNS[4].d/U273  ( .A(n4571), .B(n4574), .Z(n4393) );
  XOR \MIXCOLUMNS[4].d/U272  ( .A(n730), .B(n4565), .Z(n4394) );
  XOR \MIXCOLUMNS[4].d/U271  ( .A(n235), .B(n726), .Z(n4576) );
  XOR \MIXCOLUMNS[4].d/U270  ( .A(n4576), .B(n4395), .Z(\w0[5][45] ) );
  XOR \MIXCOLUMNS[4].d/U269  ( .A(n728), .B(n4573), .Z(n4395) );
  XOR \MIXCOLUMNS[4].d/U268  ( .A(n233), .B(n724), .Z(n4578) );
  XOR \MIXCOLUMNS[4].d/U267  ( .A(n4397), .B(n4396), .Z(\w0[5][46] ) );
  XOR \MIXCOLUMNS[4].d/U266  ( .A(n4575), .B(n4578), .Z(n4396) );
  XOR \MIXCOLUMNS[4].d/U265  ( .A(n726), .B(n4565), .Z(n4397) );
  XOR \MIXCOLUMNS[4].d/U264  ( .A(n4577), .B(n4398), .Z(\w0[5][47] ) );
  XOR \MIXCOLUMNS[4].d/U263  ( .A(n724), .B(n4565), .Z(n4398) );
  XOR \MIXCOLUMNS[4].d/U262  ( .A(n4400), .B(n4399), .Z(\w0[5][48] ) );
  XOR \MIXCOLUMNS[4].d/U261  ( .A(n244), .B(n4565), .Z(n4399) );
  XOR \MIXCOLUMNS[4].d/U260  ( .A(n735), .B(n245), .Z(n4400) );
  XOR \MIXCOLUMNS[4].d/U259  ( .A(n4402), .B(n4401), .Z(\w0[5][49] ) );
  XOR \MIXCOLUMNS[4].d/U258  ( .A(\w3[4][42] ), .B(n4566), .Z(n4401) );
  XOR \MIXCOLUMNS[4].d/U257  ( .A(n733), .B(\w3[4][50] ), .Z(n4402) );
  XOR \MIXCOLUMNS[4].d/U256  ( .A(n4404), .B(n4403), .Z(\w0[5][50] ) );
  XOR \MIXCOLUMNS[4].d/U255  ( .A(n241), .B(n4568), .Z(n4403) );
  XOR \MIXCOLUMNS[4].d/U254  ( .A(\w3[4][58] ), .B(n242), .Z(n4404) );
  XOR \MIXCOLUMNS[4].d/U253  ( .A(n246), .B(n15), .Z(n4563) );
  XOR \MIXCOLUMNS[4].d/U252  ( .A(n4406), .B(n4405), .Z(\w0[5][51] ) );
  XOR \MIXCOLUMNS[4].d/U251  ( .A(n4570), .B(n4407), .Z(n4405) );
  XOR \MIXCOLUMNS[4].d/U250  ( .A(n239), .B(n4563), .Z(n4406) );
  XOR \MIXCOLUMNS[4].d/U249  ( .A(n731), .B(n240), .Z(n4407) );
  XOR \MIXCOLUMNS[4].d/U248  ( .A(n4409), .B(n4408), .Z(\w0[5][52] ) );
  XOR \MIXCOLUMNS[4].d/U247  ( .A(n4572), .B(n4410), .Z(n4408) );
  XOR \MIXCOLUMNS[4].d/U246  ( .A(n237), .B(n4563), .Z(n4409) );
  XOR \MIXCOLUMNS[4].d/U245  ( .A(n729), .B(n238), .Z(n4410) );
  XOR \MIXCOLUMNS[4].d/U244  ( .A(n4412), .B(n4411), .Z(\w0[5][53] ) );
  XOR \MIXCOLUMNS[4].d/U243  ( .A(n235), .B(n4574), .Z(n4411) );
  XOR \MIXCOLUMNS[4].d/U242  ( .A(n727), .B(n236), .Z(n4412) );
  XOR \MIXCOLUMNS[4].d/U241  ( .A(n4414), .B(n4413), .Z(\w0[5][54] ) );
  XOR \MIXCOLUMNS[4].d/U240  ( .A(n4576), .B(n4415), .Z(n4413) );
  XOR \MIXCOLUMNS[4].d/U239  ( .A(n233), .B(n4563), .Z(n4414) );
  XOR \MIXCOLUMNS[4].d/U238  ( .A(n725), .B(n234), .Z(n4415) );
  XOR \MIXCOLUMNS[4].d/U237  ( .A(n4578), .B(n4416), .Z(\w0[5][55] ) );
  XOR \MIXCOLUMNS[4].d/U236  ( .A(n723), .B(n4563), .Z(n4416) );
  XOR \MIXCOLUMNS[4].d/U235  ( .A(n4564), .B(n4417), .Z(\w0[5][56] ) );
  XOR \MIXCOLUMNS[4].d/U234  ( .A(n246), .B(n4565), .Z(n4417) );
  XOR \MIXCOLUMNS[4].d/U233  ( .A(n4566), .B(n4418), .Z(\w0[5][57] ) );
  XOR \MIXCOLUMNS[4].d/U232  ( .A(n245), .B(n4567), .Z(n4418) );
  XOR \MIXCOLUMNS[4].d/U231  ( .A(n4568), .B(n4419), .Z(\w0[5][58] ) );
  XOR \MIXCOLUMNS[4].d/U230  ( .A(\w3[4][50] ), .B(n4569), .Z(n4419) );
  XOR \MIXCOLUMNS[4].d/U229  ( .A(n4421), .B(n4420), .Z(\w0[5][59] ) );
  XOR \MIXCOLUMNS[4].d/U228  ( .A(n4571), .B(n4570), .Z(n4420) );
  XOR \MIXCOLUMNS[4].d/U227  ( .A(n242), .B(n4579), .Z(n4421) );
  XOR \MIXCOLUMNS[4].d/U226  ( .A(n4423), .B(n4422), .Z(\w0[5][60] ) );
  XOR \MIXCOLUMNS[4].d/U225  ( .A(n4573), .B(n4572), .Z(n4422) );
  XOR \MIXCOLUMNS[4].d/U224  ( .A(n240), .B(n4579), .Z(n4423) );
  XOR \MIXCOLUMNS[4].d/U223  ( .A(n4574), .B(n4424), .Z(\w0[5][61] ) );
  XOR \MIXCOLUMNS[4].d/U222  ( .A(n238), .B(n4575), .Z(n4424) );
  XOR \MIXCOLUMNS[4].d/U221  ( .A(n4426), .B(n4425), .Z(\w0[5][62] ) );
  XOR \MIXCOLUMNS[4].d/U220  ( .A(n4577), .B(n4576), .Z(n4425) );
  XOR \MIXCOLUMNS[4].d/U219  ( .A(n236), .B(n4579), .Z(n4426) );
  XOR \MIXCOLUMNS[4].d/U218  ( .A(n4578), .B(n4427), .Z(\w0[5][63] ) );
  XOR \MIXCOLUMNS[4].d/U217  ( .A(n234), .B(n4579), .Z(n4427) );
  XOR \MIXCOLUMNS[4].d/U216  ( .A(n722), .B(n232), .Z(n4597) );
  XOR \MIXCOLUMNS[4].d/U215  ( .A(n4429), .B(n4428), .Z(\w0[5][64] ) );
  XOR \MIXCOLUMNS[4].d/U214  ( .A(n721), .B(n4597), .Z(n4428) );
  XOR \MIXCOLUMNS[4].d/U213  ( .A(n720), .B(n14), .Z(n4429) );
  XOR \MIXCOLUMNS[4].d/U212  ( .A(n720), .B(n231), .Z(n4582) );
  XOR \MIXCOLUMNS[4].d/U211  ( .A(n4431), .B(n4430), .Z(\w0[5][65] ) );
  XOR \MIXCOLUMNS[4].d/U210  ( .A(\w3[4][66] ), .B(n4582), .Z(n4430) );
  XOR \MIXCOLUMNS[4].d/U209  ( .A(\w3[4][90] ), .B(n230), .Z(n4431) );
  XOR \MIXCOLUMNS[4].d/U208  ( .A(\w3[4][90] ), .B(\w3[4][82] ), .Z(n4585) );
  XOR \MIXCOLUMNS[4].d/U207  ( .A(n4433), .B(n4432), .Z(\w0[5][66] ) );
  XOR \MIXCOLUMNS[4].d/U206  ( .A(n719), .B(n4585), .Z(n4432) );
  XOR \MIXCOLUMNS[4].d/U205  ( .A(n718), .B(\w3[4][74] ), .Z(n4433) );
  XOR \MIXCOLUMNS[4].d/U204  ( .A(n722), .B(n229), .Z(n4580) );
  XOR \MIXCOLUMNS[4].d/U203  ( .A(n718), .B(n228), .Z(n4587) );
  XOR \MIXCOLUMNS[4].d/U202  ( .A(n4435), .B(n4434), .Z(\w0[5][67] ) );
  XOR \MIXCOLUMNS[4].d/U201  ( .A(n4587), .B(n4436), .Z(n4434) );
  XOR \MIXCOLUMNS[4].d/U200  ( .A(n717), .B(n4580), .Z(n4435) );
  XOR \MIXCOLUMNS[4].d/U199  ( .A(n716), .B(n227), .Z(n4436) );
  XOR \MIXCOLUMNS[4].d/U198  ( .A(n716), .B(n226), .Z(n4589) );
  XOR \MIXCOLUMNS[4].d/U197  ( .A(n4438), .B(n4437), .Z(\w0[5][68] ) );
  XOR \MIXCOLUMNS[4].d/U196  ( .A(n4589), .B(n4439), .Z(n4437) );
  XOR \MIXCOLUMNS[4].d/U195  ( .A(n715), .B(n4580), .Z(n4438) );
  XOR \MIXCOLUMNS[4].d/U194  ( .A(n714), .B(n225), .Z(n4439) );
  XOR \MIXCOLUMNS[4].d/U193  ( .A(n714), .B(n224), .Z(n4591) );
  XOR \MIXCOLUMNS[4].d/U192  ( .A(n4441), .B(n4440), .Z(\w0[5][69] ) );
  XOR \MIXCOLUMNS[4].d/U191  ( .A(n713), .B(n4591), .Z(n4440) );
  XOR \MIXCOLUMNS[4].d/U190  ( .A(n712), .B(n223), .Z(n4441) );
  XOR \MIXCOLUMNS[4].d/U189  ( .A(n712), .B(n222), .Z(n4593) );
  XOR \MIXCOLUMNS[4].d/U188  ( .A(n4443), .B(n4442), .Z(\w0[5][70] ) );
  XOR \MIXCOLUMNS[4].d/U187  ( .A(n4593), .B(n4444), .Z(n4442) );
  XOR \MIXCOLUMNS[4].d/U186  ( .A(n711), .B(n4580), .Z(n4443) );
  XOR \MIXCOLUMNS[4].d/U185  ( .A(n710), .B(n221), .Z(n4444) );
  XOR \MIXCOLUMNS[4].d/U184  ( .A(n710), .B(n220), .Z(n4595) );
  XOR \MIXCOLUMNS[4].d/U183  ( .A(n4595), .B(n4445), .Z(\w0[5][71] ) );
  XOR \MIXCOLUMNS[4].d/U182  ( .A(n219), .B(n4580), .Z(n4445) );
  XOR \MIXCOLUMNS[4].d/U181  ( .A(n230), .B(n721), .Z(n4584) );
  XOR \MIXCOLUMNS[4].d/U180  ( .A(n4584), .B(n4446), .Z(\w0[5][72] ) );
  XOR \MIXCOLUMNS[4].d/U179  ( .A(n229), .B(n4597), .Z(n4446) );
  XOR \MIXCOLUMNS[4].d/U178  ( .A(\w3[4][74] ), .B(\w3[4][66] ), .Z(n4586) );
  XOR \MIXCOLUMNS[4].d/U177  ( .A(n4586), .B(n4447), .Z(\w0[5][73] ) );
  XOR \MIXCOLUMNS[4].d/U176  ( .A(n721), .B(n4582), .Z(n4447) );
  XOR \MIXCOLUMNS[4].d/U175  ( .A(n227), .B(n719), .Z(n4588) );
  XOR \MIXCOLUMNS[4].d/U174  ( .A(n4588), .B(n4448), .Z(\w0[5][74] ) );
  XOR \MIXCOLUMNS[4].d/U173  ( .A(\w3[4][66] ), .B(n4585), .Z(n4448) );
  XOR \MIXCOLUMNS[4].d/U172  ( .A(n14), .B(n229), .Z(n4583) );
  XOR \MIXCOLUMNS[4].d/U171  ( .A(n225), .B(n717), .Z(n4590) );
  XOR \MIXCOLUMNS[4].d/U170  ( .A(n4450), .B(n4449), .Z(\w0[5][75] ) );
  XOR \MIXCOLUMNS[4].d/U169  ( .A(n4587), .B(n4590), .Z(n4449) );
  XOR \MIXCOLUMNS[4].d/U168  ( .A(n719), .B(n4583), .Z(n4450) );
  XOR \MIXCOLUMNS[4].d/U167  ( .A(n223), .B(n715), .Z(n4592) );
  XOR \MIXCOLUMNS[4].d/U166  ( .A(n4452), .B(n4451), .Z(\w0[5][76] ) );
  XOR \MIXCOLUMNS[4].d/U165  ( .A(n4589), .B(n4592), .Z(n4451) );
  XOR \MIXCOLUMNS[4].d/U164  ( .A(n717), .B(n4583), .Z(n4452) );
  XOR \MIXCOLUMNS[4].d/U163  ( .A(n221), .B(n713), .Z(n4594) );
  XOR \MIXCOLUMNS[4].d/U162  ( .A(n4594), .B(n4453), .Z(\w0[5][77] ) );
  XOR \MIXCOLUMNS[4].d/U161  ( .A(n715), .B(n4591), .Z(n4453) );
  XOR \MIXCOLUMNS[4].d/U160  ( .A(n219), .B(n711), .Z(n4596) );
  XOR \MIXCOLUMNS[4].d/U159  ( .A(n4455), .B(n4454), .Z(\w0[5][78] ) );
  XOR \MIXCOLUMNS[4].d/U158  ( .A(n4593), .B(n4596), .Z(n4454) );
  XOR \MIXCOLUMNS[4].d/U157  ( .A(n713), .B(n4583), .Z(n4455) );
  XOR \MIXCOLUMNS[4].d/U156  ( .A(n4595), .B(n4456), .Z(\w0[5][79] ) );
  XOR \MIXCOLUMNS[4].d/U155  ( .A(n711), .B(n4583), .Z(n4456) );
  XOR \MIXCOLUMNS[4].d/U154  ( .A(n4458), .B(n4457), .Z(\w0[5][80] ) );
  XOR \MIXCOLUMNS[4].d/U153  ( .A(n230), .B(n4583), .Z(n4457) );
  XOR \MIXCOLUMNS[4].d/U152  ( .A(n722), .B(n231), .Z(n4458) );
  XOR \MIXCOLUMNS[4].d/U151  ( .A(n4460), .B(n4459), .Z(\w0[5][81] ) );
  XOR \MIXCOLUMNS[4].d/U150  ( .A(\w3[4][74] ), .B(n4584), .Z(n4459) );
  XOR \MIXCOLUMNS[4].d/U149  ( .A(n720), .B(\w3[4][82] ), .Z(n4460) );
  XOR \MIXCOLUMNS[4].d/U148  ( .A(n4462), .B(n4461), .Z(\w0[5][82] ) );
  XOR \MIXCOLUMNS[4].d/U147  ( .A(n227), .B(n4586), .Z(n4461) );
  XOR \MIXCOLUMNS[4].d/U146  ( .A(\w3[4][90] ), .B(n228), .Z(n4462) );
  XOR \MIXCOLUMNS[4].d/U145  ( .A(n232), .B(n14), .Z(n4581) );
  XOR \MIXCOLUMNS[4].d/U144  ( .A(n4464), .B(n4463), .Z(\w0[5][83] ) );
  XOR \MIXCOLUMNS[4].d/U143  ( .A(n4588), .B(n4465), .Z(n4463) );
  XOR \MIXCOLUMNS[4].d/U142  ( .A(n225), .B(n4581), .Z(n4464) );
  XOR \MIXCOLUMNS[4].d/U141  ( .A(n718), .B(n226), .Z(n4465) );
  XOR \MIXCOLUMNS[4].d/U140  ( .A(n4467), .B(n4466), .Z(\w0[5][84] ) );
  XOR \MIXCOLUMNS[4].d/U139  ( .A(n4590), .B(n4468), .Z(n4466) );
  XOR \MIXCOLUMNS[4].d/U138  ( .A(n223), .B(n4581), .Z(n4467) );
  XOR \MIXCOLUMNS[4].d/U137  ( .A(n716), .B(n224), .Z(n4468) );
  XOR \MIXCOLUMNS[4].d/U136  ( .A(n4470), .B(n4469), .Z(\w0[5][85] ) );
  XOR \MIXCOLUMNS[4].d/U135  ( .A(n221), .B(n4592), .Z(n4469) );
  XOR \MIXCOLUMNS[4].d/U134  ( .A(n714), .B(n222), .Z(n4470) );
  XOR \MIXCOLUMNS[4].d/U133  ( .A(n4472), .B(n4471), .Z(\w0[5][86] ) );
  XOR \MIXCOLUMNS[4].d/U132  ( .A(n4594), .B(n4473), .Z(n4471) );
  XOR \MIXCOLUMNS[4].d/U131  ( .A(n219), .B(n4581), .Z(n4472) );
  XOR \MIXCOLUMNS[4].d/U130  ( .A(n712), .B(n220), .Z(n4473) );
  XOR \MIXCOLUMNS[4].d/U129  ( .A(n4596), .B(n4474), .Z(\w0[5][87] ) );
  XOR \MIXCOLUMNS[4].d/U128  ( .A(n710), .B(n4581), .Z(n4474) );
  XOR \MIXCOLUMNS[4].d/U127  ( .A(n4582), .B(n4475), .Z(\w0[5][88] ) );
  XOR \MIXCOLUMNS[4].d/U126  ( .A(n232), .B(n4583), .Z(n4475) );
  XOR \MIXCOLUMNS[4].d/U125  ( .A(n4584), .B(n4476), .Z(\w0[5][89] ) );
  XOR \MIXCOLUMNS[4].d/U124  ( .A(n231), .B(n4585), .Z(n4476) );
  XOR \MIXCOLUMNS[4].d/U123  ( .A(n4586), .B(n4477), .Z(\w0[5][90] ) );
  XOR \MIXCOLUMNS[4].d/U122  ( .A(\w3[4][82] ), .B(n4587), .Z(n4477) );
  XOR \MIXCOLUMNS[4].d/U121  ( .A(n4479), .B(n4478), .Z(\w0[5][91] ) );
  XOR \MIXCOLUMNS[4].d/U120  ( .A(n4589), .B(n4588), .Z(n4478) );
  XOR \MIXCOLUMNS[4].d/U119  ( .A(n228), .B(n4597), .Z(n4479) );
  XOR \MIXCOLUMNS[4].d/U118  ( .A(n4481), .B(n4480), .Z(\w0[5][92] ) );
  XOR \MIXCOLUMNS[4].d/U117  ( .A(n4591), .B(n4590), .Z(n4480) );
  XOR \MIXCOLUMNS[4].d/U116  ( .A(n226), .B(n4597), .Z(n4481) );
  XOR \MIXCOLUMNS[4].d/U115  ( .A(n4592), .B(n4482), .Z(\w0[5][93] ) );
  XOR \MIXCOLUMNS[4].d/U114  ( .A(n224), .B(n4593), .Z(n4482) );
  XOR \MIXCOLUMNS[4].d/U113  ( .A(n4484), .B(n4483), .Z(\w0[5][94] ) );
  XOR \MIXCOLUMNS[4].d/U112  ( .A(n4595), .B(n4594), .Z(n4483) );
  XOR \MIXCOLUMNS[4].d/U111  ( .A(n222), .B(n4597), .Z(n4484) );
  XOR \MIXCOLUMNS[4].d/U110  ( .A(n4596), .B(n4485), .Z(\w0[5][95] ) );
  XOR \MIXCOLUMNS[4].d/U109  ( .A(n220), .B(n4597), .Z(n4485) );
  XOR \MIXCOLUMNS[4].d/U108  ( .A(n709), .B(n218), .Z(n4615) );
  XOR \MIXCOLUMNS[4].d/U107  ( .A(n4487), .B(n4486), .Z(\w0[5][96] ) );
  XOR \MIXCOLUMNS[4].d/U106  ( .A(n708), .B(n4615), .Z(n4486) );
  XOR \MIXCOLUMNS[4].d/U105  ( .A(n707), .B(n13), .Z(n4487) );
  XOR \MIXCOLUMNS[4].d/U104  ( .A(n707), .B(n217), .Z(n4600) );
  XOR \MIXCOLUMNS[4].d/U103  ( .A(n4489), .B(n4488), .Z(\w0[5][97] ) );
  XOR \MIXCOLUMNS[4].d/U102  ( .A(\w3[4][98] ), .B(n4600), .Z(n4488) );
  XOR \MIXCOLUMNS[4].d/U101  ( .A(\w3[4][122] ), .B(n216), .Z(n4489) );
  XOR \MIXCOLUMNS[4].d/U100  ( .A(\w3[4][122] ), .B(\w3[4][114] ), .Z(n4603)
         );
  XOR \MIXCOLUMNS[4].d/U99  ( .A(n4491), .B(n4490), .Z(\w0[5][98] ) );
  XOR \MIXCOLUMNS[4].d/U98  ( .A(n706), .B(n4603), .Z(n4490) );
  XOR \MIXCOLUMNS[4].d/U97  ( .A(n705), .B(\w3[4][106] ), .Z(n4491) );
  XOR \MIXCOLUMNS[4].d/U96  ( .A(n709), .B(n215), .Z(n4598) );
  XOR \MIXCOLUMNS[4].d/U95  ( .A(n705), .B(n214), .Z(n4605) );
  XOR \MIXCOLUMNS[4].d/U94  ( .A(n4493), .B(n4492), .Z(\w0[5][99] ) );
  XOR \MIXCOLUMNS[4].d/U93  ( .A(n4605), .B(n4494), .Z(n4492) );
  XOR \MIXCOLUMNS[4].d/U92  ( .A(n704), .B(n4598), .Z(n4493) );
  XOR \MIXCOLUMNS[4].d/U91  ( .A(n703), .B(n213), .Z(n4494) );
  XOR \MIXCOLUMNS[4].d/U90  ( .A(n703), .B(n212), .Z(n4607) );
  XOR \MIXCOLUMNS[4].d/U89  ( .A(n4496), .B(n4495), .Z(\w0[5][100] ) );
  XOR \MIXCOLUMNS[4].d/U88  ( .A(n4607), .B(n4497), .Z(n4495) );
  XOR \MIXCOLUMNS[4].d/U87  ( .A(n702), .B(n4598), .Z(n4496) );
  XOR \MIXCOLUMNS[4].d/U86  ( .A(n701), .B(n211), .Z(n4497) );
  XOR \MIXCOLUMNS[4].d/U85  ( .A(n701), .B(n210), .Z(n4609) );
  XOR \MIXCOLUMNS[4].d/U84  ( .A(n4499), .B(n4498), .Z(\w0[5][101] ) );
  XOR \MIXCOLUMNS[4].d/U83  ( .A(n700), .B(n4609), .Z(n4498) );
  XOR \MIXCOLUMNS[4].d/U82  ( .A(n699), .B(n209), .Z(n4499) );
  XOR \MIXCOLUMNS[4].d/U81  ( .A(n699), .B(n208), .Z(n4611) );
  XOR \MIXCOLUMNS[4].d/U80  ( .A(n4501), .B(n4500), .Z(\w0[5][102] ) );
  XOR \MIXCOLUMNS[4].d/U79  ( .A(n4611), .B(n4502), .Z(n4500) );
  XOR \MIXCOLUMNS[4].d/U78  ( .A(n698), .B(n4598), .Z(n4501) );
  XOR \MIXCOLUMNS[4].d/U77  ( .A(n697), .B(n207), .Z(n4502) );
  XOR \MIXCOLUMNS[4].d/U76  ( .A(n697), .B(n206), .Z(n4613) );
  XOR \MIXCOLUMNS[4].d/U75  ( .A(n4613), .B(n4503), .Z(\w0[5][103] ) );
  XOR \MIXCOLUMNS[4].d/U74  ( .A(n205), .B(n4598), .Z(n4503) );
  XOR \MIXCOLUMNS[4].d/U73  ( .A(n216), .B(n708), .Z(n4602) );
  XOR \MIXCOLUMNS[4].d/U72  ( .A(n4602), .B(n4504), .Z(\w0[5][104] ) );
  XOR \MIXCOLUMNS[4].d/U71  ( .A(n215), .B(n4615), .Z(n4504) );
  XOR \MIXCOLUMNS[4].d/U70  ( .A(\w3[4][106] ), .B(\w3[4][98] ), .Z(n4604) );
  XOR \MIXCOLUMNS[4].d/U69  ( .A(n4604), .B(n4505), .Z(\w0[5][105] ) );
  XOR \MIXCOLUMNS[4].d/U68  ( .A(n708), .B(n4600), .Z(n4505) );
  XOR \MIXCOLUMNS[4].d/U67  ( .A(n213), .B(n706), .Z(n4606) );
  XOR \MIXCOLUMNS[4].d/U66  ( .A(n4606), .B(n4506), .Z(\w0[5][106] ) );
  XOR \MIXCOLUMNS[4].d/U65  ( .A(\w3[4][98] ), .B(n4603), .Z(n4506) );
  XOR \MIXCOLUMNS[4].d/U64  ( .A(n13), .B(n215), .Z(n4601) );
  XOR \MIXCOLUMNS[4].d/U63  ( .A(n211), .B(n704), .Z(n4608) );
  XOR \MIXCOLUMNS[4].d/U62  ( .A(n4508), .B(n4507), .Z(\w0[5][107] ) );
  XOR \MIXCOLUMNS[4].d/U61  ( .A(n4605), .B(n4608), .Z(n4507) );
  XOR \MIXCOLUMNS[4].d/U60  ( .A(n706), .B(n4601), .Z(n4508) );
  XOR \MIXCOLUMNS[4].d/U59  ( .A(n209), .B(n702), .Z(n4610) );
  XOR \MIXCOLUMNS[4].d/U58  ( .A(n4510), .B(n4509), .Z(\w0[5][108] ) );
  XOR \MIXCOLUMNS[4].d/U57  ( .A(n4607), .B(n4610), .Z(n4509) );
  XOR \MIXCOLUMNS[4].d/U56  ( .A(n704), .B(n4601), .Z(n4510) );
  XOR \MIXCOLUMNS[4].d/U55  ( .A(n207), .B(n700), .Z(n4612) );
  XOR \MIXCOLUMNS[4].d/U54  ( .A(n4612), .B(n4511), .Z(\w0[5][109] ) );
  XOR \MIXCOLUMNS[4].d/U53  ( .A(n702), .B(n4609), .Z(n4511) );
  XOR \MIXCOLUMNS[4].d/U52  ( .A(n205), .B(n698), .Z(n4614) );
  XOR \MIXCOLUMNS[4].d/U51  ( .A(n4513), .B(n4512), .Z(\w0[5][110] ) );
  XOR \MIXCOLUMNS[4].d/U50  ( .A(n4611), .B(n4614), .Z(n4512) );
  XOR \MIXCOLUMNS[4].d/U49  ( .A(n700), .B(n4601), .Z(n4513) );
  XOR \MIXCOLUMNS[4].d/U48  ( .A(n4613), .B(n4514), .Z(\w0[5][111] ) );
  XOR \MIXCOLUMNS[4].d/U47  ( .A(n698), .B(n4601), .Z(n4514) );
  XOR \MIXCOLUMNS[4].d/U46  ( .A(n4516), .B(n4515), .Z(\w0[5][112] ) );
  XOR \MIXCOLUMNS[4].d/U45  ( .A(n216), .B(n4601), .Z(n4515) );
  XOR \MIXCOLUMNS[4].d/U44  ( .A(n709), .B(n217), .Z(n4516) );
  XOR \MIXCOLUMNS[4].d/U43  ( .A(n4518), .B(n4517), .Z(\w0[5][113] ) );
  XOR \MIXCOLUMNS[4].d/U42  ( .A(\w3[4][106] ), .B(n4602), .Z(n4517) );
  XOR \MIXCOLUMNS[4].d/U41  ( .A(n707), .B(\w3[4][114] ), .Z(n4518) );
  XOR \MIXCOLUMNS[4].d/U40  ( .A(n4520), .B(n4519), .Z(\w0[5][114] ) );
  XOR \MIXCOLUMNS[4].d/U39  ( .A(n213), .B(n4604), .Z(n4519) );
  XOR \MIXCOLUMNS[4].d/U38  ( .A(\w3[4][122] ), .B(n214), .Z(n4520) );
  XOR \MIXCOLUMNS[4].d/U37  ( .A(n218), .B(n13), .Z(n4599) );
  XOR \MIXCOLUMNS[4].d/U36  ( .A(n4522), .B(n4521), .Z(\w0[5][115] ) );
  XOR \MIXCOLUMNS[4].d/U35  ( .A(n4606), .B(n4523), .Z(n4521) );
  XOR \MIXCOLUMNS[4].d/U34  ( .A(n211), .B(n4599), .Z(n4522) );
  XOR \MIXCOLUMNS[4].d/U33  ( .A(n705), .B(n212), .Z(n4523) );
  XOR \MIXCOLUMNS[4].d/U32  ( .A(n4525), .B(n4524), .Z(\w0[5][116] ) );
  XOR \MIXCOLUMNS[4].d/U31  ( .A(n4608), .B(n4526), .Z(n4524) );
  XOR \MIXCOLUMNS[4].d/U30  ( .A(n209), .B(n4599), .Z(n4525) );
  XOR \MIXCOLUMNS[4].d/U29  ( .A(n703), .B(n210), .Z(n4526) );
  XOR \MIXCOLUMNS[4].d/U28  ( .A(n4528), .B(n4527), .Z(\w0[5][117] ) );
  XOR \MIXCOLUMNS[4].d/U27  ( .A(n207), .B(n4610), .Z(n4527) );
  XOR \MIXCOLUMNS[4].d/U26  ( .A(n701), .B(n208), .Z(n4528) );
  XOR \MIXCOLUMNS[4].d/U25  ( .A(n4530), .B(n4529), .Z(\w0[5][118] ) );
  XOR \MIXCOLUMNS[4].d/U24  ( .A(n4612), .B(n4531), .Z(n4529) );
  XOR \MIXCOLUMNS[4].d/U23  ( .A(n205), .B(n4599), .Z(n4530) );
  XOR \MIXCOLUMNS[4].d/U22  ( .A(n699), .B(n206), .Z(n4531) );
  XOR \MIXCOLUMNS[4].d/U21  ( .A(n4614), .B(n4532), .Z(\w0[5][119] ) );
  XOR \MIXCOLUMNS[4].d/U20  ( .A(n697), .B(n4599), .Z(n4532) );
  XOR \MIXCOLUMNS[4].d/U19  ( .A(n4600), .B(n4533), .Z(\w0[5][120] ) );
  XOR \MIXCOLUMNS[4].d/U18  ( .A(n218), .B(n4601), .Z(n4533) );
  XOR \MIXCOLUMNS[4].d/U17  ( .A(n4602), .B(n4534), .Z(\w0[5][121] ) );
  XOR \MIXCOLUMNS[4].d/U16  ( .A(n217), .B(n4603), .Z(n4534) );
  XOR \MIXCOLUMNS[4].d/U15  ( .A(n4604), .B(n4535), .Z(\w0[5][122] ) );
  XOR \MIXCOLUMNS[4].d/U14  ( .A(\w3[4][114] ), .B(n4605), .Z(n4535) );
  XOR \MIXCOLUMNS[4].d/U13  ( .A(n4537), .B(n4536), .Z(\w0[5][123] ) );
  XOR \MIXCOLUMNS[4].d/U12  ( .A(n4607), .B(n4606), .Z(n4536) );
  XOR \MIXCOLUMNS[4].d/U11  ( .A(n214), .B(n4615), .Z(n4537) );
  XOR \MIXCOLUMNS[4].d/U10  ( .A(n4539), .B(n4538), .Z(\w0[5][124] ) );
  XOR \MIXCOLUMNS[4].d/U9  ( .A(n4609), .B(n4608), .Z(n4538) );
  XOR \MIXCOLUMNS[4].d/U8  ( .A(n212), .B(n4615), .Z(n4539) );
  XOR \MIXCOLUMNS[4].d/U7  ( .A(n4610), .B(n4540), .Z(\w0[5][125] ) );
  XOR \MIXCOLUMNS[4].d/U6  ( .A(n210), .B(n4611), .Z(n4540) );
  XOR \MIXCOLUMNS[4].d/U5  ( .A(n4542), .B(n4541), .Z(\w0[5][126] ) );
  XOR \MIXCOLUMNS[4].d/U4  ( .A(n4613), .B(n4612), .Z(n4541) );
  XOR \MIXCOLUMNS[4].d/U3  ( .A(n208), .B(n4615), .Z(n4542) );
  XOR \MIXCOLUMNS[4].d/U2  ( .A(n4614), .B(n4543), .Z(\w0[5][127] ) );
  XOR \MIXCOLUMNS[4].d/U1  ( .A(n206), .B(n4615), .Z(n4543) );
  XOR \MIXCOLUMNS[3].d/U432  ( .A(n696), .B(n204), .Z(n4257) );
  XOR \MIXCOLUMNS[3].d/U431  ( .A(n4009), .B(n4008), .Z(\w0[4][0] ) );
  XOR \MIXCOLUMNS[3].d/U430  ( .A(n695), .B(n4257), .Z(n4008) );
  XOR \MIXCOLUMNS[3].d/U429  ( .A(n694), .B(n12), .Z(n4009) );
  XOR \MIXCOLUMNS[3].d/U428  ( .A(n694), .B(n203), .Z(n4242) );
  XOR \MIXCOLUMNS[3].d/U427  ( .A(n4011), .B(n4010), .Z(\w0[4][1] ) );
  XOR \MIXCOLUMNS[3].d/U426  ( .A(\w3[3][2] ), .B(n4242), .Z(n4010) );
  XOR \MIXCOLUMNS[3].d/U425  ( .A(\w3[3][26] ), .B(n202), .Z(n4011) );
  XOR \MIXCOLUMNS[3].d/U424  ( .A(\w3[3][26] ), .B(\w3[3][18] ), .Z(n4245) );
  XOR \MIXCOLUMNS[3].d/U423  ( .A(n4013), .B(n4012), .Z(\w0[4][2] ) );
  XOR \MIXCOLUMNS[3].d/U422  ( .A(n693), .B(n4245), .Z(n4012) );
  XOR \MIXCOLUMNS[3].d/U421  ( .A(n692), .B(\w3[3][10] ), .Z(n4013) );
  XOR \MIXCOLUMNS[3].d/U420  ( .A(n696), .B(n201), .Z(n4240) );
  XOR \MIXCOLUMNS[3].d/U419  ( .A(n692), .B(n200), .Z(n4247) );
  XOR \MIXCOLUMNS[3].d/U418  ( .A(n4015), .B(n4014), .Z(\w0[4][3] ) );
  XOR \MIXCOLUMNS[3].d/U417  ( .A(n4247), .B(n4016), .Z(n4014) );
  XOR \MIXCOLUMNS[3].d/U416  ( .A(n691), .B(n4240), .Z(n4015) );
  XOR \MIXCOLUMNS[3].d/U415  ( .A(n690), .B(n199), .Z(n4016) );
  XOR \MIXCOLUMNS[3].d/U414  ( .A(n690), .B(n198), .Z(n4249) );
  XOR \MIXCOLUMNS[3].d/U413  ( .A(n4018), .B(n4017), .Z(\w0[4][4] ) );
  XOR \MIXCOLUMNS[3].d/U412  ( .A(n4249), .B(n4019), .Z(n4017) );
  XOR \MIXCOLUMNS[3].d/U411  ( .A(n689), .B(n4240), .Z(n4018) );
  XOR \MIXCOLUMNS[3].d/U410  ( .A(n688), .B(n197), .Z(n4019) );
  XOR \MIXCOLUMNS[3].d/U409  ( .A(n688), .B(n196), .Z(n4251) );
  XOR \MIXCOLUMNS[3].d/U408  ( .A(n4021), .B(n4020), .Z(\w0[4][5] ) );
  XOR \MIXCOLUMNS[3].d/U407  ( .A(n687), .B(n4251), .Z(n4020) );
  XOR \MIXCOLUMNS[3].d/U406  ( .A(n686), .B(n195), .Z(n4021) );
  XOR \MIXCOLUMNS[3].d/U405  ( .A(n686), .B(n194), .Z(n4253) );
  XOR \MIXCOLUMNS[3].d/U404  ( .A(n4023), .B(n4022), .Z(\w0[4][6] ) );
  XOR \MIXCOLUMNS[3].d/U403  ( .A(n4253), .B(n4024), .Z(n4022) );
  XOR \MIXCOLUMNS[3].d/U402  ( .A(n685), .B(n4240), .Z(n4023) );
  XOR \MIXCOLUMNS[3].d/U401  ( .A(n684), .B(n193), .Z(n4024) );
  XOR \MIXCOLUMNS[3].d/U400  ( .A(n684), .B(n192), .Z(n4255) );
  XOR \MIXCOLUMNS[3].d/U399  ( .A(n4255), .B(n4025), .Z(\w0[4][7] ) );
  XOR \MIXCOLUMNS[3].d/U398  ( .A(n191), .B(n4240), .Z(n4025) );
  XOR \MIXCOLUMNS[3].d/U397  ( .A(n202), .B(n695), .Z(n4244) );
  XOR \MIXCOLUMNS[3].d/U396  ( .A(n4244), .B(n4026), .Z(\w0[4][8] ) );
  XOR \MIXCOLUMNS[3].d/U395  ( .A(n201), .B(n4257), .Z(n4026) );
  XOR \MIXCOLUMNS[3].d/U394  ( .A(\w3[3][10] ), .B(\w3[3][2] ), .Z(n4246) );
  XOR \MIXCOLUMNS[3].d/U393  ( .A(n4246), .B(n4027), .Z(\w0[4][9] ) );
  XOR \MIXCOLUMNS[3].d/U392  ( .A(n695), .B(n4242), .Z(n4027) );
  XOR \MIXCOLUMNS[3].d/U391  ( .A(n199), .B(n693), .Z(n4248) );
  XOR \MIXCOLUMNS[3].d/U390  ( .A(n4248), .B(n4028), .Z(\w0[4][10] ) );
  XOR \MIXCOLUMNS[3].d/U389  ( .A(\w3[3][2] ), .B(n4245), .Z(n4028) );
  XOR \MIXCOLUMNS[3].d/U388  ( .A(n12), .B(n201), .Z(n4243) );
  XOR \MIXCOLUMNS[3].d/U387  ( .A(n197), .B(n691), .Z(n4250) );
  XOR \MIXCOLUMNS[3].d/U386  ( .A(n4030), .B(n4029), .Z(\w0[4][11] ) );
  XOR \MIXCOLUMNS[3].d/U385  ( .A(n4247), .B(n4250), .Z(n4029) );
  XOR \MIXCOLUMNS[3].d/U384  ( .A(n693), .B(n4243), .Z(n4030) );
  XOR \MIXCOLUMNS[3].d/U383  ( .A(n195), .B(n689), .Z(n4252) );
  XOR \MIXCOLUMNS[3].d/U382  ( .A(n4032), .B(n4031), .Z(\w0[4][12] ) );
  XOR \MIXCOLUMNS[3].d/U381  ( .A(n4249), .B(n4252), .Z(n4031) );
  XOR \MIXCOLUMNS[3].d/U380  ( .A(n691), .B(n4243), .Z(n4032) );
  XOR \MIXCOLUMNS[3].d/U379  ( .A(n193), .B(n687), .Z(n4254) );
  XOR \MIXCOLUMNS[3].d/U378  ( .A(n4254), .B(n4033), .Z(\w0[4][13] ) );
  XOR \MIXCOLUMNS[3].d/U377  ( .A(n689), .B(n4251), .Z(n4033) );
  XOR \MIXCOLUMNS[3].d/U376  ( .A(n191), .B(n685), .Z(n4256) );
  XOR \MIXCOLUMNS[3].d/U375  ( .A(n4035), .B(n4034), .Z(\w0[4][14] ) );
  XOR \MIXCOLUMNS[3].d/U374  ( .A(n4253), .B(n4256), .Z(n4034) );
  XOR \MIXCOLUMNS[3].d/U373  ( .A(n687), .B(n4243), .Z(n4035) );
  XOR \MIXCOLUMNS[3].d/U372  ( .A(n4255), .B(n4036), .Z(\w0[4][15] ) );
  XOR \MIXCOLUMNS[3].d/U371  ( .A(n685), .B(n4243), .Z(n4036) );
  XOR \MIXCOLUMNS[3].d/U370  ( .A(n4038), .B(n4037), .Z(\w0[4][16] ) );
  XOR \MIXCOLUMNS[3].d/U369  ( .A(n202), .B(n4243), .Z(n4037) );
  XOR \MIXCOLUMNS[3].d/U368  ( .A(n696), .B(n203), .Z(n4038) );
  XOR \MIXCOLUMNS[3].d/U367  ( .A(n4040), .B(n4039), .Z(\w0[4][17] ) );
  XOR \MIXCOLUMNS[3].d/U366  ( .A(\w3[3][10] ), .B(n4244), .Z(n4039) );
  XOR \MIXCOLUMNS[3].d/U365  ( .A(n694), .B(\w3[3][18] ), .Z(n4040) );
  XOR \MIXCOLUMNS[3].d/U364  ( .A(n4042), .B(n4041), .Z(\w0[4][18] ) );
  XOR \MIXCOLUMNS[3].d/U363  ( .A(n199), .B(n4246), .Z(n4041) );
  XOR \MIXCOLUMNS[3].d/U362  ( .A(\w3[3][26] ), .B(n200), .Z(n4042) );
  XOR \MIXCOLUMNS[3].d/U361  ( .A(n204), .B(n12), .Z(n4241) );
  XOR \MIXCOLUMNS[3].d/U360  ( .A(n4044), .B(n4043), .Z(\w0[4][19] ) );
  XOR \MIXCOLUMNS[3].d/U359  ( .A(n4248), .B(n4045), .Z(n4043) );
  XOR \MIXCOLUMNS[3].d/U358  ( .A(n197), .B(n4241), .Z(n4044) );
  XOR \MIXCOLUMNS[3].d/U357  ( .A(n692), .B(n198), .Z(n4045) );
  XOR \MIXCOLUMNS[3].d/U356  ( .A(n4047), .B(n4046), .Z(\w0[4][20] ) );
  XOR \MIXCOLUMNS[3].d/U355  ( .A(n4250), .B(n4048), .Z(n4046) );
  XOR \MIXCOLUMNS[3].d/U354  ( .A(n195), .B(n4241), .Z(n4047) );
  XOR \MIXCOLUMNS[3].d/U353  ( .A(n690), .B(n196), .Z(n4048) );
  XOR \MIXCOLUMNS[3].d/U352  ( .A(n4050), .B(n4049), .Z(\w0[4][21] ) );
  XOR \MIXCOLUMNS[3].d/U351  ( .A(n193), .B(n4252), .Z(n4049) );
  XOR \MIXCOLUMNS[3].d/U350  ( .A(n688), .B(n194), .Z(n4050) );
  XOR \MIXCOLUMNS[3].d/U349  ( .A(n4052), .B(n4051), .Z(\w0[4][22] ) );
  XOR \MIXCOLUMNS[3].d/U348  ( .A(n4254), .B(n4053), .Z(n4051) );
  XOR \MIXCOLUMNS[3].d/U347  ( .A(n191), .B(n4241), .Z(n4052) );
  XOR \MIXCOLUMNS[3].d/U346  ( .A(n686), .B(n192), .Z(n4053) );
  XOR \MIXCOLUMNS[3].d/U345  ( .A(n4256), .B(n4054), .Z(\w0[4][23] ) );
  XOR \MIXCOLUMNS[3].d/U344  ( .A(n684), .B(n4241), .Z(n4054) );
  XOR \MIXCOLUMNS[3].d/U343  ( .A(n4242), .B(n4055), .Z(\w0[4][24] ) );
  XOR \MIXCOLUMNS[3].d/U342  ( .A(n204), .B(n4243), .Z(n4055) );
  XOR \MIXCOLUMNS[3].d/U341  ( .A(n4244), .B(n4056), .Z(\w0[4][25] ) );
  XOR \MIXCOLUMNS[3].d/U340  ( .A(n203), .B(n4245), .Z(n4056) );
  XOR \MIXCOLUMNS[3].d/U339  ( .A(n4246), .B(n4057), .Z(\w0[4][26] ) );
  XOR \MIXCOLUMNS[3].d/U338  ( .A(\w3[3][18] ), .B(n4247), .Z(n4057) );
  XOR \MIXCOLUMNS[3].d/U337  ( .A(n4059), .B(n4058), .Z(\w0[4][27] ) );
  XOR \MIXCOLUMNS[3].d/U336  ( .A(n4249), .B(n4248), .Z(n4058) );
  XOR \MIXCOLUMNS[3].d/U335  ( .A(n200), .B(n4257), .Z(n4059) );
  XOR \MIXCOLUMNS[3].d/U334  ( .A(n4061), .B(n4060), .Z(\w0[4][28] ) );
  XOR \MIXCOLUMNS[3].d/U333  ( .A(n4251), .B(n4250), .Z(n4060) );
  XOR \MIXCOLUMNS[3].d/U332  ( .A(n198), .B(n4257), .Z(n4061) );
  XOR \MIXCOLUMNS[3].d/U331  ( .A(n4252), .B(n4062), .Z(\w0[4][29] ) );
  XOR \MIXCOLUMNS[3].d/U330  ( .A(n196), .B(n4253), .Z(n4062) );
  XOR \MIXCOLUMNS[3].d/U329  ( .A(n4064), .B(n4063), .Z(\w0[4][30] ) );
  XOR \MIXCOLUMNS[3].d/U328  ( .A(n4255), .B(n4254), .Z(n4063) );
  XOR \MIXCOLUMNS[3].d/U327  ( .A(n194), .B(n4257), .Z(n4064) );
  XOR \MIXCOLUMNS[3].d/U326  ( .A(n4256), .B(n4065), .Z(\w0[4][31] ) );
  XOR \MIXCOLUMNS[3].d/U325  ( .A(n192), .B(n4257), .Z(n4065) );
  XOR \MIXCOLUMNS[3].d/U324  ( .A(n683), .B(n190), .Z(n4275) );
  XOR \MIXCOLUMNS[3].d/U323  ( .A(n4067), .B(n4066), .Z(\w0[4][32] ) );
  XOR \MIXCOLUMNS[3].d/U322  ( .A(n682), .B(n4275), .Z(n4066) );
  XOR \MIXCOLUMNS[3].d/U321  ( .A(n681), .B(n11), .Z(n4067) );
  XOR \MIXCOLUMNS[3].d/U320  ( .A(n681), .B(n189), .Z(n4260) );
  XOR \MIXCOLUMNS[3].d/U319  ( .A(n4069), .B(n4068), .Z(\w0[4][33] ) );
  XOR \MIXCOLUMNS[3].d/U318  ( .A(\w3[3][34] ), .B(n4260), .Z(n4068) );
  XOR \MIXCOLUMNS[3].d/U317  ( .A(\w3[3][58] ), .B(n188), .Z(n4069) );
  XOR \MIXCOLUMNS[3].d/U316  ( .A(\w3[3][58] ), .B(\w3[3][50] ), .Z(n4263) );
  XOR \MIXCOLUMNS[3].d/U315  ( .A(n4071), .B(n4070), .Z(\w0[4][34] ) );
  XOR \MIXCOLUMNS[3].d/U314  ( .A(n680), .B(n4263), .Z(n4070) );
  XOR \MIXCOLUMNS[3].d/U313  ( .A(n679), .B(\w3[3][42] ), .Z(n4071) );
  XOR \MIXCOLUMNS[3].d/U312  ( .A(n683), .B(n187), .Z(n4258) );
  XOR \MIXCOLUMNS[3].d/U311  ( .A(n679), .B(n186), .Z(n4265) );
  XOR \MIXCOLUMNS[3].d/U310  ( .A(n4073), .B(n4072), .Z(\w0[4][35] ) );
  XOR \MIXCOLUMNS[3].d/U309  ( .A(n4265), .B(n4074), .Z(n4072) );
  XOR \MIXCOLUMNS[3].d/U308  ( .A(n678), .B(n4258), .Z(n4073) );
  XOR \MIXCOLUMNS[3].d/U307  ( .A(n677), .B(n185), .Z(n4074) );
  XOR \MIXCOLUMNS[3].d/U306  ( .A(n677), .B(n184), .Z(n4267) );
  XOR \MIXCOLUMNS[3].d/U305  ( .A(n4076), .B(n4075), .Z(\w0[4][36] ) );
  XOR \MIXCOLUMNS[3].d/U304  ( .A(n4267), .B(n4077), .Z(n4075) );
  XOR \MIXCOLUMNS[3].d/U303  ( .A(n676), .B(n4258), .Z(n4076) );
  XOR \MIXCOLUMNS[3].d/U302  ( .A(n675), .B(n183), .Z(n4077) );
  XOR \MIXCOLUMNS[3].d/U301  ( .A(n675), .B(n182), .Z(n4269) );
  XOR \MIXCOLUMNS[3].d/U300  ( .A(n4079), .B(n4078), .Z(\w0[4][37] ) );
  XOR \MIXCOLUMNS[3].d/U299  ( .A(n674), .B(n4269), .Z(n4078) );
  XOR \MIXCOLUMNS[3].d/U298  ( .A(n673), .B(n181), .Z(n4079) );
  XOR \MIXCOLUMNS[3].d/U297  ( .A(n673), .B(n180), .Z(n4271) );
  XOR \MIXCOLUMNS[3].d/U296  ( .A(n4081), .B(n4080), .Z(\w0[4][38] ) );
  XOR \MIXCOLUMNS[3].d/U295  ( .A(n4271), .B(n4082), .Z(n4080) );
  XOR \MIXCOLUMNS[3].d/U294  ( .A(n672), .B(n4258), .Z(n4081) );
  XOR \MIXCOLUMNS[3].d/U293  ( .A(n671), .B(n179), .Z(n4082) );
  XOR \MIXCOLUMNS[3].d/U292  ( .A(n671), .B(n178), .Z(n4273) );
  XOR \MIXCOLUMNS[3].d/U291  ( .A(n4273), .B(n4083), .Z(\w0[4][39] ) );
  XOR \MIXCOLUMNS[3].d/U290  ( .A(n177), .B(n4258), .Z(n4083) );
  XOR \MIXCOLUMNS[3].d/U289  ( .A(n188), .B(n682), .Z(n4262) );
  XOR \MIXCOLUMNS[3].d/U288  ( .A(n4262), .B(n4084), .Z(\w0[4][40] ) );
  XOR \MIXCOLUMNS[3].d/U287  ( .A(n187), .B(n4275), .Z(n4084) );
  XOR \MIXCOLUMNS[3].d/U286  ( .A(\w3[3][42] ), .B(\w3[3][34] ), .Z(n4264) );
  XOR \MIXCOLUMNS[3].d/U285  ( .A(n4264), .B(n4085), .Z(\w0[4][41] ) );
  XOR \MIXCOLUMNS[3].d/U284  ( .A(n682), .B(n4260), .Z(n4085) );
  XOR \MIXCOLUMNS[3].d/U283  ( .A(n185), .B(n680), .Z(n4266) );
  XOR \MIXCOLUMNS[3].d/U282  ( .A(n4266), .B(n4086), .Z(\w0[4][42] ) );
  XOR \MIXCOLUMNS[3].d/U281  ( .A(\w3[3][34] ), .B(n4263), .Z(n4086) );
  XOR \MIXCOLUMNS[3].d/U280  ( .A(n11), .B(n187), .Z(n4261) );
  XOR \MIXCOLUMNS[3].d/U279  ( .A(n183), .B(n678), .Z(n4268) );
  XOR \MIXCOLUMNS[3].d/U278  ( .A(n4088), .B(n4087), .Z(\w0[4][43] ) );
  XOR \MIXCOLUMNS[3].d/U277  ( .A(n4265), .B(n4268), .Z(n4087) );
  XOR \MIXCOLUMNS[3].d/U276  ( .A(n680), .B(n4261), .Z(n4088) );
  XOR \MIXCOLUMNS[3].d/U275  ( .A(n181), .B(n676), .Z(n4270) );
  XOR \MIXCOLUMNS[3].d/U274  ( .A(n4090), .B(n4089), .Z(\w0[4][44] ) );
  XOR \MIXCOLUMNS[3].d/U273  ( .A(n4267), .B(n4270), .Z(n4089) );
  XOR \MIXCOLUMNS[3].d/U272  ( .A(n678), .B(n4261), .Z(n4090) );
  XOR \MIXCOLUMNS[3].d/U271  ( .A(n179), .B(n674), .Z(n4272) );
  XOR \MIXCOLUMNS[3].d/U270  ( .A(n4272), .B(n4091), .Z(\w0[4][45] ) );
  XOR \MIXCOLUMNS[3].d/U269  ( .A(n676), .B(n4269), .Z(n4091) );
  XOR \MIXCOLUMNS[3].d/U268  ( .A(n177), .B(n672), .Z(n4274) );
  XOR \MIXCOLUMNS[3].d/U267  ( .A(n4093), .B(n4092), .Z(\w0[4][46] ) );
  XOR \MIXCOLUMNS[3].d/U266  ( .A(n4271), .B(n4274), .Z(n4092) );
  XOR \MIXCOLUMNS[3].d/U265  ( .A(n674), .B(n4261), .Z(n4093) );
  XOR \MIXCOLUMNS[3].d/U264  ( .A(n4273), .B(n4094), .Z(\w0[4][47] ) );
  XOR \MIXCOLUMNS[3].d/U263  ( .A(n672), .B(n4261), .Z(n4094) );
  XOR \MIXCOLUMNS[3].d/U262  ( .A(n4096), .B(n4095), .Z(\w0[4][48] ) );
  XOR \MIXCOLUMNS[3].d/U261  ( .A(n188), .B(n4261), .Z(n4095) );
  XOR \MIXCOLUMNS[3].d/U260  ( .A(n683), .B(n189), .Z(n4096) );
  XOR \MIXCOLUMNS[3].d/U259  ( .A(n4098), .B(n4097), .Z(\w0[4][49] ) );
  XOR \MIXCOLUMNS[3].d/U258  ( .A(\w3[3][42] ), .B(n4262), .Z(n4097) );
  XOR \MIXCOLUMNS[3].d/U257  ( .A(n681), .B(\w3[3][50] ), .Z(n4098) );
  XOR \MIXCOLUMNS[3].d/U256  ( .A(n4100), .B(n4099), .Z(\w0[4][50] ) );
  XOR \MIXCOLUMNS[3].d/U255  ( .A(n185), .B(n4264), .Z(n4099) );
  XOR \MIXCOLUMNS[3].d/U254  ( .A(\w3[3][58] ), .B(n186), .Z(n4100) );
  XOR \MIXCOLUMNS[3].d/U253  ( .A(n190), .B(n11), .Z(n4259) );
  XOR \MIXCOLUMNS[3].d/U252  ( .A(n4102), .B(n4101), .Z(\w0[4][51] ) );
  XOR \MIXCOLUMNS[3].d/U251  ( .A(n4266), .B(n4103), .Z(n4101) );
  XOR \MIXCOLUMNS[3].d/U250  ( .A(n183), .B(n4259), .Z(n4102) );
  XOR \MIXCOLUMNS[3].d/U249  ( .A(n679), .B(n184), .Z(n4103) );
  XOR \MIXCOLUMNS[3].d/U248  ( .A(n4105), .B(n4104), .Z(\w0[4][52] ) );
  XOR \MIXCOLUMNS[3].d/U247  ( .A(n4268), .B(n4106), .Z(n4104) );
  XOR \MIXCOLUMNS[3].d/U246  ( .A(n181), .B(n4259), .Z(n4105) );
  XOR \MIXCOLUMNS[3].d/U245  ( .A(n677), .B(n182), .Z(n4106) );
  XOR \MIXCOLUMNS[3].d/U244  ( .A(n4108), .B(n4107), .Z(\w0[4][53] ) );
  XOR \MIXCOLUMNS[3].d/U243  ( .A(n179), .B(n4270), .Z(n4107) );
  XOR \MIXCOLUMNS[3].d/U242  ( .A(n675), .B(n180), .Z(n4108) );
  XOR \MIXCOLUMNS[3].d/U241  ( .A(n4110), .B(n4109), .Z(\w0[4][54] ) );
  XOR \MIXCOLUMNS[3].d/U240  ( .A(n4272), .B(n4111), .Z(n4109) );
  XOR \MIXCOLUMNS[3].d/U239  ( .A(n177), .B(n4259), .Z(n4110) );
  XOR \MIXCOLUMNS[3].d/U238  ( .A(n673), .B(n178), .Z(n4111) );
  XOR \MIXCOLUMNS[3].d/U237  ( .A(n4274), .B(n4112), .Z(\w0[4][55] ) );
  XOR \MIXCOLUMNS[3].d/U236  ( .A(n671), .B(n4259), .Z(n4112) );
  XOR \MIXCOLUMNS[3].d/U235  ( .A(n4260), .B(n4113), .Z(\w0[4][56] ) );
  XOR \MIXCOLUMNS[3].d/U234  ( .A(n190), .B(n4261), .Z(n4113) );
  XOR \MIXCOLUMNS[3].d/U233  ( .A(n4262), .B(n4114), .Z(\w0[4][57] ) );
  XOR \MIXCOLUMNS[3].d/U232  ( .A(n189), .B(n4263), .Z(n4114) );
  XOR \MIXCOLUMNS[3].d/U231  ( .A(n4264), .B(n4115), .Z(\w0[4][58] ) );
  XOR \MIXCOLUMNS[3].d/U230  ( .A(\w3[3][50] ), .B(n4265), .Z(n4115) );
  XOR \MIXCOLUMNS[3].d/U229  ( .A(n4117), .B(n4116), .Z(\w0[4][59] ) );
  XOR \MIXCOLUMNS[3].d/U228  ( .A(n4267), .B(n4266), .Z(n4116) );
  XOR \MIXCOLUMNS[3].d/U227  ( .A(n186), .B(n4275), .Z(n4117) );
  XOR \MIXCOLUMNS[3].d/U226  ( .A(n4119), .B(n4118), .Z(\w0[4][60] ) );
  XOR \MIXCOLUMNS[3].d/U225  ( .A(n4269), .B(n4268), .Z(n4118) );
  XOR \MIXCOLUMNS[3].d/U224  ( .A(n184), .B(n4275), .Z(n4119) );
  XOR \MIXCOLUMNS[3].d/U223  ( .A(n4270), .B(n4120), .Z(\w0[4][61] ) );
  XOR \MIXCOLUMNS[3].d/U222  ( .A(n182), .B(n4271), .Z(n4120) );
  XOR \MIXCOLUMNS[3].d/U221  ( .A(n4122), .B(n4121), .Z(\w0[4][62] ) );
  XOR \MIXCOLUMNS[3].d/U220  ( .A(n4273), .B(n4272), .Z(n4121) );
  XOR \MIXCOLUMNS[3].d/U219  ( .A(n180), .B(n4275), .Z(n4122) );
  XOR \MIXCOLUMNS[3].d/U218  ( .A(n4274), .B(n4123), .Z(\w0[4][63] ) );
  XOR \MIXCOLUMNS[3].d/U217  ( .A(n178), .B(n4275), .Z(n4123) );
  XOR \MIXCOLUMNS[3].d/U216  ( .A(n670), .B(n176), .Z(n4293) );
  XOR \MIXCOLUMNS[3].d/U215  ( .A(n4125), .B(n4124), .Z(\w0[4][64] ) );
  XOR \MIXCOLUMNS[3].d/U214  ( .A(n669), .B(n4293), .Z(n4124) );
  XOR \MIXCOLUMNS[3].d/U213  ( .A(n668), .B(n10), .Z(n4125) );
  XOR \MIXCOLUMNS[3].d/U212  ( .A(n668), .B(n175), .Z(n4278) );
  XOR \MIXCOLUMNS[3].d/U211  ( .A(n4127), .B(n4126), .Z(\w0[4][65] ) );
  XOR \MIXCOLUMNS[3].d/U210  ( .A(\w3[3][66] ), .B(n4278), .Z(n4126) );
  XOR \MIXCOLUMNS[3].d/U209  ( .A(\w3[3][90] ), .B(n174), .Z(n4127) );
  XOR \MIXCOLUMNS[3].d/U208  ( .A(\w3[3][90] ), .B(\w3[3][82] ), .Z(n4281) );
  XOR \MIXCOLUMNS[3].d/U207  ( .A(n4129), .B(n4128), .Z(\w0[4][66] ) );
  XOR \MIXCOLUMNS[3].d/U206  ( .A(n667), .B(n4281), .Z(n4128) );
  XOR \MIXCOLUMNS[3].d/U205  ( .A(n666), .B(\w3[3][74] ), .Z(n4129) );
  XOR \MIXCOLUMNS[3].d/U204  ( .A(n670), .B(n173), .Z(n4276) );
  XOR \MIXCOLUMNS[3].d/U203  ( .A(n666), .B(n172), .Z(n4283) );
  XOR \MIXCOLUMNS[3].d/U202  ( .A(n4131), .B(n4130), .Z(\w0[4][67] ) );
  XOR \MIXCOLUMNS[3].d/U201  ( .A(n4283), .B(n4132), .Z(n4130) );
  XOR \MIXCOLUMNS[3].d/U200  ( .A(n665), .B(n4276), .Z(n4131) );
  XOR \MIXCOLUMNS[3].d/U199  ( .A(n664), .B(n171), .Z(n4132) );
  XOR \MIXCOLUMNS[3].d/U198  ( .A(n664), .B(n170), .Z(n4285) );
  XOR \MIXCOLUMNS[3].d/U197  ( .A(n4134), .B(n4133), .Z(\w0[4][68] ) );
  XOR \MIXCOLUMNS[3].d/U196  ( .A(n4285), .B(n4135), .Z(n4133) );
  XOR \MIXCOLUMNS[3].d/U195  ( .A(n663), .B(n4276), .Z(n4134) );
  XOR \MIXCOLUMNS[3].d/U194  ( .A(n662), .B(n169), .Z(n4135) );
  XOR \MIXCOLUMNS[3].d/U193  ( .A(n662), .B(n168), .Z(n4287) );
  XOR \MIXCOLUMNS[3].d/U192  ( .A(n4137), .B(n4136), .Z(\w0[4][69] ) );
  XOR \MIXCOLUMNS[3].d/U191  ( .A(n661), .B(n4287), .Z(n4136) );
  XOR \MIXCOLUMNS[3].d/U190  ( .A(n660), .B(n167), .Z(n4137) );
  XOR \MIXCOLUMNS[3].d/U189  ( .A(n660), .B(n166), .Z(n4289) );
  XOR \MIXCOLUMNS[3].d/U188  ( .A(n4139), .B(n4138), .Z(\w0[4][70] ) );
  XOR \MIXCOLUMNS[3].d/U187  ( .A(n4289), .B(n4140), .Z(n4138) );
  XOR \MIXCOLUMNS[3].d/U186  ( .A(n659), .B(n4276), .Z(n4139) );
  XOR \MIXCOLUMNS[3].d/U185  ( .A(n658), .B(n165), .Z(n4140) );
  XOR \MIXCOLUMNS[3].d/U184  ( .A(n658), .B(n164), .Z(n4291) );
  XOR \MIXCOLUMNS[3].d/U183  ( .A(n4291), .B(n4141), .Z(\w0[4][71] ) );
  XOR \MIXCOLUMNS[3].d/U182  ( .A(n163), .B(n4276), .Z(n4141) );
  XOR \MIXCOLUMNS[3].d/U181  ( .A(n174), .B(n669), .Z(n4280) );
  XOR \MIXCOLUMNS[3].d/U180  ( .A(n4280), .B(n4142), .Z(\w0[4][72] ) );
  XOR \MIXCOLUMNS[3].d/U179  ( .A(n173), .B(n4293), .Z(n4142) );
  XOR \MIXCOLUMNS[3].d/U178  ( .A(\w3[3][74] ), .B(\w3[3][66] ), .Z(n4282) );
  XOR \MIXCOLUMNS[3].d/U177  ( .A(n4282), .B(n4143), .Z(\w0[4][73] ) );
  XOR \MIXCOLUMNS[3].d/U176  ( .A(n669), .B(n4278), .Z(n4143) );
  XOR \MIXCOLUMNS[3].d/U175  ( .A(n171), .B(n667), .Z(n4284) );
  XOR \MIXCOLUMNS[3].d/U174  ( .A(n4284), .B(n4144), .Z(\w0[4][74] ) );
  XOR \MIXCOLUMNS[3].d/U173  ( .A(\w3[3][66] ), .B(n4281), .Z(n4144) );
  XOR \MIXCOLUMNS[3].d/U172  ( .A(n10), .B(n173), .Z(n4279) );
  XOR \MIXCOLUMNS[3].d/U171  ( .A(n169), .B(n665), .Z(n4286) );
  XOR \MIXCOLUMNS[3].d/U170  ( .A(n4146), .B(n4145), .Z(\w0[4][75] ) );
  XOR \MIXCOLUMNS[3].d/U169  ( .A(n4283), .B(n4286), .Z(n4145) );
  XOR \MIXCOLUMNS[3].d/U168  ( .A(n667), .B(n4279), .Z(n4146) );
  XOR \MIXCOLUMNS[3].d/U167  ( .A(n167), .B(n663), .Z(n4288) );
  XOR \MIXCOLUMNS[3].d/U166  ( .A(n4148), .B(n4147), .Z(\w0[4][76] ) );
  XOR \MIXCOLUMNS[3].d/U165  ( .A(n4285), .B(n4288), .Z(n4147) );
  XOR \MIXCOLUMNS[3].d/U164  ( .A(n665), .B(n4279), .Z(n4148) );
  XOR \MIXCOLUMNS[3].d/U163  ( .A(n165), .B(n661), .Z(n4290) );
  XOR \MIXCOLUMNS[3].d/U162  ( .A(n4290), .B(n4149), .Z(\w0[4][77] ) );
  XOR \MIXCOLUMNS[3].d/U161  ( .A(n663), .B(n4287), .Z(n4149) );
  XOR \MIXCOLUMNS[3].d/U160  ( .A(n163), .B(n659), .Z(n4292) );
  XOR \MIXCOLUMNS[3].d/U159  ( .A(n4151), .B(n4150), .Z(\w0[4][78] ) );
  XOR \MIXCOLUMNS[3].d/U158  ( .A(n4289), .B(n4292), .Z(n4150) );
  XOR \MIXCOLUMNS[3].d/U157  ( .A(n661), .B(n4279), .Z(n4151) );
  XOR \MIXCOLUMNS[3].d/U156  ( .A(n4291), .B(n4152), .Z(\w0[4][79] ) );
  XOR \MIXCOLUMNS[3].d/U155  ( .A(n659), .B(n4279), .Z(n4152) );
  XOR \MIXCOLUMNS[3].d/U154  ( .A(n4154), .B(n4153), .Z(\w0[4][80] ) );
  XOR \MIXCOLUMNS[3].d/U153  ( .A(n174), .B(n4279), .Z(n4153) );
  XOR \MIXCOLUMNS[3].d/U152  ( .A(n670), .B(n175), .Z(n4154) );
  XOR \MIXCOLUMNS[3].d/U151  ( .A(n4156), .B(n4155), .Z(\w0[4][81] ) );
  XOR \MIXCOLUMNS[3].d/U150  ( .A(\w3[3][74] ), .B(n4280), .Z(n4155) );
  XOR \MIXCOLUMNS[3].d/U149  ( .A(n668), .B(\w3[3][82] ), .Z(n4156) );
  XOR \MIXCOLUMNS[3].d/U148  ( .A(n4158), .B(n4157), .Z(\w0[4][82] ) );
  XOR \MIXCOLUMNS[3].d/U147  ( .A(n171), .B(n4282), .Z(n4157) );
  XOR \MIXCOLUMNS[3].d/U146  ( .A(\w3[3][90] ), .B(n172), .Z(n4158) );
  XOR \MIXCOLUMNS[3].d/U145  ( .A(n176), .B(n10), .Z(n4277) );
  XOR \MIXCOLUMNS[3].d/U144  ( .A(n4160), .B(n4159), .Z(\w0[4][83] ) );
  XOR \MIXCOLUMNS[3].d/U143  ( .A(n4284), .B(n4161), .Z(n4159) );
  XOR \MIXCOLUMNS[3].d/U142  ( .A(n169), .B(n4277), .Z(n4160) );
  XOR \MIXCOLUMNS[3].d/U141  ( .A(n666), .B(n170), .Z(n4161) );
  XOR \MIXCOLUMNS[3].d/U140  ( .A(n4163), .B(n4162), .Z(\w0[4][84] ) );
  XOR \MIXCOLUMNS[3].d/U139  ( .A(n4286), .B(n4164), .Z(n4162) );
  XOR \MIXCOLUMNS[3].d/U138  ( .A(n167), .B(n4277), .Z(n4163) );
  XOR \MIXCOLUMNS[3].d/U137  ( .A(n664), .B(n168), .Z(n4164) );
  XOR \MIXCOLUMNS[3].d/U136  ( .A(n4166), .B(n4165), .Z(\w0[4][85] ) );
  XOR \MIXCOLUMNS[3].d/U135  ( .A(n165), .B(n4288), .Z(n4165) );
  XOR \MIXCOLUMNS[3].d/U134  ( .A(n662), .B(n166), .Z(n4166) );
  XOR \MIXCOLUMNS[3].d/U133  ( .A(n4168), .B(n4167), .Z(\w0[4][86] ) );
  XOR \MIXCOLUMNS[3].d/U132  ( .A(n4290), .B(n4169), .Z(n4167) );
  XOR \MIXCOLUMNS[3].d/U131  ( .A(n163), .B(n4277), .Z(n4168) );
  XOR \MIXCOLUMNS[3].d/U130  ( .A(n660), .B(n164), .Z(n4169) );
  XOR \MIXCOLUMNS[3].d/U129  ( .A(n4292), .B(n4170), .Z(\w0[4][87] ) );
  XOR \MIXCOLUMNS[3].d/U128  ( .A(n658), .B(n4277), .Z(n4170) );
  XOR \MIXCOLUMNS[3].d/U127  ( .A(n4278), .B(n4171), .Z(\w0[4][88] ) );
  XOR \MIXCOLUMNS[3].d/U126  ( .A(n176), .B(n4279), .Z(n4171) );
  XOR \MIXCOLUMNS[3].d/U125  ( .A(n4280), .B(n4172), .Z(\w0[4][89] ) );
  XOR \MIXCOLUMNS[3].d/U124  ( .A(n175), .B(n4281), .Z(n4172) );
  XOR \MIXCOLUMNS[3].d/U123  ( .A(n4282), .B(n4173), .Z(\w0[4][90] ) );
  XOR \MIXCOLUMNS[3].d/U122  ( .A(\w3[3][82] ), .B(n4283), .Z(n4173) );
  XOR \MIXCOLUMNS[3].d/U121  ( .A(n4175), .B(n4174), .Z(\w0[4][91] ) );
  XOR \MIXCOLUMNS[3].d/U120  ( .A(n4285), .B(n4284), .Z(n4174) );
  XOR \MIXCOLUMNS[3].d/U119  ( .A(n172), .B(n4293), .Z(n4175) );
  XOR \MIXCOLUMNS[3].d/U118  ( .A(n4177), .B(n4176), .Z(\w0[4][92] ) );
  XOR \MIXCOLUMNS[3].d/U117  ( .A(n4287), .B(n4286), .Z(n4176) );
  XOR \MIXCOLUMNS[3].d/U116  ( .A(n170), .B(n4293), .Z(n4177) );
  XOR \MIXCOLUMNS[3].d/U115  ( .A(n4288), .B(n4178), .Z(\w0[4][93] ) );
  XOR \MIXCOLUMNS[3].d/U114  ( .A(n168), .B(n4289), .Z(n4178) );
  XOR \MIXCOLUMNS[3].d/U113  ( .A(n4180), .B(n4179), .Z(\w0[4][94] ) );
  XOR \MIXCOLUMNS[3].d/U112  ( .A(n4291), .B(n4290), .Z(n4179) );
  XOR \MIXCOLUMNS[3].d/U111  ( .A(n166), .B(n4293), .Z(n4180) );
  XOR \MIXCOLUMNS[3].d/U110  ( .A(n4292), .B(n4181), .Z(\w0[4][95] ) );
  XOR \MIXCOLUMNS[3].d/U109  ( .A(n164), .B(n4293), .Z(n4181) );
  XOR \MIXCOLUMNS[3].d/U108  ( .A(n657), .B(n162), .Z(n4311) );
  XOR \MIXCOLUMNS[3].d/U107  ( .A(n4183), .B(n4182), .Z(\w0[4][96] ) );
  XOR \MIXCOLUMNS[3].d/U106  ( .A(n656), .B(n4311), .Z(n4182) );
  XOR \MIXCOLUMNS[3].d/U105  ( .A(n655), .B(n9), .Z(n4183) );
  XOR \MIXCOLUMNS[3].d/U104  ( .A(n655), .B(n161), .Z(n4296) );
  XOR \MIXCOLUMNS[3].d/U103  ( .A(n4185), .B(n4184), .Z(\w0[4][97] ) );
  XOR \MIXCOLUMNS[3].d/U102  ( .A(\w3[3][98] ), .B(n4296), .Z(n4184) );
  XOR \MIXCOLUMNS[3].d/U101  ( .A(\w3[3][122] ), .B(n160), .Z(n4185) );
  XOR \MIXCOLUMNS[3].d/U100  ( .A(\w3[3][122] ), .B(\w3[3][114] ), .Z(n4299)
         );
  XOR \MIXCOLUMNS[3].d/U99  ( .A(n4187), .B(n4186), .Z(\w0[4][98] ) );
  XOR \MIXCOLUMNS[3].d/U98  ( .A(n654), .B(n4299), .Z(n4186) );
  XOR \MIXCOLUMNS[3].d/U97  ( .A(n653), .B(\w3[3][106] ), .Z(n4187) );
  XOR \MIXCOLUMNS[3].d/U96  ( .A(n657), .B(n159), .Z(n4294) );
  XOR \MIXCOLUMNS[3].d/U95  ( .A(n653), .B(n158), .Z(n4301) );
  XOR \MIXCOLUMNS[3].d/U94  ( .A(n4189), .B(n4188), .Z(\w0[4][99] ) );
  XOR \MIXCOLUMNS[3].d/U93  ( .A(n4301), .B(n4190), .Z(n4188) );
  XOR \MIXCOLUMNS[3].d/U92  ( .A(n652), .B(n4294), .Z(n4189) );
  XOR \MIXCOLUMNS[3].d/U91  ( .A(n651), .B(n157), .Z(n4190) );
  XOR \MIXCOLUMNS[3].d/U90  ( .A(n651), .B(n156), .Z(n4303) );
  XOR \MIXCOLUMNS[3].d/U89  ( .A(n4192), .B(n4191), .Z(\w0[4][100] ) );
  XOR \MIXCOLUMNS[3].d/U88  ( .A(n4303), .B(n4193), .Z(n4191) );
  XOR \MIXCOLUMNS[3].d/U87  ( .A(n650), .B(n4294), .Z(n4192) );
  XOR \MIXCOLUMNS[3].d/U86  ( .A(n649), .B(n155), .Z(n4193) );
  XOR \MIXCOLUMNS[3].d/U85  ( .A(n649), .B(n154), .Z(n4305) );
  XOR \MIXCOLUMNS[3].d/U84  ( .A(n4195), .B(n4194), .Z(\w0[4][101] ) );
  XOR \MIXCOLUMNS[3].d/U83  ( .A(n648), .B(n4305), .Z(n4194) );
  XOR \MIXCOLUMNS[3].d/U82  ( .A(n647), .B(n153), .Z(n4195) );
  XOR \MIXCOLUMNS[3].d/U81  ( .A(n647), .B(n152), .Z(n4307) );
  XOR \MIXCOLUMNS[3].d/U80  ( .A(n4197), .B(n4196), .Z(\w0[4][102] ) );
  XOR \MIXCOLUMNS[3].d/U79  ( .A(n4307), .B(n4198), .Z(n4196) );
  XOR \MIXCOLUMNS[3].d/U78  ( .A(n646), .B(n4294), .Z(n4197) );
  XOR \MIXCOLUMNS[3].d/U77  ( .A(n645), .B(n151), .Z(n4198) );
  XOR \MIXCOLUMNS[3].d/U76  ( .A(n645), .B(n150), .Z(n4309) );
  XOR \MIXCOLUMNS[3].d/U75  ( .A(n4309), .B(n4199), .Z(\w0[4][103] ) );
  XOR \MIXCOLUMNS[3].d/U74  ( .A(n149), .B(n4294), .Z(n4199) );
  XOR \MIXCOLUMNS[3].d/U73  ( .A(n160), .B(n656), .Z(n4298) );
  XOR \MIXCOLUMNS[3].d/U72  ( .A(n4298), .B(n4200), .Z(\w0[4][104] ) );
  XOR \MIXCOLUMNS[3].d/U71  ( .A(n159), .B(n4311), .Z(n4200) );
  XOR \MIXCOLUMNS[3].d/U70  ( .A(\w3[3][106] ), .B(\w3[3][98] ), .Z(n4300) );
  XOR \MIXCOLUMNS[3].d/U69  ( .A(n4300), .B(n4201), .Z(\w0[4][105] ) );
  XOR \MIXCOLUMNS[3].d/U68  ( .A(n656), .B(n4296), .Z(n4201) );
  XOR \MIXCOLUMNS[3].d/U67  ( .A(n157), .B(n654), .Z(n4302) );
  XOR \MIXCOLUMNS[3].d/U66  ( .A(n4302), .B(n4202), .Z(\w0[4][106] ) );
  XOR \MIXCOLUMNS[3].d/U65  ( .A(\w3[3][98] ), .B(n4299), .Z(n4202) );
  XOR \MIXCOLUMNS[3].d/U64  ( .A(n9), .B(n159), .Z(n4297) );
  XOR \MIXCOLUMNS[3].d/U63  ( .A(n155), .B(n652), .Z(n4304) );
  XOR \MIXCOLUMNS[3].d/U62  ( .A(n4204), .B(n4203), .Z(\w0[4][107] ) );
  XOR \MIXCOLUMNS[3].d/U61  ( .A(n4301), .B(n4304), .Z(n4203) );
  XOR \MIXCOLUMNS[3].d/U60  ( .A(n654), .B(n4297), .Z(n4204) );
  XOR \MIXCOLUMNS[3].d/U59  ( .A(n153), .B(n650), .Z(n4306) );
  XOR \MIXCOLUMNS[3].d/U58  ( .A(n4206), .B(n4205), .Z(\w0[4][108] ) );
  XOR \MIXCOLUMNS[3].d/U57  ( .A(n4303), .B(n4306), .Z(n4205) );
  XOR \MIXCOLUMNS[3].d/U56  ( .A(n652), .B(n4297), .Z(n4206) );
  XOR \MIXCOLUMNS[3].d/U55  ( .A(n151), .B(n648), .Z(n4308) );
  XOR \MIXCOLUMNS[3].d/U54  ( .A(n4308), .B(n4207), .Z(\w0[4][109] ) );
  XOR \MIXCOLUMNS[3].d/U53  ( .A(n650), .B(n4305), .Z(n4207) );
  XOR \MIXCOLUMNS[3].d/U52  ( .A(n149), .B(n646), .Z(n4310) );
  XOR \MIXCOLUMNS[3].d/U51  ( .A(n4209), .B(n4208), .Z(\w0[4][110] ) );
  XOR \MIXCOLUMNS[3].d/U50  ( .A(n4307), .B(n4310), .Z(n4208) );
  XOR \MIXCOLUMNS[3].d/U49  ( .A(n648), .B(n4297), .Z(n4209) );
  XOR \MIXCOLUMNS[3].d/U48  ( .A(n4309), .B(n4210), .Z(\w0[4][111] ) );
  XOR \MIXCOLUMNS[3].d/U47  ( .A(n646), .B(n4297), .Z(n4210) );
  XOR \MIXCOLUMNS[3].d/U46  ( .A(n4212), .B(n4211), .Z(\w0[4][112] ) );
  XOR \MIXCOLUMNS[3].d/U45  ( .A(n160), .B(n4297), .Z(n4211) );
  XOR \MIXCOLUMNS[3].d/U44  ( .A(n657), .B(n161), .Z(n4212) );
  XOR \MIXCOLUMNS[3].d/U43  ( .A(n4214), .B(n4213), .Z(\w0[4][113] ) );
  XOR \MIXCOLUMNS[3].d/U42  ( .A(\w3[3][106] ), .B(n4298), .Z(n4213) );
  XOR \MIXCOLUMNS[3].d/U41  ( .A(n655), .B(\w3[3][114] ), .Z(n4214) );
  XOR \MIXCOLUMNS[3].d/U40  ( .A(n4216), .B(n4215), .Z(\w0[4][114] ) );
  XOR \MIXCOLUMNS[3].d/U39  ( .A(n157), .B(n4300), .Z(n4215) );
  XOR \MIXCOLUMNS[3].d/U38  ( .A(\w3[3][122] ), .B(n158), .Z(n4216) );
  XOR \MIXCOLUMNS[3].d/U37  ( .A(n162), .B(n9), .Z(n4295) );
  XOR \MIXCOLUMNS[3].d/U36  ( .A(n4218), .B(n4217), .Z(\w0[4][115] ) );
  XOR \MIXCOLUMNS[3].d/U35  ( .A(n4302), .B(n4219), .Z(n4217) );
  XOR \MIXCOLUMNS[3].d/U34  ( .A(n155), .B(n4295), .Z(n4218) );
  XOR \MIXCOLUMNS[3].d/U33  ( .A(n653), .B(n156), .Z(n4219) );
  XOR \MIXCOLUMNS[3].d/U32  ( .A(n4221), .B(n4220), .Z(\w0[4][116] ) );
  XOR \MIXCOLUMNS[3].d/U31  ( .A(n4304), .B(n4222), .Z(n4220) );
  XOR \MIXCOLUMNS[3].d/U30  ( .A(n153), .B(n4295), .Z(n4221) );
  XOR \MIXCOLUMNS[3].d/U29  ( .A(n651), .B(n154), .Z(n4222) );
  XOR \MIXCOLUMNS[3].d/U28  ( .A(n4224), .B(n4223), .Z(\w0[4][117] ) );
  XOR \MIXCOLUMNS[3].d/U27  ( .A(n151), .B(n4306), .Z(n4223) );
  XOR \MIXCOLUMNS[3].d/U26  ( .A(n649), .B(n152), .Z(n4224) );
  XOR \MIXCOLUMNS[3].d/U25  ( .A(n4226), .B(n4225), .Z(\w0[4][118] ) );
  XOR \MIXCOLUMNS[3].d/U24  ( .A(n4308), .B(n4227), .Z(n4225) );
  XOR \MIXCOLUMNS[3].d/U23  ( .A(n149), .B(n4295), .Z(n4226) );
  XOR \MIXCOLUMNS[3].d/U22  ( .A(n647), .B(n150), .Z(n4227) );
  XOR \MIXCOLUMNS[3].d/U21  ( .A(n4310), .B(n4228), .Z(\w0[4][119] ) );
  XOR \MIXCOLUMNS[3].d/U20  ( .A(n645), .B(n4295), .Z(n4228) );
  XOR \MIXCOLUMNS[3].d/U19  ( .A(n4296), .B(n4229), .Z(\w0[4][120] ) );
  XOR \MIXCOLUMNS[3].d/U18  ( .A(n162), .B(n4297), .Z(n4229) );
  XOR \MIXCOLUMNS[3].d/U17  ( .A(n4298), .B(n4230), .Z(\w0[4][121] ) );
  XOR \MIXCOLUMNS[3].d/U16  ( .A(n161), .B(n4299), .Z(n4230) );
  XOR \MIXCOLUMNS[3].d/U15  ( .A(n4300), .B(n4231), .Z(\w0[4][122] ) );
  XOR \MIXCOLUMNS[3].d/U14  ( .A(\w3[3][114] ), .B(n4301), .Z(n4231) );
  XOR \MIXCOLUMNS[3].d/U13  ( .A(n4233), .B(n4232), .Z(\w0[4][123] ) );
  XOR \MIXCOLUMNS[3].d/U12  ( .A(n4303), .B(n4302), .Z(n4232) );
  XOR \MIXCOLUMNS[3].d/U11  ( .A(n158), .B(n4311), .Z(n4233) );
  XOR \MIXCOLUMNS[3].d/U10  ( .A(n4235), .B(n4234), .Z(\w0[4][124] ) );
  XOR \MIXCOLUMNS[3].d/U9  ( .A(n4305), .B(n4304), .Z(n4234) );
  XOR \MIXCOLUMNS[3].d/U8  ( .A(n156), .B(n4311), .Z(n4235) );
  XOR \MIXCOLUMNS[3].d/U7  ( .A(n4306), .B(n4236), .Z(\w0[4][125] ) );
  XOR \MIXCOLUMNS[3].d/U6  ( .A(n154), .B(n4307), .Z(n4236) );
  XOR \MIXCOLUMNS[3].d/U5  ( .A(n4238), .B(n4237), .Z(\w0[4][126] ) );
  XOR \MIXCOLUMNS[3].d/U4  ( .A(n4309), .B(n4308), .Z(n4237) );
  XOR \MIXCOLUMNS[3].d/U3  ( .A(n152), .B(n4311), .Z(n4238) );
  XOR \MIXCOLUMNS[3].d/U2  ( .A(n4310), .B(n4239), .Z(\w0[4][127] ) );
  XOR \MIXCOLUMNS[3].d/U1  ( .A(n150), .B(n4311), .Z(n4239) );
  XOR \MIXCOLUMNS[2].d/U432  ( .A(n644), .B(n148), .Z(n3953) );
  XOR \MIXCOLUMNS[2].d/U431  ( .A(n3705), .B(n3704), .Z(\w0[3][0] ) );
  XOR \MIXCOLUMNS[2].d/U430  ( .A(n643), .B(n3953), .Z(n3704) );
  XOR \MIXCOLUMNS[2].d/U429  ( .A(n642), .B(n8), .Z(n3705) );
  XOR \MIXCOLUMNS[2].d/U428  ( .A(n642), .B(n147), .Z(n3938) );
  XOR \MIXCOLUMNS[2].d/U427  ( .A(n3707), .B(n3706), .Z(\w0[3][1] ) );
  XOR \MIXCOLUMNS[2].d/U426  ( .A(\w3[2][2] ), .B(n3938), .Z(n3706) );
  XOR \MIXCOLUMNS[2].d/U425  ( .A(\w3[2][26] ), .B(n146), .Z(n3707) );
  XOR \MIXCOLUMNS[2].d/U424  ( .A(\w3[2][26] ), .B(\w3[2][18] ), .Z(n3941) );
  XOR \MIXCOLUMNS[2].d/U423  ( .A(n3709), .B(n3708), .Z(\w0[3][2] ) );
  XOR \MIXCOLUMNS[2].d/U422  ( .A(n641), .B(n3941), .Z(n3708) );
  XOR \MIXCOLUMNS[2].d/U421  ( .A(n640), .B(\w3[2][10] ), .Z(n3709) );
  XOR \MIXCOLUMNS[2].d/U420  ( .A(n644), .B(n145), .Z(n3936) );
  XOR \MIXCOLUMNS[2].d/U419  ( .A(n640), .B(n144), .Z(n3943) );
  XOR \MIXCOLUMNS[2].d/U418  ( .A(n3711), .B(n3710), .Z(\w0[3][3] ) );
  XOR \MIXCOLUMNS[2].d/U417  ( .A(n3943), .B(n3712), .Z(n3710) );
  XOR \MIXCOLUMNS[2].d/U416  ( .A(n639), .B(n3936), .Z(n3711) );
  XOR \MIXCOLUMNS[2].d/U415  ( .A(n638), .B(n143), .Z(n3712) );
  XOR \MIXCOLUMNS[2].d/U414  ( .A(n638), .B(n142), .Z(n3945) );
  XOR \MIXCOLUMNS[2].d/U413  ( .A(n3714), .B(n3713), .Z(\w0[3][4] ) );
  XOR \MIXCOLUMNS[2].d/U412  ( .A(n3945), .B(n3715), .Z(n3713) );
  XOR \MIXCOLUMNS[2].d/U411  ( .A(n637), .B(n3936), .Z(n3714) );
  XOR \MIXCOLUMNS[2].d/U410  ( .A(n636), .B(n141), .Z(n3715) );
  XOR \MIXCOLUMNS[2].d/U409  ( .A(n636), .B(n140), .Z(n3947) );
  XOR \MIXCOLUMNS[2].d/U408  ( .A(n3717), .B(n3716), .Z(\w0[3][5] ) );
  XOR \MIXCOLUMNS[2].d/U407  ( .A(n635), .B(n3947), .Z(n3716) );
  XOR \MIXCOLUMNS[2].d/U406  ( .A(n634), .B(n139), .Z(n3717) );
  XOR \MIXCOLUMNS[2].d/U405  ( .A(n634), .B(n138), .Z(n3949) );
  XOR \MIXCOLUMNS[2].d/U404  ( .A(n3719), .B(n3718), .Z(\w0[3][6] ) );
  XOR \MIXCOLUMNS[2].d/U403  ( .A(n3949), .B(n3720), .Z(n3718) );
  XOR \MIXCOLUMNS[2].d/U402  ( .A(n633), .B(n3936), .Z(n3719) );
  XOR \MIXCOLUMNS[2].d/U401  ( .A(n632), .B(n137), .Z(n3720) );
  XOR \MIXCOLUMNS[2].d/U400  ( .A(n632), .B(n136), .Z(n3951) );
  XOR \MIXCOLUMNS[2].d/U399  ( .A(n3951), .B(n3721), .Z(\w0[3][7] ) );
  XOR \MIXCOLUMNS[2].d/U398  ( .A(n135), .B(n3936), .Z(n3721) );
  XOR \MIXCOLUMNS[2].d/U397  ( .A(n146), .B(n643), .Z(n3940) );
  XOR \MIXCOLUMNS[2].d/U396  ( .A(n3940), .B(n3722), .Z(\w0[3][8] ) );
  XOR \MIXCOLUMNS[2].d/U395  ( .A(n145), .B(n3953), .Z(n3722) );
  XOR \MIXCOLUMNS[2].d/U394  ( .A(\w3[2][10] ), .B(\w3[2][2] ), .Z(n3942) );
  XOR \MIXCOLUMNS[2].d/U393  ( .A(n3942), .B(n3723), .Z(\w0[3][9] ) );
  XOR \MIXCOLUMNS[2].d/U392  ( .A(n643), .B(n3938), .Z(n3723) );
  XOR \MIXCOLUMNS[2].d/U391  ( .A(n143), .B(n641), .Z(n3944) );
  XOR \MIXCOLUMNS[2].d/U390  ( .A(n3944), .B(n3724), .Z(\w0[3][10] ) );
  XOR \MIXCOLUMNS[2].d/U389  ( .A(\w3[2][2] ), .B(n3941), .Z(n3724) );
  XOR \MIXCOLUMNS[2].d/U388  ( .A(n8), .B(n145), .Z(n3939) );
  XOR \MIXCOLUMNS[2].d/U387  ( .A(n141), .B(n639), .Z(n3946) );
  XOR \MIXCOLUMNS[2].d/U386  ( .A(n3726), .B(n3725), .Z(\w0[3][11] ) );
  XOR \MIXCOLUMNS[2].d/U385  ( .A(n3943), .B(n3946), .Z(n3725) );
  XOR \MIXCOLUMNS[2].d/U384  ( .A(n641), .B(n3939), .Z(n3726) );
  XOR \MIXCOLUMNS[2].d/U383  ( .A(n139), .B(n637), .Z(n3948) );
  XOR \MIXCOLUMNS[2].d/U382  ( .A(n3728), .B(n3727), .Z(\w0[3][12] ) );
  XOR \MIXCOLUMNS[2].d/U381  ( .A(n3945), .B(n3948), .Z(n3727) );
  XOR \MIXCOLUMNS[2].d/U380  ( .A(n639), .B(n3939), .Z(n3728) );
  XOR \MIXCOLUMNS[2].d/U379  ( .A(n137), .B(n635), .Z(n3950) );
  XOR \MIXCOLUMNS[2].d/U378  ( .A(n3950), .B(n3729), .Z(\w0[3][13] ) );
  XOR \MIXCOLUMNS[2].d/U377  ( .A(n637), .B(n3947), .Z(n3729) );
  XOR \MIXCOLUMNS[2].d/U376  ( .A(n135), .B(n633), .Z(n3952) );
  XOR \MIXCOLUMNS[2].d/U375  ( .A(n3731), .B(n3730), .Z(\w0[3][14] ) );
  XOR \MIXCOLUMNS[2].d/U374  ( .A(n3949), .B(n3952), .Z(n3730) );
  XOR \MIXCOLUMNS[2].d/U373  ( .A(n635), .B(n3939), .Z(n3731) );
  XOR \MIXCOLUMNS[2].d/U372  ( .A(n3951), .B(n3732), .Z(\w0[3][15] ) );
  XOR \MIXCOLUMNS[2].d/U371  ( .A(n633), .B(n3939), .Z(n3732) );
  XOR \MIXCOLUMNS[2].d/U370  ( .A(n3734), .B(n3733), .Z(\w0[3][16] ) );
  XOR \MIXCOLUMNS[2].d/U369  ( .A(n146), .B(n3939), .Z(n3733) );
  XOR \MIXCOLUMNS[2].d/U368  ( .A(n644), .B(n147), .Z(n3734) );
  XOR \MIXCOLUMNS[2].d/U367  ( .A(n3736), .B(n3735), .Z(\w0[3][17] ) );
  XOR \MIXCOLUMNS[2].d/U366  ( .A(\w3[2][10] ), .B(n3940), .Z(n3735) );
  XOR \MIXCOLUMNS[2].d/U365  ( .A(n642), .B(\w3[2][18] ), .Z(n3736) );
  XOR \MIXCOLUMNS[2].d/U364  ( .A(n3738), .B(n3737), .Z(\w0[3][18] ) );
  XOR \MIXCOLUMNS[2].d/U363  ( .A(n143), .B(n3942), .Z(n3737) );
  XOR \MIXCOLUMNS[2].d/U362  ( .A(\w3[2][26] ), .B(n144), .Z(n3738) );
  XOR \MIXCOLUMNS[2].d/U361  ( .A(n148), .B(n8), .Z(n3937) );
  XOR \MIXCOLUMNS[2].d/U360  ( .A(n3740), .B(n3739), .Z(\w0[3][19] ) );
  XOR \MIXCOLUMNS[2].d/U359  ( .A(n3944), .B(n3741), .Z(n3739) );
  XOR \MIXCOLUMNS[2].d/U358  ( .A(n141), .B(n3937), .Z(n3740) );
  XOR \MIXCOLUMNS[2].d/U357  ( .A(n640), .B(n142), .Z(n3741) );
  XOR \MIXCOLUMNS[2].d/U356  ( .A(n3743), .B(n3742), .Z(\w0[3][20] ) );
  XOR \MIXCOLUMNS[2].d/U355  ( .A(n3946), .B(n3744), .Z(n3742) );
  XOR \MIXCOLUMNS[2].d/U354  ( .A(n139), .B(n3937), .Z(n3743) );
  XOR \MIXCOLUMNS[2].d/U353  ( .A(n638), .B(n140), .Z(n3744) );
  XOR \MIXCOLUMNS[2].d/U352  ( .A(n3746), .B(n3745), .Z(\w0[3][21] ) );
  XOR \MIXCOLUMNS[2].d/U351  ( .A(n137), .B(n3948), .Z(n3745) );
  XOR \MIXCOLUMNS[2].d/U350  ( .A(n636), .B(n138), .Z(n3746) );
  XOR \MIXCOLUMNS[2].d/U349  ( .A(n3748), .B(n3747), .Z(\w0[3][22] ) );
  XOR \MIXCOLUMNS[2].d/U348  ( .A(n3950), .B(n3749), .Z(n3747) );
  XOR \MIXCOLUMNS[2].d/U347  ( .A(n135), .B(n3937), .Z(n3748) );
  XOR \MIXCOLUMNS[2].d/U346  ( .A(n634), .B(n136), .Z(n3749) );
  XOR \MIXCOLUMNS[2].d/U345  ( .A(n3952), .B(n3750), .Z(\w0[3][23] ) );
  XOR \MIXCOLUMNS[2].d/U344  ( .A(n632), .B(n3937), .Z(n3750) );
  XOR \MIXCOLUMNS[2].d/U343  ( .A(n3938), .B(n3751), .Z(\w0[3][24] ) );
  XOR \MIXCOLUMNS[2].d/U342  ( .A(n148), .B(n3939), .Z(n3751) );
  XOR \MIXCOLUMNS[2].d/U341  ( .A(n3940), .B(n3752), .Z(\w0[3][25] ) );
  XOR \MIXCOLUMNS[2].d/U340  ( .A(n147), .B(n3941), .Z(n3752) );
  XOR \MIXCOLUMNS[2].d/U339  ( .A(n3942), .B(n3753), .Z(\w0[3][26] ) );
  XOR \MIXCOLUMNS[2].d/U338  ( .A(\w3[2][18] ), .B(n3943), .Z(n3753) );
  XOR \MIXCOLUMNS[2].d/U337  ( .A(n3755), .B(n3754), .Z(\w0[3][27] ) );
  XOR \MIXCOLUMNS[2].d/U336  ( .A(n3945), .B(n3944), .Z(n3754) );
  XOR \MIXCOLUMNS[2].d/U335  ( .A(n144), .B(n3953), .Z(n3755) );
  XOR \MIXCOLUMNS[2].d/U334  ( .A(n3757), .B(n3756), .Z(\w0[3][28] ) );
  XOR \MIXCOLUMNS[2].d/U333  ( .A(n3947), .B(n3946), .Z(n3756) );
  XOR \MIXCOLUMNS[2].d/U332  ( .A(n142), .B(n3953), .Z(n3757) );
  XOR \MIXCOLUMNS[2].d/U331  ( .A(n3948), .B(n3758), .Z(\w0[3][29] ) );
  XOR \MIXCOLUMNS[2].d/U330  ( .A(n140), .B(n3949), .Z(n3758) );
  XOR \MIXCOLUMNS[2].d/U329  ( .A(n3760), .B(n3759), .Z(\w0[3][30] ) );
  XOR \MIXCOLUMNS[2].d/U328  ( .A(n3951), .B(n3950), .Z(n3759) );
  XOR \MIXCOLUMNS[2].d/U327  ( .A(n138), .B(n3953), .Z(n3760) );
  XOR \MIXCOLUMNS[2].d/U326  ( .A(n3952), .B(n3761), .Z(\w0[3][31] ) );
  XOR \MIXCOLUMNS[2].d/U325  ( .A(n136), .B(n3953), .Z(n3761) );
  XOR \MIXCOLUMNS[2].d/U324  ( .A(n631), .B(n134), .Z(n3971) );
  XOR \MIXCOLUMNS[2].d/U323  ( .A(n3763), .B(n3762), .Z(\w0[3][32] ) );
  XOR \MIXCOLUMNS[2].d/U322  ( .A(n630), .B(n3971), .Z(n3762) );
  XOR \MIXCOLUMNS[2].d/U321  ( .A(n629), .B(n7), .Z(n3763) );
  XOR \MIXCOLUMNS[2].d/U320  ( .A(n629), .B(n133), .Z(n3956) );
  XOR \MIXCOLUMNS[2].d/U319  ( .A(n3765), .B(n3764), .Z(\w0[3][33] ) );
  XOR \MIXCOLUMNS[2].d/U318  ( .A(\w3[2][34] ), .B(n3956), .Z(n3764) );
  XOR \MIXCOLUMNS[2].d/U317  ( .A(\w3[2][58] ), .B(n132), .Z(n3765) );
  XOR \MIXCOLUMNS[2].d/U316  ( .A(\w3[2][58] ), .B(\w3[2][50] ), .Z(n3959) );
  XOR \MIXCOLUMNS[2].d/U315  ( .A(n3767), .B(n3766), .Z(\w0[3][34] ) );
  XOR \MIXCOLUMNS[2].d/U314  ( .A(n628), .B(n3959), .Z(n3766) );
  XOR \MIXCOLUMNS[2].d/U313  ( .A(n627), .B(\w3[2][42] ), .Z(n3767) );
  XOR \MIXCOLUMNS[2].d/U312  ( .A(n631), .B(n131), .Z(n3954) );
  XOR \MIXCOLUMNS[2].d/U311  ( .A(n627), .B(n130), .Z(n3961) );
  XOR \MIXCOLUMNS[2].d/U310  ( .A(n3769), .B(n3768), .Z(\w0[3][35] ) );
  XOR \MIXCOLUMNS[2].d/U309  ( .A(n3961), .B(n3770), .Z(n3768) );
  XOR \MIXCOLUMNS[2].d/U308  ( .A(n626), .B(n3954), .Z(n3769) );
  XOR \MIXCOLUMNS[2].d/U307  ( .A(n625), .B(n129), .Z(n3770) );
  XOR \MIXCOLUMNS[2].d/U306  ( .A(n625), .B(n128), .Z(n3963) );
  XOR \MIXCOLUMNS[2].d/U305  ( .A(n3772), .B(n3771), .Z(\w0[3][36] ) );
  XOR \MIXCOLUMNS[2].d/U304  ( .A(n3963), .B(n3773), .Z(n3771) );
  XOR \MIXCOLUMNS[2].d/U303  ( .A(n624), .B(n3954), .Z(n3772) );
  XOR \MIXCOLUMNS[2].d/U302  ( .A(n623), .B(n127), .Z(n3773) );
  XOR \MIXCOLUMNS[2].d/U301  ( .A(n623), .B(n126), .Z(n3965) );
  XOR \MIXCOLUMNS[2].d/U300  ( .A(n3775), .B(n3774), .Z(\w0[3][37] ) );
  XOR \MIXCOLUMNS[2].d/U299  ( .A(n622), .B(n3965), .Z(n3774) );
  XOR \MIXCOLUMNS[2].d/U298  ( .A(n621), .B(n125), .Z(n3775) );
  XOR \MIXCOLUMNS[2].d/U297  ( .A(n621), .B(n124), .Z(n3967) );
  XOR \MIXCOLUMNS[2].d/U296  ( .A(n3777), .B(n3776), .Z(\w0[3][38] ) );
  XOR \MIXCOLUMNS[2].d/U295  ( .A(n3967), .B(n3778), .Z(n3776) );
  XOR \MIXCOLUMNS[2].d/U294  ( .A(n620), .B(n3954), .Z(n3777) );
  XOR \MIXCOLUMNS[2].d/U293  ( .A(n619), .B(n123), .Z(n3778) );
  XOR \MIXCOLUMNS[2].d/U292  ( .A(n619), .B(n122), .Z(n3969) );
  XOR \MIXCOLUMNS[2].d/U291  ( .A(n3969), .B(n3779), .Z(\w0[3][39] ) );
  XOR \MIXCOLUMNS[2].d/U290  ( .A(n121), .B(n3954), .Z(n3779) );
  XOR \MIXCOLUMNS[2].d/U289  ( .A(n132), .B(n630), .Z(n3958) );
  XOR \MIXCOLUMNS[2].d/U288  ( .A(n3958), .B(n3780), .Z(\w0[3][40] ) );
  XOR \MIXCOLUMNS[2].d/U287  ( .A(n131), .B(n3971), .Z(n3780) );
  XOR \MIXCOLUMNS[2].d/U286  ( .A(\w3[2][42] ), .B(\w3[2][34] ), .Z(n3960) );
  XOR \MIXCOLUMNS[2].d/U285  ( .A(n3960), .B(n3781), .Z(\w0[3][41] ) );
  XOR \MIXCOLUMNS[2].d/U284  ( .A(n630), .B(n3956), .Z(n3781) );
  XOR \MIXCOLUMNS[2].d/U283  ( .A(n129), .B(n628), .Z(n3962) );
  XOR \MIXCOLUMNS[2].d/U282  ( .A(n3962), .B(n3782), .Z(\w0[3][42] ) );
  XOR \MIXCOLUMNS[2].d/U281  ( .A(\w3[2][34] ), .B(n3959), .Z(n3782) );
  XOR \MIXCOLUMNS[2].d/U280  ( .A(n7), .B(n131), .Z(n3957) );
  XOR \MIXCOLUMNS[2].d/U279  ( .A(n127), .B(n626), .Z(n3964) );
  XOR \MIXCOLUMNS[2].d/U278  ( .A(n3784), .B(n3783), .Z(\w0[3][43] ) );
  XOR \MIXCOLUMNS[2].d/U277  ( .A(n3961), .B(n3964), .Z(n3783) );
  XOR \MIXCOLUMNS[2].d/U276  ( .A(n628), .B(n3957), .Z(n3784) );
  XOR \MIXCOLUMNS[2].d/U275  ( .A(n125), .B(n624), .Z(n3966) );
  XOR \MIXCOLUMNS[2].d/U274  ( .A(n3786), .B(n3785), .Z(\w0[3][44] ) );
  XOR \MIXCOLUMNS[2].d/U273  ( .A(n3963), .B(n3966), .Z(n3785) );
  XOR \MIXCOLUMNS[2].d/U272  ( .A(n626), .B(n3957), .Z(n3786) );
  XOR \MIXCOLUMNS[2].d/U271  ( .A(n123), .B(n622), .Z(n3968) );
  XOR \MIXCOLUMNS[2].d/U270  ( .A(n3968), .B(n3787), .Z(\w0[3][45] ) );
  XOR \MIXCOLUMNS[2].d/U269  ( .A(n624), .B(n3965), .Z(n3787) );
  XOR \MIXCOLUMNS[2].d/U268  ( .A(n121), .B(n620), .Z(n3970) );
  XOR \MIXCOLUMNS[2].d/U267  ( .A(n3789), .B(n3788), .Z(\w0[3][46] ) );
  XOR \MIXCOLUMNS[2].d/U266  ( .A(n3967), .B(n3970), .Z(n3788) );
  XOR \MIXCOLUMNS[2].d/U265  ( .A(n622), .B(n3957), .Z(n3789) );
  XOR \MIXCOLUMNS[2].d/U264  ( .A(n3969), .B(n3790), .Z(\w0[3][47] ) );
  XOR \MIXCOLUMNS[2].d/U263  ( .A(n620), .B(n3957), .Z(n3790) );
  XOR \MIXCOLUMNS[2].d/U262  ( .A(n3792), .B(n3791), .Z(\w0[3][48] ) );
  XOR \MIXCOLUMNS[2].d/U261  ( .A(n132), .B(n3957), .Z(n3791) );
  XOR \MIXCOLUMNS[2].d/U260  ( .A(n631), .B(n133), .Z(n3792) );
  XOR \MIXCOLUMNS[2].d/U259  ( .A(n3794), .B(n3793), .Z(\w0[3][49] ) );
  XOR \MIXCOLUMNS[2].d/U258  ( .A(\w3[2][42] ), .B(n3958), .Z(n3793) );
  XOR \MIXCOLUMNS[2].d/U257  ( .A(n629), .B(\w3[2][50] ), .Z(n3794) );
  XOR \MIXCOLUMNS[2].d/U256  ( .A(n3796), .B(n3795), .Z(\w0[3][50] ) );
  XOR \MIXCOLUMNS[2].d/U255  ( .A(n129), .B(n3960), .Z(n3795) );
  XOR \MIXCOLUMNS[2].d/U254  ( .A(\w3[2][58] ), .B(n130), .Z(n3796) );
  XOR \MIXCOLUMNS[2].d/U253  ( .A(n134), .B(n7), .Z(n3955) );
  XOR \MIXCOLUMNS[2].d/U252  ( .A(n3798), .B(n3797), .Z(\w0[3][51] ) );
  XOR \MIXCOLUMNS[2].d/U251  ( .A(n3962), .B(n3799), .Z(n3797) );
  XOR \MIXCOLUMNS[2].d/U250  ( .A(n127), .B(n3955), .Z(n3798) );
  XOR \MIXCOLUMNS[2].d/U249  ( .A(n627), .B(n128), .Z(n3799) );
  XOR \MIXCOLUMNS[2].d/U248  ( .A(n3801), .B(n3800), .Z(\w0[3][52] ) );
  XOR \MIXCOLUMNS[2].d/U247  ( .A(n3964), .B(n3802), .Z(n3800) );
  XOR \MIXCOLUMNS[2].d/U246  ( .A(n125), .B(n3955), .Z(n3801) );
  XOR \MIXCOLUMNS[2].d/U245  ( .A(n625), .B(n126), .Z(n3802) );
  XOR \MIXCOLUMNS[2].d/U244  ( .A(n3804), .B(n3803), .Z(\w0[3][53] ) );
  XOR \MIXCOLUMNS[2].d/U243  ( .A(n123), .B(n3966), .Z(n3803) );
  XOR \MIXCOLUMNS[2].d/U242  ( .A(n623), .B(n124), .Z(n3804) );
  XOR \MIXCOLUMNS[2].d/U241  ( .A(n3806), .B(n3805), .Z(\w0[3][54] ) );
  XOR \MIXCOLUMNS[2].d/U240  ( .A(n3968), .B(n3807), .Z(n3805) );
  XOR \MIXCOLUMNS[2].d/U239  ( .A(n121), .B(n3955), .Z(n3806) );
  XOR \MIXCOLUMNS[2].d/U238  ( .A(n621), .B(n122), .Z(n3807) );
  XOR \MIXCOLUMNS[2].d/U237  ( .A(n3970), .B(n3808), .Z(\w0[3][55] ) );
  XOR \MIXCOLUMNS[2].d/U236  ( .A(n619), .B(n3955), .Z(n3808) );
  XOR \MIXCOLUMNS[2].d/U235  ( .A(n3956), .B(n3809), .Z(\w0[3][56] ) );
  XOR \MIXCOLUMNS[2].d/U234  ( .A(n134), .B(n3957), .Z(n3809) );
  XOR \MIXCOLUMNS[2].d/U233  ( .A(n3958), .B(n3810), .Z(\w0[3][57] ) );
  XOR \MIXCOLUMNS[2].d/U232  ( .A(n133), .B(n3959), .Z(n3810) );
  XOR \MIXCOLUMNS[2].d/U231  ( .A(n3960), .B(n3811), .Z(\w0[3][58] ) );
  XOR \MIXCOLUMNS[2].d/U230  ( .A(\w3[2][50] ), .B(n3961), .Z(n3811) );
  XOR \MIXCOLUMNS[2].d/U229  ( .A(n3813), .B(n3812), .Z(\w0[3][59] ) );
  XOR \MIXCOLUMNS[2].d/U228  ( .A(n3963), .B(n3962), .Z(n3812) );
  XOR \MIXCOLUMNS[2].d/U227  ( .A(n130), .B(n3971), .Z(n3813) );
  XOR \MIXCOLUMNS[2].d/U226  ( .A(n3815), .B(n3814), .Z(\w0[3][60] ) );
  XOR \MIXCOLUMNS[2].d/U225  ( .A(n3965), .B(n3964), .Z(n3814) );
  XOR \MIXCOLUMNS[2].d/U224  ( .A(n128), .B(n3971), .Z(n3815) );
  XOR \MIXCOLUMNS[2].d/U223  ( .A(n3966), .B(n3816), .Z(\w0[3][61] ) );
  XOR \MIXCOLUMNS[2].d/U222  ( .A(n126), .B(n3967), .Z(n3816) );
  XOR \MIXCOLUMNS[2].d/U221  ( .A(n3818), .B(n3817), .Z(\w0[3][62] ) );
  XOR \MIXCOLUMNS[2].d/U220  ( .A(n3969), .B(n3968), .Z(n3817) );
  XOR \MIXCOLUMNS[2].d/U219  ( .A(n124), .B(n3971), .Z(n3818) );
  XOR \MIXCOLUMNS[2].d/U218  ( .A(n3970), .B(n3819), .Z(\w0[3][63] ) );
  XOR \MIXCOLUMNS[2].d/U217  ( .A(n122), .B(n3971), .Z(n3819) );
  XOR \MIXCOLUMNS[2].d/U216  ( .A(n618), .B(n120), .Z(n3989) );
  XOR \MIXCOLUMNS[2].d/U215  ( .A(n3821), .B(n3820), .Z(\w0[3][64] ) );
  XOR \MIXCOLUMNS[2].d/U214  ( .A(n617), .B(n3989), .Z(n3820) );
  XOR \MIXCOLUMNS[2].d/U213  ( .A(n616), .B(n6), .Z(n3821) );
  XOR \MIXCOLUMNS[2].d/U212  ( .A(n616), .B(n119), .Z(n3974) );
  XOR \MIXCOLUMNS[2].d/U211  ( .A(n3823), .B(n3822), .Z(\w0[3][65] ) );
  XOR \MIXCOLUMNS[2].d/U210  ( .A(\w3[2][66] ), .B(n3974), .Z(n3822) );
  XOR \MIXCOLUMNS[2].d/U209  ( .A(\w3[2][90] ), .B(n118), .Z(n3823) );
  XOR \MIXCOLUMNS[2].d/U208  ( .A(\w3[2][90] ), .B(\w3[2][82] ), .Z(n3977) );
  XOR \MIXCOLUMNS[2].d/U207  ( .A(n3825), .B(n3824), .Z(\w0[3][66] ) );
  XOR \MIXCOLUMNS[2].d/U206  ( .A(n615), .B(n3977), .Z(n3824) );
  XOR \MIXCOLUMNS[2].d/U205  ( .A(n614), .B(\w3[2][74] ), .Z(n3825) );
  XOR \MIXCOLUMNS[2].d/U204  ( .A(n618), .B(n117), .Z(n3972) );
  XOR \MIXCOLUMNS[2].d/U203  ( .A(n614), .B(n116), .Z(n3979) );
  XOR \MIXCOLUMNS[2].d/U202  ( .A(n3827), .B(n3826), .Z(\w0[3][67] ) );
  XOR \MIXCOLUMNS[2].d/U201  ( .A(n3979), .B(n3828), .Z(n3826) );
  XOR \MIXCOLUMNS[2].d/U200  ( .A(n613), .B(n3972), .Z(n3827) );
  XOR \MIXCOLUMNS[2].d/U199  ( .A(n612), .B(n115), .Z(n3828) );
  XOR \MIXCOLUMNS[2].d/U198  ( .A(n612), .B(n114), .Z(n3981) );
  XOR \MIXCOLUMNS[2].d/U197  ( .A(n3830), .B(n3829), .Z(\w0[3][68] ) );
  XOR \MIXCOLUMNS[2].d/U196  ( .A(n3981), .B(n3831), .Z(n3829) );
  XOR \MIXCOLUMNS[2].d/U195  ( .A(n611), .B(n3972), .Z(n3830) );
  XOR \MIXCOLUMNS[2].d/U194  ( .A(n610), .B(n113), .Z(n3831) );
  XOR \MIXCOLUMNS[2].d/U193  ( .A(n610), .B(n112), .Z(n3983) );
  XOR \MIXCOLUMNS[2].d/U192  ( .A(n3833), .B(n3832), .Z(\w0[3][69] ) );
  XOR \MIXCOLUMNS[2].d/U191  ( .A(n609), .B(n3983), .Z(n3832) );
  XOR \MIXCOLUMNS[2].d/U190  ( .A(n608), .B(n111), .Z(n3833) );
  XOR \MIXCOLUMNS[2].d/U189  ( .A(n608), .B(n110), .Z(n3985) );
  XOR \MIXCOLUMNS[2].d/U188  ( .A(n3835), .B(n3834), .Z(\w0[3][70] ) );
  XOR \MIXCOLUMNS[2].d/U187  ( .A(n3985), .B(n3836), .Z(n3834) );
  XOR \MIXCOLUMNS[2].d/U186  ( .A(n607), .B(n3972), .Z(n3835) );
  XOR \MIXCOLUMNS[2].d/U185  ( .A(n606), .B(n109), .Z(n3836) );
  XOR \MIXCOLUMNS[2].d/U184  ( .A(n606), .B(n108), .Z(n3987) );
  XOR \MIXCOLUMNS[2].d/U183  ( .A(n3987), .B(n3837), .Z(\w0[3][71] ) );
  XOR \MIXCOLUMNS[2].d/U182  ( .A(n107), .B(n3972), .Z(n3837) );
  XOR \MIXCOLUMNS[2].d/U181  ( .A(n118), .B(n617), .Z(n3976) );
  XOR \MIXCOLUMNS[2].d/U180  ( .A(n3976), .B(n3838), .Z(\w0[3][72] ) );
  XOR \MIXCOLUMNS[2].d/U179  ( .A(n117), .B(n3989), .Z(n3838) );
  XOR \MIXCOLUMNS[2].d/U178  ( .A(\w3[2][74] ), .B(\w3[2][66] ), .Z(n3978) );
  XOR \MIXCOLUMNS[2].d/U177  ( .A(n3978), .B(n3839), .Z(\w0[3][73] ) );
  XOR \MIXCOLUMNS[2].d/U176  ( .A(n617), .B(n3974), .Z(n3839) );
  XOR \MIXCOLUMNS[2].d/U175  ( .A(n115), .B(n615), .Z(n3980) );
  XOR \MIXCOLUMNS[2].d/U174  ( .A(n3980), .B(n3840), .Z(\w0[3][74] ) );
  XOR \MIXCOLUMNS[2].d/U173  ( .A(\w3[2][66] ), .B(n3977), .Z(n3840) );
  XOR \MIXCOLUMNS[2].d/U172  ( .A(n6), .B(n117), .Z(n3975) );
  XOR \MIXCOLUMNS[2].d/U171  ( .A(n113), .B(n613), .Z(n3982) );
  XOR \MIXCOLUMNS[2].d/U170  ( .A(n3842), .B(n3841), .Z(\w0[3][75] ) );
  XOR \MIXCOLUMNS[2].d/U169  ( .A(n3979), .B(n3982), .Z(n3841) );
  XOR \MIXCOLUMNS[2].d/U168  ( .A(n615), .B(n3975), .Z(n3842) );
  XOR \MIXCOLUMNS[2].d/U167  ( .A(n111), .B(n611), .Z(n3984) );
  XOR \MIXCOLUMNS[2].d/U166  ( .A(n3844), .B(n3843), .Z(\w0[3][76] ) );
  XOR \MIXCOLUMNS[2].d/U165  ( .A(n3981), .B(n3984), .Z(n3843) );
  XOR \MIXCOLUMNS[2].d/U164  ( .A(n613), .B(n3975), .Z(n3844) );
  XOR \MIXCOLUMNS[2].d/U163  ( .A(n109), .B(n609), .Z(n3986) );
  XOR \MIXCOLUMNS[2].d/U162  ( .A(n3986), .B(n3845), .Z(\w0[3][77] ) );
  XOR \MIXCOLUMNS[2].d/U161  ( .A(n611), .B(n3983), .Z(n3845) );
  XOR \MIXCOLUMNS[2].d/U160  ( .A(n107), .B(n607), .Z(n3988) );
  XOR \MIXCOLUMNS[2].d/U159  ( .A(n3847), .B(n3846), .Z(\w0[3][78] ) );
  XOR \MIXCOLUMNS[2].d/U158  ( .A(n3985), .B(n3988), .Z(n3846) );
  XOR \MIXCOLUMNS[2].d/U157  ( .A(n609), .B(n3975), .Z(n3847) );
  XOR \MIXCOLUMNS[2].d/U156  ( .A(n3987), .B(n3848), .Z(\w0[3][79] ) );
  XOR \MIXCOLUMNS[2].d/U155  ( .A(n607), .B(n3975), .Z(n3848) );
  XOR \MIXCOLUMNS[2].d/U154  ( .A(n3850), .B(n3849), .Z(\w0[3][80] ) );
  XOR \MIXCOLUMNS[2].d/U153  ( .A(n118), .B(n3975), .Z(n3849) );
  XOR \MIXCOLUMNS[2].d/U152  ( .A(n618), .B(n119), .Z(n3850) );
  XOR \MIXCOLUMNS[2].d/U151  ( .A(n3852), .B(n3851), .Z(\w0[3][81] ) );
  XOR \MIXCOLUMNS[2].d/U150  ( .A(\w3[2][74] ), .B(n3976), .Z(n3851) );
  XOR \MIXCOLUMNS[2].d/U149  ( .A(n616), .B(\w3[2][82] ), .Z(n3852) );
  XOR \MIXCOLUMNS[2].d/U148  ( .A(n3854), .B(n3853), .Z(\w0[3][82] ) );
  XOR \MIXCOLUMNS[2].d/U147  ( .A(n115), .B(n3978), .Z(n3853) );
  XOR \MIXCOLUMNS[2].d/U146  ( .A(\w3[2][90] ), .B(n116), .Z(n3854) );
  XOR \MIXCOLUMNS[2].d/U145  ( .A(n120), .B(n6), .Z(n3973) );
  XOR \MIXCOLUMNS[2].d/U144  ( .A(n3856), .B(n3855), .Z(\w0[3][83] ) );
  XOR \MIXCOLUMNS[2].d/U143  ( .A(n3980), .B(n3857), .Z(n3855) );
  XOR \MIXCOLUMNS[2].d/U142  ( .A(n113), .B(n3973), .Z(n3856) );
  XOR \MIXCOLUMNS[2].d/U141  ( .A(n614), .B(n114), .Z(n3857) );
  XOR \MIXCOLUMNS[2].d/U140  ( .A(n3859), .B(n3858), .Z(\w0[3][84] ) );
  XOR \MIXCOLUMNS[2].d/U139  ( .A(n3982), .B(n3860), .Z(n3858) );
  XOR \MIXCOLUMNS[2].d/U138  ( .A(n111), .B(n3973), .Z(n3859) );
  XOR \MIXCOLUMNS[2].d/U137  ( .A(n612), .B(n112), .Z(n3860) );
  XOR \MIXCOLUMNS[2].d/U136  ( .A(n3862), .B(n3861), .Z(\w0[3][85] ) );
  XOR \MIXCOLUMNS[2].d/U135  ( .A(n109), .B(n3984), .Z(n3861) );
  XOR \MIXCOLUMNS[2].d/U134  ( .A(n610), .B(n110), .Z(n3862) );
  XOR \MIXCOLUMNS[2].d/U133  ( .A(n3864), .B(n3863), .Z(\w0[3][86] ) );
  XOR \MIXCOLUMNS[2].d/U132  ( .A(n3986), .B(n3865), .Z(n3863) );
  XOR \MIXCOLUMNS[2].d/U131  ( .A(n107), .B(n3973), .Z(n3864) );
  XOR \MIXCOLUMNS[2].d/U130  ( .A(n608), .B(n108), .Z(n3865) );
  XOR \MIXCOLUMNS[2].d/U129  ( .A(n3988), .B(n3866), .Z(\w0[3][87] ) );
  XOR \MIXCOLUMNS[2].d/U128  ( .A(n606), .B(n3973), .Z(n3866) );
  XOR \MIXCOLUMNS[2].d/U127  ( .A(n3974), .B(n3867), .Z(\w0[3][88] ) );
  XOR \MIXCOLUMNS[2].d/U126  ( .A(n120), .B(n3975), .Z(n3867) );
  XOR \MIXCOLUMNS[2].d/U125  ( .A(n3976), .B(n3868), .Z(\w0[3][89] ) );
  XOR \MIXCOLUMNS[2].d/U124  ( .A(n119), .B(n3977), .Z(n3868) );
  XOR \MIXCOLUMNS[2].d/U123  ( .A(n3978), .B(n3869), .Z(\w0[3][90] ) );
  XOR \MIXCOLUMNS[2].d/U122  ( .A(\w3[2][82] ), .B(n3979), .Z(n3869) );
  XOR \MIXCOLUMNS[2].d/U121  ( .A(n3871), .B(n3870), .Z(\w0[3][91] ) );
  XOR \MIXCOLUMNS[2].d/U120  ( .A(n3981), .B(n3980), .Z(n3870) );
  XOR \MIXCOLUMNS[2].d/U119  ( .A(n116), .B(n3989), .Z(n3871) );
  XOR \MIXCOLUMNS[2].d/U118  ( .A(n3873), .B(n3872), .Z(\w0[3][92] ) );
  XOR \MIXCOLUMNS[2].d/U117  ( .A(n3983), .B(n3982), .Z(n3872) );
  XOR \MIXCOLUMNS[2].d/U116  ( .A(n114), .B(n3989), .Z(n3873) );
  XOR \MIXCOLUMNS[2].d/U115  ( .A(n3984), .B(n3874), .Z(\w0[3][93] ) );
  XOR \MIXCOLUMNS[2].d/U114  ( .A(n112), .B(n3985), .Z(n3874) );
  XOR \MIXCOLUMNS[2].d/U113  ( .A(n3876), .B(n3875), .Z(\w0[3][94] ) );
  XOR \MIXCOLUMNS[2].d/U112  ( .A(n3987), .B(n3986), .Z(n3875) );
  XOR \MIXCOLUMNS[2].d/U111  ( .A(n110), .B(n3989), .Z(n3876) );
  XOR \MIXCOLUMNS[2].d/U110  ( .A(n3988), .B(n3877), .Z(\w0[3][95] ) );
  XOR \MIXCOLUMNS[2].d/U109  ( .A(n108), .B(n3989), .Z(n3877) );
  XOR \MIXCOLUMNS[2].d/U108  ( .A(n605), .B(n106), .Z(n4007) );
  XOR \MIXCOLUMNS[2].d/U107  ( .A(n3879), .B(n3878), .Z(\w0[3][96] ) );
  XOR \MIXCOLUMNS[2].d/U106  ( .A(n604), .B(n4007), .Z(n3878) );
  XOR \MIXCOLUMNS[2].d/U105  ( .A(n603), .B(n5), .Z(n3879) );
  XOR \MIXCOLUMNS[2].d/U104  ( .A(n603), .B(n105), .Z(n3992) );
  XOR \MIXCOLUMNS[2].d/U103  ( .A(n3881), .B(n3880), .Z(\w0[3][97] ) );
  XOR \MIXCOLUMNS[2].d/U102  ( .A(\w3[2][98] ), .B(n3992), .Z(n3880) );
  XOR \MIXCOLUMNS[2].d/U101  ( .A(\w3[2][122] ), .B(n104), .Z(n3881) );
  XOR \MIXCOLUMNS[2].d/U100  ( .A(\w3[2][122] ), .B(\w3[2][114] ), .Z(n3995)
         );
  XOR \MIXCOLUMNS[2].d/U99  ( .A(n3883), .B(n3882), .Z(\w0[3][98] ) );
  XOR \MIXCOLUMNS[2].d/U98  ( .A(n602), .B(n3995), .Z(n3882) );
  XOR \MIXCOLUMNS[2].d/U97  ( .A(n601), .B(\w3[2][106] ), .Z(n3883) );
  XOR \MIXCOLUMNS[2].d/U96  ( .A(n605), .B(n103), .Z(n3990) );
  XOR \MIXCOLUMNS[2].d/U95  ( .A(n601), .B(n102), .Z(n3997) );
  XOR \MIXCOLUMNS[2].d/U94  ( .A(n3885), .B(n3884), .Z(\w0[3][99] ) );
  XOR \MIXCOLUMNS[2].d/U93  ( .A(n3997), .B(n3886), .Z(n3884) );
  XOR \MIXCOLUMNS[2].d/U92  ( .A(n600), .B(n3990), .Z(n3885) );
  XOR \MIXCOLUMNS[2].d/U91  ( .A(n599), .B(n101), .Z(n3886) );
  XOR \MIXCOLUMNS[2].d/U90  ( .A(n599), .B(n100), .Z(n3999) );
  XOR \MIXCOLUMNS[2].d/U89  ( .A(n3888), .B(n3887), .Z(\w0[3][100] ) );
  XOR \MIXCOLUMNS[2].d/U88  ( .A(n3999), .B(n3889), .Z(n3887) );
  XOR \MIXCOLUMNS[2].d/U87  ( .A(n598), .B(n3990), .Z(n3888) );
  XOR \MIXCOLUMNS[2].d/U86  ( .A(n597), .B(n99), .Z(n3889) );
  XOR \MIXCOLUMNS[2].d/U85  ( .A(n597), .B(n98), .Z(n4001) );
  XOR \MIXCOLUMNS[2].d/U84  ( .A(n3891), .B(n3890), .Z(\w0[3][101] ) );
  XOR \MIXCOLUMNS[2].d/U83  ( .A(n596), .B(n4001), .Z(n3890) );
  XOR \MIXCOLUMNS[2].d/U82  ( .A(n595), .B(n97), .Z(n3891) );
  XOR \MIXCOLUMNS[2].d/U81  ( .A(n595), .B(n96), .Z(n4003) );
  XOR \MIXCOLUMNS[2].d/U80  ( .A(n3893), .B(n3892), .Z(\w0[3][102] ) );
  XOR \MIXCOLUMNS[2].d/U79  ( .A(n4003), .B(n3894), .Z(n3892) );
  XOR \MIXCOLUMNS[2].d/U78  ( .A(n594), .B(n3990), .Z(n3893) );
  XOR \MIXCOLUMNS[2].d/U77  ( .A(n593), .B(n95), .Z(n3894) );
  XOR \MIXCOLUMNS[2].d/U76  ( .A(n593), .B(n94), .Z(n4005) );
  XOR \MIXCOLUMNS[2].d/U75  ( .A(n4005), .B(n3895), .Z(\w0[3][103] ) );
  XOR \MIXCOLUMNS[2].d/U74  ( .A(n93), .B(n3990), .Z(n3895) );
  XOR \MIXCOLUMNS[2].d/U73  ( .A(n104), .B(n604), .Z(n3994) );
  XOR \MIXCOLUMNS[2].d/U72  ( .A(n3994), .B(n3896), .Z(\w0[3][104] ) );
  XOR \MIXCOLUMNS[2].d/U71  ( .A(n103), .B(n4007), .Z(n3896) );
  XOR \MIXCOLUMNS[2].d/U70  ( .A(\w3[2][106] ), .B(\w3[2][98] ), .Z(n3996) );
  XOR \MIXCOLUMNS[2].d/U69  ( .A(n3996), .B(n3897), .Z(\w0[3][105] ) );
  XOR \MIXCOLUMNS[2].d/U68  ( .A(n604), .B(n3992), .Z(n3897) );
  XOR \MIXCOLUMNS[2].d/U67  ( .A(n101), .B(n602), .Z(n3998) );
  XOR \MIXCOLUMNS[2].d/U66  ( .A(n3998), .B(n3898), .Z(\w0[3][106] ) );
  XOR \MIXCOLUMNS[2].d/U65  ( .A(\w3[2][98] ), .B(n3995), .Z(n3898) );
  XOR \MIXCOLUMNS[2].d/U64  ( .A(n5), .B(n103), .Z(n3993) );
  XOR \MIXCOLUMNS[2].d/U63  ( .A(n99), .B(n600), .Z(n4000) );
  XOR \MIXCOLUMNS[2].d/U62  ( .A(n3900), .B(n3899), .Z(\w0[3][107] ) );
  XOR \MIXCOLUMNS[2].d/U61  ( .A(n3997), .B(n4000), .Z(n3899) );
  XOR \MIXCOLUMNS[2].d/U60  ( .A(n602), .B(n3993), .Z(n3900) );
  XOR \MIXCOLUMNS[2].d/U59  ( .A(n97), .B(n598), .Z(n4002) );
  XOR \MIXCOLUMNS[2].d/U58  ( .A(n3902), .B(n3901), .Z(\w0[3][108] ) );
  XOR \MIXCOLUMNS[2].d/U57  ( .A(n3999), .B(n4002), .Z(n3901) );
  XOR \MIXCOLUMNS[2].d/U56  ( .A(n600), .B(n3993), .Z(n3902) );
  XOR \MIXCOLUMNS[2].d/U55  ( .A(n95), .B(n596), .Z(n4004) );
  XOR \MIXCOLUMNS[2].d/U54  ( .A(n4004), .B(n3903), .Z(\w0[3][109] ) );
  XOR \MIXCOLUMNS[2].d/U53  ( .A(n598), .B(n4001), .Z(n3903) );
  XOR \MIXCOLUMNS[2].d/U52  ( .A(n93), .B(n594), .Z(n4006) );
  XOR \MIXCOLUMNS[2].d/U51  ( .A(n3905), .B(n3904), .Z(\w0[3][110] ) );
  XOR \MIXCOLUMNS[2].d/U50  ( .A(n4003), .B(n4006), .Z(n3904) );
  XOR \MIXCOLUMNS[2].d/U49  ( .A(n596), .B(n3993), .Z(n3905) );
  XOR \MIXCOLUMNS[2].d/U48  ( .A(n4005), .B(n3906), .Z(\w0[3][111] ) );
  XOR \MIXCOLUMNS[2].d/U47  ( .A(n594), .B(n3993), .Z(n3906) );
  XOR \MIXCOLUMNS[2].d/U46  ( .A(n3908), .B(n3907), .Z(\w0[3][112] ) );
  XOR \MIXCOLUMNS[2].d/U45  ( .A(n104), .B(n3993), .Z(n3907) );
  XOR \MIXCOLUMNS[2].d/U44  ( .A(n605), .B(n105), .Z(n3908) );
  XOR \MIXCOLUMNS[2].d/U43  ( .A(n3910), .B(n3909), .Z(\w0[3][113] ) );
  XOR \MIXCOLUMNS[2].d/U42  ( .A(\w3[2][106] ), .B(n3994), .Z(n3909) );
  XOR \MIXCOLUMNS[2].d/U41  ( .A(n603), .B(\w3[2][114] ), .Z(n3910) );
  XOR \MIXCOLUMNS[2].d/U40  ( .A(n3912), .B(n3911), .Z(\w0[3][114] ) );
  XOR \MIXCOLUMNS[2].d/U39  ( .A(n101), .B(n3996), .Z(n3911) );
  XOR \MIXCOLUMNS[2].d/U38  ( .A(\w3[2][122] ), .B(n102), .Z(n3912) );
  XOR \MIXCOLUMNS[2].d/U37  ( .A(n106), .B(n5), .Z(n3991) );
  XOR \MIXCOLUMNS[2].d/U36  ( .A(n3914), .B(n3913), .Z(\w0[3][115] ) );
  XOR \MIXCOLUMNS[2].d/U35  ( .A(n3998), .B(n3915), .Z(n3913) );
  XOR \MIXCOLUMNS[2].d/U34  ( .A(n99), .B(n3991), .Z(n3914) );
  XOR \MIXCOLUMNS[2].d/U33  ( .A(n601), .B(n100), .Z(n3915) );
  XOR \MIXCOLUMNS[2].d/U32  ( .A(n3917), .B(n3916), .Z(\w0[3][116] ) );
  XOR \MIXCOLUMNS[2].d/U31  ( .A(n4000), .B(n3918), .Z(n3916) );
  XOR \MIXCOLUMNS[2].d/U30  ( .A(n97), .B(n3991), .Z(n3917) );
  XOR \MIXCOLUMNS[2].d/U29  ( .A(n599), .B(n98), .Z(n3918) );
  XOR \MIXCOLUMNS[2].d/U28  ( .A(n3920), .B(n3919), .Z(\w0[3][117] ) );
  XOR \MIXCOLUMNS[2].d/U27  ( .A(n95), .B(n4002), .Z(n3919) );
  XOR \MIXCOLUMNS[2].d/U26  ( .A(n597), .B(n96), .Z(n3920) );
  XOR \MIXCOLUMNS[2].d/U25  ( .A(n3922), .B(n3921), .Z(\w0[3][118] ) );
  XOR \MIXCOLUMNS[2].d/U24  ( .A(n4004), .B(n3923), .Z(n3921) );
  XOR \MIXCOLUMNS[2].d/U23  ( .A(n93), .B(n3991), .Z(n3922) );
  XOR \MIXCOLUMNS[2].d/U22  ( .A(n595), .B(n94), .Z(n3923) );
  XOR \MIXCOLUMNS[2].d/U21  ( .A(n4006), .B(n3924), .Z(\w0[3][119] ) );
  XOR \MIXCOLUMNS[2].d/U20  ( .A(n593), .B(n3991), .Z(n3924) );
  XOR \MIXCOLUMNS[2].d/U19  ( .A(n3992), .B(n3925), .Z(\w0[3][120] ) );
  XOR \MIXCOLUMNS[2].d/U18  ( .A(n106), .B(n3993), .Z(n3925) );
  XOR \MIXCOLUMNS[2].d/U17  ( .A(n3994), .B(n3926), .Z(\w0[3][121] ) );
  XOR \MIXCOLUMNS[2].d/U16  ( .A(n105), .B(n3995), .Z(n3926) );
  XOR \MIXCOLUMNS[2].d/U15  ( .A(n3996), .B(n3927), .Z(\w0[3][122] ) );
  XOR \MIXCOLUMNS[2].d/U14  ( .A(\w3[2][114] ), .B(n3997), .Z(n3927) );
  XOR \MIXCOLUMNS[2].d/U13  ( .A(n3929), .B(n3928), .Z(\w0[3][123] ) );
  XOR \MIXCOLUMNS[2].d/U12  ( .A(n3999), .B(n3998), .Z(n3928) );
  XOR \MIXCOLUMNS[2].d/U11  ( .A(n102), .B(n4007), .Z(n3929) );
  XOR \MIXCOLUMNS[2].d/U10  ( .A(n3931), .B(n3930), .Z(\w0[3][124] ) );
  XOR \MIXCOLUMNS[2].d/U9  ( .A(n4001), .B(n4000), .Z(n3930) );
  XOR \MIXCOLUMNS[2].d/U8  ( .A(n100), .B(n4007), .Z(n3931) );
  XOR \MIXCOLUMNS[2].d/U7  ( .A(n4002), .B(n3932), .Z(\w0[3][125] ) );
  XOR \MIXCOLUMNS[2].d/U6  ( .A(n98), .B(n4003), .Z(n3932) );
  XOR \MIXCOLUMNS[2].d/U5  ( .A(n3934), .B(n3933), .Z(\w0[3][126] ) );
  XOR \MIXCOLUMNS[2].d/U4  ( .A(n4005), .B(n4004), .Z(n3933) );
  XOR \MIXCOLUMNS[2].d/U3  ( .A(n96), .B(n4007), .Z(n3934) );
  XOR \MIXCOLUMNS[2].d/U2  ( .A(n4006), .B(n3935), .Z(\w0[3][127] ) );
  XOR \MIXCOLUMNS[2].d/U1  ( .A(n94), .B(n4007), .Z(n3935) );
  XOR \MIXCOLUMNS[1].d/U432  ( .A(n592), .B(n92), .Z(n3649) );
  XOR \MIXCOLUMNS[1].d/U431  ( .A(n3401), .B(n3400), .Z(\w0[2][0] ) );
  XOR \MIXCOLUMNS[1].d/U430  ( .A(n591), .B(n3649), .Z(n3400) );
  XOR \MIXCOLUMNS[1].d/U429  ( .A(n590), .B(n4), .Z(n3401) );
  XOR \MIXCOLUMNS[1].d/U428  ( .A(n590), .B(n91), .Z(n3634) );
  XOR \MIXCOLUMNS[1].d/U427  ( .A(n3403), .B(n3402), .Z(\w0[2][1] ) );
  XOR \MIXCOLUMNS[1].d/U426  ( .A(\w3[1][2] ), .B(n3634), .Z(n3402) );
  XOR \MIXCOLUMNS[1].d/U425  ( .A(\w3[1][26] ), .B(n90), .Z(n3403) );
  XOR \MIXCOLUMNS[1].d/U424  ( .A(\w3[1][26] ), .B(\w3[1][18] ), .Z(n3637) );
  XOR \MIXCOLUMNS[1].d/U423  ( .A(n3405), .B(n3404), .Z(\w0[2][2] ) );
  XOR \MIXCOLUMNS[1].d/U422  ( .A(n589), .B(n3637), .Z(n3404) );
  XOR \MIXCOLUMNS[1].d/U421  ( .A(n588), .B(\w3[1][10] ), .Z(n3405) );
  XOR \MIXCOLUMNS[1].d/U420  ( .A(n592), .B(n89), .Z(n3632) );
  XOR \MIXCOLUMNS[1].d/U419  ( .A(n588), .B(n88), .Z(n3639) );
  XOR \MIXCOLUMNS[1].d/U418  ( .A(n3407), .B(n3406), .Z(\w0[2][3] ) );
  XOR \MIXCOLUMNS[1].d/U417  ( .A(n3639), .B(n3408), .Z(n3406) );
  XOR \MIXCOLUMNS[1].d/U416  ( .A(n587), .B(n3632), .Z(n3407) );
  XOR \MIXCOLUMNS[1].d/U415  ( .A(n586), .B(n87), .Z(n3408) );
  XOR \MIXCOLUMNS[1].d/U414  ( .A(n586), .B(n86), .Z(n3641) );
  XOR \MIXCOLUMNS[1].d/U413  ( .A(n3410), .B(n3409), .Z(\w0[2][4] ) );
  XOR \MIXCOLUMNS[1].d/U412  ( .A(n3641), .B(n3411), .Z(n3409) );
  XOR \MIXCOLUMNS[1].d/U411  ( .A(n585), .B(n3632), .Z(n3410) );
  XOR \MIXCOLUMNS[1].d/U410  ( .A(n584), .B(n85), .Z(n3411) );
  XOR \MIXCOLUMNS[1].d/U409  ( .A(n584), .B(n84), .Z(n3643) );
  XOR \MIXCOLUMNS[1].d/U408  ( .A(n3413), .B(n3412), .Z(\w0[2][5] ) );
  XOR \MIXCOLUMNS[1].d/U407  ( .A(n583), .B(n3643), .Z(n3412) );
  XOR \MIXCOLUMNS[1].d/U406  ( .A(n582), .B(n83), .Z(n3413) );
  XOR \MIXCOLUMNS[1].d/U405  ( .A(n582), .B(n82), .Z(n3645) );
  XOR \MIXCOLUMNS[1].d/U404  ( .A(n3415), .B(n3414), .Z(\w0[2][6] ) );
  XOR \MIXCOLUMNS[1].d/U403  ( .A(n3645), .B(n3416), .Z(n3414) );
  XOR \MIXCOLUMNS[1].d/U402  ( .A(n581), .B(n3632), .Z(n3415) );
  XOR \MIXCOLUMNS[1].d/U401  ( .A(n580), .B(n81), .Z(n3416) );
  XOR \MIXCOLUMNS[1].d/U400  ( .A(n580), .B(n80), .Z(n3647) );
  XOR \MIXCOLUMNS[1].d/U399  ( .A(n3647), .B(n3417), .Z(\w0[2][7] ) );
  XOR \MIXCOLUMNS[1].d/U398  ( .A(n79), .B(n3632), .Z(n3417) );
  XOR \MIXCOLUMNS[1].d/U397  ( .A(n90), .B(n591), .Z(n3636) );
  XOR \MIXCOLUMNS[1].d/U396  ( .A(n3636), .B(n3418), .Z(\w0[2][8] ) );
  XOR \MIXCOLUMNS[1].d/U395  ( .A(n89), .B(n3649), .Z(n3418) );
  XOR \MIXCOLUMNS[1].d/U394  ( .A(\w3[1][10] ), .B(\w3[1][2] ), .Z(n3638) );
  XOR \MIXCOLUMNS[1].d/U393  ( .A(n3638), .B(n3419), .Z(\w0[2][9] ) );
  XOR \MIXCOLUMNS[1].d/U392  ( .A(n591), .B(n3634), .Z(n3419) );
  XOR \MIXCOLUMNS[1].d/U391  ( .A(n87), .B(n589), .Z(n3640) );
  XOR \MIXCOLUMNS[1].d/U390  ( .A(n3640), .B(n3420), .Z(\w0[2][10] ) );
  XOR \MIXCOLUMNS[1].d/U389  ( .A(\w3[1][2] ), .B(n3637), .Z(n3420) );
  XOR \MIXCOLUMNS[1].d/U388  ( .A(n4), .B(n89), .Z(n3635) );
  XOR \MIXCOLUMNS[1].d/U387  ( .A(n85), .B(n587), .Z(n3642) );
  XOR \MIXCOLUMNS[1].d/U386  ( .A(n3422), .B(n3421), .Z(\w0[2][11] ) );
  XOR \MIXCOLUMNS[1].d/U385  ( .A(n3639), .B(n3642), .Z(n3421) );
  XOR \MIXCOLUMNS[1].d/U384  ( .A(n589), .B(n3635), .Z(n3422) );
  XOR \MIXCOLUMNS[1].d/U383  ( .A(n83), .B(n585), .Z(n3644) );
  XOR \MIXCOLUMNS[1].d/U382  ( .A(n3424), .B(n3423), .Z(\w0[2][12] ) );
  XOR \MIXCOLUMNS[1].d/U381  ( .A(n3641), .B(n3644), .Z(n3423) );
  XOR \MIXCOLUMNS[1].d/U380  ( .A(n587), .B(n3635), .Z(n3424) );
  XOR \MIXCOLUMNS[1].d/U379  ( .A(n81), .B(n583), .Z(n3646) );
  XOR \MIXCOLUMNS[1].d/U378  ( .A(n3646), .B(n3425), .Z(\w0[2][13] ) );
  XOR \MIXCOLUMNS[1].d/U377  ( .A(n585), .B(n3643), .Z(n3425) );
  XOR \MIXCOLUMNS[1].d/U376  ( .A(n79), .B(n581), .Z(n3648) );
  XOR \MIXCOLUMNS[1].d/U375  ( .A(n3427), .B(n3426), .Z(\w0[2][14] ) );
  XOR \MIXCOLUMNS[1].d/U374  ( .A(n3645), .B(n3648), .Z(n3426) );
  XOR \MIXCOLUMNS[1].d/U373  ( .A(n583), .B(n3635), .Z(n3427) );
  XOR \MIXCOLUMNS[1].d/U372  ( .A(n3647), .B(n3428), .Z(\w0[2][15] ) );
  XOR \MIXCOLUMNS[1].d/U371  ( .A(n581), .B(n3635), .Z(n3428) );
  XOR \MIXCOLUMNS[1].d/U370  ( .A(n3430), .B(n3429), .Z(\w0[2][16] ) );
  XOR \MIXCOLUMNS[1].d/U369  ( .A(n90), .B(n3635), .Z(n3429) );
  XOR \MIXCOLUMNS[1].d/U368  ( .A(n592), .B(n91), .Z(n3430) );
  XOR \MIXCOLUMNS[1].d/U367  ( .A(n3432), .B(n3431), .Z(\w0[2][17] ) );
  XOR \MIXCOLUMNS[1].d/U366  ( .A(\w3[1][10] ), .B(n3636), .Z(n3431) );
  XOR \MIXCOLUMNS[1].d/U365  ( .A(n590), .B(\w3[1][18] ), .Z(n3432) );
  XOR \MIXCOLUMNS[1].d/U364  ( .A(n3434), .B(n3433), .Z(\w0[2][18] ) );
  XOR \MIXCOLUMNS[1].d/U363  ( .A(n87), .B(n3638), .Z(n3433) );
  XOR \MIXCOLUMNS[1].d/U362  ( .A(\w3[1][26] ), .B(n88), .Z(n3434) );
  XOR \MIXCOLUMNS[1].d/U361  ( .A(n92), .B(n4), .Z(n3633) );
  XOR \MIXCOLUMNS[1].d/U360  ( .A(n3436), .B(n3435), .Z(\w0[2][19] ) );
  XOR \MIXCOLUMNS[1].d/U359  ( .A(n3640), .B(n3437), .Z(n3435) );
  XOR \MIXCOLUMNS[1].d/U358  ( .A(n85), .B(n3633), .Z(n3436) );
  XOR \MIXCOLUMNS[1].d/U357  ( .A(n588), .B(n86), .Z(n3437) );
  XOR \MIXCOLUMNS[1].d/U356  ( .A(n3439), .B(n3438), .Z(\w0[2][20] ) );
  XOR \MIXCOLUMNS[1].d/U355  ( .A(n3642), .B(n3440), .Z(n3438) );
  XOR \MIXCOLUMNS[1].d/U354  ( .A(n83), .B(n3633), .Z(n3439) );
  XOR \MIXCOLUMNS[1].d/U353  ( .A(n586), .B(n84), .Z(n3440) );
  XOR \MIXCOLUMNS[1].d/U352  ( .A(n3442), .B(n3441), .Z(\w0[2][21] ) );
  XOR \MIXCOLUMNS[1].d/U351  ( .A(n81), .B(n3644), .Z(n3441) );
  XOR \MIXCOLUMNS[1].d/U350  ( .A(n584), .B(n82), .Z(n3442) );
  XOR \MIXCOLUMNS[1].d/U349  ( .A(n3444), .B(n3443), .Z(\w0[2][22] ) );
  XOR \MIXCOLUMNS[1].d/U348  ( .A(n3646), .B(n3445), .Z(n3443) );
  XOR \MIXCOLUMNS[1].d/U347  ( .A(n79), .B(n3633), .Z(n3444) );
  XOR \MIXCOLUMNS[1].d/U346  ( .A(n582), .B(n80), .Z(n3445) );
  XOR \MIXCOLUMNS[1].d/U345  ( .A(n3648), .B(n3446), .Z(\w0[2][23] ) );
  XOR \MIXCOLUMNS[1].d/U344  ( .A(n580), .B(n3633), .Z(n3446) );
  XOR \MIXCOLUMNS[1].d/U343  ( .A(n3634), .B(n3447), .Z(\w0[2][24] ) );
  XOR \MIXCOLUMNS[1].d/U342  ( .A(n92), .B(n3635), .Z(n3447) );
  XOR \MIXCOLUMNS[1].d/U341  ( .A(n3636), .B(n3448), .Z(\w0[2][25] ) );
  XOR \MIXCOLUMNS[1].d/U340  ( .A(n91), .B(n3637), .Z(n3448) );
  XOR \MIXCOLUMNS[1].d/U339  ( .A(n3638), .B(n3449), .Z(\w0[2][26] ) );
  XOR \MIXCOLUMNS[1].d/U338  ( .A(\w3[1][18] ), .B(n3639), .Z(n3449) );
  XOR \MIXCOLUMNS[1].d/U337  ( .A(n3451), .B(n3450), .Z(\w0[2][27] ) );
  XOR \MIXCOLUMNS[1].d/U336  ( .A(n3641), .B(n3640), .Z(n3450) );
  XOR \MIXCOLUMNS[1].d/U335  ( .A(n88), .B(n3649), .Z(n3451) );
  XOR \MIXCOLUMNS[1].d/U334  ( .A(n3453), .B(n3452), .Z(\w0[2][28] ) );
  XOR \MIXCOLUMNS[1].d/U333  ( .A(n3643), .B(n3642), .Z(n3452) );
  XOR \MIXCOLUMNS[1].d/U332  ( .A(n86), .B(n3649), .Z(n3453) );
  XOR \MIXCOLUMNS[1].d/U331  ( .A(n3644), .B(n3454), .Z(\w0[2][29] ) );
  XOR \MIXCOLUMNS[1].d/U330  ( .A(n84), .B(n3645), .Z(n3454) );
  XOR \MIXCOLUMNS[1].d/U329  ( .A(n3456), .B(n3455), .Z(\w0[2][30] ) );
  XOR \MIXCOLUMNS[1].d/U328  ( .A(n3647), .B(n3646), .Z(n3455) );
  XOR \MIXCOLUMNS[1].d/U327  ( .A(n82), .B(n3649), .Z(n3456) );
  XOR \MIXCOLUMNS[1].d/U326  ( .A(n3648), .B(n3457), .Z(\w0[2][31] ) );
  XOR \MIXCOLUMNS[1].d/U325  ( .A(n80), .B(n3649), .Z(n3457) );
  XOR \MIXCOLUMNS[1].d/U324  ( .A(n579), .B(n78), .Z(n3667) );
  XOR \MIXCOLUMNS[1].d/U323  ( .A(n3459), .B(n3458), .Z(\w0[2][32] ) );
  XOR \MIXCOLUMNS[1].d/U322  ( .A(n578), .B(n3667), .Z(n3458) );
  XOR \MIXCOLUMNS[1].d/U321  ( .A(n577), .B(n3), .Z(n3459) );
  XOR \MIXCOLUMNS[1].d/U320  ( .A(n577), .B(n77), .Z(n3652) );
  XOR \MIXCOLUMNS[1].d/U319  ( .A(n3461), .B(n3460), .Z(\w0[2][33] ) );
  XOR \MIXCOLUMNS[1].d/U318  ( .A(\w3[1][34] ), .B(n3652), .Z(n3460) );
  XOR \MIXCOLUMNS[1].d/U317  ( .A(\w3[1][58] ), .B(n76), .Z(n3461) );
  XOR \MIXCOLUMNS[1].d/U316  ( .A(\w3[1][58] ), .B(\w3[1][50] ), .Z(n3655) );
  XOR \MIXCOLUMNS[1].d/U315  ( .A(n3463), .B(n3462), .Z(\w0[2][34] ) );
  XOR \MIXCOLUMNS[1].d/U314  ( .A(n576), .B(n3655), .Z(n3462) );
  XOR \MIXCOLUMNS[1].d/U313  ( .A(n575), .B(\w3[1][42] ), .Z(n3463) );
  XOR \MIXCOLUMNS[1].d/U312  ( .A(n579), .B(n75), .Z(n3650) );
  XOR \MIXCOLUMNS[1].d/U311  ( .A(n575), .B(n74), .Z(n3657) );
  XOR \MIXCOLUMNS[1].d/U310  ( .A(n3465), .B(n3464), .Z(\w0[2][35] ) );
  XOR \MIXCOLUMNS[1].d/U309  ( .A(n3657), .B(n3466), .Z(n3464) );
  XOR \MIXCOLUMNS[1].d/U308  ( .A(n574), .B(n3650), .Z(n3465) );
  XOR \MIXCOLUMNS[1].d/U307  ( .A(n573), .B(n73), .Z(n3466) );
  XOR \MIXCOLUMNS[1].d/U306  ( .A(n573), .B(n72), .Z(n3659) );
  XOR \MIXCOLUMNS[1].d/U305  ( .A(n3468), .B(n3467), .Z(\w0[2][36] ) );
  XOR \MIXCOLUMNS[1].d/U304  ( .A(n3659), .B(n3469), .Z(n3467) );
  XOR \MIXCOLUMNS[1].d/U303  ( .A(n572), .B(n3650), .Z(n3468) );
  XOR \MIXCOLUMNS[1].d/U302  ( .A(n571), .B(n71), .Z(n3469) );
  XOR \MIXCOLUMNS[1].d/U301  ( .A(n571), .B(n70), .Z(n3661) );
  XOR \MIXCOLUMNS[1].d/U300  ( .A(n3471), .B(n3470), .Z(\w0[2][37] ) );
  XOR \MIXCOLUMNS[1].d/U299  ( .A(n570), .B(n3661), .Z(n3470) );
  XOR \MIXCOLUMNS[1].d/U298  ( .A(n569), .B(n69), .Z(n3471) );
  XOR \MIXCOLUMNS[1].d/U297  ( .A(n569), .B(n68), .Z(n3663) );
  XOR \MIXCOLUMNS[1].d/U296  ( .A(n3473), .B(n3472), .Z(\w0[2][38] ) );
  XOR \MIXCOLUMNS[1].d/U295  ( .A(n3663), .B(n3474), .Z(n3472) );
  XOR \MIXCOLUMNS[1].d/U294  ( .A(n568), .B(n3650), .Z(n3473) );
  XOR \MIXCOLUMNS[1].d/U293  ( .A(n567), .B(n67), .Z(n3474) );
  XOR \MIXCOLUMNS[1].d/U292  ( .A(n567), .B(n66), .Z(n3665) );
  XOR \MIXCOLUMNS[1].d/U291  ( .A(n3665), .B(n3475), .Z(\w0[2][39] ) );
  XOR \MIXCOLUMNS[1].d/U290  ( .A(n65), .B(n3650), .Z(n3475) );
  XOR \MIXCOLUMNS[1].d/U289  ( .A(n76), .B(n578), .Z(n3654) );
  XOR \MIXCOLUMNS[1].d/U288  ( .A(n3654), .B(n3476), .Z(\w0[2][40] ) );
  XOR \MIXCOLUMNS[1].d/U287  ( .A(n75), .B(n3667), .Z(n3476) );
  XOR \MIXCOLUMNS[1].d/U286  ( .A(\w3[1][42] ), .B(\w3[1][34] ), .Z(n3656) );
  XOR \MIXCOLUMNS[1].d/U285  ( .A(n3656), .B(n3477), .Z(\w0[2][41] ) );
  XOR \MIXCOLUMNS[1].d/U284  ( .A(n578), .B(n3652), .Z(n3477) );
  XOR \MIXCOLUMNS[1].d/U283  ( .A(n73), .B(n576), .Z(n3658) );
  XOR \MIXCOLUMNS[1].d/U282  ( .A(n3658), .B(n3478), .Z(\w0[2][42] ) );
  XOR \MIXCOLUMNS[1].d/U281  ( .A(\w3[1][34] ), .B(n3655), .Z(n3478) );
  XOR \MIXCOLUMNS[1].d/U280  ( .A(n3), .B(n75), .Z(n3653) );
  XOR \MIXCOLUMNS[1].d/U279  ( .A(n71), .B(n574), .Z(n3660) );
  XOR \MIXCOLUMNS[1].d/U278  ( .A(n3480), .B(n3479), .Z(\w0[2][43] ) );
  XOR \MIXCOLUMNS[1].d/U277  ( .A(n3657), .B(n3660), .Z(n3479) );
  XOR \MIXCOLUMNS[1].d/U276  ( .A(n576), .B(n3653), .Z(n3480) );
  XOR \MIXCOLUMNS[1].d/U275  ( .A(n69), .B(n572), .Z(n3662) );
  XOR \MIXCOLUMNS[1].d/U274  ( .A(n3482), .B(n3481), .Z(\w0[2][44] ) );
  XOR \MIXCOLUMNS[1].d/U273  ( .A(n3659), .B(n3662), .Z(n3481) );
  XOR \MIXCOLUMNS[1].d/U272  ( .A(n574), .B(n3653), .Z(n3482) );
  XOR \MIXCOLUMNS[1].d/U271  ( .A(n67), .B(n570), .Z(n3664) );
  XOR \MIXCOLUMNS[1].d/U270  ( .A(n3664), .B(n3483), .Z(\w0[2][45] ) );
  XOR \MIXCOLUMNS[1].d/U269  ( .A(n572), .B(n3661), .Z(n3483) );
  XOR \MIXCOLUMNS[1].d/U268  ( .A(n65), .B(n568), .Z(n3666) );
  XOR \MIXCOLUMNS[1].d/U267  ( .A(n3485), .B(n3484), .Z(\w0[2][46] ) );
  XOR \MIXCOLUMNS[1].d/U266  ( .A(n3663), .B(n3666), .Z(n3484) );
  XOR \MIXCOLUMNS[1].d/U265  ( .A(n570), .B(n3653), .Z(n3485) );
  XOR \MIXCOLUMNS[1].d/U264  ( .A(n3665), .B(n3486), .Z(\w0[2][47] ) );
  XOR \MIXCOLUMNS[1].d/U263  ( .A(n568), .B(n3653), .Z(n3486) );
  XOR \MIXCOLUMNS[1].d/U262  ( .A(n3488), .B(n3487), .Z(\w0[2][48] ) );
  XOR \MIXCOLUMNS[1].d/U261  ( .A(n76), .B(n3653), .Z(n3487) );
  XOR \MIXCOLUMNS[1].d/U260  ( .A(n579), .B(n77), .Z(n3488) );
  XOR \MIXCOLUMNS[1].d/U259  ( .A(n3490), .B(n3489), .Z(\w0[2][49] ) );
  XOR \MIXCOLUMNS[1].d/U258  ( .A(\w3[1][42] ), .B(n3654), .Z(n3489) );
  XOR \MIXCOLUMNS[1].d/U257  ( .A(n577), .B(\w3[1][50] ), .Z(n3490) );
  XOR \MIXCOLUMNS[1].d/U256  ( .A(n3492), .B(n3491), .Z(\w0[2][50] ) );
  XOR \MIXCOLUMNS[1].d/U255  ( .A(n73), .B(n3656), .Z(n3491) );
  XOR \MIXCOLUMNS[1].d/U254  ( .A(\w3[1][58] ), .B(n74), .Z(n3492) );
  XOR \MIXCOLUMNS[1].d/U253  ( .A(n78), .B(n3), .Z(n3651) );
  XOR \MIXCOLUMNS[1].d/U252  ( .A(n3494), .B(n3493), .Z(\w0[2][51] ) );
  XOR \MIXCOLUMNS[1].d/U251  ( .A(n3658), .B(n3495), .Z(n3493) );
  XOR \MIXCOLUMNS[1].d/U250  ( .A(n71), .B(n3651), .Z(n3494) );
  XOR \MIXCOLUMNS[1].d/U249  ( .A(n575), .B(n72), .Z(n3495) );
  XOR \MIXCOLUMNS[1].d/U248  ( .A(n3497), .B(n3496), .Z(\w0[2][52] ) );
  XOR \MIXCOLUMNS[1].d/U247  ( .A(n3660), .B(n3498), .Z(n3496) );
  XOR \MIXCOLUMNS[1].d/U246  ( .A(n69), .B(n3651), .Z(n3497) );
  XOR \MIXCOLUMNS[1].d/U245  ( .A(n573), .B(n70), .Z(n3498) );
  XOR \MIXCOLUMNS[1].d/U244  ( .A(n3500), .B(n3499), .Z(\w0[2][53] ) );
  XOR \MIXCOLUMNS[1].d/U243  ( .A(n67), .B(n3662), .Z(n3499) );
  XOR \MIXCOLUMNS[1].d/U242  ( .A(n571), .B(n68), .Z(n3500) );
  XOR \MIXCOLUMNS[1].d/U241  ( .A(n3502), .B(n3501), .Z(\w0[2][54] ) );
  XOR \MIXCOLUMNS[1].d/U240  ( .A(n3664), .B(n3503), .Z(n3501) );
  XOR \MIXCOLUMNS[1].d/U239  ( .A(n65), .B(n3651), .Z(n3502) );
  XOR \MIXCOLUMNS[1].d/U238  ( .A(n569), .B(n66), .Z(n3503) );
  XOR \MIXCOLUMNS[1].d/U237  ( .A(n3666), .B(n3504), .Z(\w0[2][55] ) );
  XOR \MIXCOLUMNS[1].d/U236  ( .A(n567), .B(n3651), .Z(n3504) );
  XOR \MIXCOLUMNS[1].d/U235  ( .A(n3652), .B(n3505), .Z(\w0[2][56] ) );
  XOR \MIXCOLUMNS[1].d/U234  ( .A(n78), .B(n3653), .Z(n3505) );
  XOR \MIXCOLUMNS[1].d/U233  ( .A(n3654), .B(n3506), .Z(\w0[2][57] ) );
  XOR \MIXCOLUMNS[1].d/U232  ( .A(n77), .B(n3655), .Z(n3506) );
  XOR \MIXCOLUMNS[1].d/U231  ( .A(n3656), .B(n3507), .Z(\w0[2][58] ) );
  XOR \MIXCOLUMNS[1].d/U230  ( .A(\w3[1][50] ), .B(n3657), .Z(n3507) );
  XOR \MIXCOLUMNS[1].d/U229  ( .A(n3509), .B(n3508), .Z(\w0[2][59] ) );
  XOR \MIXCOLUMNS[1].d/U228  ( .A(n3659), .B(n3658), .Z(n3508) );
  XOR \MIXCOLUMNS[1].d/U227  ( .A(n74), .B(n3667), .Z(n3509) );
  XOR \MIXCOLUMNS[1].d/U226  ( .A(n3511), .B(n3510), .Z(\w0[2][60] ) );
  XOR \MIXCOLUMNS[1].d/U225  ( .A(n3661), .B(n3660), .Z(n3510) );
  XOR \MIXCOLUMNS[1].d/U224  ( .A(n72), .B(n3667), .Z(n3511) );
  XOR \MIXCOLUMNS[1].d/U223  ( .A(n3662), .B(n3512), .Z(\w0[2][61] ) );
  XOR \MIXCOLUMNS[1].d/U222  ( .A(n70), .B(n3663), .Z(n3512) );
  XOR \MIXCOLUMNS[1].d/U221  ( .A(n3514), .B(n3513), .Z(\w0[2][62] ) );
  XOR \MIXCOLUMNS[1].d/U220  ( .A(n3665), .B(n3664), .Z(n3513) );
  XOR \MIXCOLUMNS[1].d/U219  ( .A(n68), .B(n3667), .Z(n3514) );
  XOR \MIXCOLUMNS[1].d/U218  ( .A(n3666), .B(n3515), .Z(\w0[2][63] ) );
  XOR \MIXCOLUMNS[1].d/U217  ( .A(n66), .B(n3667), .Z(n3515) );
  XOR \MIXCOLUMNS[1].d/U216  ( .A(n566), .B(n64), .Z(n3685) );
  XOR \MIXCOLUMNS[1].d/U215  ( .A(n3517), .B(n3516), .Z(\w0[2][64] ) );
  XOR \MIXCOLUMNS[1].d/U214  ( .A(n565), .B(n3685), .Z(n3516) );
  XOR \MIXCOLUMNS[1].d/U213  ( .A(n564), .B(n2), .Z(n3517) );
  XOR \MIXCOLUMNS[1].d/U212  ( .A(n564), .B(n63), .Z(n3670) );
  XOR \MIXCOLUMNS[1].d/U211  ( .A(n3519), .B(n3518), .Z(\w0[2][65] ) );
  XOR \MIXCOLUMNS[1].d/U210  ( .A(\w3[1][66] ), .B(n3670), .Z(n3518) );
  XOR \MIXCOLUMNS[1].d/U209  ( .A(\w3[1][90] ), .B(n62), .Z(n3519) );
  XOR \MIXCOLUMNS[1].d/U208  ( .A(\w3[1][90] ), .B(\w3[1][82] ), .Z(n3673) );
  XOR \MIXCOLUMNS[1].d/U207  ( .A(n3521), .B(n3520), .Z(\w0[2][66] ) );
  XOR \MIXCOLUMNS[1].d/U206  ( .A(n563), .B(n3673), .Z(n3520) );
  XOR \MIXCOLUMNS[1].d/U205  ( .A(n562), .B(\w3[1][74] ), .Z(n3521) );
  XOR \MIXCOLUMNS[1].d/U204  ( .A(n566), .B(n61), .Z(n3668) );
  XOR \MIXCOLUMNS[1].d/U203  ( .A(n562), .B(n60), .Z(n3675) );
  XOR \MIXCOLUMNS[1].d/U202  ( .A(n3523), .B(n3522), .Z(\w0[2][67] ) );
  XOR \MIXCOLUMNS[1].d/U201  ( .A(n3675), .B(n3524), .Z(n3522) );
  XOR \MIXCOLUMNS[1].d/U200  ( .A(n561), .B(n3668), .Z(n3523) );
  XOR \MIXCOLUMNS[1].d/U199  ( .A(n560), .B(n59), .Z(n3524) );
  XOR \MIXCOLUMNS[1].d/U198  ( .A(n560), .B(n58), .Z(n3677) );
  XOR \MIXCOLUMNS[1].d/U197  ( .A(n3526), .B(n3525), .Z(\w0[2][68] ) );
  XOR \MIXCOLUMNS[1].d/U196  ( .A(n3677), .B(n3527), .Z(n3525) );
  XOR \MIXCOLUMNS[1].d/U195  ( .A(n559), .B(n3668), .Z(n3526) );
  XOR \MIXCOLUMNS[1].d/U194  ( .A(n558), .B(n57), .Z(n3527) );
  XOR \MIXCOLUMNS[1].d/U193  ( .A(n558), .B(n56), .Z(n3679) );
  XOR \MIXCOLUMNS[1].d/U192  ( .A(n3529), .B(n3528), .Z(\w0[2][69] ) );
  XOR \MIXCOLUMNS[1].d/U191  ( .A(n557), .B(n3679), .Z(n3528) );
  XOR \MIXCOLUMNS[1].d/U190  ( .A(n556), .B(n55), .Z(n3529) );
  XOR \MIXCOLUMNS[1].d/U189  ( .A(n556), .B(n54), .Z(n3681) );
  XOR \MIXCOLUMNS[1].d/U188  ( .A(n3531), .B(n3530), .Z(\w0[2][70] ) );
  XOR \MIXCOLUMNS[1].d/U187  ( .A(n3681), .B(n3532), .Z(n3530) );
  XOR \MIXCOLUMNS[1].d/U186  ( .A(n555), .B(n3668), .Z(n3531) );
  XOR \MIXCOLUMNS[1].d/U185  ( .A(n554), .B(n53), .Z(n3532) );
  XOR \MIXCOLUMNS[1].d/U184  ( .A(n554), .B(n52), .Z(n3683) );
  XOR \MIXCOLUMNS[1].d/U183  ( .A(n3683), .B(n3533), .Z(\w0[2][71] ) );
  XOR \MIXCOLUMNS[1].d/U182  ( .A(n51), .B(n3668), .Z(n3533) );
  XOR \MIXCOLUMNS[1].d/U181  ( .A(n62), .B(n565), .Z(n3672) );
  XOR \MIXCOLUMNS[1].d/U180  ( .A(n3672), .B(n3534), .Z(\w0[2][72] ) );
  XOR \MIXCOLUMNS[1].d/U179  ( .A(n61), .B(n3685), .Z(n3534) );
  XOR \MIXCOLUMNS[1].d/U178  ( .A(\w3[1][74] ), .B(\w3[1][66] ), .Z(n3674) );
  XOR \MIXCOLUMNS[1].d/U177  ( .A(n3674), .B(n3535), .Z(\w0[2][73] ) );
  XOR \MIXCOLUMNS[1].d/U176  ( .A(n565), .B(n3670), .Z(n3535) );
  XOR \MIXCOLUMNS[1].d/U175  ( .A(n59), .B(n563), .Z(n3676) );
  XOR \MIXCOLUMNS[1].d/U174  ( .A(n3676), .B(n3536), .Z(\w0[2][74] ) );
  XOR \MIXCOLUMNS[1].d/U173  ( .A(\w3[1][66] ), .B(n3673), .Z(n3536) );
  XOR \MIXCOLUMNS[1].d/U172  ( .A(n2), .B(n61), .Z(n3671) );
  XOR \MIXCOLUMNS[1].d/U171  ( .A(n57), .B(n561), .Z(n3678) );
  XOR \MIXCOLUMNS[1].d/U170  ( .A(n3538), .B(n3537), .Z(\w0[2][75] ) );
  XOR \MIXCOLUMNS[1].d/U169  ( .A(n3675), .B(n3678), .Z(n3537) );
  XOR \MIXCOLUMNS[1].d/U168  ( .A(n563), .B(n3671), .Z(n3538) );
  XOR \MIXCOLUMNS[1].d/U167  ( .A(n55), .B(n559), .Z(n3680) );
  XOR \MIXCOLUMNS[1].d/U166  ( .A(n3540), .B(n3539), .Z(\w0[2][76] ) );
  XOR \MIXCOLUMNS[1].d/U165  ( .A(n3677), .B(n3680), .Z(n3539) );
  XOR \MIXCOLUMNS[1].d/U164  ( .A(n561), .B(n3671), .Z(n3540) );
  XOR \MIXCOLUMNS[1].d/U163  ( .A(n53), .B(n557), .Z(n3682) );
  XOR \MIXCOLUMNS[1].d/U162  ( .A(n3682), .B(n3541), .Z(\w0[2][77] ) );
  XOR \MIXCOLUMNS[1].d/U161  ( .A(n559), .B(n3679), .Z(n3541) );
  XOR \MIXCOLUMNS[1].d/U160  ( .A(n51), .B(n555), .Z(n3684) );
  XOR \MIXCOLUMNS[1].d/U159  ( .A(n3543), .B(n3542), .Z(\w0[2][78] ) );
  XOR \MIXCOLUMNS[1].d/U158  ( .A(n3681), .B(n3684), .Z(n3542) );
  XOR \MIXCOLUMNS[1].d/U157  ( .A(n557), .B(n3671), .Z(n3543) );
  XOR \MIXCOLUMNS[1].d/U156  ( .A(n3683), .B(n3544), .Z(\w0[2][79] ) );
  XOR \MIXCOLUMNS[1].d/U155  ( .A(n555), .B(n3671), .Z(n3544) );
  XOR \MIXCOLUMNS[1].d/U154  ( .A(n3546), .B(n3545), .Z(\w0[2][80] ) );
  XOR \MIXCOLUMNS[1].d/U153  ( .A(n62), .B(n3671), .Z(n3545) );
  XOR \MIXCOLUMNS[1].d/U152  ( .A(n566), .B(n63), .Z(n3546) );
  XOR \MIXCOLUMNS[1].d/U151  ( .A(n3548), .B(n3547), .Z(\w0[2][81] ) );
  XOR \MIXCOLUMNS[1].d/U150  ( .A(\w3[1][74] ), .B(n3672), .Z(n3547) );
  XOR \MIXCOLUMNS[1].d/U149  ( .A(n564), .B(\w3[1][82] ), .Z(n3548) );
  XOR \MIXCOLUMNS[1].d/U148  ( .A(n3550), .B(n3549), .Z(\w0[2][82] ) );
  XOR \MIXCOLUMNS[1].d/U147  ( .A(n59), .B(n3674), .Z(n3549) );
  XOR \MIXCOLUMNS[1].d/U146  ( .A(\w3[1][90] ), .B(n60), .Z(n3550) );
  XOR \MIXCOLUMNS[1].d/U145  ( .A(n64), .B(n2), .Z(n3669) );
  XOR \MIXCOLUMNS[1].d/U144  ( .A(n3552), .B(n3551), .Z(\w0[2][83] ) );
  XOR \MIXCOLUMNS[1].d/U143  ( .A(n3676), .B(n3553), .Z(n3551) );
  XOR \MIXCOLUMNS[1].d/U142  ( .A(n57), .B(n3669), .Z(n3552) );
  XOR \MIXCOLUMNS[1].d/U141  ( .A(n562), .B(n58), .Z(n3553) );
  XOR \MIXCOLUMNS[1].d/U140  ( .A(n3555), .B(n3554), .Z(\w0[2][84] ) );
  XOR \MIXCOLUMNS[1].d/U139  ( .A(n3678), .B(n3556), .Z(n3554) );
  XOR \MIXCOLUMNS[1].d/U138  ( .A(n55), .B(n3669), .Z(n3555) );
  XOR \MIXCOLUMNS[1].d/U137  ( .A(n560), .B(n56), .Z(n3556) );
  XOR \MIXCOLUMNS[1].d/U136  ( .A(n3558), .B(n3557), .Z(\w0[2][85] ) );
  XOR \MIXCOLUMNS[1].d/U135  ( .A(n53), .B(n3680), .Z(n3557) );
  XOR \MIXCOLUMNS[1].d/U134  ( .A(n558), .B(n54), .Z(n3558) );
  XOR \MIXCOLUMNS[1].d/U133  ( .A(n3560), .B(n3559), .Z(\w0[2][86] ) );
  XOR \MIXCOLUMNS[1].d/U132  ( .A(n3682), .B(n3561), .Z(n3559) );
  XOR \MIXCOLUMNS[1].d/U131  ( .A(n51), .B(n3669), .Z(n3560) );
  XOR \MIXCOLUMNS[1].d/U130  ( .A(n556), .B(n52), .Z(n3561) );
  XOR \MIXCOLUMNS[1].d/U129  ( .A(n3684), .B(n3562), .Z(\w0[2][87] ) );
  XOR \MIXCOLUMNS[1].d/U128  ( .A(n554), .B(n3669), .Z(n3562) );
  XOR \MIXCOLUMNS[1].d/U127  ( .A(n3670), .B(n3563), .Z(\w0[2][88] ) );
  XOR \MIXCOLUMNS[1].d/U126  ( .A(n64), .B(n3671), .Z(n3563) );
  XOR \MIXCOLUMNS[1].d/U125  ( .A(n3672), .B(n3564), .Z(\w0[2][89] ) );
  XOR \MIXCOLUMNS[1].d/U124  ( .A(n63), .B(n3673), .Z(n3564) );
  XOR \MIXCOLUMNS[1].d/U123  ( .A(n3674), .B(n3565), .Z(\w0[2][90] ) );
  XOR \MIXCOLUMNS[1].d/U122  ( .A(\w3[1][82] ), .B(n3675), .Z(n3565) );
  XOR \MIXCOLUMNS[1].d/U121  ( .A(n3567), .B(n3566), .Z(\w0[2][91] ) );
  XOR \MIXCOLUMNS[1].d/U120  ( .A(n3677), .B(n3676), .Z(n3566) );
  XOR \MIXCOLUMNS[1].d/U119  ( .A(n60), .B(n3685), .Z(n3567) );
  XOR \MIXCOLUMNS[1].d/U118  ( .A(n3569), .B(n3568), .Z(\w0[2][92] ) );
  XOR \MIXCOLUMNS[1].d/U117  ( .A(n3679), .B(n3678), .Z(n3568) );
  XOR \MIXCOLUMNS[1].d/U116  ( .A(n58), .B(n3685), .Z(n3569) );
  XOR \MIXCOLUMNS[1].d/U115  ( .A(n3680), .B(n3570), .Z(\w0[2][93] ) );
  XOR \MIXCOLUMNS[1].d/U114  ( .A(n56), .B(n3681), .Z(n3570) );
  XOR \MIXCOLUMNS[1].d/U113  ( .A(n3572), .B(n3571), .Z(\w0[2][94] ) );
  XOR \MIXCOLUMNS[1].d/U112  ( .A(n3683), .B(n3682), .Z(n3571) );
  XOR \MIXCOLUMNS[1].d/U111  ( .A(n54), .B(n3685), .Z(n3572) );
  XOR \MIXCOLUMNS[1].d/U110  ( .A(n3684), .B(n3573), .Z(\w0[2][95] ) );
  XOR \MIXCOLUMNS[1].d/U109  ( .A(n52), .B(n3685), .Z(n3573) );
  XOR \MIXCOLUMNS[1].d/U108  ( .A(n553), .B(n50), .Z(n3703) );
  XOR \MIXCOLUMNS[1].d/U107  ( .A(n3575), .B(n3574), .Z(\w0[2][96] ) );
  XOR \MIXCOLUMNS[1].d/U106  ( .A(n552), .B(n3703), .Z(n3574) );
  XOR \MIXCOLUMNS[1].d/U105  ( .A(n551), .B(n1), .Z(n3575) );
  XOR \MIXCOLUMNS[1].d/U104  ( .A(n551), .B(n49), .Z(n3688) );
  XOR \MIXCOLUMNS[1].d/U103  ( .A(n3577), .B(n3576), .Z(\w0[2][97] ) );
  XOR \MIXCOLUMNS[1].d/U102  ( .A(\w3[1][98] ), .B(n3688), .Z(n3576) );
  XOR \MIXCOLUMNS[1].d/U101  ( .A(\w3[1][122] ), .B(n48), .Z(n3577) );
  XOR \MIXCOLUMNS[1].d/U100  ( .A(\w3[1][122] ), .B(\w3[1][114] ), .Z(n3691)
         );
  XOR \MIXCOLUMNS[1].d/U99  ( .A(n3579), .B(n3578), .Z(\w0[2][98] ) );
  XOR \MIXCOLUMNS[1].d/U98  ( .A(n550), .B(n3691), .Z(n3578) );
  XOR \MIXCOLUMNS[1].d/U97  ( .A(n549), .B(\w3[1][106] ), .Z(n3579) );
  XOR \MIXCOLUMNS[1].d/U96  ( .A(n553), .B(n47), .Z(n3686) );
  XOR \MIXCOLUMNS[1].d/U95  ( .A(n549), .B(n46), .Z(n3693) );
  XOR \MIXCOLUMNS[1].d/U94  ( .A(n3581), .B(n3580), .Z(\w0[2][99] ) );
  XOR \MIXCOLUMNS[1].d/U93  ( .A(n3693), .B(n3582), .Z(n3580) );
  XOR \MIXCOLUMNS[1].d/U92  ( .A(n548), .B(n3686), .Z(n3581) );
  XOR \MIXCOLUMNS[1].d/U91  ( .A(n547), .B(n45), .Z(n3582) );
  XOR \MIXCOLUMNS[1].d/U90  ( .A(n547), .B(n44), .Z(n3695) );
  XOR \MIXCOLUMNS[1].d/U89  ( .A(n3584), .B(n3583), .Z(\w0[2][100] ) );
  XOR \MIXCOLUMNS[1].d/U88  ( .A(n3695), .B(n3585), .Z(n3583) );
  XOR \MIXCOLUMNS[1].d/U87  ( .A(n546), .B(n3686), .Z(n3584) );
  XOR \MIXCOLUMNS[1].d/U86  ( .A(n545), .B(n43), .Z(n3585) );
  XOR \MIXCOLUMNS[1].d/U85  ( .A(n545), .B(n42), .Z(n3697) );
  XOR \MIXCOLUMNS[1].d/U84  ( .A(n3587), .B(n3586), .Z(\w0[2][101] ) );
  XOR \MIXCOLUMNS[1].d/U83  ( .A(n544), .B(n3697), .Z(n3586) );
  XOR \MIXCOLUMNS[1].d/U82  ( .A(n543), .B(n41), .Z(n3587) );
  XOR \MIXCOLUMNS[1].d/U81  ( .A(n543), .B(n40), .Z(n3699) );
  XOR \MIXCOLUMNS[1].d/U80  ( .A(n3589), .B(n3588), .Z(\w0[2][102] ) );
  XOR \MIXCOLUMNS[1].d/U79  ( .A(n3699), .B(n3590), .Z(n3588) );
  XOR \MIXCOLUMNS[1].d/U78  ( .A(n542), .B(n3686), .Z(n3589) );
  XOR \MIXCOLUMNS[1].d/U77  ( .A(n541), .B(n39), .Z(n3590) );
  XOR \MIXCOLUMNS[1].d/U76  ( .A(n541), .B(n38), .Z(n3701) );
  XOR \MIXCOLUMNS[1].d/U75  ( .A(n3701), .B(n3591), .Z(\w0[2][103] ) );
  XOR \MIXCOLUMNS[1].d/U74  ( .A(n37), .B(n3686), .Z(n3591) );
  XOR \MIXCOLUMNS[1].d/U73  ( .A(n48), .B(n552), .Z(n3690) );
  XOR \MIXCOLUMNS[1].d/U72  ( .A(n3690), .B(n3592), .Z(\w0[2][104] ) );
  XOR \MIXCOLUMNS[1].d/U71  ( .A(n47), .B(n3703), .Z(n3592) );
  XOR \MIXCOLUMNS[1].d/U70  ( .A(\w3[1][106] ), .B(\w3[1][98] ), .Z(n3692) );
  XOR \MIXCOLUMNS[1].d/U69  ( .A(n3692), .B(n3593), .Z(\w0[2][105] ) );
  XOR \MIXCOLUMNS[1].d/U68  ( .A(n552), .B(n3688), .Z(n3593) );
  XOR \MIXCOLUMNS[1].d/U67  ( .A(n45), .B(n550), .Z(n3694) );
  XOR \MIXCOLUMNS[1].d/U66  ( .A(n3694), .B(n3594), .Z(\w0[2][106] ) );
  XOR \MIXCOLUMNS[1].d/U65  ( .A(\w3[1][98] ), .B(n3691), .Z(n3594) );
  XOR \MIXCOLUMNS[1].d/U64  ( .A(n1), .B(n47), .Z(n3689) );
  XOR \MIXCOLUMNS[1].d/U63  ( .A(n43), .B(n548), .Z(n3696) );
  XOR \MIXCOLUMNS[1].d/U62  ( .A(n3596), .B(n3595), .Z(\w0[2][107] ) );
  XOR \MIXCOLUMNS[1].d/U61  ( .A(n3693), .B(n3696), .Z(n3595) );
  XOR \MIXCOLUMNS[1].d/U60  ( .A(n550), .B(n3689), .Z(n3596) );
  XOR \MIXCOLUMNS[1].d/U59  ( .A(n41), .B(n546), .Z(n3698) );
  XOR \MIXCOLUMNS[1].d/U58  ( .A(n3598), .B(n3597), .Z(\w0[2][108] ) );
  XOR \MIXCOLUMNS[1].d/U57  ( .A(n3695), .B(n3698), .Z(n3597) );
  XOR \MIXCOLUMNS[1].d/U56  ( .A(n548), .B(n3689), .Z(n3598) );
  XOR \MIXCOLUMNS[1].d/U55  ( .A(n39), .B(n544), .Z(n3700) );
  XOR \MIXCOLUMNS[1].d/U54  ( .A(n3700), .B(n3599), .Z(\w0[2][109] ) );
  XOR \MIXCOLUMNS[1].d/U53  ( .A(n546), .B(n3697), .Z(n3599) );
  XOR \MIXCOLUMNS[1].d/U52  ( .A(n37), .B(n542), .Z(n3702) );
  XOR \MIXCOLUMNS[1].d/U51  ( .A(n3601), .B(n3600), .Z(\w0[2][110] ) );
  XOR \MIXCOLUMNS[1].d/U50  ( .A(n3699), .B(n3702), .Z(n3600) );
  XOR \MIXCOLUMNS[1].d/U49  ( .A(n544), .B(n3689), .Z(n3601) );
  XOR \MIXCOLUMNS[1].d/U48  ( .A(n3701), .B(n3602), .Z(\w0[2][111] ) );
  XOR \MIXCOLUMNS[1].d/U47  ( .A(n542), .B(n3689), .Z(n3602) );
  XOR \MIXCOLUMNS[1].d/U46  ( .A(n3604), .B(n3603), .Z(\w0[2][112] ) );
  XOR \MIXCOLUMNS[1].d/U45  ( .A(n48), .B(n3689), .Z(n3603) );
  XOR \MIXCOLUMNS[1].d/U44  ( .A(n553), .B(n49), .Z(n3604) );
  XOR \MIXCOLUMNS[1].d/U43  ( .A(n3606), .B(n3605), .Z(\w0[2][113] ) );
  XOR \MIXCOLUMNS[1].d/U42  ( .A(\w3[1][106] ), .B(n3690), .Z(n3605) );
  XOR \MIXCOLUMNS[1].d/U41  ( .A(n551), .B(\w3[1][114] ), .Z(n3606) );
  XOR \MIXCOLUMNS[1].d/U40  ( .A(n3608), .B(n3607), .Z(\w0[2][114] ) );
  XOR \MIXCOLUMNS[1].d/U39  ( .A(n45), .B(n3692), .Z(n3607) );
  XOR \MIXCOLUMNS[1].d/U38  ( .A(\w3[1][122] ), .B(n46), .Z(n3608) );
  XOR \MIXCOLUMNS[1].d/U37  ( .A(n50), .B(n1), .Z(n3687) );
  XOR \MIXCOLUMNS[1].d/U36  ( .A(n3610), .B(n3609), .Z(\w0[2][115] ) );
  XOR \MIXCOLUMNS[1].d/U35  ( .A(n3694), .B(n3611), .Z(n3609) );
  XOR \MIXCOLUMNS[1].d/U34  ( .A(n43), .B(n3687), .Z(n3610) );
  XOR \MIXCOLUMNS[1].d/U33  ( .A(n549), .B(n44), .Z(n3611) );
  XOR \MIXCOLUMNS[1].d/U32  ( .A(n3613), .B(n3612), .Z(\w0[2][116] ) );
  XOR \MIXCOLUMNS[1].d/U31  ( .A(n3696), .B(n3614), .Z(n3612) );
  XOR \MIXCOLUMNS[1].d/U30  ( .A(n41), .B(n3687), .Z(n3613) );
  XOR \MIXCOLUMNS[1].d/U29  ( .A(n547), .B(n42), .Z(n3614) );
  XOR \MIXCOLUMNS[1].d/U28  ( .A(n3616), .B(n3615), .Z(\w0[2][117] ) );
  XOR \MIXCOLUMNS[1].d/U27  ( .A(n39), .B(n3698), .Z(n3615) );
  XOR \MIXCOLUMNS[1].d/U26  ( .A(n545), .B(n40), .Z(n3616) );
  XOR \MIXCOLUMNS[1].d/U25  ( .A(n3618), .B(n3617), .Z(\w0[2][118] ) );
  XOR \MIXCOLUMNS[1].d/U24  ( .A(n3700), .B(n3619), .Z(n3617) );
  XOR \MIXCOLUMNS[1].d/U23  ( .A(n37), .B(n3687), .Z(n3618) );
  XOR \MIXCOLUMNS[1].d/U22  ( .A(n543), .B(n38), .Z(n3619) );
  XOR \MIXCOLUMNS[1].d/U21  ( .A(n3702), .B(n3620), .Z(\w0[2][119] ) );
  XOR \MIXCOLUMNS[1].d/U20  ( .A(n541), .B(n3687), .Z(n3620) );
  XOR \MIXCOLUMNS[1].d/U19  ( .A(n3688), .B(n3621), .Z(\w0[2][120] ) );
  XOR \MIXCOLUMNS[1].d/U18  ( .A(n50), .B(n3689), .Z(n3621) );
  XOR \MIXCOLUMNS[1].d/U17  ( .A(n3690), .B(n3622), .Z(\w0[2][121] ) );
  XOR \MIXCOLUMNS[1].d/U16  ( .A(n49), .B(n3691), .Z(n3622) );
  XOR \MIXCOLUMNS[1].d/U15  ( .A(n3692), .B(n3623), .Z(\w0[2][122] ) );
  XOR \MIXCOLUMNS[1].d/U14  ( .A(\w3[1][114] ), .B(n3693), .Z(n3623) );
  XOR \MIXCOLUMNS[1].d/U13  ( .A(n3625), .B(n3624), .Z(\w0[2][123] ) );
  XOR \MIXCOLUMNS[1].d/U12  ( .A(n3695), .B(n3694), .Z(n3624) );
  XOR \MIXCOLUMNS[1].d/U11  ( .A(n46), .B(n3703), .Z(n3625) );
  XOR \MIXCOLUMNS[1].d/U10  ( .A(n3627), .B(n3626), .Z(\w0[2][124] ) );
  XOR \MIXCOLUMNS[1].d/U9  ( .A(n3697), .B(n3696), .Z(n3626) );
  XOR \MIXCOLUMNS[1].d/U8  ( .A(n44), .B(n3703), .Z(n3627) );
  XOR \MIXCOLUMNS[1].d/U7  ( .A(n3698), .B(n3628), .Z(\w0[2][125] ) );
  XOR \MIXCOLUMNS[1].d/U6  ( .A(n42), .B(n3699), .Z(n3628) );
  XOR \MIXCOLUMNS[1].d/U5  ( .A(n3630), .B(n3629), .Z(\w0[2][126] ) );
  XOR \MIXCOLUMNS[1].d/U4  ( .A(n3701), .B(n3700), .Z(n3629) );
  XOR \MIXCOLUMNS[1].d/U3  ( .A(n40), .B(n3703), .Z(n3630) );
  XOR \MIXCOLUMNS[1].d/U2  ( .A(n3702), .B(n3631), .Z(\w0[2][127] ) );
  XOR \MIXCOLUMNS[1].d/U1  ( .A(n38), .B(n3703), .Z(n3631) );
  XNOR U1 ( .A(n6929), .B(n5985), .Z(n1) );
  XNOR U2 ( .A(n6909), .B(n5889), .Z(n2) );
  XNOR U3 ( .A(n6969), .B(n6177), .Z(n3) );
  XNOR U4 ( .A(n6949), .B(n6081), .Z(n4) );
  XNOR U5 ( .A(n8209), .B(n7265), .Z(n5) );
  XNOR U6 ( .A(n8189), .B(n7169), .Z(n6) );
  XNOR U7 ( .A(n8249), .B(n7457), .Z(n7) );
  XNOR U8 ( .A(n8229), .B(n7361), .Z(n8) );
  XNOR U9 ( .A(n9489), .B(n8545), .Z(n9) );
  XNOR U10 ( .A(n9469), .B(n8449), .Z(n10) );
  XNOR U11 ( .A(n9529), .B(n8737), .Z(n11) );
  XNOR U12 ( .A(n9509), .B(n8641), .Z(n12) );
  XNOR U13 ( .A(n10769), .B(n9825), .Z(n13) );
  XNOR U14 ( .A(n10749), .B(n9729), .Z(n14) );
  XNOR U15 ( .A(n10809), .B(n10017), .Z(n15) );
  XNOR U16 ( .A(n10789), .B(n9921), .Z(n16) );
  XNOR U17 ( .A(n12049), .B(n11105), .Z(n17) );
  XNOR U18 ( .A(n12029), .B(n11009), .Z(n18) );
  XNOR U19 ( .A(n12089), .B(n11297), .Z(n19) );
  XNOR U20 ( .A(n12069), .B(n11201), .Z(n20) );
  XNOR U21 ( .A(n13329), .B(n12385), .Z(n21) );
  XNOR U22 ( .A(n13309), .B(n12289), .Z(n22) );
  XNOR U23 ( .A(n13369), .B(n12577), .Z(n23) );
  XNOR U24 ( .A(n13349), .B(n12481), .Z(n24) );
  XNOR U25 ( .A(n14609), .B(n13665), .Z(n25) );
  XNOR U26 ( .A(n14589), .B(n13569), .Z(n26) );
  XNOR U27 ( .A(n14649), .B(n13857), .Z(n27) );
  XNOR U28 ( .A(n14629), .B(n13761), .Z(n28) );
  XNOR U29 ( .A(n15889), .B(n14945), .Z(n29) );
  XNOR U30 ( .A(n15869), .B(n14849), .Z(n30) );
  XNOR U31 ( .A(n15929), .B(n15137), .Z(n31) );
  XNOR U32 ( .A(n15909), .B(n15041), .Z(n32) );
  XNOR U33 ( .A(\SUBBYTES[0].a/n1450 ), .B(\SUBBYTES[0].a/n506 ), .Z(n33) );
  XNOR U34 ( .A(\SUBBYTES[0].a/n1430 ), .B(\SUBBYTES[0].a/n410 ), .Z(n34) );
  XNOR U35 ( .A(\SUBBYTES[0].a/n1490 ), .B(\SUBBYTES[0].a/n698 ), .Z(n35) );
  XNOR U36 ( .A(\SUBBYTES[0].a/n1470 ), .B(\SUBBYTES[0].a/n602 ), .Z(n36) );
  XNOR U37 ( .A(n6006), .B(n6005), .Z(n37) );
  XNOR U38 ( .A(n6126), .B(n6125), .Z(n38) );
  XNOR U39 ( .A(n6003), .B(n6002), .Z(n39) );
  XNOR U40 ( .A(n6123), .B(n6122), .Z(n40) );
  XNOR U41 ( .A(n5997), .B(n5996), .Z(n41) );
  XNOR U42 ( .A(n6117), .B(n6116), .Z(n42) );
  XNOR U43 ( .A(n6929), .B(n5995), .Z(n43) );
  XNOR U44 ( .A(n6954), .B(n6115), .Z(n44) );
  XNOR U45 ( .A(n6931), .B(n5994), .Z(n45) );
  XNOR U46 ( .A(n6956), .B(n6114), .Z(n46) );
  XNOR U47 ( .A(n6904), .B(n5865), .Z(n47) );
  XNOR U48 ( .A(n6932), .B(n5988), .Z(n48) );
  XNOR U49 ( .A(n6957), .B(n6108), .Z(n49) );
  XNOR U50 ( .A(n6954), .B(n6105), .Z(n50) );
  XNOR U51 ( .A(n5910), .B(n5909), .Z(n51) );
  XNOR U52 ( .A(n6030), .B(n6029), .Z(n52) );
  XNOR U53 ( .A(n5907), .B(n5906), .Z(n53) );
  XNOR U54 ( .A(n6027), .B(n6026), .Z(n54) );
  XNOR U55 ( .A(n5901), .B(n5900), .Z(n55) );
  XNOR U56 ( .A(n6021), .B(n6020), .Z(n56) );
  XNOR U57 ( .A(n6909), .B(n5899), .Z(n57) );
  XNOR U58 ( .A(n6934), .B(n6019), .Z(n58) );
  XNOR U59 ( .A(n6911), .B(n5898), .Z(n59) );
  XNOR U60 ( .A(n6936), .B(n6018), .Z(n60) );
  XNOR U61 ( .A(n6964), .B(n6153), .Z(n61) );
  XNOR U62 ( .A(n6912), .B(n5892), .Z(n62) );
  XNOR U63 ( .A(n6937), .B(n6012), .Z(n63) );
  XNOR U64 ( .A(n6934), .B(n6009), .Z(n64) );
  XNOR U65 ( .A(n6198), .B(n6197), .Z(n65) );
  XNOR U66 ( .A(n5934), .B(n5933), .Z(n66) );
  XNOR U67 ( .A(n6195), .B(n6194), .Z(n67) );
  XNOR U68 ( .A(n5931), .B(n5930), .Z(n68) );
  XNOR U69 ( .A(n6189), .B(n6188), .Z(n69) );
  XNOR U70 ( .A(n5925), .B(n5924), .Z(n70) );
  XNOR U71 ( .A(n6969), .B(n6187), .Z(n71) );
  XNOR U72 ( .A(n6914), .B(n5923), .Z(n72) );
  XNOR U73 ( .A(n6971), .B(n6186), .Z(n73) );
  XNOR U74 ( .A(n6916), .B(n5922), .Z(n74) );
  XNOR U75 ( .A(n6944), .B(n6057), .Z(n75) );
  XNOR U76 ( .A(n6972), .B(n6180), .Z(n76) );
  XNOR U77 ( .A(n6917), .B(n5916), .Z(n77) );
  XNOR U78 ( .A(n6914), .B(n5913), .Z(n78) );
  XNOR U79 ( .A(n6102), .B(n6101), .Z(n79) );
  XNOR U80 ( .A(n6222), .B(n6221), .Z(n80) );
  XNOR U81 ( .A(n6099), .B(n6098), .Z(n81) );
  XNOR U82 ( .A(n6219), .B(n6218), .Z(n82) );
  XNOR U83 ( .A(n6093), .B(n6092), .Z(n83) );
  XNOR U84 ( .A(n6213), .B(n6212), .Z(n84) );
  XNOR U85 ( .A(n6949), .B(n6091), .Z(n85) );
  XNOR U86 ( .A(n6974), .B(n6211), .Z(n86) );
  XNOR U87 ( .A(n6951), .B(n6090), .Z(n87) );
  XNOR U88 ( .A(n6976), .B(n6210), .Z(n88) );
  XNOR U89 ( .A(n6924), .B(n5961), .Z(n89) );
  XNOR U90 ( .A(n6952), .B(n6084), .Z(n90) );
  XNOR U91 ( .A(n6977), .B(n6204), .Z(n91) );
  XNOR U92 ( .A(n6974), .B(n6201), .Z(n92) );
  XNOR U93 ( .A(n7286), .B(n7285), .Z(n93) );
  XNOR U94 ( .A(n7406), .B(n7405), .Z(n94) );
  XNOR U95 ( .A(n7283), .B(n7282), .Z(n95) );
  XNOR U96 ( .A(n7403), .B(n7402), .Z(n96) );
  XNOR U97 ( .A(n7277), .B(n7276), .Z(n97) );
  XNOR U98 ( .A(n7397), .B(n7396), .Z(n98) );
  XNOR U99 ( .A(n8209), .B(n7275), .Z(n99) );
  XNOR U100 ( .A(n8234), .B(n7395), .Z(n100) );
  XNOR U101 ( .A(n8211), .B(n7274), .Z(n101) );
  XNOR U102 ( .A(n8236), .B(n7394), .Z(n102) );
  XNOR U103 ( .A(n8184), .B(n7145), .Z(n103) );
  XNOR U104 ( .A(n8212), .B(n7268), .Z(n104) );
  XNOR U105 ( .A(n8237), .B(n7388), .Z(n105) );
  XNOR U106 ( .A(n8234), .B(n7385), .Z(n106) );
  XNOR U107 ( .A(n7190), .B(n7189), .Z(n107) );
  XNOR U108 ( .A(n7310), .B(n7309), .Z(n108) );
  XNOR U109 ( .A(n7187), .B(n7186), .Z(n109) );
  XNOR U110 ( .A(n7307), .B(n7306), .Z(n110) );
  XNOR U111 ( .A(n7181), .B(n7180), .Z(n111) );
  XNOR U112 ( .A(n7301), .B(n7300), .Z(n112) );
  XNOR U113 ( .A(n8189), .B(n7179), .Z(n113) );
  XNOR U114 ( .A(n8214), .B(n7299), .Z(n114) );
  XNOR U115 ( .A(n8191), .B(n7178), .Z(n115) );
  XNOR U116 ( .A(n8216), .B(n7298), .Z(n116) );
  XNOR U117 ( .A(n8244), .B(n7433), .Z(n117) );
  XNOR U118 ( .A(n8192), .B(n7172), .Z(n118) );
  XNOR U119 ( .A(n8217), .B(n7292), .Z(n119) );
  XNOR U120 ( .A(n8214), .B(n7289), .Z(n120) );
  XNOR U121 ( .A(n7478), .B(n7477), .Z(n121) );
  XNOR U122 ( .A(n7214), .B(n7213), .Z(n122) );
  XNOR U123 ( .A(n7475), .B(n7474), .Z(n123) );
  XNOR U124 ( .A(n7211), .B(n7210), .Z(n124) );
  XNOR U125 ( .A(n7469), .B(n7468), .Z(n125) );
  XNOR U126 ( .A(n7205), .B(n7204), .Z(n126) );
  XNOR U127 ( .A(n8249), .B(n7467), .Z(n127) );
  XNOR U128 ( .A(n8194), .B(n7203), .Z(n128) );
  XNOR U129 ( .A(n8251), .B(n7466), .Z(n129) );
  XNOR U130 ( .A(n8196), .B(n7202), .Z(n130) );
  XNOR U131 ( .A(n8224), .B(n7337), .Z(n131) );
  XNOR U132 ( .A(n8252), .B(n7460), .Z(n132) );
  XNOR U133 ( .A(n8197), .B(n7196), .Z(n133) );
  XNOR U134 ( .A(n8194), .B(n7193), .Z(n134) );
  XNOR U135 ( .A(n7382), .B(n7381), .Z(n135) );
  XNOR U136 ( .A(n7502), .B(n7501), .Z(n136) );
  XNOR U137 ( .A(n7379), .B(n7378), .Z(n137) );
  XNOR U138 ( .A(n7499), .B(n7498), .Z(n138) );
  XNOR U139 ( .A(n7373), .B(n7372), .Z(n139) );
  XNOR U140 ( .A(n7493), .B(n7492), .Z(n140) );
  XNOR U141 ( .A(n8229), .B(n7371), .Z(n141) );
  XNOR U142 ( .A(n8254), .B(n7491), .Z(n142) );
  XNOR U143 ( .A(n8231), .B(n7370), .Z(n143) );
  XNOR U144 ( .A(n8256), .B(n7490), .Z(n144) );
  XNOR U145 ( .A(n8204), .B(n7241), .Z(n145) );
  XNOR U146 ( .A(n8232), .B(n7364), .Z(n146) );
  XNOR U147 ( .A(n8257), .B(n7484), .Z(n147) );
  XNOR U148 ( .A(n8254), .B(n7481), .Z(n148) );
  XNOR U149 ( .A(n8566), .B(n8565), .Z(n149) );
  XNOR U150 ( .A(n8686), .B(n8685), .Z(n150) );
  XNOR U151 ( .A(n8563), .B(n8562), .Z(n151) );
  XNOR U152 ( .A(n8683), .B(n8682), .Z(n152) );
  XNOR U153 ( .A(n8557), .B(n8556), .Z(n153) );
  XNOR U154 ( .A(n8677), .B(n8676), .Z(n154) );
  XNOR U155 ( .A(n9489), .B(n8555), .Z(n155) );
  XNOR U156 ( .A(n9514), .B(n8675), .Z(n156) );
  XNOR U157 ( .A(n9491), .B(n8554), .Z(n157) );
  XNOR U158 ( .A(n9516), .B(n8674), .Z(n158) );
  XNOR U159 ( .A(n9464), .B(n8425), .Z(n159) );
  XNOR U160 ( .A(n9492), .B(n8548), .Z(n160) );
  XNOR U161 ( .A(n9517), .B(n8668), .Z(n161) );
  XNOR U162 ( .A(n9514), .B(n8665), .Z(n162) );
  XNOR U163 ( .A(n8470), .B(n8469), .Z(n163) );
  XNOR U164 ( .A(n8590), .B(n8589), .Z(n164) );
  XNOR U165 ( .A(n8467), .B(n8466), .Z(n165) );
  XNOR U166 ( .A(n8587), .B(n8586), .Z(n166) );
  XNOR U167 ( .A(n8461), .B(n8460), .Z(n167) );
  XNOR U168 ( .A(n8581), .B(n8580), .Z(n168) );
  XNOR U169 ( .A(n9469), .B(n8459), .Z(n169) );
  XNOR U170 ( .A(n9494), .B(n8579), .Z(n170) );
  XNOR U171 ( .A(n9471), .B(n8458), .Z(n171) );
  XNOR U172 ( .A(n9496), .B(n8578), .Z(n172) );
  XNOR U173 ( .A(n9524), .B(n8713), .Z(n173) );
  XNOR U174 ( .A(n9472), .B(n8452), .Z(n174) );
  XNOR U175 ( .A(n9497), .B(n8572), .Z(n175) );
  XNOR U176 ( .A(n9494), .B(n8569), .Z(n176) );
  XNOR U177 ( .A(n8758), .B(n8757), .Z(n177) );
  XNOR U178 ( .A(n8494), .B(n8493), .Z(n178) );
  XNOR U179 ( .A(n8755), .B(n8754), .Z(n179) );
  XNOR U180 ( .A(n8491), .B(n8490), .Z(n180) );
  XNOR U181 ( .A(n8749), .B(n8748), .Z(n181) );
  XNOR U182 ( .A(n8485), .B(n8484), .Z(n182) );
  XNOR U183 ( .A(n9529), .B(n8747), .Z(n183) );
  XNOR U184 ( .A(n9474), .B(n8483), .Z(n184) );
  XNOR U185 ( .A(n9531), .B(n8746), .Z(n185) );
  XNOR U186 ( .A(n9476), .B(n8482), .Z(n186) );
  XNOR U187 ( .A(n9504), .B(n8617), .Z(n187) );
  XNOR U188 ( .A(n9532), .B(n8740), .Z(n188) );
  XNOR U189 ( .A(n9477), .B(n8476), .Z(n189) );
  XNOR U190 ( .A(n9474), .B(n8473), .Z(n190) );
  XNOR U191 ( .A(n8662), .B(n8661), .Z(n191) );
  XNOR U192 ( .A(n8782), .B(n8781), .Z(n192) );
  XNOR U193 ( .A(n8659), .B(n8658), .Z(n193) );
  XNOR U194 ( .A(n8779), .B(n8778), .Z(n194) );
  XNOR U195 ( .A(n8653), .B(n8652), .Z(n195) );
  XNOR U196 ( .A(n8773), .B(n8772), .Z(n196) );
  XNOR U197 ( .A(n9509), .B(n8651), .Z(n197) );
  XNOR U198 ( .A(n9534), .B(n8771), .Z(n198) );
  XNOR U199 ( .A(n9511), .B(n8650), .Z(n199) );
  XNOR U200 ( .A(n9536), .B(n8770), .Z(n200) );
  XNOR U201 ( .A(n9484), .B(n8521), .Z(n201) );
  XNOR U202 ( .A(n9512), .B(n8644), .Z(n202) );
  XNOR U203 ( .A(n9537), .B(n8764), .Z(n203) );
  XNOR U204 ( .A(n9534), .B(n8761), .Z(n204) );
  XNOR U205 ( .A(n9846), .B(n9845), .Z(n205) );
  XNOR U206 ( .A(n9966), .B(n9965), .Z(n206) );
  XNOR U207 ( .A(n9843), .B(n9842), .Z(n207) );
  XNOR U208 ( .A(n9963), .B(n9962), .Z(n208) );
  XNOR U209 ( .A(n9837), .B(n9836), .Z(n209) );
  XNOR U210 ( .A(n9957), .B(n9956), .Z(n210) );
  XNOR U211 ( .A(n10769), .B(n9835), .Z(n211) );
  XNOR U212 ( .A(n10794), .B(n9955), .Z(n212) );
  XNOR U213 ( .A(n10771), .B(n9834), .Z(n213) );
  XNOR U214 ( .A(n10796), .B(n9954), .Z(n214) );
  XNOR U215 ( .A(n10744), .B(n9705), .Z(n215) );
  XNOR U216 ( .A(n10772), .B(n9828), .Z(n216) );
  XNOR U217 ( .A(n10797), .B(n9948), .Z(n217) );
  XNOR U218 ( .A(n10794), .B(n9945), .Z(n218) );
  XNOR U219 ( .A(n9750), .B(n9749), .Z(n219) );
  XNOR U220 ( .A(n9870), .B(n9869), .Z(n220) );
  XNOR U221 ( .A(n9747), .B(n9746), .Z(n221) );
  XNOR U222 ( .A(n9867), .B(n9866), .Z(n222) );
  XNOR U223 ( .A(n9741), .B(n9740), .Z(n223) );
  XNOR U224 ( .A(n9861), .B(n9860), .Z(n224) );
  XNOR U225 ( .A(n10749), .B(n9739), .Z(n225) );
  XNOR U226 ( .A(n10774), .B(n9859), .Z(n226) );
  XNOR U227 ( .A(n10751), .B(n9738), .Z(n227) );
  XNOR U228 ( .A(n10776), .B(n9858), .Z(n228) );
  XNOR U229 ( .A(n10804), .B(n9993), .Z(n229) );
  XNOR U230 ( .A(n10752), .B(n9732), .Z(n230) );
  XNOR U231 ( .A(n10777), .B(n9852), .Z(n231) );
  XNOR U232 ( .A(n10774), .B(n9849), .Z(n232) );
  XNOR U233 ( .A(n10038), .B(n10037), .Z(n233) );
  XNOR U234 ( .A(n9774), .B(n9773), .Z(n234) );
  XNOR U235 ( .A(n10035), .B(n10034), .Z(n235) );
  XNOR U236 ( .A(n9771), .B(n9770), .Z(n236) );
  XNOR U237 ( .A(n10029), .B(n10028), .Z(n237) );
  XNOR U238 ( .A(n9765), .B(n9764), .Z(n238) );
  XNOR U239 ( .A(n10809), .B(n10027), .Z(n239) );
  XNOR U240 ( .A(n10754), .B(n9763), .Z(n240) );
  XNOR U241 ( .A(n10811), .B(n10026), .Z(n241) );
  XNOR U242 ( .A(n10756), .B(n9762), .Z(n242) );
  XNOR U243 ( .A(n10784), .B(n9897), .Z(n243) );
  XNOR U244 ( .A(n10812), .B(n10020), .Z(n244) );
  XNOR U245 ( .A(n10757), .B(n9756), .Z(n245) );
  XNOR U246 ( .A(n10754), .B(n9753), .Z(n246) );
  XNOR U247 ( .A(n9942), .B(n9941), .Z(n247) );
  XNOR U248 ( .A(n10062), .B(n10061), .Z(n248) );
  XNOR U249 ( .A(n9939), .B(n9938), .Z(n249) );
  XNOR U250 ( .A(n10059), .B(n10058), .Z(n250) );
  XNOR U251 ( .A(n9933), .B(n9932), .Z(n251) );
  XNOR U252 ( .A(n10053), .B(n10052), .Z(n252) );
  XNOR U253 ( .A(n10789), .B(n9931), .Z(n253) );
  XNOR U254 ( .A(n10814), .B(n10051), .Z(n254) );
  XNOR U255 ( .A(n10791), .B(n9930), .Z(n255) );
  XNOR U256 ( .A(n10816), .B(n10050), .Z(n256) );
  XNOR U257 ( .A(n10764), .B(n9801), .Z(n257) );
  XNOR U258 ( .A(n10792), .B(n9924), .Z(n258) );
  XNOR U259 ( .A(n10817), .B(n10044), .Z(n259) );
  XNOR U260 ( .A(n10814), .B(n10041), .Z(n260) );
  XNOR U261 ( .A(n11126), .B(n11125), .Z(n261) );
  XNOR U262 ( .A(n11246), .B(n11245), .Z(n262) );
  XNOR U263 ( .A(n11123), .B(n11122), .Z(n263) );
  XNOR U264 ( .A(n11243), .B(n11242), .Z(n264) );
  XNOR U265 ( .A(n11117), .B(n11116), .Z(n265) );
  XNOR U266 ( .A(n11237), .B(n11236), .Z(n266) );
  XNOR U267 ( .A(n12049), .B(n11115), .Z(n267) );
  XNOR U268 ( .A(n12074), .B(n11235), .Z(n268) );
  XNOR U269 ( .A(n12051), .B(n11114), .Z(n269) );
  XNOR U270 ( .A(n12076), .B(n11234), .Z(n270) );
  XNOR U271 ( .A(n12024), .B(n10985), .Z(n271) );
  XNOR U272 ( .A(n12052), .B(n11108), .Z(n272) );
  XNOR U273 ( .A(n12077), .B(n11228), .Z(n273) );
  XNOR U274 ( .A(n12074), .B(n11225), .Z(n274) );
  XNOR U275 ( .A(n11030), .B(n11029), .Z(n275) );
  XNOR U276 ( .A(n11150), .B(n11149), .Z(n276) );
  XNOR U277 ( .A(n11027), .B(n11026), .Z(n277) );
  XNOR U278 ( .A(n11147), .B(n11146), .Z(n278) );
  XNOR U279 ( .A(n11021), .B(n11020), .Z(n279) );
  XNOR U280 ( .A(n11141), .B(n11140), .Z(n280) );
  XNOR U281 ( .A(n12029), .B(n11019), .Z(n281) );
  XNOR U282 ( .A(n12054), .B(n11139), .Z(n282) );
  XNOR U283 ( .A(n12031), .B(n11018), .Z(n283) );
  XNOR U284 ( .A(n12056), .B(n11138), .Z(n284) );
  XNOR U285 ( .A(n12084), .B(n11273), .Z(n285) );
  XNOR U286 ( .A(n12032), .B(n11012), .Z(n286) );
  XNOR U287 ( .A(n12057), .B(n11132), .Z(n287) );
  XNOR U288 ( .A(n12054), .B(n11129), .Z(n288) );
  XNOR U289 ( .A(n11318), .B(n11317), .Z(n289) );
  XNOR U290 ( .A(n11054), .B(n11053), .Z(n290) );
  XNOR U291 ( .A(n11315), .B(n11314), .Z(n291) );
  XNOR U292 ( .A(n11051), .B(n11050), .Z(n292) );
  XNOR U293 ( .A(n11309), .B(n11308), .Z(n293) );
  XNOR U294 ( .A(n11045), .B(n11044), .Z(n294) );
  XNOR U295 ( .A(n12089), .B(n11307), .Z(n295) );
  XNOR U296 ( .A(n12034), .B(n11043), .Z(n296) );
  XNOR U297 ( .A(n12091), .B(n11306), .Z(n297) );
  XNOR U298 ( .A(n12036), .B(n11042), .Z(n298) );
  XNOR U299 ( .A(n12064), .B(n11177), .Z(n299) );
  XNOR U300 ( .A(n12092), .B(n11300), .Z(n300) );
  XNOR U301 ( .A(n12037), .B(n11036), .Z(n301) );
  XNOR U302 ( .A(n12034), .B(n11033), .Z(n302) );
  XNOR U303 ( .A(n11222), .B(n11221), .Z(n303) );
  XNOR U304 ( .A(n11342), .B(n11341), .Z(n304) );
  XNOR U305 ( .A(n11219), .B(n11218), .Z(n305) );
  XNOR U306 ( .A(n11339), .B(n11338), .Z(n306) );
  XNOR U307 ( .A(n11213), .B(n11212), .Z(n307) );
  XNOR U308 ( .A(n11333), .B(n11332), .Z(n308) );
  XNOR U309 ( .A(n12069), .B(n11211), .Z(n309) );
  XNOR U310 ( .A(n12094), .B(n11331), .Z(n310) );
  XNOR U311 ( .A(n12071), .B(n11210), .Z(n311) );
  XNOR U312 ( .A(n12096), .B(n11330), .Z(n312) );
  XNOR U313 ( .A(n12044), .B(n11081), .Z(n313) );
  XNOR U314 ( .A(n12072), .B(n11204), .Z(n314) );
  XNOR U315 ( .A(n12097), .B(n11324), .Z(n315) );
  XNOR U316 ( .A(n12094), .B(n11321), .Z(n316) );
  XNOR U317 ( .A(n12406), .B(n12405), .Z(n317) );
  XNOR U318 ( .A(n12526), .B(n12525), .Z(n318) );
  XNOR U319 ( .A(n12403), .B(n12402), .Z(n319) );
  XNOR U320 ( .A(n12523), .B(n12522), .Z(n320) );
  XNOR U321 ( .A(n12397), .B(n12396), .Z(n321) );
  XNOR U322 ( .A(n12517), .B(n12516), .Z(n322) );
  XNOR U323 ( .A(n13329), .B(n12395), .Z(n323) );
  XNOR U324 ( .A(n13354), .B(n12515), .Z(n324) );
  XNOR U325 ( .A(n13331), .B(n12394), .Z(n325) );
  XNOR U326 ( .A(n13356), .B(n12514), .Z(n326) );
  XNOR U327 ( .A(n13304), .B(n12265), .Z(n327) );
  XNOR U328 ( .A(n13332), .B(n12388), .Z(n328) );
  XNOR U329 ( .A(n13357), .B(n12508), .Z(n329) );
  XNOR U330 ( .A(n13354), .B(n12505), .Z(n330) );
  XNOR U331 ( .A(n12310), .B(n12309), .Z(n331) );
  XNOR U332 ( .A(n12430), .B(n12429), .Z(n332) );
  XNOR U333 ( .A(n12307), .B(n12306), .Z(n333) );
  XNOR U334 ( .A(n12427), .B(n12426), .Z(n334) );
  XNOR U335 ( .A(n12301), .B(n12300), .Z(n335) );
  XNOR U336 ( .A(n12421), .B(n12420), .Z(n336) );
  XNOR U337 ( .A(n13309), .B(n12299), .Z(n337) );
  XNOR U338 ( .A(n13334), .B(n12419), .Z(n338) );
  XNOR U339 ( .A(n13311), .B(n12298), .Z(n339) );
  XNOR U340 ( .A(n13336), .B(n12418), .Z(n340) );
  XNOR U341 ( .A(n13364), .B(n12553), .Z(n341) );
  XNOR U342 ( .A(n13312), .B(n12292), .Z(n342) );
  XNOR U343 ( .A(n13337), .B(n12412), .Z(n343) );
  XNOR U344 ( .A(n13334), .B(n12409), .Z(n344) );
  XNOR U345 ( .A(n12598), .B(n12597), .Z(n345) );
  XNOR U346 ( .A(n12334), .B(n12333), .Z(n346) );
  XNOR U347 ( .A(n12595), .B(n12594), .Z(n347) );
  XNOR U348 ( .A(n12331), .B(n12330), .Z(n348) );
  XNOR U349 ( .A(n12589), .B(n12588), .Z(n349) );
  XNOR U350 ( .A(n12325), .B(n12324), .Z(n350) );
  XNOR U351 ( .A(n13369), .B(n12587), .Z(n351) );
  XNOR U352 ( .A(n13314), .B(n12323), .Z(n352) );
  XNOR U353 ( .A(n13371), .B(n12586), .Z(n353) );
  XNOR U354 ( .A(n13316), .B(n12322), .Z(n354) );
  XNOR U355 ( .A(n13344), .B(n12457), .Z(n355) );
  XNOR U356 ( .A(n13372), .B(n12580), .Z(n356) );
  XNOR U357 ( .A(n13317), .B(n12316), .Z(n357) );
  XNOR U358 ( .A(n13314), .B(n12313), .Z(n358) );
  XNOR U359 ( .A(n12502), .B(n12501), .Z(n359) );
  XNOR U360 ( .A(n12622), .B(n12621), .Z(n360) );
  XNOR U361 ( .A(n12499), .B(n12498), .Z(n361) );
  XNOR U362 ( .A(n12619), .B(n12618), .Z(n362) );
  XNOR U363 ( .A(n12493), .B(n12492), .Z(n363) );
  XNOR U364 ( .A(n12613), .B(n12612), .Z(n364) );
  XNOR U365 ( .A(n13349), .B(n12491), .Z(n365) );
  XNOR U366 ( .A(n13374), .B(n12611), .Z(n366) );
  XNOR U367 ( .A(n13351), .B(n12490), .Z(n367) );
  XNOR U368 ( .A(n13376), .B(n12610), .Z(n368) );
  XNOR U369 ( .A(n13324), .B(n12361), .Z(n369) );
  XNOR U370 ( .A(n13352), .B(n12484), .Z(n370) );
  XNOR U371 ( .A(n13377), .B(n12604), .Z(n371) );
  XNOR U372 ( .A(n13374), .B(n12601), .Z(n372) );
  XNOR U373 ( .A(n13686), .B(n13685), .Z(n373) );
  XNOR U374 ( .A(n13806), .B(n13805), .Z(n374) );
  XNOR U375 ( .A(n13683), .B(n13682), .Z(n375) );
  XNOR U376 ( .A(n13803), .B(n13802), .Z(n376) );
  XNOR U377 ( .A(n13677), .B(n13676), .Z(n377) );
  XNOR U378 ( .A(n13797), .B(n13796), .Z(n378) );
  XNOR U379 ( .A(n14609), .B(n13675), .Z(n379) );
  XNOR U380 ( .A(n14634), .B(n13795), .Z(n380) );
  XNOR U381 ( .A(n14611), .B(n13674), .Z(n381) );
  XNOR U382 ( .A(n14636), .B(n13794), .Z(n382) );
  XNOR U383 ( .A(n14584), .B(n13545), .Z(n383) );
  XNOR U384 ( .A(n14612), .B(n13668), .Z(n384) );
  XNOR U385 ( .A(n14637), .B(n13788), .Z(n385) );
  XNOR U386 ( .A(n14634), .B(n13785), .Z(n386) );
  XNOR U387 ( .A(n13590), .B(n13589), .Z(n387) );
  XNOR U388 ( .A(n13710), .B(n13709), .Z(n388) );
  XNOR U389 ( .A(n13587), .B(n13586), .Z(n389) );
  XNOR U390 ( .A(n13707), .B(n13706), .Z(n390) );
  XNOR U391 ( .A(n13581), .B(n13580), .Z(n391) );
  XNOR U392 ( .A(n13701), .B(n13700), .Z(n392) );
  XNOR U393 ( .A(n14589), .B(n13579), .Z(n393) );
  XNOR U394 ( .A(n14614), .B(n13699), .Z(n394) );
  XNOR U395 ( .A(n14591), .B(n13578), .Z(n395) );
  XNOR U396 ( .A(n14616), .B(n13698), .Z(n396) );
  XNOR U397 ( .A(n14644), .B(n13833), .Z(n397) );
  XNOR U398 ( .A(n14592), .B(n13572), .Z(n398) );
  XNOR U399 ( .A(n14617), .B(n13692), .Z(n399) );
  XNOR U400 ( .A(n14614), .B(n13689), .Z(n400) );
  XNOR U401 ( .A(n13878), .B(n13877), .Z(n401) );
  XNOR U402 ( .A(n13614), .B(n13613), .Z(n402) );
  XNOR U403 ( .A(n13875), .B(n13874), .Z(n403) );
  XNOR U404 ( .A(n13611), .B(n13610), .Z(n404) );
  XNOR U405 ( .A(n13869), .B(n13868), .Z(n405) );
  XNOR U406 ( .A(n13605), .B(n13604), .Z(n406) );
  XNOR U407 ( .A(n14649), .B(n13867), .Z(n407) );
  XNOR U408 ( .A(n14594), .B(n13603), .Z(n408) );
  XNOR U409 ( .A(n14651), .B(n13866), .Z(n409) );
  XNOR U410 ( .A(n14596), .B(n13602), .Z(n410) );
  XNOR U411 ( .A(n14624), .B(n13737), .Z(n411) );
  XNOR U412 ( .A(n14652), .B(n13860), .Z(n412) );
  XNOR U413 ( .A(n14597), .B(n13596), .Z(n413) );
  XNOR U414 ( .A(n14594), .B(n13593), .Z(n414) );
  XNOR U415 ( .A(n13782), .B(n13781), .Z(n415) );
  XNOR U416 ( .A(n13902), .B(n13901), .Z(n416) );
  XNOR U417 ( .A(n13779), .B(n13778), .Z(n417) );
  XNOR U418 ( .A(n13899), .B(n13898), .Z(n418) );
  XNOR U419 ( .A(n13773), .B(n13772), .Z(n419) );
  XNOR U420 ( .A(n13893), .B(n13892), .Z(n420) );
  XNOR U421 ( .A(n14629), .B(n13771), .Z(n421) );
  XNOR U422 ( .A(n14654), .B(n13891), .Z(n422) );
  XNOR U423 ( .A(n14631), .B(n13770), .Z(n423) );
  XNOR U424 ( .A(n14656), .B(n13890), .Z(n424) );
  XNOR U425 ( .A(n14604), .B(n13641), .Z(n425) );
  XNOR U426 ( .A(n14632), .B(n13764), .Z(n426) );
  XNOR U427 ( .A(n14657), .B(n13884), .Z(n427) );
  XNOR U428 ( .A(n14654), .B(n13881), .Z(n428) );
  XNOR U429 ( .A(n14966), .B(n14965), .Z(n429) );
  XNOR U430 ( .A(n15086), .B(n15085), .Z(n430) );
  XNOR U431 ( .A(n14963), .B(n14962), .Z(n431) );
  XNOR U432 ( .A(n15083), .B(n15082), .Z(n432) );
  XNOR U433 ( .A(n14957), .B(n14956), .Z(n433) );
  XNOR U434 ( .A(n15077), .B(n15076), .Z(n434) );
  XNOR U435 ( .A(n15889), .B(n14955), .Z(n435) );
  XNOR U436 ( .A(n15914), .B(n15075), .Z(n436) );
  XNOR U437 ( .A(n15891), .B(n14954), .Z(n437) );
  XNOR U438 ( .A(n15916), .B(n15074), .Z(n438) );
  XNOR U439 ( .A(n15864), .B(n14825), .Z(n439) );
  XNOR U440 ( .A(n15892), .B(n14948), .Z(n440) );
  XNOR U441 ( .A(n15917), .B(n15068), .Z(n441) );
  XNOR U442 ( .A(n15914), .B(n15065), .Z(n442) );
  XNOR U443 ( .A(n14870), .B(n14869), .Z(n443) );
  XNOR U444 ( .A(n14990), .B(n14989), .Z(n444) );
  XNOR U445 ( .A(n14867), .B(n14866), .Z(n445) );
  XNOR U446 ( .A(n14987), .B(n14986), .Z(n446) );
  XNOR U447 ( .A(n14861), .B(n14860), .Z(n447) );
  XNOR U448 ( .A(n14981), .B(n14980), .Z(n448) );
  XNOR U449 ( .A(n15869), .B(n14859), .Z(n449) );
  XNOR U450 ( .A(n15894), .B(n14979), .Z(n450) );
  XNOR U451 ( .A(n15871), .B(n14858), .Z(n451) );
  XNOR U452 ( .A(n15896), .B(n14978), .Z(n452) );
  XNOR U453 ( .A(n15924), .B(n15113), .Z(n453) );
  XNOR U454 ( .A(n15872), .B(n14852), .Z(n454) );
  XNOR U455 ( .A(n15897), .B(n14972), .Z(n455) );
  XNOR U456 ( .A(n15894), .B(n14969), .Z(n456) );
  XNOR U457 ( .A(n15158), .B(n15157), .Z(n457) );
  XNOR U458 ( .A(n14894), .B(n14893), .Z(n458) );
  XNOR U459 ( .A(n15155), .B(n15154), .Z(n459) );
  XNOR U460 ( .A(n14891), .B(n14890), .Z(n460) );
  XNOR U461 ( .A(n15149), .B(n15148), .Z(n461) );
  XNOR U462 ( .A(n14885), .B(n14884), .Z(n462) );
  XNOR U463 ( .A(n15929), .B(n15147), .Z(n463) );
  XNOR U464 ( .A(n15874), .B(n14883), .Z(n464) );
  XNOR U465 ( .A(n15931), .B(n15146), .Z(n465) );
  XNOR U466 ( .A(n15876), .B(n14882), .Z(n466) );
  XNOR U467 ( .A(n15904), .B(n15017), .Z(n467) );
  XNOR U468 ( .A(n15932), .B(n15140), .Z(n468) );
  XNOR U469 ( .A(n15877), .B(n14876), .Z(n469) );
  XNOR U470 ( .A(n15874), .B(n14873), .Z(n470) );
  XNOR U471 ( .A(n15062), .B(n15061), .Z(n471) );
  XNOR U472 ( .A(n15182), .B(n15181), .Z(n472) );
  XNOR U473 ( .A(n15059), .B(n15058), .Z(n473) );
  XNOR U474 ( .A(n15179), .B(n15178), .Z(n474) );
  XNOR U475 ( .A(n15053), .B(n15052), .Z(n475) );
  XNOR U476 ( .A(n15173), .B(n15172), .Z(n476) );
  XNOR U477 ( .A(n15909), .B(n15051), .Z(n477) );
  XNOR U478 ( .A(n15934), .B(n15171), .Z(n478) );
  XNOR U479 ( .A(n15911), .B(n15050), .Z(n479) );
  XNOR U480 ( .A(n15936), .B(n15170), .Z(n480) );
  XNOR U481 ( .A(n15884), .B(n14921), .Z(n481) );
  XNOR U482 ( .A(n15912), .B(n15044), .Z(n482) );
  XNOR U483 ( .A(n15937), .B(n15164), .Z(n483) );
  XNOR U484 ( .A(n15934), .B(n15161), .Z(n484) );
  XNOR U485 ( .A(\SUBBYTES[0].a/n527 ), .B(\SUBBYTES[0].a/n526 ), .Z(n485) );
  XNOR U486 ( .A(\SUBBYTES[0].a/n647 ), .B(\SUBBYTES[0].a/n646 ), .Z(n486) );
  XNOR U487 ( .A(\SUBBYTES[0].a/n524 ), .B(\SUBBYTES[0].a/n523 ), .Z(n487) );
  XNOR U488 ( .A(\SUBBYTES[0].a/n644 ), .B(\SUBBYTES[0].a/n643 ), .Z(n488) );
  XNOR U489 ( .A(\SUBBYTES[0].a/n518 ), .B(\SUBBYTES[0].a/n517 ), .Z(n489) );
  XNOR U490 ( .A(\SUBBYTES[0].a/n638 ), .B(\SUBBYTES[0].a/n637 ), .Z(n490) );
  XNOR U491 ( .A(\SUBBYTES[0].a/n1450 ), .B(\SUBBYTES[0].a/n516 ), .Z(n491) );
  XNOR U492 ( .A(\SUBBYTES[0].a/n1475 ), .B(\SUBBYTES[0].a/n636 ), .Z(n492) );
  XNOR U493 ( .A(\SUBBYTES[0].a/n1452 ), .B(\SUBBYTES[0].a/n515 ), .Z(n493) );
  XNOR U494 ( .A(\SUBBYTES[0].a/n1477 ), .B(\SUBBYTES[0].a/n635 ), .Z(n494) );
  XNOR U495 ( .A(\SUBBYTES[0].a/n1425 ), .B(\SUBBYTES[0].a/n386 ), .Z(n495) );
  XNOR U496 ( .A(\SUBBYTES[0].a/n1453 ), .B(\SUBBYTES[0].a/n509 ), .Z(n496) );
  XNOR U497 ( .A(\SUBBYTES[0].a/n1478 ), .B(\SUBBYTES[0].a/n629 ), .Z(n497) );
  XNOR U498 ( .A(\SUBBYTES[0].a/n1475 ), .B(\SUBBYTES[0].a/n626 ), .Z(n498) );
  XNOR U499 ( .A(\SUBBYTES[0].a/n431 ), .B(\SUBBYTES[0].a/n430 ), .Z(n499) );
  XNOR U500 ( .A(\SUBBYTES[0].a/n551 ), .B(\SUBBYTES[0].a/n550 ), .Z(n500) );
  XNOR U501 ( .A(\SUBBYTES[0].a/n428 ), .B(\SUBBYTES[0].a/n427 ), .Z(n501) );
  XNOR U502 ( .A(\SUBBYTES[0].a/n548 ), .B(\SUBBYTES[0].a/n547 ), .Z(n502) );
  XNOR U503 ( .A(\SUBBYTES[0].a/n422 ), .B(\SUBBYTES[0].a/n421 ), .Z(n503) );
  XNOR U504 ( .A(\SUBBYTES[0].a/n542 ), .B(\SUBBYTES[0].a/n541 ), .Z(n504) );
  XNOR U505 ( .A(\SUBBYTES[0].a/n1430 ), .B(\SUBBYTES[0].a/n420 ), .Z(n505) );
  XNOR U506 ( .A(\SUBBYTES[0].a/n1455 ), .B(\SUBBYTES[0].a/n540 ), .Z(n506) );
  XNOR U507 ( .A(\SUBBYTES[0].a/n1432 ), .B(\SUBBYTES[0].a/n419 ), .Z(n507) );
  XNOR U508 ( .A(\SUBBYTES[0].a/n1457 ), .B(\SUBBYTES[0].a/n539 ), .Z(n508) );
  XNOR U509 ( .A(\SUBBYTES[0].a/n1485 ), .B(\SUBBYTES[0].a/n674 ), .Z(n509) );
  XNOR U510 ( .A(\SUBBYTES[0].a/n1433 ), .B(\SUBBYTES[0].a/n413 ), .Z(n510) );
  XNOR U511 ( .A(\SUBBYTES[0].a/n1458 ), .B(\SUBBYTES[0].a/n533 ), .Z(n511) );
  XNOR U512 ( .A(\SUBBYTES[0].a/n1455 ), .B(\SUBBYTES[0].a/n530 ), .Z(n512) );
  XNOR U513 ( .A(\SUBBYTES[0].a/n719 ), .B(\SUBBYTES[0].a/n718 ), .Z(n513) );
  XNOR U514 ( .A(\SUBBYTES[0].a/n455 ), .B(\SUBBYTES[0].a/n454 ), .Z(n514) );
  XNOR U515 ( .A(\SUBBYTES[0].a/n716 ), .B(\SUBBYTES[0].a/n715 ), .Z(n515) );
  XNOR U516 ( .A(\SUBBYTES[0].a/n452 ), .B(\SUBBYTES[0].a/n451 ), .Z(n516) );
  XNOR U517 ( .A(\SUBBYTES[0].a/n710 ), .B(\SUBBYTES[0].a/n709 ), .Z(n517) );
  XNOR U518 ( .A(\SUBBYTES[0].a/n446 ), .B(\SUBBYTES[0].a/n445 ), .Z(n518) );
  XNOR U519 ( .A(\SUBBYTES[0].a/n1490 ), .B(\SUBBYTES[0].a/n708 ), .Z(n519) );
  XNOR U520 ( .A(\SUBBYTES[0].a/n1435 ), .B(\SUBBYTES[0].a/n444 ), .Z(n520) );
  XNOR U521 ( .A(\SUBBYTES[0].a/n1492 ), .B(\SUBBYTES[0].a/n707 ), .Z(n521) );
  XNOR U522 ( .A(\SUBBYTES[0].a/n1437 ), .B(\SUBBYTES[0].a/n443 ), .Z(n522) );
  XNOR U523 ( .A(\SUBBYTES[0].a/n1465 ), .B(\SUBBYTES[0].a/n578 ), .Z(n523) );
  XNOR U524 ( .A(\SUBBYTES[0].a/n1493 ), .B(\SUBBYTES[0].a/n701 ), .Z(n524) );
  XNOR U525 ( .A(\SUBBYTES[0].a/n1438 ), .B(\SUBBYTES[0].a/n437 ), .Z(n525) );
  XNOR U526 ( .A(\SUBBYTES[0].a/n1435 ), .B(\SUBBYTES[0].a/n434 ), .Z(n526) );
  XNOR U527 ( .A(\SUBBYTES[0].a/n623 ), .B(\SUBBYTES[0].a/n622 ), .Z(n527) );
  XNOR U528 ( .A(\SUBBYTES[0].a/n743 ), .B(\SUBBYTES[0].a/n742 ), .Z(n528) );
  XNOR U529 ( .A(\SUBBYTES[0].a/n620 ), .B(\SUBBYTES[0].a/n619 ), .Z(n529) );
  XNOR U530 ( .A(\SUBBYTES[0].a/n740 ), .B(\SUBBYTES[0].a/n739 ), .Z(n530) );
  XNOR U531 ( .A(\SUBBYTES[0].a/n614 ), .B(\SUBBYTES[0].a/n613 ), .Z(n531) );
  XNOR U532 ( .A(\SUBBYTES[0].a/n734 ), .B(\SUBBYTES[0].a/n733 ), .Z(n532) );
  XNOR U533 ( .A(\SUBBYTES[0].a/n1470 ), .B(\SUBBYTES[0].a/n612 ), .Z(n533) );
  XNOR U534 ( .A(\SUBBYTES[0].a/n1495 ), .B(\SUBBYTES[0].a/n732 ), .Z(n534) );
  XNOR U535 ( .A(\SUBBYTES[0].a/n1472 ), .B(\SUBBYTES[0].a/n611 ), .Z(n535) );
  XNOR U536 ( .A(\SUBBYTES[0].a/n1497 ), .B(\SUBBYTES[0].a/n731 ), .Z(n536) );
  XNOR U537 ( .A(\SUBBYTES[0].a/n1445 ), .B(\SUBBYTES[0].a/n482 ), .Z(n537) );
  XNOR U538 ( .A(\SUBBYTES[0].a/n1473 ), .B(\SUBBYTES[0].a/n605 ), .Z(n538) );
  XNOR U539 ( .A(\SUBBYTES[0].a/n1498 ), .B(\SUBBYTES[0].a/n725 ), .Z(n539) );
  XNOR U540 ( .A(\SUBBYTES[0].a/n1495 ), .B(\SUBBYTES[0].a/n722 ), .Z(n540) );
  XNOR U541 ( .A(n6246), .B(n6245), .Z(n541) );
  XNOR U542 ( .A(n5886), .B(n5885), .Z(n542) );
  XNOR U543 ( .A(n6243), .B(n6242), .Z(n543) );
  XNOR U544 ( .A(n5883), .B(n5882), .Z(n544) );
  XNOR U545 ( .A(n6237), .B(n6236), .Z(n545) );
  XNOR U546 ( .A(n5877), .B(n5876), .Z(n546) );
  XNOR U547 ( .A(n6979), .B(n6235), .Z(n547) );
  XNOR U548 ( .A(n6904), .B(n5875), .Z(n548) );
  XNOR U549 ( .A(n6981), .B(n6234), .Z(n549) );
  XNOR U550 ( .A(n6906), .B(n5874), .Z(n550) );
  XNOR U551 ( .A(n6982), .B(n6228), .Z(n551) );
  XNOR U552 ( .A(n6907), .B(n5868), .Z(n552) );
  XNOR U553 ( .A(n6979), .B(n6225), .Z(n553) );
  XNOR U554 ( .A(n6150), .B(n6149), .Z(n554) );
  XNOR U555 ( .A(n6174), .B(n6173), .Z(n555) );
  XNOR U556 ( .A(n6147), .B(n6146), .Z(n556) );
  XNOR U557 ( .A(n6171), .B(n6170), .Z(n557) );
  XNOR U558 ( .A(n6141), .B(n6140), .Z(n558) );
  XNOR U559 ( .A(n6165), .B(n6164), .Z(n559) );
  XNOR U560 ( .A(n6959), .B(n6139), .Z(n560) );
  XNOR U561 ( .A(n6964), .B(n6163), .Z(n561) );
  XNOR U562 ( .A(n6961), .B(n6138), .Z(n562) );
  XNOR U563 ( .A(n6966), .B(n6162), .Z(n563) );
  XNOR U564 ( .A(n6962), .B(n6132), .Z(n564) );
  XNOR U565 ( .A(n6967), .B(n6156), .Z(n565) );
  XNOR U566 ( .A(n6959), .B(n6129), .Z(n566) );
  XNOR U567 ( .A(n6054), .B(n6053), .Z(n567) );
  XNOR U568 ( .A(n6078), .B(n6077), .Z(n568) );
  XNOR U569 ( .A(n6051), .B(n6050), .Z(n569) );
  XNOR U570 ( .A(n6075), .B(n6074), .Z(n570) );
  XNOR U571 ( .A(n6045), .B(n6044), .Z(n571) );
  XNOR U572 ( .A(n6069), .B(n6068), .Z(n572) );
  XNOR U573 ( .A(n6939), .B(n6043), .Z(n573) );
  XNOR U574 ( .A(n6944), .B(n6067), .Z(n574) );
  XNOR U575 ( .A(n6941), .B(n6042), .Z(n575) );
  XNOR U576 ( .A(n6946), .B(n6066), .Z(n576) );
  XNOR U577 ( .A(n6942), .B(n6036), .Z(n577) );
  XNOR U578 ( .A(n6947), .B(n6060), .Z(n578) );
  XNOR U579 ( .A(n6939), .B(n6033), .Z(n579) );
  XNOR U580 ( .A(n5958), .B(n5957), .Z(n580) );
  XNOR U581 ( .A(n5982), .B(n5981), .Z(n581) );
  XNOR U582 ( .A(n5955), .B(n5954), .Z(n582) );
  XNOR U583 ( .A(n5979), .B(n5978), .Z(n583) );
  XNOR U584 ( .A(n5949), .B(n5948), .Z(n584) );
  XNOR U585 ( .A(n5973), .B(n5972), .Z(n585) );
  XNOR U586 ( .A(n6919), .B(n5947), .Z(n586) );
  XNOR U587 ( .A(n6924), .B(n5971), .Z(n587) );
  XNOR U588 ( .A(n6921), .B(n5946), .Z(n588) );
  XNOR U589 ( .A(n6926), .B(n5970), .Z(n589) );
  XNOR U590 ( .A(n6922), .B(n5940), .Z(n590) );
  XNOR U591 ( .A(n6927), .B(n5964), .Z(n591) );
  XNOR U592 ( .A(n6919), .B(n5937), .Z(n592) );
  XNOR U593 ( .A(n7526), .B(n7525), .Z(n593) );
  XNOR U594 ( .A(n7166), .B(n7165), .Z(n594) );
  XNOR U595 ( .A(n7523), .B(n7522), .Z(n595) );
  XNOR U596 ( .A(n7163), .B(n7162), .Z(n596) );
  XNOR U597 ( .A(n7517), .B(n7516), .Z(n597) );
  XNOR U598 ( .A(n7157), .B(n7156), .Z(n598) );
  XNOR U599 ( .A(n8259), .B(n7515), .Z(n599) );
  XNOR U600 ( .A(n8184), .B(n7155), .Z(n600) );
  XNOR U601 ( .A(n8261), .B(n7514), .Z(n601) );
  XNOR U602 ( .A(n8186), .B(n7154), .Z(n602) );
  XNOR U603 ( .A(n8262), .B(n7508), .Z(n603) );
  XNOR U604 ( .A(n8187), .B(n7148), .Z(n604) );
  XNOR U605 ( .A(n8259), .B(n7505), .Z(n605) );
  XNOR U606 ( .A(n7430), .B(n7429), .Z(n606) );
  XNOR U607 ( .A(n7454), .B(n7453), .Z(n607) );
  XNOR U608 ( .A(n7427), .B(n7426), .Z(n608) );
  XNOR U609 ( .A(n7451), .B(n7450), .Z(n609) );
  XNOR U610 ( .A(n7421), .B(n7420), .Z(n610) );
  XNOR U611 ( .A(n7445), .B(n7444), .Z(n611) );
  XNOR U612 ( .A(n8239), .B(n7419), .Z(n612) );
  XNOR U613 ( .A(n8244), .B(n7443), .Z(n613) );
  XNOR U614 ( .A(n8241), .B(n7418), .Z(n614) );
  XNOR U615 ( .A(n8246), .B(n7442), .Z(n615) );
  XNOR U616 ( .A(n8242), .B(n7412), .Z(n616) );
  XNOR U617 ( .A(n8247), .B(n7436), .Z(n617) );
  XNOR U618 ( .A(n8239), .B(n7409), .Z(n618) );
  XNOR U619 ( .A(n7334), .B(n7333), .Z(n619) );
  XNOR U620 ( .A(n7358), .B(n7357), .Z(n620) );
  XNOR U621 ( .A(n7331), .B(n7330), .Z(n621) );
  XNOR U622 ( .A(n7355), .B(n7354), .Z(n622) );
  XNOR U623 ( .A(n7325), .B(n7324), .Z(n623) );
  XNOR U624 ( .A(n7349), .B(n7348), .Z(n624) );
  XNOR U625 ( .A(n8219), .B(n7323), .Z(n625) );
  XNOR U626 ( .A(n8224), .B(n7347), .Z(n626) );
  XNOR U627 ( .A(n8221), .B(n7322), .Z(n627) );
  XNOR U628 ( .A(n8226), .B(n7346), .Z(n628) );
  XNOR U629 ( .A(n8222), .B(n7316), .Z(n629) );
  XNOR U630 ( .A(n8227), .B(n7340), .Z(n630) );
  XNOR U631 ( .A(n8219), .B(n7313), .Z(n631) );
  XNOR U632 ( .A(n7238), .B(n7237), .Z(n632) );
  XNOR U633 ( .A(n7262), .B(n7261), .Z(n633) );
  XNOR U634 ( .A(n7235), .B(n7234), .Z(n634) );
  XNOR U635 ( .A(n7259), .B(n7258), .Z(n635) );
  XNOR U636 ( .A(n7229), .B(n7228), .Z(n636) );
  XNOR U637 ( .A(n7253), .B(n7252), .Z(n637) );
  XNOR U638 ( .A(n8199), .B(n7227), .Z(n638) );
  XNOR U639 ( .A(n8204), .B(n7251), .Z(n639) );
  XNOR U640 ( .A(n8201), .B(n7226), .Z(n640) );
  XNOR U641 ( .A(n8206), .B(n7250), .Z(n641) );
  XNOR U642 ( .A(n8202), .B(n7220), .Z(n642) );
  XNOR U643 ( .A(n8207), .B(n7244), .Z(n643) );
  XNOR U644 ( .A(n8199), .B(n7217), .Z(n644) );
  XNOR U645 ( .A(n8806), .B(n8805), .Z(n645) );
  XNOR U646 ( .A(n8446), .B(n8445), .Z(n646) );
  XNOR U647 ( .A(n8803), .B(n8802), .Z(n647) );
  XNOR U648 ( .A(n8443), .B(n8442), .Z(n648) );
  XNOR U649 ( .A(n8797), .B(n8796), .Z(n649) );
  XNOR U650 ( .A(n8437), .B(n8436), .Z(n650) );
  XNOR U651 ( .A(n9539), .B(n8795), .Z(n651) );
  XNOR U652 ( .A(n9464), .B(n8435), .Z(n652) );
  XNOR U653 ( .A(n9541), .B(n8794), .Z(n653) );
  XNOR U654 ( .A(n9466), .B(n8434), .Z(n654) );
  XNOR U655 ( .A(n9542), .B(n8788), .Z(n655) );
  XNOR U656 ( .A(n9467), .B(n8428), .Z(n656) );
  XNOR U657 ( .A(n9539), .B(n8785), .Z(n657) );
  XNOR U658 ( .A(n8710), .B(n8709), .Z(n658) );
  XNOR U659 ( .A(n8734), .B(n8733), .Z(n659) );
  XNOR U660 ( .A(n8707), .B(n8706), .Z(n660) );
  XNOR U661 ( .A(n8731), .B(n8730), .Z(n661) );
  XNOR U662 ( .A(n8701), .B(n8700), .Z(n662) );
  XNOR U663 ( .A(n8725), .B(n8724), .Z(n663) );
  XNOR U664 ( .A(n9519), .B(n8699), .Z(n664) );
  XNOR U665 ( .A(n9524), .B(n8723), .Z(n665) );
  XNOR U666 ( .A(n9521), .B(n8698), .Z(n666) );
  XNOR U667 ( .A(n9526), .B(n8722), .Z(n667) );
  XNOR U668 ( .A(n9522), .B(n8692), .Z(n668) );
  XNOR U669 ( .A(n9527), .B(n8716), .Z(n669) );
  XNOR U670 ( .A(n9519), .B(n8689), .Z(n670) );
  XNOR U671 ( .A(n8614), .B(n8613), .Z(n671) );
  XNOR U672 ( .A(n8638), .B(n8637), .Z(n672) );
  XNOR U673 ( .A(n8611), .B(n8610), .Z(n673) );
  XNOR U674 ( .A(n8635), .B(n8634), .Z(n674) );
  XNOR U675 ( .A(n8605), .B(n8604), .Z(n675) );
  XNOR U676 ( .A(n8629), .B(n8628), .Z(n676) );
  XNOR U677 ( .A(n9499), .B(n8603), .Z(n677) );
  XNOR U678 ( .A(n9504), .B(n8627), .Z(n678) );
  XNOR U679 ( .A(n9501), .B(n8602), .Z(n679) );
  XNOR U680 ( .A(n9506), .B(n8626), .Z(n680) );
  XNOR U681 ( .A(n9502), .B(n8596), .Z(n681) );
  XNOR U682 ( .A(n9507), .B(n8620), .Z(n682) );
  XNOR U683 ( .A(n9499), .B(n8593), .Z(n683) );
  XNOR U684 ( .A(n8518), .B(n8517), .Z(n684) );
  XNOR U685 ( .A(n8542), .B(n8541), .Z(n685) );
  XNOR U686 ( .A(n8515), .B(n8514), .Z(n686) );
  XNOR U687 ( .A(n8539), .B(n8538), .Z(n687) );
  XNOR U688 ( .A(n8509), .B(n8508), .Z(n688) );
  XNOR U689 ( .A(n8533), .B(n8532), .Z(n689) );
  XNOR U690 ( .A(n9479), .B(n8507), .Z(n690) );
  XNOR U691 ( .A(n9484), .B(n8531), .Z(n691) );
  XNOR U692 ( .A(n9481), .B(n8506), .Z(n692) );
  XNOR U693 ( .A(n9486), .B(n8530), .Z(n693) );
  XNOR U694 ( .A(n9482), .B(n8500), .Z(n694) );
  XNOR U695 ( .A(n9487), .B(n8524), .Z(n695) );
  XNOR U696 ( .A(n9479), .B(n8497), .Z(n696) );
  XNOR U697 ( .A(n10086), .B(n10085), .Z(n697) );
  XNOR U698 ( .A(n9726), .B(n9725), .Z(n698) );
  XNOR U699 ( .A(n10083), .B(n10082), .Z(n699) );
  XNOR U700 ( .A(n9723), .B(n9722), .Z(n700) );
  XNOR U701 ( .A(n10077), .B(n10076), .Z(n701) );
  XNOR U702 ( .A(n9717), .B(n9716), .Z(n702) );
  XNOR U703 ( .A(n10819), .B(n10075), .Z(n703) );
  XNOR U704 ( .A(n10744), .B(n9715), .Z(n704) );
  XNOR U705 ( .A(n10821), .B(n10074), .Z(n705) );
  XNOR U706 ( .A(n10746), .B(n9714), .Z(n706) );
  XNOR U707 ( .A(n10822), .B(n10068), .Z(n707) );
  XNOR U708 ( .A(n10747), .B(n9708), .Z(n708) );
  XNOR U709 ( .A(n10819), .B(n10065), .Z(n709) );
  XNOR U710 ( .A(n9990), .B(n9989), .Z(n710) );
  XNOR U711 ( .A(n10014), .B(n10013), .Z(n711) );
  XNOR U712 ( .A(n9987), .B(n9986), .Z(n712) );
  XNOR U713 ( .A(n10011), .B(n10010), .Z(n713) );
  XNOR U714 ( .A(n9981), .B(n9980), .Z(n714) );
  XNOR U715 ( .A(n10005), .B(n10004), .Z(n715) );
  XNOR U716 ( .A(n10799), .B(n9979), .Z(n716) );
  XNOR U717 ( .A(n10804), .B(n10003), .Z(n717) );
  XNOR U718 ( .A(n10801), .B(n9978), .Z(n718) );
  XNOR U719 ( .A(n10806), .B(n10002), .Z(n719) );
  XNOR U720 ( .A(n10802), .B(n9972), .Z(n720) );
  XNOR U721 ( .A(n10807), .B(n9996), .Z(n721) );
  XNOR U722 ( .A(n10799), .B(n9969), .Z(n722) );
  XNOR U723 ( .A(n9894), .B(n9893), .Z(n723) );
  XNOR U724 ( .A(n9918), .B(n9917), .Z(n724) );
  XNOR U725 ( .A(n9891), .B(n9890), .Z(n725) );
  XNOR U726 ( .A(n9915), .B(n9914), .Z(n726) );
  XNOR U727 ( .A(n9885), .B(n9884), .Z(n727) );
  XNOR U728 ( .A(n9909), .B(n9908), .Z(n728) );
  XNOR U729 ( .A(n10779), .B(n9883), .Z(n729) );
  XNOR U730 ( .A(n10784), .B(n9907), .Z(n730) );
  XNOR U731 ( .A(n10781), .B(n9882), .Z(n731) );
  XNOR U732 ( .A(n10786), .B(n9906), .Z(n732) );
  XNOR U733 ( .A(n10782), .B(n9876), .Z(n733) );
  XNOR U734 ( .A(n10787), .B(n9900), .Z(n734) );
  XNOR U735 ( .A(n10779), .B(n9873), .Z(n735) );
  XNOR U736 ( .A(n9798), .B(n9797), .Z(n736) );
  XNOR U737 ( .A(n9822), .B(n9821), .Z(n737) );
  XNOR U738 ( .A(n9795), .B(n9794), .Z(n738) );
  XNOR U739 ( .A(n9819), .B(n9818), .Z(n739) );
  XNOR U740 ( .A(n9789), .B(n9788), .Z(n740) );
  XNOR U741 ( .A(n9813), .B(n9812), .Z(n741) );
  XNOR U742 ( .A(n10759), .B(n9787), .Z(n742) );
  XNOR U743 ( .A(n10764), .B(n9811), .Z(n743) );
  XNOR U744 ( .A(n10761), .B(n9786), .Z(n744) );
  XNOR U745 ( .A(n10766), .B(n9810), .Z(n745) );
  XNOR U746 ( .A(n10762), .B(n9780), .Z(n746) );
  XNOR U747 ( .A(n10767), .B(n9804), .Z(n747) );
  XNOR U748 ( .A(n10759), .B(n9777), .Z(n748) );
  XNOR U749 ( .A(n11366), .B(n11365), .Z(n749) );
  XNOR U750 ( .A(n11006), .B(n11005), .Z(n750) );
  XNOR U751 ( .A(n11363), .B(n11362), .Z(n751) );
  XNOR U752 ( .A(n11003), .B(n11002), .Z(n752) );
  XNOR U753 ( .A(n11357), .B(n11356), .Z(n753) );
  XNOR U754 ( .A(n10997), .B(n10996), .Z(n754) );
  XNOR U755 ( .A(n12099), .B(n11355), .Z(n755) );
  XNOR U756 ( .A(n12024), .B(n10995), .Z(n756) );
  XNOR U757 ( .A(n12101), .B(n11354), .Z(n757) );
  XNOR U758 ( .A(n12026), .B(n10994), .Z(n758) );
  XNOR U759 ( .A(n12102), .B(n11348), .Z(n759) );
  XNOR U760 ( .A(n12027), .B(n10988), .Z(n760) );
  XNOR U761 ( .A(n12099), .B(n11345), .Z(n761) );
  XNOR U762 ( .A(n11270), .B(n11269), .Z(n762) );
  XNOR U763 ( .A(n11294), .B(n11293), .Z(n763) );
  XNOR U764 ( .A(n11267), .B(n11266), .Z(n764) );
  XNOR U765 ( .A(n11291), .B(n11290), .Z(n765) );
  XNOR U766 ( .A(n11261), .B(n11260), .Z(n766) );
  XNOR U767 ( .A(n11285), .B(n11284), .Z(n767) );
  XNOR U768 ( .A(n12079), .B(n11259), .Z(n768) );
  XNOR U769 ( .A(n12084), .B(n11283), .Z(n769) );
  XNOR U770 ( .A(n12081), .B(n11258), .Z(n770) );
  XNOR U771 ( .A(n12086), .B(n11282), .Z(n771) );
  XNOR U772 ( .A(n12082), .B(n11252), .Z(n772) );
  XNOR U773 ( .A(n12087), .B(n11276), .Z(n773) );
  XNOR U774 ( .A(n12079), .B(n11249), .Z(n774) );
  XNOR U775 ( .A(n11174), .B(n11173), .Z(n775) );
  XNOR U776 ( .A(n11198), .B(n11197), .Z(n776) );
  XNOR U777 ( .A(n11171), .B(n11170), .Z(n777) );
  XNOR U778 ( .A(n11195), .B(n11194), .Z(n778) );
  XNOR U779 ( .A(n11165), .B(n11164), .Z(n779) );
  XNOR U780 ( .A(n11189), .B(n11188), .Z(n780) );
  XNOR U781 ( .A(n12059), .B(n11163), .Z(n781) );
  XNOR U782 ( .A(n12064), .B(n11187), .Z(n782) );
  XNOR U783 ( .A(n12061), .B(n11162), .Z(n783) );
  XNOR U784 ( .A(n12066), .B(n11186), .Z(n784) );
  XNOR U785 ( .A(n12062), .B(n11156), .Z(n785) );
  XNOR U786 ( .A(n12067), .B(n11180), .Z(n786) );
  XNOR U787 ( .A(n12059), .B(n11153), .Z(n787) );
  XNOR U788 ( .A(n11078), .B(n11077), .Z(n788) );
  XNOR U789 ( .A(n11102), .B(n11101), .Z(n789) );
  XNOR U790 ( .A(n11075), .B(n11074), .Z(n790) );
  XNOR U791 ( .A(n11099), .B(n11098), .Z(n791) );
  XNOR U792 ( .A(n11069), .B(n11068), .Z(n792) );
  XNOR U793 ( .A(n11093), .B(n11092), .Z(n793) );
  XNOR U794 ( .A(n12039), .B(n11067), .Z(n794) );
  XNOR U795 ( .A(n12044), .B(n11091), .Z(n795) );
  XNOR U796 ( .A(n12041), .B(n11066), .Z(n796) );
  XNOR U797 ( .A(n12046), .B(n11090), .Z(n797) );
  XNOR U798 ( .A(n12042), .B(n11060), .Z(n798) );
  XNOR U799 ( .A(n12047), .B(n11084), .Z(n799) );
  XNOR U800 ( .A(n12039), .B(n11057), .Z(n800) );
  XNOR U801 ( .A(n12646), .B(n12645), .Z(n801) );
  XNOR U802 ( .A(n12286), .B(n12285), .Z(n802) );
  XNOR U803 ( .A(n12643), .B(n12642), .Z(n803) );
  XNOR U804 ( .A(n12283), .B(n12282), .Z(n804) );
  XNOR U805 ( .A(n12637), .B(n12636), .Z(n805) );
  XNOR U806 ( .A(n12277), .B(n12276), .Z(n806) );
  XNOR U807 ( .A(n13379), .B(n12635), .Z(n807) );
  XNOR U808 ( .A(n13304), .B(n12275), .Z(n808) );
  XNOR U809 ( .A(n13381), .B(n12634), .Z(n809) );
  XNOR U810 ( .A(n13306), .B(n12274), .Z(n810) );
  XNOR U811 ( .A(n13382), .B(n12628), .Z(n811) );
  XNOR U812 ( .A(n13307), .B(n12268), .Z(n812) );
  XNOR U813 ( .A(n13379), .B(n12625), .Z(n813) );
  XNOR U814 ( .A(n12550), .B(n12549), .Z(n814) );
  XNOR U815 ( .A(n12574), .B(n12573), .Z(n815) );
  XNOR U816 ( .A(n12547), .B(n12546), .Z(n816) );
  XNOR U817 ( .A(n12571), .B(n12570), .Z(n817) );
  XNOR U818 ( .A(n12541), .B(n12540), .Z(n818) );
  XNOR U819 ( .A(n12565), .B(n12564), .Z(n819) );
  XNOR U820 ( .A(n13359), .B(n12539), .Z(n820) );
  XNOR U821 ( .A(n13364), .B(n12563), .Z(n821) );
  XNOR U822 ( .A(n13361), .B(n12538), .Z(n822) );
  XNOR U823 ( .A(n13366), .B(n12562), .Z(n823) );
  XNOR U824 ( .A(n13362), .B(n12532), .Z(n824) );
  XNOR U825 ( .A(n13367), .B(n12556), .Z(n825) );
  XNOR U826 ( .A(n13359), .B(n12529), .Z(n826) );
  XNOR U827 ( .A(n12454), .B(n12453), .Z(n827) );
  XNOR U828 ( .A(n12478), .B(n12477), .Z(n828) );
  XNOR U829 ( .A(n12451), .B(n12450), .Z(n829) );
  XNOR U830 ( .A(n12475), .B(n12474), .Z(n830) );
  XNOR U831 ( .A(n12445), .B(n12444), .Z(n831) );
  XNOR U832 ( .A(n12469), .B(n12468), .Z(n832) );
  XNOR U833 ( .A(n13339), .B(n12443), .Z(n833) );
  XNOR U834 ( .A(n13344), .B(n12467), .Z(n834) );
  XNOR U835 ( .A(n13341), .B(n12442), .Z(n835) );
  XNOR U836 ( .A(n13346), .B(n12466), .Z(n836) );
  XNOR U837 ( .A(n13342), .B(n12436), .Z(n837) );
  XNOR U838 ( .A(n13347), .B(n12460), .Z(n838) );
  XNOR U839 ( .A(n13339), .B(n12433), .Z(n839) );
  XNOR U840 ( .A(n12358), .B(n12357), .Z(n840) );
  XNOR U841 ( .A(n12382), .B(n12381), .Z(n841) );
  XNOR U842 ( .A(n12355), .B(n12354), .Z(n842) );
  XNOR U843 ( .A(n12379), .B(n12378), .Z(n843) );
  XNOR U844 ( .A(n12349), .B(n12348), .Z(n844) );
  XNOR U845 ( .A(n12373), .B(n12372), .Z(n845) );
  XNOR U846 ( .A(n13319), .B(n12347), .Z(n846) );
  XNOR U847 ( .A(n13324), .B(n12371), .Z(n847) );
  XNOR U848 ( .A(n13321), .B(n12346), .Z(n848) );
  XNOR U849 ( .A(n13326), .B(n12370), .Z(n849) );
  XNOR U850 ( .A(n13322), .B(n12340), .Z(n850) );
  XNOR U851 ( .A(n13327), .B(n12364), .Z(n851) );
  XNOR U852 ( .A(n13319), .B(n12337), .Z(n852) );
  XNOR U853 ( .A(n13926), .B(n13925), .Z(n853) );
  XNOR U854 ( .A(n13566), .B(n13565), .Z(n854) );
  XNOR U855 ( .A(n13923), .B(n13922), .Z(n855) );
  XNOR U856 ( .A(n13563), .B(n13562), .Z(n856) );
  XNOR U857 ( .A(n13917), .B(n13916), .Z(n857) );
  XNOR U858 ( .A(n13557), .B(n13556), .Z(n858) );
  XNOR U859 ( .A(n14659), .B(n13915), .Z(n859) );
  XNOR U860 ( .A(n14584), .B(n13555), .Z(n860) );
  XNOR U861 ( .A(n14661), .B(n13914), .Z(n861) );
  XNOR U862 ( .A(n14586), .B(n13554), .Z(n862) );
  XNOR U863 ( .A(n14662), .B(n13908), .Z(n863) );
  XNOR U864 ( .A(n14587), .B(n13548), .Z(n864) );
  XNOR U865 ( .A(n14659), .B(n13905), .Z(n865) );
  XNOR U866 ( .A(n13830), .B(n13829), .Z(n866) );
  XNOR U867 ( .A(n13854), .B(n13853), .Z(n867) );
  XNOR U868 ( .A(n13827), .B(n13826), .Z(n868) );
  XNOR U869 ( .A(n13851), .B(n13850), .Z(n869) );
  XNOR U870 ( .A(n13821), .B(n13820), .Z(n870) );
  XNOR U871 ( .A(n13845), .B(n13844), .Z(n871) );
  XNOR U872 ( .A(n14639), .B(n13819), .Z(n872) );
  XNOR U873 ( .A(n14644), .B(n13843), .Z(n873) );
  XNOR U874 ( .A(n14641), .B(n13818), .Z(n874) );
  XNOR U875 ( .A(n14646), .B(n13842), .Z(n875) );
  XNOR U876 ( .A(n14642), .B(n13812), .Z(n876) );
  XNOR U877 ( .A(n14647), .B(n13836), .Z(n877) );
  XNOR U878 ( .A(n14639), .B(n13809), .Z(n878) );
  XNOR U879 ( .A(n13734), .B(n13733), .Z(n879) );
  XNOR U880 ( .A(n13758), .B(n13757), .Z(n880) );
  XNOR U881 ( .A(n13731), .B(n13730), .Z(n881) );
  XNOR U882 ( .A(n13755), .B(n13754), .Z(n882) );
  XNOR U883 ( .A(n13725), .B(n13724), .Z(n883) );
  XNOR U884 ( .A(n13749), .B(n13748), .Z(n884) );
  XNOR U885 ( .A(n14619), .B(n13723), .Z(n885) );
  XNOR U886 ( .A(n14624), .B(n13747), .Z(n886) );
  XNOR U887 ( .A(n14621), .B(n13722), .Z(n887) );
  XNOR U888 ( .A(n14626), .B(n13746), .Z(n888) );
  XNOR U889 ( .A(n14622), .B(n13716), .Z(n889) );
  XNOR U890 ( .A(n14627), .B(n13740), .Z(n890) );
  XNOR U891 ( .A(n14619), .B(n13713), .Z(n891) );
  XNOR U892 ( .A(n13638), .B(n13637), .Z(n892) );
  XNOR U893 ( .A(n13662), .B(n13661), .Z(n893) );
  XNOR U894 ( .A(n13635), .B(n13634), .Z(n894) );
  XNOR U895 ( .A(n13659), .B(n13658), .Z(n895) );
  XNOR U896 ( .A(n13629), .B(n13628), .Z(n896) );
  XNOR U897 ( .A(n13653), .B(n13652), .Z(n897) );
  XNOR U898 ( .A(n14599), .B(n13627), .Z(n898) );
  XNOR U899 ( .A(n14604), .B(n13651), .Z(n899) );
  XNOR U900 ( .A(n14601), .B(n13626), .Z(n900) );
  XNOR U901 ( .A(n14606), .B(n13650), .Z(n901) );
  XNOR U902 ( .A(n14602), .B(n13620), .Z(n902) );
  XNOR U903 ( .A(n14607), .B(n13644), .Z(n903) );
  XNOR U904 ( .A(n14599), .B(n13617), .Z(n904) );
  XNOR U905 ( .A(n15206), .B(n15205), .Z(n905) );
  XNOR U906 ( .A(n14846), .B(n14845), .Z(n906) );
  XNOR U907 ( .A(n15203), .B(n15202), .Z(n907) );
  XNOR U908 ( .A(n14843), .B(n14842), .Z(n908) );
  XNOR U909 ( .A(n15197), .B(n15196), .Z(n909) );
  XNOR U910 ( .A(n14837), .B(n14836), .Z(n910) );
  XNOR U911 ( .A(n15939), .B(n15195), .Z(n911) );
  XNOR U912 ( .A(n15864), .B(n14835), .Z(n912) );
  XNOR U913 ( .A(n15941), .B(n15194), .Z(n913) );
  XNOR U914 ( .A(n15866), .B(n14834), .Z(n914) );
  XNOR U915 ( .A(n15942), .B(n15188), .Z(n915) );
  XNOR U916 ( .A(n15867), .B(n14828), .Z(n916) );
  XNOR U917 ( .A(n15939), .B(n15185), .Z(n917) );
  XNOR U918 ( .A(n15110), .B(n15109), .Z(n918) );
  XNOR U919 ( .A(n15134), .B(n15133), .Z(n919) );
  XNOR U920 ( .A(n15107), .B(n15106), .Z(n920) );
  XNOR U921 ( .A(n15131), .B(n15130), .Z(n921) );
  XNOR U922 ( .A(n15101), .B(n15100), .Z(n922) );
  XNOR U923 ( .A(n15125), .B(n15124), .Z(n923) );
  XNOR U924 ( .A(n15919), .B(n15099), .Z(n924) );
  XNOR U925 ( .A(n15924), .B(n15123), .Z(n925) );
  XNOR U926 ( .A(n15921), .B(n15098), .Z(n926) );
  XNOR U927 ( .A(n15926), .B(n15122), .Z(n927) );
  XNOR U928 ( .A(n15922), .B(n15092), .Z(n928) );
  XNOR U929 ( .A(n15927), .B(n15116), .Z(n929) );
  XNOR U930 ( .A(n15919), .B(n15089), .Z(n930) );
  XNOR U931 ( .A(n15014), .B(n15013), .Z(n931) );
  XNOR U932 ( .A(n15038), .B(n15037), .Z(n932) );
  XNOR U933 ( .A(n15011), .B(n15010), .Z(n933) );
  XNOR U934 ( .A(n15035), .B(n15034), .Z(n934) );
  XNOR U935 ( .A(n15005), .B(n15004), .Z(n935) );
  XNOR U936 ( .A(n15029), .B(n15028), .Z(n936) );
  XNOR U937 ( .A(n15899), .B(n15003), .Z(n937) );
  XNOR U938 ( .A(n15904), .B(n15027), .Z(n938) );
  XNOR U939 ( .A(n15901), .B(n15002), .Z(n939) );
  XNOR U940 ( .A(n15906), .B(n15026), .Z(n940) );
  XNOR U941 ( .A(n15902), .B(n14996), .Z(n941) );
  XNOR U942 ( .A(n15907), .B(n15020), .Z(n942) );
  XNOR U943 ( .A(n15899), .B(n14993), .Z(n943) );
  XNOR U944 ( .A(n14918), .B(n14917), .Z(n944) );
  XNOR U945 ( .A(n14942), .B(n14941), .Z(n945) );
  XNOR U946 ( .A(n14915), .B(n14914), .Z(n946) );
  XNOR U947 ( .A(n14939), .B(n14938), .Z(n947) );
  XNOR U948 ( .A(n14909), .B(n14908), .Z(n948) );
  XNOR U949 ( .A(n14933), .B(n14932), .Z(n949) );
  XNOR U950 ( .A(n15879), .B(n14907), .Z(n950) );
  XNOR U951 ( .A(n15884), .B(n14931), .Z(n951) );
  XNOR U952 ( .A(n15881), .B(n14906), .Z(n952) );
  XNOR U953 ( .A(n15886), .B(n14930), .Z(n953) );
  XNOR U954 ( .A(n15882), .B(n14900), .Z(n954) );
  XNOR U955 ( .A(n15887), .B(n14924), .Z(n955) );
  XNOR U956 ( .A(n15879), .B(n14897), .Z(n956) );
  AND U957 ( .A(\SUBBYTES[1].a/w209 ), .B(\SUBBYTES[1].a/w222 ), .Z(n957) );
  AND U958 ( .A(\SUBBYTES[1].a/w416 ), .B(\SUBBYTES[1].a/w429 ), .Z(n958) );
  AND U959 ( .A(\SUBBYTES[1].a/w623 ), .B(\SUBBYTES[1].a/w636 ), .Z(n959) );
  AND U960 ( .A(\SUBBYTES[1].a/w830 ), .B(\SUBBYTES[1].a/w843 ), .Z(n960) );
  AND U961 ( .A(\SUBBYTES[1].a/w1037 ), .B(\SUBBYTES[1].a/w1050 ), .Z(n961) );
  AND U962 ( .A(\SUBBYTES[1].a/w1244 ), .B(\SUBBYTES[1].a/w1257 ), .Z(n962) );
  AND U963 ( .A(\SUBBYTES[1].a/w1451 ), .B(\SUBBYTES[1].a/w1464 ), .Z(n963) );
  AND U964 ( .A(\SUBBYTES[1].a/w1658 ), .B(\SUBBYTES[1].a/w1671 ), .Z(n964) );
  AND U965 ( .A(\SUBBYTES[1].a/w1865 ), .B(\SUBBYTES[1].a/w1878 ), .Z(n965) );
  AND U966 ( .A(\SUBBYTES[1].a/w2072 ), .B(\SUBBYTES[1].a/w2085 ), .Z(n966) );
  AND U967 ( .A(\SUBBYTES[1].a/w2279 ), .B(\SUBBYTES[1].a/w2292 ), .Z(n967) );
  AND U968 ( .A(\SUBBYTES[1].a/w2486 ), .B(\SUBBYTES[1].a/w2499 ), .Z(n968) );
  AND U969 ( .A(\SUBBYTES[1].a/w2693 ), .B(\SUBBYTES[1].a/w2706 ), .Z(n969) );
  AND U970 ( .A(\SUBBYTES[1].a/w2900 ), .B(\SUBBYTES[1].a/w2913 ), .Z(n970) );
  AND U971 ( .A(\SUBBYTES[1].a/w3107 ), .B(\SUBBYTES[1].a/w3120 ), .Z(n971) );
  AND U972 ( .A(\SUBBYTES[1].a/w3314 ), .B(\SUBBYTES[1].a/w3327 ), .Z(n972) );
  AND U973 ( .A(\SUBBYTES[2].a/w209 ), .B(\SUBBYTES[2].a/w222 ), .Z(n973) );
  AND U974 ( .A(\SUBBYTES[2].a/w416 ), .B(\SUBBYTES[2].a/w429 ), .Z(n974) );
  AND U975 ( .A(\SUBBYTES[2].a/w623 ), .B(\SUBBYTES[2].a/w636 ), .Z(n975) );
  AND U976 ( .A(\SUBBYTES[2].a/w830 ), .B(\SUBBYTES[2].a/w843 ), .Z(n976) );
  AND U977 ( .A(\SUBBYTES[2].a/w1037 ), .B(\SUBBYTES[2].a/w1050 ), .Z(n977) );
  AND U978 ( .A(\SUBBYTES[2].a/w1244 ), .B(\SUBBYTES[2].a/w1257 ), .Z(n978) );
  AND U979 ( .A(\SUBBYTES[2].a/w1451 ), .B(\SUBBYTES[2].a/w1464 ), .Z(n979) );
  AND U980 ( .A(\SUBBYTES[2].a/w1658 ), .B(\SUBBYTES[2].a/w1671 ), .Z(n980) );
  AND U981 ( .A(\SUBBYTES[2].a/w1865 ), .B(\SUBBYTES[2].a/w1878 ), .Z(n981) );
  AND U982 ( .A(\SUBBYTES[2].a/w2072 ), .B(\SUBBYTES[2].a/w2085 ), .Z(n982) );
  AND U983 ( .A(\SUBBYTES[2].a/w2279 ), .B(\SUBBYTES[2].a/w2292 ), .Z(n983) );
  AND U984 ( .A(\SUBBYTES[2].a/w2486 ), .B(\SUBBYTES[2].a/w2499 ), .Z(n984) );
  AND U985 ( .A(\SUBBYTES[2].a/w2693 ), .B(\SUBBYTES[2].a/w2706 ), .Z(n985) );
  AND U986 ( .A(\SUBBYTES[2].a/w2900 ), .B(\SUBBYTES[2].a/w2913 ), .Z(n986) );
  AND U987 ( .A(\SUBBYTES[2].a/w3107 ), .B(\SUBBYTES[2].a/w3120 ), .Z(n987) );
  AND U988 ( .A(\SUBBYTES[2].a/w3314 ), .B(\SUBBYTES[2].a/w3327 ), .Z(n988) );
  AND U989 ( .A(\SUBBYTES[3].a/w209 ), .B(\SUBBYTES[3].a/w222 ), .Z(n989) );
  AND U990 ( .A(\SUBBYTES[3].a/w416 ), .B(\SUBBYTES[3].a/w429 ), .Z(n990) );
  AND U991 ( .A(\SUBBYTES[3].a/w623 ), .B(\SUBBYTES[3].a/w636 ), .Z(n991) );
  AND U992 ( .A(\SUBBYTES[3].a/w830 ), .B(\SUBBYTES[3].a/w843 ), .Z(n992) );
  AND U993 ( .A(\SUBBYTES[3].a/w1037 ), .B(\SUBBYTES[3].a/w1050 ), .Z(n993) );
  AND U994 ( .A(\SUBBYTES[3].a/w1244 ), .B(\SUBBYTES[3].a/w1257 ), .Z(n994) );
  AND U995 ( .A(\SUBBYTES[3].a/w1451 ), .B(\SUBBYTES[3].a/w1464 ), .Z(n995) );
  AND U996 ( .A(\SUBBYTES[3].a/w1658 ), .B(\SUBBYTES[3].a/w1671 ), .Z(n996) );
  AND U997 ( .A(\SUBBYTES[3].a/w1865 ), .B(\SUBBYTES[3].a/w1878 ), .Z(n997) );
  AND U998 ( .A(\SUBBYTES[3].a/w2072 ), .B(\SUBBYTES[3].a/w2085 ), .Z(n998) );
  AND U999 ( .A(\SUBBYTES[3].a/w2279 ), .B(\SUBBYTES[3].a/w2292 ), .Z(n999) );
  AND U1000 ( .A(\SUBBYTES[3].a/w2486 ), .B(\SUBBYTES[3].a/w2499 ), .Z(n1000)
         );
  AND U1001 ( .A(\SUBBYTES[3].a/w2693 ), .B(\SUBBYTES[3].a/w2706 ), .Z(n1001)
         );
  AND U1002 ( .A(\SUBBYTES[3].a/w2900 ), .B(\SUBBYTES[3].a/w2913 ), .Z(n1002)
         );
  AND U1003 ( .A(\SUBBYTES[3].a/w3107 ), .B(\SUBBYTES[3].a/w3120 ), .Z(n1003)
         );
  AND U1004 ( .A(\SUBBYTES[3].a/w3314 ), .B(\SUBBYTES[3].a/w3327 ), .Z(n1004)
         );
  AND U1005 ( .A(\SUBBYTES[4].a/w209 ), .B(\SUBBYTES[4].a/w222 ), .Z(n1005) );
  AND U1006 ( .A(\SUBBYTES[4].a/w416 ), .B(\SUBBYTES[4].a/w429 ), .Z(n1006) );
  AND U1007 ( .A(\SUBBYTES[4].a/w623 ), .B(\SUBBYTES[4].a/w636 ), .Z(n1007) );
  AND U1008 ( .A(\SUBBYTES[4].a/w830 ), .B(\SUBBYTES[4].a/w843 ), .Z(n1008) );
  AND U1009 ( .A(\SUBBYTES[4].a/w1037 ), .B(\SUBBYTES[4].a/w1050 ), .Z(n1009)
         );
  AND U1010 ( .A(\SUBBYTES[4].a/w1244 ), .B(\SUBBYTES[4].a/w1257 ), .Z(n1010)
         );
  AND U1011 ( .A(\SUBBYTES[4].a/w1451 ), .B(\SUBBYTES[4].a/w1464 ), .Z(n1011)
         );
  AND U1012 ( .A(\SUBBYTES[4].a/w1658 ), .B(\SUBBYTES[4].a/w1671 ), .Z(n1012)
         );
  AND U1013 ( .A(\SUBBYTES[4].a/w1865 ), .B(\SUBBYTES[4].a/w1878 ), .Z(n1013)
         );
  AND U1014 ( .A(\SUBBYTES[4].a/w2072 ), .B(\SUBBYTES[4].a/w2085 ), .Z(n1014)
         );
  AND U1015 ( .A(\SUBBYTES[4].a/w2279 ), .B(\SUBBYTES[4].a/w2292 ), .Z(n1015)
         );
  AND U1016 ( .A(\SUBBYTES[4].a/w2486 ), .B(\SUBBYTES[4].a/w2499 ), .Z(n1016)
         );
  AND U1017 ( .A(\SUBBYTES[4].a/w2693 ), .B(\SUBBYTES[4].a/w2706 ), .Z(n1017)
         );
  AND U1018 ( .A(\SUBBYTES[4].a/w2900 ), .B(\SUBBYTES[4].a/w2913 ), .Z(n1018)
         );
  AND U1019 ( .A(\SUBBYTES[4].a/w3107 ), .B(\SUBBYTES[4].a/w3120 ), .Z(n1019)
         );
  AND U1020 ( .A(\SUBBYTES[4].a/w3314 ), .B(\SUBBYTES[4].a/w3327 ), .Z(n1020)
         );
  AND U1021 ( .A(\SUBBYTES[5].a/w209 ), .B(\SUBBYTES[5].a/w222 ), .Z(n1021) );
  AND U1022 ( .A(\SUBBYTES[5].a/w416 ), .B(\SUBBYTES[5].a/w429 ), .Z(n1022) );
  AND U1023 ( .A(\SUBBYTES[5].a/w623 ), .B(\SUBBYTES[5].a/w636 ), .Z(n1023) );
  AND U1024 ( .A(\SUBBYTES[5].a/w830 ), .B(\SUBBYTES[5].a/w843 ), .Z(n1024) );
  AND U1025 ( .A(\SUBBYTES[5].a/w1037 ), .B(\SUBBYTES[5].a/w1050 ), .Z(n1025)
         );
  AND U1026 ( .A(\SUBBYTES[5].a/w1244 ), .B(\SUBBYTES[5].a/w1257 ), .Z(n1026)
         );
  AND U1027 ( .A(\SUBBYTES[5].a/w1451 ), .B(\SUBBYTES[5].a/w1464 ), .Z(n1027)
         );
  AND U1028 ( .A(\SUBBYTES[5].a/w1658 ), .B(\SUBBYTES[5].a/w1671 ), .Z(n1028)
         );
  AND U1029 ( .A(\SUBBYTES[5].a/w1865 ), .B(\SUBBYTES[5].a/w1878 ), .Z(n1029)
         );
  AND U1030 ( .A(\SUBBYTES[5].a/w2072 ), .B(\SUBBYTES[5].a/w2085 ), .Z(n1030)
         );
  AND U1031 ( .A(\SUBBYTES[5].a/w2279 ), .B(\SUBBYTES[5].a/w2292 ), .Z(n1031)
         );
  AND U1032 ( .A(\SUBBYTES[5].a/w2486 ), .B(\SUBBYTES[5].a/w2499 ), .Z(n1032)
         );
  AND U1033 ( .A(\SUBBYTES[5].a/w2693 ), .B(\SUBBYTES[5].a/w2706 ), .Z(n1033)
         );
  AND U1034 ( .A(\SUBBYTES[5].a/w2900 ), .B(\SUBBYTES[5].a/w2913 ), .Z(n1034)
         );
  AND U1035 ( .A(\SUBBYTES[5].a/w3107 ), .B(\SUBBYTES[5].a/w3120 ), .Z(n1035)
         );
  AND U1036 ( .A(\SUBBYTES[5].a/w3314 ), .B(\SUBBYTES[5].a/w3327 ), .Z(n1036)
         );
  AND U1037 ( .A(\SUBBYTES[6].a/w209 ), .B(\SUBBYTES[6].a/w222 ), .Z(n1037) );
  AND U1038 ( .A(\SUBBYTES[6].a/w416 ), .B(\SUBBYTES[6].a/w429 ), .Z(n1038) );
  AND U1039 ( .A(\SUBBYTES[6].a/w623 ), .B(\SUBBYTES[6].a/w636 ), .Z(n1039) );
  AND U1040 ( .A(\SUBBYTES[6].a/w830 ), .B(\SUBBYTES[6].a/w843 ), .Z(n1040) );
  AND U1041 ( .A(\SUBBYTES[6].a/w1037 ), .B(\SUBBYTES[6].a/w1050 ), .Z(n1041)
         );
  AND U1042 ( .A(\SUBBYTES[6].a/w1244 ), .B(\SUBBYTES[6].a/w1257 ), .Z(n1042)
         );
  AND U1043 ( .A(\SUBBYTES[6].a/w1451 ), .B(\SUBBYTES[6].a/w1464 ), .Z(n1043)
         );
  AND U1044 ( .A(\SUBBYTES[6].a/w1658 ), .B(\SUBBYTES[6].a/w1671 ), .Z(n1044)
         );
  AND U1045 ( .A(\SUBBYTES[6].a/w1865 ), .B(\SUBBYTES[6].a/w1878 ), .Z(n1045)
         );
  AND U1046 ( .A(\SUBBYTES[6].a/w2072 ), .B(\SUBBYTES[6].a/w2085 ), .Z(n1046)
         );
  AND U1047 ( .A(\SUBBYTES[6].a/w2279 ), .B(\SUBBYTES[6].a/w2292 ), .Z(n1047)
         );
  AND U1048 ( .A(\SUBBYTES[6].a/w2486 ), .B(\SUBBYTES[6].a/w2499 ), .Z(n1048)
         );
  AND U1049 ( .A(\SUBBYTES[6].a/w2693 ), .B(\SUBBYTES[6].a/w2706 ), .Z(n1049)
         );
  AND U1050 ( .A(\SUBBYTES[6].a/w2900 ), .B(\SUBBYTES[6].a/w2913 ), .Z(n1050)
         );
  AND U1051 ( .A(\SUBBYTES[6].a/w3107 ), .B(\SUBBYTES[6].a/w3120 ), .Z(n1051)
         );
  AND U1052 ( .A(\SUBBYTES[6].a/w3314 ), .B(\SUBBYTES[6].a/w3327 ), .Z(n1052)
         );
  AND U1053 ( .A(\SUBBYTES[7].a/w209 ), .B(\SUBBYTES[7].a/w222 ), .Z(n1053) );
  AND U1054 ( .A(\SUBBYTES[7].a/w416 ), .B(\SUBBYTES[7].a/w429 ), .Z(n1054) );
  AND U1055 ( .A(\SUBBYTES[7].a/w623 ), .B(\SUBBYTES[7].a/w636 ), .Z(n1055) );
  AND U1056 ( .A(\SUBBYTES[7].a/w830 ), .B(\SUBBYTES[7].a/w843 ), .Z(n1056) );
  AND U1057 ( .A(\SUBBYTES[7].a/w1037 ), .B(\SUBBYTES[7].a/w1050 ), .Z(n1057)
         );
  AND U1058 ( .A(\SUBBYTES[7].a/w1244 ), .B(\SUBBYTES[7].a/w1257 ), .Z(n1058)
         );
  AND U1059 ( .A(\SUBBYTES[7].a/w1451 ), .B(\SUBBYTES[7].a/w1464 ), .Z(n1059)
         );
  AND U1060 ( .A(\SUBBYTES[7].a/w1658 ), .B(\SUBBYTES[7].a/w1671 ), .Z(n1060)
         );
  AND U1061 ( .A(\SUBBYTES[7].a/w1865 ), .B(\SUBBYTES[7].a/w1878 ), .Z(n1061)
         );
  AND U1062 ( .A(\SUBBYTES[7].a/w2072 ), .B(\SUBBYTES[7].a/w2085 ), .Z(n1062)
         );
  AND U1063 ( .A(\SUBBYTES[7].a/w2279 ), .B(\SUBBYTES[7].a/w2292 ), .Z(n1063)
         );
  AND U1064 ( .A(\SUBBYTES[7].a/w2486 ), .B(\SUBBYTES[7].a/w2499 ), .Z(n1064)
         );
  AND U1065 ( .A(\SUBBYTES[7].a/w2693 ), .B(\SUBBYTES[7].a/w2706 ), .Z(n1065)
         );
  AND U1066 ( .A(\SUBBYTES[7].a/w2900 ), .B(\SUBBYTES[7].a/w2913 ), .Z(n1066)
         );
  AND U1067 ( .A(\SUBBYTES[7].a/w3107 ), .B(\SUBBYTES[7].a/w3120 ), .Z(n1067)
         );
  AND U1068 ( .A(\SUBBYTES[7].a/w3314 ), .B(\SUBBYTES[7].a/w3327 ), .Z(n1068)
         );
  AND U1069 ( .A(\SUBBYTES[8].a/w209 ), .B(\SUBBYTES[8].a/w222 ), .Z(n1069) );
  AND U1070 ( .A(\SUBBYTES[8].a/w416 ), .B(\SUBBYTES[8].a/w429 ), .Z(n1070) );
  AND U1071 ( .A(\SUBBYTES[8].a/w623 ), .B(\SUBBYTES[8].a/w636 ), .Z(n1071) );
  AND U1072 ( .A(\SUBBYTES[8].a/w830 ), .B(\SUBBYTES[8].a/w843 ), .Z(n1072) );
  AND U1073 ( .A(\SUBBYTES[8].a/w1037 ), .B(\SUBBYTES[8].a/w1050 ), .Z(n1073)
         );
  AND U1074 ( .A(\SUBBYTES[8].a/w1244 ), .B(\SUBBYTES[8].a/w1257 ), .Z(n1074)
         );
  AND U1075 ( .A(\SUBBYTES[8].a/w1451 ), .B(\SUBBYTES[8].a/w1464 ), .Z(n1075)
         );
  AND U1076 ( .A(\SUBBYTES[8].a/w1658 ), .B(\SUBBYTES[8].a/w1671 ), .Z(n1076)
         );
  AND U1077 ( .A(\SUBBYTES[8].a/w1865 ), .B(\SUBBYTES[8].a/w1878 ), .Z(n1077)
         );
  AND U1078 ( .A(\SUBBYTES[8].a/w2072 ), .B(\SUBBYTES[8].a/w2085 ), .Z(n1078)
         );
  AND U1079 ( .A(\SUBBYTES[8].a/w2279 ), .B(\SUBBYTES[8].a/w2292 ), .Z(n1079)
         );
  AND U1080 ( .A(\SUBBYTES[8].a/w2486 ), .B(\SUBBYTES[8].a/w2499 ), .Z(n1080)
         );
  AND U1081 ( .A(\SUBBYTES[8].a/w2693 ), .B(\SUBBYTES[8].a/w2706 ), .Z(n1081)
         );
  AND U1082 ( .A(\SUBBYTES[8].a/w2900 ), .B(\SUBBYTES[8].a/w2913 ), .Z(n1082)
         );
  AND U1083 ( .A(\SUBBYTES[8].a/w3107 ), .B(\SUBBYTES[8].a/w3120 ), .Z(n1083)
         );
  AND U1084 ( .A(\SUBBYTES[8].a/w3314 ), .B(\SUBBYTES[8].a/w3327 ), .Z(n1084)
         );
  AND U1085 ( .A(\SUBBYTES[9].a/w209 ), .B(\SUBBYTES[9].a/w222 ), .Z(n1085) );
  AND U1086 ( .A(\SUBBYTES[9].a/w416 ), .B(\SUBBYTES[9].a/w429 ), .Z(n1086) );
  AND U1087 ( .A(\SUBBYTES[9].a/w623 ), .B(\SUBBYTES[9].a/w636 ), .Z(n1087) );
  AND U1088 ( .A(\SUBBYTES[9].a/w830 ), .B(\SUBBYTES[9].a/w843 ), .Z(n1088) );
  AND U1089 ( .A(\SUBBYTES[9].a/w1037 ), .B(\SUBBYTES[9].a/w1050 ), .Z(n1089)
         );
  AND U1090 ( .A(\SUBBYTES[9].a/w1244 ), .B(\SUBBYTES[9].a/w1257 ), .Z(n1090)
         );
  AND U1091 ( .A(\SUBBYTES[9].a/w1451 ), .B(\SUBBYTES[9].a/w1464 ), .Z(n1091)
         );
  AND U1092 ( .A(\SUBBYTES[9].a/w1658 ), .B(\SUBBYTES[9].a/w1671 ), .Z(n1092)
         );
  AND U1093 ( .A(\SUBBYTES[9].a/w1865 ), .B(\SUBBYTES[9].a/w1878 ), .Z(n1093)
         );
  AND U1094 ( .A(\SUBBYTES[9].a/w2072 ), .B(\SUBBYTES[9].a/w2085 ), .Z(n1094)
         );
  AND U1095 ( .A(\SUBBYTES[9].a/w2279 ), .B(\SUBBYTES[9].a/w2292 ), .Z(n1095)
         );
  AND U1096 ( .A(\SUBBYTES[9].a/w2486 ), .B(\SUBBYTES[9].a/w2499 ), .Z(n1096)
         );
  AND U1097 ( .A(\SUBBYTES[9].a/w2693 ), .B(\SUBBYTES[9].a/w2706 ), .Z(n1097)
         );
  AND U1098 ( .A(\SUBBYTES[9].a/w2900 ), .B(\SUBBYTES[9].a/w2913 ), .Z(n1098)
         );
  AND U1099 ( .A(\SUBBYTES[9].a/w3107 ), .B(\SUBBYTES[9].a/w3120 ), .Z(n1099)
         );
  AND U1100 ( .A(\SUBBYTES[9].a/w3314 ), .B(\SUBBYTES[9].a/w3327 ), .Z(n1100)
         );
  XNOR U1101 ( .A(\SUBBYTES[0].a/n767 ), .B(\SUBBYTES[0].a/n766 ), .Z(n1101)
         );
  XNOR U1102 ( .A(\SUBBYTES[0].a/n407 ), .B(\SUBBYTES[0].a/n406 ), .Z(n1102)
         );
  XNOR U1103 ( .A(\SUBBYTES[0].a/n764 ), .B(\SUBBYTES[0].a/n763 ), .Z(n1103)
         );
  XNOR U1104 ( .A(\SUBBYTES[0].a/n404 ), .B(\SUBBYTES[0].a/n403 ), .Z(n1104)
         );
  XNOR U1105 ( .A(\SUBBYTES[0].a/n758 ), .B(\SUBBYTES[0].a/n757 ), .Z(n1105)
         );
  XNOR U1106 ( .A(\SUBBYTES[0].a/n398 ), .B(\SUBBYTES[0].a/n397 ), .Z(n1106)
         );
  XNOR U1107 ( .A(\SUBBYTES[0].a/n1500 ), .B(\SUBBYTES[0].a/n756 ), .Z(n1107)
         );
  XNOR U1108 ( .A(\SUBBYTES[0].a/n1425 ), .B(\SUBBYTES[0].a/n396 ), .Z(n1108)
         );
  XNOR U1109 ( .A(\SUBBYTES[0].a/n1502 ), .B(\SUBBYTES[0].a/n755 ), .Z(n1109)
         );
  XNOR U1110 ( .A(\SUBBYTES[0].a/n1427 ), .B(\SUBBYTES[0].a/n395 ), .Z(n1110)
         );
  XNOR U1111 ( .A(\SUBBYTES[0].a/n1503 ), .B(\SUBBYTES[0].a/n749 ), .Z(n1111)
         );
  XNOR U1112 ( .A(\SUBBYTES[0].a/n1428 ), .B(\SUBBYTES[0].a/n389 ), .Z(n1112)
         );
  XNOR U1113 ( .A(\SUBBYTES[0].a/n1500 ), .B(\SUBBYTES[0].a/n746 ), .Z(n1113)
         );
  XNOR U1114 ( .A(\SUBBYTES[0].a/n671 ), .B(\SUBBYTES[0].a/n670 ), .Z(n1114)
         );
  XNOR U1115 ( .A(\SUBBYTES[0].a/n695 ), .B(\SUBBYTES[0].a/n694 ), .Z(n1115)
         );
  XNOR U1116 ( .A(\SUBBYTES[0].a/n668 ), .B(\SUBBYTES[0].a/n667 ), .Z(n1116)
         );
  XNOR U1117 ( .A(\SUBBYTES[0].a/n692 ), .B(\SUBBYTES[0].a/n691 ), .Z(n1117)
         );
  XNOR U1118 ( .A(\SUBBYTES[0].a/n662 ), .B(\SUBBYTES[0].a/n661 ), .Z(n1118)
         );
  XNOR U1119 ( .A(\SUBBYTES[0].a/n686 ), .B(\SUBBYTES[0].a/n685 ), .Z(n1119)
         );
  XNOR U1120 ( .A(\SUBBYTES[0].a/n1480 ), .B(\SUBBYTES[0].a/n660 ), .Z(n1120)
         );
  XNOR U1121 ( .A(\SUBBYTES[0].a/n1485 ), .B(\SUBBYTES[0].a/n684 ), .Z(n1121)
         );
  XNOR U1122 ( .A(\SUBBYTES[0].a/n1482 ), .B(\SUBBYTES[0].a/n659 ), .Z(n1122)
         );
  XNOR U1123 ( .A(\SUBBYTES[0].a/n1487 ), .B(\SUBBYTES[0].a/n683 ), .Z(n1123)
         );
  XNOR U1124 ( .A(\SUBBYTES[0].a/n1483 ), .B(\SUBBYTES[0].a/n653 ), .Z(n1124)
         );
  XNOR U1125 ( .A(\SUBBYTES[0].a/n1488 ), .B(\SUBBYTES[0].a/n677 ), .Z(n1125)
         );
  XNOR U1126 ( .A(\SUBBYTES[0].a/n1480 ), .B(\SUBBYTES[0].a/n650 ), .Z(n1126)
         );
  XNOR U1127 ( .A(\SUBBYTES[0].a/n575 ), .B(\SUBBYTES[0].a/n574 ), .Z(n1127)
         );
  XNOR U1128 ( .A(\SUBBYTES[0].a/n599 ), .B(\SUBBYTES[0].a/n598 ), .Z(n1128)
         );
  XNOR U1129 ( .A(\SUBBYTES[0].a/n572 ), .B(\SUBBYTES[0].a/n571 ), .Z(n1129)
         );
  XNOR U1130 ( .A(\SUBBYTES[0].a/n596 ), .B(\SUBBYTES[0].a/n595 ), .Z(n1130)
         );
  XNOR U1131 ( .A(\SUBBYTES[0].a/n566 ), .B(\SUBBYTES[0].a/n565 ), .Z(n1131)
         );
  XNOR U1132 ( .A(\SUBBYTES[0].a/n590 ), .B(\SUBBYTES[0].a/n589 ), .Z(n1132)
         );
  XNOR U1133 ( .A(\SUBBYTES[0].a/n1460 ), .B(\SUBBYTES[0].a/n564 ), .Z(n1133)
         );
  XNOR U1134 ( .A(\SUBBYTES[0].a/n1465 ), .B(\SUBBYTES[0].a/n588 ), .Z(n1134)
         );
  XNOR U1135 ( .A(\SUBBYTES[0].a/n1462 ), .B(\SUBBYTES[0].a/n563 ), .Z(n1135)
         );
  XNOR U1136 ( .A(\SUBBYTES[0].a/n1467 ), .B(\SUBBYTES[0].a/n587 ), .Z(n1136)
         );
  XNOR U1137 ( .A(\SUBBYTES[0].a/n1463 ), .B(\SUBBYTES[0].a/n557 ), .Z(n1137)
         );
  XNOR U1138 ( .A(\SUBBYTES[0].a/n1468 ), .B(\SUBBYTES[0].a/n581 ), .Z(n1138)
         );
  XNOR U1139 ( .A(\SUBBYTES[0].a/n1460 ), .B(\SUBBYTES[0].a/n554 ), .Z(n1139)
         );
  XNOR U1140 ( .A(\SUBBYTES[0].a/n479 ), .B(\SUBBYTES[0].a/n478 ), .Z(n1140)
         );
  XNOR U1141 ( .A(\SUBBYTES[0].a/n503 ), .B(\SUBBYTES[0].a/n502 ), .Z(n1141)
         );
  XNOR U1142 ( .A(\SUBBYTES[0].a/n476 ), .B(\SUBBYTES[0].a/n475 ), .Z(n1142)
         );
  XNOR U1143 ( .A(\SUBBYTES[0].a/n500 ), .B(\SUBBYTES[0].a/n499 ), .Z(n1143)
         );
  XNOR U1144 ( .A(\SUBBYTES[0].a/n470 ), .B(\SUBBYTES[0].a/n469 ), .Z(n1144)
         );
  XNOR U1145 ( .A(\SUBBYTES[0].a/n494 ), .B(\SUBBYTES[0].a/n493 ), .Z(n1145)
         );
  XNOR U1146 ( .A(\SUBBYTES[0].a/n1440 ), .B(\SUBBYTES[0].a/n468 ), .Z(n1146)
         );
  XNOR U1147 ( .A(\SUBBYTES[0].a/n1445 ), .B(\SUBBYTES[0].a/n492 ), .Z(n1147)
         );
  XNOR U1148 ( .A(\SUBBYTES[0].a/n1442 ), .B(\SUBBYTES[0].a/n467 ), .Z(n1148)
         );
  XNOR U1149 ( .A(\SUBBYTES[0].a/n1447 ), .B(\SUBBYTES[0].a/n491 ), .Z(n1149)
         );
  XNOR U1150 ( .A(\SUBBYTES[0].a/n1443 ), .B(\SUBBYTES[0].a/n461 ), .Z(n1150)
         );
  XNOR U1151 ( .A(\SUBBYTES[0].a/n1448 ), .B(\SUBBYTES[0].a/n485 ), .Z(n1151)
         );
  XNOR U1152 ( .A(\SUBBYTES[0].a/n1440 ), .B(\SUBBYTES[0].a/n458 ), .Z(n1152)
         );
  AND U1153 ( .A(\SUBBYTES[0].a/w209 ), .B(\SUBBYTES[0].a/w222 ), .Z(n1153) );
  AND U1154 ( .A(\SUBBYTES[0].a/w416 ), .B(\SUBBYTES[0].a/w429 ), .Z(n1154) );
  AND U1155 ( .A(\SUBBYTES[0].a/w623 ), .B(\SUBBYTES[0].a/w636 ), .Z(n1155) );
  AND U1156 ( .A(\SUBBYTES[0].a/w830 ), .B(\SUBBYTES[0].a/w843 ), .Z(n1156) );
  AND U1157 ( .A(\SUBBYTES[0].a/w1037 ), .B(\SUBBYTES[0].a/w1050 ), .Z(n1157)
         );
  AND U1158 ( .A(\SUBBYTES[0].a/w1244 ), .B(\SUBBYTES[0].a/w1257 ), .Z(n1158)
         );
  AND U1159 ( .A(\SUBBYTES[0].a/w1451 ), .B(\SUBBYTES[0].a/w1464 ), .Z(n1159)
         );
  AND U1160 ( .A(\SUBBYTES[0].a/w1658 ), .B(\SUBBYTES[0].a/w1671 ), .Z(n1160)
         );
  AND U1161 ( .A(\SUBBYTES[0].a/w1865 ), .B(\SUBBYTES[0].a/w1878 ), .Z(n1161)
         );
  AND U1162 ( .A(\SUBBYTES[0].a/w2072 ), .B(\SUBBYTES[0].a/w2085 ), .Z(n1162)
         );
  AND U1163 ( .A(\SUBBYTES[0].a/w2279 ), .B(\SUBBYTES[0].a/w2292 ), .Z(n1163)
         );
  AND U1164 ( .A(\SUBBYTES[0].a/w2486 ), .B(\SUBBYTES[0].a/w2499 ), .Z(n1164)
         );
  AND U1165 ( .A(\SUBBYTES[0].a/w2693 ), .B(\SUBBYTES[0].a/w2706 ), .Z(n1165)
         );
  AND U1166 ( .A(\SUBBYTES[0].a/w2900 ), .B(\SUBBYTES[0].a/w2913 ), .Z(n1166)
         );
  AND U1167 ( .A(\SUBBYTES[0].a/w3107 ), .B(\SUBBYTES[0].a/w3120 ), .Z(n1167)
         );
  AND U1168 ( .A(\SUBBYTES[0].a/w3314 ), .B(\SUBBYTES[0].a/w3327 ), .Z(n1168)
         );
  IV U1169 ( .A(n16056), .Z(\w3[8][98] ) );
  IV U1170 ( .A(n16067), .Z(\w3[8][90] ) );
  IV U1171 ( .A(n16062), .Z(\w3[8][82] ) );
  IV U1172 ( .A(n16057), .Z(\w3[8][74] ) );
  IV U1173 ( .A(n16068), .Z(\w3[8][66] ) );
  IV U1174 ( .A(n16063), .Z(\w3[8][58] ) );
  IV U1175 ( .A(n16058), .Z(\w3[8][50] ) );
  IV U1176 ( .A(n16069), .Z(\w3[8][42] ) );
  IV U1177 ( .A(n16064), .Z(\w3[8][34] ) );
  IV U1178 ( .A(n16060), .Z(\w3[8][2] ) );
  IV U1179 ( .A(n16059), .Z(\w3[8][26] ) );
  IV U1180 ( .A(n16070), .Z(\w3[8][18] ) );
  IV U1181 ( .A(n16071), .Z(\w3[8][122] ) );
  IV U1182 ( .A(n16066), .Z(\w3[8][114] ) );
  IV U1183 ( .A(n16065), .Z(\w3[8][10] ) );
  IV U1184 ( .A(n16061), .Z(\w3[8][106] ) );
  IV U1185 ( .A(n14776), .Z(\w3[7][98] ) );
  IV U1186 ( .A(n14787), .Z(\w3[7][90] ) );
  IV U1187 ( .A(n14782), .Z(\w3[7][82] ) );
  IV U1188 ( .A(n14777), .Z(\w3[7][74] ) );
  IV U1189 ( .A(n14788), .Z(\w3[7][66] ) );
  IV U1190 ( .A(n14783), .Z(\w3[7][58] ) );
  IV U1191 ( .A(n14778), .Z(\w3[7][50] ) );
  IV U1192 ( .A(n14789), .Z(\w3[7][42] ) );
  IV U1193 ( .A(n14784), .Z(\w3[7][34] ) );
  IV U1194 ( .A(n14780), .Z(\w3[7][2] ) );
  IV U1195 ( .A(n14779), .Z(\w3[7][26] ) );
  IV U1196 ( .A(n14790), .Z(\w3[7][18] ) );
  IV U1197 ( .A(n14791), .Z(\w3[7][122] ) );
  IV U1198 ( .A(n14786), .Z(\w3[7][114] ) );
  IV U1199 ( .A(n14785), .Z(\w3[7][10] ) );
  IV U1200 ( .A(n14781), .Z(\w3[7][106] ) );
  IV U1201 ( .A(n13496), .Z(\w3[6][98] ) );
  IV U1202 ( .A(n13507), .Z(\w3[6][90] ) );
  IV U1203 ( .A(n13502), .Z(\w3[6][82] ) );
  IV U1204 ( .A(n13497), .Z(\w3[6][74] ) );
  IV U1205 ( .A(n13508), .Z(\w3[6][66] ) );
  IV U1206 ( .A(n13503), .Z(\w3[6][58] ) );
  IV U1207 ( .A(n13498), .Z(\w3[6][50] ) );
  IV U1208 ( .A(n13509), .Z(\w3[6][42] ) );
  IV U1209 ( .A(n13504), .Z(\w3[6][34] ) );
  IV U1210 ( .A(n13500), .Z(\w3[6][2] ) );
  IV U1211 ( .A(n13499), .Z(\w3[6][26] ) );
  IV U1212 ( .A(n13510), .Z(\w3[6][18] ) );
  IV U1213 ( .A(n13511), .Z(\w3[6][122] ) );
  IV U1214 ( .A(n13506), .Z(\w3[6][114] ) );
  IV U1215 ( .A(n13505), .Z(\w3[6][10] ) );
  IV U1216 ( .A(n13501), .Z(\w3[6][106] ) );
  IV U1217 ( .A(n12216), .Z(\w3[5][98] ) );
  IV U1218 ( .A(n12227), .Z(\w3[5][90] ) );
  IV U1219 ( .A(n12222), .Z(\w3[5][82] ) );
  IV U1220 ( .A(n12217), .Z(\w3[5][74] ) );
  IV U1221 ( .A(n12228), .Z(\w3[5][66] ) );
  IV U1222 ( .A(n12223), .Z(\w3[5][58] ) );
  IV U1223 ( .A(n12218), .Z(\w3[5][50] ) );
  IV U1224 ( .A(n12229), .Z(\w3[5][42] ) );
  IV U1225 ( .A(n12224), .Z(\w3[5][34] ) );
  IV U1226 ( .A(n12220), .Z(\w3[5][2] ) );
  IV U1227 ( .A(n12219), .Z(\w3[5][26] ) );
  IV U1228 ( .A(n12230), .Z(\w3[5][18] ) );
  IV U1229 ( .A(n12231), .Z(\w3[5][122] ) );
  IV U1230 ( .A(n12226), .Z(\w3[5][114] ) );
  IV U1231 ( .A(n12225), .Z(\w3[5][10] ) );
  IV U1232 ( .A(n12221), .Z(\w3[5][106] ) );
  IV U1233 ( .A(n10936), .Z(\w3[4][98] ) );
  IV U1234 ( .A(n10947), .Z(\w3[4][90] ) );
  IV U1235 ( .A(n10942), .Z(\w3[4][82] ) );
  IV U1236 ( .A(n10937), .Z(\w3[4][74] ) );
  IV U1237 ( .A(n10948), .Z(\w3[4][66] ) );
  IV U1238 ( .A(n10943), .Z(\w3[4][58] ) );
  IV U1239 ( .A(n10938), .Z(\w3[4][50] ) );
  IV U1240 ( .A(n10949), .Z(\w3[4][42] ) );
  IV U1241 ( .A(n10944), .Z(\w3[4][34] ) );
  IV U1242 ( .A(n10940), .Z(\w3[4][2] ) );
  IV U1243 ( .A(n10939), .Z(\w3[4][26] ) );
  IV U1244 ( .A(n10950), .Z(\w3[4][18] ) );
  IV U1245 ( .A(n10951), .Z(\w3[4][122] ) );
  IV U1246 ( .A(n10946), .Z(\w3[4][114] ) );
  IV U1247 ( .A(n10945), .Z(\w3[4][10] ) );
  IV U1248 ( .A(n10941), .Z(\w3[4][106] ) );
  IV U1249 ( .A(n9656), .Z(\w3[3][98] ) );
  IV U1250 ( .A(n9667), .Z(\w3[3][90] ) );
  IV U1251 ( .A(n9662), .Z(\w3[3][82] ) );
  IV U1252 ( .A(n9657), .Z(\w3[3][74] ) );
  IV U1253 ( .A(n9668), .Z(\w3[3][66] ) );
  IV U1254 ( .A(n9663), .Z(\w3[3][58] ) );
  IV U1255 ( .A(n9658), .Z(\w3[3][50] ) );
  IV U1256 ( .A(n9669), .Z(\w3[3][42] ) );
  IV U1257 ( .A(n9664), .Z(\w3[3][34] ) );
  IV U1258 ( .A(n9660), .Z(\w3[3][2] ) );
  IV U1259 ( .A(n9659), .Z(\w3[3][26] ) );
  IV U1260 ( .A(n9670), .Z(\w3[3][18] ) );
  IV U1261 ( .A(n9671), .Z(\w3[3][122] ) );
  IV U1262 ( .A(n9666), .Z(\w3[3][114] ) );
  IV U1263 ( .A(n9665), .Z(\w3[3][10] ) );
  IV U1264 ( .A(n9661), .Z(\w3[3][106] ) );
  IV U1265 ( .A(n8376), .Z(\w3[2][98] ) );
  IV U1266 ( .A(n8387), .Z(\w3[2][90] ) );
  IV U1267 ( .A(n8382), .Z(\w3[2][82] ) );
  IV U1268 ( .A(n8377), .Z(\w3[2][74] ) );
  IV U1269 ( .A(n8388), .Z(\w3[2][66] ) );
  IV U1270 ( .A(n8383), .Z(\w3[2][58] ) );
  IV U1271 ( .A(n8378), .Z(\w3[2][50] ) );
  IV U1272 ( .A(n8389), .Z(\w3[2][42] ) );
  IV U1273 ( .A(n8384), .Z(\w3[2][34] ) );
  IV U1274 ( .A(n8380), .Z(\w3[2][2] ) );
  IV U1275 ( .A(n8379), .Z(\w3[2][26] ) );
  IV U1276 ( .A(n8390), .Z(\w3[2][18] ) );
  IV U1277 ( .A(n8391), .Z(\w3[2][122] ) );
  IV U1278 ( .A(n8386), .Z(\w3[2][114] ) );
  IV U1279 ( .A(n8385), .Z(\w3[2][10] ) );
  IV U1280 ( .A(n8381), .Z(\w3[2][106] ) );
  IV U1281 ( .A(n7096), .Z(\w3[1][98] ) );
  IV U1282 ( .A(n7107), .Z(\w3[1][90] ) );
  IV U1283 ( .A(n7102), .Z(\w3[1][82] ) );
  IV U1284 ( .A(n7097), .Z(\w3[1][74] ) );
  IV U1285 ( .A(n7108), .Z(\w3[1][66] ) );
  IV U1286 ( .A(n7103), .Z(\w3[1][58] ) );
  IV U1287 ( .A(n7098), .Z(\w3[1][50] ) );
  IV U1288 ( .A(n7109), .Z(\w3[1][42] ) );
  IV U1289 ( .A(n7104), .Z(\w3[1][34] ) );
  IV U1290 ( .A(n7100), .Z(\w3[1][2] ) );
  IV U1291 ( .A(n7099), .Z(\w3[1][26] ) );
  IV U1292 ( .A(n7110), .Z(\w3[1][18] ) );
  IV U1293 ( .A(n7111), .Z(\w3[1][122] ) );
  IV U1294 ( .A(n7106), .Z(\w3[1][114] ) );
  IV U1295 ( .A(n7105), .Z(\w3[1][10] ) );
  IV U1296 ( .A(n7101), .Z(\w3[1][106] ) );
  IV U1297 ( .A(\SUBBYTES[0].a/n1619 ), .Z(\w3[0][98] ) );
  IV U1298 ( .A(\SUBBYTES[0].a/n1707 ), .Z(\w3[0][90] ) );
  IV U1299 ( .A(\SUBBYTES[0].a/n1667 ), .Z(\w3[0][82] ) );
  IV U1300 ( .A(\SUBBYTES[0].a/n1627 ), .Z(\w3[0][74] ) );
  IV U1301 ( .A(\SUBBYTES[0].a/n1715 ), .Z(\w3[0][66] ) );
  IV U1302 ( .A(\SUBBYTES[0].a/n1675 ), .Z(\w3[0][58] ) );
  IV U1303 ( .A(\SUBBYTES[0].a/n1635 ), .Z(\w3[0][50] ) );
  IV U1304 ( .A(\SUBBYTES[0].a/n1723 ), .Z(\w3[0][42] ) );
  IV U1305 ( .A(\SUBBYTES[0].a/n1683 ), .Z(\w3[0][34] ) );
  IV U1306 ( .A(\SUBBYTES[0].a/n1651 ), .Z(\w3[0][2] ) );
  IV U1307 ( .A(\SUBBYTES[0].a/n1643 ), .Z(\w3[0][26] ) );
  IV U1308 ( .A(\SUBBYTES[0].a/n1731 ), .Z(\w3[0][18] ) );
  IV U1309 ( .A(\SUBBYTES[0].a/n1739 ), .Z(\w3[0][122] ) );
  IV U1310 ( .A(\SUBBYTES[0].a/n1699 ), .Z(\w3[0][114] ) );
  IV U1311 ( .A(\SUBBYTES[0].a/n1691 ), .Z(\w3[0][10] ) );
  IV U1312 ( .A(\SUBBYTES[0].a/n1659 ), .Z(\w3[0][106] ) );
  XOR U1313 ( .A(\w0[9][99] ), .B(g_input[1251]), .Z(\w1[9][99] ) );
  XOR U1314 ( .A(\w0[9][94] ), .B(g_input[1246]), .Z(\w1[9][94] ) );
  XOR U1315 ( .A(\w0[9][93] ), .B(g_input[1245]), .Z(\w1[9][93] ) );
  XOR U1316 ( .A(\w0[9][91] ), .B(g_input[1243]), .Z(\w1[9][91] ) );
  XOR U1317 ( .A(\w0[9][86] ), .B(g_input[1238]), .Z(\w1[9][86] ) );
  XOR U1318 ( .A(\w0[9][85] ), .B(g_input[1237]), .Z(\w1[9][85] ) );
  XOR U1319 ( .A(\w0[9][83] ), .B(g_input[1235]), .Z(\w1[9][83] ) );
  XOR U1320 ( .A(\w0[9][78] ), .B(g_input[1230]), .Z(\w1[9][78] ) );
  XOR U1321 ( .A(\w0[9][77] ), .B(g_input[1229]), .Z(\w1[9][77] ) );
  XOR U1322 ( .A(\w0[9][75] ), .B(g_input[1227]), .Z(\w1[9][75] ) );
  XOR U1323 ( .A(\w0[9][70] ), .B(g_input[1222]), .Z(\w1[9][70] ) );
  XOR U1324 ( .A(\w0[9][6] ), .B(g_input[1158]), .Z(\w1[9][6] ) );
  XOR U1325 ( .A(\w0[9][69] ), .B(g_input[1221]), .Z(\w1[9][69] ) );
  XOR U1326 ( .A(\w0[9][67] ), .B(g_input[1219]), .Z(\w1[9][67] ) );
  XOR U1327 ( .A(\w0[9][62] ), .B(g_input[1214]), .Z(\w1[9][62] ) );
  XOR U1328 ( .A(\w0[9][61] ), .B(g_input[1213]), .Z(\w1[9][61] ) );
  XOR U1329 ( .A(\w0[9][5] ), .B(g_input[1157]), .Z(\w1[9][5] ) );
  XOR U1330 ( .A(\w0[9][59] ), .B(g_input[1211]), .Z(\w1[9][59] ) );
  XOR U1331 ( .A(\w0[9][54] ), .B(g_input[1206]), .Z(\w1[9][54] ) );
  XOR U1332 ( .A(\w0[9][53] ), .B(g_input[1205]), .Z(\w1[9][53] ) );
  XOR U1333 ( .A(\w0[9][51] ), .B(g_input[1203]), .Z(\w1[9][51] ) );
  XOR U1334 ( .A(\w0[9][46] ), .B(g_input[1198]), .Z(\w1[9][46] ) );
  XOR U1335 ( .A(\w0[9][45] ), .B(g_input[1197]), .Z(\w1[9][45] ) );
  XOR U1336 ( .A(\w0[9][43] ), .B(g_input[1195]), .Z(\w1[9][43] ) );
  XOR U1337 ( .A(\w0[9][3] ), .B(g_input[1155]), .Z(\w1[9][3] ) );
  XOR U1338 ( .A(\w0[9][38] ), .B(g_input[1190]), .Z(\w1[9][38] ) );
  XOR U1339 ( .A(\w0[9][37] ), .B(g_input[1189]), .Z(\w1[9][37] ) );
  XOR U1340 ( .A(\w0[9][35] ), .B(g_input[1187]), .Z(\w1[9][35] ) );
  XOR U1341 ( .A(\w0[9][30] ), .B(g_input[1182]), .Z(\w1[9][30] ) );
  XOR U1342 ( .A(\w0[9][29] ), .B(g_input[1181]), .Z(\w1[9][29] ) );
  XOR U1343 ( .A(\w0[9][27] ), .B(g_input[1179]), .Z(\w1[9][27] ) );
  XOR U1344 ( .A(\w0[9][22] ), .B(g_input[1174]), .Z(\w1[9][22] ) );
  XOR U1345 ( .A(\w0[9][21] ), .B(g_input[1173]), .Z(\w1[9][21] ) );
  XOR U1346 ( .A(\w0[9][19] ), .B(g_input[1171]), .Z(\w1[9][19] ) );
  XOR U1347 ( .A(\w0[9][14] ), .B(g_input[1166]), .Z(\w1[9][14] ) );
  XOR U1348 ( .A(\w0[9][13] ), .B(g_input[1165]), .Z(\w1[9][13] ) );
  XOR U1349 ( .A(\w0[9][126] ), .B(g_input[1278]), .Z(\w1[9][126] ) );
  XOR U1350 ( .A(\w0[9][125] ), .B(g_input[1277]), .Z(\w1[9][125] ) );
  XOR U1351 ( .A(\w0[9][123] ), .B(g_input[1275]), .Z(\w1[9][123] ) );
  XOR U1352 ( .A(\w0[9][11] ), .B(g_input[1163]), .Z(\w1[9][11] ) );
  XOR U1353 ( .A(\w0[9][118] ), .B(g_input[1270]), .Z(\w1[9][118] ) );
  XOR U1354 ( .A(\w0[9][117] ), .B(g_input[1269]), .Z(\w1[9][117] ) );
  XOR U1355 ( .A(\w0[9][115] ), .B(g_input[1267]), .Z(\w1[9][115] ) );
  XOR U1356 ( .A(\w0[9][110] ), .B(g_input[1262]), .Z(\w1[9][110] ) );
  XOR U1357 ( .A(\w0[9][109] ), .B(g_input[1261]), .Z(\w1[9][109] ) );
  XOR U1358 ( .A(\w0[9][107] ), .B(g_input[1259]), .Z(\w1[9][107] ) );
  XOR U1359 ( .A(\w0[9][102] ), .B(g_input[1254]), .Z(\w1[9][102] ) );
  XOR U1360 ( .A(\w0[9][101] ), .B(g_input[1253]), .Z(\w1[9][101] ) );
  XOR U1361 ( .A(\w0[8][99] ), .B(g_input[1123]), .Z(\w1[8][99] ) );
  XOR U1362 ( .A(\w0[8][94] ), .B(g_input[1118]), .Z(\w1[8][94] ) );
  XOR U1363 ( .A(\w0[8][93] ), .B(g_input[1117]), .Z(\w1[8][93] ) );
  XOR U1364 ( .A(\w0[8][91] ), .B(g_input[1115]), .Z(\w1[8][91] ) );
  XOR U1365 ( .A(\w0[8][86] ), .B(g_input[1110]), .Z(\w1[8][86] ) );
  XOR U1366 ( .A(\w0[8][85] ), .B(g_input[1109]), .Z(\w1[8][85] ) );
  XOR U1367 ( .A(\w0[8][83] ), .B(g_input[1107]), .Z(\w1[8][83] ) );
  XOR U1368 ( .A(\w0[8][78] ), .B(g_input[1102]), .Z(\w1[8][78] ) );
  XOR U1369 ( .A(\w0[8][77] ), .B(g_input[1101]), .Z(\w1[8][77] ) );
  XOR U1370 ( .A(\w0[8][75] ), .B(g_input[1099]), .Z(\w1[8][75] ) );
  XOR U1371 ( .A(\w0[8][70] ), .B(g_input[1094]), .Z(\w1[8][70] ) );
  XOR U1372 ( .A(\w0[8][6] ), .B(g_input[1030]), .Z(\w1[8][6] ) );
  XOR U1373 ( .A(\w0[8][69] ), .B(g_input[1093]), .Z(\w1[8][69] ) );
  XOR U1374 ( .A(\w0[8][67] ), .B(g_input[1091]), .Z(\w1[8][67] ) );
  XOR U1375 ( .A(\w0[8][62] ), .B(g_input[1086]), .Z(\w1[8][62] ) );
  XOR U1376 ( .A(\w0[8][61] ), .B(g_input[1085]), .Z(\w1[8][61] ) );
  XOR U1377 ( .A(\w0[8][5] ), .B(g_input[1029]), .Z(\w1[8][5] ) );
  XOR U1378 ( .A(\w0[8][59] ), .B(g_input[1083]), .Z(\w1[8][59] ) );
  XOR U1379 ( .A(\w0[8][54] ), .B(g_input[1078]), .Z(\w1[8][54] ) );
  XOR U1380 ( .A(\w0[8][53] ), .B(g_input[1077]), .Z(\w1[8][53] ) );
  XOR U1381 ( .A(\w0[8][51] ), .B(g_input[1075]), .Z(\w1[8][51] ) );
  XOR U1382 ( .A(\w0[8][46] ), .B(g_input[1070]), .Z(\w1[8][46] ) );
  XOR U1383 ( .A(\w0[8][45] ), .B(g_input[1069]), .Z(\w1[8][45] ) );
  XOR U1384 ( .A(\w0[8][43] ), .B(g_input[1067]), .Z(\w1[8][43] ) );
  XOR U1385 ( .A(\w0[8][3] ), .B(g_input[1027]), .Z(\w1[8][3] ) );
  XOR U1386 ( .A(\w0[8][38] ), .B(g_input[1062]), .Z(\w1[8][38] ) );
  XOR U1387 ( .A(\w0[8][37] ), .B(g_input[1061]), .Z(\w1[8][37] ) );
  XOR U1388 ( .A(\w0[8][35] ), .B(g_input[1059]), .Z(\w1[8][35] ) );
  XOR U1389 ( .A(\w0[8][30] ), .B(g_input[1054]), .Z(\w1[8][30] ) );
  XOR U1390 ( .A(\w0[8][29] ), .B(g_input[1053]), .Z(\w1[8][29] ) );
  XOR U1391 ( .A(\w0[8][27] ), .B(g_input[1051]), .Z(\w1[8][27] ) );
  XOR U1392 ( .A(\w0[8][22] ), .B(g_input[1046]), .Z(\w1[8][22] ) );
  XOR U1393 ( .A(\w0[8][21] ), .B(g_input[1045]), .Z(\w1[8][21] ) );
  XOR U1394 ( .A(\w0[8][19] ), .B(g_input[1043]), .Z(\w1[8][19] ) );
  XOR U1395 ( .A(\w0[8][14] ), .B(g_input[1038]), .Z(\w1[8][14] ) );
  XOR U1396 ( .A(\w0[8][13] ), .B(g_input[1037]), .Z(\w1[8][13] ) );
  XOR U1397 ( .A(\w0[8][126] ), .B(g_input[1150]), .Z(\w1[8][126] ) );
  XOR U1398 ( .A(\w0[8][125] ), .B(g_input[1149]), .Z(\w1[8][125] ) );
  XOR U1399 ( .A(\w0[8][123] ), .B(g_input[1147]), .Z(\w1[8][123] ) );
  XOR U1400 ( .A(\w0[8][11] ), .B(g_input[1035]), .Z(\w1[8][11] ) );
  XOR U1401 ( .A(\w0[8][118] ), .B(g_input[1142]), .Z(\w1[8][118] ) );
  XOR U1402 ( .A(\w0[8][117] ), .B(g_input[1141]), .Z(\w1[8][117] ) );
  XOR U1403 ( .A(\w0[8][115] ), .B(g_input[1139]), .Z(\w1[8][115] ) );
  XOR U1404 ( .A(\w0[8][110] ), .B(g_input[1134]), .Z(\w1[8][110] ) );
  XOR U1405 ( .A(\w0[8][109] ), .B(g_input[1133]), .Z(\w1[8][109] ) );
  XOR U1406 ( .A(\w0[8][107] ), .B(g_input[1131]), .Z(\w1[8][107] ) );
  XOR U1407 ( .A(\w0[8][102] ), .B(g_input[1126]), .Z(\w1[8][102] ) );
  XOR U1408 ( .A(\w0[8][101] ), .B(g_input[1125]), .Z(\w1[8][101] ) );
  XOR U1409 ( .A(\w0[7][99] ), .B(g_input[995]), .Z(\w1[7][99] ) );
  XOR U1410 ( .A(\w0[7][94] ), .B(g_input[990]), .Z(\w1[7][94] ) );
  XOR U1411 ( .A(\w0[7][93] ), .B(g_input[989]), .Z(\w1[7][93] ) );
  XOR U1412 ( .A(\w0[7][91] ), .B(g_input[987]), .Z(\w1[7][91] ) );
  XOR U1413 ( .A(\w0[7][86] ), .B(g_input[982]), .Z(\w1[7][86] ) );
  XOR U1414 ( .A(\w0[7][85] ), .B(g_input[981]), .Z(\w1[7][85] ) );
  XOR U1415 ( .A(\w0[7][83] ), .B(g_input[979]), .Z(\w1[7][83] ) );
  XOR U1416 ( .A(\w0[7][78] ), .B(g_input[974]), .Z(\w1[7][78] ) );
  XOR U1417 ( .A(\w0[7][77] ), .B(g_input[973]), .Z(\w1[7][77] ) );
  XOR U1418 ( .A(\w0[7][75] ), .B(g_input[971]), .Z(\w1[7][75] ) );
  XOR U1419 ( .A(\w0[7][70] ), .B(g_input[966]), .Z(\w1[7][70] ) );
  XOR U1420 ( .A(\w0[7][6] ), .B(g_input[902]), .Z(\w1[7][6] ) );
  XOR U1421 ( .A(\w0[7][69] ), .B(g_input[965]), .Z(\w1[7][69] ) );
  XOR U1422 ( .A(\w0[7][67] ), .B(g_input[963]), .Z(\w1[7][67] ) );
  XOR U1423 ( .A(\w0[7][62] ), .B(g_input[958]), .Z(\w1[7][62] ) );
  XOR U1424 ( .A(\w0[7][61] ), .B(g_input[957]), .Z(\w1[7][61] ) );
  XOR U1425 ( .A(\w0[7][5] ), .B(g_input[901]), .Z(\w1[7][5] ) );
  XOR U1426 ( .A(\w0[7][59] ), .B(g_input[955]), .Z(\w1[7][59] ) );
  XOR U1427 ( .A(\w0[7][54] ), .B(g_input[950]), .Z(\w1[7][54] ) );
  XOR U1428 ( .A(\w0[7][53] ), .B(g_input[949]), .Z(\w1[7][53] ) );
  XOR U1429 ( .A(\w0[7][51] ), .B(g_input[947]), .Z(\w1[7][51] ) );
  XOR U1430 ( .A(\w0[7][46] ), .B(g_input[942]), .Z(\w1[7][46] ) );
  XOR U1431 ( .A(\w0[7][45] ), .B(g_input[941]), .Z(\w1[7][45] ) );
  XOR U1432 ( .A(\w0[7][43] ), .B(g_input[939]), .Z(\w1[7][43] ) );
  XOR U1433 ( .A(\w0[7][3] ), .B(g_input[899]), .Z(\w1[7][3] ) );
  XOR U1434 ( .A(\w0[7][38] ), .B(g_input[934]), .Z(\w1[7][38] ) );
  XOR U1435 ( .A(\w0[7][37] ), .B(g_input[933]), .Z(\w1[7][37] ) );
  XOR U1436 ( .A(\w0[7][35] ), .B(g_input[931]), .Z(\w1[7][35] ) );
  XOR U1437 ( .A(\w0[7][30] ), .B(g_input[926]), .Z(\w1[7][30] ) );
  XOR U1438 ( .A(\w0[7][29] ), .B(g_input[925]), .Z(\w1[7][29] ) );
  XOR U1439 ( .A(\w0[7][27] ), .B(g_input[923]), .Z(\w1[7][27] ) );
  XOR U1440 ( .A(\w0[7][22] ), .B(g_input[918]), .Z(\w1[7][22] ) );
  XOR U1441 ( .A(\w0[7][21] ), .B(g_input[917]), .Z(\w1[7][21] ) );
  XOR U1442 ( .A(\w0[7][19] ), .B(g_input[915]), .Z(\w1[7][19] ) );
  XOR U1443 ( .A(\w0[7][14] ), .B(g_input[910]), .Z(\w1[7][14] ) );
  XOR U1444 ( .A(\w0[7][13] ), .B(g_input[909]), .Z(\w1[7][13] ) );
  XOR U1445 ( .A(\w0[7][126] ), .B(g_input[1022]), .Z(\w1[7][126] ) );
  XOR U1446 ( .A(\w0[7][125] ), .B(g_input[1021]), .Z(\w1[7][125] ) );
  XOR U1447 ( .A(\w0[7][123] ), .B(g_input[1019]), .Z(\w1[7][123] ) );
  XOR U1448 ( .A(\w0[7][11] ), .B(g_input[907]), .Z(\w1[7][11] ) );
  XOR U1449 ( .A(\w0[7][118] ), .B(g_input[1014]), .Z(\w1[7][118] ) );
  XOR U1450 ( .A(\w0[7][117] ), .B(g_input[1013]), .Z(\w1[7][117] ) );
  XOR U1451 ( .A(\w0[7][115] ), .B(g_input[1011]), .Z(\w1[7][115] ) );
  XOR U1452 ( .A(\w0[7][110] ), .B(g_input[1006]), .Z(\w1[7][110] ) );
  XOR U1453 ( .A(\w0[7][109] ), .B(g_input[1005]), .Z(\w1[7][109] ) );
  XOR U1454 ( .A(\w0[7][107] ), .B(g_input[1003]), .Z(\w1[7][107] ) );
  XOR U1455 ( .A(\w0[7][102] ), .B(g_input[998]), .Z(\w1[7][102] ) );
  XOR U1456 ( .A(\w0[7][101] ), .B(g_input[997]), .Z(\w1[7][101] ) );
  XOR U1457 ( .A(\w0[6][99] ), .B(g_input[867]), .Z(\w1[6][99] ) );
  XOR U1458 ( .A(\w0[6][94] ), .B(g_input[862]), .Z(\w1[6][94] ) );
  XOR U1459 ( .A(\w0[6][93] ), .B(g_input[861]), .Z(\w1[6][93] ) );
  XOR U1460 ( .A(\w0[6][91] ), .B(g_input[859]), .Z(\w1[6][91] ) );
  XOR U1461 ( .A(\w0[6][86] ), .B(g_input[854]), .Z(\w1[6][86] ) );
  XOR U1462 ( .A(\w0[6][85] ), .B(g_input[853]), .Z(\w1[6][85] ) );
  XOR U1463 ( .A(\w0[6][83] ), .B(g_input[851]), .Z(\w1[6][83] ) );
  XOR U1464 ( .A(\w0[6][78] ), .B(g_input[846]), .Z(\w1[6][78] ) );
  XOR U1465 ( .A(\w0[6][77] ), .B(g_input[845]), .Z(\w1[6][77] ) );
  XOR U1466 ( .A(\w0[6][75] ), .B(g_input[843]), .Z(\w1[6][75] ) );
  XOR U1467 ( .A(\w0[6][70] ), .B(g_input[838]), .Z(\w1[6][70] ) );
  XOR U1468 ( .A(\w0[6][6] ), .B(g_input[774]), .Z(\w1[6][6] ) );
  XOR U1469 ( .A(\w0[6][69] ), .B(g_input[837]), .Z(\w1[6][69] ) );
  XOR U1470 ( .A(\w0[6][67] ), .B(g_input[835]), .Z(\w1[6][67] ) );
  XOR U1471 ( .A(\w0[6][62] ), .B(g_input[830]), .Z(\w1[6][62] ) );
  XOR U1472 ( .A(\w0[6][61] ), .B(g_input[829]), .Z(\w1[6][61] ) );
  XOR U1473 ( .A(\w0[6][5] ), .B(g_input[773]), .Z(\w1[6][5] ) );
  XOR U1474 ( .A(\w0[6][59] ), .B(g_input[827]), .Z(\w1[6][59] ) );
  XOR U1475 ( .A(\w0[6][54] ), .B(g_input[822]), .Z(\w1[6][54] ) );
  XOR U1476 ( .A(\w0[6][53] ), .B(g_input[821]), .Z(\w1[6][53] ) );
  XOR U1477 ( .A(\w0[6][51] ), .B(g_input[819]), .Z(\w1[6][51] ) );
  XOR U1478 ( .A(\w0[6][46] ), .B(g_input[814]), .Z(\w1[6][46] ) );
  XOR U1479 ( .A(\w0[6][45] ), .B(g_input[813]), .Z(\w1[6][45] ) );
  XOR U1480 ( .A(\w0[6][43] ), .B(g_input[811]), .Z(\w1[6][43] ) );
  XOR U1481 ( .A(\w0[6][3] ), .B(g_input[771]), .Z(\w1[6][3] ) );
  XOR U1482 ( .A(\w0[6][38] ), .B(g_input[806]), .Z(\w1[6][38] ) );
  XOR U1483 ( .A(\w0[6][37] ), .B(g_input[805]), .Z(\w1[6][37] ) );
  XOR U1484 ( .A(\w0[6][35] ), .B(g_input[803]), .Z(\w1[6][35] ) );
  XOR U1485 ( .A(\w0[6][30] ), .B(g_input[798]), .Z(\w1[6][30] ) );
  XOR U1486 ( .A(\w0[6][29] ), .B(g_input[797]), .Z(\w1[6][29] ) );
  XOR U1487 ( .A(\w0[6][27] ), .B(g_input[795]), .Z(\w1[6][27] ) );
  XOR U1488 ( .A(\w0[6][22] ), .B(g_input[790]), .Z(\w1[6][22] ) );
  XOR U1489 ( .A(\w0[6][21] ), .B(g_input[789]), .Z(\w1[6][21] ) );
  XOR U1490 ( .A(\w0[6][19] ), .B(g_input[787]), .Z(\w1[6][19] ) );
  XOR U1491 ( .A(\w0[6][14] ), .B(g_input[782]), .Z(\w1[6][14] ) );
  XOR U1492 ( .A(\w0[6][13] ), .B(g_input[781]), .Z(\w1[6][13] ) );
  XOR U1493 ( .A(\w0[6][126] ), .B(g_input[894]), .Z(\w1[6][126] ) );
  XOR U1494 ( .A(\w0[6][125] ), .B(g_input[893]), .Z(\w1[6][125] ) );
  XOR U1495 ( .A(\w0[6][123] ), .B(g_input[891]), .Z(\w1[6][123] ) );
  XOR U1496 ( .A(\w0[6][11] ), .B(g_input[779]), .Z(\w1[6][11] ) );
  XOR U1497 ( .A(\w0[6][118] ), .B(g_input[886]), .Z(\w1[6][118] ) );
  XOR U1498 ( .A(\w0[6][117] ), .B(g_input[885]), .Z(\w1[6][117] ) );
  XOR U1499 ( .A(\w0[6][115] ), .B(g_input[883]), .Z(\w1[6][115] ) );
  XOR U1500 ( .A(\w0[6][110] ), .B(g_input[878]), .Z(\w1[6][110] ) );
  XOR U1501 ( .A(\w0[6][109] ), .B(g_input[877]), .Z(\w1[6][109] ) );
  XOR U1502 ( .A(\w0[6][107] ), .B(g_input[875]), .Z(\w1[6][107] ) );
  XOR U1503 ( .A(\w0[6][102] ), .B(g_input[870]), .Z(\w1[6][102] ) );
  XOR U1504 ( .A(\w0[6][101] ), .B(g_input[869]), .Z(\w1[6][101] ) );
  XOR U1505 ( .A(\w0[5][99] ), .B(g_input[739]), .Z(\w1[5][99] ) );
  XOR U1506 ( .A(\w0[5][94] ), .B(g_input[734]), .Z(\w1[5][94] ) );
  XOR U1507 ( .A(\w0[5][93] ), .B(g_input[733]), .Z(\w1[5][93] ) );
  XOR U1508 ( .A(\w0[5][91] ), .B(g_input[731]), .Z(\w1[5][91] ) );
  XOR U1509 ( .A(\w0[5][86] ), .B(g_input[726]), .Z(\w1[5][86] ) );
  XOR U1510 ( .A(\w0[5][85] ), .B(g_input[725]), .Z(\w1[5][85] ) );
  XOR U1511 ( .A(\w0[5][83] ), .B(g_input[723]), .Z(\w1[5][83] ) );
  XOR U1512 ( .A(\w0[5][78] ), .B(g_input[718]), .Z(\w1[5][78] ) );
  XOR U1513 ( .A(\w0[5][77] ), .B(g_input[717]), .Z(\w1[5][77] ) );
  XOR U1514 ( .A(\w0[5][75] ), .B(g_input[715]), .Z(\w1[5][75] ) );
  XOR U1515 ( .A(\w0[5][70] ), .B(g_input[710]), .Z(\w1[5][70] ) );
  XOR U1516 ( .A(\w0[5][6] ), .B(g_input[646]), .Z(\w1[5][6] ) );
  XOR U1517 ( .A(\w0[5][69] ), .B(g_input[709]), .Z(\w1[5][69] ) );
  XOR U1518 ( .A(\w0[5][67] ), .B(g_input[707]), .Z(\w1[5][67] ) );
  XOR U1519 ( .A(\w0[5][62] ), .B(g_input[702]), .Z(\w1[5][62] ) );
  XOR U1520 ( .A(\w0[5][61] ), .B(g_input[701]), .Z(\w1[5][61] ) );
  XOR U1521 ( .A(\w0[5][5] ), .B(g_input[645]), .Z(\w1[5][5] ) );
  XOR U1522 ( .A(\w0[5][59] ), .B(g_input[699]), .Z(\w1[5][59] ) );
  XOR U1523 ( .A(\w0[5][54] ), .B(g_input[694]), .Z(\w1[5][54] ) );
  XOR U1524 ( .A(\w0[5][53] ), .B(g_input[693]), .Z(\w1[5][53] ) );
  XOR U1525 ( .A(\w0[5][51] ), .B(g_input[691]), .Z(\w1[5][51] ) );
  XOR U1526 ( .A(\w0[5][46] ), .B(g_input[686]), .Z(\w1[5][46] ) );
  XOR U1527 ( .A(\w0[5][45] ), .B(g_input[685]), .Z(\w1[5][45] ) );
  XOR U1528 ( .A(\w0[5][43] ), .B(g_input[683]), .Z(\w1[5][43] ) );
  XOR U1529 ( .A(\w0[5][3] ), .B(g_input[643]), .Z(\w1[5][3] ) );
  XOR U1530 ( .A(\w0[5][38] ), .B(g_input[678]), .Z(\w1[5][38] ) );
  XOR U1531 ( .A(\w0[5][37] ), .B(g_input[677]), .Z(\w1[5][37] ) );
  XOR U1532 ( .A(\w0[5][35] ), .B(g_input[675]), .Z(\w1[5][35] ) );
  XOR U1533 ( .A(\w0[5][30] ), .B(g_input[670]), .Z(\w1[5][30] ) );
  XOR U1534 ( .A(\w0[5][29] ), .B(g_input[669]), .Z(\w1[5][29] ) );
  XOR U1535 ( .A(\w0[5][27] ), .B(g_input[667]), .Z(\w1[5][27] ) );
  XOR U1536 ( .A(\w0[5][22] ), .B(g_input[662]), .Z(\w1[5][22] ) );
  XOR U1537 ( .A(\w0[5][21] ), .B(g_input[661]), .Z(\w1[5][21] ) );
  XOR U1538 ( .A(\w0[5][19] ), .B(g_input[659]), .Z(\w1[5][19] ) );
  XOR U1539 ( .A(\w0[5][14] ), .B(g_input[654]), .Z(\w1[5][14] ) );
  XOR U1540 ( .A(\w0[5][13] ), .B(g_input[653]), .Z(\w1[5][13] ) );
  XOR U1541 ( .A(\w0[5][126] ), .B(g_input[766]), .Z(\w1[5][126] ) );
  XOR U1542 ( .A(\w0[5][125] ), .B(g_input[765]), .Z(\w1[5][125] ) );
  XOR U1543 ( .A(\w0[5][123] ), .B(g_input[763]), .Z(\w1[5][123] ) );
  XOR U1544 ( .A(\w0[5][11] ), .B(g_input[651]), .Z(\w1[5][11] ) );
  XOR U1545 ( .A(\w0[5][118] ), .B(g_input[758]), .Z(\w1[5][118] ) );
  XOR U1546 ( .A(\w0[5][117] ), .B(g_input[757]), .Z(\w1[5][117] ) );
  XOR U1547 ( .A(\w0[5][115] ), .B(g_input[755]), .Z(\w1[5][115] ) );
  XOR U1548 ( .A(\w0[5][110] ), .B(g_input[750]), .Z(\w1[5][110] ) );
  XOR U1549 ( .A(\w0[5][109] ), .B(g_input[749]), .Z(\w1[5][109] ) );
  XOR U1550 ( .A(\w0[5][107] ), .B(g_input[747]), .Z(\w1[5][107] ) );
  XOR U1551 ( .A(\w0[5][102] ), .B(g_input[742]), .Z(\w1[5][102] ) );
  XOR U1552 ( .A(\w0[5][101] ), .B(g_input[741]), .Z(\w1[5][101] ) );
  XOR U1553 ( .A(\w0[4][99] ), .B(g_input[611]), .Z(\w1[4][99] ) );
  XOR U1554 ( .A(\w0[4][94] ), .B(g_input[606]), .Z(\w1[4][94] ) );
  XOR U1555 ( .A(\w0[4][93] ), .B(g_input[605]), .Z(\w1[4][93] ) );
  XOR U1556 ( .A(\w0[4][91] ), .B(g_input[603]), .Z(\w1[4][91] ) );
  XOR U1557 ( .A(\w0[4][86] ), .B(g_input[598]), .Z(\w1[4][86] ) );
  XOR U1558 ( .A(\w0[4][85] ), .B(g_input[597]), .Z(\w1[4][85] ) );
  XOR U1559 ( .A(\w0[4][83] ), .B(g_input[595]), .Z(\w1[4][83] ) );
  XOR U1560 ( .A(\w0[4][78] ), .B(g_input[590]), .Z(\w1[4][78] ) );
  XOR U1561 ( .A(\w0[4][77] ), .B(g_input[589]), .Z(\w1[4][77] ) );
  XOR U1562 ( .A(\w0[4][75] ), .B(g_input[587]), .Z(\w1[4][75] ) );
  XOR U1563 ( .A(\w0[4][70] ), .B(g_input[582]), .Z(\w1[4][70] ) );
  XOR U1564 ( .A(\w0[4][6] ), .B(g_input[518]), .Z(\w1[4][6] ) );
  XOR U1565 ( .A(\w0[4][69] ), .B(g_input[581]), .Z(\w1[4][69] ) );
  XOR U1566 ( .A(\w0[4][67] ), .B(g_input[579]), .Z(\w1[4][67] ) );
  XOR U1567 ( .A(\w0[4][62] ), .B(g_input[574]), .Z(\w1[4][62] ) );
  XOR U1568 ( .A(\w0[4][61] ), .B(g_input[573]), .Z(\w1[4][61] ) );
  XOR U1569 ( .A(\w0[4][5] ), .B(g_input[517]), .Z(\w1[4][5] ) );
  XOR U1570 ( .A(\w0[4][59] ), .B(g_input[571]), .Z(\w1[4][59] ) );
  XOR U1571 ( .A(\w0[4][54] ), .B(g_input[566]), .Z(\w1[4][54] ) );
  XOR U1572 ( .A(\w0[4][53] ), .B(g_input[565]), .Z(\w1[4][53] ) );
  XOR U1573 ( .A(\w0[4][51] ), .B(g_input[563]), .Z(\w1[4][51] ) );
  XOR U1574 ( .A(\w0[4][46] ), .B(g_input[558]), .Z(\w1[4][46] ) );
  XOR U1575 ( .A(\w0[4][45] ), .B(g_input[557]), .Z(\w1[4][45] ) );
  XOR U1576 ( .A(\w0[4][43] ), .B(g_input[555]), .Z(\w1[4][43] ) );
  XOR U1577 ( .A(\w0[4][3] ), .B(g_input[515]), .Z(\w1[4][3] ) );
  XOR U1578 ( .A(\w0[4][38] ), .B(g_input[550]), .Z(\w1[4][38] ) );
  XOR U1579 ( .A(\w0[4][37] ), .B(g_input[549]), .Z(\w1[4][37] ) );
  XOR U1580 ( .A(\w0[4][35] ), .B(g_input[547]), .Z(\w1[4][35] ) );
  XOR U1581 ( .A(\w0[4][30] ), .B(g_input[542]), .Z(\w1[4][30] ) );
  XOR U1582 ( .A(\w0[4][29] ), .B(g_input[541]), .Z(\w1[4][29] ) );
  XOR U1583 ( .A(\w0[4][27] ), .B(g_input[539]), .Z(\w1[4][27] ) );
  XOR U1584 ( .A(\w0[4][22] ), .B(g_input[534]), .Z(\w1[4][22] ) );
  XOR U1585 ( .A(\w0[4][21] ), .B(g_input[533]), .Z(\w1[4][21] ) );
  XOR U1586 ( .A(\w0[4][19] ), .B(g_input[531]), .Z(\w1[4][19] ) );
  XOR U1587 ( .A(\w0[4][14] ), .B(g_input[526]), .Z(\w1[4][14] ) );
  XOR U1588 ( .A(\w0[4][13] ), .B(g_input[525]), .Z(\w1[4][13] ) );
  XOR U1589 ( .A(\w0[4][126] ), .B(g_input[638]), .Z(\w1[4][126] ) );
  XOR U1590 ( .A(\w0[4][125] ), .B(g_input[637]), .Z(\w1[4][125] ) );
  XOR U1591 ( .A(\w0[4][123] ), .B(g_input[635]), .Z(\w1[4][123] ) );
  XOR U1592 ( .A(\w0[4][11] ), .B(g_input[523]), .Z(\w1[4][11] ) );
  XOR U1593 ( .A(\w0[4][118] ), .B(g_input[630]), .Z(\w1[4][118] ) );
  XOR U1594 ( .A(\w0[4][117] ), .B(g_input[629]), .Z(\w1[4][117] ) );
  XOR U1595 ( .A(\w0[4][115] ), .B(g_input[627]), .Z(\w1[4][115] ) );
  XOR U1596 ( .A(\w0[4][110] ), .B(g_input[622]), .Z(\w1[4][110] ) );
  XOR U1597 ( .A(\w0[4][109] ), .B(g_input[621]), .Z(\w1[4][109] ) );
  XOR U1598 ( .A(\w0[4][107] ), .B(g_input[619]), .Z(\w1[4][107] ) );
  XOR U1599 ( .A(\w0[4][102] ), .B(g_input[614]), .Z(\w1[4][102] ) );
  XOR U1600 ( .A(\w0[4][101] ), .B(g_input[613]), .Z(\w1[4][101] ) );
  XOR U1601 ( .A(\w0[3][99] ), .B(g_input[483]), .Z(\w1[3][99] ) );
  XOR U1602 ( .A(\w0[3][94] ), .B(g_input[478]), .Z(\w1[3][94] ) );
  XOR U1603 ( .A(\w0[3][93] ), .B(g_input[477]), .Z(\w1[3][93] ) );
  XOR U1604 ( .A(\w0[3][91] ), .B(g_input[475]), .Z(\w1[3][91] ) );
  XOR U1605 ( .A(\w0[3][86] ), .B(g_input[470]), .Z(\w1[3][86] ) );
  XOR U1606 ( .A(\w0[3][85] ), .B(g_input[469]), .Z(\w1[3][85] ) );
  XOR U1607 ( .A(\w0[3][83] ), .B(g_input[467]), .Z(\w1[3][83] ) );
  XOR U1608 ( .A(\w0[3][78] ), .B(g_input[462]), .Z(\w1[3][78] ) );
  XOR U1609 ( .A(\w0[3][77] ), .B(g_input[461]), .Z(\w1[3][77] ) );
  XOR U1610 ( .A(\w0[3][75] ), .B(g_input[459]), .Z(\w1[3][75] ) );
  XOR U1611 ( .A(\w0[3][70] ), .B(g_input[454]), .Z(\w1[3][70] ) );
  XOR U1612 ( .A(\w0[3][6] ), .B(g_input[390]), .Z(\w1[3][6] ) );
  XOR U1613 ( .A(\w0[3][69] ), .B(g_input[453]), .Z(\w1[3][69] ) );
  XOR U1614 ( .A(\w0[3][67] ), .B(g_input[451]), .Z(\w1[3][67] ) );
  XOR U1615 ( .A(\w0[3][62] ), .B(g_input[446]), .Z(\w1[3][62] ) );
  XOR U1616 ( .A(\w0[3][61] ), .B(g_input[445]), .Z(\w1[3][61] ) );
  XOR U1617 ( .A(\w0[3][5] ), .B(g_input[389]), .Z(\w1[3][5] ) );
  XOR U1618 ( .A(\w0[3][59] ), .B(g_input[443]), .Z(\w1[3][59] ) );
  XOR U1619 ( .A(\w0[3][54] ), .B(g_input[438]), .Z(\w1[3][54] ) );
  XOR U1620 ( .A(\w0[3][53] ), .B(g_input[437]), .Z(\w1[3][53] ) );
  XOR U1621 ( .A(\w0[3][51] ), .B(g_input[435]), .Z(\w1[3][51] ) );
  XOR U1622 ( .A(\w0[3][46] ), .B(g_input[430]), .Z(\w1[3][46] ) );
  XOR U1623 ( .A(\w0[3][45] ), .B(g_input[429]), .Z(\w1[3][45] ) );
  XOR U1624 ( .A(\w0[3][43] ), .B(g_input[427]), .Z(\w1[3][43] ) );
  XOR U1625 ( .A(\w0[3][3] ), .B(g_input[387]), .Z(\w1[3][3] ) );
  XOR U1626 ( .A(\w0[3][38] ), .B(g_input[422]), .Z(\w1[3][38] ) );
  XOR U1627 ( .A(\w0[3][37] ), .B(g_input[421]), .Z(\w1[3][37] ) );
  XOR U1628 ( .A(\w0[3][35] ), .B(g_input[419]), .Z(\w1[3][35] ) );
  XOR U1629 ( .A(\w0[3][30] ), .B(g_input[414]), .Z(\w1[3][30] ) );
  XOR U1630 ( .A(\w0[3][29] ), .B(g_input[413]), .Z(\w1[3][29] ) );
  XOR U1631 ( .A(\w0[3][27] ), .B(g_input[411]), .Z(\w1[3][27] ) );
  XOR U1632 ( .A(\w0[3][22] ), .B(g_input[406]), .Z(\w1[3][22] ) );
  XOR U1633 ( .A(\w0[3][21] ), .B(g_input[405]), .Z(\w1[3][21] ) );
  XOR U1634 ( .A(\w0[3][19] ), .B(g_input[403]), .Z(\w1[3][19] ) );
  XOR U1635 ( .A(\w0[3][14] ), .B(g_input[398]), .Z(\w1[3][14] ) );
  XOR U1636 ( .A(\w0[3][13] ), .B(g_input[397]), .Z(\w1[3][13] ) );
  XOR U1637 ( .A(\w0[3][126] ), .B(g_input[510]), .Z(\w1[3][126] ) );
  XOR U1638 ( .A(\w0[3][125] ), .B(g_input[509]), .Z(\w1[3][125] ) );
  XOR U1639 ( .A(\w0[3][123] ), .B(g_input[507]), .Z(\w1[3][123] ) );
  XOR U1640 ( .A(\w0[3][11] ), .B(g_input[395]), .Z(\w1[3][11] ) );
  XOR U1641 ( .A(\w0[3][118] ), .B(g_input[502]), .Z(\w1[3][118] ) );
  XOR U1642 ( .A(\w0[3][117] ), .B(g_input[501]), .Z(\w1[3][117] ) );
  XOR U1643 ( .A(\w0[3][115] ), .B(g_input[499]), .Z(\w1[3][115] ) );
  XOR U1644 ( .A(\w0[3][110] ), .B(g_input[494]), .Z(\w1[3][110] ) );
  XOR U1645 ( .A(\w0[3][109] ), .B(g_input[493]), .Z(\w1[3][109] ) );
  XOR U1646 ( .A(\w0[3][107] ), .B(g_input[491]), .Z(\w1[3][107] ) );
  XOR U1647 ( .A(\w0[3][102] ), .B(g_input[486]), .Z(\w1[3][102] ) );
  XOR U1648 ( .A(\w0[3][101] ), .B(g_input[485]), .Z(\w1[3][101] ) );
  XOR U1649 ( .A(\w0[2][99] ), .B(g_input[355]), .Z(\w1[2][99] ) );
  XOR U1650 ( .A(\w0[2][94] ), .B(g_input[350]), .Z(\w1[2][94] ) );
  XOR U1651 ( .A(\w0[2][93] ), .B(g_input[349]), .Z(\w1[2][93] ) );
  XOR U1652 ( .A(\w0[2][91] ), .B(g_input[347]), .Z(\w1[2][91] ) );
  XOR U1653 ( .A(\w0[2][86] ), .B(g_input[342]), .Z(\w1[2][86] ) );
  XOR U1654 ( .A(\w0[2][85] ), .B(g_input[341]), .Z(\w1[2][85] ) );
  XOR U1655 ( .A(\w0[2][83] ), .B(g_input[339]), .Z(\w1[2][83] ) );
  XOR U1656 ( .A(\w0[2][78] ), .B(g_input[334]), .Z(\w1[2][78] ) );
  XOR U1657 ( .A(\w0[2][77] ), .B(g_input[333]), .Z(\w1[2][77] ) );
  XOR U1658 ( .A(\w0[2][75] ), .B(g_input[331]), .Z(\w1[2][75] ) );
  XOR U1659 ( .A(\w0[2][70] ), .B(g_input[326]), .Z(\w1[2][70] ) );
  XOR U1660 ( .A(\w0[2][6] ), .B(g_input[262]), .Z(\w1[2][6] ) );
  XOR U1661 ( .A(\w0[2][69] ), .B(g_input[325]), .Z(\w1[2][69] ) );
  XOR U1662 ( .A(\w0[2][67] ), .B(g_input[323]), .Z(\w1[2][67] ) );
  XOR U1663 ( .A(\w0[2][62] ), .B(g_input[318]), .Z(\w1[2][62] ) );
  XOR U1664 ( .A(\w0[2][61] ), .B(g_input[317]), .Z(\w1[2][61] ) );
  XOR U1665 ( .A(\w0[2][5] ), .B(g_input[261]), .Z(\w1[2][5] ) );
  XOR U1666 ( .A(\w0[2][59] ), .B(g_input[315]), .Z(\w1[2][59] ) );
  XOR U1667 ( .A(\w0[2][54] ), .B(g_input[310]), .Z(\w1[2][54] ) );
  XOR U1668 ( .A(\w0[2][53] ), .B(g_input[309]), .Z(\w1[2][53] ) );
  XOR U1669 ( .A(\w0[2][51] ), .B(g_input[307]), .Z(\w1[2][51] ) );
  XOR U1670 ( .A(\w0[2][46] ), .B(g_input[302]), .Z(\w1[2][46] ) );
  XOR U1671 ( .A(\w0[2][45] ), .B(g_input[301]), .Z(\w1[2][45] ) );
  XOR U1672 ( .A(\w0[2][43] ), .B(g_input[299]), .Z(\w1[2][43] ) );
  XOR U1673 ( .A(\w0[2][3] ), .B(g_input[259]), .Z(\w1[2][3] ) );
  XOR U1674 ( .A(\w0[2][38] ), .B(g_input[294]), .Z(\w1[2][38] ) );
  XOR U1675 ( .A(\w0[2][37] ), .B(g_input[293]), .Z(\w1[2][37] ) );
  XOR U1676 ( .A(\w0[2][35] ), .B(g_input[291]), .Z(\w1[2][35] ) );
  XOR U1677 ( .A(\w0[2][30] ), .B(g_input[286]), .Z(\w1[2][30] ) );
  XOR U1678 ( .A(\w0[2][29] ), .B(g_input[285]), .Z(\w1[2][29] ) );
  XOR U1679 ( .A(\w0[2][27] ), .B(g_input[283]), .Z(\w1[2][27] ) );
  XOR U1680 ( .A(\w0[2][22] ), .B(g_input[278]), .Z(\w1[2][22] ) );
  XOR U1681 ( .A(\w0[2][21] ), .B(g_input[277]), .Z(\w1[2][21] ) );
  XOR U1682 ( .A(\w0[2][19] ), .B(g_input[275]), .Z(\w1[2][19] ) );
  XOR U1683 ( .A(\w0[2][14] ), .B(g_input[270]), .Z(\w1[2][14] ) );
  XOR U1684 ( .A(\w0[2][13] ), .B(g_input[269]), .Z(\w1[2][13] ) );
  XOR U1685 ( .A(\w0[2][126] ), .B(g_input[382]), .Z(\w1[2][126] ) );
  XOR U1686 ( .A(\w0[2][125] ), .B(g_input[381]), .Z(\w1[2][125] ) );
  XOR U1687 ( .A(\w0[2][123] ), .B(g_input[379]), .Z(\w1[2][123] ) );
  XOR U1688 ( .A(\w0[2][11] ), .B(g_input[267]), .Z(\w1[2][11] ) );
  XOR U1689 ( .A(\w0[2][118] ), .B(g_input[374]), .Z(\w1[2][118] ) );
  XOR U1690 ( .A(\w0[2][117] ), .B(g_input[373]), .Z(\w1[2][117] ) );
  XOR U1691 ( .A(\w0[2][115] ), .B(g_input[371]), .Z(\w1[2][115] ) );
  XOR U1692 ( .A(\w0[2][110] ), .B(g_input[366]), .Z(\w1[2][110] ) );
  XOR U1693 ( .A(\w0[2][109] ), .B(g_input[365]), .Z(\w1[2][109] ) );
  XOR U1694 ( .A(\w0[2][107] ), .B(g_input[363]), .Z(\w1[2][107] ) );
  XOR U1695 ( .A(\w0[2][102] ), .B(g_input[358]), .Z(\w1[2][102] ) );
  XOR U1696 ( .A(\w0[2][101] ), .B(g_input[357]), .Z(\w1[2][101] ) );
  XOR U1697 ( .A(\w0[1][99] ), .B(g_input[227]), .Z(\w1[1][99] ) );
  XOR U1698 ( .A(\w0[1][94] ), .B(g_input[222]), .Z(\w1[1][94] ) );
  XOR U1699 ( .A(\w0[1][93] ), .B(g_input[221]), .Z(\w1[1][93] ) );
  XOR U1700 ( .A(\w0[1][91] ), .B(g_input[219]), .Z(\w1[1][91] ) );
  XOR U1701 ( .A(\w0[1][86] ), .B(g_input[214]), .Z(\w1[1][86] ) );
  XOR U1702 ( .A(\w0[1][85] ), .B(g_input[213]), .Z(\w1[1][85] ) );
  XOR U1703 ( .A(\w0[1][83] ), .B(g_input[211]), .Z(\w1[1][83] ) );
  XOR U1704 ( .A(\w0[1][78] ), .B(g_input[206]), .Z(\w1[1][78] ) );
  XOR U1705 ( .A(\w0[1][77] ), .B(g_input[205]), .Z(\w1[1][77] ) );
  XOR U1706 ( .A(\w0[1][75] ), .B(g_input[203]), .Z(\w1[1][75] ) );
  XOR U1707 ( .A(\w0[1][70] ), .B(g_input[198]), .Z(\w1[1][70] ) );
  XOR U1708 ( .A(\w0[1][6] ), .B(g_input[134]), .Z(\w1[1][6] ) );
  XOR U1709 ( .A(\w0[1][69] ), .B(g_input[197]), .Z(\w1[1][69] ) );
  XOR U1710 ( .A(\w0[1][67] ), .B(g_input[195]), .Z(\w1[1][67] ) );
  XOR U1711 ( .A(\w0[1][62] ), .B(g_input[190]), .Z(\w1[1][62] ) );
  XOR U1712 ( .A(\w0[1][61] ), .B(g_input[189]), .Z(\w1[1][61] ) );
  XOR U1713 ( .A(\w0[1][5] ), .B(g_input[133]), .Z(\w1[1][5] ) );
  XOR U1714 ( .A(\w0[1][59] ), .B(g_input[187]), .Z(\w1[1][59] ) );
  XOR U1715 ( .A(\w0[1][54] ), .B(g_input[182]), .Z(\w1[1][54] ) );
  XOR U1716 ( .A(\w0[1][53] ), .B(g_input[181]), .Z(\w1[1][53] ) );
  XOR U1717 ( .A(\w0[1][51] ), .B(g_input[179]), .Z(\w1[1][51] ) );
  XOR U1718 ( .A(\w0[1][46] ), .B(g_input[174]), .Z(\w1[1][46] ) );
  XOR U1719 ( .A(\w0[1][45] ), .B(g_input[173]), .Z(\w1[1][45] ) );
  XOR U1720 ( .A(\w0[1][43] ), .B(g_input[171]), .Z(\w1[1][43] ) );
  XOR U1721 ( .A(\w0[1][3] ), .B(g_input[131]), .Z(\w1[1][3] ) );
  XOR U1722 ( .A(\w0[1][38] ), .B(g_input[166]), .Z(\w1[1][38] ) );
  XOR U1723 ( .A(\w0[1][37] ), .B(g_input[165]), .Z(\w1[1][37] ) );
  XOR U1724 ( .A(\w0[1][35] ), .B(g_input[163]), .Z(\w1[1][35] ) );
  XOR U1725 ( .A(\w0[1][30] ), .B(g_input[158]), .Z(\w1[1][30] ) );
  XOR U1726 ( .A(\w0[1][29] ), .B(g_input[157]), .Z(\w1[1][29] ) );
  XOR U1727 ( .A(\w0[1][27] ), .B(g_input[155]), .Z(\w1[1][27] ) );
  XOR U1728 ( .A(\w0[1][22] ), .B(g_input[150]), .Z(\w1[1][22] ) );
  XOR U1729 ( .A(\w0[1][21] ), .B(g_input[149]), .Z(\w1[1][21] ) );
  XOR U1730 ( .A(\w0[1][19] ), .B(g_input[147]), .Z(\w1[1][19] ) );
  XOR U1731 ( .A(\w0[1][14] ), .B(g_input[142]), .Z(\w1[1][14] ) );
  XOR U1732 ( .A(\w0[1][13] ), .B(g_input[141]), .Z(\w1[1][13] ) );
  XOR U1733 ( .A(\w0[1][126] ), .B(g_input[254]), .Z(\w1[1][126] ) );
  XOR U1734 ( .A(\w0[1][125] ), .B(g_input[253]), .Z(\w1[1][125] ) );
  XOR U1735 ( .A(\w0[1][123] ), .B(g_input[251]), .Z(\w1[1][123] ) );
  XOR U1736 ( .A(\w0[1][11] ), .B(g_input[139]), .Z(\w1[1][11] ) );
  XOR U1737 ( .A(\w0[1][118] ), .B(g_input[246]), .Z(\w1[1][118] ) );
  XOR U1738 ( .A(\w0[1][117] ), .B(g_input[245]), .Z(\w1[1][117] ) );
  XOR U1739 ( .A(\w0[1][115] ), .B(g_input[243]), .Z(\w1[1][115] ) );
  XOR U1740 ( .A(\w0[1][110] ), .B(g_input[238]), .Z(\w1[1][110] ) );
  XOR U1741 ( .A(\w0[1][109] ), .B(g_input[237]), .Z(\w1[1][109] ) );
  XOR U1742 ( .A(\w0[1][107] ), .B(g_input[235]), .Z(\w1[1][107] ) );
  XOR U1743 ( .A(\w0[1][102] ), .B(g_input[230]), .Z(\w1[1][102] ) );
  XOR U1744 ( .A(\w0[1][101] ), .B(g_input[229]), .Z(\w1[1][101] ) );
  XOR U1745 ( .A(g_input[99]), .B(e_input[99]), .Z(\w1[0][99] ) );
  XOR U1746 ( .A(g_input[94]), .B(e_input[94]), .Z(\w1[0][94] ) );
  XOR U1747 ( .A(g_input[93]), .B(e_input[93]), .Z(\w1[0][93] ) );
  XOR U1748 ( .A(g_input[91]), .B(e_input[91]), .Z(\w1[0][91] ) );
  XOR U1749 ( .A(g_input[86]), .B(e_input[86]), .Z(\w1[0][86] ) );
  XOR U1750 ( .A(g_input[85]), .B(e_input[85]), .Z(\w1[0][85] ) );
  XOR U1751 ( .A(g_input[83]), .B(e_input[83]), .Z(\w1[0][83] ) );
  XOR U1752 ( .A(g_input[78]), .B(e_input[78]), .Z(\w1[0][78] ) );
  XOR U1753 ( .A(g_input[77]), .B(e_input[77]), .Z(\w1[0][77] ) );
  XOR U1754 ( .A(g_input[75]), .B(e_input[75]), .Z(\w1[0][75] ) );
  XOR U1755 ( .A(g_input[70]), .B(e_input[70]), .Z(\w1[0][70] ) );
  XOR U1756 ( .A(g_input[6]), .B(e_input[6]), .Z(\w1[0][6] ) );
  XOR U1757 ( .A(g_input[69]), .B(e_input[69]), .Z(\w1[0][69] ) );
  XOR U1758 ( .A(g_input[67]), .B(e_input[67]), .Z(\w1[0][67] ) );
  XOR U1759 ( .A(g_input[62]), .B(e_input[62]), .Z(\w1[0][62] ) );
  XOR U1760 ( .A(g_input[61]), .B(e_input[61]), .Z(\w1[0][61] ) );
  XOR U1761 ( .A(g_input[5]), .B(e_input[5]), .Z(\w1[0][5] ) );
  XOR U1762 ( .A(g_input[59]), .B(e_input[59]), .Z(\w1[0][59] ) );
  XOR U1763 ( .A(g_input[54]), .B(e_input[54]), .Z(\w1[0][54] ) );
  XOR U1764 ( .A(g_input[53]), .B(e_input[53]), .Z(\w1[0][53] ) );
  XOR U1765 ( .A(g_input[51]), .B(e_input[51]), .Z(\w1[0][51] ) );
  XOR U1766 ( .A(g_input[46]), .B(e_input[46]), .Z(\w1[0][46] ) );
  XOR U1767 ( .A(g_input[45]), .B(e_input[45]), .Z(\w1[0][45] ) );
  XOR U1768 ( .A(g_input[43]), .B(e_input[43]), .Z(\w1[0][43] ) );
  XOR U1769 ( .A(g_input[3]), .B(e_input[3]), .Z(\w1[0][3] ) );
  XOR U1770 ( .A(g_input[38]), .B(e_input[38]), .Z(\w1[0][38] ) );
  XOR U1771 ( .A(g_input[37]), .B(e_input[37]), .Z(\w1[0][37] ) );
  XOR U1772 ( .A(g_input[35]), .B(e_input[35]), .Z(\w1[0][35] ) );
  XOR U1773 ( .A(g_input[30]), .B(e_input[30]), .Z(\w1[0][30] ) );
  XOR U1774 ( .A(g_input[29]), .B(e_input[29]), .Z(\w1[0][29] ) );
  XOR U1775 ( .A(g_input[27]), .B(e_input[27]), .Z(\w1[0][27] ) );
  XOR U1776 ( .A(g_input[22]), .B(e_input[22]), .Z(\w1[0][22] ) );
  XOR U1777 ( .A(g_input[21]), .B(e_input[21]), .Z(\w1[0][21] ) );
  XOR U1778 ( .A(g_input[19]), .B(e_input[19]), .Z(\w1[0][19] ) );
  XOR U1779 ( .A(g_input[14]), .B(e_input[14]), .Z(\w1[0][14] ) );
  XOR U1780 ( .A(g_input[13]), .B(e_input[13]), .Z(\w1[0][13] ) );
  XOR U1781 ( .A(g_input[126]), .B(e_input[126]), .Z(\w1[0][126] ) );
  XOR U1782 ( .A(g_input[125]), .B(e_input[125]), .Z(\w1[0][125] ) );
  XOR U1783 ( .A(g_input[123]), .B(e_input[123]), .Z(\w1[0][123] ) );
  XOR U1784 ( .A(g_input[11]), .B(e_input[11]), .Z(\w1[0][11] ) );
  XOR U1785 ( .A(g_input[118]), .B(e_input[118]), .Z(\w1[0][118] ) );
  XOR U1786 ( .A(g_input[117]), .B(e_input[117]), .Z(\w1[0][117] ) );
  XOR U1787 ( .A(g_input[115]), .B(e_input[115]), .Z(\w1[0][115] ) );
  XOR U1788 ( .A(g_input[110]), .B(e_input[110]), .Z(\w1[0][110] ) );
  XOR U1789 ( .A(g_input[109]), .B(e_input[109]), .Z(\w1[0][109] ) );
  XOR U1790 ( .A(g_input[107]), .B(e_input[107]), .Z(\w1[0][107] ) );
  XOR U1791 ( .A(g_input[102]), .B(e_input[102]), .Z(\w1[0][102] ) );
  XOR U1792 ( .A(g_input[101]), .B(e_input[101]), .Z(\w1[0][101] ) );
  XNOR U1793 ( .A(g_input[1161]), .B(n17409), .Z(o[9]) );
  XNOR U1794 ( .A(g_input[1251]), .B(n17339), .Z(o[99]) );
  XNOR U1795 ( .A(g_input[1250]), .B(n17338), .Z(o[98]) );
  XNOR U1796 ( .A(g_input[1249]), .B(n17337), .Z(o[97]) );
  XNOR U1797 ( .A(g_input[1248]), .B(n17336), .Z(o[96]) );
  XNOR U1798 ( .A(g_input[1247]), .B(n17431), .Z(o[95]) );
  XNOR U1799 ( .A(g_input[1246]), .B(n17430), .Z(o[94]) );
  XNOR U1800 ( .A(g_input[1245]), .B(n17429), .Z(o[93]) );
  XNOR U1801 ( .A(g_input[1244]), .B(n17428), .Z(o[92]) );
  XNOR U1802 ( .A(g_input[1243]), .B(n17427), .Z(o[91]) );
  XNOR U1803 ( .A(g_input[1242]), .B(n17426), .Z(o[90]) );
  XNOR U1804 ( .A(g_input[1160]), .B(n17408), .Z(o[8]) );
  XNOR U1805 ( .A(g_input[1241]), .B(n17425), .Z(o[89]) );
  XNOR U1806 ( .A(g_input[1240]), .B(n17424), .Z(o[88]) );
  XNOR U1807 ( .A(g_input[1239]), .B(n17391), .Z(o[87]) );
  XNOR U1808 ( .A(g_input[1238]), .B(n17390), .Z(o[86]) );
  XNOR U1809 ( .A(g_input[1237]), .B(n17389), .Z(o[85]) );
  XNOR U1810 ( .A(g_input[1236]), .B(n17388), .Z(o[84]) );
  XNOR U1811 ( .A(g_input[1235]), .B(n17387), .Z(o[83]) );
  XNOR U1812 ( .A(g_input[1234]), .B(n17386), .Z(o[82]) );
  XNOR U1813 ( .A(g_input[1233]), .B(n17385), .Z(o[81]) );
  XNOR U1814 ( .A(g_input[1232]), .B(n17384), .Z(o[80]) );
  XNOR U1815 ( .A(g_input[1159]), .B(n17375), .Z(o[7]) );
  XNOR U1816 ( .A(g_input[1231]), .B(n17351), .Z(o[79]) );
  XNOR U1817 ( .A(g_input[1230]), .B(n17350), .Z(o[78]) );
  XNOR U1818 ( .A(g_input[1229]), .B(n17349), .Z(o[77]) );
  XNOR U1819 ( .A(g_input[1228]), .B(n17348), .Z(o[76]) );
  XNOR U1820 ( .A(g_input[1227]), .B(n17347), .Z(o[75]) );
  XNOR U1821 ( .A(g_input[1226]), .B(n17346), .Z(o[74]) );
  XNOR U1822 ( .A(g_input[1225]), .B(n17345), .Z(o[73]) );
  XNOR U1823 ( .A(g_input[1224]), .B(n17344), .Z(o[72]) );
  XNOR U1824 ( .A(g_input[1223]), .B(n17439), .Z(o[71]) );
  XNOR U1825 ( .A(g_input[1222]), .B(n17438), .Z(o[70]) );
  XNOR U1826 ( .A(g_input[1158]), .B(n17374), .Z(o[6]) );
  XNOR U1827 ( .A(g_input[1221]), .B(n17437), .Z(o[69]) );
  XNOR U1828 ( .A(g_input[1220]), .B(n17436), .Z(o[68]) );
  XNOR U1829 ( .A(g_input[1219]), .B(n17435), .Z(o[67]) );
  XNOR U1830 ( .A(g_input[1218]), .B(n17434), .Z(o[66]) );
  XNOR U1831 ( .A(g_input[1217]), .B(n17433), .Z(o[65]) );
  XNOR U1832 ( .A(g_input[1216]), .B(n17432), .Z(o[64]) );
  XNOR U1833 ( .A(g_input[1215]), .B(n17399), .Z(o[63]) );
  XNOR U1834 ( .A(g_input[1214]), .B(n17398), .Z(o[62]) );
  XNOR U1835 ( .A(g_input[1213]), .B(n17397), .Z(o[61]) );
  XNOR U1836 ( .A(g_input[1212]), .B(n17396), .Z(o[60]) );
  XNOR U1837 ( .A(g_input[1157]), .B(n17373), .Z(o[5]) );
  XNOR U1838 ( .A(g_input[1211]), .B(n17395), .Z(o[59]) );
  XNOR U1839 ( .A(g_input[1210]), .B(n17394), .Z(o[58]) );
  XNOR U1840 ( .A(g_input[1209]), .B(n17393), .Z(o[57]) );
  XNOR U1841 ( .A(g_input[1208]), .B(n17392), .Z(o[56]) );
  XNOR U1842 ( .A(g_input[1207]), .B(n17359), .Z(o[55]) );
  XNOR U1843 ( .A(g_input[1206]), .B(n17358), .Z(o[54]) );
  XNOR U1844 ( .A(g_input[1205]), .B(n17357), .Z(o[53]) );
  XNOR U1845 ( .A(g_input[1204]), .B(n17356), .Z(o[52]) );
  XNOR U1846 ( .A(g_input[1203]), .B(n17355), .Z(o[51]) );
  XNOR U1847 ( .A(g_input[1202]), .B(n17354), .Z(o[50]) );
  XNOR U1848 ( .A(g_input[1156]), .B(n17372), .Z(o[4]) );
  XNOR U1849 ( .A(g_input[1201]), .B(n17353), .Z(o[49]) );
  XNOR U1850 ( .A(g_input[1200]), .B(n17352), .Z(o[48]) );
  XNOR U1851 ( .A(g_input[1199]), .B(n17447), .Z(o[47]) );
  XNOR U1852 ( .A(g_input[1198]), .B(n17446), .Z(o[46]) );
  XNOR U1853 ( .A(g_input[1197]), .B(n17445), .Z(o[45]) );
  XNOR U1854 ( .A(g_input[1196]), .B(n17444), .Z(o[44]) );
  XNOR U1855 ( .A(g_input[1195]), .B(n17443), .Z(o[43]) );
  XNOR U1856 ( .A(g_input[1194]), .B(n17442), .Z(o[42]) );
  XNOR U1857 ( .A(g_input[1193]), .B(n17441), .Z(o[41]) );
  XNOR U1858 ( .A(g_input[1192]), .B(n17440), .Z(o[40]) );
  XNOR U1859 ( .A(g_input[1155]), .B(n17371), .Z(o[3]) );
  XNOR U1860 ( .A(g_input[1191]), .B(n17407), .Z(o[39]) );
  XNOR U1861 ( .A(g_input[1190]), .B(n17406), .Z(o[38]) );
  XNOR U1862 ( .A(g_input[1189]), .B(n17405), .Z(o[37]) );
  XNOR U1863 ( .A(g_input[1188]), .B(n17404), .Z(o[36]) );
  XNOR U1864 ( .A(g_input[1187]), .B(n17403), .Z(o[35]) );
  XNOR U1865 ( .A(g_input[1186]), .B(n17402), .Z(o[34]) );
  XNOR U1866 ( .A(g_input[1185]), .B(n17401), .Z(o[33]) );
  XNOR U1867 ( .A(g_input[1184]), .B(n17400), .Z(o[32]) );
  XNOR U1868 ( .A(g_input[1183]), .B(n17367), .Z(o[31]) );
  XNOR U1869 ( .A(g_input[1182]), .B(n17366), .Z(o[30]) );
  XNOR U1870 ( .A(g_input[1154]), .B(n17370), .Z(o[2]) );
  XNOR U1871 ( .A(g_input[1181]), .B(n17365), .Z(o[29]) );
  XNOR U1872 ( .A(g_input[1180]), .B(n17364), .Z(o[28]) );
  XNOR U1873 ( .A(g_input[1179]), .B(n17363), .Z(o[27]) );
  XNOR U1874 ( .A(g_input[1178]), .B(n17362), .Z(o[26]) );
  XNOR U1875 ( .A(g_input[1177]), .B(n17361), .Z(o[25]) );
  XNOR U1876 ( .A(g_input[1176]), .B(n17360), .Z(o[24]) );
  XNOR U1877 ( .A(g_input[1175]), .B(n17455), .Z(o[23]) );
  XNOR U1878 ( .A(g_input[1174]), .B(n17454), .Z(o[22]) );
  XNOR U1879 ( .A(g_input[1173]), .B(n17453), .Z(o[21]) );
  XNOR U1880 ( .A(g_input[1172]), .B(n17452), .Z(o[20]) );
  XNOR U1881 ( .A(g_input[1153]), .B(n17369), .Z(o[1]) );
  XNOR U1882 ( .A(g_input[1171]), .B(n17451), .Z(o[19]) );
  XNOR U1883 ( .A(g_input[1170]), .B(n17450), .Z(o[18]) );
  XNOR U1884 ( .A(g_input[1169]), .B(n17449), .Z(o[17]) );
  XNOR U1885 ( .A(g_input[1168]), .B(n17448), .Z(o[16]) );
  XNOR U1886 ( .A(g_input[1167]), .B(n17415), .Z(o[15]) );
  XNOR U1887 ( .A(g_input[1166]), .B(n17414), .Z(o[14]) );
  XNOR U1888 ( .A(g_input[1165]), .B(n17413), .Z(o[13]) );
  XNOR U1889 ( .A(g_input[1164]), .B(n17412), .Z(o[12]) );
  XNOR U1890 ( .A(g_input[1279]), .B(n17463), .Z(o[127]) );
  XNOR U1891 ( .A(g_input[1278]), .B(n17462), .Z(o[126]) );
  XNOR U1892 ( .A(g_input[1277]), .B(n17461), .Z(o[125]) );
  XNOR U1893 ( .A(g_input[1276]), .B(n17460), .Z(o[124]) );
  XNOR U1894 ( .A(g_input[1275]), .B(n17459), .Z(o[123]) );
  XNOR U1895 ( .A(g_input[1274]), .B(n17458), .Z(o[122]) );
  XNOR U1896 ( .A(g_input[1273]), .B(n17457), .Z(o[121]) );
  XNOR U1897 ( .A(g_input[1272]), .B(n17456), .Z(o[120]) );
  XNOR U1898 ( .A(g_input[1163]), .B(n17411), .Z(o[11]) );
  XNOR U1899 ( .A(g_input[1271]), .B(n17423), .Z(o[119]) );
  XNOR U1900 ( .A(g_input[1270]), .B(n17422), .Z(o[118]) );
  XNOR U1901 ( .A(g_input[1269]), .B(n17421), .Z(o[117]) );
  XNOR U1902 ( .A(g_input[1268]), .B(n17420), .Z(o[116]) );
  XNOR U1903 ( .A(g_input[1267]), .B(n17419), .Z(o[115]) );
  XNOR U1904 ( .A(g_input[1266]), .B(n17418), .Z(o[114]) );
  XNOR U1905 ( .A(g_input[1265]), .B(n17417), .Z(o[113]) );
  XNOR U1906 ( .A(g_input[1264]), .B(n17416), .Z(o[112]) );
  XNOR U1907 ( .A(g_input[1263]), .B(n17383), .Z(o[111]) );
  XNOR U1908 ( .A(g_input[1262]), .B(n17382), .Z(o[110]) );
  XNOR U1909 ( .A(g_input[1162]), .B(n17410), .Z(o[10]) );
  XNOR U1910 ( .A(g_input[1261]), .B(n17381), .Z(o[109]) );
  XNOR U1911 ( .A(g_input[1260]), .B(n17380), .Z(o[108]) );
  XNOR U1912 ( .A(g_input[1259]), .B(n17379), .Z(o[107]) );
  XNOR U1913 ( .A(g_input[1258]), .B(n17378), .Z(o[106]) );
  XNOR U1914 ( .A(g_input[1257]), .B(n17377), .Z(o[105]) );
  XNOR U1915 ( .A(g_input[1256]), .B(n17376), .Z(o[104]) );
  XNOR U1916 ( .A(g_input[1255]), .B(n17343), .Z(o[103]) );
  XNOR U1917 ( .A(g_input[1254]), .B(n17342), .Z(o[102]) );
  XNOR U1918 ( .A(g_input[1253]), .B(n17341), .Z(o[101]) );
  XNOR U1919 ( .A(g_input[1252]), .B(n17340), .Z(o[100]) );
  XNOR U1920 ( .A(g_input[1152]), .B(n17368), .Z(o[0]) );
  AND U1921 ( .A(n1169), .B(\SUBBYTES[9].a/w781 ), .Z(\SUBBYTES[9].a/w916 ) );
  AND U1922 ( .A(n1170), .B(\SUBBYTES[9].a/w782 ), .Z(\SUBBYTES[9].a/w914 ) );
  AND U1923 ( .A(\SUBBYTES[9].a/w912 ), .B(n1171), .Z(\SUBBYTES[9].a/w913 ) );
  ANDN U1924 ( .A(\w1[9][96] ), .B(n1172), .Z(\SUBBYTES[9].a/w909 ) );
  AND U1925 ( .A(n1173), .B(\SUBBYTES[9].a/w784 ), .Z(\SUBBYTES[9].a/w907 ) );
  AND U1926 ( .A(\SUBBYTES[9].a/w905 ), .B(n1174), .Z(\SUBBYTES[9].a/w906 ) );
  XOR U1927 ( .A(\SUBBYTES[9].a/w849 ), .B(n16078), .Z(n1174) );
  AND U1928 ( .A(\SUBBYTES[9].a/w892 ), .B(\SUBBYTES[9].a/w894 ), .Z(
        \SUBBYTES[9].a/w901 ) );
  AND U1929 ( .A(\SUBBYTES[9].a/w893 ), .B(\SUBBYTES[9].a/w895 ), .Z(
        \SUBBYTES[9].a/w899 ) );
  AND U1930 ( .A(\SUBBYTES[9].a/w896 ), .B(\SUBBYTES[9].a/w897 ), .Z(
        \SUBBYTES[9].a/w898 ) );
  AND U1931 ( .A(\SUBBYTES[9].a/w785 ), .B(n1169), .Z(\SUBBYTES[9].a/w884 ) );
  XOR U1932 ( .A(\SUBBYTES[9].a/w853 ), .B(n1088), .Z(n1169) );
  AND U1933 ( .A(\SUBBYTES[9].a/w786 ), .B(n1170), .Z(\SUBBYTES[9].a/w882 ) );
  XOR U1934 ( .A(n16079), .B(\SUBBYTES[9].a/w853 ), .Z(n1170) );
  ANDN U1935 ( .A(n1171), .B(n1175), .Z(\SUBBYTES[9].a/w881 ) );
  XOR U1936 ( .A(n1088), .B(n16079), .Z(n1171) );
  ANDN U1937 ( .A(\SUBBYTES[9].a/w787 ), .B(n1172), .Z(\SUBBYTES[9].a/w877 )
         );
  XNOR U1938 ( .A(\SUBBYTES[9].a/w846 ), .B(\SUBBYTES[9].a/w849 ), .Z(n1172)
         );
  AND U1939 ( .A(\SUBBYTES[9].a/w788 ), .B(n1173), .Z(\SUBBYTES[9].a/w875 ) );
  XNOR U1940 ( .A(n1176), .B(\SUBBYTES[9].a/w846 ), .Z(n1173) );
  AND U1941 ( .A(\SUBBYTES[9].a/w873 ), .B(n1177), .Z(\SUBBYTES[9].a/w874 ) );
  XOR U1942 ( .A(n1178), .B(n1176), .Z(n1177) );
  IV U1943 ( .A(n16078), .Z(n1176) );
  ANDN U1944 ( .A(\SUBBYTES[9].a/w892 ), .B(n1179), .Z(\SUBBYTES[9].a/w869 )
         );
  ANDN U1945 ( .A(\SUBBYTES[9].a/w893 ), .B(n1180), .Z(\SUBBYTES[9].a/w867 )
         );
  AND U1946 ( .A(n1181), .B(\SUBBYTES[9].a/w896 ), .Z(\SUBBYTES[9].a/w866 ) );
  AND U1947 ( .A(\SUBBYTES[9].a/w852 ), .B(\SUBBYTES[9].a/w851 ), .Z(
        \SUBBYTES[9].a/w853 ) );
  IV U1948 ( .A(n1178), .Z(\SUBBYTES[9].a/w849 ) );
  NAND U1949 ( .A(\SUBBYTES[9].a/w828 ), .B(\SUBBYTES[9].a/w843 ), .Z(n1178)
         );
  AND U1950 ( .A(\SUBBYTES[9].a/w845 ), .B(\SUBBYTES[9].a/w851 ), .Z(
        \SUBBYTES[9].a/w846 ) );
  AND U1951 ( .A(\SUBBYTES[9].a/w830 ), .B(\SUBBYTES[9].a/w828 ), .Z(
        \SUBBYTES[9].a/w840 ) );
  AND U1952 ( .A(\SUBBYTES[9].a/w831 ), .B(\SUBBYTES[9].a/w829 ), .Z(
        \SUBBYTES[9].a/w838 ) );
  AND U1953 ( .A(\SUBBYTES[9].a/w845 ), .B(\SUBBYTES[9].a/w852 ), .Z(
        \SUBBYTES[9].a/w837 ) );
  AND U1954 ( .A(\SUBBYTES[9].a/w785 ), .B(\SUBBYTES[9].a/w781 ), .Z(
        \SUBBYTES[9].a/w822 ) );
  AND U1955 ( .A(\SUBBYTES[9].a/w786 ), .B(\SUBBYTES[9].a/w782 ), .Z(
        \SUBBYTES[9].a/w820 ) );
  ANDN U1956 ( .A(\SUBBYTES[9].a/w912 ), .B(n1175), .Z(\SUBBYTES[9].a/w819 )
         );
  XNOR U1957 ( .A(\w1[9][103] ), .B(\w1[9][97] ), .Z(n1175) );
  XOR U1958 ( .A(g_input[1249]), .B(\w0[9][97] ), .Z(\w1[9][97] ) );
  IV U1959 ( .A(n1182), .Z(\w1[9][103] ) );
  AND U1960 ( .A(\w1[9][96] ), .B(\SUBBYTES[9].a/w787 ), .Z(
        \SUBBYTES[9].a/w815 ) );
  XOR U1961 ( .A(g_input[1248]), .B(\w0[9][96] ), .Z(\w1[9][96] ) );
  AND U1962 ( .A(\SUBBYTES[9].a/w788 ), .B(\SUBBYTES[9].a/w784 ), .Z(
        \SUBBYTES[9].a/w813 ) );
  AND U1963 ( .A(\SUBBYTES[9].a/w873 ), .B(\SUBBYTES[9].a/w905 ), .Z(
        \SUBBYTES[9].a/w812 ) );
  ANDN U1964 ( .A(\SUBBYTES[9].a/w894 ), .B(n1179), .Z(\SUBBYTES[9].a/w807 )
         );
  XOR U1965 ( .A(\w1[9][100] ), .B(n1182), .Z(n1179) );
  ANDN U1966 ( .A(\SUBBYTES[9].a/w895 ), .B(n1180), .Z(\SUBBYTES[9].a/w805 )
         );
  XOR U1967 ( .A(n1182), .B(\w1[9][98] ), .Z(n1180) );
  XNOR U1968 ( .A(g_input[1255]), .B(\w0[9][103] ), .Z(n1182) );
  AND U1969 ( .A(\SUBBYTES[9].a/w897 ), .B(n1181), .Z(\SUBBYTES[9].a/w804 ) );
  XOR U1970 ( .A(\w1[9][100] ), .B(\w1[9][98] ), .Z(n1181) );
  XOR U1971 ( .A(g_input[1250]), .B(\w0[9][98] ), .Z(\w1[9][98] ) );
  XOR U1972 ( .A(g_input[1252]), .B(\w0[9][100] ), .Z(\w1[9][100] ) );
  AND U1973 ( .A(n1183), .B(\SUBBYTES[9].a/w574 ), .Z(\SUBBYTES[9].a/w709 ) );
  AND U1974 ( .A(n1184), .B(\SUBBYTES[9].a/w575 ), .Z(\SUBBYTES[9].a/w707 ) );
  AND U1975 ( .A(\SUBBYTES[9].a/w705 ), .B(n1185), .Z(\SUBBYTES[9].a/w706 ) );
  ANDN U1976 ( .A(\w1[9][104] ), .B(n1186), .Z(\SUBBYTES[9].a/w702 ) );
  AND U1977 ( .A(n1187), .B(\SUBBYTES[9].a/w577 ), .Z(\SUBBYTES[9].a/w700 ) );
  AND U1978 ( .A(\SUBBYTES[9].a/w698 ), .B(n1188), .Z(\SUBBYTES[9].a/w699 ) );
  XOR U1979 ( .A(\SUBBYTES[9].a/w642 ), .B(n16076), .Z(n1188) );
  AND U1980 ( .A(\SUBBYTES[9].a/w685 ), .B(\SUBBYTES[9].a/w687 ), .Z(
        \SUBBYTES[9].a/w694 ) );
  AND U1981 ( .A(\SUBBYTES[9].a/w686 ), .B(\SUBBYTES[9].a/w688 ), .Z(
        \SUBBYTES[9].a/w692 ) );
  AND U1982 ( .A(\SUBBYTES[9].a/w689 ), .B(\SUBBYTES[9].a/w690 ), .Z(
        \SUBBYTES[9].a/w691 ) );
  AND U1983 ( .A(\SUBBYTES[9].a/w578 ), .B(n1183), .Z(\SUBBYTES[9].a/w677 ) );
  XOR U1984 ( .A(\SUBBYTES[9].a/w646 ), .B(n1087), .Z(n1183) );
  AND U1985 ( .A(\SUBBYTES[9].a/w579 ), .B(n1184), .Z(\SUBBYTES[9].a/w675 ) );
  XOR U1986 ( .A(n16077), .B(\SUBBYTES[9].a/w646 ), .Z(n1184) );
  AND U1987 ( .A(n1189), .B(n1185), .Z(\SUBBYTES[9].a/w674 ) );
  XOR U1988 ( .A(n1087), .B(n16077), .Z(n1185) );
  ANDN U1989 ( .A(\SUBBYTES[9].a/w580 ), .B(n1186), .Z(\SUBBYTES[9].a/w670 )
         );
  XNOR U1990 ( .A(\SUBBYTES[9].a/w639 ), .B(\SUBBYTES[9].a/w642 ), .Z(n1186)
         );
  AND U1991 ( .A(\SUBBYTES[9].a/w581 ), .B(n1187), .Z(\SUBBYTES[9].a/w668 ) );
  XNOR U1992 ( .A(n1190), .B(\SUBBYTES[9].a/w639 ), .Z(n1187) );
  AND U1993 ( .A(\SUBBYTES[9].a/w666 ), .B(n1191), .Z(\SUBBYTES[9].a/w667 ) );
  XOR U1994 ( .A(n1192), .B(n1190), .Z(n1191) );
  IV U1995 ( .A(n16076), .Z(n1190) );
  AND U1996 ( .A(n1193), .B(\SUBBYTES[9].a/w685 ), .Z(\SUBBYTES[9].a/w662 ) );
  ANDN U1997 ( .A(\SUBBYTES[9].a/w686 ), .B(n1194), .Z(\SUBBYTES[9].a/w660 )
         );
  AND U1998 ( .A(n1195), .B(\SUBBYTES[9].a/w689 ), .Z(\SUBBYTES[9].a/w659 ) );
  AND U1999 ( .A(\SUBBYTES[9].a/w645 ), .B(\SUBBYTES[9].a/w644 ), .Z(
        \SUBBYTES[9].a/w646 ) );
  IV U2000 ( .A(n1192), .Z(\SUBBYTES[9].a/w642 ) );
  NAND U2001 ( .A(\SUBBYTES[9].a/w621 ), .B(\SUBBYTES[9].a/w636 ), .Z(n1192)
         );
  AND U2002 ( .A(\SUBBYTES[9].a/w638 ), .B(\SUBBYTES[9].a/w644 ), .Z(
        \SUBBYTES[9].a/w639 ) );
  AND U2003 ( .A(\SUBBYTES[9].a/w623 ), .B(\SUBBYTES[9].a/w621 ), .Z(
        \SUBBYTES[9].a/w633 ) );
  AND U2004 ( .A(\SUBBYTES[9].a/w624 ), .B(\SUBBYTES[9].a/w622 ), .Z(
        \SUBBYTES[9].a/w631 ) );
  AND U2005 ( .A(\SUBBYTES[9].a/w638 ), .B(\SUBBYTES[9].a/w645 ), .Z(
        \SUBBYTES[9].a/w630 ) );
  AND U2006 ( .A(\SUBBYTES[9].a/w578 ), .B(\SUBBYTES[9].a/w574 ), .Z(
        \SUBBYTES[9].a/w615 ) );
  AND U2007 ( .A(\SUBBYTES[9].a/w579 ), .B(\SUBBYTES[9].a/w575 ), .Z(
        \SUBBYTES[9].a/w613 ) );
  AND U2008 ( .A(\SUBBYTES[9].a/w705 ), .B(n1189), .Z(\SUBBYTES[9].a/w612 ) );
  XNOR U2009 ( .A(\w1[9][105] ), .B(n1196), .Z(n1189) );
  XOR U2010 ( .A(g_input[1257]), .B(\w0[9][105] ), .Z(\w1[9][105] ) );
  AND U2011 ( .A(\w1[9][104] ), .B(\SUBBYTES[9].a/w580 ), .Z(
        \SUBBYTES[9].a/w608 ) );
  XOR U2012 ( .A(g_input[1256]), .B(\w0[9][104] ), .Z(\w1[9][104] ) );
  AND U2013 ( .A(\SUBBYTES[9].a/w581 ), .B(\SUBBYTES[9].a/w577 ), .Z(
        \SUBBYTES[9].a/w606 ) );
  AND U2014 ( .A(\SUBBYTES[9].a/w666 ), .B(\SUBBYTES[9].a/w698 ), .Z(
        \SUBBYTES[9].a/w605 ) );
  AND U2015 ( .A(\SUBBYTES[9].a/w687 ), .B(n1193), .Z(\SUBBYTES[9].a/w600 ) );
  XOR U2016 ( .A(\w1[9][108] ), .B(\w1[9][111] ), .Z(n1193) );
  ANDN U2017 ( .A(\SUBBYTES[9].a/w688 ), .B(n1194), .Z(\SUBBYTES[9].a/w598 )
         );
  XNOR U2018 ( .A(\w1[9][106] ), .B(\w1[9][111] ), .Z(n1194) );
  IV U2019 ( .A(n1196), .Z(\w1[9][111] ) );
  XNOR U2020 ( .A(g_input[1263]), .B(\w0[9][111] ), .Z(n1196) );
  AND U2021 ( .A(\SUBBYTES[9].a/w690 ), .B(n1195), .Z(\SUBBYTES[9].a/w597 ) );
  XOR U2022 ( .A(\w1[9][106] ), .B(\w1[9][108] ), .Z(n1195) );
  XOR U2023 ( .A(g_input[1260]), .B(\w0[9][108] ), .Z(\w1[9][108] ) );
  XOR U2024 ( .A(g_input[1258]), .B(\w0[9][106] ), .Z(\w1[9][106] ) );
  AND U2025 ( .A(n1197), .B(\SUBBYTES[9].a/w367 ), .Z(\SUBBYTES[9].a/w502 ) );
  AND U2026 ( .A(n1198), .B(\SUBBYTES[9].a/w368 ), .Z(\SUBBYTES[9].a/w500 ) );
  AND U2027 ( .A(\SUBBYTES[9].a/w498 ), .B(n1199), .Z(\SUBBYTES[9].a/w499 ) );
  ANDN U2028 ( .A(\w1[9][112] ), .B(n1200), .Z(\SUBBYTES[9].a/w495 ) );
  AND U2029 ( .A(n1201), .B(\SUBBYTES[9].a/w370 ), .Z(\SUBBYTES[9].a/w493 ) );
  AND U2030 ( .A(\SUBBYTES[9].a/w491 ), .B(n1202), .Z(\SUBBYTES[9].a/w492 ) );
  XOR U2031 ( .A(\SUBBYTES[9].a/w435 ), .B(n16074), .Z(n1202) );
  AND U2032 ( .A(\SUBBYTES[9].a/w478 ), .B(\SUBBYTES[9].a/w480 ), .Z(
        \SUBBYTES[9].a/w487 ) );
  AND U2033 ( .A(\SUBBYTES[9].a/w479 ), .B(\SUBBYTES[9].a/w481 ), .Z(
        \SUBBYTES[9].a/w485 ) );
  AND U2034 ( .A(\SUBBYTES[9].a/w482 ), .B(\SUBBYTES[9].a/w483 ), .Z(
        \SUBBYTES[9].a/w484 ) );
  AND U2035 ( .A(\SUBBYTES[9].a/w371 ), .B(n1197), .Z(\SUBBYTES[9].a/w470 ) );
  XOR U2036 ( .A(\SUBBYTES[9].a/w439 ), .B(n1086), .Z(n1197) );
  AND U2037 ( .A(\SUBBYTES[9].a/w372 ), .B(n1198), .Z(\SUBBYTES[9].a/w468 ) );
  XOR U2038 ( .A(n16075), .B(\SUBBYTES[9].a/w439 ), .Z(n1198) );
  AND U2039 ( .A(n1203), .B(n1199), .Z(\SUBBYTES[9].a/w467 ) );
  XOR U2040 ( .A(n1086), .B(n16075), .Z(n1199) );
  ANDN U2041 ( .A(\SUBBYTES[9].a/w373 ), .B(n1200), .Z(\SUBBYTES[9].a/w463 )
         );
  XNOR U2042 ( .A(\SUBBYTES[9].a/w432 ), .B(\SUBBYTES[9].a/w435 ), .Z(n1200)
         );
  AND U2043 ( .A(\SUBBYTES[9].a/w374 ), .B(n1201), .Z(\SUBBYTES[9].a/w461 ) );
  XNOR U2044 ( .A(n1204), .B(\SUBBYTES[9].a/w432 ), .Z(n1201) );
  AND U2045 ( .A(\SUBBYTES[9].a/w459 ), .B(n1205), .Z(\SUBBYTES[9].a/w460 ) );
  XOR U2046 ( .A(n1206), .B(n1204), .Z(n1205) );
  IV U2047 ( .A(n16074), .Z(n1204) );
  AND U2048 ( .A(n1207), .B(\SUBBYTES[9].a/w478 ), .Z(\SUBBYTES[9].a/w455 ) );
  ANDN U2049 ( .A(\SUBBYTES[9].a/w479 ), .B(n1208), .Z(\SUBBYTES[9].a/w453 )
         );
  AND U2050 ( .A(n1209), .B(\SUBBYTES[9].a/w482 ), .Z(\SUBBYTES[9].a/w452 ) );
  AND U2051 ( .A(\SUBBYTES[9].a/w438 ), .B(\SUBBYTES[9].a/w437 ), .Z(
        \SUBBYTES[9].a/w439 ) );
  IV U2052 ( .A(n1206), .Z(\SUBBYTES[9].a/w435 ) );
  NAND U2053 ( .A(\SUBBYTES[9].a/w414 ), .B(\SUBBYTES[9].a/w429 ), .Z(n1206)
         );
  AND U2054 ( .A(\SUBBYTES[9].a/w431 ), .B(\SUBBYTES[9].a/w437 ), .Z(
        \SUBBYTES[9].a/w432 ) );
  AND U2055 ( .A(\SUBBYTES[9].a/w416 ), .B(\SUBBYTES[9].a/w414 ), .Z(
        \SUBBYTES[9].a/w426 ) );
  AND U2056 ( .A(\SUBBYTES[9].a/w417 ), .B(\SUBBYTES[9].a/w415 ), .Z(
        \SUBBYTES[9].a/w424 ) );
  AND U2057 ( .A(\SUBBYTES[9].a/w431 ), .B(\SUBBYTES[9].a/w438 ), .Z(
        \SUBBYTES[9].a/w423 ) );
  AND U2058 ( .A(\SUBBYTES[9].a/w371 ), .B(\SUBBYTES[9].a/w367 ), .Z(
        \SUBBYTES[9].a/w408 ) );
  AND U2059 ( .A(\SUBBYTES[9].a/w372 ), .B(\SUBBYTES[9].a/w368 ), .Z(
        \SUBBYTES[9].a/w406 ) );
  AND U2060 ( .A(\SUBBYTES[9].a/w498 ), .B(n1203), .Z(\SUBBYTES[9].a/w405 ) );
  XNOR U2061 ( .A(\w1[9][113] ), .B(n1210), .Z(n1203) );
  XOR U2062 ( .A(g_input[1265]), .B(\w0[9][113] ), .Z(\w1[9][113] ) );
  AND U2063 ( .A(\w1[9][112] ), .B(\SUBBYTES[9].a/w373 ), .Z(
        \SUBBYTES[9].a/w401 ) );
  XOR U2064 ( .A(g_input[1264]), .B(\w0[9][112] ), .Z(\w1[9][112] ) );
  AND U2065 ( .A(\SUBBYTES[9].a/w374 ), .B(\SUBBYTES[9].a/w370 ), .Z(
        \SUBBYTES[9].a/w399 ) );
  AND U2066 ( .A(\SUBBYTES[9].a/w459 ), .B(\SUBBYTES[9].a/w491 ), .Z(
        \SUBBYTES[9].a/w398 ) );
  AND U2067 ( .A(\SUBBYTES[9].a/w480 ), .B(n1207), .Z(\SUBBYTES[9].a/w393 ) );
  XOR U2068 ( .A(\w1[9][116] ), .B(\w1[9][119] ), .Z(n1207) );
  ANDN U2069 ( .A(\SUBBYTES[9].a/w481 ), .B(n1208), .Z(\SUBBYTES[9].a/w391 )
         );
  XNOR U2070 ( .A(\w1[9][114] ), .B(\w1[9][119] ), .Z(n1208) );
  IV U2071 ( .A(n1210), .Z(\w1[9][119] ) );
  XNOR U2072 ( .A(g_input[1271]), .B(\w0[9][119] ), .Z(n1210) );
  AND U2073 ( .A(\SUBBYTES[9].a/w483 ), .B(n1209), .Z(\SUBBYTES[9].a/w390 ) );
  XOR U2074 ( .A(\w1[9][114] ), .B(\w1[9][116] ), .Z(n1209) );
  XOR U2075 ( .A(g_input[1268]), .B(\w0[9][116] ), .Z(\w1[9][116] ) );
  XOR U2076 ( .A(g_input[1266]), .B(\w0[9][114] ), .Z(\w1[9][114] ) );
  AND U2077 ( .A(n1211), .B(\SUBBYTES[9].a/w3265 ), .Z(\SUBBYTES[9].a/w3400 )
         );
  AND U2078 ( .A(n1212), .B(\SUBBYTES[9].a/w3266 ), .Z(\SUBBYTES[9].a/w3398 )
         );
  AND U2079 ( .A(\SUBBYTES[9].a/w3396 ), .B(n1213), .Z(\SUBBYTES[9].a/w3397 )
         );
  ANDN U2080 ( .A(\w1[9][0] ), .B(n1214), .Z(\SUBBYTES[9].a/w3393 ) );
  AND U2081 ( .A(n1215), .B(\SUBBYTES[9].a/w3268 ), .Z(\SUBBYTES[9].a/w3391 )
         );
  AND U2082 ( .A(\SUBBYTES[9].a/w3389 ), .B(n1216), .Z(\SUBBYTES[9].a/w3390 )
         );
  XOR U2083 ( .A(\SUBBYTES[9].a/w3333 ), .B(n16102), .Z(n1216) );
  AND U2084 ( .A(\SUBBYTES[9].a/w3376 ), .B(\SUBBYTES[9].a/w3378 ), .Z(
        \SUBBYTES[9].a/w3385 ) );
  AND U2085 ( .A(\SUBBYTES[9].a/w3377 ), .B(\SUBBYTES[9].a/w3379 ), .Z(
        \SUBBYTES[9].a/w3383 ) );
  AND U2086 ( .A(\SUBBYTES[9].a/w3380 ), .B(\SUBBYTES[9].a/w3381 ), .Z(
        \SUBBYTES[9].a/w3382 ) );
  AND U2087 ( .A(\SUBBYTES[9].a/w3269 ), .B(n1211), .Z(\SUBBYTES[9].a/w3368 )
         );
  XOR U2088 ( .A(\SUBBYTES[9].a/w3337 ), .B(n1100), .Z(n1211) );
  AND U2089 ( .A(\SUBBYTES[9].a/w3270 ), .B(n1212), .Z(\SUBBYTES[9].a/w3366 )
         );
  XOR U2090 ( .A(n16103), .B(\SUBBYTES[9].a/w3337 ), .Z(n1212) );
  AND U2091 ( .A(n1217), .B(n1213), .Z(\SUBBYTES[9].a/w3365 ) );
  XOR U2092 ( .A(n1100), .B(n16103), .Z(n1213) );
  ANDN U2093 ( .A(\SUBBYTES[9].a/w3271 ), .B(n1214), .Z(\SUBBYTES[9].a/w3361 )
         );
  XNOR U2094 ( .A(\SUBBYTES[9].a/w3330 ), .B(\SUBBYTES[9].a/w3333 ), .Z(n1214)
         );
  AND U2095 ( .A(\SUBBYTES[9].a/w3272 ), .B(n1215), .Z(\SUBBYTES[9].a/w3359 )
         );
  XNOR U2096 ( .A(n1218), .B(\SUBBYTES[9].a/w3330 ), .Z(n1215) );
  AND U2097 ( .A(\SUBBYTES[9].a/w3357 ), .B(n1219), .Z(\SUBBYTES[9].a/w3358 )
         );
  XOR U2098 ( .A(n1220), .B(n1218), .Z(n1219) );
  IV U2099 ( .A(n16102), .Z(n1218) );
  AND U2100 ( .A(n1221), .B(\SUBBYTES[9].a/w3376 ), .Z(\SUBBYTES[9].a/w3353 )
         );
  ANDN U2101 ( .A(\SUBBYTES[9].a/w3377 ), .B(n1222), .Z(\SUBBYTES[9].a/w3351 )
         );
  AND U2102 ( .A(n1223), .B(\SUBBYTES[9].a/w3380 ), .Z(\SUBBYTES[9].a/w3350 )
         );
  AND U2103 ( .A(\SUBBYTES[9].a/w3336 ), .B(\SUBBYTES[9].a/w3335 ), .Z(
        \SUBBYTES[9].a/w3337 ) );
  IV U2104 ( .A(n1220), .Z(\SUBBYTES[9].a/w3333 ) );
  NAND U2105 ( .A(\SUBBYTES[9].a/w3312 ), .B(\SUBBYTES[9].a/w3327 ), .Z(n1220)
         );
  AND U2106 ( .A(\SUBBYTES[9].a/w3329 ), .B(\SUBBYTES[9].a/w3335 ), .Z(
        \SUBBYTES[9].a/w3330 ) );
  AND U2107 ( .A(\SUBBYTES[9].a/w3314 ), .B(\SUBBYTES[9].a/w3312 ), .Z(
        \SUBBYTES[9].a/w3324 ) );
  AND U2108 ( .A(\SUBBYTES[9].a/w3315 ), .B(\SUBBYTES[9].a/w3313 ), .Z(
        \SUBBYTES[9].a/w3322 ) );
  AND U2109 ( .A(\SUBBYTES[9].a/w3329 ), .B(\SUBBYTES[9].a/w3336 ), .Z(
        \SUBBYTES[9].a/w3321 ) );
  AND U2110 ( .A(\SUBBYTES[9].a/w3269 ), .B(\SUBBYTES[9].a/w3265 ), .Z(
        \SUBBYTES[9].a/w3306 ) );
  AND U2111 ( .A(\SUBBYTES[9].a/w3270 ), .B(\SUBBYTES[9].a/w3266 ), .Z(
        \SUBBYTES[9].a/w3304 ) );
  AND U2112 ( .A(\SUBBYTES[9].a/w3396 ), .B(n1217), .Z(\SUBBYTES[9].a/w3303 )
         );
  XNOR U2113 ( .A(\w1[9][1] ), .B(n1224), .Z(n1217) );
  XOR U2114 ( .A(g_input[1153]), .B(\w0[9][1] ), .Z(\w1[9][1] ) );
  AND U2115 ( .A(\w1[9][0] ), .B(\SUBBYTES[9].a/w3271 ), .Z(
        \SUBBYTES[9].a/w3299 ) );
  XOR U2116 ( .A(g_input[1152]), .B(\w0[9][0] ), .Z(\w1[9][0] ) );
  AND U2117 ( .A(\SUBBYTES[9].a/w3272 ), .B(\SUBBYTES[9].a/w3268 ), .Z(
        \SUBBYTES[9].a/w3297 ) );
  AND U2118 ( .A(\SUBBYTES[9].a/w3357 ), .B(\SUBBYTES[9].a/w3389 ), .Z(
        \SUBBYTES[9].a/w3296 ) );
  AND U2119 ( .A(\SUBBYTES[9].a/w3378 ), .B(n1221), .Z(\SUBBYTES[9].a/w3291 )
         );
  XOR U2120 ( .A(\w1[9][4] ), .B(\w1[9][7] ), .Z(n1221) );
  ANDN U2121 ( .A(\SUBBYTES[9].a/w3379 ), .B(n1222), .Z(\SUBBYTES[9].a/w3289 )
         );
  XNOR U2122 ( .A(\w1[9][2] ), .B(\w1[9][7] ), .Z(n1222) );
  IV U2123 ( .A(n1224), .Z(\w1[9][7] ) );
  XNOR U2124 ( .A(g_input[1159]), .B(\w0[9][7] ), .Z(n1224) );
  AND U2125 ( .A(\SUBBYTES[9].a/w3381 ), .B(n1223), .Z(\SUBBYTES[9].a/w3288 )
         );
  XOR U2126 ( .A(\w1[9][2] ), .B(\w1[9][4] ), .Z(n1223) );
  XOR U2127 ( .A(g_input[1156]), .B(\w0[9][4] ), .Z(\w1[9][4] ) );
  XOR U2128 ( .A(g_input[1154]), .B(\w0[9][2] ), .Z(\w1[9][2] ) );
  AND U2129 ( .A(n1225), .B(\SUBBYTES[9].a/w3058 ), .Z(\SUBBYTES[9].a/w3193 )
         );
  AND U2130 ( .A(n1226), .B(\SUBBYTES[9].a/w3059 ), .Z(\SUBBYTES[9].a/w3191 )
         );
  AND U2131 ( .A(\SUBBYTES[9].a/w3189 ), .B(n1227), .Z(\SUBBYTES[9].a/w3190 )
         );
  ANDN U2132 ( .A(\w1[9][8] ), .B(n1228), .Z(\SUBBYTES[9].a/w3186 ) );
  AND U2133 ( .A(n1229), .B(\SUBBYTES[9].a/w3061 ), .Z(\SUBBYTES[9].a/w3184 )
         );
  AND U2134 ( .A(\SUBBYTES[9].a/w3182 ), .B(n1230), .Z(\SUBBYTES[9].a/w3183 )
         );
  XOR U2135 ( .A(\SUBBYTES[9].a/w3126 ), .B(n16100), .Z(n1230) );
  AND U2136 ( .A(\SUBBYTES[9].a/w3169 ), .B(\SUBBYTES[9].a/w3171 ), .Z(
        \SUBBYTES[9].a/w3178 ) );
  AND U2137 ( .A(\SUBBYTES[9].a/w3170 ), .B(\SUBBYTES[9].a/w3172 ), .Z(
        \SUBBYTES[9].a/w3176 ) );
  AND U2138 ( .A(\SUBBYTES[9].a/w3173 ), .B(\SUBBYTES[9].a/w3174 ), .Z(
        \SUBBYTES[9].a/w3175 ) );
  AND U2139 ( .A(\SUBBYTES[9].a/w3062 ), .B(n1225), .Z(\SUBBYTES[9].a/w3161 )
         );
  XOR U2140 ( .A(\SUBBYTES[9].a/w3130 ), .B(n1099), .Z(n1225) );
  AND U2141 ( .A(\SUBBYTES[9].a/w3063 ), .B(n1226), .Z(\SUBBYTES[9].a/w3159 )
         );
  XOR U2142 ( .A(n16101), .B(\SUBBYTES[9].a/w3130 ), .Z(n1226) );
  AND U2143 ( .A(n1231), .B(n1227), .Z(\SUBBYTES[9].a/w3158 ) );
  XOR U2144 ( .A(n1099), .B(n16101), .Z(n1227) );
  ANDN U2145 ( .A(\SUBBYTES[9].a/w3064 ), .B(n1228), .Z(\SUBBYTES[9].a/w3154 )
         );
  XNOR U2146 ( .A(\SUBBYTES[9].a/w3123 ), .B(\SUBBYTES[9].a/w3126 ), .Z(n1228)
         );
  AND U2147 ( .A(\SUBBYTES[9].a/w3065 ), .B(n1229), .Z(\SUBBYTES[9].a/w3152 )
         );
  XNOR U2148 ( .A(n1232), .B(\SUBBYTES[9].a/w3123 ), .Z(n1229) );
  AND U2149 ( .A(\SUBBYTES[9].a/w3150 ), .B(n1233), .Z(\SUBBYTES[9].a/w3151 )
         );
  XOR U2150 ( .A(n1234), .B(n1232), .Z(n1233) );
  IV U2151 ( .A(n16100), .Z(n1232) );
  AND U2152 ( .A(n1235), .B(\SUBBYTES[9].a/w3169 ), .Z(\SUBBYTES[9].a/w3146 )
         );
  ANDN U2153 ( .A(\SUBBYTES[9].a/w3170 ), .B(n1236), .Z(\SUBBYTES[9].a/w3144 )
         );
  AND U2154 ( .A(n1237), .B(\SUBBYTES[9].a/w3173 ), .Z(\SUBBYTES[9].a/w3143 )
         );
  AND U2155 ( .A(\SUBBYTES[9].a/w3129 ), .B(\SUBBYTES[9].a/w3128 ), .Z(
        \SUBBYTES[9].a/w3130 ) );
  IV U2156 ( .A(n1234), .Z(\SUBBYTES[9].a/w3126 ) );
  NAND U2157 ( .A(\SUBBYTES[9].a/w3105 ), .B(\SUBBYTES[9].a/w3120 ), .Z(n1234)
         );
  AND U2158 ( .A(\SUBBYTES[9].a/w3122 ), .B(\SUBBYTES[9].a/w3128 ), .Z(
        \SUBBYTES[9].a/w3123 ) );
  AND U2159 ( .A(\SUBBYTES[9].a/w3107 ), .B(\SUBBYTES[9].a/w3105 ), .Z(
        \SUBBYTES[9].a/w3117 ) );
  AND U2160 ( .A(\SUBBYTES[9].a/w3108 ), .B(\SUBBYTES[9].a/w3106 ), .Z(
        \SUBBYTES[9].a/w3115 ) );
  AND U2161 ( .A(\SUBBYTES[9].a/w3122 ), .B(\SUBBYTES[9].a/w3129 ), .Z(
        \SUBBYTES[9].a/w3114 ) );
  AND U2162 ( .A(\SUBBYTES[9].a/w3062 ), .B(\SUBBYTES[9].a/w3058 ), .Z(
        \SUBBYTES[9].a/w3099 ) );
  AND U2163 ( .A(\SUBBYTES[9].a/w3063 ), .B(\SUBBYTES[9].a/w3059 ), .Z(
        \SUBBYTES[9].a/w3097 ) );
  AND U2164 ( .A(\SUBBYTES[9].a/w3189 ), .B(n1231), .Z(\SUBBYTES[9].a/w3096 )
         );
  XNOR U2165 ( .A(n1238), .B(\w1[9][9] ), .Z(n1231) );
  XOR U2166 ( .A(g_input[1161]), .B(\w0[9][9] ), .Z(\w1[9][9] ) );
  AND U2167 ( .A(\w1[9][8] ), .B(\SUBBYTES[9].a/w3064 ), .Z(
        \SUBBYTES[9].a/w3092 ) );
  XOR U2168 ( .A(g_input[1160]), .B(\w0[9][8] ), .Z(\w1[9][8] ) );
  AND U2169 ( .A(\SUBBYTES[9].a/w3065 ), .B(\SUBBYTES[9].a/w3061 ), .Z(
        \SUBBYTES[9].a/w3090 ) );
  AND U2170 ( .A(\SUBBYTES[9].a/w3150 ), .B(\SUBBYTES[9].a/w3182 ), .Z(
        \SUBBYTES[9].a/w3089 ) );
  AND U2171 ( .A(\SUBBYTES[9].a/w3171 ), .B(n1235), .Z(\SUBBYTES[9].a/w3084 )
         );
  XOR U2172 ( .A(\w1[9][12] ), .B(\w1[9][15] ), .Z(n1235) );
  ANDN U2173 ( .A(\SUBBYTES[9].a/w3172 ), .B(n1236), .Z(\SUBBYTES[9].a/w3082 )
         );
  XNOR U2174 ( .A(\w1[9][10] ), .B(\w1[9][15] ), .Z(n1236) );
  IV U2175 ( .A(n1238), .Z(\w1[9][15] ) );
  XNOR U2176 ( .A(g_input[1167]), .B(\w0[9][15] ), .Z(n1238) );
  AND U2177 ( .A(\SUBBYTES[9].a/w3174 ), .B(n1237), .Z(\SUBBYTES[9].a/w3081 )
         );
  XOR U2178 ( .A(\w1[9][10] ), .B(\w1[9][12] ), .Z(n1237) );
  XOR U2179 ( .A(g_input[1164]), .B(\w0[9][12] ), .Z(\w1[9][12] ) );
  XOR U2180 ( .A(g_input[1162]), .B(\w0[9][10] ), .Z(\w1[9][10] ) );
  AND U2181 ( .A(n1239), .B(\SUBBYTES[9].a/w2851 ), .Z(\SUBBYTES[9].a/w2986 )
         );
  AND U2182 ( .A(n1240), .B(\SUBBYTES[9].a/w2852 ), .Z(\SUBBYTES[9].a/w2984 )
         );
  AND U2183 ( .A(\SUBBYTES[9].a/w2982 ), .B(n1241), .Z(\SUBBYTES[9].a/w2983 )
         );
  ANDN U2184 ( .A(\w1[9][16] ), .B(n1242), .Z(\SUBBYTES[9].a/w2979 ) );
  AND U2185 ( .A(n1243), .B(\SUBBYTES[9].a/w2854 ), .Z(\SUBBYTES[9].a/w2977 )
         );
  AND U2186 ( .A(\SUBBYTES[9].a/w2975 ), .B(n1244), .Z(\SUBBYTES[9].a/w2976 )
         );
  XOR U2187 ( .A(\SUBBYTES[9].a/w2919 ), .B(n16098), .Z(n1244) );
  AND U2188 ( .A(\SUBBYTES[9].a/w2962 ), .B(\SUBBYTES[9].a/w2964 ), .Z(
        \SUBBYTES[9].a/w2971 ) );
  AND U2189 ( .A(\SUBBYTES[9].a/w2963 ), .B(\SUBBYTES[9].a/w2965 ), .Z(
        \SUBBYTES[9].a/w2969 ) );
  AND U2190 ( .A(\SUBBYTES[9].a/w2966 ), .B(\SUBBYTES[9].a/w2967 ), .Z(
        \SUBBYTES[9].a/w2968 ) );
  AND U2191 ( .A(\SUBBYTES[9].a/w2855 ), .B(n1239), .Z(\SUBBYTES[9].a/w2954 )
         );
  XOR U2192 ( .A(\SUBBYTES[9].a/w2923 ), .B(n1098), .Z(n1239) );
  AND U2193 ( .A(\SUBBYTES[9].a/w2856 ), .B(n1240), .Z(\SUBBYTES[9].a/w2952 )
         );
  XOR U2194 ( .A(n16099), .B(\SUBBYTES[9].a/w2923 ), .Z(n1240) );
  AND U2195 ( .A(n1245), .B(n1241), .Z(\SUBBYTES[9].a/w2951 ) );
  XOR U2196 ( .A(n1098), .B(n16099), .Z(n1241) );
  AND U2197 ( .A(n1246), .B(\SUBBYTES[9].a/w160 ), .Z(\SUBBYTES[9].a/w295 ) );
  ANDN U2198 ( .A(\SUBBYTES[9].a/w2857 ), .B(n1242), .Z(\SUBBYTES[9].a/w2947 )
         );
  XNOR U2199 ( .A(\SUBBYTES[9].a/w2916 ), .B(\SUBBYTES[9].a/w2919 ), .Z(n1242)
         );
  AND U2200 ( .A(\SUBBYTES[9].a/w2858 ), .B(n1243), .Z(\SUBBYTES[9].a/w2945 )
         );
  XNOR U2201 ( .A(n1247), .B(\SUBBYTES[9].a/w2916 ), .Z(n1243) );
  AND U2202 ( .A(\SUBBYTES[9].a/w2943 ), .B(n1248), .Z(\SUBBYTES[9].a/w2944 )
         );
  XOR U2203 ( .A(n1249), .B(n1247), .Z(n1248) );
  IV U2204 ( .A(n16098), .Z(n1247) );
  AND U2205 ( .A(n1250), .B(\SUBBYTES[9].a/w2962 ), .Z(\SUBBYTES[9].a/w2939 )
         );
  ANDN U2206 ( .A(\SUBBYTES[9].a/w2963 ), .B(n1251), .Z(\SUBBYTES[9].a/w2937 )
         );
  AND U2207 ( .A(n1252), .B(\SUBBYTES[9].a/w2966 ), .Z(\SUBBYTES[9].a/w2936 )
         );
  AND U2208 ( .A(n1253), .B(\SUBBYTES[9].a/w161 ), .Z(\SUBBYTES[9].a/w293 ) );
  AND U2209 ( .A(\SUBBYTES[9].a/w2922 ), .B(\SUBBYTES[9].a/w2921 ), .Z(
        \SUBBYTES[9].a/w2923 ) );
  AND U2210 ( .A(\SUBBYTES[9].a/w291 ), .B(n1254), .Z(\SUBBYTES[9].a/w292 ) );
  IV U2211 ( .A(n1249), .Z(\SUBBYTES[9].a/w2919 ) );
  NAND U2212 ( .A(\SUBBYTES[9].a/w2898 ), .B(\SUBBYTES[9].a/w2913 ), .Z(n1249)
         );
  AND U2213 ( .A(\SUBBYTES[9].a/w2915 ), .B(\SUBBYTES[9].a/w2921 ), .Z(
        \SUBBYTES[9].a/w2916 ) );
  AND U2214 ( .A(\SUBBYTES[9].a/w2900 ), .B(\SUBBYTES[9].a/w2898 ), .Z(
        \SUBBYTES[9].a/w2910 ) );
  AND U2215 ( .A(\SUBBYTES[9].a/w2901 ), .B(\SUBBYTES[9].a/w2899 ), .Z(
        \SUBBYTES[9].a/w2908 ) );
  AND U2216 ( .A(\SUBBYTES[9].a/w2915 ), .B(\SUBBYTES[9].a/w2922 ), .Z(
        \SUBBYTES[9].a/w2907 ) );
  AND U2217 ( .A(\SUBBYTES[9].a/w2855 ), .B(\SUBBYTES[9].a/w2851 ), .Z(
        \SUBBYTES[9].a/w2892 ) );
  AND U2218 ( .A(\SUBBYTES[9].a/w2856 ), .B(\SUBBYTES[9].a/w2852 ), .Z(
        \SUBBYTES[9].a/w2890 ) );
  AND U2219 ( .A(\SUBBYTES[9].a/w2982 ), .B(n1245), .Z(\SUBBYTES[9].a/w2889 )
         );
  XNOR U2220 ( .A(\w1[9][17] ), .B(n1255), .Z(n1245) );
  XOR U2221 ( .A(g_input[1169]), .B(\w0[9][17] ), .Z(\w1[9][17] ) );
  AND U2222 ( .A(\w1[9][16] ), .B(\SUBBYTES[9].a/w2857 ), .Z(
        \SUBBYTES[9].a/w2885 ) );
  XOR U2223 ( .A(g_input[1168]), .B(\w0[9][16] ), .Z(\w1[9][16] ) );
  AND U2224 ( .A(\SUBBYTES[9].a/w2858 ), .B(\SUBBYTES[9].a/w2854 ), .Z(
        \SUBBYTES[9].a/w2883 ) );
  AND U2225 ( .A(\SUBBYTES[9].a/w2943 ), .B(\SUBBYTES[9].a/w2975 ), .Z(
        \SUBBYTES[9].a/w2882 ) );
  ANDN U2226 ( .A(\w1[9][120] ), .B(n1256), .Z(\SUBBYTES[9].a/w288 ) );
  AND U2227 ( .A(\SUBBYTES[9].a/w2964 ), .B(n1250), .Z(\SUBBYTES[9].a/w2877 )
         );
  XOR U2228 ( .A(\w1[9][20] ), .B(\w1[9][23] ), .Z(n1250) );
  ANDN U2229 ( .A(\SUBBYTES[9].a/w2965 ), .B(n1251), .Z(\SUBBYTES[9].a/w2875 )
         );
  XNOR U2230 ( .A(\w1[9][18] ), .B(\w1[9][23] ), .Z(n1251) );
  IV U2231 ( .A(n1255), .Z(\w1[9][23] ) );
  XNOR U2232 ( .A(g_input[1175]), .B(\w0[9][23] ), .Z(n1255) );
  AND U2233 ( .A(\SUBBYTES[9].a/w2967 ), .B(n1252), .Z(\SUBBYTES[9].a/w2874 )
         );
  XOR U2234 ( .A(\w1[9][18] ), .B(\w1[9][20] ), .Z(n1252) );
  XOR U2235 ( .A(g_input[1172]), .B(\w0[9][20] ), .Z(\w1[9][20] ) );
  XOR U2236 ( .A(g_input[1170]), .B(\w0[9][18] ), .Z(\w1[9][18] ) );
  AND U2237 ( .A(n1257), .B(\SUBBYTES[9].a/w163 ), .Z(\SUBBYTES[9].a/w286 ) );
  AND U2238 ( .A(\SUBBYTES[9].a/w284 ), .B(n1258), .Z(\SUBBYTES[9].a/w285 ) );
  XOR U2239 ( .A(\SUBBYTES[9].a/w228 ), .B(n16072), .Z(n1258) );
  AND U2240 ( .A(\SUBBYTES[9].a/w271 ), .B(\SUBBYTES[9].a/w273 ), .Z(
        \SUBBYTES[9].a/w280 ) );
  AND U2241 ( .A(\SUBBYTES[9].a/w272 ), .B(\SUBBYTES[9].a/w274 ), .Z(
        \SUBBYTES[9].a/w278 ) );
  AND U2242 ( .A(n1259), .B(\SUBBYTES[9].a/w2644 ), .Z(\SUBBYTES[9].a/w2779 )
         );
  AND U2243 ( .A(n1260), .B(\SUBBYTES[9].a/w2645 ), .Z(\SUBBYTES[9].a/w2777 )
         );
  AND U2244 ( .A(\SUBBYTES[9].a/w2775 ), .B(n1261), .Z(\SUBBYTES[9].a/w2776 )
         );
  ANDN U2245 ( .A(\w1[9][24] ), .B(n1262), .Z(\SUBBYTES[9].a/w2772 ) );
  AND U2246 ( .A(n1263), .B(\SUBBYTES[9].a/w2647 ), .Z(\SUBBYTES[9].a/w2770 )
         );
  AND U2247 ( .A(\SUBBYTES[9].a/w275 ), .B(\SUBBYTES[9].a/w276 ), .Z(
        \SUBBYTES[9].a/w277 ) );
  AND U2248 ( .A(\SUBBYTES[9].a/w2768 ), .B(n1264), .Z(\SUBBYTES[9].a/w2769 )
         );
  XOR U2249 ( .A(\SUBBYTES[9].a/w2712 ), .B(n16096), .Z(n1264) );
  AND U2250 ( .A(\SUBBYTES[9].a/w2755 ), .B(\SUBBYTES[9].a/w2757 ), .Z(
        \SUBBYTES[9].a/w2764 ) );
  AND U2251 ( .A(\SUBBYTES[9].a/w2756 ), .B(\SUBBYTES[9].a/w2758 ), .Z(
        \SUBBYTES[9].a/w2762 ) );
  AND U2252 ( .A(\SUBBYTES[9].a/w2759 ), .B(\SUBBYTES[9].a/w2760 ), .Z(
        \SUBBYTES[9].a/w2761 ) );
  AND U2253 ( .A(\SUBBYTES[9].a/w2648 ), .B(n1259), .Z(\SUBBYTES[9].a/w2747 )
         );
  XOR U2254 ( .A(\SUBBYTES[9].a/w2716 ), .B(n1097), .Z(n1259) );
  AND U2255 ( .A(\SUBBYTES[9].a/w2649 ), .B(n1260), .Z(\SUBBYTES[9].a/w2745 )
         );
  XOR U2256 ( .A(n16097), .B(\SUBBYTES[9].a/w2716 ), .Z(n1260) );
  AND U2257 ( .A(n1265), .B(n1261), .Z(\SUBBYTES[9].a/w2744 ) );
  XOR U2258 ( .A(n1097), .B(n16097), .Z(n1261) );
  ANDN U2259 ( .A(\SUBBYTES[9].a/w2650 ), .B(n1262), .Z(\SUBBYTES[9].a/w2740 )
         );
  XNOR U2260 ( .A(\SUBBYTES[9].a/w2709 ), .B(\SUBBYTES[9].a/w2712 ), .Z(n1262)
         );
  AND U2261 ( .A(\SUBBYTES[9].a/w2651 ), .B(n1263), .Z(\SUBBYTES[9].a/w2738 )
         );
  XNOR U2262 ( .A(n1266), .B(\SUBBYTES[9].a/w2709 ), .Z(n1263) );
  AND U2263 ( .A(\SUBBYTES[9].a/w2736 ), .B(n1267), .Z(\SUBBYTES[9].a/w2737 )
         );
  XOR U2264 ( .A(n1268), .B(n1266), .Z(n1267) );
  IV U2265 ( .A(n16096), .Z(n1266) );
  AND U2266 ( .A(n1269), .B(\SUBBYTES[9].a/w2755 ), .Z(\SUBBYTES[9].a/w2732 )
         );
  ANDN U2267 ( .A(\SUBBYTES[9].a/w2756 ), .B(n1270), .Z(\SUBBYTES[9].a/w2730 )
         );
  AND U2268 ( .A(n1271), .B(\SUBBYTES[9].a/w2759 ), .Z(\SUBBYTES[9].a/w2729 )
         );
  AND U2269 ( .A(\SUBBYTES[9].a/w2715 ), .B(\SUBBYTES[9].a/w2714 ), .Z(
        \SUBBYTES[9].a/w2716 ) );
  IV U2270 ( .A(n1268), .Z(\SUBBYTES[9].a/w2712 ) );
  NAND U2271 ( .A(\SUBBYTES[9].a/w2691 ), .B(\SUBBYTES[9].a/w2706 ), .Z(n1268)
         );
  AND U2272 ( .A(\SUBBYTES[9].a/w2708 ), .B(\SUBBYTES[9].a/w2714 ), .Z(
        \SUBBYTES[9].a/w2709 ) );
  AND U2273 ( .A(\SUBBYTES[9].a/w2693 ), .B(\SUBBYTES[9].a/w2691 ), .Z(
        \SUBBYTES[9].a/w2703 ) );
  AND U2274 ( .A(\SUBBYTES[9].a/w2694 ), .B(\SUBBYTES[9].a/w2692 ), .Z(
        \SUBBYTES[9].a/w2701 ) );
  AND U2275 ( .A(\SUBBYTES[9].a/w2708 ), .B(\SUBBYTES[9].a/w2715 ), .Z(
        \SUBBYTES[9].a/w2700 ) );
  AND U2276 ( .A(\SUBBYTES[9].a/w2648 ), .B(\SUBBYTES[9].a/w2644 ), .Z(
        \SUBBYTES[9].a/w2685 ) );
  AND U2277 ( .A(\SUBBYTES[9].a/w2649 ), .B(\SUBBYTES[9].a/w2645 ), .Z(
        \SUBBYTES[9].a/w2683 ) );
  AND U2278 ( .A(\SUBBYTES[9].a/w2775 ), .B(n1265), .Z(\SUBBYTES[9].a/w2682 )
         );
  XNOR U2279 ( .A(\w1[9][25] ), .B(n1272), .Z(n1265) );
  XOR U2280 ( .A(g_input[1177]), .B(\w0[9][25] ), .Z(\w1[9][25] ) );
  AND U2281 ( .A(\w1[9][24] ), .B(\SUBBYTES[9].a/w2650 ), .Z(
        \SUBBYTES[9].a/w2678 ) );
  XOR U2282 ( .A(g_input[1176]), .B(\w0[9][24] ), .Z(\w1[9][24] ) );
  AND U2283 ( .A(\SUBBYTES[9].a/w2651 ), .B(\SUBBYTES[9].a/w2647 ), .Z(
        \SUBBYTES[9].a/w2676 ) );
  AND U2284 ( .A(\SUBBYTES[9].a/w2736 ), .B(\SUBBYTES[9].a/w2768 ), .Z(
        \SUBBYTES[9].a/w2675 ) );
  AND U2285 ( .A(\SUBBYTES[9].a/w2757 ), .B(n1269), .Z(\SUBBYTES[9].a/w2670 )
         );
  XOR U2286 ( .A(\w1[9][28] ), .B(\w1[9][31] ), .Z(n1269) );
  ANDN U2287 ( .A(\SUBBYTES[9].a/w2758 ), .B(n1270), .Z(\SUBBYTES[9].a/w2668 )
         );
  XNOR U2288 ( .A(\w1[9][26] ), .B(\w1[9][31] ), .Z(n1270) );
  IV U2289 ( .A(n1272), .Z(\w1[9][31] ) );
  XNOR U2290 ( .A(g_input[1183]), .B(\w0[9][31] ), .Z(n1272) );
  AND U2291 ( .A(\SUBBYTES[9].a/w2760 ), .B(n1271), .Z(\SUBBYTES[9].a/w2667 )
         );
  XOR U2292 ( .A(\w1[9][26] ), .B(\w1[9][28] ), .Z(n1271) );
  XOR U2293 ( .A(g_input[1180]), .B(\w0[9][28] ), .Z(\w1[9][28] ) );
  XOR U2294 ( .A(g_input[1178]), .B(\w0[9][26] ), .Z(\w1[9][26] ) );
  AND U2295 ( .A(\SUBBYTES[9].a/w164 ), .B(n1246), .Z(\SUBBYTES[9].a/w263 ) );
  XOR U2296 ( .A(\SUBBYTES[9].a/w232 ), .B(n1085), .Z(n1246) );
  AND U2297 ( .A(\SUBBYTES[9].a/w165 ), .B(n1253), .Z(\SUBBYTES[9].a/w261 ) );
  XOR U2298 ( .A(n16073), .B(\SUBBYTES[9].a/w232 ), .Z(n1253) );
  AND U2299 ( .A(n1273), .B(n1254), .Z(\SUBBYTES[9].a/w260 ) );
  XOR U2300 ( .A(n1085), .B(n16073), .Z(n1254) );
  AND U2301 ( .A(n1274), .B(\SUBBYTES[9].a/w2437 ), .Z(\SUBBYTES[9].a/w2572 )
         );
  AND U2302 ( .A(n1275), .B(\SUBBYTES[9].a/w2438 ), .Z(\SUBBYTES[9].a/w2570 )
         );
  AND U2303 ( .A(\SUBBYTES[9].a/w2568 ), .B(n1276), .Z(\SUBBYTES[9].a/w2569 )
         );
  ANDN U2304 ( .A(\w1[9][32] ), .B(n1277), .Z(\SUBBYTES[9].a/w2565 ) );
  AND U2305 ( .A(n1278), .B(\SUBBYTES[9].a/w2440 ), .Z(\SUBBYTES[9].a/w2563 )
         );
  AND U2306 ( .A(\SUBBYTES[9].a/w2561 ), .B(n1279), .Z(\SUBBYTES[9].a/w2562 )
         );
  XOR U2307 ( .A(\SUBBYTES[9].a/w2505 ), .B(n16094), .Z(n1279) );
  ANDN U2308 ( .A(\SUBBYTES[9].a/w166 ), .B(n1256), .Z(\SUBBYTES[9].a/w256 )
         );
  XNOR U2309 ( .A(\SUBBYTES[9].a/w225 ), .B(\SUBBYTES[9].a/w228 ), .Z(n1256)
         );
  AND U2310 ( .A(\SUBBYTES[9].a/w2548 ), .B(\SUBBYTES[9].a/w2550 ), .Z(
        \SUBBYTES[9].a/w2557 ) );
  AND U2311 ( .A(\SUBBYTES[9].a/w2549 ), .B(\SUBBYTES[9].a/w2551 ), .Z(
        \SUBBYTES[9].a/w2555 ) );
  AND U2312 ( .A(\SUBBYTES[9].a/w2552 ), .B(\SUBBYTES[9].a/w2553 ), .Z(
        \SUBBYTES[9].a/w2554 ) );
  AND U2313 ( .A(\SUBBYTES[9].a/w2441 ), .B(n1274), .Z(\SUBBYTES[9].a/w2540 )
         );
  XOR U2314 ( .A(\SUBBYTES[9].a/w2509 ), .B(n1096), .Z(n1274) );
  AND U2315 ( .A(\SUBBYTES[9].a/w167 ), .B(n1257), .Z(\SUBBYTES[9].a/w254 ) );
  XNOR U2316 ( .A(n1280), .B(\SUBBYTES[9].a/w225 ), .Z(n1257) );
  AND U2317 ( .A(\SUBBYTES[9].a/w2442 ), .B(n1275), .Z(\SUBBYTES[9].a/w2538 )
         );
  XOR U2318 ( .A(n16095), .B(\SUBBYTES[9].a/w2509 ), .Z(n1275) );
  AND U2319 ( .A(n1281), .B(n1276), .Z(\SUBBYTES[9].a/w2537 ) );
  XOR U2320 ( .A(n1096), .B(n16095), .Z(n1276) );
  ANDN U2321 ( .A(\SUBBYTES[9].a/w2443 ), .B(n1277), .Z(\SUBBYTES[9].a/w2533 )
         );
  XNOR U2322 ( .A(\SUBBYTES[9].a/w2502 ), .B(\SUBBYTES[9].a/w2505 ), .Z(n1277)
         );
  AND U2323 ( .A(\SUBBYTES[9].a/w2444 ), .B(n1278), .Z(\SUBBYTES[9].a/w2531 )
         );
  XNOR U2324 ( .A(n1282), .B(\SUBBYTES[9].a/w2502 ), .Z(n1278) );
  AND U2325 ( .A(\SUBBYTES[9].a/w2529 ), .B(n1283), .Z(\SUBBYTES[9].a/w2530 )
         );
  XOR U2326 ( .A(n1284), .B(n1282), .Z(n1283) );
  IV U2327 ( .A(n16094), .Z(n1282) );
  AND U2328 ( .A(\SUBBYTES[9].a/w252 ), .B(n1285), .Z(\SUBBYTES[9].a/w253 ) );
  XOR U2329 ( .A(n1286), .B(n1280), .Z(n1285) );
  IV U2330 ( .A(n16072), .Z(n1280) );
  AND U2331 ( .A(n1287), .B(\SUBBYTES[9].a/w2548 ), .Z(\SUBBYTES[9].a/w2525 )
         );
  ANDN U2332 ( .A(\SUBBYTES[9].a/w2549 ), .B(n1288), .Z(\SUBBYTES[9].a/w2523 )
         );
  AND U2333 ( .A(n1289), .B(\SUBBYTES[9].a/w2552 ), .Z(\SUBBYTES[9].a/w2522 )
         );
  AND U2334 ( .A(\SUBBYTES[9].a/w2508 ), .B(\SUBBYTES[9].a/w2507 ), .Z(
        \SUBBYTES[9].a/w2509 ) );
  IV U2335 ( .A(n1284), .Z(\SUBBYTES[9].a/w2505 ) );
  NAND U2336 ( .A(\SUBBYTES[9].a/w2484 ), .B(\SUBBYTES[9].a/w2499 ), .Z(n1284)
         );
  AND U2337 ( .A(\SUBBYTES[9].a/w2501 ), .B(\SUBBYTES[9].a/w2507 ), .Z(
        \SUBBYTES[9].a/w2502 ) );
  AND U2338 ( .A(\SUBBYTES[9].a/w2486 ), .B(\SUBBYTES[9].a/w2484 ), .Z(
        \SUBBYTES[9].a/w2496 ) );
  AND U2339 ( .A(\SUBBYTES[9].a/w2487 ), .B(\SUBBYTES[9].a/w2485 ), .Z(
        \SUBBYTES[9].a/w2494 ) );
  AND U2340 ( .A(\SUBBYTES[9].a/w2501 ), .B(\SUBBYTES[9].a/w2508 ), .Z(
        \SUBBYTES[9].a/w2493 ) );
  AND U2341 ( .A(n1290), .B(\SUBBYTES[9].a/w271 ), .Z(\SUBBYTES[9].a/w248 ) );
  AND U2342 ( .A(\SUBBYTES[9].a/w2441 ), .B(\SUBBYTES[9].a/w2437 ), .Z(
        \SUBBYTES[9].a/w2478 ) );
  AND U2343 ( .A(\SUBBYTES[9].a/w2442 ), .B(\SUBBYTES[9].a/w2438 ), .Z(
        \SUBBYTES[9].a/w2476 ) );
  AND U2344 ( .A(\SUBBYTES[9].a/w2568 ), .B(n1281), .Z(\SUBBYTES[9].a/w2475 )
         );
  XNOR U2345 ( .A(\w1[9][33] ), .B(n1291), .Z(n1281) );
  XOR U2346 ( .A(g_input[1185]), .B(\w0[9][33] ), .Z(\w1[9][33] ) );
  AND U2347 ( .A(\w1[9][32] ), .B(\SUBBYTES[9].a/w2443 ), .Z(
        \SUBBYTES[9].a/w2471 ) );
  XOR U2348 ( .A(g_input[1184]), .B(\w0[9][32] ), .Z(\w1[9][32] ) );
  AND U2349 ( .A(\SUBBYTES[9].a/w2444 ), .B(\SUBBYTES[9].a/w2440 ), .Z(
        \SUBBYTES[9].a/w2469 ) );
  AND U2350 ( .A(\SUBBYTES[9].a/w2529 ), .B(\SUBBYTES[9].a/w2561 ), .Z(
        \SUBBYTES[9].a/w2468 ) );
  AND U2351 ( .A(\SUBBYTES[9].a/w2550 ), .B(n1287), .Z(\SUBBYTES[9].a/w2463 )
         );
  XOR U2352 ( .A(\w1[9][36] ), .B(\w1[9][39] ), .Z(n1287) );
  ANDN U2353 ( .A(\SUBBYTES[9].a/w2551 ), .B(n1288), .Z(\SUBBYTES[9].a/w2461 )
         );
  XNOR U2354 ( .A(\w1[9][34] ), .B(\w1[9][39] ), .Z(n1288) );
  IV U2355 ( .A(n1291), .Z(\w1[9][39] ) );
  XNOR U2356 ( .A(g_input[1191]), .B(\w0[9][39] ), .Z(n1291) );
  AND U2357 ( .A(\SUBBYTES[9].a/w2553 ), .B(n1289), .Z(\SUBBYTES[9].a/w2460 )
         );
  XOR U2358 ( .A(\w1[9][34] ), .B(\w1[9][36] ), .Z(n1289) );
  XOR U2359 ( .A(g_input[1188]), .B(\w0[9][36] ), .Z(\w1[9][36] ) );
  XOR U2360 ( .A(g_input[1186]), .B(\w0[9][34] ), .Z(\w1[9][34] ) );
  ANDN U2361 ( .A(\SUBBYTES[9].a/w272 ), .B(n1292), .Z(\SUBBYTES[9].a/w246 )
         );
  AND U2362 ( .A(n1293), .B(\SUBBYTES[9].a/w275 ), .Z(\SUBBYTES[9].a/w245 ) );
  AND U2363 ( .A(n1294), .B(\SUBBYTES[9].a/w2230 ), .Z(\SUBBYTES[9].a/w2365 )
         );
  AND U2364 ( .A(n1295), .B(\SUBBYTES[9].a/w2231 ), .Z(\SUBBYTES[9].a/w2363 )
         );
  AND U2365 ( .A(\SUBBYTES[9].a/w2361 ), .B(n1296), .Z(\SUBBYTES[9].a/w2362 )
         );
  ANDN U2366 ( .A(\w1[9][40] ), .B(n1297), .Z(\SUBBYTES[9].a/w2358 ) );
  AND U2367 ( .A(n1298), .B(\SUBBYTES[9].a/w2233 ), .Z(\SUBBYTES[9].a/w2356 )
         );
  AND U2368 ( .A(\SUBBYTES[9].a/w2354 ), .B(n1299), .Z(\SUBBYTES[9].a/w2355 )
         );
  XOR U2369 ( .A(\SUBBYTES[9].a/w2298 ), .B(n16092), .Z(n1299) );
  AND U2370 ( .A(\SUBBYTES[9].a/w2341 ), .B(\SUBBYTES[9].a/w2343 ), .Z(
        \SUBBYTES[9].a/w2350 ) );
  AND U2371 ( .A(\SUBBYTES[9].a/w2342 ), .B(\SUBBYTES[9].a/w2344 ), .Z(
        \SUBBYTES[9].a/w2348 ) );
  AND U2372 ( .A(\SUBBYTES[9].a/w2345 ), .B(\SUBBYTES[9].a/w2346 ), .Z(
        \SUBBYTES[9].a/w2347 ) );
  AND U2373 ( .A(\SUBBYTES[9].a/w2234 ), .B(n1294), .Z(\SUBBYTES[9].a/w2333 )
         );
  XOR U2374 ( .A(\SUBBYTES[9].a/w2302 ), .B(n1095), .Z(n1294) );
  AND U2375 ( .A(\SUBBYTES[9].a/w2235 ), .B(n1295), .Z(\SUBBYTES[9].a/w2331 )
         );
  XOR U2376 ( .A(n16093), .B(\SUBBYTES[9].a/w2302 ), .Z(n1295) );
  AND U2377 ( .A(n1300), .B(n1296), .Z(\SUBBYTES[9].a/w2330 ) );
  XOR U2378 ( .A(n1095), .B(n16093), .Z(n1296) );
  ANDN U2379 ( .A(\SUBBYTES[9].a/w2236 ), .B(n1297), .Z(\SUBBYTES[9].a/w2326 )
         );
  XNOR U2380 ( .A(\SUBBYTES[9].a/w2295 ), .B(\SUBBYTES[9].a/w2298 ), .Z(n1297)
         );
  AND U2381 ( .A(\SUBBYTES[9].a/w2237 ), .B(n1298), .Z(\SUBBYTES[9].a/w2324 )
         );
  XNOR U2382 ( .A(n1301), .B(\SUBBYTES[9].a/w2295 ), .Z(n1298) );
  AND U2383 ( .A(\SUBBYTES[9].a/w2322 ), .B(n1302), .Z(\SUBBYTES[9].a/w2323 )
         );
  XOR U2384 ( .A(n1303), .B(n1301), .Z(n1302) );
  IV U2385 ( .A(n16092), .Z(n1301) );
  AND U2386 ( .A(\SUBBYTES[9].a/w231 ), .B(\SUBBYTES[9].a/w230 ), .Z(
        \SUBBYTES[9].a/w232 ) );
  AND U2387 ( .A(n1304), .B(\SUBBYTES[9].a/w2341 ), .Z(\SUBBYTES[9].a/w2318 )
         );
  ANDN U2388 ( .A(\SUBBYTES[9].a/w2342 ), .B(n1305), .Z(\SUBBYTES[9].a/w2316 )
         );
  AND U2389 ( .A(n1306), .B(\SUBBYTES[9].a/w2345 ), .Z(\SUBBYTES[9].a/w2315 )
         );
  AND U2390 ( .A(\SUBBYTES[9].a/w2301 ), .B(\SUBBYTES[9].a/w2300 ), .Z(
        \SUBBYTES[9].a/w2302 ) );
  IV U2391 ( .A(n1303), .Z(\SUBBYTES[9].a/w2298 ) );
  NAND U2392 ( .A(\SUBBYTES[9].a/w2277 ), .B(\SUBBYTES[9].a/w2292 ), .Z(n1303)
         );
  AND U2393 ( .A(\SUBBYTES[9].a/w2294 ), .B(\SUBBYTES[9].a/w2300 ), .Z(
        \SUBBYTES[9].a/w2295 ) );
  AND U2394 ( .A(\SUBBYTES[9].a/w2279 ), .B(\SUBBYTES[9].a/w2277 ), .Z(
        \SUBBYTES[9].a/w2289 ) );
  AND U2395 ( .A(\SUBBYTES[9].a/w2280 ), .B(\SUBBYTES[9].a/w2278 ), .Z(
        \SUBBYTES[9].a/w2287 ) );
  AND U2396 ( .A(\SUBBYTES[9].a/w2294 ), .B(\SUBBYTES[9].a/w2301 ), .Z(
        \SUBBYTES[9].a/w2286 ) );
  IV U2397 ( .A(n1286), .Z(\SUBBYTES[9].a/w228 ) );
  NAND U2398 ( .A(\SUBBYTES[9].a/w207 ), .B(\SUBBYTES[9].a/w222 ), .Z(n1286)
         );
  AND U2399 ( .A(\SUBBYTES[9].a/w2234 ), .B(\SUBBYTES[9].a/w2230 ), .Z(
        \SUBBYTES[9].a/w2271 ) );
  AND U2400 ( .A(\SUBBYTES[9].a/w2235 ), .B(\SUBBYTES[9].a/w2231 ), .Z(
        \SUBBYTES[9].a/w2269 ) );
  AND U2401 ( .A(\SUBBYTES[9].a/w2361 ), .B(n1300), .Z(\SUBBYTES[9].a/w2268 )
         );
  XNOR U2402 ( .A(\w1[9][41] ), .B(n1307), .Z(n1300) );
  XOR U2403 ( .A(g_input[1193]), .B(\w0[9][41] ), .Z(\w1[9][41] ) );
  AND U2404 ( .A(\w1[9][40] ), .B(\SUBBYTES[9].a/w2236 ), .Z(
        \SUBBYTES[9].a/w2264 ) );
  XOR U2405 ( .A(g_input[1192]), .B(\w0[9][40] ), .Z(\w1[9][40] ) );
  AND U2406 ( .A(\SUBBYTES[9].a/w2237 ), .B(\SUBBYTES[9].a/w2233 ), .Z(
        \SUBBYTES[9].a/w2262 ) );
  AND U2407 ( .A(\SUBBYTES[9].a/w2322 ), .B(\SUBBYTES[9].a/w2354 ), .Z(
        \SUBBYTES[9].a/w2261 ) );
  AND U2408 ( .A(\SUBBYTES[9].a/w2343 ), .B(n1304), .Z(\SUBBYTES[9].a/w2256 )
         );
  XOR U2409 ( .A(\w1[9][44] ), .B(\w1[9][47] ), .Z(n1304) );
  ANDN U2410 ( .A(\SUBBYTES[9].a/w2344 ), .B(n1305), .Z(\SUBBYTES[9].a/w2254 )
         );
  XNOR U2411 ( .A(\w1[9][42] ), .B(\w1[9][47] ), .Z(n1305) );
  IV U2412 ( .A(n1307), .Z(\w1[9][47] ) );
  XNOR U2413 ( .A(g_input[1199]), .B(\w0[9][47] ), .Z(n1307) );
  AND U2414 ( .A(\SUBBYTES[9].a/w2346 ), .B(n1306), .Z(\SUBBYTES[9].a/w2253 )
         );
  XOR U2415 ( .A(\w1[9][42] ), .B(\w1[9][44] ), .Z(n1306) );
  XOR U2416 ( .A(g_input[1196]), .B(\w0[9][44] ), .Z(\w1[9][44] ) );
  XOR U2417 ( .A(g_input[1194]), .B(\w0[9][42] ), .Z(\w1[9][42] ) );
  AND U2418 ( .A(\SUBBYTES[9].a/w224 ), .B(\SUBBYTES[9].a/w230 ), .Z(
        \SUBBYTES[9].a/w225 ) );
  AND U2419 ( .A(\SUBBYTES[9].a/w209 ), .B(\SUBBYTES[9].a/w207 ), .Z(
        \SUBBYTES[9].a/w219 ) );
  AND U2420 ( .A(\SUBBYTES[9].a/w210 ), .B(\SUBBYTES[9].a/w208 ), .Z(
        \SUBBYTES[9].a/w217 ) );
  AND U2421 ( .A(\SUBBYTES[9].a/w224 ), .B(\SUBBYTES[9].a/w231 ), .Z(
        \SUBBYTES[9].a/w216 ) );
  AND U2422 ( .A(n1308), .B(\SUBBYTES[9].a/w2023 ), .Z(\SUBBYTES[9].a/w2158 )
         );
  AND U2423 ( .A(n1309), .B(\SUBBYTES[9].a/w2024 ), .Z(\SUBBYTES[9].a/w2156 )
         );
  AND U2424 ( .A(\SUBBYTES[9].a/w2154 ), .B(n1310), .Z(\SUBBYTES[9].a/w2155 )
         );
  ANDN U2425 ( .A(\w1[9][48] ), .B(n1311), .Z(\SUBBYTES[9].a/w2151 ) );
  AND U2426 ( .A(n1312), .B(\SUBBYTES[9].a/w2026 ), .Z(\SUBBYTES[9].a/w2149 )
         );
  AND U2427 ( .A(\SUBBYTES[9].a/w2147 ), .B(n1313), .Z(\SUBBYTES[9].a/w2148 )
         );
  XOR U2428 ( .A(\SUBBYTES[9].a/w2091 ), .B(n16090), .Z(n1313) );
  AND U2429 ( .A(\SUBBYTES[9].a/w2134 ), .B(\SUBBYTES[9].a/w2136 ), .Z(
        \SUBBYTES[9].a/w2143 ) );
  AND U2430 ( .A(\SUBBYTES[9].a/w2135 ), .B(\SUBBYTES[9].a/w2137 ), .Z(
        \SUBBYTES[9].a/w2141 ) );
  AND U2431 ( .A(\SUBBYTES[9].a/w2138 ), .B(\SUBBYTES[9].a/w2139 ), .Z(
        \SUBBYTES[9].a/w2140 ) );
  AND U2432 ( .A(\SUBBYTES[9].a/w2027 ), .B(n1308), .Z(\SUBBYTES[9].a/w2126 )
         );
  XOR U2433 ( .A(\SUBBYTES[9].a/w2095 ), .B(n1094), .Z(n1308) );
  AND U2434 ( .A(\SUBBYTES[9].a/w2028 ), .B(n1309), .Z(\SUBBYTES[9].a/w2124 )
         );
  XOR U2435 ( .A(n16091), .B(\SUBBYTES[9].a/w2095 ), .Z(n1309) );
  AND U2436 ( .A(n1314), .B(n1310), .Z(\SUBBYTES[9].a/w2123 ) );
  XOR U2437 ( .A(n1094), .B(n16091), .Z(n1310) );
  ANDN U2438 ( .A(\SUBBYTES[9].a/w2029 ), .B(n1311), .Z(\SUBBYTES[9].a/w2119 )
         );
  XNOR U2439 ( .A(\SUBBYTES[9].a/w2088 ), .B(\SUBBYTES[9].a/w2091 ), .Z(n1311)
         );
  AND U2440 ( .A(\SUBBYTES[9].a/w2030 ), .B(n1312), .Z(\SUBBYTES[9].a/w2117 )
         );
  XNOR U2441 ( .A(n1315), .B(\SUBBYTES[9].a/w2088 ), .Z(n1312) );
  AND U2442 ( .A(\SUBBYTES[9].a/w2115 ), .B(n1316), .Z(\SUBBYTES[9].a/w2116 )
         );
  XOR U2443 ( .A(n1317), .B(n1315), .Z(n1316) );
  IV U2444 ( .A(n16090), .Z(n1315) );
  AND U2445 ( .A(n1318), .B(\SUBBYTES[9].a/w2134 ), .Z(\SUBBYTES[9].a/w2111 )
         );
  ANDN U2446 ( .A(\SUBBYTES[9].a/w2135 ), .B(n1319), .Z(\SUBBYTES[9].a/w2109 )
         );
  AND U2447 ( .A(n1320), .B(\SUBBYTES[9].a/w2138 ), .Z(\SUBBYTES[9].a/w2108 )
         );
  AND U2448 ( .A(\SUBBYTES[9].a/w2094 ), .B(\SUBBYTES[9].a/w2093 ), .Z(
        \SUBBYTES[9].a/w2095 ) );
  IV U2449 ( .A(n1317), .Z(\SUBBYTES[9].a/w2091 ) );
  NAND U2450 ( .A(\SUBBYTES[9].a/w2070 ), .B(\SUBBYTES[9].a/w2085 ), .Z(n1317)
         );
  AND U2451 ( .A(\SUBBYTES[9].a/w2087 ), .B(\SUBBYTES[9].a/w2093 ), .Z(
        \SUBBYTES[9].a/w2088 ) );
  AND U2452 ( .A(\SUBBYTES[9].a/w2072 ), .B(\SUBBYTES[9].a/w2070 ), .Z(
        \SUBBYTES[9].a/w2082 ) );
  AND U2453 ( .A(\SUBBYTES[9].a/w2073 ), .B(\SUBBYTES[9].a/w2071 ), .Z(
        \SUBBYTES[9].a/w2080 ) );
  AND U2454 ( .A(\SUBBYTES[9].a/w2087 ), .B(\SUBBYTES[9].a/w2094 ), .Z(
        \SUBBYTES[9].a/w2079 ) );
  AND U2455 ( .A(\SUBBYTES[9].a/w2027 ), .B(\SUBBYTES[9].a/w2023 ), .Z(
        \SUBBYTES[9].a/w2064 ) );
  AND U2456 ( .A(\SUBBYTES[9].a/w2028 ), .B(\SUBBYTES[9].a/w2024 ), .Z(
        \SUBBYTES[9].a/w2062 ) );
  AND U2457 ( .A(\SUBBYTES[9].a/w2154 ), .B(n1314), .Z(\SUBBYTES[9].a/w2061 )
         );
  XNOR U2458 ( .A(\w1[9][49] ), .B(n1321), .Z(n1314) );
  XOR U2459 ( .A(g_input[1201]), .B(\w0[9][49] ), .Z(\w1[9][49] ) );
  AND U2460 ( .A(\w1[9][48] ), .B(\SUBBYTES[9].a/w2029 ), .Z(
        \SUBBYTES[9].a/w2057 ) );
  XOR U2461 ( .A(g_input[1200]), .B(\w0[9][48] ), .Z(\w1[9][48] ) );
  AND U2462 ( .A(\SUBBYTES[9].a/w2030 ), .B(\SUBBYTES[9].a/w2026 ), .Z(
        \SUBBYTES[9].a/w2055 ) );
  AND U2463 ( .A(\SUBBYTES[9].a/w2115 ), .B(\SUBBYTES[9].a/w2147 ), .Z(
        \SUBBYTES[9].a/w2054 ) );
  AND U2464 ( .A(\SUBBYTES[9].a/w2136 ), .B(n1318), .Z(\SUBBYTES[9].a/w2049 )
         );
  XOR U2465 ( .A(\w1[9][52] ), .B(\w1[9][55] ), .Z(n1318) );
  ANDN U2466 ( .A(\SUBBYTES[9].a/w2137 ), .B(n1319), .Z(\SUBBYTES[9].a/w2047 )
         );
  XNOR U2467 ( .A(\w1[9][50] ), .B(\w1[9][55] ), .Z(n1319) );
  IV U2468 ( .A(n1321), .Z(\w1[9][55] ) );
  XNOR U2469 ( .A(g_input[1207]), .B(\w0[9][55] ), .Z(n1321) );
  AND U2470 ( .A(\SUBBYTES[9].a/w2139 ), .B(n1320), .Z(\SUBBYTES[9].a/w2046 )
         );
  XOR U2471 ( .A(\w1[9][50] ), .B(\w1[9][52] ), .Z(n1320) );
  XOR U2472 ( .A(g_input[1204]), .B(\w0[9][52] ), .Z(\w1[9][52] ) );
  XOR U2473 ( .A(g_input[1202]), .B(\w0[9][50] ), .Z(\w1[9][50] ) );
  AND U2474 ( .A(\SUBBYTES[9].a/w164 ), .B(\SUBBYTES[9].a/w160 ), .Z(
        \SUBBYTES[9].a/w201 ) );
  AND U2475 ( .A(\SUBBYTES[9].a/w165 ), .B(\SUBBYTES[9].a/w161 ), .Z(
        \SUBBYTES[9].a/w199 ) );
  AND U2476 ( .A(\SUBBYTES[9].a/w291 ), .B(n1273), .Z(\SUBBYTES[9].a/w198 ) );
  XNOR U2477 ( .A(\w1[9][121] ), .B(n1322), .Z(n1273) );
  XOR U2478 ( .A(g_input[1273]), .B(\w0[9][121] ), .Z(\w1[9][121] ) );
  AND U2479 ( .A(n1323), .B(\SUBBYTES[9].a/w1816 ), .Z(\SUBBYTES[9].a/w1951 )
         );
  AND U2480 ( .A(n1324), .B(\SUBBYTES[9].a/w1817 ), .Z(\SUBBYTES[9].a/w1949 )
         );
  AND U2481 ( .A(\SUBBYTES[9].a/w1947 ), .B(n1325), .Z(\SUBBYTES[9].a/w1948 )
         );
  ANDN U2482 ( .A(\w1[9][56] ), .B(n1326), .Z(\SUBBYTES[9].a/w1944 ) );
  AND U2483 ( .A(n1327), .B(\SUBBYTES[9].a/w1819 ), .Z(\SUBBYTES[9].a/w1942 )
         );
  AND U2484 ( .A(\SUBBYTES[9].a/w1940 ), .B(n1328), .Z(\SUBBYTES[9].a/w1941 )
         );
  XOR U2485 ( .A(\SUBBYTES[9].a/w1884 ), .B(n16088), .Z(n1328) );
  AND U2486 ( .A(\w1[9][120] ), .B(\SUBBYTES[9].a/w166 ), .Z(
        \SUBBYTES[9].a/w194 ) );
  XOR U2487 ( .A(g_input[1272]), .B(\w0[9][120] ), .Z(\w1[9][120] ) );
  AND U2488 ( .A(\SUBBYTES[9].a/w1927 ), .B(\SUBBYTES[9].a/w1929 ), .Z(
        \SUBBYTES[9].a/w1936 ) );
  AND U2489 ( .A(\SUBBYTES[9].a/w1928 ), .B(\SUBBYTES[9].a/w1930 ), .Z(
        \SUBBYTES[9].a/w1934 ) );
  AND U2490 ( .A(\SUBBYTES[9].a/w1931 ), .B(\SUBBYTES[9].a/w1932 ), .Z(
        \SUBBYTES[9].a/w1933 ) );
  AND U2491 ( .A(\SUBBYTES[9].a/w167 ), .B(\SUBBYTES[9].a/w163 ), .Z(
        \SUBBYTES[9].a/w192 ) );
  AND U2492 ( .A(\SUBBYTES[9].a/w1820 ), .B(n1323), .Z(\SUBBYTES[9].a/w1919 )
         );
  XOR U2493 ( .A(\SUBBYTES[9].a/w1888 ), .B(n1093), .Z(n1323) );
  AND U2494 ( .A(\SUBBYTES[9].a/w1821 ), .B(n1324), .Z(\SUBBYTES[9].a/w1917 )
         );
  XOR U2495 ( .A(n16089), .B(\SUBBYTES[9].a/w1888 ), .Z(n1324) );
  AND U2496 ( .A(n1329), .B(n1325), .Z(\SUBBYTES[9].a/w1916 ) );
  XOR U2497 ( .A(n1093), .B(n16089), .Z(n1325) );
  ANDN U2498 ( .A(\SUBBYTES[9].a/w1822 ), .B(n1326), .Z(\SUBBYTES[9].a/w1912 )
         );
  XNOR U2499 ( .A(\SUBBYTES[9].a/w1881 ), .B(\SUBBYTES[9].a/w1884 ), .Z(n1326)
         );
  AND U2500 ( .A(\SUBBYTES[9].a/w1823 ), .B(n1327), .Z(\SUBBYTES[9].a/w1910 )
         );
  XNOR U2501 ( .A(n1330), .B(\SUBBYTES[9].a/w1881 ), .Z(n1327) );
  AND U2502 ( .A(\SUBBYTES[9].a/w252 ), .B(\SUBBYTES[9].a/w284 ), .Z(
        \SUBBYTES[9].a/w191 ) );
  AND U2503 ( .A(\SUBBYTES[9].a/w1908 ), .B(n1331), .Z(\SUBBYTES[9].a/w1909 )
         );
  XOR U2504 ( .A(n1332), .B(n1330), .Z(n1331) );
  IV U2505 ( .A(n16088), .Z(n1330) );
  AND U2506 ( .A(n1333), .B(\SUBBYTES[9].a/w1927 ), .Z(\SUBBYTES[9].a/w1904 )
         );
  ANDN U2507 ( .A(\SUBBYTES[9].a/w1928 ), .B(n1334), .Z(\SUBBYTES[9].a/w1902 )
         );
  AND U2508 ( .A(n1335), .B(\SUBBYTES[9].a/w1931 ), .Z(\SUBBYTES[9].a/w1901 )
         );
  AND U2509 ( .A(\SUBBYTES[9].a/w1887 ), .B(\SUBBYTES[9].a/w1886 ), .Z(
        \SUBBYTES[9].a/w1888 ) );
  IV U2510 ( .A(n1332), .Z(\SUBBYTES[9].a/w1884 ) );
  NAND U2511 ( .A(\SUBBYTES[9].a/w1863 ), .B(\SUBBYTES[9].a/w1878 ), .Z(n1332)
         );
  AND U2512 ( .A(\SUBBYTES[9].a/w1880 ), .B(\SUBBYTES[9].a/w1886 ), .Z(
        \SUBBYTES[9].a/w1881 ) );
  AND U2513 ( .A(\SUBBYTES[9].a/w1865 ), .B(\SUBBYTES[9].a/w1863 ), .Z(
        \SUBBYTES[9].a/w1875 ) );
  AND U2514 ( .A(\SUBBYTES[9].a/w1866 ), .B(\SUBBYTES[9].a/w1864 ), .Z(
        \SUBBYTES[9].a/w1873 ) );
  AND U2515 ( .A(\SUBBYTES[9].a/w1880 ), .B(\SUBBYTES[9].a/w1887 ), .Z(
        \SUBBYTES[9].a/w1872 ) );
  AND U2516 ( .A(\SUBBYTES[9].a/w273 ), .B(n1290), .Z(\SUBBYTES[9].a/w186 ) );
  XOR U2517 ( .A(\w1[9][124] ), .B(\w1[9][127] ), .Z(n1290) );
  AND U2518 ( .A(\SUBBYTES[9].a/w1820 ), .B(\SUBBYTES[9].a/w1816 ), .Z(
        \SUBBYTES[9].a/w1857 ) );
  AND U2519 ( .A(\SUBBYTES[9].a/w1821 ), .B(\SUBBYTES[9].a/w1817 ), .Z(
        \SUBBYTES[9].a/w1855 ) );
  AND U2520 ( .A(\SUBBYTES[9].a/w1947 ), .B(n1329), .Z(\SUBBYTES[9].a/w1854 )
         );
  XNOR U2521 ( .A(\w1[9][57] ), .B(n1336), .Z(n1329) );
  XOR U2522 ( .A(g_input[1209]), .B(\w0[9][57] ), .Z(\w1[9][57] ) );
  AND U2523 ( .A(\w1[9][56] ), .B(\SUBBYTES[9].a/w1822 ), .Z(
        \SUBBYTES[9].a/w1850 ) );
  XOR U2524 ( .A(g_input[1208]), .B(\w0[9][56] ), .Z(\w1[9][56] ) );
  AND U2525 ( .A(\SUBBYTES[9].a/w1823 ), .B(\SUBBYTES[9].a/w1819 ), .Z(
        \SUBBYTES[9].a/w1848 ) );
  AND U2526 ( .A(\SUBBYTES[9].a/w1908 ), .B(\SUBBYTES[9].a/w1940 ), .Z(
        \SUBBYTES[9].a/w1847 ) );
  AND U2527 ( .A(\SUBBYTES[9].a/w1929 ), .B(n1333), .Z(\SUBBYTES[9].a/w1842 )
         );
  XOR U2528 ( .A(\w1[9][60] ), .B(\w1[9][63] ), .Z(n1333) );
  ANDN U2529 ( .A(\SUBBYTES[9].a/w1930 ), .B(n1334), .Z(\SUBBYTES[9].a/w1840 )
         );
  XNOR U2530 ( .A(\w1[9][58] ), .B(\w1[9][63] ), .Z(n1334) );
  IV U2531 ( .A(n1336), .Z(\w1[9][63] ) );
  XNOR U2532 ( .A(g_input[1215]), .B(\w0[9][63] ), .Z(n1336) );
  ANDN U2533 ( .A(\SUBBYTES[9].a/w274 ), .B(n1292), .Z(\SUBBYTES[9].a/w184 )
         );
  XNOR U2534 ( .A(\w1[9][122] ), .B(\w1[9][127] ), .Z(n1292) );
  IV U2535 ( .A(n1322), .Z(\w1[9][127] ) );
  XNOR U2536 ( .A(g_input[1279]), .B(\w0[9][127] ), .Z(n1322) );
  AND U2537 ( .A(\SUBBYTES[9].a/w1932 ), .B(n1335), .Z(\SUBBYTES[9].a/w1839 )
         );
  XOR U2538 ( .A(\w1[9][58] ), .B(\w1[9][60] ), .Z(n1335) );
  XOR U2539 ( .A(g_input[1212]), .B(\w0[9][60] ), .Z(\w1[9][60] ) );
  XOR U2540 ( .A(g_input[1210]), .B(\w0[9][58] ), .Z(\w1[9][58] ) );
  AND U2541 ( .A(\SUBBYTES[9].a/w276 ), .B(n1293), .Z(\SUBBYTES[9].a/w183 ) );
  XOR U2542 ( .A(\w1[9][122] ), .B(\w1[9][124] ), .Z(n1293) );
  XOR U2543 ( .A(g_input[1276]), .B(\w0[9][124] ), .Z(\w1[9][124] ) );
  XOR U2544 ( .A(g_input[1274]), .B(\w0[9][122] ), .Z(\w1[9][122] ) );
  AND U2545 ( .A(n1337), .B(\SUBBYTES[9].a/w1609 ), .Z(\SUBBYTES[9].a/w1744 )
         );
  AND U2546 ( .A(n1338), .B(\SUBBYTES[9].a/w1610 ), .Z(\SUBBYTES[9].a/w1742 )
         );
  AND U2547 ( .A(\SUBBYTES[9].a/w1740 ), .B(n1339), .Z(\SUBBYTES[9].a/w1741 )
         );
  ANDN U2548 ( .A(\w1[9][64] ), .B(n1340), .Z(\SUBBYTES[9].a/w1737 ) );
  AND U2549 ( .A(n1341), .B(\SUBBYTES[9].a/w1612 ), .Z(\SUBBYTES[9].a/w1735 )
         );
  AND U2550 ( .A(\SUBBYTES[9].a/w1733 ), .B(n1342), .Z(\SUBBYTES[9].a/w1734 )
         );
  XOR U2551 ( .A(\SUBBYTES[9].a/w1677 ), .B(n16086), .Z(n1342) );
  AND U2552 ( .A(\SUBBYTES[9].a/w1720 ), .B(\SUBBYTES[9].a/w1722 ), .Z(
        \SUBBYTES[9].a/w1729 ) );
  AND U2553 ( .A(\SUBBYTES[9].a/w1721 ), .B(\SUBBYTES[9].a/w1723 ), .Z(
        \SUBBYTES[9].a/w1727 ) );
  AND U2554 ( .A(\SUBBYTES[9].a/w1724 ), .B(\SUBBYTES[9].a/w1725 ), .Z(
        \SUBBYTES[9].a/w1726 ) );
  AND U2555 ( .A(\SUBBYTES[9].a/w1613 ), .B(n1337), .Z(\SUBBYTES[9].a/w1712 )
         );
  XOR U2556 ( .A(\SUBBYTES[9].a/w1681 ), .B(n1092), .Z(n1337) );
  AND U2557 ( .A(\SUBBYTES[9].a/w1614 ), .B(n1338), .Z(\SUBBYTES[9].a/w1710 )
         );
  XOR U2558 ( .A(n16087), .B(\SUBBYTES[9].a/w1681 ), .Z(n1338) );
  AND U2559 ( .A(n1343), .B(n1339), .Z(\SUBBYTES[9].a/w1709 ) );
  XOR U2560 ( .A(n1092), .B(n16087), .Z(n1339) );
  ANDN U2561 ( .A(\SUBBYTES[9].a/w1615 ), .B(n1340), .Z(\SUBBYTES[9].a/w1705 )
         );
  XNOR U2562 ( .A(\SUBBYTES[9].a/w1674 ), .B(\SUBBYTES[9].a/w1677 ), .Z(n1340)
         );
  AND U2563 ( .A(\SUBBYTES[9].a/w1616 ), .B(n1341), .Z(\SUBBYTES[9].a/w1703 )
         );
  XNOR U2564 ( .A(n1344), .B(\SUBBYTES[9].a/w1674 ), .Z(n1341) );
  AND U2565 ( .A(\SUBBYTES[9].a/w1701 ), .B(n1345), .Z(\SUBBYTES[9].a/w1702 )
         );
  XOR U2566 ( .A(n1346), .B(n1344), .Z(n1345) );
  IV U2567 ( .A(n16086), .Z(n1344) );
  AND U2568 ( .A(n1347), .B(\SUBBYTES[9].a/w1720 ), .Z(\SUBBYTES[9].a/w1697 )
         );
  ANDN U2569 ( .A(\SUBBYTES[9].a/w1721 ), .B(n1348), .Z(\SUBBYTES[9].a/w1695 )
         );
  AND U2570 ( .A(n1349), .B(\SUBBYTES[9].a/w1724 ), .Z(\SUBBYTES[9].a/w1694 )
         );
  AND U2571 ( .A(\SUBBYTES[9].a/w1680 ), .B(\SUBBYTES[9].a/w1679 ), .Z(
        \SUBBYTES[9].a/w1681 ) );
  IV U2572 ( .A(n1346), .Z(\SUBBYTES[9].a/w1677 ) );
  NAND U2573 ( .A(\SUBBYTES[9].a/w1656 ), .B(\SUBBYTES[9].a/w1671 ), .Z(n1346)
         );
  AND U2574 ( .A(\SUBBYTES[9].a/w1673 ), .B(\SUBBYTES[9].a/w1679 ), .Z(
        \SUBBYTES[9].a/w1674 ) );
  AND U2575 ( .A(\SUBBYTES[9].a/w1658 ), .B(\SUBBYTES[9].a/w1656 ), .Z(
        \SUBBYTES[9].a/w1668 ) );
  AND U2576 ( .A(\SUBBYTES[9].a/w1659 ), .B(\SUBBYTES[9].a/w1657 ), .Z(
        \SUBBYTES[9].a/w1666 ) );
  AND U2577 ( .A(\SUBBYTES[9].a/w1673 ), .B(\SUBBYTES[9].a/w1680 ), .Z(
        \SUBBYTES[9].a/w1665 ) );
  AND U2578 ( .A(\SUBBYTES[9].a/w1613 ), .B(\SUBBYTES[9].a/w1609 ), .Z(
        \SUBBYTES[9].a/w1650 ) );
  AND U2579 ( .A(\SUBBYTES[9].a/w1614 ), .B(\SUBBYTES[9].a/w1610 ), .Z(
        \SUBBYTES[9].a/w1648 ) );
  AND U2580 ( .A(\SUBBYTES[9].a/w1740 ), .B(n1343), .Z(\SUBBYTES[9].a/w1647 )
         );
  XNOR U2581 ( .A(\w1[9][65] ), .B(n1350), .Z(n1343) );
  XOR U2582 ( .A(g_input[1217]), .B(\w0[9][65] ), .Z(\w1[9][65] ) );
  AND U2583 ( .A(\w1[9][64] ), .B(\SUBBYTES[9].a/w1615 ), .Z(
        \SUBBYTES[9].a/w1643 ) );
  XOR U2584 ( .A(g_input[1216]), .B(\w0[9][64] ), .Z(\w1[9][64] ) );
  AND U2585 ( .A(\SUBBYTES[9].a/w1616 ), .B(\SUBBYTES[9].a/w1612 ), .Z(
        \SUBBYTES[9].a/w1641 ) );
  AND U2586 ( .A(\SUBBYTES[9].a/w1701 ), .B(\SUBBYTES[9].a/w1733 ), .Z(
        \SUBBYTES[9].a/w1640 ) );
  AND U2587 ( .A(\SUBBYTES[9].a/w1722 ), .B(n1347), .Z(\SUBBYTES[9].a/w1635 )
         );
  XOR U2588 ( .A(\w1[9][68] ), .B(\w1[9][71] ), .Z(n1347) );
  ANDN U2589 ( .A(\SUBBYTES[9].a/w1723 ), .B(n1348), .Z(\SUBBYTES[9].a/w1633 )
         );
  XNOR U2590 ( .A(\w1[9][66] ), .B(\w1[9][71] ), .Z(n1348) );
  IV U2591 ( .A(n1350), .Z(\w1[9][71] ) );
  XNOR U2592 ( .A(g_input[1223]), .B(\w0[9][71] ), .Z(n1350) );
  AND U2593 ( .A(\SUBBYTES[9].a/w1725 ), .B(n1349), .Z(\SUBBYTES[9].a/w1632 )
         );
  XOR U2594 ( .A(\w1[9][66] ), .B(\w1[9][68] ), .Z(n1349) );
  XOR U2595 ( .A(g_input[1220]), .B(\w0[9][68] ), .Z(\w1[9][68] ) );
  XOR U2596 ( .A(g_input[1218]), .B(\w0[9][66] ), .Z(\w1[9][66] ) );
  AND U2597 ( .A(n1351), .B(\SUBBYTES[9].a/w1402 ), .Z(\SUBBYTES[9].a/w1537 )
         );
  AND U2598 ( .A(n1352), .B(\SUBBYTES[9].a/w1403 ), .Z(\SUBBYTES[9].a/w1535 )
         );
  AND U2599 ( .A(\SUBBYTES[9].a/w1533 ), .B(n1353), .Z(\SUBBYTES[9].a/w1534 )
         );
  ANDN U2600 ( .A(\w1[9][72] ), .B(n1354), .Z(\SUBBYTES[9].a/w1530 ) );
  AND U2601 ( .A(n1355), .B(\SUBBYTES[9].a/w1405 ), .Z(\SUBBYTES[9].a/w1528 )
         );
  AND U2602 ( .A(\SUBBYTES[9].a/w1526 ), .B(n1356), .Z(\SUBBYTES[9].a/w1527 )
         );
  XOR U2603 ( .A(\SUBBYTES[9].a/w1470 ), .B(n16084), .Z(n1356) );
  AND U2604 ( .A(\SUBBYTES[9].a/w1513 ), .B(\SUBBYTES[9].a/w1515 ), .Z(
        \SUBBYTES[9].a/w1522 ) );
  AND U2605 ( .A(\SUBBYTES[9].a/w1514 ), .B(\SUBBYTES[9].a/w1516 ), .Z(
        \SUBBYTES[9].a/w1520 ) );
  AND U2606 ( .A(\SUBBYTES[9].a/w1517 ), .B(\SUBBYTES[9].a/w1518 ), .Z(
        \SUBBYTES[9].a/w1519 ) );
  AND U2607 ( .A(\SUBBYTES[9].a/w1406 ), .B(n1351), .Z(\SUBBYTES[9].a/w1505 )
         );
  XOR U2608 ( .A(\SUBBYTES[9].a/w1474 ), .B(n1091), .Z(n1351) );
  AND U2609 ( .A(\SUBBYTES[9].a/w1407 ), .B(n1352), .Z(\SUBBYTES[9].a/w1503 )
         );
  XOR U2610 ( .A(n16085), .B(\SUBBYTES[9].a/w1474 ), .Z(n1352) );
  AND U2611 ( .A(n1357), .B(n1353), .Z(\SUBBYTES[9].a/w1502 ) );
  XOR U2612 ( .A(n1091), .B(n16085), .Z(n1353) );
  ANDN U2613 ( .A(\SUBBYTES[9].a/w1408 ), .B(n1354), .Z(\SUBBYTES[9].a/w1498 )
         );
  XNOR U2614 ( .A(\SUBBYTES[9].a/w1467 ), .B(\SUBBYTES[9].a/w1470 ), .Z(n1354)
         );
  AND U2615 ( .A(\SUBBYTES[9].a/w1409 ), .B(n1355), .Z(\SUBBYTES[9].a/w1496 )
         );
  XNOR U2616 ( .A(n1358), .B(\SUBBYTES[9].a/w1467 ), .Z(n1355) );
  AND U2617 ( .A(\SUBBYTES[9].a/w1494 ), .B(n1359), .Z(\SUBBYTES[9].a/w1495 )
         );
  XOR U2618 ( .A(n1360), .B(n1358), .Z(n1359) );
  IV U2619 ( .A(n16084), .Z(n1358) );
  AND U2620 ( .A(n1361), .B(\SUBBYTES[9].a/w1513 ), .Z(\SUBBYTES[9].a/w1490 )
         );
  ANDN U2621 ( .A(\SUBBYTES[9].a/w1514 ), .B(n1362), .Z(\SUBBYTES[9].a/w1488 )
         );
  AND U2622 ( .A(n1363), .B(\SUBBYTES[9].a/w1517 ), .Z(\SUBBYTES[9].a/w1487 )
         );
  AND U2623 ( .A(\SUBBYTES[9].a/w1473 ), .B(\SUBBYTES[9].a/w1472 ), .Z(
        \SUBBYTES[9].a/w1474 ) );
  IV U2624 ( .A(n1360), .Z(\SUBBYTES[9].a/w1470 ) );
  NAND U2625 ( .A(\SUBBYTES[9].a/w1449 ), .B(\SUBBYTES[9].a/w1464 ), .Z(n1360)
         );
  AND U2626 ( .A(\SUBBYTES[9].a/w1466 ), .B(\SUBBYTES[9].a/w1472 ), .Z(
        \SUBBYTES[9].a/w1467 ) );
  AND U2627 ( .A(\SUBBYTES[9].a/w1451 ), .B(\SUBBYTES[9].a/w1449 ), .Z(
        \SUBBYTES[9].a/w1461 ) );
  AND U2628 ( .A(\SUBBYTES[9].a/w1452 ), .B(\SUBBYTES[9].a/w1450 ), .Z(
        \SUBBYTES[9].a/w1459 ) );
  AND U2629 ( .A(\SUBBYTES[9].a/w1466 ), .B(\SUBBYTES[9].a/w1473 ), .Z(
        \SUBBYTES[9].a/w1458 ) );
  AND U2630 ( .A(\SUBBYTES[9].a/w1406 ), .B(\SUBBYTES[9].a/w1402 ), .Z(
        \SUBBYTES[9].a/w1443 ) );
  AND U2631 ( .A(\SUBBYTES[9].a/w1407 ), .B(\SUBBYTES[9].a/w1403 ), .Z(
        \SUBBYTES[9].a/w1441 ) );
  AND U2632 ( .A(\SUBBYTES[9].a/w1533 ), .B(n1357), .Z(\SUBBYTES[9].a/w1440 )
         );
  XNOR U2633 ( .A(\w1[9][73] ), .B(n1364), .Z(n1357) );
  XOR U2634 ( .A(g_input[1225]), .B(\w0[9][73] ), .Z(\w1[9][73] ) );
  AND U2635 ( .A(\w1[9][72] ), .B(\SUBBYTES[9].a/w1408 ), .Z(
        \SUBBYTES[9].a/w1436 ) );
  XOR U2636 ( .A(g_input[1224]), .B(\w0[9][72] ), .Z(\w1[9][72] ) );
  AND U2637 ( .A(\SUBBYTES[9].a/w1409 ), .B(\SUBBYTES[9].a/w1405 ), .Z(
        \SUBBYTES[9].a/w1434 ) );
  AND U2638 ( .A(\SUBBYTES[9].a/w1494 ), .B(\SUBBYTES[9].a/w1526 ), .Z(
        \SUBBYTES[9].a/w1433 ) );
  AND U2639 ( .A(\SUBBYTES[9].a/w1515 ), .B(n1361), .Z(\SUBBYTES[9].a/w1428 )
         );
  XOR U2640 ( .A(\w1[9][76] ), .B(\w1[9][79] ), .Z(n1361) );
  ANDN U2641 ( .A(\SUBBYTES[9].a/w1516 ), .B(n1362), .Z(\SUBBYTES[9].a/w1426 )
         );
  XNOR U2642 ( .A(\w1[9][74] ), .B(\w1[9][79] ), .Z(n1362) );
  IV U2643 ( .A(n1364), .Z(\w1[9][79] ) );
  XNOR U2644 ( .A(g_input[1231]), .B(\w0[9][79] ), .Z(n1364) );
  AND U2645 ( .A(\SUBBYTES[9].a/w1518 ), .B(n1363), .Z(\SUBBYTES[9].a/w1425 )
         );
  XOR U2646 ( .A(\w1[9][74] ), .B(\w1[9][76] ), .Z(n1363) );
  XOR U2647 ( .A(g_input[1228]), .B(\w0[9][76] ), .Z(\w1[9][76] ) );
  XOR U2648 ( .A(g_input[1226]), .B(\w0[9][74] ), .Z(\w1[9][74] ) );
  AND U2649 ( .A(n1365), .B(\SUBBYTES[9].a/w1195 ), .Z(\SUBBYTES[9].a/w1330 )
         );
  AND U2650 ( .A(n1366), .B(\SUBBYTES[9].a/w1196 ), .Z(\SUBBYTES[9].a/w1328 )
         );
  AND U2651 ( .A(\SUBBYTES[9].a/w1326 ), .B(n1367), .Z(\SUBBYTES[9].a/w1327 )
         );
  ANDN U2652 ( .A(\w1[9][80] ), .B(n1368), .Z(\SUBBYTES[9].a/w1323 ) );
  AND U2653 ( .A(n1369), .B(\SUBBYTES[9].a/w1198 ), .Z(\SUBBYTES[9].a/w1321 )
         );
  AND U2654 ( .A(\SUBBYTES[9].a/w1319 ), .B(n1370), .Z(\SUBBYTES[9].a/w1320 )
         );
  XOR U2655 ( .A(\SUBBYTES[9].a/w1263 ), .B(n16082), .Z(n1370) );
  AND U2656 ( .A(\SUBBYTES[9].a/w1306 ), .B(\SUBBYTES[9].a/w1308 ), .Z(
        \SUBBYTES[9].a/w1315 ) );
  AND U2657 ( .A(\SUBBYTES[9].a/w1307 ), .B(\SUBBYTES[9].a/w1309 ), .Z(
        \SUBBYTES[9].a/w1313 ) );
  AND U2658 ( .A(\SUBBYTES[9].a/w1310 ), .B(\SUBBYTES[9].a/w1311 ), .Z(
        \SUBBYTES[9].a/w1312 ) );
  AND U2659 ( .A(\SUBBYTES[9].a/w1199 ), .B(n1365), .Z(\SUBBYTES[9].a/w1298 )
         );
  XOR U2660 ( .A(\SUBBYTES[9].a/w1267 ), .B(n1090), .Z(n1365) );
  AND U2661 ( .A(\SUBBYTES[9].a/w1200 ), .B(n1366), .Z(\SUBBYTES[9].a/w1296 )
         );
  XOR U2662 ( .A(n16083), .B(\SUBBYTES[9].a/w1267 ), .Z(n1366) );
  AND U2663 ( .A(n1371), .B(n1367), .Z(\SUBBYTES[9].a/w1295 ) );
  XOR U2664 ( .A(n1090), .B(n16083), .Z(n1367) );
  ANDN U2665 ( .A(\SUBBYTES[9].a/w1201 ), .B(n1368), .Z(\SUBBYTES[9].a/w1291 )
         );
  XNOR U2666 ( .A(\SUBBYTES[9].a/w1260 ), .B(\SUBBYTES[9].a/w1263 ), .Z(n1368)
         );
  AND U2667 ( .A(\SUBBYTES[9].a/w1202 ), .B(n1369), .Z(\SUBBYTES[9].a/w1289 )
         );
  XNOR U2668 ( .A(n1372), .B(\SUBBYTES[9].a/w1260 ), .Z(n1369) );
  AND U2669 ( .A(\SUBBYTES[9].a/w1287 ), .B(n1373), .Z(\SUBBYTES[9].a/w1288 )
         );
  XOR U2670 ( .A(n1374), .B(n1372), .Z(n1373) );
  IV U2671 ( .A(n16082), .Z(n1372) );
  AND U2672 ( .A(n1375), .B(\SUBBYTES[9].a/w1306 ), .Z(\SUBBYTES[9].a/w1283 )
         );
  ANDN U2673 ( .A(\SUBBYTES[9].a/w1307 ), .B(n1376), .Z(\SUBBYTES[9].a/w1281 )
         );
  AND U2674 ( .A(n1377), .B(\SUBBYTES[9].a/w1310 ), .Z(\SUBBYTES[9].a/w1280 )
         );
  AND U2675 ( .A(\SUBBYTES[9].a/w1266 ), .B(\SUBBYTES[9].a/w1265 ), .Z(
        \SUBBYTES[9].a/w1267 ) );
  IV U2676 ( .A(n1374), .Z(\SUBBYTES[9].a/w1263 ) );
  NAND U2677 ( .A(\SUBBYTES[9].a/w1242 ), .B(\SUBBYTES[9].a/w1257 ), .Z(n1374)
         );
  AND U2678 ( .A(\SUBBYTES[9].a/w1259 ), .B(\SUBBYTES[9].a/w1265 ), .Z(
        \SUBBYTES[9].a/w1260 ) );
  AND U2679 ( .A(\SUBBYTES[9].a/w1244 ), .B(\SUBBYTES[9].a/w1242 ), .Z(
        \SUBBYTES[9].a/w1254 ) );
  AND U2680 ( .A(\SUBBYTES[9].a/w1245 ), .B(\SUBBYTES[9].a/w1243 ), .Z(
        \SUBBYTES[9].a/w1252 ) );
  AND U2681 ( .A(\SUBBYTES[9].a/w1259 ), .B(\SUBBYTES[9].a/w1266 ), .Z(
        \SUBBYTES[9].a/w1251 ) );
  AND U2682 ( .A(\SUBBYTES[9].a/w1199 ), .B(\SUBBYTES[9].a/w1195 ), .Z(
        \SUBBYTES[9].a/w1236 ) );
  AND U2683 ( .A(\SUBBYTES[9].a/w1200 ), .B(\SUBBYTES[9].a/w1196 ), .Z(
        \SUBBYTES[9].a/w1234 ) );
  AND U2684 ( .A(\SUBBYTES[9].a/w1326 ), .B(n1371), .Z(\SUBBYTES[9].a/w1233 )
         );
  XNOR U2685 ( .A(\w1[9][81] ), .B(n1378), .Z(n1371) );
  XOR U2686 ( .A(g_input[1233]), .B(\w0[9][81] ), .Z(\w1[9][81] ) );
  AND U2687 ( .A(\w1[9][80] ), .B(\SUBBYTES[9].a/w1201 ), .Z(
        \SUBBYTES[9].a/w1229 ) );
  XOR U2688 ( .A(g_input[1232]), .B(\w0[9][80] ), .Z(\w1[9][80] ) );
  AND U2689 ( .A(\SUBBYTES[9].a/w1202 ), .B(\SUBBYTES[9].a/w1198 ), .Z(
        \SUBBYTES[9].a/w1227 ) );
  AND U2690 ( .A(\SUBBYTES[9].a/w1287 ), .B(\SUBBYTES[9].a/w1319 ), .Z(
        \SUBBYTES[9].a/w1226 ) );
  AND U2691 ( .A(\SUBBYTES[9].a/w1308 ), .B(n1375), .Z(\SUBBYTES[9].a/w1221 )
         );
  XOR U2692 ( .A(\w1[9][84] ), .B(\w1[9][87] ), .Z(n1375) );
  ANDN U2693 ( .A(\SUBBYTES[9].a/w1309 ), .B(n1376), .Z(\SUBBYTES[9].a/w1219 )
         );
  XNOR U2694 ( .A(\w1[9][82] ), .B(\w1[9][87] ), .Z(n1376) );
  IV U2695 ( .A(n1378), .Z(\w1[9][87] ) );
  XNOR U2696 ( .A(g_input[1239]), .B(\w0[9][87] ), .Z(n1378) );
  AND U2697 ( .A(\SUBBYTES[9].a/w1311 ), .B(n1377), .Z(\SUBBYTES[9].a/w1218 )
         );
  XOR U2698 ( .A(\w1[9][82] ), .B(\w1[9][84] ), .Z(n1377) );
  XOR U2699 ( .A(g_input[1236]), .B(\w0[9][84] ), .Z(\w1[9][84] ) );
  XOR U2700 ( .A(g_input[1234]), .B(\w0[9][82] ), .Z(\w1[9][82] ) );
  AND U2701 ( .A(n1379), .B(\SUBBYTES[9].a/w988 ), .Z(\SUBBYTES[9].a/w1123 )
         );
  AND U2702 ( .A(n1380), .B(\SUBBYTES[9].a/w989 ), .Z(\SUBBYTES[9].a/w1121 )
         );
  AND U2703 ( .A(\SUBBYTES[9].a/w1119 ), .B(n1381), .Z(\SUBBYTES[9].a/w1120 )
         );
  ANDN U2704 ( .A(\w1[9][88] ), .B(n1382), .Z(\SUBBYTES[9].a/w1116 ) );
  AND U2705 ( .A(n1383), .B(\SUBBYTES[9].a/w991 ), .Z(\SUBBYTES[9].a/w1114 )
         );
  AND U2706 ( .A(\SUBBYTES[9].a/w1112 ), .B(n1384), .Z(\SUBBYTES[9].a/w1113 )
         );
  XOR U2707 ( .A(\SUBBYTES[9].a/w1056 ), .B(n16080), .Z(n1384) );
  AND U2708 ( .A(\SUBBYTES[9].a/w1099 ), .B(\SUBBYTES[9].a/w1101 ), .Z(
        \SUBBYTES[9].a/w1108 ) );
  AND U2709 ( .A(\SUBBYTES[9].a/w1100 ), .B(\SUBBYTES[9].a/w1102 ), .Z(
        \SUBBYTES[9].a/w1106 ) );
  AND U2710 ( .A(\SUBBYTES[9].a/w1103 ), .B(\SUBBYTES[9].a/w1104 ), .Z(
        \SUBBYTES[9].a/w1105 ) );
  AND U2711 ( .A(\SUBBYTES[9].a/w992 ), .B(n1379), .Z(\SUBBYTES[9].a/w1091 )
         );
  XOR U2712 ( .A(\SUBBYTES[9].a/w1060 ), .B(n1089), .Z(n1379) );
  AND U2713 ( .A(\SUBBYTES[9].a/w993 ), .B(n1380), .Z(\SUBBYTES[9].a/w1089 )
         );
  XOR U2714 ( .A(n16081), .B(\SUBBYTES[9].a/w1060 ), .Z(n1380) );
  AND U2715 ( .A(n1385), .B(n1381), .Z(\SUBBYTES[9].a/w1088 ) );
  XOR U2716 ( .A(n1089), .B(n16081), .Z(n1381) );
  ANDN U2717 ( .A(\SUBBYTES[9].a/w994 ), .B(n1382), .Z(\SUBBYTES[9].a/w1084 )
         );
  XNOR U2718 ( .A(\SUBBYTES[9].a/w1053 ), .B(\SUBBYTES[9].a/w1056 ), .Z(n1382)
         );
  AND U2719 ( .A(\SUBBYTES[9].a/w995 ), .B(n1383), .Z(\SUBBYTES[9].a/w1082 )
         );
  XNOR U2720 ( .A(n1386), .B(\SUBBYTES[9].a/w1053 ), .Z(n1383) );
  AND U2721 ( .A(\SUBBYTES[9].a/w1080 ), .B(n1387), .Z(\SUBBYTES[9].a/w1081 )
         );
  XOR U2722 ( .A(n1388), .B(n1386), .Z(n1387) );
  IV U2723 ( .A(n16080), .Z(n1386) );
  AND U2724 ( .A(n1389), .B(\SUBBYTES[9].a/w1099 ), .Z(\SUBBYTES[9].a/w1076 )
         );
  ANDN U2725 ( .A(\SUBBYTES[9].a/w1100 ), .B(n1390), .Z(\SUBBYTES[9].a/w1074 )
         );
  AND U2726 ( .A(n1391), .B(\SUBBYTES[9].a/w1103 ), .Z(\SUBBYTES[9].a/w1073 )
         );
  AND U2727 ( .A(\SUBBYTES[9].a/w1059 ), .B(\SUBBYTES[9].a/w1058 ), .Z(
        \SUBBYTES[9].a/w1060 ) );
  IV U2728 ( .A(n1388), .Z(\SUBBYTES[9].a/w1056 ) );
  NAND U2729 ( .A(\SUBBYTES[9].a/w1035 ), .B(\SUBBYTES[9].a/w1050 ), .Z(n1388)
         );
  AND U2730 ( .A(\SUBBYTES[9].a/w1052 ), .B(\SUBBYTES[9].a/w1058 ), .Z(
        \SUBBYTES[9].a/w1053 ) );
  AND U2731 ( .A(\SUBBYTES[9].a/w1037 ), .B(\SUBBYTES[9].a/w1035 ), .Z(
        \SUBBYTES[9].a/w1047 ) );
  AND U2732 ( .A(\SUBBYTES[9].a/w1038 ), .B(\SUBBYTES[9].a/w1036 ), .Z(
        \SUBBYTES[9].a/w1045 ) );
  AND U2733 ( .A(\SUBBYTES[9].a/w1052 ), .B(\SUBBYTES[9].a/w1059 ), .Z(
        \SUBBYTES[9].a/w1044 ) );
  AND U2734 ( .A(\SUBBYTES[9].a/w992 ), .B(\SUBBYTES[9].a/w988 ), .Z(
        \SUBBYTES[9].a/w1029 ) );
  AND U2735 ( .A(\SUBBYTES[9].a/w993 ), .B(\SUBBYTES[9].a/w989 ), .Z(
        \SUBBYTES[9].a/w1027 ) );
  AND U2736 ( .A(\SUBBYTES[9].a/w1119 ), .B(n1385), .Z(\SUBBYTES[9].a/w1026 )
         );
  XNOR U2737 ( .A(\w1[9][89] ), .B(n1392), .Z(n1385) );
  XOR U2738 ( .A(g_input[1241]), .B(\w0[9][89] ), .Z(\w1[9][89] ) );
  AND U2739 ( .A(\w1[9][88] ), .B(\SUBBYTES[9].a/w994 ), .Z(
        \SUBBYTES[9].a/w1022 ) );
  XOR U2740 ( .A(g_input[1240]), .B(\w0[9][88] ), .Z(\w1[9][88] ) );
  AND U2741 ( .A(\SUBBYTES[9].a/w995 ), .B(\SUBBYTES[9].a/w991 ), .Z(
        \SUBBYTES[9].a/w1020 ) );
  AND U2742 ( .A(\SUBBYTES[9].a/w1080 ), .B(\SUBBYTES[9].a/w1112 ), .Z(
        \SUBBYTES[9].a/w1019 ) );
  AND U2743 ( .A(\SUBBYTES[9].a/w1101 ), .B(n1389), .Z(\SUBBYTES[9].a/w1014 )
         );
  XOR U2744 ( .A(\w1[9][92] ), .B(\w1[9][95] ), .Z(n1389) );
  ANDN U2745 ( .A(\SUBBYTES[9].a/w1102 ), .B(n1390), .Z(\SUBBYTES[9].a/w1012 )
         );
  XNOR U2746 ( .A(\w1[9][90] ), .B(\w1[9][95] ), .Z(n1390) );
  IV U2747 ( .A(n1392), .Z(\w1[9][95] ) );
  XNOR U2748 ( .A(g_input[1247]), .B(\w0[9][95] ), .Z(n1392) );
  AND U2749 ( .A(\SUBBYTES[9].a/w1104 ), .B(n1391), .Z(\SUBBYTES[9].a/w1011 )
         );
  XOR U2750 ( .A(\w1[9][90] ), .B(\w1[9][92] ), .Z(n1391) );
  XOR U2751 ( .A(g_input[1244]), .B(\w0[9][92] ), .Z(\w1[9][92] ) );
  XOR U2752 ( .A(g_input[1242]), .B(\w0[9][90] ), .Z(\w1[9][90] ) );
  AND U2753 ( .A(\SUBBYTES[9].a/w2084 ), .B(\SUBBYTES[9].a/w2071 ), .Z(n16090)
         );
  AND U2754 ( .A(\SUBBYTES[9].a/w1877 ), .B(\SUBBYTES[9].a/w1866 ), .Z(n16089)
         );
  AND U2755 ( .A(\SUBBYTES[9].a/w221 ), .B(\SUBBYTES[9].a/w208 ), .Z(n16072)
         );
  AND U2756 ( .A(\SUBBYTES[9].a/w1877 ), .B(\SUBBYTES[9].a/w1864 ), .Z(n16088)
         );
  AND U2757 ( .A(\SUBBYTES[9].a/w1670 ), .B(\SUBBYTES[9].a/w1659 ), .Z(n16087)
         );
  AND U2758 ( .A(\SUBBYTES[9].a/w1670 ), .B(\SUBBYTES[9].a/w1657 ), .Z(n16086)
         );
  AND U2759 ( .A(\SUBBYTES[9].a/w1463 ), .B(\SUBBYTES[9].a/w1452 ), .Z(n16085)
         );
  AND U2760 ( .A(\SUBBYTES[9].a/w1463 ), .B(\SUBBYTES[9].a/w1450 ), .Z(n16084)
         );
  AND U2761 ( .A(\SUBBYTES[9].a/w1256 ), .B(\SUBBYTES[9].a/w1245 ), .Z(n16083)
         );
  AND U2762 ( .A(\SUBBYTES[9].a/w1256 ), .B(\SUBBYTES[9].a/w1243 ), .Z(n16082)
         );
  AND U2763 ( .A(\SUBBYTES[9].a/w1049 ), .B(\SUBBYTES[9].a/w1038 ), .Z(n16081)
         );
  AND U2764 ( .A(\SUBBYTES[9].a/w1049 ), .B(\SUBBYTES[9].a/w1036 ), .Z(n16080)
         );
  AND U2765 ( .A(\SUBBYTES[9].a/w842 ), .B(\SUBBYTES[9].a/w831 ), .Z(n16079)
         );
  AND U2766 ( .A(\SUBBYTES[9].a/w842 ), .B(\SUBBYTES[9].a/w829 ), .Z(n16078)
         );
  AND U2767 ( .A(\SUBBYTES[9].a/w635 ), .B(\SUBBYTES[9].a/w624 ), .Z(n16077)
         );
  AND U2768 ( .A(\SUBBYTES[9].a/w635 ), .B(\SUBBYTES[9].a/w622 ), .Z(n16076)
         );
  AND U2769 ( .A(\SUBBYTES[9].a/w428 ), .B(\SUBBYTES[9].a/w417 ), .Z(n16075)
         );
  AND U2770 ( .A(\SUBBYTES[9].a/w428 ), .B(\SUBBYTES[9].a/w415 ), .Z(n16074)
         );
  AND U2771 ( .A(\SUBBYTES[9].a/w3326 ), .B(\SUBBYTES[9].a/w3315 ), .Z(n16103)
         );
  AND U2772 ( .A(\SUBBYTES[9].a/w3326 ), .B(\SUBBYTES[9].a/w3313 ), .Z(n16102)
         );
  AND U2773 ( .A(\SUBBYTES[9].a/w3119 ), .B(\SUBBYTES[9].a/w3108 ), .Z(n16101)
         );
  AND U2774 ( .A(\SUBBYTES[9].a/w3119 ), .B(\SUBBYTES[9].a/w3106 ), .Z(n16100)
         );
  AND U2775 ( .A(\SUBBYTES[9].a/w2912 ), .B(\SUBBYTES[9].a/w2901 ), .Z(n16099)
         );
  AND U2776 ( .A(\SUBBYTES[9].a/w2912 ), .B(\SUBBYTES[9].a/w2899 ), .Z(n16098)
         );
  AND U2777 ( .A(\SUBBYTES[9].a/w2705 ), .B(\SUBBYTES[9].a/w2694 ), .Z(n16097)
         );
  AND U2778 ( .A(\SUBBYTES[9].a/w2705 ), .B(\SUBBYTES[9].a/w2692 ), .Z(n16096)
         );
  AND U2779 ( .A(\SUBBYTES[9].a/w2498 ), .B(\SUBBYTES[9].a/w2487 ), .Z(n16095)
         );
  AND U2780 ( .A(\SUBBYTES[9].a/w2498 ), .B(\SUBBYTES[9].a/w2485 ), .Z(n16094)
         );
  AND U2781 ( .A(\SUBBYTES[9].a/w2291 ), .B(\SUBBYTES[9].a/w2280 ), .Z(n16093)
         );
  AND U2782 ( .A(\SUBBYTES[9].a/w2291 ), .B(\SUBBYTES[9].a/w2278 ), .Z(n16092)
         );
  AND U2783 ( .A(\SUBBYTES[9].a/w2084 ), .B(\SUBBYTES[9].a/w2073 ), .Z(n16091)
         );
  AND U2784 ( .A(\SUBBYTES[9].a/w221 ), .B(\SUBBYTES[9].a/w210 ), .Z(n16073)
         );
  AND U2785 ( .A(n1393), .B(\SUBBYTES[8].a/w781 ), .Z(\SUBBYTES[8].a/w916 ) );
  AND U2786 ( .A(n1394), .B(\SUBBYTES[8].a/w782 ), .Z(\SUBBYTES[8].a/w914 ) );
  AND U2787 ( .A(\SUBBYTES[8].a/w912 ), .B(n1395), .Z(\SUBBYTES[8].a/w913 ) );
  ANDN U2788 ( .A(\w1[8][96] ), .B(n1396), .Z(\SUBBYTES[8].a/w909 ) );
  AND U2789 ( .A(n1397), .B(\SUBBYTES[8].a/w784 ), .Z(\SUBBYTES[8].a/w907 ) );
  AND U2790 ( .A(\SUBBYTES[8].a/w905 ), .B(n1398), .Z(\SUBBYTES[8].a/w906 ) );
  XOR U2791 ( .A(\SUBBYTES[8].a/w849 ), .B(n14798), .Z(n1398) );
  AND U2792 ( .A(\SUBBYTES[8].a/w892 ), .B(\SUBBYTES[8].a/w894 ), .Z(
        \SUBBYTES[8].a/w901 ) );
  AND U2793 ( .A(\SUBBYTES[8].a/w893 ), .B(\SUBBYTES[8].a/w895 ), .Z(
        \SUBBYTES[8].a/w899 ) );
  AND U2794 ( .A(\SUBBYTES[8].a/w896 ), .B(\SUBBYTES[8].a/w897 ), .Z(
        \SUBBYTES[8].a/w898 ) );
  AND U2795 ( .A(\SUBBYTES[8].a/w785 ), .B(n1393), .Z(\SUBBYTES[8].a/w884 ) );
  XOR U2796 ( .A(\SUBBYTES[8].a/w853 ), .B(n1072), .Z(n1393) );
  AND U2797 ( .A(\SUBBYTES[8].a/w786 ), .B(n1394), .Z(\SUBBYTES[8].a/w882 ) );
  XOR U2798 ( .A(n14799), .B(\SUBBYTES[8].a/w853 ), .Z(n1394) );
  ANDN U2799 ( .A(n1395), .B(n1399), .Z(\SUBBYTES[8].a/w881 ) );
  XOR U2800 ( .A(n1072), .B(n14799), .Z(n1395) );
  ANDN U2801 ( .A(\SUBBYTES[8].a/w787 ), .B(n1396), .Z(\SUBBYTES[8].a/w877 )
         );
  XNOR U2802 ( .A(\SUBBYTES[8].a/w846 ), .B(\SUBBYTES[8].a/w849 ), .Z(n1396)
         );
  AND U2803 ( .A(\SUBBYTES[8].a/w788 ), .B(n1397), .Z(\SUBBYTES[8].a/w875 ) );
  XNOR U2804 ( .A(n1400), .B(\SUBBYTES[8].a/w846 ), .Z(n1397) );
  AND U2805 ( .A(\SUBBYTES[8].a/w873 ), .B(n1401), .Z(\SUBBYTES[8].a/w874 ) );
  XOR U2806 ( .A(n1402), .B(n1400), .Z(n1401) );
  IV U2807 ( .A(n14798), .Z(n1400) );
  ANDN U2808 ( .A(\SUBBYTES[8].a/w892 ), .B(n1403), .Z(\SUBBYTES[8].a/w869 )
         );
  ANDN U2809 ( .A(\SUBBYTES[8].a/w893 ), .B(n1404), .Z(\SUBBYTES[8].a/w867 )
         );
  ANDN U2810 ( .A(\SUBBYTES[8].a/w896 ), .B(n1405), .Z(\SUBBYTES[8].a/w866 )
         );
  AND U2811 ( .A(\SUBBYTES[8].a/w852 ), .B(\SUBBYTES[8].a/w851 ), .Z(
        \SUBBYTES[8].a/w853 ) );
  IV U2812 ( .A(n1402), .Z(\SUBBYTES[8].a/w849 ) );
  NAND U2813 ( .A(\SUBBYTES[8].a/w828 ), .B(\SUBBYTES[8].a/w843 ), .Z(n1402)
         );
  AND U2814 ( .A(\SUBBYTES[8].a/w845 ), .B(\SUBBYTES[8].a/w851 ), .Z(
        \SUBBYTES[8].a/w846 ) );
  AND U2815 ( .A(\SUBBYTES[8].a/w830 ), .B(\SUBBYTES[8].a/w828 ), .Z(
        \SUBBYTES[8].a/w840 ) );
  AND U2816 ( .A(\SUBBYTES[8].a/w831 ), .B(\SUBBYTES[8].a/w829 ), .Z(
        \SUBBYTES[8].a/w838 ) );
  AND U2817 ( .A(\SUBBYTES[8].a/w845 ), .B(\SUBBYTES[8].a/w852 ), .Z(
        \SUBBYTES[8].a/w837 ) );
  AND U2818 ( .A(\SUBBYTES[8].a/w785 ), .B(\SUBBYTES[8].a/w781 ), .Z(
        \SUBBYTES[8].a/w822 ) );
  AND U2819 ( .A(\SUBBYTES[8].a/w786 ), .B(\SUBBYTES[8].a/w782 ), .Z(
        \SUBBYTES[8].a/w820 ) );
  ANDN U2820 ( .A(\SUBBYTES[8].a/w912 ), .B(n1399), .Z(\SUBBYTES[8].a/w819 )
         );
  XNOR U2821 ( .A(\w1[8][103] ), .B(\w1[8][97] ), .Z(n1399) );
  XOR U2822 ( .A(\w0[8][97] ), .B(g_input[1121]), .Z(\w1[8][97] ) );
  IV U2823 ( .A(n1406), .Z(\w1[8][103] ) );
  AND U2824 ( .A(\w1[8][96] ), .B(\SUBBYTES[8].a/w787 ), .Z(
        \SUBBYTES[8].a/w815 ) );
  XOR U2825 ( .A(\w0[8][96] ), .B(g_input[1120]), .Z(\w1[8][96] ) );
  AND U2826 ( .A(\SUBBYTES[8].a/w788 ), .B(\SUBBYTES[8].a/w784 ), .Z(
        \SUBBYTES[8].a/w813 ) );
  AND U2827 ( .A(\SUBBYTES[8].a/w873 ), .B(\SUBBYTES[8].a/w905 ), .Z(
        \SUBBYTES[8].a/w812 ) );
  ANDN U2828 ( .A(\SUBBYTES[8].a/w894 ), .B(n1403), .Z(\SUBBYTES[8].a/w807 )
         );
  XOR U2829 ( .A(\w1[8][100] ), .B(n1406), .Z(n1403) );
  ANDN U2830 ( .A(\SUBBYTES[8].a/w895 ), .B(n1404), .Z(\SUBBYTES[8].a/w805 )
         );
  XOR U2831 ( .A(n1406), .B(\w1[8][98] ), .Z(n1404) );
  XNOR U2832 ( .A(\w0[8][103] ), .B(g_input[1127]), .Z(n1406) );
  ANDN U2833 ( .A(\SUBBYTES[8].a/w897 ), .B(n1405), .Z(\SUBBYTES[8].a/w804 )
         );
  XNOR U2834 ( .A(\w1[8][100] ), .B(\w1[8][98] ), .Z(n1405) );
  XOR U2835 ( .A(\w0[8][98] ), .B(g_input[1122]), .Z(\w1[8][98] ) );
  XOR U2836 ( .A(\w0[8][100] ), .B(g_input[1124]), .Z(\w1[8][100] ) );
  AND U2837 ( .A(n1407), .B(\SUBBYTES[8].a/w574 ), .Z(\SUBBYTES[8].a/w709 ) );
  AND U2838 ( .A(n1408), .B(\SUBBYTES[8].a/w575 ), .Z(\SUBBYTES[8].a/w707 ) );
  AND U2839 ( .A(\SUBBYTES[8].a/w705 ), .B(n1409), .Z(\SUBBYTES[8].a/w706 ) );
  ANDN U2840 ( .A(\w1[8][104] ), .B(n1410), .Z(\SUBBYTES[8].a/w702 ) );
  AND U2841 ( .A(n1411), .B(\SUBBYTES[8].a/w577 ), .Z(\SUBBYTES[8].a/w700 ) );
  AND U2842 ( .A(\SUBBYTES[8].a/w698 ), .B(n1412), .Z(\SUBBYTES[8].a/w699 ) );
  XOR U2843 ( .A(\SUBBYTES[8].a/w642 ), .B(n14796), .Z(n1412) );
  AND U2844 ( .A(\SUBBYTES[8].a/w685 ), .B(\SUBBYTES[8].a/w687 ), .Z(
        \SUBBYTES[8].a/w694 ) );
  AND U2845 ( .A(\SUBBYTES[8].a/w686 ), .B(\SUBBYTES[8].a/w688 ), .Z(
        \SUBBYTES[8].a/w692 ) );
  AND U2846 ( .A(\SUBBYTES[8].a/w689 ), .B(\SUBBYTES[8].a/w690 ), .Z(
        \SUBBYTES[8].a/w691 ) );
  AND U2847 ( .A(\SUBBYTES[8].a/w578 ), .B(n1407), .Z(\SUBBYTES[8].a/w677 ) );
  XOR U2848 ( .A(\SUBBYTES[8].a/w646 ), .B(n1071), .Z(n1407) );
  AND U2849 ( .A(\SUBBYTES[8].a/w579 ), .B(n1408), .Z(\SUBBYTES[8].a/w675 ) );
  XOR U2850 ( .A(n14797), .B(\SUBBYTES[8].a/w646 ), .Z(n1408) );
  ANDN U2851 ( .A(n1409), .B(n1413), .Z(\SUBBYTES[8].a/w674 ) );
  XOR U2852 ( .A(n1071), .B(n14797), .Z(n1409) );
  ANDN U2853 ( .A(\SUBBYTES[8].a/w580 ), .B(n1410), .Z(\SUBBYTES[8].a/w670 )
         );
  XNOR U2854 ( .A(\SUBBYTES[8].a/w639 ), .B(\SUBBYTES[8].a/w642 ), .Z(n1410)
         );
  AND U2855 ( .A(\SUBBYTES[8].a/w581 ), .B(n1411), .Z(\SUBBYTES[8].a/w668 ) );
  XNOR U2856 ( .A(n1414), .B(\SUBBYTES[8].a/w639 ), .Z(n1411) );
  AND U2857 ( .A(\SUBBYTES[8].a/w666 ), .B(n1415), .Z(\SUBBYTES[8].a/w667 ) );
  XOR U2858 ( .A(n1416), .B(n1414), .Z(n1415) );
  IV U2859 ( .A(n14796), .Z(n1414) );
  ANDN U2860 ( .A(\SUBBYTES[8].a/w685 ), .B(n1417), .Z(\SUBBYTES[8].a/w662 )
         );
  ANDN U2861 ( .A(\SUBBYTES[8].a/w686 ), .B(n1418), .Z(\SUBBYTES[8].a/w660 )
         );
  ANDN U2862 ( .A(\SUBBYTES[8].a/w689 ), .B(n1419), .Z(\SUBBYTES[8].a/w659 )
         );
  AND U2863 ( .A(\SUBBYTES[8].a/w645 ), .B(\SUBBYTES[8].a/w644 ), .Z(
        \SUBBYTES[8].a/w646 ) );
  IV U2864 ( .A(n1416), .Z(\SUBBYTES[8].a/w642 ) );
  NAND U2865 ( .A(\SUBBYTES[8].a/w621 ), .B(\SUBBYTES[8].a/w636 ), .Z(n1416)
         );
  AND U2866 ( .A(\SUBBYTES[8].a/w638 ), .B(\SUBBYTES[8].a/w644 ), .Z(
        \SUBBYTES[8].a/w639 ) );
  AND U2867 ( .A(\SUBBYTES[8].a/w623 ), .B(\SUBBYTES[8].a/w621 ), .Z(
        \SUBBYTES[8].a/w633 ) );
  AND U2868 ( .A(\SUBBYTES[8].a/w624 ), .B(\SUBBYTES[8].a/w622 ), .Z(
        \SUBBYTES[8].a/w631 ) );
  AND U2869 ( .A(\SUBBYTES[8].a/w638 ), .B(\SUBBYTES[8].a/w645 ), .Z(
        \SUBBYTES[8].a/w630 ) );
  AND U2870 ( .A(\SUBBYTES[8].a/w578 ), .B(\SUBBYTES[8].a/w574 ), .Z(
        \SUBBYTES[8].a/w615 ) );
  AND U2871 ( .A(\SUBBYTES[8].a/w579 ), .B(\SUBBYTES[8].a/w575 ), .Z(
        \SUBBYTES[8].a/w613 ) );
  ANDN U2872 ( .A(\SUBBYTES[8].a/w705 ), .B(n1413), .Z(\SUBBYTES[8].a/w612 )
         );
  XNOR U2873 ( .A(\w1[8][105] ), .B(\w1[8][111] ), .Z(n1413) );
  XOR U2874 ( .A(\w0[8][105] ), .B(g_input[1129]), .Z(\w1[8][105] ) );
  AND U2875 ( .A(\w1[8][104] ), .B(\SUBBYTES[8].a/w580 ), .Z(
        \SUBBYTES[8].a/w608 ) );
  XOR U2876 ( .A(\w0[8][104] ), .B(g_input[1128]), .Z(\w1[8][104] ) );
  AND U2877 ( .A(\SUBBYTES[8].a/w581 ), .B(\SUBBYTES[8].a/w577 ), .Z(
        \SUBBYTES[8].a/w606 ) );
  AND U2878 ( .A(\SUBBYTES[8].a/w666 ), .B(\SUBBYTES[8].a/w698 ), .Z(
        \SUBBYTES[8].a/w605 ) );
  ANDN U2879 ( .A(\SUBBYTES[8].a/w687 ), .B(n1417), .Z(\SUBBYTES[8].a/w600 )
         );
  XNOR U2880 ( .A(\w1[8][108] ), .B(\w1[8][111] ), .Z(n1417) );
  ANDN U2881 ( .A(\SUBBYTES[8].a/w688 ), .B(n1418), .Z(\SUBBYTES[8].a/w598 )
         );
  XNOR U2882 ( .A(\w1[8][106] ), .B(\w1[8][111] ), .Z(n1418) );
  XOR U2883 ( .A(\w0[8][111] ), .B(g_input[1135]), .Z(\w1[8][111] ) );
  IV U2884 ( .A(n1420), .Z(\w1[8][106] ) );
  ANDN U2885 ( .A(\SUBBYTES[8].a/w690 ), .B(n1419), .Z(\SUBBYTES[8].a/w597 )
         );
  XOR U2886 ( .A(n1420), .B(\w1[8][108] ), .Z(n1419) );
  XOR U2887 ( .A(\w0[8][108] ), .B(g_input[1132]), .Z(\w1[8][108] ) );
  XNOR U2888 ( .A(\w0[8][106] ), .B(g_input[1130]), .Z(n1420) );
  AND U2889 ( .A(n1421), .B(\SUBBYTES[8].a/w367 ), .Z(\SUBBYTES[8].a/w502 ) );
  AND U2890 ( .A(n1422), .B(\SUBBYTES[8].a/w368 ), .Z(\SUBBYTES[8].a/w500 ) );
  AND U2891 ( .A(\SUBBYTES[8].a/w498 ), .B(n1423), .Z(\SUBBYTES[8].a/w499 ) );
  ANDN U2892 ( .A(\w1[8][112] ), .B(n1424), .Z(\SUBBYTES[8].a/w495 ) );
  AND U2893 ( .A(n1425), .B(\SUBBYTES[8].a/w370 ), .Z(\SUBBYTES[8].a/w493 ) );
  AND U2894 ( .A(\SUBBYTES[8].a/w491 ), .B(n1426), .Z(\SUBBYTES[8].a/w492 ) );
  XOR U2895 ( .A(\SUBBYTES[8].a/w435 ), .B(n14794), .Z(n1426) );
  AND U2896 ( .A(\SUBBYTES[8].a/w478 ), .B(\SUBBYTES[8].a/w480 ), .Z(
        \SUBBYTES[8].a/w487 ) );
  AND U2897 ( .A(\SUBBYTES[8].a/w479 ), .B(\SUBBYTES[8].a/w481 ), .Z(
        \SUBBYTES[8].a/w485 ) );
  AND U2898 ( .A(\SUBBYTES[8].a/w482 ), .B(\SUBBYTES[8].a/w483 ), .Z(
        \SUBBYTES[8].a/w484 ) );
  AND U2899 ( .A(\SUBBYTES[8].a/w371 ), .B(n1421), .Z(\SUBBYTES[8].a/w470 ) );
  XOR U2900 ( .A(\SUBBYTES[8].a/w439 ), .B(n1070), .Z(n1421) );
  AND U2901 ( .A(\SUBBYTES[8].a/w372 ), .B(n1422), .Z(\SUBBYTES[8].a/w468 ) );
  XOR U2902 ( .A(n14795), .B(\SUBBYTES[8].a/w439 ), .Z(n1422) );
  ANDN U2903 ( .A(n1423), .B(n1427), .Z(\SUBBYTES[8].a/w467 ) );
  XOR U2904 ( .A(n1070), .B(n14795), .Z(n1423) );
  ANDN U2905 ( .A(\SUBBYTES[8].a/w373 ), .B(n1424), .Z(\SUBBYTES[8].a/w463 )
         );
  XNOR U2906 ( .A(\SUBBYTES[8].a/w432 ), .B(\SUBBYTES[8].a/w435 ), .Z(n1424)
         );
  AND U2907 ( .A(\SUBBYTES[8].a/w374 ), .B(n1425), .Z(\SUBBYTES[8].a/w461 ) );
  XNOR U2908 ( .A(n1428), .B(\SUBBYTES[8].a/w432 ), .Z(n1425) );
  AND U2909 ( .A(\SUBBYTES[8].a/w459 ), .B(n1429), .Z(\SUBBYTES[8].a/w460 ) );
  XOR U2910 ( .A(n1430), .B(n1428), .Z(n1429) );
  IV U2911 ( .A(n14794), .Z(n1428) );
  ANDN U2912 ( .A(\SUBBYTES[8].a/w478 ), .B(n1431), .Z(\SUBBYTES[8].a/w455 )
         );
  ANDN U2913 ( .A(\SUBBYTES[8].a/w479 ), .B(n1432), .Z(\SUBBYTES[8].a/w453 )
         );
  ANDN U2914 ( .A(\SUBBYTES[8].a/w482 ), .B(n1433), .Z(\SUBBYTES[8].a/w452 )
         );
  AND U2915 ( .A(\SUBBYTES[8].a/w438 ), .B(\SUBBYTES[8].a/w437 ), .Z(
        \SUBBYTES[8].a/w439 ) );
  IV U2916 ( .A(n1430), .Z(\SUBBYTES[8].a/w435 ) );
  NAND U2917 ( .A(\SUBBYTES[8].a/w414 ), .B(\SUBBYTES[8].a/w429 ), .Z(n1430)
         );
  AND U2918 ( .A(\SUBBYTES[8].a/w431 ), .B(\SUBBYTES[8].a/w437 ), .Z(
        \SUBBYTES[8].a/w432 ) );
  AND U2919 ( .A(\SUBBYTES[8].a/w416 ), .B(\SUBBYTES[8].a/w414 ), .Z(
        \SUBBYTES[8].a/w426 ) );
  AND U2920 ( .A(\SUBBYTES[8].a/w417 ), .B(\SUBBYTES[8].a/w415 ), .Z(
        \SUBBYTES[8].a/w424 ) );
  AND U2921 ( .A(\SUBBYTES[8].a/w431 ), .B(\SUBBYTES[8].a/w438 ), .Z(
        \SUBBYTES[8].a/w423 ) );
  AND U2922 ( .A(\SUBBYTES[8].a/w371 ), .B(\SUBBYTES[8].a/w367 ), .Z(
        \SUBBYTES[8].a/w408 ) );
  AND U2923 ( .A(\SUBBYTES[8].a/w372 ), .B(\SUBBYTES[8].a/w368 ), .Z(
        \SUBBYTES[8].a/w406 ) );
  ANDN U2924 ( .A(\SUBBYTES[8].a/w498 ), .B(n1427), .Z(\SUBBYTES[8].a/w405 )
         );
  XNOR U2925 ( .A(\w1[8][113] ), .B(\w1[8][119] ), .Z(n1427) );
  XOR U2926 ( .A(\w0[8][113] ), .B(g_input[1137]), .Z(\w1[8][113] ) );
  AND U2927 ( .A(\w1[8][112] ), .B(\SUBBYTES[8].a/w373 ), .Z(
        \SUBBYTES[8].a/w401 ) );
  XOR U2928 ( .A(\w0[8][112] ), .B(g_input[1136]), .Z(\w1[8][112] ) );
  AND U2929 ( .A(\SUBBYTES[8].a/w374 ), .B(\SUBBYTES[8].a/w370 ), .Z(
        \SUBBYTES[8].a/w399 ) );
  AND U2930 ( .A(\SUBBYTES[8].a/w459 ), .B(\SUBBYTES[8].a/w491 ), .Z(
        \SUBBYTES[8].a/w398 ) );
  ANDN U2931 ( .A(\SUBBYTES[8].a/w480 ), .B(n1431), .Z(\SUBBYTES[8].a/w393 )
         );
  XNOR U2932 ( .A(\w1[8][116] ), .B(\w1[8][119] ), .Z(n1431) );
  ANDN U2933 ( .A(\SUBBYTES[8].a/w481 ), .B(n1432), .Z(\SUBBYTES[8].a/w391 )
         );
  XNOR U2934 ( .A(\w1[8][114] ), .B(\w1[8][119] ), .Z(n1432) );
  XOR U2935 ( .A(\w0[8][119] ), .B(g_input[1143]), .Z(\w1[8][119] ) );
  IV U2936 ( .A(n1434), .Z(\w1[8][114] ) );
  ANDN U2937 ( .A(\SUBBYTES[8].a/w483 ), .B(n1433), .Z(\SUBBYTES[8].a/w390 )
         );
  XOR U2938 ( .A(n1434), .B(\w1[8][116] ), .Z(n1433) );
  XOR U2939 ( .A(\w0[8][116] ), .B(g_input[1140]), .Z(\w1[8][116] ) );
  XNOR U2940 ( .A(\w0[8][114] ), .B(g_input[1138]), .Z(n1434) );
  AND U2941 ( .A(n1435), .B(\SUBBYTES[8].a/w3265 ), .Z(\SUBBYTES[8].a/w3400 )
         );
  AND U2942 ( .A(n1436), .B(\SUBBYTES[8].a/w3266 ), .Z(\SUBBYTES[8].a/w3398 )
         );
  AND U2943 ( .A(\SUBBYTES[8].a/w3396 ), .B(n1437), .Z(\SUBBYTES[8].a/w3397 )
         );
  ANDN U2944 ( .A(\w1[8][0] ), .B(n1438), .Z(\SUBBYTES[8].a/w3393 ) );
  AND U2945 ( .A(n1439), .B(\SUBBYTES[8].a/w3268 ), .Z(\SUBBYTES[8].a/w3391 )
         );
  AND U2946 ( .A(\SUBBYTES[8].a/w3389 ), .B(n1440), .Z(\SUBBYTES[8].a/w3390 )
         );
  XOR U2947 ( .A(\SUBBYTES[8].a/w3333 ), .B(n14822), .Z(n1440) );
  AND U2948 ( .A(\SUBBYTES[8].a/w3376 ), .B(\SUBBYTES[8].a/w3378 ), .Z(
        \SUBBYTES[8].a/w3385 ) );
  AND U2949 ( .A(\SUBBYTES[8].a/w3377 ), .B(\SUBBYTES[8].a/w3379 ), .Z(
        \SUBBYTES[8].a/w3383 ) );
  AND U2950 ( .A(\SUBBYTES[8].a/w3380 ), .B(\SUBBYTES[8].a/w3381 ), .Z(
        \SUBBYTES[8].a/w3382 ) );
  AND U2951 ( .A(\SUBBYTES[8].a/w3269 ), .B(n1435), .Z(\SUBBYTES[8].a/w3368 )
         );
  XOR U2952 ( .A(\SUBBYTES[8].a/w3337 ), .B(n1084), .Z(n1435) );
  AND U2953 ( .A(\SUBBYTES[8].a/w3270 ), .B(n1436), .Z(\SUBBYTES[8].a/w3366 )
         );
  XOR U2954 ( .A(n14823), .B(\SUBBYTES[8].a/w3337 ), .Z(n1436) );
  ANDN U2955 ( .A(n1437), .B(n1441), .Z(\SUBBYTES[8].a/w3365 ) );
  XOR U2956 ( .A(n1084), .B(n14823), .Z(n1437) );
  ANDN U2957 ( .A(\SUBBYTES[8].a/w3271 ), .B(n1438), .Z(\SUBBYTES[8].a/w3361 )
         );
  XNOR U2958 ( .A(\SUBBYTES[8].a/w3330 ), .B(\SUBBYTES[8].a/w3333 ), .Z(n1438)
         );
  AND U2959 ( .A(\SUBBYTES[8].a/w3272 ), .B(n1439), .Z(\SUBBYTES[8].a/w3359 )
         );
  XNOR U2960 ( .A(n1442), .B(\SUBBYTES[8].a/w3330 ), .Z(n1439) );
  AND U2961 ( .A(\SUBBYTES[8].a/w3357 ), .B(n1443), .Z(\SUBBYTES[8].a/w3358 )
         );
  XOR U2962 ( .A(n1444), .B(n1442), .Z(n1443) );
  IV U2963 ( .A(n14822), .Z(n1442) );
  ANDN U2964 ( .A(\SUBBYTES[8].a/w3376 ), .B(n1445), .Z(\SUBBYTES[8].a/w3353 )
         );
  ANDN U2965 ( .A(\SUBBYTES[8].a/w3377 ), .B(n1446), .Z(\SUBBYTES[8].a/w3351 )
         );
  ANDN U2966 ( .A(\SUBBYTES[8].a/w3380 ), .B(n1447), .Z(\SUBBYTES[8].a/w3350 )
         );
  AND U2967 ( .A(\SUBBYTES[8].a/w3336 ), .B(\SUBBYTES[8].a/w3335 ), .Z(
        \SUBBYTES[8].a/w3337 ) );
  IV U2968 ( .A(n1444), .Z(\SUBBYTES[8].a/w3333 ) );
  NAND U2969 ( .A(\SUBBYTES[8].a/w3312 ), .B(\SUBBYTES[8].a/w3327 ), .Z(n1444)
         );
  AND U2970 ( .A(\SUBBYTES[8].a/w3329 ), .B(\SUBBYTES[8].a/w3335 ), .Z(
        \SUBBYTES[8].a/w3330 ) );
  AND U2971 ( .A(\SUBBYTES[8].a/w3314 ), .B(\SUBBYTES[8].a/w3312 ), .Z(
        \SUBBYTES[8].a/w3324 ) );
  AND U2972 ( .A(\SUBBYTES[8].a/w3315 ), .B(\SUBBYTES[8].a/w3313 ), .Z(
        \SUBBYTES[8].a/w3322 ) );
  AND U2973 ( .A(\SUBBYTES[8].a/w3329 ), .B(\SUBBYTES[8].a/w3336 ), .Z(
        \SUBBYTES[8].a/w3321 ) );
  AND U2974 ( .A(\SUBBYTES[8].a/w3269 ), .B(\SUBBYTES[8].a/w3265 ), .Z(
        \SUBBYTES[8].a/w3306 ) );
  AND U2975 ( .A(\SUBBYTES[8].a/w3270 ), .B(\SUBBYTES[8].a/w3266 ), .Z(
        \SUBBYTES[8].a/w3304 ) );
  ANDN U2976 ( .A(\SUBBYTES[8].a/w3396 ), .B(n1441), .Z(\SUBBYTES[8].a/w3303 )
         );
  XNOR U2977 ( .A(\w1[8][1] ), .B(\w1[8][7] ), .Z(n1441) );
  XOR U2978 ( .A(\w0[8][1] ), .B(g_input[1025]), .Z(\w1[8][1] ) );
  AND U2979 ( .A(\w1[8][0] ), .B(\SUBBYTES[8].a/w3271 ), .Z(
        \SUBBYTES[8].a/w3299 ) );
  XOR U2980 ( .A(\w0[8][0] ), .B(g_input[1024]), .Z(\w1[8][0] ) );
  AND U2981 ( .A(\SUBBYTES[8].a/w3272 ), .B(\SUBBYTES[8].a/w3268 ), .Z(
        \SUBBYTES[8].a/w3297 ) );
  AND U2982 ( .A(\SUBBYTES[8].a/w3357 ), .B(\SUBBYTES[8].a/w3389 ), .Z(
        \SUBBYTES[8].a/w3296 ) );
  ANDN U2983 ( .A(\SUBBYTES[8].a/w3378 ), .B(n1445), .Z(\SUBBYTES[8].a/w3291 )
         );
  XNOR U2984 ( .A(\w1[8][4] ), .B(\w1[8][7] ), .Z(n1445) );
  ANDN U2985 ( .A(\SUBBYTES[8].a/w3379 ), .B(n1446), .Z(\SUBBYTES[8].a/w3289 )
         );
  XNOR U2986 ( .A(\w1[8][2] ), .B(\w1[8][7] ), .Z(n1446) );
  XOR U2987 ( .A(\w0[8][7] ), .B(g_input[1031]), .Z(\w1[8][7] ) );
  IV U2988 ( .A(n1448), .Z(\w1[8][2] ) );
  ANDN U2989 ( .A(\SUBBYTES[8].a/w3381 ), .B(n1447), .Z(\SUBBYTES[8].a/w3288 )
         );
  XOR U2990 ( .A(n1448), .B(\w1[8][4] ), .Z(n1447) );
  XOR U2991 ( .A(\w0[8][4] ), .B(g_input[1028]), .Z(\w1[8][4] ) );
  XNOR U2992 ( .A(\w0[8][2] ), .B(g_input[1026]), .Z(n1448) );
  AND U2993 ( .A(n1449), .B(\SUBBYTES[8].a/w3058 ), .Z(\SUBBYTES[8].a/w3193 )
         );
  AND U2994 ( .A(n1450), .B(\SUBBYTES[8].a/w3059 ), .Z(\SUBBYTES[8].a/w3191 )
         );
  AND U2995 ( .A(\SUBBYTES[8].a/w3189 ), .B(n1451), .Z(\SUBBYTES[8].a/w3190 )
         );
  ANDN U2996 ( .A(\w1[8][8] ), .B(n1452), .Z(\SUBBYTES[8].a/w3186 ) );
  AND U2997 ( .A(n1453), .B(\SUBBYTES[8].a/w3061 ), .Z(\SUBBYTES[8].a/w3184 )
         );
  AND U2998 ( .A(\SUBBYTES[8].a/w3182 ), .B(n1454), .Z(\SUBBYTES[8].a/w3183 )
         );
  XOR U2999 ( .A(\SUBBYTES[8].a/w3126 ), .B(n14820), .Z(n1454) );
  AND U3000 ( .A(\SUBBYTES[8].a/w3169 ), .B(\SUBBYTES[8].a/w3171 ), .Z(
        \SUBBYTES[8].a/w3178 ) );
  AND U3001 ( .A(\SUBBYTES[8].a/w3170 ), .B(\SUBBYTES[8].a/w3172 ), .Z(
        \SUBBYTES[8].a/w3176 ) );
  AND U3002 ( .A(\SUBBYTES[8].a/w3173 ), .B(\SUBBYTES[8].a/w3174 ), .Z(
        \SUBBYTES[8].a/w3175 ) );
  AND U3003 ( .A(\SUBBYTES[8].a/w3062 ), .B(n1449), .Z(\SUBBYTES[8].a/w3161 )
         );
  XOR U3004 ( .A(\SUBBYTES[8].a/w3130 ), .B(n1083), .Z(n1449) );
  AND U3005 ( .A(\SUBBYTES[8].a/w3063 ), .B(n1450), .Z(\SUBBYTES[8].a/w3159 )
         );
  XOR U3006 ( .A(n14821), .B(\SUBBYTES[8].a/w3130 ), .Z(n1450) );
  ANDN U3007 ( .A(n1451), .B(n1455), .Z(\SUBBYTES[8].a/w3158 ) );
  XOR U3008 ( .A(n1083), .B(n14821), .Z(n1451) );
  ANDN U3009 ( .A(\SUBBYTES[8].a/w3064 ), .B(n1452), .Z(\SUBBYTES[8].a/w3154 )
         );
  XNOR U3010 ( .A(\SUBBYTES[8].a/w3123 ), .B(\SUBBYTES[8].a/w3126 ), .Z(n1452)
         );
  AND U3011 ( .A(\SUBBYTES[8].a/w3065 ), .B(n1453), .Z(\SUBBYTES[8].a/w3152 )
         );
  XNOR U3012 ( .A(n1456), .B(\SUBBYTES[8].a/w3123 ), .Z(n1453) );
  AND U3013 ( .A(\SUBBYTES[8].a/w3150 ), .B(n1457), .Z(\SUBBYTES[8].a/w3151 )
         );
  XOR U3014 ( .A(n1458), .B(n1456), .Z(n1457) );
  IV U3015 ( .A(n14820), .Z(n1456) );
  ANDN U3016 ( .A(\SUBBYTES[8].a/w3169 ), .B(n1459), .Z(\SUBBYTES[8].a/w3146 )
         );
  ANDN U3017 ( .A(\SUBBYTES[8].a/w3170 ), .B(n1460), .Z(\SUBBYTES[8].a/w3144 )
         );
  ANDN U3018 ( .A(\SUBBYTES[8].a/w3173 ), .B(n1461), .Z(\SUBBYTES[8].a/w3143 )
         );
  AND U3019 ( .A(\SUBBYTES[8].a/w3129 ), .B(\SUBBYTES[8].a/w3128 ), .Z(
        \SUBBYTES[8].a/w3130 ) );
  IV U3020 ( .A(n1458), .Z(\SUBBYTES[8].a/w3126 ) );
  NAND U3021 ( .A(\SUBBYTES[8].a/w3105 ), .B(\SUBBYTES[8].a/w3120 ), .Z(n1458)
         );
  AND U3022 ( .A(\SUBBYTES[8].a/w3122 ), .B(\SUBBYTES[8].a/w3128 ), .Z(
        \SUBBYTES[8].a/w3123 ) );
  AND U3023 ( .A(\SUBBYTES[8].a/w3107 ), .B(\SUBBYTES[8].a/w3105 ), .Z(
        \SUBBYTES[8].a/w3117 ) );
  AND U3024 ( .A(\SUBBYTES[8].a/w3108 ), .B(\SUBBYTES[8].a/w3106 ), .Z(
        \SUBBYTES[8].a/w3115 ) );
  AND U3025 ( .A(\SUBBYTES[8].a/w3122 ), .B(\SUBBYTES[8].a/w3129 ), .Z(
        \SUBBYTES[8].a/w3114 ) );
  AND U3026 ( .A(\SUBBYTES[8].a/w3062 ), .B(\SUBBYTES[8].a/w3058 ), .Z(
        \SUBBYTES[8].a/w3099 ) );
  AND U3027 ( .A(\SUBBYTES[8].a/w3063 ), .B(\SUBBYTES[8].a/w3059 ), .Z(
        \SUBBYTES[8].a/w3097 ) );
  ANDN U3028 ( .A(\SUBBYTES[8].a/w3189 ), .B(n1455), .Z(\SUBBYTES[8].a/w3096 )
         );
  XNOR U3029 ( .A(\w1[8][15] ), .B(\w1[8][9] ), .Z(n1455) );
  XOR U3030 ( .A(\w0[8][9] ), .B(g_input[1033]), .Z(\w1[8][9] ) );
  AND U3031 ( .A(\w1[8][8] ), .B(\SUBBYTES[8].a/w3064 ), .Z(
        \SUBBYTES[8].a/w3092 ) );
  XOR U3032 ( .A(\w0[8][8] ), .B(g_input[1032]), .Z(\w1[8][8] ) );
  AND U3033 ( .A(\SUBBYTES[8].a/w3065 ), .B(\SUBBYTES[8].a/w3061 ), .Z(
        \SUBBYTES[8].a/w3090 ) );
  AND U3034 ( .A(\SUBBYTES[8].a/w3150 ), .B(\SUBBYTES[8].a/w3182 ), .Z(
        \SUBBYTES[8].a/w3089 ) );
  ANDN U3035 ( .A(\SUBBYTES[8].a/w3171 ), .B(n1459), .Z(\SUBBYTES[8].a/w3084 )
         );
  XNOR U3036 ( .A(\w1[8][12] ), .B(\w1[8][15] ), .Z(n1459) );
  ANDN U3037 ( .A(\SUBBYTES[8].a/w3172 ), .B(n1460), .Z(\SUBBYTES[8].a/w3082 )
         );
  XNOR U3038 ( .A(\w1[8][10] ), .B(\w1[8][15] ), .Z(n1460) );
  XOR U3039 ( .A(\w0[8][15] ), .B(g_input[1039]), .Z(\w1[8][15] ) );
  ANDN U3040 ( .A(\SUBBYTES[8].a/w3174 ), .B(n1461), .Z(\SUBBYTES[8].a/w3081 )
         );
  XNOR U3041 ( .A(\w1[8][10] ), .B(\w1[8][12] ), .Z(n1461) );
  XOR U3042 ( .A(\w0[8][12] ), .B(g_input[1036]), .Z(\w1[8][12] ) );
  XOR U3043 ( .A(\w0[8][10] ), .B(g_input[1034]), .Z(\w1[8][10] ) );
  AND U3044 ( .A(n1462), .B(\SUBBYTES[8].a/w2851 ), .Z(\SUBBYTES[8].a/w2986 )
         );
  AND U3045 ( .A(n1463), .B(\SUBBYTES[8].a/w2852 ), .Z(\SUBBYTES[8].a/w2984 )
         );
  AND U3046 ( .A(\SUBBYTES[8].a/w2982 ), .B(n1464), .Z(\SUBBYTES[8].a/w2983 )
         );
  ANDN U3047 ( .A(\w1[8][16] ), .B(n1465), .Z(\SUBBYTES[8].a/w2979 ) );
  AND U3048 ( .A(n1466), .B(\SUBBYTES[8].a/w2854 ), .Z(\SUBBYTES[8].a/w2977 )
         );
  AND U3049 ( .A(\SUBBYTES[8].a/w2975 ), .B(n1467), .Z(\SUBBYTES[8].a/w2976 )
         );
  XOR U3050 ( .A(\SUBBYTES[8].a/w2919 ), .B(n14818), .Z(n1467) );
  AND U3051 ( .A(\SUBBYTES[8].a/w2962 ), .B(\SUBBYTES[8].a/w2964 ), .Z(
        \SUBBYTES[8].a/w2971 ) );
  AND U3052 ( .A(\SUBBYTES[8].a/w2963 ), .B(\SUBBYTES[8].a/w2965 ), .Z(
        \SUBBYTES[8].a/w2969 ) );
  AND U3053 ( .A(\SUBBYTES[8].a/w2966 ), .B(\SUBBYTES[8].a/w2967 ), .Z(
        \SUBBYTES[8].a/w2968 ) );
  AND U3054 ( .A(\SUBBYTES[8].a/w2855 ), .B(n1462), .Z(\SUBBYTES[8].a/w2954 )
         );
  XOR U3055 ( .A(\SUBBYTES[8].a/w2923 ), .B(n1082), .Z(n1462) );
  AND U3056 ( .A(\SUBBYTES[8].a/w2856 ), .B(n1463), .Z(\SUBBYTES[8].a/w2952 )
         );
  XOR U3057 ( .A(n14819), .B(\SUBBYTES[8].a/w2923 ), .Z(n1463) );
  ANDN U3058 ( .A(n1464), .B(n1468), .Z(\SUBBYTES[8].a/w2951 ) );
  XOR U3059 ( .A(n1082), .B(n14819), .Z(n1464) );
  AND U3060 ( .A(n1469), .B(\SUBBYTES[8].a/w160 ), .Z(\SUBBYTES[8].a/w295 ) );
  ANDN U3061 ( .A(\SUBBYTES[8].a/w2857 ), .B(n1465), .Z(\SUBBYTES[8].a/w2947 )
         );
  XNOR U3062 ( .A(\SUBBYTES[8].a/w2916 ), .B(\SUBBYTES[8].a/w2919 ), .Z(n1465)
         );
  AND U3063 ( .A(\SUBBYTES[8].a/w2858 ), .B(n1466), .Z(\SUBBYTES[8].a/w2945 )
         );
  XNOR U3064 ( .A(n1470), .B(\SUBBYTES[8].a/w2916 ), .Z(n1466) );
  AND U3065 ( .A(\SUBBYTES[8].a/w2943 ), .B(n1471), .Z(\SUBBYTES[8].a/w2944 )
         );
  XOR U3066 ( .A(n1472), .B(n1470), .Z(n1471) );
  IV U3067 ( .A(n14818), .Z(n1470) );
  ANDN U3068 ( .A(\SUBBYTES[8].a/w2962 ), .B(n1473), .Z(\SUBBYTES[8].a/w2939 )
         );
  ANDN U3069 ( .A(\SUBBYTES[8].a/w2963 ), .B(n1474), .Z(\SUBBYTES[8].a/w2937 )
         );
  ANDN U3070 ( .A(\SUBBYTES[8].a/w2966 ), .B(n1475), .Z(\SUBBYTES[8].a/w2936 )
         );
  AND U3071 ( .A(n1476), .B(\SUBBYTES[8].a/w161 ), .Z(\SUBBYTES[8].a/w293 ) );
  AND U3072 ( .A(\SUBBYTES[8].a/w2922 ), .B(\SUBBYTES[8].a/w2921 ), .Z(
        \SUBBYTES[8].a/w2923 ) );
  AND U3073 ( .A(\SUBBYTES[8].a/w291 ), .B(n1477), .Z(\SUBBYTES[8].a/w292 ) );
  IV U3074 ( .A(n1472), .Z(\SUBBYTES[8].a/w2919 ) );
  NAND U3075 ( .A(\SUBBYTES[8].a/w2898 ), .B(\SUBBYTES[8].a/w2913 ), .Z(n1472)
         );
  AND U3076 ( .A(\SUBBYTES[8].a/w2915 ), .B(\SUBBYTES[8].a/w2921 ), .Z(
        \SUBBYTES[8].a/w2916 ) );
  AND U3077 ( .A(\SUBBYTES[8].a/w2900 ), .B(\SUBBYTES[8].a/w2898 ), .Z(
        \SUBBYTES[8].a/w2910 ) );
  AND U3078 ( .A(\SUBBYTES[8].a/w2901 ), .B(\SUBBYTES[8].a/w2899 ), .Z(
        \SUBBYTES[8].a/w2908 ) );
  AND U3079 ( .A(\SUBBYTES[8].a/w2915 ), .B(\SUBBYTES[8].a/w2922 ), .Z(
        \SUBBYTES[8].a/w2907 ) );
  AND U3080 ( .A(\SUBBYTES[8].a/w2855 ), .B(\SUBBYTES[8].a/w2851 ), .Z(
        \SUBBYTES[8].a/w2892 ) );
  AND U3081 ( .A(\SUBBYTES[8].a/w2856 ), .B(\SUBBYTES[8].a/w2852 ), .Z(
        \SUBBYTES[8].a/w2890 ) );
  ANDN U3082 ( .A(\SUBBYTES[8].a/w2982 ), .B(n1468), .Z(\SUBBYTES[8].a/w2889 )
         );
  XNOR U3083 ( .A(\w1[8][17] ), .B(\w1[8][23] ), .Z(n1468) );
  XOR U3084 ( .A(\w0[8][17] ), .B(g_input[1041]), .Z(\w1[8][17] ) );
  AND U3085 ( .A(\w1[8][16] ), .B(\SUBBYTES[8].a/w2857 ), .Z(
        \SUBBYTES[8].a/w2885 ) );
  XOR U3086 ( .A(\w0[8][16] ), .B(g_input[1040]), .Z(\w1[8][16] ) );
  AND U3087 ( .A(\SUBBYTES[8].a/w2858 ), .B(\SUBBYTES[8].a/w2854 ), .Z(
        \SUBBYTES[8].a/w2883 ) );
  AND U3088 ( .A(\SUBBYTES[8].a/w2943 ), .B(\SUBBYTES[8].a/w2975 ), .Z(
        \SUBBYTES[8].a/w2882 ) );
  ANDN U3089 ( .A(\w1[8][120] ), .B(n1478), .Z(\SUBBYTES[8].a/w288 ) );
  ANDN U3090 ( .A(\SUBBYTES[8].a/w2964 ), .B(n1473), .Z(\SUBBYTES[8].a/w2877 )
         );
  XNOR U3091 ( .A(\w1[8][20] ), .B(\w1[8][23] ), .Z(n1473) );
  ANDN U3092 ( .A(\SUBBYTES[8].a/w2965 ), .B(n1474), .Z(\SUBBYTES[8].a/w2875 )
         );
  XNOR U3093 ( .A(\w1[8][18] ), .B(\w1[8][23] ), .Z(n1474) );
  XOR U3094 ( .A(\w0[8][23] ), .B(g_input[1047]), .Z(\w1[8][23] ) );
  IV U3095 ( .A(n1479), .Z(\w1[8][18] ) );
  ANDN U3096 ( .A(\SUBBYTES[8].a/w2967 ), .B(n1475), .Z(\SUBBYTES[8].a/w2874 )
         );
  XOR U3097 ( .A(n1479), .B(\w1[8][20] ), .Z(n1475) );
  XOR U3098 ( .A(\w0[8][20] ), .B(g_input[1044]), .Z(\w1[8][20] ) );
  XNOR U3099 ( .A(\w0[8][18] ), .B(g_input[1042]), .Z(n1479) );
  AND U3100 ( .A(n1480), .B(\SUBBYTES[8].a/w163 ), .Z(\SUBBYTES[8].a/w286 ) );
  AND U3101 ( .A(\SUBBYTES[8].a/w284 ), .B(n1481), .Z(\SUBBYTES[8].a/w285 ) );
  XOR U3102 ( .A(\SUBBYTES[8].a/w228 ), .B(n14792), .Z(n1481) );
  AND U3103 ( .A(\SUBBYTES[8].a/w271 ), .B(\SUBBYTES[8].a/w273 ), .Z(
        \SUBBYTES[8].a/w280 ) );
  AND U3104 ( .A(\SUBBYTES[8].a/w272 ), .B(\SUBBYTES[8].a/w274 ), .Z(
        \SUBBYTES[8].a/w278 ) );
  AND U3105 ( .A(n1482), .B(\SUBBYTES[8].a/w2644 ), .Z(\SUBBYTES[8].a/w2779 )
         );
  AND U3106 ( .A(n1483), .B(\SUBBYTES[8].a/w2645 ), .Z(\SUBBYTES[8].a/w2777 )
         );
  AND U3107 ( .A(\SUBBYTES[8].a/w2775 ), .B(n1484), .Z(\SUBBYTES[8].a/w2776 )
         );
  ANDN U3108 ( .A(\w1[8][24] ), .B(n1485), .Z(\SUBBYTES[8].a/w2772 ) );
  AND U3109 ( .A(n1486), .B(\SUBBYTES[8].a/w2647 ), .Z(\SUBBYTES[8].a/w2770 )
         );
  AND U3110 ( .A(\SUBBYTES[8].a/w275 ), .B(\SUBBYTES[8].a/w276 ), .Z(
        \SUBBYTES[8].a/w277 ) );
  AND U3111 ( .A(\SUBBYTES[8].a/w2768 ), .B(n1487), .Z(\SUBBYTES[8].a/w2769 )
         );
  XOR U3112 ( .A(\SUBBYTES[8].a/w2712 ), .B(n14816), .Z(n1487) );
  AND U3113 ( .A(\SUBBYTES[8].a/w2755 ), .B(\SUBBYTES[8].a/w2757 ), .Z(
        \SUBBYTES[8].a/w2764 ) );
  AND U3114 ( .A(\SUBBYTES[8].a/w2756 ), .B(\SUBBYTES[8].a/w2758 ), .Z(
        \SUBBYTES[8].a/w2762 ) );
  AND U3115 ( .A(\SUBBYTES[8].a/w2759 ), .B(\SUBBYTES[8].a/w2760 ), .Z(
        \SUBBYTES[8].a/w2761 ) );
  AND U3116 ( .A(\SUBBYTES[8].a/w2648 ), .B(n1482), .Z(\SUBBYTES[8].a/w2747 )
         );
  XOR U3117 ( .A(\SUBBYTES[8].a/w2716 ), .B(n1081), .Z(n1482) );
  AND U3118 ( .A(\SUBBYTES[8].a/w2649 ), .B(n1483), .Z(\SUBBYTES[8].a/w2745 )
         );
  XOR U3119 ( .A(n14817), .B(\SUBBYTES[8].a/w2716 ), .Z(n1483) );
  ANDN U3120 ( .A(n1484), .B(n1488), .Z(\SUBBYTES[8].a/w2744 ) );
  XOR U3121 ( .A(n1081), .B(n14817), .Z(n1484) );
  ANDN U3122 ( .A(\SUBBYTES[8].a/w2650 ), .B(n1485), .Z(\SUBBYTES[8].a/w2740 )
         );
  XNOR U3123 ( .A(\SUBBYTES[8].a/w2709 ), .B(\SUBBYTES[8].a/w2712 ), .Z(n1485)
         );
  AND U3124 ( .A(\SUBBYTES[8].a/w2651 ), .B(n1486), .Z(\SUBBYTES[8].a/w2738 )
         );
  XNOR U3125 ( .A(n1489), .B(\SUBBYTES[8].a/w2709 ), .Z(n1486) );
  AND U3126 ( .A(\SUBBYTES[8].a/w2736 ), .B(n1490), .Z(\SUBBYTES[8].a/w2737 )
         );
  XOR U3127 ( .A(n1491), .B(n1489), .Z(n1490) );
  IV U3128 ( .A(n14816), .Z(n1489) );
  ANDN U3129 ( .A(\SUBBYTES[8].a/w2755 ), .B(n1492), .Z(\SUBBYTES[8].a/w2732 )
         );
  ANDN U3130 ( .A(\SUBBYTES[8].a/w2756 ), .B(n1493), .Z(\SUBBYTES[8].a/w2730 )
         );
  ANDN U3131 ( .A(\SUBBYTES[8].a/w2759 ), .B(n1494), .Z(\SUBBYTES[8].a/w2729 )
         );
  AND U3132 ( .A(\SUBBYTES[8].a/w2715 ), .B(\SUBBYTES[8].a/w2714 ), .Z(
        \SUBBYTES[8].a/w2716 ) );
  IV U3133 ( .A(n1491), .Z(\SUBBYTES[8].a/w2712 ) );
  NAND U3134 ( .A(\SUBBYTES[8].a/w2691 ), .B(\SUBBYTES[8].a/w2706 ), .Z(n1491)
         );
  AND U3135 ( .A(\SUBBYTES[8].a/w2708 ), .B(\SUBBYTES[8].a/w2714 ), .Z(
        \SUBBYTES[8].a/w2709 ) );
  AND U3136 ( .A(\SUBBYTES[8].a/w2693 ), .B(\SUBBYTES[8].a/w2691 ), .Z(
        \SUBBYTES[8].a/w2703 ) );
  AND U3137 ( .A(\SUBBYTES[8].a/w2694 ), .B(\SUBBYTES[8].a/w2692 ), .Z(
        \SUBBYTES[8].a/w2701 ) );
  AND U3138 ( .A(\SUBBYTES[8].a/w2708 ), .B(\SUBBYTES[8].a/w2715 ), .Z(
        \SUBBYTES[8].a/w2700 ) );
  AND U3139 ( .A(\SUBBYTES[8].a/w2648 ), .B(\SUBBYTES[8].a/w2644 ), .Z(
        \SUBBYTES[8].a/w2685 ) );
  AND U3140 ( .A(\SUBBYTES[8].a/w2649 ), .B(\SUBBYTES[8].a/w2645 ), .Z(
        \SUBBYTES[8].a/w2683 ) );
  ANDN U3141 ( .A(\SUBBYTES[8].a/w2775 ), .B(n1488), .Z(\SUBBYTES[8].a/w2682 )
         );
  XNOR U3142 ( .A(\w1[8][25] ), .B(\w1[8][31] ), .Z(n1488) );
  XOR U3143 ( .A(\w0[8][25] ), .B(g_input[1049]), .Z(\w1[8][25] ) );
  AND U3144 ( .A(\w1[8][24] ), .B(\SUBBYTES[8].a/w2650 ), .Z(
        \SUBBYTES[8].a/w2678 ) );
  XOR U3145 ( .A(\w0[8][24] ), .B(g_input[1048]), .Z(\w1[8][24] ) );
  AND U3146 ( .A(\SUBBYTES[8].a/w2651 ), .B(\SUBBYTES[8].a/w2647 ), .Z(
        \SUBBYTES[8].a/w2676 ) );
  AND U3147 ( .A(\SUBBYTES[8].a/w2736 ), .B(\SUBBYTES[8].a/w2768 ), .Z(
        \SUBBYTES[8].a/w2675 ) );
  ANDN U3148 ( .A(\SUBBYTES[8].a/w2757 ), .B(n1492), .Z(\SUBBYTES[8].a/w2670 )
         );
  XNOR U3149 ( .A(\w1[8][28] ), .B(\w1[8][31] ), .Z(n1492) );
  ANDN U3150 ( .A(\SUBBYTES[8].a/w2758 ), .B(n1493), .Z(\SUBBYTES[8].a/w2668 )
         );
  XNOR U3151 ( .A(\w1[8][26] ), .B(\w1[8][31] ), .Z(n1493) );
  XOR U3152 ( .A(\w0[8][31] ), .B(g_input[1055]), .Z(\w1[8][31] ) );
  IV U3153 ( .A(n1495), .Z(\w1[8][26] ) );
  ANDN U3154 ( .A(\SUBBYTES[8].a/w2760 ), .B(n1494), .Z(\SUBBYTES[8].a/w2667 )
         );
  XOR U3155 ( .A(n1495), .B(\w1[8][28] ), .Z(n1494) );
  XOR U3156 ( .A(\w0[8][28] ), .B(g_input[1052]), .Z(\w1[8][28] ) );
  XNOR U3157 ( .A(\w0[8][26] ), .B(g_input[1050]), .Z(n1495) );
  AND U3158 ( .A(\SUBBYTES[8].a/w164 ), .B(n1469), .Z(\SUBBYTES[8].a/w263 ) );
  XOR U3159 ( .A(\SUBBYTES[8].a/w232 ), .B(n1069), .Z(n1469) );
  AND U3160 ( .A(\SUBBYTES[8].a/w165 ), .B(n1476), .Z(\SUBBYTES[8].a/w261 ) );
  XOR U3161 ( .A(n14793), .B(\SUBBYTES[8].a/w232 ), .Z(n1476) );
  ANDN U3162 ( .A(n1477), .B(n1496), .Z(\SUBBYTES[8].a/w260 ) );
  XOR U3163 ( .A(n1069), .B(n14793), .Z(n1477) );
  AND U3164 ( .A(n1497), .B(\SUBBYTES[8].a/w2437 ), .Z(\SUBBYTES[8].a/w2572 )
         );
  AND U3165 ( .A(n1498), .B(\SUBBYTES[8].a/w2438 ), .Z(\SUBBYTES[8].a/w2570 )
         );
  AND U3166 ( .A(\SUBBYTES[8].a/w2568 ), .B(n1499), .Z(\SUBBYTES[8].a/w2569 )
         );
  ANDN U3167 ( .A(\w1[8][32] ), .B(n1500), .Z(\SUBBYTES[8].a/w2565 ) );
  AND U3168 ( .A(n1501), .B(\SUBBYTES[8].a/w2440 ), .Z(\SUBBYTES[8].a/w2563 )
         );
  AND U3169 ( .A(\SUBBYTES[8].a/w2561 ), .B(n1502), .Z(\SUBBYTES[8].a/w2562 )
         );
  XOR U3170 ( .A(\SUBBYTES[8].a/w2505 ), .B(n14814), .Z(n1502) );
  ANDN U3171 ( .A(\SUBBYTES[8].a/w166 ), .B(n1478), .Z(\SUBBYTES[8].a/w256 )
         );
  XNOR U3172 ( .A(\SUBBYTES[8].a/w225 ), .B(\SUBBYTES[8].a/w228 ), .Z(n1478)
         );
  AND U3173 ( .A(\SUBBYTES[8].a/w2548 ), .B(\SUBBYTES[8].a/w2550 ), .Z(
        \SUBBYTES[8].a/w2557 ) );
  AND U3174 ( .A(\SUBBYTES[8].a/w2549 ), .B(\SUBBYTES[8].a/w2551 ), .Z(
        \SUBBYTES[8].a/w2555 ) );
  AND U3175 ( .A(\SUBBYTES[8].a/w2552 ), .B(\SUBBYTES[8].a/w2553 ), .Z(
        \SUBBYTES[8].a/w2554 ) );
  AND U3176 ( .A(\SUBBYTES[8].a/w2441 ), .B(n1497), .Z(\SUBBYTES[8].a/w2540 )
         );
  XOR U3177 ( .A(\SUBBYTES[8].a/w2509 ), .B(n1080), .Z(n1497) );
  AND U3178 ( .A(\SUBBYTES[8].a/w167 ), .B(n1480), .Z(\SUBBYTES[8].a/w254 ) );
  XNOR U3179 ( .A(n1503), .B(\SUBBYTES[8].a/w225 ), .Z(n1480) );
  AND U3180 ( .A(\SUBBYTES[8].a/w2442 ), .B(n1498), .Z(\SUBBYTES[8].a/w2538 )
         );
  XOR U3181 ( .A(n14815), .B(\SUBBYTES[8].a/w2509 ), .Z(n1498) );
  ANDN U3182 ( .A(n1499), .B(n1504), .Z(\SUBBYTES[8].a/w2537 ) );
  XOR U3183 ( .A(n1080), .B(n14815), .Z(n1499) );
  ANDN U3184 ( .A(\SUBBYTES[8].a/w2443 ), .B(n1500), .Z(\SUBBYTES[8].a/w2533 )
         );
  XNOR U3185 ( .A(\SUBBYTES[8].a/w2502 ), .B(\SUBBYTES[8].a/w2505 ), .Z(n1500)
         );
  AND U3186 ( .A(\SUBBYTES[8].a/w2444 ), .B(n1501), .Z(\SUBBYTES[8].a/w2531 )
         );
  XNOR U3187 ( .A(n1505), .B(\SUBBYTES[8].a/w2502 ), .Z(n1501) );
  AND U3188 ( .A(\SUBBYTES[8].a/w2529 ), .B(n1506), .Z(\SUBBYTES[8].a/w2530 )
         );
  XOR U3189 ( .A(n1507), .B(n1505), .Z(n1506) );
  IV U3190 ( .A(n14814), .Z(n1505) );
  AND U3191 ( .A(\SUBBYTES[8].a/w252 ), .B(n1508), .Z(\SUBBYTES[8].a/w253 ) );
  XOR U3192 ( .A(n1509), .B(n1503), .Z(n1508) );
  IV U3193 ( .A(n14792), .Z(n1503) );
  ANDN U3194 ( .A(\SUBBYTES[8].a/w2548 ), .B(n1510), .Z(\SUBBYTES[8].a/w2525 )
         );
  ANDN U3195 ( .A(\SUBBYTES[8].a/w2549 ), .B(n1511), .Z(\SUBBYTES[8].a/w2523 )
         );
  ANDN U3196 ( .A(\SUBBYTES[8].a/w2552 ), .B(n1512), .Z(\SUBBYTES[8].a/w2522 )
         );
  AND U3197 ( .A(\SUBBYTES[8].a/w2508 ), .B(\SUBBYTES[8].a/w2507 ), .Z(
        \SUBBYTES[8].a/w2509 ) );
  IV U3198 ( .A(n1507), .Z(\SUBBYTES[8].a/w2505 ) );
  NAND U3199 ( .A(\SUBBYTES[8].a/w2484 ), .B(\SUBBYTES[8].a/w2499 ), .Z(n1507)
         );
  AND U3200 ( .A(\SUBBYTES[8].a/w2501 ), .B(\SUBBYTES[8].a/w2507 ), .Z(
        \SUBBYTES[8].a/w2502 ) );
  AND U3201 ( .A(\SUBBYTES[8].a/w2486 ), .B(\SUBBYTES[8].a/w2484 ), .Z(
        \SUBBYTES[8].a/w2496 ) );
  AND U3202 ( .A(\SUBBYTES[8].a/w2487 ), .B(\SUBBYTES[8].a/w2485 ), .Z(
        \SUBBYTES[8].a/w2494 ) );
  AND U3203 ( .A(\SUBBYTES[8].a/w2501 ), .B(\SUBBYTES[8].a/w2508 ), .Z(
        \SUBBYTES[8].a/w2493 ) );
  ANDN U3204 ( .A(\SUBBYTES[8].a/w271 ), .B(n1513), .Z(\SUBBYTES[8].a/w248 )
         );
  AND U3205 ( .A(\SUBBYTES[8].a/w2441 ), .B(\SUBBYTES[8].a/w2437 ), .Z(
        \SUBBYTES[8].a/w2478 ) );
  AND U3206 ( .A(\SUBBYTES[8].a/w2442 ), .B(\SUBBYTES[8].a/w2438 ), .Z(
        \SUBBYTES[8].a/w2476 ) );
  ANDN U3207 ( .A(\SUBBYTES[8].a/w2568 ), .B(n1504), .Z(\SUBBYTES[8].a/w2475 )
         );
  XNOR U3208 ( .A(\w1[8][33] ), .B(\w1[8][39] ), .Z(n1504) );
  XOR U3209 ( .A(\w0[8][33] ), .B(g_input[1057]), .Z(\w1[8][33] ) );
  AND U3210 ( .A(\w1[8][32] ), .B(\SUBBYTES[8].a/w2443 ), .Z(
        \SUBBYTES[8].a/w2471 ) );
  XOR U3211 ( .A(\w0[8][32] ), .B(g_input[1056]), .Z(\w1[8][32] ) );
  AND U3212 ( .A(\SUBBYTES[8].a/w2444 ), .B(\SUBBYTES[8].a/w2440 ), .Z(
        \SUBBYTES[8].a/w2469 ) );
  AND U3213 ( .A(\SUBBYTES[8].a/w2529 ), .B(\SUBBYTES[8].a/w2561 ), .Z(
        \SUBBYTES[8].a/w2468 ) );
  ANDN U3214 ( .A(\SUBBYTES[8].a/w2550 ), .B(n1510), .Z(\SUBBYTES[8].a/w2463 )
         );
  XNOR U3215 ( .A(\w1[8][36] ), .B(\w1[8][39] ), .Z(n1510) );
  ANDN U3216 ( .A(\SUBBYTES[8].a/w2551 ), .B(n1511), .Z(\SUBBYTES[8].a/w2461 )
         );
  XNOR U3217 ( .A(\w1[8][34] ), .B(\w1[8][39] ), .Z(n1511) );
  XOR U3218 ( .A(\w0[8][39] ), .B(g_input[1063]), .Z(\w1[8][39] ) );
  IV U3219 ( .A(n1514), .Z(\w1[8][34] ) );
  ANDN U3220 ( .A(\SUBBYTES[8].a/w2553 ), .B(n1512), .Z(\SUBBYTES[8].a/w2460 )
         );
  XOR U3221 ( .A(n1514), .B(\w1[8][36] ), .Z(n1512) );
  XOR U3222 ( .A(\w0[8][36] ), .B(g_input[1060]), .Z(\w1[8][36] ) );
  XNOR U3223 ( .A(\w0[8][34] ), .B(g_input[1058]), .Z(n1514) );
  ANDN U3224 ( .A(\SUBBYTES[8].a/w272 ), .B(n1515), .Z(\SUBBYTES[8].a/w246 )
         );
  ANDN U3225 ( .A(\SUBBYTES[8].a/w275 ), .B(n1516), .Z(\SUBBYTES[8].a/w245 )
         );
  AND U3226 ( .A(n1517), .B(\SUBBYTES[8].a/w2230 ), .Z(\SUBBYTES[8].a/w2365 )
         );
  AND U3227 ( .A(n1518), .B(\SUBBYTES[8].a/w2231 ), .Z(\SUBBYTES[8].a/w2363 )
         );
  AND U3228 ( .A(\SUBBYTES[8].a/w2361 ), .B(n1519), .Z(\SUBBYTES[8].a/w2362 )
         );
  ANDN U3229 ( .A(\w1[8][40] ), .B(n1520), .Z(\SUBBYTES[8].a/w2358 ) );
  AND U3230 ( .A(n1521), .B(\SUBBYTES[8].a/w2233 ), .Z(\SUBBYTES[8].a/w2356 )
         );
  AND U3231 ( .A(\SUBBYTES[8].a/w2354 ), .B(n1522), .Z(\SUBBYTES[8].a/w2355 )
         );
  XOR U3232 ( .A(\SUBBYTES[8].a/w2298 ), .B(n14812), .Z(n1522) );
  AND U3233 ( .A(\SUBBYTES[8].a/w2341 ), .B(\SUBBYTES[8].a/w2343 ), .Z(
        \SUBBYTES[8].a/w2350 ) );
  AND U3234 ( .A(\SUBBYTES[8].a/w2342 ), .B(\SUBBYTES[8].a/w2344 ), .Z(
        \SUBBYTES[8].a/w2348 ) );
  AND U3235 ( .A(\SUBBYTES[8].a/w2345 ), .B(\SUBBYTES[8].a/w2346 ), .Z(
        \SUBBYTES[8].a/w2347 ) );
  AND U3236 ( .A(\SUBBYTES[8].a/w2234 ), .B(n1517), .Z(\SUBBYTES[8].a/w2333 )
         );
  XOR U3237 ( .A(\SUBBYTES[8].a/w2302 ), .B(n1079), .Z(n1517) );
  AND U3238 ( .A(\SUBBYTES[8].a/w2235 ), .B(n1518), .Z(\SUBBYTES[8].a/w2331 )
         );
  XOR U3239 ( .A(n14813), .B(\SUBBYTES[8].a/w2302 ), .Z(n1518) );
  ANDN U3240 ( .A(n1519), .B(n1523), .Z(\SUBBYTES[8].a/w2330 ) );
  XOR U3241 ( .A(n1079), .B(n14813), .Z(n1519) );
  ANDN U3242 ( .A(\SUBBYTES[8].a/w2236 ), .B(n1520), .Z(\SUBBYTES[8].a/w2326 )
         );
  XNOR U3243 ( .A(\SUBBYTES[8].a/w2295 ), .B(\SUBBYTES[8].a/w2298 ), .Z(n1520)
         );
  AND U3244 ( .A(\SUBBYTES[8].a/w2237 ), .B(n1521), .Z(\SUBBYTES[8].a/w2324 )
         );
  XNOR U3245 ( .A(n1524), .B(\SUBBYTES[8].a/w2295 ), .Z(n1521) );
  AND U3246 ( .A(\SUBBYTES[8].a/w2322 ), .B(n1525), .Z(\SUBBYTES[8].a/w2323 )
         );
  XOR U3247 ( .A(n1526), .B(n1524), .Z(n1525) );
  IV U3248 ( .A(n14812), .Z(n1524) );
  AND U3249 ( .A(\SUBBYTES[8].a/w231 ), .B(\SUBBYTES[8].a/w230 ), .Z(
        \SUBBYTES[8].a/w232 ) );
  ANDN U3250 ( .A(\SUBBYTES[8].a/w2341 ), .B(n1527), .Z(\SUBBYTES[8].a/w2318 )
         );
  ANDN U3251 ( .A(\SUBBYTES[8].a/w2342 ), .B(n1528), .Z(\SUBBYTES[8].a/w2316 )
         );
  ANDN U3252 ( .A(\SUBBYTES[8].a/w2345 ), .B(n1529), .Z(\SUBBYTES[8].a/w2315 )
         );
  AND U3253 ( .A(\SUBBYTES[8].a/w2301 ), .B(\SUBBYTES[8].a/w2300 ), .Z(
        \SUBBYTES[8].a/w2302 ) );
  IV U3254 ( .A(n1526), .Z(\SUBBYTES[8].a/w2298 ) );
  NAND U3255 ( .A(\SUBBYTES[8].a/w2277 ), .B(\SUBBYTES[8].a/w2292 ), .Z(n1526)
         );
  AND U3256 ( .A(\SUBBYTES[8].a/w2294 ), .B(\SUBBYTES[8].a/w2300 ), .Z(
        \SUBBYTES[8].a/w2295 ) );
  AND U3257 ( .A(\SUBBYTES[8].a/w2279 ), .B(\SUBBYTES[8].a/w2277 ), .Z(
        \SUBBYTES[8].a/w2289 ) );
  AND U3258 ( .A(\SUBBYTES[8].a/w2280 ), .B(\SUBBYTES[8].a/w2278 ), .Z(
        \SUBBYTES[8].a/w2287 ) );
  AND U3259 ( .A(\SUBBYTES[8].a/w2294 ), .B(\SUBBYTES[8].a/w2301 ), .Z(
        \SUBBYTES[8].a/w2286 ) );
  IV U3260 ( .A(n1509), .Z(\SUBBYTES[8].a/w228 ) );
  NAND U3261 ( .A(\SUBBYTES[8].a/w207 ), .B(\SUBBYTES[8].a/w222 ), .Z(n1509)
         );
  AND U3262 ( .A(\SUBBYTES[8].a/w2234 ), .B(\SUBBYTES[8].a/w2230 ), .Z(
        \SUBBYTES[8].a/w2271 ) );
  AND U3263 ( .A(\SUBBYTES[8].a/w2235 ), .B(\SUBBYTES[8].a/w2231 ), .Z(
        \SUBBYTES[8].a/w2269 ) );
  ANDN U3264 ( .A(\SUBBYTES[8].a/w2361 ), .B(n1523), .Z(\SUBBYTES[8].a/w2268 )
         );
  XNOR U3265 ( .A(\w1[8][41] ), .B(\w1[8][47] ), .Z(n1523) );
  XOR U3266 ( .A(\w0[8][41] ), .B(g_input[1065]), .Z(\w1[8][41] ) );
  AND U3267 ( .A(\w1[8][40] ), .B(\SUBBYTES[8].a/w2236 ), .Z(
        \SUBBYTES[8].a/w2264 ) );
  XOR U3268 ( .A(\w0[8][40] ), .B(g_input[1064]), .Z(\w1[8][40] ) );
  AND U3269 ( .A(\SUBBYTES[8].a/w2237 ), .B(\SUBBYTES[8].a/w2233 ), .Z(
        \SUBBYTES[8].a/w2262 ) );
  AND U3270 ( .A(\SUBBYTES[8].a/w2322 ), .B(\SUBBYTES[8].a/w2354 ), .Z(
        \SUBBYTES[8].a/w2261 ) );
  ANDN U3271 ( .A(\SUBBYTES[8].a/w2343 ), .B(n1527), .Z(\SUBBYTES[8].a/w2256 )
         );
  XNOR U3272 ( .A(\w1[8][44] ), .B(\w1[8][47] ), .Z(n1527) );
  ANDN U3273 ( .A(\SUBBYTES[8].a/w2344 ), .B(n1528), .Z(\SUBBYTES[8].a/w2254 )
         );
  XNOR U3274 ( .A(\w1[8][42] ), .B(\w1[8][47] ), .Z(n1528) );
  XOR U3275 ( .A(\w0[8][47] ), .B(g_input[1071]), .Z(\w1[8][47] ) );
  IV U3276 ( .A(n1530), .Z(\w1[8][42] ) );
  ANDN U3277 ( .A(\SUBBYTES[8].a/w2346 ), .B(n1529), .Z(\SUBBYTES[8].a/w2253 )
         );
  XOR U3278 ( .A(n1530), .B(\w1[8][44] ), .Z(n1529) );
  XOR U3279 ( .A(\w0[8][44] ), .B(g_input[1068]), .Z(\w1[8][44] ) );
  XNOR U3280 ( .A(\w0[8][42] ), .B(g_input[1066]), .Z(n1530) );
  AND U3281 ( .A(\SUBBYTES[8].a/w224 ), .B(\SUBBYTES[8].a/w230 ), .Z(
        \SUBBYTES[8].a/w225 ) );
  AND U3282 ( .A(\SUBBYTES[8].a/w209 ), .B(\SUBBYTES[8].a/w207 ), .Z(
        \SUBBYTES[8].a/w219 ) );
  AND U3283 ( .A(\SUBBYTES[8].a/w210 ), .B(\SUBBYTES[8].a/w208 ), .Z(
        \SUBBYTES[8].a/w217 ) );
  AND U3284 ( .A(\SUBBYTES[8].a/w224 ), .B(\SUBBYTES[8].a/w231 ), .Z(
        \SUBBYTES[8].a/w216 ) );
  AND U3285 ( .A(n1531), .B(\SUBBYTES[8].a/w2023 ), .Z(\SUBBYTES[8].a/w2158 )
         );
  AND U3286 ( .A(n1532), .B(\SUBBYTES[8].a/w2024 ), .Z(\SUBBYTES[8].a/w2156 )
         );
  AND U3287 ( .A(\SUBBYTES[8].a/w2154 ), .B(n1533), .Z(\SUBBYTES[8].a/w2155 )
         );
  ANDN U3288 ( .A(\w1[8][48] ), .B(n1534), .Z(\SUBBYTES[8].a/w2151 ) );
  AND U3289 ( .A(n1535), .B(\SUBBYTES[8].a/w2026 ), .Z(\SUBBYTES[8].a/w2149 )
         );
  AND U3290 ( .A(\SUBBYTES[8].a/w2147 ), .B(n1536), .Z(\SUBBYTES[8].a/w2148 )
         );
  XOR U3291 ( .A(\SUBBYTES[8].a/w2091 ), .B(n14810), .Z(n1536) );
  AND U3292 ( .A(\SUBBYTES[8].a/w2134 ), .B(\SUBBYTES[8].a/w2136 ), .Z(
        \SUBBYTES[8].a/w2143 ) );
  AND U3293 ( .A(\SUBBYTES[8].a/w2135 ), .B(\SUBBYTES[8].a/w2137 ), .Z(
        \SUBBYTES[8].a/w2141 ) );
  AND U3294 ( .A(\SUBBYTES[8].a/w2138 ), .B(\SUBBYTES[8].a/w2139 ), .Z(
        \SUBBYTES[8].a/w2140 ) );
  AND U3295 ( .A(\SUBBYTES[8].a/w2027 ), .B(n1531), .Z(\SUBBYTES[8].a/w2126 )
         );
  XOR U3296 ( .A(\SUBBYTES[8].a/w2095 ), .B(n1078), .Z(n1531) );
  AND U3297 ( .A(\SUBBYTES[8].a/w2028 ), .B(n1532), .Z(\SUBBYTES[8].a/w2124 )
         );
  XOR U3298 ( .A(n14811), .B(\SUBBYTES[8].a/w2095 ), .Z(n1532) );
  ANDN U3299 ( .A(n1533), .B(n1537), .Z(\SUBBYTES[8].a/w2123 ) );
  XOR U3300 ( .A(n1078), .B(n14811), .Z(n1533) );
  ANDN U3301 ( .A(\SUBBYTES[8].a/w2029 ), .B(n1534), .Z(\SUBBYTES[8].a/w2119 )
         );
  XNOR U3302 ( .A(\SUBBYTES[8].a/w2088 ), .B(\SUBBYTES[8].a/w2091 ), .Z(n1534)
         );
  AND U3303 ( .A(\SUBBYTES[8].a/w2030 ), .B(n1535), .Z(\SUBBYTES[8].a/w2117 )
         );
  XNOR U3304 ( .A(n1538), .B(\SUBBYTES[8].a/w2088 ), .Z(n1535) );
  AND U3305 ( .A(\SUBBYTES[8].a/w2115 ), .B(n1539), .Z(\SUBBYTES[8].a/w2116 )
         );
  XOR U3306 ( .A(n1540), .B(n1538), .Z(n1539) );
  IV U3307 ( .A(n14810), .Z(n1538) );
  ANDN U3308 ( .A(\SUBBYTES[8].a/w2134 ), .B(n1541), .Z(\SUBBYTES[8].a/w2111 )
         );
  ANDN U3309 ( .A(\SUBBYTES[8].a/w2135 ), .B(n1542), .Z(\SUBBYTES[8].a/w2109 )
         );
  ANDN U3310 ( .A(\SUBBYTES[8].a/w2138 ), .B(n1543), .Z(\SUBBYTES[8].a/w2108 )
         );
  AND U3311 ( .A(\SUBBYTES[8].a/w2094 ), .B(\SUBBYTES[8].a/w2093 ), .Z(
        \SUBBYTES[8].a/w2095 ) );
  IV U3312 ( .A(n1540), .Z(\SUBBYTES[8].a/w2091 ) );
  NAND U3313 ( .A(\SUBBYTES[8].a/w2070 ), .B(\SUBBYTES[8].a/w2085 ), .Z(n1540)
         );
  AND U3314 ( .A(\SUBBYTES[8].a/w2087 ), .B(\SUBBYTES[8].a/w2093 ), .Z(
        \SUBBYTES[8].a/w2088 ) );
  AND U3315 ( .A(\SUBBYTES[8].a/w2072 ), .B(\SUBBYTES[8].a/w2070 ), .Z(
        \SUBBYTES[8].a/w2082 ) );
  AND U3316 ( .A(\SUBBYTES[8].a/w2073 ), .B(\SUBBYTES[8].a/w2071 ), .Z(
        \SUBBYTES[8].a/w2080 ) );
  AND U3317 ( .A(\SUBBYTES[8].a/w2087 ), .B(\SUBBYTES[8].a/w2094 ), .Z(
        \SUBBYTES[8].a/w2079 ) );
  AND U3318 ( .A(\SUBBYTES[8].a/w2027 ), .B(\SUBBYTES[8].a/w2023 ), .Z(
        \SUBBYTES[8].a/w2064 ) );
  AND U3319 ( .A(\SUBBYTES[8].a/w2028 ), .B(\SUBBYTES[8].a/w2024 ), .Z(
        \SUBBYTES[8].a/w2062 ) );
  ANDN U3320 ( .A(\SUBBYTES[8].a/w2154 ), .B(n1537), .Z(\SUBBYTES[8].a/w2061 )
         );
  XNOR U3321 ( .A(\w1[8][49] ), .B(\w1[8][55] ), .Z(n1537) );
  XOR U3322 ( .A(\w0[8][49] ), .B(g_input[1073]), .Z(\w1[8][49] ) );
  AND U3323 ( .A(\w1[8][48] ), .B(\SUBBYTES[8].a/w2029 ), .Z(
        \SUBBYTES[8].a/w2057 ) );
  XOR U3324 ( .A(\w0[8][48] ), .B(g_input[1072]), .Z(\w1[8][48] ) );
  AND U3325 ( .A(\SUBBYTES[8].a/w2030 ), .B(\SUBBYTES[8].a/w2026 ), .Z(
        \SUBBYTES[8].a/w2055 ) );
  AND U3326 ( .A(\SUBBYTES[8].a/w2115 ), .B(\SUBBYTES[8].a/w2147 ), .Z(
        \SUBBYTES[8].a/w2054 ) );
  ANDN U3327 ( .A(\SUBBYTES[8].a/w2136 ), .B(n1541), .Z(\SUBBYTES[8].a/w2049 )
         );
  XNOR U3328 ( .A(\w1[8][52] ), .B(\w1[8][55] ), .Z(n1541) );
  ANDN U3329 ( .A(\SUBBYTES[8].a/w2137 ), .B(n1542), .Z(\SUBBYTES[8].a/w2047 )
         );
  XNOR U3330 ( .A(\w1[8][50] ), .B(\w1[8][55] ), .Z(n1542) );
  XOR U3331 ( .A(\w0[8][55] ), .B(g_input[1079]), .Z(\w1[8][55] ) );
  IV U3332 ( .A(n1544), .Z(\w1[8][50] ) );
  ANDN U3333 ( .A(\SUBBYTES[8].a/w2139 ), .B(n1543), .Z(\SUBBYTES[8].a/w2046 )
         );
  XOR U3334 ( .A(n1544), .B(\w1[8][52] ), .Z(n1543) );
  XOR U3335 ( .A(\w0[8][52] ), .B(g_input[1076]), .Z(\w1[8][52] ) );
  XNOR U3336 ( .A(\w0[8][50] ), .B(g_input[1074]), .Z(n1544) );
  AND U3337 ( .A(\SUBBYTES[8].a/w164 ), .B(\SUBBYTES[8].a/w160 ), .Z(
        \SUBBYTES[8].a/w201 ) );
  AND U3338 ( .A(\SUBBYTES[8].a/w165 ), .B(\SUBBYTES[8].a/w161 ), .Z(
        \SUBBYTES[8].a/w199 ) );
  ANDN U3339 ( .A(\SUBBYTES[8].a/w291 ), .B(n1496), .Z(\SUBBYTES[8].a/w198 )
         );
  XNOR U3340 ( .A(\w1[8][121] ), .B(\w1[8][127] ), .Z(n1496) );
  XOR U3341 ( .A(\w0[8][121] ), .B(g_input[1145]), .Z(\w1[8][121] ) );
  AND U3342 ( .A(n1545), .B(\SUBBYTES[8].a/w1816 ), .Z(\SUBBYTES[8].a/w1951 )
         );
  AND U3343 ( .A(n1546), .B(\SUBBYTES[8].a/w1817 ), .Z(\SUBBYTES[8].a/w1949 )
         );
  AND U3344 ( .A(\SUBBYTES[8].a/w1947 ), .B(n1547), .Z(\SUBBYTES[8].a/w1948 )
         );
  ANDN U3345 ( .A(\w1[8][56] ), .B(n1548), .Z(\SUBBYTES[8].a/w1944 ) );
  AND U3346 ( .A(n1549), .B(\SUBBYTES[8].a/w1819 ), .Z(\SUBBYTES[8].a/w1942 )
         );
  AND U3347 ( .A(\SUBBYTES[8].a/w1940 ), .B(n1550), .Z(\SUBBYTES[8].a/w1941 )
         );
  XOR U3348 ( .A(\SUBBYTES[8].a/w1884 ), .B(n14808), .Z(n1550) );
  AND U3349 ( .A(\w1[8][120] ), .B(\SUBBYTES[8].a/w166 ), .Z(
        \SUBBYTES[8].a/w194 ) );
  XOR U3350 ( .A(\w0[8][120] ), .B(g_input[1144]), .Z(\w1[8][120] ) );
  AND U3351 ( .A(\SUBBYTES[8].a/w1927 ), .B(\SUBBYTES[8].a/w1929 ), .Z(
        \SUBBYTES[8].a/w1936 ) );
  AND U3352 ( .A(\SUBBYTES[8].a/w1928 ), .B(\SUBBYTES[8].a/w1930 ), .Z(
        \SUBBYTES[8].a/w1934 ) );
  AND U3353 ( .A(\SUBBYTES[8].a/w1931 ), .B(\SUBBYTES[8].a/w1932 ), .Z(
        \SUBBYTES[8].a/w1933 ) );
  AND U3354 ( .A(\SUBBYTES[8].a/w167 ), .B(\SUBBYTES[8].a/w163 ), .Z(
        \SUBBYTES[8].a/w192 ) );
  AND U3355 ( .A(\SUBBYTES[8].a/w1820 ), .B(n1545), .Z(\SUBBYTES[8].a/w1919 )
         );
  XOR U3356 ( .A(\SUBBYTES[8].a/w1888 ), .B(n1077), .Z(n1545) );
  AND U3357 ( .A(\SUBBYTES[8].a/w1821 ), .B(n1546), .Z(\SUBBYTES[8].a/w1917 )
         );
  XOR U3358 ( .A(n14809), .B(\SUBBYTES[8].a/w1888 ), .Z(n1546) );
  ANDN U3359 ( .A(n1547), .B(n1551), .Z(\SUBBYTES[8].a/w1916 ) );
  XOR U3360 ( .A(n1077), .B(n14809), .Z(n1547) );
  ANDN U3361 ( .A(\SUBBYTES[8].a/w1822 ), .B(n1548), .Z(\SUBBYTES[8].a/w1912 )
         );
  XNOR U3362 ( .A(\SUBBYTES[8].a/w1881 ), .B(\SUBBYTES[8].a/w1884 ), .Z(n1548)
         );
  AND U3363 ( .A(\SUBBYTES[8].a/w1823 ), .B(n1549), .Z(\SUBBYTES[8].a/w1910 )
         );
  XNOR U3364 ( .A(n1552), .B(\SUBBYTES[8].a/w1881 ), .Z(n1549) );
  AND U3365 ( .A(\SUBBYTES[8].a/w252 ), .B(\SUBBYTES[8].a/w284 ), .Z(
        \SUBBYTES[8].a/w191 ) );
  AND U3366 ( .A(\SUBBYTES[8].a/w1908 ), .B(n1553), .Z(\SUBBYTES[8].a/w1909 )
         );
  XOR U3367 ( .A(n1554), .B(n1552), .Z(n1553) );
  IV U3368 ( .A(n14808), .Z(n1552) );
  ANDN U3369 ( .A(\SUBBYTES[8].a/w1927 ), .B(n1555), .Z(\SUBBYTES[8].a/w1904 )
         );
  ANDN U3370 ( .A(\SUBBYTES[8].a/w1928 ), .B(n1556), .Z(\SUBBYTES[8].a/w1902 )
         );
  ANDN U3371 ( .A(\SUBBYTES[8].a/w1931 ), .B(n1557), .Z(\SUBBYTES[8].a/w1901 )
         );
  AND U3372 ( .A(\SUBBYTES[8].a/w1887 ), .B(\SUBBYTES[8].a/w1886 ), .Z(
        \SUBBYTES[8].a/w1888 ) );
  IV U3373 ( .A(n1554), .Z(\SUBBYTES[8].a/w1884 ) );
  NAND U3374 ( .A(\SUBBYTES[8].a/w1863 ), .B(\SUBBYTES[8].a/w1878 ), .Z(n1554)
         );
  AND U3375 ( .A(\SUBBYTES[8].a/w1880 ), .B(\SUBBYTES[8].a/w1886 ), .Z(
        \SUBBYTES[8].a/w1881 ) );
  AND U3376 ( .A(\SUBBYTES[8].a/w1865 ), .B(\SUBBYTES[8].a/w1863 ), .Z(
        \SUBBYTES[8].a/w1875 ) );
  AND U3377 ( .A(\SUBBYTES[8].a/w1866 ), .B(\SUBBYTES[8].a/w1864 ), .Z(
        \SUBBYTES[8].a/w1873 ) );
  AND U3378 ( .A(\SUBBYTES[8].a/w1880 ), .B(\SUBBYTES[8].a/w1887 ), .Z(
        \SUBBYTES[8].a/w1872 ) );
  ANDN U3379 ( .A(\SUBBYTES[8].a/w273 ), .B(n1513), .Z(\SUBBYTES[8].a/w186 )
         );
  XNOR U3380 ( .A(\w1[8][124] ), .B(\w1[8][127] ), .Z(n1513) );
  AND U3381 ( .A(\SUBBYTES[8].a/w1820 ), .B(\SUBBYTES[8].a/w1816 ), .Z(
        \SUBBYTES[8].a/w1857 ) );
  AND U3382 ( .A(\SUBBYTES[8].a/w1821 ), .B(\SUBBYTES[8].a/w1817 ), .Z(
        \SUBBYTES[8].a/w1855 ) );
  ANDN U3383 ( .A(\SUBBYTES[8].a/w1947 ), .B(n1551), .Z(\SUBBYTES[8].a/w1854 )
         );
  XNOR U3384 ( .A(\w1[8][57] ), .B(\w1[8][63] ), .Z(n1551) );
  XOR U3385 ( .A(\w0[8][57] ), .B(g_input[1081]), .Z(\w1[8][57] ) );
  AND U3386 ( .A(\w1[8][56] ), .B(\SUBBYTES[8].a/w1822 ), .Z(
        \SUBBYTES[8].a/w1850 ) );
  XOR U3387 ( .A(\w0[8][56] ), .B(g_input[1080]), .Z(\w1[8][56] ) );
  AND U3388 ( .A(\SUBBYTES[8].a/w1823 ), .B(\SUBBYTES[8].a/w1819 ), .Z(
        \SUBBYTES[8].a/w1848 ) );
  AND U3389 ( .A(\SUBBYTES[8].a/w1908 ), .B(\SUBBYTES[8].a/w1940 ), .Z(
        \SUBBYTES[8].a/w1847 ) );
  ANDN U3390 ( .A(\SUBBYTES[8].a/w1929 ), .B(n1555), .Z(\SUBBYTES[8].a/w1842 )
         );
  XNOR U3391 ( .A(\w1[8][60] ), .B(\w1[8][63] ), .Z(n1555) );
  ANDN U3392 ( .A(\SUBBYTES[8].a/w1930 ), .B(n1556), .Z(\SUBBYTES[8].a/w1840 )
         );
  XNOR U3393 ( .A(\w1[8][58] ), .B(\w1[8][63] ), .Z(n1556) );
  XOR U3394 ( .A(\w0[8][63] ), .B(g_input[1087]), .Z(\w1[8][63] ) );
  IV U3395 ( .A(n1558), .Z(\w1[8][58] ) );
  ANDN U3396 ( .A(\SUBBYTES[8].a/w274 ), .B(n1515), .Z(\SUBBYTES[8].a/w184 )
         );
  XNOR U3397 ( .A(\w1[8][122] ), .B(\w1[8][127] ), .Z(n1515) );
  XOR U3398 ( .A(\w0[8][127] ), .B(g_input[1151]), .Z(\w1[8][127] ) );
  IV U3399 ( .A(n1559), .Z(\w1[8][122] ) );
  ANDN U3400 ( .A(\SUBBYTES[8].a/w1932 ), .B(n1557), .Z(\SUBBYTES[8].a/w1839 )
         );
  XOR U3401 ( .A(n1558), .B(\w1[8][60] ), .Z(n1557) );
  XOR U3402 ( .A(\w0[8][60] ), .B(g_input[1084]), .Z(\w1[8][60] ) );
  XNOR U3403 ( .A(\w0[8][58] ), .B(g_input[1082]), .Z(n1558) );
  ANDN U3404 ( .A(\SUBBYTES[8].a/w276 ), .B(n1516), .Z(\SUBBYTES[8].a/w183 )
         );
  XOR U3405 ( .A(n1559), .B(\w1[8][124] ), .Z(n1516) );
  XOR U3406 ( .A(\w0[8][124] ), .B(g_input[1148]), .Z(\w1[8][124] ) );
  XNOR U3407 ( .A(\w0[8][122] ), .B(g_input[1146]), .Z(n1559) );
  AND U3408 ( .A(n1560), .B(\SUBBYTES[8].a/w1609 ), .Z(\SUBBYTES[8].a/w1744 )
         );
  AND U3409 ( .A(n1561), .B(\SUBBYTES[8].a/w1610 ), .Z(\SUBBYTES[8].a/w1742 )
         );
  AND U3410 ( .A(\SUBBYTES[8].a/w1740 ), .B(n1562), .Z(\SUBBYTES[8].a/w1741 )
         );
  ANDN U3411 ( .A(\w1[8][64] ), .B(n1563), .Z(\SUBBYTES[8].a/w1737 ) );
  AND U3412 ( .A(n1564), .B(\SUBBYTES[8].a/w1612 ), .Z(\SUBBYTES[8].a/w1735 )
         );
  AND U3413 ( .A(\SUBBYTES[8].a/w1733 ), .B(n1565), .Z(\SUBBYTES[8].a/w1734 )
         );
  XOR U3414 ( .A(\SUBBYTES[8].a/w1677 ), .B(n14806), .Z(n1565) );
  AND U3415 ( .A(\SUBBYTES[8].a/w1720 ), .B(\SUBBYTES[8].a/w1722 ), .Z(
        \SUBBYTES[8].a/w1729 ) );
  AND U3416 ( .A(\SUBBYTES[8].a/w1721 ), .B(\SUBBYTES[8].a/w1723 ), .Z(
        \SUBBYTES[8].a/w1727 ) );
  AND U3417 ( .A(\SUBBYTES[8].a/w1724 ), .B(\SUBBYTES[8].a/w1725 ), .Z(
        \SUBBYTES[8].a/w1726 ) );
  AND U3418 ( .A(\SUBBYTES[8].a/w1613 ), .B(n1560), .Z(\SUBBYTES[8].a/w1712 )
         );
  XOR U3419 ( .A(\SUBBYTES[8].a/w1681 ), .B(n1076), .Z(n1560) );
  AND U3420 ( .A(\SUBBYTES[8].a/w1614 ), .B(n1561), .Z(\SUBBYTES[8].a/w1710 )
         );
  XOR U3421 ( .A(n14807), .B(\SUBBYTES[8].a/w1681 ), .Z(n1561) );
  ANDN U3422 ( .A(n1562), .B(n1566), .Z(\SUBBYTES[8].a/w1709 ) );
  XOR U3423 ( .A(n1076), .B(n14807), .Z(n1562) );
  ANDN U3424 ( .A(\SUBBYTES[8].a/w1615 ), .B(n1563), .Z(\SUBBYTES[8].a/w1705 )
         );
  XNOR U3425 ( .A(\SUBBYTES[8].a/w1674 ), .B(\SUBBYTES[8].a/w1677 ), .Z(n1563)
         );
  AND U3426 ( .A(\SUBBYTES[8].a/w1616 ), .B(n1564), .Z(\SUBBYTES[8].a/w1703 )
         );
  XNOR U3427 ( .A(n1567), .B(\SUBBYTES[8].a/w1674 ), .Z(n1564) );
  AND U3428 ( .A(\SUBBYTES[8].a/w1701 ), .B(n1568), .Z(\SUBBYTES[8].a/w1702 )
         );
  XOR U3429 ( .A(n1569), .B(n1567), .Z(n1568) );
  IV U3430 ( .A(n14806), .Z(n1567) );
  ANDN U3431 ( .A(\SUBBYTES[8].a/w1720 ), .B(n1570), .Z(\SUBBYTES[8].a/w1697 )
         );
  ANDN U3432 ( .A(\SUBBYTES[8].a/w1721 ), .B(n1571), .Z(\SUBBYTES[8].a/w1695 )
         );
  ANDN U3433 ( .A(\SUBBYTES[8].a/w1724 ), .B(n1572), .Z(\SUBBYTES[8].a/w1694 )
         );
  AND U3434 ( .A(\SUBBYTES[8].a/w1680 ), .B(\SUBBYTES[8].a/w1679 ), .Z(
        \SUBBYTES[8].a/w1681 ) );
  IV U3435 ( .A(n1569), .Z(\SUBBYTES[8].a/w1677 ) );
  NAND U3436 ( .A(\SUBBYTES[8].a/w1656 ), .B(\SUBBYTES[8].a/w1671 ), .Z(n1569)
         );
  AND U3437 ( .A(\SUBBYTES[8].a/w1673 ), .B(\SUBBYTES[8].a/w1679 ), .Z(
        \SUBBYTES[8].a/w1674 ) );
  AND U3438 ( .A(\SUBBYTES[8].a/w1658 ), .B(\SUBBYTES[8].a/w1656 ), .Z(
        \SUBBYTES[8].a/w1668 ) );
  AND U3439 ( .A(\SUBBYTES[8].a/w1659 ), .B(\SUBBYTES[8].a/w1657 ), .Z(
        \SUBBYTES[8].a/w1666 ) );
  AND U3440 ( .A(\SUBBYTES[8].a/w1673 ), .B(\SUBBYTES[8].a/w1680 ), .Z(
        \SUBBYTES[8].a/w1665 ) );
  AND U3441 ( .A(\SUBBYTES[8].a/w1613 ), .B(\SUBBYTES[8].a/w1609 ), .Z(
        \SUBBYTES[8].a/w1650 ) );
  AND U3442 ( .A(\SUBBYTES[8].a/w1614 ), .B(\SUBBYTES[8].a/w1610 ), .Z(
        \SUBBYTES[8].a/w1648 ) );
  ANDN U3443 ( .A(\SUBBYTES[8].a/w1740 ), .B(n1566), .Z(\SUBBYTES[8].a/w1647 )
         );
  XNOR U3444 ( .A(\w1[8][65] ), .B(\w1[8][71] ), .Z(n1566) );
  XOR U3445 ( .A(\w0[8][65] ), .B(g_input[1089]), .Z(\w1[8][65] ) );
  AND U3446 ( .A(\w1[8][64] ), .B(\SUBBYTES[8].a/w1615 ), .Z(
        \SUBBYTES[8].a/w1643 ) );
  XOR U3447 ( .A(\w0[8][64] ), .B(g_input[1088]), .Z(\w1[8][64] ) );
  AND U3448 ( .A(\SUBBYTES[8].a/w1616 ), .B(\SUBBYTES[8].a/w1612 ), .Z(
        \SUBBYTES[8].a/w1641 ) );
  AND U3449 ( .A(\SUBBYTES[8].a/w1701 ), .B(\SUBBYTES[8].a/w1733 ), .Z(
        \SUBBYTES[8].a/w1640 ) );
  ANDN U3450 ( .A(\SUBBYTES[8].a/w1722 ), .B(n1570), .Z(\SUBBYTES[8].a/w1635 )
         );
  XNOR U3451 ( .A(\w1[8][68] ), .B(\w1[8][71] ), .Z(n1570) );
  ANDN U3452 ( .A(\SUBBYTES[8].a/w1723 ), .B(n1571), .Z(\SUBBYTES[8].a/w1633 )
         );
  XNOR U3453 ( .A(\w1[8][66] ), .B(\w1[8][71] ), .Z(n1571) );
  XOR U3454 ( .A(\w0[8][71] ), .B(g_input[1095]), .Z(\w1[8][71] ) );
  IV U3455 ( .A(n1573), .Z(\w1[8][66] ) );
  ANDN U3456 ( .A(\SUBBYTES[8].a/w1725 ), .B(n1572), .Z(\SUBBYTES[8].a/w1632 )
         );
  XOR U3457 ( .A(n1573), .B(\w1[8][68] ), .Z(n1572) );
  XOR U3458 ( .A(\w0[8][68] ), .B(g_input[1092]), .Z(\w1[8][68] ) );
  XNOR U3459 ( .A(\w0[8][66] ), .B(g_input[1090]), .Z(n1573) );
  AND U3460 ( .A(n1574), .B(\SUBBYTES[8].a/w1402 ), .Z(\SUBBYTES[8].a/w1537 )
         );
  AND U3461 ( .A(n1575), .B(\SUBBYTES[8].a/w1403 ), .Z(\SUBBYTES[8].a/w1535 )
         );
  AND U3462 ( .A(\SUBBYTES[8].a/w1533 ), .B(n1576), .Z(\SUBBYTES[8].a/w1534 )
         );
  ANDN U3463 ( .A(\w1[8][72] ), .B(n1577), .Z(\SUBBYTES[8].a/w1530 ) );
  AND U3464 ( .A(n1578), .B(\SUBBYTES[8].a/w1405 ), .Z(\SUBBYTES[8].a/w1528 )
         );
  AND U3465 ( .A(\SUBBYTES[8].a/w1526 ), .B(n1579), .Z(\SUBBYTES[8].a/w1527 )
         );
  XOR U3466 ( .A(\SUBBYTES[8].a/w1470 ), .B(n14804), .Z(n1579) );
  AND U3467 ( .A(\SUBBYTES[8].a/w1513 ), .B(\SUBBYTES[8].a/w1515 ), .Z(
        \SUBBYTES[8].a/w1522 ) );
  AND U3468 ( .A(\SUBBYTES[8].a/w1514 ), .B(\SUBBYTES[8].a/w1516 ), .Z(
        \SUBBYTES[8].a/w1520 ) );
  AND U3469 ( .A(\SUBBYTES[8].a/w1517 ), .B(\SUBBYTES[8].a/w1518 ), .Z(
        \SUBBYTES[8].a/w1519 ) );
  AND U3470 ( .A(\SUBBYTES[8].a/w1406 ), .B(n1574), .Z(\SUBBYTES[8].a/w1505 )
         );
  XOR U3471 ( .A(\SUBBYTES[8].a/w1474 ), .B(n1075), .Z(n1574) );
  AND U3472 ( .A(\SUBBYTES[8].a/w1407 ), .B(n1575), .Z(\SUBBYTES[8].a/w1503 )
         );
  XOR U3473 ( .A(n14805), .B(\SUBBYTES[8].a/w1474 ), .Z(n1575) );
  ANDN U3474 ( .A(n1576), .B(n1580), .Z(\SUBBYTES[8].a/w1502 ) );
  XOR U3475 ( .A(n1075), .B(n14805), .Z(n1576) );
  ANDN U3476 ( .A(\SUBBYTES[8].a/w1408 ), .B(n1577), .Z(\SUBBYTES[8].a/w1498 )
         );
  XNOR U3477 ( .A(\SUBBYTES[8].a/w1467 ), .B(\SUBBYTES[8].a/w1470 ), .Z(n1577)
         );
  AND U3478 ( .A(\SUBBYTES[8].a/w1409 ), .B(n1578), .Z(\SUBBYTES[8].a/w1496 )
         );
  XNOR U3479 ( .A(n1581), .B(\SUBBYTES[8].a/w1467 ), .Z(n1578) );
  AND U3480 ( .A(\SUBBYTES[8].a/w1494 ), .B(n1582), .Z(\SUBBYTES[8].a/w1495 )
         );
  XOR U3481 ( .A(n1583), .B(n1581), .Z(n1582) );
  IV U3482 ( .A(n14804), .Z(n1581) );
  ANDN U3483 ( .A(\SUBBYTES[8].a/w1513 ), .B(n1584), .Z(\SUBBYTES[8].a/w1490 )
         );
  ANDN U3484 ( .A(\SUBBYTES[8].a/w1514 ), .B(n1585), .Z(\SUBBYTES[8].a/w1488 )
         );
  ANDN U3485 ( .A(\SUBBYTES[8].a/w1517 ), .B(n1586), .Z(\SUBBYTES[8].a/w1487 )
         );
  AND U3486 ( .A(\SUBBYTES[8].a/w1473 ), .B(\SUBBYTES[8].a/w1472 ), .Z(
        \SUBBYTES[8].a/w1474 ) );
  IV U3487 ( .A(n1583), .Z(\SUBBYTES[8].a/w1470 ) );
  NAND U3488 ( .A(\SUBBYTES[8].a/w1449 ), .B(\SUBBYTES[8].a/w1464 ), .Z(n1583)
         );
  AND U3489 ( .A(\SUBBYTES[8].a/w1466 ), .B(\SUBBYTES[8].a/w1472 ), .Z(
        \SUBBYTES[8].a/w1467 ) );
  AND U3490 ( .A(\SUBBYTES[8].a/w1451 ), .B(\SUBBYTES[8].a/w1449 ), .Z(
        \SUBBYTES[8].a/w1461 ) );
  AND U3491 ( .A(\SUBBYTES[8].a/w1452 ), .B(\SUBBYTES[8].a/w1450 ), .Z(
        \SUBBYTES[8].a/w1459 ) );
  AND U3492 ( .A(\SUBBYTES[8].a/w1466 ), .B(\SUBBYTES[8].a/w1473 ), .Z(
        \SUBBYTES[8].a/w1458 ) );
  AND U3493 ( .A(\SUBBYTES[8].a/w1406 ), .B(\SUBBYTES[8].a/w1402 ), .Z(
        \SUBBYTES[8].a/w1443 ) );
  AND U3494 ( .A(\SUBBYTES[8].a/w1407 ), .B(\SUBBYTES[8].a/w1403 ), .Z(
        \SUBBYTES[8].a/w1441 ) );
  ANDN U3495 ( .A(\SUBBYTES[8].a/w1533 ), .B(n1580), .Z(\SUBBYTES[8].a/w1440 )
         );
  XNOR U3496 ( .A(\w1[8][73] ), .B(\w1[8][79] ), .Z(n1580) );
  XOR U3497 ( .A(\w0[8][73] ), .B(g_input[1097]), .Z(\w1[8][73] ) );
  AND U3498 ( .A(\w1[8][72] ), .B(\SUBBYTES[8].a/w1408 ), .Z(
        \SUBBYTES[8].a/w1436 ) );
  XOR U3499 ( .A(\w0[8][72] ), .B(g_input[1096]), .Z(\w1[8][72] ) );
  AND U3500 ( .A(\SUBBYTES[8].a/w1409 ), .B(\SUBBYTES[8].a/w1405 ), .Z(
        \SUBBYTES[8].a/w1434 ) );
  AND U3501 ( .A(\SUBBYTES[8].a/w1494 ), .B(\SUBBYTES[8].a/w1526 ), .Z(
        \SUBBYTES[8].a/w1433 ) );
  ANDN U3502 ( .A(\SUBBYTES[8].a/w1515 ), .B(n1584), .Z(\SUBBYTES[8].a/w1428 )
         );
  XNOR U3503 ( .A(\w1[8][76] ), .B(\w1[8][79] ), .Z(n1584) );
  ANDN U3504 ( .A(\SUBBYTES[8].a/w1516 ), .B(n1585), .Z(\SUBBYTES[8].a/w1426 )
         );
  XNOR U3505 ( .A(\w1[8][74] ), .B(\w1[8][79] ), .Z(n1585) );
  XOR U3506 ( .A(\w0[8][79] ), .B(g_input[1103]), .Z(\w1[8][79] ) );
  IV U3507 ( .A(n1587), .Z(\w1[8][74] ) );
  ANDN U3508 ( .A(\SUBBYTES[8].a/w1518 ), .B(n1586), .Z(\SUBBYTES[8].a/w1425 )
         );
  XOR U3509 ( .A(n1587), .B(\w1[8][76] ), .Z(n1586) );
  XOR U3510 ( .A(\w0[8][76] ), .B(g_input[1100]), .Z(\w1[8][76] ) );
  XNOR U3511 ( .A(\w0[8][74] ), .B(g_input[1098]), .Z(n1587) );
  AND U3512 ( .A(n1588), .B(\SUBBYTES[8].a/w1195 ), .Z(\SUBBYTES[8].a/w1330 )
         );
  AND U3513 ( .A(n1589), .B(\SUBBYTES[8].a/w1196 ), .Z(\SUBBYTES[8].a/w1328 )
         );
  AND U3514 ( .A(\SUBBYTES[8].a/w1326 ), .B(n1590), .Z(\SUBBYTES[8].a/w1327 )
         );
  ANDN U3515 ( .A(\w1[8][80] ), .B(n1591), .Z(\SUBBYTES[8].a/w1323 ) );
  AND U3516 ( .A(n1592), .B(\SUBBYTES[8].a/w1198 ), .Z(\SUBBYTES[8].a/w1321 )
         );
  AND U3517 ( .A(\SUBBYTES[8].a/w1319 ), .B(n1593), .Z(\SUBBYTES[8].a/w1320 )
         );
  XOR U3518 ( .A(\SUBBYTES[8].a/w1263 ), .B(n14802), .Z(n1593) );
  AND U3519 ( .A(\SUBBYTES[8].a/w1306 ), .B(\SUBBYTES[8].a/w1308 ), .Z(
        \SUBBYTES[8].a/w1315 ) );
  AND U3520 ( .A(\SUBBYTES[8].a/w1307 ), .B(\SUBBYTES[8].a/w1309 ), .Z(
        \SUBBYTES[8].a/w1313 ) );
  AND U3521 ( .A(\SUBBYTES[8].a/w1310 ), .B(\SUBBYTES[8].a/w1311 ), .Z(
        \SUBBYTES[8].a/w1312 ) );
  AND U3522 ( .A(\SUBBYTES[8].a/w1199 ), .B(n1588), .Z(\SUBBYTES[8].a/w1298 )
         );
  XOR U3523 ( .A(\SUBBYTES[8].a/w1267 ), .B(n1074), .Z(n1588) );
  AND U3524 ( .A(\SUBBYTES[8].a/w1200 ), .B(n1589), .Z(\SUBBYTES[8].a/w1296 )
         );
  XOR U3525 ( .A(n14803), .B(\SUBBYTES[8].a/w1267 ), .Z(n1589) );
  ANDN U3526 ( .A(n1590), .B(n1594), .Z(\SUBBYTES[8].a/w1295 ) );
  XOR U3527 ( .A(n1074), .B(n14803), .Z(n1590) );
  ANDN U3528 ( .A(\SUBBYTES[8].a/w1201 ), .B(n1591), .Z(\SUBBYTES[8].a/w1291 )
         );
  XNOR U3529 ( .A(\SUBBYTES[8].a/w1260 ), .B(\SUBBYTES[8].a/w1263 ), .Z(n1591)
         );
  AND U3530 ( .A(\SUBBYTES[8].a/w1202 ), .B(n1592), .Z(\SUBBYTES[8].a/w1289 )
         );
  XNOR U3531 ( .A(n1595), .B(\SUBBYTES[8].a/w1260 ), .Z(n1592) );
  AND U3532 ( .A(\SUBBYTES[8].a/w1287 ), .B(n1596), .Z(\SUBBYTES[8].a/w1288 )
         );
  XOR U3533 ( .A(n1597), .B(n1595), .Z(n1596) );
  IV U3534 ( .A(n14802), .Z(n1595) );
  ANDN U3535 ( .A(\SUBBYTES[8].a/w1306 ), .B(n1598), .Z(\SUBBYTES[8].a/w1283 )
         );
  ANDN U3536 ( .A(\SUBBYTES[8].a/w1307 ), .B(n1599), .Z(\SUBBYTES[8].a/w1281 )
         );
  ANDN U3537 ( .A(\SUBBYTES[8].a/w1310 ), .B(n1600), .Z(\SUBBYTES[8].a/w1280 )
         );
  AND U3538 ( .A(\SUBBYTES[8].a/w1266 ), .B(\SUBBYTES[8].a/w1265 ), .Z(
        \SUBBYTES[8].a/w1267 ) );
  IV U3539 ( .A(n1597), .Z(\SUBBYTES[8].a/w1263 ) );
  NAND U3540 ( .A(\SUBBYTES[8].a/w1242 ), .B(\SUBBYTES[8].a/w1257 ), .Z(n1597)
         );
  AND U3541 ( .A(\SUBBYTES[8].a/w1259 ), .B(\SUBBYTES[8].a/w1265 ), .Z(
        \SUBBYTES[8].a/w1260 ) );
  AND U3542 ( .A(\SUBBYTES[8].a/w1244 ), .B(\SUBBYTES[8].a/w1242 ), .Z(
        \SUBBYTES[8].a/w1254 ) );
  AND U3543 ( .A(\SUBBYTES[8].a/w1245 ), .B(\SUBBYTES[8].a/w1243 ), .Z(
        \SUBBYTES[8].a/w1252 ) );
  AND U3544 ( .A(\SUBBYTES[8].a/w1259 ), .B(\SUBBYTES[8].a/w1266 ), .Z(
        \SUBBYTES[8].a/w1251 ) );
  AND U3545 ( .A(\SUBBYTES[8].a/w1199 ), .B(\SUBBYTES[8].a/w1195 ), .Z(
        \SUBBYTES[8].a/w1236 ) );
  AND U3546 ( .A(\SUBBYTES[8].a/w1200 ), .B(\SUBBYTES[8].a/w1196 ), .Z(
        \SUBBYTES[8].a/w1234 ) );
  ANDN U3547 ( .A(\SUBBYTES[8].a/w1326 ), .B(n1594), .Z(\SUBBYTES[8].a/w1233 )
         );
  XNOR U3548 ( .A(\w1[8][81] ), .B(\w1[8][87] ), .Z(n1594) );
  XOR U3549 ( .A(\w0[8][81] ), .B(g_input[1105]), .Z(\w1[8][81] ) );
  AND U3550 ( .A(\w1[8][80] ), .B(\SUBBYTES[8].a/w1201 ), .Z(
        \SUBBYTES[8].a/w1229 ) );
  XOR U3551 ( .A(\w0[8][80] ), .B(g_input[1104]), .Z(\w1[8][80] ) );
  AND U3552 ( .A(\SUBBYTES[8].a/w1202 ), .B(\SUBBYTES[8].a/w1198 ), .Z(
        \SUBBYTES[8].a/w1227 ) );
  AND U3553 ( .A(\SUBBYTES[8].a/w1287 ), .B(\SUBBYTES[8].a/w1319 ), .Z(
        \SUBBYTES[8].a/w1226 ) );
  ANDN U3554 ( .A(\SUBBYTES[8].a/w1308 ), .B(n1598), .Z(\SUBBYTES[8].a/w1221 )
         );
  XNOR U3555 ( .A(\w1[8][84] ), .B(\w1[8][87] ), .Z(n1598) );
  ANDN U3556 ( .A(\SUBBYTES[8].a/w1309 ), .B(n1599), .Z(\SUBBYTES[8].a/w1219 )
         );
  XNOR U3557 ( .A(\w1[8][82] ), .B(\w1[8][87] ), .Z(n1599) );
  XOR U3558 ( .A(\w0[8][87] ), .B(g_input[1111]), .Z(\w1[8][87] ) );
  IV U3559 ( .A(n1601), .Z(\w1[8][82] ) );
  ANDN U3560 ( .A(\SUBBYTES[8].a/w1311 ), .B(n1600), .Z(\SUBBYTES[8].a/w1218 )
         );
  XOR U3561 ( .A(n1601), .B(\w1[8][84] ), .Z(n1600) );
  XOR U3562 ( .A(\w0[8][84] ), .B(g_input[1108]), .Z(\w1[8][84] ) );
  XNOR U3563 ( .A(\w0[8][82] ), .B(g_input[1106]), .Z(n1601) );
  AND U3564 ( .A(n1602), .B(\SUBBYTES[8].a/w988 ), .Z(\SUBBYTES[8].a/w1123 )
         );
  AND U3565 ( .A(n1603), .B(\SUBBYTES[8].a/w989 ), .Z(\SUBBYTES[8].a/w1121 )
         );
  AND U3566 ( .A(\SUBBYTES[8].a/w1119 ), .B(n1604), .Z(\SUBBYTES[8].a/w1120 )
         );
  ANDN U3567 ( .A(\w1[8][88] ), .B(n1605), .Z(\SUBBYTES[8].a/w1116 ) );
  AND U3568 ( .A(n1606), .B(\SUBBYTES[8].a/w991 ), .Z(\SUBBYTES[8].a/w1114 )
         );
  AND U3569 ( .A(\SUBBYTES[8].a/w1112 ), .B(n1607), .Z(\SUBBYTES[8].a/w1113 )
         );
  XOR U3570 ( .A(\SUBBYTES[8].a/w1056 ), .B(n14800), .Z(n1607) );
  AND U3571 ( .A(\SUBBYTES[8].a/w1099 ), .B(\SUBBYTES[8].a/w1101 ), .Z(
        \SUBBYTES[8].a/w1108 ) );
  AND U3572 ( .A(\SUBBYTES[8].a/w1100 ), .B(\SUBBYTES[8].a/w1102 ), .Z(
        \SUBBYTES[8].a/w1106 ) );
  AND U3573 ( .A(\SUBBYTES[8].a/w1103 ), .B(\SUBBYTES[8].a/w1104 ), .Z(
        \SUBBYTES[8].a/w1105 ) );
  AND U3574 ( .A(\SUBBYTES[8].a/w992 ), .B(n1602), .Z(\SUBBYTES[8].a/w1091 )
         );
  XOR U3575 ( .A(\SUBBYTES[8].a/w1060 ), .B(n1073), .Z(n1602) );
  AND U3576 ( .A(\SUBBYTES[8].a/w993 ), .B(n1603), .Z(\SUBBYTES[8].a/w1089 )
         );
  XOR U3577 ( .A(n14801), .B(\SUBBYTES[8].a/w1060 ), .Z(n1603) );
  ANDN U3578 ( .A(n1604), .B(n1608), .Z(\SUBBYTES[8].a/w1088 ) );
  XOR U3579 ( .A(n1073), .B(n14801), .Z(n1604) );
  ANDN U3580 ( .A(\SUBBYTES[8].a/w994 ), .B(n1605), .Z(\SUBBYTES[8].a/w1084 )
         );
  XNOR U3581 ( .A(\SUBBYTES[8].a/w1053 ), .B(\SUBBYTES[8].a/w1056 ), .Z(n1605)
         );
  AND U3582 ( .A(\SUBBYTES[8].a/w995 ), .B(n1606), .Z(\SUBBYTES[8].a/w1082 )
         );
  XNOR U3583 ( .A(n1609), .B(\SUBBYTES[8].a/w1053 ), .Z(n1606) );
  AND U3584 ( .A(\SUBBYTES[8].a/w1080 ), .B(n1610), .Z(\SUBBYTES[8].a/w1081 )
         );
  XOR U3585 ( .A(n1611), .B(n1609), .Z(n1610) );
  IV U3586 ( .A(n14800), .Z(n1609) );
  ANDN U3587 ( .A(\SUBBYTES[8].a/w1099 ), .B(n1612), .Z(\SUBBYTES[8].a/w1076 )
         );
  ANDN U3588 ( .A(\SUBBYTES[8].a/w1100 ), .B(n1613), .Z(\SUBBYTES[8].a/w1074 )
         );
  ANDN U3589 ( .A(\SUBBYTES[8].a/w1103 ), .B(n1614), .Z(\SUBBYTES[8].a/w1073 )
         );
  AND U3590 ( .A(\SUBBYTES[8].a/w1059 ), .B(\SUBBYTES[8].a/w1058 ), .Z(
        \SUBBYTES[8].a/w1060 ) );
  IV U3591 ( .A(n1611), .Z(\SUBBYTES[8].a/w1056 ) );
  NAND U3592 ( .A(\SUBBYTES[8].a/w1035 ), .B(\SUBBYTES[8].a/w1050 ), .Z(n1611)
         );
  AND U3593 ( .A(\SUBBYTES[8].a/w1052 ), .B(\SUBBYTES[8].a/w1058 ), .Z(
        \SUBBYTES[8].a/w1053 ) );
  AND U3594 ( .A(\SUBBYTES[8].a/w1037 ), .B(\SUBBYTES[8].a/w1035 ), .Z(
        \SUBBYTES[8].a/w1047 ) );
  AND U3595 ( .A(\SUBBYTES[8].a/w1038 ), .B(\SUBBYTES[8].a/w1036 ), .Z(
        \SUBBYTES[8].a/w1045 ) );
  AND U3596 ( .A(\SUBBYTES[8].a/w1052 ), .B(\SUBBYTES[8].a/w1059 ), .Z(
        \SUBBYTES[8].a/w1044 ) );
  AND U3597 ( .A(\SUBBYTES[8].a/w992 ), .B(\SUBBYTES[8].a/w988 ), .Z(
        \SUBBYTES[8].a/w1029 ) );
  AND U3598 ( .A(\SUBBYTES[8].a/w993 ), .B(\SUBBYTES[8].a/w989 ), .Z(
        \SUBBYTES[8].a/w1027 ) );
  ANDN U3599 ( .A(\SUBBYTES[8].a/w1119 ), .B(n1608), .Z(\SUBBYTES[8].a/w1026 )
         );
  XNOR U3600 ( .A(\w1[8][89] ), .B(\w1[8][95] ), .Z(n1608) );
  XOR U3601 ( .A(\w0[8][89] ), .B(g_input[1113]), .Z(\w1[8][89] ) );
  AND U3602 ( .A(\w1[8][88] ), .B(\SUBBYTES[8].a/w994 ), .Z(
        \SUBBYTES[8].a/w1022 ) );
  XOR U3603 ( .A(\w0[8][88] ), .B(g_input[1112]), .Z(\w1[8][88] ) );
  AND U3604 ( .A(\SUBBYTES[8].a/w995 ), .B(\SUBBYTES[8].a/w991 ), .Z(
        \SUBBYTES[8].a/w1020 ) );
  AND U3605 ( .A(\SUBBYTES[8].a/w1080 ), .B(\SUBBYTES[8].a/w1112 ), .Z(
        \SUBBYTES[8].a/w1019 ) );
  ANDN U3606 ( .A(\SUBBYTES[8].a/w1101 ), .B(n1612), .Z(\SUBBYTES[8].a/w1014 )
         );
  XNOR U3607 ( .A(\w1[8][92] ), .B(\w1[8][95] ), .Z(n1612) );
  ANDN U3608 ( .A(\SUBBYTES[8].a/w1102 ), .B(n1613), .Z(\SUBBYTES[8].a/w1012 )
         );
  XNOR U3609 ( .A(\w1[8][90] ), .B(\w1[8][95] ), .Z(n1613) );
  XOR U3610 ( .A(\w0[8][95] ), .B(g_input[1119]), .Z(\w1[8][95] ) );
  IV U3611 ( .A(n1615), .Z(\w1[8][90] ) );
  ANDN U3612 ( .A(\SUBBYTES[8].a/w1104 ), .B(n1614), .Z(\SUBBYTES[8].a/w1011 )
         );
  XOR U3613 ( .A(n1615), .B(\w1[8][92] ), .Z(n1614) );
  XOR U3614 ( .A(\w0[8][92] ), .B(g_input[1116]), .Z(\w1[8][92] ) );
  XNOR U3615 ( .A(\w0[8][90] ), .B(g_input[1114]), .Z(n1615) );
  AND U3616 ( .A(\SUBBYTES[8].a/w2084 ), .B(\SUBBYTES[8].a/w2071 ), .Z(n14810)
         );
  AND U3617 ( .A(\SUBBYTES[8].a/w1877 ), .B(\SUBBYTES[8].a/w1866 ), .Z(n14809)
         );
  AND U3618 ( .A(\SUBBYTES[8].a/w221 ), .B(\SUBBYTES[8].a/w208 ), .Z(n14792)
         );
  AND U3619 ( .A(\SUBBYTES[8].a/w1877 ), .B(\SUBBYTES[8].a/w1864 ), .Z(n14808)
         );
  AND U3620 ( .A(\SUBBYTES[8].a/w1670 ), .B(\SUBBYTES[8].a/w1659 ), .Z(n14807)
         );
  AND U3621 ( .A(\SUBBYTES[8].a/w1670 ), .B(\SUBBYTES[8].a/w1657 ), .Z(n14806)
         );
  AND U3622 ( .A(\SUBBYTES[8].a/w1463 ), .B(\SUBBYTES[8].a/w1452 ), .Z(n14805)
         );
  AND U3623 ( .A(\SUBBYTES[8].a/w1463 ), .B(\SUBBYTES[8].a/w1450 ), .Z(n14804)
         );
  AND U3624 ( .A(\SUBBYTES[8].a/w1256 ), .B(\SUBBYTES[8].a/w1245 ), .Z(n14803)
         );
  AND U3625 ( .A(\SUBBYTES[8].a/w1256 ), .B(\SUBBYTES[8].a/w1243 ), .Z(n14802)
         );
  AND U3626 ( .A(\SUBBYTES[8].a/w1049 ), .B(\SUBBYTES[8].a/w1038 ), .Z(n14801)
         );
  AND U3627 ( .A(\SUBBYTES[8].a/w1049 ), .B(\SUBBYTES[8].a/w1036 ), .Z(n14800)
         );
  AND U3628 ( .A(\SUBBYTES[8].a/w842 ), .B(\SUBBYTES[8].a/w831 ), .Z(n14799)
         );
  AND U3629 ( .A(\SUBBYTES[8].a/w842 ), .B(\SUBBYTES[8].a/w829 ), .Z(n14798)
         );
  AND U3630 ( .A(\SUBBYTES[8].a/w635 ), .B(\SUBBYTES[8].a/w624 ), .Z(n14797)
         );
  AND U3631 ( .A(\SUBBYTES[8].a/w635 ), .B(\SUBBYTES[8].a/w622 ), .Z(n14796)
         );
  AND U3632 ( .A(\SUBBYTES[8].a/w428 ), .B(\SUBBYTES[8].a/w417 ), .Z(n14795)
         );
  AND U3633 ( .A(\SUBBYTES[8].a/w428 ), .B(\SUBBYTES[8].a/w415 ), .Z(n14794)
         );
  AND U3634 ( .A(\SUBBYTES[8].a/w3326 ), .B(\SUBBYTES[8].a/w3315 ), .Z(n14823)
         );
  AND U3635 ( .A(\SUBBYTES[8].a/w3326 ), .B(\SUBBYTES[8].a/w3313 ), .Z(n14822)
         );
  AND U3636 ( .A(\SUBBYTES[8].a/w3119 ), .B(\SUBBYTES[8].a/w3108 ), .Z(n14821)
         );
  AND U3637 ( .A(\SUBBYTES[8].a/w3119 ), .B(\SUBBYTES[8].a/w3106 ), .Z(n14820)
         );
  AND U3638 ( .A(\SUBBYTES[8].a/w2912 ), .B(\SUBBYTES[8].a/w2901 ), .Z(n14819)
         );
  AND U3639 ( .A(\SUBBYTES[8].a/w2912 ), .B(\SUBBYTES[8].a/w2899 ), .Z(n14818)
         );
  AND U3640 ( .A(\SUBBYTES[8].a/w2705 ), .B(\SUBBYTES[8].a/w2694 ), .Z(n14817)
         );
  AND U3641 ( .A(\SUBBYTES[8].a/w2705 ), .B(\SUBBYTES[8].a/w2692 ), .Z(n14816)
         );
  AND U3642 ( .A(\SUBBYTES[8].a/w2498 ), .B(\SUBBYTES[8].a/w2487 ), .Z(n14815)
         );
  AND U3643 ( .A(\SUBBYTES[8].a/w2498 ), .B(\SUBBYTES[8].a/w2485 ), .Z(n14814)
         );
  AND U3644 ( .A(\SUBBYTES[8].a/w2291 ), .B(\SUBBYTES[8].a/w2280 ), .Z(n14813)
         );
  AND U3645 ( .A(\SUBBYTES[8].a/w2291 ), .B(\SUBBYTES[8].a/w2278 ), .Z(n14812)
         );
  AND U3646 ( .A(\SUBBYTES[8].a/w2084 ), .B(\SUBBYTES[8].a/w2073 ), .Z(n14811)
         );
  AND U3647 ( .A(\SUBBYTES[8].a/w221 ), .B(\SUBBYTES[8].a/w210 ), .Z(n14793)
         );
  AND U3648 ( .A(n1616), .B(\SUBBYTES[7].a/w781 ), .Z(\SUBBYTES[7].a/w916 ) );
  AND U3649 ( .A(n1617), .B(\SUBBYTES[7].a/w782 ), .Z(\SUBBYTES[7].a/w914 ) );
  AND U3650 ( .A(\SUBBYTES[7].a/w912 ), .B(n1618), .Z(\SUBBYTES[7].a/w913 ) );
  ANDN U3651 ( .A(\w1[7][96] ), .B(n1619), .Z(\SUBBYTES[7].a/w909 ) );
  AND U3652 ( .A(n1620), .B(\SUBBYTES[7].a/w784 ), .Z(\SUBBYTES[7].a/w907 ) );
  AND U3653 ( .A(\SUBBYTES[7].a/w905 ), .B(n1621), .Z(\SUBBYTES[7].a/w906 ) );
  XOR U3654 ( .A(\SUBBYTES[7].a/w849 ), .B(n13518), .Z(n1621) );
  AND U3655 ( .A(\SUBBYTES[7].a/w892 ), .B(\SUBBYTES[7].a/w894 ), .Z(
        \SUBBYTES[7].a/w901 ) );
  AND U3656 ( .A(\SUBBYTES[7].a/w893 ), .B(\SUBBYTES[7].a/w895 ), .Z(
        \SUBBYTES[7].a/w899 ) );
  AND U3657 ( .A(\SUBBYTES[7].a/w896 ), .B(\SUBBYTES[7].a/w897 ), .Z(
        \SUBBYTES[7].a/w898 ) );
  AND U3658 ( .A(\SUBBYTES[7].a/w785 ), .B(n1616), .Z(\SUBBYTES[7].a/w884 ) );
  XOR U3659 ( .A(\SUBBYTES[7].a/w853 ), .B(n1056), .Z(n1616) );
  AND U3660 ( .A(\SUBBYTES[7].a/w786 ), .B(n1617), .Z(\SUBBYTES[7].a/w882 ) );
  XOR U3661 ( .A(n13519), .B(\SUBBYTES[7].a/w853 ), .Z(n1617) );
  ANDN U3662 ( .A(n1618), .B(n1622), .Z(\SUBBYTES[7].a/w881 ) );
  XOR U3663 ( .A(n1056), .B(n13519), .Z(n1618) );
  ANDN U3664 ( .A(\SUBBYTES[7].a/w787 ), .B(n1619), .Z(\SUBBYTES[7].a/w877 )
         );
  XNOR U3665 ( .A(\SUBBYTES[7].a/w846 ), .B(\SUBBYTES[7].a/w849 ), .Z(n1619)
         );
  AND U3666 ( .A(\SUBBYTES[7].a/w788 ), .B(n1620), .Z(\SUBBYTES[7].a/w875 ) );
  XNOR U3667 ( .A(n1623), .B(\SUBBYTES[7].a/w846 ), .Z(n1620) );
  AND U3668 ( .A(\SUBBYTES[7].a/w873 ), .B(n1624), .Z(\SUBBYTES[7].a/w874 ) );
  XOR U3669 ( .A(n1625), .B(n1623), .Z(n1624) );
  IV U3670 ( .A(n13518), .Z(n1623) );
  ANDN U3671 ( .A(\SUBBYTES[7].a/w892 ), .B(n1626), .Z(\SUBBYTES[7].a/w869 )
         );
  ANDN U3672 ( .A(\SUBBYTES[7].a/w893 ), .B(n1627), .Z(\SUBBYTES[7].a/w867 )
         );
  ANDN U3673 ( .A(\SUBBYTES[7].a/w896 ), .B(n1628), .Z(\SUBBYTES[7].a/w866 )
         );
  AND U3674 ( .A(\SUBBYTES[7].a/w852 ), .B(\SUBBYTES[7].a/w851 ), .Z(
        \SUBBYTES[7].a/w853 ) );
  IV U3675 ( .A(n1625), .Z(\SUBBYTES[7].a/w849 ) );
  NAND U3676 ( .A(\SUBBYTES[7].a/w828 ), .B(\SUBBYTES[7].a/w843 ), .Z(n1625)
         );
  AND U3677 ( .A(\SUBBYTES[7].a/w845 ), .B(\SUBBYTES[7].a/w851 ), .Z(
        \SUBBYTES[7].a/w846 ) );
  AND U3678 ( .A(\SUBBYTES[7].a/w830 ), .B(\SUBBYTES[7].a/w828 ), .Z(
        \SUBBYTES[7].a/w840 ) );
  AND U3679 ( .A(\SUBBYTES[7].a/w831 ), .B(\SUBBYTES[7].a/w829 ), .Z(
        \SUBBYTES[7].a/w838 ) );
  AND U3680 ( .A(\SUBBYTES[7].a/w845 ), .B(\SUBBYTES[7].a/w852 ), .Z(
        \SUBBYTES[7].a/w837 ) );
  AND U3681 ( .A(\SUBBYTES[7].a/w785 ), .B(\SUBBYTES[7].a/w781 ), .Z(
        \SUBBYTES[7].a/w822 ) );
  AND U3682 ( .A(\SUBBYTES[7].a/w786 ), .B(\SUBBYTES[7].a/w782 ), .Z(
        \SUBBYTES[7].a/w820 ) );
  ANDN U3683 ( .A(\SUBBYTES[7].a/w912 ), .B(n1622), .Z(\SUBBYTES[7].a/w819 )
         );
  XNOR U3684 ( .A(\w1[7][103] ), .B(\w1[7][97] ), .Z(n1622) );
  XOR U3685 ( .A(\w0[7][97] ), .B(g_input[993]), .Z(\w1[7][97] ) );
  IV U3686 ( .A(n1629), .Z(\w1[7][103] ) );
  AND U3687 ( .A(\w1[7][96] ), .B(\SUBBYTES[7].a/w787 ), .Z(
        \SUBBYTES[7].a/w815 ) );
  XOR U3688 ( .A(\w0[7][96] ), .B(g_input[992]), .Z(\w1[7][96] ) );
  AND U3689 ( .A(\SUBBYTES[7].a/w788 ), .B(\SUBBYTES[7].a/w784 ), .Z(
        \SUBBYTES[7].a/w813 ) );
  AND U3690 ( .A(\SUBBYTES[7].a/w873 ), .B(\SUBBYTES[7].a/w905 ), .Z(
        \SUBBYTES[7].a/w812 ) );
  ANDN U3691 ( .A(\SUBBYTES[7].a/w894 ), .B(n1626), .Z(\SUBBYTES[7].a/w807 )
         );
  XOR U3692 ( .A(\w1[7][100] ), .B(n1629), .Z(n1626) );
  ANDN U3693 ( .A(\SUBBYTES[7].a/w895 ), .B(n1627), .Z(\SUBBYTES[7].a/w805 )
         );
  XOR U3694 ( .A(n1629), .B(\w1[7][98] ), .Z(n1627) );
  XNOR U3695 ( .A(\w0[7][103] ), .B(g_input[999]), .Z(n1629) );
  ANDN U3696 ( .A(\SUBBYTES[7].a/w897 ), .B(n1628), .Z(\SUBBYTES[7].a/w804 )
         );
  XNOR U3697 ( .A(\w1[7][100] ), .B(\w1[7][98] ), .Z(n1628) );
  XOR U3698 ( .A(\w0[7][98] ), .B(g_input[994]), .Z(\w1[7][98] ) );
  XOR U3699 ( .A(\w0[7][100] ), .B(g_input[996]), .Z(\w1[7][100] ) );
  AND U3700 ( .A(n1630), .B(\SUBBYTES[7].a/w574 ), .Z(\SUBBYTES[7].a/w709 ) );
  AND U3701 ( .A(n1631), .B(\SUBBYTES[7].a/w575 ), .Z(\SUBBYTES[7].a/w707 ) );
  AND U3702 ( .A(\SUBBYTES[7].a/w705 ), .B(n1632), .Z(\SUBBYTES[7].a/w706 ) );
  ANDN U3703 ( .A(\w1[7][104] ), .B(n1633), .Z(\SUBBYTES[7].a/w702 ) );
  AND U3704 ( .A(n1634), .B(\SUBBYTES[7].a/w577 ), .Z(\SUBBYTES[7].a/w700 ) );
  AND U3705 ( .A(\SUBBYTES[7].a/w698 ), .B(n1635), .Z(\SUBBYTES[7].a/w699 ) );
  XOR U3706 ( .A(\SUBBYTES[7].a/w642 ), .B(n13516), .Z(n1635) );
  AND U3707 ( .A(\SUBBYTES[7].a/w685 ), .B(\SUBBYTES[7].a/w687 ), .Z(
        \SUBBYTES[7].a/w694 ) );
  AND U3708 ( .A(\SUBBYTES[7].a/w686 ), .B(\SUBBYTES[7].a/w688 ), .Z(
        \SUBBYTES[7].a/w692 ) );
  AND U3709 ( .A(\SUBBYTES[7].a/w689 ), .B(\SUBBYTES[7].a/w690 ), .Z(
        \SUBBYTES[7].a/w691 ) );
  AND U3710 ( .A(\SUBBYTES[7].a/w578 ), .B(n1630), .Z(\SUBBYTES[7].a/w677 ) );
  XOR U3711 ( .A(\SUBBYTES[7].a/w646 ), .B(n1055), .Z(n1630) );
  AND U3712 ( .A(\SUBBYTES[7].a/w579 ), .B(n1631), .Z(\SUBBYTES[7].a/w675 ) );
  XOR U3713 ( .A(n13517), .B(\SUBBYTES[7].a/w646 ), .Z(n1631) );
  ANDN U3714 ( .A(n1632), .B(n1636), .Z(\SUBBYTES[7].a/w674 ) );
  XOR U3715 ( .A(n1055), .B(n13517), .Z(n1632) );
  ANDN U3716 ( .A(\SUBBYTES[7].a/w580 ), .B(n1633), .Z(\SUBBYTES[7].a/w670 )
         );
  XNOR U3717 ( .A(\SUBBYTES[7].a/w639 ), .B(\SUBBYTES[7].a/w642 ), .Z(n1633)
         );
  AND U3718 ( .A(\SUBBYTES[7].a/w581 ), .B(n1634), .Z(\SUBBYTES[7].a/w668 ) );
  XNOR U3719 ( .A(n1637), .B(\SUBBYTES[7].a/w639 ), .Z(n1634) );
  AND U3720 ( .A(\SUBBYTES[7].a/w666 ), .B(n1638), .Z(\SUBBYTES[7].a/w667 ) );
  XOR U3721 ( .A(n1639), .B(n1637), .Z(n1638) );
  IV U3722 ( .A(n13516), .Z(n1637) );
  ANDN U3723 ( .A(\SUBBYTES[7].a/w685 ), .B(n1640), .Z(\SUBBYTES[7].a/w662 )
         );
  ANDN U3724 ( .A(\SUBBYTES[7].a/w686 ), .B(n1641), .Z(\SUBBYTES[7].a/w660 )
         );
  ANDN U3725 ( .A(\SUBBYTES[7].a/w689 ), .B(n1642), .Z(\SUBBYTES[7].a/w659 )
         );
  AND U3726 ( .A(\SUBBYTES[7].a/w645 ), .B(\SUBBYTES[7].a/w644 ), .Z(
        \SUBBYTES[7].a/w646 ) );
  IV U3727 ( .A(n1639), .Z(\SUBBYTES[7].a/w642 ) );
  NAND U3728 ( .A(\SUBBYTES[7].a/w621 ), .B(\SUBBYTES[7].a/w636 ), .Z(n1639)
         );
  AND U3729 ( .A(\SUBBYTES[7].a/w638 ), .B(\SUBBYTES[7].a/w644 ), .Z(
        \SUBBYTES[7].a/w639 ) );
  AND U3730 ( .A(\SUBBYTES[7].a/w623 ), .B(\SUBBYTES[7].a/w621 ), .Z(
        \SUBBYTES[7].a/w633 ) );
  AND U3731 ( .A(\SUBBYTES[7].a/w624 ), .B(\SUBBYTES[7].a/w622 ), .Z(
        \SUBBYTES[7].a/w631 ) );
  AND U3732 ( .A(\SUBBYTES[7].a/w638 ), .B(\SUBBYTES[7].a/w645 ), .Z(
        \SUBBYTES[7].a/w630 ) );
  AND U3733 ( .A(\SUBBYTES[7].a/w578 ), .B(\SUBBYTES[7].a/w574 ), .Z(
        \SUBBYTES[7].a/w615 ) );
  AND U3734 ( .A(\SUBBYTES[7].a/w579 ), .B(\SUBBYTES[7].a/w575 ), .Z(
        \SUBBYTES[7].a/w613 ) );
  ANDN U3735 ( .A(\SUBBYTES[7].a/w705 ), .B(n1636), .Z(\SUBBYTES[7].a/w612 )
         );
  XNOR U3736 ( .A(\w1[7][105] ), .B(\w1[7][111] ), .Z(n1636) );
  XOR U3737 ( .A(\w0[7][105] ), .B(g_input[1001]), .Z(\w1[7][105] ) );
  AND U3738 ( .A(\w1[7][104] ), .B(\SUBBYTES[7].a/w580 ), .Z(
        \SUBBYTES[7].a/w608 ) );
  XOR U3739 ( .A(\w0[7][104] ), .B(g_input[1000]), .Z(\w1[7][104] ) );
  AND U3740 ( .A(\SUBBYTES[7].a/w581 ), .B(\SUBBYTES[7].a/w577 ), .Z(
        \SUBBYTES[7].a/w606 ) );
  AND U3741 ( .A(\SUBBYTES[7].a/w666 ), .B(\SUBBYTES[7].a/w698 ), .Z(
        \SUBBYTES[7].a/w605 ) );
  ANDN U3742 ( .A(\SUBBYTES[7].a/w687 ), .B(n1640), .Z(\SUBBYTES[7].a/w600 )
         );
  XNOR U3743 ( .A(\w1[7][108] ), .B(\w1[7][111] ), .Z(n1640) );
  ANDN U3744 ( .A(\SUBBYTES[7].a/w688 ), .B(n1641), .Z(\SUBBYTES[7].a/w598 )
         );
  XNOR U3745 ( .A(\w1[7][106] ), .B(\w1[7][111] ), .Z(n1641) );
  XOR U3746 ( .A(\w0[7][111] ), .B(g_input[1007]), .Z(\w1[7][111] ) );
  IV U3747 ( .A(n1643), .Z(\w1[7][106] ) );
  ANDN U3748 ( .A(\SUBBYTES[7].a/w690 ), .B(n1642), .Z(\SUBBYTES[7].a/w597 )
         );
  XOR U3749 ( .A(n1643), .B(\w1[7][108] ), .Z(n1642) );
  XOR U3750 ( .A(\w0[7][108] ), .B(g_input[1004]), .Z(\w1[7][108] ) );
  XNOR U3751 ( .A(\w0[7][106] ), .B(g_input[1002]), .Z(n1643) );
  AND U3752 ( .A(n1644), .B(\SUBBYTES[7].a/w367 ), .Z(\SUBBYTES[7].a/w502 ) );
  AND U3753 ( .A(n1645), .B(\SUBBYTES[7].a/w368 ), .Z(\SUBBYTES[7].a/w500 ) );
  AND U3754 ( .A(\SUBBYTES[7].a/w498 ), .B(n1646), .Z(\SUBBYTES[7].a/w499 ) );
  ANDN U3755 ( .A(\w1[7][112] ), .B(n1647), .Z(\SUBBYTES[7].a/w495 ) );
  AND U3756 ( .A(n1648), .B(\SUBBYTES[7].a/w370 ), .Z(\SUBBYTES[7].a/w493 ) );
  AND U3757 ( .A(\SUBBYTES[7].a/w491 ), .B(n1649), .Z(\SUBBYTES[7].a/w492 ) );
  XOR U3758 ( .A(\SUBBYTES[7].a/w435 ), .B(n13514), .Z(n1649) );
  AND U3759 ( .A(\SUBBYTES[7].a/w478 ), .B(\SUBBYTES[7].a/w480 ), .Z(
        \SUBBYTES[7].a/w487 ) );
  AND U3760 ( .A(\SUBBYTES[7].a/w479 ), .B(\SUBBYTES[7].a/w481 ), .Z(
        \SUBBYTES[7].a/w485 ) );
  AND U3761 ( .A(\SUBBYTES[7].a/w482 ), .B(\SUBBYTES[7].a/w483 ), .Z(
        \SUBBYTES[7].a/w484 ) );
  AND U3762 ( .A(\SUBBYTES[7].a/w371 ), .B(n1644), .Z(\SUBBYTES[7].a/w470 ) );
  XOR U3763 ( .A(\SUBBYTES[7].a/w439 ), .B(n1054), .Z(n1644) );
  AND U3764 ( .A(\SUBBYTES[7].a/w372 ), .B(n1645), .Z(\SUBBYTES[7].a/w468 ) );
  XOR U3765 ( .A(n13515), .B(\SUBBYTES[7].a/w439 ), .Z(n1645) );
  ANDN U3766 ( .A(n1646), .B(n1650), .Z(\SUBBYTES[7].a/w467 ) );
  XOR U3767 ( .A(n1054), .B(n13515), .Z(n1646) );
  ANDN U3768 ( .A(\SUBBYTES[7].a/w373 ), .B(n1647), .Z(\SUBBYTES[7].a/w463 )
         );
  XNOR U3769 ( .A(\SUBBYTES[7].a/w432 ), .B(\SUBBYTES[7].a/w435 ), .Z(n1647)
         );
  AND U3770 ( .A(\SUBBYTES[7].a/w374 ), .B(n1648), .Z(\SUBBYTES[7].a/w461 ) );
  XNOR U3771 ( .A(n1651), .B(\SUBBYTES[7].a/w432 ), .Z(n1648) );
  AND U3772 ( .A(\SUBBYTES[7].a/w459 ), .B(n1652), .Z(\SUBBYTES[7].a/w460 ) );
  XOR U3773 ( .A(n1653), .B(n1651), .Z(n1652) );
  IV U3774 ( .A(n13514), .Z(n1651) );
  ANDN U3775 ( .A(\SUBBYTES[7].a/w478 ), .B(n1654), .Z(\SUBBYTES[7].a/w455 )
         );
  ANDN U3776 ( .A(\SUBBYTES[7].a/w479 ), .B(n1655), .Z(\SUBBYTES[7].a/w453 )
         );
  ANDN U3777 ( .A(\SUBBYTES[7].a/w482 ), .B(n1656), .Z(\SUBBYTES[7].a/w452 )
         );
  AND U3778 ( .A(\SUBBYTES[7].a/w438 ), .B(\SUBBYTES[7].a/w437 ), .Z(
        \SUBBYTES[7].a/w439 ) );
  IV U3779 ( .A(n1653), .Z(\SUBBYTES[7].a/w435 ) );
  NAND U3780 ( .A(\SUBBYTES[7].a/w414 ), .B(\SUBBYTES[7].a/w429 ), .Z(n1653)
         );
  AND U3781 ( .A(\SUBBYTES[7].a/w431 ), .B(\SUBBYTES[7].a/w437 ), .Z(
        \SUBBYTES[7].a/w432 ) );
  AND U3782 ( .A(\SUBBYTES[7].a/w416 ), .B(\SUBBYTES[7].a/w414 ), .Z(
        \SUBBYTES[7].a/w426 ) );
  AND U3783 ( .A(\SUBBYTES[7].a/w417 ), .B(\SUBBYTES[7].a/w415 ), .Z(
        \SUBBYTES[7].a/w424 ) );
  AND U3784 ( .A(\SUBBYTES[7].a/w431 ), .B(\SUBBYTES[7].a/w438 ), .Z(
        \SUBBYTES[7].a/w423 ) );
  AND U3785 ( .A(\SUBBYTES[7].a/w371 ), .B(\SUBBYTES[7].a/w367 ), .Z(
        \SUBBYTES[7].a/w408 ) );
  AND U3786 ( .A(\SUBBYTES[7].a/w372 ), .B(\SUBBYTES[7].a/w368 ), .Z(
        \SUBBYTES[7].a/w406 ) );
  ANDN U3787 ( .A(\SUBBYTES[7].a/w498 ), .B(n1650), .Z(\SUBBYTES[7].a/w405 )
         );
  XNOR U3788 ( .A(\w1[7][113] ), .B(\w1[7][119] ), .Z(n1650) );
  XOR U3789 ( .A(\w0[7][113] ), .B(g_input[1009]), .Z(\w1[7][113] ) );
  AND U3790 ( .A(\w1[7][112] ), .B(\SUBBYTES[7].a/w373 ), .Z(
        \SUBBYTES[7].a/w401 ) );
  XOR U3791 ( .A(\w0[7][112] ), .B(g_input[1008]), .Z(\w1[7][112] ) );
  AND U3792 ( .A(\SUBBYTES[7].a/w374 ), .B(\SUBBYTES[7].a/w370 ), .Z(
        \SUBBYTES[7].a/w399 ) );
  AND U3793 ( .A(\SUBBYTES[7].a/w459 ), .B(\SUBBYTES[7].a/w491 ), .Z(
        \SUBBYTES[7].a/w398 ) );
  ANDN U3794 ( .A(\SUBBYTES[7].a/w480 ), .B(n1654), .Z(\SUBBYTES[7].a/w393 )
         );
  XNOR U3795 ( .A(\w1[7][116] ), .B(\w1[7][119] ), .Z(n1654) );
  ANDN U3796 ( .A(\SUBBYTES[7].a/w481 ), .B(n1655), .Z(\SUBBYTES[7].a/w391 )
         );
  XNOR U3797 ( .A(\w1[7][114] ), .B(\w1[7][119] ), .Z(n1655) );
  XOR U3798 ( .A(\w0[7][119] ), .B(g_input[1015]), .Z(\w1[7][119] ) );
  IV U3799 ( .A(n1657), .Z(\w1[7][114] ) );
  ANDN U3800 ( .A(\SUBBYTES[7].a/w483 ), .B(n1656), .Z(\SUBBYTES[7].a/w390 )
         );
  XOR U3801 ( .A(n1657), .B(\w1[7][116] ), .Z(n1656) );
  XOR U3802 ( .A(\w0[7][116] ), .B(g_input[1012]), .Z(\w1[7][116] ) );
  XNOR U3803 ( .A(\w0[7][114] ), .B(g_input[1010]), .Z(n1657) );
  AND U3804 ( .A(n1658), .B(\SUBBYTES[7].a/w3265 ), .Z(\SUBBYTES[7].a/w3400 )
         );
  AND U3805 ( .A(n1659), .B(\SUBBYTES[7].a/w3266 ), .Z(\SUBBYTES[7].a/w3398 )
         );
  AND U3806 ( .A(\SUBBYTES[7].a/w3396 ), .B(n1660), .Z(\SUBBYTES[7].a/w3397 )
         );
  ANDN U3807 ( .A(\w1[7][0] ), .B(n1661), .Z(\SUBBYTES[7].a/w3393 ) );
  AND U3808 ( .A(n1662), .B(\SUBBYTES[7].a/w3268 ), .Z(\SUBBYTES[7].a/w3391 )
         );
  AND U3809 ( .A(\SUBBYTES[7].a/w3389 ), .B(n1663), .Z(\SUBBYTES[7].a/w3390 )
         );
  XOR U3810 ( .A(\SUBBYTES[7].a/w3333 ), .B(n13542), .Z(n1663) );
  AND U3811 ( .A(\SUBBYTES[7].a/w3376 ), .B(\SUBBYTES[7].a/w3378 ), .Z(
        \SUBBYTES[7].a/w3385 ) );
  AND U3812 ( .A(\SUBBYTES[7].a/w3377 ), .B(\SUBBYTES[7].a/w3379 ), .Z(
        \SUBBYTES[7].a/w3383 ) );
  AND U3813 ( .A(\SUBBYTES[7].a/w3380 ), .B(\SUBBYTES[7].a/w3381 ), .Z(
        \SUBBYTES[7].a/w3382 ) );
  AND U3814 ( .A(\SUBBYTES[7].a/w3269 ), .B(n1658), .Z(\SUBBYTES[7].a/w3368 )
         );
  XOR U3815 ( .A(\SUBBYTES[7].a/w3337 ), .B(n1068), .Z(n1658) );
  AND U3816 ( .A(\SUBBYTES[7].a/w3270 ), .B(n1659), .Z(\SUBBYTES[7].a/w3366 )
         );
  XOR U3817 ( .A(n13543), .B(\SUBBYTES[7].a/w3337 ), .Z(n1659) );
  ANDN U3818 ( .A(n1660), .B(n1664), .Z(\SUBBYTES[7].a/w3365 ) );
  XOR U3819 ( .A(n1068), .B(n13543), .Z(n1660) );
  ANDN U3820 ( .A(\SUBBYTES[7].a/w3271 ), .B(n1661), .Z(\SUBBYTES[7].a/w3361 )
         );
  XNOR U3821 ( .A(\SUBBYTES[7].a/w3330 ), .B(\SUBBYTES[7].a/w3333 ), .Z(n1661)
         );
  AND U3822 ( .A(\SUBBYTES[7].a/w3272 ), .B(n1662), .Z(\SUBBYTES[7].a/w3359 )
         );
  XNOR U3823 ( .A(n1665), .B(\SUBBYTES[7].a/w3330 ), .Z(n1662) );
  AND U3824 ( .A(\SUBBYTES[7].a/w3357 ), .B(n1666), .Z(\SUBBYTES[7].a/w3358 )
         );
  XOR U3825 ( .A(n1667), .B(n1665), .Z(n1666) );
  IV U3826 ( .A(n13542), .Z(n1665) );
  ANDN U3827 ( .A(\SUBBYTES[7].a/w3376 ), .B(n1668), .Z(\SUBBYTES[7].a/w3353 )
         );
  ANDN U3828 ( .A(\SUBBYTES[7].a/w3377 ), .B(n1669), .Z(\SUBBYTES[7].a/w3351 )
         );
  ANDN U3829 ( .A(\SUBBYTES[7].a/w3380 ), .B(n1670), .Z(\SUBBYTES[7].a/w3350 )
         );
  AND U3830 ( .A(\SUBBYTES[7].a/w3336 ), .B(\SUBBYTES[7].a/w3335 ), .Z(
        \SUBBYTES[7].a/w3337 ) );
  IV U3831 ( .A(n1667), .Z(\SUBBYTES[7].a/w3333 ) );
  NAND U3832 ( .A(\SUBBYTES[7].a/w3312 ), .B(\SUBBYTES[7].a/w3327 ), .Z(n1667)
         );
  AND U3833 ( .A(\SUBBYTES[7].a/w3329 ), .B(\SUBBYTES[7].a/w3335 ), .Z(
        \SUBBYTES[7].a/w3330 ) );
  AND U3834 ( .A(\SUBBYTES[7].a/w3314 ), .B(\SUBBYTES[7].a/w3312 ), .Z(
        \SUBBYTES[7].a/w3324 ) );
  AND U3835 ( .A(\SUBBYTES[7].a/w3315 ), .B(\SUBBYTES[7].a/w3313 ), .Z(
        \SUBBYTES[7].a/w3322 ) );
  AND U3836 ( .A(\SUBBYTES[7].a/w3329 ), .B(\SUBBYTES[7].a/w3336 ), .Z(
        \SUBBYTES[7].a/w3321 ) );
  AND U3837 ( .A(\SUBBYTES[7].a/w3269 ), .B(\SUBBYTES[7].a/w3265 ), .Z(
        \SUBBYTES[7].a/w3306 ) );
  AND U3838 ( .A(\SUBBYTES[7].a/w3270 ), .B(\SUBBYTES[7].a/w3266 ), .Z(
        \SUBBYTES[7].a/w3304 ) );
  ANDN U3839 ( .A(\SUBBYTES[7].a/w3396 ), .B(n1664), .Z(\SUBBYTES[7].a/w3303 )
         );
  XNOR U3840 ( .A(\w1[7][1] ), .B(\w1[7][7] ), .Z(n1664) );
  XOR U3841 ( .A(\w0[7][1] ), .B(g_input[897]), .Z(\w1[7][1] ) );
  AND U3842 ( .A(\w1[7][0] ), .B(\SUBBYTES[7].a/w3271 ), .Z(
        \SUBBYTES[7].a/w3299 ) );
  XOR U3843 ( .A(\w0[7][0] ), .B(g_input[896]), .Z(\w1[7][0] ) );
  AND U3844 ( .A(\SUBBYTES[7].a/w3272 ), .B(\SUBBYTES[7].a/w3268 ), .Z(
        \SUBBYTES[7].a/w3297 ) );
  AND U3845 ( .A(\SUBBYTES[7].a/w3357 ), .B(\SUBBYTES[7].a/w3389 ), .Z(
        \SUBBYTES[7].a/w3296 ) );
  ANDN U3846 ( .A(\SUBBYTES[7].a/w3378 ), .B(n1668), .Z(\SUBBYTES[7].a/w3291 )
         );
  XNOR U3847 ( .A(\w1[7][4] ), .B(\w1[7][7] ), .Z(n1668) );
  ANDN U3848 ( .A(\SUBBYTES[7].a/w3379 ), .B(n1669), .Z(\SUBBYTES[7].a/w3289 )
         );
  XNOR U3849 ( .A(\w1[7][2] ), .B(\w1[7][7] ), .Z(n1669) );
  XOR U3850 ( .A(\w0[7][7] ), .B(g_input[903]), .Z(\w1[7][7] ) );
  IV U3851 ( .A(n1671), .Z(\w1[7][2] ) );
  ANDN U3852 ( .A(\SUBBYTES[7].a/w3381 ), .B(n1670), .Z(\SUBBYTES[7].a/w3288 )
         );
  XOR U3853 ( .A(n1671), .B(\w1[7][4] ), .Z(n1670) );
  XOR U3854 ( .A(\w0[7][4] ), .B(g_input[900]), .Z(\w1[7][4] ) );
  XNOR U3855 ( .A(\w0[7][2] ), .B(g_input[898]), .Z(n1671) );
  AND U3856 ( .A(n1672), .B(\SUBBYTES[7].a/w3058 ), .Z(\SUBBYTES[7].a/w3193 )
         );
  AND U3857 ( .A(n1673), .B(\SUBBYTES[7].a/w3059 ), .Z(\SUBBYTES[7].a/w3191 )
         );
  AND U3858 ( .A(\SUBBYTES[7].a/w3189 ), .B(n1674), .Z(\SUBBYTES[7].a/w3190 )
         );
  ANDN U3859 ( .A(\w1[7][8] ), .B(n1675), .Z(\SUBBYTES[7].a/w3186 ) );
  AND U3860 ( .A(n1676), .B(\SUBBYTES[7].a/w3061 ), .Z(\SUBBYTES[7].a/w3184 )
         );
  AND U3861 ( .A(\SUBBYTES[7].a/w3182 ), .B(n1677), .Z(\SUBBYTES[7].a/w3183 )
         );
  XOR U3862 ( .A(\SUBBYTES[7].a/w3126 ), .B(n13540), .Z(n1677) );
  AND U3863 ( .A(\SUBBYTES[7].a/w3169 ), .B(\SUBBYTES[7].a/w3171 ), .Z(
        \SUBBYTES[7].a/w3178 ) );
  AND U3864 ( .A(\SUBBYTES[7].a/w3170 ), .B(\SUBBYTES[7].a/w3172 ), .Z(
        \SUBBYTES[7].a/w3176 ) );
  AND U3865 ( .A(\SUBBYTES[7].a/w3173 ), .B(\SUBBYTES[7].a/w3174 ), .Z(
        \SUBBYTES[7].a/w3175 ) );
  AND U3866 ( .A(\SUBBYTES[7].a/w3062 ), .B(n1672), .Z(\SUBBYTES[7].a/w3161 )
         );
  XOR U3867 ( .A(\SUBBYTES[7].a/w3130 ), .B(n1067), .Z(n1672) );
  AND U3868 ( .A(\SUBBYTES[7].a/w3063 ), .B(n1673), .Z(\SUBBYTES[7].a/w3159 )
         );
  XOR U3869 ( .A(n13541), .B(\SUBBYTES[7].a/w3130 ), .Z(n1673) );
  ANDN U3870 ( .A(n1674), .B(n1678), .Z(\SUBBYTES[7].a/w3158 ) );
  XOR U3871 ( .A(n1067), .B(n13541), .Z(n1674) );
  ANDN U3872 ( .A(\SUBBYTES[7].a/w3064 ), .B(n1675), .Z(\SUBBYTES[7].a/w3154 )
         );
  XNOR U3873 ( .A(\SUBBYTES[7].a/w3123 ), .B(\SUBBYTES[7].a/w3126 ), .Z(n1675)
         );
  AND U3874 ( .A(\SUBBYTES[7].a/w3065 ), .B(n1676), .Z(\SUBBYTES[7].a/w3152 )
         );
  XNOR U3875 ( .A(n1679), .B(\SUBBYTES[7].a/w3123 ), .Z(n1676) );
  AND U3876 ( .A(\SUBBYTES[7].a/w3150 ), .B(n1680), .Z(\SUBBYTES[7].a/w3151 )
         );
  XOR U3877 ( .A(n1681), .B(n1679), .Z(n1680) );
  IV U3878 ( .A(n13540), .Z(n1679) );
  ANDN U3879 ( .A(\SUBBYTES[7].a/w3169 ), .B(n1682), .Z(\SUBBYTES[7].a/w3146 )
         );
  ANDN U3880 ( .A(\SUBBYTES[7].a/w3170 ), .B(n1683), .Z(\SUBBYTES[7].a/w3144 )
         );
  ANDN U3881 ( .A(\SUBBYTES[7].a/w3173 ), .B(n1684), .Z(\SUBBYTES[7].a/w3143 )
         );
  AND U3882 ( .A(\SUBBYTES[7].a/w3129 ), .B(\SUBBYTES[7].a/w3128 ), .Z(
        \SUBBYTES[7].a/w3130 ) );
  IV U3883 ( .A(n1681), .Z(\SUBBYTES[7].a/w3126 ) );
  NAND U3884 ( .A(\SUBBYTES[7].a/w3105 ), .B(\SUBBYTES[7].a/w3120 ), .Z(n1681)
         );
  AND U3885 ( .A(\SUBBYTES[7].a/w3122 ), .B(\SUBBYTES[7].a/w3128 ), .Z(
        \SUBBYTES[7].a/w3123 ) );
  AND U3886 ( .A(\SUBBYTES[7].a/w3107 ), .B(\SUBBYTES[7].a/w3105 ), .Z(
        \SUBBYTES[7].a/w3117 ) );
  AND U3887 ( .A(\SUBBYTES[7].a/w3108 ), .B(\SUBBYTES[7].a/w3106 ), .Z(
        \SUBBYTES[7].a/w3115 ) );
  AND U3888 ( .A(\SUBBYTES[7].a/w3122 ), .B(\SUBBYTES[7].a/w3129 ), .Z(
        \SUBBYTES[7].a/w3114 ) );
  AND U3889 ( .A(\SUBBYTES[7].a/w3062 ), .B(\SUBBYTES[7].a/w3058 ), .Z(
        \SUBBYTES[7].a/w3099 ) );
  AND U3890 ( .A(\SUBBYTES[7].a/w3063 ), .B(\SUBBYTES[7].a/w3059 ), .Z(
        \SUBBYTES[7].a/w3097 ) );
  ANDN U3891 ( .A(\SUBBYTES[7].a/w3189 ), .B(n1678), .Z(\SUBBYTES[7].a/w3096 )
         );
  XNOR U3892 ( .A(\w1[7][15] ), .B(\w1[7][9] ), .Z(n1678) );
  XOR U3893 ( .A(\w0[7][9] ), .B(g_input[905]), .Z(\w1[7][9] ) );
  AND U3894 ( .A(\w1[7][8] ), .B(\SUBBYTES[7].a/w3064 ), .Z(
        \SUBBYTES[7].a/w3092 ) );
  XOR U3895 ( .A(\w0[7][8] ), .B(g_input[904]), .Z(\w1[7][8] ) );
  AND U3896 ( .A(\SUBBYTES[7].a/w3065 ), .B(\SUBBYTES[7].a/w3061 ), .Z(
        \SUBBYTES[7].a/w3090 ) );
  AND U3897 ( .A(\SUBBYTES[7].a/w3150 ), .B(\SUBBYTES[7].a/w3182 ), .Z(
        \SUBBYTES[7].a/w3089 ) );
  ANDN U3898 ( .A(\SUBBYTES[7].a/w3171 ), .B(n1682), .Z(\SUBBYTES[7].a/w3084 )
         );
  XNOR U3899 ( .A(\w1[7][12] ), .B(\w1[7][15] ), .Z(n1682) );
  ANDN U3900 ( .A(\SUBBYTES[7].a/w3172 ), .B(n1683), .Z(\SUBBYTES[7].a/w3082 )
         );
  XNOR U3901 ( .A(\w1[7][10] ), .B(\w1[7][15] ), .Z(n1683) );
  XOR U3902 ( .A(\w0[7][15] ), .B(g_input[911]), .Z(\w1[7][15] ) );
  ANDN U3903 ( .A(\SUBBYTES[7].a/w3174 ), .B(n1684), .Z(\SUBBYTES[7].a/w3081 )
         );
  XNOR U3904 ( .A(\w1[7][10] ), .B(\w1[7][12] ), .Z(n1684) );
  XOR U3905 ( .A(\w0[7][12] ), .B(g_input[908]), .Z(\w1[7][12] ) );
  XOR U3906 ( .A(\w0[7][10] ), .B(g_input[906]), .Z(\w1[7][10] ) );
  AND U3907 ( .A(n1685), .B(\SUBBYTES[7].a/w2851 ), .Z(\SUBBYTES[7].a/w2986 )
         );
  AND U3908 ( .A(n1686), .B(\SUBBYTES[7].a/w2852 ), .Z(\SUBBYTES[7].a/w2984 )
         );
  AND U3909 ( .A(\SUBBYTES[7].a/w2982 ), .B(n1687), .Z(\SUBBYTES[7].a/w2983 )
         );
  ANDN U3910 ( .A(\w1[7][16] ), .B(n1688), .Z(\SUBBYTES[7].a/w2979 ) );
  AND U3911 ( .A(n1689), .B(\SUBBYTES[7].a/w2854 ), .Z(\SUBBYTES[7].a/w2977 )
         );
  AND U3912 ( .A(\SUBBYTES[7].a/w2975 ), .B(n1690), .Z(\SUBBYTES[7].a/w2976 )
         );
  XOR U3913 ( .A(\SUBBYTES[7].a/w2919 ), .B(n13538), .Z(n1690) );
  AND U3914 ( .A(\SUBBYTES[7].a/w2962 ), .B(\SUBBYTES[7].a/w2964 ), .Z(
        \SUBBYTES[7].a/w2971 ) );
  AND U3915 ( .A(\SUBBYTES[7].a/w2963 ), .B(\SUBBYTES[7].a/w2965 ), .Z(
        \SUBBYTES[7].a/w2969 ) );
  AND U3916 ( .A(\SUBBYTES[7].a/w2966 ), .B(\SUBBYTES[7].a/w2967 ), .Z(
        \SUBBYTES[7].a/w2968 ) );
  AND U3917 ( .A(\SUBBYTES[7].a/w2855 ), .B(n1685), .Z(\SUBBYTES[7].a/w2954 )
         );
  XOR U3918 ( .A(\SUBBYTES[7].a/w2923 ), .B(n1066), .Z(n1685) );
  AND U3919 ( .A(\SUBBYTES[7].a/w2856 ), .B(n1686), .Z(\SUBBYTES[7].a/w2952 )
         );
  XOR U3920 ( .A(n13539), .B(\SUBBYTES[7].a/w2923 ), .Z(n1686) );
  ANDN U3921 ( .A(n1687), .B(n1691), .Z(\SUBBYTES[7].a/w2951 ) );
  XOR U3922 ( .A(n1066), .B(n13539), .Z(n1687) );
  AND U3923 ( .A(n1692), .B(\SUBBYTES[7].a/w160 ), .Z(\SUBBYTES[7].a/w295 ) );
  ANDN U3924 ( .A(\SUBBYTES[7].a/w2857 ), .B(n1688), .Z(\SUBBYTES[7].a/w2947 )
         );
  XNOR U3925 ( .A(\SUBBYTES[7].a/w2916 ), .B(\SUBBYTES[7].a/w2919 ), .Z(n1688)
         );
  AND U3926 ( .A(\SUBBYTES[7].a/w2858 ), .B(n1689), .Z(\SUBBYTES[7].a/w2945 )
         );
  XNOR U3927 ( .A(n1693), .B(\SUBBYTES[7].a/w2916 ), .Z(n1689) );
  AND U3928 ( .A(\SUBBYTES[7].a/w2943 ), .B(n1694), .Z(\SUBBYTES[7].a/w2944 )
         );
  XOR U3929 ( .A(n1695), .B(n1693), .Z(n1694) );
  IV U3930 ( .A(n13538), .Z(n1693) );
  ANDN U3931 ( .A(\SUBBYTES[7].a/w2962 ), .B(n1696), .Z(\SUBBYTES[7].a/w2939 )
         );
  ANDN U3932 ( .A(\SUBBYTES[7].a/w2963 ), .B(n1697), .Z(\SUBBYTES[7].a/w2937 )
         );
  ANDN U3933 ( .A(\SUBBYTES[7].a/w2966 ), .B(n1698), .Z(\SUBBYTES[7].a/w2936 )
         );
  AND U3934 ( .A(n1699), .B(\SUBBYTES[7].a/w161 ), .Z(\SUBBYTES[7].a/w293 ) );
  AND U3935 ( .A(\SUBBYTES[7].a/w2922 ), .B(\SUBBYTES[7].a/w2921 ), .Z(
        \SUBBYTES[7].a/w2923 ) );
  AND U3936 ( .A(\SUBBYTES[7].a/w291 ), .B(n1700), .Z(\SUBBYTES[7].a/w292 ) );
  IV U3937 ( .A(n1695), .Z(\SUBBYTES[7].a/w2919 ) );
  NAND U3938 ( .A(\SUBBYTES[7].a/w2898 ), .B(\SUBBYTES[7].a/w2913 ), .Z(n1695)
         );
  AND U3939 ( .A(\SUBBYTES[7].a/w2915 ), .B(\SUBBYTES[7].a/w2921 ), .Z(
        \SUBBYTES[7].a/w2916 ) );
  AND U3940 ( .A(\SUBBYTES[7].a/w2900 ), .B(\SUBBYTES[7].a/w2898 ), .Z(
        \SUBBYTES[7].a/w2910 ) );
  AND U3941 ( .A(\SUBBYTES[7].a/w2901 ), .B(\SUBBYTES[7].a/w2899 ), .Z(
        \SUBBYTES[7].a/w2908 ) );
  AND U3942 ( .A(\SUBBYTES[7].a/w2915 ), .B(\SUBBYTES[7].a/w2922 ), .Z(
        \SUBBYTES[7].a/w2907 ) );
  AND U3943 ( .A(\SUBBYTES[7].a/w2855 ), .B(\SUBBYTES[7].a/w2851 ), .Z(
        \SUBBYTES[7].a/w2892 ) );
  AND U3944 ( .A(\SUBBYTES[7].a/w2856 ), .B(\SUBBYTES[7].a/w2852 ), .Z(
        \SUBBYTES[7].a/w2890 ) );
  ANDN U3945 ( .A(\SUBBYTES[7].a/w2982 ), .B(n1691), .Z(\SUBBYTES[7].a/w2889 )
         );
  XNOR U3946 ( .A(\w1[7][17] ), .B(\w1[7][23] ), .Z(n1691) );
  XOR U3947 ( .A(\w0[7][17] ), .B(g_input[913]), .Z(\w1[7][17] ) );
  AND U3948 ( .A(\w1[7][16] ), .B(\SUBBYTES[7].a/w2857 ), .Z(
        \SUBBYTES[7].a/w2885 ) );
  XOR U3949 ( .A(\w0[7][16] ), .B(g_input[912]), .Z(\w1[7][16] ) );
  AND U3950 ( .A(\SUBBYTES[7].a/w2858 ), .B(\SUBBYTES[7].a/w2854 ), .Z(
        \SUBBYTES[7].a/w2883 ) );
  AND U3951 ( .A(\SUBBYTES[7].a/w2943 ), .B(\SUBBYTES[7].a/w2975 ), .Z(
        \SUBBYTES[7].a/w2882 ) );
  ANDN U3952 ( .A(\w1[7][120] ), .B(n1701), .Z(\SUBBYTES[7].a/w288 ) );
  ANDN U3953 ( .A(\SUBBYTES[7].a/w2964 ), .B(n1696), .Z(\SUBBYTES[7].a/w2877 )
         );
  XNOR U3954 ( .A(\w1[7][20] ), .B(\w1[7][23] ), .Z(n1696) );
  ANDN U3955 ( .A(\SUBBYTES[7].a/w2965 ), .B(n1697), .Z(\SUBBYTES[7].a/w2875 )
         );
  XNOR U3956 ( .A(\w1[7][18] ), .B(\w1[7][23] ), .Z(n1697) );
  XOR U3957 ( .A(\w0[7][23] ), .B(g_input[919]), .Z(\w1[7][23] ) );
  IV U3958 ( .A(n1702), .Z(\w1[7][18] ) );
  ANDN U3959 ( .A(\SUBBYTES[7].a/w2967 ), .B(n1698), .Z(\SUBBYTES[7].a/w2874 )
         );
  XOR U3960 ( .A(n1702), .B(\w1[7][20] ), .Z(n1698) );
  XOR U3961 ( .A(\w0[7][20] ), .B(g_input[916]), .Z(\w1[7][20] ) );
  XNOR U3962 ( .A(\w0[7][18] ), .B(g_input[914]), .Z(n1702) );
  AND U3963 ( .A(n1703), .B(\SUBBYTES[7].a/w163 ), .Z(\SUBBYTES[7].a/w286 ) );
  AND U3964 ( .A(\SUBBYTES[7].a/w284 ), .B(n1704), .Z(\SUBBYTES[7].a/w285 ) );
  XOR U3965 ( .A(\SUBBYTES[7].a/w228 ), .B(n13512), .Z(n1704) );
  AND U3966 ( .A(\SUBBYTES[7].a/w271 ), .B(\SUBBYTES[7].a/w273 ), .Z(
        \SUBBYTES[7].a/w280 ) );
  AND U3967 ( .A(\SUBBYTES[7].a/w272 ), .B(\SUBBYTES[7].a/w274 ), .Z(
        \SUBBYTES[7].a/w278 ) );
  AND U3968 ( .A(n1705), .B(\SUBBYTES[7].a/w2644 ), .Z(\SUBBYTES[7].a/w2779 )
         );
  AND U3969 ( .A(n1706), .B(\SUBBYTES[7].a/w2645 ), .Z(\SUBBYTES[7].a/w2777 )
         );
  AND U3970 ( .A(\SUBBYTES[7].a/w2775 ), .B(n1707), .Z(\SUBBYTES[7].a/w2776 )
         );
  ANDN U3971 ( .A(\w1[7][24] ), .B(n1708), .Z(\SUBBYTES[7].a/w2772 ) );
  AND U3972 ( .A(n1709), .B(\SUBBYTES[7].a/w2647 ), .Z(\SUBBYTES[7].a/w2770 )
         );
  AND U3973 ( .A(\SUBBYTES[7].a/w275 ), .B(\SUBBYTES[7].a/w276 ), .Z(
        \SUBBYTES[7].a/w277 ) );
  AND U3974 ( .A(\SUBBYTES[7].a/w2768 ), .B(n1710), .Z(\SUBBYTES[7].a/w2769 )
         );
  XOR U3975 ( .A(\SUBBYTES[7].a/w2712 ), .B(n13536), .Z(n1710) );
  AND U3976 ( .A(\SUBBYTES[7].a/w2755 ), .B(\SUBBYTES[7].a/w2757 ), .Z(
        \SUBBYTES[7].a/w2764 ) );
  AND U3977 ( .A(\SUBBYTES[7].a/w2756 ), .B(\SUBBYTES[7].a/w2758 ), .Z(
        \SUBBYTES[7].a/w2762 ) );
  AND U3978 ( .A(\SUBBYTES[7].a/w2759 ), .B(\SUBBYTES[7].a/w2760 ), .Z(
        \SUBBYTES[7].a/w2761 ) );
  AND U3979 ( .A(\SUBBYTES[7].a/w2648 ), .B(n1705), .Z(\SUBBYTES[7].a/w2747 )
         );
  XOR U3980 ( .A(\SUBBYTES[7].a/w2716 ), .B(n1065), .Z(n1705) );
  AND U3981 ( .A(\SUBBYTES[7].a/w2649 ), .B(n1706), .Z(\SUBBYTES[7].a/w2745 )
         );
  XOR U3982 ( .A(n13537), .B(\SUBBYTES[7].a/w2716 ), .Z(n1706) );
  ANDN U3983 ( .A(n1707), .B(n1711), .Z(\SUBBYTES[7].a/w2744 ) );
  XOR U3984 ( .A(n1065), .B(n13537), .Z(n1707) );
  ANDN U3985 ( .A(\SUBBYTES[7].a/w2650 ), .B(n1708), .Z(\SUBBYTES[7].a/w2740 )
         );
  XNOR U3986 ( .A(\SUBBYTES[7].a/w2709 ), .B(\SUBBYTES[7].a/w2712 ), .Z(n1708)
         );
  AND U3987 ( .A(\SUBBYTES[7].a/w2651 ), .B(n1709), .Z(\SUBBYTES[7].a/w2738 )
         );
  XNOR U3988 ( .A(n1712), .B(\SUBBYTES[7].a/w2709 ), .Z(n1709) );
  AND U3989 ( .A(\SUBBYTES[7].a/w2736 ), .B(n1713), .Z(\SUBBYTES[7].a/w2737 )
         );
  XOR U3990 ( .A(n1714), .B(n1712), .Z(n1713) );
  IV U3991 ( .A(n13536), .Z(n1712) );
  ANDN U3992 ( .A(\SUBBYTES[7].a/w2755 ), .B(n1715), .Z(\SUBBYTES[7].a/w2732 )
         );
  ANDN U3993 ( .A(\SUBBYTES[7].a/w2756 ), .B(n1716), .Z(\SUBBYTES[7].a/w2730 )
         );
  ANDN U3994 ( .A(\SUBBYTES[7].a/w2759 ), .B(n1717), .Z(\SUBBYTES[7].a/w2729 )
         );
  AND U3995 ( .A(\SUBBYTES[7].a/w2715 ), .B(\SUBBYTES[7].a/w2714 ), .Z(
        \SUBBYTES[7].a/w2716 ) );
  IV U3996 ( .A(n1714), .Z(\SUBBYTES[7].a/w2712 ) );
  NAND U3997 ( .A(\SUBBYTES[7].a/w2691 ), .B(\SUBBYTES[7].a/w2706 ), .Z(n1714)
         );
  AND U3998 ( .A(\SUBBYTES[7].a/w2708 ), .B(\SUBBYTES[7].a/w2714 ), .Z(
        \SUBBYTES[7].a/w2709 ) );
  AND U3999 ( .A(\SUBBYTES[7].a/w2693 ), .B(\SUBBYTES[7].a/w2691 ), .Z(
        \SUBBYTES[7].a/w2703 ) );
  AND U4000 ( .A(\SUBBYTES[7].a/w2694 ), .B(\SUBBYTES[7].a/w2692 ), .Z(
        \SUBBYTES[7].a/w2701 ) );
  AND U4001 ( .A(\SUBBYTES[7].a/w2708 ), .B(\SUBBYTES[7].a/w2715 ), .Z(
        \SUBBYTES[7].a/w2700 ) );
  AND U4002 ( .A(\SUBBYTES[7].a/w2648 ), .B(\SUBBYTES[7].a/w2644 ), .Z(
        \SUBBYTES[7].a/w2685 ) );
  AND U4003 ( .A(\SUBBYTES[7].a/w2649 ), .B(\SUBBYTES[7].a/w2645 ), .Z(
        \SUBBYTES[7].a/w2683 ) );
  ANDN U4004 ( .A(\SUBBYTES[7].a/w2775 ), .B(n1711), .Z(\SUBBYTES[7].a/w2682 )
         );
  XNOR U4005 ( .A(\w1[7][25] ), .B(\w1[7][31] ), .Z(n1711) );
  XOR U4006 ( .A(\w0[7][25] ), .B(g_input[921]), .Z(\w1[7][25] ) );
  AND U4007 ( .A(\w1[7][24] ), .B(\SUBBYTES[7].a/w2650 ), .Z(
        \SUBBYTES[7].a/w2678 ) );
  XOR U4008 ( .A(\w0[7][24] ), .B(g_input[920]), .Z(\w1[7][24] ) );
  AND U4009 ( .A(\SUBBYTES[7].a/w2651 ), .B(\SUBBYTES[7].a/w2647 ), .Z(
        \SUBBYTES[7].a/w2676 ) );
  AND U4010 ( .A(\SUBBYTES[7].a/w2736 ), .B(\SUBBYTES[7].a/w2768 ), .Z(
        \SUBBYTES[7].a/w2675 ) );
  ANDN U4011 ( .A(\SUBBYTES[7].a/w2757 ), .B(n1715), .Z(\SUBBYTES[7].a/w2670 )
         );
  XNOR U4012 ( .A(\w1[7][28] ), .B(\w1[7][31] ), .Z(n1715) );
  ANDN U4013 ( .A(\SUBBYTES[7].a/w2758 ), .B(n1716), .Z(\SUBBYTES[7].a/w2668 )
         );
  XNOR U4014 ( .A(\w1[7][26] ), .B(\w1[7][31] ), .Z(n1716) );
  XOR U4015 ( .A(\w0[7][31] ), .B(g_input[927]), .Z(\w1[7][31] ) );
  IV U4016 ( .A(n1718), .Z(\w1[7][26] ) );
  ANDN U4017 ( .A(\SUBBYTES[7].a/w2760 ), .B(n1717), .Z(\SUBBYTES[7].a/w2667 )
         );
  XOR U4018 ( .A(n1718), .B(\w1[7][28] ), .Z(n1717) );
  XOR U4019 ( .A(\w0[7][28] ), .B(g_input[924]), .Z(\w1[7][28] ) );
  XNOR U4020 ( .A(\w0[7][26] ), .B(g_input[922]), .Z(n1718) );
  AND U4021 ( .A(\SUBBYTES[7].a/w164 ), .B(n1692), .Z(\SUBBYTES[7].a/w263 ) );
  XOR U4022 ( .A(\SUBBYTES[7].a/w232 ), .B(n1053), .Z(n1692) );
  AND U4023 ( .A(\SUBBYTES[7].a/w165 ), .B(n1699), .Z(\SUBBYTES[7].a/w261 ) );
  XOR U4024 ( .A(n13513), .B(\SUBBYTES[7].a/w232 ), .Z(n1699) );
  ANDN U4025 ( .A(n1700), .B(n1719), .Z(\SUBBYTES[7].a/w260 ) );
  XOR U4026 ( .A(n1053), .B(n13513), .Z(n1700) );
  AND U4027 ( .A(n1720), .B(\SUBBYTES[7].a/w2437 ), .Z(\SUBBYTES[7].a/w2572 )
         );
  AND U4028 ( .A(n1721), .B(\SUBBYTES[7].a/w2438 ), .Z(\SUBBYTES[7].a/w2570 )
         );
  AND U4029 ( .A(\SUBBYTES[7].a/w2568 ), .B(n1722), .Z(\SUBBYTES[7].a/w2569 )
         );
  ANDN U4030 ( .A(\w1[7][32] ), .B(n1723), .Z(\SUBBYTES[7].a/w2565 ) );
  AND U4031 ( .A(n1724), .B(\SUBBYTES[7].a/w2440 ), .Z(\SUBBYTES[7].a/w2563 )
         );
  AND U4032 ( .A(\SUBBYTES[7].a/w2561 ), .B(n1725), .Z(\SUBBYTES[7].a/w2562 )
         );
  XOR U4033 ( .A(\SUBBYTES[7].a/w2505 ), .B(n13534), .Z(n1725) );
  ANDN U4034 ( .A(\SUBBYTES[7].a/w166 ), .B(n1701), .Z(\SUBBYTES[7].a/w256 )
         );
  XNOR U4035 ( .A(\SUBBYTES[7].a/w225 ), .B(\SUBBYTES[7].a/w228 ), .Z(n1701)
         );
  AND U4036 ( .A(\SUBBYTES[7].a/w2548 ), .B(\SUBBYTES[7].a/w2550 ), .Z(
        \SUBBYTES[7].a/w2557 ) );
  AND U4037 ( .A(\SUBBYTES[7].a/w2549 ), .B(\SUBBYTES[7].a/w2551 ), .Z(
        \SUBBYTES[7].a/w2555 ) );
  AND U4038 ( .A(\SUBBYTES[7].a/w2552 ), .B(\SUBBYTES[7].a/w2553 ), .Z(
        \SUBBYTES[7].a/w2554 ) );
  AND U4039 ( .A(\SUBBYTES[7].a/w2441 ), .B(n1720), .Z(\SUBBYTES[7].a/w2540 )
         );
  XOR U4040 ( .A(\SUBBYTES[7].a/w2509 ), .B(n1064), .Z(n1720) );
  AND U4041 ( .A(\SUBBYTES[7].a/w167 ), .B(n1703), .Z(\SUBBYTES[7].a/w254 ) );
  XNOR U4042 ( .A(n1726), .B(\SUBBYTES[7].a/w225 ), .Z(n1703) );
  AND U4043 ( .A(\SUBBYTES[7].a/w2442 ), .B(n1721), .Z(\SUBBYTES[7].a/w2538 )
         );
  XOR U4044 ( .A(n13535), .B(\SUBBYTES[7].a/w2509 ), .Z(n1721) );
  ANDN U4045 ( .A(n1722), .B(n1727), .Z(\SUBBYTES[7].a/w2537 ) );
  XOR U4046 ( .A(n1064), .B(n13535), .Z(n1722) );
  ANDN U4047 ( .A(\SUBBYTES[7].a/w2443 ), .B(n1723), .Z(\SUBBYTES[7].a/w2533 )
         );
  XNOR U4048 ( .A(\SUBBYTES[7].a/w2502 ), .B(\SUBBYTES[7].a/w2505 ), .Z(n1723)
         );
  AND U4049 ( .A(\SUBBYTES[7].a/w2444 ), .B(n1724), .Z(\SUBBYTES[7].a/w2531 )
         );
  XNOR U4050 ( .A(n1728), .B(\SUBBYTES[7].a/w2502 ), .Z(n1724) );
  AND U4051 ( .A(\SUBBYTES[7].a/w2529 ), .B(n1729), .Z(\SUBBYTES[7].a/w2530 )
         );
  XOR U4052 ( .A(n1730), .B(n1728), .Z(n1729) );
  IV U4053 ( .A(n13534), .Z(n1728) );
  AND U4054 ( .A(\SUBBYTES[7].a/w252 ), .B(n1731), .Z(\SUBBYTES[7].a/w253 ) );
  XOR U4055 ( .A(n1732), .B(n1726), .Z(n1731) );
  IV U4056 ( .A(n13512), .Z(n1726) );
  ANDN U4057 ( .A(\SUBBYTES[7].a/w2548 ), .B(n1733), .Z(\SUBBYTES[7].a/w2525 )
         );
  ANDN U4058 ( .A(\SUBBYTES[7].a/w2549 ), .B(n1734), .Z(\SUBBYTES[7].a/w2523 )
         );
  ANDN U4059 ( .A(\SUBBYTES[7].a/w2552 ), .B(n1735), .Z(\SUBBYTES[7].a/w2522 )
         );
  AND U4060 ( .A(\SUBBYTES[7].a/w2508 ), .B(\SUBBYTES[7].a/w2507 ), .Z(
        \SUBBYTES[7].a/w2509 ) );
  IV U4061 ( .A(n1730), .Z(\SUBBYTES[7].a/w2505 ) );
  NAND U4062 ( .A(\SUBBYTES[7].a/w2484 ), .B(\SUBBYTES[7].a/w2499 ), .Z(n1730)
         );
  AND U4063 ( .A(\SUBBYTES[7].a/w2501 ), .B(\SUBBYTES[7].a/w2507 ), .Z(
        \SUBBYTES[7].a/w2502 ) );
  AND U4064 ( .A(\SUBBYTES[7].a/w2486 ), .B(\SUBBYTES[7].a/w2484 ), .Z(
        \SUBBYTES[7].a/w2496 ) );
  AND U4065 ( .A(\SUBBYTES[7].a/w2487 ), .B(\SUBBYTES[7].a/w2485 ), .Z(
        \SUBBYTES[7].a/w2494 ) );
  AND U4066 ( .A(\SUBBYTES[7].a/w2501 ), .B(\SUBBYTES[7].a/w2508 ), .Z(
        \SUBBYTES[7].a/w2493 ) );
  ANDN U4067 ( .A(\SUBBYTES[7].a/w271 ), .B(n1736), .Z(\SUBBYTES[7].a/w248 )
         );
  AND U4068 ( .A(\SUBBYTES[7].a/w2441 ), .B(\SUBBYTES[7].a/w2437 ), .Z(
        \SUBBYTES[7].a/w2478 ) );
  AND U4069 ( .A(\SUBBYTES[7].a/w2442 ), .B(\SUBBYTES[7].a/w2438 ), .Z(
        \SUBBYTES[7].a/w2476 ) );
  ANDN U4070 ( .A(\SUBBYTES[7].a/w2568 ), .B(n1727), .Z(\SUBBYTES[7].a/w2475 )
         );
  XNOR U4071 ( .A(\w1[7][33] ), .B(\w1[7][39] ), .Z(n1727) );
  XOR U4072 ( .A(\w0[7][33] ), .B(g_input[929]), .Z(\w1[7][33] ) );
  AND U4073 ( .A(\w1[7][32] ), .B(\SUBBYTES[7].a/w2443 ), .Z(
        \SUBBYTES[7].a/w2471 ) );
  XOR U4074 ( .A(\w0[7][32] ), .B(g_input[928]), .Z(\w1[7][32] ) );
  AND U4075 ( .A(\SUBBYTES[7].a/w2444 ), .B(\SUBBYTES[7].a/w2440 ), .Z(
        \SUBBYTES[7].a/w2469 ) );
  AND U4076 ( .A(\SUBBYTES[7].a/w2529 ), .B(\SUBBYTES[7].a/w2561 ), .Z(
        \SUBBYTES[7].a/w2468 ) );
  ANDN U4077 ( .A(\SUBBYTES[7].a/w2550 ), .B(n1733), .Z(\SUBBYTES[7].a/w2463 )
         );
  XNOR U4078 ( .A(\w1[7][36] ), .B(\w1[7][39] ), .Z(n1733) );
  ANDN U4079 ( .A(\SUBBYTES[7].a/w2551 ), .B(n1734), .Z(\SUBBYTES[7].a/w2461 )
         );
  XNOR U4080 ( .A(\w1[7][34] ), .B(\w1[7][39] ), .Z(n1734) );
  XOR U4081 ( .A(\w0[7][39] ), .B(g_input[935]), .Z(\w1[7][39] ) );
  IV U4082 ( .A(n1737), .Z(\w1[7][34] ) );
  ANDN U4083 ( .A(\SUBBYTES[7].a/w2553 ), .B(n1735), .Z(\SUBBYTES[7].a/w2460 )
         );
  XOR U4084 ( .A(n1737), .B(\w1[7][36] ), .Z(n1735) );
  XOR U4085 ( .A(\w0[7][36] ), .B(g_input[932]), .Z(\w1[7][36] ) );
  XNOR U4086 ( .A(\w0[7][34] ), .B(g_input[930]), .Z(n1737) );
  ANDN U4087 ( .A(\SUBBYTES[7].a/w272 ), .B(n1738), .Z(\SUBBYTES[7].a/w246 )
         );
  ANDN U4088 ( .A(\SUBBYTES[7].a/w275 ), .B(n1739), .Z(\SUBBYTES[7].a/w245 )
         );
  AND U4089 ( .A(n1740), .B(\SUBBYTES[7].a/w2230 ), .Z(\SUBBYTES[7].a/w2365 )
         );
  AND U4090 ( .A(n1741), .B(\SUBBYTES[7].a/w2231 ), .Z(\SUBBYTES[7].a/w2363 )
         );
  AND U4091 ( .A(\SUBBYTES[7].a/w2361 ), .B(n1742), .Z(\SUBBYTES[7].a/w2362 )
         );
  ANDN U4092 ( .A(\w1[7][40] ), .B(n1743), .Z(\SUBBYTES[7].a/w2358 ) );
  AND U4093 ( .A(n1744), .B(\SUBBYTES[7].a/w2233 ), .Z(\SUBBYTES[7].a/w2356 )
         );
  AND U4094 ( .A(\SUBBYTES[7].a/w2354 ), .B(n1745), .Z(\SUBBYTES[7].a/w2355 )
         );
  XOR U4095 ( .A(\SUBBYTES[7].a/w2298 ), .B(n13532), .Z(n1745) );
  AND U4096 ( .A(\SUBBYTES[7].a/w2341 ), .B(\SUBBYTES[7].a/w2343 ), .Z(
        \SUBBYTES[7].a/w2350 ) );
  AND U4097 ( .A(\SUBBYTES[7].a/w2342 ), .B(\SUBBYTES[7].a/w2344 ), .Z(
        \SUBBYTES[7].a/w2348 ) );
  AND U4098 ( .A(\SUBBYTES[7].a/w2345 ), .B(\SUBBYTES[7].a/w2346 ), .Z(
        \SUBBYTES[7].a/w2347 ) );
  AND U4099 ( .A(\SUBBYTES[7].a/w2234 ), .B(n1740), .Z(\SUBBYTES[7].a/w2333 )
         );
  XOR U4100 ( .A(\SUBBYTES[7].a/w2302 ), .B(n1063), .Z(n1740) );
  AND U4101 ( .A(\SUBBYTES[7].a/w2235 ), .B(n1741), .Z(\SUBBYTES[7].a/w2331 )
         );
  XOR U4102 ( .A(n13533), .B(\SUBBYTES[7].a/w2302 ), .Z(n1741) );
  ANDN U4103 ( .A(n1742), .B(n1746), .Z(\SUBBYTES[7].a/w2330 ) );
  XOR U4104 ( .A(n1063), .B(n13533), .Z(n1742) );
  ANDN U4105 ( .A(\SUBBYTES[7].a/w2236 ), .B(n1743), .Z(\SUBBYTES[7].a/w2326 )
         );
  XNOR U4106 ( .A(\SUBBYTES[7].a/w2295 ), .B(\SUBBYTES[7].a/w2298 ), .Z(n1743)
         );
  AND U4107 ( .A(\SUBBYTES[7].a/w2237 ), .B(n1744), .Z(\SUBBYTES[7].a/w2324 )
         );
  XNOR U4108 ( .A(n1747), .B(\SUBBYTES[7].a/w2295 ), .Z(n1744) );
  AND U4109 ( .A(\SUBBYTES[7].a/w2322 ), .B(n1748), .Z(\SUBBYTES[7].a/w2323 )
         );
  XOR U4110 ( .A(n1749), .B(n1747), .Z(n1748) );
  IV U4111 ( .A(n13532), .Z(n1747) );
  AND U4112 ( .A(\SUBBYTES[7].a/w231 ), .B(\SUBBYTES[7].a/w230 ), .Z(
        \SUBBYTES[7].a/w232 ) );
  ANDN U4113 ( .A(\SUBBYTES[7].a/w2341 ), .B(n1750), .Z(\SUBBYTES[7].a/w2318 )
         );
  ANDN U4114 ( .A(\SUBBYTES[7].a/w2342 ), .B(n1751), .Z(\SUBBYTES[7].a/w2316 )
         );
  ANDN U4115 ( .A(\SUBBYTES[7].a/w2345 ), .B(n1752), .Z(\SUBBYTES[7].a/w2315 )
         );
  AND U4116 ( .A(\SUBBYTES[7].a/w2301 ), .B(\SUBBYTES[7].a/w2300 ), .Z(
        \SUBBYTES[7].a/w2302 ) );
  IV U4117 ( .A(n1749), .Z(\SUBBYTES[7].a/w2298 ) );
  NAND U4118 ( .A(\SUBBYTES[7].a/w2277 ), .B(\SUBBYTES[7].a/w2292 ), .Z(n1749)
         );
  AND U4119 ( .A(\SUBBYTES[7].a/w2294 ), .B(\SUBBYTES[7].a/w2300 ), .Z(
        \SUBBYTES[7].a/w2295 ) );
  AND U4120 ( .A(\SUBBYTES[7].a/w2279 ), .B(\SUBBYTES[7].a/w2277 ), .Z(
        \SUBBYTES[7].a/w2289 ) );
  AND U4121 ( .A(\SUBBYTES[7].a/w2280 ), .B(\SUBBYTES[7].a/w2278 ), .Z(
        \SUBBYTES[7].a/w2287 ) );
  AND U4122 ( .A(\SUBBYTES[7].a/w2294 ), .B(\SUBBYTES[7].a/w2301 ), .Z(
        \SUBBYTES[7].a/w2286 ) );
  IV U4123 ( .A(n1732), .Z(\SUBBYTES[7].a/w228 ) );
  NAND U4124 ( .A(\SUBBYTES[7].a/w207 ), .B(\SUBBYTES[7].a/w222 ), .Z(n1732)
         );
  AND U4125 ( .A(\SUBBYTES[7].a/w2234 ), .B(\SUBBYTES[7].a/w2230 ), .Z(
        \SUBBYTES[7].a/w2271 ) );
  AND U4126 ( .A(\SUBBYTES[7].a/w2235 ), .B(\SUBBYTES[7].a/w2231 ), .Z(
        \SUBBYTES[7].a/w2269 ) );
  ANDN U4127 ( .A(\SUBBYTES[7].a/w2361 ), .B(n1746), .Z(\SUBBYTES[7].a/w2268 )
         );
  XNOR U4128 ( .A(\w1[7][41] ), .B(\w1[7][47] ), .Z(n1746) );
  XOR U4129 ( .A(\w0[7][41] ), .B(g_input[937]), .Z(\w1[7][41] ) );
  AND U4130 ( .A(\w1[7][40] ), .B(\SUBBYTES[7].a/w2236 ), .Z(
        \SUBBYTES[7].a/w2264 ) );
  XOR U4131 ( .A(\w0[7][40] ), .B(g_input[936]), .Z(\w1[7][40] ) );
  AND U4132 ( .A(\SUBBYTES[7].a/w2237 ), .B(\SUBBYTES[7].a/w2233 ), .Z(
        \SUBBYTES[7].a/w2262 ) );
  AND U4133 ( .A(\SUBBYTES[7].a/w2322 ), .B(\SUBBYTES[7].a/w2354 ), .Z(
        \SUBBYTES[7].a/w2261 ) );
  ANDN U4134 ( .A(\SUBBYTES[7].a/w2343 ), .B(n1750), .Z(\SUBBYTES[7].a/w2256 )
         );
  XNOR U4135 ( .A(\w1[7][44] ), .B(\w1[7][47] ), .Z(n1750) );
  ANDN U4136 ( .A(\SUBBYTES[7].a/w2344 ), .B(n1751), .Z(\SUBBYTES[7].a/w2254 )
         );
  XNOR U4137 ( .A(\w1[7][42] ), .B(\w1[7][47] ), .Z(n1751) );
  XOR U4138 ( .A(\w0[7][47] ), .B(g_input[943]), .Z(\w1[7][47] ) );
  IV U4139 ( .A(n1753), .Z(\w1[7][42] ) );
  ANDN U4140 ( .A(\SUBBYTES[7].a/w2346 ), .B(n1752), .Z(\SUBBYTES[7].a/w2253 )
         );
  XOR U4141 ( .A(n1753), .B(\w1[7][44] ), .Z(n1752) );
  XOR U4142 ( .A(\w0[7][44] ), .B(g_input[940]), .Z(\w1[7][44] ) );
  XNOR U4143 ( .A(\w0[7][42] ), .B(g_input[938]), .Z(n1753) );
  AND U4144 ( .A(\SUBBYTES[7].a/w224 ), .B(\SUBBYTES[7].a/w230 ), .Z(
        \SUBBYTES[7].a/w225 ) );
  AND U4145 ( .A(\SUBBYTES[7].a/w209 ), .B(\SUBBYTES[7].a/w207 ), .Z(
        \SUBBYTES[7].a/w219 ) );
  AND U4146 ( .A(\SUBBYTES[7].a/w210 ), .B(\SUBBYTES[7].a/w208 ), .Z(
        \SUBBYTES[7].a/w217 ) );
  AND U4147 ( .A(\SUBBYTES[7].a/w224 ), .B(\SUBBYTES[7].a/w231 ), .Z(
        \SUBBYTES[7].a/w216 ) );
  AND U4148 ( .A(n1754), .B(\SUBBYTES[7].a/w2023 ), .Z(\SUBBYTES[7].a/w2158 )
         );
  AND U4149 ( .A(n1755), .B(\SUBBYTES[7].a/w2024 ), .Z(\SUBBYTES[7].a/w2156 )
         );
  AND U4150 ( .A(\SUBBYTES[7].a/w2154 ), .B(n1756), .Z(\SUBBYTES[7].a/w2155 )
         );
  ANDN U4151 ( .A(\w1[7][48] ), .B(n1757), .Z(\SUBBYTES[7].a/w2151 ) );
  AND U4152 ( .A(n1758), .B(\SUBBYTES[7].a/w2026 ), .Z(\SUBBYTES[7].a/w2149 )
         );
  AND U4153 ( .A(\SUBBYTES[7].a/w2147 ), .B(n1759), .Z(\SUBBYTES[7].a/w2148 )
         );
  XOR U4154 ( .A(\SUBBYTES[7].a/w2091 ), .B(n13530), .Z(n1759) );
  AND U4155 ( .A(\SUBBYTES[7].a/w2134 ), .B(\SUBBYTES[7].a/w2136 ), .Z(
        \SUBBYTES[7].a/w2143 ) );
  AND U4156 ( .A(\SUBBYTES[7].a/w2135 ), .B(\SUBBYTES[7].a/w2137 ), .Z(
        \SUBBYTES[7].a/w2141 ) );
  AND U4157 ( .A(\SUBBYTES[7].a/w2138 ), .B(\SUBBYTES[7].a/w2139 ), .Z(
        \SUBBYTES[7].a/w2140 ) );
  AND U4158 ( .A(\SUBBYTES[7].a/w2027 ), .B(n1754), .Z(\SUBBYTES[7].a/w2126 )
         );
  XOR U4159 ( .A(\SUBBYTES[7].a/w2095 ), .B(n1062), .Z(n1754) );
  AND U4160 ( .A(\SUBBYTES[7].a/w2028 ), .B(n1755), .Z(\SUBBYTES[7].a/w2124 )
         );
  XOR U4161 ( .A(n13531), .B(\SUBBYTES[7].a/w2095 ), .Z(n1755) );
  ANDN U4162 ( .A(n1756), .B(n1760), .Z(\SUBBYTES[7].a/w2123 ) );
  XOR U4163 ( .A(n1062), .B(n13531), .Z(n1756) );
  ANDN U4164 ( .A(\SUBBYTES[7].a/w2029 ), .B(n1757), .Z(\SUBBYTES[7].a/w2119 )
         );
  XNOR U4165 ( .A(\SUBBYTES[7].a/w2088 ), .B(\SUBBYTES[7].a/w2091 ), .Z(n1757)
         );
  AND U4166 ( .A(\SUBBYTES[7].a/w2030 ), .B(n1758), .Z(\SUBBYTES[7].a/w2117 )
         );
  XNOR U4167 ( .A(n1761), .B(\SUBBYTES[7].a/w2088 ), .Z(n1758) );
  AND U4168 ( .A(\SUBBYTES[7].a/w2115 ), .B(n1762), .Z(\SUBBYTES[7].a/w2116 )
         );
  XOR U4169 ( .A(n1763), .B(n1761), .Z(n1762) );
  IV U4170 ( .A(n13530), .Z(n1761) );
  ANDN U4171 ( .A(\SUBBYTES[7].a/w2134 ), .B(n1764), .Z(\SUBBYTES[7].a/w2111 )
         );
  ANDN U4172 ( .A(\SUBBYTES[7].a/w2135 ), .B(n1765), .Z(\SUBBYTES[7].a/w2109 )
         );
  ANDN U4173 ( .A(\SUBBYTES[7].a/w2138 ), .B(n1766), .Z(\SUBBYTES[7].a/w2108 )
         );
  AND U4174 ( .A(\SUBBYTES[7].a/w2094 ), .B(\SUBBYTES[7].a/w2093 ), .Z(
        \SUBBYTES[7].a/w2095 ) );
  IV U4175 ( .A(n1763), .Z(\SUBBYTES[7].a/w2091 ) );
  NAND U4176 ( .A(\SUBBYTES[7].a/w2070 ), .B(\SUBBYTES[7].a/w2085 ), .Z(n1763)
         );
  AND U4177 ( .A(\SUBBYTES[7].a/w2087 ), .B(\SUBBYTES[7].a/w2093 ), .Z(
        \SUBBYTES[7].a/w2088 ) );
  AND U4178 ( .A(\SUBBYTES[7].a/w2072 ), .B(\SUBBYTES[7].a/w2070 ), .Z(
        \SUBBYTES[7].a/w2082 ) );
  AND U4179 ( .A(\SUBBYTES[7].a/w2073 ), .B(\SUBBYTES[7].a/w2071 ), .Z(
        \SUBBYTES[7].a/w2080 ) );
  AND U4180 ( .A(\SUBBYTES[7].a/w2087 ), .B(\SUBBYTES[7].a/w2094 ), .Z(
        \SUBBYTES[7].a/w2079 ) );
  AND U4181 ( .A(\SUBBYTES[7].a/w2027 ), .B(\SUBBYTES[7].a/w2023 ), .Z(
        \SUBBYTES[7].a/w2064 ) );
  AND U4182 ( .A(\SUBBYTES[7].a/w2028 ), .B(\SUBBYTES[7].a/w2024 ), .Z(
        \SUBBYTES[7].a/w2062 ) );
  ANDN U4183 ( .A(\SUBBYTES[7].a/w2154 ), .B(n1760), .Z(\SUBBYTES[7].a/w2061 )
         );
  XNOR U4184 ( .A(\w1[7][49] ), .B(\w1[7][55] ), .Z(n1760) );
  XOR U4185 ( .A(\w0[7][49] ), .B(g_input[945]), .Z(\w1[7][49] ) );
  AND U4186 ( .A(\w1[7][48] ), .B(\SUBBYTES[7].a/w2029 ), .Z(
        \SUBBYTES[7].a/w2057 ) );
  XOR U4187 ( .A(\w0[7][48] ), .B(g_input[944]), .Z(\w1[7][48] ) );
  AND U4188 ( .A(\SUBBYTES[7].a/w2030 ), .B(\SUBBYTES[7].a/w2026 ), .Z(
        \SUBBYTES[7].a/w2055 ) );
  AND U4189 ( .A(\SUBBYTES[7].a/w2115 ), .B(\SUBBYTES[7].a/w2147 ), .Z(
        \SUBBYTES[7].a/w2054 ) );
  ANDN U4190 ( .A(\SUBBYTES[7].a/w2136 ), .B(n1764), .Z(\SUBBYTES[7].a/w2049 )
         );
  XNOR U4191 ( .A(\w1[7][52] ), .B(\w1[7][55] ), .Z(n1764) );
  ANDN U4192 ( .A(\SUBBYTES[7].a/w2137 ), .B(n1765), .Z(\SUBBYTES[7].a/w2047 )
         );
  XNOR U4193 ( .A(\w1[7][50] ), .B(\w1[7][55] ), .Z(n1765) );
  XOR U4194 ( .A(\w0[7][55] ), .B(g_input[951]), .Z(\w1[7][55] ) );
  IV U4195 ( .A(n1767), .Z(\w1[7][50] ) );
  ANDN U4196 ( .A(\SUBBYTES[7].a/w2139 ), .B(n1766), .Z(\SUBBYTES[7].a/w2046 )
         );
  XOR U4197 ( .A(n1767), .B(\w1[7][52] ), .Z(n1766) );
  XOR U4198 ( .A(\w0[7][52] ), .B(g_input[948]), .Z(\w1[7][52] ) );
  XNOR U4199 ( .A(\w0[7][50] ), .B(g_input[946]), .Z(n1767) );
  AND U4200 ( .A(\SUBBYTES[7].a/w164 ), .B(\SUBBYTES[7].a/w160 ), .Z(
        \SUBBYTES[7].a/w201 ) );
  AND U4201 ( .A(\SUBBYTES[7].a/w165 ), .B(\SUBBYTES[7].a/w161 ), .Z(
        \SUBBYTES[7].a/w199 ) );
  ANDN U4202 ( .A(\SUBBYTES[7].a/w291 ), .B(n1719), .Z(\SUBBYTES[7].a/w198 )
         );
  XNOR U4203 ( .A(\w1[7][121] ), .B(\w1[7][127] ), .Z(n1719) );
  XOR U4204 ( .A(\w0[7][121] ), .B(g_input[1017]), .Z(\w1[7][121] ) );
  AND U4205 ( .A(n1768), .B(\SUBBYTES[7].a/w1816 ), .Z(\SUBBYTES[7].a/w1951 )
         );
  AND U4206 ( .A(n1769), .B(\SUBBYTES[7].a/w1817 ), .Z(\SUBBYTES[7].a/w1949 )
         );
  AND U4207 ( .A(\SUBBYTES[7].a/w1947 ), .B(n1770), .Z(\SUBBYTES[7].a/w1948 )
         );
  ANDN U4208 ( .A(\w1[7][56] ), .B(n1771), .Z(\SUBBYTES[7].a/w1944 ) );
  AND U4209 ( .A(n1772), .B(\SUBBYTES[7].a/w1819 ), .Z(\SUBBYTES[7].a/w1942 )
         );
  AND U4210 ( .A(\SUBBYTES[7].a/w1940 ), .B(n1773), .Z(\SUBBYTES[7].a/w1941 )
         );
  XOR U4211 ( .A(\SUBBYTES[7].a/w1884 ), .B(n13528), .Z(n1773) );
  AND U4212 ( .A(\w1[7][120] ), .B(\SUBBYTES[7].a/w166 ), .Z(
        \SUBBYTES[7].a/w194 ) );
  XOR U4213 ( .A(\w0[7][120] ), .B(g_input[1016]), .Z(\w1[7][120] ) );
  AND U4214 ( .A(\SUBBYTES[7].a/w1927 ), .B(\SUBBYTES[7].a/w1929 ), .Z(
        \SUBBYTES[7].a/w1936 ) );
  AND U4215 ( .A(\SUBBYTES[7].a/w1928 ), .B(\SUBBYTES[7].a/w1930 ), .Z(
        \SUBBYTES[7].a/w1934 ) );
  AND U4216 ( .A(\SUBBYTES[7].a/w1931 ), .B(\SUBBYTES[7].a/w1932 ), .Z(
        \SUBBYTES[7].a/w1933 ) );
  AND U4217 ( .A(\SUBBYTES[7].a/w167 ), .B(\SUBBYTES[7].a/w163 ), .Z(
        \SUBBYTES[7].a/w192 ) );
  AND U4218 ( .A(\SUBBYTES[7].a/w1820 ), .B(n1768), .Z(\SUBBYTES[7].a/w1919 )
         );
  XOR U4219 ( .A(\SUBBYTES[7].a/w1888 ), .B(n1061), .Z(n1768) );
  AND U4220 ( .A(\SUBBYTES[7].a/w1821 ), .B(n1769), .Z(\SUBBYTES[7].a/w1917 )
         );
  XOR U4221 ( .A(n13529), .B(\SUBBYTES[7].a/w1888 ), .Z(n1769) );
  ANDN U4222 ( .A(n1770), .B(n1774), .Z(\SUBBYTES[7].a/w1916 ) );
  XOR U4223 ( .A(n1061), .B(n13529), .Z(n1770) );
  ANDN U4224 ( .A(\SUBBYTES[7].a/w1822 ), .B(n1771), .Z(\SUBBYTES[7].a/w1912 )
         );
  XNOR U4225 ( .A(\SUBBYTES[7].a/w1881 ), .B(\SUBBYTES[7].a/w1884 ), .Z(n1771)
         );
  AND U4226 ( .A(\SUBBYTES[7].a/w1823 ), .B(n1772), .Z(\SUBBYTES[7].a/w1910 )
         );
  XNOR U4227 ( .A(n1775), .B(\SUBBYTES[7].a/w1881 ), .Z(n1772) );
  AND U4228 ( .A(\SUBBYTES[7].a/w252 ), .B(\SUBBYTES[7].a/w284 ), .Z(
        \SUBBYTES[7].a/w191 ) );
  AND U4229 ( .A(\SUBBYTES[7].a/w1908 ), .B(n1776), .Z(\SUBBYTES[7].a/w1909 )
         );
  XOR U4230 ( .A(n1777), .B(n1775), .Z(n1776) );
  IV U4231 ( .A(n13528), .Z(n1775) );
  ANDN U4232 ( .A(\SUBBYTES[7].a/w1927 ), .B(n1778), .Z(\SUBBYTES[7].a/w1904 )
         );
  ANDN U4233 ( .A(\SUBBYTES[7].a/w1928 ), .B(n1779), .Z(\SUBBYTES[7].a/w1902 )
         );
  ANDN U4234 ( .A(\SUBBYTES[7].a/w1931 ), .B(n1780), .Z(\SUBBYTES[7].a/w1901 )
         );
  AND U4235 ( .A(\SUBBYTES[7].a/w1887 ), .B(\SUBBYTES[7].a/w1886 ), .Z(
        \SUBBYTES[7].a/w1888 ) );
  IV U4236 ( .A(n1777), .Z(\SUBBYTES[7].a/w1884 ) );
  NAND U4237 ( .A(\SUBBYTES[7].a/w1863 ), .B(\SUBBYTES[7].a/w1878 ), .Z(n1777)
         );
  AND U4238 ( .A(\SUBBYTES[7].a/w1880 ), .B(\SUBBYTES[7].a/w1886 ), .Z(
        \SUBBYTES[7].a/w1881 ) );
  AND U4239 ( .A(\SUBBYTES[7].a/w1865 ), .B(\SUBBYTES[7].a/w1863 ), .Z(
        \SUBBYTES[7].a/w1875 ) );
  AND U4240 ( .A(\SUBBYTES[7].a/w1866 ), .B(\SUBBYTES[7].a/w1864 ), .Z(
        \SUBBYTES[7].a/w1873 ) );
  AND U4241 ( .A(\SUBBYTES[7].a/w1880 ), .B(\SUBBYTES[7].a/w1887 ), .Z(
        \SUBBYTES[7].a/w1872 ) );
  ANDN U4242 ( .A(\SUBBYTES[7].a/w273 ), .B(n1736), .Z(\SUBBYTES[7].a/w186 )
         );
  XNOR U4243 ( .A(\w1[7][124] ), .B(\w1[7][127] ), .Z(n1736) );
  AND U4244 ( .A(\SUBBYTES[7].a/w1820 ), .B(\SUBBYTES[7].a/w1816 ), .Z(
        \SUBBYTES[7].a/w1857 ) );
  AND U4245 ( .A(\SUBBYTES[7].a/w1821 ), .B(\SUBBYTES[7].a/w1817 ), .Z(
        \SUBBYTES[7].a/w1855 ) );
  ANDN U4246 ( .A(\SUBBYTES[7].a/w1947 ), .B(n1774), .Z(\SUBBYTES[7].a/w1854 )
         );
  XNOR U4247 ( .A(\w1[7][57] ), .B(\w1[7][63] ), .Z(n1774) );
  XOR U4248 ( .A(\w0[7][57] ), .B(g_input[953]), .Z(\w1[7][57] ) );
  AND U4249 ( .A(\w1[7][56] ), .B(\SUBBYTES[7].a/w1822 ), .Z(
        \SUBBYTES[7].a/w1850 ) );
  XOR U4250 ( .A(\w0[7][56] ), .B(g_input[952]), .Z(\w1[7][56] ) );
  AND U4251 ( .A(\SUBBYTES[7].a/w1823 ), .B(\SUBBYTES[7].a/w1819 ), .Z(
        \SUBBYTES[7].a/w1848 ) );
  AND U4252 ( .A(\SUBBYTES[7].a/w1908 ), .B(\SUBBYTES[7].a/w1940 ), .Z(
        \SUBBYTES[7].a/w1847 ) );
  ANDN U4253 ( .A(\SUBBYTES[7].a/w1929 ), .B(n1778), .Z(\SUBBYTES[7].a/w1842 )
         );
  XNOR U4254 ( .A(\w1[7][60] ), .B(\w1[7][63] ), .Z(n1778) );
  ANDN U4255 ( .A(\SUBBYTES[7].a/w1930 ), .B(n1779), .Z(\SUBBYTES[7].a/w1840 )
         );
  XNOR U4256 ( .A(\w1[7][58] ), .B(\w1[7][63] ), .Z(n1779) );
  XOR U4257 ( .A(\w0[7][63] ), .B(g_input[959]), .Z(\w1[7][63] ) );
  IV U4258 ( .A(n1781), .Z(\w1[7][58] ) );
  ANDN U4259 ( .A(\SUBBYTES[7].a/w274 ), .B(n1738), .Z(\SUBBYTES[7].a/w184 )
         );
  XNOR U4260 ( .A(\w1[7][122] ), .B(\w1[7][127] ), .Z(n1738) );
  XOR U4261 ( .A(\w0[7][127] ), .B(g_input[1023]), .Z(\w1[7][127] ) );
  IV U4262 ( .A(n1782), .Z(\w1[7][122] ) );
  ANDN U4263 ( .A(\SUBBYTES[7].a/w1932 ), .B(n1780), .Z(\SUBBYTES[7].a/w1839 )
         );
  XOR U4264 ( .A(n1781), .B(\w1[7][60] ), .Z(n1780) );
  XOR U4265 ( .A(\w0[7][60] ), .B(g_input[956]), .Z(\w1[7][60] ) );
  XNOR U4266 ( .A(\w0[7][58] ), .B(g_input[954]), .Z(n1781) );
  ANDN U4267 ( .A(\SUBBYTES[7].a/w276 ), .B(n1739), .Z(\SUBBYTES[7].a/w183 )
         );
  XOR U4268 ( .A(n1782), .B(\w1[7][124] ), .Z(n1739) );
  XOR U4269 ( .A(\w0[7][124] ), .B(g_input[1020]), .Z(\w1[7][124] ) );
  XNOR U4270 ( .A(\w0[7][122] ), .B(g_input[1018]), .Z(n1782) );
  AND U4271 ( .A(n1783), .B(\SUBBYTES[7].a/w1609 ), .Z(\SUBBYTES[7].a/w1744 )
         );
  AND U4272 ( .A(n1784), .B(\SUBBYTES[7].a/w1610 ), .Z(\SUBBYTES[7].a/w1742 )
         );
  AND U4273 ( .A(\SUBBYTES[7].a/w1740 ), .B(n1785), .Z(\SUBBYTES[7].a/w1741 )
         );
  ANDN U4274 ( .A(\w1[7][64] ), .B(n1786), .Z(\SUBBYTES[7].a/w1737 ) );
  AND U4275 ( .A(n1787), .B(\SUBBYTES[7].a/w1612 ), .Z(\SUBBYTES[7].a/w1735 )
         );
  AND U4276 ( .A(\SUBBYTES[7].a/w1733 ), .B(n1788), .Z(\SUBBYTES[7].a/w1734 )
         );
  XOR U4277 ( .A(\SUBBYTES[7].a/w1677 ), .B(n13526), .Z(n1788) );
  AND U4278 ( .A(\SUBBYTES[7].a/w1720 ), .B(\SUBBYTES[7].a/w1722 ), .Z(
        \SUBBYTES[7].a/w1729 ) );
  AND U4279 ( .A(\SUBBYTES[7].a/w1721 ), .B(\SUBBYTES[7].a/w1723 ), .Z(
        \SUBBYTES[7].a/w1727 ) );
  AND U4280 ( .A(\SUBBYTES[7].a/w1724 ), .B(\SUBBYTES[7].a/w1725 ), .Z(
        \SUBBYTES[7].a/w1726 ) );
  AND U4281 ( .A(\SUBBYTES[7].a/w1613 ), .B(n1783), .Z(\SUBBYTES[7].a/w1712 )
         );
  XOR U4282 ( .A(\SUBBYTES[7].a/w1681 ), .B(n1060), .Z(n1783) );
  AND U4283 ( .A(\SUBBYTES[7].a/w1614 ), .B(n1784), .Z(\SUBBYTES[7].a/w1710 )
         );
  XOR U4284 ( .A(n13527), .B(\SUBBYTES[7].a/w1681 ), .Z(n1784) );
  ANDN U4285 ( .A(n1785), .B(n1789), .Z(\SUBBYTES[7].a/w1709 ) );
  XOR U4286 ( .A(n1060), .B(n13527), .Z(n1785) );
  ANDN U4287 ( .A(\SUBBYTES[7].a/w1615 ), .B(n1786), .Z(\SUBBYTES[7].a/w1705 )
         );
  XNOR U4288 ( .A(\SUBBYTES[7].a/w1674 ), .B(\SUBBYTES[7].a/w1677 ), .Z(n1786)
         );
  AND U4289 ( .A(\SUBBYTES[7].a/w1616 ), .B(n1787), .Z(\SUBBYTES[7].a/w1703 )
         );
  XNOR U4290 ( .A(n1790), .B(\SUBBYTES[7].a/w1674 ), .Z(n1787) );
  AND U4291 ( .A(\SUBBYTES[7].a/w1701 ), .B(n1791), .Z(\SUBBYTES[7].a/w1702 )
         );
  XOR U4292 ( .A(n1792), .B(n1790), .Z(n1791) );
  IV U4293 ( .A(n13526), .Z(n1790) );
  ANDN U4294 ( .A(\SUBBYTES[7].a/w1720 ), .B(n1793), .Z(\SUBBYTES[7].a/w1697 )
         );
  ANDN U4295 ( .A(\SUBBYTES[7].a/w1721 ), .B(n1794), .Z(\SUBBYTES[7].a/w1695 )
         );
  ANDN U4296 ( .A(\SUBBYTES[7].a/w1724 ), .B(n1795), .Z(\SUBBYTES[7].a/w1694 )
         );
  AND U4297 ( .A(\SUBBYTES[7].a/w1680 ), .B(\SUBBYTES[7].a/w1679 ), .Z(
        \SUBBYTES[7].a/w1681 ) );
  IV U4298 ( .A(n1792), .Z(\SUBBYTES[7].a/w1677 ) );
  NAND U4299 ( .A(\SUBBYTES[7].a/w1656 ), .B(\SUBBYTES[7].a/w1671 ), .Z(n1792)
         );
  AND U4300 ( .A(\SUBBYTES[7].a/w1673 ), .B(\SUBBYTES[7].a/w1679 ), .Z(
        \SUBBYTES[7].a/w1674 ) );
  AND U4301 ( .A(\SUBBYTES[7].a/w1658 ), .B(\SUBBYTES[7].a/w1656 ), .Z(
        \SUBBYTES[7].a/w1668 ) );
  AND U4302 ( .A(\SUBBYTES[7].a/w1659 ), .B(\SUBBYTES[7].a/w1657 ), .Z(
        \SUBBYTES[7].a/w1666 ) );
  AND U4303 ( .A(\SUBBYTES[7].a/w1673 ), .B(\SUBBYTES[7].a/w1680 ), .Z(
        \SUBBYTES[7].a/w1665 ) );
  AND U4304 ( .A(\SUBBYTES[7].a/w1613 ), .B(\SUBBYTES[7].a/w1609 ), .Z(
        \SUBBYTES[7].a/w1650 ) );
  AND U4305 ( .A(\SUBBYTES[7].a/w1614 ), .B(\SUBBYTES[7].a/w1610 ), .Z(
        \SUBBYTES[7].a/w1648 ) );
  ANDN U4306 ( .A(\SUBBYTES[7].a/w1740 ), .B(n1789), .Z(\SUBBYTES[7].a/w1647 )
         );
  XNOR U4307 ( .A(\w1[7][65] ), .B(\w1[7][71] ), .Z(n1789) );
  XOR U4308 ( .A(\w0[7][65] ), .B(g_input[961]), .Z(\w1[7][65] ) );
  AND U4309 ( .A(\w1[7][64] ), .B(\SUBBYTES[7].a/w1615 ), .Z(
        \SUBBYTES[7].a/w1643 ) );
  XOR U4310 ( .A(\w0[7][64] ), .B(g_input[960]), .Z(\w1[7][64] ) );
  AND U4311 ( .A(\SUBBYTES[7].a/w1616 ), .B(\SUBBYTES[7].a/w1612 ), .Z(
        \SUBBYTES[7].a/w1641 ) );
  AND U4312 ( .A(\SUBBYTES[7].a/w1701 ), .B(\SUBBYTES[7].a/w1733 ), .Z(
        \SUBBYTES[7].a/w1640 ) );
  ANDN U4313 ( .A(\SUBBYTES[7].a/w1722 ), .B(n1793), .Z(\SUBBYTES[7].a/w1635 )
         );
  XNOR U4314 ( .A(\w1[7][68] ), .B(\w1[7][71] ), .Z(n1793) );
  ANDN U4315 ( .A(\SUBBYTES[7].a/w1723 ), .B(n1794), .Z(\SUBBYTES[7].a/w1633 )
         );
  XNOR U4316 ( .A(\w1[7][66] ), .B(\w1[7][71] ), .Z(n1794) );
  XOR U4317 ( .A(\w0[7][71] ), .B(g_input[967]), .Z(\w1[7][71] ) );
  IV U4318 ( .A(n1796), .Z(\w1[7][66] ) );
  ANDN U4319 ( .A(\SUBBYTES[7].a/w1725 ), .B(n1795), .Z(\SUBBYTES[7].a/w1632 )
         );
  XOR U4320 ( .A(n1796), .B(\w1[7][68] ), .Z(n1795) );
  XOR U4321 ( .A(\w0[7][68] ), .B(g_input[964]), .Z(\w1[7][68] ) );
  XNOR U4322 ( .A(\w0[7][66] ), .B(g_input[962]), .Z(n1796) );
  AND U4323 ( .A(n1797), .B(\SUBBYTES[7].a/w1402 ), .Z(\SUBBYTES[7].a/w1537 )
         );
  AND U4324 ( .A(n1798), .B(\SUBBYTES[7].a/w1403 ), .Z(\SUBBYTES[7].a/w1535 )
         );
  AND U4325 ( .A(\SUBBYTES[7].a/w1533 ), .B(n1799), .Z(\SUBBYTES[7].a/w1534 )
         );
  ANDN U4326 ( .A(\w1[7][72] ), .B(n1800), .Z(\SUBBYTES[7].a/w1530 ) );
  AND U4327 ( .A(n1801), .B(\SUBBYTES[7].a/w1405 ), .Z(\SUBBYTES[7].a/w1528 )
         );
  AND U4328 ( .A(\SUBBYTES[7].a/w1526 ), .B(n1802), .Z(\SUBBYTES[7].a/w1527 )
         );
  XOR U4329 ( .A(\SUBBYTES[7].a/w1470 ), .B(n13524), .Z(n1802) );
  AND U4330 ( .A(\SUBBYTES[7].a/w1513 ), .B(\SUBBYTES[7].a/w1515 ), .Z(
        \SUBBYTES[7].a/w1522 ) );
  AND U4331 ( .A(\SUBBYTES[7].a/w1514 ), .B(\SUBBYTES[7].a/w1516 ), .Z(
        \SUBBYTES[7].a/w1520 ) );
  AND U4332 ( .A(\SUBBYTES[7].a/w1517 ), .B(\SUBBYTES[7].a/w1518 ), .Z(
        \SUBBYTES[7].a/w1519 ) );
  AND U4333 ( .A(\SUBBYTES[7].a/w1406 ), .B(n1797), .Z(\SUBBYTES[7].a/w1505 )
         );
  XOR U4334 ( .A(\SUBBYTES[7].a/w1474 ), .B(n1059), .Z(n1797) );
  AND U4335 ( .A(\SUBBYTES[7].a/w1407 ), .B(n1798), .Z(\SUBBYTES[7].a/w1503 )
         );
  XOR U4336 ( .A(n13525), .B(\SUBBYTES[7].a/w1474 ), .Z(n1798) );
  ANDN U4337 ( .A(n1799), .B(n1803), .Z(\SUBBYTES[7].a/w1502 ) );
  XOR U4338 ( .A(n1059), .B(n13525), .Z(n1799) );
  ANDN U4339 ( .A(\SUBBYTES[7].a/w1408 ), .B(n1800), .Z(\SUBBYTES[7].a/w1498 )
         );
  XNOR U4340 ( .A(\SUBBYTES[7].a/w1467 ), .B(\SUBBYTES[7].a/w1470 ), .Z(n1800)
         );
  AND U4341 ( .A(\SUBBYTES[7].a/w1409 ), .B(n1801), .Z(\SUBBYTES[7].a/w1496 )
         );
  XNOR U4342 ( .A(n1804), .B(\SUBBYTES[7].a/w1467 ), .Z(n1801) );
  AND U4343 ( .A(\SUBBYTES[7].a/w1494 ), .B(n1805), .Z(\SUBBYTES[7].a/w1495 )
         );
  XOR U4344 ( .A(n1806), .B(n1804), .Z(n1805) );
  IV U4345 ( .A(n13524), .Z(n1804) );
  ANDN U4346 ( .A(\SUBBYTES[7].a/w1513 ), .B(n1807), .Z(\SUBBYTES[7].a/w1490 )
         );
  ANDN U4347 ( .A(\SUBBYTES[7].a/w1514 ), .B(n1808), .Z(\SUBBYTES[7].a/w1488 )
         );
  ANDN U4348 ( .A(\SUBBYTES[7].a/w1517 ), .B(n1809), .Z(\SUBBYTES[7].a/w1487 )
         );
  AND U4349 ( .A(\SUBBYTES[7].a/w1473 ), .B(\SUBBYTES[7].a/w1472 ), .Z(
        \SUBBYTES[7].a/w1474 ) );
  IV U4350 ( .A(n1806), .Z(\SUBBYTES[7].a/w1470 ) );
  NAND U4351 ( .A(\SUBBYTES[7].a/w1449 ), .B(\SUBBYTES[7].a/w1464 ), .Z(n1806)
         );
  AND U4352 ( .A(\SUBBYTES[7].a/w1466 ), .B(\SUBBYTES[7].a/w1472 ), .Z(
        \SUBBYTES[7].a/w1467 ) );
  AND U4353 ( .A(\SUBBYTES[7].a/w1451 ), .B(\SUBBYTES[7].a/w1449 ), .Z(
        \SUBBYTES[7].a/w1461 ) );
  AND U4354 ( .A(\SUBBYTES[7].a/w1452 ), .B(\SUBBYTES[7].a/w1450 ), .Z(
        \SUBBYTES[7].a/w1459 ) );
  AND U4355 ( .A(\SUBBYTES[7].a/w1466 ), .B(\SUBBYTES[7].a/w1473 ), .Z(
        \SUBBYTES[7].a/w1458 ) );
  AND U4356 ( .A(\SUBBYTES[7].a/w1406 ), .B(\SUBBYTES[7].a/w1402 ), .Z(
        \SUBBYTES[7].a/w1443 ) );
  AND U4357 ( .A(\SUBBYTES[7].a/w1407 ), .B(\SUBBYTES[7].a/w1403 ), .Z(
        \SUBBYTES[7].a/w1441 ) );
  ANDN U4358 ( .A(\SUBBYTES[7].a/w1533 ), .B(n1803), .Z(\SUBBYTES[7].a/w1440 )
         );
  XNOR U4359 ( .A(\w1[7][73] ), .B(\w1[7][79] ), .Z(n1803) );
  XOR U4360 ( .A(\w0[7][73] ), .B(g_input[969]), .Z(\w1[7][73] ) );
  AND U4361 ( .A(\w1[7][72] ), .B(\SUBBYTES[7].a/w1408 ), .Z(
        \SUBBYTES[7].a/w1436 ) );
  XOR U4362 ( .A(\w0[7][72] ), .B(g_input[968]), .Z(\w1[7][72] ) );
  AND U4363 ( .A(\SUBBYTES[7].a/w1409 ), .B(\SUBBYTES[7].a/w1405 ), .Z(
        \SUBBYTES[7].a/w1434 ) );
  AND U4364 ( .A(\SUBBYTES[7].a/w1494 ), .B(\SUBBYTES[7].a/w1526 ), .Z(
        \SUBBYTES[7].a/w1433 ) );
  ANDN U4365 ( .A(\SUBBYTES[7].a/w1515 ), .B(n1807), .Z(\SUBBYTES[7].a/w1428 )
         );
  XNOR U4366 ( .A(\w1[7][76] ), .B(\w1[7][79] ), .Z(n1807) );
  ANDN U4367 ( .A(\SUBBYTES[7].a/w1516 ), .B(n1808), .Z(\SUBBYTES[7].a/w1426 )
         );
  XNOR U4368 ( .A(\w1[7][74] ), .B(\w1[7][79] ), .Z(n1808) );
  XOR U4369 ( .A(\w0[7][79] ), .B(g_input[975]), .Z(\w1[7][79] ) );
  IV U4370 ( .A(n1810), .Z(\w1[7][74] ) );
  ANDN U4371 ( .A(\SUBBYTES[7].a/w1518 ), .B(n1809), .Z(\SUBBYTES[7].a/w1425 )
         );
  XOR U4372 ( .A(n1810), .B(\w1[7][76] ), .Z(n1809) );
  XOR U4373 ( .A(\w0[7][76] ), .B(g_input[972]), .Z(\w1[7][76] ) );
  XNOR U4374 ( .A(\w0[7][74] ), .B(g_input[970]), .Z(n1810) );
  AND U4375 ( .A(n1811), .B(\SUBBYTES[7].a/w1195 ), .Z(\SUBBYTES[7].a/w1330 )
         );
  AND U4376 ( .A(n1812), .B(\SUBBYTES[7].a/w1196 ), .Z(\SUBBYTES[7].a/w1328 )
         );
  AND U4377 ( .A(\SUBBYTES[7].a/w1326 ), .B(n1813), .Z(\SUBBYTES[7].a/w1327 )
         );
  ANDN U4378 ( .A(\w1[7][80] ), .B(n1814), .Z(\SUBBYTES[7].a/w1323 ) );
  AND U4379 ( .A(n1815), .B(\SUBBYTES[7].a/w1198 ), .Z(\SUBBYTES[7].a/w1321 )
         );
  AND U4380 ( .A(\SUBBYTES[7].a/w1319 ), .B(n1816), .Z(\SUBBYTES[7].a/w1320 )
         );
  XOR U4381 ( .A(\SUBBYTES[7].a/w1263 ), .B(n13522), .Z(n1816) );
  AND U4382 ( .A(\SUBBYTES[7].a/w1306 ), .B(\SUBBYTES[7].a/w1308 ), .Z(
        \SUBBYTES[7].a/w1315 ) );
  AND U4383 ( .A(\SUBBYTES[7].a/w1307 ), .B(\SUBBYTES[7].a/w1309 ), .Z(
        \SUBBYTES[7].a/w1313 ) );
  AND U4384 ( .A(\SUBBYTES[7].a/w1310 ), .B(\SUBBYTES[7].a/w1311 ), .Z(
        \SUBBYTES[7].a/w1312 ) );
  AND U4385 ( .A(\SUBBYTES[7].a/w1199 ), .B(n1811), .Z(\SUBBYTES[7].a/w1298 )
         );
  XOR U4386 ( .A(\SUBBYTES[7].a/w1267 ), .B(n1058), .Z(n1811) );
  AND U4387 ( .A(\SUBBYTES[7].a/w1200 ), .B(n1812), .Z(\SUBBYTES[7].a/w1296 )
         );
  XOR U4388 ( .A(n13523), .B(\SUBBYTES[7].a/w1267 ), .Z(n1812) );
  ANDN U4389 ( .A(n1813), .B(n1817), .Z(\SUBBYTES[7].a/w1295 ) );
  XOR U4390 ( .A(n1058), .B(n13523), .Z(n1813) );
  ANDN U4391 ( .A(\SUBBYTES[7].a/w1201 ), .B(n1814), .Z(\SUBBYTES[7].a/w1291 )
         );
  XNOR U4392 ( .A(\SUBBYTES[7].a/w1260 ), .B(\SUBBYTES[7].a/w1263 ), .Z(n1814)
         );
  AND U4393 ( .A(\SUBBYTES[7].a/w1202 ), .B(n1815), .Z(\SUBBYTES[7].a/w1289 )
         );
  XNOR U4394 ( .A(n1818), .B(\SUBBYTES[7].a/w1260 ), .Z(n1815) );
  AND U4395 ( .A(\SUBBYTES[7].a/w1287 ), .B(n1819), .Z(\SUBBYTES[7].a/w1288 )
         );
  XOR U4396 ( .A(n1820), .B(n1818), .Z(n1819) );
  IV U4397 ( .A(n13522), .Z(n1818) );
  ANDN U4398 ( .A(\SUBBYTES[7].a/w1306 ), .B(n1821), .Z(\SUBBYTES[7].a/w1283 )
         );
  ANDN U4399 ( .A(\SUBBYTES[7].a/w1307 ), .B(n1822), .Z(\SUBBYTES[7].a/w1281 )
         );
  ANDN U4400 ( .A(\SUBBYTES[7].a/w1310 ), .B(n1823), .Z(\SUBBYTES[7].a/w1280 )
         );
  AND U4401 ( .A(\SUBBYTES[7].a/w1266 ), .B(\SUBBYTES[7].a/w1265 ), .Z(
        \SUBBYTES[7].a/w1267 ) );
  IV U4402 ( .A(n1820), .Z(\SUBBYTES[7].a/w1263 ) );
  NAND U4403 ( .A(\SUBBYTES[7].a/w1242 ), .B(\SUBBYTES[7].a/w1257 ), .Z(n1820)
         );
  AND U4404 ( .A(\SUBBYTES[7].a/w1259 ), .B(\SUBBYTES[7].a/w1265 ), .Z(
        \SUBBYTES[7].a/w1260 ) );
  AND U4405 ( .A(\SUBBYTES[7].a/w1244 ), .B(\SUBBYTES[7].a/w1242 ), .Z(
        \SUBBYTES[7].a/w1254 ) );
  AND U4406 ( .A(\SUBBYTES[7].a/w1245 ), .B(\SUBBYTES[7].a/w1243 ), .Z(
        \SUBBYTES[7].a/w1252 ) );
  AND U4407 ( .A(\SUBBYTES[7].a/w1259 ), .B(\SUBBYTES[7].a/w1266 ), .Z(
        \SUBBYTES[7].a/w1251 ) );
  AND U4408 ( .A(\SUBBYTES[7].a/w1199 ), .B(\SUBBYTES[7].a/w1195 ), .Z(
        \SUBBYTES[7].a/w1236 ) );
  AND U4409 ( .A(\SUBBYTES[7].a/w1200 ), .B(\SUBBYTES[7].a/w1196 ), .Z(
        \SUBBYTES[7].a/w1234 ) );
  ANDN U4410 ( .A(\SUBBYTES[7].a/w1326 ), .B(n1817), .Z(\SUBBYTES[7].a/w1233 )
         );
  XNOR U4411 ( .A(\w1[7][81] ), .B(\w1[7][87] ), .Z(n1817) );
  XOR U4412 ( .A(\w0[7][81] ), .B(g_input[977]), .Z(\w1[7][81] ) );
  AND U4413 ( .A(\w1[7][80] ), .B(\SUBBYTES[7].a/w1201 ), .Z(
        \SUBBYTES[7].a/w1229 ) );
  XOR U4414 ( .A(\w0[7][80] ), .B(g_input[976]), .Z(\w1[7][80] ) );
  AND U4415 ( .A(\SUBBYTES[7].a/w1202 ), .B(\SUBBYTES[7].a/w1198 ), .Z(
        \SUBBYTES[7].a/w1227 ) );
  AND U4416 ( .A(\SUBBYTES[7].a/w1287 ), .B(\SUBBYTES[7].a/w1319 ), .Z(
        \SUBBYTES[7].a/w1226 ) );
  ANDN U4417 ( .A(\SUBBYTES[7].a/w1308 ), .B(n1821), .Z(\SUBBYTES[7].a/w1221 )
         );
  XNOR U4418 ( .A(\w1[7][84] ), .B(\w1[7][87] ), .Z(n1821) );
  ANDN U4419 ( .A(\SUBBYTES[7].a/w1309 ), .B(n1822), .Z(\SUBBYTES[7].a/w1219 )
         );
  XNOR U4420 ( .A(\w1[7][82] ), .B(\w1[7][87] ), .Z(n1822) );
  XOR U4421 ( .A(\w0[7][87] ), .B(g_input[983]), .Z(\w1[7][87] ) );
  IV U4422 ( .A(n1824), .Z(\w1[7][82] ) );
  ANDN U4423 ( .A(\SUBBYTES[7].a/w1311 ), .B(n1823), .Z(\SUBBYTES[7].a/w1218 )
         );
  XOR U4424 ( .A(n1824), .B(\w1[7][84] ), .Z(n1823) );
  XOR U4425 ( .A(\w0[7][84] ), .B(g_input[980]), .Z(\w1[7][84] ) );
  XNOR U4426 ( .A(\w0[7][82] ), .B(g_input[978]), .Z(n1824) );
  AND U4427 ( .A(n1825), .B(\SUBBYTES[7].a/w988 ), .Z(\SUBBYTES[7].a/w1123 )
         );
  AND U4428 ( .A(n1826), .B(\SUBBYTES[7].a/w989 ), .Z(\SUBBYTES[7].a/w1121 )
         );
  AND U4429 ( .A(\SUBBYTES[7].a/w1119 ), .B(n1827), .Z(\SUBBYTES[7].a/w1120 )
         );
  ANDN U4430 ( .A(\w1[7][88] ), .B(n1828), .Z(\SUBBYTES[7].a/w1116 ) );
  AND U4431 ( .A(n1829), .B(\SUBBYTES[7].a/w991 ), .Z(\SUBBYTES[7].a/w1114 )
         );
  AND U4432 ( .A(\SUBBYTES[7].a/w1112 ), .B(n1830), .Z(\SUBBYTES[7].a/w1113 )
         );
  XOR U4433 ( .A(\SUBBYTES[7].a/w1056 ), .B(n13520), .Z(n1830) );
  AND U4434 ( .A(\SUBBYTES[7].a/w1099 ), .B(\SUBBYTES[7].a/w1101 ), .Z(
        \SUBBYTES[7].a/w1108 ) );
  AND U4435 ( .A(\SUBBYTES[7].a/w1100 ), .B(\SUBBYTES[7].a/w1102 ), .Z(
        \SUBBYTES[7].a/w1106 ) );
  AND U4436 ( .A(\SUBBYTES[7].a/w1103 ), .B(\SUBBYTES[7].a/w1104 ), .Z(
        \SUBBYTES[7].a/w1105 ) );
  AND U4437 ( .A(\SUBBYTES[7].a/w992 ), .B(n1825), .Z(\SUBBYTES[7].a/w1091 )
         );
  XOR U4438 ( .A(\SUBBYTES[7].a/w1060 ), .B(n1057), .Z(n1825) );
  AND U4439 ( .A(\SUBBYTES[7].a/w993 ), .B(n1826), .Z(\SUBBYTES[7].a/w1089 )
         );
  XOR U4440 ( .A(n13521), .B(\SUBBYTES[7].a/w1060 ), .Z(n1826) );
  ANDN U4441 ( .A(n1827), .B(n1831), .Z(\SUBBYTES[7].a/w1088 ) );
  XOR U4442 ( .A(n1057), .B(n13521), .Z(n1827) );
  ANDN U4443 ( .A(\SUBBYTES[7].a/w994 ), .B(n1828), .Z(\SUBBYTES[7].a/w1084 )
         );
  XNOR U4444 ( .A(\SUBBYTES[7].a/w1053 ), .B(\SUBBYTES[7].a/w1056 ), .Z(n1828)
         );
  AND U4445 ( .A(\SUBBYTES[7].a/w995 ), .B(n1829), .Z(\SUBBYTES[7].a/w1082 )
         );
  XNOR U4446 ( .A(n1832), .B(\SUBBYTES[7].a/w1053 ), .Z(n1829) );
  AND U4447 ( .A(\SUBBYTES[7].a/w1080 ), .B(n1833), .Z(\SUBBYTES[7].a/w1081 )
         );
  XOR U4448 ( .A(n1834), .B(n1832), .Z(n1833) );
  IV U4449 ( .A(n13520), .Z(n1832) );
  ANDN U4450 ( .A(\SUBBYTES[7].a/w1099 ), .B(n1835), .Z(\SUBBYTES[7].a/w1076 )
         );
  ANDN U4451 ( .A(\SUBBYTES[7].a/w1100 ), .B(n1836), .Z(\SUBBYTES[7].a/w1074 )
         );
  ANDN U4452 ( .A(\SUBBYTES[7].a/w1103 ), .B(n1837), .Z(\SUBBYTES[7].a/w1073 )
         );
  AND U4453 ( .A(\SUBBYTES[7].a/w1059 ), .B(\SUBBYTES[7].a/w1058 ), .Z(
        \SUBBYTES[7].a/w1060 ) );
  IV U4454 ( .A(n1834), .Z(\SUBBYTES[7].a/w1056 ) );
  NAND U4455 ( .A(\SUBBYTES[7].a/w1035 ), .B(\SUBBYTES[7].a/w1050 ), .Z(n1834)
         );
  AND U4456 ( .A(\SUBBYTES[7].a/w1052 ), .B(\SUBBYTES[7].a/w1058 ), .Z(
        \SUBBYTES[7].a/w1053 ) );
  AND U4457 ( .A(\SUBBYTES[7].a/w1037 ), .B(\SUBBYTES[7].a/w1035 ), .Z(
        \SUBBYTES[7].a/w1047 ) );
  AND U4458 ( .A(\SUBBYTES[7].a/w1038 ), .B(\SUBBYTES[7].a/w1036 ), .Z(
        \SUBBYTES[7].a/w1045 ) );
  AND U4459 ( .A(\SUBBYTES[7].a/w1052 ), .B(\SUBBYTES[7].a/w1059 ), .Z(
        \SUBBYTES[7].a/w1044 ) );
  AND U4460 ( .A(\SUBBYTES[7].a/w992 ), .B(\SUBBYTES[7].a/w988 ), .Z(
        \SUBBYTES[7].a/w1029 ) );
  AND U4461 ( .A(\SUBBYTES[7].a/w993 ), .B(\SUBBYTES[7].a/w989 ), .Z(
        \SUBBYTES[7].a/w1027 ) );
  ANDN U4462 ( .A(\SUBBYTES[7].a/w1119 ), .B(n1831), .Z(\SUBBYTES[7].a/w1026 )
         );
  XNOR U4463 ( .A(\w1[7][89] ), .B(\w1[7][95] ), .Z(n1831) );
  XOR U4464 ( .A(\w0[7][89] ), .B(g_input[985]), .Z(\w1[7][89] ) );
  AND U4465 ( .A(\w1[7][88] ), .B(\SUBBYTES[7].a/w994 ), .Z(
        \SUBBYTES[7].a/w1022 ) );
  XOR U4466 ( .A(\w0[7][88] ), .B(g_input[984]), .Z(\w1[7][88] ) );
  AND U4467 ( .A(\SUBBYTES[7].a/w995 ), .B(\SUBBYTES[7].a/w991 ), .Z(
        \SUBBYTES[7].a/w1020 ) );
  AND U4468 ( .A(\SUBBYTES[7].a/w1080 ), .B(\SUBBYTES[7].a/w1112 ), .Z(
        \SUBBYTES[7].a/w1019 ) );
  ANDN U4469 ( .A(\SUBBYTES[7].a/w1101 ), .B(n1835), .Z(\SUBBYTES[7].a/w1014 )
         );
  XNOR U4470 ( .A(\w1[7][92] ), .B(\w1[7][95] ), .Z(n1835) );
  ANDN U4471 ( .A(\SUBBYTES[7].a/w1102 ), .B(n1836), .Z(\SUBBYTES[7].a/w1012 )
         );
  XNOR U4472 ( .A(\w1[7][90] ), .B(\w1[7][95] ), .Z(n1836) );
  XOR U4473 ( .A(\w0[7][95] ), .B(g_input[991]), .Z(\w1[7][95] ) );
  IV U4474 ( .A(n1838), .Z(\w1[7][90] ) );
  ANDN U4475 ( .A(\SUBBYTES[7].a/w1104 ), .B(n1837), .Z(\SUBBYTES[7].a/w1011 )
         );
  XOR U4476 ( .A(n1838), .B(\w1[7][92] ), .Z(n1837) );
  XOR U4477 ( .A(\w0[7][92] ), .B(g_input[988]), .Z(\w1[7][92] ) );
  XNOR U4478 ( .A(\w0[7][90] ), .B(g_input[986]), .Z(n1838) );
  AND U4479 ( .A(\SUBBYTES[7].a/w2084 ), .B(\SUBBYTES[7].a/w2071 ), .Z(n13530)
         );
  AND U4480 ( .A(\SUBBYTES[7].a/w1877 ), .B(\SUBBYTES[7].a/w1866 ), .Z(n13529)
         );
  AND U4481 ( .A(\SUBBYTES[7].a/w221 ), .B(\SUBBYTES[7].a/w208 ), .Z(n13512)
         );
  AND U4482 ( .A(\SUBBYTES[7].a/w1877 ), .B(\SUBBYTES[7].a/w1864 ), .Z(n13528)
         );
  AND U4483 ( .A(\SUBBYTES[7].a/w1670 ), .B(\SUBBYTES[7].a/w1659 ), .Z(n13527)
         );
  AND U4484 ( .A(\SUBBYTES[7].a/w1670 ), .B(\SUBBYTES[7].a/w1657 ), .Z(n13526)
         );
  AND U4485 ( .A(\SUBBYTES[7].a/w1463 ), .B(\SUBBYTES[7].a/w1452 ), .Z(n13525)
         );
  AND U4486 ( .A(\SUBBYTES[7].a/w1463 ), .B(\SUBBYTES[7].a/w1450 ), .Z(n13524)
         );
  AND U4487 ( .A(\SUBBYTES[7].a/w1256 ), .B(\SUBBYTES[7].a/w1245 ), .Z(n13523)
         );
  AND U4488 ( .A(\SUBBYTES[7].a/w1256 ), .B(\SUBBYTES[7].a/w1243 ), .Z(n13522)
         );
  AND U4489 ( .A(\SUBBYTES[7].a/w1049 ), .B(\SUBBYTES[7].a/w1038 ), .Z(n13521)
         );
  AND U4490 ( .A(\SUBBYTES[7].a/w1049 ), .B(\SUBBYTES[7].a/w1036 ), .Z(n13520)
         );
  AND U4491 ( .A(\SUBBYTES[7].a/w842 ), .B(\SUBBYTES[7].a/w831 ), .Z(n13519)
         );
  AND U4492 ( .A(\SUBBYTES[7].a/w842 ), .B(\SUBBYTES[7].a/w829 ), .Z(n13518)
         );
  AND U4493 ( .A(\SUBBYTES[7].a/w635 ), .B(\SUBBYTES[7].a/w624 ), .Z(n13517)
         );
  AND U4494 ( .A(\SUBBYTES[7].a/w635 ), .B(\SUBBYTES[7].a/w622 ), .Z(n13516)
         );
  AND U4495 ( .A(\SUBBYTES[7].a/w428 ), .B(\SUBBYTES[7].a/w417 ), .Z(n13515)
         );
  AND U4496 ( .A(\SUBBYTES[7].a/w428 ), .B(\SUBBYTES[7].a/w415 ), .Z(n13514)
         );
  AND U4497 ( .A(\SUBBYTES[7].a/w3326 ), .B(\SUBBYTES[7].a/w3315 ), .Z(n13543)
         );
  AND U4498 ( .A(\SUBBYTES[7].a/w3326 ), .B(\SUBBYTES[7].a/w3313 ), .Z(n13542)
         );
  AND U4499 ( .A(\SUBBYTES[7].a/w3119 ), .B(\SUBBYTES[7].a/w3108 ), .Z(n13541)
         );
  AND U4500 ( .A(\SUBBYTES[7].a/w3119 ), .B(\SUBBYTES[7].a/w3106 ), .Z(n13540)
         );
  AND U4501 ( .A(\SUBBYTES[7].a/w2912 ), .B(\SUBBYTES[7].a/w2901 ), .Z(n13539)
         );
  AND U4502 ( .A(\SUBBYTES[7].a/w2912 ), .B(\SUBBYTES[7].a/w2899 ), .Z(n13538)
         );
  AND U4503 ( .A(\SUBBYTES[7].a/w2705 ), .B(\SUBBYTES[7].a/w2694 ), .Z(n13537)
         );
  AND U4504 ( .A(\SUBBYTES[7].a/w2705 ), .B(\SUBBYTES[7].a/w2692 ), .Z(n13536)
         );
  AND U4505 ( .A(\SUBBYTES[7].a/w2498 ), .B(\SUBBYTES[7].a/w2487 ), .Z(n13535)
         );
  AND U4506 ( .A(\SUBBYTES[7].a/w2498 ), .B(\SUBBYTES[7].a/w2485 ), .Z(n13534)
         );
  AND U4507 ( .A(\SUBBYTES[7].a/w2291 ), .B(\SUBBYTES[7].a/w2280 ), .Z(n13533)
         );
  AND U4508 ( .A(\SUBBYTES[7].a/w2291 ), .B(\SUBBYTES[7].a/w2278 ), .Z(n13532)
         );
  AND U4509 ( .A(\SUBBYTES[7].a/w2084 ), .B(\SUBBYTES[7].a/w2073 ), .Z(n13531)
         );
  AND U4510 ( .A(\SUBBYTES[7].a/w221 ), .B(\SUBBYTES[7].a/w210 ), .Z(n13513)
         );
  AND U4511 ( .A(n1839), .B(\SUBBYTES[6].a/w781 ), .Z(\SUBBYTES[6].a/w916 ) );
  AND U4512 ( .A(n1840), .B(\SUBBYTES[6].a/w782 ), .Z(\SUBBYTES[6].a/w914 ) );
  AND U4513 ( .A(\SUBBYTES[6].a/w912 ), .B(n1841), .Z(\SUBBYTES[6].a/w913 ) );
  ANDN U4514 ( .A(\w1[6][96] ), .B(n1842), .Z(\SUBBYTES[6].a/w909 ) );
  AND U4515 ( .A(n1843), .B(\SUBBYTES[6].a/w784 ), .Z(\SUBBYTES[6].a/w907 ) );
  AND U4516 ( .A(\SUBBYTES[6].a/w905 ), .B(n1844), .Z(\SUBBYTES[6].a/w906 ) );
  XOR U4517 ( .A(\SUBBYTES[6].a/w849 ), .B(n12238), .Z(n1844) );
  AND U4518 ( .A(\SUBBYTES[6].a/w892 ), .B(\SUBBYTES[6].a/w894 ), .Z(
        \SUBBYTES[6].a/w901 ) );
  AND U4519 ( .A(\SUBBYTES[6].a/w893 ), .B(\SUBBYTES[6].a/w895 ), .Z(
        \SUBBYTES[6].a/w899 ) );
  AND U4520 ( .A(\SUBBYTES[6].a/w896 ), .B(\SUBBYTES[6].a/w897 ), .Z(
        \SUBBYTES[6].a/w898 ) );
  AND U4521 ( .A(\SUBBYTES[6].a/w785 ), .B(n1839), .Z(\SUBBYTES[6].a/w884 ) );
  XOR U4522 ( .A(\SUBBYTES[6].a/w853 ), .B(n1040), .Z(n1839) );
  AND U4523 ( .A(\SUBBYTES[6].a/w786 ), .B(n1840), .Z(\SUBBYTES[6].a/w882 ) );
  XOR U4524 ( .A(n12239), .B(\SUBBYTES[6].a/w853 ), .Z(n1840) );
  ANDN U4525 ( .A(n1841), .B(n1845), .Z(\SUBBYTES[6].a/w881 ) );
  XOR U4526 ( .A(n1040), .B(n12239), .Z(n1841) );
  ANDN U4527 ( .A(\SUBBYTES[6].a/w787 ), .B(n1842), .Z(\SUBBYTES[6].a/w877 )
         );
  XNOR U4528 ( .A(\SUBBYTES[6].a/w846 ), .B(\SUBBYTES[6].a/w849 ), .Z(n1842)
         );
  AND U4529 ( .A(\SUBBYTES[6].a/w788 ), .B(n1843), .Z(\SUBBYTES[6].a/w875 ) );
  XNOR U4530 ( .A(n1846), .B(\SUBBYTES[6].a/w846 ), .Z(n1843) );
  AND U4531 ( .A(\SUBBYTES[6].a/w873 ), .B(n1847), .Z(\SUBBYTES[6].a/w874 ) );
  XOR U4532 ( .A(n1848), .B(n1846), .Z(n1847) );
  IV U4533 ( .A(n12238), .Z(n1846) );
  ANDN U4534 ( .A(\SUBBYTES[6].a/w892 ), .B(n1849), .Z(\SUBBYTES[6].a/w869 )
         );
  ANDN U4535 ( .A(\SUBBYTES[6].a/w893 ), .B(n1850), .Z(\SUBBYTES[6].a/w867 )
         );
  ANDN U4536 ( .A(\SUBBYTES[6].a/w896 ), .B(n1851), .Z(\SUBBYTES[6].a/w866 )
         );
  AND U4537 ( .A(\SUBBYTES[6].a/w852 ), .B(\SUBBYTES[6].a/w851 ), .Z(
        \SUBBYTES[6].a/w853 ) );
  IV U4538 ( .A(n1848), .Z(\SUBBYTES[6].a/w849 ) );
  NAND U4539 ( .A(\SUBBYTES[6].a/w828 ), .B(\SUBBYTES[6].a/w843 ), .Z(n1848)
         );
  AND U4540 ( .A(\SUBBYTES[6].a/w845 ), .B(\SUBBYTES[6].a/w851 ), .Z(
        \SUBBYTES[6].a/w846 ) );
  AND U4541 ( .A(\SUBBYTES[6].a/w830 ), .B(\SUBBYTES[6].a/w828 ), .Z(
        \SUBBYTES[6].a/w840 ) );
  AND U4542 ( .A(\SUBBYTES[6].a/w831 ), .B(\SUBBYTES[6].a/w829 ), .Z(
        \SUBBYTES[6].a/w838 ) );
  AND U4543 ( .A(\SUBBYTES[6].a/w845 ), .B(\SUBBYTES[6].a/w852 ), .Z(
        \SUBBYTES[6].a/w837 ) );
  AND U4544 ( .A(\SUBBYTES[6].a/w785 ), .B(\SUBBYTES[6].a/w781 ), .Z(
        \SUBBYTES[6].a/w822 ) );
  AND U4545 ( .A(\SUBBYTES[6].a/w786 ), .B(\SUBBYTES[6].a/w782 ), .Z(
        \SUBBYTES[6].a/w820 ) );
  ANDN U4546 ( .A(\SUBBYTES[6].a/w912 ), .B(n1845), .Z(\SUBBYTES[6].a/w819 )
         );
  XNOR U4547 ( .A(\w1[6][103] ), .B(\w1[6][97] ), .Z(n1845) );
  XOR U4548 ( .A(\w0[6][97] ), .B(g_input[865]), .Z(\w1[6][97] ) );
  IV U4549 ( .A(n1852), .Z(\w1[6][103] ) );
  AND U4550 ( .A(\w1[6][96] ), .B(\SUBBYTES[6].a/w787 ), .Z(
        \SUBBYTES[6].a/w815 ) );
  XOR U4551 ( .A(\w0[6][96] ), .B(g_input[864]), .Z(\w1[6][96] ) );
  AND U4552 ( .A(\SUBBYTES[6].a/w788 ), .B(\SUBBYTES[6].a/w784 ), .Z(
        \SUBBYTES[6].a/w813 ) );
  AND U4553 ( .A(\SUBBYTES[6].a/w873 ), .B(\SUBBYTES[6].a/w905 ), .Z(
        \SUBBYTES[6].a/w812 ) );
  ANDN U4554 ( .A(\SUBBYTES[6].a/w894 ), .B(n1849), .Z(\SUBBYTES[6].a/w807 )
         );
  XOR U4555 ( .A(\w1[6][100] ), .B(n1852), .Z(n1849) );
  ANDN U4556 ( .A(\SUBBYTES[6].a/w895 ), .B(n1850), .Z(\SUBBYTES[6].a/w805 )
         );
  XOR U4557 ( .A(n1852), .B(\w1[6][98] ), .Z(n1850) );
  XNOR U4558 ( .A(\w0[6][103] ), .B(g_input[871]), .Z(n1852) );
  ANDN U4559 ( .A(\SUBBYTES[6].a/w897 ), .B(n1851), .Z(\SUBBYTES[6].a/w804 )
         );
  XNOR U4560 ( .A(\w1[6][100] ), .B(\w1[6][98] ), .Z(n1851) );
  XOR U4561 ( .A(\w0[6][98] ), .B(g_input[866]), .Z(\w1[6][98] ) );
  XOR U4562 ( .A(\w0[6][100] ), .B(g_input[868]), .Z(\w1[6][100] ) );
  AND U4563 ( .A(n1853), .B(\SUBBYTES[6].a/w574 ), .Z(\SUBBYTES[6].a/w709 ) );
  AND U4564 ( .A(n1854), .B(\SUBBYTES[6].a/w575 ), .Z(\SUBBYTES[6].a/w707 ) );
  AND U4565 ( .A(\SUBBYTES[6].a/w705 ), .B(n1855), .Z(\SUBBYTES[6].a/w706 ) );
  ANDN U4566 ( .A(\w1[6][104] ), .B(n1856), .Z(\SUBBYTES[6].a/w702 ) );
  AND U4567 ( .A(n1857), .B(\SUBBYTES[6].a/w577 ), .Z(\SUBBYTES[6].a/w700 ) );
  AND U4568 ( .A(\SUBBYTES[6].a/w698 ), .B(n1858), .Z(\SUBBYTES[6].a/w699 ) );
  XOR U4569 ( .A(\SUBBYTES[6].a/w642 ), .B(n12236), .Z(n1858) );
  AND U4570 ( .A(\SUBBYTES[6].a/w685 ), .B(\SUBBYTES[6].a/w687 ), .Z(
        \SUBBYTES[6].a/w694 ) );
  AND U4571 ( .A(\SUBBYTES[6].a/w686 ), .B(\SUBBYTES[6].a/w688 ), .Z(
        \SUBBYTES[6].a/w692 ) );
  AND U4572 ( .A(\SUBBYTES[6].a/w689 ), .B(\SUBBYTES[6].a/w690 ), .Z(
        \SUBBYTES[6].a/w691 ) );
  AND U4573 ( .A(\SUBBYTES[6].a/w578 ), .B(n1853), .Z(\SUBBYTES[6].a/w677 ) );
  XOR U4574 ( .A(\SUBBYTES[6].a/w646 ), .B(n1039), .Z(n1853) );
  AND U4575 ( .A(\SUBBYTES[6].a/w579 ), .B(n1854), .Z(\SUBBYTES[6].a/w675 ) );
  XOR U4576 ( .A(n12237), .B(\SUBBYTES[6].a/w646 ), .Z(n1854) );
  ANDN U4577 ( .A(n1855), .B(n1859), .Z(\SUBBYTES[6].a/w674 ) );
  XOR U4578 ( .A(n1039), .B(n12237), .Z(n1855) );
  ANDN U4579 ( .A(\SUBBYTES[6].a/w580 ), .B(n1856), .Z(\SUBBYTES[6].a/w670 )
         );
  XNOR U4580 ( .A(\SUBBYTES[6].a/w639 ), .B(\SUBBYTES[6].a/w642 ), .Z(n1856)
         );
  AND U4581 ( .A(\SUBBYTES[6].a/w581 ), .B(n1857), .Z(\SUBBYTES[6].a/w668 ) );
  XNOR U4582 ( .A(n1860), .B(\SUBBYTES[6].a/w639 ), .Z(n1857) );
  AND U4583 ( .A(\SUBBYTES[6].a/w666 ), .B(n1861), .Z(\SUBBYTES[6].a/w667 ) );
  XOR U4584 ( .A(n1862), .B(n1860), .Z(n1861) );
  IV U4585 ( .A(n12236), .Z(n1860) );
  ANDN U4586 ( .A(\SUBBYTES[6].a/w685 ), .B(n1863), .Z(\SUBBYTES[6].a/w662 )
         );
  ANDN U4587 ( .A(\SUBBYTES[6].a/w686 ), .B(n1864), .Z(\SUBBYTES[6].a/w660 )
         );
  ANDN U4588 ( .A(\SUBBYTES[6].a/w689 ), .B(n1865), .Z(\SUBBYTES[6].a/w659 )
         );
  AND U4589 ( .A(\SUBBYTES[6].a/w645 ), .B(\SUBBYTES[6].a/w644 ), .Z(
        \SUBBYTES[6].a/w646 ) );
  IV U4590 ( .A(n1862), .Z(\SUBBYTES[6].a/w642 ) );
  NAND U4591 ( .A(\SUBBYTES[6].a/w621 ), .B(\SUBBYTES[6].a/w636 ), .Z(n1862)
         );
  AND U4592 ( .A(\SUBBYTES[6].a/w638 ), .B(\SUBBYTES[6].a/w644 ), .Z(
        \SUBBYTES[6].a/w639 ) );
  AND U4593 ( .A(\SUBBYTES[6].a/w623 ), .B(\SUBBYTES[6].a/w621 ), .Z(
        \SUBBYTES[6].a/w633 ) );
  AND U4594 ( .A(\SUBBYTES[6].a/w624 ), .B(\SUBBYTES[6].a/w622 ), .Z(
        \SUBBYTES[6].a/w631 ) );
  AND U4595 ( .A(\SUBBYTES[6].a/w638 ), .B(\SUBBYTES[6].a/w645 ), .Z(
        \SUBBYTES[6].a/w630 ) );
  AND U4596 ( .A(\SUBBYTES[6].a/w578 ), .B(\SUBBYTES[6].a/w574 ), .Z(
        \SUBBYTES[6].a/w615 ) );
  AND U4597 ( .A(\SUBBYTES[6].a/w579 ), .B(\SUBBYTES[6].a/w575 ), .Z(
        \SUBBYTES[6].a/w613 ) );
  ANDN U4598 ( .A(\SUBBYTES[6].a/w705 ), .B(n1859), .Z(\SUBBYTES[6].a/w612 )
         );
  XNOR U4599 ( .A(\w1[6][105] ), .B(\w1[6][111] ), .Z(n1859) );
  XOR U4600 ( .A(\w0[6][105] ), .B(g_input[873]), .Z(\w1[6][105] ) );
  AND U4601 ( .A(\w1[6][104] ), .B(\SUBBYTES[6].a/w580 ), .Z(
        \SUBBYTES[6].a/w608 ) );
  XOR U4602 ( .A(\w0[6][104] ), .B(g_input[872]), .Z(\w1[6][104] ) );
  AND U4603 ( .A(\SUBBYTES[6].a/w581 ), .B(\SUBBYTES[6].a/w577 ), .Z(
        \SUBBYTES[6].a/w606 ) );
  AND U4604 ( .A(\SUBBYTES[6].a/w666 ), .B(\SUBBYTES[6].a/w698 ), .Z(
        \SUBBYTES[6].a/w605 ) );
  ANDN U4605 ( .A(\SUBBYTES[6].a/w687 ), .B(n1863), .Z(\SUBBYTES[6].a/w600 )
         );
  XNOR U4606 ( .A(\w1[6][108] ), .B(\w1[6][111] ), .Z(n1863) );
  ANDN U4607 ( .A(\SUBBYTES[6].a/w688 ), .B(n1864), .Z(\SUBBYTES[6].a/w598 )
         );
  XNOR U4608 ( .A(\w1[6][106] ), .B(\w1[6][111] ), .Z(n1864) );
  XOR U4609 ( .A(\w0[6][111] ), .B(g_input[879]), .Z(\w1[6][111] ) );
  IV U4610 ( .A(n1866), .Z(\w1[6][106] ) );
  ANDN U4611 ( .A(\SUBBYTES[6].a/w690 ), .B(n1865), .Z(\SUBBYTES[6].a/w597 )
         );
  XOR U4612 ( .A(n1866), .B(\w1[6][108] ), .Z(n1865) );
  XOR U4613 ( .A(\w0[6][108] ), .B(g_input[876]), .Z(\w1[6][108] ) );
  XNOR U4614 ( .A(\w0[6][106] ), .B(g_input[874]), .Z(n1866) );
  AND U4615 ( .A(n1867), .B(\SUBBYTES[6].a/w367 ), .Z(\SUBBYTES[6].a/w502 ) );
  AND U4616 ( .A(n1868), .B(\SUBBYTES[6].a/w368 ), .Z(\SUBBYTES[6].a/w500 ) );
  AND U4617 ( .A(\SUBBYTES[6].a/w498 ), .B(n1869), .Z(\SUBBYTES[6].a/w499 ) );
  ANDN U4618 ( .A(\w1[6][112] ), .B(n1870), .Z(\SUBBYTES[6].a/w495 ) );
  AND U4619 ( .A(n1871), .B(\SUBBYTES[6].a/w370 ), .Z(\SUBBYTES[6].a/w493 ) );
  AND U4620 ( .A(\SUBBYTES[6].a/w491 ), .B(n1872), .Z(\SUBBYTES[6].a/w492 ) );
  XOR U4621 ( .A(\SUBBYTES[6].a/w435 ), .B(n12234), .Z(n1872) );
  AND U4622 ( .A(\SUBBYTES[6].a/w478 ), .B(\SUBBYTES[6].a/w480 ), .Z(
        \SUBBYTES[6].a/w487 ) );
  AND U4623 ( .A(\SUBBYTES[6].a/w479 ), .B(\SUBBYTES[6].a/w481 ), .Z(
        \SUBBYTES[6].a/w485 ) );
  AND U4624 ( .A(\SUBBYTES[6].a/w482 ), .B(\SUBBYTES[6].a/w483 ), .Z(
        \SUBBYTES[6].a/w484 ) );
  AND U4625 ( .A(\SUBBYTES[6].a/w371 ), .B(n1867), .Z(\SUBBYTES[6].a/w470 ) );
  XOR U4626 ( .A(\SUBBYTES[6].a/w439 ), .B(n1038), .Z(n1867) );
  AND U4627 ( .A(\SUBBYTES[6].a/w372 ), .B(n1868), .Z(\SUBBYTES[6].a/w468 ) );
  XOR U4628 ( .A(n12235), .B(\SUBBYTES[6].a/w439 ), .Z(n1868) );
  ANDN U4629 ( .A(n1869), .B(n1873), .Z(\SUBBYTES[6].a/w467 ) );
  XOR U4630 ( .A(n1038), .B(n12235), .Z(n1869) );
  ANDN U4631 ( .A(\SUBBYTES[6].a/w373 ), .B(n1870), .Z(\SUBBYTES[6].a/w463 )
         );
  XNOR U4632 ( .A(\SUBBYTES[6].a/w432 ), .B(\SUBBYTES[6].a/w435 ), .Z(n1870)
         );
  AND U4633 ( .A(\SUBBYTES[6].a/w374 ), .B(n1871), .Z(\SUBBYTES[6].a/w461 ) );
  XNOR U4634 ( .A(n1874), .B(\SUBBYTES[6].a/w432 ), .Z(n1871) );
  AND U4635 ( .A(\SUBBYTES[6].a/w459 ), .B(n1875), .Z(\SUBBYTES[6].a/w460 ) );
  XOR U4636 ( .A(n1876), .B(n1874), .Z(n1875) );
  IV U4637 ( .A(n12234), .Z(n1874) );
  ANDN U4638 ( .A(\SUBBYTES[6].a/w478 ), .B(n1877), .Z(\SUBBYTES[6].a/w455 )
         );
  ANDN U4639 ( .A(\SUBBYTES[6].a/w479 ), .B(n1878), .Z(\SUBBYTES[6].a/w453 )
         );
  ANDN U4640 ( .A(\SUBBYTES[6].a/w482 ), .B(n1879), .Z(\SUBBYTES[6].a/w452 )
         );
  AND U4641 ( .A(\SUBBYTES[6].a/w438 ), .B(\SUBBYTES[6].a/w437 ), .Z(
        \SUBBYTES[6].a/w439 ) );
  IV U4642 ( .A(n1876), .Z(\SUBBYTES[6].a/w435 ) );
  NAND U4643 ( .A(\SUBBYTES[6].a/w414 ), .B(\SUBBYTES[6].a/w429 ), .Z(n1876)
         );
  AND U4644 ( .A(\SUBBYTES[6].a/w431 ), .B(\SUBBYTES[6].a/w437 ), .Z(
        \SUBBYTES[6].a/w432 ) );
  AND U4645 ( .A(\SUBBYTES[6].a/w416 ), .B(\SUBBYTES[6].a/w414 ), .Z(
        \SUBBYTES[6].a/w426 ) );
  AND U4646 ( .A(\SUBBYTES[6].a/w417 ), .B(\SUBBYTES[6].a/w415 ), .Z(
        \SUBBYTES[6].a/w424 ) );
  AND U4647 ( .A(\SUBBYTES[6].a/w431 ), .B(\SUBBYTES[6].a/w438 ), .Z(
        \SUBBYTES[6].a/w423 ) );
  AND U4648 ( .A(\SUBBYTES[6].a/w371 ), .B(\SUBBYTES[6].a/w367 ), .Z(
        \SUBBYTES[6].a/w408 ) );
  AND U4649 ( .A(\SUBBYTES[6].a/w372 ), .B(\SUBBYTES[6].a/w368 ), .Z(
        \SUBBYTES[6].a/w406 ) );
  ANDN U4650 ( .A(\SUBBYTES[6].a/w498 ), .B(n1873), .Z(\SUBBYTES[6].a/w405 )
         );
  XNOR U4651 ( .A(\w1[6][113] ), .B(\w1[6][119] ), .Z(n1873) );
  XOR U4652 ( .A(\w0[6][113] ), .B(g_input[881]), .Z(\w1[6][113] ) );
  AND U4653 ( .A(\w1[6][112] ), .B(\SUBBYTES[6].a/w373 ), .Z(
        \SUBBYTES[6].a/w401 ) );
  XOR U4654 ( .A(\w0[6][112] ), .B(g_input[880]), .Z(\w1[6][112] ) );
  AND U4655 ( .A(\SUBBYTES[6].a/w374 ), .B(\SUBBYTES[6].a/w370 ), .Z(
        \SUBBYTES[6].a/w399 ) );
  AND U4656 ( .A(\SUBBYTES[6].a/w459 ), .B(\SUBBYTES[6].a/w491 ), .Z(
        \SUBBYTES[6].a/w398 ) );
  ANDN U4657 ( .A(\SUBBYTES[6].a/w480 ), .B(n1877), .Z(\SUBBYTES[6].a/w393 )
         );
  XNOR U4658 ( .A(\w1[6][116] ), .B(\w1[6][119] ), .Z(n1877) );
  ANDN U4659 ( .A(\SUBBYTES[6].a/w481 ), .B(n1878), .Z(\SUBBYTES[6].a/w391 )
         );
  XNOR U4660 ( .A(\w1[6][114] ), .B(\w1[6][119] ), .Z(n1878) );
  XOR U4661 ( .A(\w0[6][119] ), .B(g_input[887]), .Z(\w1[6][119] ) );
  IV U4662 ( .A(n1880), .Z(\w1[6][114] ) );
  ANDN U4663 ( .A(\SUBBYTES[6].a/w483 ), .B(n1879), .Z(\SUBBYTES[6].a/w390 )
         );
  XOR U4664 ( .A(n1880), .B(\w1[6][116] ), .Z(n1879) );
  XOR U4665 ( .A(\w0[6][116] ), .B(g_input[884]), .Z(\w1[6][116] ) );
  XNOR U4666 ( .A(\w0[6][114] ), .B(g_input[882]), .Z(n1880) );
  AND U4667 ( .A(n1881), .B(\SUBBYTES[6].a/w3265 ), .Z(\SUBBYTES[6].a/w3400 )
         );
  AND U4668 ( .A(n1882), .B(\SUBBYTES[6].a/w3266 ), .Z(\SUBBYTES[6].a/w3398 )
         );
  AND U4669 ( .A(\SUBBYTES[6].a/w3396 ), .B(n1883), .Z(\SUBBYTES[6].a/w3397 )
         );
  ANDN U4670 ( .A(\w1[6][0] ), .B(n1884), .Z(\SUBBYTES[6].a/w3393 ) );
  AND U4671 ( .A(n1885), .B(\SUBBYTES[6].a/w3268 ), .Z(\SUBBYTES[6].a/w3391 )
         );
  AND U4672 ( .A(\SUBBYTES[6].a/w3389 ), .B(n1886), .Z(\SUBBYTES[6].a/w3390 )
         );
  XOR U4673 ( .A(\SUBBYTES[6].a/w3333 ), .B(n12262), .Z(n1886) );
  AND U4674 ( .A(\SUBBYTES[6].a/w3376 ), .B(\SUBBYTES[6].a/w3378 ), .Z(
        \SUBBYTES[6].a/w3385 ) );
  AND U4675 ( .A(\SUBBYTES[6].a/w3377 ), .B(\SUBBYTES[6].a/w3379 ), .Z(
        \SUBBYTES[6].a/w3383 ) );
  AND U4676 ( .A(\SUBBYTES[6].a/w3380 ), .B(\SUBBYTES[6].a/w3381 ), .Z(
        \SUBBYTES[6].a/w3382 ) );
  AND U4677 ( .A(\SUBBYTES[6].a/w3269 ), .B(n1881), .Z(\SUBBYTES[6].a/w3368 )
         );
  XOR U4678 ( .A(\SUBBYTES[6].a/w3337 ), .B(n1052), .Z(n1881) );
  AND U4679 ( .A(\SUBBYTES[6].a/w3270 ), .B(n1882), .Z(\SUBBYTES[6].a/w3366 )
         );
  XOR U4680 ( .A(n12263), .B(\SUBBYTES[6].a/w3337 ), .Z(n1882) );
  ANDN U4681 ( .A(n1883), .B(n1887), .Z(\SUBBYTES[6].a/w3365 ) );
  XOR U4682 ( .A(n1052), .B(n12263), .Z(n1883) );
  ANDN U4683 ( .A(\SUBBYTES[6].a/w3271 ), .B(n1884), .Z(\SUBBYTES[6].a/w3361 )
         );
  XNOR U4684 ( .A(\SUBBYTES[6].a/w3330 ), .B(\SUBBYTES[6].a/w3333 ), .Z(n1884)
         );
  AND U4685 ( .A(\SUBBYTES[6].a/w3272 ), .B(n1885), .Z(\SUBBYTES[6].a/w3359 )
         );
  XNOR U4686 ( .A(n1888), .B(\SUBBYTES[6].a/w3330 ), .Z(n1885) );
  AND U4687 ( .A(\SUBBYTES[6].a/w3357 ), .B(n1889), .Z(\SUBBYTES[6].a/w3358 )
         );
  XOR U4688 ( .A(n1890), .B(n1888), .Z(n1889) );
  IV U4689 ( .A(n12262), .Z(n1888) );
  ANDN U4690 ( .A(\SUBBYTES[6].a/w3376 ), .B(n1891), .Z(\SUBBYTES[6].a/w3353 )
         );
  ANDN U4691 ( .A(\SUBBYTES[6].a/w3377 ), .B(n1892), .Z(\SUBBYTES[6].a/w3351 )
         );
  ANDN U4692 ( .A(\SUBBYTES[6].a/w3380 ), .B(n1893), .Z(\SUBBYTES[6].a/w3350 )
         );
  AND U4693 ( .A(\SUBBYTES[6].a/w3336 ), .B(\SUBBYTES[6].a/w3335 ), .Z(
        \SUBBYTES[6].a/w3337 ) );
  IV U4694 ( .A(n1890), .Z(\SUBBYTES[6].a/w3333 ) );
  NAND U4695 ( .A(\SUBBYTES[6].a/w3312 ), .B(\SUBBYTES[6].a/w3327 ), .Z(n1890)
         );
  AND U4696 ( .A(\SUBBYTES[6].a/w3329 ), .B(\SUBBYTES[6].a/w3335 ), .Z(
        \SUBBYTES[6].a/w3330 ) );
  AND U4697 ( .A(\SUBBYTES[6].a/w3314 ), .B(\SUBBYTES[6].a/w3312 ), .Z(
        \SUBBYTES[6].a/w3324 ) );
  AND U4698 ( .A(\SUBBYTES[6].a/w3315 ), .B(\SUBBYTES[6].a/w3313 ), .Z(
        \SUBBYTES[6].a/w3322 ) );
  AND U4699 ( .A(\SUBBYTES[6].a/w3329 ), .B(\SUBBYTES[6].a/w3336 ), .Z(
        \SUBBYTES[6].a/w3321 ) );
  AND U4700 ( .A(\SUBBYTES[6].a/w3269 ), .B(\SUBBYTES[6].a/w3265 ), .Z(
        \SUBBYTES[6].a/w3306 ) );
  AND U4701 ( .A(\SUBBYTES[6].a/w3270 ), .B(\SUBBYTES[6].a/w3266 ), .Z(
        \SUBBYTES[6].a/w3304 ) );
  ANDN U4702 ( .A(\SUBBYTES[6].a/w3396 ), .B(n1887), .Z(\SUBBYTES[6].a/w3303 )
         );
  XNOR U4703 ( .A(\w1[6][1] ), .B(\w1[6][7] ), .Z(n1887) );
  XOR U4704 ( .A(\w0[6][1] ), .B(g_input[769]), .Z(\w1[6][1] ) );
  AND U4705 ( .A(\w1[6][0] ), .B(\SUBBYTES[6].a/w3271 ), .Z(
        \SUBBYTES[6].a/w3299 ) );
  XOR U4706 ( .A(\w0[6][0] ), .B(g_input[768]), .Z(\w1[6][0] ) );
  AND U4707 ( .A(\SUBBYTES[6].a/w3272 ), .B(\SUBBYTES[6].a/w3268 ), .Z(
        \SUBBYTES[6].a/w3297 ) );
  AND U4708 ( .A(\SUBBYTES[6].a/w3357 ), .B(\SUBBYTES[6].a/w3389 ), .Z(
        \SUBBYTES[6].a/w3296 ) );
  ANDN U4709 ( .A(\SUBBYTES[6].a/w3378 ), .B(n1891), .Z(\SUBBYTES[6].a/w3291 )
         );
  XNOR U4710 ( .A(\w1[6][4] ), .B(\w1[6][7] ), .Z(n1891) );
  ANDN U4711 ( .A(\SUBBYTES[6].a/w3379 ), .B(n1892), .Z(\SUBBYTES[6].a/w3289 )
         );
  XNOR U4712 ( .A(\w1[6][2] ), .B(\w1[6][7] ), .Z(n1892) );
  XOR U4713 ( .A(\w0[6][7] ), .B(g_input[775]), .Z(\w1[6][7] ) );
  IV U4714 ( .A(n1894), .Z(\w1[6][2] ) );
  ANDN U4715 ( .A(\SUBBYTES[6].a/w3381 ), .B(n1893), .Z(\SUBBYTES[6].a/w3288 )
         );
  XOR U4716 ( .A(n1894), .B(\w1[6][4] ), .Z(n1893) );
  XOR U4717 ( .A(\w0[6][4] ), .B(g_input[772]), .Z(\w1[6][4] ) );
  XNOR U4718 ( .A(\w0[6][2] ), .B(g_input[770]), .Z(n1894) );
  AND U4719 ( .A(n1895), .B(\SUBBYTES[6].a/w3058 ), .Z(\SUBBYTES[6].a/w3193 )
         );
  AND U4720 ( .A(n1896), .B(\SUBBYTES[6].a/w3059 ), .Z(\SUBBYTES[6].a/w3191 )
         );
  AND U4721 ( .A(\SUBBYTES[6].a/w3189 ), .B(n1897), .Z(\SUBBYTES[6].a/w3190 )
         );
  ANDN U4722 ( .A(\w1[6][8] ), .B(n1898), .Z(\SUBBYTES[6].a/w3186 ) );
  AND U4723 ( .A(n1899), .B(\SUBBYTES[6].a/w3061 ), .Z(\SUBBYTES[6].a/w3184 )
         );
  AND U4724 ( .A(\SUBBYTES[6].a/w3182 ), .B(n1900), .Z(\SUBBYTES[6].a/w3183 )
         );
  XOR U4725 ( .A(\SUBBYTES[6].a/w3126 ), .B(n12260), .Z(n1900) );
  AND U4726 ( .A(\SUBBYTES[6].a/w3169 ), .B(\SUBBYTES[6].a/w3171 ), .Z(
        \SUBBYTES[6].a/w3178 ) );
  AND U4727 ( .A(\SUBBYTES[6].a/w3170 ), .B(\SUBBYTES[6].a/w3172 ), .Z(
        \SUBBYTES[6].a/w3176 ) );
  AND U4728 ( .A(\SUBBYTES[6].a/w3173 ), .B(\SUBBYTES[6].a/w3174 ), .Z(
        \SUBBYTES[6].a/w3175 ) );
  AND U4729 ( .A(\SUBBYTES[6].a/w3062 ), .B(n1895), .Z(\SUBBYTES[6].a/w3161 )
         );
  XOR U4730 ( .A(\SUBBYTES[6].a/w3130 ), .B(n1051), .Z(n1895) );
  AND U4731 ( .A(\SUBBYTES[6].a/w3063 ), .B(n1896), .Z(\SUBBYTES[6].a/w3159 )
         );
  XOR U4732 ( .A(n12261), .B(\SUBBYTES[6].a/w3130 ), .Z(n1896) );
  ANDN U4733 ( .A(n1897), .B(n1901), .Z(\SUBBYTES[6].a/w3158 ) );
  XOR U4734 ( .A(n1051), .B(n12261), .Z(n1897) );
  ANDN U4735 ( .A(\SUBBYTES[6].a/w3064 ), .B(n1898), .Z(\SUBBYTES[6].a/w3154 )
         );
  XNOR U4736 ( .A(\SUBBYTES[6].a/w3123 ), .B(\SUBBYTES[6].a/w3126 ), .Z(n1898)
         );
  AND U4737 ( .A(\SUBBYTES[6].a/w3065 ), .B(n1899), .Z(\SUBBYTES[6].a/w3152 )
         );
  XNOR U4738 ( .A(n1902), .B(\SUBBYTES[6].a/w3123 ), .Z(n1899) );
  AND U4739 ( .A(\SUBBYTES[6].a/w3150 ), .B(n1903), .Z(\SUBBYTES[6].a/w3151 )
         );
  XOR U4740 ( .A(n1904), .B(n1902), .Z(n1903) );
  IV U4741 ( .A(n12260), .Z(n1902) );
  ANDN U4742 ( .A(\SUBBYTES[6].a/w3169 ), .B(n1905), .Z(\SUBBYTES[6].a/w3146 )
         );
  ANDN U4743 ( .A(\SUBBYTES[6].a/w3170 ), .B(n1906), .Z(\SUBBYTES[6].a/w3144 )
         );
  ANDN U4744 ( .A(\SUBBYTES[6].a/w3173 ), .B(n1907), .Z(\SUBBYTES[6].a/w3143 )
         );
  AND U4745 ( .A(\SUBBYTES[6].a/w3129 ), .B(\SUBBYTES[6].a/w3128 ), .Z(
        \SUBBYTES[6].a/w3130 ) );
  IV U4746 ( .A(n1904), .Z(\SUBBYTES[6].a/w3126 ) );
  NAND U4747 ( .A(\SUBBYTES[6].a/w3105 ), .B(\SUBBYTES[6].a/w3120 ), .Z(n1904)
         );
  AND U4748 ( .A(\SUBBYTES[6].a/w3122 ), .B(\SUBBYTES[6].a/w3128 ), .Z(
        \SUBBYTES[6].a/w3123 ) );
  AND U4749 ( .A(\SUBBYTES[6].a/w3107 ), .B(\SUBBYTES[6].a/w3105 ), .Z(
        \SUBBYTES[6].a/w3117 ) );
  AND U4750 ( .A(\SUBBYTES[6].a/w3108 ), .B(\SUBBYTES[6].a/w3106 ), .Z(
        \SUBBYTES[6].a/w3115 ) );
  AND U4751 ( .A(\SUBBYTES[6].a/w3122 ), .B(\SUBBYTES[6].a/w3129 ), .Z(
        \SUBBYTES[6].a/w3114 ) );
  AND U4752 ( .A(\SUBBYTES[6].a/w3062 ), .B(\SUBBYTES[6].a/w3058 ), .Z(
        \SUBBYTES[6].a/w3099 ) );
  AND U4753 ( .A(\SUBBYTES[6].a/w3063 ), .B(\SUBBYTES[6].a/w3059 ), .Z(
        \SUBBYTES[6].a/w3097 ) );
  ANDN U4754 ( .A(\SUBBYTES[6].a/w3189 ), .B(n1901), .Z(\SUBBYTES[6].a/w3096 )
         );
  XNOR U4755 ( .A(\w1[6][15] ), .B(\w1[6][9] ), .Z(n1901) );
  XOR U4756 ( .A(\w0[6][9] ), .B(g_input[777]), .Z(\w1[6][9] ) );
  AND U4757 ( .A(\w1[6][8] ), .B(\SUBBYTES[6].a/w3064 ), .Z(
        \SUBBYTES[6].a/w3092 ) );
  XOR U4758 ( .A(\w0[6][8] ), .B(g_input[776]), .Z(\w1[6][8] ) );
  AND U4759 ( .A(\SUBBYTES[6].a/w3065 ), .B(\SUBBYTES[6].a/w3061 ), .Z(
        \SUBBYTES[6].a/w3090 ) );
  AND U4760 ( .A(\SUBBYTES[6].a/w3150 ), .B(\SUBBYTES[6].a/w3182 ), .Z(
        \SUBBYTES[6].a/w3089 ) );
  ANDN U4761 ( .A(\SUBBYTES[6].a/w3171 ), .B(n1905), .Z(\SUBBYTES[6].a/w3084 )
         );
  XNOR U4762 ( .A(\w1[6][12] ), .B(\w1[6][15] ), .Z(n1905) );
  ANDN U4763 ( .A(\SUBBYTES[6].a/w3172 ), .B(n1906), .Z(\SUBBYTES[6].a/w3082 )
         );
  XNOR U4764 ( .A(\w1[6][10] ), .B(\w1[6][15] ), .Z(n1906) );
  XOR U4765 ( .A(\w0[6][15] ), .B(g_input[783]), .Z(\w1[6][15] ) );
  ANDN U4766 ( .A(\SUBBYTES[6].a/w3174 ), .B(n1907), .Z(\SUBBYTES[6].a/w3081 )
         );
  XNOR U4767 ( .A(\w1[6][10] ), .B(\w1[6][12] ), .Z(n1907) );
  XOR U4768 ( .A(\w0[6][12] ), .B(g_input[780]), .Z(\w1[6][12] ) );
  XOR U4769 ( .A(\w0[6][10] ), .B(g_input[778]), .Z(\w1[6][10] ) );
  AND U4770 ( .A(n1908), .B(\SUBBYTES[6].a/w2851 ), .Z(\SUBBYTES[6].a/w2986 )
         );
  AND U4771 ( .A(n1909), .B(\SUBBYTES[6].a/w2852 ), .Z(\SUBBYTES[6].a/w2984 )
         );
  AND U4772 ( .A(\SUBBYTES[6].a/w2982 ), .B(n1910), .Z(\SUBBYTES[6].a/w2983 )
         );
  ANDN U4773 ( .A(\w1[6][16] ), .B(n1911), .Z(\SUBBYTES[6].a/w2979 ) );
  AND U4774 ( .A(n1912), .B(\SUBBYTES[6].a/w2854 ), .Z(\SUBBYTES[6].a/w2977 )
         );
  AND U4775 ( .A(\SUBBYTES[6].a/w2975 ), .B(n1913), .Z(\SUBBYTES[6].a/w2976 )
         );
  XOR U4776 ( .A(\SUBBYTES[6].a/w2919 ), .B(n12258), .Z(n1913) );
  AND U4777 ( .A(\SUBBYTES[6].a/w2962 ), .B(\SUBBYTES[6].a/w2964 ), .Z(
        \SUBBYTES[6].a/w2971 ) );
  AND U4778 ( .A(\SUBBYTES[6].a/w2963 ), .B(\SUBBYTES[6].a/w2965 ), .Z(
        \SUBBYTES[6].a/w2969 ) );
  AND U4779 ( .A(\SUBBYTES[6].a/w2966 ), .B(\SUBBYTES[6].a/w2967 ), .Z(
        \SUBBYTES[6].a/w2968 ) );
  AND U4780 ( .A(\SUBBYTES[6].a/w2855 ), .B(n1908), .Z(\SUBBYTES[6].a/w2954 )
         );
  XOR U4781 ( .A(\SUBBYTES[6].a/w2923 ), .B(n1050), .Z(n1908) );
  AND U4782 ( .A(\SUBBYTES[6].a/w2856 ), .B(n1909), .Z(\SUBBYTES[6].a/w2952 )
         );
  XOR U4783 ( .A(n12259), .B(\SUBBYTES[6].a/w2923 ), .Z(n1909) );
  ANDN U4784 ( .A(n1910), .B(n1914), .Z(\SUBBYTES[6].a/w2951 ) );
  XOR U4785 ( .A(n1050), .B(n12259), .Z(n1910) );
  AND U4786 ( .A(n1915), .B(\SUBBYTES[6].a/w160 ), .Z(\SUBBYTES[6].a/w295 ) );
  ANDN U4787 ( .A(\SUBBYTES[6].a/w2857 ), .B(n1911), .Z(\SUBBYTES[6].a/w2947 )
         );
  XNOR U4788 ( .A(\SUBBYTES[6].a/w2916 ), .B(\SUBBYTES[6].a/w2919 ), .Z(n1911)
         );
  AND U4789 ( .A(\SUBBYTES[6].a/w2858 ), .B(n1912), .Z(\SUBBYTES[6].a/w2945 )
         );
  XNOR U4790 ( .A(n1916), .B(\SUBBYTES[6].a/w2916 ), .Z(n1912) );
  AND U4791 ( .A(\SUBBYTES[6].a/w2943 ), .B(n1917), .Z(\SUBBYTES[6].a/w2944 )
         );
  XOR U4792 ( .A(n1918), .B(n1916), .Z(n1917) );
  IV U4793 ( .A(n12258), .Z(n1916) );
  ANDN U4794 ( .A(\SUBBYTES[6].a/w2962 ), .B(n1919), .Z(\SUBBYTES[6].a/w2939 )
         );
  ANDN U4795 ( .A(\SUBBYTES[6].a/w2963 ), .B(n1920), .Z(\SUBBYTES[6].a/w2937 )
         );
  ANDN U4796 ( .A(\SUBBYTES[6].a/w2966 ), .B(n1921), .Z(\SUBBYTES[6].a/w2936 )
         );
  AND U4797 ( .A(n1922), .B(\SUBBYTES[6].a/w161 ), .Z(\SUBBYTES[6].a/w293 ) );
  AND U4798 ( .A(\SUBBYTES[6].a/w2922 ), .B(\SUBBYTES[6].a/w2921 ), .Z(
        \SUBBYTES[6].a/w2923 ) );
  AND U4799 ( .A(\SUBBYTES[6].a/w291 ), .B(n1923), .Z(\SUBBYTES[6].a/w292 ) );
  IV U4800 ( .A(n1918), .Z(\SUBBYTES[6].a/w2919 ) );
  NAND U4801 ( .A(\SUBBYTES[6].a/w2898 ), .B(\SUBBYTES[6].a/w2913 ), .Z(n1918)
         );
  AND U4802 ( .A(\SUBBYTES[6].a/w2915 ), .B(\SUBBYTES[6].a/w2921 ), .Z(
        \SUBBYTES[6].a/w2916 ) );
  AND U4803 ( .A(\SUBBYTES[6].a/w2900 ), .B(\SUBBYTES[6].a/w2898 ), .Z(
        \SUBBYTES[6].a/w2910 ) );
  AND U4804 ( .A(\SUBBYTES[6].a/w2901 ), .B(\SUBBYTES[6].a/w2899 ), .Z(
        \SUBBYTES[6].a/w2908 ) );
  AND U4805 ( .A(\SUBBYTES[6].a/w2915 ), .B(\SUBBYTES[6].a/w2922 ), .Z(
        \SUBBYTES[6].a/w2907 ) );
  AND U4806 ( .A(\SUBBYTES[6].a/w2855 ), .B(\SUBBYTES[6].a/w2851 ), .Z(
        \SUBBYTES[6].a/w2892 ) );
  AND U4807 ( .A(\SUBBYTES[6].a/w2856 ), .B(\SUBBYTES[6].a/w2852 ), .Z(
        \SUBBYTES[6].a/w2890 ) );
  ANDN U4808 ( .A(\SUBBYTES[6].a/w2982 ), .B(n1914), .Z(\SUBBYTES[6].a/w2889 )
         );
  XNOR U4809 ( .A(\w1[6][17] ), .B(\w1[6][23] ), .Z(n1914) );
  XOR U4810 ( .A(\w0[6][17] ), .B(g_input[785]), .Z(\w1[6][17] ) );
  AND U4811 ( .A(\w1[6][16] ), .B(\SUBBYTES[6].a/w2857 ), .Z(
        \SUBBYTES[6].a/w2885 ) );
  XOR U4812 ( .A(\w0[6][16] ), .B(g_input[784]), .Z(\w1[6][16] ) );
  AND U4813 ( .A(\SUBBYTES[6].a/w2858 ), .B(\SUBBYTES[6].a/w2854 ), .Z(
        \SUBBYTES[6].a/w2883 ) );
  AND U4814 ( .A(\SUBBYTES[6].a/w2943 ), .B(\SUBBYTES[6].a/w2975 ), .Z(
        \SUBBYTES[6].a/w2882 ) );
  ANDN U4815 ( .A(\w1[6][120] ), .B(n1924), .Z(\SUBBYTES[6].a/w288 ) );
  ANDN U4816 ( .A(\SUBBYTES[6].a/w2964 ), .B(n1919), .Z(\SUBBYTES[6].a/w2877 )
         );
  XNOR U4817 ( .A(\w1[6][20] ), .B(\w1[6][23] ), .Z(n1919) );
  ANDN U4818 ( .A(\SUBBYTES[6].a/w2965 ), .B(n1920), .Z(\SUBBYTES[6].a/w2875 )
         );
  XNOR U4819 ( .A(\w1[6][18] ), .B(\w1[6][23] ), .Z(n1920) );
  XOR U4820 ( .A(\w0[6][23] ), .B(g_input[791]), .Z(\w1[6][23] ) );
  IV U4821 ( .A(n1925), .Z(\w1[6][18] ) );
  ANDN U4822 ( .A(\SUBBYTES[6].a/w2967 ), .B(n1921), .Z(\SUBBYTES[6].a/w2874 )
         );
  XOR U4823 ( .A(n1925), .B(\w1[6][20] ), .Z(n1921) );
  XOR U4824 ( .A(\w0[6][20] ), .B(g_input[788]), .Z(\w1[6][20] ) );
  XNOR U4825 ( .A(\w0[6][18] ), .B(g_input[786]), .Z(n1925) );
  AND U4826 ( .A(n1926), .B(\SUBBYTES[6].a/w163 ), .Z(\SUBBYTES[6].a/w286 ) );
  AND U4827 ( .A(\SUBBYTES[6].a/w284 ), .B(n1927), .Z(\SUBBYTES[6].a/w285 ) );
  XOR U4828 ( .A(\SUBBYTES[6].a/w228 ), .B(n12232), .Z(n1927) );
  AND U4829 ( .A(\SUBBYTES[6].a/w271 ), .B(\SUBBYTES[6].a/w273 ), .Z(
        \SUBBYTES[6].a/w280 ) );
  AND U4830 ( .A(\SUBBYTES[6].a/w272 ), .B(\SUBBYTES[6].a/w274 ), .Z(
        \SUBBYTES[6].a/w278 ) );
  AND U4831 ( .A(n1928), .B(\SUBBYTES[6].a/w2644 ), .Z(\SUBBYTES[6].a/w2779 )
         );
  AND U4832 ( .A(n1929), .B(\SUBBYTES[6].a/w2645 ), .Z(\SUBBYTES[6].a/w2777 )
         );
  AND U4833 ( .A(\SUBBYTES[6].a/w2775 ), .B(n1930), .Z(\SUBBYTES[6].a/w2776 )
         );
  ANDN U4834 ( .A(\w1[6][24] ), .B(n1931), .Z(\SUBBYTES[6].a/w2772 ) );
  AND U4835 ( .A(n1932), .B(\SUBBYTES[6].a/w2647 ), .Z(\SUBBYTES[6].a/w2770 )
         );
  AND U4836 ( .A(\SUBBYTES[6].a/w275 ), .B(\SUBBYTES[6].a/w276 ), .Z(
        \SUBBYTES[6].a/w277 ) );
  AND U4837 ( .A(\SUBBYTES[6].a/w2768 ), .B(n1933), .Z(\SUBBYTES[6].a/w2769 )
         );
  XOR U4838 ( .A(\SUBBYTES[6].a/w2712 ), .B(n12256), .Z(n1933) );
  AND U4839 ( .A(\SUBBYTES[6].a/w2755 ), .B(\SUBBYTES[6].a/w2757 ), .Z(
        \SUBBYTES[6].a/w2764 ) );
  AND U4840 ( .A(\SUBBYTES[6].a/w2756 ), .B(\SUBBYTES[6].a/w2758 ), .Z(
        \SUBBYTES[6].a/w2762 ) );
  AND U4841 ( .A(\SUBBYTES[6].a/w2759 ), .B(\SUBBYTES[6].a/w2760 ), .Z(
        \SUBBYTES[6].a/w2761 ) );
  AND U4842 ( .A(\SUBBYTES[6].a/w2648 ), .B(n1928), .Z(\SUBBYTES[6].a/w2747 )
         );
  XOR U4843 ( .A(\SUBBYTES[6].a/w2716 ), .B(n1049), .Z(n1928) );
  AND U4844 ( .A(\SUBBYTES[6].a/w2649 ), .B(n1929), .Z(\SUBBYTES[6].a/w2745 )
         );
  XOR U4845 ( .A(n12257), .B(\SUBBYTES[6].a/w2716 ), .Z(n1929) );
  ANDN U4846 ( .A(n1930), .B(n1934), .Z(\SUBBYTES[6].a/w2744 ) );
  XOR U4847 ( .A(n1049), .B(n12257), .Z(n1930) );
  ANDN U4848 ( .A(\SUBBYTES[6].a/w2650 ), .B(n1931), .Z(\SUBBYTES[6].a/w2740 )
         );
  XNOR U4849 ( .A(\SUBBYTES[6].a/w2709 ), .B(\SUBBYTES[6].a/w2712 ), .Z(n1931)
         );
  AND U4850 ( .A(\SUBBYTES[6].a/w2651 ), .B(n1932), .Z(\SUBBYTES[6].a/w2738 )
         );
  XNOR U4851 ( .A(n1935), .B(\SUBBYTES[6].a/w2709 ), .Z(n1932) );
  AND U4852 ( .A(\SUBBYTES[6].a/w2736 ), .B(n1936), .Z(\SUBBYTES[6].a/w2737 )
         );
  XOR U4853 ( .A(n1937), .B(n1935), .Z(n1936) );
  IV U4854 ( .A(n12256), .Z(n1935) );
  ANDN U4855 ( .A(\SUBBYTES[6].a/w2755 ), .B(n1938), .Z(\SUBBYTES[6].a/w2732 )
         );
  ANDN U4856 ( .A(\SUBBYTES[6].a/w2756 ), .B(n1939), .Z(\SUBBYTES[6].a/w2730 )
         );
  ANDN U4857 ( .A(\SUBBYTES[6].a/w2759 ), .B(n1940), .Z(\SUBBYTES[6].a/w2729 )
         );
  AND U4858 ( .A(\SUBBYTES[6].a/w2715 ), .B(\SUBBYTES[6].a/w2714 ), .Z(
        \SUBBYTES[6].a/w2716 ) );
  IV U4859 ( .A(n1937), .Z(\SUBBYTES[6].a/w2712 ) );
  NAND U4860 ( .A(\SUBBYTES[6].a/w2691 ), .B(\SUBBYTES[6].a/w2706 ), .Z(n1937)
         );
  AND U4861 ( .A(\SUBBYTES[6].a/w2708 ), .B(\SUBBYTES[6].a/w2714 ), .Z(
        \SUBBYTES[6].a/w2709 ) );
  AND U4862 ( .A(\SUBBYTES[6].a/w2693 ), .B(\SUBBYTES[6].a/w2691 ), .Z(
        \SUBBYTES[6].a/w2703 ) );
  AND U4863 ( .A(\SUBBYTES[6].a/w2694 ), .B(\SUBBYTES[6].a/w2692 ), .Z(
        \SUBBYTES[6].a/w2701 ) );
  AND U4864 ( .A(\SUBBYTES[6].a/w2708 ), .B(\SUBBYTES[6].a/w2715 ), .Z(
        \SUBBYTES[6].a/w2700 ) );
  AND U4865 ( .A(\SUBBYTES[6].a/w2648 ), .B(\SUBBYTES[6].a/w2644 ), .Z(
        \SUBBYTES[6].a/w2685 ) );
  AND U4866 ( .A(\SUBBYTES[6].a/w2649 ), .B(\SUBBYTES[6].a/w2645 ), .Z(
        \SUBBYTES[6].a/w2683 ) );
  ANDN U4867 ( .A(\SUBBYTES[6].a/w2775 ), .B(n1934), .Z(\SUBBYTES[6].a/w2682 )
         );
  XNOR U4868 ( .A(\w1[6][25] ), .B(\w1[6][31] ), .Z(n1934) );
  XOR U4869 ( .A(\w0[6][25] ), .B(g_input[793]), .Z(\w1[6][25] ) );
  AND U4870 ( .A(\w1[6][24] ), .B(\SUBBYTES[6].a/w2650 ), .Z(
        \SUBBYTES[6].a/w2678 ) );
  XOR U4871 ( .A(\w0[6][24] ), .B(g_input[792]), .Z(\w1[6][24] ) );
  AND U4872 ( .A(\SUBBYTES[6].a/w2651 ), .B(\SUBBYTES[6].a/w2647 ), .Z(
        \SUBBYTES[6].a/w2676 ) );
  AND U4873 ( .A(\SUBBYTES[6].a/w2736 ), .B(\SUBBYTES[6].a/w2768 ), .Z(
        \SUBBYTES[6].a/w2675 ) );
  ANDN U4874 ( .A(\SUBBYTES[6].a/w2757 ), .B(n1938), .Z(\SUBBYTES[6].a/w2670 )
         );
  XNOR U4875 ( .A(\w1[6][28] ), .B(\w1[6][31] ), .Z(n1938) );
  ANDN U4876 ( .A(\SUBBYTES[6].a/w2758 ), .B(n1939), .Z(\SUBBYTES[6].a/w2668 )
         );
  XNOR U4877 ( .A(\w1[6][26] ), .B(\w1[6][31] ), .Z(n1939) );
  XOR U4878 ( .A(\w0[6][31] ), .B(g_input[799]), .Z(\w1[6][31] ) );
  IV U4879 ( .A(n1941), .Z(\w1[6][26] ) );
  ANDN U4880 ( .A(\SUBBYTES[6].a/w2760 ), .B(n1940), .Z(\SUBBYTES[6].a/w2667 )
         );
  XOR U4881 ( .A(n1941), .B(\w1[6][28] ), .Z(n1940) );
  XOR U4882 ( .A(\w0[6][28] ), .B(g_input[796]), .Z(\w1[6][28] ) );
  XNOR U4883 ( .A(\w0[6][26] ), .B(g_input[794]), .Z(n1941) );
  AND U4884 ( .A(\SUBBYTES[6].a/w164 ), .B(n1915), .Z(\SUBBYTES[6].a/w263 ) );
  XOR U4885 ( .A(\SUBBYTES[6].a/w232 ), .B(n1037), .Z(n1915) );
  AND U4886 ( .A(\SUBBYTES[6].a/w165 ), .B(n1922), .Z(\SUBBYTES[6].a/w261 ) );
  XOR U4887 ( .A(n12233), .B(\SUBBYTES[6].a/w232 ), .Z(n1922) );
  ANDN U4888 ( .A(n1923), .B(n1942), .Z(\SUBBYTES[6].a/w260 ) );
  XOR U4889 ( .A(n1037), .B(n12233), .Z(n1923) );
  AND U4890 ( .A(n1943), .B(\SUBBYTES[6].a/w2437 ), .Z(\SUBBYTES[6].a/w2572 )
         );
  AND U4891 ( .A(n1944), .B(\SUBBYTES[6].a/w2438 ), .Z(\SUBBYTES[6].a/w2570 )
         );
  AND U4892 ( .A(\SUBBYTES[6].a/w2568 ), .B(n1945), .Z(\SUBBYTES[6].a/w2569 )
         );
  ANDN U4893 ( .A(\w1[6][32] ), .B(n1946), .Z(\SUBBYTES[6].a/w2565 ) );
  AND U4894 ( .A(n1947), .B(\SUBBYTES[6].a/w2440 ), .Z(\SUBBYTES[6].a/w2563 )
         );
  AND U4895 ( .A(\SUBBYTES[6].a/w2561 ), .B(n1948), .Z(\SUBBYTES[6].a/w2562 )
         );
  XOR U4896 ( .A(\SUBBYTES[6].a/w2505 ), .B(n12254), .Z(n1948) );
  ANDN U4897 ( .A(\SUBBYTES[6].a/w166 ), .B(n1924), .Z(\SUBBYTES[6].a/w256 )
         );
  XNOR U4898 ( .A(\SUBBYTES[6].a/w225 ), .B(\SUBBYTES[6].a/w228 ), .Z(n1924)
         );
  AND U4899 ( .A(\SUBBYTES[6].a/w2548 ), .B(\SUBBYTES[6].a/w2550 ), .Z(
        \SUBBYTES[6].a/w2557 ) );
  AND U4900 ( .A(\SUBBYTES[6].a/w2549 ), .B(\SUBBYTES[6].a/w2551 ), .Z(
        \SUBBYTES[6].a/w2555 ) );
  AND U4901 ( .A(\SUBBYTES[6].a/w2552 ), .B(\SUBBYTES[6].a/w2553 ), .Z(
        \SUBBYTES[6].a/w2554 ) );
  AND U4902 ( .A(\SUBBYTES[6].a/w2441 ), .B(n1943), .Z(\SUBBYTES[6].a/w2540 )
         );
  XOR U4903 ( .A(\SUBBYTES[6].a/w2509 ), .B(n1048), .Z(n1943) );
  AND U4904 ( .A(\SUBBYTES[6].a/w167 ), .B(n1926), .Z(\SUBBYTES[6].a/w254 ) );
  XNOR U4905 ( .A(n1949), .B(\SUBBYTES[6].a/w225 ), .Z(n1926) );
  AND U4906 ( .A(\SUBBYTES[6].a/w2442 ), .B(n1944), .Z(\SUBBYTES[6].a/w2538 )
         );
  XOR U4907 ( .A(n12255), .B(\SUBBYTES[6].a/w2509 ), .Z(n1944) );
  ANDN U4908 ( .A(n1945), .B(n1950), .Z(\SUBBYTES[6].a/w2537 ) );
  XOR U4909 ( .A(n1048), .B(n12255), .Z(n1945) );
  ANDN U4910 ( .A(\SUBBYTES[6].a/w2443 ), .B(n1946), .Z(\SUBBYTES[6].a/w2533 )
         );
  XNOR U4911 ( .A(\SUBBYTES[6].a/w2502 ), .B(\SUBBYTES[6].a/w2505 ), .Z(n1946)
         );
  AND U4912 ( .A(\SUBBYTES[6].a/w2444 ), .B(n1947), .Z(\SUBBYTES[6].a/w2531 )
         );
  XNOR U4913 ( .A(n1951), .B(\SUBBYTES[6].a/w2502 ), .Z(n1947) );
  AND U4914 ( .A(\SUBBYTES[6].a/w2529 ), .B(n1952), .Z(\SUBBYTES[6].a/w2530 )
         );
  XOR U4915 ( .A(n1953), .B(n1951), .Z(n1952) );
  IV U4916 ( .A(n12254), .Z(n1951) );
  AND U4917 ( .A(\SUBBYTES[6].a/w252 ), .B(n1954), .Z(\SUBBYTES[6].a/w253 ) );
  XOR U4918 ( .A(n1955), .B(n1949), .Z(n1954) );
  IV U4919 ( .A(n12232), .Z(n1949) );
  ANDN U4920 ( .A(\SUBBYTES[6].a/w2548 ), .B(n1956), .Z(\SUBBYTES[6].a/w2525 )
         );
  ANDN U4921 ( .A(\SUBBYTES[6].a/w2549 ), .B(n1957), .Z(\SUBBYTES[6].a/w2523 )
         );
  ANDN U4922 ( .A(\SUBBYTES[6].a/w2552 ), .B(n1958), .Z(\SUBBYTES[6].a/w2522 )
         );
  AND U4923 ( .A(\SUBBYTES[6].a/w2508 ), .B(\SUBBYTES[6].a/w2507 ), .Z(
        \SUBBYTES[6].a/w2509 ) );
  IV U4924 ( .A(n1953), .Z(\SUBBYTES[6].a/w2505 ) );
  NAND U4925 ( .A(\SUBBYTES[6].a/w2484 ), .B(\SUBBYTES[6].a/w2499 ), .Z(n1953)
         );
  AND U4926 ( .A(\SUBBYTES[6].a/w2501 ), .B(\SUBBYTES[6].a/w2507 ), .Z(
        \SUBBYTES[6].a/w2502 ) );
  AND U4927 ( .A(\SUBBYTES[6].a/w2486 ), .B(\SUBBYTES[6].a/w2484 ), .Z(
        \SUBBYTES[6].a/w2496 ) );
  AND U4928 ( .A(\SUBBYTES[6].a/w2487 ), .B(\SUBBYTES[6].a/w2485 ), .Z(
        \SUBBYTES[6].a/w2494 ) );
  AND U4929 ( .A(\SUBBYTES[6].a/w2501 ), .B(\SUBBYTES[6].a/w2508 ), .Z(
        \SUBBYTES[6].a/w2493 ) );
  ANDN U4930 ( .A(\SUBBYTES[6].a/w271 ), .B(n1959), .Z(\SUBBYTES[6].a/w248 )
         );
  AND U4931 ( .A(\SUBBYTES[6].a/w2441 ), .B(\SUBBYTES[6].a/w2437 ), .Z(
        \SUBBYTES[6].a/w2478 ) );
  AND U4932 ( .A(\SUBBYTES[6].a/w2442 ), .B(\SUBBYTES[6].a/w2438 ), .Z(
        \SUBBYTES[6].a/w2476 ) );
  ANDN U4933 ( .A(\SUBBYTES[6].a/w2568 ), .B(n1950), .Z(\SUBBYTES[6].a/w2475 )
         );
  XNOR U4934 ( .A(\w1[6][33] ), .B(\w1[6][39] ), .Z(n1950) );
  XOR U4935 ( .A(\w0[6][33] ), .B(g_input[801]), .Z(\w1[6][33] ) );
  AND U4936 ( .A(\w1[6][32] ), .B(\SUBBYTES[6].a/w2443 ), .Z(
        \SUBBYTES[6].a/w2471 ) );
  XOR U4937 ( .A(\w0[6][32] ), .B(g_input[800]), .Z(\w1[6][32] ) );
  AND U4938 ( .A(\SUBBYTES[6].a/w2444 ), .B(\SUBBYTES[6].a/w2440 ), .Z(
        \SUBBYTES[6].a/w2469 ) );
  AND U4939 ( .A(\SUBBYTES[6].a/w2529 ), .B(\SUBBYTES[6].a/w2561 ), .Z(
        \SUBBYTES[6].a/w2468 ) );
  ANDN U4940 ( .A(\SUBBYTES[6].a/w2550 ), .B(n1956), .Z(\SUBBYTES[6].a/w2463 )
         );
  XNOR U4941 ( .A(\w1[6][36] ), .B(\w1[6][39] ), .Z(n1956) );
  ANDN U4942 ( .A(\SUBBYTES[6].a/w2551 ), .B(n1957), .Z(\SUBBYTES[6].a/w2461 )
         );
  XNOR U4943 ( .A(\w1[6][34] ), .B(\w1[6][39] ), .Z(n1957) );
  XOR U4944 ( .A(\w0[6][39] ), .B(g_input[807]), .Z(\w1[6][39] ) );
  IV U4945 ( .A(n1960), .Z(\w1[6][34] ) );
  ANDN U4946 ( .A(\SUBBYTES[6].a/w2553 ), .B(n1958), .Z(\SUBBYTES[6].a/w2460 )
         );
  XOR U4947 ( .A(n1960), .B(\w1[6][36] ), .Z(n1958) );
  XOR U4948 ( .A(\w0[6][36] ), .B(g_input[804]), .Z(\w1[6][36] ) );
  XNOR U4949 ( .A(\w0[6][34] ), .B(g_input[802]), .Z(n1960) );
  ANDN U4950 ( .A(\SUBBYTES[6].a/w272 ), .B(n1961), .Z(\SUBBYTES[6].a/w246 )
         );
  ANDN U4951 ( .A(\SUBBYTES[6].a/w275 ), .B(n1962), .Z(\SUBBYTES[6].a/w245 )
         );
  AND U4952 ( .A(n1963), .B(\SUBBYTES[6].a/w2230 ), .Z(\SUBBYTES[6].a/w2365 )
         );
  AND U4953 ( .A(n1964), .B(\SUBBYTES[6].a/w2231 ), .Z(\SUBBYTES[6].a/w2363 )
         );
  AND U4954 ( .A(\SUBBYTES[6].a/w2361 ), .B(n1965), .Z(\SUBBYTES[6].a/w2362 )
         );
  ANDN U4955 ( .A(\w1[6][40] ), .B(n1966), .Z(\SUBBYTES[6].a/w2358 ) );
  AND U4956 ( .A(n1967), .B(\SUBBYTES[6].a/w2233 ), .Z(\SUBBYTES[6].a/w2356 )
         );
  AND U4957 ( .A(\SUBBYTES[6].a/w2354 ), .B(n1968), .Z(\SUBBYTES[6].a/w2355 )
         );
  XOR U4958 ( .A(\SUBBYTES[6].a/w2298 ), .B(n12252), .Z(n1968) );
  AND U4959 ( .A(\SUBBYTES[6].a/w2341 ), .B(\SUBBYTES[6].a/w2343 ), .Z(
        \SUBBYTES[6].a/w2350 ) );
  AND U4960 ( .A(\SUBBYTES[6].a/w2342 ), .B(\SUBBYTES[6].a/w2344 ), .Z(
        \SUBBYTES[6].a/w2348 ) );
  AND U4961 ( .A(\SUBBYTES[6].a/w2345 ), .B(\SUBBYTES[6].a/w2346 ), .Z(
        \SUBBYTES[6].a/w2347 ) );
  AND U4962 ( .A(\SUBBYTES[6].a/w2234 ), .B(n1963), .Z(\SUBBYTES[6].a/w2333 )
         );
  XOR U4963 ( .A(\SUBBYTES[6].a/w2302 ), .B(n1047), .Z(n1963) );
  AND U4964 ( .A(\SUBBYTES[6].a/w2235 ), .B(n1964), .Z(\SUBBYTES[6].a/w2331 )
         );
  XOR U4965 ( .A(n12253), .B(\SUBBYTES[6].a/w2302 ), .Z(n1964) );
  ANDN U4966 ( .A(n1965), .B(n1969), .Z(\SUBBYTES[6].a/w2330 ) );
  XOR U4967 ( .A(n1047), .B(n12253), .Z(n1965) );
  ANDN U4968 ( .A(\SUBBYTES[6].a/w2236 ), .B(n1966), .Z(\SUBBYTES[6].a/w2326 )
         );
  XNOR U4969 ( .A(\SUBBYTES[6].a/w2295 ), .B(\SUBBYTES[6].a/w2298 ), .Z(n1966)
         );
  AND U4970 ( .A(\SUBBYTES[6].a/w2237 ), .B(n1967), .Z(\SUBBYTES[6].a/w2324 )
         );
  XNOR U4971 ( .A(n1970), .B(\SUBBYTES[6].a/w2295 ), .Z(n1967) );
  AND U4972 ( .A(\SUBBYTES[6].a/w2322 ), .B(n1971), .Z(\SUBBYTES[6].a/w2323 )
         );
  XOR U4973 ( .A(n1972), .B(n1970), .Z(n1971) );
  IV U4974 ( .A(n12252), .Z(n1970) );
  AND U4975 ( .A(\SUBBYTES[6].a/w231 ), .B(\SUBBYTES[6].a/w230 ), .Z(
        \SUBBYTES[6].a/w232 ) );
  ANDN U4976 ( .A(\SUBBYTES[6].a/w2341 ), .B(n1973), .Z(\SUBBYTES[6].a/w2318 )
         );
  ANDN U4977 ( .A(\SUBBYTES[6].a/w2342 ), .B(n1974), .Z(\SUBBYTES[6].a/w2316 )
         );
  ANDN U4978 ( .A(\SUBBYTES[6].a/w2345 ), .B(n1975), .Z(\SUBBYTES[6].a/w2315 )
         );
  AND U4979 ( .A(\SUBBYTES[6].a/w2301 ), .B(\SUBBYTES[6].a/w2300 ), .Z(
        \SUBBYTES[6].a/w2302 ) );
  IV U4980 ( .A(n1972), .Z(\SUBBYTES[6].a/w2298 ) );
  NAND U4981 ( .A(\SUBBYTES[6].a/w2277 ), .B(\SUBBYTES[6].a/w2292 ), .Z(n1972)
         );
  AND U4982 ( .A(\SUBBYTES[6].a/w2294 ), .B(\SUBBYTES[6].a/w2300 ), .Z(
        \SUBBYTES[6].a/w2295 ) );
  AND U4983 ( .A(\SUBBYTES[6].a/w2279 ), .B(\SUBBYTES[6].a/w2277 ), .Z(
        \SUBBYTES[6].a/w2289 ) );
  AND U4984 ( .A(\SUBBYTES[6].a/w2280 ), .B(\SUBBYTES[6].a/w2278 ), .Z(
        \SUBBYTES[6].a/w2287 ) );
  AND U4985 ( .A(\SUBBYTES[6].a/w2294 ), .B(\SUBBYTES[6].a/w2301 ), .Z(
        \SUBBYTES[6].a/w2286 ) );
  IV U4986 ( .A(n1955), .Z(\SUBBYTES[6].a/w228 ) );
  NAND U4987 ( .A(\SUBBYTES[6].a/w207 ), .B(\SUBBYTES[6].a/w222 ), .Z(n1955)
         );
  AND U4988 ( .A(\SUBBYTES[6].a/w2234 ), .B(\SUBBYTES[6].a/w2230 ), .Z(
        \SUBBYTES[6].a/w2271 ) );
  AND U4989 ( .A(\SUBBYTES[6].a/w2235 ), .B(\SUBBYTES[6].a/w2231 ), .Z(
        \SUBBYTES[6].a/w2269 ) );
  ANDN U4990 ( .A(\SUBBYTES[6].a/w2361 ), .B(n1969), .Z(\SUBBYTES[6].a/w2268 )
         );
  XNOR U4991 ( .A(\w1[6][41] ), .B(\w1[6][47] ), .Z(n1969) );
  XOR U4992 ( .A(\w0[6][41] ), .B(g_input[809]), .Z(\w1[6][41] ) );
  AND U4993 ( .A(\w1[6][40] ), .B(\SUBBYTES[6].a/w2236 ), .Z(
        \SUBBYTES[6].a/w2264 ) );
  XOR U4994 ( .A(\w0[6][40] ), .B(g_input[808]), .Z(\w1[6][40] ) );
  AND U4995 ( .A(\SUBBYTES[6].a/w2237 ), .B(\SUBBYTES[6].a/w2233 ), .Z(
        \SUBBYTES[6].a/w2262 ) );
  AND U4996 ( .A(\SUBBYTES[6].a/w2322 ), .B(\SUBBYTES[6].a/w2354 ), .Z(
        \SUBBYTES[6].a/w2261 ) );
  ANDN U4997 ( .A(\SUBBYTES[6].a/w2343 ), .B(n1973), .Z(\SUBBYTES[6].a/w2256 )
         );
  XNOR U4998 ( .A(\w1[6][44] ), .B(\w1[6][47] ), .Z(n1973) );
  ANDN U4999 ( .A(\SUBBYTES[6].a/w2344 ), .B(n1974), .Z(\SUBBYTES[6].a/w2254 )
         );
  XNOR U5000 ( .A(\w1[6][42] ), .B(\w1[6][47] ), .Z(n1974) );
  XOR U5001 ( .A(\w0[6][47] ), .B(g_input[815]), .Z(\w1[6][47] ) );
  IV U5002 ( .A(n1976), .Z(\w1[6][42] ) );
  ANDN U5003 ( .A(\SUBBYTES[6].a/w2346 ), .B(n1975), .Z(\SUBBYTES[6].a/w2253 )
         );
  XOR U5004 ( .A(n1976), .B(\w1[6][44] ), .Z(n1975) );
  XOR U5005 ( .A(\w0[6][44] ), .B(g_input[812]), .Z(\w1[6][44] ) );
  XNOR U5006 ( .A(\w0[6][42] ), .B(g_input[810]), .Z(n1976) );
  AND U5007 ( .A(\SUBBYTES[6].a/w224 ), .B(\SUBBYTES[6].a/w230 ), .Z(
        \SUBBYTES[6].a/w225 ) );
  AND U5008 ( .A(\SUBBYTES[6].a/w209 ), .B(\SUBBYTES[6].a/w207 ), .Z(
        \SUBBYTES[6].a/w219 ) );
  AND U5009 ( .A(\SUBBYTES[6].a/w210 ), .B(\SUBBYTES[6].a/w208 ), .Z(
        \SUBBYTES[6].a/w217 ) );
  AND U5010 ( .A(\SUBBYTES[6].a/w224 ), .B(\SUBBYTES[6].a/w231 ), .Z(
        \SUBBYTES[6].a/w216 ) );
  AND U5011 ( .A(n1977), .B(\SUBBYTES[6].a/w2023 ), .Z(\SUBBYTES[6].a/w2158 )
         );
  AND U5012 ( .A(n1978), .B(\SUBBYTES[6].a/w2024 ), .Z(\SUBBYTES[6].a/w2156 )
         );
  AND U5013 ( .A(\SUBBYTES[6].a/w2154 ), .B(n1979), .Z(\SUBBYTES[6].a/w2155 )
         );
  ANDN U5014 ( .A(\w1[6][48] ), .B(n1980), .Z(\SUBBYTES[6].a/w2151 ) );
  AND U5015 ( .A(n1981), .B(\SUBBYTES[6].a/w2026 ), .Z(\SUBBYTES[6].a/w2149 )
         );
  AND U5016 ( .A(\SUBBYTES[6].a/w2147 ), .B(n1982), .Z(\SUBBYTES[6].a/w2148 )
         );
  XOR U5017 ( .A(\SUBBYTES[6].a/w2091 ), .B(n12250), .Z(n1982) );
  AND U5018 ( .A(\SUBBYTES[6].a/w2134 ), .B(\SUBBYTES[6].a/w2136 ), .Z(
        \SUBBYTES[6].a/w2143 ) );
  AND U5019 ( .A(\SUBBYTES[6].a/w2135 ), .B(\SUBBYTES[6].a/w2137 ), .Z(
        \SUBBYTES[6].a/w2141 ) );
  AND U5020 ( .A(\SUBBYTES[6].a/w2138 ), .B(\SUBBYTES[6].a/w2139 ), .Z(
        \SUBBYTES[6].a/w2140 ) );
  AND U5021 ( .A(\SUBBYTES[6].a/w2027 ), .B(n1977), .Z(\SUBBYTES[6].a/w2126 )
         );
  XOR U5022 ( .A(\SUBBYTES[6].a/w2095 ), .B(n1046), .Z(n1977) );
  AND U5023 ( .A(\SUBBYTES[6].a/w2028 ), .B(n1978), .Z(\SUBBYTES[6].a/w2124 )
         );
  XOR U5024 ( .A(n12251), .B(\SUBBYTES[6].a/w2095 ), .Z(n1978) );
  ANDN U5025 ( .A(n1979), .B(n1983), .Z(\SUBBYTES[6].a/w2123 ) );
  XOR U5026 ( .A(n1046), .B(n12251), .Z(n1979) );
  ANDN U5027 ( .A(\SUBBYTES[6].a/w2029 ), .B(n1980), .Z(\SUBBYTES[6].a/w2119 )
         );
  XNOR U5028 ( .A(\SUBBYTES[6].a/w2088 ), .B(\SUBBYTES[6].a/w2091 ), .Z(n1980)
         );
  AND U5029 ( .A(\SUBBYTES[6].a/w2030 ), .B(n1981), .Z(\SUBBYTES[6].a/w2117 )
         );
  XNOR U5030 ( .A(n1984), .B(\SUBBYTES[6].a/w2088 ), .Z(n1981) );
  AND U5031 ( .A(\SUBBYTES[6].a/w2115 ), .B(n1985), .Z(\SUBBYTES[6].a/w2116 )
         );
  XOR U5032 ( .A(n1986), .B(n1984), .Z(n1985) );
  IV U5033 ( .A(n12250), .Z(n1984) );
  ANDN U5034 ( .A(\SUBBYTES[6].a/w2134 ), .B(n1987), .Z(\SUBBYTES[6].a/w2111 )
         );
  ANDN U5035 ( .A(\SUBBYTES[6].a/w2135 ), .B(n1988), .Z(\SUBBYTES[6].a/w2109 )
         );
  ANDN U5036 ( .A(\SUBBYTES[6].a/w2138 ), .B(n1989), .Z(\SUBBYTES[6].a/w2108 )
         );
  AND U5037 ( .A(\SUBBYTES[6].a/w2094 ), .B(\SUBBYTES[6].a/w2093 ), .Z(
        \SUBBYTES[6].a/w2095 ) );
  IV U5038 ( .A(n1986), .Z(\SUBBYTES[6].a/w2091 ) );
  NAND U5039 ( .A(\SUBBYTES[6].a/w2070 ), .B(\SUBBYTES[6].a/w2085 ), .Z(n1986)
         );
  AND U5040 ( .A(\SUBBYTES[6].a/w2087 ), .B(\SUBBYTES[6].a/w2093 ), .Z(
        \SUBBYTES[6].a/w2088 ) );
  AND U5041 ( .A(\SUBBYTES[6].a/w2072 ), .B(\SUBBYTES[6].a/w2070 ), .Z(
        \SUBBYTES[6].a/w2082 ) );
  AND U5042 ( .A(\SUBBYTES[6].a/w2073 ), .B(\SUBBYTES[6].a/w2071 ), .Z(
        \SUBBYTES[6].a/w2080 ) );
  AND U5043 ( .A(\SUBBYTES[6].a/w2087 ), .B(\SUBBYTES[6].a/w2094 ), .Z(
        \SUBBYTES[6].a/w2079 ) );
  AND U5044 ( .A(\SUBBYTES[6].a/w2027 ), .B(\SUBBYTES[6].a/w2023 ), .Z(
        \SUBBYTES[6].a/w2064 ) );
  AND U5045 ( .A(\SUBBYTES[6].a/w2028 ), .B(\SUBBYTES[6].a/w2024 ), .Z(
        \SUBBYTES[6].a/w2062 ) );
  ANDN U5046 ( .A(\SUBBYTES[6].a/w2154 ), .B(n1983), .Z(\SUBBYTES[6].a/w2061 )
         );
  XNOR U5047 ( .A(\w1[6][49] ), .B(\w1[6][55] ), .Z(n1983) );
  XOR U5048 ( .A(\w0[6][49] ), .B(g_input[817]), .Z(\w1[6][49] ) );
  AND U5049 ( .A(\w1[6][48] ), .B(\SUBBYTES[6].a/w2029 ), .Z(
        \SUBBYTES[6].a/w2057 ) );
  XOR U5050 ( .A(\w0[6][48] ), .B(g_input[816]), .Z(\w1[6][48] ) );
  AND U5051 ( .A(\SUBBYTES[6].a/w2030 ), .B(\SUBBYTES[6].a/w2026 ), .Z(
        \SUBBYTES[6].a/w2055 ) );
  AND U5052 ( .A(\SUBBYTES[6].a/w2115 ), .B(\SUBBYTES[6].a/w2147 ), .Z(
        \SUBBYTES[6].a/w2054 ) );
  ANDN U5053 ( .A(\SUBBYTES[6].a/w2136 ), .B(n1987), .Z(\SUBBYTES[6].a/w2049 )
         );
  XNOR U5054 ( .A(\w1[6][52] ), .B(\w1[6][55] ), .Z(n1987) );
  ANDN U5055 ( .A(\SUBBYTES[6].a/w2137 ), .B(n1988), .Z(\SUBBYTES[6].a/w2047 )
         );
  XNOR U5056 ( .A(\w1[6][50] ), .B(\w1[6][55] ), .Z(n1988) );
  XOR U5057 ( .A(\w0[6][55] ), .B(g_input[823]), .Z(\w1[6][55] ) );
  IV U5058 ( .A(n1990), .Z(\w1[6][50] ) );
  ANDN U5059 ( .A(\SUBBYTES[6].a/w2139 ), .B(n1989), .Z(\SUBBYTES[6].a/w2046 )
         );
  XOR U5060 ( .A(n1990), .B(\w1[6][52] ), .Z(n1989) );
  XOR U5061 ( .A(\w0[6][52] ), .B(g_input[820]), .Z(\w1[6][52] ) );
  XNOR U5062 ( .A(\w0[6][50] ), .B(g_input[818]), .Z(n1990) );
  AND U5063 ( .A(\SUBBYTES[6].a/w164 ), .B(\SUBBYTES[6].a/w160 ), .Z(
        \SUBBYTES[6].a/w201 ) );
  AND U5064 ( .A(\SUBBYTES[6].a/w165 ), .B(\SUBBYTES[6].a/w161 ), .Z(
        \SUBBYTES[6].a/w199 ) );
  ANDN U5065 ( .A(\SUBBYTES[6].a/w291 ), .B(n1942), .Z(\SUBBYTES[6].a/w198 )
         );
  XNOR U5066 ( .A(\w1[6][121] ), .B(\w1[6][127] ), .Z(n1942) );
  XOR U5067 ( .A(\w0[6][121] ), .B(g_input[889]), .Z(\w1[6][121] ) );
  AND U5068 ( .A(n1991), .B(\SUBBYTES[6].a/w1816 ), .Z(\SUBBYTES[6].a/w1951 )
         );
  AND U5069 ( .A(n1992), .B(\SUBBYTES[6].a/w1817 ), .Z(\SUBBYTES[6].a/w1949 )
         );
  AND U5070 ( .A(\SUBBYTES[6].a/w1947 ), .B(n1993), .Z(\SUBBYTES[6].a/w1948 )
         );
  ANDN U5071 ( .A(\w1[6][56] ), .B(n1994), .Z(\SUBBYTES[6].a/w1944 ) );
  AND U5072 ( .A(n1995), .B(\SUBBYTES[6].a/w1819 ), .Z(\SUBBYTES[6].a/w1942 )
         );
  AND U5073 ( .A(\SUBBYTES[6].a/w1940 ), .B(n1996), .Z(\SUBBYTES[6].a/w1941 )
         );
  XOR U5074 ( .A(\SUBBYTES[6].a/w1884 ), .B(n12248), .Z(n1996) );
  AND U5075 ( .A(\w1[6][120] ), .B(\SUBBYTES[6].a/w166 ), .Z(
        \SUBBYTES[6].a/w194 ) );
  XOR U5076 ( .A(\w0[6][120] ), .B(g_input[888]), .Z(\w1[6][120] ) );
  AND U5077 ( .A(\SUBBYTES[6].a/w1927 ), .B(\SUBBYTES[6].a/w1929 ), .Z(
        \SUBBYTES[6].a/w1936 ) );
  AND U5078 ( .A(\SUBBYTES[6].a/w1928 ), .B(\SUBBYTES[6].a/w1930 ), .Z(
        \SUBBYTES[6].a/w1934 ) );
  AND U5079 ( .A(\SUBBYTES[6].a/w1931 ), .B(\SUBBYTES[6].a/w1932 ), .Z(
        \SUBBYTES[6].a/w1933 ) );
  AND U5080 ( .A(\SUBBYTES[6].a/w167 ), .B(\SUBBYTES[6].a/w163 ), .Z(
        \SUBBYTES[6].a/w192 ) );
  AND U5081 ( .A(\SUBBYTES[6].a/w1820 ), .B(n1991), .Z(\SUBBYTES[6].a/w1919 )
         );
  XOR U5082 ( .A(\SUBBYTES[6].a/w1888 ), .B(n1045), .Z(n1991) );
  AND U5083 ( .A(\SUBBYTES[6].a/w1821 ), .B(n1992), .Z(\SUBBYTES[6].a/w1917 )
         );
  XOR U5084 ( .A(n12249), .B(\SUBBYTES[6].a/w1888 ), .Z(n1992) );
  ANDN U5085 ( .A(n1993), .B(n1997), .Z(\SUBBYTES[6].a/w1916 ) );
  XOR U5086 ( .A(n1045), .B(n12249), .Z(n1993) );
  ANDN U5087 ( .A(\SUBBYTES[6].a/w1822 ), .B(n1994), .Z(\SUBBYTES[6].a/w1912 )
         );
  XNOR U5088 ( .A(\SUBBYTES[6].a/w1881 ), .B(\SUBBYTES[6].a/w1884 ), .Z(n1994)
         );
  AND U5089 ( .A(\SUBBYTES[6].a/w1823 ), .B(n1995), .Z(\SUBBYTES[6].a/w1910 )
         );
  XNOR U5090 ( .A(n1998), .B(\SUBBYTES[6].a/w1881 ), .Z(n1995) );
  AND U5091 ( .A(\SUBBYTES[6].a/w252 ), .B(\SUBBYTES[6].a/w284 ), .Z(
        \SUBBYTES[6].a/w191 ) );
  AND U5092 ( .A(\SUBBYTES[6].a/w1908 ), .B(n1999), .Z(\SUBBYTES[6].a/w1909 )
         );
  XOR U5093 ( .A(n2000), .B(n1998), .Z(n1999) );
  IV U5094 ( .A(n12248), .Z(n1998) );
  ANDN U5095 ( .A(\SUBBYTES[6].a/w1927 ), .B(n2001), .Z(\SUBBYTES[6].a/w1904 )
         );
  ANDN U5096 ( .A(\SUBBYTES[6].a/w1928 ), .B(n2002), .Z(\SUBBYTES[6].a/w1902 )
         );
  ANDN U5097 ( .A(\SUBBYTES[6].a/w1931 ), .B(n2003), .Z(\SUBBYTES[6].a/w1901 )
         );
  AND U5098 ( .A(\SUBBYTES[6].a/w1887 ), .B(\SUBBYTES[6].a/w1886 ), .Z(
        \SUBBYTES[6].a/w1888 ) );
  IV U5099 ( .A(n2000), .Z(\SUBBYTES[6].a/w1884 ) );
  NAND U5100 ( .A(\SUBBYTES[6].a/w1863 ), .B(\SUBBYTES[6].a/w1878 ), .Z(n2000)
         );
  AND U5101 ( .A(\SUBBYTES[6].a/w1880 ), .B(\SUBBYTES[6].a/w1886 ), .Z(
        \SUBBYTES[6].a/w1881 ) );
  AND U5102 ( .A(\SUBBYTES[6].a/w1865 ), .B(\SUBBYTES[6].a/w1863 ), .Z(
        \SUBBYTES[6].a/w1875 ) );
  AND U5103 ( .A(\SUBBYTES[6].a/w1866 ), .B(\SUBBYTES[6].a/w1864 ), .Z(
        \SUBBYTES[6].a/w1873 ) );
  AND U5104 ( .A(\SUBBYTES[6].a/w1880 ), .B(\SUBBYTES[6].a/w1887 ), .Z(
        \SUBBYTES[6].a/w1872 ) );
  ANDN U5105 ( .A(\SUBBYTES[6].a/w273 ), .B(n1959), .Z(\SUBBYTES[6].a/w186 )
         );
  XNOR U5106 ( .A(\w1[6][124] ), .B(\w1[6][127] ), .Z(n1959) );
  AND U5107 ( .A(\SUBBYTES[6].a/w1820 ), .B(\SUBBYTES[6].a/w1816 ), .Z(
        \SUBBYTES[6].a/w1857 ) );
  AND U5108 ( .A(\SUBBYTES[6].a/w1821 ), .B(\SUBBYTES[6].a/w1817 ), .Z(
        \SUBBYTES[6].a/w1855 ) );
  ANDN U5109 ( .A(\SUBBYTES[6].a/w1947 ), .B(n1997), .Z(\SUBBYTES[6].a/w1854 )
         );
  XNOR U5110 ( .A(\w1[6][57] ), .B(\w1[6][63] ), .Z(n1997) );
  XOR U5111 ( .A(\w0[6][57] ), .B(g_input[825]), .Z(\w1[6][57] ) );
  AND U5112 ( .A(\w1[6][56] ), .B(\SUBBYTES[6].a/w1822 ), .Z(
        \SUBBYTES[6].a/w1850 ) );
  XOR U5113 ( .A(\w0[6][56] ), .B(g_input[824]), .Z(\w1[6][56] ) );
  AND U5114 ( .A(\SUBBYTES[6].a/w1823 ), .B(\SUBBYTES[6].a/w1819 ), .Z(
        \SUBBYTES[6].a/w1848 ) );
  AND U5115 ( .A(\SUBBYTES[6].a/w1908 ), .B(\SUBBYTES[6].a/w1940 ), .Z(
        \SUBBYTES[6].a/w1847 ) );
  ANDN U5116 ( .A(\SUBBYTES[6].a/w1929 ), .B(n2001), .Z(\SUBBYTES[6].a/w1842 )
         );
  XNOR U5117 ( .A(\w1[6][60] ), .B(\w1[6][63] ), .Z(n2001) );
  ANDN U5118 ( .A(\SUBBYTES[6].a/w1930 ), .B(n2002), .Z(\SUBBYTES[6].a/w1840 )
         );
  XNOR U5119 ( .A(\w1[6][58] ), .B(\w1[6][63] ), .Z(n2002) );
  XOR U5120 ( .A(\w0[6][63] ), .B(g_input[831]), .Z(\w1[6][63] ) );
  IV U5121 ( .A(n2004), .Z(\w1[6][58] ) );
  ANDN U5122 ( .A(\SUBBYTES[6].a/w274 ), .B(n1961), .Z(\SUBBYTES[6].a/w184 )
         );
  XNOR U5123 ( .A(\w1[6][122] ), .B(\w1[6][127] ), .Z(n1961) );
  XOR U5124 ( .A(\w0[6][127] ), .B(g_input[895]), .Z(\w1[6][127] ) );
  IV U5125 ( .A(n2005), .Z(\w1[6][122] ) );
  ANDN U5126 ( .A(\SUBBYTES[6].a/w1932 ), .B(n2003), .Z(\SUBBYTES[6].a/w1839 )
         );
  XOR U5127 ( .A(n2004), .B(\w1[6][60] ), .Z(n2003) );
  XOR U5128 ( .A(\w0[6][60] ), .B(g_input[828]), .Z(\w1[6][60] ) );
  XNOR U5129 ( .A(\w0[6][58] ), .B(g_input[826]), .Z(n2004) );
  ANDN U5130 ( .A(\SUBBYTES[6].a/w276 ), .B(n1962), .Z(\SUBBYTES[6].a/w183 )
         );
  XOR U5131 ( .A(n2005), .B(\w1[6][124] ), .Z(n1962) );
  XOR U5132 ( .A(\w0[6][124] ), .B(g_input[892]), .Z(\w1[6][124] ) );
  XNOR U5133 ( .A(\w0[6][122] ), .B(g_input[890]), .Z(n2005) );
  AND U5134 ( .A(n2006), .B(\SUBBYTES[6].a/w1609 ), .Z(\SUBBYTES[6].a/w1744 )
         );
  AND U5135 ( .A(n2007), .B(\SUBBYTES[6].a/w1610 ), .Z(\SUBBYTES[6].a/w1742 )
         );
  AND U5136 ( .A(\SUBBYTES[6].a/w1740 ), .B(n2008), .Z(\SUBBYTES[6].a/w1741 )
         );
  ANDN U5137 ( .A(\w1[6][64] ), .B(n2009), .Z(\SUBBYTES[6].a/w1737 ) );
  AND U5138 ( .A(n2010), .B(\SUBBYTES[6].a/w1612 ), .Z(\SUBBYTES[6].a/w1735 )
         );
  AND U5139 ( .A(\SUBBYTES[6].a/w1733 ), .B(n2011), .Z(\SUBBYTES[6].a/w1734 )
         );
  XOR U5140 ( .A(\SUBBYTES[6].a/w1677 ), .B(n12246), .Z(n2011) );
  AND U5141 ( .A(\SUBBYTES[6].a/w1720 ), .B(\SUBBYTES[6].a/w1722 ), .Z(
        \SUBBYTES[6].a/w1729 ) );
  AND U5142 ( .A(\SUBBYTES[6].a/w1721 ), .B(\SUBBYTES[6].a/w1723 ), .Z(
        \SUBBYTES[6].a/w1727 ) );
  AND U5143 ( .A(\SUBBYTES[6].a/w1724 ), .B(\SUBBYTES[6].a/w1725 ), .Z(
        \SUBBYTES[6].a/w1726 ) );
  AND U5144 ( .A(\SUBBYTES[6].a/w1613 ), .B(n2006), .Z(\SUBBYTES[6].a/w1712 )
         );
  XOR U5145 ( .A(\SUBBYTES[6].a/w1681 ), .B(n1044), .Z(n2006) );
  AND U5146 ( .A(\SUBBYTES[6].a/w1614 ), .B(n2007), .Z(\SUBBYTES[6].a/w1710 )
         );
  XOR U5147 ( .A(n12247), .B(\SUBBYTES[6].a/w1681 ), .Z(n2007) );
  ANDN U5148 ( .A(n2008), .B(n2012), .Z(\SUBBYTES[6].a/w1709 ) );
  XOR U5149 ( .A(n1044), .B(n12247), .Z(n2008) );
  ANDN U5150 ( .A(\SUBBYTES[6].a/w1615 ), .B(n2009), .Z(\SUBBYTES[6].a/w1705 )
         );
  XNOR U5151 ( .A(\SUBBYTES[6].a/w1674 ), .B(\SUBBYTES[6].a/w1677 ), .Z(n2009)
         );
  AND U5152 ( .A(\SUBBYTES[6].a/w1616 ), .B(n2010), .Z(\SUBBYTES[6].a/w1703 )
         );
  XNOR U5153 ( .A(n2013), .B(\SUBBYTES[6].a/w1674 ), .Z(n2010) );
  AND U5154 ( .A(\SUBBYTES[6].a/w1701 ), .B(n2014), .Z(\SUBBYTES[6].a/w1702 )
         );
  XOR U5155 ( .A(n2015), .B(n2013), .Z(n2014) );
  IV U5156 ( .A(n12246), .Z(n2013) );
  ANDN U5157 ( .A(\SUBBYTES[6].a/w1720 ), .B(n2016), .Z(\SUBBYTES[6].a/w1697 )
         );
  ANDN U5158 ( .A(\SUBBYTES[6].a/w1721 ), .B(n2017), .Z(\SUBBYTES[6].a/w1695 )
         );
  ANDN U5159 ( .A(\SUBBYTES[6].a/w1724 ), .B(n2018), .Z(\SUBBYTES[6].a/w1694 )
         );
  AND U5160 ( .A(\SUBBYTES[6].a/w1680 ), .B(\SUBBYTES[6].a/w1679 ), .Z(
        \SUBBYTES[6].a/w1681 ) );
  IV U5161 ( .A(n2015), .Z(\SUBBYTES[6].a/w1677 ) );
  NAND U5162 ( .A(\SUBBYTES[6].a/w1656 ), .B(\SUBBYTES[6].a/w1671 ), .Z(n2015)
         );
  AND U5163 ( .A(\SUBBYTES[6].a/w1673 ), .B(\SUBBYTES[6].a/w1679 ), .Z(
        \SUBBYTES[6].a/w1674 ) );
  AND U5164 ( .A(\SUBBYTES[6].a/w1658 ), .B(\SUBBYTES[6].a/w1656 ), .Z(
        \SUBBYTES[6].a/w1668 ) );
  AND U5165 ( .A(\SUBBYTES[6].a/w1659 ), .B(\SUBBYTES[6].a/w1657 ), .Z(
        \SUBBYTES[6].a/w1666 ) );
  AND U5166 ( .A(\SUBBYTES[6].a/w1673 ), .B(\SUBBYTES[6].a/w1680 ), .Z(
        \SUBBYTES[6].a/w1665 ) );
  AND U5167 ( .A(\SUBBYTES[6].a/w1613 ), .B(\SUBBYTES[6].a/w1609 ), .Z(
        \SUBBYTES[6].a/w1650 ) );
  AND U5168 ( .A(\SUBBYTES[6].a/w1614 ), .B(\SUBBYTES[6].a/w1610 ), .Z(
        \SUBBYTES[6].a/w1648 ) );
  ANDN U5169 ( .A(\SUBBYTES[6].a/w1740 ), .B(n2012), .Z(\SUBBYTES[6].a/w1647 )
         );
  XNOR U5170 ( .A(\w1[6][65] ), .B(\w1[6][71] ), .Z(n2012) );
  XOR U5171 ( .A(\w0[6][65] ), .B(g_input[833]), .Z(\w1[6][65] ) );
  AND U5172 ( .A(\w1[6][64] ), .B(\SUBBYTES[6].a/w1615 ), .Z(
        \SUBBYTES[6].a/w1643 ) );
  XOR U5173 ( .A(\w0[6][64] ), .B(g_input[832]), .Z(\w1[6][64] ) );
  AND U5174 ( .A(\SUBBYTES[6].a/w1616 ), .B(\SUBBYTES[6].a/w1612 ), .Z(
        \SUBBYTES[6].a/w1641 ) );
  AND U5175 ( .A(\SUBBYTES[6].a/w1701 ), .B(\SUBBYTES[6].a/w1733 ), .Z(
        \SUBBYTES[6].a/w1640 ) );
  ANDN U5176 ( .A(\SUBBYTES[6].a/w1722 ), .B(n2016), .Z(\SUBBYTES[6].a/w1635 )
         );
  XNOR U5177 ( .A(\w1[6][68] ), .B(\w1[6][71] ), .Z(n2016) );
  ANDN U5178 ( .A(\SUBBYTES[6].a/w1723 ), .B(n2017), .Z(\SUBBYTES[6].a/w1633 )
         );
  XNOR U5179 ( .A(\w1[6][66] ), .B(\w1[6][71] ), .Z(n2017) );
  XOR U5180 ( .A(\w0[6][71] ), .B(g_input[839]), .Z(\w1[6][71] ) );
  IV U5181 ( .A(n2019), .Z(\w1[6][66] ) );
  ANDN U5182 ( .A(\SUBBYTES[6].a/w1725 ), .B(n2018), .Z(\SUBBYTES[6].a/w1632 )
         );
  XOR U5183 ( .A(n2019), .B(\w1[6][68] ), .Z(n2018) );
  XOR U5184 ( .A(\w0[6][68] ), .B(g_input[836]), .Z(\w1[6][68] ) );
  XNOR U5185 ( .A(\w0[6][66] ), .B(g_input[834]), .Z(n2019) );
  AND U5186 ( .A(n2020), .B(\SUBBYTES[6].a/w1402 ), .Z(\SUBBYTES[6].a/w1537 )
         );
  AND U5187 ( .A(n2021), .B(\SUBBYTES[6].a/w1403 ), .Z(\SUBBYTES[6].a/w1535 )
         );
  AND U5188 ( .A(\SUBBYTES[6].a/w1533 ), .B(n2022), .Z(\SUBBYTES[6].a/w1534 )
         );
  ANDN U5189 ( .A(\w1[6][72] ), .B(n2023), .Z(\SUBBYTES[6].a/w1530 ) );
  AND U5190 ( .A(n2024), .B(\SUBBYTES[6].a/w1405 ), .Z(\SUBBYTES[6].a/w1528 )
         );
  AND U5191 ( .A(\SUBBYTES[6].a/w1526 ), .B(n2025), .Z(\SUBBYTES[6].a/w1527 )
         );
  XOR U5192 ( .A(\SUBBYTES[6].a/w1470 ), .B(n12244), .Z(n2025) );
  AND U5193 ( .A(\SUBBYTES[6].a/w1513 ), .B(\SUBBYTES[6].a/w1515 ), .Z(
        \SUBBYTES[6].a/w1522 ) );
  AND U5194 ( .A(\SUBBYTES[6].a/w1514 ), .B(\SUBBYTES[6].a/w1516 ), .Z(
        \SUBBYTES[6].a/w1520 ) );
  AND U5195 ( .A(\SUBBYTES[6].a/w1517 ), .B(\SUBBYTES[6].a/w1518 ), .Z(
        \SUBBYTES[6].a/w1519 ) );
  AND U5196 ( .A(\SUBBYTES[6].a/w1406 ), .B(n2020), .Z(\SUBBYTES[6].a/w1505 )
         );
  XOR U5197 ( .A(\SUBBYTES[6].a/w1474 ), .B(n1043), .Z(n2020) );
  AND U5198 ( .A(\SUBBYTES[6].a/w1407 ), .B(n2021), .Z(\SUBBYTES[6].a/w1503 )
         );
  XOR U5199 ( .A(n12245), .B(\SUBBYTES[6].a/w1474 ), .Z(n2021) );
  ANDN U5200 ( .A(n2022), .B(n2026), .Z(\SUBBYTES[6].a/w1502 ) );
  XOR U5201 ( .A(n1043), .B(n12245), .Z(n2022) );
  ANDN U5202 ( .A(\SUBBYTES[6].a/w1408 ), .B(n2023), .Z(\SUBBYTES[6].a/w1498 )
         );
  XNOR U5203 ( .A(\SUBBYTES[6].a/w1467 ), .B(\SUBBYTES[6].a/w1470 ), .Z(n2023)
         );
  AND U5204 ( .A(\SUBBYTES[6].a/w1409 ), .B(n2024), .Z(\SUBBYTES[6].a/w1496 )
         );
  XNOR U5205 ( .A(n2027), .B(\SUBBYTES[6].a/w1467 ), .Z(n2024) );
  AND U5206 ( .A(\SUBBYTES[6].a/w1494 ), .B(n2028), .Z(\SUBBYTES[6].a/w1495 )
         );
  XOR U5207 ( .A(n2029), .B(n2027), .Z(n2028) );
  IV U5208 ( .A(n12244), .Z(n2027) );
  ANDN U5209 ( .A(\SUBBYTES[6].a/w1513 ), .B(n2030), .Z(\SUBBYTES[6].a/w1490 )
         );
  ANDN U5210 ( .A(\SUBBYTES[6].a/w1514 ), .B(n2031), .Z(\SUBBYTES[6].a/w1488 )
         );
  ANDN U5211 ( .A(\SUBBYTES[6].a/w1517 ), .B(n2032), .Z(\SUBBYTES[6].a/w1487 )
         );
  AND U5212 ( .A(\SUBBYTES[6].a/w1473 ), .B(\SUBBYTES[6].a/w1472 ), .Z(
        \SUBBYTES[6].a/w1474 ) );
  IV U5213 ( .A(n2029), .Z(\SUBBYTES[6].a/w1470 ) );
  NAND U5214 ( .A(\SUBBYTES[6].a/w1449 ), .B(\SUBBYTES[6].a/w1464 ), .Z(n2029)
         );
  AND U5215 ( .A(\SUBBYTES[6].a/w1466 ), .B(\SUBBYTES[6].a/w1472 ), .Z(
        \SUBBYTES[6].a/w1467 ) );
  AND U5216 ( .A(\SUBBYTES[6].a/w1451 ), .B(\SUBBYTES[6].a/w1449 ), .Z(
        \SUBBYTES[6].a/w1461 ) );
  AND U5217 ( .A(\SUBBYTES[6].a/w1452 ), .B(\SUBBYTES[6].a/w1450 ), .Z(
        \SUBBYTES[6].a/w1459 ) );
  AND U5218 ( .A(\SUBBYTES[6].a/w1466 ), .B(\SUBBYTES[6].a/w1473 ), .Z(
        \SUBBYTES[6].a/w1458 ) );
  AND U5219 ( .A(\SUBBYTES[6].a/w1406 ), .B(\SUBBYTES[6].a/w1402 ), .Z(
        \SUBBYTES[6].a/w1443 ) );
  AND U5220 ( .A(\SUBBYTES[6].a/w1407 ), .B(\SUBBYTES[6].a/w1403 ), .Z(
        \SUBBYTES[6].a/w1441 ) );
  ANDN U5221 ( .A(\SUBBYTES[6].a/w1533 ), .B(n2026), .Z(\SUBBYTES[6].a/w1440 )
         );
  XNOR U5222 ( .A(\w1[6][73] ), .B(\w1[6][79] ), .Z(n2026) );
  XOR U5223 ( .A(\w0[6][73] ), .B(g_input[841]), .Z(\w1[6][73] ) );
  AND U5224 ( .A(\w1[6][72] ), .B(\SUBBYTES[6].a/w1408 ), .Z(
        \SUBBYTES[6].a/w1436 ) );
  XOR U5225 ( .A(\w0[6][72] ), .B(g_input[840]), .Z(\w1[6][72] ) );
  AND U5226 ( .A(\SUBBYTES[6].a/w1409 ), .B(\SUBBYTES[6].a/w1405 ), .Z(
        \SUBBYTES[6].a/w1434 ) );
  AND U5227 ( .A(\SUBBYTES[6].a/w1494 ), .B(\SUBBYTES[6].a/w1526 ), .Z(
        \SUBBYTES[6].a/w1433 ) );
  ANDN U5228 ( .A(\SUBBYTES[6].a/w1515 ), .B(n2030), .Z(\SUBBYTES[6].a/w1428 )
         );
  XNOR U5229 ( .A(\w1[6][76] ), .B(\w1[6][79] ), .Z(n2030) );
  ANDN U5230 ( .A(\SUBBYTES[6].a/w1516 ), .B(n2031), .Z(\SUBBYTES[6].a/w1426 )
         );
  XNOR U5231 ( .A(\w1[6][74] ), .B(\w1[6][79] ), .Z(n2031) );
  XOR U5232 ( .A(\w0[6][79] ), .B(g_input[847]), .Z(\w1[6][79] ) );
  IV U5233 ( .A(n2033), .Z(\w1[6][74] ) );
  ANDN U5234 ( .A(\SUBBYTES[6].a/w1518 ), .B(n2032), .Z(\SUBBYTES[6].a/w1425 )
         );
  XOR U5235 ( .A(n2033), .B(\w1[6][76] ), .Z(n2032) );
  XOR U5236 ( .A(\w0[6][76] ), .B(g_input[844]), .Z(\w1[6][76] ) );
  XNOR U5237 ( .A(\w0[6][74] ), .B(g_input[842]), .Z(n2033) );
  AND U5238 ( .A(n2034), .B(\SUBBYTES[6].a/w1195 ), .Z(\SUBBYTES[6].a/w1330 )
         );
  AND U5239 ( .A(n2035), .B(\SUBBYTES[6].a/w1196 ), .Z(\SUBBYTES[6].a/w1328 )
         );
  AND U5240 ( .A(\SUBBYTES[6].a/w1326 ), .B(n2036), .Z(\SUBBYTES[6].a/w1327 )
         );
  ANDN U5241 ( .A(\w1[6][80] ), .B(n2037), .Z(\SUBBYTES[6].a/w1323 ) );
  AND U5242 ( .A(n2038), .B(\SUBBYTES[6].a/w1198 ), .Z(\SUBBYTES[6].a/w1321 )
         );
  AND U5243 ( .A(\SUBBYTES[6].a/w1319 ), .B(n2039), .Z(\SUBBYTES[6].a/w1320 )
         );
  XOR U5244 ( .A(\SUBBYTES[6].a/w1263 ), .B(n12242), .Z(n2039) );
  AND U5245 ( .A(\SUBBYTES[6].a/w1306 ), .B(\SUBBYTES[6].a/w1308 ), .Z(
        \SUBBYTES[6].a/w1315 ) );
  AND U5246 ( .A(\SUBBYTES[6].a/w1307 ), .B(\SUBBYTES[6].a/w1309 ), .Z(
        \SUBBYTES[6].a/w1313 ) );
  AND U5247 ( .A(\SUBBYTES[6].a/w1310 ), .B(\SUBBYTES[6].a/w1311 ), .Z(
        \SUBBYTES[6].a/w1312 ) );
  AND U5248 ( .A(\SUBBYTES[6].a/w1199 ), .B(n2034), .Z(\SUBBYTES[6].a/w1298 )
         );
  XOR U5249 ( .A(\SUBBYTES[6].a/w1267 ), .B(n1042), .Z(n2034) );
  AND U5250 ( .A(\SUBBYTES[6].a/w1200 ), .B(n2035), .Z(\SUBBYTES[6].a/w1296 )
         );
  XOR U5251 ( .A(n12243), .B(\SUBBYTES[6].a/w1267 ), .Z(n2035) );
  ANDN U5252 ( .A(n2036), .B(n2040), .Z(\SUBBYTES[6].a/w1295 ) );
  XOR U5253 ( .A(n1042), .B(n12243), .Z(n2036) );
  ANDN U5254 ( .A(\SUBBYTES[6].a/w1201 ), .B(n2037), .Z(\SUBBYTES[6].a/w1291 )
         );
  XNOR U5255 ( .A(\SUBBYTES[6].a/w1260 ), .B(\SUBBYTES[6].a/w1263 ), .Z(n2037)
         );
  AND U5256 ( .A(\SUBBYTES[6].a/w1202 ), .B(n2038), .Z(\SUBBYTES[6].a/w1289 )
         );
  XNOR U5257 ( .A(n2041), .B(\SUBBYTES[6].a/w1260 ), .Z(n2038) );
  AND U5258 ( .A(\SUBBYTES[6].a/w1287 ), .B(n2042), .Z(\SUBBYTES[6].a/w1288 )
         );
  XOR U5259 ( .A(n2043), .B(n2041), .Z(n2042) );
  IV U5260 ( .A(n12242), .Z(n2041) );
  ANDN U5261 ( .A(\SUBBYTES[6].a/w1306 ), .B(n2044), .Z(\SUBBYTES[6].a/w1283 )
         );
  ANDN U5262 ( .A(\SUBBYTES[6].a/w1307 ), .B(n2045), .Z(\SUBBYTES[6].a/w1281 )
         );
  ANDN U5263 ( .A(\SUBBYTES[6].a/w1310 ), .B(n2046), .Z(\SUBBYTES[6].a/w1280 )
         );
  AND U5264 ( .A(\SUBBYTES[6].a/w1266 ), .B(\SUBBYTES[6].a/w1265 ), .Z(
        \SUBBYTES[6].a/w1267 ) );
  IV U5265 ( .A(n2043), .Z(\SUBBYTES[6].a/w1263 ) );
  NAND U5266 ( .A(\SUBBYTES[6].a/w1242 ), .B(\SUBBYTES[6].a/w1257 ), .Z(n2043)
         );
  AND U5267 ( .A(\SUBBYTES[6].a/w1259 ), .B(\SUBBYTES[6].a/w1265 ), .Z(
        \SUBBYTES[6].a/w1260 ) );
  AND U5268 ( .A(\SUBBYTES[6].a/w1244 ), .B(\SUBBYTES[6].a/w1242 ), .Z(
        \SUBBYTES[6].a/w1254 ) );
  AND U5269 ( .A(\SUBBYTES[6].a/w1245 ), .B(\SUBBYTES[6].a/w1243 ), .Z(
        \SUBBYTES[6].a/w1252 ) );
  AND U5270 ( .A(\SUBBYTES[6].a/w1259 ), .B(\SUBBYTES[6].a/w1266 ), .Z(
        \SUBBYTES[6].a/w1251 ) );
  AND U5271 ( .A(\SUBBYTES[6].a/w1199 ), .B(\SUBBYTES[6].a/w1195 ), .Z(
        \SUBBYTES[6].a/w1236 ) );
  AND U5272 ( .A(\SUBBYTES[6].a/w1200 ), .B(\SUBBYTES[6].a/w1196 ), .Z(
        \SUBBYTES[6].a/w1234 ) );
  ANDN U5273 ( .A(\SUBBYTES[6].a/w1326 ), .B(n2040), .Z(\SUBBYTES[6].a/w1233 )
         );
  XNOR U5274 ( .A(\w1[6][81] ), .B(\w1[6][87] ), .Z(n2040) );
  XOR U5275 ( .A(\w0[6][81] ), .B(g_input[849]), .Z(\w1[6][81] ) );
  AND U5276 ( .A(\w1[6][80] ), .B(\SUBBYTES[6].a/w1201 ), .Z(
        \SUBBYTES[6].a/w1229 ) );
  XOR U5277 ( .A(\w0[6][80] ), .B(g_input[848]), .Z(\w1[6][80] ) );
  AND U5278 ( .A(\SUBBYTES[6].a/w1202 ), .B(\SUBBYTES[6].a/w1198 ), .Z(
        \SUBBYTES[6].a/w1227 ) );
  AND U5279 ( .A(\SUBBYTES[6].a/w1287 ), .B(\SUBBYTES[6].a/w1319 ), .Z(
        \SUBBYTES[6].a/w1226 ) );
  ANDN U5280 ( .A(\SUBBYTES[6].a/w1308 ), .B(n2044), .Z(\SUBBYTES[6].a/w1221 )
         );
  XNOR U5281 ( .A(\w1[6][84] ), .B(\w1[6][87] ), .Z(n2044) );
  ANDN U5282 ( .A(\SUBBYTES[6].a/w1309 ), .B(n2045), .Z(\SUBBYTES[6].a/w1219 )
         );
  XNOR U5283 ( .A(\w1[6][82] ), .B(\w1[6][87] ), .Z(n2045) );
  XOR U5284 ( .A(\w0[6][87] ), .B(g_input[855]), .Z(\w1[6][87] ) );
  IV U5285 ( .A(n2047), .Z(\w1[6][82] ) );
  ANDN U5286 ( .A(\SUBBYTES[6].a/w1311 ), .B(n2046), .Z(\SUBBYTES[6].a/w1218 )
         );
  XOR U5287 ( .A(n2047), .B(\w1[6][84] ), .Z(n2046) );
  XOR U5288 ( .A(\w0[6][84] ), .B(g_input[852]), .Z(\w1[6][84] ) );
  XNOR U5289 ( .A(\w0[6][82] ), .B(g_input[850]), .Z(n2047) );
  AND U5290 ( .A(n2048), .B(\SUBBYTES[6].a/w988 ), .Z(\SUBBYTES[6].a/w1123 )
         );
  AND U5291 ( .A(n2049), .B(\SUBBYTES[6].a/w989 ), .Z(\SUBBYTES[6].a/w1121 )
         );
  AND U5292 ( .A(\SUBBYTES[6].a/w1119 ), .B(n2050), .Z(\SUBBYTES[6].a/w1120 )
         );
  ANDN U5293 ( .A(\w1[6][88] ), .B(n2051), .Z(\SUBBYTES[6].a/w1116 ) );
  AND U5294 ( .A(n2052), .B(\SUBBYTES[6].a/w991 ), .Z(\SUBBYTES[6].a/w1114 )
         );
  AND U5295 ( .A(\SUBBYTES[6].a/w1112 ), .B(n2053), .Z(\SUBBYTES[6].a/w1113 )
         );
  XOR U5296 ( .A(\SUBBYTES[6].a/w1056 ), .B(n12240), .Z(n2053) );
  AND U5297 ( .A(\SUBBYTES[6].a/w1099 ), .B(\SUBBYTES[6].a/w1101 ), .Z(
        \SUBBYTES[6].a/w1108 ) );
  AND U5298 ( .A(\SUBBYTES[6].a/w1100 ), .B(\SUBBYTES[6].a/w1102 ), .Z(
        \SUBBYTES[6].a/w1106 ) );
  AND U5299 ( .A(\SUBBYTES[6].a/w1103 ), .B(\SUBBYTES[6].a/w1104 ), .Z(
        \SUBBYTES[6].a/w1105 ) );
  AND U5300 ( .A(\SUBBYTES[6].a/w992 ), .B(n2048), .Z(\SUBBYTES[6].a/w1091 )
         );
  XOR U5301 ( .A(\SUBBYTES[6].a/w1060 ), .B(n1041), .Z(n2048) );
  AND U5302 ( .A(\SUBBYTES[6].a/w993 ), .B(n2049), .Z(\SUBBYTES[6].a/w1089 )
         );
  XOR U5303 ( .A(n12241), .B(\SUBBYTES[6].a/w1060 ), .Z(n2049) );
  ANDN U5304 ( .A(n2050), .B(n2054), .Z(\SUBBYTES[6].a/w1088 ) );
  XOR U5305 ( .A(n1041), .B(n12241), .Z(n2050) );
  ANDN U5306 ( .A(\SUBBYTES[6].a/w994 ), .B(n2051), .Z(\SUBBYTES[6].a/w1084 )
         );
  XNOR U5307 ( .A(\SUBBYTES[6].a/w1053 ), .B(\SUBBYTES[6].a/w1056 ), .Z(n2051)
         );
  AND U5308 ( .A(\SUBBYTES[6].a/w995 ), .B(n2052), .Z(\SUBBYTES[6].a/w1082 )
         );
  XNOR U5309 ( .A(n2055), .B(\SUBBYTES[6].a/w1053 ), .Z(n2052) );
  AND U5310 ( .A(\SUBBYTES[6].a/w1080 ), .B(n2056), .Z(\SUBBYTES[6].a/w1081 )
         );
  XOR U5311 ( .A(n2057), .B(n2055), .Z(n2056) );
  IV U5312 ( .A(n12240), .Z(n2055) );
  ANDN U5313 ( .A(\SUBBYTES[6].a/w1099 ), .B(n2058), .Z(\SUBBYTES[6].a/w1076 )
         );
  ANDN U5314 ( .A(\SUBBYTES[6].a/w1100 ), .B(n2059), .Z(\SUBBYTES[6].a/w1074 )
         );
  ANDN U5315 ( .A(\SUBBYTES[6].a/w1103 ), .B(n2060), .Z(\SUBBYTES[6].a/w1073 )
         );
  AND U5316 ( .A(\SUBBYTES[6].a/w1059 ), .B(\SUBBYTES[6].a/w1058 ), .Z(
        \SUBBYTES[6].a/w1060 ) );
  IV U5317 ( .A(n2057), .Z(\SUBBYTES[6].a/w1056 ) );
  NAND U5318 ( .A(\SUBBYTES[6].a/w1035 ), .B(\SUBBYTES[6].a/w1050 ), .Z(n2057)
         );
  AND U5319 ( .A(\SUBBYTES[6].a/w1052 ), .B(\SUBBYTES[6].a/w1058 ), .Z(
        \SUBBYTES[6].a/w1053 ) );
  AND U5320 ( .A(\SUBBYTES[6].a/w1037 ), .B(\SUBBYTES[6].a/w1035 ), .Z(
        \SUBBYTES[6].a/w1047 ) );
  AND U5321 ( .A(\SUBBYTES[6].a/w1038 ), .B(\SUBBYTES[6].a/w1036 ), .Z(
        \SUBBYTES[6].a/w1045 ) );
  AND U5322 ( .A(\SUBBYTES[6].a/w1052 ), .B(\SUBBYTES[6].a/w1059 ), .Z(
        \SUBBYTES[6].a/w1044 ) );
  AND U5323 ( .A(\SUBBYTES[6].a/w992 ), .B(\SUBBYTES[6].a/w988 ), .Z(
        \SUBBYTES[6].a/w1029 ) );
  AND U5324 ( .A(\SUBBYTES[6].a/w993 ), .B(\SUBBYTES[6].a/w989 ), .Z(
        \SUBBYTES[6].a/w1027 ) );
  ANDN U5325 ( .A(\SUBBYTES[6].a/w1119 ), .B(n2054), .Z(\SUBBYTES[6].a/w1026 )
         );
  XNOR U5326 ( .A(\w1[6][89] ), .B(\w1[6][95] ), .Z(n2054) );
  XOR U5327 ( .A(\w0[6][89] ), .B(g_input[857]), .Z(\w1[6][89] ) );
  AND U5328 ( .A(\w1[6][88] ), .B(\SUBBYTES[6].a/w994 ), .Z(
        \SUBBYTES[6].a/w1022 ) );
  XOR U5329 ( .A(\w0[6][88] ), .B(g_input[856]), .Z(\w1[6][88] ) );
  AND U5330 ( .A(\SUBBYTES[6].a/w995 ), .B(\SUBBYTES[6].a/w991 ), .Z(
        \SUBBYTES[6].a/w1020 ) );
  AND U5331 ( .A(\SUBBYTES[6].a/w1080 ), .B(\SUBBYTES[6].a/w1112 ), .Z(
        \SUBBYTES[6].a/w1019 ) );
  ANDN U5332 ( .A(\SUBBYTES[6].a/w1101 ), .B(n2058), .Z(\SUBBYTES[6].a/w1014 )
         );
  XNOR U5333 ( .A(\w1[6][92] ), .B(\w1[6][95] ), .Z(n2058) );
  ANDN U5334 ( .A(\SUBBYTES[6].a/w1102 ), .B(n2059), .Z(\SUBBYTES[6].a/w1012 )
         );
  XNOR U5335 ( .A(\w1[6][90] ), .B(\w1[6][95] ), .Z(n2059) );
  XOR U5336 ( .A(\w0[6][95] ), .B(g_input[863]), .Z(\w1[6][95] ) );
  IV U5337 ( .A(n2061), .Z(\w1[6][90] ) );
  ANDN U5338 ( .A(\SUBBYTES[6].a/w1104 ), .B(n2060), .Z(\SUBBYTES[6].a/w1011 )
         );
  XOR U5339 ( .A(n2061), .B(\w1[6][92] ), .Z(n2060) );
  XOR U5340 ( .A(\w0[6][92] ), .B(g_input[860]), .Z(\w1[6][92] ) );
  XNOR U5341 ( .A(\w0[6][90] ), .B(g_input[858]), .Z(n2061) );
  AND U5342 ( .A(\SUBBYTES[6].a/w2084 ), .B(\SUBBYTES[6].a/w2071 ), .Z(n12250)
         );
  AND U5343 ( .A(\SUBBYTES[6].a/w1877 ), .B(\SUBBYTES[6].a/w1866 ), .Z(n12249)
         );
  AND U5344 ( .A(\SUBBYTES[6].a/w221 ), .B(\SUBBYTES[6].a/w208 ), .Z(n12232)
         );
  AND U5345 ( .A(\SUBBYTES[6].a/w1877 ), .B(\SUBBYTES[6].a/w1864 ), .Z(n12248)
         );
  AND U5346 ( .A(\SUBBYTES[6].a/w1670 ), .B(\SUBBYTES[6].a/w1659 ), .Z(n12247)
         );
  AND U5347 ( .A(\SUBBYTES[6].a/w1670 ), .B(\SUBBYTES[6].a/w1657 ), .Z(n12246)
         );
  AND U5348 ( .A(\SUBBYTES[6].a/w1463 ), .B(\SUBBYTES[6].a/w1452 ), .Z(n12245)
         );
  AND U5349 ( .A(\SUBBYTES[6].a/w1463 ), .B(\SUBBYTES[6].a/w1450 ), .Z(n12244)
         );
  AND U5350 ( .A(\SUBBYTES[6].a/w1256 ), .B(\SUBBYTES[6].a/w1245 ), .Z(n12243)
         );
  AND U5351 ( .A(\SUBBYTES[6].a/w1256 ), .B(\SUBBYTES[6].a/w1243 ), .Z(n12242)
         );
  AND U5352 ( .A(\SUBBYTES[6].a/w1049 ), .B(\SUBBYTES[6].a/w1038 ), .Z(n12241)
         );
  AND U5353 ( .A(\SUBBYTES[6].a/w1049 ), .B(\SUBBYTES[6].a/w1036 ), .Z(n12240)
         );
  AND U5354 ( .A(\SUBBYTES[6].a/w842 ), .B(\SUBBYTES[6].a/w831 ), .Z(n12239)
         );
  AND U5355 ( .A(\SUBBYTES[6].a/w842 ), .B(\SUBBYTES[6].a/w829 ), .Z(n12238)
         );
  AND U5356 ( .A(\SUBBYTES[6].a/w635 ), .B(\SUBBYTES[6].a/w624 ), .Z(n12237)
         );
  AND U5357 ( .A(\SUBBYTES[6].a/w635 ), .B(\SUBBYTES[6].a/w622 ), .Z(n12236)
         );
  AND U5358 ( .A(\SUBBYTES[6].a/w428 ), .B(\SUBBYTES[6].a/w417 ), .Z(n12235)
         );
  AND U5359 ( .A(\SUBBYTES[6].a/w428 ), .B(\SUBBYTES[6].a/w415 ), .Z(n12234)
         );
  AND U5360 ( .A(\SUBBYTES[6].a/w3326 ), .B(\SUBBYTES[6].a/w3315 ), .Z(n12263)
         );
  AND U5361 ( .A(\SUBBYTES[6].a/w3326 ), .B(\SUBBYTES[6].a/w3313 ), .Z(n12262)
         );
  AND U5362 ( .A(\SUBBYTES[6].a/w3119 ), .B(\SUBBYTES[6].a/w3108 ), .Z(n12261)
         );
  AND U5363 ( .A(\SUBBYTES[6].a/w3119 ), .B(\SUBBYTES[6].a/w3106 ), .Z(n12260)
         );
  AND U5364 ( .A(\SUBBYTES[6].a/w2912 ), .B(\SUBBYTES[6].a/w2901 ), .Z(n12259)
         );
  AND U5365 ( .A(\SUBBYTES[6].a/w2912 ), .B(\SUBBYTES[6].a/w2899 ), .Z(n12258)
         );
  AND U5366 ( .A(\SUBBYTES[6].a/w2705 ), .B(\SUBBYTES[6].a/w2694 ), .Z(n12257)
         );
  AND U5367 ( .A(\SUBBYTES[6].a/w2705 ), .B(\SUBBYTES[6].a/w2692 ), .Z(n12256)
         );
  AND U5368 ( .A(\SUBBYTES[6].a/w2498 ), .B(\SUBBYTES[6].a/w2487 ), .Z(n12255)
         );
  AND U5369 ( .A(\SUBBYTES[6].a/w2498 ), .B(\SUBBYTES[6].a/w2485 ), .Z(n12254)
         );
  AND U5370 ( .A(\SUBBYTES[6].a/w2291 ), .B(\SUBBYTES[6].a/w2280 ), .Z(n12253)
         );
  AND U5371 ( .A(\SUBBYTES[6].a/w2291 ), .B(\SUBBYTES[6].a/w2278 ), .Z(n12252)
         );
  AND U5372 ( .A(\SUBBYTES[6].a/w2084 ), .B(\SUBBYTES[6].a/w2073 ), .Z(n12251)
         );
  AND U5373 ( .A(\SUBBYTES[6].a/w221 ), .B(\SUBBYTES[6].a/w210 ), .Z(n12233)
         );
  AND U5374 ( .A(n2062), .B(\SUBBYTES[5].a/w781 ), .Z(\SUBBYTES[5].a/w916 ) );
  AND U5375 ( .A(n2063), .B(\SUBBYTES[5].a/w782 ), .Z(\SUBBYTES[5].a/w914 ) );
  AND U5376 ( .A(\SUBBYTES[5].a/w912 ), .B(n2064), .Z(\SUBBYTES[5].a/w913 ) );
  ANDN U5377 ( .A(\w1[5][96] ), .B(n2065), .Z(\SUBBYTES[5].a/w909 ) );
  AND U5378 ( .A(n2066), .B(\SUBBYTES[5].a/w784 ), .Z(\SUBBYTES[5].a/w907 ) );
  AND U5379 ( .A(\SUBBYTES[5].a/w905 ), .B(n2067), .Z(\SUBBYTES[5].a/w906 ) );
  XOR U5380 ( .A(\SUBBYTES[5].a/w849 ), .B(n10958), .Z(n2067) );
  AND U5381 ( .A(\SUBBYTES[5].a/w892 ), .B(\SUBBYTES[5].a/w894 ), .Z(
        \SUBBYTES[5].a/w901 ) );
  AND U5382 ( .A(\SUBBYTES[5].a/w893 ), .B(\SUBBYTES[5].a/w895 ), .Z(
        \SUBBYTES[5].a/w899 ) );
  AND U5383 ( .A(\SUBBYTES[5].a/w896 ), .B(\SUBBYTES[5].a/w897 ), .Z(
        \SUBBYTES[5].a/w898 ) );
  AND U5384 ( .A(\SUBBYTES[5].a/w785 ), .B(n2062), .Z(\SUBBYTES[5].a/w884 ) );
  XOR U5385 ( .A(\SUBBYTES[5].a/w853 ), .B(n1024), .Z(n2062) );
  AND U5386 ( .A(\SUBBYTES[5].a/w786 ), .B(n2063), .Z(\SUBBYTES[5].a/w882 ) );
  XOR U5387 ( .A(n10959), .B(\SUBBYTES[5].a/w853 ), .Z(n2063) );
  ANDN U5388 ( .A(n2064), .B(n2068), .Z(\SUBBYTES[5].a/w881 ) );
  XOR U5389 ( .A(n1024), .B(n10959), .Z(n2064) );
  ANDN U5390 ( .A(\SUBBYTES[5].a/w787 ), .B(n2065), .Z(\SUBBYTES[5].a/w877 )
         );
  XNOR U5391 ( .A(\SUBBYTES[5].a/w846 ), .B(\SUBBYTES[5].a/w849 ), .Z(n2065)
         );
  AND U5392 ( .A(\SUBBYTES[5].a/w788 ), .B(n2066), .Z(\SUBBYTES[5].a/w875 ) );
  XNOR U5393 ( .A(n2069), .B(\SUBBYTES[5].a/w846 ), .Z(n2066) );
  AND U5394 ( .A(\SUBBYTES[5].a/w873 ), .B(n2070), .Z(\SUBBYTES[5].a/w874 ) );
  XOR U5395 ( .A(n2071), .B(n2069), .Z(n2070) );
  IV U5396 ( .A(n10958), .Z(n2069) );
  ANDN U5397 ( .A(\SUBBYTES[5].a/w892 ), .B(n2072), .Z(\SUBBYTES[5].a/w869 )
         );
  ANDN U5398 ( .A(\SUBBYTES[5].a/w893 ), .B(n2073), .Z(\SUBBYTES[5].a/w867 )
         );
  ANDN U5399 ( .A(\SUBBYTES[5].a/w896 ), .B(n2074), .Z(\SUBBYTES[5].a/w866 )
         );
  AND U5400 ( .A(\SUBBYTES[5].a/w852 ), .B(\SUBBYTES[5].a/w851 ), .Z(
        \SUBBYTES[5].a/w853 ) );
  IV U5401 ( .A(n2071), .Z(\SUBBYTES[5].a/w849 ) );
  NAND U5402 ( .A(\SUBBYTES[5].a/w828 ), .B(\SUBBYTES[5].a/w843 ), .Z(n2071)
         );
  AND U5403 ( .A(\SUBBYTES[5].a/w845 ), .B(\SUBBYTES[5].a/w851 ), .Z(
        \SUBBYTES[5].a/w846 ) );
  AND U5404 ( .A(\SUBBYTES[5].a/w830 ), .B(\SUBBYTES[5].a/w828 ), .Z(
        \SUBBYTES[5].a/w840 ) );
  AND U5405 ( .A(\SUBBYTES[5].a/w831 ), .B(\SUBBYTES[5].a/w829 ), .Z(
        \SUBBYTES[5].a/w838 ) );
  AND U5406 ( .A(\SUBBYTES[5].a/w845 ), .B(\SUBBYTES[5].a/w852 ), .Z(
        \SUBBYTES[5].a/w837 ) );
  AND U5407 ( .A(\SUBBYTES[5].a/w785 ), .B(\SUBBYTES[5].a/w781 ), .Z(
        \SUBBYTES[5].a/w822 ) );
  AND U5408 ( .A(\SUBBYTES[5].a/w786 ), .B(\SUBBYTES[5].a/w782 ), .Z(
        \SUBBYTES[5].a/w820 ) );
  ANDN U5409 ( .A(\SUBBYTES[5].a/w912 ), .B(n2068), .Z(\SUBBYTES[5].a/w819 )
         );
  XNOR U5410 ( .A(\w1[5][103] ), .B(\w1[5][97] ), .Z(n2068) );
  XOR U5411 ( .A(\w0[5][97] ), .B(g_input[737]), .Z(\w1[5][97] ) );
  IV U5412 ( .A(n2075), .Z(\w1[5][103] ) );
  AND U5413 ( .A(\w1[5][96] ), .B(\SUBBYTES[5].a/w787 ), .Z(
        \SUBBYTES[5].a/w815 ) );
  XOR U5414 ( .A(\w0[5][96] ), .B(g_input[736]), .Z(\w1[5][96] ) );
  AND U5415 ( .A(\SUBBYTES[5].a/w788 ), .B(\SUBBYTES[5].a/w784 ), .Z(
        \SUBBYTES[5].a/w813 ) );
  AND U5416 ( .A(\SUBBYTES[5].a/w873 ), .B(\SUBBYTES[5].a/w905 ), .Z(
        \SUBBYTES[5].a/w812 ) );
  ANDN U5417 ( .A(\SUBBYTES[5].a/w894 ), .B(n2072), .Z(\SUBBYTES[5].a/w807 )
         );
  XOR U5418 ( .A(\w1[5][100] ), .B(n2075), .Z(n2072) );
  ANDN U5419 ( .A(\SUBBYTES[5].a/w895 ), .B(n2073), .Z(\SUBBYTES[5].a/w805 )
         );
  XOR U5420 ( .A(n2075), .B(\w1[5][98] ), .Z(n2073) );
  XNOR U5421 ( .A(\w0[5][103] ), .B(g_input[743]), .Z(n2075) );
  ANDN U5422 ( .A(\SUBBYTES[5].a/w897 ), .B(n2074), .Z(\SUBBYTES[5].a/w804 )
         );
  XNOR U5423 ( .A(\w1[5][100] ), .B(\w1[5][98] ), .Z(n2074) );
  XOR U5424 ( .A(\w0[5][98] ), .B(g_input[738]), .Z(\w1[5][98] ) );
  XOR U5425 ( .A(\w0[5][100] ), .B(g_input[740]), .Z(\w1[5][100] ) );
  AND U5426 ( .A(n2076), .B(\SUBBYTES[5].a/w574 ), .Z(\SUBBYTES[5].a/w709 ) );
  AND U5427 ( .A(n2077), .B(\SUBBYTES[5].a/w575 ), .Z(\SUBBYTES[5].a/w707 ) );
  AND U5428 ( .A(\SUBBYTES[5].a/w705 ), .B(n2078), .Z(\SUBBYTES[5].a/w706 ) );
  ANDN U5429 ( .A(\w1[5][104] ), .B(n2079), .Z(\SUBBYTES[5].a/w702 ) );
  AND U5430 ( .A(n2080), .B(\SUBBYTES[5].a/w577 ), .Z(\SUBBYTES[5].a/w700 ) );
  AND U5431 ( .A(\SUBBYTES[5].a/w698 ), .B(n2081), .Z(\SUBBYTES[5].a/w699 ) );
  XOR U5432 ( .A(\SUBBYTES[5].a/w642 ), .B(n10956), .Z(n2081) );
  AND U5433 ( .A(\SUBBYTES[5].a/w685 ), .B(\SUBBYTES[5].a/w687 ), .Z(
        \SUBBYTES[5].a/w694 ) );
  AND U5434 ( .A(\SUBBYTES[5].a/w686 ), .B(\SUBBYTES[5].a/w688 ), .Z(
        \SUBBYTES[5].a/w692 ) );
  AND U5435 ( .A(\SUBBYTES[5].a/w689 ), .B(\SUBBYTES[5].a/w690 ), .Z(
        \SUBBYTES[5].a/w691 ) );
  AND U5436 ( .A(\SUBBYTES[5].a/w578 ), .B(n2076), .Z(\SUBBYTES[5].a/w677 ) );
  XOR U5437 ( .A(\SUBBYTES[5].a/w646 ), .B(n1023), .Z(n2076) );
  AND U5438 ( .A(\SUBBYTES[5].a/w579 ), .B(n2077), .Z(\SUBBYTES[5].a/w675 ) );
  XOR U5439 ( .A(n10957), .B(\SUBBYTES[5].a/w646 ), .Z(n2077) );
  ANDN U5440 ( .A(n2078), .B(n2082), .Z(\SUBBYTES[5].a/w674 ) );
  XOR U5441 ( .A(n1023), .B(n10957), .Z(n2078) );
  ANDN U5442 ( .A(\SUBBYTES[5].a/w580 ), .B(n2079), .Z(\SUBBYTES[5].a/w670 )
         );
  XNOR U5443 ( .A(\SUBBYTES[5].a/w639 ), .B(\SUBBYTES[5].a/w642 ), .Z(n2079)
         );
  AND U5444 ( .A(\SUBBYTES[5].a/w581 ), .B(n2080), .Z(\SUBBYTES[5].a/w668 ) );
  XNOR U5445 ( .A(n2083), .B(\SUBBYTES[5].a/w639 ), .Z(n2080) );
  AND U5446 ( .A(\SUBBYTES[5].a/w666 ), .B(n2084), .Z(\SUBBYTES[5].a/w667 ) );
  XOR U5447 ( .A(n2085), .B(n2083), .Z(n2084) );
  IV U5448 ( .A(n10956), .Z(n2083) );
  ANDN U5449 ( .A(\SUBBYTES[5].a/w685 ), .B(n2086), .Z(\SUBBYTES[5].a/w662 )
         );
  ANDN U5450 ( .A(\SUBBYTES[5].a/w686 ), .B(n2087), .Z(\SUBBYTES[5].a/w660 )
         );
  ANDN U5451 ( .A(\SUBBYTES[5].a/w689 ), .B(n2088), .Z(\SUBBYTES[5].a/w659 )
         );
  AND U5452 ( .A(\SUBBYTES[5].a/w645 ), .B(\SUBBYTES[5].a/w644 ), .Z(
        \SUBBYTES[5].a/w646 ) );
  IV U5453 ( .A(n2085), .Z(\SUBBYTES[5].a/w642 ) );
  NAND U5454 ( .A(\SUBBYTES[5].a/w621 ), .B(\SUBBYTES[5].a/w636 ), .Z(n2085)
         );
  AND U5455 ( .A(\SUBBYTES[5].a/w638 ), .B(\SUBBYTES[5].a/w644 ), .Z(
        \SUBBYTES[5].a/w639 ) );
  AND U5456 ( .A(\SUBBYTES[5].a/w623 ), .B(\SUBBYTES[5].a/w621 ), .Z(
        \SUBBYTES[5].a/w633 ) );
  AND U5457 ( .A(\SUBBYTES[5].a/w624 ), .B(\SUBBYTES[5].a/w622 ), .Z(
        \SUBBYTES[5].a/w631 ) );
  AND U5458 ( .A(\SUBBYTES[5].a/w638 ), .B(\SUBBYTES[5].a/w645 ), .Z(
        \SUBBYTES[5].a/w630 ) );
  AND U5459 ( .A(\SUBBYTES[5].a/w578 ), .B(\SUBBYTES[5].a/w574 ), .Z(
        \SUBBYTES[5].a/w615 ) );
  AND U5460 ( .A(\SUBBYTES[5].a/w579 ), .B(\SUBBYTES[5].a/w575 ), .Z(
        \SUBBYTES[5].a/w613 ) );
  ANDN U5461 ( .A(\SUBBYTES[5].a/w705 ), .B(n2082), .Z(\SUBBYTES[5].a/w612 )
         );
  XNOR U5462 ( .A(\w1[5][105] ), .B(\w1[5][111] ), .Z(n2082) );
  XOR U5463 ( .A(\w0[5][105] ), .B(g_input[745]), .Z(\w1[5][105] ) );
  AND U5464 ( .A(\w1[5][104] ), .B(\SUBBYTES[5].a/w580 ), .Z(
        \SUBBYTES[5].a/w608 ) );
  XOR U5465 ( .A(\w0[5][104] ), .B(g_input[744]), .Z(\w1[5][104] ) );
  AND U5466 ( .A(\SUBBYTES[5].a/w581 ), .B(\SUBBYTES[5].a/w577 ), .Z(
        \SUBBYTES[5].a/w606 ) );
  AND U5467 ( .A(\SUBBYTES[5].a/w666 ), .B(\SUBBYTES[5].a/w698 ), .Z(
        \SUBBYTES[5].a/w605 ) );
  ANDN U5468 ( .A(\SUBBYTES[5].a/w687 ), .B(n2086), .Z(\SUBBYTES[5].a/w600 )
         );
  XNOR U5469 ( .A(\w1[5][108] ), .B(\w1[5][111] ), .Z(n2086) );
  ANDN U5470 ( .A(\SUBBYTES[5].a/w688 ), .B(n2087), .Z(\SUBBYTES[5].a/w598 )
         );
  XNOR U5471 ( .A(\w1[5][106] ), .B(\w1[5][111] ), .Z(n2087) );
  XOR U5472 ( .A(\w0[5][111] ), .B(g_input[751]), .Z(\w1[5][111] ) );
  IV U5473 ( .A(n2089), .Z(\w1[5][106] ) );
  ANDN U5474 ( .A(\SUBBYTES[5].a/w690 ), .B(n2088), .Z(\SUBBYTES[5].a/w597 )
         );
  XOR U5475 ( .A(n2089), .B(\w1[5][108] ), .Z(n2088) );
  XOR U5476 ( .A(\w0[5][108] ), .B(g_input[748]), .Z(\w1[5][108] ) );
  XNOR U5477 ( .A(\w0[5][106] ), .B(g_input[746]), .Z(n2089) );
  AND U5478 ( .A(n2090), .B(\SUBBYTES[5].a/w367 ), .Z(\SUBBYTES[5].a/w502 ) );
  AND U5479 ( .A(n2091), .B(\SUBBYTES[5].a/w368 ), .Z(\SUBBYTES[5].a/w500 ) );
  AND U5480 ( .A(\SUBBYTES[5].a/w498 ), .B(n2092), .Z(\SUBBYTES[5].a/w499 ) );
  ANDN U5481 ( .A(\w1[5][112] ), .B(n2093), .Z(\SUBBYTES[5].a/w495 ) );
  AND U5482 ( .A(n2094), .B(\SUBBYTES[5].a/w370 ), .Z(\SUBBYTES[5].a/w493 ) );
  AND U5483 ( .A(\SUBBYTES[5].a/w491 ), .B(n2095), .Z(\SUBBYTES[5].a/w492 ) );
  XOR U5484 ( .A(\SUBBYTES[5].a/w435 ), .B(n10954), .Z(n2095) );
  AND U5485 ( .A(\SUBBYTES[5].a/w478 ), .B(\SUBBYTES[5].a/w480 ), .Z(
        \SUBBYTES[5].a/w487 ) );
  AND U5486 ( .A(\SUBBYTES[5].a/w479 ), .B(\SUBBYTES[5].a/w481 ), .Z(
        \SUBBYTES[5].a/w485 ) );
  AND U5487 ( .A(\SUBBYTES[5].a/w482 ), .B(\SUBBYTES[5].a/w483 ), .Z(
        \SUBBYTES[5].a/w484 ) );
  AND U5488 ( .A(\SUBBYTES[5].a/w371 ), .B(n2090), .Z(\SUBBYTES[5].a/w470 ) );
  XOR U5489 ( .A(\SUBBYTES[5].a/w439 ), .B(n1022), .Z(n2090) );
  AND U5490 ( .A(\SUBBYTES[5].a/w372 ), .B(n2091), .Z(\SUBBYTES[5].a/w468 ) );
  XOR U5491 ( .A(n10955), .B(\SUBBYTES[5].a/w439 ), .Z(n2091) );
  ANDN U5492 ( .A(n2092), .B(n2096), .Z(\SUBBYTES[5].a/w467 ) );
  XOR U5493 ( .A(n1022), .B(n10955), .Z(n2092) );
  ANDN U5494 ( .A(\SUBBYTES[5].a/w373 ), .B(n2093), .Z(\SUBBYTES[5].a/w463 )
         );
  XNOR U5495 ( .A(\SUBBYTES[5].a/w432 ), .B(\SUBBYTES[5].a/w435 ), .Z(n2093)
         );
  AND U5496 ( .A(\SUBBYTES[5].a/w374 ), .B(n2094), .Z(\SUBBYTES[5].a/w461 ) );
  XNOR U5497 ( .A(n2097), .B(\SUBBYTES[5].a/w432 ), .Z(n2094) );
  AND U5498 ( .A(\SUBBYTES[5].a/w459 ), .B(n2098), .Z(\SUBBYTES[5].a/w460 ) );
  XOR U5499 ( .A(n2099), .B(n2097), .Z(n2098) );
  IV U5500 ( .A(n10954), .Z(n2097) );
  ANDN U5501 ( .A(\SUBBYTES[5].a/w478 ), .B(n2100), .Z(\SUBBYTES[5].a/w455 )
         );
  ANDN U5502 ( .A(\SUBBYTES[5].a/w479 ), .B(n2101), .Z(\SUBBYTES[5].a/w453 )
         );
  ANDN U5503 ( .A(\SUBBYTES[5].a/w482 ), .B(n2102), .Z(\SUBBYTES[5].a/w452 )
         );
  AND U5504 ( .A(\SUBBYTES[5].a/w438 ), .B(\SUBBYTES[5].a/w437 ), .Z(
        \SUBBYTES[5].a/w439 ) );
  IV U5505 ( .A(n2099), .Z(\SUBBYTES[5].a/w435 ) );
  NAND U5506 ( .A(\SUBBYTES[5].a/w414 ), .B(\SUBBYTES[5].a/w429 ), .Z(n2099)
         );
  AND U5507 ( .A(\SUBBYTES[5].a/w431 ), .B(\SUBBYTES[5].a/w437 ), .Z(
        \SUBBYTES[5].a/w432 ) );
  AND U5508 ( .A(\SUBBYTES[5].a/w416 ), .B(\SUBBYTES[5].a/w414 ), .Z(
        \SUBBYTES[5].a/w426 ) );
  AND U5509 ( .A(\SUBBYTES[5].a/w417 ), .B(\SUBBYTES[5].a/w415 ), .Z(
        \SUBBYTES[5].a/w424 ) );
  AND U5510 ( .A(\SUBBYTES[5].a/w431 ), .B(\SUBBYTES[5].a/w438 ), .Z(
        \SUBBYTES[5].a/w423 ) );
  AND U5511 ( .A(\SUBBYTES[5].a/w371 ), .B(\SUBBYTES[5].a/w367 ), .Z(
        \SUBBYTES[5].a/w408 ) );
  AND U5512 ( .A(\SUBBYTES[5].a/w372 ), .B(\SUBBYTES[5].a/w368 ), .Z(
        \SUBBYTES[5].a/w406 ) );
  ANDN U5513 ( .A(\SUBBYTES[5].a/w498 ), .B(n2096), .Z(\SUBBYTES[5].a/w405 )
         );
  XNOR U5514 ( .A(\w1[5][113] ), .B(\w1[5][119] ), .Z(n2096) );
  XOR U5515 ( .A(\w0[5][113] ), .B(g_input[753]), .Z(\w1[5][113] ) );
  AND U5516 ( .A(\w1[5][112] ), .B(\SUBBYTES[5].a/w373 ), .Z(
        \SUBBYTES[5].a/w401 ) );
  XOR U5517 ( .A(\w0[5][112] ), .B(g_input[752]), .Z(\w1[5][112] ) );
  AND U5518 ( .A(\SUBBYTES[5].a/w374 ), .B(\SUBBYTES[5].a/w370 ), .Z(
        \SUBBYTES[5].a/w399 ) );
  AND U5519 ( .A(\SUBBYTES[5].a/w459 ), .B(\SUBBYTES[5].a/w491 ), .Z(
        \SUBBYTES[5].a/w398 ) );
  ANDN U5520 ( .A(\SUBBYTES[5].a/w480 ), .B(n2100), .Z(\SUBBYTES[5].a/w393 )
         );
  XNOR U5521 ( .A(\w1[5][116] ), .B(\w1[5][119] ), .Z(n2100) );
  ANDN U5522 ( .A(\SUBBYTES[5].a/w481 ), .B(n2101), .Z(\SUBBYTES[5].a/w391 )
         );
  XNOR U5523 ( .A(\w1[5][114] ), .B(\w1[5][119] ), .Z(n2101) );
  XOR U5524 ( .A(\w0[5][119] ), .B(g_input[759]), .Z(\w1[5][119] ) );
  IV U5525 ( .A(n2103), .Z(\w1[5][114] ) );
  ANDN U5526 ( .A(\SUBBYTES[5].a/w483 ), .B(n2102), .Z(\SUBBYTES[5].a/w390 )
         );
  XOR U5527 ( .A(n2103), .B(\w1[5][116] ), .Z(n2102) );
  XOR U5528 ( .A(\w0[5][116] ), .B(g_input[756]), .Z(\w1[5][116] ) );
  XNOR U5529 ( .A(\w0[5][114] ), .B(g_input[754]), .Z(n2103) );
  AND U5530 ( .A(n2104), .B(\SUBBYTES[5].a/w3265 ), .Z(\SUBBYTES[5].a/w3400 )
         );
  AND U5531 ( .A(n2105), .B(\SUBBYTES[5].a/w3266 ), .Z(\SUBBYTES[5].a/w3398 )
         );
  AND U5532 ( .A(\SUBBYTES[5].a/w3396 ), .B(n2106), .Z(\SUBBYTES[5].a/w3397 )
         );
  ANDN U5533 ( .A(\w1[5][0] ), .B(n2107), .Z(\SUBBYTES[5].a/w3393 ) );
  AND U5534 ( .A(n2108), .B(\SUBBYTES[5].a/w3268 ), .Z(\SUBBYTES[5].a/w3391 )
         );
  AND U5535 ( .A(\SUBBYTES[5].a/w3389 ), .B(n2109), .Z(\SUBBYTES[5].a/w3390 )
         );
  XOR U5536 ( .A(\SUBBYTES[5].a/w3333 ), .B(n10982), .Z(n2109) );
  AND U5537 ( .A(\SUBBYTES[5].a/w3376 ), .B(\SUBBYTES[5].a/w3378 ), .Z(
        \SUBBYTES[5].a/w3385 ) );
  AND U5538 ( .A(\SUBBYTES[5].a/w3377 ), .B(\SUBBYTES[5].a/w3379 ), .Z(
        \SUBBYTES[5].a/w3383 ) );
  AND U5539 ( .A(\SUBBYTES[5].a/w3380 ), .B(\SUBBYTES[5].a/w3381 ), .Z(
        \SUBBYTES[5].a/w3382 ) );
  AND U5540 ( .A(\SUBBYTES[5].a/w3269 ), .B(n2104), .Z(\SUBBYTES[5].a/w3368 )
         );
  XOR U5541 ( .A(\SUBBYTES[5].a/w3337 ), .B(n1036), .Z(n2104) );
  AND U5542 ( .A(\SUBBYTES[5].a/w3270 ), .B(n2105), .Z(\SUBBYTES[5].a/w3366 )
         );
  XOR U5543 ( .A(n10983), .B(\SUBBYTES[5].a/w3337 ), .Z(n2105) );
  ANDN U5544 ( .A(n2106), .B(n2110), .Z(\SUBBYTES[5].a/w3365 ) );
  XOR U5545 ( .A(n1036), .B(n10983), .Z(n2106) );
  ANDN U5546 ( .A(\SUBBYTES[5].a/w3271 ), .B(n2107), .Z(\SUBBYTES[5].a/w3361 )
         );
  XNOR U5547 ( .A(\SUBBYTES[5].a/w3330 ), .B(\SUBBYTES[5].a/w3333 ), .Z(n2107)
         );
  AND U5548 ( .A(\SUBBYTES[5].a/w3272 ), .B(n2108), .Z(\SUBBYTES[5].a/w3359 )
         );
  XNOR U5549 ( .A(n2111), .B(\SUBBYTES[5].a/w3330 ), .Z(n2108) );
  AND U5550 ( .A(\SUBBYTES[5].a/w3357 ), .B(n2112), .Z(\SUBBYTES[5].a/w3358 )
         );
  XOR U5551 ( .A(n2113), .B(n2111), .Z(n2112) );
  IV U5552 ( .A(n10982), .Z(n2111) );
  ANDN U5553 ( .A(\SUBBYTES[5].a/w3376 ), .B(n2114), .Z(\SUBBYTES[5].a/w3353 )
         );
  ANDN U5554 ( .A(\SUBBYTES[5].a/w3377 ), .B(n2115), .Z(\SUBBYTES[5].a/w3351 )
         );
  ANDN U5555 ( .A(\SUBBYTES[5].a/w3380 ), .B(n2116), .Z(\SUBBYTES[5].a/w3350 )
         );
  AND U5556 ( .A(\SUBBYTES[5].a/w3336 ), .B(\SUBBYTES[5].a/w3335 ), .Z(
        \SUBBYTES[5].a/w3337 ) );
  IV U5557 ( .A(n2113), .Z(\SUBBYTES[5].a/w3333 ) );
  NAND U5558 ( .A(\SUBBYTES[5].a/w3312 ), .B(\SUBBYTES[5].a/w3327 ), .Z(n2113)
         );
  AND U5559 ( .A(\SUBBYTES[5].a/w3329 ), .B(\SUBBYTES[5].a/w3335 ), .Z(
        \SUBBYTES[5].a/w3330 ) );
  AND U5560 ( .A(\SUBBYTES[5].a/w3314 ), .B(\SUBBYTES[5].a/w3312 ), .Z(
        \SUBBYTES[5].a/w3324 ) );
  AND U5561 ( .A(\SUBBYTES[5].a/w3315 ), .B(\SUBBYTES[5].a/w3313 ), .Z(
        \SUBBYTES[5].a/w3322 ) );
  AND U5562 ( .A(\SUBBYTES[5].a/w3329 ), .B(\SUBBYTES[5].a/w3336 ), .Z(
        \SUBBYTES[5].a/w3321 ) );
  AND U5563 ( .A(\SUBBYTES[5].a/w3269 ), .B(\SUBBYTES[5].a/w3265 ), .Z(
        \SUBBYTES[5].a/w3306 ) );
  AND U5564 ( .A(\SUBBYTES[5].a/w3270 ), .B(\SUBBYTES[5].a/w3266 ), .Z(
        \SUBBYTES[5].a/w3304 ) );
  ANDN U5565 ( .A(\SUBBYTES[5].a/w3396 ), .B(n2110), .Z(\SUBBYTES[5].a/w3303 )
         );
  XNOR U5566 ( .A(\w1[5][1] ), .B(\w1[5][7] ), .Z(n2110) );
  XOR U5567 ( .A(\w0[5][1] ), .B(g_input[641]), .Z(\w1[5][1] ) );
  AND U5568 ( .A(\w1[5][0] ), .B(\SUBBYTES[5].a/w3271 ), .Z(
        \SUBBYTES[5].a/w3299 ) );
  XOR U5569 ( .A(\w0[5][0] ), .B(g_input[640]), .Z(\w1[5][0] ) );
  AND U5570 ( .A(\SUBBYTES[5].a/w3272 ), .B(\SUBBYTES[5].a/w3268 ), .Z(
        \SUBBYTES[5].a/w3297 ) );
  AND U5571 ( .A(\SUBBYTES[5].a/w3357 ), .B(\SUBBYTES[5].a/w3389 ), .Z(
        \SUBBYTES[5].a/w3296 ) );
  ANDN U5572 ( .A(\SUBBYTES[5].a/w3378 ), .B(n2114), .Z(\SUBBYTES[5].a/w3291 )
         );
  XNOR U5573 ( .A(\w1[5][4] ), .B(\w1[5][7] ), .Z(n2114) );
  ANDN U5574 ( .A(\SUBBYTES[5].a/w3379 ), .B(n2115), .Z(\SUBBYTES[5].a/w3289 )
         );
  XNOR U5575 ( .A(\w1[5][2] ), .B(\w1[5][7] ), .Z(n2115) );
  XOR U5576 ( .A(\w0[5][7] ), .B(g_input[647]), .Z(\w1[5][7] ) );
  IV U5577 ( .A(n2117), .Z(\w1[5][2] ) );
  ANDN U5578 ( .A(\SUBBYTES[5].a/w3381 ), .B(n2116), .Z(\SUBBYTES[5].a/w3288 )
         );
  XOR U5579 ( .A(n2117), .B(\w1[5][4] ), .Z(n2116) );
  XOR U5580 ( .A(\w0[5][4] ), .B(g_input[644]), .Z(\w1[5][4] ) );
  XNOR U5581 ( .A(\w0[5][2] ), .B(g_input[642]), .Z(n2117) );
  AND U5582 ( .A(n2118), .B(\SUBBYTES[5].a/w3058 ), .Z(\SUBBYTES[5].a/w3193 )
         );
  AND U5583 ( .A(n2119), .B(\SUBBYTES[5].a/w3059 ), .Z(\SUBBYTES[5].a/w3191 )
         );
  AND U5584 ( .A(\SUBBYTES[5].a/w3189 ), .B(n2120), .Z(\SUBBYTES[5].a/w3190 )
         );
  ANDN U5585 ( .A(\w1[5][8] ), .B(n2121), .Z(\SUBBYTES[5].a/w3186 ) );
  AND U5586 ( .A(n2122), .B(\SUBBYTES[5].a/w3061 ), .Z(\SUBBYTES[5].a/w3184 )
         );
  AND U5587 ( .A(\SUBBYTES[5].a/w3182 ), .B(n2123), .Z(\SUBBYTES[5].a/w3183 )
         );
  XOR U5588 ( .A(\SUBBYTES[5].a/w3126 ), .B(n10980), .Z(n2123) );
  AND U5589 ( .A(\SUBBYTES[5].a/w3169 ), .B(\SUBBYTES[5].a/w3171 ), .Z(
        \SUBBYTES[5].a/w3178 ) );
  AND U5590 ( .A(\SUBBYTES[5].a/w3170 ), .B(\SUBBYTES[5].a/w3172 ), .Z(
        \SUBBYTES[5].a/w3176 ) );
  AND U5591 ( .A(\SUBBYTES[5].a/w3173 ), .B(\SUBBYTES[5].a/w3174 ), .Z(
        \SUBBYTES[5].a/w3175 ) );
  AND U5592 ( .A(\SUBBYTES[5].a/w3062 ), .B(n2118), .Z(\SUBBYTES[5].a/w3161 )
         );
  XOR U5593 ( .A(\SUBBYTES[5].a/w3130 ), .B(n1035), .Z(n2118) );
  AND U5594 ( .A(\SUBBYTES[5].a/w3063 ), .B(n2119), .Z(\SUBBYTES[5].a/w3159 )
         );
  XOR U5595 ( .A(n10981), .B(\SUBBYTES[5].a/w3130 ), .Z(n2119) );
  ANDN U5596 ( .A(n2120), .B(n2124), .Z(\SUBBYTES[5].a/w3158 ) );
  XOR U5597 ( .A(n1035), .B(n10981), .Z(n2120) );
  ANDN U5598 ( .A(\SUBBYTES[5].a/w3064 ), .B(n2121), .Z(\SUBBYTES[5].a/w3154 )
         );
  XNOR U5599 ( .A(\SUBBYTES[5].a/w3123 ), .B(\SUBBYTES[5].a/w3126 ), .Z(n2121)
         );
  AND U5600 ( .A(\SUBBYTES[5].a/w3065 ), .B(n2122), .Z(\SUBBYTES[5].a/w3152 )
         );
  XNOR U5601 ( .A(n2125), .B(\SUBBYTES[5].a/w3123 ), .Z(n2122) );
  AND U5602 ( .A(\SUBBYTES[5].a/w3150 ), .B(n2126), .Z(\SUBBYTES[5].a/w3151 )
         );
  XOR U5603 ( .A(n2127), .B(n2125), .Z(n2126) );
  IV U5604 ( .A(n10980), .Z(n2125) );
  ANDN U5605 ( .A(\SUBBYTES[5].a/w3169 ), .B(n2128), .Z(\SUBBYTES[5].a/w3146 )
         );
  ANDN U5606 ( .A(\SUBBYTES[5].a/w3170 ), .B(n2129), .Z(\SUBBYTES[5].a/w3144 )
         );
  ANDN U5607 ( .A(\SUBBYTES[5].a/w3173 ), .B(n2130), .Z(\SUBBYTES[5].a/w3143 )
         );
  AND U5608 ( .A(\SUBBYTES[5].a/w3129 ), .B(\SUBBYTES[5].a/w3128 ), .Z(
        \SUBBYTES[5].a/w3130 ) );
  IV U5609 ( .A(n2127), .Z(\SUBBYTES[5].a/w3126 ) );
  NAND U5610 ( .A(\SUBBYTES[5].a/w3105 ), .B(\SUBBYTES[5].a/w3120 ), .Z(n2127)
         );
  AND U5611 ( .A(\SUBBYTES[5].a/w3122 ), .B(\SUBBYTES[5].a/w3128 ), .Z(
        \SUBBYTES[5].a/w3123 ) );
  AND U5612 ( .A(\SUBBYTES[5].a/w3107 ), .B(\SUBBYTES[5].a/w3105 ), .Z(
        \SUBBYTES[5].a/w3117 ) );
  AND U5613 ( .A(\SUBBYTES[5].a/w3108 ), .B(\SUBBYTES[5].a/w3106 ), .Z(
        \SUBBYTES[5].a/w3115 ) );
  AND U5614 ( .A(\SUBBYTES[5].a/w3122 ), .B(\SUBBYTES[5].a/w3129 ), .Z(
        \SUBBYTES[5].a/w3114 ) );
  AND U5615 ( .A(\SUBBYTES[5].a/w3062 ), .B(\SUBBYTES[5].a/w3058 ), .Z(
        \SUBBYTES[5].a/w3099 ) );
  AND U5616 ( .A(\SUBBYTES[5].a/w3063 ), .B(\SUBBYTES[5].a/w3059 ), .Z(
        \SUBBYTES[5].a/w3097 ) );
  ANDN U5617 ( .A(\SUBBYTES[5].a/w3189 ), .B(n2124), .Z(\SUBBYTES[5].a/w3096 )
         );
  XNOR U5618 ( .A(\w1[5][15] ), .B(\w1[5][9] ), .Z(n2124) );
  XOR U5619 ( .A(\w0[5][9] ), .B(g_input[649]), .Z(\w1[5][9] ) );
  AND U5620 ( .A(\w1[5][8] ), .B(\SUBBYTES[5].a/w3064 ), .Z(
        \SUBBYTES[5].a/w3092 ) );
  XOR U5621 ( .A(\w0[5][8] ), .B(g_input[648]), .Z(\w1[5][8] ) );
  AND U5622 ( .A(\SUBBYTES[5].a/w3065 ), .B(\SUBBYTES[5].a/w3061 ), .Z(
        \SUBBYTES[5].a/w3090 ) );
  AND U5623 ( .A(\SUBBYTES[5].a/w3150 ), .B(\SUBBYTES[5].a/w3182 ), .Z(
        \SUBBYTES[5].a/w3089 ) );
  ANDN U5624 ( .A(\SUBBYTES[5].a/w3171 ), .B(n2128), .Z(\SUBBYTES[5].a/w3084 )
         );
  XNOR U5625 ( .A(\w1[5][12] ), .B(\w1[5][15] ), .Z(n2128) );
  ANDN U5626 ( .A(\SUBBYTES[5].a/w3172 ), .B(n2129), .Z(\SUBBYTES[5].a/w3082 )
         );
  XNOR U5627 ( .A(\w1[5][10] ), .B(\w1[5][15] ), .Z(n2129) );
  XOR U5628 ( .A(\w0[5][15] ), .B(g_input[655]), .Z(\w1[5][15] ) );
  ANDN U5629 ( .A(\SUBBYTES[5].a/w3174 ), .B(n2130), .Z(\SUBBYTES[5].a/w3081 )
         );
  XNOR U5630 ( .A(\w1[5][10] ), .B(\w1[5][12] ), .Z(n2130) );
  XOR U5631 ( .A(\w0[5][12] ), .B(g_input[652]), .Z(\w1[5][12] ) );
  XOR U5632 ( .A(\w0[5][10] ), .B(g_input[650]), .Z(\w1[5][10] ) );
  AND U5633 ( .A(n2131), .B(\SUBBYTES[5].a/w2851 ), .Z(\SUBBYTES[5].a/w2986 )
         );
  AND U5634 ( .A(n2132), .B(\SUBBYTES[5].a/w2852 ), .Z(\SUBBYTES[5].a/w2984 )
         );
  AND U5635 ( .A(\SUBBYTES[5].a/w2982 ), .B(n2133), .Z(\SUBBYTES[5].a/w2983 )
         );
  ANDN U5636 ( .A(\w1[5][16] ), .B(n2134), .Z(\SUBBYTES[5].a/w2979 ) );
  AND U5637 ( .A(n2135), .B(\SUBBYTES[5].a/w2854 ), .Z(\SUBBYTES[5].a/w2977 )
         );
  AND U5638 ( .A(\SUBBYTES[5].a/w2975 ), .B(n2136), .Z(\SUBBYTES[5].a/w2976 )
         );
  XOR U5639 ( .A(\SUBBYTES[5].a/w2919 ), .B(n10978), .Z(n2136) );
  AND U5640 ( .A(\SUBBYTES[5].a/w2962 ), .B(\SUBBYTES[5].a/w2964 ), .Z(
        \SUBBYTES[5].a/w2971 ) );
  AND U5641 ( .A(\SUBBYTES[5].a/w2963 ), .B(\SUBBYTES[5].a/w2965 ), .Z(
        \SUBBYTES[5].a/w2969 ) );
  AND U5642 ( .A(\SUBBYTES[5].a/w2966 ), .B(\SUBBYTES[5].a/w2967 ), .Z(
        \SUBBYTES[5].a/w2968 ) );
  AND U5643 ( .A(\SUBBYTES[5].a/w2855 ), .B(n2131), .Z(\SUBBYTES[5].a/w2954 )
         );
  XOR U5644 ( .A(\SUBBYTES[5].a/w2923 ), .B(n1034), .Z(n2131) );
  AND U5645 ( .A(\SUBBYTES[5].a/w2856 ), .B(n2132), .Z(\SUBBYTES[5].a/w2952 )
         );
  XOR U5646 ( .A(n10979), .B(\SUBBYTES[5].a/w2923 ), .Z(n2132) );
  ANDN U5647 ( .A(n2133), .B(n2137), .Z(\SUBBYTES[5].a/w2951 ) );
  XOR U5648 ( .A(n1034), .B(n10979), .Z(n2133) );
  AND U5649 ( .A(n2138), .B(\SUBBYTES[5].a/w160 ), .Z(\SUBBYTES[5].a/w295 ) );
  ANDN U5650 ( .A(\SUBBYTES[5].a/w2857 ), .B(n2134), .Z(\SUBBYTES[5].a/w2947 )
         );
  XNOR U5651 ( .A(\SUBBYTES[5].a/w2916 ), .B(\SUBBYTES[5].a/w2919 ), .Z(n2134)
         );
  AND U5652 ( .A(\SUBBYTES[5].a/w2858 ), .B(n2135), .Z(\SUBBYTES[5].a/w2945 )
         );
  XNOR U5653 ( .A(n2139), .B(\SUBBYTES[5].a/w2916 ), .Z(n2135) );
  AND U5654 ( .A(\SUBBYTES[5].a/w2943 ), .B(n2140), .Z(\SUBBYTES[5].a/w2944 )
         );
  XOR U5655 ( .A(n2141), .B(n2139), .Z(n2140) );
  IV U5656 ( .A(n10978), .Z(n2139) );
  ANDN U5657 ( .A(\SUBBYTES[5].a/w2962 ), .B(n2142), .Z(\SUBBYTES[5].a/w2939 )
         );
  ANDN U5658 ( .A(\SUBBYTES[5].a/w2963 ), .B(n2143), .Z(\SUBBYTES[5].a/w2937 )
         );
  ANDN U5659 ( .A(\SUBBYTES[5].a/w2966 ), .B(n2144), .Z(\SUBBYTES[5].a/w2936 )
         );
  AND U5660 ( .A(n2145), .B(\SUBBYTES[5].a/w161 ), .Z(\SUBBYTES[5].a/w293 ) );
  AND U5661 ( .A(\SUBBYTES[5].a/w2922 ), .B(\SUBBYTES[5].a/w2921 ), .Z(
        \SUBBYTES[5].a/w2923 ) );
  AND U5662 ( .A(\SUBBYTES[5].a/w291 ), .B(n2146), .Z(\SUBBYTES[5].a/w292 ) );
  IV U5663 ( .A(n2141), .Z(\SUBBYTES[5].a/w2919 ) );
  NAND U5664 ( .A(\SUBBYTES[5].a/w2898 ), .B(\SUBBYTES[5].a/w2913 ), .Z(n2141)
         );
  AND U5665 ( .A(\SUBBYTES[5].a/w2915 ), .B(\SUBBYTES[5].a/w2921 ), .Z(
        \SUBBYTES[5].a/w2916 ) );
  AND U5666 ( .A(\SUBBYTES[5].a/w2900 ), .B(\SUBBYTES[5].a/w2898 ), .Z(
        \SUBBYTES[5].a/w2910 ) );
  AND U5667 ( .A(\SUBBYTES[5].a/w2901 ), .B(\SUBBYTES[5].a/w2899 ), .Z(
        \SUBBYTES[5].a/w2908 ) );
  AND U5668 ( .A(\SUBBYTES[5].a/w2915 ), .B(\SUBBYTES[5].a/w2922 ), .Z(
        \SUBBYTES[5].a/w2907 ) );
  AND U5669 ( .A(\SUBBYTES[5].a/w2855 ), .B(\SUBBYTES[5].a/w2851 ), .Z(
        \SUBBYTES[5].a/w2892 ) );
  AND U5670 ( .A(\SUBBYTES[5].a/w2856 ), .B(\SUBBYTES[5].a/w2852 ), .Z(
        \SUBBYTES[5].a/w2890 ) );
  ANDN U5671 ( .A(\SUBBYTES[5].a/w2982 ), .B(n2137), .Z(\SUBBYTES[5].a/w2889 )
         );
  XNOR U5672 ( .A(\w1[5][17] ), .B(\w1[5][23] ), .Z(n2137) );
  XOR U5673 ( .A(\w0[5][17] ), .B(g_input[657]), .Z(\w1[5][17] ) );
  AND U5674 ( .A(\w1[5][16] ), .B(\SUBBYTES[5].a/w2857 ), .Z(
        \SUBBYTES[5].a/w2885 ) );
  XOR U5675 ( .A(\w0[5][16] ), .B(g_input[656]), .Z(\w1[5][16] ) );
  AND U5676 ( .A(\SUBBYTES[5].a/w2858 ), .B(\SUBBYTES[5].a/w2854 ), .Z(
        \SUBBYTES[5].a/w2883 ) );
  AND U5677 ( .A(\SUBBYTES[5].a/w2943 ), .B(\SUBBYTES[5].a/w2975 ), .Z(
        \SUBBYTES[5].a/w2882 ) );
  ANDN U5678 ( .A(\w1[5][120] ), .B(n2147), .Z(\SUBBYTES[5].a/w288 ) );
  ANDN U5679 ( .A(\SUBBYTES[5].a/w2964 ), .B(n2142), .Z(\SUBBYTES[5].a/w2877 )
         );
  XNOR U5680 ( .A(\w1[5][20] ), .B(\w1[5][23] ), .Z(n2142) );
  ANDN U5681 ( .A(\SUBBYTES[5].a/w2965 ), .B(n2143), .Z(\SUBBYTES[5].a/w2875 )
         );
  XNOR U5682 ( .A(\w1[5][18] ), .B(\w1[5][23] ), .Z(n2143) );
  XOR U5683 ( .A(\w0[5][23] ), .B(g_input[663]), .Z(\w1[5][23] ) );
  IV U5684 ( .A(n2148), .Z(\w1[5][18] ) );
  ANDN U5685 ( .A(\SUBBYTES[5].a/w2967 ), .B(n2144), .Z(\SUBBYTES[5].a/w2874 )
         );
  XOR U5686 ( .A(n2148), .B(\w1[5][20] ), .Z(n2144) );
  XOR U5687 ( .A(\w0[5][20] ), .B(g_input[660]), .Z(\w1[5][20] ) );
  XNOR U5688 ( .A(\w0[5][18] ), .B(g_input[658]), .Z(n2148) );
  AND U5689 ( .A(n2149), .B(\SUBBYTES[5].a/w163 ), .Z(\SUBBYTES[5].a/w286 ) );
  AND U5690 ( .A(\SUBBYTES[5].a/w284 ), .B(n2150), .Z(\SUBBYTES[5].a/w285 ) );
  XOR U5691 ( .A(\SUBBYTES[5].a/w228 ), .B(n10952), .Z(n2150) );
  AND U5692 ( .A(\SUBBYTES[5].a/w271 ), .B(\SUBBYTES[5].a/w273 ), .Z(
        \SUBBYTES[5].a/w280 ) );
  AND U5693 ( .A(\SUBBYTES[5].a/w272 ), .B(\SUBBYTES[5].a/w274 ), .Z(
        \SUBBYTES[5].a/w278 ) );
  AND U5694 ( .A(n2151), .B(\SUBBYTES[5].a/w2644 ), .Z(\SUBBYTES[5].a/w2779 )
         );
  AND U5695 ( .A(n2152), .B(\SUBBYTES[5].a/w2645 ), .Z(\SUBBYTES[5].a/w2777 )
         );
  AND U5696 ( .A(\SUBBYTES[5].a/w2775 ), .B(n2153), .Z(\SUBBYTES[5].a/w2776 )
         );
  ANDN U5697 ( .A(\w1[5][24] ), .B(n2154), .Z(\SUBBYTES[5].a/w2772 ) );
  AND U5698 ( .A(n2155), .B(\SUBBYTES[5].a/w2647 ), .Z(\SUBBYTES[5].a/w2770 )
         );
  AND U5699 ( .A(\SUBBYTES[5].a/w275 ), .B(\SUBBYTES[5].a/w276 ), .Z(
        \SUBBYTES[5].a/w277 ) );
  AND U5700 ( .A(\SUBBYTES[5].a/w2768 ), .B(n2156), .Z(\SUBBYTES[5].a/w2769 )
         );
  XOR U5701 ( .A(\SUBBYTES[5].a/w2712 ), .B(n10976), .Z(n2156) );
  AND U5702 ( .A(\SUBBYTES[5].a/w2755 ), .B(\SUBBYTES[5].a/w2757 ), .Z(
        \SUBBYTES[5].a/w2764 ) );
  AND U5703 ( .A(\SUBBYTES[5].a/w2756 ), .B(\SUBBYTES[5].a/w2758 ), .Z(
        \SUBBYTES[5].a/w2762 ) );
  AND U5704 ( .A(\SUBBYTES[5].a/w2759 ), .B(\SUBBYTES[5].a/w2760 ), .Z(
        \SUBBYTES[5].a/w2761 ) );
  AND U5705 ( .A(\SUBBYTES[5].a/w2648 ), .B(n2151), .Z(\SUBBYTES[5].a/w2747 )
         );
  XOR U5706 ( .A(\SUBBYTES[5].a/w2716 ), .B(n1033), .Z(n2151) );
  AND U5707 ( .A(\SUBBYTES[5].a/w2649 ), .B(n2152), .Z(\SUBBYTES[5].a/w2745 )
         );
  XOR U5708 ( .A(n10977), .B(\SUBBYTES[5].a/w2716 ), .Z(n2152) );
  ANDN U5709 ( .A(n2153), .B(n2157), .Z(\SUBBYTES[5].a/w2744 ) );
  XOR U5710 ( .A(n1033), .B(n10977), .Z(n2153) );
  ANDN U5711 ( .A(\SUBBYTES[5].a/w2650 ), .B(n2154), .Z(\SUBBYTES[5].a/w2740 )
         );
  XNOR U5712 ( .A(\SUBBYTES[5].a/w2709 ), .B(\SUBBYTES[5].a/w2712 ), .Z(n2154)
         );
  AND U5713 ( .A(\SUBBYTES[5].a/w2651 ), .B(n2155), .Z(\SUBBYTES[5].a/w2738 )
         );
  XNOR U5714 ( .A(n2158), .B(\SUBBYTES[5].a/w2709 ), .Z(n2155) );
  AND U5715 ( .A(\SUBBYTES[5].a/w2736 ), .B(n2159), .Z(\SUBBYTES[5].a/w2737 )
         );
  XOR U5716 ( .A(n2160), .B(n2158), .Z(n2159) );
  IV U5717 ( .A(n10976), .Z(n2158) );
  ANDN U5718 ( .A(\SUBBYTES[5].a/w2755 ), .B(n2161), .Z(\SUBBYTES[5].a/w2732 )
         );
  ANDN U5719 ( .A(\SUBBYTES[5].a/w2756 ), .B(n2162), .Z(\SUBBYTES[5].a/w2730 )
         );
  ANDN U5720 ( .A(\SUBBYTES[5].a/w2759 ), .B(n2163), .Z(\SUBBYTES[5].a/w2729 )
         );
  AND U5721 ( .A(\SUBBYTES[5].a/w2715 ), .B(\SUBBYTES[5].a/w2714 ), .Z(
        \SUBBYTES[5].a/w2716 ) );
  IV U5722 ( .A(n2160), .Z(\SUBBYTES[5].a/w2712 ) );
  NAND U5723 ( .A(\SUBBYTES[5].a/w2691 ), .B(\SUBBYTES[5].a/w2706 ), .Z(n2160)
         );
  AND U5724 ( .A(\SUBBYTES[5].a/w2708 ), .B(\SUBBYTES[5].a/w2714 ), .Z(
        \SUBBYTES[5].a/w2709 ) );
  AND U5725 ( .A(\SUBBYTES[5].a/w2693 ), .B(\SUBBYTES[5].a/w2691 ), .Z(
        \SUBBYTES[5].a/w2703 ) );
  AND U5726 ( .A(\SUBBYTES[5].a/w2694 ), .B(\SUBBYTES[5].a/w2692 ), .Z(
        \SUBBYTES[5].a/w2701 ) );
  AND U5727 ( .A(\SUBBYTES[5].a/w2708 ), .B(\SUBBYTES[5].a/w2715 ), .Z(
        \SUBBYTES[5].a/w2700 ) );
  AND U5728 ( .A(\SUBBYTES[5].a/w2648 ), .B(\SUBBYTES[5].a/w2644 ), .Z(
        \SUBBYTES[5].a/w2685 ) );
  AND U5729 ( .A(\SUBBYTES[5].a/w2649 ), .B(\SUBBYTES[5].a/w2645 ), .Z(
        \SUBBYTES[5].a/w2683 ) );
  ANDN U5730 ( .A(\SUBBYTES[5].a/w2775 ), .B(n2157), .Z(\SUBBYTES[5].a/w2682 )
         );
  XNOR U5731 ( .A(\w1[5][25] ), .B(\w1[5][31] ), .Z(n2157) );
  XOR U5732 ( .A(\w0[5][25] ), .B(g_input[665]), .Z(\w1[5][25] ) );
  AND U5733 ( .A(\w1[5][24] ), .B(\SUBBYTES[5].a/w2650 ), .Z(
        \SUBBYTES[5].a/w2678 ) );
  XOR U5734 ( .A(\w0[5][24] ), .B(g_input[664]), .Z(\w1[5][24] ) );
  AND U5735 ( .A(\SUBBYTES[5].a/w2651 ), .B(\SUBBYTES[5].a/w2647 ), .Z(
        \SUBBYTES[5].a/w2676 ) );
  AND U5736 ( .A(\SUBBYTES[5].a/w2736 ), .B(\SUBBYTES[5].a/w2768 ), .Z(
        \SUBBYTES[5].a/w2675 ) );
  ANDN U5737 ( .A(\SUBBYTES[5].a/w2757 ), .B(n2161), .Z(\SUBBYTES[5].a/w2670 )
         );
  XNOR U5738 ( .A(\w1[5][28] ), .B(\w1[5][31] ), .Z(n2161) );
  ANDN U5739 ( .A(\SUBBYTES[5].a/w2758 ), .B(n2162), .Z(\SUBBYTES[5].a/w2668 )
         );
  XNOR U5740 ( .A(\w1[5][26] ), .B(\w1[5][31] ), .Z(n2162) );
  XOR U5741 ( .A(\w0[5][31] ), .B(g_input[671]), .Z(\w1[5][31] ) );
  IV U5742 ( .A(n2164), .Z(\w1[5][26] ) );
  ANDN U5743 ( .A(\SUBBYTES[5].a/w2760 ), .B(n2163), .Z(\SUBBYTES[5].a/w2667 )
         );
  XOR U5744 ( .A(n2164), .B(\w1[5][28] ), .Z(n2163) );
  XOR U5745 ( .A(\w0[5][28] ), .B(g_input[668]), .Z(\w1[5][28] ) );
  XNOR U5746 ( .A(\w0[5][26] ), .B(g_input[666]), .Z(n2164) );
  AND U5747 ( .A(\SUBBYTES[5].a/w164 ), .B(n2138), .Z(\SUBBYTES[5].a/w263 ) );
  XOR U5748 ( .A(\SUBBYTES[5].a/w232 ), .B(n1021), .Z(n2138) );
  AND U5749 ( .A(\SUBBYTES[5].a/w165 ), .B(n2145), .Z(\SUBBYTES[5].a/w261 ) );
  XOR U5750 ( .A(n10953), .B(\SUBBYTES[5].a/w232 ), .Z(n2145) );
  ANDN U5751 ( .A(n2146), .B(n2165), .Z(\SUBBYTES[5].a/w260 ) );
  XOR U5752 ( .A(n1021), .B(n10953), .Z(n2146) );
  AND U5753 ( .A(n2166), .B(\SUBBYTES[5].a/w2437 ), .Z(\SUBBYTES[5].a/w2572 )
         );
  AND U5754 ( .A(n2167), .B(\SUBBYTES[5].a/w2438 ), .Z(\SUBBYTES[5].a/w2570 )
         );
  AND U5755 ( .A(\SUBBYTES[5].a/w2568 ), .B(n2168), .Z(\SUBBYTES[5].a/w2569 )
         );
  ANDN U5756 ( .A(\w1[5][32] ), .B(n2169), .Z(\SUBBYTES[5].a/w2565 ) );
  AND U5757 ( .A(n2170), .B(\SUBBYTES[5].a/w2440 ), .Z(\SUBBYTES[5].a/w2563 )
         );
  AND U5758 ( .A(\SUBBYTES[5].a/w2561 ), .B(n2171), .Z(\SUBBYTES[5].a/w2562 )
         );
  XOR U5759 ( .A(\SUBBYTES[5].a/w2505 ), .B(n10974), .Z(n2171) );
  ANDN U5760 ( .A(\SUBBYTES[5].a/w166 ), .B(n2147), .Z(\SUBBYTES[5].a/w256 )
         );
  XNOR U5761 ( .A(\SUBBYTES[5].a/w225 ), .B(\SUBBYTES[5].a/w228 ), .Z(n2147)
         );
  AND U5762 ( .A(\SUBBYTES[5].a/w2548 ), .B(\SUBBYTES[5].a/w2550 ), .Z(
        \SUBBYTES[5].a/w2557 ) );
  AND U5763 ( .A(\SUBBYTES[5].a/w2549 ), .B(\SUBBYTES[5].a/w2551 ), .Z(
        \SUBBYTES[5].a/w2555 ) );
  AND U5764 ( .A(\SUBBYTES[5].a/w2552 ), .B(\SUBBYTES[5].a/w2553 ), .Z(
        \SUBBYTES[5].a/w2554 ) );
  AND U5765 ( .A(\SUBBYTES[5].a/w2441 ), .B(n2166), .Z(\SUBBYTES[5].a/w2540 )
         );
  XOR U5766 ( .A(\SUBBYTES[5].a/w2509 ), .B(n1032), .Z(n2166) );
  AND U5767 ( .A(\SUBBYTES[5].a/w167 ), .B(n2149), .Z(\SUBBYTES[5].a/w254 ) );
  XNOR U5768 ( .A(n2172), .B(\SUBBYTES[5].a/w225 ), .Z(n2149) );
  AND U5769 ( .A(\SUBBYTES[5].a/w2442 ), .B(n2167), .Z(\SUBBYTES[5].a/w2538 )
         );
  XOR U5770 ( .A(n10975), .B(\SUBBYTES[5].a/w2509 ), .Z(n2167) );
  ANDN U5771 ( .A(n2168), .B(n2173), .Z(\SUBBYTES[5].a/w2537 ) );
  XOR U5772 ( .A(n1032), .B(n10975), .Z(n2168) );
  ANDN U5773 ( .A(\SUBBYTES[5].a/w2443 ), .B(n2169), .Z(\SUBBYTES[5].a/w2533 )
         );
  XNOR U5774 ( .A(\SUBBYTES[5].a/w2502 ), .B(\SUBBYTES[5].a/w2505 ), .Z(n2169)
         );
  AND U5775 ( .A(\SUBBYTES[5].a/w2444 ), .B(n2170), .Z(\SUBBYTES[5].a/w2531 )
         );
  XNOR U5776 ( .A(n2174), .B(\SUBBYTES[5].a/w2502 ), .Z(n2170) );
  AND U5777 ( .A(\SUBBYTES[5].a/w2529 ), .B(n2175), .Z(\SUBBYTES[5].a/w2530 )
         );
  XOR U5778 ( .A(n2176), .B(n2174), .Z(n2175) );
  IV U5779 ( .A(n10974), .Z(n2174) );
  AND U5780 ( .A(\SUBBYTES[5].a/w252 ), .B(n2177), .Z(\SUBBYTES[5].a/w253 ) );
  XOR U5781 ( .A(n2178), .B(n2172), .Z(n2177) );
  IV U5782 ( .A(n10952), .Z(n2172) );
  ANDN U5783 ( .A(\SUBBYTES[5].a/w2548 ), .B(n2179), .Z(\SUBBYTES[5].a/w2525 )
         );
  ANDN U5784 ( .A(\SUBBYTES[5].a/w2549 ), .B(n2180), .Z(\SUBBYTES[5].a/w2523 )
         );
  ANDN U5785 ( .A(\SUBBYTES[5].a/w2552 ), .B(n2181), .Z(\SUBBYTES[5].a/w2522 )
         );
  AND U5786 ( .A(\SUBBYTES[5].a/w2508 ), .B(\SUBBYTES[5].a/w2507 ), .Z(
        \SUBBYTES[5].a/w2509 ) );
  IV U5787 ( .A(n2176), .Z(\SUBBYTES[5].a/w2505 ) );
  NAND U5788 ( .A(\SUBBYTES[5].a/w2484 ), .B(\SUBBYTES[5].a/w2499 ), .Z(n2176)
         );
  AND U5789 ( .A(\SUBBYTES[5].a/w2501 ), .B(\SUBBYTES[5].a/w2507 ), .Z(
        \SUBBYTES[5].a/w2502 ) );
  AND U5790 ( .A(\SUBBYTES[5].a/w2486 ), .B(\SUBBYTES[5].a/w2484 ), .Z(
        \SUBBYTES[5].a/w2496 ) );
  AND U5791 ( .A(\SUBBYTES[5].a/w2487 ), .B(\SUBBYTES[5].a/w2485 ), .Z(
        \SUBBYTES[5].a/w2494 ) );
  AND U5792 ( .A(\SUBBYTES[5].a/w2501 ), .B(\SUBBYTES[5].a/w2508 ), .Z(
        \SUBBYTES[5].a/w2493 ) );
  ANDN U5793 ( .A(\SUBBYTES[5].a/w271 ), .B(n2182), .Z(\SUBBYTES[5].a/w248 )
         );
  AND U5794 ( .A(\SUBBYTES[5].a/w2441 ), .B(\SUBBYTES[5].a/w2437 ), .Z(
        \SUBBYTES[5].a/w2478 ) );
  AND U5795 ( .A(\SUBBYTES[5].a/w2442 ), .B(\SUBBYTES[5].a/w2438 ), .Z(
        \SUBBYTES[5].a/w2476 ) );
  ANDN U5796 ( .A(\SUBBYTES[5].a/w2568 ), .B(n2173), .Z(\SUBBYTES[5].a/w2475 )
         );
  XNOR U5797 ( .A(\w1[5][33] ), .B(\w1[5][39] ), .Z(n2173) );
  XOR U5798 ( .A(\w0[5][33] ), .B(g_input[673]), .Z(\w1[5][33] ) );
  AND U5799 ( .A(\w1[5][32] ), .B(\SUBBYTES[5].a/w2443 ), .Z(
        \SUBBYTES[5].a/w2471 ) );
  XOR U5800 ( .A(\w0[5][32] ), .B(g_input[672]), .Z(\w1[5][32] ) );
  AND U5801 ( .A(\SUBBYTES[5].a/w2444 ), .B(\SUBBYTES[5].a/w2440 ), .Z(
        \SUBBYTES[5].a/w2469 ) );
  AND U5802 ( .A(\SUBBYTES[5].a/w2529 ), .B(\SUBBYTES[5].a/w2561 ), .Z(
        \SUBBYTES[5].a/w2468 ) );
  ANDN U5803 ( .A(\SUBBYTES[5].a/w2550 ), .B(n2179), .Z(\SUBBYTES[5].a/w2463 )
         );
  XNOR U5804 ( .A(\w1[5][36] ), .B(\w1[5][39] ), .Z(n2179) );
  ANDN U5805 ( .A(\SUBBYTES[5].a/w2551 ), .B(n2180), .Z(\SUBBYTES[5].a/w2461 )
         );
  XNOR U5806 ( .A(\w1[5][34] ), .B(\w1[5][39] ), .Z(n2180) );
  XOR U5807 ( .A(\w0[5][39] ), .B(g_input[679]), .Z(\w1[5][39] ) );
  IV U5808 ( .A(n2183), .Z(\w1[5][34] ) );
  ANDN U5809 ( .A(\SUBBYTES[5].a/w2553 ), .B(n2181), .Z(\SUBBYTES[5].a/w2460 )
         );
  XOR U5810 ( .A(n2183), .B(\w1[5][36] ), .Z(n2181) );
  XOR U5811 ( .A(\w0[5][36] ), .B(g_input[676]), .Z(\w1[5][36] ) );
  XNOR U5812 ( .A(\w0[5][34] ), .B(g_input[674]), .Z(n2183) );
  ANDN U5813 ( .A(\SUBBYTES[5].a/w272 ), .B(n2184), .Z(\SUBBYTES[5].a/w246 )
         );
  ANDN U5814 ( .A(\SUBBYTES[5].a/w275 ), .B(n2185), .Z(\SUBBYTES[5].a/w245 )
         );
  AND U5815 ( .A(n2186), .B(\SUBBYTES[5].a/w2230 ), .Z(\SUBBYTES[5].a/w2365 )
         );
  AND U5816 ( .A(n2187), .B(\SUBBYTES[5].a/w2231 ), .Z(\SUBBYTES[5].a/w2363 )
         );
  AND U5817 ( .A(\SUBBYTES[5].a/w2361 ), .B(n2188), .Z(\SUBBYTES[5].a/w2362 )
         );
  ANDN U5818 ( .A(\w1[5][40] ), .B(n2189), .Z(\SUBBYTES[5].a/w2358 ) );
  AND U5819 ( .A(n2190), .B(\SUBBYTES[5].a/w2233 ), .Z(\SUBBYTES[5].a/w2356 )
         );
  AND U5820 ( .A(\SUBBYTES[5].a/w2354 ), .B(n2191), .Z(\SUBBYTES[5].a/w2355 )
         );
  XOR U5821 ( .A(\SUBBYTES[5].a/w2298 ), .B(n10972), .Z(n2191) );
  AND U5822 ( .A(\SUBBYTES[5].a/w2341 ), .B(\SUBBYTES[5].a/w2343 ), .Z(
        \SUBBYTES[5].a/w2350 ) );
  AND U5823 ( .A(\SUBBYTES[5].a/w2342 ), .B(\SUBBYTES[5].a/w2344 ), .Z(
        \SUBBYTES[5].a/w2348 ) );
  AND U5824 ( .A(\SUBBYTES[5].a/w2345 ), .B(\SUBBYTES[5].a/w2346 ), .Z(
        \SUBBYTES[5].a/w2347 ) );
  AND U5825 ( .A(\SUBBYTES[5].a/w2234 ), .B(n2186), .Z(\SUBBYTES[5].a/w2333 )
         );
  XOR U5826 ( .A(\SUBBYTES[5].a/w2302 ), .B(n1031), .Z(n2186) );
  AND U5827 ( .A(\SUBBYTES[5].a/w2235 ), .B(n2187), .Z(\SUBBYTES[5].a/w2331 )
         );
  XOR U5828 ( .A(n10973), .B(\SUBBYTES[5].a/w2302 ), .Z(n2187) );
  ANDN U5829 ( .A(n2188), .B(n2192), .Z(\SUBBYTES[5].a/w2330 ) );
  XOR U5830 ( .A(n1031), .B(n10973), .Z(n2188) );
  ANDN U5831 ( .A(\SUBBYTES[5].a/w2236 ), .B(n2189), .Z(\SUBBYTES[5].a/w2326 )
         );
  XNOR U5832 ( .A(\SUBBYTES[5].a/w2295 ), .B(\SUBBYTES[5].a/w2298 ), .Z(n2189)
         );
  AND U5833 ( .A(\SUBBYTES[5].a/w2237 ), .B(n2190), .Z(\SUBBYTES[5].a/w2324 )
         );
  XNOR U5834 ( .A(n2193), .B(\SUBBYTES[5].a/w2295 ), .Z(n2190) );
  AND U5835 ( .A(\SUBBYTES[5].a/w2322 ), .B(n2194), .Z(\SUBBYTES[5].a/w2323 )
         );
  XOR U5836 ( .A(n2195), .B(n2193), .Z(n2194) );
  IV U5837 ( .A(n10972), .Z(n2193) );
  AND U5838 ( .A(\SUBBYTES[5].a/w231 ), .B(\SUBBYTES[5].a/w230 ), .Z(
        \SUBBYTES[5].a/w232 ) );
  ANDN U5839 ( .A(\SUBBYTES[5].a/w2341 ), .B(n2196), .Z(\SUBBYTES[5].a/w2318 )
         );
  ANDN U5840 ( .A(\SUBBYTES[5].a/w2342 ), .B(n2197), .Z(\SUBBYTES[5].a/w2316 )
         );
  ANDN U5841 ( .A(\SUBBYTES[5].a/w2345 ), .B(n2198), .Z(\SUBBYTES[5].a/w2315 )
         );
  AND U5842 ( .A(\SUBBYTES[5].a/w2301 ), .B(\SUBBYTES[5].a/w2300 ), .Z(
        \SUBBYTES[5].a/w2302 ) );
  IV U5843 ( .A(n2195), .Z(\SUBBYTES[5].a/w2298 ) );
  NAND U5844 ( .A(\SUBBYTES[5].a/w2277 ), .B(\SUBBYTES[5].a/w2292 ), .Z(n2195)
         );
  AND U5845 ( .A(\SUBBYTES[5].a/w2294 ), .B(\SUBBYTES[5].a/w2300 ), .Z(
        \SUBBYTES[5].a/w2295 ) );
  AND U5846 ( .A(\SUBBYTES[5].a/w2279 ), .B(\SUBBYTES[5].a/w2277 ), .Z(
        \SUBBYTES[5].a/w2289 ) );
  AND U5847 ( .A(\SUBBYTES[5].a/w2280 ), .B(\SUBBYTES[5].a/w2278 ), .Z(
        \SUBBYTES[5].a/w2287 ) );
  AND U5848 ( .A(\SUBBYTES[5].a/w2294 ), .B(\SUBBYTES[5].a/w2301 ), .Z(
        \SUBBYTES[5].a/w2286 ) );
  IV U5849 ( .A(n2178), .Z(\SUBBYTES[5].a/w228 ) );
  NAND U5850 ( .A(\SUBBYTES[5].a/w207 ), .B(\SUBBYTES[5].a/w222 ), .Z(n2178)
         );
  AND U5851 ( .A(\SUBBYTES[5].a/w2234 ), .B(\SUBBYTES[5].a/w2230 ), .Z(
        \SUBBYTES[5].a/w2271 ) );
  AND U5852 ( .A(\SUBBYTES[5].a/w2235 ), .B(\SUBBYTES[5].a/w2231 ), .Z(
        \SUBBYTES[5].a/w2269 ) );
  ANDN U5853 ( .A(\SUBBYTES[5].a/w2361 ), .B(n2192), .Z(\SUBBYTES[5].a/w2268 )
         );
  XNOR U5854 ( .A(\w1[5][41] ), .B(\w1[5][47] ), .Z(n2192) );
  XOR U5855 ( .A(\w0[5][41] ), .B(g_input[681]), .Z(\w1[5][41] ) );
  AND U5856 ( .A(\w1[5][40] ), .B(\SUBBYTES[5].a/w2236 ), .Z(
        \SUBBYTES[5].a/w2264 ) );
  XOR U5857 ( .A(\w0[5][40] ), .B(g_input[680]), .Z(\w1[5][40] ) );
  AND U5858 ( .A(\SUBBYTES[5].a/w2237 ), .B(\SUBBYTES[5].a/w2233 ), .Z(
        \SUBBYTES[5].a/w2262 ) );
  AND U5859 ( .A(\SUBBYTES[5].a/w2322 ), .B(\SUBBYTES[5].a/w2354 ), .Z(
        \SUBBYTES[5].a/w2261 ) );
  ANDN U5860 ( .A(\SUBBYTES[5].a/w2343 ), .B(n2196), .Z(\SUBBYTES[5].a/w2256 )
         );
  XNOR U5861 ( .A(\w1[5][44] ), .B(\w1[5][47] ), .Z(n2196) );
  ANDN U5862 ( .A(\SUBBYTES[5].a/w2344 ), .B(n2197), .Z(\SUBBYTES[5].a/w2254 )
         );
  XNOR U5863 ( .A(\w1[5][42] ), .B(\w1[5][47] ), .Z(n2197) );
  XOR U5864 ( .A(\w0[5][47] ), .B(g_input[687]), .Z(\w1[5][47] ) );
  IV U5865 ( .A(n2199), .Z(\w1[5][42] ) );
  ANDN U5866 ( .A(\SUBBYTES[5].a/w2346 ), .B(n2198), .Z(\SUBBYTES[5].a/w2253 )
         );
  XOR U5867 ( .A(n2199), .B(\w1[5][44] ), .Z(n2198) );
  XOR U5868 ( .A(\w0[5][44] ), .B(g_input[684]), .Z(\w1[5][44] ) );
  XNOR U5869 ( .A(\w0[5][42] ), .B(g_input[682]), .Z(n2199) );
  AND U5870 ( .A(\SUBBYTES[5].a/w224 ), .B(\SUBBYTES[5].a/w230 ), .Z(
        \SUBBYTES[5].a/w225 ) );
  AND U5871 ( .A(\SUBBYTES[5].a/w209 ), .B(\SUBBYTES[5].a/w207 ), .Z(
        \SUBBYTES[5].a/w219 ) );
  AND U5872 ( .A(\SUBBYTES[5].a/w210 ), .B(\SUBBYTES[5].a/w208 ), .Z(
        \SUBBYTES[5].a/w217 ) );
  AND U5873 ( .A(\SUBBYTES[5].a/w224 ), .B(\SUBBYTES[5].a/w231 ), .Z(
        \SUBBYTES[5].a/w216 ) );
  AND U5874 ( .A(n2200), .B(\SUBBYTES[5].a/w2023 ), .Z(\SUBBYTES[5].a/w2158 )
         );
  AND U5875 ( .A(n2201), .B(\SUBBYTES[5].a/w2024 ), .Z(\SUBBYTES[5].a/w2156 )
         );
  AND U5876 ( .A(\SUBBYTES[5].a/w2154 ), .B(n2202), .Z(\SUBBYTES[5].a/w2155 )
         );
  ANDN U5877 ( .A(\w1[5][48] ), .B(n2203), .Z(\SUBBYTES[5].a/w2151 ) );
  AND U5878 ( .A(n2204), .B(\SUBBYTES[5].a/w2026 ), .Z(\SUBBYTES[5].a/w2149 )
         );
  AND U5879 ( .A(\SUBBYTES[5].a/w2147 ), .B(n2205), .Z(\SUBBYTES[5].a/w2148 )
         );
  XOR U5880 ( .A(\SUBBYTES[5].a/w2091 ), .B(n10970), .Z(n2205) );
  AND U5881 ( .A(\SUBBYTES[5].a/w2134 ), .B(\SUBBYTES[5].a/w2136 ), .Z(
        \SUBBYTES[5].a/w2143 ) );
  AND U5882 ( .A(\SUBBYTES[5].a/w2135 ), .B(\SUBBYTES[5].a/w2137 ), .Z(
        \SUBBYTES[5].a/w2141 ) );
  AND U5883 ( .A(\SUBBYTES[5].a/w2138 ), .B(\SUBBYTES[5].a/w2139 ), .Z(
        \SUBBYTES[5].a/w2140 ) );
  AND U5884 ( .A(\SUBBYTES[5].a/w2027 ), .B(n2200), .Z(\SUBBYTES[5].a/w2126 )
         );
  XOR U5885 ( .A(\SUBBYTES[5].a/w2095 ), .B(n1030), .Z(n2200) );
  AND U5886 ( .A(\SUBBYTES[5].a/w2028 ), .B(n2201), .Z(\SUBBYTES[5].a/w2124 )
         );
  XOR U5887 ( .A(n10971), .B(\SUBBYTES[5].a/w2095 ), .Z(n2201) );
  ANDN U5888 ( .A(n2202), .B(n2206), .Z(\SUBBYTES[5].a/w2123 ) );
  XOR U5889 ( .A(n1030), .B(n10971), .Z(n2202) );
  ANDN U5890 ( .A(\SUBBYTES[5].a/w2029 ), .B(n2203), .Z(\SUBBYTES[5].a/w2119 )
         );
  XNOR U5891 ( .A(\SUBBYTES[5].a/w2088 ), .B(\SUBBYTES[5].a/w2091 ), .Z(n2203)
         );
  AND U5892 ( .A(\SUBBYTES[5].a/w2030 ), .B(n2204), .Z(\SUBBYTES[5].a/w2117 )
         );
  XNOR U5893 ( .A(n2207), .B(\SUBBYTES[5].a/w2088 ), .Z(n2204) );
  AND U5894 ( .A(\SUBBYTES[5].a/w2115 ), .B(n2208), .Z(\SUBBYTES[5].a/w2116 )
         );
  XOR U5895 ( .A(n2209), .B(n2207), .Z(n2208) );
  IV U5896 ( .A(n10970), .Z(n2207) );
  ANDN U5897 ( .A(\SUBBYTES[5].a/w2134 ), .B(n2210), .Z(\SUBBYTES[5].a/w2111 )
         );
  ANDN U5898 ( .A(\SUBBYTES[5].a/w2135 ), .B(n2211), .Z(\SUBBYTES[5].a/w2109 )
         );
  ANDN U5899 ( .A(\SUBBYTES[5].a/w2138 ), .B(n2212), .Z(\SUBBYTES[5].a/w2108 )
         );
  AND U5900 ( .A(\SUBBYTES[5].a/w2094 ), .B(\SUBBYTES[5].a/w2093 ), .Z(
        \SUBBYTES[5].a/w2095 ) );
  IV U5901 ( .A(n2209), .Z(\SUBBYTES[5].a/w2091 ) );
  NAND U5902 ( .A(\SUBBYTES[5].a/w2070 ), .B(\SUBBYTES[5].a/w2085 ), .Z(n2209)
         );
  AND U5903 ( .A(\SUBBYTES[5].a/w2087 ), .B(\SUBBYTES[5].a/w2093 ), .Z(
        \SUBBYTES[5].a/w2088 ) );
  AND U5904 ( .A(\SUBBYTES[5].a/w2072 ), .B(\SUBBYTES[5].a/w2070 ), .Z(
        \SUBBYTES[5].a/w2082 ) );
  AND U5905 ( .A(\SUBBYTES[5].a/w2073 ), .B(\SUBBYTES[5].a/w2071 ), .Z(
        \SUBBYTES[5].a/w2080 ) );
  AND U5906 ( .A(\SUBBYTES[5].a/w2087 ), .B(\SUBBYTES[5].a/w2094 ), .Z(
        \SUBBYTES[5].a/w2079 ) );
  AND U5907 ( .A(\SUBBYTES[5].a/w2027 ), .B(\SUBBYTES[5].a/w2023 ), .Z(
        \SUBBYTES[5].a/w2064 ) );
  AND U5908 ( .A(\SUBBYTES[5].a/w2028 ), .B(\SUBBYTES[5].a/w2024 ), .Z(
        \SUBBYTES[5].a/w2062 ) );
  ANDN U5909 ( .A(\SUBBYTES[5].a/w2154 ), .B(n2206), .Z(\SUBBYTES[5].a/w2061 )
         );
  XNOR U5910 ( .A(\w1[5][49] ), .B(\w1[5][55] ), .Z(n2206) );
  XOR U5911 ( .A(\w0[5][49] ), .B(g_input[689]), .Z(\w1[5][49] ) );
  AND U5912 ( .A(\w1[5][48] ), .B(\SUBBYTES[5].a/w2029 ), .Z(
        \SUBBYTES[5].a/w2057 ) );
  XOR U5913 ( .A(\w0[5][48] ), .B(g_input[688]), .Z(\w1[5][48] ) );
  AND U5914 ( .A(\SUBBYTES[5].a/w2030 ), .B(\SUBBYTES[5].a/w2026 ), .Z(
        \SUBBYTES[5].a/w2055 ) );
  AND U5915 ( .A(\SUBBYTES[5].a/w2115 ), .B(\SUBBYTES[5].a/w2147 ), .Z(
        \SUBBYTES[5].a/w2054 ) );
  ANDN U5916 ( .A(\SUBBYTES[5].a/w2136 ), .B(n2210), .Z(\SUBBYTES[5].a/w2049 )
         );
  XNOR U5917 ( .A(\w1[5][52] ), .B(\w1[5][55] ), .Z(n2210) );
  ANDN U5918 ( .A(\SUBBYTES[5].a/w2137 ), .B(n2211), .Z(\SUBBYTES[5].a/w2047 )
         );
  XNOR U5919 ( .A(\w1[5][50] ), .B(\w1[5][55] ), .Z(n2211) );
  XOR U5920 ( .A(\w0[5][55] ), .B(g_input[695]), .Z(\w1[5][55] ) );
  IV U5921 ( .A(n2213), .Z(\w1[5][50] ) );
  ANDN U5922 ( .A(\SUBBYTES[5].a/w2139 ), .B(n2212), .Z(\SUBBYTES[5].a/w2046 )
         );
  XOR U5923 ( .A(n2213), .B(\w1[5][52] ), .Z(n2212) );
  XOR U5924 ( .A(\w0[5][52] ), .B(g_input[692]), .Z(\w1[5][52] ) );
  XNOR U5925 ( .A(\w0[5][50] ), .B(g_input[690]), .Z(n2213) );
  AND U5926 ( .A(\SUBBYTES[5].a/w164 ), .B(\SUBBYTES[5].a/w160 ), .Z(
        \SUBBYTES[5].a/w201 ) );
  AND U5927 ( .A(\SUBBYTES[5].a/w165 ), .B(\SUBBYTES[5].a/w161 ), .Z(
        \SUBBYTES[5].a/w199 ) );
  ANDN U5928 ( .A(\SUBBYTES[5].a/w291 ), .B(n2165), .Z(\SUBBYTES[5].a/w198 )
         );
  XNOR U5929 ( .A(\w1[5][121] ), .B(\w1[5][127] ), .Z(n2165) );
  XOR U5930 ( .A(\w0[5][121] ), .B(g_input[761]), .Z(\w1[5][121] ) );
  AND U5931 ( .A(n2214), .B(\SUBBYTES[5].a/w1816 ), .Z(\SUBBYTES[5].a/w1951 )
         );
  AND U5932 ( .A(n2215), .B(\SUBBYTES[5].a/w1817 ), .Z(\SUBBYTES[5].a/w1949 )
         );
  AND U5933 ( .A(\SUBBYTES[5].a/w1947 ), .B(n2216), .Z(\SUBBYTES[5].a/w1948 )
         );
  ANDN U5934 ( .A(\w1[5][56] ), .B(n2217), .Z(\SUBBYTES[5].a/w1944 ) );
  AND U5935 ( .A(n2218), .B(\SUBBYTES[5].a/w1819 ), .Z(\SUBBYTES[5].a/w1942 )
         );
  AND U5936 ( .A(\SUBBYTES[5].a/w1940 ), .B(n2219), .Z(\SUBBYTES[5].a/w1941 )
         );
  XOR U5937 ( .A(\SUBBYTES[5].a/w1884 ), .B(n10968), .Z(n2219) );
  AND U5938 ( .A(\w1[5][120] ), .B(\SUBBYTES[5].a/w166 ), .Z(
        \SUBBYTES[5].a/w194 ) );
  XOR U5939 ( .A(\w0[5][120] ), .B(g_input[760]), .Z(\w1[5][120] ) );
  AND U5940 ( .A(\SUBBYTES[5].a/w1927 ), .B(\SUBBYTES[5].a/w1929 ), .Z(
        \SUBBYTES[5].a/w1936 ) );
  AND U5941 ( .A(\SUBBYTES[5].a/w1928 ), .B(\SUBBYTES[5].a/w1930 ), .Z(
        \SUBBYTES[5].a/w1934 ) );
  AND U5942 ( .A(\SUBBYTES[5].a/w1931 ), .B(\SUBBYTES[5].a/w1932 ), .Z(
        \SUBBYTES[5].a/w1933 ) );
  AND U5943 ( .A(\SUBBYTES[5].a/w167 ), .B(\SUBBYTES[5].a/w163 ), .Z(
        \SUBBYTES[5].a/w192 ) );
  AND U5944 ( .A(\SUBBYTES[5].a/w1820 ), .B(n2214), .Z(\SUBBYTES[5].a/w1919 )
         );
  XOR U5945 ( .A(\SUBBYTES[5].a/w1888 ), .B(n1029), .Z(n2214) );
  AND U5946 ( .A(\SUBBYTES[5].a/w1821 ), .B(n2215), .Z(\SUBBYTES[5].a/w1917 )
         );
  XOR U5947 ( .A(n10969), .B(\SUBBYTES[5].a/w1888 ), .Z(n2215) );
  ANDN U5948 ( .A(n2216), .B(n2220), .Z(\SUBBYTES[5].a/w1916 ) );
  XOR U5949 ( .A(n1029), .B(n10969), .Z(n2216) );
  ANDN U5950 ( .A(\SUBBYTES[5].a/w1822 ), .B(n2217), .Z(\SUBBYTES[5].a/w1912 )
         );
  XNOR U5951 ( .A(\SUBBYTES[5].a/w1881 ), .B(\SUBBYTES[5].a/w1884 ), .Z(n2217)
         );
  AND U5952 ( .A(\SUBBYTES[5].a/w1823 ), .B(n2218), .Z(\SUBBYTES[5].a/w1910 )
         );
  XNOR U5953 ( .A(n2221), .B(\SUBBYTES[5].a/w1881 ), .Z(n2218) );
  AND U5954 ( .A(\SUBBYTES[5].a/w252 ), .B(\SUBBYTES[5].a/w284 ), .Z(
        \SUBBYTES[5].a/w191 ) );
  AND U5955 ( .A(\SUBBYTES[5].a/w1908 ), .B(n2222), .Z(\SUBBYTES[5].a/w1909 )
         );
  XOR U5956 ( .A(n2223), .B(n2221), .Z(n2222) );
  IV U5957 ( .A(n10968), .Z(n2221) );
  ANDN U5958 ( .A(\SUBBYTES[5].a/w1927 ), .B(n2224), .Z(\SUBBYTES[5].a/w1904 )
         );
  ANDN U5959 ( .A(\SUBBYTES[5].a/w1928 ), .B(n2225), .Z(\SUBBYTES[5].a/w1902 )
         );
  ANDN U5960 ( .A(\SUBBYTES[5].a/w1931 ), .B(n2226), .Z(\SUBBYTES[5].a/w1901 )
         );
  AND U5961 ( .A(\SUBBYTES[5].a/w1887 ), .B(\SUBBYTES[5].a/w1886 ), .Z(
        \SUBBYTES[5].a/w1888 ) );
  IV U5962 ( .A(n2223), .Z(\SUBBYTES[5].a/w1884 ) );
  NAND U5963 ( .A(\SUBBYTES[5].a/w1863 ), .B(\SUBBYTES[5].a/w1878 ), .Z(n2223)
         );
  AND U5964 ( .A(\SUBBYTES[5].a/w1880 ), .B(\SUBBYTES[5].a/w1886 ), .Z(
        \SUBBYTES[5].a/w1881 ) );
  AND U5965 ( .A(\SUBBYTES[5].a/w1865 ), .B(\SUBBYTES[5].a/w1863 ), .Z(
        \SUBBYTES[5].a/w1875 ) );
  AND U5966 ( .A(\SUBBYTES[5].a/w1866 ), .B(\SUBBYTES[5].a/w1864 ), .Z(
        \SUBBYTES[5].a/w1873 ) );
  AND U5967 ( .A(\SUBBYTES[5].a/w1880 ), .B(\SUBBYTES[5].a/w1887 ), .Z(
        \SUBBYTES[5].a/w1872 ) );
  ANDN U5968 ( .A(\SUBBYTES[5].a/w273 ), .B(n2182), .Z(\SUBBYTES[5].a/w186 )
         );
  XNOR U5969 ( .A(\w1[5][124] ), .B(\w1[5][127] ), .Z(n2182) );
  AND U5970 ( .A(\SUBBYTES[5].a/w1820 ), .B(\SUBBYTES[5].a/w1816 ), .Z(
        \SUBBYTES[5].a/w1857 ) );
  AND U5971 ( .A(\SUBBYTES[5].a/w1821 ), .B(\SUBBYTES[5].a/w1817 ), .Z(
        \SUBBYTES[5].a/w1855 ) );
  ANDN U5972 ( .A(\SUBBYTES[5].a/w1947 ), .B(n2220), .Z(\SUBBYTES[5].a/w1854 )
         );
  XNOR U5973 ( .A(\w1[5][57] ), .B(\w1[5][63] ), .Z(n2220) );
  XOR U5974 ( .A(\w0[5][57] ), .B(g_input[697]), .Z(\w1[5][57] ) );
  AND U5975 ( .A(\w1[5][56] ), .B(\SUBBYTES[5].a/w1822 ), .Z(
        \SUBBYTES[5].a/w1850 ) );
  XOR U5976 ( .A(\w0[5][56] ), .B(g_input[696]), .Z(\w1[5][56] ) );
  AND U5977 ( .A(\SUBBYTES[5].a/w1823 ), .B(\SUBBYTES[5].a/w1819 ), .Z(
        \SUBBYTES[5].a/w1848 ) );
  AND U5978 ( .A(\SUBBYTES[5].a/w1908 ), .B(\SUBBYTES[5].a/w1940 ), .Z(
        \SUBBYTES[5].a/w1847 ) );
  ANDN U5979 ( .A(\SUBBYTES[5].a/w1929 ), .B(n2224), .Z(\SUBBYTES[5].a/w1842 )
         );
  XNOR U5980 ( .A(\w1[5][60] ), .B(\w1[5][63] ), .Z(n2224) );
  ANDN U5981 ( .A(\SUBBYTES[5].a/w1930 ), .B(n2225), .Z(\SUBBYTES[5].a/w1840 )
         );
  XNOR U5982 ( .A(\w1[5][58] ), .B(\w1[5][63] ), .Z(n2225) );
  XOR U5983 ( .A(\w0[5][63] ), .B(g_input[703]), .Z(\w1[5][63] ) );
  IV U5984 ( .A(n2227), .Z(\w1[5][58] ) );
  ANDN U5985 ( .A(\SUBBYTES[5].a/w274 ), .B(n2184), .Z(\SUBBYTES[5].a/w184 )
         );
  XNOR U5986 ( .A(\w1[5][122] ), .B(\w1[5][127] ), .Z(n2184) );
  XOR U5987 ( .A(\w0[5][127] ), .B(g_input[767]), .Z(\w1[5][127] ) );
  IV U5988 ( .A(n2228), .Z(\w1[5][122] ) );
  ANDN U5989 ( .A(\SUBBYTES[5].a/w1932 ), .B(n2226), .Z(\SUBBYTES[5].a/w1839 )
         );
  XOR U5990 ( .A(n2227), .B(\w1[5][60] ), .Z(n2226) );
  XOR U5991 ( .A(\w0[5][60] ), .B(g_input[700]), .Z(\w1[5][60] ) );
  XNOR U5992 ( .A(\w0[5][58] ), .B(g_input[698]), .Z(n2227) );
  ANDN U5993 ( .A(\SUBBYTES[5].a/w276 ), .B(n2185), .Z(\SUBBYTES[5].a/w183 )
         );
  XOR U5994 ( .A(n2228), .B(\w1[5][124] ), .Z(n2185) );
  XOR U5995 ( .A(\w0[5][124] ), .B(g_input[764]), .Z(\w1[5][124] ) );
  XNOR U5996 ( .A(\w0[5][122] ), .B(g_input[762]), .Z(n2228) );
  AND U5997 ( .A(n2229), .B(\SUBBYTES[5].a/w1609 ), .Z(\SUBBYTES[5].a/w1744 )
         );
  AND U5998 ( .A(n2230), .B(\SUBBYTES[5].a/w1610 ), .Z(\SUBBYTES[5].a/w1742 )
         );
  AND U5999 ( .A(\SUBBYTES[5].a/w1740 ), .B(n2231), .Z(\SUBBYTES[5].a/w1741 )
         );
  ANDN U6000 ( .A(\w1[5][64] ), .B(n2232), .Z(\SUBBYTES[5].a/w1737 ) );
  AND U6001 ( .A(n2233), .B(\SUBBYTES[5].a/w1612 ), .Z(\SUBBYTES[5].a/w1735 )
         );
  AND U6002 ( .A(\SUBBYTES[5].a/w1733 ), .B(n2234), .Z(\SUBBYTES[5].a/w1734 )
         );
  XOR U6003 ( .A(\SUBBYTES[5].a/w1677 ), .B(n10966), .Z(n2234) );
  AND U6004 ( .A(\SUBBYTES[5].a/w1720 ), .B(\SUBBYTES[5].a/w1722 ), .Z(
        \SUBBYTES[5].a/w1729 ) );
  AND U6005 ( .A(\SUBBYTES[5].a/w1721 ), .B(\SUBBYTES[5].a/w1723 ), .Z(
        \SUBBYTES[5].a/w1727 ) );
  AND U6006 ( .A(\SUBBYTES[5].a/w1724 ), .B(\SUBBYTES[5].a/w1725 ), .Z(
        \SUBBYTES[5].a/w1726 ) );
  AND U6007 ( .A(\SUBBYTES[5].a/w1613 ), .B(n2229), .Z(\SUBBYTES[5].a/w1712 )
         );
  XOR U6008 ( .A(\SUBBYTES[5].a/w1681 ), .B(n1028), .Z(n2229) );
  AND U6009 ( .A(\SUBBYTES[5].a/w1614 ), .B(n2230), .Z(\SUBBYTES[5].a/w1710 )
         );
  XOR U6010 ( .A(n10967), .B(\SUBBYTES[5].a/w1681 ), .Z(n2230) );
  ANDN U6011 ( .A(n2231), .B(n2235), .Z(\SUBBYTES[5].a/w1709 ) );
  XOR U6012 ( .A(n1028), .B(n10967), .Z(n2231) );
  ANDN U6013 ( .A(\SUBBYTES[5].a/w1615 ), .B(n2232), .Z(\SUBBYTES[5].a/w1705 )
         );
  XNOR U6014 ( .A(\SUBBYTES[5].a/w1674 ), .B(\SUBBYTES[5].a/w1677 ), .Z(n2232)
         );
  AND U6015 ( .A(\SUBBYTES[5].a/w1616 ), .B(n2233), .Z(\SUBBYTES[5].a/w1703 )
         );
  XNOR U6016 ( .A(n2236), .B(\SUBBYTES[5].a/w1674 ), .Z(n2233) );
  AND U6017 ( .A(\SUBBYTES[5].a/w1701 ), .B(n2237), .Z(\SUBBYTES[5].a/w1702 )
         );
  XOR U6018 ( .A(n2238), .B(n2236), .Z(n2237) );
  IV U6019 ( .A(n10966), .Z(n2236) );
  ANDN U6020 ( .A(\SUBBYTES[5].a/w1720 ), .B(n2239), .Z(\SUBBYTES[5].a/w1697 )
         );
  ANDN U6021 ( .A(\SUBBYTES[5].a/w1721 ), .B(n2240), .Z(\SUBBYTES[5].a/w1695 )
         );
  ANDN U6022 ( .A(\SUBBYTES[5].a/w1724 ), .B(n2241), .Z(\SUBBYTES[5].a/w1694 )
         );
  AND U6023 ( .A(\SUBBYTES[5].a/w1680 ), .B(\SUBBYTES[5].a/w1679 ), .Z(
        \SUBBYTES[5].a/w1681 ) );
  IV U6024 ( .A(n2238), .Z(\SUBBYTES[5].a/w1677 ) );
  NAND U6025 ( .A(\SUBBYTES[5].a/w1656 ), .B(\SUBBYTES[5].a/w1671 ), .Z(n2238)
         );
  AND U6026 ( .A(\SUBBYTES[5].a/w1673 ), .B(\SUBBYTES[5].a/w1679 ), .Z(
        \SUBBYTES[5].a/w1674 ) );
  AND U6027 ( .A(\SUBBYTES[5].a/w1658 ), .B(\SUBBYTES[5].a/w1656 ), .Z(
        \SUBBYTES[5].a/w1668 ) );
  AND U6028 ( .A(\SUBBYTES[5].a/w1659 ), .B(\SUBBYTES[5].a/w1657 ), .Z(
        \SUBBYTES[5].a/w1666 ) );
  AND U6029 ( .A(\SUBBYTES[5].a/w1673 ), .B(\SUBBYTES[5].a/w1680 ), .Z(
        \SUBBYTES[5].a/w1665 ) );
  AND U6030 ( .A(\SUBBYTES[5].a/w1613 ), .B(\SUBBYTES[5].a/w1609 ), .Z(
        \SUBBYTES[5].a/w1650 ) );
  AND U6031 ( .A(\SUBBYTES[5].a/w1614 ), .B(\SUBBYTES[5].a/w1610 ), .Z(
        \SUBBYTES[5].a/w1648 ) );
  ANDN U6032 ( .A(\SUBBYTES[5].a/w1740 ), .B(n2235), .Z(\SUBBYTES[5].a/w1647 )
         );
  XNOR U6033 ( .A(\w1[5][65] ), .B(\w1[5][71] ), .Z(n2235) );
  XOR U6034 ( .A(\w0[5][65] ), .B(g_input[705]), .Z(\w1[5][65] ) );
  AND U6035 ( .A(\w1[5][64] ), .B(\SUBBYTES[5].a/w1615 ), .Z(
        \SUBBYTES[5].a/w1643 ) );
  XOR U6036 ( .A(\w0[5][64] ), .B(g_input[704]), .Z(\w1[5][64] ) );
  AND U6037 ( .A(\SUBBYTES[5].a/w1616 ), .B(\SUBBYTES[5].a/w1612 ), .Z(
        \SUBBYTES[5].a/w1641 ) );
  AND U6038 ( .A(\SUBBYTES[5].a/w1701 ), .B(\SUBBYTES[5].a/w1733 ), .Z(
        \SUBBYTES[5].a/w1640 ) );
  ANDN U6039 ( .A(\SUBBYTES[5].a/w1722 ), .B(n2239), .Z(\SUBBYTES[5].a/w1635 )
         );
  XNOR U6040 ( .A(\w1[5][68] ), .B(\w1[5][71] ), .Z(n2239) );
  ANDN U6041 ( .A(\SUBBYTES[5].a/w1723 ), .B(n2240), .Z(\SUBBYTES[5].a/w1633 )
         );
  XNOR U6042 ( .A(\w1[5][66] ), .B(\w1[5][71] ), .Z(n2240) );
  XOR U6043 ( .A(\w0[5][71] ), .B(g_input[711]), .Z(\w1[5][71] ) );
  IV U6044 ( .A(n2242), .Z(\w1[5][66] ) );
  ANDN U6045 ( .A(\SUBBYTES[5].a/w1725 ), .B(n2241), .Z(\SUBBYTES[5].a/w1632 )
         );
  XOR U6046 ( .A(n2242), .B(\w1[5][68] ), .Z(n2241) );
  XOR U6047 ( .A(\w0[5][68] ), .B(g_input[708]), .Z(\w1[5][68] ) );
  XNOR U6048 ( .A(\w0[5][66] ), .B(g_input[706]), .Z(n2242) );
  AND U6049 ( .A(n2243), .B(\SUBBYTES[5].a/w1402 ), .Z(\SUBBYTES[5].a/w1537 )
         );
  AND U6050 ( .A(n2244), .B(\SUBBYTES[5].a/w1403 ), .Z(\SUBBYTES[5].a/w1535 )
         );
  AND U6051 ( .A(\SUBBYTES[5].a/w1533 ), .B(n2245), .Z(\SUBBYTES[5].a/w1534 )
         );
  ANDN U6052 ( .A(\w1[5][72] ), .B(n2246), .Z(\SUBBYTES[5].a/w1530 ) );
  AND U6053 ( .A(n2247), .B(\SUBBYTES[5].a/w1405 ), .Z(\SUBBYTES[5].a/w1528 )
         );
  AND U6054 ( .A(\SUBBYTES[5].a/w1526 ), .B(n2248), .Z(\SUBBYTES[5].a/w1527 )
         );
  XOR U6055 ( .A(\SUBBYTES[5].a/w1470 ), .B(n10964), .Z(n2248) );
  AND U6056 ( .A(\SUBBYTES[5].a/w1513 ), .B(\SUBBYTES[5].a/w1515 ), .Z(
        \SUBBYTES[5].a/w1522 ) );
  AND U6057 ( .A(\SUBBYTES[5].a/w1514 ), .B(\SUBBYTES[5].a/w1516 ), .Z(
        \SUBBYTES[5].a/w1520 ) );
  AND U6058 ( .A(\SUBBYTES[5].a/w1517 ), .B(\SUBBYTES[5].a/w1518 ), .Z(
        \SUBBYTES[5].a/w1519 ) );
  AND U6059 ( .A(\SUBBYTES[5].a/w1406 ), .B(n2243), .Z(\SUBBYTES[5].a/w1505 )
         );
  XOR U6060 ( .A(\SUBBYTES[5].a/w1474 ), .B(n1027), .Z(n2243) );
  AND U6061 ( .A(\SUBBYTES[5].a/w1407 ), .B(n2244), .Z(\SUBBYTES[5].a/w1503 )
         );
  XOR U6062 ( .A(n10965), .B(\SUBBYTES[5].a/w1474 ), .Z(n2244) );
  ANDN U6063 ( .A(n2245), .B(n2249), .Z(\SUBBYTES[5].a/w1502 ) );
  XOR U6064 ( .A(n1027), .B(n10965), .Z(n2245) );
  ANDN U6065 ( .A(\SUBBYTES[5].a/w1408 ), .B(n2246), .Z(\SUBBYTES[5].a/w1498 )
         );
  XNOR U6066 ( .A(\SUBBYTES[5].a/w1467 ), .B(\SUBBYTES[5].a/w1470 ), .Z(n2246)
         );
  AND U6067 ( .A(\SUBBYTES[5].a/w1409 ), .B(n2247), .Z(\SUBBYTES[5].a/w1496 )
         );
  XNOR U6068 ( .A(n2250), .B(\SUBBYTES[5].a/w1467 ), .Z(n2247) );
  AND U6069 ( .A(\SUBBYTES[5].a/w1494 ), .B(n2251), .Z(\SUBBYTES[5].a/w1495 )
         );
  XOR U6070 ( .A(n2252), .B(n2250), .Z(n2251) );
  IV U6071 ( .A(n10964), .Z(n2250) );
  ANDN U6072 ( .A(\SUBBYTES[5].a/w1513 ), .B(n2253), .Z(\SUBBYTES[5].a/w1490 )
         );
  ANDN U6073 ( .A(\SUBBYTES[5].a/w1514 ), .B(n2254), .Z(\SUBBYTES[5].a/w1488 )
         );
  ANDN U6074 ( .A(\SUBBYTES[5].a/w1517 ), .B(n2255), .Z(\SUBBYTES[5].a/w1487 )
         );
  AND U6075 ( .A(\SUBBYTES[5].a/w1473 ), .B(\SUBBYTES[5].a/w1472 ), .Z(
        \SUBBYTES[5].a/w1474 ) );
  IV U6076 ( .A(n2252), .Z(\SUBBYTES[5].a/w1470 ) );
  NAND U6077 ( .A(\SUBBYTES[5].a/w1449 ), .B(\SUBBYTES[5].a/w1464 ), .Z(n2252)
         );
  AND U6078 ( .A(\SUBBYTES[5].a/w1466 ), .B(\SUBBYTES[5].a/w1472 ), .Z(
        \SUBBYTES[5].a/w1467 ) );
  AND U6079 ( .A(\SUBBYTES[5].a/w1451 ), .B(\SUBBYTES[5].a/w1449 ), .Z(
        \SUBBYTES[5].a/w1461 ) );
  AND U6080 ( .A(\SUBBYTES[5].a/w1452 ), .B(\SUBBYTES[5].a/w1450 ), .Z(
        \SUBBYTES[5].a/w1459 ) );
  AND U6081 ( .A(\SUBBYTES[5].a/w1466 ), .B(\SUBBYTES[5].a/w1473 ), .Z(
        \SUBBYTES[5].a/w1458 ) );
  AND U6082 ( .A(\SUBBYTES[5].a/w1406 ), .B(\SUBBYTES[5].a/w1402 ), .Z(
        \SUBBYTES[5].a/w1443 ) );
  AND U6083 ( .A(\SUBBYTES[5].a/w1407 ), .B(\SUBBYTES[5].a/w1403 ), .Z(
        \SUBBYTES[5].a/w1441 ) );
  ANDN U6084 ( .A(\SUBBYTES[5].a/w1533 ), .B(n2249), .Z(\SUBBYTES[5].a/w1440 )
         );
  XNOR U6085 ( .A(\w1[5][73] ), .B(\w1[5][79] ), .Z(n2249) );
  XOR U6086 ( .A(\w0[5][73] ), .B(g_input[713]), .Z(\w1[5][73] ) );
  AND U6087 ( .A(\w1[5][72] ), .B(\SUBBYTES[5].a/w1408 ), .Z(
        \SUBBYTES[5].a/w1436 ) );
  XOR U6088 ( .A(\w0[5][72] ), .B(g_input[712]), .Z(\w1[5][72] ) );
  AND U6089 ( .A(\SUBBYTES[5].a/w1409 ), .B(\SUBBYTES[5].a/w1405 ), .Z(
        \SUBBYTES[5].a/w1434 ) );
  AND U6090 ( .A(\SUBBYTES[5].a/w1494 ), .B(\SUBBYTES[5].a/w1526 ), .Z(
        \SUBBYTES[5].a/w1433 ) );
  ANDN U6091 ( .A(\SUBBYTES[5].a/w1515 ), .B(n2253), .Z(\SUBBYTES[5].a/w1428 )
         );
  XNOR U6092 ( .A(\w1[5][76] ), .B(\w1[5][79] ), .Z(n2253) );
  ANDN U6093 ( .A(\SUBBYTES[5].a/w1516 ), .B(n2254), .Z(\SUBBYTES[5].a/w1426 )
         );
  XNOR U6094 ( .A(\w1[5][74] ), .B(\w1[5][79] ), .Z(n2254) );
  XOR U6095 ( .A(\w0[5][79] ), .B(g_input[719]), .Z(\w1[5][79] ) );
  IV U6096 ( .A(n2256), .Z(\w1[5][74] ) );
  ANDN U6097 ( .A(\SUBBYTES[5].a/w1518 ), .B(n2255), .Z(\SUBBYTES[5].a/w1425 )
         );
  XOR U6098 ( .A(n2256), .B(\w1[5][76] ), .Z(n2255) );
  XOR U6099 ( .A(\w0[5][76] ), .B(g_input[716]), .Z(\w1[5][76] ) );
  XNOR U6100 ( .A(\w0[5][74] ), .B(g_input[714]), .Z(n2256) );
  AND U6101 ( .A(n2257), .B(\SUBBYTES[5].a/w1195 ), .Z(\SUBBYTES[5].a/w1330 )
         );
  AND U6102 ( .A(n2258), .B(\SUBBYTES[5].a/w1196 ), .Z(\SUBBYTES[5].a/w1328 )
         );
  AND U6103 ( .A(\SUBBYTES[5].a/w1326 ), .B(n2259), .Z(\SUBBYTES[5].a/w1327 )
         );
  ANDN U6104 ( .A(\w1[5][80] ), .B(n2260), .Z(\SUBBYTES[5].a/w1323 ) );
  AND U6105 ( .A(n2261), .B(\SUBBYTES[5].a/w1198 ), .Z(\SUBBYTES[5].a/w1321 )
         );
  AND U6106 ( .A(\SUBBYTES[5].a/w1319 ), .B(n2262), .Z(\SUBBYTES[5].a/w1320 )
         );
  XOR U6107 ( .A(\SUBBYTES[5].a/w1263 ), .B(n10962), .Z(n2262) );
  AND U6108 ( .A(\SUBBYTES[5].a/w1306 ), .B(\SUBBYTES[5].a/w1308 ), .Z(
        \SUBBYTES[5].a/w1315 ) );
  AND U6109 ( .A(\SUBBYTES[5].a/w1307 ), .B(\SUBBYTES[5].a/w1309 ), .Z(
        \SUBBYTES[5].a/w1313 ) );
  AND U6110 ( .A(\SUBBYTES[5].a/w1310 ), .B(\SUBBYTES[5].a/w1311 ), .Z(
        \SUBBYTES[5].a/w1312 ) );
  AND U6111 ( .A(\SUBBYTES[5].a/w1199 ), .B(n2257), .Z(\SUBBYTES[5].a/w1298 )
         );
  XOR U6112 ( .A(\SUBBYTES[5].a/w1267 ), .B(n1026), .Z(n2257) );
  AND U6113 ( .A(\SUBBYTES[5].a/w1200 ), .B(n2258), .Z(\SUBBYTES[5].a/w1296 )
         );
  XOR U6114 ( .A(n10963), .B(\SUBBYTES[5].a/w1267 ), .Z(n2258) );
  ANDN U6115 ( .A(n2259), .B(n2263), .Z(\SUBBYTES[5].a/w1295 ) );
  XOR U6116 ( .A(n1026), .B(n10963), .Z(n2259) );
  ANDN U6117 ( .A(\SUBBYTES[5].a/w1201 ), .B(n2260), .Z(\SUBBYTES[5].a/w1291 )
         );
  XNOR U6118 ( .A(\SUBBYTES[5].a/w1260 ), .B(\SUBBYTES[5].a/w1263 ), .Z(n2260)
         );
  AND U6119 ( .A(\SUBBYTES[5].a/w1202 ), .B(n2261), .Z(\SUBBYTES[5].a/w1289 )
         );
  XNOR U6120 ( .A(n2264), .B(\SUBBYTES[5].a/w1260 ), .Z(n2261) );
  AND U6121 ( .A(\SUBBYTES[5].a/w1287 ), .B(n2265), .Z(\SUBBYTES[5].a/w1288 )
         );
  XOR U6122 ( .A(n2266), .B(n2264), .Z(n2265) );
  IV U6123 ( .A(n10962), .Z(n2264) );
  ANDN U6124 ( .A(\SUBBYTES[5].a/w1306 ), .B(n2267), .Z(\SUBBYTES[5].a/w1283 )
         );
  ANDN U6125 ( .A(\SUBBYTES[5].a/w1307 ), .B(n2268), .Z(\SUBBYTES[5].a/w1281 )
         );
  ANDN U6126 ( .A(\SUBBYTES[5].a/w1310 ), .B(n2269), .Z(\SUBBYTES[5].a/w1280 )
         );
  AND U6127 ( .A(\SUBBYTES[5].a/w1266 ), .B(\SUBBYTES[5].a/w1265 ), .Z(
        \SUBBYTES[5].a/w1267 ) );
  IV U6128 ( .A(n2266), .Z(\SUBBYTES[5].a/w1263 ) );
  NAND U6129 ( .A(\SUBBYTES[5].a/w1242 ), .B(\SUBBYTES[5].a/w1257 ), .Z(n2266)
         );
  AND U6130 ( .A(\SUBBYTES[5].a/w1259 ), .B(\SUBBYTES[5].a/w1265 ), .Z(
        \SUBBYTES[5].a/w1260 ) );
  AND U6131 ( .A(\SUBBYTES[5].a/w1244 ), .B(\SUBBYTES[5].a/w1242 ), .Z(
        \SUBBYTES[5].a/w1254 ) );
  AND U6132 ( .A(\SUBBYTES[5].a/w1245 ), .B(\SUBBYTES[5].a/w1243 ), .Z(
        \SUBBYTES[5].a/w1252 ) );
  AND U6133 ( .A(\SUBBYTES[5].a/w1259 ), .B(\SUBBYTES[5].a/w1266 ), .Z(
        \SUBBYTES[5].a/w1251 ) );
  AND U6134 ( .A(\SUBBYTES[5].a/w1199 ), .B(\SUBBYTES[5].a/w1195 ), .Z(
        \SUBBYTES[5].a/w1236 ) );
  AND U6135 ( .A(\SUBBYTES[5].a/w1200 ), .B(\SUBBYTES[5].a/w1196 ), .Z(
        \SUBBYTES[5].a/w1234 ) );
  ANDN U6136 ( .A(\SUBBYTES[5].a/w1326 ), .B(n2263), .Z(\SUBBYTES[5].a/w1233 )
         );
  XNOR U6137 ( .A(\w1[5][81] ), .B(\w1[5][87] ), .Z(n2263) );
  XOR U6138 ( .A(\w0[5][81] ), .B(g_input[721]), .Z(\w1[5][81] ) );
  AND U6139 ( .A(\w1[5][80] ), .B(\SUBBYTES[5].a/w1201 ), .Z(
        \SUBBYTES[5].a/w1229 ) );
  XOR U6140 ( .A(\w0[5][80] ), .B(g_input[720]), .Z(\w1[5][80] ) );
  AND U6141 ( .A(\SUBBYTES[5].a/w1202 ), .B(\SUBBYTES[5].a/w1198 ), .Z(
        \SUBBYTES[5].a/w1227 ) );
  AND U6142 ( .A(\SUBBYTES[5].a/w1287 ), .B(\SUBBYTES[5].a/w1319 ), .Z(
        \SUBBYTES[5].a/w1226 ) );
  ANDN U6143 ( .A(\SUBBYTES[5].a/w1308 ), .B(n2267), .Z(\SUBBYTES[5].a/w1221 )
         );
  XNOR U6144 ( .A(\w1[5][84] ), .B(\w1[5][87] ), .Z(n2267) );
  ANDN U6145 ( .A(\SUBBYTES[5].a/w1309 ), .B(n2268), .Z(\SUBBYTES[5].a/w1219 )
         );
  XNOR U6146 ( .A(\w1[5][82] ), .B(\w1[5][87] ), .Z(n2268) );
  XOR U6147 ( .A(\w0[5][87] ), .B(g_input[727]), .Z(\w1[5][87] ) );
  IV U6148 ( .A(n2270), .Z(\w1[5][82] ) );
  ANDN U6149 ( .A(\SUBBYTES[5].a/w1311 ), .B(n2269), .Z(\SUBBYTES[5].a/w1218 )
         );
  XOR U6150 ( .A(n2270), .B(\w1[5][84] ), .Z(n2269) );
  XOR U6151 ( .A(\w0[5][84] ), .B(g_input[724]), .Z(\w1[5][84] ) );
  XNOR U6152 ( .A(\w0[5][82] ), .B(g_input[722]), .Z(n2270) );
  AND U6153 ( .A(n2271), .B(\SUBBYTES[5].a/w988 ), .Z(\SUBBYTES[5].a/w1123 )
         );
  AND U6154 ( .A(n2272), .B(\SUBBYTES[5].a/w989 ), .Z(\SUBBYTES[5].a/w1121 )
         );
  AND U6155 ( .A(\SUBBYTES[5].a/w1119 ), .B(n2273), .Z(\SUBBYTES[5].a/w1120 )
         );
  ANDN U6156 ( .A(\w1[5][88] ), .B(n2274), .Z(\SUBBYTES[5].a/w1116 ) );
  AND U6157 ( .A(n2275), .B(\SUBBYTES[5].a/w991 ), .Z(\SUBBYTES[5].a/w1114 )
         );
  AND U6158 ( .A(\SUBBYTES[5].a/w1112 ), .B(n2276), .Z(\SUBBYTES[5].a/w1113 )
         );
  XOR U6159 ( .A(\SUBBYTES[5].a/w1056 ), .B(n10960), .Z(n2276) );
  AND U6160 ( .A(\SUBBYTES[5].a/w1099 ), .B(\SUBBYTES[5].a/w1101 ), .Z(
        \SUBBYTES[5].a/w1108 ) );
  AND U6161 ( .A(\SUBBYTES[5].a/w1100 ), .B(\SUBBYTES[5].a/w1102 ), .Z(
        \SUBBYTES[5].a/w1106 ) );
  AND U6162 ( .A(\SUBBYTES[5].a/w1103 ), .B(\SUBBYTES[5].a/w1104 ), .Z(
        \SUBBYTES[5].a/w1105 ) );
  AND U6163 ( .A(\SUBBYTES[5].a/w992 ), .B(n2271), .Z(\SUBBYTES[5].a/w1091 )
         );
  XOR U6164 ( .A(\SUBBYTES[5].a/w1060 ), .B(n1025), .Z(n2271) );
  AND U6165 ( .A(\SUBBYTES[5].a/w993 ), .B(n2272), .Z(\SUBBYTES[5].a/w1089 )
         );
  XOR U6166 ( .A(n10961), .B(\SUBBYTES[5].a/w1060 ), .Z(n2272) );
  ANDN U6167 ( .A(n2273), .B(n2277), .Z(\SUBBYTES[5].a/w1088 ) );
  XOR U6168 ( .A(n1025), .B(n10961), .Z(n2273) );
  ANDN U6169 ( .A(\SUBBYTES[5].a/w994 ), .B(n2274), .Z(\SUBBYTES[5].a/w1084 )
         );
  XNOR U6170 ( .A(\SUBBYTES[5].a/w1053 ), .B(\SUBBYTES[5].a/w1056 ), .Z(n2274)
         );
  AND U6171 ( .A(\SUBBYTES[5].a/w995 ), .B(n2275), .Z(\SUBBYTES[5].a/w1082 )
         );
  XNOR U6172 ( .A(n2278), .B(\SUBBYTES[5].a/w1053 ), .Z(n2275) );
  AND U6173 ( .A(\SUBBYTES[5].a/w1080 ), .B(n2279), .Z(\SUBBYTES[5].a/w1081 )
         );
  XOR U6174 ( .A(n2280), .B(n2278), .Z(n2279) );
  IV U6175 ( .A(n10960), .Z(n2278) );
  ANDN U6176 ( .A(\SUBBYTES[5].a/w1099 ), .B(n2281), .Z(\SUBBYTES[5].a/w1076 )
         );
  ANDN U6177 ( .A(\SUBBYTES[5].a/w1100 ), .B(n2282), .Z(\SUBBYTES[5].a/w1074 )
         );
  ANDN U6178 ( .A(\SUBBYTES[5].a/w1103 ), .B(n2283), .Z(\SUBBYTES[5].a/w1073 )
         );
  AND U6179 ( .A(\SUBBYTES[5].a/w1059 ), .B(\SUBBYTES[5].a/w1058 ), .Z(
        \SUBBYTES[5].a/w1060 ) );
  IV U6180 ( .A(n2280), .Z(\SUBBYTES[5].a/w1056 ) );
  NAND U6181 ( .A(\SUBBYTES[5].a/w1035 ), .B(\SUBBYTES[5].a/w1050 ), .Z(n2280)
         );
  AND U6182 ( .A(\SUBBYTES[5].a/w1052 ), .B(\SUBBYTES[5].a/w1058 ), .Z(
        \SUBBYTES[5].a/w1053 ) );
  AND U6183 ( .A(\SUBBYTES[5].a/w1037 ), .B(\SUBBYTES[5].a/w1035 ), .Z(
        \SUBBYTES[5].a/w1047 ) );
  AND U6184 ( .A(\SUBBYTES[5].a/w1038 ), .B(\SUBBYTES[5].a/w1036 ), .Z(
        \SUBBYTES[5].a/w1045 ) );
  AND U6185 ( .A(\SUBBYTES[5].a/w1052 ), .B(\SUBBYTES[5].a/w1059 ), .Z(
        \SUBBYTES[5].a/w1044 ) );
  AND U6186 ( .A(\SUBBYTES[5].a/w992 ), .B(\SUBBYTES[5].a/w988 ), .Z(
        \SUBBYTES[5].a/w1029 ) );
  AND U6187 ( .A(\SUBBYTES[5].a/w993 ), .B(\SUBBYTES[5].a/w989 ), .Z(
        \SUBBYTES[5].a/w1027 ) );
  ANDN U6188 ( .A(\SUBBYTES[5].a/w1119 ), .B(n2277), .Z(\SUBBYTES[5].a/w1026 )
         );
  XNOR U6189 ( .A(\w1[5][89] ), .B(\w1[5][95] ), .Z(n2277) );
  XOR U6190 ( .A(\w0[5][89] ), .B(g_input[729]), .Z(\w1[5][89] ) );
  AND U6191 ( .A(\w1[5][88] ), .B(\SUBBYTES[5].a/w994 ), .Z(
        \SUBBYTES[5].a/w1022 ) );
  XOR U6192 ( .A(\w0[5][88] ), .B(g_input[728]), .Z(\w1[5][88] ) );
  AND U6193 ( .A(\SUBBYTES[5].a/w995 ), .B(\SUBBYTES[5].a/w991 ), .Z(
        \SUBBYTES[5].a/w1020 ) );
  AND U6194 ( .A(\SUBBYTES[5].a/w1080 ), .B(\SUBBYTES[5].a/w1112 ), .Z(
        \SUBBYTES[5].a/w1019 ) );
  ANDN U6195 ( .A(\SUBBYTES[5].a/w1101 ), .B(n2281), .Z(\SUBBYTES[5].a/w1014 )
         );
  XNOR U6196 ( .A(\w1[5][92] ), .B(\w1[5][95] ), .Z(n2281) );
  ANDN U6197 ( .A(\SUBBYTES[5].a/w1102 ), .B(n2282), .Z(\SUBBYTES[5].a/w1012 )
         );
  XNOR U6198 ( .A(\w1[5][90] ), .B(\w1[5][95] ), .Z(n2282) );
  XOR U6199 ( .A(\w0[5][95] ), .B(g_input[735]), .Z(\w1[5][95] ) );
  IV U6200 ( .A(n2284), .Z(\w1[5][90] ) );
  ANDN U6201 ( .A(\SUBBYTES[5].a/w1104 ), .B(n2283), .Z(\SUBBYTES[5].a/w1011 )
         );
  XOR U6202 ( .A(n2284), .B(\w1[5][92] ), .Z(n2283) );
  XOR U6203 ( .A(\w0[5][92] ), .B(g_input[732]), .Z(\w1[5][92] ) );
  XNOR U6204 ( .A(\w0[5][90] ), .B(g_input[730]), .Z(n2284) );
  AND U6205 ( .A(\SUBBYTES[5].a/w2084 ), .B(\SUBBYTES[5].a/w2071 ), .Z(n10970)
         );
  AND U6206 ( .A(\SUBBYTES[5].a/w1877 ), .B(\SUBBYTES[5].a/w1866 ), .Z(n10969)
         );
  AND U6207 ( .A(\SUBBYTES[5].a/w221 ), .B(\SUBBYTES[5].a/w208 ), .Z(n10952)
         );
  AND U6208 ( .A(\SUBBYTES[5].a/w1877 ), .B(\SUBBYTES[5].a/w1864 ), .Z(n10968)
         );
  AND U6209 ( .A(\SUBBYTES[5].a/w1670 ), .B(\SUBBYTES[5].a/w1659 ), .Z(n10967)
         );
  AND U6210 ( .A(\SUBBYTES[5].a/w1670 ), .B(\SUBBYTES[5].a/w1657 ), .Z(n10966)
         );
  AND U6211 ( .A(\SUBBYTES[5].a/w1463 ), .B(\SUBBYTES[5].a/w1452 ), .Z(n10965)
         );
  AND U6212 ( .A(\SUBBYTES[5].a/w1463 ), .B(\SUBBYTES[5].a/w1450 ), .Z(n10964)
         );
  AND U6213 ( .A(\SUBBYTES[5].a/w1256 ), .B(\SUBBYTES[5].a/w1245 ), .Z(n10963)
         );
  AND U6214 ( .A(\SUBBYTES[5].a/w1256 ), .B(\SUBBYTES[5].a/w1243 ), .Z(n10962)
         );
  AND U6215 ( .A(\SUBBYTES[5].a/w1049 ), .B(\SUBBYTES[5].a/w1038 ), .Z(n10961)
         );
  AND U6216 ( .A(\SUBBYTES[5].a/w1049 ), .B(\SUBBYTES[5].a/w1036 ), .Z(n10960)
         );
  AND U6217 ( .A(\SUBBYTES[5].a/w842 ), .B(\SUBBYTES[5].a/w831 ), .Z(n10959)
         );
  AND U6218 ( .A(\SUBBYTES[5].a/w842 ), .B(\SUBBYTES[5].a/w829 ), .Z(n10958)
         );
  AND U6219 ( .A(\SUBBYTES[5].a/w635 ), .B(\SUBBYTES[5].a/w624 ), .Z(n10957)
         );
  AND U6220 ( .A(\SUBBYTES[5].a/w635 ), .B(\SUBBYTES[5].a/w622 ), .Z(n10956)
         );
  AND U6221 ( .A(\SUBBYTES[5].a/w428 ), .B(\SUBBYTES[5].a/w417 ), .Z(n10955)
         );
  AND U6222 ( .A(\SUBBYTES[5].a/w428 ), .B(\SUBBYTES[5].a/w415 ), .Z(n10954)
         );
  AND U6223 ( .A(\SUBBYTES[5].a/w3326 ), .B(\SUBBYTES[5].a/w3315 ), .Z(n10983)
         );
  AND U6224 ( .A(\SUBBYTES[5].a/w3326 ), .B(\SUBBYTES[5].a/w3313 ), .Z(n10982)
         );
  AND U6225 ( .A(\SUBBYTES[5].a/w3119 ), .B(\SUBBYTES[5].a/w3108 ), .Z(n10981)
         );
  AND U6226 ( .A(\SUBBYTES[5].a/w3119 ), .B(\SUBBYTES[5].a/w3106 ), .Z(n10980)
         );
  AND U6227 ( .A(\SUBBYTES[5].a/w2912 ), .B(\SUBBYTES[5].a/w2901 ), .Z(n10979)
         );
  AND U6228 ( .A(\SUBBYTES[5].a/w2912 ), .B(\SUBBYTES[5].a/w2899 ), .Z(n10978)
         );
  AND U6229 ( .A(\SUBBYTES[5].a/w2705 ), .B(\SUBBYTES[5].a/w2694 ), .Z(n10977)
         );
  AND U6230 ( .A(\SUBBYTES[5].a/w2705 ), .B(\SUBBYTES[5].a/w2692 ), .Z(n10976)
         );
  AND U6231 ( .A(\SUBBYTES[5].a/w2498 ), .B(\SUBBYTES[5].a/w2487 ), .Z(n10975)
         );
  AND U6232 ( .A(\SUBBYTES[5].a/w2498 ), .B(\SUBBYTES[5].a/w2485 ), .Z(n10974)
         );
  AND U6233 ( .A(\SUBBYTES[5].a/w2291 ), .B(\SUBBYTES[5].a/w2280 ), .Z(n10973)
         );
  AND U6234 ( .A(\SUBBYTES[5].a/w2291 ), .B(\SUBBYTES[5].a/w2278 ), .Z(n10972)
         );
  AND U6235 ( .A(\SUBBYTES[5].a/w2084 ), .B(\SUBBYTES[5].a/w2073 ), .Z(n10971)
         );
  AND U6236 ( .A(\SUBBYTES[5].a/w221 ), .B(\SUBBYTES[5].a/w210 ), .Z(n10953)
         );
  AND U6237 ( .A(n2285), .B(\SUBBYTES[4].a/w781 ), .Z(\SUBBYTES[4].a/w916 ) );
  AND U6238 ( .A(n2286), .B(\SUBBYTES[4].a/w782 ), .Z(\SUBBYTES[4].a/w914 ) );
  AND U6239 ( .A(\SUBBYTES[4].a/w912 ), .B(n2287), .Z(\SUBBYTES[4].a/w913 ) );
  ANDN U6240 ( .A(\w1[4][96] ), .B(n2288), .Z(\SUBBYTES[4].a/w909 ) );
  AND U6241 ( .A(n2289), .B(\SUBBYTES[4].a/w784 ), .Z(\SUBBYTES[4].a/w907 ) );
  AND U6242 ( .A(\SUBBYTES[4].a/w905 ), .B(n2290), .Z(\SUBBYTES[4].a/w906 ) );
  XOR U6243 ( .A(\SUBBYTES[4].a/w849 ), .B(n9678), .Z(n2290) );
  AND U6244 ( .A(\SUBBYTES[4].a/w892 ), .B(\SUBBYTES[4].a/w894 ), .Z(
        \SUBBYTES[4].a/w901 ) );
  AND U6245 ( .A(\SUBBYTES[4].a/w893 ), .B(\SUBBYTES[4].a/w895 ), .Z(
        \SUBBYTES[4].a/w899 ) );
  AND U6246 ( .A(\SUBBYTES[4].a/w896 ), .B(\SUBBYTES[4].a/w897 ), .Z(
        \SUBBYTES[4].a/w898 ) );
  AND U6247 ( .A(\SUBBYTES[4].a/w785 ), .B(n2285), .Z(\SUBBYTES[4].a/w884 ) );
  XOR U6248 ( .A(\SUBBYTES[4].a/w853 ), .B(n1008), .Z(n2285) );
  AND U6249 ( .A(\SUBBYTES[4].a/w786 ), .B(n2286), .Z(\SUBBYTES[4].a/w882 ) );
  XOR U6250 ( .A(n9679), .B(\SUBBYTES[4].a/w853 ), .Z(n2286) );
  ANDN U6251 ( .A(n2287), .B(n2291), .Z(\SUBBYTES[4].a/w881 ) );
  XOR U6252 ( .A(n1008), .B(n9679), .Z(n2287) );
  ANDN U6253 ( .A(\SUBBYTES[4].a/w787 ), .B(n2288), .Z(\SUBBYTES[4].a/w877 )
         );
  XNOR U6254 ( .A(\SUBBYTES[4].a/w846 ), .B(\SUBBYTES[4].a/w849 ), .Z(n2288)
         );
  AND U6255 ( .A(\SUBBYTES[4].a/w788 ), .B(n2289), .Z(\SUBBYTES[4].a/w875 ) );
  XNOR U6256 ( .A(n2292), .B(\SUBBYTES[4].a/w846 ), .Z(n2289) );
  AND U6257 ( .A(\SUBBYTES[4].a/w873 ), .B(n2293), .Z(\SUBBYTES[4].a/w874 ) );
  XOR U6258 ( .A(n2294), .B(n2292), .Z(n2293) );
  IV U6259 ( .A(n9678), .Z(n2292) );
  ANDN U6260 ( .A(\SUBBYTES[4].a/w892 ), .B(n2295), .Z(\SUBBYTES[4].a/w869 )
         );
  ANDN U6261 ( .A(\SUBBYTES[4].a/w893 ), .B(n2296), .Z(\SUBBYTES[4].a/w867 )
         );
  ANDN U6262 ( .A(\SUBBYTES[4].a/w896 ), .B(n2297), .Z(\SUBBYTES[4].a/w866 )
         );
  AND U6263 ( .A(\SUBBYTES[4].a/w852 ), .B(\SUBBYTES[4].a/w851 ), .Z(
        \SUBBYTES[4].a/w853 ) );
  IV U6264 ( .A(n2294), .Z(\SUBBYTES[4].a/w849 ) );
  NAND U6265 ( .A(\SUBBYTES[4].a/w828 ), .B(\SUBBYTES[4].a/w843 ), .Z(n2294)
         );
  AND U6266 ( .A(\SUBBYTES[4].a/w845 ), .B(\SUBBYTES[4].a/w851 ), .Z(
        \SUBBYTES[4].a/w846 ) );
  AND U6267 ( .A(\SUBBYTES[4].a/w830 ), .B(\SUBBYTES[4].a/w828 ), .Z(
        \SUBBYTES[4].a/w840 ) );
  AND U6268 ( .A(\SUBBYTES[4].a/w831 ), .B(\SUBBYTES[4].a/w829 ), .Z(
        \SUBBYTES[4].a/w838 ) );
  AND U6269 ( .A(\SUBBYTES[4].a/w845 ), .B(\SUBBYTES[4].a/w852 ), .Z(
        \SUBBYTES[4].a/w837 ) );
  AND U6270 ( .A(\SUBBYTES[4].a/w785 ), .B(\SUBBYTES[4].a/w781 ), .Z(
        \SUBBYTES[4].a/w822 ) );
  AND U6271 ( .A(\SUBBYTES[4].a/w786 ), .B(\SUBBYTES[4].a/w782 ), .Z(
        \SUBBYTES[4].a/w820 ) );
  ANDN U6272 ( .A(\SUBBYTES[4].a/w912 ), .B(n2291), .Z(\SUBBYTES[4].a/w819 )
         );
  XNOR U6273 ( .A(\w1[4][103] ), .B(\w1[4][97] ), .Z(n2291) );
  XOR U6274 ( .A(\w0[4][97] ), .B(g_input[609]), .Z(\w1[4][97] ) );
  IV U6275 ( .A(n2298), .Z(\w1[4][103] ) );
  AND U6276 ( .A(\w1[4][96] ), .B(\SUBBYTES[4].a/w787 ), .Z(
        \SUBBYTES[4].a/w815 ) );
  XOR U6277 ( .A(\w0[4][96] ), .B(g_input[608]), .Z(\w1[4][96] ) );
  AND U6278 ( .A(\SUBBYTES[4].a/w788 ), .B(\SUBBYTES[4].a/w784 ), .Z(
        \SUBBYTES[4].a/w813 ) );
  AND U6279 ( .A(\SUBBYTES[4].a/w873 ), .B(\SUBBYTES[4].a/w905 ), .Z(
        \SUBBYTES[4].a/w812 ) );
  ANDN U6280 ( .A(\SUBBYTES[4].a/w894 ), .B(n2295), .Z(\SUBBYTES[4].a/w807 )
         );
  XOR U6281 ( .A(\w1[4][100] ), .B(n2298), .Z(n2295) );
  ANDN U6282 ( .A(\SUBBYTES[4].a/w895 ), .B(n2296), .Z(\SUBBYTES[4].a/w805 )
         );
  XOR U6283 ( .A(n2298), .B(\w1[4][98] ), .Z(n2296) );
  XNOR U6284 ( .A(\w0[4][103] ), .B(g_input[615]), .Z(n2298) );
  ANDN U6285 ( .A(\SUBBYTES[4].a/w897 ), .B(n2297), .Z(\SUBBYTES[4].a/w804 )
         );
  XNOR U6286 ( .A(\w1[4][100] ), .B(\w1[4][98] ), .Z(n2297) );
  XOR U6287 ( .A(\w0[4][98] ), .B(g_input[610]), .Z(\w1[4][98] ) );
  XOR U6288 ( .A(\w0[4][100] ), .B(g_input[612]), .Z(\w1[4][100] ) );
  AND U6289 ( .A(n2299), .B(\SUBBYTES[4].a/w574 ), .Z(\SUBBYTES[4].a/w709 ) );
  AND U6290 ( .A(n2300), .B(\SUBBYTES[4].a/w575 ), .Z(\SUBBYTES[4].a/w707 ) );
  AND U6291 ( .A(\SUBBYTES[4].a/w705 ), .B(n2301), .Z(\SUBBYTES[4].a/w706 ) );
  ANDN U6292 ( .A(\w1[4][104] ), .B(n2302), .Z(\SUBBYTES[4].a/w702 ) );
  AND U6293 ( .A(n2303), .B(\SUBBYTES[4].a/w577 ), .Z(\SUBBYTES[4].a/w700 ) );
  AND U6294 ( .A(\SUBBYTES[4].a/w698 ), .B(n2304), .Z(\SUBBYTES[4].a/w699 ) );
  XOR U6295 ( .A(\SUBBYTES[4].a/w642 ), .B(n9676), .Z(n2304) );
  AND U6296 ( .A(\SUBBYTES[4].a/w685 ), .B(\SUBBYTES[4].a/w687 ), .Z(
        \SUBBYTES[4].a/w694 ) );
  AND U6297 ( .A(\SUBBYTES[4].a/w686 ), .B(\SUBBYTES[4].a/w688 ), .Z(
        \SUBBYTES[4].a/w692 ) );
  AND U6298 ( .A(\SUBBYTES[4].a/w689 ), .B(\SUBBYTES[4].a/w690 ), .Z(
        \SUBBYTES[4].a/w691 ) );
  AND U6299 ( .A(\SUBBYTES[4].a/w578 ), .B(n2299), .Z(\SUBBYTES[4].a/w677 ) );
  XOR U6300 ( .A(\SUBBYTES[4].a/w646 ), .B(n1007), .Z(n2299) );
  AND U6301 ( .A(\SUBBYTES[4].a/w579 ), .B(n2300), .Z(\SUBBYTES[4].a/w675 ) );
  XOR U6302 ( .A(n9677), .B(\SUBBYTES[4].a/w646 ), .Z(n2300) );
  ANDN U6303 ( .A(n2301), .B(n2305), .Z(\SUBBYTES[4].a/w674 ) );
  XOR U6304 ( .A(n1007), .B(n9677), .Z(n2301) );
  ANDN U6305 ( .A(\SUBBYTES[4].a/w580 ), .B(n2302), .Z(\SUBBYTES[4].a/w670 )
         );
  XNOR U6306 ( .A(\SUBBYTES[4].a/w639 ), .B(\SUBBYTES[4].a/w642 ), .Z(n2302)
         );
  AND U6307 ( .A(\SUBBYTES[4].a/w581 ), .B(n2303), .Z(\SUBBYTES[4].a/w668 ) );
  XNOR U6308 ( .A(n2306), .B(\SUBBYTES[4].a/w639 ), .Z(n2303) );
  AND U6309 ( .A(\SUBBYTES[4].a/w666 ), .B(n2307), .Z(\SUBBYTES[4].a/w667 ) );
  XOR U6310 ( .A(n2308), .B(n2306), .Z(n2307) );
  IV U6311 ( .A(n9676), .Z(n2306) );
  ANDN U6312 ( .A(\SUBBYTES[4].a/w685 ), .B(n2309), .Z(\SUBBYTES[4].a/w662 )
         );
  ANDN U6313 ( .A(\SUBBYTES[4].a/w686 ), .B(n2310), .Z(\SUBBYTES[4].a/w660 )
         );
  ANDN U6314 ( .A(\SUBBYTES[4].a/w689 ), .B(n2311), .Z(\SUBBYTES[4].a/w659 )
         );
  AND U6315 ( .A(\SUBBYTES[4].a/w645 ), .B(\SUBBYTES[4].a/w644 ), .Z(
        \SUBBYTES[4].a/w646 ) );
  IV U6316 ( .A(n2308), .Z(\SUBBYTES[4].a/w642 ) );
  NAND U6317 ( .A(\SUBBYTES[4].a/w621 ), .B(\SUBBYTES[4].a/w636 ), .Z(n2308)
         );
  AND U6318 ( .A(\SUBBYTES[4].a/w638 ), .B(\SUBBYTES[4].a/w644 ), .Z(
        \SUBBYTES[4].a/w639 ) );
  AND U6319 ( .A(\SUBBYTES[4].a/w623 ), .B(\SUBBYTES[4].a/w621 ), .Z(
        \SUBBYTES[4].a/w633 ) );
  AND U6320 ( .A(\SUBBYTES[4].a/w624 ), .B(\SUBBYTES[4].a/w622 ), .Z(
        \SUBBYTES[4].a/w631 ) );
  AND U6321 ( .A(\SUBBYTES[4].a/w638 ), .B(\SUBBYTES[4].a/w645 ), .Z(
        \SUBBYTES[4].a/w630 ) );
  AND U6322 ( .A(\SUBBYTES[4].a/w578 ), .B(\SUBBYTES[4].a/w574 ), .Z(
        \SUBBYTES[4].a/w615 ) );
  AND U6323 ( .A(\SUBBYTES[4].a/w579 ), .B(\SUBBYTES[4].a/w575 ), .Z(
        \SUBBYTES[4].a/w613 ) );
  ANDN U6324 ( .A(\SUBBYTES[4].a/w705 ), .B(n2305), .Z(\SUBBYTES[4].a/w612 )
         );
  XNOR U6325 ( .A(\w1[4][105] ), .B(\w1[4][111] ), .Z(n2305) );
  XOR U6326 ( .A(\w0[4][105] ), .B(g_input[617]), .Z(\w1[4][105] ) );
  AND U6327 ( .A(\w1[4][104] ), .B(\SUBBYTES[4].a/w580 ), .Z(
        \SUBBYTES[4].a/w608 ) );
  XOR U6328 ( .A(\w0[4][104] ), .B(g_input[616]), .Z(\w1[4][104] ) );
  AND U6329 ( .A(\SUBBYTES[4].a/w581 ), .B(\SUBBYTES[4].a/w577 ), .Z(
        \SUBBYTES[4].a/w606 ) );
  AND U6330 ( .A(\SUBBYTES[4].a/w666 ), .B(\SUBBYTES[4].a/w698 ), .Z(
        \SUBBYTES[4].a/w605 ) );
  ANDN U6331 ( .A(\SUBBYTES[4].a/w687 ), .B(n2309), .Z(\SUBBYTES[4].a/w600 )
         );
  XNOR U6332 ( .A(\w1[4][108] ), .B(\w1[4][111] ), .Z(n2309) );
  ANDN U6333 ( .A(\SUBBYTES[4].a/w688 ), .B(n2310), .Z(\SUBBYTES[4].a/w598 )
         );
  XNOR U6334 ( .A(\w1[4][106] ), .B(\w1[4][111] ), .Z(n2310) );
  XOR U6335 ( .A(\w0[4][111] ), .B(g_input[623]), .Z(\w1[4][111] ) );
  IV U6336 ( .A(n2312), .Z(\w1[4][106] ) );
  ANDN U6337 ( .A(\SUBBYTES[4].a/w690 ), .B(n2311), .Z(\SUBBYTES[4].a/w597 )
         );
  XOR U6338 ( .A(n2312), .B(\w1[4][108] ), .Z(n2311) );
  XOR U6339 ( .A(\w0[4][108] ), .B(g_input[620]), .Z(\w1[4][108] ) );
  XNOR U6340 ( .A(\w0[4][106] ), .B(g_input[618]), .Z(n2312) );
  AND U6341 ( .A(n2313), .B(\SUBBYTES[4].a/w367 ), .Z(\SUBBYTES[4].a/w502 ) );
  AND U6342 ( .A(n2314), .B(\SUBBYTES[4].a/w368 ), .Z(\SUBBYTES[4].a/w500 ) );
  AND U6343 ( .A(\SUBBYTES[4].a/w498 ), .B(n2315), .Z(\SUBBYTES[4].a/w499 ) );
  ANDN U6344 ( .A(\w1[4][112] ), .B(n2316), .Z(\SUBBYTES[4].a/w495 ) );
  AND U6345 ( .A(n2317), .B(\SUBBYTES[4].a/w370 ), .Z(\SUBBYTES[4].a/w493 ) );
  AND U6346 ( .A(\SUBBYTES[4].a/w491 ), .B(n2318), .Z(\SUBBYTES[4].a/w492 ) );
  XOR U6347 ( .A(\SUBBYTES[4].a/w435 ), .B(n9674), .Z(n2318) );
  AND U6348 ( .A(\SUBBYTES[4].a/w478 ), .B(\SUBBYTES[4].a/w480 ), .Z(
        \SUBBYTES[4].a/w487 ) );
  AND U6349 ( .A(\SUBBYTES[4].a/w479 ), .B(\SUBBYTES[4].a/w481 ), .Z(
        \SUBBYTES[4].a/w485 ) );
  AND U6350 ( .A(\SUBBYTES[4].a/w482 ), .B(\SUBBYTES[4].a/w483 ), .Z(
        \SUBBYTES[4].a/w484 ) );
  AND U6351 ( .A(\SUBBYTES[4].a/w371 ), .B(n2313), .Z(\SUBBYTES[4].a/w470 ) );
  XOR U6352 ( .A(\SUBBYTES[4].a/w439 ), .B(n1006), .Z(n2313) );
  AND U6353 ( .A(\SUBBYTES[4].a/w372 ), .B(n2314), .Z(\SUBBYTES[4].a/w468 ) );
  XOR U6354 ( .A(n9675), .B(\SUBBYTES[4].a/w439 ), .Z(n2314) );
  ANDN U6355 ( .A(n2315), .B(n2319), .Z(\SUBBYTES[4].a/w467 ) );
  XOR U6356 ( .A(n1006), .B(n9675), .Z(n2315) );
  ANDN U6357 ( .A(\SUBBYTES[4].a/w373 ), .B(n2316), .Z(\SUBBYTES[4].a/w463 )
         );
  XNOR U6358 ( .A(\SUBBYTES[4].a/w432 ), .B(\SUBBYTES[4].a/w435 ), .Z(n2316)
         );
  AND U6359 ( .A(\SUBBYTES[4].a/w374 ), .B(n2317), .Z(\SUBBYTES[4].a/w461 ) );
  XNOR U6360 ( .A(n2320), .B(\SUBBYTES[4].a/w432 ), .Z(n2317) );
  AND U6361 ( .A(\SUBBYTES[4].a/w459 ), .B(n2321), .Z(\SUBBYTES[4].a/w460 ) );
  XOR U6362 ( .A(n2322), .B(n2320), .Z(n2321) );
  IV U6363 ( .A(n9674), .Z(n2320) );
  ANDN U6364 ( .A(\SUBBYTES[4].a/w478 ), .B(n2323), .Z(\SUBBYTES[4].a/w455 )
         );
  ANDN U6365 ( .A(\SUBBYTES[4].a/w479 ), .B(n2324), .Z(\SUBBYTES[4].a/w453 )
         );
  ANDN U6366 ( .A(\SUBBYTES[4].a/w482 ), .B(n2325), .Z(\SUBBYTES[4].a/w452 )
         );
  AND U6367 ( .A(\SUBBYTES[4].a/w438 ), .B(\SUBBYTES[4].a/w437 ), .Z(
        \SUBBYTES[4].a/w439 ) );
  IV U6368 ( .A(n2322), .Z(\SUBBYTES[4].a/w435 ) );
  NAND U6369 ( .A(\SUBBYTES[4].a/w414 ), .B(\SUBBYTES[4].a/w429 ), .Z(n2322)
         );
  AND U6370 ( .A(\SUBBYTES[4].a/w431 ), .B(\SUBBYTES[4].a/w437 ), .Z(
        \SUBBYTES[4].a/w432 ) );
  AND U6371 ( .A(\SUBBYTES[4].a/w416 ), .B(\SUBBYTES[4].a/w414 ), .Z(
        \SUBBYTES[4].a/w426 ) );
  AND U6372 ( .A(\SUBBYTES[4].a/w417 ), .B(\SUBBYTES[4].a/w415 ), .Z(
        \SUBBYTES[4].a/w424 ) );
  AND U6373 ( .A(\SUBBYTES[4].a/w431 ), .B(\SUBBYTES[4].a/w438 ), .Z(
        \SUBBYTES[4].a/w423 ) );
  AND U6374 ( .A(\SUBBYTES[4].a/w371 ), .B(\SUBBYTES[4].a/w367 ), .Z(
        \SUBBYTES[4].a/w408 ) );
  AND U6375 ( .A(\SUBBYTES[4].a/w372 ), .B(\SUBBYTES[4].a/w368 ), .Z(
        \SUBBYTES[4].a/w406 ) );
  ANDN U6376 ( .A(\SUBBYTES[4].a/w498 ), .B(n2319), .Z(\SUBBYTES[4].a/w405 )
         );
  XNOR U6377 ( .A(\w1[4][113] ), .B(\w1[4][119] ), .Z(n2319) );
  XOR U6378 ( .A(\w0[4][113] ), .B(g_input[625]), .Z(\w1[4][113] ) );
  AND U6379 ( .A(\w1[4][112] ), .B(\SUBBYTES[4].a/w373 ), .Z(
        \SUBBYTES[4].a/w401 ) );
  XOR U6380 ( .A(\w0[4][112] ), .B(g_input[624]), .Z(\w1[4][112] ) );
  AND U6381 ( .A(\SUBBYTES[4].a/w374 ), .B(\SUBBYTES[4].a/w370 ), .Z(
        \SUBBYTES[4].a/w399 ) );
  AND U6382 ( .A(\SUBBYTES[4].a/w459 ), .B(\SUBBYTES[4].a/w491 ), .Z(
        \SUBBYTES[4].a/w398 ) );
  ANDN U6383 ( .A(\SUBBYTES[4].a/w480 ), .B(n2323), .Z(\SUBBYTES[4].a/w393 )
         );
  XNOR U6384 ( .A(\w1[4][116] ), .B(\w1[4][119] ), .Z(n2323) );
  ANDN U6385 ( .A(\SUBBYTES[4].a/w481 ), .B(n2324), .Z(\SUBBYTES[4].a/w391 )
         );
  XNOR U6386 ( .A(\w1[4][114] ), .B(\w1[4][119] ), .Z(n2324) );
  XOR U6387 ( .A(\w0[4][119] ), .B(g_input[631]), .Z(\w1[4][119] ) );
  IV U6388 ( .A(n2326), .Z(\w1[4][114] ) );
  ANDN U6389 ( .A(\SUBBYTES[4].a/w483 ), .B(n2325), .Z(\SUBBYTES[4].a/w390 )
         );
  XOR U6390 ( .A(n2326), .B(\w1[4][116] ), .Z(n2325) );
  XOR U6391 ( .A(\w0[4][116] ), .B(g_input[628]), .Z(\w1[4][116] ) );
  XNOR U6392 ( .A(\w0[4][114] ), .B(g_input[626]), .Z(n2326) );
  AND U6393 ( .A(n2327), .B(\SUBBYTES[4].a/w3265 ), .Z(\SUBBYTES[4].a/w3400 )
         );
  AND U6394 ( .A(n2328), .B(\SUBBYTES[4].a/w3266 ), .Z(\SUBBYTES[4].a/w3398 )
         );
  AND U6395 ( .A(\SUBBYTES[4].a/w3396 ), .B(n2329), .Z(\SUBBYTES[4].a/w3397 )
         );
  ANDN U6396 ( .A(\w1[4][0] ), .B(n2330), .Z(\SUBBYTES[4].a/w3393 ) );
  AND U6397 ( .A(n2331), .B(\SUBBYTES[4].a/w3268 ), .Z(\SUBBYTES[4].a/w3391 )
         );
  AND U6398 ( .A(\SUBBYTES[4].a/w3389 ), .B(n2332), .Z(\SUBBYTES[4].a/w3390 )
         );
  XOR U6399 ( .A(\SUBBYTES[4].a/w3333 ), .B(n9702), .Z(n2332) );
  AND U6400 ( .A(\SUBBYTES[4].a/w3376 ), .B(\SUBBYTES[4].a/w3378 ), .Z(
        \SUBBYTES[4].a/w3385 ) );
  AND U6401 ( .A(\SUBBYTES[4].a/w3377 ), .B(\SUBBYTES[4].a/w3379 ), .Z(
        \SUBBYTES[4].a/w3383 ) );
  AND U6402 ( .A(\SUBBYTES[4].a/w3380 ), .B(\SUBBYTES[4].a/w3381 ), .Z(
        \SUBBYTES[4].a/w3382 ) );
  AND U6403 ( .A(\SUBBYTES[4].a/w3269 ), .B(n2327), .Z(\SUBBYTES[4].a/w3368 )
         );
  XOR U6404 ( .A(\SUBBYTES[4].a/w3337 ), .B(n1020), .Z(n2327) );
  AND U6405 ( .A(\SUBBYTES[4].a/w3270 ), .B(n2328), .Z(\SUBBYTES[4].a/w3366 )
         );
  XOR U6406 ( .A(n9703), .B(\SUBBYTES[4].a/w3337 ), .Z(n2328) );
  ANDN U6407 ( .A(n2329), .B(n2333), .Z(\SUBBYTES[4].a/w3365 ) );
  XOR U6408 ( .A(n1020), .B(n9703), .Z(n2329) );
  ANDN U6409 ( .A(\SUBBYTES[4].a/w3271 ), .B(n2330), .Z(\SUBBYTES[4].a/w3361 )
         );
  XNOR U6410 ( .A(\SUBBYTES[4].a/w3330 ), .B(\SUBBYTES[4].a/w3333 ), .Z(n2330)
         );
  AND U6411 ( .A(\SUBBYTES[4].a/w3272 ), .B(n2331), .Z(\SUBBYTES[4].a/w3359 )
         );
  XNOR U6412 ( .A(n2334), .B(\SUBBYTES[4].a/w3330 ), .Z(n2331) );
  AND U6413 ( .A(\SUBBYTES[4].a/w3357 ), .B(n2335), .Z(\SUBBYTES[4].a/w3358 )
         );
  XOR U6414 ( .A(n2336), .B(n2334), .Z(n2335) );
  IV U6415 ( .A(n9702), .Z(n2334) );
  ANDN U6416 ( .A(\SUBBYTES[4].a/w3376 ), .B(n2337), .Z(\SUBBYTES[4].a/w3353 )
         );
  ANDN U6417 ( .A(\SUBBYTES[4].a/w3377 ), .B(n2338), .Z(\SUBBYTES[4].a/w3351 )
         );
  ANDN U6418 ( .A(\SUBBYTES[4].a/w3380 ), .B(n2339), .Z(\SUBBYTES[4].a/w3350 )
         );
  AND U6419 ( .A(\SUBBYTES[4].a/w3336 ), .B(\SUBBYTES[4].a/w3335 ), .Z(
        \SUBBYTES[4].a/w3337 ) );
  IV U6420 ( .A(n2336), .Z(\SUBBYTES[4].a/w3333 ) );
  NAND U6421 ( .A(\SUBBYTES[4].a/w3312 ), .B(\SUBBYTES[4].a/w3327 ), .Z(n2336)
         );
  AND U6422 ( .A(\SUBBYTES[4].a/w3329 ), .B(\SUBBYTES[4].a/w3335 ), .Z(
        \SUBBYTES[4].a/w3330 ) );
  AND U6423 ( .A(\SUBBYTES[4].a/w3314 ), .B(\SUBBYTES[4].a/w3312 ), .Z(
        \SUBBYTES[4].a/w3324 ) );
  AND U6424 ( .A(\SUBBYTES[4].a/w3315 ), .B(\SUBBYTES[4].a/w3313 ), .Z(
        \SUBBYTES[4].a/w3322 ) );
  AND U6425 ( .A(\SUBBYTES[4].a/w3329 ), .B(\SUBBYTES[4].a/w3336 ), .Z(
        \SUBBYTES[4].a/w3321 ) );
  AND U6426 ( .A(\SUBBYTES[4].a/w3269 ), .B(\SUBBYTES[4].a/w3265 ), .Z(
        \SUBBYTES[4].a/w3306 ) );
  AND U6427 ( .A(\SUBBYTES[4].a/w3270 ), .B(\SUBBYTES[4].a/w3266 ), .Z(
        \SUBBYTES[4].a/w3304 ) );
  ANDN U6428 ( .A(\SUBBYTES[4].a/w3396 ), .B(n2333), .Z(\SUBBYTES[4].a/w3303 )
         );
  XNOR U6429 ( .A(\w1[4][1] ), .B(\w1[4][7] ), .Z(n2333) );
  XOR U6430 ( .A(\w0[4][1] ), .B(g_input[513]), .Z(\w1[4][1] ) );
  AND U6431 ( .A(\w1[4][0] ), .B(\SUBBYTES[4].a/w3271 ), .Z(
        \SUBBYTES[4].a/w3299 ) );
  XOR U6432 ( .A(\w0[4][0] ), .B(g_input[512]), .Z(\w1[4][0] ) );
  AND U6433 ( .A(\SUBBYTES[4].a/w3272 ), .B(\SUBBYTES[4].a/w3268 ), .Z(
        \SUBBYTES[4].a/w3297 ) );
  AND U6434 ( .A(\SUBBYTES[4].a/w3357 ), .B(\SUBBYTES[4].a/w3389 ), .Z(
        \SUBBYTES[4].a/w3296 ) );
  ANDN U6435 ( .A(\SUBBYTES[4].a/w3378 ), .B(n2337), .Z(\SUBBYTES[4].a/w3291 )
         );
  XNOR U6436 ( .A(\w1[4][4] ), .B(\w1[4][7] ), .Z(n2337) );
  ANDN U6437 ( .A(\SUBBYTES[4].a/w3379 ), .B(n2338), .Z(\SUBBYTES[4].a/w3289 )
         );
  XNOR U6438 ( .A(\w1[4][2] ), .B(\w1[4][7] ), .Z(n2338) );
  XOR U6439 ( .A(\w0[4][7] ), .B(g_input[519]), .Z(\w1[4][7] ) );
  IV U6440 ( .A(n2340), .Z(\w1[4][2] ) );
  ANDN U6441 ( .A(\SUBBYTES[4].a/w3381 ), .B(n2339), .Z(\SUBBYTES[4].a/w3288 )
         );
  XOR U6442 ( .A(n2340), .B(\w1[4][4] ), .Z(n2339) );
  XOR U6443 ( .A(\w0[4][4] ), .B(g_input[516]), .Z(\w1[4][4] ) );
  XNOR U6444 ( .A(\w0[4][2] ), .B(g_input[514]), .Z(n2340) );
  AND U6445 ( .A(n2341), .B(\SUBBYTES[4].a/w3058 ), .Z(\SUBBYTES[4].a/w3193 )
         );
  AND U6446 ( .A(n2342), .B(\SUBBYTES[4].a/w3059 ), .Z(\SUBBYTES[4].a/w3191 )
         );
  AND U6447 ( .A(\SUBBYTES[4].a/w3189 ), .B(n2343), .Z(\SUBBYTES[4].a/w3190 )
         );
  ANDN U6448 ( .A(\w1[4][8] ), .B(n2344), .Z(\SUBBYTES[4].a/w3186 ) );
  AND U6449 ( .A(n2345), .B(\SUBBYTES[4].a/w3061 ), .Z(\SUBBYTES[4].a/w3184 )
         );
  AND U6450 ( .A(\SUBBYTES[4].a/w3182 ), .B(n2346), .Z(\SUBBYTES[4].a/w3183 )
         );
  XOR U6451 ( .A(\SUBBYTES[4].a/w3126 ), .B(n9700), .Z(n2346) );
  AND U6452 ( .A(\SUBBYTES[4].a/w3169 ), .B(\SUBBYTES[4].a/w3171 ), .Z(
        \SUBBYTES[4].a/w3178 ) );
  AND U6453 ( .A(\SUBBYTES[4].a/w3170 ), .B(\SUBBYTES[4].a/w3172 ), .Z(
        \SUBBYTES[4].a/w3176 ) );
  AND U6454 ( .A(\SUBBYTES[4].a/w3173 ), .B(\SUBBYTES[4].a/w3174 ), .Z(
        \SUBBYTES[4].a/w3175 ) );
  AND U6455 ( .A(\SUBBYTES[4].a/w3062 ), .B(n2341), .Z(\SUBBYTES[4].a/w3161 )
         );
  XOR U6456 ( .A(\SUBBYTES[4].a/w3130 ), .B(n1019), .Z(n2341) );
  AND U6457 ( .A(\SUBBYTES[4].a/w3063 ), .B(n2342), .Z(\SUBBYTES[4].a/w3159 )
         );
  XOR U6458 ( .A(n9701), .B(\SUBBYTES[4].a/w3130 ), .Z(n2342) );
  ANDN U6459 ( .A(n2343), .B(n2347), .Z(\SUBBYTES[4].a/w3158 ) );
  XOR U6460 ( .A(n1019), .B(n9701), .Z(n2343) );
  ANDN U6461 ( .A(\SUBBYTES[4].a/w3064 ), .B(n2344), .Z(\SUBBYTES[4].a/w3154 )
         );
  XNOR U6462 ( .A(\SUBBYTES[4].a/w3123 ), .B(\SUBBYTES[4].a/w3126 ), .Z(n2344)
         );
  AND U6463 ( .A(\SUBBYTES[4].a/w3065 ), .B(n2345), .Z(\SUBBYTES[4].a/w3152 )
         );
  XNOR U6464 ( .A(n2348), .B(\SUBBYTES[4].a/w3123 ), .Z(n2345) );
  AND U6465 ( .A(\SUBBYTES[4].a/w3150 ), .B(n2349), .Z(\SUBBYTES[4].a/w3151 )
         );
  XOR U6466 ( .A(n2350), .B(n2348), .Z(n2349) );
  IV U6467 ( .A(n9700), .Z(n2348) );
  ANDN U6468 ( .A(\SUBBYTES[4].a/w3169 ), .B(n2351), .Z(\SUBBYTES[4].a/w3146 )
         );
  ANDN U6469 ( .A(\SUBBYTES[4].a/w3170 ), .B(n2352), .Z(\SUBBYTES[4].a/w3144 )
         );
  ANDN U6470 ( .A(\SUBBYTES[4].a/w3173 ), .B(n2353), .Z(\SUBBYTES[4].a/w3143 )
         );
  AND U6471 ( .A(\SUBBYTES[4].a/w3129 ), .B(\SUBBYTES[4].a/w3128 ), .Z(
        \SUBBYTES[4].a/w3130 ) );
  IV U6472 ( .A(n2350), .Z(\SUBBYTES[4].a/w3126 ) );
  NAND U6473 ( .A(\SUBBYTES[4].a/w3105 ), .B(\SUBBYTES[4].a/w3120 ), .Z(n2350)
         );
  AND U6474 ( .A(\SUBBYTES[4].a/w3122 ), .B(\SUBBYTES[4].a/w3128 ), .Z(
        \SUBBYTES[4].a/w3123 ) );
  AND U6475 ( .A(\SUBBYTES[4].a/w3107 ), .B(\SUBBYTES[4].a/w3105 ), .Z(
        \SUBBYTES[4].a/w3117 ) );
  AND U6476 ( .A(\SUBBYTES[4].a/w3108 ), .B(\SUBBYTES[4].a/w3106 ), .Z(
        \SUBBYTES[4].a/w3115 ) );
  AND U6477 ( .A(\SUBBYTES[4].a/w3122 ), .B(\SUBBYTES[4].a/w3129 ), .Z(
        \SUBBYTES[4].a/w3114 ) );
  AND U6478 ( .A(\SUBBYTES[4].a/w3062 ), .B(\SUBBYTES[4].a/w3058 ), .Z(
        \SUBBYTES[4].a/w3099 ) );
  AND U6479 ( .A(\SUBBYTES[4].a/w3063 ), .B(\SUBBYTES[4].a/w3059 ), .Z(
        \SUBBYTES[4].a/w3097 ) );
  ANDN U6480 ( .A(\SUBBYTES[4].a/w3189 ), .B(n2347), .Z(\SUBBYTES[4].a/w3096 )
         );
  XNOR U6481 ( .A(\w1[4][15] ), .B(\w1[4][9] ), .Z(n2347) );
  XOR U6482 ( .A(\w0[4][9] ), .B(g_input[521]), .Z(\w1[4][9] ) );
  AND U6483 ( .A(\w1[4][8] ), .B(\SUBBYTES[4].a/w3064 ), .Z(
        \SUBBYTES[4].a/w3092 ) );
  XOR U6484 ( .A(\w0[4][8] ), .B(g_input[520]), .Z(\w1[4][8] ) );
  AND U6485 ( .A(\SUBBYTES[4].a/w3065 ), .B(\SUBBYTES[4].a/w3061 ), .Z(
        \SUBBYTES[4].a/w3090 ) );
  AND U6486 ( .A(\SUBBYTES[4].a/w3150 ), .B(\SUBBYTES[4].a/w3182 ), .Z(
        \SUBBYTES[4].a/w3089 ) );
  ANDN U6487 ( .A(\SUBBYTES[4].a/w3171 ), .B(n2351), .Z(\SUBBYTES[4].a/w3084 )
         );
  XNOR U6488 ( .A(\w1[4][12] ), .B(\w1[4][15] ), .Z(n2351) );
  ANDN U6489 ( .A(\SUBBYTES[4].a/w3172 ), .B(n2352), .Z(\SUBBYTES[4].a/w3082 )
         );
  XNOR U6490 ( .A(\w1[4][10] ), .B(\w1[4][15] ), .Z(n2352) );
  XOR U6491 ( .A(\w0[4][15] ), .B(g_input[527]), .Z(\w1[4][15] ) );
  ANDN U6492 ( .A(\SUBBYTES[4].a/w3174 ), .B(n2353), .Z(\SUBBYTES[4].a/w3081 )
         );
  XNOR U6493 ( .A(\w1[4][10] ), .B(\w1[4][12] ), .Z(n2353) );
  XOR U6494 ( .A(\w0[4][12] ), .B(g_input[524]), .Z(\w1[4][12] ) );
  XOR U6495 ( .A(\w0[4][10] ), .B(g_input[522]), .Z(\w1[4][10] ) );
  AND U6496 ( .A(n2354), .B(\SUBBYTES[4].a/w2851 ), .Z(\SUBBYTES[4].a/w2986 )
         );
  AND U6497 ( .A(n2355), .B(\SUBBYTES[4].a/w2852 ), .Z(\SUBBYTES[4].a/w2984 )
         );
  AND U6498 ( .A(\SUBBYTES[4].a/w2982 ), .B(n2356), .Z(\SUBBYTES[4].a/w2983 )
         );
  ANDN U6499 ( .A(\w1[4][16] ), .B(n2357), .Z(\SUBBYTES[4].a/w2979 ) );
  AND U6500 ( .A(n2358), .B(\SUBBYTES[4].a/w2854 ), .Z(\SUBBYTES[4].a/w2977 )
         );
  AND U6501 ( .A(\SUBBYTES[4].a/w2975 ), .B(n2359), .Z(\SUBBYTES[4].a/w2976 )
         );
  XOR U6502 ( .A(\SUBBYTES[4].a/w2919 ), .B(n9698), .Z(n2359) );
  AND U6503 ( .A(\SUBBYTES[4].a/w2962 ), .B(\SUBBYTES[4].a/w2964 ), .Z(
        \SUBBYTES[4].a/w2971 ) );
  AND U6504 ( .A(\SUBBYTES[4].a/w2963 ), .B(\SUBBYTES[4].a/w2965 ), .Z(
        \SUBBYTES[4].a/w2969 ) );
  AND U6505 ( .A(\SUBBYTES[4].a/w2966 ), .B(\SUBBYTES[4].a/w2967 ), .Z(
        \SUBBYTES[4].a/w2968 ) );
  AND U6506 ( .A(\SUBBYTES[4].a/w2855 ), .B(n2354), .Z(\SUBBYTES[4].a/w2954 )
         );
  XOR U6507 ( .A(\SUBBYTES[4].a/w2923 ), .B(n1018), .Z(n2354) );
  AND U6508 ( .A(\SUBBYTES[4].a/w2856 ), .B(n2355), .Z(\SUBBYTES[4].a/w2952 )
         );
  XOR U6509 ( .A(n9699), .B(\SUBBYTES[4].a/w2923 ), .Z(n2355) );
  ANDN U6510 ( .A(n2356), .B(n2360), .Z(\SUBBYTES[4].a/w2951 ) );
  XOR U6511 ( .A(n1018), .B(n9699), .Z(n2356) );
  AND U6512 ( .A(n2361), .B(\SUBBYTES[4].a/w160 ), .Z(\SUBBYTES[4].a/w295 ) );
  ANDN U6513 ( .A(\SUBBYTES[4].a/w2857 ), .B(n2357), .Z(\SUBBYTES[4].a/w2947 )
         );
  XNOR U6514 ( .A(\SUBBYTES[4].a/w2916 ), .B(\SUBBYTES[4].a/w2919 ), .Z(n2357)
         );
  AND U6515 ( .A(\SUBBYTES[4].a/w2858 ), .B(n2358), .Z(\SUBBYTES[4].a/w2945 )
         );
  XNOR U6516 ( .A(n2362), .B(\SUBBYTES[4].a/w2916 ), .Z(n2358) );
  AND U6517 ( .A(\SUBBYTES[4].a/w2943 ), .B(n2363), .Z(\SUBBYTES[4].a/w2944 )
         );
  XOR U6518 ( .A(n2364), .B(n2362), .Z(n2363) );
  IV U6519 ( .A(n9698), .Z(n2362) );
  ANDN U6520 ( .A(\SUBBYTES[4].a/w2962 ), .B(n2365), .Z(\SUBBYTES[4].a/w2939 )
         );
  ANDN U6521 ( .A(\SUBBYTES[4].a/w2963 ), .B(n2366), .Z(\SUBBYTES[4].a/w2937 )
         );
  ANDN U6522 ( .A(\SUBBYTES[4].a/w2966 ), .B(n2367), .Z(\SUBBYTES[4].a/w2936 )
         );
  AND U6523 ( .A(n2368), .B(\SUBBYTES[4].a/w161 ), .Z(\SUBBYTES[4].a/w293 ) );
  AND U6524 ( .A(\SUBBYTES[4].a/w2922 ), .B(\SUBBYTES[4].a/w2921 ), .Z(
        \SUBBYTES[4].a/w2923 ) );
  AND U6525 ( .A(\SUBBYTES[4].a/w291 ), .B(n2369), .Z(\SUBBYTES[4].a/w292 ) );
  IV U6526 ( .A(n2364), .Z(\SUBBYTES[4].a/w2919 ) );
  NAND U6527 ( .A(\SUBBYTES[4].a/w2898 ), .B(\SUBBYTES[4].a/w2913 ), .Z(n2364)
         );
  AND U6528 ( .A(\SUBBYTES[4].a/w2915 ), .B(\SUBBYTES[4].a/w2921 ), .Z(
        \SUBBYTES[4].a/w2916 ) );
  AND U6529 ( .A(\SUBBYTES[4].a/w2900 ), .B(\SUBBYTES[4].a/w2898 ), .Z(
        \SUBBYTES[4].a/w2910 ) );
  AND U6530 ( .A(\SUBBYTES[4].a/w2901 ), .B(\SUBBYTES[4].a/w2899 ), .Z(
        \SUBBYTES[4].a/w2908 ) );
  AND U6531 ( .A(\SUBBYTES[4].a/w2915 ), .B(\SUBBYTES[4].a/w2922 ), .Z(
        \SUBBYTES[4].a/w2907 ) );
  AND U6532 ( .A(\SUBBYTES[4].a/w2855 ), .B(\SUBBYTES[4].a/w2851 ), .Z(
        \SUBBYTES[4].a/w2892 ) );
  AND U6533 ( .A(\SUBBYTES[4].a/w2856 ), .B(\SUBBYTES[4].a/w2852 ), .Z(
        \SUBBYTES[4].a/w2890 ) );
  ANDN U6534 ( .A(\SUBBYTES[4].a/w2982 ), .B(n2360), .Z(\SUBBYTES[4].a/w2889 )
         );
  XNOR U6535 ( .A(\w1[4][17] ), .B(\w1[4][23] ), .Z(n2360) );
  XOR U6536 ( .A(\w0[4][17] ), .B(g_input[529]), .Z(\w1[4][17] ) );
  AND U6537 ( .A(\w1[4][16] ), .B(\SUBBYTES[4].a/w2857 ), .Z(
        \SUBBYTES[4].a/w2885 ) );
  XOR U6538 ( .A(\w0[4][16] ), .B(g_input[528]), .Z(\w1[4][16] ) );
  AND U6539 ( .A(\SUBBYTES[4].a/w2858 ), .B(\SUBBYTES[4].a/w2854 ), .Z(
        \SUBBYTES[4].a/w2883 ) );
  AND U6540 ( .A(\SUBBYTES[4].a/w2943 ), .B(\SUBBYTES[4].a/w2975 ), .Z(
        \SUBBYTES[4].a/w2882 ) );
  ANDN U6541 ( .A(\w1[4][120] ), .B(n2370), .Z(\SUBBYTES[4].a/w288 ) );
  ANDN U6542 ( .A(\SUBBYTES[4].a/w2964 ), .B(n2365), .Z(\SUBBYTES[4].a/w2877 )
         );
  XNOR U6543 ( .A(\w1[4][20] ), .B(\w1[4][23] ), .Z(n2365) );
  ANDN U6544 ( .A(\SUBBYTES[4].a/w2965 ), .B(n2366), .Z(\SUBBYTES[4].a/w2875 )
         );
  XNOR U6545 ( .A(\w1[4][18] ), .B(\w1[4][23] ), .Z(n2366) );
  XOR U6546 ( .A(\w0[4][23] ), .B(g_input[535]), .Z(\w1[4][23] ) );
  IV U6547 ( .A(n2371), .Z(\w1[4][18] ) );
  ANDN U6548 ( .A(\SUBBYTES[4].a/w2967 ), .B(n2367), .Z(\SUBBYTES[4].a/w2874 )
         );
  XOR U6549 ( .A(n2371), .B(\w1[4][20] ), .Z(n2367) );
  XOR U6550 ( .A(\w0[4][20] ), .B(g_input[532]), .Z(\w1[4][20] ) );
  XNOR U6551 ( .A(\w0[4][18] ), .B(g_input[530]), .Z(n2371) );
  AND U6552 ( .A(n2372), .B(\SUBBYTES[4].a/w163 ), .Z(\SUBBYTES[4].a/w286 ) );
  AND U6553 ( .A(\SUBBYTES[4].a/w284 ), .B(n2373), .Z(\SUBBYTES[4].a/w285 ) );
  XOR U6554 ( .A(\SUBBYTES[4].a/w228 ), .B(n9672), .Z(n2373) );
  AND U6555 ( .A(\SUBBYTES[4].a/w271 ), .B(\SUBBYTES[4].a/w273 ), .Z(
        \SUBBYTES[4].a/w280 ) );
  AND U6556 ( .A(\SUBBYTES[4].a/w272 ), .B(\SUBBYTES[4].a/w274 ), .Z(
        \SUBBYTES[4].a/w278 ) );
  AND U6557 ( .A(n2374), .B(\SUBBYTES[4].a/w2644 ), .Z(\SUBBYTES[4].a/w2779 )
         );
  AND U6558 ( .A(n2375), .B(\SUBBYTES[4].a/w2645 ), .Z(\SUBBYTES[4].a/w2777 )
         );
  AND U6559 ( .A(\SUBBYTES[4].a/w2775 ), .B(n2376), .Z(\SUBBYTES[4].a/w2776 )
         );
  ANDN U6560 ( .A(\w1[4][24] ), .B(n2377), .Z(\SUBBYTES[4].a/w2772 ) );
  AND U6561 ( .A(n2378), .B(\SUBBYTES[4].a/w2647 ), .Z(\SUBBYTES[4].a/w2770 )
         );
  AND U6562 ( .A(\SUBBYTES[4].a/w275 ), .B(\SUBBYTES[4].a/w276 ), .Z(
        \SUBBYTES[4].a/w277 ) );
  AND U6563 ( .A(\SUBBYTES[4].a/w2768 ), .B(n2379), .Z(\SUBBYTES[4].a/w2769 )
         );
  XOR U6564 ( .A(\SUBBYTES[4].a/w2712 ), .B(n9696), .Z(n2379) );
  AND U6565 ( .A(\SUBBYTES[4].a/w2755 ), .B(\SUBBYTES[4].a/w2757 ), .Z(
        \SUBBYTES[4].a/w2764 ) );
  AND U6566 ( .A(\SUBBYTES[4].a/w2756 ), .B(\SUBBYTES[4].a/w2758 ), .Z(
        \SUBBYTES[4].a/w2762 ) );
  AND U6567 ( .A(\SUBBYTES[4].a/w2759 ), .B(\SUBBYTES[4].a/w2760 ), .Z(
        \SUBBYTES[4].a/w2761 ) );
  AND U6568 ( .A(\SUBBYTES[4].a/w2648 ), .B(n2374), .Z(\SUBBYTES[4].a/w2747 )
         );
  XOR U6569 ( .A(\SUBBYTES[4].a/w2716 ), .B(n1017), .Z(n2374) );
  AND U6570 ( .A(\SUBBYTES[4].a/w2649 ), .B(n2375), .Z(\SUBBYTES[4].a/w2745 )
         );
  XOR U6571 ( .A(n9697), .B(\SUBBYTES[4].a/w2716 ), .Z(n2375) );
  ANDN U6572 ( .A(n2376), .B(n2380), .Z(\SUBBYTES[4].a/w2744 ) );
  XOR U6573 ( .A(n1017), .B(n9697), .Z(n2376) );
  ANDN U6574 ( .A(\SUBBYTES[4].a/w2650 ), .B(n2377), .Z(\SUBBYTES[4].a/w2740 )
         );
  XNOR U6575 ( .A(\SUBBYTES[4].a/w2709 ), .B(\SUBBYTES[4].a/w2712 ), .Z(n2377)
         );
  AND U6576 ( .A(\SUBBYTES[4].a/w2651 ), .B(n2378), .Z(\SUBBYTES[4].a/w2738 )
         );
  XNOR U6577 ( .A(n2381), .B(\SUBBYTES[4].a/w2709 ), .Z(n2378) );
  AND U6578 ( .A(\SUBBYTES[4].a/w2736 ), .B(n2382), .Z(\SUBBYTES[4].a/w2737 )
         );
  XOR U6579 ( .A(n2383), .B(n2381), .Z(n2382) );
  IV U6580 ( .A(n9696), .Z(n2381) );
  ANDN U6581 ( .A(\SUBBYTES[4].a/w2755 ), .B(n2384), .Z(\SUBBYTES[4].a/w2732 )
         );
  ANDN U6582 ( .A(\SUBBYTES[4].a/w2756 ), .B(n2385), .Z(\SUBBYTES[4].a/w2730 )
         );
  ANDN U6583 ( .A(\SUBBYTES[4].a/w2759 ), .B(n2386), .Z(\SUBBYTES[4].a/w2729 )
         );
  AND U6584 ( .A(\SUBBYTES[4].a/w2715 ), .B(\SUBBYTES[4].a/w2714 ), .Z(
        \SUBBYTES[4].a/w2716 ) );
  IV U6585 ( .A(n2383), .Z(\SUBBYTES[4].a/w2712 ) );
  NAND U6586 ( .A(\SUBBYTES[4].a/w2691 ), .B(\SUBBYTES[4].a/w2706 ), .Z(n2383)
         );
  AND U6587 ( .A(\SUBBYTES[4].a/w2708 ), .B(\SUBBYTES[4].a/w2714 ), .Z(
        \SUBBYTES[4].a/w2709 ) );
  AND U6588 ( .A(\SUBBYTES[4].a/w2693 ), .B(\SUBBYTES[4].a/w2691 ), .Z(
        \SUBBYTES[4].a/w2703 ) );
  AND U6589 ( .A(\SUBBYTES[4].a/w2694 ), .B(\SUBBYTES[4].a/w2692 ), .Z(
        \SUBBYTES[4].a/w2701 ) );
  AND U6590 ( .A(\SUBBYTES[4].a/w2708 ), .B(\SUBBYTES[4].a/w2715 ), .Z(
        \SUBBYTES[4].a/w2700 ) );
  AND U6591 ( .A(\SUBBYTES[4].a/w2648 ), .B(\SUBBYTES[4].a/w2644 ), .Z(
        \SUBBYTES[4].a/w2685 ) );
  AND U6592 ( .A(\SUBBYTES[4].a/w2649 ), .B(\SUBBYTES[4].a/w2645 ), .Z(
        \SUBBYTES[4].a/w2683 ) );
  ANDN U6593 ( .A(\SUBBYTES[4].a/w2775 ), .B(n2380), .Z(\SUBBYTES[4].a/w2682 )
         );
  XNOR U6594 ( .A(\w1[4][25] ), .B(\w1[4][31] ), .Z(n2380) );
  XOR U6595 ( .A(\w0[4][25] ), .B(g_input[537]), .Z(\w1[4][25] ) );
  AND U6596 ( .A(\w1[4][24] ), .B(\SUBBYTES[4].a/w2650 ), .Z(
        \SUBBYTES[4].a/w2678 ) );
  XOR U6597 ( .A(\w0[4][24] ), .B(g_input[536]), .Z(\w1[4][24] ) );
  AND U6598 ( .A(\SUBBYTES[4].a/w2651 ), .B(\SUBBYTES[4].a/w2647 ), .Z(
        \SUBBYTES[4].a/w2676 ) );
  AND U6599 ( .A(\SUBBYTES[4].a/w2736 ), .B(\SUBBYTES[4].a/w2768 ), .Z(
        \SUBBYTES[4].a/w2675 ) );
  ANDN U6600 ( .A(\SUBBYTES[4].a/w2757 ), .B(n2384), .Z(\SUBBYTES[4].a/w2670 )
         );
  XNOR U6601 ( .A(\w1[4][28] ), .B(\w1[4][31] ), .Z(n2384) );
  ANDN U6602 ( .A(\SUBBYTES[4].a/w2758 ), .B(n2385), .Z(\SUBBYTES[4].a/w2668 )
         );
  XNOR U6603 ( .A(\w1[4][26] ), .B(\w1[4][31] ), .Z(n2385) );
  XOR U6604 ( .A(\w0[4][31] ), .B(g_input[543]), .Z(\w1[4][31] ) );
  IV U6605 ( .A(n2387), .Z(\w1[4][26] ) );
  ANDN U6606 ( .A(\SUBBYTES[4].a/w2760 ), .B(n2386), .Z(\SUBBYTES[4].a/w2667 )
         );
  XOR U6607 ( .A(n2387), .B(\w1[4][28] ), .Z(n2386) );
  XOR U6608 ( .A(\w0[4][28] ), .B(g_input[540]), .Z(\w1[4][28] ) );
  XNOR U6609 ( .A(\w0[4][26] ), .B(g_input[538]), .Z(n2387) );
  AND U6610 ( .A(\SUBBYTES[4].a/w164 ), .B(n2361), .Z(\SUBBYTES[4].a/w263 ) );
  XOR U6611 ( .A(\SUBBYTES[4].a/w232 ), .B(n1005), .Z(n2361) );
  AND U6612 ( .A(\SUBBYTES[4].a/w165 ), .B(n2368), .Z(\SUBBYTES[4].a/w261 ) );
  XOR U6613 ( .A(n9673), .B(\SUBBYTES[4].a/w232 ), .Z(n2368) );
  ANDN U6614 ( .A(n2369), .B(n2388), .Z(\SUBBYTES[4].a/w260 ) );
  XOR U6615 ( .A(n1005), .B(n9673), .Z(n2369) );
  AND U6616 ( .A(n2389), .B(\SUBBYTES[4].a/w2437 ), .Z(\SUBBYTES[4].a/w2572 )
         );
  AND U6617 ( .A(n2390), .B(\SUBBYTES[4].a/w2438 ), .Z(\SUBBYTES[4].a/w2570 )
         );
  AND U6618 ( .A(\SUBBYTES[4].a/w2568 ), .B(n2391), .Z(\SUBBYTES[4].a/w2569 )
         );
  ANDN U6619 ( .A(\w1[4][32] ), .B(n2392), .Z(\SUBBYTES[4].a/w2565 ) );
  AND U6620 ( .A(n2393), .B(\SUBBYTES[4].a/w2440 ), .Z(\SUBBYTES[4].a/w2563 )
         );
  AND U6621 ( .A(\SUBBYTES[4].a/w2561 ), .B(n2394), .Z(\SUBBYTES[4].a/w2562 )
         );
  XOR U6622 ( .A(\SUBBYTES[4].a/w2505 ), .B(n9694), .Z(n2394) );
  ANDN U6623 ( .A(\SUBBYTES[4].a/w166 ), .B(n2370), .Z(\SUBBYTES[4].a/w256 )
         );
  XNOR U6624 ( .A(\SUBBYTES[4].a/w225 ), .B(\SUBBYTES[4].a/w228 ), .Z(n2370)
         );
  AND U6625 ( .A(\SUBBYTES[4].a/w2548 ), .B(\SUBBYTES[4].a/w2550 ), .Z(
        \SUBBYTES[4].a/w2557 ) );
  AND U6626 ( .A(\SUBBYTES[4].a/w2549 ), .B(\SUBBYTES[4].a/w2551 ), .Z(
        \SUBBYTES[4].a/w2555 ) );
  AND U6627 ( .A(\SUBBYTES[4].a/w2552 ), .B(\SUBBYTES[4].a/w2553 ), .Z(
        \SUBBYTES[4].a/w2554 ) );
  AND U6628 ( .A(\SUBBYTES[4].a/w2441 ), .B(n2389), .Z(\SUBBYTES[4].a/w2540 )
         );
  XOR U6629 ( .A(\SUBBYTES[4].a/w2509 ), .B(n1016), .Z(n2389) );
  AND U6630 ( .A(\SUBBYTES[4].a/w167 ), .B(n2372), .Z(\SUBBYTES[4].a/w254 ) );
  XNOR U6631 ( .A(n2395), .B(\SUBBYTES[4].a/w225 ), .Z(n2372) );
  AND U6632 ( .A(\SUBBYTES[4].a/w2442 ), .B(n2390), .Z(\SUBBYTES[4].a/w2538 )
         );
  XOR U6633 ( .A(n9695), .B(\SUBBYTES[4].a/w2509 ), .Z(n2390) );
  ANDN U6634 ( .A(n2391), .B(n2396), .Z(\SUBBYTES[4].a/w2537 ) );
  XOR U6635 ( .A(n1016), .B(n9695), .Z(n2391) );
  ANDN U6636 ( .A(\SUBBYTES[4].a/w2443 ), .B(n2392), .Z(\SUBBYTES[4].a/w2533 )
         );
  XNOR U6637 ( .A(\SUBBYTES[4].a/w2502 ), .B(\SUBBYTES[4].a/w2505 ), .Z(n2392)
         );
  AND U6638 ( .A(\SUBBYTES[4].a/w2444 ), .B(n2393), .Z(\SUBBYTES[4].a/w2531 )
         );
  XNOR U6639 ( .A(n2397), .B(\SUBBYTES[4].a/w2502 ), .Z(n2393) );
  AND U6640 ( .A(\SUBBYTES[4].a/w2529 ), .B(n2398), .Z(\SUBBYTES[4].a/w2530 )
         );
  XOR U6641 ( .A(n2399), .B(n2397), .Z(n2398) );
  IV U6642 ( .A(n9694), .Z(n2397) );
  AND U6643 ( .A(\SUBBYTES[4].a/w252 ), .B(n2400), .Z(\SUBBYTES[4].a/w253 ) );
  XOR U6644 ( .A(n2401), .B(n2395), .Z(n2400) );
  IV U6645 ( .A(n9672), .Z(n2395) );
  ANDN U6646 ( .A(\SUBBYTES[4].a/w2548 ), .B(n2402), .Z(\SUBBYTES[4].a/w2525 )
         );
  ANDN U6647 ( .A(\SUBBYTES[4].a/w2549 ), .B(n2403), .Z(\SUBBYTES[4].a/w2523 )
         );
  ANDN U6648 ( .A(\SUBBYTES[4].a/w2552 ), .B(n2404), .Z(\SUBBYTES[4].a/w2522 )
         );
  AND U6649 ( .A(\SUBBYTES[4].a/w2508 ), .B(\SUBBYTES[4].a/w2507 ), .Z(
        \SUBBYTES[4].a/w2509 ) );
  IV U6650 ( .A(n2399), .Z(\SUBBYTES[4].a/w2505 ) );
  NAND U6651 ( .A(\SUBBYTES[4].a/w2484 ), .B(\SUBBYTES[4].a/w2499 ), .Z(n2399)
         );
  AND U6652 ( .A(\SUBBYTES[4].a/w2501 ), .B(\SUBBYTES[4].a/w2507 ), .Z(
        \SUBBYTES[4].a/w2502 ) );
  AND U6653 ( .A(\SUBBYTES[4].a/w2486 ), .B(\SUBBYTES[4].a/w2484 ), .Z(
        \SUBBYTES[4].a/w2496 ) );
  AND U6654 ( .A(\SUBBYTES[4].a/w2487 ), .B(\SUBBYTES[4].a/w2485 ), .Z(
        \SUBBYTES[4].a/w2494 ) );
  AND U6655 ( .A(\SUBBYTES[4].a/w2501 ), .B(\SUBBYTES[4].a/w2508 ), .Z(
        \SUBBYTES[4].a/w2493 ) );
  ANDN U6656 ( .A(\SUBBYTES[4].a/w271 ), .B(n2405), .Z(\SUBBYTES[4].a/w248 )
         );
  AND U6657 ( .A(\SUBBYTES[4].a/w2441 ), .B(\SUBBYTES[4].a/w2437 ), .Z(
        \SUBBYTES[4].a/w2478 ) );
  AND U6658 ( .A(\SUBBYTES[4].a/w2442 ), .B(\SUBBYTES[4].a/w2438 ), .Z(
        \SUBBYTES[4].a/w2476 ) );
  ANDN U6659 ( .A(\SUBBYTES[4].a/w2568 ), .B(n2396), .Z(\SUBBYTES[4].a/w2475 )
         );
  XNOR U6660 ( .A(\w1[4][33] ), .B(\w1[4][39] ), .Z(n2396) );
  XOR U6661 ( .A(\w0[4][33] ), .B(g_input[545]), .Z(\w1[4][33] ) );
  AND U6662 ( .A(\w1[4][32] ), .B(\SUBBYTES[4].a/w2443 ), .Z(
        \SUBBYTES[4].a/w2471 ) );
  XOR U6663 ( .A(\w0[4][32] ), .B(g_input[544]), .Z(\w1[4][32] ) );
  AND U6664 ( .A(\SUBBYTES[4].a/w2444 ), .B(\SUBBYTES[4].a/w2440 ), .Z(
        \SUBBYTES[4].a/w2469 ) );
  AND U6665 ( .A(\SUBBYTES[4].a/w2529 ), .B(\SUBBYTES[4].a/w2561 ), .Z(
        \SUBBYTES[4].a/w2468 ) );
  ANDN U6666 ( .A(\SUBBYTES[4].a/w2550 ), .B(n2402), .Z(\SUBBYTES[4].a/w2463 )
         );
  XNOR U6667 ( .A(\w1[4][36] ), .B(\w1[4][39] ), .Z(n2402) );
  ANDN U6668 ( .A(\SUBBYTES[4].a/w2551 ), .B(n2403), .Z(\SUBBYTES[4].a/w2461 )
         );
  XNOR U6669 ( .A(\w1[4][34] ), .B(\w1[4][39] ), .Z(n2403) );
  XOR U6670 ( .A(\w0[4][39] ), .B(g_input[551]), .Z(\w1[4][39] ) );
  IV U6671 ( .A(n2406), .Z(\w1[4][34] ) );
  ANDN U6672 ( .A(\SUBBYTES[4].a/w2553 ), .B(n2404), .Z(\SUBBYTES[4].a/w2460 )
         );
  XOR U6673 ( .A(n2406), .B(\w1[4][36] ), .Z(n2404) );
  XOR U6674 ( .A(\w0[4][36] ), .B(g_input[548]), .Z(\w1[4][36] ) );
  XNOR U6675 ( .A(\w0[4][34] ), .B(g_input[546]), .Z(n2406) );
  ANDN U6676 ( .A(\SUBBYTES[4].a/w272 ), .B(n2407), .Z(\SUBBYTES[4].a/w246 )
         );
  ANDN U6677 ( .A(\SUBBYTES[4].a/w275 ), .B(n2408), .Z(\SUBBYTES[4].a/w245 )
         );
  AND U6678 ( .A(n2409), .B(\SUBBYTES[4].a/w2230 ), .Z(\SUBBYTES[4].a/w2365 )
         );
  AND U6679 ( .A(n2410), .B(\SUBBYTES[4].a/w2231 ), .Z(\SUBBYTES[4].a/w2363 )
         );
  AND U6680 ( .A(\SUBBYTES[4].a/w2361 ), .B(n2411), .Z(\SUBBYTES[4].a/w2362 )
         );
  ANDN U6681 ( .A(\w1[4][40] ), .B(n2412), .Z(\SUBBYTES[4].a/w2358 ) );
  AND U6682 ( .A(n2413), .B(\SUBBYTES[4].a/w2233 ), .Z(\SUBBYTES[4].a/w2356 )
         );
  AND U6683 ( .A(\SUBBYTES[4].a/w2354 ), .B(n2414), .Z(\SUBBYTES[4].a/w2355 )
         );
  XOR U6684 ( .A(\SUBBYTES[4].a/w2298 ), .B(n9692), .Z(n2414) );
  AND U6685 ( .A(\SUBBYTES[4].a/w2341 ), .B(\SUBBYTES[4].a/w2343 ), .Z(
        \SUBBYTES[4].a/w2350 ) );
  AND U6686 ( .A(\SUBBYTES[4].a/w2342 ), .B(\SUBBYTES[4].a/w2344 ), .Z(
        \SUBBYTES[4].a/w2348 ) );
  AND U6687 ( .A(\SUBBYTES[4].a/w2345 ), .B(\SUBBYTES[4].a/w2346 ), .Z(
        \SUBBYTES[4].a/w2347 ) );
  AND U6688 ( .A(\SUBBYTES[4].a/w2234 ), .B(n2409), .Z(\SUBBYTES[4].a/w2333 )
         );
  XOR U6689 ( .A(\SUBBYTES[4].a/w2302 ), .B(n1015), .Z(n2409) );
  AND U6690 ( .A(\SUBBYTES[4].a/w2235 ), .B(n2410), .Z(\SUBBYTES[4].a/w2331 )
         );
  XOR U6691 ( .A(n9693), .B(\SUBBYTES[4].a/w2302 ), .Z(n2410) );
  ANDN U6692 ( .A(n2411), .B(n2415), .Z(\SUBBYTES[4].a/w2330 ) );
  XOR U6693 ( .A(n1015), .B(n9693), .Z(n2411) );
  ANDN U6694 ( .A(\SUBBYTES[4].a/w2236 ), .B(n2412), .Z(\SUBBYTES[4].a/w2326 )
         );
  XNOR U6695 ( .A(\SUBBYTES[4].a/w2295 ), .B(\SUBBYTES[4].a/w2298 ), .Z(n2412)
         );
  AND U6696 ( .A(\SUBBYTES[4].a/w2237 ), .B(n2413), .Z(\SUBBYTES[4].a/w2324 )
         );
  XNOR U6697 ( .A(n2416), .B(\SUBBYTES[4].a/w2295 ), .Z(n2413) );
  AND U6698 ( .A(\SUBBYTES[4].a/w2322 ), .B(n2417), .Z(\SUBBYTES[4].a/w2323 )
         );
  XOR U6699 ( .A(n2418), .B(n2416), .Z(n2417) );
  IV U6700 ( .A(n9692), .Z(n2416) );
  AND U6701 ( .A(\SUBBYTES[4].a/w231 ), .B(\SUBBYTES[4].a/w230 ), .Z(
        \SUBBYTES[4].a/w232 ) );
  ANDN U6702 ( .A(\SUBBYTES[4].a/w2341 ), .B(n2419), .Z(\SUBBYTES[4].a/w2318 )
         );
  ANDN U6703 ( .A(\SUBBYTES[4].a/w2342 ), .B(n2420), .Z(\SUBBYTES[4].a/w2316 )
         );
  ANDN U6704 ( .A(\SUBBYTES[4].a/w2345 ), .B(n2421), .Z(\SUBBYTES[4].a/w2315 )
         );
  AND U6705 ( .A(\SUBBYTES[4].a/w2301 ), .B(\SUBBYTES[4].a/w2300 ), .Z(
        \SUBBYTES[4].a/w2302 ) );
  IV U6706 ( .A(n2418), .Z(\SUBBYTES[4].a/w2298 ) );
  NAND U6707 ( .A(\SUBBYTES[4].a/w2277 ), .B(\SUBBYTES[4].a/w2292 ), .Z(n2418)
         );
  AND U6708 ( .A(\SUBBYTES[4].a/w2294 ), .B(\SUBBYTES[4].a/w2300 ), .Z(
        \SUBBYTES[4].a/w2295 ) );
  AND U6709 ( .A(\SUBBYTES[4].a/w2279 ), .B(\SUBBYTES[4].a/w2277 ), .Z(
        \SUBBYTES[4].a/w2289 ) );
  AND U6710 ( .A(\SUBBYTES[4].a/w2280 ), .B(\SUBBYTES[4].a/w2278 ), .Z(
        \SUBBYTES[4].a/w2287 ) );
  AND U6711 ( .A(\SUBBYTES[4].a/w2294 ), .B(\SUBBYTES[4].a/w2301 ), .Z(
        \SUBBYTES[4].a/w2286 ) );
  IV U6712 ( .A(n2401), .Z(\SUBBYTES[4].a/w228 ) );
  NAND U6713 ( .A(\SUBBYTES[4].a/w207 ), .B(\SUBBYTES[4].a/w222 ), .Z(n2401)
         );
  AND U6714 ( .A(\SUBBYTES[4].a/w2234 ), .B(\SUBBYTES[4].a/w2230 ), .Z(
        \SUBBYTES[4].a/w2271 ) );
  AND U6715 ( .A(\SUBBYTES[4].a/w2235 ), .B(\SUBBYTES[4].a/w2231 ), .Z(
        \SUBBYTES[4].a/w2269 ) );
  ANDN U6716 ( .A(\SUBBYTES[4].a/w2361 ), .B(n2415), .Z(\SUBBYTES[4].a/w2268 )
         );
  XNOR U6717 ( .A(\w1[4][41] ), .B(\w1[4][47] ), .Z(n2415) );
  XOR U6718 ( .A(\w0[4][41] ), .B(g_input[553]), .Z(\w1[4][41] ) );
  AND U6719 ( .A(\w1[4][40] ), .B(\SUBBYTES[4].a/w2236 ), .Z(
        \SUBBYTES[4].a/w2264 ) );
  XOR U6720 ( .A(\w0[4][40] ), .B(g_input[552]), .Z(\w1[4][40] ) );
  AND U6721 ( .A(\SUBBYTES[4].a/w2237 ), .B(\SUBBYTES[4].a/w2233 ), .Z(
        \SUBBYTES[4].a/w2262 ) );
  AND U6722 ( .A(\SUBBYTES[4].a/w2322 ), .B(\SUBBYTES[4].a/w2354 ), .Z(
        \SUBBYTES[4].a/w2261 ) );
  ANDN U6723 ( .A(\SUBBYTES[4].a/w2343 ), .B(n2419), .Z(\SUBBYTES[4].a/w2256 )
         );
  XNOR U6724 ( .A(\w1[4][44] ), .B(\w1[4][47] ), .Z(n2419) );
  ANDN U6725 ( .A(\SUBBYTES[4].a/w2344 ), .B(n2420), .Z(\SUBBYTES[4].a/w2254 )
         );
  XNOR U6726 ( .A(\w1[4][42] ), .B(\w1[4][47] ), .Z(n2420) );
  XOR U6727 ( .A(\w0[4][47] ), .B(g_input[559]), .Z(\w1[4][47] ) );
  IV U6728 ( .A(n2422), .Z(\w1[4][42] ) );
  ANDN U6729 ( .A(\SUBBYTES[4].a/w2346 ), .B(n2421), .Z(\SUBBYTES[4].a/w2253 )
         );
  XOR U6730 ( .A(n2422), .B(\w1[4][44] ), .Z(n2421) );
  XOR U6731 ( .A(\w0[4][44] ), .B(g_input[556]), .Z(\w1[4][44] ) );
  XNOR U6732 ( .A(\w0[4][42] ), .B(g_input[554]), .Z(n2422) );
  AND U6733 ( .A(\SUBBYTES[4].a/w224 ), .B(\SUBBYTES[4].a/w230 ), .Z(
        \SUBBYTES[4].a/w225 ) );
  AND U6734 ( .A(\SUBBYTES[4].a/w209 ), .B(\SUBBYTES[4].a/w207 ), .Z(
        \SUBBYTES[4].a/w219 ) );
  AND U6735 ( .A(\SUBBYTES[4].a/w210 ), .B(\SUBBYTES[4].a/w208 ), .Z(
        \SUBBYTES[4].a/w217 ) );
  AND U6736 ( .A(\SUBBYTES[4].a/w224 ), .B(\SUBBYTES[4].a/w231 ), .Z(
        \SUBBYTES[4].a/w216 ) );
  AND U6737 ( .A(n2423), .B(\SUBBYTES[4].a/w2023 ), .Z(\SUBBYTES[4].a/w2158 )
         );
  AND U6738 ( .A(n2424), .B(\SUBBYTES[4].a/w2024 ), .Z(\SUBBYTES[4].a/w2156 )
         );
  AND U6739 ( .A(\SUBBYTES[4].a/w2154 ), .B(n2425), .Z(\SUBBYTES[4].a/w2155 )
         );
  ANDN U6740 ( .A(\w1[4][48] ), .B(n2426), .Z(\SUBBYTES[4].a/w2151 ) );
  AND U6741 ( .A(n2427), .B(\SUBBYTES[4].a/w2026 ), .Z(\SUBBYTES[4].a/w2149 )
         );
  AND U6742 ( .A(\SUBBYTES[4].a/w2147 ), .B(n2428), .Z(\SUBBYTES[4].a/w2148 )
         );
  XOR U6743 ( .A(\SUBBYTES[4].a/w2091 ), .B(n9690), .Z(n2428) );
  AND U6744 ( .A(\SUBBYTES[4].a/w2134 ), .B(\SUBBYTES[4].a/w2136 ), .Z(
        \SUBBYTES[4].a/w2143 ) );
  AND U6745 ( .A(\SUBBYTES[4].a/w2135 ), .B(\SUBBYTES[4].a/w2137 ), .Z(
        \SUBBYTES[4].a/w2141 ) );
  AND U6746 ( .A(\SUBBYTES[4].a/w2138 ), .B(\SUBBYTES[4].a/w2139 ), .Z(
        \SUBBYTES[4].a/w2140 ) );
  AND U6747 ( .A(\SUBBYTES[4].a/w2027 ), .B(n2423), .Z(\SUBBYTES[4].a/w2126 )
         );
  XOR U6748 ( .A(\SUBBYTES[4].a/w2095 ), .B(n1014), .Z(n2423) );
  AND U6749 ( .A(\SUBBYTES[4].a/w2028 ), .B(n2424), .Z(\SUBBYTES[4].a/w2124 )
         );
  XOR U6750 ( .A(n9691), .B(\SUBBYTES[4].a/w2095 ), .Z(n2424) );
  ANDN U6751 ( .A(n2425), .B(n2429), .Z(\SUBBYTES[4].a/w2123 ) );
  XOR U6752 ( .A(n1014), .B(n9691), .Z(n2425) );
  ANDN U6753 ( .A(\SUBBYTES[4].a/w2029 ), .B(n2426), .Z(\SUBBYTES[4].a/w2119 )
         );
  XNOR U6754 ( .A(\SUBBYTES[4].a/w2088 ), .B(\SUBBYTES[4].a/w2091 ), .Z(n2426)
         );
  AND U6755 ( .A(\SUBBYTES[4].a/w2030 ), .B(n2427), .Z(\SUBBYTES[4].a/w2117 )
         );
  XNOR U6756 ( .A(n2430), .B(\SUBBYTES[4].a/w2088 ), .Z(n2427) );
  AND U6757 ( .A(\SUBBYTES[4].a/w2115 ), .B(n2431), .Z(\SUBBYTES[4].a/w2116 )
         );
  XOR U6758 ( .A(n2432), .B(n2430), .Z(n2431) );
  IV U6759 ( .A(n9690), .Z(n2430) );
  ANDN U6760 ( .A(\SUBBYTES[4].a/w2134 ), .B(n2433), .Z(\SUBBYTES[4].a/w2111 )
         );
  ANDN U6761 ( .A(\SUBBYTES[4].a/w2135 ), .B(n2434), .Z(\SUBBYTES[4].a/w2109 )
         );
  ANDN U6762 ( .A(\SUBBYTES[4].a/w2138 ), .B(n2435), .Z(\SUBBYTES[4].a/w2108 )
         );
  AND U6763 ( .A(\SUBBYTES[4].a/w2094 ), .B(\SUBBYTES[4].a/w2093 ), .Z(
        \SUBBYTES[4].a/w2095 ) );
  IV U6764 ( .A(n2432), .Z(\SUBBYTES[4].a/w2091 ) );
  NAND U6765 ( .A(\SUBBYTES[4].a/w2070 ), .B(\SUBBYTES[4].a/w2085 ), .Z(n2432)
         );
  AND U6766 ( .A(\SUBBYTES[4].a/w2087 ), .B(\SUBBYTES[4].a/w2093 ), .Z(
        \SUBBYTES[4].a/w2088 ) );
  AND U6767 ( .A(\SUBBYTES[4].a/w2072 ), .B(\SUBBYTES[4].a/w2070 ), .Z(
        \SUBBYTES[4].a/w2082 ) );
  AND U6768 ( .A(\SUBBYTES[4].a/w2073 ), .B(\SUBBYTES[4].a/w2071 ), .Z(
        \SUBBYTES[4].a/w2080 ) );
  AND U6769 ( .A(\SUBBYTES[4].a/w2087 ), .B(\SUBBYTES[4].a/w2094 ), .Z(
        \SUBBYTES[4].a/w2079 ) );
  AND U6770 ( .A(\SUBBYTES[4].a/w2027 ), .B(\SUBBYTES[4].a/w2023 ), .Z(
        \SUBBYTES[4].a/w2064 ) );
  AND U6771 ( .A(\SUBBYTES[4].a/w2028 ), .B(\SUBBYTES[4].a/w2024 ), .Z(
        \SUBBYTES[4].a/w2062 ) );
  ANDN U6772 ( .A(\SUBBYTES[4].a/w2154 ), .B(n2429), .Z(\SUBBYTES[4].a/w2061 )
         );
  XNOR U6773 ( .A(\w1[4][49] ), .B(\w1[4][55] ), .Z(n2429) );
  XOR U6774 ( .A(\w0[4][49] ), .B(g_input[561]), .Z(\w1[4][49] ) );
  AND U6775 ( .A(\w1[4][48] ), .B(\SUBBYTES[4].a/w2029 ), .Z(
        \SUBBYTES[4].a/w2057 ) );
  XOR U6776 ( .A(\w0[4][48] ), .B(g_input[560]), .Z(\w1[4][48] ) );
  AND U6777 ( .A(\SUBBYTES[4].a/w2030 ), .B(\SUBBYTES[4].a/w2026 ), .Z(
        \SUBBYTES[4].a/w2055 ) );
  AND U6778 ( .A(\SUBBYTES[4].a/w2115 ), .B(\SUBBYTES[4].a/w2147 ), .Z(
        \SUBBYTES[4].a/w2054 ) );
  ANDN U6779 ( .A(\SUBBYTES[4].a/w2136 ), .B(n2433), .Z(\SUBBYTES[4].a/w2049 )
         );
  XNOR U6780 ( .A(\w1[4][52] ), .B(\w1[4][55] ), .Z(n2433) );
  ANDN U6781 ( .A(\SUBBYTES[4].a/w2137 ), .B(n2434), .Z(\SUBBYTES[4].a/w2047 )
         );
  XNOR U6782 ( .A(\w1[4][50] ), .B(\w1[4][55] ), .Z(n2434) );
  XOR U6783 ( .A(\w0[4][55] ), .B(g_input[567]), .Z(\w1[4][55] ) );
  IV U6784 ( .A(n2436), .Z(\w1[4][50] ) );
  ANDN U6785 ( .A(\SUBBYTES[4].a/w2139 ), .B(n2435), .Z(\SUBBYTES[4].a/w2046 )
         );
  XOR U6786 ( .A(n2436), .B(\w1[4][52] ), .Z(n2435) );
  XOR U6787 ( .A(\w0[4][52] ), .B(g_input[564]), .Z(\w1[4][52] ) );
  XNOR U6788 ( .A(\w0[4][50] ), .B(g_input[562]), .Z(n2436) );
  AND U6789 ( .A(\SUBBYTES[4].a/w164 ), .B(\SUBBYTES[4].a/w160 ), .Z(
        \SUBBYTES[4].a/w201 ) );
  AND U6790 ( .A(\SUBBYTES[4].a/w165 ), .B(\SUBBYTES[4].a/w161 ), .Z(
        \SUBBYTES[4].a/w199 ) );
  ANDN U6791 ( .A(\SUBBYTES[4].a/w291 ), .B(n2388), .Z(\SUBBYTES[4].a/w198 )
         );
  XNOR U6792 ( .A(\w1[4][121] ), .B(\w1[4][127] ), .Z(n2388) );
  XOR U6793 ( .A(\w0[4][121] ), .B(g_input[633]), .Z(\w1[4][121] ) );
  AND U6794 ( .A(n2437), .B(\SUBBYTES[4].a/w1816 ), .Z(\SUBBYTES[4].a/w1951 )
         );
  AND U6795 ( .A(n2438), .B(\SUBBYTES[4].a/w1817 ), .Z(\SUBBYTES[4].a/w1949 )
         );
  AND U6796 ( .A(\SUBBYTES[4].a/w1947 ), .B(n2439), .Z(\SUBBYTES[4].a/w1948 )
         );
  ANDN U6797 ( .A(\w1[4][56] ), .B(n2440), .Z(\SUBBYTES[4].a/w1944 ) );
  AND U6798 ( .A(n2441), .B(\SUBBYTES[4].a/w1819 ), .Z(\SUBBYTES[4].a/w1942 )
         );
  AND U6799 ( .A(\SUBBYTES[4].a/w1940 ), .B(n2442), .Z(\SUBBYTES[4].a/w1941 )
         );
  XOR U6800 ( .A(\SUBBYTES[4].a/w1884 ), .B(n9688), .Z(n2442) );
  AND U6801 ( .A(\w1[4][120] ), .B(\SUBBYTES[4].a/w166 ), .Z(
        \SUBBYTES[4].a/w194 ) );
  XOR U6802 ( .A(\w0[4][120] ), .B(g_input[632]), .Z(\w1[4][120] ) );
  AND U6803 ( .A(\SUBBYTES[4].a/w1927 ), .B(\SUBBYTES[4].a/w1929 ), .Z(
        \SUBBYTES[4].a/w1936 ) );
  AND U6804 ( .A(\SUBBYTES[4].a/w1928 ), .B(\SUBBYTES[4].a/w1930 ), .Z(
        \SUBBYTES[4].a/w1934 ) );
  AND U6805 ( .A(\SUBBYTES[4].a/w1931 ), .B(\SUBBYTES[4].a/w1932 ), .Z(
        \SUBBYTES[4].a/w1933 ) );
  AND U6806 ( .A(\SUBBYTES[4].a/w167 ), .B(\SUBBYTES[4].a/w163 ), .Z(
        \SUBBYTES[4].a/w192 ) );
  AND U6807 ( .A(\SUBBYTES[4].a/w1820 ), .B(n2437), .Z(\SUBBYTES[4].a/w1919 )
         );
  XOR U6808 ( .A(\SUBBYTES[4].a/w1888 ), .B(n1013), .Z(n2437) );
  AND U6809 ( .A(\SUBBYTES[4].a/w1821 ), .B(n2438), .Z(\SUBBYTES[4].a/w1917 )
         );
  XOR U6810 ( .A(n9689), .B(\SUBBYTES[4].a/w1888 ), .Z(n2438) );
  ANDN U6811 ( .A(n2439), .B(n2443), .Z(\SUBBYTES[4].a/w1916 ) );
  XOR U6812 ( .A(n1013), .B(n9689), .Z(n2439) );
  ANDN U6813 ( .A(\SUBBYTES[4].a/w1822 ), .B(n2440), .Z(\SUBBYTES[4].a/w1912 )
         );
  XNOR U6814 ( .A(\SUBBYTES[4].a/w1881 ), .B(\SUBBYTES[4].a/w1884 ), .Z(n2440)
         );
  AND U6815 ( .A(\SUBBYTES[4].a/w1823 ), .B(n2441), .Z(\SUBBYTES[4].a/w1910 )
         );
  XNOR U6816 ( .A(n2444), .B(\SUBBYTES[4].a/w1881 ), .Z(n2441) );
  AND U6817 ( .A(\SUBBYTES[4].a/w252 ), .B(\SUBBYTES[4].a/w284 ), .Z(
        \SUBBYTES[4].a/w191 ) );
  AND U6818 ( .A(\SUBBYTES[4].a/w1908 ), .B(n2445), .Z(\SUBBYTES[4].a/w1909 )
         );
  XOR U6819 ( .A(n2446), .B(n2444), .Z(n2445) );
  IV U6820 ( .A(n9688), .Z(n2444) );
  ANDN U6821 ( .A(\SUBBYTES[4].a/w1927 ), .B(n2447), .Z(\SUBBYTES[4].a/w1904 )
         );
  ANDN U6822 ( .A(\SUBBYTES[4].a/w1928 ), .B(n2448), .Z(\SUBBYTES[4].a/w1902 )
         );
  ANDN U6823 ( .A(\SUBBYTES[4].a/w1931 ), .B(n2449), .Z(\SUBBYTES[4].a/w1901 )
         );
  AND U6824 ( .A(\SUBBYTES[4].a/w1887 ), .B(\SUBBYTES[4].a/w1886 ), .Z(
        \SUBBYTES[4].a/w1888 ) );
  IV U6825 ( .A(n2446), .Z(\SUBBYTES[4].a/w1884 ) );
  NAND U6826 ( .A(\SUBBYTES[4].a/w1863 ), .B(\SUBBYTES[4].a/w1878 ), .Z(n2446)
         );
  AND U6827 ( .A(\SUBBYTES[4].a/w1880 ), .B(\SUBBYTES[4].a/w1886 ), .Z(
        \SUBBYTES[4].a/w1881 ) );
  AND U6828 ( .A(\SUBBYTES[4].a/w1865 ), .B(\SUBBYTES[4].a/w1863 ), .Z(
        \SUBBYTES[4].a/w1875 ) );
  AND U6829 ( .A(\SUBBYTES[4].a/w1866 ), .B(\SUBBYTES[4].a/w1864 ), .Z(
        \SUBBYTES[4].a/w1873 ) );
  AND U6830 ( .A(\SUBBYTES[4].a/w1880 ), .B(\SUBBYTES[4].a/w1887 ), .Z(
        \SUBBYTES[4].a/w1872 ) );
  ANDN U6831 ( .A(\SUBBYTES[4].a/w273 ), .B(n2405), .Z(\SUBBYTES[4].a/w186 )
         );
  XNOR U6832 ( .A(\w1[4][124] ), .B(\w1[4][127] ), .Z(n2405) );
  AND U6833 ( .A(\SUBBYTES[4].a/w1820 ), .B(\SUBBYTES[4].a/w1816 ), .Z(
        \SUBBYTES[4].a/w1857 ) );
  AND U6834 ( .A(\SUBBYTES[4].a/w1821 ), .B(\SUBBYTES[4].a/w1817 ), .Z(
        \SUBBYTES[4].a/w1855 ) );
  ANDN U6835 ( .A(\SUBBYTES[4].a/w1947 ), .B(n2443), .Z(\SUBBYTES[4].a/w1854 )
         );
  XNOR U6836 ( .A(\w1[4][57] ), .B(\w1[4][63] ), .Z(n2443) );
  XOR U6837 ( .A(\w0[4][57] ), .B(g_input[569]), .Z(\w1[4][57] ) );
  AND U6838 ( .A(\w1[4][56] ), .B(\SUBBYTES[4].a/w1822 ), .Z(
        \SUBBYTES[4].a/w1850 ) );
  XOR U6839 ( .A(\w0[4][56] ), .B(g_input[568]), .Z(\w1[4][56] ) );
  AND U6840 ( .A(\SUBBYTES[4].a/w1823 ), .B(\SUBBYTES[4].a/w1819 ), .Z(
        \SUBBYTES[4].a/w1848 ) );
  AND U6841 ( .A(\SUBBYTES[4].a/w1908 ), .B(\SUBBYTES[4].a/w1940 ), .Z(
        \SUBBYTES[4].a/w1847 ) );
  ANDN U6842 ( .A(\SUBBYTES[4].a/w1929 ), .B(n2447), .Z(\SUBBYTES[4].a/w1842 )
         );
  XNOR U6843 ( .A(\w1[4][60] ), .B(\w1[4][63] ), .Z(n2447) );
  ANDN U6844 ( .A(\SUBBYTES[4].a/w1930 ), .B(n2448), .Z(\SUBBYTES[4].a/w1840 )
         );
  XNOR U6845 ( .A(\w1[4][58] ), .B(\w1[4][63] ), .Z(n2448) );
  XOR U6846 ( .A(\w0[4][63] ), .B(g_input[575]), .Z(\w1[4][63] ) );
  IV U6847 ( .A(n2450), .Z(\w1[4][58] ) );
  ANDN U6848 ( .A(\SUBBYTES[4].a/w274 ), .B(n2407), .Z(\SUBBYTES[4].a/w184 )
         );
  XNOR U6849 ( .A(\w1[4][122] ), .B(\w1[4][127] ), .Z(n2407) );
  XOR U6850 ( .A(\w0[4][127] ), .B(g_input[639]), .Z(\w1[4][127] ) );
  IV U6851 ( .A(n2451), .Z(\w1[4][122] ) );
  ANDN U6852 ( .A(\SUBBYTES[4].a/w1932 ), .B(n2449), .Z(\SUBBYTES[4].a/w1839 )
         );
  XOR U6853 ( .A(n2450), .B(\w1[4][60] ), .Z(n2449) );
  XOR U6854 ( .A(\w0[4][60] ), .B(g_input[572]), .Z(\w1[4][60] ) );
  XNOR U6855 ( .A(\w0[4][58] ), .B(g_input[570]), .Z(n2450) );
  ANDN U6856 ( .A(\SUBBYTES[4].a/w276 ), .B(n2408), .Z(\SUBBYTES[4].a/w183 )
         );
  XOR U6857 ( .A(n2451), .B(\w1[4][124] ), .Z(n2408) );
  XOR U6858 ( .A(\w0[4][124] ), .B(g_input[636]), .Z(\w1[4][124] ) );
  XNOR U6859 ( .A(\w0[4][122] ), .B(g_input[634]), .Z(n2451) );
  AND U6860 ( .A(n2452), .B(\SUBBYTES[4].a/w1609 ), .Z(\SUBBYTES[4].a/w1744 )
         );
  AND U6861 ( .A(n2453), .B(\SUBBYTES[4].a/w1610 ), .Z(\SUBBYTES[4].a/w1742 )
         );
  AND U6862 ( .A(\SUBBYTES[4].a/w1740 ), .B(n2454), .Z(\SUBBYTES[4].a/w1741 )
         );
  ANDN U6863 ( .A(\w1[4][64] ), .B(n2455), .Z(\SUBBYTES[4].a/w1737 ) );
  AND U6864 ( .A(n2456), .B(\SUBBYTES[4].a/w1612 ), .Z(\SUBBYTES[4].a/w1735 )
         );
  AND U6865 ( .A(\SUBBYTES[4].a/w1733 ), .B(n2457), .Z(\SUBBYTES[4].a/w1734 )
         );
  XOR U6866 ( .A(\SUBBYTES[4].a/w1677 ), .B(n9686), .Z(n2457) );
  AND U6867 ( .A(\SUBBYTES[4].a/w1720 ), .B(\SUBBYTES[4].a/w1722 ), .Z(
        \SUBBYTES[4].a/w1729 ) );
  AND U6868 ( .A(\SUBBYTES[4].a/w1721 ), .B(\SUBBYTES[4].a/w1723 ), .Z(
        \SUBBYTES[4].a/w1727 ) );
  AND U6869 ( .A(\SUBBYTES[4].a/w1724 ), .B(\SUBBYTES[4].a/w1725 ), .Z(
        \SUBBYTES[4].a/w1726 ) );
  AND U6870 ( .A(\SUBBYTES[4].a/w1613 ), .B(n2452), .Z(\SUBBYTES[4].a/w1712 )
         );
  XOR U6871 ( .A(\SUBBYTES[4].a/w1681 ), .B(n1012), .Z(n2452) );
  AND U6872 ( .A(\SUBBYTES[4].a/w1614 ), .B(n2453), .Z(\SUBBYTES[4].a/w1710 )
         );
  XOR U6873 ( .A(n9687), .B(\SUBBYTES[4].a/w1681 ), .Z(n2453) );
  ANDN U6874 ( .A(n2454), .B(n2458), .Z(\SUBBYTES[4].a/w1709 ) );
  XOR U6875 ( .A(n1012), .B(n9687), .Z(n2454) );
  ANDN U6876 ( .A(\SUBBYTES[4].a/w1615 ), .B(n2455), .Z(\SUBBYTES[4].a/w1705 )
         );
  XNOR U6877 ( .A(\SUBBYTES[4].a/w1674 ), .B(\SUBBYTES[4].a/w1677 ), .Z(n2455)
         );
  AND U6878 ( .A(\SUBBYTES[4].a/w1616 ), .B(n2456), .Z(\SUBBYTES[4].a/w1703 )
         );
  XNOR U6879 ( .A(n2459), .B(\SUBBYTES[4].a/w1674 ), .Z(n2456) );
  AND U6880 ( .A(\SUBBYTES[4].a/w1701 ), .B(n2460), .Z(\SUBBYTES[4].a/w1702 )
         );
  XOR U6881 ( .A(n2461), .B(n2459), .Z(n2460) );
  IV U6882 ( .A(n9686), .Z(n2459) );
  ANDN U6883 ( .A(\SUBBYTES[4].a/w1720 ), .B(n2462), .Z(\SUBBYTES[4].a/w1697 )
         );
  ANDN U6884 ( .A(\SUBBYTES[4].a/w1721 ), .B(n2463), .Z(\SUBBYTES[4].a/w1695 )
         );
  ANDN U6885 ( .A(\SUBBYTES[4].a/w1724 ), .B(n2464), .Z(\SUBBYTES[4].a/w1694 )
         );
  AND U6886 ( .A(\SUBBYTES[4].a/w1680 ), .B(\SUBBYTES[4].a/w1679 ), .Z(
        \SUBBYTES[4].a/w1681 ) );
  IV U6887 ( .A(n2461), .Z(\SUBBYTES[4].a/w1677 ) );
  NAND U6888 ( .A(\SUBBYTES[4].a/w1656 ), .B(\SUBBYTES[4].a/w1671 ), .Z(n2461)
         );
  AND U6889 ( .A(\SUBBYTES[4].a/w1673 ), .B(\SUBBYTES[4].a/w1679 ), .Z(
        \SUBBYTES[4].a/w1674 ) );
  AND U6890 ( .A(\SUBBYTES[4].a/w1658 ), .B(\SUBBYTES[4].a/w1656 ), .Z(
        \SUBBYTES[4].a/w1668 ) );
  AND U6891 ( .A(\SUBBYTES[4].a/w1659 ), .B(\SUBBYTES[4].a/w1657 ), .Z(
        \SUBBYTES[4].a/w1666 ) );
  AND U6892 ( .A(\SUBBYTES[4].a/w1673 ), .B(\SUBBYTES[4].a/w1680 ), .Z(
        \SUBBYTES[4].a/w1665 ) );
  AND U6893 ( .A(\SUBBYTES[4].a/w1613 ), .B(\SUBBYTES[4].a/w1609 ), .Z(
        \SUBBYTES[4].a/w1650 ) );
  AND U6894 ( .A(\SUBBYTES[4].a/w1614 ), .B(\SUBBYTES[4].a/w1610 ), .Z(
        \SUBBYTES[4].a/w1648 ) );
  ANDN U6895 ( .A(\SUBBYTES[4].a/w1740 ), .B(n2458), .Z(\SUBBYTES[4].a/w1647 )
         );
  XNOR U6896 ( .A(\w1[4][65] ), .B(\w1[4][71] ), .Z(n2458) );
  XOR U6897 ( .A(\w0[4][65] ), .B(g_input[577]), .Z(\w1[4][65] ) );
  AND U6898 ( .A(\w1[4][64] ), .B(\SUBBYTES[4].a/w1615 ), .Z(
        \SUBBYTES[4].a/w1643 ) );
  XOR U6899 ( .A(\w0[4][64] ), .B(g_input[576]), .Z(\w1[4][64] ) );
  AND U6900 ( .A(\SUBBYTES[4].a/w1616 ), .B(\SUBBYTES[4].a/w1612 ), .Z(
        \SUBBYTES[4].a/w1641 ) );
  AND U6901 ( .A(\SUBBYTES[4].a/w1701 ), .B(\SUBBYTES[4].a/w1733 ), .Z(
        \SUBBYTES[4].a/w1640 ) );
  ANDN U6902 ( .A(\SUBBYTES[4].a/w1722 ), .B(n2462), .Z(\SUBBYTES[4].a/w1635 )
         );
  XNOR U6903 ( .A(\w1[4][68] ), .B(\w1[4][71] ), .Z(n2462) );
  ANDN U6904 ( .A(\SUBBYTES[4].a/w1723 ), .B(n2463), .Z(\SUBBYTES[4].a/w1633 )
         );
  XNOR U6905 ( .A(\w1[4][66] ), .B(\w1[4][71] ), .Z(n2463) );
  XOR U6906 ( .A(\w0[4][71] ), .B(g_input[583]), .Z(\w1[4][71] ) );
  IV U6907 ( .A(n2465), .Z(\w1[4][66] ) );
  ANDN U6908 ( .A(\SUBBYTES[4].a/w1725 ), .B(n2464), .Z(\SUBBYTES[4].a/w1632 )
         );
  XOR U6909 ( .A(n2465), .B(\w1[4][68] ), .Z(n2464) );
  XOR U6910 ( .A(\w0[4][68] ), .B(g_input[580]), .Z(\w1[4][68] ) );
  XNOR U6911 ( .A(\w0[4][66] ), .B(g_input[578]), .Z(n2465) );
  AND U6912 ( .A(n2466), .B(\SUBBYTES[4].a/w1402 ), .Z(\SUBBYTES[4].a/w1537 )
         );
  AND U6913 ( .A(n2467), .B(\SUBBYTES[4].a/w1403 ), .Z(\SUBBYTES[4].a/w1535 )
         );
  AND U6914 ( .A(\SUBBYTES[4].a/w1533 ), .B(n2468), .Z(\SUBBYTES[4].a/w1534 )
         );
  ANDN U6915 ( .A(\w1[4][72] ), .B(n2469), .Z(\SUBBYTES[4].a/w1530 ) );
  AND U6916 ( .A(n2470), .B(\SUBBYTES[4].a/w1405 ), .Z(\SUBBYTES[4].a/w1528 )
         );
  AND U6917 ( .A(\SUBBYTES[4].a/w1526 ), .B(n2471), .Z(\SUBBYTES[4].a/w1527 )
         );
  XOR U6918 ( .A(\SUBBYTES[4].a/w1470 ), .B(n9684), .Z(n2471) );
  AND U6919 ( .A(\SUBBYTES[4].a/w1513 ), .B(\SUBBYTES[4].a/w1515 ), .Z(
        \SUBBYTES[4].a/w1522 ) );
  AND U6920 ( .A(\SUBBYTES[4].a/w1514 ), .B(\SUBBYTES[4].a/w1516 ), .Z(
        \SUBBYTES[4].a/w1520 ) );
  AND U6921 ( .A(\SUBBYTES[4].a/w1517 ), .B(\SUBBYTES[4].a/w1518 ), .Z(
        \SUBBYTES[4].a/w1519 ) );
  AND U6922 ( .A(\SUBBYTES[4].a/w1406 ), .B(n2466), .Z(\SUBBYTES[4].a/w1505 )
         );
  XOR U6923 ( .A(\SUBBYTES[4].a/w1474 ), .B(n1011), .Z(n2466) );
  AND U6924 ( .A(\SUBBYTES[4].a/w1407 ), .B(n2467), .Z(\SUBBYTES[4].a/w1503 )
         );
  XOR U6925 ( .A(n9685), .B(\SUBBYTES[4].a/w1474 ), .Z(n2467) );
  ANDN U6926 ( .A(n2468), .B(n2472), .Z(\SUBBYTES[4].a/w1502 ) );
  XOR U6927 ( .A(n1011), .B(n9685), .Z(n2468) );
  ANDN U6928 ( .A(\SUBBYTES[4].a/w1408 ), .B(n2469), .Z(\SUBBYTES[4].a/w1498 )
         );
  XNOR U6929 ( .A(\SUBBYTES[4].a/w1467 ), .B(\SUBBYTES[4].a/w1470 ), .Z(n2469)
         );
  AND U6930 ( .A(\SUBBYTES[4].a/w1409 ), .B(n2470), .Z(\SUBBYTES[4].a/w1496 )
         );
  XNOR U6931 ( .A(n2473), .B(\SUBBYTES[4].a/w1467 ), .Z(n2470) );
  AND U6932 ( .A(\SUBBYTES[4].a/w1494 ), .B(n2474), .Z(\SUBBYTES[4].a/w1495 )
         );
  XOR U6933 ( .A(n2475), .B(n2473), .Z(n2474) );
  IV U6934 ( .A(n9684), .Z(n2473) );
  ANDN U6935 ( .A(\SUBBYTES[4].a/w1513 ), .B(n2476), .Z(\SUBBYTES[4].a/w1490 )
         );
  ANDN U6936 ( .A(\SUBBYTES[4].a/w1514 ), .B(n2477), .Z(\SUBBYTES[4].a/w1488 )
         );
  ANDN U6937 ( .A(\SUBBYTES[4].a/w1517 ), .B(n2478), .Z(\SUBBYTES[4].a/w1487 )
         );
  AND U6938 ( .A(\SUBBYTES[4].a/w1473 ), .B(\SUBBYTES[4].a/w1472 ), .Z(
        \SUBBYTES[4].a/w1474 ) );
  IV U6939 ( .A(n2475), .Z(\SUBBYTES[4].a/w1470 ) );
  NAND U6940 ( .A(\SUBBYTES[4].a/w1449 ), .B(\SUBBYTES[4].a/w1464 ), .Z(n2475)
         );
  AND U6941 ( .A(\SUBBYTES[4].a/w1466 ), .B(\SUBBYTES[4].a/w1472 ), .Z(
        \SUBBYTES[4].a/w1467 ) );
  AND U6942 ( .A(\SUBBYTES[4].a/w1451 ), .B(\SUBBYTES[4].a/w1449 ), .Z(
        \SUBBYTES[4].a/w1461 ) );
  AND U6943 ( .A(\SUBBYTES[4].a/w1452 ), .B(\SUBBYTES[4].a/w1450 ), .Z(
        \SUBBYTES[4].a/w1459 ) );
  AND U6944 ( .A(\SUBBYTES[4].a/w1466 ), .B(\SUBBYTES[4].a/w1473 ), .Z(
        \SUBBYTES[4].a/w1458 ) );
  AND U6945 ( .A(\SUBBYTES[4].a/w1406 ), .B(\SUBBYTES[4].a/w1402 ), .Z(
        \SUBBYTES[4].a/w1443 ) );
  AND U6946 ( .A(\SUBBYTES[4].a/w1407 ), .B(\SUBBYTES[4].a/w1403 ), .Z(
        \SUBBYTES[4].a/w1441 ) );
  ANDN U6947 ( .A(\SUBBYTES[4].a/w1533 ), .B(n2472), .Z(\SUBBYTES[4].a/w1440 )
         );
  XNOR U6948 ( .A(\w1[4][73] ), .B(\w1[4][79] ), .Z(n2472) );
  XOR U6949 ( .A(\w0[4][73] ), .B(g_input[585]), .Z(\w1[4][73] ) );
  AND U6950 ( .A(\w1[4][72] ), .B(\SUBBYTES[4].a/w1408 ), .Z(
        \SUBBYTES[4].a/w1436 ) );
  XOR U6951 ( .A(\w0[4][72] ), .B(g_input[584]), .Z(\w1[4][72] ) );
  AND U6952 ( .A(\SUBBYTES[4].a/w1409 ), .B(\SUBBYTES[4].a/w1405 ), .Z(
        \SUBBYTES[4].a/w1434 ) );
  AND U6953 ( .A(\SUBBYTES[4].a/w1494 ), .B(\SUBBYTES[4].a/w1526 ), .Z(
        \SUBBYTES[4].a/w1433 ) );
  ANDN U6954 ( .A(\SUBBYTES[4].a/w1515 ), .B(n2476), .Z(\SUBBYTES[4].a/w1428 )
         );
  XNOR U6955 ( .A(\w1[4][76] ), .B(\w1[4][79] ), .Z(n2476) );
  ANDN U6956 ( .A(\SUBBYTES[4].a/w1516 ), .B(n2477), .Z(\SUBBYTES[4].a/w1426 )
         );
  XNOR U6957 ( .A(\w1[4][74] ), .B(\w1[4][79] ), .Z(n2477) );
  XOR U6958 ( .A(\w0[4][79] ), .B(g_input[591]), .Z(\w1[4][79] ) );
  IV U6959 ( .A(n2479), .Z(\w1[4][74] ) );
  ANDN U6960 ( .A(\SUBBYTES[4].a/w1518 ), .B(n2478), .Z(\SUBBYTES[4].a/w1425 )
         );
  XOR U6961 ( .A(n2479), .B(\w1[4][76] ), .Z(n2478) );
  XOR U6962 ( .A(\w0[4][76] ), .B(g_input[588]), .Z(\w1[4][76] ) );
  XNOR U6963 ( .A(\w0[4][74] ), .B(g_input[586]), .Z(n2479) );
  AND U6964 ( .A(n2480), .B(\SUBBYTES[4].a/w1195 ), .Z(\SUBBYTES[4].a/w1330 )
         );
  AND U6965 ( .A(n2481), .B(\SUBBYTES[4].a/w1196 ), .Z(\SUBBYTES[4].a/w1328 )
         );
  AND U6966 ( .A(\SUBBYTES[4].a/w1326 ), .B(n2482), .Z(\SUBBYTES[4].a/w1327 )
         );
  ANDN U6967 ( .A(\w1[4][80] ), .B(n2483), .Z(\SUBBYTES[4].a/w1323 ) );
  AND U6968 ( .A(n2484), .B(\SUBBYTES[4].a/w1198 ), .Z(\SUBBYTES[4].a/w1321 )
         );
  AND U6969 ( .A(\SUBBYTES[4].a/w1319 ), .B(n2485), .Z(\SUBBYTES[4].a/w1320 )
         );
  XOR U6970 ( .A(\SUBBYTES[4].a/w1263 ), .B(n9682), .Z(n2485) );
  AND U6971 ( .A(\SUBBYTES[4].a/w1306 ), .B(\SUBBYTES[4].a/w1308 ), .Z(
        \SUBBYTES[4].a/w1315 ) );
  AND U6972 ( .A(\SUBBYTES[4].a/w1307 ), .B(\SUBBYTES[4].a/w1309 ), .Z(
        \SUBBYTES[4].a/w1313 ) );
  AND U6973 ( .A(\SUBBYTES[4].a/w1310 ), .B(\SUBBYTES[4].a/w1311 ), .Z(
        \SUBBYTES[4].a/w1312 ) );
  AND U6974 ( .A(\SUBBYTES[4].a/w1199 ), .B(n2480), .Z(\SUBBYTES[4].a/w1298 )
         );
  XOR U6975 ( .A(\SUBBYTES[4].a/w1267 ), .B(n1010), .Z(n2480) );
  AND U6976 ( .A(\SUBBYTES[4].a/w1200 ), .B(n2481), .Z(\SUBBYTES[4].a/w1296 )
         );
  XOR U6977 ( .A(n9683), .B(\SUBBYTES[4].a/w1267 ), .Z(n2481) );
  ANDN U6978 ( .A(n2482), .B(n2486), .Z(\SUBBYTES[4].a/w1295 ) );
  XOR U6979 ( .A(n1010), .B(n9683), .Z(n2482) );
  ANDN U6980 ( .A(\SUBBYTES[4].a/w1201 ), .B(n2483), .Z(\SUBBYTES[4].a/w1291 )
         );
  XNOR U6981 ( .A(\SUBBYTES[4].a/w1260 ), .B(\SUBBYTES[4].a/w1263 ), .Z(n2483)
         );
  AND U6982 ( .A(\SUBBYTES[4].a/w1202 ), .B(n2484), .Z(\SUBBYTES[4].a/w1289 )
         );
  XNOR U6983 ( .A(n2487), .B(\SUBBYTES[4].a/w1260 ), .Z(n2484) );
  AND U6984 ( .A(\SUBBYTES[4].a/w1287 ), .B(n2488), .Z(\SUBBYTES[4].a/w1288 )
         );
  XOR U6985 ( .A(n2489), .B(n2487), .Z(n2488) );
  IV U6986 ( .A(n9682), .Z(n2487) );
  ANDN U6987 ( .A(\SUBBYTES[4].a/w1306 ), .B(n2490), .Z(\SUBBYTES[4].a/w1283 )
         );
  ANDN U6988 ( .A(\SUBBYTES[4].a/w1307 ), .B(n2491), .Z(\SUBBYTES[4].a/w1281 )
         );
  ANDN U6989 ( .A(\SUBBYTES[4].a/w1310 ), .B(n2492), .Z(\SUBBYTES[4].a/w1280 )
         );
  AND U6990 ( .A(\SUBBYTES[4].a/w1266 ), .B(\SUBBYTES[4].a/w1265 ), .Z(
        \SUBBYTES[4].a/w1267 ) );
  IV U6991 ( .A(n2489), .Z(\SUBBYTES[4].a/w1263 ) );
  NAND U6992 ( .A(\SUBBYTES[4].a/w1242 ), .B(\SUBBYTES[4].a/w1257 ), .Z(n2489)
         );
  AND U6993 ( .A(\SUBBYTES[4].a/w1259 ), .B(\SUBBYTES[4].a/w1265 ), .Z(
        \SUBBYTES[4].a/w1260 ) );
  AND U6994 ( .A(\SUBBYTES[4].a/w1244 ), .B(\SUBBYTES[4].a/w1242 ), .Z(
        \SUBBYTES[4].a/w1254 ) );
  AND U6995 ( .A(\SUBBYTES[4].a/w1245 ), .B(\SUBBYTES[4].a/w1243 ), .Z(
        \SUBBYTES[4].a/w1252 ) );
  AND U6996 ( .A(\SUBBYTES[4].a/w1259 ), .B(\SUBBYTES[4].a/w1266 ), .Z(
        \SUBBYTES[4].a/w1251 ) );
  AND U6997 ( .A(\SUBBYTES[4].a/w1199 ), .B(\SUBBYTES[4].a/w1195 ), .Z(
        \SUBBYTES[4].a/w1236 ) );
  AND U6998 ( .A(\SUBBYTES[4].a/w1200 ), .B(\SUBBYTES[4].a/w1196 ), .Z(
        \SUBBYTES[4].a/w1234 ) );
  ANDN U6999 ( .A(\SUBBYTES[4].a/w1326 ), .B(n2486), .Z(\SUBBYTES[4].a/w1233 )
         );
  XNOR U7000 ( .A(\w1[4][81] ), .B(\w1[4][87] ), .Z(n2486) );
  XOR U7001 ( .A(\w0[4][81] ), .B(g_input[593]), .Z(\w1[4][81] ) );
  AND U7002 ( .A(\w1[4][80] ), .B(\SUBBYTES[4].a/w1201 ), .Z(
        \SUBBYTES[4].a/w1229 ) );
  XOR U7003 ( .A(\w0[4][80] ), .B(g_input[592]), .Z(\w1[4][80] ) );
  AND U7004 ( .A(\SUBBYTES[4].a/w1202 ), .B(\SUBBYTES[4].a/w1198 ), .Z(
        \SUBBYTES[4].a/w1227 ) );
  AND U7005 ( .A(\SUBBYTES[4].a/w1287 ), .B(\SUBBYTES[4].a/w1319 ), .Z(
        \SUBBYTES[4].a/w1226 ) );
  ANDN U7006 ( .A(\SUBBYTES[4].a/w1308 ), .B(n2490), .Z(\SUBBYTES[4].a/w1221 )
         );
  XNOR U7007 ( .A(\w1[4][84] ), .B(\w1[4][87] ), .Z(n2490) );
  ANDN U7008 ( .A(\SUBBYTES[4].a/w1309 ), .B(n2491), .Z(\SUBBYTES[4].a/w1219 )
         );
  XNOR U7009 ( .A(\w1[4][82] ), .B(\w1[4][87] ), .Z(n2491) );
  XOR U7010 ( .A(\w0[4][87] ), .B(g_input[599]), .Z(\w1[4][87] ) );
  IV U7011 ( .A(n2493), .Z(\w1[4][82] ) );
  ANDN U7012 ( .A(\SUBBYTES[4].a/w1311 ), .B(n2492), .Z(\SUBBYTES[4].a/w1218 )
         );
  XOR U7013 ( .A(n2493), .B(\w1[4][84] ), .Z(n2492) );
  XOR U7014 ( .A(\w0[4][84] ), .B(g_input[596]), .Z(\w1[4][84] ) );
  XNOR U7015 ( .A(\w0[4][82] ), .B(g_input[594]), .Z(n2493) );
  AND U7016 ( .A(n2494), .B(\SUBBYTES[4].a/w988 ), .Z(\SUBBYTES[4].a/w1123 )
         );
  AND U7017 ( .A(n2495), .B(\SUBBYTES[4].a/w989 ), .Z(\SUBBYTES[4].a/w1121 )
         );
  AND U7018 ( .A(\SUBBYTES[4].a/w1119 ), .B(n2496), .Z(\SUBBYTES[4].a/w1120 )
         );
  ANDN U7019 ( .A(\w1[4][88] ), .B(n2497), .Z(\SUBBYTES[4].a/w1116 ) );
  AND U7020 ( .A(n2498), .B(\SUBBYTES[4].a/w991 ), .Z(\SUBBYTES[4].a/w1114 )
         );
  AND U7021 ( .A(\SUBBYTES[4].a/w1112 ), .B(n2499), .Z(\SUBBYTES[4].a/w1113 )
         );
  XOR U7022 ( .A(\SUBBYTES[4].a/w1056 ), .B(n9680), .Z(n2499) );
  AND U7023 ( .A(\SUBBYTES[4].a/w1099 ), .B(\SUBBYTES[4].a/w1101 ), .Z(
        \SUBBYTES[4].a/w1108 ) );
  AND U7024 ( .A(\SUBBYTES[4].a/w1100 ), .B(\SUBBYTES[4].a/w1102 ), .Z(
        \SUBBYTES[4].a/w1106 ) );
  AND U7025 ( .A(\SUBBYTES[4].a/w1103 ), .B(\SUBBYTES[4].a/w1104 ), .Z(
        \SUBBYTES[4].a/w1105 ) );
  AND U7026 ( .A(\SUBBYTES[4].a/w992 ), .B(n2494), .Z(\SUBBYTES[4].a/w1091 )
         );
  XOR U7027 ( .A(\SUBBYTES[4].a/w1060 ), .B(n1009), .Z(n2494) );
  AND U7028 ( .A(\SUBBYTES[4].a/w993 ), .B(n2495), .Z(\SUBBYTES[4].a/w1089 )
         );
  XOR U7029 ( .A(n9681), .B(\SUBBYTES[4].a/w1060 ), .Z(n2495) );
  ANDN U7030 ( .A(n2496), .B(n2500), .Z(\SUBBYTES[4].a/w1088 ) );
  XOR U7031 ( .A(n1009), .B(n9681), .Z(n2496) );
  ANDN U7032 ( .A(\SUBBYTES[4].a/w994 ), .B(n2497), .Z(\SUBBYTES[4].a/w1084 )
         );
  XNOR U7033 ( .A(\SUBBYTES[4].a/w1053 ), .B(\SUBBYTES[4].a/w1056 ), .Z(n2497)
         );
  AND U7034 ( .A(\SUBBYTES[4].a/w995 ), .B(n2498), .Z(\SUBBYTES[4].a/w1082 )
         );
  XNOR U7035 ( .A(n2501), .B(\SUBBYTES[4].a/w1053 ), .Z(n2498) );
  AND U7036 ( .A(\SUBBYTES[4].a/w1080 ), .B(n2502), .Z(\SUBBYTES[4].a/w1081 )
         );
  XOR U7037 ( .A(n2503), .B(n2501), .Z(n2502) );
  IV U7038 ( .A(n9680), .Z(n2501) );
  ANDN U7039 ( .A(\SUBBYTES[4].a/w1099 ), .B(n2504), .Z(\SUBBYTES[4].a/w1076 )
         );
  ANDN U7040 ( .A(\SUBBYTES[4].a/w1100 ), .B(n2505), .Z(\SUBBYTES[4].a/w1074 )
         );
  ANDN U7041 ( .A(\SUBBYTES[4].a/w1103 ), .B(n2506), .Z(\SUBBYTES[4].a/w1073 )
         );
  AND U7042 ( .A(\SUBBYTES[4].a/w1059 ), .B(\SUBBYTES[4].a/w1058 ), .Z(
        \SUBBYTES[4].a/w1060 ) );
  IV U7043 ( .A(n2503), .Z(\SUBBYTES[4].a/w1056 ) );
  NAND U7044 ( .A(\SUBBYTES[4].a/w1035 ), .B(\SUBBYTES[4].a/w1050 ), .Z(n2503)
         );
  AND U7045 ( .A(\SUBBYTES[4].a/w1052 ), .B(\SUBBYTES[4].a/w1058 ), .Z(
        \SUBBYTES[4].a/w1053 ) );
  AND U7046 ( .A(\SUBBYTES[4].a/w1037 ), .B(\SUBBYTES[4].a/w1035 ), .Z(
        \SUBBYTES[4].a/w1047 ) );
  AND U7047 ( .A(\SUBBYTES[4].a/w1038 ), .B(\SUBBYTES[4].a/w1036 ), .Z(
        \SUBBYTES[4].a/w1045 ) );
  AND U7048 ( .A(\SUBBYTES[4].a/w1052 ), .B(\SUBBYTES[4].a/w1059 ), .Z(
        \SUBBYTES[4].a/w1044 ) );
  AND U7049 ( .A(\SUBBYTES[4].a/w992 ), .B(\SUBBYTES[4].a/w988 ), .Z(
        \SUBBYTES[4].a/w1029 ) );
  AND U7050 ( .A(\SUBBYTES[4].a/w993 ), .B(\SUBBYTES[4].a/w989 ), .Z(
        \SUBBYTES[4].a/w1027 ) );
  ANDN U7051 ( .A(\SUBBYTES[4].a/w1119 ), .B(n2500), .Z(\SUBBYTES[4].a/w1026 )
         );
  XNOR U7052 ( .A(\w1[4][89] ), .B(\w1[4][95] ), .Z(n2500) );
  XOR U7053 ( .A(\w0[4][89] ), .B(g_input[601]), .Z(\w1[4][89] ) );
  AND U7054 ( .A(\w1[4][88] ), .B(\SUBBYTES[4].a/w994 ), .Z(
        \SUBBYTES[4].a/w1022 ) );
  XOR U7055 ( .A(\w0[4][88] ), .B(g_input[600]), .Z(\w1[4][88] ) );
  AND U7056 ( .A(\SUBBYTES[4].a/w995 ), .B(\SUBBYTES[4].a/w991 ), .Z(
        \SUBBYTES[4].a/w1020 ) );
  AND U7057 ( .A(\SUBBYTES[4].a/w1080 ), .B(\SUBBYTES[4].a/w1112 ), .Z(
        \SUBBYTES[4].a/w1019 ) );
  ANDN U7058 ( .A(\SUBBYTES[4].a/w1101 ), .B(n2504), .Z(\SUBBYTES[4].a/w1014 )
         );
  XNOR U7059 ( .A(\w1[4][92] ), .B(\w1[4][95] ), .Z(n2504) );
  ANDN U7060 ( .A(\SUBBYTES[4].a/w1102 ), .B(n2505), .Z(\SUBBYTES[4].a/w1012 )
         );
  XNOR U7061 ( .A(\w1[4][90] ), .B(\w1[4][95] ), .Z(n2505) );
  XOR U7062 ( .A(\w0[4][95] ), .B(g_input[607]), .Z(\w1[4][95] ) );
  IV U7063 ( .A(n2507), .Z(\w1[4][90] ) );
  ANDN U7064 ( .A(\SUBBYTES[4].a/w1104 ), .B(n2506), .Z(\SUBBYTES[4].a/w1011 )
         );
  XOR U7065 ( .A(n2507), .B(\w1[4][92] ), .Z(n2506) );
  XOR U7066 ( .A(\w0[4][92] ), .B(g_input[604]), .Z(\w1[4][92] ) );
  XNOR U7067 ( .A(\w0[4][90] ), .B(g_input[602]), .Z(n2507) );
  AND U7068 ( .A(\SUBBYTES[4].a/w2084 ), .B(\SUBBYTES[4].a/w2071 ), .Z(n9690)
         );
  AND U7069 ( .A(\SUBBYTES[4].a/w1877 ), .B(\SUBBYTES[4].a/w1866 ), .Z(n9689)
         );
  AND U7070 ( .A(\SUBBYTES[4].a/w221 ), .B(\SUBBYTES[4].a/w208 ), .Z(n9672) );
  AND U7071 ( .A(\SUBBYTES[4].a/w1877 ), .B(\SUBBYTES[4].a/w1864 ), .Z(n9688)
         );
  AND U7072 ( .A(\SUBBYTES[4].a/w1670 ), .B(\SUBBYTES[4].a/w1659 ), .Z(n9687)
         );
  AND U7073 ( .A(\SUBBYTES[4].a/w1670 ), .B(\SUBBYTES[4].a/w1657 ), .Z(n9686)
         );
  AND U7074 ( .A(\SUBBYTES[4].a/w1463 ), .B(\SUBBYTES[4].a/w1452 ), .Z(n9685)
         );
  AND U7075 ( .A(\SUBBYTES[4].a/w1463 ), .B(\SUBBYTES[4].a/w1450 ), .Z(n9684)
         );
  AND U7076 ( .A(\SUBBYTES[4].a/w1256 ), .B(\SUBBYTES[4].a/w1245 ), .Z(n9683)
         );
  AND U7077 ( .A(\SUBBYTES[4].a/w1256 ), .B(\SUBBYTES[4].a/w1243 ), .Z(n9682)
         );
  AND U7078 ( .A(\SUBBYTES[4].a/w1049 ), .B(\SUBBYTES[4].a/w1038 ), .Z(n9681)
         );
  AND U7079 ( .A(\SUBBYTES[4].a/w1049 ), .B(\SUBBYTES[4].a/w1036 ), .Z(n9680)
         );
  AND U7080 ( .A(\SUBBYTES[4].a/w842 ), .B(\SUBBYTES[4].a/w831 ), .Z(n9679) );
  AND U7081 ( .A(\SUBBYTES[4].a/w842 ), .B(\SUBBYTES[4].a/w829 ), .Z(n9678) );
  AND U7082 ( .A(\SUBBYTES[4].a/w635 ), .B(\SUBBYTES[4].a/w624 ), .Z(n9677) );
  AND U7083 ( .A(\SUBBYTES[4].a/w635 ), .B(\SUBBYTES[4].a/w622 ), .Z(n9676) );
  AND U7084 ( .A(\SUBBYTES[4].a/w428 ), .B(\SUBBYTES[4].a/w417 ), .Z(n9675) );
  AND U7085 ( .A(\SUBBYTES[4].a/w428 ), .B(\SUBBYTES[4].a/w415 ), .Z(n9674) );
  AND U7086 ( .A(\SUBBYTES[4].a/w3326 ), .B(\SUBBYTES[4].a/w3315 ), .Z(n9703)
         );
  AND U7087 ( .A(\SUBBYTES[4].a/w3326 ), .B(\SUBBYTES[4].a/w3313 ), .Z(n9702)
         );
  AND U7088 ( .A(\SUBBYTES[4].a/w3119 ), .B(\SUBBYTES[4].a/w3108 ), .Z(n9701)
         );
  AND U7089 ( .A(\SUBBYTES[4].a/w3119 ), .B(\SUBBYTES[4].a/w3106 ), .Z(n9700)
         );
  AND U7090 ( .A(\SUBBYTES[4].a/w2912 ), .B(\SUBBYTES[4].a/w2901 ), .Z(n9699)
         );
  AND U7091 ( .A(\SUBBYTES[4].a/w2912 ), .B(\SUBBYTES[4].a/w2899 ), .Z(n9698)
         );
  AND U7092 ( .A(\SUBBYTES[4].a/w2705 ), .B(\SUBBYTES[4].a/w2694 ), .Z(n9697)
         );
  AND U7093 ( .A(\SUBBYTES[4].a/w2705 ), .B(\SUBBYTES[4].a/w2692 ), .Z(n9696)
         );
  AND U7094 ( .A(\SUBBYTES[4].a/w2498 ), .B(\SUBBYTES[4].a/w2487 ), .Z(n9695)
         );
  AND U7095 ( .A(\SUBBYTES[4].a/w2498 ), .B(\SUBBYTES[4].a/w2485 ), .Z(n9694)
         );
  AND U7096 ( .A(\SUBBYTES[4].a/w2291 ), .B(\SUBBYTES[4].a/w2280 ), .Z(n9693)
         );
  AND U7097 ( .A(\SUBBYTES[4].a/w2291 ), .B(\SUBBYTES[4].a/w2278 ), .Z(n9692)
         );
  AND U7098 ( .A(\SUBBYTES[4].a/w2084 ), .B(\SUBBYTES[4].a/w2073 ), .Z(n9691)
         );
  AND U7099 ( .A(\SUBBYTES[4].a/w221 ), .B(\SUBBYTES[4].a/w210 ), .Z(n9673) );
  AND U7100 ( .A(n2508), .B(\SUBBYTES[3].a/w781 ), .Z(\SUBBYTES[3].a/w916 ) );
  AND U7101 ( .A(n2509), .B(\SUBBYTES[3].a/w782 ), .Z(\SUBBYTES[3].a/w914 ) );
  AND U7102 ( .A(\SUBBYTES[3].a/w912 ), .B(n2510), .Z(\SUBBYTES[3].a/w913 ) );
  ANDN U7103 ( .A(\w1[3][96] ), .B(n2511), .Z(\SUBBYTES[3].a/w909 ) );
  AND U7104 ( .A(n2512), .B(\SUBBYTES[3].a/w784 ), .Z(\SUBBYTES[3].a/w907 ) );
  AND U7105 ( .A(\SUBBYTES[3].a/w905 ), .B(n2513), .Z(\SUBBYTES[3].a/w906 ) );
  XOR U7106 ( .A(\SUBBYTES[3].a/w849 ), .B(n8398), .Z(n2513) );
  AND U7107 ( .A(\SUBBYTES[3].a/w892 ), .B(\SUBBYTES[3].a/w894 ), .Z(
        \SUBBYTES[3].a/w901 ) );
  AND U7108 ( .A(\SUBBYTES[3].a/w893 ), .B(\SUBBYTES[3].a/w895 ), .Z(
        \SUBBYTES[3].a/w899 ) );
  AND U7109 ( .A(\SUBBYTES[3].a/w896 ), .B(\SUBBYTES[3].a/w897 ), .Z(
        \SUBBYTES[3].a/w898 ) );
  AND U7110 ( .A(\SUBBYTES[3].a/w785 ), .B(n2508), .Z(\SUBBYTES[3].a/w884 ) );
  XOR U7111 ( .A(\SUBBYTES[3].a/w853 ), .B(n992), .Z(n2508) );
  AND U7112 ( .A(\SUBBYTES[3].a/w786 ), .B(n2509), .Z(\SUBBYTES[3].a/w882 ) );
  XOR U7113 ( .A(n8399), .B(\SUBBYTES[3].a/w853 ), .Z(n2509) );
  ANDN U7114 ( .A(n2510), .B(n2514), .Z(\SUBBYTES[3].a/w881 ) );
  XOR U7115 ( .A(n992), .B(n8399), .Z(n2510) );
  ANDN U7116 ( .A(\SUBBYTES[3].a/w787 ), .B(n2511), .Z(\SUBBYTES[3].a/w877 )
         );
  XNOR U7117 ( .A(\SUBBYTES[3].a/w846 ), .B(\SUBBYTES[3].a/w849 ), .Z(n2511)
         );
  AND U7118 ( .A(\SUBBYTES[3].a/w788 ), .B(n2512), .Z(\SUBBYTES[3].a/w875 ) );
  XNOR U7119 ( .A(n2515), .B(\SUBBYTES[3].a/w846 ), .Z(n2512) );
  AND U7120 ( .A(\SUBBYTES[3].a/w873 ), .B(n2516), .Z(\SUBBYTES[3].a/w874 ) );
  XOR U7121 ( .A(n2517), .B(n2515), .Z(n2516) );
  IV U7122 ( .A(n8398), .Z(n2515) );
  ANDN U7123 ( .A(\SUBBYTES[3].a/w892 ), .B(n2518), .Z(\SUBBYTES[3].a/w869 )
         );
  ANDN U7124 ( .A(\SUBBYTES[3].a/w893 ), .B(n2519), .Z(\SUBBYTES[3].a/w867 )
         );
  ANDN U7125 ( .A(\SUBBYTES[3].a/w896 ), .B(n2520), .Z(\SUBBYTES[3].a/w866 )
         );
  AND U7126 ( .A(\SUBBYTES[3].a/w852 ), .B(\SUBBYTES[3].a/w851 ), .Z(
        \SUBBYTES[3].a/w853 ) );
  IV U7127 ( .A(n2517), .Z(\SUBBYTES[3].a/w849 ) );
  NAND U7128 ( .A(\SUBBYTES[3].a/w828 ), .B(\SUBBYTES[3].a/w843 ), .Z(n2517)
         );
  AND U7129 ( .A(\SUBBYTES[3].a/w845 ), .B(\SUBBYTES[3].a/w851 ), .Z(
        \SUBBYTES[3].a/w846 ) );
  AND U7130 ( .A(\SUBBYTES[3].a/w830 ), .B(\SUBBYTES[3].a/w828 ), .Z(
        \SUBBYTES[3].a/w840 ) );
  AND U7131 ( .A(\SUBBYTES[3].a/w831 ), .B(\SUBBYTES[3].a/w829 ), .Z(
        \SUBBYTES[3].a/w838 ) );
  AND U7132 ( .A(\SUBBYTES[3].a/w845 ), .B(\SUBBYTES[3].a/w852 ), .Z(
        \SUBBYTES[3].a/w837 ) );
  AND U7133 ( .A(\SUBBYTES[3].a/w785 ), .B(\SUBBYTES[3].a/w781 ), .Z(
        \SUBBYTES[3].a/w822 ) );
  AND U7134 ( .A(\SUBBYTES[3].a/w786 ), .B(\SUBBYTES[3].a/w782 ), .Z(
        \SUBBYTES[3].a/w820 ) );
  ANDN U7135 ( .A(\SUBBYTES[3].a/w912 ), .B(n2514), .Z(\SUBBYTES[3].a/w819 )
         );
  XNOR U7136 ( .A(\w1[3][103] ), .B(\w1[3][97] ), .Z(n2514) );
  XOR U7137 ( .A(\w0[3][97] ), .B(g_input[481]), .Z(\w1[3][97] ) );
  IV U7138 ( .A(n2521), .Z(\w1[3][103] ) );
  AND U7139 ( .A(\w1[3][96] ), .B(\SUBBYTES[3].a/w787 ), .Z(
        \SUBBYTES[3].a/w815 ) );
  XOR U7140 ( .A(\w0[3][96] ), .B(g_input[480]), .Z(\w1[3][96] ) );
  AND U7141 ( .A(\SUBBYTES[3].a/w788 ), .B(\SUBBYTES[3].a/w784 ), .Z(
        \SUBBYTES[3].a/w813 ) );
  AND U7142 ( .A(\SUBBYTES[3].a/w873 ), .B(\SUBBYTES[3].a/w905 ), .Z(
        \SUBBYTES[3].a/w812 ) );
  ANDN U7143 ( .A(\SUBBYTES[3].a/w894 ), .B(n2518), .Z(\SUBBYTES[3].a/w807 )
         );
  XOR U7144 ( .A(\w1[3][100] ), .B(n2521), .Z(n2518) );
  ANDN U7145 ( .A(\SUBBYTES[3].a/w895 ), .B(n2519), .Z(\SUBBYTES[3].a/w805 )
         );
  XOR U7146 ( .A(n2521), .B(\w1[3][98] ), .Z(n2519) );
  XNOR U7147 ( .A(\w0[3][103] ), .B(g_input[487]), .Z(n2521) );
  ANDN U7148 ( .A(\SUBBYTES[3].a/w897 ), .B(n2520), .Z(\SUBBYTES[3].a/w804 )
         );
  XNOR U7149 ( .A(\w1[3][100] ), .B(\w1[3][98] ), .Z(n2520) );
  XOR U7150 ( .A(\w0[3][98] ), .B(g_input[482]), .Z(\w1[3][98] ) );
  XOR U7151 ( .A(\w0[3][100] ), .B(g_input[484]), .Z(\w1[3][100] ) );
  AND U7152 ( .A(n2522), .B(\SUBBYTES[3].a/w574 ), .Z(\SUBBYTES[3].a/w709 ) );
  AND U7153 ( .A(n2523), .B(\SUBBYTES[3].a/w575 ), .Z(\SUBBYTES[3].a/w707 ) );
  AND U7154 ( .A(\SUBBYTES[3].a/w705 ), .B(n2524), .Z(\SUBBYTES[3].a/w706 ) );
  ANDN U7155 ( .A(\w1[3][104] ), .B(n2525), .Z(\SUBBYTES[3].a/w702 ) );
  AND U7156 ( .A(n2526), .B(\SUBBYTES[3].a/w577 ), .Z(\SUBBYTES[3].a/w700 ) );
  AND U7157 ( .A(\SUBBYTES[3].a/w698 ), .B(n2527), .Z(\SUBBYTES[3].a/w699 ) );
  XOR U7158 ( .A(\SUBBYTES[3].a/w642 ), .B(n8396), .Z(n2527) );
  AND U7159 ( .A(\SUBBYTES[3].a/w685 ), .B(\SUBBYTES[3].a/w687 ), .Z(
        \SUBBYTES[3].a/w694 ) );
  AND U7160 ( .A(\SUBBYTES[3].a/w686 ), .B(\SUBBYTES[3].a/w688 ), .Z(
        \SUBBYTES[3].a/w692 ) );
  AND U7161 ( .A(\SUBBYTES[3].a/w689 ), .B(\SUBBYTES[3].a/w690 ), .Z(
        \SUBBYTES[3].a/w691 ) );
  AND U7162 ( .A(\SUBBYTES[3].a/w578 ), .B(n2522), .Z(\SUBBYTES[3].a/w677 ) );
  XOR U7163 ( .A(\SUBBYTES[3].a/w646 ), .B(n991), .Z(n2522) );
  AND U7164 ( .A(\SUBBYTES[3].a/w579 ), .B(n2523), .Z(\SUBBYTES[3].a/w675 ) );
  XOR U7165 ( .A(n8397), .B(\SUBBYTES[3].a/w646 ), .Z(n2523) );
  ANDN U7166 ( .A(n2524), .B(n2528), .Z(\SUBBYTES[3].a/w674 ) );
  XOR U7167 ( .A(n991), .B(n8397), .Z(n2524) );
  ANDN U7168 ( .A(\SUBBYTES[3].a/w580 ), .B(n2525), .Z(\SUBBYTES[3].a/w670 )
         );
  XNOR U7169 ( .A(\SUBBYTES[3].a/w639 ), .B(\SUBBYTES[3].a/w642 ), .Z(n2525)
         );
  AND U7170 ( .A(\SUBBYTES[3].a/w581 ), .B(n2526), .Z(\SUBBYTES[3].a/w668 ) );
  XNOR U7171 ( .A(n2529), .B(\SUBBYTES[3].a/w639 ), .Z(n2526) );
  AND U7172 ( .A(\SUBBYTES[3].a/w666 ), .B(n2530), .Z(\SUBBYTES[3].a/w667 ) );
  XOR U7173 ( .A(n2531), .B(n2529), .Z(n2530) );
  IV U7174 ( .A(n8396), .Z(n2529) );
  ANDN U7175 ( .A(\SUBBYTES[3].a/w685 ), .B(n2532), .Z(\SUBBYTES[3].a/w662 )
         );
  ANDN U7176 ( .A(\SUBBYTES[3].a/w686 ), .B(n2533), .Z(\SUBBYTES[3].a/w660 )
         );
  ANDN U7177 ( .A(\SUBBYTES[3].a/w689 ), .B(n2534), .Z(\SUBBYTES[3].a/w659 )
         );
  AND U7178 ( .A(\SUBBYTES[3].a/w645 ), .B(\SUBBYTES[3].a/w644 ), .Z(
        \SUBBYTES[3].a/w646 ) );
  IV U7179 ( .A(n2531), .Z(\SUBBYTES[3].a/w642 ) );
  NAND U7180 ( .A(\SUBBYTES[3].a/w621 ), .B(\SUBBYTES[3].a/w636 ), .Z(n2531)
         );
  AND U7181 ( .A(\SUBBYTES[3].a/w638 ), .B(\SUBBYTES[3].a/w644 ), .Z(
        \SUBBYTES[3].a/w639 ) );
  AND U7182 ( .A(\SUBBYTES[3].a/w623 ), .B(\SUBBYTES[3].a/w621 ), .Z(
        \SUBBYTES[3].a/w633 ) );
  AND U7183 ( .A(\SUBBYTES[3].a/w624 ), .B(\SUBBYTES[3].a/w622 ), .Z(
        \SUBBYTES[3].a/w631 ) );
  AND U7184 ( .A(\SUBBYTES[3].a/w638 ), .B(\SUBBYTES[3].a/w645 ), .Z(
        \SUBBYTES[3].a/w630 ) );
  AND U7185 ( .A(\SUBBYTES[3].a/w578 ), .B(\SUBBYTES[3].a/w574 ), .Z(
        \SUBBYTES[3].a/w615 ) );
  AND U7186 ( .A(\SUBBYTES[3].a/w579 ), .B(\SUBBYTES[3].a/w575 ), .Z(
        \SUBBYTES[3].a/w613 ) );
  ANDN U7187 ( .A(\SUBBYTES[3].a/w705 ), .B(n2528), .Z(\SUBBYTES[3].a/w612 )
         );
  XNOR U7188 ( .A(\w1[3][105] ), .B(\w1[3][111] ), .Z(n2528) );
  XOR U7189 ( .A(\w0[3][105] ), .B(g_input[489]), .Z(\w1[3][105] ) );
  AND U7190 ( .A(\w1[3][104] ), .B(\SUBBYTES[3].a/w580 ), .Z(
        \SUBBYTES[3].a/w608 ) );
  XOR U7191 ( .A(\w0[3][104] ), .B(g_input[488]), .Z(\w1[3][104] ) );
  AND U7192 ( .A(\SUBBYTES[3].a/w581 ), .B(\SUBBYTES[3].a/w577 ), .Z(
        \SUBBYTES[3].a/w606 ) );
  AND U7193 ( .A(\SUBBYTES[3].a/w666 ), .B(\SUBBYTES[3].a/w698 ), .Z(
        \SUBBYTES[3].a/w605 ) );
  ANDN U7194 ( .A(\SUBBYTES[3].a/w687 ), .B(n2532), .Z(\SUBBYTES[3].a/w600 )
         );
  XNOR U7195 ( .A(\w1[3][108] ), .B(\w1[3][111] ), .Z(n2532) );
  ANDN U7196 ( .A(\SUBBYTES[3].a/w688 ), .B(n2533), .Z(\SUBBYTES[3].a/w598 )
         );
  XNOR U7197 ( .A(\w1[3][106] ), .B(\w1[3][111] ), .Z(n2533) );
  XOR U7198 ( .A(\w0[3][111] ), .B(g_input[495]), .Z(\w1[3][111] ) );
  IV U7199 ( .A(n2535), .Z(\w1[3][106] ) );
  ANDN U7200 ( .A(\SUBBYTES[3].a/w690 ), .B(n2534), .Z(\SUBBYTES[3].a/w597 )
         );
  XOR U7201 ( .A(n2535), .B(\w1[3][108] ), .Z(n2534) );
  XOR U7202 ( .A(\w0[3][108] ), .B(g_input[492]), .Z(\w1[3][108] ) );
  XNOR U7203 ( .A(\w0[3][106] ), .B(g_input[490]), .Z(n2535) );
  AND U7204 ( .A(n2536), .B(\SUBBYTES[3].a/w367 ), .Z(\SUBBYTES[3].a/w502 ) );
  AND U7205 ( .A(n2537), .B(\SUBBYTES[3].a/w368 ), .Z(\SUBBYTES[3].a/w500 ) );
  AND U7206 ( .A(\SUBBYTES[3].a/w498 ), .B(n2538), .Z(\SUBBYTES[3].a/w499 ) );
  ANDN U7207 ( .A(\w1[3][112] ), .B(n2539), .Z(\SUBBYTES[3].a/w495 ) );
  AND U7208 ( .A(n2540), .B(\SUBBYTES[3].a/w370 ), .Z(\SUBBYTES[3].a/w493 ) );
  AND U7209 ( .A(\SUBBYTES[3].a/w491 ), .B(n2541), .Z(\SUBBYTES[3].a/w492 ) );
  XOR U7210 ( .A(\SUBBYTES[3].a/w435 ), .B(n8394), .Z(n2541) );
  AND U7211 ( .A(\SUBBYTES[3].a/w478 ), .B(\SUBBYTES[3].a/w480 ), .Z(
        \SUBBYTES[3].a/w487 ) );
  AND U7212 ( .A(\SUBBYTES[3].a/w479 ), .B(\SUBBYTES[3].a/w481 ), .Z(
        \SUBBYTES[3].a/w485 ) );
  AND U7213 ( .A(\SUBBYTES[3].a/w482 ), .B(\SUBBYTES[3].a/w483 ), .Z(
        \SUBBYTES[3].a/w484 ) );
  AND U7214 ( .A(\SUBBYTES[3].a/w371 ), .B(n2536), .Z(\SUBBYTES[3].a/w470 ) );
  XOR U7215 ( .A(\SUBBYTES[3].a/w439 ), .B(n990), .Z(n2536) );
  AND U7216 ( .A(\SUBBYTES[3].a/w372 ), .B(n2537), .Z(\SUBBYTES[3].a/w468 ) );
  XOR U7217 ( .A(n8395), .B(\SUBBYTES[3].a/w439 ), .Z(n2537) );
  ANDN U7218 ( .A(n2538), .B(n2542), .Z(\SUBBYTES[3].a/w467 ) );
  XOR U7219 ( .A(n990), .B(n8395), .Z(n2538) );
  ANDN U7220 ( .A(\SUBBYTES[3].a/w373 ), .B(n2539), .Z(\SUBBYTES[3].a/w463 )
         );
  XNOR U7221 ( .A(\SUBBYTES[3].a/w432 ), .B(\SUBBYTES[3].a/w435 ), .Z(n2539)
         );
  AND U7222 ( .A(\SUBBYTES[3].a/w374 ), .B(n2540), .Z(\SUBBYTES[3].a/w461 ) );
  XNOR U7223 ( .A(n2543), .B(\SUBBYTES[3].a/w432 ), .Z(n2540) );
  AND U7224 ( .A(\SUBBYTES[3].a/w459 ), .B(n2544), .Z(\SUBBYTES[3].a/w460 ) );
  XOR U7225 ( .A(n2545), .B(n2543), .Z(n2544) );
  IV U7226 ( .A(n8394), .Z(n2543) );
  ANDN U7227 ( .A(\SUBBYTES[3].a/w478 ), .B(n2546), .Z(\SUBBYTES[3].a/w455 )
         );
  ANDN U7228 ( .A(\SUBBYTES[3].a/w479 ), .B(n2547), .Z(\SUBBYTES[3].a/w453 )
         );
  ANDN U7229 ( .A(\SUBBYTES[3].a/w482 ), .B(n2548), .Z(\SUBBYTES[3].a/w452 )
         );
  AND U7230 ( .A(\SUBBYTES[3].a/w438 ), .B(\SUBBYTES[3].a/w437 ), .Z(
        \SUBBYTES[3].a/w439 ) );
  IV U7231 ( .A(n2545), .Z(\SUBBYTES[3].a/w435 ) );
  NAND U7232 ( .A(\SUBBYTES[3].a/w414 ), .B(\SUBBYTES[3].a/w429 ), .Z(n2545)
         );
  AND U7233 ( .A(\SUBBYTES[3].a/w431 ), .B(\SUBBYTES[3].a/w437 ), .Z(
        \SUBBYTES[3].a/w432 ) );
  AND U7234 ( .A(\SUBBYTES[3].a/w416 ), .B(\SUBBYTES[3].a/w414 ), .Z(
        \SUBBYTES[3].a/w426 ) );
  AND U7235 ( .A(\SUBBYTES[3].a/w417 ), .B(\SUBBYTES[3].a/w415 ), .Z(
        \SUBBYTES[3].a/w424 ) );
  AND U7236 ( .A(\SUBBYTES[3].a/w431 ), .B(\SUBBYTES[3].a/w438 ), .Z(
        \SUBBYTES[3].a/w423 ) );
  AND U7237 ( .A(\SUBBYTES[3].a/w371 ), .B(\SUBBYTES[3].a/w367 ), .Z(
        \SUBBYTES[3].a/w408 ) );
  AND U7238 ( .A(\SUBBYTES[3].a/w372 ), .B(\SUBBYTES[3].a/w368 ), .Z(
        \SUBBYTES[3].a/w406 ) );
  ANDN U7239 ( .A(\SUBBYTES[3].a/w498 ), .B(n2542), .Z(\SUBBYTES[3].a/w405 )
         );
  XNOR U7240 ( .A(\w1[3][113] ), .B(\w1[3][119] ), .Z(n2542) );
  XOR U7241 ( .A(\w0[3][113] ), .B(g_input[497]), .Z(\w1[3][113] ) );
  AND U7242 ( .A(\w1[3][112] ), .B(\SUBBYTES[3].a/w373 ), .Z(
        \SUBBYTES[3].a/w401 ) );
  XOR U7243 ( .A(\w0[3][112] ), .B(g_input[496]), .Z(\w1[3][112] ) );
  AND U7244 ( .A(\SUBBYTES[3].a/w374 ), .B(\SUBBYTES[3].a/w370 ), .Z(
        \SUBBYTES[3].a/w399 ) );
  AND U7245 ( .A(\SUBBYTES[3].a/w459 ), .B(\SUBBYTES[3].a/w491 ), .Z(
        \SUBBYTES[3].a/w398 ) );
  ANDN U7246 ( .A(\SUBBYTES[3].a/w480 ), .B(n2546), .Z(\SUBBYTES[3].a/w393 )
         );
  XNOR U7247 ( .A(\w1[3][116] ), .B(\w1[3][119] ), .Z(n2546) );
  ANDN U7248 ( .A(\SUBBYTES[3].a/w481 ), .B(n2547), .Z(\SUBBYTES[3].a/w391 )
         );
  XNOR U7249 ( .A(\w1[3][114] ), .B(\w1[3][119] ), .Z(n2547) );
  XOR U7250 ( .A(\w0[3][119] ), .B(g_input[503]), .Z(\w1[3][119] ) );
  IV U7251 ( .A(n2549), .Z(\w1[3][114] ) );
  ANDN U7252 ( .A(\SUBBYTES[3].a/w483 ), .B(n2548), .Z(\SUBBYTES[3].a/w390 )
         );
  XOR U7253 ( .A(n2549), .B(\w1[3][116] ), .Z(n2548) );
  XOR U7254 ( .A(\w0[3][116] ), .B(g_input[500]), .Z(\w1[3][116] ) );
  XNOR U7255 ( .A(\w0[3][114] ), .B(g_input[498]), .Z(n2549) );
  AND U7256 ( .A(n2550), .B(\SUBBYTES[3].a/w3265 ), .Z(\SUBBYTES[3].a/w3400 )
         );
  AND U7257 ( .A(n2551), .B(\SUBBYTES[3].a/w3266 ), .Z(\SUBBYTES[3].a/w3398 )
         );
  AND U7258 ( .A(\SUBBYTES[3].a/w3396 ), .B(n2552), .Z(\SUBBYTES[3].a/w3397 )
         );
  ANDN U7259 ( .A(\w1[3][0] ), .B(n2553), .Z(\SUBBYTES[3].a/w3393 ) );
  AND U7260 ( .A(n2554), .B(\SUBBYTES[3].a/w3268 ), .Z(\SUBBYTES[3].a/w3391 )
         );
  AND U7261 ( .A(\SUBBYTES[3].a/w3389 ), .B(n2555), .Z(\SUBBYTES[3].a/w3390 )
         );
  XOR U7262 ( .A(\SUBBYTES[3].a/w3333 ), .B(n8422), .Z(n2555) );
  AND U7263 ( .A(\SUBBYTES[3].a/w3376 ), .B(\SUBBYTES[3].a/w3378 ), .Z(
        \SUBBYTES[3].a/w3385 ) );
  AND U7264 ( .A(\SUBBYTES[3].a/w3377 ), .B(\SUBBYTES[3].a/w3379 ), .Z(
        \SUBBYTES[3].a/w3383 ) );
  AND U7265 ( .A(\SUBBYTES[3].a/w3380 ), .B(\SUBBYTES[3].a/w3381 ), .Z(
        \SUBBYTES[3].a/w3382 ) );
  AND U7266 ( .A(\SUBBYTES[3].a/w3269 ), .B(n2550), .Z(\SUBBYTES[3].a/w3368 )
         );
  XOR U7267 ( .A(\SUBBYTES[3].a/w3337 ), .B(n1004), .Z(n2550) );
  AND U7268 ( .A(\SUBBYTES[3].a/w3270 ), .B(n2551), .Z(\SUBBYTES[3].a/w3366 )
         );
  XOR U7269 ( .A(n8423), .B(\SUBBYTES[3].a/w3337 ), .Z(n2551) );
  ANDN U7270 ( .A(n2552), .B(n2556), .Z(\SUBBYTES[3].a/w3365 ) );
  XOR U7271 ( .A(n1004), .B(n8423), .Z(n2552) );
  ANDN U7272 ( .A(\SUBBYTES[3].a/w3271 ), .B(n2553), .Z(\SUBBYTES[3].a/w3361 )
         );
  XNOR U7273 ( .A(\SUBBYTES[3].a/w3330 ), .B(\SUBBYTES[3].a/w3333 ), .Z(n2553)
         );
  AND U7274 ( .A(\SUBBYTES[3].a/w3272 ), .B(n2554), .Z(\SUBBYTES[3].a/w3359 )
         );
  XNOR U7275 ( .A(n2557), .B(\SUBBYTES[3].a/w3330 ), .Z(n2554) );
  AND U7276 ( .A(\SUBBYTES[3].a/w3357 ), .B(n2558), .Z(\SUBBYTES[3].a/w3358 )
         );
  XOR U7277 ( .A(n2559), .B(n2557), .Z(n2558) );
  IV U7278 ( .A(n8422), .Z(n2557) );
  ANDN U7279 ( .A(\SUBBYTES[3].a/w3376 ), .B(n2560), .Z(\SUBBYTES[3].a/w3353 )
         );
  ANDN U7280 ( .A(\SUBBYTES[3].a/w3377 ), .B(n2561), .Z(\SUBBYTES[3].a/w3351 )
         );
  ANDN U7281 ( .A(\SUBBYTES[3].a/w3380 ), .B(n2562), .Z(\SUBBYTES[3].a/w3350 )
         );
  AND U7282 ( .A(\SUBBYTES[3].a/w3336 ), .B(\SUBBYTES[3].a/w3335 ), .Z(
        \SUBBYTES[3].a/w3337 ) );
  IV U7283 ( .A(n2559), .Z(\SUBBYTES[3].a/w3333 ) );
  NAND U7284 ( .A(\SUBBYTES[3].a/w3312 ), .B(\SUBBYTES[3].a/w3327 ), .Z(n2559)
         );
  AND U7285 ( .A(\SUBBYTES[3].a/w3329 ), .B(\SUBBYTES[3].a/w3335 ), .Z(
        \SUBBYTES[3].a/w3330 ) );
  AND U7286 ( .A(\SUBBYTES[3].a/w3314 ), .B(\SUBBYTES[3].a/w3312 ), .Z(
        \SUBBYTES[3].a/w3324 ) );
  AND U7287 ( .A(\SUBBYTES[3].a/w3315 ), .B(\SUBBYTES[3].a/w3313 ), .Z(
        \SUBBYTES[3].a/w3322 ) );
  AND U7288 ( .A(\SUBBYTES[3].a/w3329 ), .B(\SUBBYTES[3].a/w3336 ), .Z(
        \SUBBYTES[3].a/w3321 ) );
  AND U7289 ( .A(\SUBBYTES[3].a/w3269 ), .B(\SUBBYTES[3].a/w3265 ), .Z(
        \SUBBYTES[3].a/w3306 ) );
  AND U7290 ( .A(\SUBBYTES[3].a/w3270 ), .B(\SUBBYTES[3].a/w3266 ), .Z(
        \SUBBYTES[3].a/w3304 ) );
  ANDN U7291 ( .A(\SUBBYTES[3].a/w3396 ), .B(n2556), .Z(\SUBBYTES[3].a/w3303 )
         );
  XNOR U7292 ( .A(\w1[3][1] ), .B(\w1[3][7] ), .Z(n2556) );
  XOR U7293 ( .A(\w0[3][1] ), .B(g_input[385]), .Z(\w1[3][1] ) );
  AND U7294 ( .A(\w1[3][0] ), .B(\SUBBYTES[3].a/w3271 ), .Z(
        \SUBBYTES[3].a/w3299 ) );
  XOR U7295 ( .A(\w0[3][0] ), .B(g_input[384]), .Z(\w1[3][0] ) );
  AND U7296 ( .A(\SUBBYTES[3].a/w3272 ), .B(\SUBBYTES[3].a/w3268 ), .Z(
        \SUBBYTES[3].a/w3297 ) );
  AND U7297 ( .A(\SUBBYTES[3].a/w3357 ), .B(\SUBBYTES[3].a/w3389 ), .Z(
        \SUBBYTES[3].a/w3296 ) );
  ANDN U7298 ( .A(\SUBBYTES[3].a/w3378 ), .B(n2560), .Z(\SUBBYTES[3].a/w3291 )
         );
  XNOR U7299 ( .A(\w1[3][4] ), .B(\w1[3][7] ), .Z(n2560) );
  ANDN U7300 ( .A(\SUBBYTES[3].a/w3379 ), .B(n2561), .Z(\SUBBYTES[3].a/w3289 )
         );
  XNOR U7301 ( .A(\w1[3][2] ), .B(\w1[3][7] ), .Z(n2561) );
  XOR U7302 ( .A(\w0[3][7] ), .B(g_input[391]), .Z(\w1[3][7] ) );
  IV U7303 ( .A(n2563), .Z(\w1[3][2] ) );
  ANDN U7304 ( .A(\SUBBYTES[3].a/w3381 ), .B(n2562), .Z(\SUBBYTES[3].a/w3288 )
         );
  XOR U7305 ( .A(n2563), .B(\w1[3][4] ), .Z(n2562) );
  XOR U7306 ( .A(\w0[3][4] ), .B(g_input[388]), .Z(\w1[3][4] ) );
  XNOR U7307 ( .A(\w0[3][2] ), .B(g_input[386]), .Z(n2563) );
  AND U7308 ( .A(n2564), .B(\SUBBYTES[3].a/w3058 ), .Z(\SUBBYTES[3].a/w3193 )
         );
  AND U7309 ( .A(n2565), .B(\SUBBYTES[3].a/w3059 ), .Z(\SUBBYTES[3].a/w3191 )
         );
  AND U7310 ( .A(\SUBBYTES[3].a/w3189 ), .B(n2566), .Z(\SUBBYTES[3].a/w3190 )
         );
  ANDN U7311 ( .A(\w1[3][8] ), .B(n2567), .Z(\SUBBYTES[3].a/w3186 ) );
  AND U7312 ( .A(n2568), .B(\SUBBYTES[3].a/w3061 ), .Z(\SUBBYTES[3].a/w3184 )
         );
  AND U7313 ( .A(\SUBBYTES[3].a/w3182 ), .B(n2569), .Z(\SUBBYTES[3].a/w3183 )
         );
  XOR U7314 ( .A(\SUBBYTES[3].a/w3126 ), .B(n8420), .Z(n2569) );
  AND U7315 ( .A(\SUBBYTES[3].a/w3169 ), .B(\SUBBYTES[3].a/w3171 ), .Z(
        \SUBBYTES[3].a/w3178 ) );
  AND U7316 ( .A(\SUBBYTES[3].a/w3170 ), .B(\SUBBYTES[3].a/w3172 ), .Z(
        \SUBBYTES[3].a/w3176 ) );
  AND U7317 ( .A(\SUBBYTES[3].a/w3173 ), .B(\SUBBYTES[3].a/w3174 ), .Z(
        \SUBBYTES[3].a/w3175 ) );
  AND U7318 ( .A(\SUBBYTES[3].a/w3062 ), .B(n2564), .Z(\SUBBYTES[3].a/w3161 )
         );
  XOR U7319 ( .A(\SUBBYTES[3].a/w3130 ), .B(n1003), .Z(n2564) );
  AND U7320 ( .A(\SUBBYTES[3].a/w3063 ), .B(n2565), .Z(\SUBBYTES[3].a/w3159 )
         );
  XOR U7321 ( .A(n8421), .B(\SUBBYTES[3].a/w3130 ), .Z(n2565) );
  ANDN U7322 ( .A(n2566), .B(n2570), .Z(\SUBBYTES[3].a/w3158 ) );
  XOR U7323 ( .A(n1003), .B(n8421), .Z(n2566) );
  ANDN U7324 ( .A(\SUBBYTES[3].a/w3064 ), .B(n2567), .Z(\SUBBYTES[3].a/w3154 )
         );
  XNOR U7325 ( .A(\SUBBYTES[3].a/w3123 ), .B(\SUBBYTES[3].a/w3126 ), .Z(n2567)
         );
  AND U7326 ( .A(\SUBBYTES[3].a/w3065 ), .B(n2568), .Z(\SUBBYTES[3].a/w3152 )
         );
  XNOR U7327 ( .A(n2571), .B(\SUBBYTES[3].a/w3123 ), .Z(n2568) );
  AND U7328 ( .A(\SUBBYTES[3].a/w3150 ), .B(n2572), .Z(\SUBBYTES[3].a/w3151 )
         );
  XOR U7329 ( .A(n2573), .B(n2571), .Z(n2572) );
  IV U7330 ( .A(n8420), .Z(n2571) );
  ANDN U7331 ( .A(\SUBBYTES[3].a/w3169 ), .B(n2574), .Z(\SUBBYTES[3].a/w3146 )
         );
  ANDN U7332 ( .A(\SUBBYTES[3].a/w3170 ), .B(n2575), .Z(\SUBBYTES[3].a/w3144 )
         );
  ANDN U7333 ( .A(\SUBBYTES[3].a/w3173 ), .B(n2576), .Z(\SUBBYTES[3].a/w3143 )
         );
  AND U7334 ( .A(\SUBBYTES[3].a/w3129 ), .B(\SUBBYTES[3].a/w3128 ), .Z(
        \SUBBYTES[3].a/w3130 ) );
  IV U7335 ( .A(n2573), .Z(\SUBBYTES[3].a/w3126 ) );
  NAND U7336 ( .A(\SUBBYTES[3].a/w3105 ), .B(\SUBBYTES[3].a/w3120 ), .Z(n2573)
         );
  AND U7337 ( .A(\SUBBYTES[3].a/w3122 ), .B(\SUBBYTES[3].a/w3128 ), .Z(
        \SUBBYTES[3].a/w3123 ) );
  AND U7338 ( .A(\SUBBYTES[3].a/w3107 ), .B(\SUBBYTES[3].a/w3105 ), .Z(
        \SUBBYTES[3].a/w3117 ) );
  AND U7339 ( .A(\SUBBYTES[3].a/w3108 ), .B(\SUBBYTES[3].a/w3106 ), .Z(
        \SUBBYTES[3].a/w3115 ) );
  AND U7340 ( .A(\SUBBYTES[3].a/w3122 ), .B(\SUBBYTES[3].a/w3129 ), .Z(
        \SUBBYTES[3].a/w3114 ) );
  AND U7341 ( .A(\SUBBYTES[3].a/w3062 ), .B(\SUBBYTES[3].a/w3058 ), .Z(
        \SUBBYTES[3].a/w3099 ) );
  AND U7342 ( .A(\SUBBYTES[3].a/w3063 ), .B(\SUBBYTES[3].a/w3059 ), .Z(
        \SUBBYTES[3].a/w3097 ) );
  ANDN U7343 ( .A(\SUBBYTES[3].a/w3189 ), .B(n2570), .Z(\SUBBYTES[3].a/w3096 )
         );
  XNOR U7344 ( .A(\w1[3][15] ), .B(\w1[3][9] ), .Z(n2570) );
  XOR U7345 ( .A(\w0[3][9] ), .B(g_input[393]), .Z(\w1[3][9] ) );
  AND U7346 ( .A(\w1[3][8] ), .B(\SUBBYTES[3].a/w3064 ), .Z(
        \SUBBYTES[3].a/w3092 ) );
  XOR U7347 ( .A(\w0[3][8] ), .B(g_input[392]), .Z(\w1[3][8] ) );
  AND U7348 ( .A(\SUBBYTES[3].a/w3065 ), .B(\SUBBYTES[3].a/w3061 ), .Z(
        \SUBBYTES[3].a/w3090 ) );
  AND U7349 ( .A(\SUBBYTES[3].a/w3150 ), .B(\SUBBYTES[3].a/w3182 ), .Z(
        \SUBBYTES[3].a/w3089 ) );
  ANDN U7350 ( .A(\SUBBYTES[3].a/w3171 ), .B(n2574), .Z(\SUBBYTES[3].a/w3084 )
         );
  XNOR U7351 ( .A(\w1[3][12] ), .B(\w1[3][15] ), .Z(n2574) );
  ANDN U7352 ( .A(\SUBBYTES[3].a/w3172 ), .B(n2575), .Z(\SUBBYTES[3].a/w3082 )
         );
  XNOR U7353 ( .A(\w1[3][10] ), .B(\w1[3][15] ), .Z(n2575) );
  XOR U7354 ( .A(\w0[3][15] ), .B(g_input[399]), .Z(\w1[3][15] ) );
  ANDN U7355 ( .A(\SUBBYTES[3].a/w3174 ), .B(n2576), .Z(\SUBBYTES[3].a/w3081 )
         );
  XNOR U7356 ( .A(\w1[3][10] ), .B(\w1[3][12] ), .Z(n2576) );
  XOR U7357 ( .A(\w0[3][12] ), .B(g_input[396]), .Z(\w1[3][12] ) );
  XOR U7358 ( .A(\w0[3][10] ), .B(g_input[394]), .Z(\w1[3][10] ) );
  AND U7359 ( .A(n2577), .B(\SUBBYTES[3].a/w2851 ), .Z(\SUBBYTES[3].a/w2986 )
         );
  AND U7360 ( .A(n2578), .B(\SUBBYTES[3].a/w2852 ), .Z(\SUBBYTES[3].a/w2984 )
         );
  AND U7361 ( .A(\SUBBYTES[3].a/w2982 ), .B(n2579), .Z(\SUBBYTES[3].a/w2983 )
         );
  ANDN U7362 ( .A(\w1[3][16] ), .B(n2580), .Z(\SUBBYTES[3].a/w2979 ) );
  AND U7363 ( .A(n2581), .B(\SUBBYTES[3].a/w2854 ), .Z(\SUBBYTES[3].a/w2977 )
         );
  AND U7364 ( .A(\SUBBYTES[3].a/w2975 ), .B(n2582), .Z(\SUBBYTES[3].a/w2976 )
         );
  XOR U7365 ( .A(\SUBBYTES[3].a/w2919 ), .B(n8418), .Z(n2582) );
  AND U7366 ( .A(\SUBBYTES[3].a/w2962 ), .B(\SUBBYTES[3].a/w2964 ), .Z(
        \SUBBYTES[3].a/w2971 ) );
  AND U7367 ( .A(\SUBBYTES[3].a/w2963 ), .B(\SUBBYTES[3].a/w2965 ), .Z(
        \SUBBYTES[3].a/w2969 ) );
  AND U7368 ( .A(\SUBBYTES[3].a/w2966 ), .B(\SUBBYTES[3].a/w2967 ), .Z(
        \SUBBYTES[3].a/w2968 ) );
  AND U7369 ( .A(\SUBBYTES[3].a/w2855 ), .B(n2577), .Z(\SUBBYTES[3].a/w2954 )
         );
  XOR U7370 ( .A(\SUBBYTES[3].a/w2923 ), .B(n1002), .Z(n2577) );
  AND U7371 ( .A(\SUBBYTES[3].a/w2856 ), .B(n2578), .Z(\SUBBYTES[3].a/w2952 )
         );
  XOR U7372 ( .A(n8419), .B(\SUBBYTES[3].a/w2923 ), .Z(n2578) );
  ANDN U7373 ( .A(n2579), .B(n2583), .Z(\SUBBYTES[3].a/w2951 ) );
  XOR U7374 ( .A(n1002), .B(n8419), .Z(n2579) );
  AND U7375 ( .A(n2584), .B(\SUBBYTES[3].a/w160 ), .Z(\SUBBYTES[3].a/w295 ) );
  ANDN U7376 ( .A(\SUBBYTES[3].a/w2857 ), .B(n2580), .Z(\SUBBYTES[3].a/w2947 )
         );
  XNOR U7377 ( .A(\SUBBYTES[3].a/w2916 ), .B(\SUBBYTES[3].a/w2919 ), .Z(n2580)
         );
  AND U7378 ( .A(\SUBBYTES[3].a/w2858 ), .B(n2581), .Z(\SUBBYTES[3].a/w2945 )
         );
  XNOR U7379 ( .A(n2585), .B(\SUBBYTES[3].a/w2916 ), .Z(n2581) );
  AND U7380 ( .A(\SUBBYTES[3].a/w2943 ), .B(n2586), .Z(\SUBBYTES[3].a/w2944 )
         );
  XOR U7381 ( .A(n2587), .B(n2585), .Z(n2586) );
  IV U7382 ( .A(n8418), .Z(n2585) );
  ANDN U7383 ( .A(\SUBBYTES[3].a/w2962 ), .B(n2588), .Z(\SUBBYTES[3].a/w2939 )
         );
  ANDN U7384 ( .A(\SUBBYTES[3].a/w2963 ), .B(n2589), .Z(\SUBBYTES[3].a/w2937 )
         );
  ANDN U7385 ( .A(\SUBBYTES[3].a/w2966 ), .B(n2590), .Z(\SUBBYTES[3].a/w2936 )
         );
  AND U7386 ( .A(n2591), .B(\SUBBYTES[3].a/w161 ), .Z(\SUBBYTES[3].a/w293 ) );
  AND U7387 ( .A(\SUBBYTES[3].a/w2922 ), .B(\SUBBYTES[3].a/w2921 ), .Z(
        \SUBBYTES[3].a/w2923 ) );
  AND U7388 ( .A(\SUBBYTES[3].a/w291 ), .B(n2592), .Z(\SUBBYTES[3].a/w292 ) );
  IV U7389 ( .A(n2587), .Z(\SUBBYTES[3].a/w2919 ) );
  NAND U7390 ( .A(\SUBBYTES[3].a/w2898 ), .B(\SUBBYTES[3].a/w2913 ), .Z(n2587)
         );
  AND U7391 ( .A(\SUBBYTES[3].a/w2915 ), .B(\SUBBYTES[3].a/w2921 ), .Z(
        \SUBBYTES[3].a/w2916 ) );
  AND U7392 ( .A(\SUBBYTES[3].a/w2900 ), .B(\SUBBYTES[3].a/w2898 ), .Z(
        \SUBBYTES[3].a/w2910 ) );
  AND U7393 ( .A(\SUBBYTES[3].a/w2901 ), .B(\SUBBYTES[3].a/w2899 ), .Z(
        \SUBBYTES[3].a/w2908 ) );
  AND U7394 ( .A(\SUBBYTES[3].a/w2915 ), .B(\SUBBYTES[3].a/w2922 ), .Z(
        \SUBBYTES[3].a/w2907 ) );
  AND U7395 ( .A(\SUBBYTES[3].a/w2855 ), .B(\SUBBYTES[3].a/w2851 ), .Z(
        \SUBBYTES[3].a/w2892 ) );
  AND U7396 ( .A(\SUBBYTES[3].a/w2856 ), .B(\SUBBYTES[3].a/w2852 ), .Z(
        \SUBBYTES[3].a/w2890 ) );
  ANDN U7397 ( .A(\SUBBYTES[3].a/w2982 ), .B(n2583), .Z(\SUBBYTES[3].a/w2889 )
         );
  XNOR U7398 ( .A(\w1[3][17] ), .B(\w1[3][23] ), .Z(n2583) );
  XOR U7399 ( .A(\w0[3][17] ), .B(g_input[401]), .Z(\w1[3][17] ) );
  AND U7400 ( .A(\w1[3][16] ), .B(\SUBBYTES[3].a/w2857 ), .Z(
        \SUBBYTES[3].a/w2885 ) );
  XOR U7401 ( .A(\w0[3][16] ), .B(g_input[400]), .Z(\w1[3][16] ) );
  AND U7402 ( .A(\SUBBYTES[3].a/w2858 ), .B(\SUBBYTES[3].a/w2854 ), .Z(
        \SUBBYTES[3].a/w2883 ) );
  AND U7403 ( .A(\SUBBYTES[3].a/w2943 ), .B(\SUBBYTES[3].a/w2975 ), .Z(
        \SUBBYTES[3].a/w2882 ) );
  ANDN U7404 ( .A(\w1[3][120] ), .B(n2593), .Z(\SUBBYTES[3].a/w288 ) );
  ANDN U7405 ( .A(\SUBBYTES[3].a/w2964 ), .B(n2588), .Z(\SUBBYTES[3].a/w2877 )
         );
  XNOR U7406 ( .A(\w1[3][20] ), .B(\w1[3][23] ), .Z(n2588) );
  ANDN U7407 ( .A(\SUBBYTES[3].a/w2965 ), .B(n2589), .Z(\SUBBYTES[3].a/w2875 )
         );
  XNOR U7408 ( .A(\w1[3][18] ), .B(\w1[3][23] ), .Z(n2589) );
  XOR U7409 ( .A(\w0[3][23] ), .B(g_input[407]), .Z(\w1[3][23] ) );
  IV U7410 ( .A(n2594), .Z(\w1[3][18] ) );
  ANDN U7411 ( .A(\SUBBYTES[3].a/w2967 ), .B(n2590), .Z(\SUBBYTES[3].a/w2874 )
         );
  XOR U7412 ( .A(n2594), .B(\w1[3][20] ), .Z(n2590) );
  XOR U7413 ( .A(\w0[3][20] ), .B(g_input[404]), .Z(\w1[3][20] ) );
  XNOR U7414 ( .A(\w0[3][18] ), .B(g_input[402]), .Z(n2594) );
  AND U7415 ( .A(n2595), .B(\SUBBYTES[3].a/w163 ), .Z(\SUBBYTES[3].a/w286 ) );
  AND U7416 ( .A(\SUBBYTES[3].a/w284 ), .B(n2596), .Z(\SUBBYTES[3].a/w285 ) );
  XOR U7417 ( .A(\SUBBYTES[3].a/w228 ), .B(n8392), .Z(n2596) );
  AND U7418 ( .A(\SUBBYTES[3].a/w271 ), .B(\SUBBYTES[3].a/w273 ), .Z(
        \SUBBYTES[3].a/w280 ) );
  AND U7419 ( .A(\SUBBYTES[3].a/w272 ), .B(\SUBBYTES[3].a/w274 ), .Z(
        \SUBBYTES[3].a/w278 ) );
  AND U7420 ( .A(n2597), .B(\SUBBYTES[3].a/w2644 ), .Z(\SUBBYTES[3].a/w2779 )
         );
  AND U7421 ( .A(n2598), .B(\SUBBYTES[3].a/w2645 ), .Z(\SUBBYTES[3].a/w2777 )
         );
  AND U7422 ( .A(\SUBBYTES[3].a/w2775 ), .B(n2599), .Z(\SUBBYTES[3].a/w2776 )
         );
  ANDN U7423 ( .A(\w1[3][24] ), .B(n2600), .Z(\SUBBYTES[3].a/w2772 ) );
  AND U7424 ( .A(n2601), .B(\SUBBYTES[3].a/w2647 ), .Z(\SUBBYTES[3].a/w2770 )
         );
  AND U7425 ( .A(\SUBBYTES[3].a/w275 ), .B(\SUBBYTES[3].a/w276 ), .Z(
        \SUBBYTES[3].a/w277 ) );
  AND U7426 ( .A(\SUBBYTES[3].a/w2768 ), .B(n2602), .Z(\SUBBYTES[3].a/w2769 )
         );
  XOR U7427 ( .A(\SUBBYTES[3].a/w2712 ), .B(n8416), .Z(n2602) );
  AND U7428 ( .A(\SUBBYTES[3].a/w2755 ), .B(\SUBBYTES[3].a/w2757 ), .Z(
        \SUBBYTES[3].a/w2764 ) );
  AND U7429 ( .A(\SUBBYTES[3].a/w2756 ), .B(\SUBBYTES[3].a/w2758 ), .Z(
        \SUBBYTES[3].a/w2762 ) );
  AND U7430 ( .A(\SUBBYTES[3].a/w2759 ), .B(\SUBBYTES[3].a/w2760 ), .Z(
        \SUBBYTES[3].a/w2761 ) );
  AND U7431 ( .A(\SUBBYTES[3].a/w2648 ), .B(n2597), .Z(\SUBBYTES[3].a/w2747 )
         );
  XOR U7432 ( .A(\SUBBYTES[3].a/w2716 ), .B(n1001), .Z(n2597) );
  AND U7433 ( .A(\SUBBYTES[3].a/w2649 ), .B(n2598), .Z(\SUBBYTES[3].a/w2745 )
         );
  XOR U7434 ( .A(n8417), .B(\SUBBYTES[3].a/w2716 ), .Z(n2598) );
  ANDN U7435 ( .A(n2599), .B(n2603), .Z(\SUBBYTES[3].a/w2744 ) );
  XOR U7436 ( .A(n1001), .B(n8417), .Z(n2599) );
  ANDN U7437 ( .A(\SUBBYTES[3].a/w2650 ), .B(n2600), .Z(\SUBBYTES[3].a/w2740 )
         );
  XNOR U7438 ( .A(\SUBBYTES[3].a/w2709 ), .B(\SUBBYTES[3].a/w2712 ), .Z(n2600)
         );
  AND U7439 ( .A(\SUBBYTES[3].a/w2651 ), .B(n2601), .Z(\SUBBYTES[3].a/w2738 )
         );
  XNOR U7440 ( .A(n2604), .B(\SUBBYTES[3].a/w2709 ), .Z(n2601) );
  AND U7441 ( .A(\SUBBYTES[3].a/w2736 ), .B(n2605), .Z(\SUBBYTES[3].a/w2737 )
         );
  XOR U7442 ( .A(n2606), .B(n2604), .Z(n2605) );
  IV U7443 ( .A(n8416), .Z(n2604) );
  ANDN U7444 ( .A(\SUBBYTES[3].a/w2755 ), .B(n2607), .Z(\SUBBYTES[3].a/w2732 )
         );
  ANDN U7445 ( .A(\SUBBYTES[3].a/w2756 ), .B(n2608), .Z(\SUBBYTES[3].a/w2730 )
         );
  ANDN U7446 ( .A(\SUBBYTES[3].a/w2759 ), .B(n2609), .Z(\SUBBYTES[3].a/w2729 )
         );
  AND U7447 ( .A(\SUBBYTES[3].a/w2715 ), .B(\SUBBYTES[3].a/w2714 ), .Z(
        \SUBBYTES[3].a/w2716 ) );
  IV U7448 ( .A(n2606), .Z(\SUBBYTES[3].a/w2712 ) );
  NAND U7449 ( .A(\SUBBYTES[3].a/w2691 ), .B(\SUBBYTES[3].a/w2706 ), .Z(n2606)
         );
  AND U7450 ( .A(\SUBBYTES[3].a/w2708 ), .B(\SUBBYTES[3].a/w2714 ), .Z(
        \SUBBYTES[3].a/w2709 ) );
  AND U7451 ( .A(\SUBBYTES[3].a/w2693 ), .B(\SUBBYTES[3].a/w2691 ), .Z(
        \SUBBYTES[3].a/w2703 ) );
  AND U7452 ( .A(\SUBBYTES[3].a/w2694 ), .B(\SUBBYTES[3].a/w2692 ), .Z(
        \SUBBYTES[3].a/w2701 ) );
  AND U7453 ( .A(\SUBBYTES[3].a/w2708 ), .B(\SUBBYTES[3].a/w2715 ), .Z(
        \SUBBYTES[3].a/w2700 ) );
  AND U7454 ( .A(\SUBBYTES[3].a/w2648 ), .B(\SUBBYTES[3].a/w2644 ), .Z(
        \SUBBYTES[3].a/w2685 ) );
  AND U7455 ( .A(\SUBBYTES[3].a/w2649 ), .B(\SUBBYTES[3].a/w2645 ), .Z(
        \SUBBYTES[3].a/w2683 ) );
  ANDN U7456 ( .A(\SUBBYTES[3].a/w2775 ), .B(n2603), .Z(\SUBBYTES[3].a/w2682 )
         );
  XNOR U7457 ( .A(\w1[3][25] ), .B(\w1[3][31] ), .Z(n2603) );
  XOR U7458 ( .A(\w0[3][25] ), .B(g_input[409]), .Z(\w1[3][25] ) );
  AND U7459 ( .A(\w1[3][24] ), .B(\SUBBYTES[3].a/w2650 ), .Z(
        \SUBBYTES[3].a/w2678 ) );
  XOR U7460 ( .A(\w0[3][24] ), .B(g_input[408]), .Z(\w1[3][24] ) );
  AND U7461 ( .A(\SUBBYTES[3].a/w2651 ), .B(\SUBBYTES[3].a/w2647 ), .Z(
        \SUBBYTES[3].a/w2676 ) );
  AND U7462 ( .A(\SUBBYTES[3].a/w2736 ), .B(\SUBBYTES[3].a/w2768 ), .Z(
        \SUBBYTES[3].a/w2675 ) );
  ANDN U7463 ( .A(\SUBBYTES[3].a/w2757 ), .B(n2607), .Z(\SUBBYTES[3].a/w2670 )
         );
  XNOR U7464 ( .A(\w1[3][28] ), .B(\w1[3][31] ), .Z(n2607) );
  ANDN U7465 ( .A(\SUBBYTES[3].a/w2758 ), .B(n2608), .Z(\SUBBYTES[3].a/w2668 )
         );
  XNOR U7466 ( .A(\w1[3][26] ), .B(\w1[3][31] ), .Z(n2608) );
  XOR U7467 ( .A(\w0[3][31] ), .B(g_input[415]), .Z(\w1[3][31] ) );
  IV U7468 ( .A(n2610), .Z(\w1[3][26] ) );
  ANDN U7469 ( .A(\SUBBYTES[3].a/w2760 ), .B(n2609), .Z(\SUBBYTES[3].a/w2667 )
         );
  XOR U7470 ( .A(n2610), .B(\w1[3][28] ), .Z(n2609) );
  XOR U7471 ( .A(\w0[3][28] ), .B(g_input[412]), .Z(\w1[3][28] ) );
  XNOR U7472 ( .A(\w0[3][26] ), .B(g_input[410]), .Z(n2610) );
  AND U7473 ( .A(\SUBBYTES[3].a/w164 ), .B(n2584), .Z(\SUBBYTES[3].a/w263 ) );
  XOR U7474 ( .A(\SUBBYTES[3].a/w232 ), .B(n989), .Z(n2584) );
  AND U7475 ( .A(\SUBBYTES[3].a/w165 ), .B(n2591), .Z(\SUBBYTES[3].a/w261 ) );
  XOR U7476 ( .A(n8393), .B(\SUBBYTES[3].a/w232 ), .Z(n2591) );
  ANDN U7477 ( .A(n2592), .B(n2611), .Z(\SUBBYTES[3].a/w260 ) );
  XOR U7478 ( .A(n989), .B(n8393), .Z(n2592) );
  AND U7479 ( .A(n2612), .B(\SUBBYTES[3].a/w2437 ), .Z(\SUBBYTES[3].a/w2572 )
         );
  AND U7480 ( .A(n2613), .B(\SUBBYTES[3].a/w2438 ), .Z(\SUBBYTES[3].a/w2570 )
         );
  AND U7481 ( .A(\SUBBYTES[3].a/w2568 ), .B(n2614), .Z(\SUBBYTES[3].a/w2569 )
         );
  ANDN U7482 ( .A(\w1[3][32] ), .B(n2615), .Z(\SUBBYTES[3].a/w2565 ) );
  AND U7483 ( .A(n2616), .B(\SUBBYTES[3].a/w2440 ), .Z(\SUBBYTES[3].a/w2563 )
         );
  AND U7484 ( .A(\SUBBYTES[3].a/w2561 ), .B(n2617), .Z(\SUBBYTES[3].a/w2562 )
         );
  XOR U7485 ( .A(\SUBBYTES[3].a/w2505 ), .B(n8414), .Z(n2617) );
  ANDN U7486 ( .A(\SUBBYTES[3].a/w166 ), .B(n2593), .Z(\SUBBYTES[3].a/w256 )
         );
  XNOR U7487 ( .A(\SUBBYTES[3].a/w225 ), .B(\SUBBYTES[3].a/w228 ), .Z(n2593)
         );
  AND U7488 ( .A(\SUBBYTES[3].a/w2548 ), .B(\SUBBYTES[3].a/w2550 ), .Z(
        \SUBBYTES[3].a/w2557 ) );
  AND U7489 ( .A(\SUBBYTES[3].a/w2549 ), .B(\SUBBYTES[3].a/w2551 ), .Z(
        \SUBBYTES[3].a/w2555 ) );
  AND U7490 ( .A(\SUBBYTES[3].a/w2552 ), .B(\SUBBYTES[3].a/w2553 ), .Z(
        \SUBBYTES[3].a/w2554 ) );
  AND U7491 ( .A(\SUBBYTES[3].a/w2441 ), .B(n2612), .Z(\SUBBYTES[3].a/w2540 )
         );
  XOR U7492 ( .A(\SUBBYTES[3].a/w2509 ), .B(n1000), .Z(n2612) );
  AND U7493 ( .A(\SUBBYTES[3].a/w167 ), .B(n2595), .Z(\SUBBYTES[3].a/w254 ) );
  XNOR U7494 ( .A(n2618), .B(\SUBBYTES[3].a/w225 ), .Z(n2595) );
  AND U7495 ( .A(\SUBBYTES[3].a/w2442 ), .B(n2613), .Z(\SUBBYTES[3].a/w2538 )
         );
  XOR U7496 ( .A(n8415), .B(\SUBBYTES[3].a/w2509 ), .Z(n2613) );
  ANDN U7497 ( .A(n2614), .B(n2619), .Z(\SUBBYTES[3].a/w2537 ) );
  XOR U7498 ( .A(n1000), .B(n8415), .Z(n2614) );
  ANDN U7499 ( .A(\SUBBYTES[3].a/w2443 ), .B(n2615), .Z(\SUBBYTES[3].a/w2533 )
         );
  XNOR U7500 ( .A(\SUBBYTES[3].a/w2502 ), .B(\SUBBYTES[3].a/w2505 ), .Z(n2615)
         );
  AND U7501 ( .A(\SUBBYTES[3].a/w2444 ), .B(n2616), .Z(\SUBBYTES[3].a/w2531 )
         );
  XNOR U7502 ( .A(n2620), .B(\SUBBYTES[3].a/w2502 ), .Z(n2616) );
  AND U7503 ( .A(\SUBBYTES[3].a/w2529 ), .B(n2621), .Z(\SUBBYTES[3].a/w2530 )
         );
  XOR U7504 ( .A(n2622), .B(n2620), .Z(n2621) );
  IV U7505 ( .A(n8414), .Z(n2620) );
  AND U7506 ( .A(\SUBBYTES[3].a/w252 ), .B(n2623), .Z(\SUBBYTES[3].a/w253 ) );
  XOR U7507 ( .A(n2624), .B(n2618), .Z(n2623) );
  IV U7508 ( .A(n8392), .Z(n2618) );
  ANDN U7509 ( .A(\SUBBYTES[3].a/w2548 ), .B(n2625), .Z(\SUBBYTES[3].a/w2525 )
         );
  ANDN U7510 ( .A(\SUBBYTES[3].a/w2549 ), .B(n2626), .Z(\SUBBYTES[3].a/w2523 )
         );
  ANDN U7511 ( .A(\SUBBYTES[3].a/w2552 ), .B(n2627), .Z(\SUBBYTES[3].a/w2522 )
         );
  AND U7512 ( .A(\SUBBYTES[3].a/w2508 ), .B(\SUBBYTES[3].a/w2507 ), .Z(
        \SUBBYTES[3].a/w2509 ) );
  IV U7513 ( .A(n2622), .Z(\SUBBYTES[3].a/w2505 ) );
  NAND U7514 ( .A(\SUBBYTES[3].a/w2484 ), .B(\SUBBYTES[3].a/w2499 ), .Z(n2622)
         );
  AND U7515 ( .A(\SUBBYTES[3].a/w2501 ), .B(\SUBBYTES[3].a/w2507 ), .Z(
        \SUBBYTES[3].a/w2502 ) );
  AND U7516 ( .A(\SUBBYTES[3].a/w2486 ), .B(\SUBBYTES[3].a/w2484 ), .Z(
        \SUBBYTES[3].a/w2496 ) );
  AND U7517 ( .A(\SUBBYTES[3].a/w2487 ), .B(\SUBBYTES[3].a/w2485 ), .Z(
        \SUBBYTES[3].a/w2494 ) );
  AND U7518 ( .A(\SUBBYTES[3].a/w2501 ), .B(\SUBBYTES[3].a/w2508 ), .Z(
        \SUBBYTES[3].a/w2493 ) );
  ANDN U7519 ( .A(\SUBBYTES[3].a/w271 ), .B(n2628), .Z(\SUBBYTES[3].a/w248 )
         );
  AND U7520 ( .A(\SUBBYTES[3].a/w2441 ), .B(\SUBBYTES[3].a/w2437 ), .Z(
        \SUBBYTES[3].a/w2478 ) );
  AND U7521 ( .A(\SUBBYTES[3].a/w2442 ), .B(\SUBBYTES[3].a/w2438 ), .Z(
        \SUBBYTES[3].a/w2476 ) );
  ANDN U7522 ( .A(\SUBBYTES[3].a/w2568 ), .B(n2619), .Z(\SUBBYTES[3].a/w2475 )
         );
  XNOR U7523 ( .A(\w1[3][33] ), .B(\w1[3][39] ), .Z(n2619) );
  XOR U7524 ( .A(\w0[3][33] ), .B(g_input[417]), .Z(\w1[3][33] ) );
  AND U7525 ( .A(\w1[3][32] ), .B(\SUBBYTES[3].a/w2443 ), .Z(
        \SUBBYTES[3].a/w2471 ) );
  XOR U7526 ( .A(\w0[3][32] ), .B(g_input[416]), .Z(\w1[3][32] ) );
  AND U7527 ( .A(\SUBBYTES[3].a/w2444 ), .B(\SUBBYTES[3].a/w2440 ), .Z(
        \SUBBYTES[3].a/w2469 ) );
  AND U7528 ( .A(\SUBBYTES[3].a/w2529 ), .B(\SUBBYTES[3].a/w2561 ), .Z(
        \SUBBYTES[3].a/w2468 ) );
  ANDN U7529 ( .A(\SUBBYTES[3].a/w2550 ), .B(n2625), .Z(\SUBBYTES[3].a/w2463 )
         );
  XNOR U7530 ( .A(\w1[3][36] ), .B(\w1[3][39] ), .Z(n2625) );
  ANDN U7531 ( .A(\SUBBYTES[3].a/w2551 ), .B(n2626), .Z(\SUBBYTES[3].a/w2461 )
         );
  XNOR U7532 ( .A(\w1[3][34] ), .B(\w1[3][39] ), .Z(n2626) );
  XOR U7533 ( .A(\w0[3][39] ), .B(g_input[423]), .Z(\w1[3][39] ) );
  IV U7534 ( .A(n2629), .Z(\w1[3][34] ) );
  ANDN U7535 ( .A(\SUBBYTES[3].a/w2553 ), .B(n2627), .Z(\SUBBYTES[3].a/w2460 )
         );
  XOR U7536 ( .A(n2629), .B(\w1[3][36] ), .Z(n2627) );
  XOR U7537 ( .A(\w0[3][36] ), .B(g_input[420]), .Z(\w1[3][36] ) );
  XNOR U7538 ( .A(\w0[3][34] ), .B(g_input[418]), .Z(n2629) );
  ANDN U7539 ( .A(\SUBBYTES[3].a/w272 ), .B(n2630), .Z(\SUBBYTES[3].a/w246 )
         );
  ANDN U7540 ( .A(\SUBBYTES[3].a/w275 ), .B(n2631), .Z(\SUBBYTES[3].a/w245 )
         );
  AND U7541 ( .A(n2632), .B(\SUBBYTES[3].a/w2230 ), .Z(\SUBBYTES[3].a/w2365 )
         );
  AND U7542 ( .A(n2633), .B(\SUBBYTES[3].a/w2231 ), .Z(\SUBBYTES[3].a/w2363 )
         );
  AND U7543 ( .A(\SUBBYTES[3].a/w2361 ), .B(n2634), .Z(\SUBBYTES[3].a/w2362 )
         );
  ANDN U7544 ( .A(\w1[3][40] ), .B(n2635), .Z(\SUBBYTES[3].a/w2358 ) );
  AND U7545 ( .A(n2636), .B(\SUBBYTES[3].a/w2233 ), .Z(\SUBBYTES[3].a/w2356 )
         );
  AND U7546 ( .A(\SUBBYTES[3].a/w2354 ), .B(n2637), .Z(\SUBBYTES[3].a/w2355 )
         );
  XOR U7547 ( .A(\SUBBYTES[3].a/w2298 ), .B(n8412), .Z(n2637) );
  AND U7548 ( .A(\SUBBYTES[3].a/w2341 ), .B(\SUBBYTES[3].a/w2343 ), .Z(
        \SUBBYTES[3].a/w2350 ) );
  AND U7549 ( .A(\SUBBYTES[3].a/w2342 ), .B(\SUBBYTES[3].a/w2344 ), .Z(
        \SUBBYTES[3].a/w2348 ) );
  AND U7550 ( .A(\SUBBYTES[3].a/w2345 ), .B(\SUBBYTES[3].a/w2346 ), .Z(
        \SUBBYTES[3].a/w2347 ) );
  AND U7551 ( .A(\SUBBYTES[3].a/w2234 ), .B(n2632), .Z(\SUBBYTES[3].a/w2333 )
         );
  XOR U7552 ( .A(\SUBBYTES[3].a/w2302 ), .B(n999), .Z(n2632) );
  AND U7553 ( .A(\SUBBYTES[3].a/w2235 ), .B(n2633), .Z(\SUBBYTES[3].a/w2331 )
         );
  XOR U7554 ( .A(n8413), .B(\SUBBYTES[3].a/w2302 ), .Z(n2633) );
  ANDN U7555 ( .A(n2634), .B(n2638), .Z(\SUBBYTES[3].a/w2330 ) );
  XOR U7556 ( .A(n999), .B(n8413), .Z(n2634) );
  ANDN U7557 ( .A(\SUBBYTES[3].a/w2236 ), .B(n2635), .Z(\SUBBYTES[3].a/w2326 )
         );
  XNOR U7558 ( .A(\SUBBYTES[3].a/w2295 ), .B(\SUBBYTES[3].a/w2298 ), .Z(n2635)
         );
  AND U7559 ( .A(\SUBBYTES[3].a/w2237 ), .B(n2636), .Z(\SUBBYTES[3].a/w2324 )
         );
  XNOR U7560 ( .A(n2639), .B(\SUBBYTES[3].a/w2295 ), .Z(n2636) );
  AND U7561 ( .A(\SUBBYTES[3].a/w2322 ), .B(n2640), .Z(\SUBBYTES[3].a/w2323 )
         );
  XOR U7562 ( .A(n2641), .B(n2639), .Z(n2640) );
  IV U7563 ( .A(n8412), .Z(n2639) );
  AND U7564 ( .A(\SUBBYTES[3].a/w231 ), .B(\SUBBYTES[3].a/w230 ), .Z(
        \SUBBYTES[3].a/w232 ) );
  ANDN U7565 ( .A(\SUBBYTES[3].a/w2341 ), .B(n2642), .Z(\SUBBYTES[3].a/w2318 )
         );
  ANDN U7566 ( .A(\SUBBYTES[3].a/w2342 ), .B(n2643), .Z(\SUBBYTES[3].a/w2316 )
         );
  ANDN U7567 ( .A(\SUBBYTES[3].a/w2345 ), .B(n2644), .Z(\SUBBYTES[3].a/w2315 )
         );
  AND U7568 ( .A(\SUBBYTES[3].a/w2301 ), .B(\SUBBYTES[3].a/w2300 ), .Z(
        \SUBBYTES[3].a/w2302 ) );
  IV U7569 ( .A(n2641), .Z(\SUBBYTES[3].a/w2298 ) );
  NAND U7570 ( .A(\SUBBYTES[3].a/w2277 ), .B(\SUBBYTES[3].a/w2292 ), .Z(n2641)
         );
  AND U7571 ( .A(\SUBBYTES[3].a/w2294 ), .B(\SUBBYTES[3].a/w2300 ), .Z(
        \SUBBYTES[3].a/w2295 ) );
  AND U7572 ( .A(\SUBBYTES[3].a/w2279 ), .B(\SUBBYTES[3].a/w2277 ), .Z(
        \SUBBYTES[3].a/w2289 ) );
  AND U7573 ( .A(\SUBBYTES[3].a/w2280 ), .B(\SUBBYTES[3].a/w2278 ), .Z(
        \SUBBYTES[3].a/w2287 ) );
  AND U7574 ( .A(\SUBBYTES[3].a/w2294 ), .B(\SUBBYTES[3].a/w2301 ), .Z(
        \SUBBYTES[3].a/w2286 ) );
  IV U7575 ( .A(n2624), .Z(\SUBBYTES[3].a/w228 ) );
  NAND U7576 ( .A(\SUBBYTES[3].a/w207 ), .B(\SUBBYTES[3].a/w222 ), .Z(n2624)
         );
  AND U7577 ( .A(\SUBBYTES[3].a/w2234 ), .B(\SUBBYTES[3].a/w2230 ), .Z(
        \SUBBYTES[3].a/w2271 ) );
  AND U7578 ( .A(\SUBBYTES[3].a/w2235 ), .B(\SUBBYTES[3].a/w2231 ), .Z(
        \SUBBYTES[3].a/w2269 ) );
  ANDN U7579 ( .A(\SUBBYTES[3].a/w2361 ), .B(n2638), .Z(\SUBBYTES[3].a/w2268 )
         );
  XNOR U7580 ( .A(\w1[3][41] ), .B(\w1[3][47] ), .Z(n2638) );
  XOR U7581 ( .A(\w0[3][41] ), .B(g_input[425]), .Z(\w1[3][41] ) );
  AND U7582 ( .A(\w1[3][40] ), .B(\SUBBYTES[3].a/w2236 ), .Z(
        \SUBBYTES[3].a/w2264 ) );
  XOR U7583 ( .A(\w0[3][40] ), .B(g_input[424]), .Z(\w1[3][40] ) );
  AND U7584 ( .A(\SUBBYTES[3].a/w2237 ), .B(\SUBBYTES[3].a/w2233 ), .Z(
        \SUBBYTES[3].a/w2262 ) );
  AND U7585 ( .A(\SUBBYTES[3].a/w2322 ), .B(\SUBBYTES[3].a/w2354 ), .Z(
        \SUBBYTES[3].a/w2261 ) );
  ANDN U7586 ( .A(\SUBBYTES[3].a/w2343 ), .B(n2642), .Z(\SUBBYTES[3].a/w2256 )
         );
  XNOR U7587 ( .A(\w1[3][44] ), .B(\w1[3][47] ), .Z(n2642) );
  ANDN U7588 ( .A(\SUBBYTES[3].a/w2344 ), .B(n2643), .Z(\SUBBYTES[3].a/w2254 )
         );
  XNOR U7589 ( .A(\w1[3][42] ), .B(\w1[3][47] ), .Z(n2643) );
  XOR U7590 ( .A(\w0[3][47] ), .B(g_input[431]), .Z(\w1[3][47] ) );
  IV U7591 ( .A(n2645), .Z(\w1[3][42] ) );
  ANDN U7592 ( .A(\SUBBYTES[3].a/w2346 ), .B(n2644), .Z(\SUBBYTES[3].a/w2253 )
         );
  XOR U7593 ( .A(n2645), .B(\w1[3][44] ), .Z(n2644) );
  XOR U7594 ( .A(\w0[3][44] ), .B(g_input[428]), .Z(\w1[3][44] ) );
  XNOR U7595 ( .A(\w0[3][42] ), .B(g_input[426]), .Z(n2645) );
  AND U7596 ( .A(\SUBBYTES[3].a/w224 ), .B(\SUBBYTES[3].a/w230 ), .Z(
        \SUBBYTES[3].a/w225 ) );
  AND U7597 ( .A(\SUBBYTES[3].a/w209 ), .B(\SUBBYTES[3].a/w207 ), .Z(
        \SUBBYTES[3].a/w219 ) );
  AND U7598 ( .A(\SUBBYTES[3].a/w210 ), .B(\SUBBYTES[3].a/w208 ), .Z(
        \SUBBYTES[3].a/w217 ) );
  AND U7599 ( .A(\SUBBYTES[3].a/w224 ), .B(\SUBBYTES[3].a/w231 ), .Z(
        \SUBBYTES[3].a/w216 ) );
  AND U7600 ( .A(n2646), .B(\SUBBYTES[3].a/w2023 ), .Z(\SUBBYTES[3].a/w2158 )
         );
  AND U7601 ( .A(n2647), .B(\SUBBYTES[3].a/w2024 ), .Z(\SUBBYTES[3].a/w2156 )
         );
  AND U7602 ( .A(\SUBBYTES[3].a/w2154 ), .B(n2648), .Z(\SUBBYTES[3].a/w2155 )
         );
  ANDN U7603 ( .A(\w1[3][48] ), .B(n2649), .Z(\SUBBYTES[3].a/w2151 ) );
  AND U7604 ( .A(n2650), .B(\SUBBYTES[3].a/w2026 ), .Z(\SUBBYTES[3].a/w2149 )
         );
  AND U7605 ( .A(\SUBBYTES[3].a/w2147 ), .B(n2651), .Z(\SUBBYTES[3].a/w2148 )
         );
  XOR U7606 ( .A(\SUBBYTES[3].a/w2091 ), .B(n8410), .Z(n2651) );
  AND U7607 ( .A(\SUBBYTES[3].a/w2134 ), .B(\SUBBYTES[3].a/w2136 ), .Z(
        \SUBBYTES[3].a/w2143 ) );
  AND U7608 ( .A(\SUBBYTES[3].a/w2135 ), .B(\SUBBYTES[3].a/w2137 ), .Z(
        \SUBBYTES[3].a/w2141 ) );
  AND U7609 ( .A(\SUBBYTES[3].a/w2138 ), .B(\SUBBYTES[3].a/w2139 ), .Z(
        \SUBBYTES[3].a/w2140 ) );
  AND U7610 ( .A(\SUBBYTES[3].a/w2027 ), .B(n2646), .Z(\SUBBYTES[3].a/w2126 )
         );
  XOR U7611 ( .A(\SUBBYTES[3].a/w2095 ), .B(n998), .Z(n2646) );
  AND U7612 ( .A(\SUBBYTES[3].a/w2028 ), .B(n2647), .Z(\SUBBYTES[3].a/w2124 )
         );
  XOR U7613 ( .A(n8411), .B(\SUBBYTES[3].a/w2095 ), .Z(n2647) );
  ANDN U7614 ( .A(n2648), .B(n2652), .Z(\SUBBYTES[3].a/w2123 ) );
  XOR U7615 ( .A(n998), .B(n8411), .Z(n2648) );
  ANDN U7616 ( .A(\SUBBYTES[3].a/w2029 ), .B(n2649), .Z(\SUBBYTES[3].a/w2119 )
         );
  XNOR U7617 ( .A(\SUBBYTES[3].a/w2088 ), .B(\SUBBYTES[3].a/w2091 ), .Z(n2649)
         );
  AND U7618 ( .A(\SUBBYTES[3].a/w2030 ), .B(n2650), .Z(\SUBBYTES[3].a/w2117 )
         );
  XNOR U7619 ( .A(n2653), .B(\SUBBYTES[3].a/w2088 ), .Z(n2650) );
  AND U7620 ( .A(\SUBBYTES[3].a/w2115 ), .B(n2654), .Z(\SUBBYTES[3].a/w2116 )
         );
  XOR U7621 ( .A(n2655), .B(n2653), .Z(n2654) );
  IV U7622 ( .A(n8410), .Z(n2653) );
  ANDN U7623 ( .A(\SUBBYTES[3].a/w2134 ), .B(n2656), .Z(\SUBBYTES[3].a/w2111 )
         );
  ANDN U7624 ( .A(\SUBBYTES[3].a/w2135 ), .B(n2657), .Z(\SUBBYTES[3].a/w2109 )
         );
  ANDN U7625 ( .A(\SUBBYTES[3].a/w2138 ), .B(n2658), .Z(\SUBBYTES[3].a/w2108 )
         );
  AND U7626 ( .A(\SUBBYTES[3].a/w2094 ), .B(\SUBBYTES[3].a/w2093 ), .Z(
        \SUBBYTES[3].a/w2095 ) );
  IV U7627 ( .A(n2655), .Z(\SUBBYTES[3].a/w2091 ) );
  NAND U7628 ( .A(\SUBBYTES[3].a/w2070 ), .B(\SUBBYTES[3].a/w2085 ), .Z(n2655)
         );
  AND U7629 ( .A(\SUBBYTES[3].a/w2087 ), .B(\SUBBYTES[3].a/w2093 ), .Z(
        \SUBBYTES[3].a/w2088 ) );
  AND U7630 ( .A(\SUBBYTES[3].a/w2072 ), .B(\SUBBYTES[3].a/w2070 ), .Z(
        \SUBBYTES[3].a/w2082 ) );
  AND U7631 ( .A(\SUBBYTES[3].a/w2073 ), .B(\SUBBYTES[3].a/w2071 ), .Z(
        \SUBBYTES[3].a/w2080 ) );
  AND U7632 ( .A(\SUBBYTES[3].a/w2087 ), .B(\SUBBYTES[3].a/w2094 ), .Z(
        \SUBBYTES[3].a/w2079 ) );
  AND U7633 ( .A(\SUBBYTES[3].a/w2027 ), .B(\SUBBYTES[3].a/w2023 ), .Z(
        \SUBBYTES[3].a/w2064 ) );
  AND U7634 ( .A(\SUBBYTES[3].a/w2028 ), .B(\SUBBYTES[3].a/w2024 ), .Z(
        \SUBBYTES[3].a/w2062 ) );
  ANDN U7635 ( .A(\SUBBYTES[3].a/w2154 ), .B(n2652), .Z(\SUBBYTES[3].a/w2061 )
         );
  XNOR U7636 ( .A(\w1[3][49] ), .B(\w1[3][55] ), .Z(n2652) );
  XOR U7637 ( .A(\w0[3][49] ), .B(g_input[433]), .Z(\w1[3][49] ) );
  AND U7638 ( .A(\w1[3][48] ), .B(\SUBBYTES[3].a/w2029 ), .Z(
        \SUBBYTES[3].a/w2057 ) );
  XOR U7639 ( .A(\w0[3][48] ), .B(g_input[432]), .Z(\w1[3][48] ) );
  AND U7640 ( .A(\SUBBYTES[3].a/w2030 ), .B(\SUBBYTES[3].a/w2026 ), .Z(
        \SUBBYTES[3].a/w2055 ) );
  AND U7641 ( .A(\SUBBYTES[3].a/w2115 ), .B(\SUBBYTES[3].a/w2147 ), .Z(
        \SUBBYTES[3].a/w2054 ) );
  ANDN U7642 ( .A(\SUBBYTES[3].a/w2136 ), .B(n2656), .Z(\SUBBYTES[3].a/w2049 )
         );
  XNOR U7643 ( .A(\w1[3][52] ), .B(\w1[3][55] ), .Z(n2656) );
  ANDN U7644 ( .A(\SUBBYTES[3].a/w2137 ), .B(n2657), .Z(\SUBBYTES[3].a/w2047 )
         );
  XNOR U7645 ( .A(\w1[3][50] ), .B(\w1[3][55] ), .Z(n2657) );
  XOR U7646 ( .A(\w0[3][55] ), .B(g_input[439]), .Z(\w1[3][55] ) );
  IV U7647 ( .A(n2659), .Z(\w1[3][50] ) );
  ANDN U7648 ( .A(\SUBBYTES[3].a/w2139 ), .B(n2658), .Z(\SUBBYTES[3].a/w2046 )
         );
  XOR U7649 ( .A(n2659), .B(\w1[3][52] ), .Z(n2658) );
  XOR U7650 ( .A(\w0[3][52] ), .B(g_input[436]), .Z(\w1[3][52] ) );
  XNOR U7651 ( .A(\w0[3][50] ), .B(g_input[434]), .Z(n2659) );
  AND U7652 ( .A(\SUBBYTES[3].a/w164 ), .B(\SUBBYTES[3].a/w160 ), .Z(
        \SUBBYTES[3].a/w201 ) );
  AND U7653 ( .A(\SUBBYTES[3].a/w165 ), .B(\SUBBYTES[3].a/w161 ), .Z(
        \SUBBYTES[3].a/w199 ) );
  ANDN U7654 ( .A(\SUBBYTES[3].a/w291 ), .B(n2611), .Z(\SUBBYTES[3].a/w198 )
         );
  XNOR U7655 ( .A(\w1[3][121] ), .B(\w1[3][127] ), .Z(n2611) );
  XOR U7656 ( .A(\w0[3][121] ), .B(g_input[505]), .Z(\w1[3][121] ) );
  AND U7657 ( .A(n2660), .B(\SUBBYTES[3].a/w1816 ), .Z(\SUBBYTES[3].a/w1951 )
         );
  AND U7658 ( .A(n2661), .B(\SUBBYTES[3].a/w1817 ), .Z(\SUBBYTES[3].a/w1949 )
         );
  AND U7659 ( .A(\SUBBYTES[3].a/w1947 ), .B(n2662), .Z(\SUBBYTES[3].a/w1948 )
         );
  ANDN U7660 ( .A(\w1[3][56] ), .B(n2663), .Z(\SUBBYTES[3].a/w1944 ) );
  AND U7661 ( .A(n2664), .B(\SUBBYTES[3].a/w1819 ), .Z(\SUBBYTES[3].a/w1942 )
         );
  AND U7662 ( .A(\SUBBYTES[3].a/w1940 ), .B(n2665), .Z(\SUBBYTES[3].a/w1941 )
         );
  XOR U7663 ( .A(\SUBBYTES[3].a/w1884 ), .B(n8408), .Z(n2665) );
  AND U7664 ( .A(\w1[3][120] ), .B(\SUBBYTES[3].a/w166 ), .Z(
        \SUBBYTES[3].a/w194 ) );
  XOR U7665 ( .A(\w0[3][120] ), .B(g_input[504]), .Z(\w1[3][120] ) );
  AND U7666 ( .A(\SUBBYTES[3].a/w1927 ), .B(\SUBBYTES[3].a/w1929 ), .Z(
        \SUBBYTES[3].a/w1936 ) );
  AND U7667 ( .A(\SUBBYTES[3].a/w1928 ), .B(\SUBBYTES[3].a/w1930 ), .Z(
        \SUBBYTES[3].a/w1934 ) );
  AND U7668 ( .A(\SUBBYTES[3].a/w1931 ), .B(\SUBBYTES[3].a/w1932 ), .Z(
        \SUBBYTES[3].a/w1933 ) );
  AND U7669 ( .A(\SUBBYTES[3].a/w167 ), .B(\SUBBYTES[3].a/w163 ), .Z(
        \SUBBYTES[3].a/w192 ) );
  AND U7670 ( .A(\SUBBYTES[3].a/w1820 ), .B(n2660), .Z(\SUBBYTES[3].a/w1919 )
         );
  XOR U7671 ( .A(\SUBBYTES[3].a/w1888 ), .B(n997), .Z(n2660) );
  AND U7672 ( .A(\SUBBYTES[3].a/w1821 ), .B(n2661), .Z(\SUBBYTES[3].a/w1917 )
         );
  XOR U7673 ( .A(n8409), .B(\SUBBYTES[3].a/w1888 ), .Z(n2661) );
  ANDN U7674 ( .A(n2662), .B(n2666), .Z(\SUBBYTES[3].a/w1916 ) );
  XOR U7675 ( .A(n997), .B(n8409), .Z(n2662) );
  ANDN U7676 ( .A(\SUBBYTES[3].a/w1822 ), .B(n2663), .Z(\SUBBYTES[3].a/w1912 )
         );
  XNOR U7677 ( .A(\SUBBYTES[3].a/w1881 ), .B(\SUBBYTES[3].a/w1884 ), .Z(n2663)
         );
  AND U7678 ( .A(\SUBBYTES[3].a/w1823 ), .B(n2664), .Z(\SUBBYTES[3].a/w1910 )
         );
  XNOR U7679 ( .A(n2667), .B(\SUBBYTES[3].a/w1881 ), .Z(n2664) );
  AND U7680 ( .A(\SUBBYTES[3].a/w252 ), .B(\SUBBYTES[3].a/w284 ), .Z(
        \SUBBYTES[3].a/w191 ) );
  AND U7681 ( .A(\SUBBYTES[3].a/w1908 ), .B(n2668), .Z(\SUBBYTES[3].a/w1909 )
         );
  XOR U7682 ( .A(n2669), .B(n2667), .Z(n2668) );
  IV U7683 ( .A(n8408), .Z(n2667) );
  ANDN U7684 ( .A(\SUBBYTES[3].a/w1927 ), .B(n2670), .Z(\SUBBYTES[3].a/w1904 )
         );
  ANDN U7685 ( .A(\SUBBYTES[3].a/w1928 ), .B(n2671), .Z(\SUBBYTES[3].a/w1902 )
         );
  ANDN U7686 ( .A(\SUBBYTES[3].a/w1931 ), .B(n2672), .Z(\SUBBYTES[3].a/w1901 )
         );
  AND U7687 ( .A(\SUBBYTES[3].a/w1887 ), .B(\SUBBYTES[3].a/w1886 ), .Z(
        \SUBBYTES[3].a/w1888 ) );
  IV U7688 ( .A(n2669), .Z(\SUBBYTES[3].a/w1884 ) );
  NAND U7689 ( .A(\SUBBYTES[3].a/w1863 ), .B(\SUBBYTES[3].a/w1878 ), .Z(n2669)
         );
  AND U7690 ( .A(\SUBBYTES[3].a/w1880 ), .B(\SUBBYTES[3].a/w1886 ), .Z(
        \SUBBYTES[3].a/w1881 ) );
  AND U7691 ( .A(\SUBBYTES[3].a/w1865 ), .B(\SUBBYTES[3].a/w1863 ), .Z(
        \SUBBYTES[3].a/w1875 ) );
  AND U7692 ( .A(\SUBBYTES[3].a/w1866 ), .B(\SUBBYTES[3].a/w1864 ), .Z(
        \SUBBYTES[3].a/w1873 ) );
  AND U7693 ( .A(\SUBBYTES[3].a/w1880 ), .B(\SUBBYTES[3].a/w1887 ), .Z(
        \SUBBYTES[3].a/w1872 ) );
  ANDN U7694 ( .A(\SUBBYTES[3].a/w273 ), .B(n2628), .Z(\SUBBYTES[3].a/w186 )
         );
  XNOR U7695 ( .A(\w1[3][124] ), .B(\w1[3][127] ), .Z(n2628) );
  AND U7696 ( .A(\SUBBYTES[3].a/w1820 ), .B(\SUBBYTES[3].a/w1816 ), .Z(
        \SUBBYTES[3].a/w1857 ) );
  AND U7697 ( .A(\SUBBYTES[3].a/w1821 ), .B(\SUBBYTES[3].a/w1817 ), .Z(
        \SUBBYTES[3].a/w1855 ) );
  ANDN U7698 ( .A(\SUBBYTES[3].a/w1947 ), .B(n2666), .Z(\SUBBYTES[3].a/w1854 )
         );
  XNOR U7699 ( .A(\w1[3][57] ), .B(\w1[3][63] ), .Z(n2666) );
  XOR U7700 ( .A(\w0[3][57] ), .B(g_input[441]), .Z(\w1[3][57] ) );
  AND U7701 ( .A(\w1[3][56] ), .B(\SUBBYTES[3].a/w1822 ), .Z(
        \SUBBYTES[3].a/w1850 ) );
  XOR U7702 ( .A(\w0[3][56] ), .B(g_input[440]), .Z(\w1[3][56] ) );
  AND U7703 ( .A(\SUBBYTES[3].a/w1823 ), .B(\SUBBYTES[3].a/w1819 ), .Z(
        \SUBBYTES[3].a/w1848 ) );
  AND U7704 ( .A(\SUBBYTES[3].a/w1908 ), .B(\SUBBYTES[3].a/w1940 ), .Z(
        \SUBBYTES[3].a/w1847 ) );
  ANDN U7705 ( .A(\SUBBYTES[3].a/w1929 ), .B(n2670), .Z(\SUBBYTES[3].a/w1842 )
         );
  XNOR U7706 ( .A(\w1[3][60] ), .B(\w1[3][63] ), .Z(n2670) );
  ANDN U7707 ( .A(\SUBBYTES[3].a/w1930 ), .B(n2671), .Z(\SUBBYTES[3].a/w1840 )
         );
  XNOR U7708 ( .A(\w1[3][58] ), .B(\w1[3][63] ), .Z(n2671) );
  XOR U7709 ( .A(\w0[3][63] ), .B(g_input[447]), .Z(\w1[3][63] ) );
  IV U7710 ( .A(n2673), .Z(\w1[3][58] ) );
  ANDN U7711 ( .A(\SUBBYTES[3].a/w274 ), .B(n2630), .Z(\SUBBYTES[3].a/w184 )
         );
  XNOR U7712 ( .A(\w1[3][122] ), .B(\w1[3][127] ), .Z(n2630) );
  XOR U7713 ( .A(\w0[3][127] ), .B(g_input[511]), .Z(\w1[3][127] ) );
  IV U7714 ( .A(n2674), .Z(\w1[3][122] ) );
  ANDN U7715 ( .A(\SUBBYTES[3].a/w1932 ), .B(n2672), .Z(\SUBBYTES[3].a/w1839 )
         );
  XOR U7716 ( .A(n2673), .B(\w1[3][60] ), .Z(n2672) );
  XOR U7717 ( .A(\w0[3][60] ), .B(g_input[444]), .Z(\w1[3][60] ) );
  XNOR U7718 ( .A(\w0[3][58] ), .B(g_input[442]), .Z(n2673) );
  ANDN U7719 ( .A(\SUBBYTES[3].a/w276 ), .B(n2631), .Z(\SUBBYTES[3].a/w183 )
         );
  XOR U7720 ( .A(n2674), .B(\w1[3][124] ), .Z(n2631) );
  XOR U7721 ( .A(\w0[3][124] ), .B(g_input[508]), .Z(\w1[3][124] ) );
  XNOR U7722 ( .A(\w0[3][122] ), .B(g_input[506]), .Z(n2674) );
  AND U7723 ( .A(n2675), .B(\SUBBYTES[3].a/w1609 ), .Z(\SUBBYTES[3].a/w1744 )
         );
  AND U7724 ( .A(n2676), .B(\SUBBYTES[3].a/w1610 ), .Z(\SUBBYTES[3].a/w1742 )
         );
  AND U7725 ( .A(\SUBBYTES[3].a/w1740 ), .B(n2677), .Z(\SUBBYTES[3].a/w1741 )
         );
  ANDN U7726 ( .A(\w1[3][64] ), .B(n2678), .Z(\SUBBYTES[3].a/w1737 ) );
  AND U7727 ( .A(n2679), .B(\SUBBYTES[3].a/w1612 ), .Z(\SUBBYTES[3].a/w1735 )
         );
  AND U7728 ( .A(\SUBBYTES[3].a/w1733 ), .B(n2680), .Z(\SUBBYTES[3].a/w1734 )
         );
  XOR U7729 ( .A(\SUBBYTES[3].a/w1677 ), .B(n8406), .Z(n2680) );
  AND U7730 ( .A(\SUBBYTES[3].a/w1720 ), .B(\SUBBYTES[3].a/w1722 ), .Z(
        \SUBBYTES[3].a/w1729 ) );
  AND U7731 ( .A(\SUBBYTES[3].a/w1721 ), .B(\SUBBYTES[3].a/w1723 ), .Z(
        \SUBBYTES[3].a/w1727 ) );
  AND U7732 ( .A(\SUBBYTES[3].a/w1724 ), .B(\SUBBYTES[3].a/w1725 ), .Z(
        \SUBBYTES[3].a/w1726 ) );
  AND U7733 ( .A(\SUBBYTES[3].a/w1613 ), .B(n2675), .Z(\SUBBYTES[3].a/w1712 )
         );
  XOR U7734 ( .A(\SUBBYTES[3].a/w1681 ), .B(n996), .Z(n2675) );
  AND U7735 ( .A(\SUBBYTES[3].a/w1614 ), .B(n2676), .Z(\SUBBYTES[3].a/w1710 )
         );
  XOR U7736 ( .A(n8407), .B(\SUBBYTES[3].a/w1681 ), .Z(n2676) );
  ANDN U7737 ( .A(n2677), .B(n2681), .Z(\SUBBYTES[3].a/w1709 ) );
  XOR U7738 ( .A(n996), .B(n8407), .Z(n2677) );
  ANDN U7739 ( .A(\SUBBYTES[3].a/w1615 ), .B(n2678), .Z(\SUBBYTES[3].a/w1705 )
         );
  XNOR U7740 ( .A(\SUBBYTES[3].a/w1674 ), .B(\SUBBYTES[3].a/w1677 ), .Z(n2678)
         );
  AND U7741 ( .A(\SUBBYTES[3].a/w1616 ), .B(n2679), .Z(\SUBBYTES[3].a/w1703 )
         );
  XNOR U7742 ( .A(n2682), .B(\SUBBYTES[3].a/w1674 ), .Z(n2679) );
  AND U7743 ( .A(\SUBBYTES[3].a/w1701 ), .B(n2683), .Z(\SUBBYTES[3].a/w1702 )
         );
  XOR U7744 ( .A(n2684), .B(n2682), .Z(n2683) );
  IV U7745 ( .A(n8406), .Z(n2682) );
  ANDN U7746 ( .A(\SUBBYTES[3].a/w1720 ), .B(n2685), .Z(\SUBBYTES[3].a/w1697 )
         );
  ANDN U7747 ( .A(\SUBBYTES[3].a/w1721 ), .B(n2686), .Z(\SUBBYTES[3].a/w1695 )
         );
  ANDN U7748 ( .A(\SUBBYTES[3].a/w1724 ), .B(n2687), .Z(\SUBBYTES[3].a/w1694 )
         );
  AND U7749 ( .A(\SUBBYTES[3].a/w1680 ), .B(\SUBBYTES[3].a/w1679 ), .Z(
        \SUBBYTES[3].a/w1681 ) );
  IV U7750 ( .A(n2684), .Z(\SUBBYTES[3].a/w1677 ) );
  NAND U7751 ( .A(\SUBBYTES[3].a/w1656 ), .B(\SUBBYTES[3].a/w1671 ), .Z(n2684)
         );
  AND U7752 ( .A(\SUBBYTES[3].a/w1673 ), .B(\SUBBYTES[3].a/w1679 ), .Z(
        \SUBBYTES[3].a/w1674 ) );
  AND U7753 ( .A(\SUBBYTES[3].a/w1658 ), .B(\SUBBYTES[3].a/w1656 ), .Z(
        \SUBBYTES[3].a/w1668 ) );
  AND U7754 ( .A(\SUBBYTES[3].a/w1659 ), .B(\SUBBYTES[3].a/w1657 ), .Z(
        \SUBBYTES[3].a/w1666 ) );
  AND U7755 ( .A(\SUBBYTES[3].a/w1673 ), .B(\SUBBYTES[3].a/w1680 ), .Z(
        \SUBBYTES[3].a/w1665 ) );
  AND U7756 ( .A(\SUBBYTES[3].a/w1613 ), .B(\SUBBYTES[3].a/w1609 ), .Z(
        \SUBBYTES[3].a/w1650 ) );
  AND U7757 ( .A(\SUBBYTES[3].a/w1614 ), .B(\SUBBYTES[3].a/w1610 ), .Z(
        \SUBBYTES[3].a/w1648 ) );
  ANDN U7758 ( .A(\SUBBYTES[3].a/w1740 ), .B(n2681), .Z(\SUBBYTES[3].a/w1647 )
         );
  XNOR U7759 ( .A(\w1[3][65] ), .B(\w1[3][71] ), .Z(n2681) );
  XOR U7760 ( .A(\w0[3][65] ), .B(g_input[449]), .Z(\w1[3][65] ) );
  AND U7761 ( .A(\w1[3][64] ), .B(\SUBBYTES[3].a/w1615 ), .Z(
        \SUBBYTES[3].a/w1643 ) );
  XOR U7762 ( .A(\w0[3][64] ), .B(g_input[448]), .Z(\w1[3][64] ) );
  AND U7763 ( .A(\SUBBYTES[3].a/w1616 ), .B(\SUBBYTES[3].a/w1612 ), .Z(
        \SUBBYTES[3].a/w1641 ) );
  AND U7764 ( .A(\SUBBYTES[3].a/w1701 ), .B(\SUBBYTES[3].a/w1733 ), .Z(
        \SUBBYTES[3].a/w1640 ) );
  ANDN U7765 ( .A(\SUBBYTES[3].a/w1722 ), .B(n2685), .Z(\SUBBYTES[3].a/w1635 )
         );
  XNOR U7766 ( .A(\w1[3][68] ), .B(\w1[3][71] ), .Z(n2685) );
  ANDN U7767 ( .A(\SUBBYTES[3].a/w1723 ), .B(n2686), .Z(\SUBBYTES[3].a/w1633 )
         );
  XNOR U7768 ( .A(\w1[3][66] ), .B(\w1[3][71] ), .Z(n2686) );
  XOR U7769 ( .A(\w0[3][71] ), .B(g_input[455]), .Z(\w1[3][71] ) );
  IV U7770 ( .A(n2688), .Z(\w1[3][66] ) );
  ANDN U7771 ( .A(\SUBBYTES[3].a/w1725 ), .B(n2687), .Z(\SUBBYTES[3].a/w1632 )
         );
  XOR U7772 ( .A(n2688), .B(\w1[3][68] ), .Z(n2687) );
  XOR U7773 ( .A(\w0[3][68] ), .B(g_input[452]), .Z(\w1[3][68] ) );
  XNOR U7774 ( .A(\w0[3][66] ), .B(g_input[450]), .Z(n2688) );
  AND U7775 ( .A(n2689), .B(\SUBBYTES[3].a/w1402 ), .Z(\SUBBYTES[3].a/w1537 )
         );
  AND U7776 ( .A(n2690), .B(\SUBBYTES[3].a/w1403 ), .Z(\SUBBYTES[3].a/w1535 )
         );
  AND U7777 ( .A(\SUBBYTES[3].a/w1533 ), .B(n2691), .Z(\SUBBYTES[3].a/w1534 )
         );
  ANDN U7778 ( .A(\w1[3][72] ), .B(n2692), .Z(\SUBBYTES[3].a/w1530 ) );
  AND U7779 ( .A(n2693), .B(\SUBBYTES[3].a/w1405 ), .Z(\SUBBYTES[3].a/w1528 )
         );
  AND U7780 ( .A(\SUBBYTES[3].a/w1526 ), .B(n2694), .Z(\SUBBYTES[3].a/w1527 )
         );
  XOR U7781 ( .A(\SUBBYTES[3].a/w1470 ), .B(n8404), .Z(n2694) );
  AND U7782 ( .A(\SUBBYTES[3].a/w1513 ), .B(\SUBBYTES[3].a/w1515 ), .Z(
        \SUBBYTES[3].a/w1522 ) );
  AND U7783 ( .A(\SUBBYTES[3].a/w1514 ), .B(\SUBBYTES[3].a/w1516 ), .Z(
        \SUBBYTES[3].a/w1520 ) );
  AND U7784 ( .A(\SUBBYTES[3].a/w1517 ), .B(\SUBBYTES[3].a/w1518 ), .Z(
        \SUBBYTES[3].a/w1519 ) );
  AND U7785 ( .A(\SUBBYTES[3].a/w1406 ), .B(n2689), .Z(\SUBBYTES[3].a/w1505 )
         );
  XOR U7786 ( .A(\SUBBYTES[3].a/w1474 ), .B(n995), .Z(n2689) );
  AND U7787 ( .A(\SUBBYTES[3].a/w1407 ), .B(n2690), .Z(\SUBBYTES[3].a/w1503 )
         );
  XOR U7788 ( .A(n8405), .B(\SUBBYTES[3].a/w1474 ), .Z(n2690) );
  ANDN U7789 ( .A(n2691), .B(n2695), .Z(\SUBBYTES[3].a/w1502 ) );
  XOR U7790 ( .A(n995), .B(n8405), .Z(n2691) );
  ANDN U7791 ( .A(\SUBBYTES[3].a/w1408 ), .B(n2692), .Z(\SUBBYTES[3].a/w1498 )
         );
  XNOR U7792 ( .A(\SUBBYTES[3].a/w1467 ), .B(\SUBBYTES[3].a/w1470 ), .Z(n2692)
         );
  AND U7793 ( .A(\SUBBYTES[3].a/w1409 ), .B(n2693), .Z(\SUBBYTES[3].a/w1496 )
         );
  XNOR U7794 ( .A(n2696), .B(\SUBBYTES[3].a/w1467 ), .Z(n2693) );
  AND U7795 ( .A(\SUBBYTES[3].a/w1494 ), .B(n2697), .Z(\SUBBYTES[3].a/w1495 )
         );
  XOR U7796 ( .A(n2698), .B(n2696), .Z(n2697) );
  IV U7797 ( .A(n8404), .Z(n2696) );
  ANDN U7798 ( .A(\SUBBYTES[3].a/w1513 ), .B(n2699), .Z(\SUBBYTES[3].a/w1490 )
         );
  ANDN U7799 ( .A(\SUBBYTES[3].a/w1514 ), .B(n2700), .Z(\SUBBYTES[3].a/w1488 )
         );
  ANDN U7800 ( .A(\SUBBYTES[3].a/w1517 ), .B(n2701), .Z(\SUBBYTES[3].a/w1487 )
         );
  AND U7801 ( .A(\SUBBYTES[3].a/w1473 ), .B(\SUBBYTES[3].a/w1472 ), .Z(
        \SUBBYTES[3].a/w1474 ) );
  IV U7802 ( .A(n2698), .Z(\SUBBYTES[3].a/w1470 ) );
  NAND U7803 ( .A(\SUBBYTES[3].a/w1449 ), .B(\SUBBYTES[3].a/w1464 ), .Z(n2698)
         );
  AND U7804 ( .A(\SUBBYTES[3].a/w1466 ), .B(\SUBBYTES[3].a/w1472 ), .Z(
        \SUBBYTES[3].a/w1467 ) );
  AND U7805 ( .A(\SUBBYTES[3].a/w1451 ), .B(\SUBBYTES[3].a/w1449 ), .Z(
        \SUBBYTES[3].a/w1461 ) );
  AND U7806 ( .A(\SUBBYTES[3].a/w1452 ), .B(\SUBBYTES[3].a/w1450 ), .Z(
        \SUBBYTES[3].a/w1459 ) );
  AND U7807 ( .A(\SUBBYTES[3].a/w1466 ), .B(\SUBBYTES[3].a/w1473 ), .Z(
        \SUBBYTES[3].a/w1458 ) );
  AND U7808 ( .A(\SUBBYTES[3].a/w1406 ), .B(\SUBBYTES[3].a/w1402 ), .Z(
        \SUBBYTES[3].a/w1443 ) );
  AND U7809 ( .A(\SUBBYTES[3].a/w1407 ), .B(\SUBBYTES[3].a/w1403 ), .Z(
        \SUBBYTES[3].a/w1441 ) );
  ANDN U7810 ( .A(\SUBBYTES[3].a/w1533 ), .B(n2695), .Z(\SUBBYTES[3].a/w1440 )
         );
  XNOR U7811 ( .A(\w1[3][73] ), .B(\w1[3][79] ), .Z(n2695) );
  XOR U7812 ( .A(\w0[3][73] ), .B(g_input[457]), .Z(\w1[3][73] ) );
  AND U7813 ( .A(\w1[3][72] ), .B(\SUBBYTES[3].a/w1408 ), .Z(
        \SUBBYTES[3].a/w1436 ) );
  XOR U7814 ( .A(\w0[3][72] ), .B(g_input[456]), .Z(\w1[3][72] ) );
  AND U7815 ( .A(\SUBBYTES[3].a/w1409 ), .B(\SUBBYTES[3].a/w1405 ), .Z(
        \SUBBYTES[3].a/w1434 ) );
  AND U7816 ( .A(\SUBBYTES[3].a/w1494 ), .B(\SUBBYTES[3].a/w1526 ), .Z(
        \SUBBYTES[3].a/w1433 ) );
  ANDN U7817 ( .A(\SUBBYTES[3].a/w1515 ), .B(n2699), .Z(\SUBBYTES[3].a/w1428 )
         );
  XNOR U7818 ( .A(\w1[3][76] ), .B(\w1[3][79] ), .Z(n2699) );
  ANDN U7819 ( .A(\SUBBYTES[3].a/w1516 ), .B(n2700), .Z(\SUBBYTES[3].a/w1426 )
         );
  XNOR U7820 ( .A(\w1[3][74] ), .B(\w1[3][79] ), .Z(n2700) );
  XOR U7821 ( .A(\w0[3][79] ), .B(g_input[463]), .Z(\w1[3][79] ) );
  IV U7822 ( .A(n2702), .Z(\w1[3][74] ) );
  ANDN U7823 ( .A(\SUBBYTES[3].a/w1518 ), .B(n2701), .Z(\SUBBYTES[3].a/w1425 )
         );
  XOR U7824 ( .A(n2702), .B(\w1[3][76] ), .Z(n2701) );
  XOR U7825 ( .A(\w0[3][76] ), .B(g_input[460]), .Z(\w1[3][76] ) );
  XNOR U7826 ( .A(\w0[3][74] ), .B(g_input[458]), .Z(n2702) );
  AND U7827 ( .A(n2703), .B(\SUBBYTES[3].a/w1195 ), .Z(\SUBBYTES[3].a/w1330 )
         );
  AND U7828 ( .A(n2704), .B(\SUBBYTES[3].a/w1196 ), .Z(\SUBBYTES[3].a/w1328 )
         );
  AND U7829 ( .A(\SUBBYTES[3].a/w1326 ), .B(n2705), .Z(\SUBBYTES[3].a/w1327 )
         );
  ANDN U7830 ( .A(\w1[3][80] ), .B(n2706), .Z(\SUBBYTES[3].a/w1323 ) );
  AND U7831 ( .A(n2707), .B(\SUBBYTES[3].a/w1198 ), .Z(\SUBBYTES[3].a/w1321 )
         );
  AND U7832 ( .A(\SUBBYTES[3].a/w1319 ), .B(n2708), .Z(\SUBBYTES[3].a/w1320 )
         );
  XOR U7833 ( .A(\SUBBYTES[3].a/w1263 ), .B(n8402), .Z(n2708) );
  AND U7834 ( .A(\SUBBYTES[3].a/w1306 ), .B(\SUBBYTES[3].a/w1308 ), .Z(
        \SUBBYTES[3].a/w1315 ) );
  AND U7835 ( .A(\SUBBYTES[3].a/w1307 ), .B(\SUBBYTES[3].a/w1309 ), .Z(
        \SUBBYTES[3].a/w1313 ) );
  AND U7836 ( .A(\SUBBYTES[3].a/w1310 ), .B(\SUBBYTES[3].a/w1311 ), .Z(
        \SUBBYTES[3].a/w1312 ) );
  AND U7837 ( .A(\SUBBYTES[3].a/w1199 ), .B(n2703), .Z(\SUBBYTES[3].a/w1298 )
         );
  XOR U7838 ( .A(\SUBBYTES[3].a/w1267 ), .B(n994), .Z(n2703) );
  AND U7839 ( .A(\SUBBYTES[3].a/w1200 ), .B(n2704), .Z(\SUBBYTES[3].a/w1296 )
         );
  XOR U7840 ( .A(n8403), .B(\SUBBYTES[3].a/w1267 ), .Z(n2704) );
  ANDN U7841 ( .A(n2705), .B(n2709), .Z(\SUBBYTES[3].a/w1295 ) );
  XOR U7842 ( .A(n994), .B(n8403), .Z(n2705) );
  ANDN U7843 ( .A(\SUBBYTES[3].a/w1201 ), .B(n2706), .Z(\SUBBYTES[3].a/w1291 )
         );
  XNOR U7844 ( .A(\SUBBYTES[3].a/w1260 ), .B(\SUBBYTES[3].a/w1263 ), .Z(n2706)
         );
  AND U7845 ( .A(\SUBBYTES[3].a/w1202 ), .B(n2707), .Z(\SUBBYTES[3].a/w1289 )
         );
  XNOR U7846 ( .A(n2710), .B(\SUBBYTES[3].a/w1260 ), .Z(n2707) );
  AND U7847 ( .A(\SUBBYTES[3].a/w1287 ), .B(n2711), .Z(\SUBBYTES[3].a/w1288 )
         );
  XOR U7848 ( .A(n2712), .B(n2710), .Z(n2711) );
  IV U7849 ( .A(n8402), .Z(n2710) );
  ANDN U7850 ( .A(\SUBBYTES[3].a/w1306 ), .B(n2713), .Z(\SUBBYTES[3].a/w1283 )
         );
  ANDN U7851 ( .A(\SUBBYTES[3].a/w1307 ), .B(n2714), .Z(\SUBBYTES[3].a/w1281 )
         );
  ANDN U7852 ( .A(\SUBBYTES[3].a/w1310 ), .B(n2715), .Z(\SUBBYTES[3].a/w1280 )
         );
  AND U7853 ( .A(\SUBBYTES[3].a/w1266 ), .B(\SUBBYTES[3].a/w1265 ), .Z(
        \SUBBYTES[3].a/w1267 ) );
  IV U7854 ( .A(n2712), .Z(\SUBBYTES[3].a/w1263 ) );
  NAND U7855 ( .A(\SUBBYTES[3].a/w1242 ), .B(\SUBBYTES[3].a/w1257 ), .Z(n2712)
         );
  AND U7856 ( .A(\SUBBYTES[3].a/w1259 ), .B(\SUBBYTES[3].a/w1265 ), .Z(
        \SUBBYTES[3].a/w1260 ) );
  AND U7857 ( .A(\SUBBYTES[3].a/w1244 ), .B(\SUBBYTES[3].a/w1242 ), .Z(
        \SUBBYTES[3].a/w1254 ) );
  AND U7858 ( .A(\SUBBYTES[3].a/w1245 ), .B(\SUBBYTES[3].a/w1243 ), .Z(
        \SUBBYTES[3].a/w1252 ) );
  AND U7859 ( .A(\SUBBYTES[3].a/w1259 ), .B(\SUBBYTES[3].a/w1266 ), .Z(
        \SUBBYTES[3].a/w1251 ) );
  AND U7860 ( .A(\SUBBYTES[3].a/w1199 ), .B(\SUBBYTES[3].a/w1195 ), .Z(
        \SUBBYTES[3].a/w1236 ) );
  AND U7861 ( .A(\SUBBYTES[3].a/w1200 ), .B(\SUBBYTES[3].a/w1196 ), .Z(
        \SUBBYTES[3].a/w1234 ) );
  ANDN U7862 ( .A(\SUBBYTES[3].a/w1326 ), .B(n2709), .Z(\SUBBYTES[3].a/w1233 )
         );
  XNOR U7863 ( .A(\w1[3][81] ), .B(\w1[3][87] ), .Z(n2709) );
  XOR U7864 ( .A(\w0[3][81] ), .B(g_input[465]), .Z(\w1[3][81] ) );
  AND U7865 ( .A(\w1[3][80] ), .B(\SUBBYTES[3].a/w1201 ), .Z(
        \SUBBYTES[3].a/w1229 ) );
  XOR U7866 ( .A(\w0[3][80] ), .B(g_input[464]), .Z(\w1[3][80] ) );
  AND U7867 ( .A(\SUBBYTES[3].a/w1202 ), .B(\SUBBYTES[3].a/w1198 ), .Z(
        \SUBBYTES[3].a/w1227 ) );
  AND U7868 ( .A(\SUBBYTES[3].a/w1287 ), .B(\SUBBYTES[3].a/w1319 ), .Z(
        \SUBBYTES[3].a/w1226 ) );
  ANDN U7869 ( .A(\SUBBYTES[3].a/w1308 ), .B(n2713), .Z(\SUBBYTES[3].a/w1221 )
         );
  XNOR U7870 ( .A(\w1[3][84] ), .B(\w1[3][87] ), .Z(n2713) );
  ANDN U7871 ( .A(\SUBBYTES[3].a/w1309 ), .B(n2714), .Z(\SUBBYTES[3].a/w1219 )
         );
  XNOR U7872 ( .A(\w1[3][82] ), .B(\w1[3][87] ), .Z(n2714) );
  XOR U7873 ( .A(\w0[3][87] ), .B(g_input[471]), .Z(\w1[3][87] ) );
  IV U7874 ( .A(n2716), .Z(\w1[3][82] ) );
  ANDN U7875 ( .A(\SUBBYTES[3].a/w1311 ), .B(n2715), .Z(\SUBBYTES[3].a/w1218 )
         );
  XOR U7876 ( .A(n2716), .B(\w1[3][84] ), .Z(n2715) );
  XOR U7877 ( .A(\w0[3][84] ), .B(g_input[468]), .Z(\w1[3][84] ) );
  XNOR U7878 ( .A(\w0[3][82] ), .B(g_input[466]), .Z(n2716) );
  AND U7879 ( .A(n2717), .B(\SUBBYTES[3].a/w988 ), .Z(\SUBBYTES[3].a/w1123 )
         );
  AND U7880 ( .A(n2718), .B(\SUBBYTES[3].a/w989 ), .Z(\SUBBYTES[3].a/w1121 )
         );
  AND U7881 ( .A(\SUBBYTES[3].a/w1119 ), .B(n2719), .Z(\SUBBYTES[3].a/w1120 )
         );
  ANDN U7882 ( .A(\w1[3][88] ), .B(n2720), .Z(\SUBBYTES[3].a/w1116 ) );
  AND U7883 ( .A(n2721), .B(\SUBBYTES[3].a/w991 ), .Z(\SUBBYTES[3].a/w1114 )
         );
  AND U7884 ( .A(\SUBBYTES[3].a/w1112 ), .B(n2722), .Z(\SUBBYTES[3].a/w1113 )
         );
  XOR U7885 ( .A(\SUBBYTES[3].a/w1056 ), .B(n8400), .Z(n2722) );
  AND U7886 ( .A(\SUBBYTES[3].a/w1099 ), .B(\SUBBYTES[3].a/w1101 ), .Z(
        \SUBBYTES[3].a/w1108 ) );
  AND U7887 ( .A(\SUBBYTES[3].a/w1100 ), .B(\SUBBYTES[3].a/w1102 ), .Z(
        \SUBBYTES[3].a/w1106 ) );
  AND U7888 ( .A(\SUBBYTES[3].a/w1103 ), .B(\SUBBYTES[3].a/w1104 ), .Z(
        \SUBBYTES[3].a/w1105 ) );
  AND U7889 ( .A(\SUBBYTES[3].a/w992 ), .B(n2717), .Z(\SUBBYTES[3].a/w1091 )
         );
  XOR U7890 ( .A(\SUBBYTES[3].a/w1060 ), .B(n993), .Z(n2717) );
  AND U7891 ( .A(\SUBBYTES[3].a/w993 ), .B(n2718), .Z(\SUBBYTES[3].a/w1089 )
         );
  XOR U7892 ( .A(n8401), .B(\SUBBYTES[3].a/w1060 ), .Z(n2718) );
  ANDN U7893 ( .A(n2719), .B(n2723), .Z(\SUBBYTES[3].a/w1088 ) );
  XOR U7894 ( .A(n993), .B(n8401), .Z(n2719) );
  ANDN U7895 ( .A(\SUBBYTES[3].a/w994 ), .B(n2720), .Z(\SUBBYTES[3].a/w1084 )
         );
  XNOR U7896 ( .A(\SUBBYTES[3].a/w1053 ), .B(\SUBBYTES[3].a/w1056 ), .Z(n2720)
         );
  AND U7897 ( .A(\SUBBYTES[3].a/w995 ), .B(n2721), .Z(\SUBBYTES[3].a/w1082 )
         );
  XNOR U7898 ( .A(n2724), .B(\SUBBYTES[3].a/w1053 ), .Z(n2721) );
  AND U7899 ( .A(\SUBBYTES[3].a/w1080 ), .B(n2725), .Z(\SUBBYTES[3].a/w1081 )
         );
  XOR U7900 ( .A(n2726), .B(n2724), .Z(n2725) );
  IV U7901 ( .A(n8400), .Z(n2724) );
  ANDN U7902 ( .A(\SUBBYTES[3].a/w1099 ), .B(n2727), .Z(\SUBBYTES[3].a/w1076 )
         );
  ANDN U7903 ( .A(\SUBBYTES[3].a/w1100 ), .B(n2728), .Z(\SUBBYTES[3].a/w1074 )
         );
  ANDN U7904 ( .A(\SUBBYTES[3].a/w1103 ), .B(n2729), .Z(\SUBBYTES[3].a/w1073 )
         );
  AND U7905 ( .A(\SUBBYTES[3].a/w1059 ), .B(\SUBBYTES[3].a/w1058 ), .Z(
        \SUBBYTES[3].a/w1060 ) );
  IV U7906 ( .A(n2726), .Z(\SUBBYTES[3].a/w1056 ) );
  NAND U7907 ( .A(\SUBBYTES[3].a/w1035 ), .B(\SUBBYTES[3].a/w1050 ), .Z(n2726)
         );
  AND U7908 ( .A(\SUBBYTES[3].a/w1052 ), .B(\SUBBYTES[3].a/w1058 ), .Z(
        \SUBBYTES[3].a/w1053 ) );
  AND U7909 ( .A(\SUBBYTES[3].a/w1037 ), .B(\SUBBYTES[3].a/w1035 ), .Z(
        \SUBBYTES[3].a/w1047 ) );
  AND U7910 ( .A(\SUBBYTES[3].a/w1038 ), .B(\SUBBYTES[3].a/w1036 ), .Z(
        \SUBBYTES[3].a/w1045 ) );
  AND U7911 ( .A(\SUBBYTES[3].a/w1052 ), .B(\SUBBYTES[3].a/w1059 ), .Z(
        \SUBBYTES[3].a/w1044 ) );
  AND U7912 ( .A(\SUBBYTES[3].a/w992 ), .B(\SUBBYTES[3].a/w988 ), .Z(
        \SUBBYTES[3].a/w1029 ) );
  AND U7913 ( .A(\SUBBYTES[3].a/w993 ), .B(\SUBBYTES[3].a/w989 ), .Z(
        \SUBBYTES[3].a/w1027 ) );
  ANDN U7914 ( .A(\SUBBYTES[3].a/w1119 ), .B(n2723), .Z(\SUBBYTES[3].a/w1026 )
         );
  XNOR U7915 ( .A(\w1[3][89] ), .B(\w1[3][95] ), .Z(n2723) );
  XOR U7916 ( .A(\w0[3][89] ), .B(g_input[473]), .Z(\w1[3][89] ) );
  AND U7917 ( .A(\w1[3][88] ), .B(\SUBBYTES[3].a/w994 ), .Z(
        \SUBBYTES[3].a/w1022 ) );
  XOR U7918 ( .A(\w0[3][88] ), .B(g_input[472]), .Z(\w1[3][88] ) );
  AND U7919 ( .A(\SUBBYTES[3].a/w995 ), .B(\SUBBYTES[3].a/w991 ), .Z(
        \SUBBYTES[3].a/w1020 ) );
  AND U7920 ( .A(\SUBBYTES[3].a/w1080 ), .B(\SUBBYTES[3].a/w1112 ), .Z(
        \SUBBYTES[3].a/w1019 ) );
  ANDN U7921 ( .A(\SUBBYTES[3].a/w1101 ), .B(n2727), .Z(\SUBBYTES[3].a/w1014 )
         );
  XNOR U7922 ( .A(\w1[3][92] ), .B(\w1[3][95] ), .Z(n2727) );
  ANDN U7923 ( .A(\SUBBYTES[3].a/w1102 ), .B(n2728), .Z(\SUBBYTES[3].a/w1012 )
         );
  XNOR U7924 ( .A(\w1[3][90] ), .B(\w1[3][95] ), .Z(n2728) );
  XOR U7925 ( .A(\w0[3][95] ), .B(g_input[479]), .Z(\w1[3][95] ) );
  IV U7926 ( .A(n2730), .Z(\w1[3][90] ) );
  ANDN U7927 ( .A(\SUBBYTES[3].a/w1104 ), .B(n2729), .Z(\SUBBYTES[3].a/w1011 )
         );
  XOR U7928 ( .A(n2730), .B(\w1[3][92] ), .Z(n2729) );
  XOR U7929 ( .A(\w0[3][92] ), .B(g_input[476]), .Z(\w1[3][92] ) );
  XNOR U7930 ( .A(\w0[3][90] ), .B(g_input[474]), .Z(n2730) );
  AND U7931 ( .A(\SUBBYTES[3].a/w2084 ), .B(\SUBBYTES[3].a/w2071 ), .Z(n8410)
         );
  AND U7932 ( .A(\SUBBYTES[3].a/w1877 ), .B(\SUBBYTES[3].a/w1866 ), .Z(n8409)
         );
  AND U7933 ( .A(\SUBBYTES[3].a/w221 ), .B(\SUBBYTES[3].a/w208 ), .Z(n8392) );
  AND U7934 ( .A(\SUBBYTES[3].a/w1877 ), .B(\SUBBYTES[3].a/w1864 ), .Z(n8408)
         );
  AND U7935 ( .A(\SUBBYTES[3].a/w1670 ), .B(\SUBBYTES[3].a/w1659 ), .Z(n8407)
         );
  AND U7936 ( .A(\SUBBYTES[3].a/w1670 ), .B(\SUBBYTES[3].a/w1657 ), .Z(n8406)
         );
  AND U7937 ( .A(\SUBBYTES[3].a/w1463 ), .B(\SUBBYTES[3].a/w1452 ), .Z(n8405)
         );
  AND U7938 ( .A(\SUBBYTES[3].a/w1463 ), .B(\SUBBYTES[3].a/w1450 ), .Z(n8404)
         );
  AND U7939 ( .A(\SUBBYTES[3].a/w1256 ), .B(\SUBBYTES[3].a/w1245 ), .Z(n8403)
         );
  AND U7940 ( .A(\SUBBYTES[3].a/w1256 ), .B(\SUBBYTES[3].a/w1243 ), .Z(n8402)
         );
  AND U7941 ( .A(\SUBBYTES[3].a/w1049 ), .B(\SUBBYTES[3].a/w1038 ), .Z(n8401)
         );
  AND U7942 ( .A(\SUBBYTES[3].a/w1049 ), .B(\SUBBYTES[3].a/w1036 ), .Z(n8400)
         );
  AND U7943 ( .A(\SUBBYTES[3].a/w842 ), .B(\SUBBYTES[3].a/w831 ), .Z(n8399) );
  AND U7944 ( .A(\SUBBYTES[3].a/w842 ), .B(\SUBBYTES[3].a/w829 ), .Z(n8398) );
  AND U7945 ( .A(\SUBBYTES[3].a/w635 ), .B(\SUBBYTES[3].a/w624 ), .Z(n8397) );
  AND U7946 ( .A(\SUBBYTES[3].a/w635 ), .B(\SUBBYTES[3].a/w622 ), .Z(n8396) );
  AND U7947 ( .A(\SUBBYTES[3].a/w428 ), .B(\SUBBYTES[3].a/w417 ), .Z(n8395) );
  AND U7948 ( .A(\SUBBYTES[3].a/w428 ), .B(\SUBBYTES[3].a/w415 ), .Z(n8394) );
  AND U7949 ( .A(\SUBBYTES[3].a/w3326 ), .B(\SUBBYTES[3].a/w3315 ), .Z(n8423)
         );
  AND U7950 ( .A(\SUBBYTES[3].a/w3326 ), .B(\SUBBYTES[3].a/w3313 ), .Z(n8422)
         );
  AND U7951 ( .A(\SUBBYTES[3].a/w3119 ), .B(\SUBBYTES[3].a/w3108 ), .Z(n8421)
         );
  AND U7952 ( .A(\SUBBYTES[3].a/w3119 ), .B(\SUBBYTES[3].a/w3106 ), .Z(n8420)
         );
  AND U7953 ( .A(\SUBBYTES[3].a/w2912 ), .B(\SUBBYTES[3].a/w2901 ), .Z(n8419)
         );
  AND U7954 ( .A(\SUBBYTES[3].a/w2912 ), .B(\SUBBYTES[3].a/w2899 ), .Z(n8418)
         );
  AND U7955 ( .A(\SUBBYTES[3].a/w2705 ), .B(\SUBBYTES[3].a/w2694 ), .Z(n8417)
         );
  AND U7956 ( .A(\SUBBYTES[3].a/w2705 ), .B(\SUBBYTES[3].a/w2692 ), .Z(n8416)
         );
  AND U7957 ( .A(\SUBBYTES[3].a/w2498 ), .B(\SUBBYTES[3].a/w2487 ), .Z(n8415)
         );
  AND U7958 ( .A(\SUBBYTES[3].a/w2498 ), .B(\SUBBYTES[3].a/w2485 ), .Z(n8414)
         );
  AND U7959 ( .A(\SUBBYTES[3].a/w2291 ), .B(\SUBBYTES[3].a/w2280 ), .Z(n8413)
         );
  AND U7960 ( .A(\SUBBYTES[3].a/w2291 ), .B(\SUBBYTES[3].a/w2278 ), .Z(n8412)
         );
  AND U7961 ( .A(\SUBBYTES[3].a/w2084 ), .B(\SUBBYTES[3].a/w2073 ), .Z(n8411)
         );
  AND U7962 ( .A(\SUBBYTES[3].a/w221 ), .B(\SUBBYTES[3].a/w210 ), .Z(n8393) );
  AND U7963 ( .A(n2731), .B(\SUBBYTES[2].a/w781 ), .Z(\SUBBYTES[2].a/w916 ) );
  AND U7964 ( .A(n2732), .B(\SUBBYTES[2].a/w782 ), .Z(\SUBBYTES[2].a/w914 ) );
  AND U7965 ( .A(\SUBBYTES[2].a/w912 ), .B(n2733), .Z(\SUBBYTES[2].a/w913 ) );
  ANDN U7966 ( .A(\w1[2][96] ), .B(n2734), .Z(\SUBBYTES[2].a/w909 ) );
  AND U7967 ( .A(n2735), .B(\SUBBYTES[2].a/w784 ), .Z(\SUBBYTES[2].a/w907 ) );
  AND U7968 ( .A(\SUBBYTES[2].a/w905 ), .B(n2736), .Z(\SUBBYTES[2].a/w906 ) );
  XOR U7969 ( .A(\SUBBYTES[2].a/w849 ), .B(n7118), .Z(n2736) );
  AND U7970 ( .A(\SUBBYTES[2].a/w892 ), .B(\SUBBYTES[2].a/w894 ), .Z(
        \SUBBYTES[2].a/w901 ) );
  AND U7971 ( .A(\SUBBYTES[2].a/w893 ), .B(\SUBBYTES[2].a/w895 ), .Z(
        \SUBBYTES[2].a/w899 ) );
  AND U7972 ( .A(\SUBBYTES[2].a/w896 ), .B(\SUBBYTES[2].a/w897 ), .Z(
        \SUBBYTES[2].a/w898 ) );
  AND U7973 ( .A(\SUBBYTES[2].a/w785 ), .B(n2731), .Z(\SUBBYTES[2].a/w884 ) );
  XOR U7974 ( .A(\SUBBYTES[2].a/w853 ), .B(n976), .Z(n2731) );
  AND U7975 ( .A(\SUBBYTES[2].a/w786 ), .B(n2732), .Z(\SUBBYTES[2].a/w882 ) );
  XOR U7976 ( .A(n7119), .B(\SUBBYTES[2].a/w853 ), .Z(n2732) );
  ANDN U7977 ( .A(n2733), .B(n2737), .Z(\SUBBYTES[2].a/w881 ) );
  XOR U7978 ( .A(n976), .B(n7119), .Z(n2733) );
  ANDN U7979 ( .A(\SUBBYTES[2].a/w787 ), .B(n2734), .Z(\SUBBYTES[2].a/w877 )
         );
  XNOR U7980 ( .A(\SUBBYTES[2].a/w846 ), .B(\SUBBYTES[2].a/w849 ), .Z(n2734)
         );
  AND U7981 ( .A(\SUBBYTES[2].a/w788 ), .B(n2735), .Z(\SUBBYTES[2].a/w875 ) );
  XNOR U7982 ( .A(n2738), .B(\SUBBYTES[2].a/w846 ), .Z(n2735) );
  AND U7983 ( .A(\SUBBYTES[2].a/w873 ), .B(n2739), .Z(\SUBBYTES[2].a/w874 ) );
  XOR U7984 ( .A(n2740), .B(n2738), .Z(n2739) );
  IV U7985 ( .A(n7118), .Z(n2738) );
  ANDN U7986 ( .A(\SUBBYTES[2].a/w892 ), .B(n2741), .Z(\SUBBYTES[2].a/w869 )
         );
  ANDN U7987 ( .A(\SUBBYTES[2].a/w893 ), .B(n2742), .Z(\SUBBYTES[2].a/w867 )
         );
  ANDN U7988 ( .A(\SUBBYTES[2].a/w896 ), .B(n2743), .Z(\SUBBYTES[2].a/w866 )
         );
  AND U7989 ( .A(\SUBBYTES[2].a/w852 ), .B(\SUBBYTES[2].a/w851 ), .Z(
        \SUBBYTES[2].a/w853 ) );
  IV U7990 ( .A(n2740), .Z(\SUBBYTES[2].a/w849 ) );
  NAND U7991 ( .A(\SUBBYTES[2].a/w828 ), .B(\SUBBYTES[2].a/w843 ), .Z(n2740)
         );
  AND U7992 ( .A(\SUBBYTES[2].a/w845 ), .B(\SUBBYTES[2].a/w851 ), .Z(
        \SUBBYTES[2].a/w846 ) );
  AND U7993 ( .A(\SUBBYTES[2].a/w830 ), .B(\SUBBYTES[2].a/w828 ), .Z(
        \SUBBYTES[2].a/w840 ) );
  AND U7994 ( .A(\SUBBYTES[2].a/w831 ), .B(\SUBBYTES[2].a/w829 ), .Z(
        \SUBBYTES[2].a/w838 ) );
  AND U7995 ( .A(\SUBBYTES[2].a/w845 ), .B(\SUBBYTES[2].a/w852 ), .Z(
        \SUBBYTES[2].a/w837 ) );
  AND U7996 ( .A(\SUBBYTES[2].a/w785 ), .B(\SUBBYTES[2].a/w781 ), .Z(
        \SUBBYTES[2].a/w822 ) );
  AND U7997 ( .A(\SUBBYTES[2].a/w786 ), .B(\SUBBYTES[2].a/w782 ), .Z(
        \SUBBYTES[2].a/w820 ) );
  ANDN U7998 ( .A(\SUBBYTES[2].a/w912 ), .B(n2737), .Z(\SUBBYTES[2].a/w819 )
         );
  XNOR U7999 ( .A(\w1[2][103] ), .B(\w1[2][97] ), .Z(n2737) );
  XOR U8000 ( .A(\w0[2][97] ), .B(g_input[353]), .Z(\w1[2][97] ) );
  IV U8001 ( .A(n2744), .Z(\w1[2][103] ) );
  AND U8002 ( .A(\w1[2][96] ), .B(\SUBBYTES[2].a/w787 ), .Z(
        \SUBBYTES[2].a/w815 ) );
  XOR U8003 ( .A(\w0[2][96] ), .B(g_input[352]), .Z(\w1[2][96] ) );
  AND U8004 ( .A(\SUBBYTES[2].a/w788 ), .B(\SUBBYTES[2].a/w784 ), .Z(
        \SUBBYTES[2].a/w813 ) );
  AND U8005 ( .A(\SUBBYTES[2].a/w873 ), .B(\SUBBYTES[2].a/w905 ), .Z(
        \SUBBYTES[2].a/w812 ) );
  ANDN U8006 ( .A(\SUBBYTES[2].a/w894 ), .B(n2741), .Z(\SUBBYTES[2].a/w807 )
         );
  XOR U8007 ( .A(\w1[2][100] ), .B(n2744), .Z(n2741) );
  ANDN U8008 ( .A(\SUBBYTES[2].a/w895 ), .B(n2742), .Z(\SUBBYTES[2].a/w805 )
         );
  XOR U8009 ( .A(n2744), .B(\w1[2][98] ), .Z(n2742) );
  XNOR U8010 ( .A(\w0[2][103] ), .B(g_input[359]), .Z(n2744) );
  ANDN U8011 ( .A(\SUBBYTES[2].a/w897 ), .B(n2743), .Z(\SUBBYTES[2].a/w804 )
         );
  XNOR U8012 ( .A(\w1[2][100] ), .B(\w1[2][98] ), .Z(n2743) );
  XOR U8013 ( .A(\w0[2][98] ), .B(g_input[354]), .Z(\w1[2][98] ) );
  XOR U8014 ( .A(\w0[2][100] ), .B(g_input[356]), .Z(\w1[2][100] ) );
  AND U8015 ( .A(n2745), .B(\SUBBYTES[2].a/w574 ), .Z(\SUBBYTES[2].a/w709 ) );
  AND U8016 ( .A(n2746), .B(\SUBBYTES[2].a/w575 ), .Z(\SUBBYTES[2].a/w707 ) );
  AND U8017 ( .A(\SUBBYTES[2].a/w705 ), .B(n2747), .Z(\SUBBYTES[2].a/w706 ) );
  ANDN U8018 ( .A(\w1[2][104] ), .B(n2748), .Z(\SUBBYTES[2].a/w702 ) );
  AND U8019 ( .A(n2749), .B(\SUBBYTES[2].a/w577 ), .Z(\SUBBYTES[2].a/w700 ) );
  AND U8020 ( .A(\SUBBYTES[2].a/w698 ), .B(n2750), .Z(\SUBBYTES[2].a/w699 ) );
  XOR U8021 ( .A(\SUBBYTES[2].a/w642 ), .B(n7116), .Z(n2750) );
  AND U8022 ( .A(\SUBBYTES[2].a/w685 ), .B(\SUBBYTES[2].a/w687 ), .Z(
        \SUBBYTES[2].a/w694 ) );
  AND U8023 ( .A(\SUBBYTES[2].a/w686 ), .B(\SUBBYTES[2].a/w688 ), .Z(
        \SUBBYTES[2].a/w692 ) );
  AND U8024 ( .A(\SUBBYTES[2].a/w689 ), .B(\SUBBYTES[2].a/w690 ), .Z(
        \SUBBYTES[2].a/w691 ) );
  AND U8025 ( .A(\SUBBYTES[2].a/w578 ), .B(n2745), .Z(\SUBBYTES[2].a/w677 ) );
  XOR U8026 ( .A(\SUBBYTES[2].a/w646 ), .B(n975), .Z(n2745) );
  AND U8027 ( .A(\SUBBYTES[2].a/w579 ), .B(n2746), .Z(\SUBBYTES[2].a/w675 ) );
  XOR U8028 ( .A(n7117), .B(\SUBBYTES[2].a/w646 ), .Z(n2746) );
  ANDN U8029 ( .A(n2747), .B(n2751), .Z(\SUBBYTES[2].a/w674 ) );
  XOR U8030 ( .A(n975), .B(n7117), .Z(n2747) );
  ANDN U8031 ( .A(\SUBBYTES[2].a/w580 ), .B(n2748), .Z(\SUBBYTES[2].a/w670 )
         );
  XNOR U8032 ( .A(\SUBBYTES[2].a/w639 ), .B(\SUBBYTES[2].a/w642 ), .Z(n2748)
         );
  AND U8033 ( .A(\SUBBYTES[2].a/w581 ), .B(n2749), .Z(\SUBBYTES[2].a/w668 ) );
  XNOR U8034 ( .A(n2752), .B(\SUBBYTES[2].a/w639 ), .Z(n2749) );
  AND U8035 ( .A(\SUBBYTES[2].a/w666 ), .B(n2753), .Z(\SUBBYTES[2].a/w667 ) );
  XOR U8036 ( .A(n2754), .B(n2752), .Z(n2753) );
  IV U8037 ( .A(n7116), .Z(n2752) );
  ANDN U8038 ( .A(\SUBBYTES[2].a/w685 ), .B(n2755), .Z(\SUBBYTES[2].a/w662 )
         );
  ANDN U8039 ( .A(\SUBBYTES[2].a/w686 ), .B(n2756), .Z(\SUBBYTES[2].a/w660 )
         );
  ANDN U8040 ( .A(\SUBBYTES[2].a/w689 ), .B(n2757), .Z(\SUBBYTES[2].a/w659 )
         );
  AND U8041 ( .A(\SUBBYTES[2].a/w645 ), .B(\SUBBYTES[2].a/w644 ), .Z(
        \SUBBYTES[2].a/w646 ) );
  IV U8042 ( .A(n2754), .Z(\SUBBYTES[2].a/w642 ) );
  NAND U8043 ( .A(\SUBBYTES[2].a/w621 ), .B(\SUBBYTES[2].a/w636 ), .Z(n2754)
         );
  AND U8044 ( .A(\SUBBYTES[2].a/w638 ), .B(\SUBBYTES[2].a/w644 ), .Z(
        \SUBBYTES[2].a/w639 ) );
  AND U8045 ( .A(\SUBBYTES[2].a/w623 ), .B(\SUBBYTES[2].a/w621 ), .Z(
        \SUBBYTES[2].a/w633 ) );
  AND U8046 ( .A(\SUBBYTES[2].a/w624 ), .B(\SUBBYTES[2].a/w622 ), .Z(
        \SUBBYTES[2].a/w631 ) );
  AND U8047 ( .A(\SUBBYTES[2].a/w638 ), .B(\SUBBYTES[2].a/w645 ), .Z(
        \SUBBYTES[2].a/w630 ) );
  AND U8048 ( .A(\SUBBYTES[2].a/w578 ), .B(\SUBBYTES[2].a/w574 ), .Z(
        \SUBBYTES[2].a/w615 ) );
  AND U8049 ( .A(\SUBBYTES[2].a/w579 ), .B(\SUBBYTES[2].a/w575 ), .Z(
        \SUBBYTES[2].a/w613 ) );
  ANDN U8050 ( .A(\SUBBYTES[2].a/w705 ), .B(n2751), .Z(\SUBBYTES[2].a/w612 )
         );
  XNOR U8051 ( .A(\w1[2][105] ), .B(\w1[2][111] ), .Z(n2751) );
  XOR U8052 ( .A(\w0[2][105] ), .B(g_input[361]), .Z(\w1[2][105] ) );
  AND U8053 ( .A(\w1[2][104] ), .B(\SUBBYTES[2].a/w580 ), .Z(
        \SUBBYTES[2].a/w608 ) );
  XOR U8054 ( .A(\w0[2][104] ), .B(g_input[360]), .Z(\w1[2][104] ) );
  AND U8055 ( .A(\SUBBYTES[2].a/w581 ), .B(\SUBBYTES[2].a/w577 ), .Z(
        \SUBBYTES[2].a/w606 ) );
  AND U8056 ( .A(\SUBBYTES[2].a/w666 ), .B(\SUBBYTES[2].a/w698 ), .Z(
        \SUBBYTES[2].a/w605 ) );
  ANDN U8057 ( .A(\SUBBYTES[2].a/w687 ), .B(n2755), .Z(\SUBBYTES[2].a/w600 )
         );
  XNOR U8058 ( .A(\w1[2][108] ), .B(\w1[2][111] ), .Z(n2755) );
  ANDN U8059 ( .A(\SUBBYTES[2].a/w688 ), .B(n2756), .Z(\SUBBYTES[2].a/w598 )
         );
  XNOR U8060 ( .A(\w1[2][106] ), .B(\w1[2][111] ), .Z(n2756) );
  XOR U8061 ( .A(\w0[2][111] ), .B(g_input[367]), .Z(\w1[2][111] ) );
  IV U8062 ( .A(n2758), .Z(\w1[2][106] ) );
  ANDN U8063 ( .A(\SUBBYTES[2].a/w690 ), .B(n2757), .Z(\SUBBYTES[2].a/w597 )
         );
  XOR U8064 ( .A(n2758), .B(\w1[2][108] ), .Z(n2757) );
  XOR U8065 ( .A(\w0[2][108] ), .B(g_input[364]), .Z(\w1[2][108] ) );
  XNOR U8066 ( .A(\w0[2][106] ), .B(g_input[362]), .Z(n2758) );
  AND U8067 ( .A(n2759), .B(\SUBBYTES[2].a/w367 ), .Z(\SUBBYTES[2].a/w502 ) );
  AND U8068 ( .A(n2760), .B(\SUBBYTES[2].a/w368 ), .Z(\SUBBYTES[2].a/w500 ) );
  AND U8069 ( .A(\SUBBYTES[2].a/w498 ), .B(n2761), .Z(\SUBBYTES[2].a/w499 ) );
  ANDN U8070 ( .A(\w1[2][112] ), .B(n2762), .Z(\SUBBYTES[2].a/w495 ) );
  AND U8071 ( .A(n2763), .B(\SUBBYTES[2].a/w370 ), .Z(\SUBBYTES[2].a/w493 ) );
  AND U8072 ( .A(\SUBBYTES[2].a/w491 ), .B(n2764), .Z(\SUBBYTES[2].a/w492 ) );
  XOR U8073 ( .A(\SUBBYTES[2].a/w435 ), .B(n7114), .Z(n2764) );
  AND U8074 ( .A(\SUBBYTES[2].a/w478 ), .B(\SUBBYTES[2].a/w480 ), .Z(
        \SUBBYTES[2].a/w487 ) );
  AND U8075 ( .A(\SUBBYTES[2].a/w479 ), .B(\SUBBYTES[2].a/w481 ), .Z(
        \SUBBYTES[2].a/w485 ) );
  AND U8076 ( .A(\SUBBYTES[2].a/w482 ), .B(\SUBBYTES[2].a/w483 ), .Z(
        \SUBBYTES[2].a/w484 ) );
  AND U8077 ( .A(\SUBBYTES[2].a/w371 ), .B(n2759), .Z(\SUBBYTES[2].a/w470 ) );
  XOR U8078 ( .A(\SUBBYTES[2].a/w439 ), .B(n974), .Z(n2759) );
  AND U8079 ( .A(\SUBBYTES[2].a/w372 ), .B(n2760), .Z(\SUBBYTES[2].a/w468 ) );
  XOR U8080 ( .A(n7115), .B(\SUBBYTES[2].a/w439 ), .Z(n2760) );
  ANDN U8081 ( .A(n2761), .B(n2765), .Z(\SUBBYTES[2].a/w467 ) );
  XOR U8082 ( .A(n974), .B(n7115), .Z(n2761) );
  ANDN U8083 ( .A(\SUBBYTES[2].a/w373 ), .B(n2762), .Z(\SUBBYTES[2].a/w463 )
         );
  XNOR U8084 ( .A(\SUBBYTES[2].a/w432 ), .B(\SUBBYTES[2].a/w435 ), .Z(n2762)
         );
  AND U8085 ( .A(\SUBBYTES[2].a/w374 ), .B(n2763), .Z(\SUBBYTES[2].a/w461 ) );
  XNOR U8086 ( .A(n2766), .B(\SUBBYTES[2].a/w432 ), .Z(n2763) );
  AND U8087 ( .A(\SUBBYTES[2].a/w459 ), .B(n2767), .Z(\SUBBYTES[2].a/w460 ) );
  XOR U8088 ( .A(n2768), .B(n2766), .Z(n2767) );
  IV U8089 ( .A(n7114), .Z(n2766) );
  ANDN U8090 ( .A(\SUBBYTES[2].a/w478 ), .B(n2769), .Z(\SUBBYTES[2].a/w455 )
         );
  ANDN U8091 ( .A(\SUBBYTES[2].a/w479 ), .B(n2770), .Z(\SUBBYTES[2].a/w453 )
         );
  ANDN U8092 ( .A(\SUBBYTES[2].a/w482 ), .B(n2771), .Z(\SUBBYTES[2].a/w452 )
         );
  AND U8093 ( .A(\SUBBYTES[2].a/w438 ), .B(\SUBBYTES[2].a/w437 ), .Z(
        \SUBBYTES[2].a/w439 ) );
  IV U8094 ( .A(n2768), .Z(\SUBBYTES[2].a/w435 ) );
  NAND U8095 ( .A(\SUBBYTES[2].a/w414 ), .B(\SUBBYTES[2].a/w429 ), .Z(n2768)
         );
  AND U8096 ( .A(\SUBBYTES[2].a/w431 ), .B(\SUBBYTES[2].a/w437 ), .Z(
        \SUBBYTES[2].a/w432 ) );
  AND U8097 ( .A(\SUBBYTES[2].a/w416 ), .B(\SUBBYTES[2].a/w414 ), .Z(
        \SUBBYTES[2].a/w426 ) );
  AND U8098 ( .A(\SUBBYTES[2].a/w417 ), .B(\SUBBYTES[2].a/w415 ), .Z(
        \SUBBYTES[2].a/w424 ) );
  AND U8099 ( .A(\SUBBYTES[2].a/w431 ), .B(\SUBBYTES[2].a/w438 ), .Z(
        \SUBBYTES[2].a/w423 ) );
  AND U8100 ( .A(\SUBBYTES[2].a/w371 ), .B(\SUBBYTES[2].a/w367 ), .Z(
        \SUBBYTES[2].a/w408 ) );
  AND U8101 ( .A(\SUBBYTES[2].a/w372 ), .B(\SUBBYTES[2].a/w368 ), .Z(
        \SUBBYTES[2].a/w406 ) );
  ANDN U8102 ( .A(\SUBBYTES[2].a/w498 ), .B(n2765), .Z(\SUBBYTES[2].a/w405 )
         );
  XNOR U8103 ( .A(\w1[2][113] ), .B(\w1[2][119] ), .Z(n2765) );
  XOR U8104 ( .A(\w0[2][113] ), .B(g_input[369]), .Z(\w1[2][113] ) );
  AND U8105 ( .A(\w1[2][112] ), .B(\SUBBYTES[2].a/w373 ), .Z(
        \SUBBYTES[2].a/w401 ) );
  XOR U8106 ( .A(\w0[2][112] ), .B(g_input[368]), .Z(\w1[2][112] ) );
  AND U8107 ( .A(\SUBBYTES[2].a/w374 ), .B(\SUBBYTES[2].a/w370 ), .Z(
        \SUBBYTES[2].a/w399 ) );
  AND U8108 ( .A(\SUBBYTES[2].a/w459 ), .B(\SUBBYTES[2].a/w491 ), .Z(
        \SUBBYTES[2].a/w398 ) );
  ANDN U8109 ( .A(\SUBBYTES[2].a/w480 ), .B(n2769), .Z(\SUBBYTES[2].a/w393 )
         );
  XNOR U8110 ( .A(\w1[2][116] ), .B(\w1[2][119] ), .Z(n2769) );
  ANDN U8111 ( .A(\SUBBYTES[2].a/w481 ), .B(n2770), .Z(\SUBBYTES[2].a/w391 )
         );
  XNOR U8112 ( .A(\w1[2][114] ), .B(\w1[2][119] ), .Z(n2770) );
  XOR U8113 ( .A(\w0[2][119] ), .B(g_input[375]), .Z(\w1[2][119] ) );
  IV U8114 ( .A(n2772), .Z(\w1[2][114] ) );
  ANDN U8115 ( .A(\SUBBYTES[2].a/w483 ), .B(n2771), .Z(\SUBBYTES[2].a/w390 )
         );
  XOR U8116 ( .A(n2772), .B(\w1[2][116] ), .Z(n2771) );
  XOR U8117 ( .A(\w0[2][116] ), .B(g_input[372]), .Z(\w1[2][116] ) );
  XNOR U8118 ( .A(\w0[2][114] ), .B(g_input[370]), .Z(n2772) );
  AND U8119 ( .A(n2773), .B(\SUBBYTES[2].a/w3265 ), .Z(\SUBBYTES[2].a/w3400 )
         );
  AND U8120 ( .A(n2774), .B(\SUBBYTES[2].a/w3266 ), .Z(\SUBBYTES[2].a/w3398 )
         );
  AND U8121 ( .A(\SUBBYTES[2].a/w3396 ), .B(n2775), .Z(\SUBBYTES[2].a/w3397 )
         );
  ANDN U8122 ( .A(\w1[2][0] ), .B(n2776), .Z(\SUBBYTES[2].a/w3393 ) );
  AND U8123 ( .A(n2777), .B(\SUBBYTES[2].a/w3268 ), .Z(\SUBBYTES[2].a/w3391 )
         );
  AND U8124 ( .A(\SUBBYTES[2].a/w3389 ), .B(n2778), .Z(\SUBBYTES[2].a/w3390 )
         );
  XOR U8125 ( .A(\SUBBYTES[2].a/w3333 ), .B(n7142), .Z(n2778) );
  AND U8126 ( .A(\SUBBYTES[2].a/w3376 ), .B(\SUBBYTES[2].a/w3378 ), .Z(
        \SUBBYTES[2].a/w3385 ) );
  AND U8127 ( .A(\SUBBYTES[2].a/w3377 ), .B(\SUBBYTES[2].a/w3379 ), .Z(
        \SUBBYTES[2].a/w3383 ) );
  AND U8128 ( .A(\SUBBYTES[2].a/w3380 ), .B(\SUBBYTES[2].a/w3381 ), .Z(
        \SUBBYTES[2].a/w3382 ) );
  AND U8129 ( .A(\SUBBYTES[2].a/w3269 ), .B(n2773), .Z(\SUBBYTES[2].a/w3368 )
         );
  XOR U8130 ( .A(\SUBBYTES[2].a/w3337 ), .B(n988), .Z(n2773) );
  AND U8131 ( .A(\SUBBYTES[2].a/w3270 ), .B(n2774), .Z(\SUBBYTES[2].a/w3366 )
         );
  XOR U8132 ( .A(n7143), .B(\SUBBYTES[2].a/w3337 ), .Z(n2774) );
  ANDN U8133 ( .A(n2775), .B(n2779), .Z(\SUBBYTES[2].a/w3365 ) );
  XOR U8134 ( .A(n988), .B(n7143), .Z(n2775) );
  ANDN U8135 ( .A(\SUBBYTES[2].a/w3271 ), .B(n2776), .Z(\SUBBYTES[2].a/w3361 )
         );
  XNOR U8136 ( .A(\SUBBYTES[2].a/w3330 ), .B(\SUBBYTES[2].a/w3333 ), .Z(n2776)
         );
  AND U8137 ( .A(\SUBBYTES[2].a/w3272 ), .B(n2777), .Z(\SUBBYTES[2].a/w3359 )
         );
  XNOR U8138 ( .A(n2780), .B(\SUBBYTES[2].a/w3330 ), .Z(n2777) );
  AND U8139 ( .A(\SUBBYTES[2].a/w3357 ), .B(n2781), .Z(\SUBBYTES[2].a/w3358 )
         );
  XOR U8140 ( .A(n2782), .B(n2780), .Z(n2781) );
  IV U8141 ( .A(n7142), .Z(n2780) );
  ANDN U8142 ( .A(\SUBBYTES[2].a/w3376 ), .B(n2783), .Z(\SUBBYTES[2].a/w3353 )
         );
  ANDN U8143 ( .A(\SUBBYTES[2].a/w3377 ), .B(n2784), .Z(\SUBBYTES[2].a/w3351 )
         );
  ANDN U8144 ( .A(\SUBBYTES[2].a/w3380 ), .B(n2785), .Z(\SUBBYTES[2].a/w3350 )
         );
  AND U8145 ( .A(\SUBBYTES[2].a/w3336 ), .B(\SUBBYTES[2].a/w3335 ), .Z(
        \SUBBYTES[2].a/w3337 ) );
  IV U8146 ( .A(n2782), .Z(\SUBBYTES[2].a/w3333 ) );
  NAND U8147 ( .A(\SUBBYTES[2].a/w3312 ), .B(\SUBBYTES[2].a/w3327 ), .Z(n2782)
         );
  AND U8148 ( .A(\SUBBYTES[2].a/w3329 ), .B(\SUBBYTES[2].a/w3335 ), .Z(
        \SUBBYTES[2].a/w3330 ) );
  AND U8149 ( .A(\SUBBYTES[2].a/w3314 ), .B(\SUBBYTES[2].a/w3312 ), .Z(
        \SUBBYTES[2].a/w3324 ) );
  AND U8150 ( .A(\SUBBYTES[2].a/w3315 ), .B(\SUBBYTES[2].a/w3313 ), .Z(
        \SUBBYTES[2].a/w3322 ) );
  AND U8151 ( .A(\SUBBYTES[2].a/w3329 ), .B(\SUBBYTES[2].a/w3336 ), .Z(
        \SUBBYTES[2].a/w3321 ) );
  AND U8152 ( .A(\SUBBYTES[2].a/w3269 ), .B(\SUBBYTES[2].a/w3265 ), .Z(
        \SUBBYTES[2].a/w3306 ) );
  AND U8153 ( .A(\SUBBYTES[2].a/w3270 ), .B(\SUBBYTES[2].a/w3266 ), .Z(
        \SUBBYTES[2].a/w3304 ) );
  ANDN U8154 ( .A(\SUBBYTES[2].a/w3396 ), .B(n2779), .Z(\SUBBYTES[2].a/w3303 )
         );
  XNOR U8155 ( .A(\w1[2][1] ), .B(\w1[2][7] ), .Z(n2779) );
  XOR U8156 ( .A(\w0[2][1] ), .B(g_input[257]), .Z(\w1[2][1] ) );
  AND U8157 ( .A(\w1[2][0] ), .B(\SUBBYTES[2].a/w3271 ), .Z(
        \SUBBYTES[2].a/w3299 ) );
  XOR U8158 ( .A(\w0[2][0] ), .B(g_input[256]), .Z(\w1[2][0] ) );
  AND U8159 ( .A(\SUBBYTES[2].a/w3272 ), .B(\SUBBYTES[2].a/w3268 ), .Z(
        \SUBBYTES[2].a/w3297 ) );
  AND U8160 ( .A(\SUBBYTES[2].a/w3357 ), .B(\SUBBYTES[2].a/w3389 ), .Z(
        \SUBBYTES[2].a/w3296 ) );
  ANDN U8161 ( .A(\SUBBYTES[2].a/w3378 ), .B(n2783), .Z(\SUBBYTES[2].a/w3291 )
         );
  XNOR U8162 ( .A(\w1[2][4] ), .B(\w1[2][7] ), .Z(n2783) );
  ANDN U8163 ( .A(\SUBBYTES[2].a/w3379 ), .B(n2784), .Z(\SUBBYTES[2].a/w3289 )
         );
  XNOR U8164 ( .A(\w1[2][2] ), .B(\w1[2][7] ), .Z(n2784) );
  XOR U8165 ( .A(\w0[2][7] ), .B(g_input[263]), .Z(\w1[2][7] ) );
  IV U8166 ( .A(n2786), .Z(\w1[2][2] ) );
  ANDN U8167 ( .A(\SUBBYTES[2].a/w3381 ), .B(n2785), .Z(\SUBBYTES[2].a/w3288 )
         );
  XOR U8168 ( .A(n2786), .B(\w1[2][4] ), .Z(n2785) );
  XOR U8169 ( .A(\w0[2][4] ), .B(g_input[260]), .Z(\w1[2][4] ) );
  XNOR U8170 ( .A(\w0[2][2] ), .B(g_input[258]), .Z(n2786) );
  AND U8171 ( .A(n2787), .B(\SUBBYTES[2].a/w3058 ), .Z(\SUBBYTES[2].a/w3193 )
         );
  AND U8172 ( .A(n2788), .B(\SUBBYTES[2].a/w3059 ), .Z(\SUBBYTES[2].a/w3191 )
         );
  AND U8173 ( .A(\SUBBYTES[2].a/w3189 ), .B(n2789), .Z(\SUBBYTES[2].a/w3190 )
         );
  ANDN U8174 ( .A(\w1[2][8] ), .B(n2790), .Z(\SUBBYTES[2].a/w3186 ) );
  AND U8175 ( .A(n2791), .B(\SUBBYTES[2].a/w3061 ), .Z(\SUBBYTES[2].a/w3184 )
         );
  AND U8176 ( .A(\SUBBYTES[2].a/w3182 ), .B(n2792), .Z(\SUBBYTES[2].a/w3183 )
         );
  XOR U8177 ( .A(\SUBBYTES[2].a/w3126 ), .B(n7140), .Z(n2792) );
  AND U8178 ( .A(\SUBBYTES[2].a/w3169 ), .B(\SUBBYTES[2].a/w3171 ), .Z(
        \SUBBYTES[2].a/w3178 ) );
  AND U8179 ( .A(\SUBBYTES[2].a/w3170 ), .B(\SUBBYTES[2].a/w3172 ), .Z(
        \SUBBYTES[2].a/w3176 ) );
  AND U8180 ( .A(\SUBBYTES[2].a/w3173 ), .B(\SUBBYTES[2].a/w3174 ), .Z(
        \SUBBYTES[2].a/w3175 ) );
  AND U8181 ( .A(\SUBBYTES[2].a/w3062 ), .B(n2787), .Z(\SUBBYTES[2].a/w3161 )
         );
  XOR U8182 ( .A(\SUBBYTES[2].a/w3130 ), .B(n987), .Z(n2787) );
  AND U8183 ( .A(\SUBBYTES[2].a/w3063 ), .B(n2788), .Z(\SUBBYTES[2].a/w3159 )
         );
  XOR U8184 ( .A(n7141), .B(\SUBBYTES[2].a/w3130 ), .Z(n2788) );
  ANDN U8185 ( .A(n2789), .B(n2793), .Z(\SUBBYTES[2].a/w3158 ) );
  XOR U8186 ( .A(n987), .B(n7141), .Z(n2789) );
  ANDN U8187 ( .A(\SUBBYTES[2].a/w3064 ), .B(n2790), .Z(\SUBBYTES[2].a/w3154 )
         );
  XNOR U8188 ( .A(\SUBBYTES[2].a/w3123 ), .B(\SUBBYTES[2].a/w3126 ), .Z(n2790)
         );
  AND U8189 ( .A(\SUBBYTES[2].a/w3065 ), .B(n2791), .Z(\SUBBYTES[2].a/w3152 )
         );
  XNOR U8190 ( .A(n2794), .B(\SUBBYTES[2].a/w3123 ), .Z(n2791) );
  AND U8191 ( .A(\SUBBYTES[2].a/w3150 ), .B(n2795), .Z(\SUBBYTES[2].a/w3151 )
         );
  XOR U8192 ( .A(n2796), .B(n2794), .Z(n2795) );
  IV U8193 ( .A(n7140), .Z(n2794) );
  ANDN U8194 ( .A(\SUBBYTES[2].a/w3169 ), .B(n2797), .Z(\SUBBYTES[2].a/w3146 )
         );
  ANDN U8195 ( .A(\SUBBYTES[2].a/w3170 ), .B(n2798), .Z(\SUBBYTES[2].a/w3144 )
         );
  ANDN U8196 ( .A(\SUBBYTES[2].a/w3173 ), .B(n2799), .Z(\SUBBYTES[2].a/w3143 )
         );
  AND U8197 ( .A(\SUBBYTES[2].a/w3129 ), .B(\SUBBYTES[2].a/w3128 ), .Z(
        \SUBBYTES[2].a/w3130 ) );
  IV U8198 ( .A(n2796), .Z(\SUBBYTES[2].a/w3126 ) );
  NAND U8199 ( .A(\SUBBYTES[2].a/w3105 ), .B(\SUBBYTES[2].a/w3120 ), .Z(n2796)
         );
  AND U8200 ( .A(\SUBBYTES[2].a/w3122 ), .B(\SUBBYTES[2].a/w3128 ), .Z(
        \SUBBYTES[2].a/w3123 ) );
  AND U8201 ( .A(\SUBBYTES[2].a/w3107 ), .B(\SUBBYTES[2].a/w3105 ), .Z(
        \SUBBYTES[2].a/w3117 ) );
  AND U8202 ( .A(\SUBBYTES[2].a/w3108 ), .B(\SUBBYTES[2].a/w3106 ), .Z(
        \SUBBYTES[2].a/w3115 ) );
  AND U8203 ( .A(\SUBBYTES[2].a/w3122 ), .B(\SUBBYTES[2].a/w3129 ), .Z(
        \SUBBYTES[2].a/w3114 ) );
  AND U8204 ( .A(\SUBBYTES[2].a/w3062 ), .B(\SUBBYTES[2].a/w3058 ), .Z(
        \SUBBYTES[2].a/w3099 ) );
  AND U8205 ( .A(\SUBBYTES[2].a/w3063 ), .B(\SUBBYTES[2].a/w3059 ), .Z(
        \SUBBYTES[2].a/w3097 ) );
  ANDN U8206 ( .A(\SUBBYTES[2].a/w3189 ), .B(n2793), .Z(\SUBBYTES[2].a/w3096 )
         );
  XNOR U8207 ( .A(\w1[2][15] ), .B(\w1[2][9] ), .Z(n2793) );
  XOR U8208 ( .A(\w0[2][9] ), .B(g_input[265]), .Z(\w1[2][9] ) );
  AND U8209 ( .A(\w1[2][8] ), .B(\SUBBYTES[2].a/w3064 ), .Z(
        \SUBBYTES[2].a/w3092 ) );
  XOR U8210 ( .A(\w0[2][8] ), .B(g_input[264]), .Z(\w1[2][8] ) );
  AND U8211 ( .A(\SUBBYTES[2].a/w3065 ), .B(\SUBBYTES[2].a/w3061 ), .Z(
        \SUBBYTES[2].a/w3090 ) );
  AND U8212 ( .A(\SUBBYTES[2].a/w3150 ), .B(\SUBBYTES[2].a/w3182 ), .Z(
        \SUBBYTES[2].a/w3089 ) );
  ANDN U8213 ( .A(\SUBBYTES[2].a/w3171 ), .B(n2797), .Z(\SUBBYTES[2].a/w3084 )
         );
  XNOR U8214 ( .A(\w1[2][12] ), .B(\w1[2][15] ), .Z(n2797) );
  ANDN U8215 ( .A(\SUBBYTES[2].a/w3172 ), .B(n2798), .Z(\SUBBYTES[2].a/w3082 )
         );
  XNOR U8216 ( .A(\w1[2][10] ), .B(\w1[2][15] ), .Z(n2798) );
  XOR U8217 ( .A(\w0[2][15] ), .B(g_input[271]), .Z(\w1[2][15] ) );
  ANDN U8218 ( .A(\SUBBYTES[2].a/w3174 ), .B(n2799), .Z(\SUBBYTES[2].a/w3081 )
         );
  XNOR U8219 ( .A(\w1[2][10] ), .B(\w1[2][12] ), .Z(n2799) );
  XOR U8220 ( .A(\w0[2][12] ), .B(g_input[268]), .Z(\w1[2][12] ) );
  XOR U8221 ( .A(\w0[2][10] ), .B(g_input[266]), .Z(\w1[2][10] ) );
  AND U8222 ( .A(n2800), .B(\SUBBYTES[2].a/w2851 ), .Z(\SUBBYTES[2].a/w2986 )
         );
  AND U8223 ( .A(n2801), .B(\SUBBYTES[2].a/w2852 ), .Z(\SUBBYTES[2].a/w2984 )
         );
  AND U8224 ( .A(\SUBBYTES[2].a/w2982 ), .B(n2802), .Z(\SUBBYTES[2].a/w2983 )
         );
  ANDN U8225 ( .A(\w1[2][16] ), .B(n2803), .Z(\SUBBYTES[2].a/w2979 ) );
  AND U8226 ( .A(n2804), .B(\SUBBYTES[2].a/w2854 ), .Z(\SUBBYTES[2].a/w2977 )
         );
  AND U8227 ( .A(\SUBBYTES[2].a/w2975 ), .B(n2805), .Z(\SUBBYTES[2].a/w2976 )
         );
  XOR U8228 ( .A(\SUBBYTES[2].a/w2919 ), .B(n7138), .Z(n2805) );
  AND U8229 ( .A(\SUBBYTES[2].a/w2962 ), .B(\SUBBYTES[2].a/w2964 ), .Z(
        \SUBBYTES[2].a/w2971 ) );
  AND U8230 ( .A(\SUBBYTES[2].a/w2963 ), .B(\SUBBYTES[2].a/w2965 ), .Z(
        \SUBBYTES[2].a/w2969 ) );
  AND U8231 ( .A(\SUBBYTES[2].a/w2966 ), .B(\SUBBYTES[2].a/w2967 ), .Z(
        \SUBBYTES[2].a/w2968 ) );
  AND U8232 ( .A(\SUBBYTES[2].a/w2855 ), .B(n2800), .Z(\SUBBYTES[2].a/w2954 )
         );
  XOR U8233 ( .A(\SUBBYTES[2].a/w2923 ), .B(n986), .Z(n2800) );
  AND U8234 ( .A(\SUBBYTES[2].a/w2856 ), .B(n2801), .Z(\SUBBYTES[2].a/w2952 )
         );
  XOR U8235 ( .A(n7139), .B(\SUBBYTES[2].a/w2923 ), .Z(n2801) );
  ANDN U8236 ( .A(n2802), .B(n2806), .Z(\SUBBYTES[2].a/w2951 ) );
  XOR U8237 ( .A(n986), .B(n7139), .Z(n2802) );
  AND U8238 ( .A(n2807), .B(\SUBBYTES[2].a/w160 ), .Z(\SUBBYTES[2].a/w295 ) );
  ANDN U8239 ( .A(\SUBBYTES[2].a/w2857 ), .B(n2803), .Z(\SUBBYTES[2].a/w2947 )
         );
  XNOR U8240 ( .A(\SUBBYTES[2].a/w2916 ), .B(\SUBBYTES[2].a/w2919 ), .Z(n2803)
         );
  AND U8241 ( .A(\SUBBYTES[2].a/w2858 ), .B(n2804), .Z(\SUBBYTES[2].a/w2945 )
         );
  XNOR U8242 ( .A(n2808), .B(\SUBBYTES[2].a/w2916 ), .Z(n2804) );
  AND U8243 ( .A(\SUBBYTES[2].a/w2943 ), .B(n2809), .Z(\SUBBYTES[2].a/w2944 )
         );
  XOR U8244 ( .A(n2810), .B(n2808), .Z(n2809) );
  IV U8245 ( .A(n7138), .Z(n2808) );
  ANDN U8246 ( .A(\SUBBYTES[2].a/w2962 ), .B(n2811), .Z(\SUBBYTES[2].a/w2939 )
         );
  ANDN U8247 ( .A(\SUBBYTES[2].a/w2963 ), .B(n2812), .Z(\SUBBYTES[2].a/w2937 )
         );
  ANDN U8248 ( .A(\SUBBYTES[2].a/w2966 ), .B(n2813), .Z(\SUBBYTES[2].a/w2936 )
         );
  AND U8249 ( .A(n2814), .B(\SUBBYTES[2].a/w161 ), .Z(\SUBBYTES[2].a/w293 ) );
  AND U8250 ( .A(\SUBBYTES[2].a/w2922 ), .B(\SUBBYTES[2].a/w2921 ), .Z(
        \SUBBYTES[2].a/w2923 ) );
  AND U8251 ( .A(\SUBBYTES[2].a/w291 ), .B(n2815), .Z(\SUBBYTES[2].a/w292 ) );
  IV U8252 ( .A(n2810), .Z(\SUBBYTES[2].a/w2919 ) );
  NAND U8253 ( .A(\SUBBYTES[2].a/w2898 ), .B(\SUBBYTES[2].a/w2913 ), .Z(n2810)
         );
  AND U8254 ( .A(\SUBBYTES[2].a/w2915 ), .B(\SUBBYTES[2].a/w2921 ), .Z(
        \SUBBYTES[2].a/w2916 ) );
  AND U8255 ( .A(\SUBBYTES[2].a/w2900 ), .B(\SUBBYTES[2].a/w2898 ), .Z(
        \SUBBYTES[2].a/w2910 ) );
  AND U8256 ( .A(\SUBBYTES[2].a/w2901 ), .B(\SUBBYTES[2].a/w2899 ), .Z(
        \SUBBYTES[2].a/w2908 ) );
  AND U8257 ( .A(\SUBBYTES[2].a/w2915 ), .B(\SUBBYTES[2].a/w2922 ), .Z(
        \SUBBYTES[2].a/w2907 ) );
  AND U8258 ( .A(\SUBBYTES[2].a/w2855 ), .B(\SUBBYTES[2].a/w2851 ), .Z(
        \SUBBYTES[2].a/w2892 ) );
  AND U8259 ( .A(\SUBBYTES[2].a/w2856 ), .B(\SUBBYTES[2].a/w2852 ), .Z(
        \SUBBYTES[2].a/w2890 ) );
  ANDN U8260 ( .A(\SUBBYTES[2].a/w2982 ), .B(n2806), .Z(\SUBBYTES[2].a/w2889 )
         );
  XNOR U8261 ( .A(\w1[2][17] ), .B(\w1[2][23] ), .Z(n2806) );
  XOR U8262 ( .A(\w0[2][17] ), .B(g_input[273]), .Z(\w1[2][17] ) );
  AND U8263 ( .A(\w1[2][16] ), .B(\SUBBYTES[2].a/w2857 ), .Z(
        \SUBBYTES[2].a/w2885 ) );
  XOR U8264 ( .A(\w0[2][16] ), .B(g_input[272]), .Z(\w1[2][16] ) );
  AND U8265 ( .A(\SUBBYTES[2].a/w2858 ), .B(\SUBBYTES[2].a/w2854 ), .Z(
        \SUBBYTES[2].a/w2883 ) );
  AND U8266 ( .A(\SUBBYTES[2].a/w2943 ), .B(\SUBBYTES[2].a/w2975 ), .Z(
        \SUBBYTES[2].a/w2882 ) );
  ANDN U8267 ( .A(\w1[2][120] ), .B(n2816), .Z(\SUBBYTES[2].a/w288 ) );
  ANDN U8268 ( .A(\SUBBYTES[2].a/w2964 ), .B(n2811), .Z(\SUBBYTES[2].a/w2877 )
         );
  XNOR U8269 ( .A(\w1[2][20] ), .B(\w1[2][23] ), .Z(n2811) );
  ANDN U8270 ( .A(\SUBBYTES[2].a/w2965 ), .B(n2812), .Z(\SUBBYTES[2].a/w2875 )
         );
  XNOR U8271 ( .A(\w1[2][18] ), .B(\w1[2][23] ), .Z(n2812) );
  XOR U8272 ( .A(\w0[2][23] ), .B(g_input[279]), .Z(\w1[2][23] ) );
  IV U8273 ( .A(n2817), .Z(\w1[2][18] ) );
  ANDN U8274 ( .A(\SUBBYTES[2].a/w2967 ), .B(n2813), .Z(\SUBBYTES[2].a/w2874 )
         );
  XOR U8275 ( .A(n2817), .B(\w1[2][20] ), .Z(n2813) );
  XOR U8276 ( .A(\w0[2][20] ), .B(g_input[276]), .Z(\w1[2][20] ) );
  XNOR U8277 ( .A(\w0[2][18] ), .B(g_input[274]), .Z(n2817) );
  AND U8278 ( .A(n2818), .B(\SUBBYTES[2].a/w163 ), .Z(\SUBBYTES[2].a/w286 ) );
  AND U8279 ( .A(\SUBBYTES[2].a/w284 ), .B(n2819), .Z(\SUBBYTES[2].a/w285 ) );
  XOR U8280 ( .A(\SUBBYTES[2].a/w228 ), .B(n7112), .Z(n2819) );
  AND U8281 ( .A(\SUBBYTES[2].a/w271 ), .B(\SUBBYTES[2].a/w273 ), .Z(
        \SUBBYTES[2].a/w280 ) );
  AND U8282 ( .A(\SUBBYTES[2].a/w272 ), .B(\SUBBYTES[2].a/w274 ), .Z(
        \SUBBYTES[2].a/w278 ) );
  AND U8283 ( .A(n2820), .B(\SUBBYTES[2].a/w2644 ), .Z(\SUBBYTES[2].a/w2779 )
         );
  AND U8284 ( .A(n2821), .B(\SUBBYTES[2].a/w2645 ), .Z(\SUBBYTES[2].a/w2777 )
         );
  AND U8285 ( .A(\SUBBYTES[2].a/w2775 ), .B(n2822), .Z(\SUBBYTES[2].a/w2776 )
         );
  ANDN U8286 ( .A(\w1[2][24] ), .B(n2823), .Z(\SUBBYTES[2].a/w2772 ) );
  AND U8287 ( .A(n2824), .B(\SUBBYTES[2].a/w2647 ), .Z(\SUBBYTES[2].a/w2770 )
         );
  AND U8288 ( .A(\SUBBYTES[2].a/w275 ), .B(\SUBBYTES[2].a/w276 ), .Z(
        \SUBBYTES[2].a/w277 ) );
  AND U8289 ( .A(\SUBBYTES[2].a/w2768 ), .B(n2825), .Z(\SUBBYTES[2].a/w2769 )
         );
  XOR U8290 ( .A(\SUBBYTES[2].a/w2712 ), .B(n7136), .Z(n2825) );
  AND U8291 ( .A(\SUBBYTES[2].a/w2755 ), .B(\SUBBYTES[2].a/w2757 ), .Z(
        \SUBBYTES[2].a/w2764 ) );
  AND U8292 ( .A(\SUBBYTES[2].a/w2756 ), .B(\SUBBYTES[2].a/w2758 ), .Z(
        \SUBBYTES[2].a/w2762 ) );
  AND U8293 ( .A(\SUBBYTES[2].a/w2759 ), .B(\SUBBYTES[2].a/w2760 ), .Z(
        \SUBBYTES[2].a/w2761 ) );
  AND U8294 ( .A(\SUBBYTES[2].a/w2648 ), .B(n2820), .Z(\SUBBYTES[2].a/w2747 )
         );
  XOR U8295 ( .A(\SUBBYTES[2].a/w2716 ), .B(n985), .Z(n2820) );
  AND U8296 ( .A(\SUBBYTES[2].a/w2649 ), .B(n2821), .Z(\SUBBYTES[2].a/w2745 )
         );
  XOR U8297 ( .A(n7137), .B(\SUBBYTES[2].a/w2716 ), .Z(n2821) );
  ANDN U8298 ( .A(n2822), .B(n2826), .Z(\SUBBYTES[2].a/w2744 ) );
  XOR U8299 ( .A(n985), .B(n7137), .Z(n2822) );
  ANDN U8300 ( .A(\SUBBYTES[2].a/w2650 ), .B(n2823), .Z(\SUBBYTES[2].a/w2740 )
         );
  XNOR U8301 ( .A(\SUBBYTES[2].a/w2709 ), .B(\SUBBYTES[2].a/w2712 ), .Z(n2823)
         );
  AND U8302 ( .A(\SUBBYTES[2].a/w2651 ), .B(n2824), .Z(\SUBBYTES[2].a/w2738 )
         );
  XNOR U8303 ( .A(n2827), .B(\SUBBYTES[2].a/w2709 ), .Z(n2824) );
  AND U8304 ( .A(\SUBBYTES[2].a/w2736 ), .B(n2828), .Z(\SUBBYTES[2].a/w2737 )
         );
  XOR U8305 ( .A(n2829), .B(n2827), .Z(n2828) );
  IV U8306 ( .A(n7136), .Z(n2827) );
  ANDN U8307 ( .A(\SUBBYTES[2].a/w2755 ), .B(n2830), .Z(\SUBBYTES[2].a/w2732 )
         );
  ANDN U8308 ( .A(\SUBBYTES[2].a/w2756 ), .B(n2831), .Z(\SUBBYTES[2].a/w2730 )
         );
  ANDN U8309 ( .A(\SUBBYTES[2].a/w2759 ), .B(n2832), .Z(\SUBBYTES[2].a/w2729 )
         );
  AND U8310 ( .A(\SUBBYTES[2].a/w2715 ), .B(\SUBBYTES[2].a/w2714 ), .Z(
        \SUBBYTES[2].a/w2716 ) );
  IV U8311 ( .A(n2829), .Z(\SUBBYTES[2].a/w2712 ) );
  NAND U8312 ( .A(\SUBBYTES[2].a/w2691 ), .B(\SUBBYTES[2].a/w2706 ), .Z(n2829)
         );
  AND U8313 ( .A(\SUBBYTES[2].a/w2708 ), .B(\SUBBYTES[2].a/w2714 ), .Z(
        \SUBBYTES[2].a/w2709 ) );
  AND U8314 ( .A(\SUBBYTES[2].a/w2693 ), .B(\SUBBYTES[2].a/w2691 ), .Z(
        \SUBBYTES[2].a/w2703 ) );
  AND U8315 ( .A(\SUBBYTES[2].a/w2694 ), .B(\SUBBYTES[2].a/w2692 ), .Z(
        \SUBBYTES[2].a/w2701 ) );
  AND U8316 ( .A(\SUBBYTES[2].a/w2708 ), .B(\SUBBYTES[2].a/w2715 ), .Z(
        \SUBBYTES[2].a/w2700 ) );
  AND U8317 ( .A(\SUBBYTES[2].a/w2648 ), .B(\SUBBYTES[2].a/w2644 ), .Z(
        \SUBBYTES[2].a/w2685 ) );
  AND U8318 ( .A(\SUBBYTES[2].a/w2649 ), .B(\SUBBYTES[2].a/w2645 ), .Z(
        \SUBBYTES[2].a/w2683 ) );
  ANDN U8319 ( .A(\SUBBYTES[2].a/w2775 ), .B(n2826), .Z(\SUBBYTES[2].a/w2682 )
         );
  XNOR U8320 ( .A(\w1[2][25] ), .B(\w1[2][31] ), .Z(n2826) );
  XOR U8321 ( .A(\w0[2][25] ), .B(g_input[281]), .Z(\w1[2][25] ) );
  AND U8322 ( .A(\w1[2][24] ), .B(\SUBBYTES[2].a/w2650 ), .Z(
        \SUBBYTES[2].a/w2678 ) );
  XOR U8323 ( .A(\w0[2][24] ), .B(g_input[280]), .Z(\w1[2][24] ) );
  AND U8324 ( .A(\SUBBYTES[2].a/w2651 ), .B(\SUBBYTES[2].a/w2647 ), .Z(
        \SUBBYTES[2].a/w2676 ) );
  AND U8325 ( .A(\SUBBYTES[2].a/w2736 ), .B(\SUBBYTES[2].a/w2768 ), .Z(
        \SUBBYTES[2].a/w2675 ) );
  ANDN U8326 ( .A(\SUBBYTES[2].a/w2757 ), .B(n2830), .Z(\SUBBYTES[2].a/w2670 )
         );
  XNOR U8327 ( .A(\w1[2][28] ), .B(\w1[2][31] ), .Z(n2830) );
  ANDN U8328 ( .A(\SUBBYTES[2].a/w2758 ), .B(n2831), .Z(\SUBBYTES[2].a/w2668 )
         );
  XNOR U8329 ( .A(\w1[2][26] ), .B(\w1[2][31] ), .Z(n2831) );
  XOR U8330 ( .A(\w0[2][31] ), .B(g_input[287]), .Z(\w1[2][31] ) );
  IV U8331 ( .A(n2833), .Z(\w1[2][26] ) );
  ANDN U8332 ( .A(\SUBBYTES[2].a/w2760 ), .B(n2832), .Z(\SUBBYTES[2].a/w2667 )
         );
  XOR U8333 ( .A(n2833), .B(\w1[2][28] ), .Z(n2832) );
  XOR U8334 ( .A(\w0[2][28] ), .B(g_input[284]), .Z(\w1[2][28] ) );
  XNOR U8335 ( .A(\w0[2][26] ), .B(g_input[282]), .Z(n2833) );
  AND U8336 ( .A(\SUBBYTES[2].a/w164 ), .B(n2807), .Z(\SUBBYTES[2].a/w263 ) );
  XOR U8337 ( .A(\SUBBYTES[2].a/w232 ), .B(n973), .Z(n2807) );
  AND U8338 ( .A(\SUBBYTES[2].a/w165 ), .B(n2814), .Z(\SUBBYTES[2].a/w261 ) );
  XOR U8339 ( .A(n7113), .B(\SUBBYTES[2].a/w232 ), .Z(n2814) );
  ANDN U8340 ( .A(n2815), .B(n2834), .Z(\SUBBYTES[2].a/w260 ) );
  XOR U8341 ( .A(n973), .B(n7113), .Z(n2815) );
  AND U8342 ( .A(n2835), .B(\SUBBYTES[2].a/w2437 ), .Z(\SUBBYTES[2].a/w2572 )
         );
  AND U8343 ( .A(n2836), .B(\SUBBYTES[2].a/w2438 ), .Z(\SUBBYTES[2].a/w2570 )
         );
  AND U8344 ( .A(\SUBBYTES[2].a/w2568 ), .B(n2837), .Z(\SUBBYTES[2].a/w2569 )
         );
  ANDN U8345 ( .A(\w1[2][32] ), .B(n2838), .Z(\SUBBYTES[2].a/w2565 ) );
  AND U8346 ( .A(n2839), .B(\SUBBYTES[2].a/w2440 ), .Z(\SUBBYTES[2].a/w2563 )
         );
  AND U8347 ( .A(\SUBBYTES[2].a/w2561 ), .B(n2840), .Z(\SUBBYTES[2].a/w2562 )
         );
  XOR U8348 ( .A(\SUBBYTES[2].a/w2505 ), .B(n7134), .Z(n2840) );
  ANDN U8349 ( .A(\SUBBYTES[2].a/w166 ), .B(n2816), .Z(\SUBBYTES[2].a/w256 )
         );
  XNOR U8350 ( .A(\SUBBYTES[2].a/w225 ), .B(\SUBBYTES[2].a/w228 ), .Z(n2816)
         );
  AND U8351 ( .A(\SUBBYTES[2].a/w2548 ), .B(\SUBBYTES[2].a/w2550 ), .Z(
        \SUBBYTES[2].a/w2557 ) );
  AND U8352 ( .A(\SUBBYTES[2].a/w2549 ), .B(\SUBBYTES[2].a/w2551 ), .Z(
        \SUBBYTES[2].a/w2555 ) );
  AND U8353 ( .A(\SUBBYTES[2].a/w2552 ), .B(\SUBBYTES[2].a/w2553 ), .Z(
        \SUBBYTES[2].a/w2554 ) );
  AND U8354 ( .A(\SUBBYTES[2].a/w2441 ), .B(n2835), .Z(\SUBBYTES[2].a/w2540 )
         );
  XOR U8355 ( .A(\SUBBYTES[2].a/w2509 ), .B(n984), .Z(n2835) );
  AND U8356 ( .A(\SUBBYTES[2].a/w167 ), .B(n2818), .Z(\SUBBYTES[2].a/w254 ) );
  XNOR U8357 ( .A(n2841), .B(\SUBBYTES[2].a/w225 ), .Z(n2818) );
  AND U8358 ( .A(\SUBBYTES[2].a/w2442 ), .B(n2836), .Z(\SUBBYTES[2].a/w2538 )
         );
  XOR U8359 ( .A(n7135), .B(\SUBBYTES[2].a/w2509 ), .Z(n2836) );
  ANDN U8360 ( .A(n2837), .B(n2842), .Z(\SUBBYTES[2].a/w2537 ) );
  XOR U8361 ( .A(n984), .B(n7135), .Z(n2837) );
  ANDN U8362 ( .A(\SUBBYTES[2].a/w2443 ), .B(n2838), .Z(\SUBBYTES[2].a/w2533 )
         );
  XNOR U8363 ( .A(\SUBBYTES[2].a/w2502 ), .B(\SUBBYTES[2].a/w2505 ), .Z(n2838)
         );
  AND U8364 ( .A(\SUBBYTES[2].a/w2444 ), .B(n2839), .Z(\SUBBYTES[2].a/w2531 )
         );
  XNOR U8365 ( .A(n2843), .B(\SUBBYTES[2].a/w2502 ), .Z(n2839) );
  AND U8366 ( .A(\SUBBYTES[2].a/w2529 ), .B(n2844), .Z(\SUBBYTES[2].a/w2530 )
         );
  XOR U8367 ( .A(n2845), .B(n2843), .Z(n2844) );
  IV U8368 ( .A(n7134), .Z(n2843) );
  AND U8369 ( .A(\SUBBYTES[2].a/w252 ), .B(n2846), .Z(\SUBBYTES[2].a/w253 ) );
  XOR U8370 ( .A(n2847), .B(n2841), .Z(n2846) );
  IV U8371 ( .A(n7112), .Z(n2841) );
  ANDN U8372 ( .A(\SUBBYTES[2].a/w2548 ), .B(n2848), .Z(\SUBBYTES[2].a/w2525 )
         );
  ANDN U8373 ( .A(\SUBBYTES[2].a/w2549 ), .B(n2849), .Z(\SUBBYTES[2].a/w2523 )
         );
  ANDN U8374 ( .A(\SUBBYTES[2].a/w2552 ), .B(n2850), .Z(\SUBBYTES[2].a/w2522 )
         );
  AND U8375 ( .A(\SUBBYTES[2].a/w2508 ), .B(\SUBBYTES[2].a/w2507 ), .Z(
        \SUBBYTES[2].a/w2509 ) );
  IV U8376 ( .A(n2845), .Z(\SUBBYTES[2].a/w2505 ) );
  NAND U8377 ( .A(\SUBBYTES[2].a/w2484 ), .B(\SUBBYTES[2].a/w2499 ), .Z(n2845)
         );
  AND U8378 ( .A(\SUBBYTES[2].a/w2501 ), .B(\SUBBYTES[2].a/w2507 ), .Z(
        \SUBBYTES[2].a/w2502 ) );
  AND U8379 ( .A(\SUBBYTES[2].a/w2486 ), .B(\SUBBYTES[2].a/w2484 ), .Z(
        \SUBBYTES[2].a/w2496 ) );
  AND U8380 ( .A(\SUBBYTES[2].a/w2487 ), .B(\SUBBYTES[2].a/w2485 ), .Z(
        \SUBBYTES[2].a/w2494 ) );
  AND U8381 ( .A(\SUBBYTES[2].a/w2501 ), .B(\SUBBYTES[2].a/w2508 ), .Z(
        \SUBBYTES[2].a/w2493 ) );
  ANDN U8382 ( .A(\SUBBYTES[2].a/w271 ), .B(n2851), .Z(\SUBBYTES[2].a/w248 )
         );
  AND U8383 ( .A(\SUBBYTES[2].a/w2441 ), .B(\SUBBYTES[2].a/w2437 ), .Z(
        \SUBBYTES[2].a/w2478 ) );
  AND U8384 ( .A(\SUBBYTES[2].a/w2442 ), .B(\SUBBYTES[2].a/w2438 ), .Z(
        \SUBBYTES[2].a/w2476 ) );
  ANDN U8385 ( .A(\SUBBYTES[2].a/w2568 ), .B(n2842), .Z(\SUBBYTES[2].a/w2475 )
         );
  XNOR U8386 ( .A(\w1[2][33] ), .B(\w1[2][39] ), .Z(n2842) );
  XOR U8387 ( .A(\w0[2][33] ), .B(g_input[289]), .Z(\w1[2][33] ) );
  AND U8388 ( .A(\w1[2][32] ), .B(\SUBBYTES[2].a/w2443 ), .Z(
        \SUBBYTES[2].a/w2471 ) );
  XOR U8389 ( .A(\w0[2][32] ), .B(g_input[288]), .Z(\w1[2][32] ) );
  AND U8390 ( .A(\SUBBYTES[2].a/w2444 ), .B(\SUBBYTES[2].a/w2440 ), .Z(
        \SUBBYTES[2].a/w2469 ) );
  AND U8391 ( .A(\SUBBYTES[2].a/w2529 ), .B(\SUBBYTES[2].a/w2561 ), .Z(
        \SUBBYTES[2].a/w2468 ) );
  ANDN U8392 ( .A(\SUBBYTES[2].a/w2550 ), .B(n2848), .Z(\SUBBYTES[2].a/w2463 )
         );
  XNOR U8393 ( .A(\w1[2][36] ), .B(\w1[2][39] ), .Z(n2848) );
  ANDN U8394 ( .A(\SUBBYTES[2].a/w2551 ), .B(n2849), .Z(\SUBBYTES[2].a/w2461 )
         );
  XNOR U8395 ( .A(\w1[2][34] ), .B(\w1[2][39] ), .Z(n2849) );
  XOR U8396 ( .A(\w0[2][39] ), .B(g_input[295]), .Z(\w1[2][39] ) );
  IV U8397 ( .A(n2852), .Z(\w1[2][34] ) );
  ANDN U8398 ( .A(\SUBBYTES[2].a/w2553 ), .B(n2850), .Z(\SUBBYTES[2].a/w2460 )
         );
  XOR U8399 ( .A(n2852), .B(\w1[2][36] ), .Z(n2850) );
  XOR U8400 ( .A(\w0[2][36] ), .B(g_input[292]), .Z(\w1[2][36] ) );
  XNOR U8401 ( .A(\w0[2][34] ), .B(g_input[290]), .Z(n2852) );
  ANDN U8402 ( .A(\SUBBYTES[2].a/w272 ), .B(n2853), .Z(\SUBBYTES[2].a/w246 )
         );
  ANDN U8403 ( .A(\SUBBYTES[2].a/w275 ), .B(n2854), .Z(\SUBBYTES[2].a/w245 )
         );
  AND U8404 ( .A(n2855), .B(\SUBBYTES[2].a/w2230 ), .Z(\SUBBYTES[2].a/w2365 )
         );
  AND U8405 ( .A(n2856), .B(\SUBBYTES[2].a/w2231 ), .Z(\SUBBYTES[2].a/w2363 )
         );
  AND U8406 ( .A(\SUBBYTES[2].a/w2361 ), .B(n2857), .Z(\SUBBYTES[2].a/w2362 )
         );
  ANDN U8407 ( .A(\w1[2][40] ), .B(n2858), .Z(\SUBBYTES[2].a/w2358 ) );
  AND U8408 ( .A(n2859), .B(\SUBBYTES[2].a/w2233 ), .Z(\SUBBYTES[2].a/w2356 )
         );
  AND U8409 ( .A(\SUBBYTES[2].a/w2354 ), .B(n2860), .Z(\SUBBYTES[2].a/w2355 )
         );
  XOR U8410 ( .A(\SUBBYTES[2].a/w2298 ), .B(n7132), .Z(n2860) );
  AND U8411 ( .A(\SUBBYTES[2].a/w2341 ), .B(\SUBBYTES[2].a/w2343 ), .Z(
        \SUBBYTES[2].a/w2350 ) );
  AND U8412 ( .A(\SUBBYTES[2].a/w2342 ), .B(\SUBBYTES[2].a/w2344 ), .Z(
        \SUBBYTES[2].a/w2348 ) );
  AND U8413 ( .A(\SUBBYTES[2].a/w2345 ), .B(\SUBBYTES[2].a/w2346 ), .Z(
        \SUBBYTES[2].a/w2347 ) );
  AND U8414 ( .A(\SUBBYTES[2].a/w2234 ), .B(n2855), .Z(\SUBBYTES[2].a/w2333 )
         );
  XOR U8415 ( .A(\SUBBYTES[2].a/w2302 ), .B(n983), .Z(n2855) );
  AND U8416 ( .A(\SUBBYTES[2].a/w2235 ), .B(n2856), .Z(\SUBBYTES[2].a/w2331 )
         );
  XOR U8417 ( .A(n7133), .B(\SUBBYTES[2].a/w2302 ), .Z(n2856) );
  ANDN U8418 ( .A(n2857), .B(n2861), .Z(\SUBBYTES[2].a/w2330 ) );
  XOR U8419 ( .A(n983), .B(n7133), .Z(n2857) );
  ANDN U8420 ( .A(\SUBBYTES[2].a/w2236 ), .B(n2858), .Z(\SUBBYTES[2].a/w2326 )
         );
  XNOR U8421 ( .A(\SUBBYTES[2].a/w2295 ), .B(\SUBBYTES[2].a/w2298 ), .Z(n2858)
         );
  AND U8422 ( .A(\SUBBYTES[2].a/w2237 ), .B(n2859), .Z(\SUBBYTES[2].a/w2324 )
         );
  XNOR U8423 ( .A(n2862), .B(\SUBBYTES[2].a/w2295 ), .Z(n2859) );
  AND U8424 ( .A(\SUBBYTES[2].a/w2322 ), .B(n2863), .Z(\SUBBYTES[2].a/w2323 )
         );
  XOR U8425 ( .A(n2864), .B(n2862), .Z(n2863) );
  IV U8426 ( .A(n7132), .Z(n2862) );
  AND U8427 ( .A(\SUBBYTES[2].a/w231 ), .B(\SUBBYTES[2].a/w230 ), .Z(
        \SUBBYTES[2].a/w232 ) );
  ANDN U8428 ( .A(\SUBBYTES[2].a/w2341 ), .B(n2865), .Z(\SUBBYTES[2].a/w2318 )
         );
  ANDN U8429 ( .A(\SUBBYTES[2].a/w2342 ), .B(n2866), .Z(\SUBBYTES[2].a/w2316 )
         );
  ANDN U8430 ( .A(\SUBBYTES[2].a/w2345 ), .B(n2867), .Z(\SUBBYTES[2].a/w2315 )
         );
  AND U8431 ( .A(\SUBBYTES[2].a/w2301 ), .B(\SUBBYTES[2].a/w2300 ), .Z(
        \SUBBYTES[2].a/w2302 ) );
  IV U8432 ( .A(n2864), .Z(\SUBBYTES[2].a/w2298 ) );
  NAND U8433 ( .A(\SUBBYTES[2].a/w2277 ), .B(\SUBBYTES[2].a/w2292 ), .Z(n2864)
         );
  AND U8434 ( .A(\SUBBYTES[2].a/w2294 ), .B(\SUBBYTES[2].a/w2300 ), .Z(
        \SUBBYTES[2].a/w2295 ) );
  AND U8435 ( .A(\SUBBYTES[2].a/w2279 ), .B(\SUBBYTES[2].a/w2277 ), .Z(
        \SUBBYTES[2].a/w2289 ) );
  AND U8436 ( .A(\SUBBYTES[2].a/w2280 ), .B(\SUBBYTES[2].a/w2278 ), .Z(
        \SUBBYTES[2].a/w2287 ) );
  AND U8437 ( .A(\SUBBYTES[2].a/w2294 ), .B(\SUBBYTES[2].a/w2301 ), .Z(
        \SUBBYTES[2].a/w2286 ) );
  IV U8438 ( .A(n2847), .Z(\SUBBYTES[2].a/w228 ) );
  NAND U8439 ( .A(\SUBBYTES[2].a/w207 ), .B(\SUBBYTES[2].a/w222 ), .Z(n2847)
         );
  AND U8440 ( .A(\SUBBYTES[2].a/w2234 ), .B(\SUBBYTES[2].a/w2230 ), .Z(
        \SUBBYTES[2].a/w2271 ) );
  AND U8441 ( .A(\SUBBYTES[2].a/w2235 ), .B(\SUBBYTES[2].a/w2231 ), .Z(
        \SUBBYTES[2].a/w2269 ) );
  ANDN U8442 ( .A(\SUBBYTES[2].a/w2361 ), .B(n2861), .Z(\SUBBYTES[2].a/w2268 )
         );
  XNOR U8443 ( .A(\w1[2][41] ), .B(\w1[2][47] ), .Z(n2861) );
  XOR U8444 ( .A(\w0[2][41] ), .B(g_input[297]), .Z(\w1[2][41] ) );
  AND U8445 ( .A(\w1[2][40] ), .B(\SUBBYTES[2].a/w2236 ), .Z(
        \SUBBYTES[2].a/w2264 ) );
  XOR U8446 ( .A(\w0[2][40] ), .B(g_input[296]), .Z(\w1[2][40] ) );
  AND U8447 ( .A(\SUBBYTES[2].a/w2237 ), .B(\SUBBYTES[2].a/w2233 ), .Z(
        \SUBBYTES[2].a/w2262 ) );
  AND U8448 ( .A(\SUBBYTES[2].a/w2322 ), .B(\SUBBYTES[2].a/w2354 ), .Z(
        \SUBBYTES[2].a/w2261 ) );
  ANDN U8449 ( .A(\SUBBYTES[2].a/w2343 ), .B(n2865), .Z(\SUBBYTES[2].a/w2256 )
         );
  XNOR U8450 ( .A(\w1[2][44] ), .B(\w1[2][47] ), .Z(n2865) );
  ANDN U8451 ( .A(\SUBBYTES[2].a/w2344 ), .B(n2866), .Z(\SUBBYTES[2].a/w2254 )
         );
  XNOR U8452 ( .A(\w1[2][42] ), .B(\w1[2][47] ), .Z(n2866) );
  XOR U8453 ( .A(\w0[2][47] ), .B(g_input[303]), .Z(\w1[2][47] ) );
  IV U8454 ( .A(n2868), .Z(\w1[2][42] ) );
  ANDN U8455 ( .A(\SUBBYTES[2].a/w2346 ), .B(n2867), .Z(\SUBBYTES[2].a/w2253 )
         );
  XOR U8456 ( .A(n2868), .B(\w1[2][44] ), .Z(n2867) );
  XOR U8457 ( .A(\w0[2][44] ), .B(g_input[300]), .Z(\w1[2][44] ) );
  XNOR U8458 ( .A(\w0[2][42] ), .B(g_input[298]), .Z(n2868) );
  AND U8459 ( .A(\SUBBYTES[2].a/w224 ), .B(\SUBBYTES[2].a/w230 ), .Z(
        \SUBBYTES[2].a/w225 ) );
  AND U8460 ( .A(\SUBBYTES[2].a/w209 ), .B(\SUBBYTES[2].a/w207 ), .Z(
        \SUBBYTES[2].a/w219 ) );
  AND U8461 ( .A(\SUBBYTES[2].a/w210 ), .B(\SUBBYTES[2].a/w208 ), .Z(
        \SUBBYTES[2].a/w217 ) );
  AND U8462 ( .A(\SUBBYTES[2].a/w224 ), .B(\SUBBYTES[2].a/w231 ), .Z(
        \SUBBYTES[2].a/w216 ) );
  AND U8463 ( .A(n2869), .B(\SUBBYTES[2].a/w2023 ), .Z(\SUBBYTES[2].a/w2158 )
         );
  AND U8464 ( .A(n2870), .B(\SUBBYTES[2].a/w2024 ), .Z(\SUBBYTES[2].a/w2156 )
         );
  AND U8465 ( .A(\SUBBYTES[2].a/w2154 ), .B(n2871), .Z(\SUBBYTES[2].a/w2155 )
         );
  ANDN U8466 ( .A(\w1[2][48] ), .B(n2872), .Z(\SUBBYTES[2].a/w2151 ) );
  AND U8467 ( .A(n2873), .B(\SUBBYTES[2].a/w2026 ), .Z(\SUBBYTES[2].a/w2149 )
         );
  AND U8468 ( .A(\SUBBYTES[2].a/w2147 ), .B(n2874), .Z(\SUBBYTES[2].a/w2148 )
         );
  XOR U8469 ( .A(\SUBBYTES[2].a/w2091 ), .B(n7130), .Z(n2874) );
  AND U8470 ( .A(\SUBBYTES[2].a/w2134 ), .B(\SUBBYTES[2].a/w2136 ), .Z(
        \SUBBYTES[2].a/w2143 ) );
  AND U8471 ( .A(\SUBBYTES[2].a/w2135 ), .B(\SUBBYTES[2].a/w2137 ), .Z(
        \SUBBYTES[2].a/w2141 ) );
  AND U8472 ( .A(\SUBBYTES[2].a/w2138 ), .B(\SUBBYTES[2].a/w2139 ), .Z(
        \SUBBYTES[2].a/w2140 ) );
  AND U8473 ( .A(\SUBBYTES[2].a/w2027 ), .B(n2869), .Z(\SUBBYTES[2].a/w2126 )
         );
  XOR U8474 ( .A(\SUBBYTES[2].a/w2095 ), .B(n982), .Z(n2869) );
  AND U8475 ( .A(\SUBBYTES[2].a/w2028 ), .B(n2870), .Z(\SUBBYTES[2].a/w2124 )
         );
  XOR U8476 ( .A(n7131), .B(\SUBBYTES[2].a/w2095 ), .Z(n2870) );
  ANDN U8477 ( .A(n2871), .B(n2875), .Z(\SUBBYTES[2].a/w2123 ) );
  XOR U8478 ( .A(n982), .B(n7131), .Z(n2871) );
  ANDN U8479 ( .A(\SUBBYTES[2].a/w2029 ), .B(n2872), .Z(\SUBBYTES[2].a/w2119 )
         );
  XNOR U8480 ( .A(\SUBBYTES[2].a/w2088 ), .B(\SUBBYTES[2].a/w2091 ), .Z(n2872)
         );
  AND U8481 ( .A(\SUBBYTES[2].a/w2030 ), .B(n2873), .Z(\SUBBYTES[2].a/w2117 )
         );
  XNOR U8482 ( .A(n2876), .B(\SUBBYTES[2].a/w2088 ), .Z(n2873) );
  AND U8483 ( .A(\SUBBYTES[2].a/w2115 ), .B(n2877), .Z(\SUBBYTES[2].a/w2116 )
         );
  XOR U8484 ( .A(n2878), .B(n2876), .Z(n2877) );
  IV U8485 ( .A(n7130), .Z(n2876) );
  ANDN U8486 ( .A(\SUBBYTES[2].a/w2134 ), .B(n2879), .Z(\SUBBYTES[2].a/w2111 )
         );
  ANDN U8487 ( .A(\SUBBYTES[2].a/w2135 ), .B(n2880), .Z(\SUBBYTES[2].a/w2109 )
         );
  ANDN U8488 ( .A(\SUBBYTES[2].a/w2138 ), .B(n2881), .Z(\SUBBYTES[2].a/w2108 )
         );
  AND U8489 ( .A(\SUBBYTES[2].a/w2094 ), .B(\SUBBYTES[2].a/w2093 ), .Z(
        \SUBBYTES[2].a/w2095 ) );
  IV U8490 ( .A(n2878), .Z(\SUBBYTES[2].a/w2091 ) );
  NAND U8491 ( .A(\SUBBYTES[2].a/w2070 ), .B(\SUBBYTES[2].a/w2085 ), .Z(n2878)
         );
  AND U8492 ( .A(\SUBBYTES[2].a/w2087 ), .B(\SUBBYTES[2].a/w2093 ), .Z(
        \SUBBYTES[2].a/w2088 ) );
  AND U8493 ( .A(\SUBBYTES[2].a/w2072 ), .B(\SUBBYTES[2].a/w2070 ), .Z(
        \SUBBYTES[2].a/w2082 ) );
  AND U8494 ( .A(\SUBBYTES[2].a/w2073 ), .B(\SUBBYTES[2].a/w2071 ), .Z(
        \SUBBYTES[2].a/w2080 ) );
  AND U8495 ( .A(\SUBBYTES[2].a/w2087 ), .B(\SUBBYTES[2].a/w2094 ), .Z(
        \SUBBYTES[2].a/w2079 ) );
  AND U8496 ( .A(\SUBBYTES[2].a/w2027 ), .B(\SUBBYTES[2].a/w2023 ), .Z(
        \SUBBYTES[2].a/w2064 ) );
  AND U8497 ( .A(\SUBBYTES[2].a/w2028 ), .B(\SUBBYTES[2].a/w2024 ), .Z(
        \SUBBYTES[2].a/w2062 ) );
  ANDN U8498 ( .A(\SUBBYTES[2].a/w2154 ), .B(n2875), .Z(\SUBBYTES[2].a/w2061 )
         );
  XNOR U8499 ( .A(\w1[2][49] ), .B(\w1[2][55] ), .Z(n2875) );
  XOR U8500 ( .A(\w0[2][49] ), .B(g_input[305]), .Z(\w1[2][49] ) );
  AND U8501 ( .A(\w1[2][48] ), .B(\SUBBYTES[2].a/w2029 ), .Z(
        \SUBBYTES[2].a/w2057 ) );
  XOR U8502 ( .A(\w0[2][48] ), .B(g_input[304]), .Z(\w1[2][48] ) );
  AND U8503 ( .A(\SUBBYTES[2].a/w2030 ), .B(\SUBBYTES[2].a/w2026 ), .Z(
        \SUBBYTES[2].a/w2055 ) );
  AND U8504 ( .A(\SUBBYTES[2].a/w2115 ), .B(\SUBBYTES[2].a/w2147 ), .Z(
        \SUBBYTES[2].a/w2054 ) );
  ANDN U8505 ( .A(\SUBBYTES[2].a/w2136 ), .B(n2879), .Z(\SUBBYTES[2].a/w2049 )
         );
  XNOR U8506 ( .A(\w1[2][52] ), .B(\w1[2][55] ), .Z(n2879) );
  ANDN U8507 ( .A(\SUBBYTES[2].a/w2137 ), .B(n2880), .Z(\SUBBYTES[2].a/w2047 )
         );
  XNOR U8508 ( .A(\w1[2][50] ), .B(\w1[2][55] ), .Z(n2880) );
  XOR U8509 ( .A(\w0[2][55] ), .B(g_input[311]), .Z(\w1[2][55] ) );
  IV U8510 ( .A(n2882), .Z(\w1[2][50] ) );
  ANDN U8511 ( .A(\SUBBYTES[2].a/w2139 ), .B(n2881), .Z(\SUBBYTES[2].a/w2046 )
         );
  XOR U8512 ( .A(n2882), .B(\w1[2][52] ), .Z(n2881) );
  XOR U8513 ( .A(\w0[2][52] ), .B(g_input[308]), .Z(\w1[2][52] ) );
  XNOR U8514 ( .A(\w0[2][50] ), .B(g_input[306]), .Z(n2882) );
  AND U8515 ( .A(\SUBBYTES[2].a/w164 ), .B(\SUBBYTES[2].a/w160 ), .Z(
        \SUBBYTES[2].a/w201 ) );
  AND U8516 ( .A(\SUBBYTES[2].a/w165 ), .B(\SUBBYTES[2].a/w161 ), .Z(
        \SUBBYTES[2].a/w199 ) );
  ANDN U8517 ( .A(\SUBBYTES[2].a/w291 ), .B(n2834), .Z(\SUBBYTES[2].a/w198 )
         );
  XNOR U8518 ( .A(\w1[2][121] ), .B(\w1[2][127] ), .Z(n2834) );
  XOR U8519 ( .A(\w0[2][121] ), .B(g_input[377]), .Z(\w1[2][121] ) );
  AND U8520 ( .A(n2883), .B(\SUBBYTES[2].a/w1816 ), .Z(\SUBBYTES[2].a/w1951 )
         );
  AND U8521 ( .A(n2884), .B(\SUBBYTES[2].a/w1817 ), .Z(\SUBBYTES[2].a/w1949 )
         );
  AND U8522 ( .A(\SUBBYTES[2].a/w1947 ), .B(n2885), .Z(\SUBBYTES[2].a/w1948 )
         );
  ANDN U8523 ( .A(\w1[2][56] ), .B(n2886), .Z(\SUBBYTES[2].a/w1944 ) );
  AND U8524 ( .A(n2887), .B(\SUBBYTES[2].a/w1819 ), .Z(\SUBBYTES[2].a/w1942 )
         );
  AND U8525 ( .A(\SUBBYTES[2].a/w1940 ), .B(n2888), .Z(\SUBBYTES[2].a/w1941 )
         );
  XOR U8526 ( .A(\SUBBYTES[2].a/w1884 ), .B(n7128), .Z(n2888) );
  AND U8527 ( .A(\w1[2][120] ), .B(\SUBBYTES[2].a/w166 ), .Z(
        \SUBBYTES[2].a/w194 ) );
  XOR U8528 ( .A(\w0[2][120] ), .B(g_input[376]), .Z(\w1[2][120] ) );
  AND U8529 ( .A(\SUBBYTES[2].a/w1927 ), .B(\SUBBYTES[2].a/w1929 ), .Z(
        \SUBBYTES[2].a/w1936 ) );
  AND U8530 ( .A(\SUBBYTES[2].a/w1928 ), .B(\SUBBYTES[2].a/w1930 ), .Z(
        \SUBBYTES[2].a/w1934 ) );
  AND U8531 ( .A(\SUBBYTES[2].a/w1931 ), .B(\SUBBYTES[2].a/w1932 ), .Z(
        \SUBBYTES[2].a/w1933 ) );
  AND U8532 ( .A(\SUBBYTES[2].a/w167 ), .B(\SUBBYTES[2].a/w163 ), .Z(
        \SUBBYTES[2].a/w192 ) );
  AND U8533 ( .A(\SUBBYTES[2].a/w1820 ), .B(n2883), .Z(\SUBBYTES[2].a/w1919 )
         );
  XOR U8534 ( .A(\SUBBYTES[2].a/w1888 ), .B(n981), .Z(n2883) );
  AND U8535 ( .A(\SUBBYTES[2].a/w1821 ), .B(n2884), .Z(\SUBBYTES[2].a/w1917 )
         );
  XOR U8536 ( .A(n7129), .B(\SUBBYTES[2].a/w1888 ), .Z(n2884) );
  ANDN U8537 ( .A(n2885), .B(n2889), .Z(\SUBBYTES[2].a/w1916 ) );
  XOR U8538 ( .A(n981), .B(n7129), .Z(n2885) );
  ANDN U8539 ( .A(\SUBBYTES[2].a/w1822 ), .B(n2886), .Z(\SUBBYTES[2].a/w1912 )
         );
  XNOR U8540 ( .A(\SUBBYTES[2].a/w1881 ), .B(\SUBBYTES[2].a/w1884 ), .Z(n2886)
         );
  AND U8541 ( .A(\SUBBYTES[2].a/w1823 ), .B(n2887), .Z(\SUBBYTES[2].a/w1910 )
         );
  XNOR U8542 ( .A(n2890), .B(\SUBBYTES[2].a/w1881 ), .Z(n2887) );
  AND U8543 ( .A(\SUBBYTES[2].a/w252 ), .B(\SUBBYTES[2].a/w284 ), .Z(
        \SUBBYTES[2].a/w191 ) );
  AND U8544 ( .A(\SUBBYTES[2].a/w1908 ), .B(n2891), .Z(\SUBBYTES[2].a/w1909 )
         );
  XOR U8545 ( .A(n2892), .B(n2890), .Z(n2891) );
  IV U8546 ( .A(n7128), .Z(n2890) );
  ANDN U8547 ( .A(\SUBBYTES[2].a/w1927 ), .B(n2893), .Z(\SUBBYTES[2].a/w1904 )
         );
  ANDN U8548 ( .A(\SUBBYTES[2].a/w1928 ), .B(n2894), .Z(\SUBBYTES[2].a/w1902 )
         );
  ANDN U8549 ( .A(\SUBBYTES[2].a/w1931 ), .B(n2895), .Z(\SUBBYTES[2].a/w1901 )
         );
  AND U8550 ( .A(\SUBBYTES[2].a/w1887 ), .B(\SUBBYTES[2].a/w1886 ), .Z(
        \SUBBYTES[2].a/w1888 ) );
  IV U8551 ( .A(n2892), .Z(\SUBBYTES[2].a/w1884 ) );
  NAND U8552 ( .A(\SUBBYTES[2].a/w1863 ), .B(\SUBBYTES[2].a/w1878 ), .Z(n2892)
         );
  AND U8553 ( .A(\SUBBYTES[2].a/w1880 ), .B(\SUBBYTES[2].a/w1886 ), .Z(
        \SUBBYTES[2].a/w1881 ) );
  AND U8554 ( .A(\SUBBYTES[2].a/w1865 ), .B(\SUBBYTES[2].a/w1863 ), .Z(
        \SUBBYTES[2].a/w1875 ) );
  AND U8555 ( .A(\SUBBYTES[2].a/w1866 ), .B(\SUBBYTES[2].a/w1864 ), .Z(
        \SUBBYTES[2].a/w1873 ) );
  AND U8556 ( .A(\SUBBYTES[2].a/w1880 ), .B(\SUBBYTES[2].a/w1887 ), .Z(
        \SUBBYTES[2].a/w1872 ) );
  ANDN U8557 ( .A(\SUBBYTES[2].a/w273 ), .B(n2851), .Z(\SUBBYTES[2].a/w186 )
         );
  XNOR U8558 ( .A(\w1[2][124] ), .B(\w1[2][127] ), .Z(n2851) );
  AND U8559 ( .A(\SUBBYTES[2].a/w1820 ), .B(\SUBBYTES[2].a/w1816 ), .Z(
        \SUBBYTES[2].a/w1857 ) );
  AND U8560 ( .A(\SUBBYTES[2].a/w1821 ), .B(\SUBBYTES[2].a/w1817 ), .Z(
        \SUBBYTES[2].a/w1855 ) );
  ANDN U8561 ( .A(\SUBBYTES[2].a/w1947 ), .B(n2889), .Z(\SUBBYTES[2].a/w1854 )
         );
  XNOR U8562 ( .A(\w1[2][57] ), .B(\w1[2][63] ), .Z(n2889) );
  XOR U8563 ( .A(\w0[2][57] ), .B(g_input[313]), .Z(\w1[2][57] ) );
  AND U8564 ( .A(\w1[2][56] ), .B(\SUBBYTES[2].a/w1822 ), .Z(
        \SUBBYTES[2].a/w1850 ) );
  XOR U8565 ( .A(\w0[2][56] ), .B(g_input[312]), .Z(\w1[2][56] ) );
  AND U8566 ( .A(\SUBBYTES[2].a/w1823 ), .B(\SUBBYTES[2].a/w1819 ), .Z(
        \SUBBYTES[2].a/w1848 ) );
  AND U8567 ( .A(\SUBBYTES[2].a/w1908 ), .B(\SUBBYTES[2].a/w1940 ), .Z(
        \SUBBYTES[2].a/w1847 ) );
  ANDN U8568 ( .A(\SUBBYTES[2].a/w1929 ), .B(n2893), .Z(\SUBBYTES[2].a/w1842 )
         );
  XNOR U8569 ( .A(\w1[2][60] ), .B(\w1[2][63] ), .Z(n2893) );
  ANDN U8570 ( .A(\SUBBYTES[2].a/w1930 ), .B(n2894), .Z(\SUBBYTES[2].a/w1840 )
         );
  XNOR U8571 ( .A(\w1[2][58] ), .B(\w1[2][63] ), .Z(n2894) );
  XOR U8572 ( .A(\w0[2][63] ), .B(g_input[319]), .Z(\w1[2][63] ) );
  IV U8573 ( .A(n2896), .Z(\w1[2][58] ) );
  ANDN U8574 ( .A(\SUBBYTES[2].a/w274 ), .B(n2853), .Z(\SUBBYTES[2].a/w184 )
         );
  XNOR U8575 ( .A(\w1[2][122] ), .B(\w1[2][127] ), .Z(n2853) );
  XOR U8576 ( .A(\w0[2][127] ), .B(g_input[383]), .Z(\w1[2][127] ) );
  IV U8577 ( .A(n2897), .Z(\w1[2][122] ) );
  ANDN U8578 ( .A(\SUBBYTES[2].a/w1932 ), .B(n2895), .Z(\SUBBYTES[2].a/w1839 )
         );
  XOR U8579 ( .A(n2896), .B(\w1[2][60] ), .Z(n2895) );
  XOR U8580 ( .A(\w0[2][60] ), .B(g_input[316]), .Z(\w1[2][60] ) );
  XNOR U8581 ( .A(\w0[2][58] ), .B(g_input[314]), .Z(n2896) );
  ANDN U8582 ( .A(\SUBBYTES[2].a/w276 ), .B(n2854), .Z(\SUBBYTES[2].a/w183 )
         );
  XOR U8583 ( .A(n2897), .B(\w1[2][124] ), .Z(n2854) );
  XOR U8584 ( .A(\w0[2][124] ), .B(g_input[380]), .Z(\w1[2][124] ) );
  XNOR U8585 ( .A(\w0[2][122] ), .B(g_input[378]), .Z(n2897) );
  AND U8586 ( .A(n2898), .B(\SUBBYTES[2].a/w1609 ), .Z(\SUBBYTES[2].a/w1744 )
         );
  AND U8587 ( .A(n2899), .B(\SUBBYTES[2].a/w1610 ), .Z(\SUBBYTES[2].a/w1742 )
         );
  AND U8588 ( .A(\SUBBYTES[2].a/w1740 ), .B(n2900), .Z(\SUBBYTES[2].a/w1741 )
         );
  ANDN U8589 ( .A(\w1[2][64] ), .B(n2901), .Z(\SUBBYTES[2].a/w1737 ) );
  AND U8590 ( .A(n2902), .B(\SUBBYTES[2].a/w1612 ), .Z(\SUBBYTES[2].a/w1735 )
         );
  AND U8591 ( .A(\SUBBYTES[2].a/w1733 ), .B(n2903), .Z(\SUBBYTES[2].a/w1734 )
         );
  XOR U8592 ( .A(\SUBBYTES[2].a/w1677 ), .B(n7126), .Z(n2903) );
  AND U8593 ( .A(\SUBBYTES[2].a/w1720 ), .B(\SUBBYTES[2].a/w1722 ), .Z(
        \SUBBYTES[2].a/w1729 ) );
  AND U8594 ( .A(\SUBBYTES[2].a/w1721 ), .B(\SUBBYTES[2].a/w1723 ), .Z(
        \SUBBYTES[2].a/w1727 ) );
  AND U8595 ( .A(\SUBBYTES[2].a/w1724 ), .B(\SUBBYTES[2].a/w1725 ), .Z(
        \SUBBYTES[2].a/w1726 ) );
  AND U8596 ( .A(\SUBBYTES[2].a/w1613 ), .B(n2898), .Z(\SUBBYTES[2].a/w1712 )
         );
  XOR U8597 ( .A(\SUBBYTES[2].a/w1681 ), .B(n980), .Z(n2898) );
  AND U8598 ( .A(\SUBBYTES[2].a/w1614 ), .B(n2899), .Z(\SUBBYTES[2].a/w1710 )
         );
  XOR U8599 ( .A(n7127), .B(\SUBBYTES[2].a/w1681 ), .Z(n2899) );
  ANDN U8600 ( .A(n2900), .B(n2904), .Z(\SUBBYTES[2].a/w1709 ) );
  XOR U8601 ( .A(n980), .B(n7127), .Z(n2900) );
  ANDN U8602 ( .A(\SUBBYTES[2].a/w1615 ), .B(n2901), .Z(\SUBBYTES[2].a/w1705 )
         );
  XNOR U8603 ( .A(\SUBBYTES[2].a/w1674 ), .B(\SUBBYTES[2].a/w1677 ), .Z(n2901)
         );
  AND U8604 ( .A(\SUBBYTES[2].a/w1616 ), .B(n2902), .Z(\SUBBYTES[2].a/w1703 )
         );
  XNOR U8605 ( .A(n2905), .B(\SUBBYTES[2].a/w1674 ), .Z(n2902) );
  AND U8606 ( .A(\SUBBYTES[2].a/w1701 ), .B(n2906), .Z(\SUBBYTES[2].a/w1702 )
         );
  XOR U8607 ( .A(n2907), .B(n2905), .Z(n2906) );
  IV U8608 ( .A(n7126), .Z(n2905) );
  ANDN U8609 ( .A(\SUBBYTES[2].a/w1720 ), .B(n2908), .Z(\SUBBYTES[2].a/w1697 )
         );
  ANDN U8610 ( .A(\SUBBYTES[2].a/w1721 ), .B(n2909), .Z(\SUBBYTES[2].a/w1695 )
         );
  ANDN U8611 ( .A(\SUBBYTES[2].a/w1724 ), .B(n2910), .Z(\SUBBYTES[2].a/w1694 )
         );
  AND U8612 ( .A(\SUBBYTES[2].a/w1680 ), .B(\SUBBYTES[2].a/w1679 ), .Z(
        \SUBBYTES[2].a/w1681 ) );
  IV U8613 ( .A(n2907), .Z(\SUBBYTES[2].a/w1677 ) );
  NAND U8614 ( .A(\SUBBYTES[2].a/w1656 ), .B(\SUBBYTES[2].a/w1671 ), .Z(n2907)
         );
  AND U8615 ( .A(\SUBBYTES[2].a/w1673 ), .B(\SUBBYTES[2].a/w1679 ), .Z(
        \SUBBYTES[2].a/w1674 ) );
  AND U8616 ( .A(\SUBBYTES[2].a/w1658 ), .B(\SUBBYTES[2].a/w1656 ), .Z(
        \SUBBYTES[2].a/w1668 ) );
  AND U8617 ( .A(\SUBBYTES[2].a/w1659 ), .B(\SUBBYTES[2].a/w1657 ), .Z(
        \SUBBYTES[2].a/w1666 ) );
  AND U8618 ( .A(\SUBBYTES[2].a/w1673 ), .B(\SUBBYTES[2].a/w1680 ), .Z(
        \SUBBYTES[2].a/w1665 ) );
  AND U8619 ( .A(\SUBBYTES[2].a/w1613 ), .B(\SUBBYTES[2].a/w1609 ), .Z(
        \SUBBYTES[2].a/w1650 ) );
  AND U8620 ( .A(\SUBBYTES[2].a/w1614 ), .B(\SUBBYTES[2].a/w1610 ), .Z(
        \SUBBYTES[2].a/w1648 ) );
  ANDN U8621 ( .A(\SUBBYTES[2].a/w1740 ), .B(n2904), .Z(\SUBBYTES[2].a/w1647 )
         );
  XNOR U8622 ( .A(\w1[2][65] ), .B(\w1[2][71] ), .Z(n2904) );
  XOR U8623 ( .A(\w0[2][65] ), .B(g_input[321]), .Z(\w1[2][65] ) );
  AND U8624 ( .A(\w1[2][64] ), .B(\SUBBYTES[2].a/w1615 ), .Z(
        \SUBBYTES[2].a/w1643 ) );
  XOR U8625 ( .A(\w0[2][64] ), .B(g_input[320]), .Z(\w1[2][64] ) );
  AND U8626 ( .A(\SUBBYTES[2].a/w1616 ), .B(\SUBBYTES[2].a/w1612 ), .Z(
        \SUBBYTES[2].a/w1641 ) );
  AND U8627 ( .A(\SUBBYTES[2].a/w1701 ), .B(\SUBBYTES[2].a/w1733 ), .Z(
        \SUBBYTES[2].a/w1640 ) );
  ANDN U8628 ( .A(\SUBBYTES[2].a/w1722 ), .B(n2908), .Z(\SUBBYTES[2].a/w1635 )
         );
  XNOR U8629 ( .A(\w1[2][68] ), .B(\w1[2][71] ), .Z(n2908) );
  ANDN U8630 ( .A(\SUBBYTES[2].a/w1723 ), .B(n2909), .Z(\SUBBYTES[2].a/w1633 )
         );
  XNOR U8631 ( .A(\w1[2][66] ), .B(\w1[2][71] ), .Z(n2909) );
  XOR U8632 ( .A(\w0[2][71] ), .B(g_input[327]), .Z(\w1[2][71] ) );
  IV U8633 ( .A(n2911), .Z(\w1[2][66] ) );
  ANDN U8634 ( .A(\SUBBYTES[2].a/w1725 ), .B(n2910), .Z(\SUBBYTES[2].a/w1632 )
         );
  XOR U8635 ( .A(n2911), .B(\w1[2][68] ), .Z(n2910) );
  XOR U8636 ( .A(\w0[2][68] ), .B(g_input[324]), .Z(\w1[2][68] ) );
  XNOR U8637 ( .A(\w0[2][66] ), .B(g_input[322]), .Z(n2911) );
  AND U8638 ( .A(n2912), .B(\SUBBYTES[2].a/w1402 ), .Z(\SUBBYTES[2].a/w1537 )
         );
  AND U8639 ( .A(n2913), .B(\SUBBYTES[2].a/w1403 ), .Z(\SUBBYTES[2].a/w1535 )
         );
  AND U8640 ( .A(\SUBBYTES[2].a/w1533 ), .B(n2914), .Z(\SUBBYTES[2].a/w1534 )
         );
  ANDN U8641 ( .A(\w1[2][72] ), .B(n2915), .Z(\SUBBYTES[2].a/w1530 ) );
  AND U8642 ( .A(n2916), .B(\SUBBYTES[2].a/w1405 ), .Z(\SUBBYTES[2].a/w1528 )
         );
  AND U8643 ( .A(\SUBBYTES[2].a/w1526 ), .B(n2917), .Z(\SUBBYTES[2].a/w1527 )
         );
  XOR U8644 ( .A(\SUBBYTES[2].a/w1470 ), .B(n7124), .Z(n2917) );
  AND U8645 ( .A(\SUBBYTES[2].a/w1513 ), .B(\SUBBYTES[2].a/w1515 ), .Z(
        \SUBBYTES[2].a/w1522 ) );
  AND U8646 ( .A(\SUBBYTES[2].a/w1514 ), .B(\SUBBYTES[2].a/w1516 ), .Z(
        \SUBBYTES[2].a/w1520 ) );
  AND U8647 ( .A(\SUBBYTES[2].a/w1517 ), .B(\SUBBYTES[2].a/w1518 ), .Z(
        \SUBBYTES[2].a/w1519 ) );
  AND U8648 ( .A(\SUBBYTES[2].a/w1406 ), .B(n2912), .Z(\SUBBYTES[2].a/w1505 )
         );
  XOR U8649 ( .A(\SUBBYTES[2].a/w1474 ), .B(n979), .Z(n2912) );
  AND U8650 ( .A(\SUBBYTES[2].a/w1407 ), .B(n2913), .Z(\SUBBYTES[2].a/w1503 )
         );
  XOR U8651 ( .A(n7125), .B(\SUBBYTES[2].a/w1474 ), .Z(n2913) );
  ANDN U8652 ( .A(n2914), .B(n2918), .Z(\SUBBYTES[2].a/w1502 ) );
  XOR U8653 ( .A(n979), .B(n7125), .Z(n2914) );
  ANDN U8654 ( .A(\SUBBYTES[2].a/w1408 ), .B(n2915), .Z(\SUBBYTES[2].a/w1498 )
         );
  XNOR U8655 ( .A(\SUBBYTES[2].a/w1467 ), .B(\SUBBYTES[2].a/w1470 ), .Z(n2915)
         );
  AND U8656 ( .A(\SUBBYTES[2].a/w1409 ), .B(n2916), .Z(\SUBBYTES[2].a/w1496 )
         );
  XNOR U8657 ( .A(n2919), .B(\SUBBYTES[2].a/w1467 ), .Z(n2916) );
  AND U8658 ( .A(\SUBBYTES[2].a/w1494 ), .B(n2920), .Z(\SUBBYTES[2].a/w1495 )
         );
  XOR U8659 ( .A(n2921), .B(n2919), .Z(n2920) );
  IV U8660 ( .A(n7124), .Z(n2919) );
  ANDN U8661 ( .A(\SUBBYTES[2].a/w1513 ), .B(n2922), .Z(\SUBBYTES[2].a/w1490 )
         );
  ANDN U8662 ( .A(\SUBBYTES[2].a/w1514 ), .B(n2923), .Z(\SUBBYTES[2].a/w1488 )
         );
  ANDN U8663 ( .A(\SUBBYTES[2].a/w1517 ), .B(n2924), .Z(\SUBBYTES[2].a/w1487 )
         );
  AND U8664 ( .A(\SUBBYTES[2].a/w1473 ), .B(\SUBBYTES[2].a/w1472 ), .Z(
        \SUBBYTES[2].a/w1474 ) );
  IV U8665 ( .A(n2921), .Z(\SUBBYTES[2].a/w1470 ) );
  NAND U8666 ( .A(\SUBBYTES[2].a/w1449 ), .B(\SUBBYTES[2].a/w1464 ), .Z(n2921)
         );
  AND U8667 ( .A(\SUBBYTES[2].a/w1466 ), .B(\SUBBYTES[2].a/w1472 ), .Z(
        \SUBBYTES[2].a/w1467 ) );
  AND U8668 ( .A(\SUBBYTES[2].a/w1451 ), .B(\SUBBYTES[2].a/w1449 ), .Z(
        \SUBBYTES[2].a/w1461 ) );
  AND U8669 ( .A(\SUBBYTES[2].a/w1452 ), .B(\SUBBYTES[2].a/w1450 ), .Z(
        \SUBBYTES[2].a/w1459 ) );
  AND U8670 ( .A(\SUBBYTES[2].a/w1466 ), .B(\SUBBYTES[2].a/w1473 ), .Z(
        \SUBBYTES[2].a/w1458 ) );
  AND U8671 ( .A(\SUBBYTES[2].a/w1406 ), .B(\SUBBYTES[2].a/w1402 ), .Z(
        \SUBBYTES[2].a/w1443 ) );
  AND U8672 ( .A(\SUBBYTES[2].a/w1407 ), .B(\SUBBYTES[2].a/w1403 ), .Z(
        \SUBBYTES[2].a/w1441 ) );
  ANDN U8673 ( .A(\SUBBYTES[2].a/w1533 ), .B(n2918), .Z(\SUBBYTES[2].a/w1440 )
         );
  XNOR U8674 ( .A(\w1[2][73] ), .B(\w1[2][79] ), .Z(n2918) );
  XOR U8675 ( .A(\w0[2][73] ), .B(g_input[329]), .Z(\w1[2][73] ) );
  AND U8676 ( .A(\w1[2][72] ), .B(\SUBBYTES[2].a/w1408 ), .Z(
        \SUBBYTES[2].a/w1436 ) );
  XOR U8677 ( .A(\w0[2][72] ), .B(g_input[328]), .Z(\w1[2][72] ) );
  AND U8678 ( .A(\SUBBYTES[2].a/w1409 ), .B(\SUBBYTES[2].a/w1405 ), .Z(
        \SUBBYTES[2].a/w1434 ) );
  AND U8679 ( .A(\SUBBYTES[2].a/w1494 ), .B(\SUBBYTES[2].a/w1526 ), .Z(
        \SUBBYTES[2].a/w1433 ) );
  ANDN U8680 ( .A(\SUBBYTES[2].a/w1515 ), .B(n2922), .Z(\SUBBYTES[2].a/w1428 )
         );
  XNOR U8681 ( .A(\w1[2][76] ), .B(\w1[2][79] ), .Z(n2922) );
  ANDN U8682 ( .A(\SUBBYTES[2].a/w1516 ), .B(n2923), .Z(\SUBBYTES[2].a/w1426 )
         );
  XNOR U8683 ( .A(\w1[2][74] ), .B(\w1[2][79] ), .Z(n2923) );
  XOR U8684 ( .A(\w0[2][79] ), .B(g_input[335]), .Z(\w1[2][79] ) );
  IV U8685 ( .A(n2925), .Z(\w1[2][74] ) );
  ANDN U8686 ( .A(\SUBBYTES[2].a/w1518 ), .B(n2924), .Z(\SUBBYTES[2].a/w1425 )
         );
  XOR U8687 ( .A(n2925), .B(\w1[2][76] ), .Z(n2924) );
  XOR U8688 ( .A(\w0[2][76] ), .B(g_input[332]), .Z(\w1[2][76] ) );
  XNOR U8689 ( .A(\w0[2][74] ), .B(g_input[330]), .Z(n2925) );
  AND U8690 ( .A(n2926), .B(\SUBBYTES[2].a/w1195 ), .Z(\SUBBYTES[2].a/w1330 )
         );
  AND U8691 ( .A(n2927), .B(\SUBBYTES[2].a/w1196 ), .Z(\SUBBYTES[2].a/w1328 )
         );
  AND U8692 ( .A(\SUBBYTES[2].a/w1326 ), .B(n2928), .Z(\SUBBYTES[2].a/w1327 )
         );
  ANDN U8693 ( .A(\w1[2][80] ), .B(n2929), .Z(\SUBBYTES[2].a/w1323 ) );
  AND U8694 ( .A(n2930), .B(\SUBBYTES[2].a/w1198 ), .Z(\SUBBYTES[2].a/w1321 )
         );
  AND U8695 ( .A(\SUBBYTES[2].a/w1319 ), .B(n2931), .Z(\SUBBYTES[2].a/w1320 )
         );
  XOR U8696 ( .A(\SUBBYTES[2].a/w1263 ), .B(n7122), .Z(n2931) );
  AND U8697 ( .A(\SUBBYTES[2].a/w1306 ), .B(\SUBBYTES[2].a/w1308 ), .Z(
        \SUBBYTES[2].a/w1315 ) );
  AND U8698 ( .A(\SUBBYTES[2].a/w1307 ), .B(\SUBBYTES[2].a/w1309 ), .Z(
        \SUBBYTES[2].a/w1313 ) );
  AND U8699 ( .A(\SUBBYTES[2].a/w1310 ), .B(\SUBBYTES[2].a/w1311 ), .Z(
        \SUBBYTES[2].a/w1312 ) );
  AND U8700 ( .A(\SUBBYTES[2].a/w1199 ), .B(n2926), .Z(\SUBBYTES[2].a/w1298 )
         );
  XOR U8701 ( .A(\SUBBYTES[2].a/w1267 ), .B(n978), .Z(n2926) );
  AND U8702 ( .A(\SUBBYTES[2].a/w1200 ), .B(n2927), .Z(\SUBBYTES[2].a/w1296 )
         );
  XOR U8703 ( .A(n7123), .B(\SUBBYTES[2].a/w1267 ), .Z(n2927) );
  ANDN U8704 ( .A(n2928), .B(n2932), .Z(\SUBBYTES[2].a/w1295 ) );
  XOR U8705 ( .A(n978), .B(n7123), .Z(n2928) );
  ANDN U8706 ( .A(\SUBBYTES[2].a/w1201 ), .B(n2929), .Z(\SUBBYTES[2].a/w1291 )
         );
  XNOR U8707 ( .A(\SUBBYTES[2].a/w1260 ), .B(\SUBBYTES[2].a/w1263 ), .Z(n2929)
         );
  AND U8708 ( .A(\SUBBYTES[2].a/w1202 ), .B(n2930), .Z(\SUBBYTES[2].a/w1289 )
         );
  XNOR U8709 ( .A(n2933), .B(\SUBBYTES[2].a/w1260 ), .Z(n2930) );
  AND U8710 ( .A(\SUBBYTES[2].a/w1287 ), .B(n2934), .Z(\SUBBYTES[2].a/w1288 )
         );
  XOR U8711 ( .A(n2935), .B(n2933), .Z(n2934) );
  IV U8712 ( .A(n7122), .Z(n2933) );
  ANDN U8713 ( .A(\SUBBYTES[2].a/w1306 ), .B(n2936), .Z(\SUBBYTES[2].a/w1283 )
         );
  ANDN U8714 ( .A(\SUBBYTES[2].a/w1307 ), .B(n2937), .Z(\SUBBYTES[2].a/w1281 )
         );
  ANDN U8715 ( .A(\SUBBYTES[2].a/w1310 ), .B(n2938), .Z(\SUBBYTES[2].a/w1280 )
         );
  AND U8716 ( .A(\SUBBYTES[2].a/w1266 ), .B(\SUBBYTES[2].a/w1265 ), .Z(
        \SUBBYTES[2].a/w1267 ) );
  IV U8717 ( .A(n2935), .Z(\SUBBYTES[2].a/w1263 ) );
  NAND U8718 ( .A(\SUBBYTES[2].a/w1242 ), .B(\SUBBYTES[2].a/w1257 ), .Z(n2935)
         );
  AND U8719 ( .A(\SUBBYTES[2].a/w1259 ), .B(\SUBBYTES[2].a/w1265 ), .Z(
        \SUBBYTES[2].a/w1260 ) );
  AND U8720 ( .A(\SUBBYTES[2].a/w1244 ), .B(\SUBBYTES[2].a/w1242 ), .Z(
        \SUBBYTES[2].a/w1254 ) );
  AND U8721 ( .A(\SUBBYTES[2].a/w1245 ), .B(\SUBBYTES[2].a/w1243 ), .Z(
        \SUBBYTES[2].a/w1252 ) );
  AND U8722 ( .A(\SUBBYTES[2].a/w1259 ), .B(\SUBBYTES[2].a/w1266 ), .Z(
        \SUBBYTES[2].a/w1251 ) );
  AND U8723 ( .A(\SUBBYTES[2].a/w1199 ), .B(\SUBBYTES[2].a/w1195 ), .Z(
        \SUBBYTES[2].a/w1236 ) );
  AND U8724 ( .A(\SUBBYTES[2].a/w1200 ), .B(\SUBBYTES[2].a/w1196 ), .Z(
        \SUBBYTES[2].a/w1234 ) );
  ANDN U8725 ( .A(\SUBBYTES[2].a/w1326 ), .B(n2932), .Z(\SUBBYTES[2].a/w1233 )
         );
  XNOR U8726 ( .A(\w1[2][81] ), .B(\w1[2][87] ), .Z(n2932) );
  XOR U8727 ( .A(\w0[2][81] ), .B(g_input[337]), .Z(\w1[2][81] ) );
  AND U8728 ( .A(\w1[2][80] ), .B(\SUBBYTES[2].a/w1201 ), .Z(
        \SUBBYTES[2].a/w1229 ) );
  XOR U8729 ( .A(\w0[2][80] ), .B(g_input[336]), .Z(\w1[2][80] ) );
  AND U8730 ( .A(\SUBBYTES[2].a/w1202 ), .B(\SUBBYTES[2].a/w1198 ), .Z(
        \SUBBYTES[2].a/w1227 ) );
  AND U8731 ( .A(\SUBBYTES[2].a/w1287 ), .B(\SUBBYTES[2].a/w1319 ), .Z(
        \SUBBYTES[2].a/w1226 ) );
  ANDN U8732 ( .A(\SUBBYTES[2].a/w1308 ), .B(n2936), .Z(\SUBBYTES[2].a/w1221 )
         );
  XNOR U8733 ( .A(\w1[2][84] ), .B(\w1[2][87] ), .Z(n2936) );
  ANDN U8734 ( .A(\SUBBYTES[2].a/w1309 ), .B(n2937), .Z(\SUBBYTES[2].a/w1219 )
         );
  XNOR U8735 ( .A(\w1[2][82] ), .B(\w1[2][87] ), .Z(n2937) );
  XOR U8736 ( .A(\w0[2][87] ), .B(g_input[343]), .Z(\w1[2][87] ) );
  IV U8737 ( .A(n2939), .Z(\w1[2][82] ) );
  ANDN U8738 ( .A(\SUBBYTES[2].a/w1311 ), .B(n2938), .Z(\SUBBYTES[2].a/w1218 )
         );
  XOR U8739 ( .A(n2939), .B(\w1[2][84] ), .Z(n2938) );
  XOR U8740 ( .A(\w0[2][84] ), .B(g_input[340]), .Z(\w1[2][84] ) );
  XNOR U8741 ( .A(\w0[2][82] ), .B(g_input[338]), .Z(n2939) );
  AND U8742 ( .A(n2940), .B(\SUBBYTES[2].a/w988 ), .Z(\SUBBYTES[2].a/w1123 )
         );
  AND U8743 ( .A(n2941), .B(\SUBBYTES[2].a/w989 ), .Z(\SUBBYTES[2].a/w1121 )
         );
  AND U8744 ( .A(\SUBBYTES[2].a/w1119 ), .B(n2942), .Z(\SUBBYTES[2].a/w1120 )
         );
  ANDN U8745 ( .A(\w1[2][88] ), .B(n2943), .Z(\SUBBYTES[2].a/w1116 ) );
  AND U8746 ( .A(n2944), .B(\SUBBYTES[2].a/w991 ), .Z(\SUBBYTES[2].a/w1114 )
         );
  AND U8747 ( .A(\SUBBYTES[2].a/w1112 ), .B(n2945), .Z(\SUBBYTES[2].a/w1113 )
         );
  XOR U8748 ( .A(\SUBBYTES[2].a/w1056 ), .B(n7120), .Z(n2945) );
  AND U8749 ( .A(\SUBBYTES[2].a/w1099 ), .B(\SUBBYTES[2].a/w1101 ), .Z(
        \SUBBYTES[2].a/w1108 ) );
  AND U8750 ( .A(\SUBBYTES[2].a/w1100 ), .B(\SUBBYTES[2].a/w1102 ), .Z(
        \SUBBYTES[2].a/w1106 ) );
  AND U8751 ( .A(\SUBBYTES[2].a/w1103 ), .B(\SUBBYTES[2].a/w1104 ), .Z(
        \SUBBYTES[2].a/w1105 ) );
  AND U8752 ( .A(\SUBBYTES[2].a/w992 ), .B(n2940), .Z(\SUBBYTES[2].a/w1091 )
         );
  XOR U8753 ( .A(\SUBBYTES[2].a/w1060 ), .B(n977), .Z(n2940) );
  AND U8754 ( .A(\SUBBYTES[2].a/w993 ), .B(n2941), .Z(\SUBBYTES[2].a/w1089 )
         );
  XOR U8755 ( .A(n7121), .B(\SUBBYTES[2].a/w1060 ), .Z(n2941) );
  ANDN U8756 ( .A(n2942), .B(n2946), .Z(\SUBBYTES[2].a/w1088 ) );
  XOR U8757 ( .A(n977), .B(n7121), .Z(n2942) );
  ANDN U8758 ( .A(\SUBBYTES[2].a/w994 ), .B(n2943), .Z(\SUBBYTES[2].a/w1084 )
         );
  XNOR U8759 ( .A(\SUBBYTES[2].a/w1053 ), .B(\SUBBYTES[2].a/w1056 ), .Z(n2943)
         );
  AND U8760 ( .A(\SUBBYTES[2].a/w995 ), .B(n2944), .Z(\SUBBYTES[2].a/w1082 )
         );
  XNOR U8761 ( .A(n2947), .B(\SUBBYTES[2].a/w1053 ), .Z(n2944) );
  AND U8762 ( .A(\SUBBYTES[2].a/w1080 ), .B(n2948), .Z(\SUBBYTES[2].a/w1081 )
         );
  XOR U8763 ( .A(n2949), .B(n2947), .Z(n2948) );
  IV U8764 ( .A(n7120), .Z(n2947) );
  ANDN U8765 ( .A(\SUBBYTES[2].a/w1099 ), .B(n2950), .Z(\SUBBYTES[2].a/w1076 )
         );
  ANDN U8766 ( .A(\SUBBYTES[2].a/w1100 ), .B(n2951), .Z(\SUBBYTES[2].a/w1074 )
         );
  ANDN U8767 ( .A(\SUBBYTES[2].a/w1103 ), .B(n2952), .Z(\SUBBYTES[2].a/w1073 )
         );
  AND U8768 ( .A(\SUBBYTES[2].a/w1059 ), .B(\SUBBYTES[2].a/w1058 ), .Z(
        \SUBBYTES[2].a/w1060 ) );
  IV U8769 ( .A(n2949), .Z(\SUBBYTES[2].a/w1056 ) );
  NAND U8770 ( .A(\SUBBYTES[2].a/w1035 ), .B(\SUBBYTES[2].a/w1050 ), .Z(n2949)
         );
  AND U8771 ( .A(\SUBBYTES[2].a/w1052 ), .B(\SUBBYTES[2].a/w1058 ), .Z(
        \SUBBYTES[2].a/w1053 ) );
  AND U8772 ( .A(\SUBBYTES[2].a/w1037 ), .B(\SUBBYTES[2].a/w1035 ), .Z(
        \SUBBYTES[2].a/w1047 ) );
  AND U8773 ( .A(\SUBBYTES[2].a/w1038 ), .B(\SUBBYTES[2].a/w1036 ), .Z(
        \SUBBYTES[2].a/w1045 ) );
  AND U8774 ( .A(\SUBBYTES[2].a/w1052 ), .B(\SUBBYTES[2].a/w1059 ), .Z(
        \SUBBYTES[2].a/w1044 ) );
  AND U8775 ( .A(\SUBBYTES[2].a/w992 ), .B(\SUBBYTES[2].a/w988 ), .Z(
        \SUBBYTES[2].a/w1029 ) );
  AND U8776 ( .A(\SUBBYTES[2].a/w993 ), .B(\SUBBYTES[2].a/w989 ), .Z(
        \SUBBYTES[2].a/w1027 ) );
  ANDN U8777 ( .A(\SUBBYTES[2].a/w1119 ), .B(n2946), .Z(\SUBBYTES[2].a/w1026 )
         );
  XNOR U8778 ( .A(\w1[2][89] ), .B(\w1[2][95] ), .Z(n2946) );
  XOR U8779 ( .A(\w0[2][89] ), .B(g_input[345]), .Z(\w1[2][89] ) );
  AND U8780 ( .A(\w1[2][88] ), .B(\SUBBYTES[2].a/w994 ), .Z(
        \SUBBYTES[2].a/w1022 ) );
  XOR U8781 ( .A(\w0[2][88] ), .B(g_input[344]), .Z(\w1[2][88] ) );
  AND U8782 ( .A(\SUBBYTES[2].a/w995 ), .B(\SUBBYTES[2].a/w991 ), .Z(
        \SUBBYTES[2].a/w1020 ) );
  AND U8783 ( .A(\SUBBYTES[2].a/w1080 ), .B(\SUBBYTES[2].a/w1112 ), .Z(
        \SUBBYTES[2].a/w1019 ) );
  ANDN U8784 ( .A(\SUBBYTES[2].a/w1101 ), .B(n2950), .Z(\SUBBYTES[2].a/w1014 )
         );
  XNOR U8785 ( .A(\w1[2][92] ), .B(\w1[2][95] ), .Z(n2950) );
  ANDN U8786 ( .A(\SUBBYTES[2].a/w1102 ), .B(n2951), .Z(\SUBBYTES[2].a/w1012 )
         );
  XNOR U8787 ( .A(\w1[2][90] ), .B(\w1[2][95] ), .Z(n2951) );
  XOR U8788 ( .A(\w0[2][95] ), .B(g_input[351]), .Z(\w1[2][95] ) );
  IV U8789 ( .A(n2953), .Z(\w1[2][90] ) );
  ANDN U8790 ( .A(\SUBBYTES[2].a/w1104 ), .B(n2952), .Z(\SUBBYTES[2].a/w1011 )
         );
  XOR U8791 ( .A(n2953), .B(\w1[2][92] ), .Z(n2952) );
  XOR U8792 ( .A(\w0[2][92] ), .B(g_input[348]), .Z(\w1[2][92] ) );
  XNOR U8793 ( .A(\w0[2][90] ), .B(g_input[346]), .Z(n2953) );
  AND U8794 ( .A(\SUBBYTES[2].a/w2084 ), .B(\SUBBYTES[2].a/w2071 ), .Z(n7130)
         );
  AND U8795 ( .A(\SUBBYTES[2].a/w1877 ), .B(\SUBBYTES[2].a/w1866 ), .Z(n7129)
         );
  AND U8796 ( .A(\SUBBYTES[2].a/w221 ), .B(\SUBBYTES[2].a/w208 ), .Z(n7112) );
  AND U8797 ( .A(\SUBBYTES[2].a/w1877 ), .B(\SUBBYTES[2].a/w1864 ), .Z(n7128)
         );
  AND U8798 ( .A(\SUBBYTES[2].a/w1670 ), .B(\SUBBYTES[2].a/w1659 ), .Z(n7127)
         );
  AND U8799 ( .A(\SUBBYTES[2].a/w1670 ), .B(\SUBBYTES[2].a/w1657 ), .Z(n7126)
         );
  AND U8800 ( .A(\SUBBYTES[2].a/w1463 ), .B(\SUBBYTES[2].a/w1452 ), .Z(n7125)
         );
  AND U8801 ( .A(\SUBBYTES[2].a/w1463 ), .B(\SUBBYTES[2].a/w1450 ), .Z(n7124)
         );
  AND U8802 ( .A(\SUBBYTES[2].a/w1256 ), .B(\SUBBYTES[2].a/w1245 ), .Z(n7123)
         );
  AND U8803 ( .A(\SUBBYTES[2].a/w1256 ), .B(\SUBBYTES[2].a/w1243 ), .Z(n7122)
         );
  AND U8804 ( .A(\SUBBYTES[2].a/w1049 ), .B(\SUBBYTES[2].a/w1038 ), .Z(n7121)
         );
  AND U8805 ( .A(\SUBBYTES[2].a/w1049 ), .B(\SUBBYTES[2].a/w1036 ), .Z(n7120)
         );
  AND U8806 ( .A(\SUBBYTES[2].a/w842 ), .B(\SUBBYTES[2].a/w831 ), .Z(n7119) );
  AND U8807 ( .A(\SUBBYTES[2].a/w842 ), .B(\SUBBYTES[2].a/w829 ), .Z(n7118) );
  AND U8808 ( .A(\SUBBYTES[2].a/w635 ), .B(\SUBBYTES[2].a/w624 ), .Z(n7117) );
  AND U8809 ( .A(\SUBBYTES[2].a/w635 ), .B(\SUBBYTES[2].a/w622 ), .Z(n7116) );
  AND U8810 ( .A(\SUBBYTES[2].a/w428 ), .B(\SUBBYTES[2].a/w417 ), .Z(n7115) );
  AND U8811 ( .A(\SUBBYTES[2].a/w428 ), .B(\SUBBYTES[2].a/w415 ), .Z(n7114) );
  AND U8812 ( .A(\SUBBYTES[2].a/w3326 ), .B(\SUBBYTES[2].a/w3315 ), .Z(n7143)
         );
  AND U8813 ( .A(\SUBBYTES[2].a/w3326 ), .B(\SUBBYTES[2].a/w3313 ), .Z(n7142)
         );
  AND U8814 ( .A(\SUBBYTES[2].a/w3119 ), .B(\SUBBYTES[2].a/w3108 ), .Z(n7141)
         );
  AND U8815 ( .A(\SUBBYTES[2].a/w3119 ), .B(\SUBBYTES[2].a/w3106 ), .Z(n7140)
         );
  AND U8816 ( .A(\SUBBYTES[2].a/w2912 ), .B(\SUBBYTES[2].a/w2901 ), .Z(n7139)
         );
  AND U8817 ( .A(\SUBBYTES[2].a/w2912 ), .B(\SUBBYTES[2].a/w2899 ), .Z(n7138)
         );
  AND U8818 ( .A(\SUBBYTES[2].a/w2705 ), .B(\SUBBYTES[2].a/w2694 ), .Z(n7137)
         );
  AND U8819 ( .A(\SUBBYTES[2].a/w2705 ), .B(\SUBBYTES[2].a/w2692 ), .Z(n7136)
         );
  AND U8820 ( .A(\SUBBYTES[2].a/w2498 ), .B(\SUBBYTES[2].a/w2487 ), .Z(n7135)
         );
  AND U8821 ( .A(\SUBBYTES[2].a/w2498 ), .B(\SUBBYTES[2].a/w2485 ), .Z(n7134)
         );
  AND U8822 ( .A(\SUBBYTES[2].a/w2291 ), .B(\SUBBYTES[2].a/w2280 ), .Z(n7133)
         );
  AND U8823 ( .A(\SUBBYTES[2].a/w2291 ), .B(\SUBBYTES[2].a/w2278 ), .Z(n7132)
         );
  AND U8824 ( .A(\SUBBYTES[2].a/w2084 ), .B(\SUBBYTES[2].a/w2073 ), .Z(n7131)
         );
  AND U8825 ( .A(\SUBBYTES[2].a/w221 ), .B(\SUBBYTES[2].a/w210 ), .Z(n7113) );
  AND U8826 ( .A(n2954), .B(\SUBBYTES[1].a/w781 ), .Z(\SUBBYTES[1].a/w916 ) );
  AND U8827 ( .A(n2955), .B(\SUBBYTES[1].a/w782 ), .Z(\SUBBYTES[1].a/w914 ) );
  AND U8828 ( .A(\SUBBYTES[1].a/w912 ), .B(n2956), .Z(\SUBBYTES[1].a/w913 ) );
  ANDN U8829 ( .A(\w1[1][96] ), .B(n2957), .Z(\SUBBYTES[1].a/w909 ) );
  AND U8830 ( .A(n2958), .B(\SUBBYTES[1].a/w784 ), .Z(\SUBBYTES[1].a/w907 ) );
  AND U8831 ( .A(\SUBBYTES[1].a/w905 ), .B(n2959), .Z(\SUBBYTES[1].a/w906 ) );
  XOR U8832 ( .A(\SUBBYTES[1].a/w849 ), .B(n5838), .Z(n2959) );
  AND U8833 ( .A(\SUBBYTES[1].a/w892 ), .B(\SUBBYTES[1].a/w894 ), .Z(
        \SUBBYTES[1].a/w901 ) );
  AND U8834 ( .A(\SUBBYTES[1].a/w893 ), .B(\SUBBYTES[1].a/w895 ), .Z(
        \SUBBYTES[1].a/w899 ) );
  AND U8835 ( .A(\SUBBYTES[1].a/w896 ), .B(\SUBBYTES[1].a/w897 ), .Z(
        \SUBBYTES[1].a/w898 ) );
  AND U8836 ( .A(\SUBBYTES[1].a/w785 ), .B(n2954), .Z(\SUBBYTES[1].a/w884 ) );
  XOR U8837 ( .A(\SUBBYTES[1].a/w853 ), .B(n960), .Z(n2954) );
  AND U8838 ( .A(\SUBBYTES[1].a/w786 ), .B(n2955), .Z(\SUBBYTES[1].a/w882 ) );
  XOR U8839 ( .A(n5839), .B(\SUBBYTES[1].a/w853 ), .Z(n2955) );
  ANDN U8840 ( .A(n2956), .B(n2960), .Z(\SUBBYTES[1].a/w881 ) );
  XOR U8841 ( .A(n960), .B(n5839), .Z(n2956) );
  ANDN U8842 ( .A(\SUBBYTES[1].a/w787 ), .B(n2957), .Z(\SUBBYTES[1].a/w877 )
         );
  XNOR U8843 ( .A(\SUBBYTES[1].a/w846 ), .B(\SUBBYTES[1].a/w849 ), .Z(n2957)
         );
  AND U8844 ( .A(\SUBBYTES[1].a/w788 ), .B(n2958), .Z(\SUBBYTES[1].a/w875 ) );
  XNOR U8845 ( .A(n2961), .B(\SUBBYTES[1].a/w846 ), .Z(n2958) );
  AND U8846 ( .A(\SUBBYTES[1].a/w873 ), .B(n2962), .Z(\SUBBYTES[1].a/w874 ) );
  XOR U8847 ( .A(n2963), .B(n2961), .Z(n2962) );
  IV U8848 ( .A(n5838), .Z(n2961) );
  ANDN U8849 ( .A(\SUBBYTES[1].a/w892 ), .B(n2964), .Z(\SUBBYTES[1].a/w869 )
         );
  ANDN U8850 ( .A(\SUBBYTES[1].a/w893 ), .B(n2965), .Z(\SUBBYTES[1].a/w867 )
         );
  ANDN U8851 ( .A(\SUBBYTES[1].a/w896 ), .B(n2966), .Z(\SUBBYTES[1].a/w866 )
         );
  AND U8852 ( .A(\SUBBYTES[1].a/w852 ), .B(\SUBBYTES[1].a/w851 ), .Z(
        \SUBBYTES[1].a/w853 ) );
  IV U8853 ( .A(n2963), .Z(\SUBBYTES[1].a/w849 ) );
  NAND U8854 ( .A(\SUBBYTES[1].a/w828 ), .B(\SUBBYTES[1].a/w843 ), .Z(n2963)
         );
  AND U8855 ( .A(\SUBBYTES[1].a/w845 ), .B(\SUBBYTES[1].a/w851 ), .Z(
        \SUBBYTES[1].a/w846 ) );
  AND U8856 ( .A(\SUBBYTES[1].a/w830 ), .B(\SUBBYTES[1].a/w828 ), .Z(
        \SUBBYTES[1].a/w840 ) );
  AND U8857 ( .A(\SUBBYTES[1].a/w831 ), .B(\SUBBYTES[1].a/w829 ), .Z(
        \SUBBYTES[1].a/w838 ) );
  AND U8858 ( .A(\SUBBYTES[1].a/w845 ), .B(\SUBBYTES[1].a/w852 ), .Z(
        \SUBBYTES[1].a/w837 ) );
  AND U8859 ( .A(\SUBBYTES[1].a/w785 ), .B(\SUBBYTES[1].a/w781 ), .Z(
        \SUBBYTES[1].a/w822 ) );
  AND U8860 ( .A(\SUBBYTES[1].a/w786 ), .B(\SUBBYTES[1].a/w782 ), .Z(
        \SUBBYTES[1].a/w820 ) );
  ANDN U8861 ( .A(\SUBBYTES[1].a/w912 ), .B(n2960), .Z(\SUBBYTES[1].a/w819 )
         );
  XNOR U8862 ( .A(\w1[1][103] ), .B(\w1[1][97] ), .Z(n2960) );
  XOR U8863 ( .A(\w0[1][97] ), .B(g_input[225]), .Z(\w1[1][97] ) );
  IV U8864 ( .A(n2967), .Z(\w1[1][103] ) );
  AND U8865 ( .A(\w1[1][96] ), .B(\SUBBYTES[1].a/w787 ), .Z(
        \SUBBYTES[1].a/w815 ) );
  XOR U8866 ( .A(\w0[1][96] ), .B(g_input[224]), .Z(\w1[1][96] ) );
  AND U8867 ( .A(\SUBBYTES[1].a/w788 ), .B(\SUBBYTES[1].a/w784 ), .Z(
        \SUBBYTES[1].a/w813 ) );
  AND U8868 ( .A(\SUBBYTES[1].a/w873 ), .B(\SUBBYTES[1].a/w905 ), .Z(
        \SUBBYTES[1].a/w812 ) );
  ANDN U8869 ( .A(\SUBBYTES[1].a/w894 ), .B(n2964), .Z(\SUBBYTES[1].a/w807 )
         );
  XOR U8870 ( .A(\w1[1][100] ), .B(n2967), .Z(n2964) );
  ANDN U8871 ( .A(\SUBBYTES[1].a/w895 ), .B(n2965), .Z(\SUBBYTES[1].a/w805 )
         );
  XOR U8872 ( .A(n2967), .B(\w1[1][98] ), .Z(n2965) );
  XNOR U8873 ( .A(\w0[1][103] ), .B(g_input[231]), .Z(n2967) );
  ANDN U8874 ( .A(\SUBBYTES[1].a/w897 ), .B(n2966), .Z(\SUBBYTES[1].a/w804 )
         );
  XNOR U8875 ( .A(\w1[1][100] ), .B(\w1[1][98] ), .Z(n2966) );
  XOR U8876 ( .A(\w0[1][98] ), .B(g_input[226]), .Z(\w1[1][98] ) );
  XOR U8877 ( .A(\w0[1][100] ), .B(g_input[228]), .Z(\w1[1][100] ) );
  AND U8878 ( .A(n2968), .B(\SUBBYTES[1].a/w574 ), .Z(\SUBBYTES[1].a/w709 ) );
  AND U8879 ( .A(n2969), .B(\SUBBYTES[1].a/w575 ), .Z(\SUBBYTES[1].a/w707 ) );
  AND U8880 ( .A(\SUBBYTES[1].a/w705 ), .B(n2970), .Z(\SUBBYTES[1].a/w706 ) );
  ANDN U8881 ( .A(\w1[1][104] ), .B(n2971), .Z(\SUBBYTES[1].a/w702 ) );
  AND U8882 ( .A(n2972), .B(\SUBBYTES[1].a/w577 ), .Z(\SUBBYTES[1].a/w700 ) );
  AND U8883 ( .A(\SUBBYTES[1].a/w698 ), .B(n2973), .Z(\SUBBYTES[1].a/w699 ) );
  XOR U8884 ( .A(\SUBBYTES[1].a/w642 ), .B(n5836), .Z(n2973) );
  AND U8885 ( .A(\SUBBYTES[1].a/w685 ), .B(\SUBBYTES[1].a/w687 ), .Z(
        \SUBBYTES[1].a/w694 ) );
  AND U8886 ( .A(\SUBBYTES[1].a/w686 ), .B(\SUBBYTES[1].a/w688 ), .Z(
        \SUBBYTES[1].a/w692 ) );
  AND U8887 ( .A(\SUBBYTES[1].a/w689 ), .B(\SUBBYTES[1].a/w690 ), .Z(
        \SUBBYTES[1].a/w691 ) );
  AND U8888 ( .A(\SUBBYTES[1].a/w578 ), .B(n2968), .Z(\SUBBYTES[1].a/w677 ) );
  XOR U8889 ( .A(\SUBBYTES[1].a/w646 ), .B(n959), .Z(n2968) );
  AND U8890 ( .A(\SUBBYTES[1].a/w579 ), .B(n2969), .Z(\SUBBYTES[1].a/w675 ) );
  XOR U8891 ( .A(n5837), .B(\SUBBYTES[1].a/w646 ), .Z(n2969) );
  ANDN U8892 ( .A(n2970), .B(n2974), .Z(\SUBBYTES[1].a/w674 ) );
  XOR U8893 ( .A(n959), .B(n5837), .Z(n2970) );
  ANDN U8894 ( .A(\SUBBYTES[1].a/w580 ), .B(n2971), .Z(\SUBBYTES[1].a/w670 )
         );
  XNOR U8895 ( .A(\SUBBYTES[1].a/w639 ), .B(\SUBBYTES[1].a/w642 ), .Z(n2971)
         );
  AND U8896 ( .A(\SUBBYTES[1].a/w581 ), .B(n2972), .Z(\SUBBYTES[1].a/w668 ) );
  XNOR U8897 ( .A(n2975), .B(\SUBBYTES[1].a/w639 ), .Z(n2972) );
  AND U8898 ( .A(\SUBBYTES[1].a/w666 ), .B(n2976), .Z(\SUBBYTES[1].a/w667 ) );
  XOR U8899 ( .A(n2977), .B(n2975), .Z(n2976) );
  IV U8900 ( .A(n5836), .Z(n2975) );
  ANDN U8901 ( .A(\SUBBYTES[1].a/w685 ), .B(n2978), .Z(\SUBBYTES[1].a/w662 )
         );
  ANDN U8902 ( .A(\SUBBYTES[1].a/w686 ), .B(n2979), .Z(\SUBBYTES[1].a/w660 )
         );
  ANDN U8903 ( .A(\SUBBYTES[1].a/w689 ), .B(n2980), .Z(\SUBBYTES[1].a/w659 )
         );
  AND U8904 ( .A(\SUBBYTES[1].a/w645 ), .B(\SUBBYTES[1].a/w644 ), .Z(
        \SUBBYTES[1].a/w646 ) );
  IV U8905 ( .A(n2977), .Z(\SUBBYTES[1].a/w642 ) );
  NAND U8906 ( .A(\SUBBYTES[1].a/w621 ), .B(\SUBBYTES[1].a/w636 ), .Z(n2977)
         );
  AND U8907 ( .A(\SUBBYTES[1].a/w638 ), .B(\SUBBYTES[1].a/w644 ), .Z(
        \SUBBYTES[1].a/w639 ) );
  AND U8908 ( .A(\SUBBYTES[1].a/w623 ), .B(\SUBBYTES[1].a/w621 ), .Z(
        \SUBBYTES[1].a/w633 ) );
  AND U8909 ( .A(\SUBBYTES[1].a/w624 ), .B(\SUBBYTES[1].a/w622 ), .Z(
        \SUBBYTES[1].a/w631 ) );
  AND U8910 ( .A(\SUBBYTES[1].a/w638 ), .B(\SUBBYTES[1].a/w645 ), .Z(
        \SUBBYTES[1].a/w630 ) );
  AND U8911 ( .A(\SUBBYTES[1].a/w578 ), .B(\SUBBYTES[1].a/w574 ), .Z(
        \SUBBYTES[1].a/w615 ) );
  AND U8912 ( .A(\SUBBYTES[1].a/w579 ), .B(\SUBBYTES[1].a/w575 ), .Z(
        \SUBBYTES[1].a/w613 ) );
  ANDN U8913 ( .A(\SUBBYTES[1].a/w705 ), .B(n2974), .Z(\SUBBYTES[1].a/w612 )
         );
  XNOR U8914 ( .A(\w1[1][105] ), .B(\w1[1][111] ), .Z(n2974) );
  XOR U8915 ( .A(\w0[1][105] ), .B(g_input[233]), .Z(\w1[1][105] ) );
  AND U8916 ( .A(\w1[1][104] ), .B(\SUBBYTES[1].a/w580 ), .Z(
        \SUBBYTES[1].a/w608 ) );
  XOR U8917 ( .A(\w0[1][104] ), .B(g_input[232]), .Z(\w1[1][104] ) );
  AND U8918 ( .A(\SUBBYTES[1].a/w581 ), .B(\SUBBYTES[1].a/w577 ), .Z(
        \SUBBYTES[1].a/w606 ) );
  AND U8919 ( .A(\SUBBYTES[1].a/w666 ), .B(\SUBBYTES[1].a/w698 ), .Z(
        \SUBBYTES[1].a/w605 ) );
  ANDN U8920 ( .A(\SUBBYTES[1].a/w687 ), .B(n2978), .Z(\SUBBYTES[1].a/w600 )
         );
  XNOR U8921 ( .A(\w1[1][108] ), .B(\w1[1][111] ), .Z(n2978) );
  ANDN U8922 ( .A(\SUBBYTES[1].a/w688 ), .B(n2979), .Z(\SUBBYTES[1].a/w598 )
         );
  XNOR U8923 ( .A(\w1[1][106] ), .B(\w1[1][111] ), .Z(n2979) );
  XOR U8924 ( .A(\w0[1][111] ), .B(g_input[239]), .Z(\w1[1][111] ) );
  IV U8925 ( .A(n2981), .Z(\w1[1][106] ) );
  ANDN U8926 ( .A(\SUBBYTES[1].a/w690 ), .B(n2980), .Z(\SUBBYTES[1].a/w597 )
         );
  XOR U8927 ( .A(n2981), .B(\w1[1][108] ), .Z(n2980) );
  XOR U8928 ( .A(\w0[1][108] ), .B(g_input[236]), .Z(\w1[1][108] ) );
  XNOR U8929 ( .A(\w0[1][106] ), .B(g_input[234]), .Z(n2981) );
  AND U8930 ( .A(n2982), .B(\SUBBYTES[1].a/w367 ), .Z(\SUBBYTES[1].a/w502 ) );
  AND U8931 ( .A(n2983), .B(\SUBBYTES[1].a/w368 ), .Z(\SUBBYTES[1].a/w500 ) );
  AND U8932 ( .A(\SUBBYTES[1].a/w498 ), .B(n2984), .Z(\SUBBYTES[1].a/w499 ) );
  ANDN U8933 ( .A(\w1[1][112] ), .B(n2985), .Z(\SUBBYTES[1].a/w495 ) );
  AND U8934 ( .A(n2986), .B(\SUBBYTES[1].a/w370 ), .Z(\SUBBYTES[1].a/w493 ) );
  AND U8935 ( .A(\SUBBYTES[1].a/w491 ), .B(n2987), .Z(\SUBBYTES[1].a/w492 ) );
  XOR U8936 ( .A(\SUBBYTES[1].a/w435 ), .B(n5834), .Z(n2987) );
  AND U8937 ( .A(\SUBBYTES[1].a/w478 ), .B(\SUBBYTES[1].a/w480 ), .Z(
        \SUBBYTES[1].a/w487 ) );
  AND U8938 ( .A(\SUBBYTES[1].a/w479 ), .B(\SUBBYTES[1].a/w481 ), .Z(
        \SUBBYTES[1].a/w485 ) );
  AND U8939 ( .A(\SUBBYTES[1].a/w482 ), .B(\SUBBYTES[1].a/w483 ), .Z(
        \SUBBYTES[1].a/w484 ) );
  AND U8940 ( .A(\SUBBYTES[1].a/w371 ), .B(n2982), .Z(\SUBBYTES[1].a/w470 ) );
  XOR U8941 ( .A(\SUBBYTES[1].a/w439 ), .B(n958), .Z(n2982) );
  AND U8942 ( .A(\SUBBYTES[1].a/w372 ), .B(n2983), .Z(\SUBBYTES[1].a/w468 ) );
  XOR U8943 ( .A(n5835), .B(\SUBBYTES[1].a/w439 ), .Z(n2983) );
  ANDN U8944 ( .A(n2984), .B(n2988), .Z(\SUBBYTES[1].a/w467 ) );
  XOR U8945 ( .A(n958), .B(n5835), .Z(n2984) );
  ANDN U8946 ( .A(\SUBBYTES[1].a/w373 ), .B(n2985), .Z(\SUBBYTES[1].a/w463 )
         );
  XNOR U8947 ( .A(\SUBBYTES[1].a/w432 ), .B(\SUBBYTES[1].a/w435 ), .Z(n2985)
         );
  AND U8948 ( .A(\SUBBYTES[1].a/w374 ), .B(n2986), .Z(\SUBBYTES[1].a/w461 ) );
  XNOR U8949 ( .A(n2989), .B(\SUBBYTES[1].a/w432 ), .Z(n2986) );
  AND U8950 ( .A(\SUBBYTES[1].a/w459 ), .B(n2990), .Z(\SUBBYTES[1].a/w460 ) );
  XOR U8951 ( .A(n2991), .B(n2989), .Z(n2990) );
  IV U8952 ( .A(n5834), .Z(n2989) );
  ANDN U8953 ( .A(\SUBBYTES[1].a/w478 ), .B(n2992), .Z(\SUBBYTES[1].a/w455 )
         );
  ANDN U8954 ( .A(\SUBBYTES[1].a/w479 ), .B(n2993), .Z(\SUBBYTES[1].a/w453 )
         );
  ANDN U8955 ( .A(\SUBBYTES[1].a/w482 ), .B(n2994), .Z(\SUBBYTES[1].a/w452 )
         );
  AND U8956 ( .A(\SUBBYTES[1].a/w438 ), .B(\SUBBYTES[1].a/w437 ), .Z(
        \SUBBYTES[1].a/w439 ) );
  IV U8957 ( .A(n2991), .Z(\SUBBYTES[1].a/w435 ) );
  NAND U8958 ( .A(\SUBBYTES[1].a/w414 ), .B(\SUBBYTES[1].a/w429 ), .Z(n2991)
         );
  AND U8959 ( .A(\SUBBYTES[1].a/w431 ), .B(\SUBBYTES[1].a/w437 ), .Z(
        \SUBBYTES[1].a/w432 ) );
  AND U8960 ( .A(\SUBBYTES[1].a/w416 ), .B(\SUBBYTES[1].a/w414 ), .Z(
        \SUBBYTES[1].a/w426 ) );
  AND U8961 ( .A(\SUBBYTES[1].a/w417 ), .B(\SUBBYTES[1].a/w415 ), .Z(
        \SUBBYTES[1].a/w424 ) );
  AND U8962 ( .A(\SUBBYTES[1].a/w431 ), .B(\SUBBYTES[1].a/w438 ), .Z(
        \SUBBYTES[1].a/w423 ) );
  AND U8963 ( .A(\SUBBYTES[1].a/w371 ), .B(\SUBBYTES[1].a/w367 ), .Z(
        \SUBBYTES[1].a/w408 ) );
  AND U8964 ( .A(\SUBBYTES[1].a/w372 ), .B(\SUBBYTES[1].a/w368 ), .Z(
        \SUBBYTES[1].a/w406 ) );
  ANDN U8965 ( .A(\SUBBYTES[1].a/w498 ), .B(n2988), .Z(\SUBBYTES[1].a/w405 )
         );
  XNOR U8966 ( .A(\w1[1][113] ), .B(\w1[1][119] ), .Z(n2988) );
  XOR U8967 ( .A(\w0[1][113] ), .B(g_input[241]), .Z(\w1[1][113] ) );
  AND U8968 ( .A(\w1[1][112] ), .B(\SUBBYTES[1].a/w373 ), .Z(
        \SUBBYTES[1].a/w401 ) );
  XOR U8969 ( .A(\w0[1][112] ), .B(g_input[240]), .Z(\w1[1][112] ) );
  AND U8970 ( .A(\SUBBYTES[1].a/w374 ), .B(\SUBBYTES[1].a/w370 ), .Z(
        \SUBBYTES[1].a/w399 ) );
  AND U8971 ( .A(\SUBBYTES[1].a/w459 ), .B(\SUBBYTES[1].a/w491 ), .Z(
        \SUBBYTES[1].a/w398 ) );
  ANDN U8972 ( .A(\SUBBYTES[1].a/w480 ), .B(n2992), .Z(\SUBBYTES[1].a/w393 )
         );
  XNOR U8973 ( .A(\w1[1][116] ), .B(\w1[1][119] ), .Z(n2992) );
  ANDN U8974 ( .A(\SUBBYTES[1].a/w481 ), .B(n2993), .Z(\SUBBYTES[1].a/w391 )
         );
  XNOR U8975 ( .A(\w1[1][114] ), .B(\w1[1][119] ), .Z(n2993) );
  XOR U8976 ( .A(\w0[1][119] ), .B(g_input[247]), .Z(\w1[1][119] ) );
  IV U8977 ( .A(n2995), .Z(\w1[1][114] ) );
  ANDN U8978 ( .A(\SUBBYTES[1].a/w483 ), .B(n2994), .Z(\SUBBYTES[1].a/w390 )
         );
  XOR U8979 ( .A(n2995), .B(\w1[1][116] ), .Z(n2994) );
  XOR U8980 ( .A(\w0[1][116] ), .B(g_input[244]), .Z(\w1[1][116] ) );
  XNOR U8981 ( .A(\w0[1][114] ), .B(g_input[242]), .Z(n2995) );
  AND U8982 ( .A(n2996), .B(\SUBBYTES[1].a/w3265 ), .Z(\SUBBYTES[1].a/w3400 )
         );
  AND U8983 ( .A(n2997), .B(\SUBBYTES[1].a/w3266 ), .Z(\SUBBYTES[1].a/w3398 )
         );
  AND U8984 ( .A(\SUBBYTES[1].a/w3396 ), .B(n2998), .Z(\SUBBYTES[1].a/w3397 )
         );
  ANDN U8985 ( .A(\w1[1][0] ), .B(n2999), .Z(\SUBBYTES[1].a/w3393 ) );
  AND U8986 ( .A(n3000), .B(\SUBBYTES[1].a/w3268 ), .Z(\SUBBYTES[1].a/w3391 )
         );
  AND U8987 ( .A(\SUBBYTES[1].a/w3389 ), .B(n3001), .Z(\SUBBYTES[1].a/w3390 )
         );
  XOR U8988 ( .A(\SUBBYTES[1].a/w3333 ), .B(n5862), .Z(n3001) );
  AND U8989 ( .A(\SUBBYTES[1].a/w3376 ), .B(\SUBBYTES[1].a/w3378 ), .Z(
        \SUBBYTES[1].a/w3385 ) );
  AND U8990 ( .A(\SUBBYTES[1].a/w3377 ), .B(\SUBBYTES[1].a/w3379 ), .Z(
        \SUBBYTES[1].a/w3383 ) );
  AND U8991 ( .A(\SUBBYTES[1].a/w3380 ), .B(\SUBBYTES[1].a/w3381 ), .Z(
        \SUBBYTES[1].a/w3382 ) );
  AND U8992 ( .A(\SUBBYTES[1].a/w3269 ), .B(n2996), .Z(\SUBBYTES[1].a/w3368 )
         );
  XOR U8993 ( .A(\SUBBYTES[1].a/w3337 ), .B(n972), .Z(n2996) );
  AND U8994 ( .A(\SUBBYTES[1].a/w3270 ), .B(n2997), .Z(\SUBBYTES[1].a/w3366 )
         );
  XOR U8995 ( .A(n5863), .B(\SUBBYTES[1].a/w3337 ), .Z(n2997) );
  ANDN U8996 ( .A(n2998), .B(n3002), .Z(\SUBBYTES[1].a/w3365 ) );
  XOR U8997 ( .A(n972), .B(n5863), .Z(n2998) );
  ANDN U8998 ( .A(\SUBBYTES[1].a/w3271 ), .B(n2999), .Z(\SUBBYTES[1].a/w3361 )
         );
  XNOR U8999 ( .A(\SUBBYTES[1].a/w3330 ), .B(\SUBBYTES[1].a/w3333 ), .Z(n2999)
         );
  AND U9000 ( .A(\SUBBYTES[1].a/w3272 ), .B(n3000), .Z(\SUBBYTES[1].a/w3359 )
         );
  XNOR U9001 ( .A(n3003), .B(\SUBBYTES[1].a/w3330 ), .Z(n3000) );
  AND U9002 ( .A(\SUBBYTES[1].a/w3357 ), .B(n3004), .Z(\SUBBYTES[1].a/w3358 )
         );
  XOR U9003 ( .A(n3005), .B(n3003), .Z(n3004) );
  IV U9004 ( .A(n5862), .Z(n3003) );
  ANDN U9005 ( .A(\SUBBYTES[1].a/w3376 ), .B(n3006), .Z(\SUBBYTES[1].a/w3353 )
         );
  ANDN U9006 ( .A(\SUBBYTES[1].a/w3377 ), .B(n3007), .Z(\SUBBYTES[1].a/w3351 )
         );
  ANDN U9007 ( .A(\SUBBYTES[1].a/w3380 ), .B(n3008), .Z(\SUBBYTES[1].a/w3350 )
         );
  AND U9008 ( .A(\SUBBYTES[1].a/w3336 ), .B(\SUBBYTES[1].a/w3335 ), .Z(
        \SUBBYTES[1].a/w3337 ) );
  IV U9009 ( .A(n3005), .Z(\SUBBYTES[1].a/w3333 ) );
  NAND U9010 ( .A(\SUBBYTES[1].a/w3312 ), .B(\SUBBYTES[1].a/w3327 ), .Z(n3005)
         );
  AND U9011 ( .A(\SUBBYTES[1].a/w3329 ), .B(\SUBBYTES[1].a/w3335 ), .Z(
        \SUBBYTES[1].a/w3330 ) );
  AND U9012 ( .A(\SUBBYTES[1].a/w3314 ), .B(\SUBBYTES[1].a/w3312 ), .Z(
        \SUBBYTES[1].a/w3324 ) );
  AND U9013 ( .A(\SUBBYTES[1].a/w3315 ), .B(\SUBBYTES[1].a/w3313 ), .Z(
        \SUBBYTES[1].a/w3322 ) );
  AND U9014 ( .A(\SUBBYTES[1].a/w3329 ), .B(\SUBBYTES[1].a/w3336 ), .Z(
        \SUBBYTES[1].a/w3321 ) );
  AND U9015 ( .A(\SUBBYTES[1].a/w3269 ), .B(\SUBBYTES[1].a/w3265 ), .Z(
        \SUBBYTES[1].a/w3306 ) );
  AND U9016 ( .A(\SUBBYTES[1].a/w3270 ), .B(\SUBBYTES[1].a/w3266 ), .Z(
        \SUBBYTES[1].a/w3304 ) );
  ANDN U9017 ( .A(\SUBBYTES[1].a/w3396 ), .B(n3002), .Z(\SUBBYTES[1].a/w3303 )
         );
  XNOR U9018 ( .A(\w1[1][1] ), .B(\w1[1][7] ), .Z(n3002) );
  XOR U9019 ( .A(\w0[1][1] ), .B(g_input[129]), .Z(\w1[1][1] ) );
  AND U9020 ( .A(\w1[1][0] ), .B(\SUBBYTES[1].a/w3271 ), .Z(
        \SUBBYTES[1].a/w3299 ) );
  XOR U9021 ( .A(\w0[1][0] ), .B(g_input[128]), .Z(\w1[1][0] ) );
  AND U9022 ( .A(\SUBBYTES[1].a/w3272 ), .B(\SUBBYTES[1].a/w3268 ), .Z(
        \SUBBYTES[1].a/w3297 ) );
  AND U9023 ( .A(\SUBBYTES[1].a/w3357 ), .B(\SUBBYTES[1].a/w3389 ), .Z(
        \SUBBYTES[1].a/w3296 ) );
  ANDN U9024 ( .A(\SUBBYTES[1].a/w3378 ), .B(n3006), .Z(\SUBBYTES[1].a/w3291 )
         );
  XNOR U9025 ( .A(\w1[1][4] ), .B(\w1[1][7] ), .Z(n3006) );
  ANDN U9026 ( .A(\SUBBYTES[1].a/w3379 ), .B(n3007), .Z(\SUBBYTES[1].a/w3289 )
         );
  XNOR U9027 ( .A(\w1[1][2] ), .B(\w1[1][7] ), .Z(n3007) );
  XOR U9028 ( .A(\w0[1][7] ), .B(g_input[135]), .Z(\w1[1][7] ) );
  IV U9029 ( .A(n3009), .Z(\w1[1][2] ) );
  ANDN U9030 ( .A(\SUBBYTES[1].a/w3381 ), .B(n3008), .Z(\SUBBYTES[1].a/w3288 )
         );
  XOR U9031 ( .A(n3009), .B(\w1[1][4] ), .Z(n3008) );
  XOR U9032 ( .A(\w0[1][4] ), .B(g_input[132]), .Z(\w1[1][4] ) );
  XNOR U9033 ( .A(\w0[1][2] ), .B(g_input[130]), .Z(n3009) );
  AND U9034 ( .A(n3010), .B(\SUBBYTES[1].a/w3058 ), .Z(\SUBBYTES[1].a/w3193 )
         );
  AND U9035 ( .A(n3011), .B(\SUBBYTES[1].a/w3059 ), .Z(\SUBBYTES[1].a/w3191 )
         );
  AND U9036 ( .A(\SUBBYTES[1].a/w3189 ), .B(n3012), .Z(\SUBBYTES[1].a/w3190 )
         );
  ANDN U9037 ( .A(\w1[1][8] ), .B(n3013), .Z(\SUBBYTES[1].a/w3186 ) );
  AND U9038 ( .A(n3014), .B(\SUBBYTES[1].a/w3061 ), .Z(\SUBBYTES[1].a/w3184 )
         );
  AND U9039 ( .A(\SUBBYTES[1].a/w3182 ), .B(n3015), .Z(\SUBBYTES[1].a/w3183 )
         );
  XOR U9040 ( .A(\SUBBYTES[1].a/w3126 ), .B(n5860), .Z(n3015) );
  AND U9041 ( .A(\SUBBYTES[1].a/w3169 ), .B(\SUBBYTES[1].a/w3171 ), .Z(
        \SUBBYTES[1].a/w3178 ) );
  AND U9042 ( .A(\SUBBYTES[1].a/w3170 ), .B(\SUBBYTES[1].a/w3172 ), .Z(
        \SUBBYTES[1].a/w3176 ) );
  AND U9043 ( .A(\SUBBYTES[1].a/w3173 ), .B(\SUBBYTES[1].a/w3174 ), .Z(
        \SUBBYTES[1].a/w3175 ) );
  AND U9044 ( .A(\SUBBYTES[1].a/w3062 ), .B(n3010), .Z(\SUBBYTES[1].a/w3161 )
         );
  XOR U9045 ( .A(\SUBBYTES[1].a/w3130 ), .B(n971), .Z(n3010) );
  AND U9046 ( .A(\SUBBYTES[1].a/w3063 ), .B(n3011), .Z(\SUBBYTES[1].a/w3159 )
         );
  XOR U9047 ( .A(n5861), .B(\SUBBYTES[1].a/w3130 ), .Z(n3011) );
  ANDN U9048 ( .A(n3012), .B(n3016), .Z(\SUBBYTES[1].a/w3158 ) );
  XOR U9049 ( .A(n971), .B(n5861), .Z(n3012) );
  ANDN U9050 ( .A(\SUBBYTES[1].a/w3064 ), .B(n3013), .Z(\SUBBYTES[1].a/w3154 )
         );
  XNOR U9051 ( .A(\SUBBYTES[1].a/w3123 ), .B(\SUBBYTES[1].a/w3126 ), .Z(n3013)
         );
  AND U9052 ( .A(\SUBBYTES[1].a/w3065 ), .B(n3014), .Z(\SUBBYTES[1].a/w3152 )
         );
  XNOR U9053 ( .A(n3017), .B(\SUBBYTES[1].a/w3123 ), .Z(n3014) );
  AND U9054 ( .A(\SUBBYTES[1].a/w3150 ), .B(n3018), .Z(\SUBBYTES[1].a/w3151 )
         );
  XOR U9055 ( .A(n3019), .B(n3017), .Z(n3018) );
  IV U9056 ( .A(n5860), .Z(n3017) );
  ANDN U9057 ( .A(\SUBBYTES[1].a/w3169 ), .B(n3020), .Z(\SUBBYTES[1].a/w3146 )
         );
  ANDN U9058 ( .A(\SUBBYTES[1].a/w3170 ), .B(n3021), .Z(\SUBBYTES[1].a/w3144 )
         );
  ANDN U9059 ( .A(\SUBBYTES[1].a/w3173 ), .B(n3022), .Z(\SUBBYTES[1].a/w3143 )
         );
  AND U9060 ( .A(\SUBBYTES[1].a/w3129 ), .B(\SUBBYTES[1].a/w3128 ), .Z(
        \SUBBYTES[1].a/w3130 ) );
  IV U9061 ( .A(n3019), .Z(\SUBBYTES[1].a/w3126 ) );
  NAND U9062 ( .A(\SUBBYTES[1].a/w3105 ), .B(\SUBBYTES[1].a/w3120 ), .Z(n3019)
         );
  AND U9063 ( .A(\SUBBYTES[1].a/w3122 ), .B(\SUBBYTES[1].a/w3128 ), .Z(
        \SUBBYTES[1].a/w3123 ) );
  AND U9064 ( .A(\SUBBYTES[1].a/w3107 ), .B(\SUBBYTES[1].a/w3105 ), .Z(
        \SUBBYTES[1].a/w3117 ) );
  AND U9065 ( .A(\SUBBYTES[1].a/w3108 ), .B(\SUBBYTES[1].a/w3106 ), .Z(
        \SUBBYTES[1].a/w3115 ) );
  AND U9066 ( .A(\SUBBYTES[1].a/w3122 ), .B(\SUBBYTES[1].a/w3129 ), .Z(
        \SUBBYTES[1].a/w3114 ) );
  AND U9067 ( .A(\SUBBYTES[1].a/w3062 ), .B(\SUBBYTES[1].a/w3058 ), .Z(
        \SUBBYTES[1].a/w3099 ) );
  AND U9068 ( .A(\SUBBYTES[1].a/w3063 ), .B(\SUBBYTES[1].a/w3059 ), .Z(
        \SUBBYTES[1].a/w3097 ) );
  ANDN U9069 ( .A(\SUBBYTES[1].a/w3189 ), .B(n3016), .Z(\SUBBYTES[1].a/w3096 )
         );
  XNOR U9070 ( .A(\w1[1][15] ), .B(\w1[1][9] ), .Z(n3016) );
  XOR U9071 ( .A(\w0[1][9] ), .B(g_input[137]), .Z(\w1[1][9] ) );
  AND U9072 ( .A(\w1[1][8] ), .B(\SUBBYTES[1].a/w3064 ), .Z(
        \SUBBYTES[1].a/w3092 ) );
  XOR U9073 ( .A(\w0[1][8] ), .B(g_input[136]), .Z(\w1[1][8] ) );
  AND U9074 ( .A(\SUBBYTES[1].a/w3065 ), .B(\SUBBYTES[1].a/w3061 ), .Z(
        \SUBBYTES[1].a/w3090 ) );
  AND U9075 ( .A(\SUBBYTES[1].a/w3150 ), .B(\SUBBYTES[1].a/w3182 ), .Z(
        \SUBBYTES[1].a/w3089 ) );
  ANDN U9076 ( .A(\SUBBYTES[1].a/w3171 ), .B(n3020), .Z(\SUBBYTES[1].a/w3084 )
         );
  XNOR U9077 ( .A(\w1[1][12] ), .B(\w1[1][15] ), .Z(n3020) );
  ANDN U9078 ( .A(\SUBBYTES[1].a/w3172 ), .B(n3021), .Z(\SUBBYTES[1].a/w3082 )
         );
  XNOR U9079 ( .A(\w1[1][10] ), .B(\w1[1][15] ), .Z(n3021) );
  XOR U9080 ( .A(\w0[1][15] ), .B(g_input[143]), .Z(\w1[1][15] ) );
  ANDN U9081 ( .A(\SUBBYTES[1].a/w3174 ), .B(n3022), .Z(\SUBBYTES[1].a/w3081 )
         );
  XNOR U9082 ( .A(\w1[1][10] ), .B(\w1[1][12] ), .Z(n3022) );
  XOR U9083 ( .A(\w0[1][12] ), .B(g_input[140]), .Z(\w1[1][12] ) );
  XOR U9084 ( .A(\w0[1][10] ), .B(g_input[138]), .Z(\w1[1][10] ) );
  AND U9085 ( .A(n3023), .B(\SUBBYTES[1].a/w2851 ), .Z(\SUBBYTES[1].a/w2986 )
         );
  AND U9086 ( .A(n3024), .B(\SUBBYTES[1].a/w2852 ), .Z(\SUBBYTES[1].a/w2984 )
         );
  AND U9087 ( .A(\SUBBYTES[1].a/w2982 ), .B(n3025), .Z(\SUBBYTES[1].a/w2983 )
         );
  ANDN U9088 ( .A(\w1[1][16] ), .B(n3026), .Z(\SUBBYTES[1].a/w2979 ) );
  AND U9089 ( .A(n3027), .B(\SUBBYTES[1].a/w2854 ), .Z(\SUBBYTES[1].a/w2977 )
         );
  AND U9090 ( .A(\SUBBYTES[1].a/w2975 ), .B(n3028), .Z(\SUBBYTES[1].a/w2976 )
         );
  XOR U9091 ( .A(\SUBBYTES[1].a/w2919 ), .B(n5858), .Z(n3028) );
  AND U9092 ( .A(\SUBBYTES[1].a/w2962 ), .B(\SUBBYTES[1].a/w2964 ), .Z(
        \SUBBYTES[1].a/w2971 ) );
  AND U9093 ( .A(\SUBBYTES[1].a/w2963 ), .B(\SUBBYTES[1].a/w2965 ), .Z(
        \SUBBYTES[1].a/w2969 ) );
  AND U9094 ( .A(\SUBBYTES[1].a/w2966 ), .B(\SUBBYTES[1].a/w2967 ), .Z(
        \SUBBYTES[1].a/w2968 ) );
  AND U9095 ( .A(\SUBBYTES[1].a/w2855 ), .B(n3023), .Z(\SUBBYTES[1].a/w2954 )
         );
  XOR U9096 ( .A(\SUBBYTES[1].a/w2923 ), .B(n970), .Z(n3023) );
  AND U9097 ( .A(\SUBBYTES[1].a/w2856 ), .B(n3024), .Z(\SUBBYTES[1].a/w2952 )
         );
  XOR U9098 ( .A(n5859), .B(\SUBBYTES[1].a/w2923 ), .Z(n3024) );
  ANDN U9099 ( .A(n3025), .B(n3029), .Z(\SUBBYTES[1].a/w2951 ) );
  XOR U9100 ( .A(n970), .B(n5859), .Z(n3025) );
  AND U9101 ( .A(n3030), .B(\SUBBYTES[1].a/w160 ), .Z(\SUBBYTES[1].a/w295 ) );
  ANDN U9102 ( .A(\SUBBYTES[1].a/w2857 ), .B(n3026), .Z(\SUBBYTES[1].a/w2947 )
         );
  XNOR U9103 ( .A(\SUBBYTES[1].a/w2916 ), .B(\SUBBYTES[1].a/w2919 ), .Z(n3026)
         );
  AND U9104 ( .A(\SUBBYTES[1].a/w2858 ), .B(n3027), .Z(\SUBBYTES[1].a/w2945 )
         );
  XNOR U9105 ( .A(n3031), .B(\SUBBYTES[1].a/w2916 ), .Z(n3027) );
  AND U9106 ( .A(\SUBBYTES[1].a/w2943 ), .B(n3032), .Z(\SUBBYTES[1].a/w2944 )
         );
  XOR U9107 ( .A(n3033), .B(n3031), .Z(n3032) );
  IV U9108 ( .A(n5858), .Z(n3031) );
  ANDN U9109 ( .A(\SUBBYTES[1].a/w2962 ), .B(n3034), .Z(\SUBBYTES[1].a/w2939 )
         );
  ANDN U9110 ( .A(\SUBBYTES[1].a/w2963 ), .B(n3035), .Z(\SUBBYTES[1].a/w2937 )
         );
  ANDN U9111 ( .A(\SUBBYTES[1].a/w2966 ), .B(n3036), .Z(\SUBBYTES[1].a/w2936 )
         );
  AND U9112 ( .A(n3037), .B(\SUBBYTES[1].a/w161 ), .Z(\SUBBYTES[1].a/w293 ) );
  AND U9113 ( .A(\SUBBYTES[1].a/w2922 ), .B(\SUBBYTES[1].a/w2921 ), .Z(
        \SUBBYTES[1].a/w2923 ) );
  AND U9114 ( .A(\SUBBYTES[1].a/w291 ), .B(n3038), .Z(\SUBBYTES[1].a/w292 ) );
  IV U9115 ( .A(n3033), .Z(\SUBBYTES[1].a/w2919 ) );
  NAND U9116 ( .A(\SUBBYTES[1].a/w2898 ), .B(\SUBBYTES[1].a/w2913 ), .Z(n3033)
         );
  AND U9117 ( .A(\SUBBYTES[1].a/w2915 ), .B(\SUBBYTES[1].a/w2921 ), .Z(
        \SUBBYTES[1].a/w2916 ) );
  AND U9118 ( .A(\SUBBYTES[1].a/w2900 ), .B(\SUBBYTES[1].a/w2898 ), .Z(
        \SUBBYTES[1].a/w2910 ) );
  AND U9119 ( .A(\SUBBYTES[1].a/w2901 ), .B(\SUBBYTES[1].a/w2899 ), .Z(
        \SUBBYTES[1].a/w2908 ) );
  AND U9120 ( .A(\SUBBYTES[1].a/w2915 ), .B(\SUBBYTES[1].a/w2922 ), .Z(
        \SUBBYTES[1].a/w2907 ) );
  AND U9121 ( .A(\SUBBYTES[1].a/w2855 ), .B(\SUBBYTES[1].a/w2851 ), .Z(
        \SUBBYTES[1].a/w2892 ) );
  AND U9122 ( .A(\SUBBYTES[1].a/w2856 ), .B(\SUBBYTES[1].a/w2852 ), .Z(
        \SUBBYTES[1].a/w2890 ) );
  ANDN U9123 ( .A(\SUBBYTES[1].a/w2982 ), .B(n3029), .Z(\SUBBYTES[1].a/w2889 )
         );
  XNOR U9124 ( .A(\w1[1][17] ), .B(\w1[1][23] ), .Z(n3029) );
  XOR U9125 ( .A(\w0[1][17] ), .B(g_input[145]), .Z(\w1[1][17] ) );
  AND U9126 ( .A(\w1[1][16] ), .B(\SUBBYTES[1].a/w2857 ), .Z(
        \SUBBYTES[1].a/w2885 ) );
  XOR U9127 ( .A(\w0[1][16] ), .B(g_input[144]), .Z(\w1[1][16] ) );
  AND U9128 ( .A(\SUBBYTES[1].a/w2858 ), .B(\SUBBYTES[1].a/w2854 ), .Z(
        \SUBBYTES[1].a/w2883 ) );
  AND U9129 ( .A(\SUBBYTES[1].a/w2943 ), .B(\SUBBYTES[1].a/w2975 ), .Z(
        \SUBBYTES[1].a/w2882 ) );
  ANDN U9130 ( .A(\w1[1][120] ), .B(n3039), .Z(\SUBBYTES[1].a/w288 ) );
  ANDN U9131 ( .A(\SUBBYTES[1].a/w2964 ), .B(n3034), .Z(\SUBBYTES[1].a/w2877 )
         );
  XNOR U9132 ( .A(\w1[1][20] ), .B(\w1[1][23] ), .Z(n3034) );
  ANDN U9133 ( .A(\SUBBYTES[1].a/w2965 ), .B(n3035), .Z(\SUBBYTES[1].a/w2875 )
         );
  XNOR U9134 ( .A(\w1[1][18] ), .B(\w1[1][23] ), .Z(n3035) );
  XOR U9135 ( .A(\w0[1][23] ), .B(g_input[151]), .Z(\w1[1][23] ) );
  IV U9136 ( .A(n3040), .Z(\w1[1][18] ) );
  ANDN U9137 ( .A(\SUBBYTES[1].a/w2967 ), .B(n3036), .Z(\SUBBYTES[1].a/w2874 )
         );
  XOR U9138 ( .A(n3040), .B(\w1[1][20] ), .Z(n3036) );
  XOR U9139 ( .A(\w0[1][20] ), .B(g_input[148]), .Z(\w1[1][20] ) );
  XNOR U9140 ( .A(\w0[1][18] ), .B(g_input[146]), .Z(n3040) );
  AND U9141 ( .A(n3041), .B(\SUBBYTES[1].a/w163 ), .Z(\SUBBYTES[1].a/w286 ) );
  AND U9142 ( .A(\SUBBYTES[1].a/w284 ), .B(n3042), .Z(\SUBBYTES[1].a/w285 ) );
  XOR U9143 ( .A(\SUBBYTES[1].a/w228 ), .B(n5832), .Z(n3042) );
  AND U9144 ( .A(\SUBBYTES[1].a/w271 ), .B(\SUBBYTES[1].a/w273 ), .Z(
        \SUBBYTES[1].a/w280 ) );
  AND U9145 ( .A(\SUBBYTES[1].a/w272 ), .B(\SUBBYTES[1].a/w274 ), .Z(
        \SUBBYTES[1].a/w278 ) );
  AND U9146 ( .A(n3043), .B(\SUBBYTES[1].a/w2644 ), .Z(\SUBBYTES[1].a/w2779 )
         );
  AND U9147 ( .A(n3044), .B(\SUBBYTES[1].a/w2645 ), .Z(\SUBBYTES[1].a/w2777 )
         );
  AND U9148 ( .A(\SUBBYTES[1].a/w2775 ), .B(n3045), .Z(\SUBBYTES[1].a/w2776 )
         );
  ANDN U9149 ( .A(\w1[1][24] ), .B(n3046), .Z(\SUBBYTES[1].a/w2772 ) );
  AND U9150 ( .A(n3047), .B(\SUBBYTES[1].a/w2647 ), .Z(\SUBBYTES[1].a/w2770 )
         );
  AND U9151 ( .A(\SUBBYTES[1].a/w275 ), .B(\SUBBYTES[1].a/w276 ), .Z(
        \SUBBYTES[1].a/w277 ) );
  AND U9152 ( .A(\SUBBYTES[1].a/w2768 ), .B(n3048), .Z(\SUBBYTES[1].a/w2769 )
         );
  XOR U9153 ( .A(\SUBBYTES[1].a/w2712 ), .B(n5856), .Z(n3048) );
  AND U9154 ( .A(\SUBBYTES[1].a/w2755 ), .B(\SUBBYTES[1].a/w2757 ), .Z(
        \SUBBYTES[1].a/w2764 ) );
  AND U9155 ( .A(\SUBBYTES[1].a/w2756 ), .B(\SUBBYTES[1].a/w2758 ), .Z(
        \SUBBYTES[1].a/w2762 ) );
  AND U9156 ( .A(\SUBBYTES[1].a/w2759 ), .B(\SUBBYTES[1].a/w2760 ), .Z(
        \SUBBYTES[1].a/w2761 ) );
  AND U9157 ( .A(\SUBBYTES[1].a/w2648 ), .B(n3043), .Z(\SUBBYTES[1].a/w2747 )
         );
  XOR U9158 ( .A(\SUBBYTES[1].a/w2716 ), .B(n969), .Z(n3043) );
  AND U9159 ( .A(\SUBBYTES[1].a/w2649 ), .B(n3044), .Z(\SUBBYTES[1].a/w2745 )
         );
  XOR U9160 ( .A(n5857), .B(\SUBBYTES[1].a/w2716 ), .Z(n3044) );
  ANDN U9161 ( .A(n3045), .B(n3049), .Z(\SUBBYTES[1].a/w2744 ) );
  XOR U9162 ( .A(n969), .B(n5857), .Z(n3045) );
  ANDN U9163 ( .A(\SUBBYTES[1].a/w2650 ), .B(n3046), .Z(\SUBBYTES[1].a/w2740 )
         );
  XNOR U9164 ( .A(\SUBBYTES[1].a/w2709 ), .B(\SUBBYTES[1].a/w2712 ), .Z(n3046)
         );
  AND U9165 ( .A(\SUBBYTES[1].a/w2651 ), .B(n3047), .Z(\SUBBYTES[1].a/w2738 )
         );
  XNOR U9166 ( .A(n3050), .B(\SUBBYTES[1].a/w2709 ), .Z(n3047) );
  AND U9167 ( .A(\SUBBYTES[1].a/w2736 ), .B(n3051), .Z(\SUBBYTES[1].a/w2737 )
         );
  XOR U9168 ( .A(n3052), .B(n3050), .Z(n3051) );
  IV U9169 ( .A(n5856), .Z(n3050) );
  ANDN U9170 ( .A(\SUBBYTES[1].a/w2755 ), .B(n3053), .Z(\SUBBYTES[1].a/w2732 )
         );
  ANDN U9171 ( .A(\SUBBYTES[1].a/w2756 ), .B(n3054), .Z(\SUBBYTES[1].a/w2730 )
         );
  ANDN U9172 ( .A(\SUBBYTES[1].a/w2759 ), .B(n3055), .Z(\SUBBYTES[1].a/w2729 )
         );
  AND U9173 ( .A(\SUBBYTES[1].a/w2715 ), .B(\SUBBYTES[1].a/w2714 ), .Z(
        \SUBBYTES[1].a/w2716 ) );
  IV U9174 ( .A(n3052), .Z(\SUBBYTES[1].a/w2712 ) );
  NAND U9175 ( .A(\SUBBYTES[1].a/w2691 ), .B(\SUBBYTES[1].a/w2706 ), .Z(n3052)
         );
  AND U9176 ( .A(\SUBBYTES[1].a/w2708 ), .B(\SUBBYTES[1].a/w2714 ), .Z(
        \SUBBYTES[1].a/w2709 ) );
  AND U9177 ( .A(\SUBBYTES[1].a/w2693 ), .B(\SUBBYTES[1].a/w2691 ), .Z(
        \SUBBYTES[1].a/w2703 ) );
  AND U9178 ( .A(\SUBBYTES[1].a/w2694 ), .B(\SUBBYTES[1].a/w2692 ), .Z(
        \SUBBYTES[1].a/w2701 ) );
  AND U9179 ( .A(\SUBBYTES[1].a/w2708 ), .B(\SUBBYTES[1].a/w2715 ), .Z(
        \SUBBYTES[1].a/w2700 ) );
  AND U9180 ( .A(\SUBBYTES[1].a/w2648 ), .B(\SUBBYTES[1].a/w2644 ), .Z(
        \SUBBYTES[1].a/w2685 ) );
  AND U9181 ( .A(\SUBBYTES[1].a/w2649 ), .B(\SUBBYTES[1].a/w2645 ), .Z(
        \SUBBYTES[1].a/w2683 ) );
  ANDN U9182 ( .A(\SUBBYTES[1].a/w2775 ), .B(n3049), .Z(\SUBBYTES[1].a/w2682 )
         );
  XNOR U9183 ( .A(\w1[1][25] ), .B(\w1[1][31] ), .Z(n3049) );
  XOR U9184 ( .A(\w0[1][25] ), .B(g_input[153]), .Z(\w1[1][25] ) );
  AND U9185 ( .A(\w1[1][24] ), .B(\SUBBYTES[1].a/w2650 ), .Z(
        \SUBBYTES[1].a/w2678 ) );
  XOR U9186 ( .A(\w0[1][24] ), .B(g_input[152]), .Z(\w1[1][24] ) );
  AND U9187 ( .A(\SUBBYTES[1].a/w2651 ), .B(\SUBBYTES[1].a/w2647 ), .Z(
        \SUBBYTES[1].a/w2676 ) );
  AND U9188 ( .A(\SUBBYTES[1].a/w2736 ), .B(\SUBBYTES[1].a/w2768 ), .Z(
        \SUBBYTES[1].a/w2675 ) );
  ANDN U9189 ( .A(\SUBBYTES[1].a/w2757 ), .B(n3053), .Z(\SUBBYTES[1].a/w2670 )
         );
  XNOR U9190 ( .A(\w1[1][28] ), .B(\w1[1][31] ), .Z(n3053) );
  ANDN U9191 ( .A(\SUBBYTES[1].a/w2758 ), .B(n3054), .Z(\SUBBYTES[1].a/w2668 )
         );
  XNOR U9192 ( .A(\w1[1][26] ), .B(\w1[1][31] ), .Z(n3054) );
  XOR U9193 ( .A(\w0[1][31] ), .B(g_input[159]), .Z(\w1[1][31] ) );
  IV U9194 ( .A(n3056), .Z(\w1[1][26] ) );
  ANDN U9195 ( .A(\SUBBYTES[1].a/w2760 ), .B(n3055), .Z(\SUBBYTES[1].a/w2667 )
         );
  XOR U9196 ( .A(n3056), .B(\w1[1][28] ), .Z(n3055) );
  XOR U9197 ( .A(\w0[1][28] ), .B(g_input[156]), .Z(\w1[1][28] ) );
  XNOR U9198 ( .A(\w0[1][26] ), .B(g_input[154]), .Z(n3056) );
  AND U9199 ( .A(\SUBBYTES[1].a/w164 ), .B(n3030), .Z(\SUBBYTES[1].a/w263 ) );
  XOR U9200 ( .A(\SUBBYTES[1].a/w232 ), .B(n957), .Z(n3030) );
  AND U9201 ( .A(\SUBBYTES[1].a/w165 ), .B(n3037), .Z(\SUBBYTES[1].a/w261 ) );
  XOR U9202 ( .A(n5833), .B(\SUBBYTES[1].a/w232 ), .Z(n3037) );
  ANDN U9203 ( .A(n3038), .B(n3057), .Z(\SUBBYTES[1].a/w260 ) );
  XOR U9204 ( .A(n957), .B(n5833), .Z(n3038) );
  AND U9205 ( .A(n3058), .B(\SUBBYTES[1].a/w2437 ), .Z(\SUBBYTES[1].a/w2572 )
         );
  AND U9206 ( .A(n3059), .B(\SUBBYTES[1].a/w2438 ), .Z(\SUBBYTES[1].a/w2570 )
         );
  AND U9207 ( .A(\SUBBYTES[1].a/w2568 ), .B(n3060), .Z(\SUBBYTES[1].a/w2569 )
         );
  ANDN U9208 ( .A(\w1[1][32] ), .B(n3061), .Z(\SUBBYTES[1].a/w2565 ) );
  AND U9209 ( .A(n3062), .B(\SUBBYTES[1].a/w2440 ), .Z(\SUBBYTES[1].a/w2563 )
         );
  AND U9210 ( .A(\SUBBYTES[1].a/w2561 ), .B(n3063), .Z(\SUBBYTES[1].a/w2562 )
         );
  XOR U9211 ( .A(\SUBBYTES[1].a/w2505 ), .B(n5854), .Z(n3063) );
  ANDN U9212 ( .A(\SUBBYTES[1].a/w166 ), .B(n3039), .Z(\SUBBYTES[1].a/w256 )
         );
  XNOR U9213 ( .A(\SUBBYTES[1].a/w225 ), .B(\SUBBYTES[1].a/w228 ), .Z(n3039)
         );
  AND U9214 ( .A(\SUBBYTES[1].a/w2548 ), .B(\SUBBYTES[1].a/w2550 ), .Z(
        \SUBBYTES[1].a/w2557 ) );
  AND U9215 ( .A(\SUBBYTES[1].a/w2549 ), .B(\SUBBYTES[1].a/w2551 ), .Z(
        \SUBBYTES[1].a/w2555 ) );
  AND U9216 ( .A(\SUBBYTES[1].a/w2552 ), .B(\SUBBYTES[1].a/w2553 ), .Z(
        \SUBBYTES[1].a/w2554 ) );
  AND U9217 ( .A(\SUBBYTES[1].a/w2441 ), .B(n3058), .Z(\SUBBYTES[1].a/w2540 )
         );
  XOR U9218 ( .A(\SUBBYTES[1].a/w2509 ), .B(n968), .Z(n3058) );
  AND U9219 ( .A(\SUBBYTES[1].a/w167 ), .B(n3041), .Z(\SUBBYTES[1].a/w254 ) );
  XNOR U9220 ( .A(n3064), .B(\SUBBYTES[1].a/w225 ), .Z(n3041) );
  AND U9221 ( .A(\SUBBYTES[1].a/w2442 ), .B(n3059), .Z(\SUBBYTES[1].a/w2538 )
         );
  XOR U9222 ( .A(n5855), .B(\SUBBYTES[1].a/w2509 ), .Z(n3059) );
  ANDN U9223 ( .A(n3060), .B(n3065), .Z(\SUBBYTES[1].a/w2537 ) );
  XOR U9224 ( .A(n968), .B(n5855), .Z(n3060) );
  ANDN U9225 ( .A(\SUBBYTES[1].a/w2443 ), .B(n3061), .Z(\SUBBYTES[1].a/w2533 )
         );
  XNOR U9226 ( .A(\SUBBYTES[1].a/w2502 ), .B(\SUBBYTES[1].a/w2505 ), .Z(n3061)
         );
  AND U9227 ( .A(\SUBBYTES[1].a/w2444 ), .B(n3062), .Z(\SUBBYTES[1].a/w2531 )
         );
  XNOR U9228 ( .A(n3066), .B(\SUBBYTES[1].a/w2502 ), .Z(n3062) );
  AND U9229 ( .A(\SUBBYTES[1].a/w2529 ), .B(n3067), .Z(\SUBBYTES[1].a/w2530 )
         );
  XOR U9230 ( .A(n3068), .B(n3066), .Z(n3067) );
  IV U9231 ( .A(n5854), .Z(n3066) );
  AND U9232 ( .A(\SUBBYTES[1].a/w252 ), .B(n3069), .Z(\SUBBYTES[1].a/w253 ) );
  XOR U9233 ( .A(n3070), .B(n3064), .Z(n3069) );
  IV U9234 ( .A(n5832), .Z(n3064) );
  ANDN U9235 ( .A(\SUBBYTES[1].a/w2548 ), .B(n3071), .Z(\SUBBYTES[1].a/w2525 )
         );
  ANDN U9236 ( .A(\SUBBYTES[1].a/w2549 ), .B(n3072), .Z(\SUBBYTES[1].a/w2523 )
         );
  ANDN U9237 ( .A(\SUBBYTES[1].a/w2552 ), .B(n3073), .Z(\SUBBYTES[1].a/w2522 )
         );
  AND U9238 ( .A(\SUBBYTES[1].a/w2508 ), .B(\SUBBYTES[1].a/w2507 ), .Z(
        \SUBBYTES[1].a/w2509 ) );
  IV U9239 ( .A(n3068), .Z(\SUBBYTES[1].a/w2505 ) );
  NAND U9240 ( .A(\SUBBYTES[1].a/w2484 ), .B(\SUBBYTES[1].a/w2499 ), .Z(n3068)
         );
  AND U9241 ( .A(\SUBBYTES[1].a/w2501 ), .B(\SUBBYTES[1].a/w2507 ), .Z(
        \SUBBYTES[1].a/w2502 ) );
  AND U9242 ( .A(\SUBBYTES[1].a/w2486 ), .B(\SUBBYTES[1].a/w2484 ), .Z(
        \SUBBYTES[1].a/w2496 ) );
  AND U9243 ( .A(\SUBBYTES[1].a/w2487 ), .B(\SUBBYTES[1].a/w2485 ), .Z(
        \SUBBYTES[1].a/w2494 ) );
  AND U9244 ( .A(\SUBBYTES[1].a/w2501 ), .B(\SUBBYTES[1].a/w2508 ), .Z(
        \SUBBYTES[1].a/w2493 ) );
  ANDN U9245 ( .A(\SUBBYTES[1].a/w271 ), .B(n3074), .Z(\SUBBYTES[1].a/w248 )
         );
  AND U9246 ( .A(\SUBBYTES[1].a/w2441 ), .B(\SUBBYTES[1].a/w2437 ), .Z(
        \SUBBYTES[1].a/w2478 ) );
  AND U9247 ( .A(\SUBBYTES[1].a/w2442 ), .B(\SUBBYTES[1].a/w2438 ), .Z(
        \SUBBYTES[1].a/w2476 ) );
  ANDN U9248 ( .A(\SUBBYTES[1].a/w2568 ), .B(n3065), .Z(\SUBBYTES[1].a/w2475 )
         );
  XNOR U9249 ( .A(\w1[1][33] ), .B(\w1[1][39] ), .Z(n3065) );
  XOR U9250 ( .A(\w0[1][33] ), .B(g_input[161]), .Z(\w1[1][33] ) );
  AND U9251 ( .A(\w1[1][32] ), .B(\SUBBYTES[1].a/w2443 ), .Z(
        \SUBBYTES[1].a/w2471 ) );
  XOR U9252 ( .A(\w0[1][32] ), .B(g_input[160]), .Z(\w1[1][32] ) );
  AND U9253 ( .A(\SUBBYTES[1].a/w2444 ), .B(\SUBBYTES[1].a/w2440 ), .Z(
        \SUBBYTES[1].a/w2469 ) );
  AND U9254 ( .A(\SUBBYTES[1].a/w2529 ), .B(\SUBBYTES[1].a/w2561 ), .Z(
        \SUBBYTES[1].a/w2468 ) );
  ANDN U9255 ( .A(\SUBBYTES[1].a/w2550 ), .B(n3071), .Z(\SUBBYTES[1].a/w2463 )
         );
  XNOR U9256 ( .A(\w1[1][36] ), .B(\w1[1][39] ), .Z(n3071) );
  ANDN U9257 ( .A(\SUBBYTES[1].a/w2551 ), .B(n3072), .Z(\SUBBYTES[1].a/w2461 )
         );
  XNOR U9258 ( .A(\w1[1][34] ), .B(\w1[1][39] ), .Z(n3072) );
  XOR U9259 ( .A(\w0[1][39] ), .B(g_input[167]), .Z(\w1[1][39] ) );
  IV U9260 ( .A(n3075), .Z(\w1[1][34] ) );
  ANDN U9261 ( .A(\SUBBYTES[1].a/w2553 ), .B(n3073), .Z(\SUBBYTES[1].a/w2460 )
         );
  XOR U9262 ( .A(n3075), .B(\w1[1][36] ), .Z(n3073) );
  XOR U9263 ( .A(\w0[1][36] ), .B(g_input[164]), .Z(\w1[1][36] ) );
  XNOR U9264 ( .A(\w0[1][34] ), .B(g_input[162]), .Z(n3075) );
  ANDN U9265 ( .A(\SUBBYTES[1].a/w272 ), .B(n3076), .Z(\SUBBYTES[1].a/w246 )
         );
  ANDN U9266 ( .A(\SUBBYTES[1].a/w275 ), .B(n3077), .Z(\SUBBYTES[1].a/w245 )
         );
  AND U9267 ( .A(n3078), .B(\SUBBYTES[1].a/w2230 ), .Z(\SUBBYTES[1].a/w2365 )
         );
  AND U9268 ( .A(n3079), .B(\SUBBYTES[1].a/w2231 ), .Z(\SUBBYTES[1].a/w2363 )
         );
  AND U9269 ( .A(\SUBBYTES[1].a/w2361 ), .B(n3080), .Z(\SUBBYTES[1].a/w2362 )
         );
  ANDN U9270 ( .A(\w1[1][40] ), .B(n3081), .Z(\SUBBYTES[1].a/w2358 ) );
  AND U9271 ( .A(n3082), .B(\SUBBYTES[1].a/w2233 ), .Z(\SUBBYTES[1].a/w2356 )
         );
  AND U9272 ( .A(\SUBBYTES[1].a/w2354 ), .B(n3083), .Z(\SUBBYTES[1].a/w2355 )
         );
  XOR U9273 ( .A(\SUBBYTES[1].a/w2298 ), .B(n5852), .Z(n3083) );
  AND U9274 ( .A(\SUBBYTES[1].a/w2341 ), .B(\SUBBYTES[1].a/w2343 ), .Z(
        \SUBBYTES[1].a/w2350 ) );
  AND U9275 ( .A(\SUBBYTES[1].a/w2342 ), .B(\SUBBYTES[1].a/w2344 ), .Z(
        \SUBBYTES[1].a/w2348 ) );
  AND U9276 ( .A(\SUBBYTES[1].a/w2345 ), .B(\SUBBYTES[1].a/w2346 ), .Z(
        \SUBBYTES[1].a/w2347 ) );
  AND U9277 ( .A(\SUBBYTES[1].a/w2234 ), .B(n3078), .Z(\SUBBYTES[1].a/w2333 )
         );
  XOR U9278 ( .A(\SUBBYTES[1].a/w2302 ), .B(n967), .Z(n3078) );
  AND U9279 ( .A(\SUBBYTES[1].a/w2235 ), .B(n3079), .Z(\SUBBYTES[1].a/w2331 )
         );
  XOR U9280 ( .A(n5853), .B(\SUBBYTES[1].a/w2302 ), .Z(n3079) );
  ANDN U9281 ( .A(n3080), .B(n3084), .Z(\SUBBYTES[1].a/w2330 ) );
  XOR U9282 ( .A(n967), .B(n5853), .Z(n3080) );
  ANDN U9283 ( .A(\SUBBYTES[1].a/w2236 ), .B(n3081), .Z(\SUBBYTES[1].a/w2326 )
         );
  XNOR U9284 ( .A(\SUBBYTES[1].a/w2295 ), .B(\SUBBYTES[1].a/w2298 ), .Z(n3081)
         );
  AND U9285 ( .A(\SUBBYTES[1].a/w2237 ), .B(n3082), .Z(\SUBBYTES[1].a/w2324 )
         );
  XNOR U9286 ( .A(n3085), .B(\SUBBYTES[1].a/w2295 ), .Z(n3082) );
  AND U9287 ( .A(\SUBBYTES[1].a/w2322 ), .B(n3086), .Z(\SUBBYTES[1].a/w2323 )
         );
  XOR U9288 ( .A(n3087), .B(n3085), .Z(n3086) );
  IV U9289 ( .A(n5852), .Z(n3085) );
  AND U9290 ( .A(\SUBBYTES[1].a/w231 ), .B(\SUBBYTES[1].a/w230 ), .Z(
        \SUBBYTES[1].a/w232 ) );
  ANDN U9291 ( .A(\SUBBYTES[1].a/w2341 ), .B(n3088), .Z(\SUBBYTES[1].a/w2318 )
         );
  ANDN U9292 ( .A(\SUBBYTES[1].a/w2342 ), .B(n3089), .Z(\SUBBYTES[1].a/w2316 )
         );
  ANDN U9293 ( .A(\SUBBYTES[1].a/w2345 ), .B(n3090), .Z(\SUBBYTES[1].a/w2315 )
         );
  AND U9294 ( .A(\SUBBYTES[1].a/w2301 ), .B(\SUBBYTES[1].a/w2300 ), .Z(
        \SUBBYTES[1].a/w2302 ) );
  IV U9295 ( .A(n3087), .Z(\SUBBYTES[1].a/w2298 ) );
  NAND U9296 ( .A(\SUBBYTES[1].a/w2277 ), .B(\SUBBYTES[1].a/w2292 ), .Z(n3087)
         );
  AND U9297 ( .A(\SUBBYTES[1].a/w2294 ), .B(\SUBBYTES[1].a/w2300 ), .Z(
        \SUBBYTES[1].a/w2295 ) );
  AND U9298 ( .A(\SUBBYTES[1].a/w2279 ), .B(\SUBBYTES[1].a/w2277 ), .Z(
        \SUBBYTES[1].a/w2289 ) );
  AND U9299 ( .A(\SUBBYTES[1].a/w2280 ), .B(\SUBBYTES[1].a/w2278 ), .Z(
        \SUBBYTES[1].a/w2287 ) );
  AND U9300 ( .A(\SUBBYTES[1].a/w2294 ), .B(\SUBBYTES[1].a/w2301 ), .Z(
        \SUBBYTES[1].a/w2286 ) );
  IV U9301 ( .A(n3070), .Z(\SUBBYTES[1].a/w228 ) );
  NAND U9302 ( .A(\SUBBYTES[1].a/w207 ), .B(\SUBBYTES[1].a/w222 ), .Z(n3070)
         );
  AND U9303 ( .A(\SUBBYTES[1].a/w2234 ), .B(\SUBBYTES[1].a/w2230 ), .Z(
        \SUBBYTES[1].a/w2271 ) );
  AND U9304 ( .A(\SUBBYTES[1].a/w2235 ), .B(\SUBBYTES[1].a/w2231 ), .Z(
        \SUBBYTES[1].a/w2269 ) );
  ANDN U9305 ( .A(\SUBBYTES[1].a/w2361 ), .B(n3084), .Z(\SUBBYTES[1].a/w2268 )
         );
  XNOR U9306 ( .A(\w1[1][41] ), .B(\w1[1][47] ), .Z(n3084) );
  XOR U9307 ( .A(\w0[1][41] ), .B(g_input[169]), .Z(\w1[1][41] ) );
  AND U9308 ( .A(\w1[1][40] ), .B(\SUBBYTES[1].a/w2236 ), .Z(
        \SUBBYTES[1].a/w2264 ) );
  XOR U9309 ( .A(\w0[1][40] ), .B(g_input[168]), .Z(\w1[1][40] ) );
  AND U9310 ( .A(\SUBBYTES[1].a/w2237 ), .B(\SUBBYTES[1].a/w2233 ), .Z(
        \SUBBYTES[1].a/w2262 ) );
  AND U9311 ( .A(\SUBBYTES[1].a/w2322 ), .B(\SUBBYTES[1].a/w2354 ), .Z(
        \SUBBYTES[1].a/w2261 ) );
  ANDN U9312 ( .A(\SUBBYTES[1].a/w2343 ), .B(n3088), .Z(\SUBBYTES[1].a/w2256 )
         );
  XNOR U9313 ( .A(\w1[1][44] ), .B(\w1[1][47] ), .Z(n3088) );
  ANDN U9314 ( .A(\SUBBYTES[1].a/w2344 ), .B(n3089), .Z(\SUBBYTES[1].a/w2254 )
         );
  XNOR U9315 ( .A(\w1[1][42] ), .B(\w1[1][47] ), .Z(n3089) );
  XOR U9316 ( .A(\w0[1][47] ), .B(g_input[175]), .Z(\w1[1][47] ) );
  IV U9317 ( .A(n3091), .Z(\w1[1][42] ) );
  ANDN U9318 ( .A(\SUBBYTES[1].a/w2346 ), .B(n3090), .Z(\SUBBYTES[1].a/w2253 )
         );
  XOR U9319 ( .A(n3091), .B(\w1[1][44] ), .Z(n3090) );
  XOR U9320 ( .A(\w0[1][44] ), .B(g_input[172]), .Z(\w1[1][44] ) );
  XNOR U9321 ( .A(\w0[1][42] ), .B(g_input[170]), .Z(n3091) );
  AND U9322 ( .A(\SUBBYTES[1].a/w224 ), .B(\SUBBYTES[1].a/w230 ), .Z(
        \SUBBYTES[1].a/w225 ) );
  AND U9323 ( .A(\SUBBYTES[1].a/w209 ), .B(\SUBBYTES[1].a/w207 ), .Z(
        \SUBBYTES[1].a/w219 ) );
  AND U9324 ( .A(\SUBBYTES[1].a/w210 ), .B(\SUBBYTES[1].a/w208 ), .Z(
        \SUBBYTES[1].a/w217 ) );
  AND U9325 ( .A(\SUBBYTES[1].a/w224 ), .B(\SUBBYTES[1].a/w231 ), .Z(
        \SUBBYTES[1].a/w216 ) );
  AND U9326 ( .A(n3092), .B(\SUBBYTES[1].a/w2023 ), .Z(\SUBBYTES[1].a/w2158 )
         );
  AND U9327 ( .A(n3093), .B(\SUBBYTES[1].a/w2024 ), .Z(\SUBBYTES[1].a/w2156 )
         );
  AND U9328 ( .A(\SUBBYTES[1].a/w2154 ), .B(n3094), .Z(\SUBBYTES[1].a/w2155 )
         );
  ANDN U9329 ( .A(\w1[1][48] ), .B(n3095), .Z(\SUBBYTES[1].a/w2151 ) );
  AND U9330 ( .A(n3096), .B(\SUBBYTES[1].a/w2026 ), .Z(\SUBBYTES[1].a/w2149 )
         );
  AND U9331 ( .A(\SUBBYTES[1].a/w2147 ), .B(n3097), .Z(\SUBBYTES[1].a/w2148 )
         );
  XOR U9332 ( .A(\SUBBYTES[1].a/w2091 ), .B(n5850), .Z(n3097) );
  AND U9333 ( .A(\SUBBYTES[1].a/w2134 ), .B(\SUBBYTES[1].a/w2136 ), .Z(
        \SUBBYTES[1].a/w2143 ) );
  AND U9334 ( .A(\SUBBYTES[1].a/w2135 ), .B(\SUBBYTES[1].a/w2137 ), .Z(
        \SUBBYTES[1].a/w2141 ) );
  AND U9335 ( .A(\SUBBYTES[1].a/w2138 ), .B(\SUBBYTES[1].a/w2139 ), .Z(
        \SUBBYTES[1].a/w2140 ) );
  AND U9336 ( .A(\SUBBYTES[1].a/w2027 ), .B(n3092), .Z(\SUBBYTES[1].a/w2126 )
         );
  XOR U9337 ( .A(\SUBBYTES[1].a/w2095 ), .B(n966), .Z(n3092) );
  AND U9338 ( .A(\SUBBYTES[1].a/w2028 ), .B(n3093), .Z(\SUBBYTES[1].a/w2124 )
         );
  XOR U9339 ( .A(n5851), .B(\SUBBYTES[1].a/w2095 ), .Z(n3093) );
  ANDN U9340 ( .A(n3094), .B(n3098), .Z(\SUBBYTES[1].a/w2123 ) );
  XOR U9341 ( .A(n966), .B(n5851), .Z(n3094) );
  ANDN U9342 ( .A(\SUBBYTES[1].a/w2029 ), .B(n3095), .Z(\SUBBYTES[1].a/w2119 )
         );
  XNOR U9343 ( .A(\SUBBYTES[1].a/w2088 ), .B(\SUBBYTES[1].a/w2091 ), .Z(n3095)
         );
  AND U9344 ( .A(\SUBBYTES[1].a/w2030 ), .B(n3096), .Z(\SUBBYTES[1].a/w2117 )
         );
  XNOR U9345 ( .A(n3099), .B(\SUBBYTES[1].a/w2088 ), .Z(n3096) );
  AND U9346 ( .A(\SUBBYTES[1].a/w2115 ), .B(n3100), .Z(\SUBBYTES[1].a/w2116 )
         );
  XOR U9347 ( .A(n3101), .B(n3099), .Z(n3100) );
  IV U9348 ( .A(n5850), .Z(n3099) );
  ANDN U9349 ( .A(\SUBBYTES[1].a/w2134 ), .B(n3102), .Z(\SUBBYTES[1].a/w2111 )
         );
  ANDN U9350 ( .A(\SUBBYTES[1].a/w2135 ), .B(n3103), .Z(\SUBBYTES[1].a/w2109 )
         );
  ANDN U9351 ( .A(\SUBBYTES[1].a/w2138 ), .B(n3104), .Z(\SUBBYTES[1].a/w2108 )
         );
  AND U9352 ( .A(\SUBBYTES[1].a/w2094 ), .B(\SUBBYTES[1].a/w2093 ), .Z(
        \SUBBYTES[1].a/w2095 ) );
  IV U9353 ( .A(n3101), .Z(\SUBBYTES[1].a/w2091 ) );
  NAND U9354 ( .A(\SUBBYTES[1].a/w2070 ), .B(\SUBBYTES[1].a/w2085 ), .Z(n3101)
         );
  AND U9355 ( .A(\SUBBYTES[1].a/w2087 ), .B(\SUBBYTES[1].a/w2093 ), .Z(
        \SUBBYTES[1].a/w2088 ) );
  AND U9356 ( .A(\SUBBYTES[1].a/w2072 ), .B(\SUBBYTES[1].a/w2070 ), .Z(
        \SUBBYTES[1].a/w2082 ) );
  AND U9357 ( .A(\SUBBYTES[1].a/w2073 ), .B(\SUBBYTES[1].a/w2071 ), .Z(
        \SUBBYTES[1].a/w2080 ) );
  AND U9358 ( .A(\SUBBYTES[1].a/w2087 ), .B(\SUBBYTES[1].a/w2094 ), .Z(
        \SUBBYTES[1].a/w2079 ) );
  AND U9359 ( .A(\SUBBYTES[1].a/w2027 ), .B(\SUBBYTES[1].a/w2023 ), .Z(
        \SUBBYTES[1].a/w2064 ) );
  AND U9360 ( .A(\SUBBYTES[1].a/w2028 ), .B(\SUBBYTES[1].a/w2024 ), .Z(
        \SUBBYTES[1].a/w2062 ) );
  ANDN U9361 ( .A(\SUBBYTES[1].a/w2154 ), .B(n3098), .Z(\SUBBYTES[1].a/w2061 )
         );
  XNOR U9362 ( .A(\w1[1][49] ), .B(\w1[1][55] ), .Z(n3098) );
  XOR U9363 ( .A(\w0[1][49] ), .B(g_input[177]), .Z(\w1[1][49] ) );
  AND U9364 ( .A(\w1[1][48] ), .B(\SUBBYTES[1].a/w2029 ), .Z(
        \SUBBYTES[1].a/w2057 ) );
  XOR U9365 ( .A(\w0[1][48] ), .B(g_input[176]), .Z(\w1[1][48] ) );
  AND U9366 ( .A(\SUBBYTES[1].a/w2030 ), .B(\SUBBYTES[1].a/w2026 ), .Z(
        \SUBBYTES[1].a/w2055 ) );
  AND U9367 ( .A(\SUBBYTES[1].a/w2115 ), .B(\SUBBYTES[1].a/w2147 ), .Z(
        \SUBBYTES[1].a/w2054 ) );
  ANDN U9368 ( .A(\SUBBYTES[1].a/w2136 ), .B(n3102), .Z(\SUBBYTES[1].a/w2049 )
         );
  XNOR U9369 ( .A(\w1[1][52] ), .B(\w1[1][55] ), .Z(n3102) );
  ANDN U9370 ( .A(\SUBBYTES[1].a/w2137 ), .B(n3103), .Z(\SUBBYTES[1].a/w2047 )
         );
  XNOR U9371 ( .A(\w1[1][50] ), .B(\w1[1][55] ), .Z(n3103) );
  XOR U9372 ( .A(\w0[1][55] ), .B(g_input[183]), .Z(\w1[1][55] ) );
  IV U9373 ( .A(n3105), .Z(\w1[1][50] ) );
  ANDN U9374 ( .A(\SUBBYTES[1].a/w2139 ), .B(n3104), .Z(\SUBBYTES[1].a/w2046 )
         );
  XOR U9375 ( .A(n3105), .B(\w1[1][52] ), .Z(n3104) );
  XOR U9376 ( .A(\w0[1][52] ), .B(g_input[180]), .Z(\w1[1][52] ) );
  XNOR U9377 ( .A(\w0[1][50] ), .B(g_input[178]), .Z(n3105) );
  AND U9378 ( .A(\SUBBYTES[1].a/w164 ), .B(\SUBBYTES[1].a/w160 ), .Z(
        \SUBBYTES[1].a/w201 ) );
  AND U9379 ( .A(\SUBBYTES[1].a/w165 ), .B(\SUBBYTES[1].a/w161 ), .Z(
        \SUBBYTES[1].a/w199 ) );
  ANDN U9380 ( .A(\SUBBYTES[1].a/w291 ), .B(n3057), .Z(\SUBBYTES[1].a/w198 )
         );
  XNOR U9381 ( .A(\w1[1][121] ), .B(\w1[1][127] ), .Z(n3057) );
  XOR U9382 ( .A(\w0[1][121] ), .B(g_input[249]), .Z(\w1[1][121] ) );
  AND U9383 ( .A(n3106), .B(\SUBBYTES[1].a/w1816 ), .Z(\SUBBYTES[1].a/w1951 )
         );
  AND U9384 ( .A(n3107), .B(\SUBBYTES[1].a/w1817 ), .Z(\SUBBYTES[1].a/w1949 )
         );
  AND U9385 ( .A(\SUBBYTES[1].a/w1947 ), .B(n3108), .Z(\SUBBYTES[1].a/w1948 )
         );
  ANDN U9386 ( .A(\w1[1][56] ), .B(n3109), .Z(\SUBBYTES[1].a/w1944 ) );
  AND U9387 ( .A(n3110), .B(\SUBBYTES[1].a/w1819 ), .Z(\SUBBYTES[1].a/w1942 )
         );
  AND U9388 ( .A(\SUBBYTES[1].a/w1940 ), .B(n3111), .Z(\SUBBYTES[1].a/w1941 )
         );
  XOR U9389 ( .A(\SUBBYTES[1].a/w1884 ), .B(n5848), .Z(n3111) );
  AND U9390 ( .A(\w1[1][120] ), .B(\SUBBYTES[1].a/w166 ), .Z(
        \SUBBYTES[1].a/w194 ) );
  XOR U9391 ( .A(\w0[1][120] ), .B(g_input[248]), .Z(\w1[1][120] ) );
  AND U9392 ( .A(\SUBBYTES[1].a/w1927 ), .B(\SUBBYTES[1].a/w1929 ), .Z(
        \SUBBYTES[1].a/w1936 ) );
  AND U9393 ( .A(\SUBBYTES[1].a/w1928 ), .B(\SUBBYTES[1].a/w1930 ), .Z(
        \SUBBYTES[1].a/w1934 ) );
  AND U9394 ( .A(\SUBBYTES[1].a/w1931 ), .B(\SUBBYTES[1].a/w1932 ), .Z(
        \SUBBYTES[1].a/w1933 ) );
  AND U9395 ( .A(\SUBBYTES[1].a/w167 ), .B(\SUBBYTES[1].a/w163 ), .Z(
        \SUBBYTES[1].a/w192 ) );
  AND U9396 ( .A(\SUBBYTES[1].a/w1820 ), .B(n3106), .Z(\SUBBYTES[1].a/w1919 )
         );
  XOR U9397 ( .A(\SUBBYTES[1].a/w1888 ), .B(n965), .Z(n3106) );
  AND U9398 ( .A(\SUBBYTES[1].a/w1821 ), .B(n3107), .Z(\SUBBYTES[1].a/w1917 )
         );
  XOR U9399 ( .A(n5849), .B(\SUBBYTES[1].a/w1888 ), .Z(n3107) );
  ANDN U9400 ( .A(n3108), .B(n3112), .Z(\SUBBYTES[1].a/w1916 ) );
  XOR U9401 ( .A(n965), .B(n5849), .Z(n3108) );
  ANDN U9402 ( .A(\SUBBYTES[1].a/w1822 ), .B(n3109), .Z(\SUBBYTES[1].a/w1912 )
         );
  XNOR U9403 ( .A(\SUBBYTES[1].a/w1881 ), .B(\SUBBYTES[1].a/w1884 ), .Z(n3109)
         );
  AND U9404 ( .A(\SUBBYTES[1].a/w1823 ), .B(n3110), .Z(\SUBBYTES[1].a/w1910 )
         );
  XNOR U9405 ( .A(n3113), .B(\SUBBYTES[1].a/w1881 ), .Z(n3110) );
  AND U9406 ( .A(\SUBBYTES[1].a/w252 ), .B(\SUBBYTES[1].a/w284 ), .Z(
        \SUBBYTES[1].a/w191 ) );
  AND U9407 ( .A(\SUBBYTES[1].a/w1908 ), .B(n3114), .Z(\SUBBYTES[1].a/w1909 )
         );
  XOR U9408 ( .A(n3115), .B(n3113), .Z(n3114) );
  IV U9409 ( .A(n5848), .Z(n3113) );
  ANDN U9410 ( .A(\SUBBYTES[1].a/w1927 ), .B(n3116), .Z(\SUBBYTES[1].a/w1904 )
         );
  ANDN U9411 ( .A(\SUBBYTES[1].a/w1928 ), .B(n3117), .Z(\SUBBYTES[1].a/w1902 )
         );
  ANDN U9412 ( .A(\SUBBYTES[1].a/w1931 ), .B(n3118), .Z(\SUBBYTES[1].a/w1901 )
         );
  AND U9413 ( .A(\SUBBYTES[1].a/w1887 ), .B(\SUBBYTES[1].a/w1886 ), .Z(
        \SUBBYTES[1].a/w1888 ) );
  IV U9414 ( .A(n3115), .Z(\SUBBYTES[1].a/w1884 ) );
  NAND U9415 ( .A(\SUBBYTES[1].a/w1863 ), .B(\SUBBYTES[1].a/w1878 ), .Z(n3115)
         );
  AND U9416 ( .A(\SUBBYTES[1].a/w1880 ), .B(\SUBBYTES[1].a/w1886 ), .Z(
        \SUBBYTES[1].a/w1881 ) );
  AND U9417 ( .A(\SUBBYTES[1].a/w1865 ), .B(\SUBBYTES[1].a/w1863 ), .Z(
        \SUBBYTES[1].a/w1875 ) );
  AND U9418 ( .A(\SUBBYTES[1].a/w1866 ), .B(\SUBBYTES[1].a/w1864 ), .Z(
        \SUBBYTES[1].a/w1873 ) );
  AND U9419 ( .A(\SUBBYTES[1].a/w1880 ), .B(\SUBBYTES[1].a/w1887 ), .Z(
        \SUBBYTES[1].a/w1872 ) );
  ANDN U9420 ( .A(\SUBBYTES[1].a/w273 ), .B(n3074), .Z(\SUBBYTES[1].a/w186 )
         );
  XNOR U9421 ( .A(\w1[1][124] ), .B(\w1[1][127] ), .Z(n3074) );
  AND U9422 ( .A(\SUBBYTES[1].a/w1820 ), .B(\SUBBYTES[1].a/w1816 ), .Z(
        \SUBBYTES[1].a/w1857 ) );
  AND U9423 ( .A(\SUBBYTES[1].a/w1821 ), .B(\SUBBYTES[1].a/w1817 ), .Z(
        \SUBBYTES[1].a/w1855 ) );
  ANDN U9424 ( .A(\SUBBYTES[1].a/w1947 ), .B(n3112), .Z(\SUBBYTES[1].a/w1854 )
         );
  XNOR U9425 ( .A(\w1[1][57] ), .B(\w1[1][63] ), .Z(n3112) );
  XOR U9426 ( .A(\w0[1][57] ), .B(g_input[185]), .Z(\w1[1][57] ) );
  AND U9427 ( .A(\w1[1][56] ), .B(\SUBBYTES[1].a/w1822 ), .Z(
        \SUBBYTES[1].a/w1850 ) );
  XOR U9428 ( .A(\w0[1][56] ), .B(g_input[184]), .Z(\w1[1][56] ) );
  AND U9429 ( .A(\SUBBYTES[1].a/w1823 ), .B(\SUBBYTES[1].a/w1819 ), .Z(
        \SUBBYTES[1].a/w1848 ) );
  AND U9430 ( .A(\SUBBYTES[1].a/w1908 ), .B(\SUBBYTES[1].a/w1940 ), .Z(
        \SUBBYTES[1].a/w1847 ) );
  ANDN U9431 ( .A(\SUBBYTES[1].a/w1929 ), .B(n3116), .Z(\SUBBYTES[1].a/w1842 )
         );
  XNOR U9432 ( .A(\w1[1][60] ), .B(\w1[1][63] ), .Z(n3116) );
  ANDN U9433 ( .A(\SUBBYTES[1].a/w1930 ), .B(n3117), .Z(\SUBBYTES[1].a/w1840 )
         );
  XNOR U9434 ( .A(\w1[1][58] ), .B(\w1[1][63] ), .Z(n3117) );
  XOR U9435 ( .A(\w0[1][63] ), .B(g_input[191]), .Z(\w1[1][63] ) );
  IV U9436 ( .A(n3119), .Z(\w1[1][58] ) );
  ANDN U9437 ( .A(\SUBBYTES[1].a/w274 ), .B(n3076), .Z(\SUBBYTES[1].a/w184 )
         );
  XNOR U9438 ( .A(\w1[1][122] ), .B(\w1[1][127] ), .Z(n3076) );
  XOR U9439 ( .A(\w0[1][127] ), .B(g_input[255]), .Z(\w1[1][127] ) );
  IV U9440 ( .A(n3120), .Z(\w1[1][122] ) );
  ANDN U9441 ( .A(\SUBBYTES[1].a/w1932 ), .B(n3118), .Z(\SUBBYTES[1].a/w1839 )
         );
  XOR U9442 ( .A(n3119), .B(\w1[1][60] ), .Z(n3118) );
  XOR U9443 ( .A(\w0[1][60] ), .B(g_input[188]), .Z(\w1[1][60] ) );
  XNOR U9444 ( .A(\w0[1][58] ), .B(g_input[186]), .Z(n3119) );
  ANDN U9445 ( .A(\SUBBYTES[1].a/w276 ), .B(n3077), .Z(\SUBBYTES[1].a/w183 )
         );
  XOR U9446 ( .A(n3120), .B(\w1[1][124] ), .Z(n3077) );
  XOR U9447 ( .A(\w0[1][124] ), .B(g_input[252]), .Z(\w1[1][124] ) );
  XNOR U9448 ( .A(\w0[1][122] ), .B(g_input[250]), .Z(n3120) );
  AND U9449 ( .A(n3121), .B(\SUBBYTES[1].a/w1609 ), .Z(\SUBBYTES[1].a/w1744 )
         );
  AND U9450 ( .A(n3122), .B(\SUBBYTES[1].a/w1610 ), .Z(\SUBBYTES[1].a/w1742 )
         );
  AND U9451 ( .A(\SUBBYTES[1].a/w1740 ), .B(n3123), .Z(\SUBBYTES[1].a/w1741 )
         );
  ANDN U9452 ( .A(\w1[1][64] ), .B(n3124), .Z(\SUBBYTES[1].a/w1737 ) );
  AND U9453 ( .A(n3125), .B(\SUBBYTES[1].a/w1612 ), .Z(\SUBBYTES[1].a/w1735 )
         );
  AND U9454 ( .A(\SUBBYTES[1].a/w1733 ), .B(n3126), .Z(\SUBBYTES[1].a/w1734 )
         );
  XOR U9455 ( .A(\SUBBYTES[1].a/w1677 ), .B(n5846), .Z(n3126) );
  AND U9456 ( .A(\SUBBYTES[1].a/w1720 ), .B(\SUBBYTES[1].a/w1722 ), .Z(
        \SUBBYTES[1].a/w1729 ) );
  AND U9457 ( .A(\SUBBYTES[1].a/w1721 ), .B(\SUBBYTES[1].a/w1723 ), .Z(
        \SUBBYTES[1].a/w1727 ) );
  AND U9458 ( .A(\SUBBYTES[1].a/w1724 ), .B(\SUBBYTES[1].a/w1725 ), .Z(
        \SUBBYTES[1].a/w1726 ) );
  AND U9459 ( .A(\SUBBYTES[1].a/w1613 ), .B(n3121), .Z(\SUBBYTES[1].a/w1712 )
         );
  XOR U9460 ( .A(\SUBBYTES[1].a/w1681 ), .B(n964), .Z(n3121) );
  AND U9461 ( .A(\SUBBYTES[1].a/w1614 ), .B(n3122), .Z(\SUBBYTES[1].a/w1710 )
         );
  XOR U9462 ( .A(n5847), .B(\SUBBYTES[1].a/w1681 ), .Z(n3122) );
  ANDN U9463 ( .A(n3123), .B(n3127), .Z(\SUBBYTES[1].a/w1709 ) );
  XOR U9464 ( .A(n964), .B(n5847), .Z(n3123) );
  ANDN U9465 ( .A(\SUBBYTES[1].a/w1615 ), .B(n3124), .Z(\SUBBYTES[1].a/w1705 )
         );
  XNOR U9466 ( .A(\SUBBYTES[1].a/w1674 ), .B(\SUBBYTES[1].a/w1677 ), .Z(n3124)
         );
  AND U9467 ( .A(\SUBBYTES[1].a/w1616 ), .B(n3125), .Z(\SUBBYTES[1].a/w1703 )
         );
  XNOR U9468 ( .A(n3128), .B(\SUBBYTES[1].a/w1674 ), .Z(n3125) );
  AND U9469 ( .A(\SUBBYTES[1].a/w1701 ), .B(n3129), .Z(\SUBBYTES[1].a/w1702 )
         );
  XOR U9470 ( .A(n3130), .B(n3128), .Z(n3129) );
  IV U9471 ( .A(n5846), .Z(n3128) );
  ANDN U9472 ( .A(\SUBBYTES[1].a/w1720 ), .B(n3131), .Z(\SUBBYTES[1].a/w1697 )
         );
  ANDN U9473 ( .A(\SUBBYTES[1].a/w1721 ), .B(n3132), .Z(\SUBBYTES[1].a/w1695 )
         );
  ANDN U9474 ( .A(\SUBBYTES[1].a/w1724 ), .B(n3133), .Z(\SUBBYTES[1].a/w1694 )
         );
  AND U9475 ( .A(\SUBBYTES[1].a/w1680 ), .B(\SUBBYTES[1].a/w1679 ), .Z(
        \SUBBYTES[1].a/w1681 ) );
  IV U9476 ( .A(n3130), .Z(\SUBBYTES[1].a/w1677 ) );
  NAND U9477 ( .A(\SUBBYTES[1].a/w1656 ), .B(\SUBBYTES[1].a/w1671 ), .Z(n3130)
         );
  AND U9478 ( .A(\SUBBYTES[1].a/w1673 ), .B(\SUBBYTES[1].a/w1679 ), .Z(
        \SUBBYTES[1].a/w1674 ) );
  AND U9479 ( .A(\SUBBYTES[1].a/w1658 ), .B(\SUBBYTES[1].a/w1656 ), .Z(
        \SUBBYTES[1].a/w1668 ) );
  AND U9480 ( .A(\SUBBYTES[1].a/w1659 ), .B(\SUBBYTES[1].a/w1657 ), .Z(
        \SUBBYTES[1].a/w1666 ) );
  AND U9481 ( .A(\SUBBYTES[1].a/w1673 ), .B(\SUBBYTES[1].a/w1680 ), .Z(
        \SUBBYTES[1].a/w1665 ) );
  AND U9482 ( .A(\SUBBYTES[1].a/w1613 ), .B(\SUBBYTES[1].a/w1609 ), .Z(
        \SUBBYTES[1].a/w1650 ) );
  AND U9483 ( .A(\SUBBYTES[1].a/w1614 ), .B(\SUBBYTES[1].a/w1610 ), .Z(
        \SUBBYTES[1].a/w1648 ) );
  ANDN U9484 ( .A(\SUBBYTES[1].a/w1740 ), .B(n3127), .Z(\SUBBYTES[1].a/w1647 )
         );
  XNOR U9485 ( .A(\w1[1][65] ), .B(\w1[1][71] ), .Z(n3127) );
  XOR U9486 ( .A(\w0[1][65] ), .B(g_input[193]), .Z(\w1[1][65] ) );
  AND U9487 ( .A(\w1[1][64] ), .B(\SUBBYTES[1].a/w1615 ), .Z(
        \SUBBYTES[1].a/w1643 ) );
  XOR U9488 ( .A(\w0[1][64] ), .B(g_input[192]), .Z(\w1[1][64] ) );
  AND U9489 ( .A(\SUBBYTES[1].a/w1616 ), .B(\SUBBYTES[1].a/w1612 ), .Z(
        \SUBBYTES[1].a/w1641 ) );
  AND U9490 ( .A(\SUBBYTES[1].a/w1701 ), .B(\SUBBYTES[1].a/w1733 ), .Z(
        \SUBBYTES[1].a/w1640 ) );
  ANDN U9491 ( .A(\SUBBYTES[1].a/w1722 ), .B(n3131), .Z(\SUBBYTES[1].a/w1635 )
         );
  XNOR U9492 ( .A(\w1[1][68] ), .B(\w1[1][71] ), .Z(n3131) );
  ANDN U9493 ( .A(\SUBBYTES[1].a/w1723 ), .B(n3132), .Z(\SUBBYTES[1].a/w1633 )
         );
  XNOR U9494 ( .A(\w1[1][66] ), .B(\w1[1][71] ), .Z(n3132) );
  XOR U9495 ( .A(\w0[1][71] ), .B(g_input[199]), .Z(\w1[1][71] ) );
  IV U9496 ( .A(n3134), .Z(\w1[1][66] ) );
  ANDN U9497 ( .A(\SUBBYTES[1].a/w1725 ), .B(n3133), .Z(\SUBBYTES[1].a/w1632 )
         );
  XOR U9498 ( .A(n3134), .B(\w1[1][68] ), .Z(n3133) );
  XOR U9499 ( .A(\w0[1][68] ), .B(g_input[196]), .Z(\w1[1][68] ) );
  XNOR U9500 ( .A(\w0[1][66] ), .B(g_input[194]), .Z(n3134) );
  AND U9501 ( .A(n3135), .B(\SUBBYTES[1].a/w1402 ), .Z(\SUBBYTES[1].a/w1537 )
         );
  AND U9502 ( .A(n3136), .B(\SUBBYTES[1].a/w1403 ), .Z(\SUBBYTES[1].a/w1535 )
         );
  AND U9503 ( .A(\SUBBYTES[1].a/w1533 ), .B(n3137), .Z(\SUBBYTES[1].a/w1534 )
         );
  ANDN U9504 ( .A(\w1[1][72] ), .B(n3138), .Z(\SUBBYTES[1].a/w1530 ) );
  AND U9505 ( .A(n3139), .B(\SUBBYTES[1].a/w1405 ), .Z(\SUBBYTES[1].a/w1528 )
         );
  AND U9506 ( .A(\SUBBYTES[1].a/w1526 ), .B(n3140), .Z(\SUBBYTES[1].a/w1527 )
         );
  XOR U9507 ( .A(\SUBBYTES[1].a/w1470 ), .B(n5844), .Z(n3140) );
  AND U9508 ( .A(\SUBBYTES[1].a/w1513 ), .B(\SUBBYTES[1].a/w1515 ), .Z(
        \SUBBYTES[1].a/w1522 ) );
  AND U9509 ( .A(\SUBBYTES[1].a/w1514 ), .B(\SUBBYTES[1].a/w1516 ), .Z(
        \SUBBYTES[1].a/w1520 ) );
  AND U9510 ( .A(\SUBBYTES[1].a/w1517 ), .B(\SUBBYTES[1].a/w1518 ), .Z(
        \SUBBYTES[1].a/w1519 ) );
  AND U9511 ( .A(\SUBBYTES[1].a/w1406 ), .B(n3135), .Z(\SUBBYTES[1].a/w1505 )
         );
  XOR U9512 ( .A(\SUBBYTES[1].a/w1474 ), .B(n963), .Z(n3135) );
  AND U9513 ( .A(\SUBBYTES[1].a/w1407 ), .B(n3136), .Z(\SUBBYTES[1].a/w1503 )
         );
  XOR U9514 ( .A(n5845), .B(\SUBBYTES[1].a/w1474 ), .Z(n3136) );
  ANDN U9515 ( .A(n3137), .B(n3141), .Z(\SUBBYTES[1].a/w1502 ) );
  XOR U9516 ( .A(n963), .B(n5845), .Z(n3137) );
  ANDN U9517 ( .A(\SUBBYTES[1].a/w1408 ), .B(n3138), .Z(\SUBBYTES[1].a/w1498 )
         );
  XNOR U9518 ( .A(\SUBBYTES[1].a/w1467 ), .B(\SUBBYTES[1].a/w1470 ), .Z(n3138)
         );
  AND U9519 ( .A(\SUBBYTES[1].a/w1409 ), .B(n3139), .Z(\SUBBYTES[1].a/w1496 )
         );
  XNOR U9520 ( .A(n3142), .B(\SUBBYTES[1].a/w1467 ), .Z(n3139) );
  AND U9521 ( .A(\SUBBYTES[1].a/w1494 ), .B(n3143), .Z(\SUBBYTES[1].a/w1495 )
         );
  XOR U9522 ( .A(n3144), .B(n3142), .Z(n3143) );
  IV U9523 ( .A(n5844), .Z(n3142) );
  ANDN U9524 ( .A(\SUBBYTES[1].a/w1513 ), .B(n3145), .Z(\SUBBYTES[1].a/w1490 )
         );
  ANDN U9525 ( .A(\SUBBYTES[1].a/w1514 ), .B(n3146), .Z(\SUBBYTES[1].a/w1488 )
         );
  ANDN U9526 ( .A(\SUBBYTES[1].a/w1517 ), .B(n3147), .Z(\SUBBYTES[1].a/w1487 )
         );
  AND U9527 ( .A(\SUBBYTES[1].a/w1473 ), .B(\SUBBYTES[1].a/w1472 ), .Z(
        \SUBBYTES[1].a/w1474 ) );
  IV U9528 ( .A(n3144), .Z(\SUBBYTES[1].a/w1470 ) );
  NAND U9529 ( .A(\SUBBYTES[1].a/w1449 ), .B(\SUBBYTES[1].a/w1464 ), .Z(n3144)
         );
  AND U9530 ( .A(\SUBBYTES[1].a/w1466 ), .B(\SUBBYTES[1].a/w1472 ), .Z(
        \SUBBYTES[1].a/w1467 ) );
  AND U9531 ( .A(\SUBBYTES[1].a/w1451 ), .B(\SUBBYTES[1].a/w1449 ), .Z(
        \SUBBYTES[1].a/w1461 ) );
  AND U9532 ( .A(\SUBBYTES[1].a/w1452 ), .B(\SUBBYTES[1].a/w1450 ), .Z(
        \SUBBYTES[1].a/w1459 ) );
  AND U9533 ( .A(\SUBBYTES[1].a/w1466 ), .B(\SUBBYTES[1].a/w1473 ), .Z(
        \SUBBYTES[1].a/w1458 ) );
  AND U9534 ( .A(\SUBBYTES[1].a/w1406 ), .B(\SUBBYTES[1].a/w1402 ), .Z(
        \SUBBYTES[1].a/w1443 ) );
  AND U9535 ( .A(\SUBBYTES[1].a/w1407 ), .B(\SUBBYTES[1].a/w1403 ), .Z(
        \SUBBYTES[1].a/w1441 ) );
  ANDN U9536 ( .A(\SUBBYTES[1].a/w1533 ), .B(n3141), .Z(\SUBBYTES[1].a/w1440 )
         );
  XNOR U9537 ( .A(\w1[1][73] ), .B(\w1[1][79] ), .Z(n3141) );
  XOR U9538 ( .A(\w0[1][73] ), .B(g_input[201]), .Z(\w1[1][73] ) );
  AND U9539 ( .A(\w1[1][72] ), .B(\SUBBYTES[1].a/w1408 ), .Z(
        \SUBBYTES[1].a/w1436 ) );
  XOR U9540 ( .A(\w0[1][72] ), .B(g_input[200]), .Z(\w1[1][72] ) );
  AND U9541 ( .A(\SUBBYTES[1].a/w1409 ), .B(\SUBBYTES[1].a/w1405 ), .Z(
        \SUBBYTES[1].a/w1434 ) );
  AND U9542 ( .A(\SUBBYTES[1].a/w1494 ), .B(\SUBBYTES[1].a/w1526 ), .Z(
        \SUBBYTES[1].a/w1433 ) );
  ANDN U9543 ( .A(\SUBBYTES[1].a/w1515 ), .B(n3145), .Z(\SUBBYTES[1].a/w1428 )
         );
  XNOR U9544 ( .A(\w1[1][76] ), .B(\w1[1][79] ), .Z(n3145) );
  ANDN U9545 ( .A(\SUBBYTES[1].a/w1516 ), .B(n3146), .Z(\SUBBYTES[1].a/w1426 )
         );
  XNOR U9546 ( .A(\w1[1][74] ), .B(\w1[1][79] ), .Z(n3146) );
  XOR U9547 ( .A(\w0[1][79] ), .B(g_input[207]), .Z(\w1[1][79] ) );
  IV U9548 ( .A(n3148), .Z(\w1[1][74] ) );
  ANDN U9549 ( .A(\SUBBYTES[1].a/w1518 ), .B(n3147), .Z(\SUBBYTES[1].a/w1425 )
         );
  XOR U9550 ( .A(n3148), .B(\w1[1][76] ), .Z(n3147) );
  XOR U9551 ( .A(\w0[1][76] ), .B(g_input[204]), .Z(\w1[1][76] ) );
  XNOR U9552 ( .A(\w0[1][74] ), .B(g_input[202]), .Z(n3148) );
  AND U9553 ( .A(n3149), .B(\SUBBYTES[1].a/w1195 ), .Z(\SUBBYTES[1].a/w1330 )
         );
  AND U9554 ( .A(n3150), .B(\SUBBYTES[1].a/w1196 ), .Z(\SUBBYTES[1].a/w1328 )
         );
  AND U9555 ( .A(\SUBBYTES[1].a/w1326 ), .B(n3151), .Z(\SUBBYTES[1].a/w1327 )
         );
  ANDN U9556 ( .A(\w1[1][80] ), .B(n3152), .Z(\SUBBYTES[1].a/w1323 ) );
  AND U9557 ( .A(n3153), .B(\SUBBYTES[1].a/w1198 ), .Z(\SUBBYTES[1].a/w1321 )
         );
  AND U9558 ( .A(\SUBBYTES[1].a/w1319 ), .B(n3154), .Z(\SUBBYTES[1].a/w1320 )
         );
  XOR U9559 ( .A(\SUBBYTES[1].a/w1263 ), .B(n5842), .Z(n3154) );
  AND U9560 ( .A(\SUBBYTES[1].a/w1306 ), .B(\SUBBYTES[1].a/w1308 ), .Z(
        \SUBBYTES[1].a/w1315 ) );
  AND U9561 ( .A(\SUBBYTES[1].a/w1307 ), .B(\SUBBYTES[1].a/w1309 ), .Z(
        \SUBBYTES[1].a/w1313 ) );
  AND U9562 ( .A(\SUBBYTES[1].a/w1310 ), .B(\SUBBYTES[1].a/w1311 ), .Z(
        \SUBBYTES[1].a/w1312 ) );
  AND U9563 ( .A(\SUBBYTES[1].a/w1199 ), .B(n3149), .Z(\SUBBYTES[1].a/w1298 )
         );
  XOR U9564 ( .A(\SUBBYTES[1].a/w1267 ), .B(n962), .Z(n3149) );
  AND U9565 ( .A(\SUBBYTES[1].a/w1200 ), .B(n3150), .Z(\SUBBYTES[1].a/w1296 )
         );
  XOR U9566 ( .A(n5843), .B(\SUBBYTES[1].a/w1267 ), .Z(n3150) );
  ANDN U9567 ( .A(n3151), .B(n3155), .Z(\SUBBYTES[1].a/w1295 ) );
  XOR U9568 ( .A(n962), .B(n5843), .Z(n3151) );
  ANDN U9569 ( .A(\SUBBYTES[1].a/w1201 ), .B(n3152), .Z(\SUBBYTES[1].a/w1291 )
         );
  XNOR U9570 ( .A(\SUBBYTES[1].a/w1260 ), .B(\SUBBYTES[1].a/w1263 ), .Z(n3152)
         );
  AND U9571 ( .A(\SUBBYTES[1].a/w1202 ), .B(n3153), .Z(\SUBBYTES[1].a/w1289 )
         );
  XNOR U9572 ( .A(n3156), .B(\SUBBYTES[1].a/w1260 ), .Z(n3153) );
  AND U9573 ( .A(\SUBBYTES[1].a/w1287 ), .B(n3157), .Z(\SUBBYTES[1].a/w1288 )
         );
  XOR U9574 ( .A(n3158), .B(n3156), .Z(n3157) );
  IV U9575 ( .A(n5842), .Z(n3156) );
  ANDN U9576 ( .A(\SUBBYTES[1].a/w1306 ), .B(n3159), .Z(\SUBBYTES[1].a/w1283 )
         );
  ANDN U9577 ( .A(\SUBBYTES[1].a/w1307 ), .B(n3160), .Z(\SUBBYTES[1].a/w1281 )
         );
  ANDN U9578 ( .A(\SUBBYTES[1].a/w1310 ), .B(n3161), .Z(\SUBBYTES[1].a/w1280 )
         );
  AND U9579 ( .A(\SUBBYTES[1].a/w1266 ), .B(\SUBBYTES[1].a/w1265 ), .Z(
        \SUBBYTES[1].a/w1267 ) );
  IV U9580 ( .A(n3158), .Z(\SUBBYTES[1].a/w1263 ) );
  NAND U9581 ( .A(\SUBBYTES[1].a/w1242 ), .B(\SUBBYTES[1].a/w1257 ), .Z(n3158)
         );
  AND U9582 ( .A(\SUBBYTES[1].a/w1259 ), .B(\SUBBYTES[1].a/w1265 ), .Z(
        \SUBBYTES[1].a/w1260 ) );
  AND U9583 ( .A(\SUBBYTES[1].a/w1244 ), .B(\SUBBYTES[1].a/w1242 ), .Z(
        \SUBBYTES[1].a/w1254 ) );
  AND U9584 ( .A(\SUBBYTES[1].a/w1245 ), .B(\SUBBYTES[1].a/w1243 ), .Z(
        \SUBBYTES[1].a/w1252 ) );
  AND U9585 ( .A(\SUBBYTES[1].a/w1259 ), .B(\SUBBYTES[1].a/w1266 ), .Z(
        \SUBBYTES[1].a/w1251 ) );
  AND U9586 ( .A(\SUBBYTES[1].a/w1199 ), .B(\SUBBYTES[1].a/w1195 ), .Z(
        \SUBBYTES[1].a/w1236 ) );
  AND U9587 ( .A(\SUBBYTES[1].a/w1200 ), .B(\SUBBYTES[1].a/w1196 ), .Z(
        \SUBBYTES[1].a/w1234 ) );
  ANDN U9588 ( .A(\SUBBYTES[1].a/w1326 ), .B(n3155), .Z(\SUBBYTES[1].a/w1233 )
         );
  XNOR U9589 ( .A(\w1[1][81] ), .B(\w1[1][87] ), .Z(n3155) );
  XOR U9590 ( .A(\w0[1][81] ), .B(g_input[209]), .Z(\w1[1][81] ) );
  AND U9591 ( .A(\w1[1][80] ), .B(\SUBBYTES[1].a/w1201 ), .Z(
        \SUBBYTES[1].a/w1229 ) );
  XOR U9592 ( .A(\w0[1][80] ), .B(g_input[208]), .Z(\w1[1][80] ) );
  AND U9593 ( .A(\SUBBYTES[1].a/w1202 ), .B(\SUBBYTES[1].a/w1198 ), .Z(
        \SUBBYTES[1].a/w1227 ) );
  AND U9594 ( .A(\SUBBYTES[1].a/w1287 ), .B(\SUBBYTES[1].a/w1319 ), .Z(
        \SUBBYTES[1].a/w1226 ) );
  ANDN U9595 ( .A(\SUBBYTES[1].a/w1308 ), .B(n3159), .Z(\SUBBYTES[1].a/w1221 )
         );
  XNOR U9596 ( .A(\w1[1][84] ), .B(\w1[1][87] ), .Z(n3159) );
  ANDN U9597 ( .A(\SUBBYTES[1].a/w1309 ), .B(n3160), .Z(\SUBBYTES[1].a/w1219 )
         );
  XNOR U9598 ( .A(\w1[1][82] ), .B(\w1[1][87] ), .Z(n3160) );
  XOR U9599 ( .A(\w0[1][87] ), .B(g_input[215]), .Z(\w1[1][87] ) );
  IV U9600 ( .A(n3162), .Z(\w1[1][82] ) );
  ANDN U9601 ( .A(\SUBBYTES[1].a/w1311 ), .B(n3161), .Z(\SUBBYTES[1].a/w1218 )
         );
  XOR U9602 ( .A(n3162), .B(\w1[1][84] ), .Z(n3161) );
  XOR U9603 ( .A(\w0[1][84] ), .B(g_input[212]), .Z(\w1[1][84] ) );
  XNOR U9604 ( .A(\w0[1][82] ), .B(g_input[210]), .Z(n3162) );
  AND U9605 ( .A(n3163), .B(\SUBBYTES[1].a/w988 ), .Z(\SUBBYTES[1].a/w1123 )
         );
  AND U9606 ( .A(n3164), .B(\SUBBYTES[1].a/w989 ), .Z(\SUBBYTES[1].a/w1121 )
         );
  AND U9607 ( .A(\SUBBYTES[1].a/w1119 ), .B(n3165), .Z(\SUBBYTES[1].a/w1120 )
         );
  ANDN U9608 ( .A(\w1[1][88] ), .B(n3166), .Z(\SUBBYTES[1].a/w1116 ) );
  AND U9609 ( .A(n3167), .B(\SUBBYTES[1].a/w991 ), .Z(\SUBBYTES[1].a/w1114 )
         );
  AND U9610 ( .A(\SUBBYTES[1].a/w1112 ), .B(n3168), .Z(\SUBBYTES[1].a/w1113 )
         );
  XOR U9611 ( .A(\SUBBYTES[1].a/w1056 ), .B(n5840), .Z(n3168) );
  AND U9612 ( .A(\SUBBYTES[1].a/w1099 ), .B(\SUBBYTES[1].a/w1101 ), .Z(
        \SUBBYTES[1].a/w1108 ) );
  AND U9613 ( .A(\SUBBYTES[1].a/w1100 ), .B(\SUBBYTES[1].a/w1102 ), .Z(
        \SUBBYTES[1].a/w1106 ) );
  AND U9614 ( .A(\SUBBYTES[1].a/w1103 ), .B(\SUBBYTES[1].a/w1104 ), .Z(
        \SUBBYTES[1].a/w1105 ) );
  AND U9615 ( .A(\SUBBYTES[1].a/w992 ), .B(n3163), .Z(\SUBBYTES[1].a/w1091 )
         );
  XOR U9616 ( .A(\SUBBYTES[1].a/w1060 ), .B(n961), .Z(n3163) );
  AND U9617 ( .A(\SUBBYTES[1].a/w993 ), .B(n3164), .Z(\SUBBYTES[1].a/w1089 )
         );
  XOR U9618 ( .A(n5841), .B(\SUBBYTES[1].a/w1060 ), .Z(n3164) );
  ANDN U9619 ( .A(n3165), .B(n3169), .Z(\SUBBYTES[1].a/w1088 ) );
  XOR U9620 ( .A(n961), .B(n5841), .Z(n3165) );
  ANDN U9621 ( .A(\SUBBYTES[1].a/w994 ), .B(n3166), .Z(\SUBBYTES[1].a/w1084 )
         );
  XNOR U9622 ( .A(\SUBBYTES[1].a/w1053 ), .B(\SUBBYTES[1].a/w1056 ), .Z(n3166)
         );
  AND U9623 ( .A(\SUBBYTES[1].a/w995 ), .B(n3167), .Z(\SUBBYTES[1].a/w1082 )
         );
  XNOR U9624 ( .A(n3170), .B(\SUBBYTES[1].a/w1053 ), .Z(n3167) );
  AND U9625 ( .A(\SUBBYTES[1].a/w1080 ), .B(n3171), .Z(\SUBBYTES[1].a/w1081 )
         );
  XOR U9626 ( .A(n3172), .B(n3170), .Z(n3171) );
  IV U9627 ( .A(n5840), .Z(n3170) );
  ANDN U9628 ( .A(\SUBBYTES[1].a/w1099 ), .B(n3173), .Z(\SUBBYTES[1].a/w1076 )
         );
  ANDN U9629 ( .A(\SUBBYTES[1].a/w1100 ), .B(n3174), .Z(\SUBBYTES[1].a/w1074 )
         );
  ANDN U9630 ( .A(\SUBBYTES[1].a/w1103 ), .B(n3175), .Z(\SUBBYTES[1].a/w1073 )
         );
  AND U9631 ( .A(\SUBBYTES[1].a/w1059 ), .B(\SUBBYTES[1].a/w1058 ), .Z(
        \SUBBYTES[1].a/w1060 ) );
  IV U9632 ( .A(n3172), .Z(\SUBBYTES[1].a/w1056 ) );
  NAND U9633 ( .A(\SUBBYTES[1].a/w1035 ), .B(\SUBBYTES[1].a/w1050 ), .Z(n3172)
         );
  AND U9634 ( .A(\SUBBYTES[1].a/w1052 ), .B(\SUBBYTES[1].a/w1058 ), .Z(
        \SUBBYTES[1].a/w1053 ) );
  AND U9635 ( .A(\SUBBYTES[1].a/w1037 ), .B(\SUBBYTES[1].a/w1035 ), .Z(
        \SUBBYTES[1].a/w1047 ) );
  AND U9636 ( .A(\SUBBYTES[1].a/w1038 ), .B(\SUBBYTES[1].a/w1036 ), .Z(
        \SUBBYTES[1].a/w1045 ) );
  AND U9637 ( .A(\SUBBYTES[1].a/w1052 ), .B(\SUBBYTES[1].a/w1059 ), .Z(
        \SUBBYTES[1].a/w1044 ) );
  AND U9638 ( .A(\SUBBYTES[1].a/w992 ), .B(\SUBBYTES[1].a/w988 ), .Z(
        \SUBBYTES[1].a/w1029 ) );
  AND U9639 ( .A(\SUBBYTES[1].a/w993 ), .B(\SUBBYTES[1].a/w989 ), .Z(
        \SUBBYTES[1].a/w1027 ) );
  ANDN U9640 ( .A(\SUBBYTES[1].a/w1119 ), .B(n3169), .Z(\SUBBYTES[1].a/w1026 )
         );
  XNOR U9641 ( .A(\w1[1][89] ), .B(\w1[1][95] ), .Z(n3169) );
  XOR U9642 ( .A(\w0[1][89] ), .B(g_input[217]), .Z(\w1[1][89] ) );
  AND U9643 ( .A(\w1[1][88] ), .B(\SUBBYTES[1].a/w994 ), .Z(
        \SUBBYTES[1].a/w1022 ) );
  XOR U9644 ( .A(\w0[1][88] ), .B(g_input[216]), .Z(\w1[1][88] ) );
  AND U9645 ( .A(\SUBBYTES[1].a/w995 ), .B(\SUBBYTES[1].a/w991 ), .Z(
        \SUBBYTES[1].a/w1020 ) );
  AND U9646 ( .A(\SUBBYTES[1].a/w1080 ), .B(\SUBBYTES[1].a/w1112 ), .Z(
        \SUBBYTES[1].a/w1019 ) );
  ANDN U9647 ( .A(\SUBBYTES[1].a/w1101 ), .B(n3173), .Z(\SUBBYTES[1].a/w1014 )
         );
  XNOR U9648 ( .A(\w1[1][92] ), .B(\w1[1][95] ), .Z(n3173) );
  ANDN U9649 ( .A(\SUBBYTES[1].a/w1102 ), .B(n3174), .Z(\SUBBYTES[1].a/w1012 )
         );
  XNOR U9650 ( .A(\w1[1][90] ), .B(\w1[1][95] ), .Z(n3174) );
  XOR U9651 ( .A(\w0[1][95] ), .B(g_input[223]), .Z(\w1[1][95] ) );
  IV U9652 ( .A(n3176), .Z(\w1[1][90] ) );
  ANDN U9653 ( .A(\SUBBYTES[1].a/w1104 ), .B(n3175), .Z(\SUBBYTES[1].a/w1011 )
         );
  XOR U9654 ( .A(n3176), .B(\w1[1][92] ), .Z(n3175) );
  XOR U9655 ( .A(\w0[1][92] ), .B(g_input[220]), .Z(\w1[1][92] ) );
  XNOR U9656 ( .A(\w0[1][90] ), .B(g_input[218]), .Z(n3176) );
  AND U9657 ( .A(\SUBBYTES[1].a/w2084 ), .B(\SUBBYTES[1].a/w2071 ), .Z(n5850)
         );
  AND U9658 ( .A(\SUBBYTES[1].a/w1877 ), .B(\SUBBYTES[1].a/w1866 ), .Z(n5849)
         );
  AND U9659 ( .A(\SUBBYTES[1].a/w221 ), .B(\SUBBYTES[1].a/w208 ), .Z(n5832) );
  AND U9660 ( .A(\SUBBYTES[1].a/w1877 ), .B(\SUBBYTES[1].a/w1864 ), .Z(n5848)
         );
  AND U9661 ( .A(\SUBBYTES[1].a/w1670 ), .B(\SUBBYTES[1].a/w1659 ), .Z(n5847)
         );
  AND U9662 ( .A(\SUBBYTES[1].a/w1670 ), .B(\SUBBYTES[1].a/w1657 ), .Z(n5846)
         );
  AND U9663 ( .A(\SUBBYTES[1].a/w1463 ), .B(\SUBBYTES[1].a/w1452 ), .Z(n5845)
         );
  AND U9664 ( .A(\SUBBYTES[1].a/w1463 ), .B(\SUBBYTES[1].a/w1450 ), .Z(n5844)
         );
  AND U9665 ( .A(\SUBBYTES[1].a/w1256 ), .B(\SUBBYTES[1].a/w1245 ), .Z(n5843)
         );
  AND U9666 ( .A(\SUBBYTES[1].a/w1256 ), .B(\SUBBYTES[1].a/w1243 ), .Z(n5842)
         );
  AND U9667 ( .A(\SUBBYTES[1].a/w1049 ), .B(\SUBBYTES[1].a/w1038 ), .Z(n5841)
         );
  AND U9668 ( .A(\SUBBYTES[1].a/w1049 ), .B(\SUBBYTES[1].a/w1036 ), .Z(n5840)
         );
  AND U9669 ( .A(\SUBBYTES[1].a/w842 ), .B(\SUBBYTES[1].a/w831 ), .Z(n5839) );
  AND U9670 ( .A(\SUBBYTES[1].a/w842 ), .B(\SUBBYTES[1].a/w829 ), .Z(n5838) );
  AND U9671 ( .A(\SUBBYTES[1].a/w635 ), .B(\SUBBYTES[1].a/w624 ), .Z(n5837) );
  AND U9672 ( .A(\SUBBYTES[1].a/w635 ), .B(\SUBBYTES[1].a/w622 ), .Z(n5836) );
  AND U9673 ( .A(\SUBBYTES[1].a/w428 ), .B(\SUBBYTES[1].a/w417 ), .Z(n5835) );
  AND U9674 ( .A(\SUBBYTES[1].a/w428 ), .B(\SUBBYTES[1].a/w415 ), .Z(n5834) );
  AND U9675 ( .A(\SUBBYTES[1].a/w3326 ), .B(\SUBBYTES[1].a/w3315 ), .Z(n5863)
         );
  AND U9676 ( .A(\SUBBYTES[1].a/w3326 ), .B(\SUBBYTES[1].a/w3313 ), .Z(n5862)
         );
  AND U9677 ( .A(\SUBBYTES[1].a/w3119 ), .B(\SUBBYTES[1].a/w3108 ), .Z(n5861)
         );
  AND U9678 ( .A(\SUBBYTES[1].a/w3119 ), .B(\SUBBYTES[1].a/w3106 ), .Z(n5860)
         );
  AND U9679 ( .A(\SUBBYTES[1].a/w2912 ), .B(\SUBBYTES[1].a/w2901 ), .Z(n5859)
         );
  AND U9680 ( .A(\SUBBYTES[1].a/w2912 ), .B(\SUBBYTES[1].a/w2899 ), .Z(n5858)
         );
  AND U9681 ( .A(\SUBBYTES[1].a/w2705 ), .B(\SUBBYTES[1].a/w2694 ), .Z(n5857)
         );
  AND U9682 ( .A(\SUBBYTES[1].a/w2705 ), .B(\SUBBYTES[1].a/w2692 ), .Z(n5856)
         );
  AND U9683 ( .A(\SUBBYTES[1].a/w2498 ), .B(\SUBBYTES[1].a/w2487 ), .Z(n5855)
         );
  AND U9684 ( .A(\SUBBYTES[1].a/w2498 ), .B(\SUBBYTES[1].a/w2485 ), .Z(n5854)
         );
  AND U9685 ( .A(\SUBBYTES[1].a/w2291 ), .B(\SUBBYTES[1].a/w2280 ), .Z(n5853)
         );
  AND U9686 ( .A(\SUBBYTES[1].a/w2291 ), .B(\SUBBYTES[1].a/w2278 ), .Z(n5852)
         );
  AND U9687 ( .A(\SUBBYTES[1].a/w2084 ), .B(\SUBBYTES[1].a/w2073 ), .Z(n5851)
         );
  AND U9688 ( .A(\SUBBYTES[1].a/w221 ), .B(\SUBBYTES[1].a/w210 ), .Z(n5833) );
  AND U9689 ( .A(n3177), .B(\SUBBYTES[0].a/w781 ), .Z(\SUBBYTES[0].a/w916 ) );
  AND U9690 ( .A(n3178), .B(\SUBBYTES[0].a/w782 ), .Z(\SUBBYTES[0].a/w914 ) );
  AND U9691 ( .A(\SUBBYTES[0].a/w912 ), .B(n3179), .Z(\SUBBYTES[0].a/w913 ) );
  ANDN U9692 ( .A(\w1[0][96] ), .B(n3180), .Z(\SUBBYTES[0].a/w909 ) );
  AND U9693 ( .A(n3181), .B(\SUBBYTES[0].a/w784 ), .Z(\SUBBYTES[0].a/w907 ) );
  AND U9694 ( .A(\SUBBYTES[0].a/w905 ), .B(n3182), .Z(\SUBBYTES[0].a/w906 ) );
  XOR U9695 ( .A(\SUBBYTES[0].a/w849 ), .B(\SUBBYTES[0].a/n39 ), .Z(n3182) );
  AND U9696 ( .A(\SUBBYTES[0].a/w892 ), .B(\SUBBYTES[0].a/w894 ), .Z(
        \SUBBYTES[0].a/w901 ) );
  AND U9697 ( .A(\SUBBYTES[0].a/w893 ), .B(\SUBBYTES[0].a/w895 ), .Z(
        \SUBBYTES[0].a/w899 ) );
  AND U9698 ( .A(\SUBBYTES[0].a/w896 ), .B(\SUBBYTES[0].a/w897 ), .Z(
        \SUBBYTES[0].a/w898 ) );
  AND U9699 ( .A(\SUBBYTES[0].a/w785 ), .B(n3177), .Z(\SUBBYTES[0].a/w884 ) );
  XOR U9700 ( .A(\SUBBYTES[0].a/w853 ), .B(n1156), .Z(n3177) );
  AND U9701 ( .A(\SUBBYTES[0].a/w786 ), .B(n3178), .Z(\SUBBYTES[0].a/w882 ) );
  XOR U9702 ( .A(\SUBBYTES[0].a/n40 ), .B(\SUBBYTES[0].a/w853 ), .Z(n3178) );
  ANDN U9703 ( .A(n3179), .B(n3183), .Z(\SUBBYTES[0].a/w881 ) );
  XOR U9704 ( .A(n1156), .B(\SUBBYTES[0].a/n40 ), .Z(n3179) );
  ANDN U9705 ( .A(\SUBBYTES[0].a/w787 ), .B(n3180), .Z(\SUBBYTES[0].a/w877 )
         );
  XNOR U9706 ( .A(\SUBBYTES[0].a/w846 ), .B(\SUBBYTES[0].a/w849 ), .Z(n3180)
         );
  AND U9707 ( .A(\SUBBYTES[0].a/w788 ), .B(n3181), .Z(\SUBBYTES[0].a/w875 ) );
  XNOR U9708 ( .A(n3184), .B(\SUBBYTES[0].a/w846 ), .Z(n3181) );
  AND U9709 ( .A(\SUBBYTES[0].a/w873 ), .B(n3185), .Z(\SUBBYTES[0].a/w874 ) );
  XOR U9710 ( .A(n3186), .B(n3184), .Z(n3185) );
  IV U9711 ( .A(\SUBBYTES[0].a/n39 ), .Z(n3184) );
  ANDN U9712 ( .A(\SUBBYTES[0].a/w892 ), .B(n3187), .Z(\SUBBYTES[0].a/w869 )
         );
  ANDN U9713 ( .A(\SUBBYTES[0].a/w893 ), .B(n3188), .Z(\SUBBYTES[0].a/w867 )
         );
  ANDN U9714 ( .A(\SUBBYTES[0].a/w896 ), .B(n3189), .Z(\SUBBYTES[0].a/w866 )
         );
  AND U9715 ( .A(\SUBBYTES[0].a/w852 ), .B(\SUBBYTES[0].a/w851 ), .Z(
        \SUBBYTES[0].a/w853 ) );
  IV U9716 ( .A(n3186), .Z(\SUBBYTES[0].a/w849 ) );
  NAND U9717 ( .A(\SUBBYTES[0].a/w828 ), .B(\SUBBYTES[0].a/w843 ), .Z(n3186)
         );
  AND U9718 ( .A(\SUBBYTES[0].a/w845 ), .B(\SUBBYTES[0].a/w851 ), .Z(
        \SUBBYTES[0].a/w846 ) );
  AND U9719 ( .A(\SUBBYTES[0].a/w830 ), .B(\SUBBYTES[0].a/w828 ), .Z(
        \SUBBYTES[0].a/w840 ) );
  AND U9720 ( .A(\SUBBYTES[0].a/w831 ), .B(\SUBBYTES[0].a/w829 ), .Z(
        \SUBBYTES[0].a/w838 ) );
  AND U9721 ( .A(\SUBBYTES[0].a/w845 ), .B(\SUBBYTES[0].a/w852 ), .Z(
        \SUBBYTES[0].a/w837 ) );
  AND U9722 ( .A(\SUBBYTES[0].a/w785 ), .B(\SUBBYTES[0].a/w781 ), .Z(
        \SUBBYTES[0].a/w822 ) );
  AND U9723 ( .A(\SUBBYTES[0].a/w786 ), .B(\SUBBYTES[0].a/w782 ), .Z(
        \SUBBYTES[0].a/w820 ) );
  ANDN U9724 ( .A(\SUBBYTES[0].a/w912 ), .B(n3183), .Z(\SUBBYTES[0].a/w819 )
         );
  XNOR U9725 ( .A(\w1[0][103] ), .B(\w1[0][97] ), .Z(n3183) );
  XOR U9726 ( .A(g_input[97]), .B(e_input[97]), .Z(\w1[0][97] ) );
  IV U9727 ( .A(n3190), .Z(\w1[0][103] ) );
  AND U9728 ( .A(\w1[0][96] ), .B(\SUBBYTES[0].a/w787 ), .Z(
        \SUBBYTES[0].a/w815 ) );
  XOR U9729 ( .A(g_input[96]), .B(e_input[96]), .Z(\w1[0][96] ) );
  AND U9730 ( .A(\SUBBYTES[0].a/w788 ), .B(\SUBBYTES[0].a/w784 ), .Z(
        \SUBBYTES[0].a/w813 ) );
  AND U9731 ( .A(\SUBBYTES[0].a/w873 ), .B(\SUBBYTES[0].a/w905 ), .Z(
        \SUBBYTES[0].a/w812 ) );
  ANDN U9732 ( .A(\SUBBYTES[0].a/w894 ), .B(n3187), .Z(\SUBBYTES[0].a/w807 )
         );
  XOR U9733 ( .A(\w1[0][100] ), .B(n3190), .Z(n3187) );
  ANDN U9734 ( .A(\SUBBYTES[0].a/w895 ), .B(n3188), .Z(\SUBBYTES[0].a/w805 )
         );
  XOR U9735 ( .A(n3190), .B(\w1[0][98] ), .Z(n3188) );
  XNOR U9736 ( .A(g_input[103]), .B(e_input[103]), .Z(n3190) );
  ANDN U9737 ( .A(\SUBBYTES[0].a/w897 ), .B(n3189), .Z(\SUBBYTES[0].a/w804 )
         );
  XNOR U9738 ( .A(\w1[0][100] ), .B(\w1[0][98] ), .Z(n3189) );
  XOR U9739 ( .A(g_input[98]), .B(e_input[98]), .Z(\w1[0][98] ) );
  XOR U9740 ( .A(g_input[100]), .B(e_input[100]), .Z(\w1[0][100] ) );
  AND U9741 ( .A(n3191), .B(\SUBBYTES[0].a/w574 ), .Z(\SUBBYTES[0].a/w709 ) );
  AND U9742 ( .A(n3192), .B(\SUBBYTES[0].a/w575 ), .Z(\SUBBYTES[0].a/w707 ) );
  AND U9743 ( .A(\SUBBYTES[0].a/w705 ), .B(n3193), .Z(\SUBBYTES[0].a/w706 ) );
  ANDN U9744 ( .A(\w1[0][104] ), .B(n3194), .Z(\SUBBYTES[0].a/w702 ) );
  AND U9745 ( .A(n3195), .B(\SUBBYTES[0].a/w577 ), .Z(\SUBBYTES[0].a/w700 ) );
  AND U9746 ( .A(\SUBBYTES[0].a/w698 ), .B(n3196), .Z(\SUBBYTES[0].a/w699 ) );
  XOR U9747 ( .A(\SUBBYTES[0].a/w642 ), .B(\SUBBYTES[0].a/n29 ), .Z(n3196) );
  AND U9748 ( .A(\SUBBYTES[0].a/w685 ), .B(\SUBBYTES[0].a/w687 ), .Z(
        \SUBBYTES[0].a/w694 ) );
  AND U9749 ( .A(\SUBBYTES[0].a/w686 ), .B(\SUBBYTES[0].a/w688 ), .Z(
        \SUBBYTES[0].a/w692 ) );
  AND U9750 ( .A(\SUBBYTES[0].a/w689 ), .B(\SUBBYTES[0].a/w690 ), .Z(
        \SUBBYTES[0].a/w691 ) );
  AND U9751 ( .A(\SUBBYTES[0].a/w578 ), .B(n3191), .Z(\SUBBYTES[0].a/w677 ) );
  XOR U9752 ( .A(\SUBBYTES[0].a/w646 ), .B(n1155), .Z(n3191) );
  AND U9753 ( .A(\SUBBYTES[0].a/w579 ), .B(n3192), .Z(\SUBBYTES[0].a/w675 ) );
  XOR U9754 ( .A(\SUBBYTES[0].a/n30 ), .B(\SUBBYTES[0].a/w646 ), .Z(n3192) );
  ANDN U9755 ( .A(n3193), .B(n3197), .Z(\SUBBYTES[0].a/w674 ) );
  XOR U9756 ( .A(n1155), .B(\SUBBYTES[0].a/n30 ), .Z(n3193) );
  ANDN U9757 ( .A(\SUBBYTES[0].a/w580 ), .B(n3194), .Z(\SUBBYTES[0].a/w670 )
         );
  XNOR U9758 ( .A(\SUBBYTES[0].a/w639 ), .B(\SUBBYTES[0].a/w642 ), .Z(n3194)
         );
  AND U9759 ( .A(\SUBBYTES[0].a/w581 ), .B(n3195), .Z(\SUBBYTES[0].a/w668 ) );
  XNOR U9760 ( .A(n3198), .B(\SUBBYTES[0].a/w639 ), .Z(n3195) );
  AND U9761 ( .A(\SUBBYTES[0].a/w666 ), .B(n3199), .Z(\SUBBYTES[0].a/w667 ) );
  XOR U9762 ( .A(n3200), .B(n3198), .Z(n3199) );
  IV U9763 ( .A(\SUBBYTES[0].a/n29 ), .Z(n3198) );
  ANDN U9764 ( .A(\SUBBYTES[0].a/w685 ), .B(n3201), .Z(\SUBBYTES[0].a/w662 )
         );
  ANDN U9765 ( .A(\SUBBYTES[0].a/w686 ), .B(n3202), .Z(\SUBBYTES[0].a/w660 )
         );
  ANDN U9766 ( .A(\SUBBYTES[0].a/w689 ), .B(n3203), .Z(\SUBBYTES[0].a/w659 )
         );
  AND U9767 ( .A(\SUBBYTES[0].a/w645 ), .B(\SUBBYTES[0].a/w644 ), .Z(
        \SUBBYTES[0].a/w646 ) );
  IV U9768 ( .A(n3200), .Z(\SUBBYTES[0].a/w642 ) );
  NAND U9769 ( .A(\SUBBYTES[0].a/w621 ), .B(\SUBBYTES[0].a/w636 ), .Z(n3200)
         );
  AND U9770 ( .A(\SUBBYTES[0].a/w638 ), .B(\SUBBYTES[0].a/w644 ), .Z(
        \SUBBYTES[0].a/w639 ) );
  AND U9771 ( .A(\SUBBYTES[0].a/w623 ), .B(\SUBBYTES[0].a/w621 ), .Z(
        \SUBBYTES[0].a/w633 ) );
  AND U9772 ( .A(\SUBBYTES[0].a/w624 ), .B(\SUBBYTES[0].a/w622 ), .Z(
        \SUBBYTES[0].a/w631 ) );
  AND U9773 ( .A(\SUBBYTES[0].a/w638 ), .B(\SUBBYTES[0].a/w645 ), .Z(
        \SUBBYTES[0].a/w630 ) );
  AND U9774 ( .A(\SUBBYTES[0].a/w578 ), .B(\SUBBYTES[0].a/w574 ), .Z(
        \SUBBYTES[0].a/w615 ) );
  AND U9775 ( .A(\SUBBYTES[0].a/w579 ), .B(\SUBBYTES[0].a/w575 ), .Z(
        \SUBBYTES[0].a/w613 ) );
  ANDN U9776 ( .A(\SUBBYTES[0].a/w705 ), .B(n3197), .Z(\SUBBYTES[0].a/w612 )
         );
  XNOR U9777 ( .A(\w1[0][105] ), .B(\w1[0][111] ), .Z(n3197) );
  XOR U9778 ( .A(g_input[105]), .B(e_input[105]), .Z(\w1[0][105] ) );
  AND U9779 ( .A(\w1[0][104] ), .B(\SUBBYTES[0].a/w580 ), .Z(
        \SUBBYTES[0].a/w608 ) );
  XOR U9780 ( .A(g_input[104]), .B(e_input[104]), .Z(\w1[0][104] ) );
  AND U9781 ( .A(\SUBBYTES[0].a/w581 ), .B(\SUBBYTES[0].a/w577 ), .Z(
        \SUBBYTES[0].a/w606 ) );
  AND U9782 ( .A(\SUBBYTES[0].a/w666 ), .B(\SUBBYTES[0].a/w698 ), .Z(
        \SUBBYTES[0].a/w605 ) );
  ANDN U9783 ( .A(\SUBBYTES[0].a/w687 ), .B(n3201), .Z(\SUBBYTES[0].a/w600 )
         );
  XNOR U9784 ( .A(\w1[0][108] ), .B(\w1[0][111] ), .Z(n3201) );
  ANDN U9785 ( .A(\SUBBYTES[0].a/w688 ), .B(n3202), .Z(\SUBBYTES[0].a/w598 )
         );
  XNOR U9786 ( .A(\w1[0][106] ), .B(\w1[0][111] ), .Z(n3202) );
  XOR U9787 ( .A(g_input[111]), .B(e_input[111]), .Z(\w1[0][111] ) );
  IV U9788 ( .A(n3204), .Z(\w1[0][106] ) );
  ANDN U9789 ( .A(\SUBBYTES[0].a/w690 ), .B(n3203), .Z(\SUBBYTES[0].a/w597 )
         );
  XOR U9790 ( .A(n3204), .B(\w1[0][108] ), .Z(n3203) );
  XOR U9791 ( .A(g_input[108]), .B(e_input[108]), .Z(\w1[0][108] ) );
  XNOR U9792 ( .A(g_input[106]), .B(e_input[106]), .Z(n3204) );
  AND U9793 ( .A(n3205), .B(\SUBBYTES[0].a/w367 ), .Z(\SUBBYTES[0].a/w502 ) );
  AND U9794 ( .A(n3206), .B(\SUBBYTES[0].a/w368 ), .Z(\SUBBYTES[0].a/w500 ) );
  AND U9795 ( .A(\SUBBYTES[0].a/w498 ), .B(n3207), .Z(\SUBBYTES[0].a/w499 ) );
  ANDN U9796 ( .A(\w1[0][112] ), .B(n3208), .Z(\SUBBYTES[0].a/w495 ) );
  AND U9797 ( .A(n3209), .B(\SUBBYTES[0].a/w370 ), .Z(\SUBBYTES[0].a/w493 ) );
  AND U9798 ( .A(\SUBBYTES[0].a/w491 ), .B(n3210), .Z(\SUBBYTES[0].a/w492 ) );
  XOR U9799 ( .A(\SUBBYTES[0].a/w435 ), .B(\SUBBYTES[0].a/n19 ), .Z(n3210) );
  AND U9800 ( .A(\SUBBYTES[0].a/w478 ), .B(\SUBBYTES[0].a/w480 ), .Z(
        \SUBBYTES[0].a/w487 ) );
  AND U9801 ( .A(\SUBBYTES[0].a/w479 ), .B(\SUBBYTES[0].a/w481 ), .Z(
        \SUBBYTES[0].a/w485 ) );
  AND U9802 ( .A(\SUBBYTES[0].a/w482 ), .B(\SUBBYTES[0].a/w483 ), .Z(
        \SUBBYTES[0].a/w484 ) );
  AND U9803 ( .A(\SUBBYTES[0].a/w371 ), .B(n3205), .Z(\SUBBYTES[0].a/w470 ) );
  XOR U9804 ( .A(\SUBBYTES[0].a/w439 ), .B(n1154), .Z(n3205) );
  AND U9805 ( .A(\SUBBYTES[0].a/w372 ), .B(n3206), .Z(\SUBBYTES[0].a/w468 ) );
  XOR U9806 ( .A(\SUBBYTES[0].a/n20 ), .B(\SUBBYTES[0].a/w439 ), .Z(n3206) );
  ANDN U9807 ( .A(n3207), .B(n3211), .Z(\SUBBYTES[0].a/w467 ) );
  XOR U9808 ( .A(n1154), .B(\SUBBYTES[0].a/n20 ), .Z(n3207) );
  ANDN U9809 ( .A(\SUBBYTES[0].a/w373 ), .B(n3208), .Z(\SUBBYTES[0].a/w463 )
         );
  XNOR U9810 ( .A(\SUBBYTES[0].a/w432 ), .B(\SUBBYTES[0].a/w435 ), .Z(n3208)
         );
  AND U9811 ( .A(\SUBBYTES[0].a/w374 ), .B(n3209), .Z(\SUBBYTES[0].a/w461 ) );
  XNOR U9812 ( .A(n3212), .B(\SUBBYTES[0].a/w432 ), .Z(n3209) );
  AND U9813 ( .A(\SUBBYTES[0].a/w459 ), .B(n3213), .Z(\SUBBYTES[0].a/w460 ) );
  XOR U9814 ( .A(n3214), .B(n3212), .Z(n3213) );
  IV U9815 ( .A(\SUBBYTES[0].a/n19 ), .Z(n3212) );
  ANDN U9816 ( .A(\SUBBYTES[0].a/w478 ), .B(n3215), .Z(\SUBBYTES[0].a/w455 )
         );
  ANDN U9817 ( .A(\SUBBYTES[0].a/w479 ), .B(n3216), .Z(\SUBBYTES[0].a/w453 )
         );
  ANDN U9818 ( .A(\SUBBYTES[0].a/w482 ), .B(n3217), .Z(\SUBBYTES[0].a/w452 )
         );
  AND U9819 ( .A(\SUBBYTES[0].a/w438 ), .B(\SUBBYTES[0].a/w437 ), .Z(
        \SUBBYTES[0].a/w439 ) );
  IV U9820 ( .A(n3214), .Z(\SUBBYTES[0].a/w435 ) );
  NAND U9821 ( .A(\SUBBYTES[0].a/w414 ), .B(\SUBBYTES[0].a/w429 ), .Z(n3214)
         );
  AND U9822 ( .A(\SUBBYTES[0].a/w431 ), .B(\SUBBYTES[0].a/w437 ), .Z(
        \SUBBYTES[0].a/w432 ) );
  AND U9823 ( .A(\SUBBYTES[0].a/w416 ), .B(\SUBBYTES[0].a/w414 ), .Z(
        \SUBBYTES[0].a/w426 ) );
  AND U9824 ( .A(\SUBBYTES[0].a/w417 ), .B(\SUBBYTES[0].a/w415 ), .Z(
        \SUBBYTES[0].a/w424 ) );
  AND U9825 ( .A(\SUBBYTES[0].a/w431 ), .B(\SUBBYTES[0].a/w438 ), .Z(
        \SUBBYTES[0].a/w423 ) );
  AND U9826 ( .A(\SUBBYTES[0].a/w371 ), .B(\SUBBYTES[0].a/w367 ), .Z(
        \SUBBYTES[0].a/w408 ) );
  AND U9827 ( .A(\SUBBYTES[0].a/w372 ), .B(\SUBBYTES[0].a/w368 ), .Z(
        \SUBBYTES[0].a/w406 ) );
  ANDN U9828 ( .A(\SUBBYTES[0].a/w498 ), .B(n3211), .Z(\SUBBYTES[0].a/w405 )
         );
  XNOR U9829 ( .A(\w1[0][113] ), .B(\w1[0][119] ), .Z(n3211) );
  XOR U9830 ( .A(g_input[113]), .B(e_input[113]), .Z(\w1[0][113] ) );
  AND U9831 ( .A(\w1[0][112] ), .B(\SUBBYTES[0].a/w373 ), .Z(
        \SUBBYTES[0].a/w401 ) );
  XOR U9832 ( .A(g_input[112]), .B(e_input[112]), .Z(\w1[0][112] ) );
  AND U9833 ( .A(\SUBBYTES[0].a/w374 ), .B(\SUBBYTES[0].a/w370 ), .Z(
        \SUBBYTES[0].a/w399 ) );
  AND U9834 ( .A(\SUBBYTES[0].a/w459 ), .B(\SUBBYTES[0].a/w491 ), .Z(
        \SUBBYTES[0].a/w398 ) );
  ANDN U9835 ( .A(\SUBBYTES[0].a/w480 ), .B(n3215), .Z(\SUBBYTES[0].a/w393 )
         );
  XNOR U9836 ( .A(\w1[0][116] ), .B(\w1[0][119] ), .Z(n3215) );
  ANDN U9837 ( .A(\SUBBYTES[0].a/w481 ), .B(n3216), .Z(\SUBBYTES[0].a/w391 )
         );
  XNOR U9838 ( .A(\w1[0][114] ), .B(\w1[0][119] ), .Z(n3216) );
  XOR U9839 ( .A(g_input[119]), .B(e_input[119]), .Z(\w1[0][119] ) );
  IV U9840 ( .A(n3218), .Z(\w1[0][114] ) );
  ANDN U9841 ( .A(\SUBBYTES[0].a/w483 ), .B(n3217), .Z(\SUBBYTES[0].a/w390 )
         );
  XOR U9842 ( .A(n3218), .B(\w1[0][116] ), .Z(n3217) );
  XOR U9843 ( .A(g_input[116]), .B(e_input[116]), .Z(\w1[0][116] ) );
  XNOR U9844 ( .A(g_input[114]), .B(e_input[114]), .Z(n3218) );
  AND U9845 ( .A(n3219), .B(\SUBBYTES[0].a/w3265 ), .Z(\SUBBYTES[0].a/w3400 )
         );
  AND U9846 ( .A(n3220), .B(\SUBBYTES[0].a/w3266 ), .Z(\SUBBYTES[0].a/w3398 )
         );
  AND U9847 ( .A(\SUBBYTES[0].a/w3396 ), .B(n3221), .Z(\SUBBYTES[0].a/w3397 )
         );
  ANDN U9848 ( .A(\w1[0][0] ), .B(n3222), .Z(\SUBBYTES[0].a/w3393 ) );
  AND U9849 ( .A(n3223), .B(\SUBBYTES[0].a/w3268 ), .Z(\SUBBYTES[0].a/w3391 )
         );
  AND U9850 ( .A(\SUBBYTES[0].a/w3389 ), .B(n3224), .Z(\SUBBYTES[0].a/w3390 )
         );
  XOR U9851 ( .A(\SUBBYTES[0].a/w3333 ), .B(\SUBBYTES[0].a/n159 ), .Z(n3224)
         );
  AND U9852 ( .A(\SUBBYTES[0].a/w3376 ), .B(\SUBBYTES[0].a/w3378 ), .Z(
        \SUBBYTES[0].a/w3385 ) );
  AND U9853 ( .A(\SUBBYTES[0].a/w3377 ), .B(\SUBBYTES[0].a/w3379 ), .Z(
        \SUBBYTES[0].a/w3383 ) );
  AND U9854 ( .A(\SUBBYTES[0].a/w3380 ), .B(\SUBBYTES[0].a/w3381 ), .Z(
        \SUBBYTES[0].a/w3382 ) );
  AND U9855 ( .A(\SUBBYTES[0].a/w3269 ), .B(n3219), .Z(\SUBBYTES[0].a/w3368 )
         );
  XOR U9856 ( .A(\SUBBYTES[0].a/w3337 ), .B(n1168), .Z(n3219) );
  AND U9857 ( .A(\SUBBYTES[0].a/w3270 ), .B(n3220), .Z(\SUBBYTES[0].a/w3366 )
         );
  XOR U9858 ( .A(\SUBBYTES[0].a/n160 ), .B(\SUBBYTES[0].a/w3337 ), .Z(n3220)
         );
  ANDN U9859 ( .A(n3221), .B(n3225), .Z(\SUBBYTES[0].a/w3365 ) );
  XOR U9860 ( .A(n1168), .B(\SUBBYTES[0].a/n160 ), .Z(n3221) );
  ANDN U9861 ( .A(\SUBBYTES[0].a/w3271 ), .B(n3222), .Z(\SUBBYTES[0].a/w3361 )
         );
  XNOR U9862 ( .A(\SUBBYTES[0].a/w3330 ), .B(\SUBBYTES[0].a/w3333 ), .Z(n3222)
         );
  AND U9863 ( .A(\SUBBYTES[0].a/w3272 ), .B(n3223), .Z(\SUBBYTES[0].a/w3359 )
         );
  XNOR U9864 ( .A(n3226), .B(\SUBBYTES[0].a/w3330 ), .Z(n3223) );
  AND U9865 ( .A(\SUBBYTES[0].a/w3357 ), .B(n3227), .Z(\SUBBYTES[0].a/w3358 )
         );
  XOR U9866 ( .A(n3228), .B(n3226), .Z(n3227) );
  IV U9867 ( .A(\SUBBYTES[0].a/n159 ), .Z(n3226) );
  ANDN U9868 ( .A(\SUBBYTES[0].a/w3376 ), .B(n3229), .Z(\SUBBYTES[0].a/w3353 )
         );
  ANDN U9869 ( .A(\SUBBYTES[0].a/w3377 ), .B(n3230), .Z(\SUBBYTES[0].a/w3351 )
         );
  ANDN U9870 ( .A(\SUBBYTES[0].a/w3380 ), .B(n3231), .Z(\SUBBYTES[0].a/w3350 )
         );
  AND U9871 ( .A(\SUBBYTES[0].a/w3336 ), .B(\SUBBYTES[0].a/w3335 ), .Z(
        \SUBBYTES[0].a/w3337 ) );
  IV U9872 ( .A(n3228), .Z(\SUBBYTES[0].a/w3333 ) );
  NAND U9873 ( .A(\SUBBYTES[0].a/w3312 ), .B(\SUBBYTES[0].a/w3327 ), .Z(n3228)
         );
  AND U9874 ( .A(\SUBBYTES[0].a/w3329 ), .B(\SUBBYTES[0].a/w3335 ), .Z(
        \SUBBYTES[0].a/w3330 ) );
  AND U9875 ( .A(\SUBBYTES[0].a/w3314 ), .B(\SUBBYTES[0].a/w3312 ), .Z(
        \SUBBYTES[0].a/w3324 ) );
  AND U9876 ( .A(\SUBBYTES[0].a/w3315 ), .B(\SUBBYTES[0].a/w3313 ), .Z(
        \SUBBYTES[0].a/w3322 ) );
  AND U9877 ( .A(\SUBBYTES[0].a/w3329 ), .B(\SUBBYTES[0].a/w3336 ), .Z(
        \SUBBYTES[0].a/w3321 ) );
  AND U9878 ( .A(\SUBBYTES[0].a/w3269 ), .B(\SUBBYTES[0].a/w3265 ), .Z(
        \SUBBYTES[0].a/w3306 ) );
  AND U9879 ( .A(\SUBBYTES[0].a/w3270 ), .B(\SUBBYTES[0].a/w3266 ), .Z(
        \SUBBYTES[0].a/w3304 ) );
  ANDN U9880 ( .A(\SUBBYTES[0].a/w3396 ), .B(n3225), .Z(\SUBBYTES[0].a/w3303 )
         );
  XNOR U9881 ( .A(\w1[0][1] ), .B(\w1[0][7] ), .Z(n3225) );
  XOR U9882 ( .A(g_input[1]), .B(e_input[1]), .Z(\w1[0][1] ) );
  AND U9883 ( .A(\w1[0][0] ), .B(\SUBBYTES[0].a/w3271 ), .Z(
        \SUBBYTES[0].a/w3299 ) );
  XOR U9884 ( .A(g_input[0]), .B(e_input[0]), .Z(\w1[0][0] ) );
  AND U9885 ( .A(\SUBBYTES[0].a/w3272 ), .B(\SUBBYTES[0].a/w3268 ), .Z(
        \SUBBYTES[0].a/w3297 ) );
  AND U9886 ( .A(\SUBBYTES[0].a/w3357 ), .B(\SUBBYTES[0].a/w3389 ), .Z(
        \SUBBYTES[0].a/w3296 ) );
  ANDN U9887 ( .A(\SUBBYTES[0].a/w3378 ), .B(n3229), .Z(\SUBBYTES[0].a/w3291 )
         );
  XNOR U9888 ( .A(\w1[0][4] ), .B(\w1[0][7] ), .Z(n3229) );
  ANDN U9889 ( .A(\SUBBYTES[0].a/w3379 ), .B(n3230), .Z(\SUBBYTES[0].a/w3289 )
         );
  XNOR U9890 ( .A(\w1[0][2] ), .B(\w1[0][7] ), .Z(n3230) );
  XOR U9891 ( .A(g_input[7]), .B(e_input[7]), .Z(\w1[0][7] ) );
  IV U9892 ( .A(n3232), .Z(\w1[0][2] ) );
  ANDN U9893 ( .A(\SUBBYTES[0].a/w3381 ), .B(n3231), .Z(\SUBBYTES[0].a/w3288 )
         );
  XOR U9894 ( .A(n3232), .B(\w1[0][4] ), .Z(n3231) );
  XOR U9895 ( .A(g_input[4]), .B(e_input[4]), .Z(\w1[0][4] ) );
  XNOR U9896 ( .A(g_input[2]), .B(e_input[2]), .Z(n3232) );
  AND U9897 ( .A(n3233), .B(\SUBBYTES[0].a/w3058 ), .Z(\SUBBYTES[0].a/w3193 )
         );
  AND U9898 ( .A(n3234), .B(\SUBBYTES[0].a/w3059 ), .Z(\SUBBYTES[0].a/w3191 )
         );
  AND U9899 ( .A(\SUBBYTES[0].a/w3189 ), .B(n3235), .Z(\SUBBYTES[0].a/w3190 )
         );
  ANDN U9900 ( .A(\w1[0][8] ), .B(n3236), .Z(\SUBBYTES[0].a/w3186 ) );
  AND U9901 ( .A(n3237), .B(\SUBBYTES[0].a/w3061 ), .Z(\SUBBYTES[0].a/w3184 )
         );
  AND U9902 ( .A(\SUBBYTES[0].a/w3182 ), .B(n3238), .Z(\SUBBYTES[0].a/w3183 )
         );
  XOR U9903 ( .A(\SUBBYTES[0].a/w3126 ), .B(\SUBBYTES[0].a/n149 ), .Z(n3238)
         );
  AND U9904 ( .A(\SUBBYTES[0].a/w3169 ), .B(\SUBBYTES[0].a/w3171 ), .Z(
        \SUBBYTES[0].a/w3178 ) );
  AND U9905 ( .A(\SUBBYTES[0].a/w3170 ), .B(\SUBBYTES[0].a/w3172 ), .Z(
        \SUBBYTES[0].a/w3176 ) );
  AND U9906 ( .A(\SUBBYTES[0].a/w3173 ), .B(\SUBBYTES[0].a/w3174 ), .Z(
        \SUBBYTES[0].a/w3175 ) );
  AND U9907 ( .A(\SUBBYTES[0].a/w3062 ), .B(n3233), .Z(\SUBBYTES[0].a/w3161 )
         );
  XOR U9908 ( .A(\SUBBYTES[0].a/w3130 ), .B(n1167), .Z(n3233) );
  AND U9909 ( .A(\SUBBYTES[0].a/w3063 ), .B(n3234), .Z(\SUBBYTES[0].a/w3159 )
         );
  XOR U9910 ( .A(\SUBBYTES[0].a/n150 ), .B(\SUBBYTES[0].a/w3130 ), .Z(n3234)
         );
  ANDN U9911 ( .A(n3235), .B(n3239), .Z(\SUBBYTES[0].a/w3158 ) );
  XOR U9912 ( .A(n1167), .B(\SUBBYTES[0].a/n150 ), .Z(n3235) );
  ANDN U9913 ( .A(\SUBBYTES[0].a/w3064 ), .B(n3236), .Z(\SUBBYTES[0].a/w3154 )
         );
  XNOR U9914 ( .A(\SUBBYTES[0].a/w3123 ), .B(\SUBBYTES[0].a/w3126 ), .Z(n3236)
         );
  AND U9915 ( .A(\SUBBYTES[0].a/w3065 ), .B(n3237), .Z(\SUBBYTES[0].a/w3152 )
         );
  XNOR U9916 ( .A(n3240), .B(\SUBBYTES[0].a/w3123 ), .Z(n3237) );
  AND U9917 ( .A(\SUBBYTES[0].a/w3150 ), .B(n3241), .Z(\SUBBYTES[0].a/w3151 )
         );
  XOR U9918 ( .A(n3242), .B(n3240), .Z(n3241) );
  IV U9919 ( .A(\SUBBYTES[0].a/n149 ), .Z(n3240) );
  ANDN U9920 ( .A(\SUBBYTES[0].a/w3169 ), .B(n3243), .Z(\SUBBYTES[0].a/w3146 )
         );
  ANDN U9921 ( .A(\SUBBYTES[0].a/w3170 ), .B(n3244), .Z(\SUBBYTES[0].a/w3144 )
         );
  ANDN U9922 ( .A(\SUBBYTES[0].a/w3173 ), .B(n3245), .Z(\SUBBYTES[0].a/w3143 )
         );
  AND U9923 ( .A(\SUBBYTES[0].a/w3129 ), .B(\SUBBYTES[0].a/w3128 ), .Z(
        \SUBBYTES[0].a/w3130 ) );
  IV U9924 ( .A(n3242), .Z(\SUBBYTES[0].a/w3126 ) );
  NAND U9925 ( .A(\SUBBYTES[0].a/w3105 ), .B(\SUBBYTES[0].a/w3120 ), .Z(n3242)
         );
  AND U9926 ( .A(\SUBBYTES[0].a/w3122 ), .B(\SUBBYTES[0].a/w3128 ), .Z(
        \SUBBYTES[0].a/w3123 ) );
  AND U9927 ( .A(\SUBBYTES[0].a/w3107 ), .B(\SUBBYTES[0].a/w3105 ), .Z(
        \SUBBYTES[0].a/w3117 ) );
  AND U9928 ( .A(\SUBBYTES[0].a/w3108 ), .B(\SUBBYTES[0].a/w3106 ), .Z(
        \SUBBYTES[0].a/w3115 ) );
  AND U9929 ( .A(\SUBBYTES[0].a/w3122 ), .B(\SUBBYTES[0].a/w3129 ), .Z(
        \SUBBYTES[0].a/w3114 ) );
  AND U9930 ( .A(\SUBBYTES[0].a/w3062 ), .B(\SUBBYTES[0].a/w3058 ), .Z(
        \SUBBYTES[0].a/w3099 ) );
  AND U9931 ( .A(\SUBBYTES[0].a/w3063 ), .B(\SUBBYTES[0].a/w3059 ), .Z(
        \SUBBYTES[0].a/w3097 ) );
  ANDN U9932 ( .A(\SUBBYTES[0].a/w3189 ), .B(n3239), .Z(\SUBBYTES[0].a/w3096 )
         );
  XNOR U9933 ( .A(\w1[0][15] ), .B(\w1[0][9] ), .Z(n3239) );
  XOR U9934 ( .A(g_input[9]), .B(e_input[9]), .Z(\w1[0][9] ) );
  AND U9935 ( .A(\w1[0][8] ), .B(\SUBBYTES[0].a/w3064 ), .Z(
        \SUBBYTES[0].a/w3092 ) );
  XOR U9936 ( .A(g_input[8]), .B(e_input[8]), .Z(\w1[0][8] ) );
  AND U9937 ( .A(\SUBBYTES[0].a/w3065 ), .B(\SUBBYTES[0].a/w3061 ), .Z(
        \SUBBYTES[0].a/w3090 ) );
  AND U9938 ( .A(\SUBBYTES[0].a/w3150 ), .B(\SUBBYTES[0].a/w3182 ), .Z(
        \SUBBYTES[0].a/w3089 ) );
  ANDN U9939 ( .A(\SUBBYTES[0].a/w3171 ), .B(n3243), .Z(\SUBBYTES[0].a/w3084 )
         );
  XNOR U9940 ( .A(\w1[0][12] ), .B(\w1[0][15] ), .Z(n3243) );
  ANDN U9941 ( .A(\SUBBYTES[0].a/w3172 ), .B(n3244), .Z(\SUBBYTES[0].a/w3082 )
         );
  XNOR U9942 ( .A(\w1[0][10] ), .B(\w1[0][15] ), .Z(n3244) );
  XOR U9943 ( .A(g_input[15]), .B(e_input[15]), .Z(\w1[0][15] ) );
  ANDN U9944 ( .A(\SUBBYTES[0].a/w3174 ), .B(n3245), .Z(\SUBBYTES[0].a/w3081 )
         );
  XNOR U9945 ( .A(\w1[0][10] ), .B(\w1[0][12] ), .Z(n3245) );
  XOR U9946 ( .A(g_input[12]), .B(e_input[12]), .Z(\w1[0][12] ) );
  XOR U9947 ( .A(g_input[10]), .B(e_input[10]), .Z(\w1[0][10] ) );
  AND U9948 ( .A(n3246), .B(\SUBBYTES[0].a/w2851 ), .Z(\SUBBYTES[0].a/w2986 )
         );
  AND U9949 ( .A(n3247), .B(\SUBBYTES[0].a/w2852 ), .Z(\SUBBYTES[0].a/w2984 )
         );
  AND U9950 ( .A(\SUBBYTES[0].a/w2982 ), .B(n3248), .Z(\SUBBYTES[0].a/w2983 )
         );
  ANDN U9951 ( .A(\w1[0][16] ), .B(n3249), .Z(\SUBBYTES[0].a/w2979 ) );
  AND U9952 ( .A(n3250), .B(\SUBBYTES[0].a/w2854 ), .Z(\SUBBYTES[0].a/w2977 )
         );
  AND U9953 ( .A(\SUBBYTES[0].a/w2975 ), .B(n3251), .Z(\SUBBYTES[0].a/w2976 )
         );
  XOR U9954 ( .A(\SUBBYTES[0].a/w2919 ), .B(\SUBBYTES[0].a/n139 ), .Z(n3251)
         );
  AND U9955 ( .A(\SUBBYTES[0].a/w2962 ), .B(\SUBBYTES[0].a/w2964 ), .Z(
        \SUBBYTES[0].a/w2971 ) );
  AND U9956 ( .A(\SUBBYTES[0].a/w2963 ), .B(\SUBBYTES[0].a/w2965 ), .Z(
        \SUBBYTES[0].a/w2969 ) );
  AND U9957 ( .A(\SUBBYTES[0].a/w2966 ), .B(\SUBBYTES[0].a/w2967 ), .Z(
        \SUBBYTES[0].a/w2968 ) );
  AND U9958 ( .A(\SUBBYTES[0].a/w2855 ), .B(n3246), .Z(\SUBBYTES[0].a/w2954 )
         );
  XOR U9959 ( .A(\SUBBYTES[0].a/w2923 ), .B(n1166), .Z(n3246) );
  AND U9960 ( .A(\SUBBYTES[0].a/w2856 ), .B(n3247), .Z(\SUBBYTES[0].a/w2952 )
         );
  XOR U9961 ( .A(\SUBBYTES[0].a/n140 ), .B(\SUBBYTES[0].a/w2923 ), .Z(n3247)
         );
  ANDN U9962 ( .A(n3248), .B(n3252), .Z(\SUBBYTES[0].a/w2951 ) );
  XOR U9963 ( .A(n1166), .B(\SUBBYTES[0].a/n140 ), .Z(n3248) );
  AND U9964 ( .A(n3253), .B(\SUBBYTES[0].a/w160 ), .Z(\SUBBYTES[0].a/w295 ) );
  ANDN U9965 ( .A(\SUBBYTES[0].a/w2857 ), .B(n3249), .Z(\SUBBYTES[0].a/w2947 )
         );
  XNOR U9966 ( .A(\SUBBYTES[0].a/w2916 ), .B(\SUBBYTES[0].a/w2919 ), .Z(n3249)
         );
  AND U9967 ( .A(\SUBBYTES[0].a/w2858 ), .B(n3250), .Z(\SUBBYTES[0].a/w2945 )
         );
  XNOR U9968 ( .A(n3254), .B(\SUBBYTES[0].a/w2916 ), .Z(n3250) );
  AND U9969 ( .A(\SUBBYTES[0].a/w2943 ), .B(n3255), .Z(\SUBBYTES[0].a/w2944 )
         );
  XOR U9970 ( .A(n3256), .B(n3254), .Z(n3255) );
  IV U9971 ( .A(\SUBBYTES[0].a/n139 ), .Z(n3254) );
  ANDN U9972 ( .A(\SUBBYTES[0].a/w2962 ), .B(n3257), .Z(\SUBBYTES[0].a/w2939 )
         );
  ANDN U9973 ( .A(\SUBBYTES[0].a/w2963 ), .B(n3258), .Z(\SUBBYTES[0].a/w2937 )
         );
  ANDN U9974 ( .A(\SUBBYTES[0].a/w2966 ), .B(n3259), .Z(\SUBBYTES[0].a/w2936 )
         );
  AND U9975 ( .A(n3260), .B(\SUBBYTES[0].a/w161 ), .Z(\SUBBYTES[0].a/w293 ) );
  AND U9976 ( .A(\SUBBYTES[0].a/w2922 ), .B(\SUBBYTES[0].a/w2921 ), .Z(
        \SUBBYTES[0].a/w2923 ) );
  AND U9977 ( .A(\SUBBYTES[0].a/w291 ), .B(n3261), .Z(\SUBBYTES[0].a/w292 ) );
  IV U9978 ( .A(n3256), .Z(\SUBBYTES[0].a/w2919 ) );
  NAND U9979 ( .A(\SUBBYTES[0].a/w2898 ), .B(\SUBBYTES[0].a/w2913 ), .Z(n3256)
         );
  AND U9980 ( .A(\SUBBYTES[0].a/w2915 ), .B(\SUBBYTES[0].a/w2921 ), .Z(
        \SUBBYTES[0].a/w2916 ) );
  AND U9981 ( .A(\SUBBYTES[0].a/w2900 ), .B(\SUBBYTES[0].a/w2898 ), .Z(
        \SUBBYTES[0].a/w2910 ) );
  AND U9982 ( .A(\SUBBYTES[0].a/w2901 ), .B(\SUBBYTES[0].a/w2899 ), .Z(
        \SUBBYTES[0].a/w2908 ) );
  AND U9983 ( .A(\SUBBYTES[0].a/w2915 ), .B(\SUBBYTES[0].a/w2922 ), .Z(
        \SUBBYTES[0].a/w2907 ) );
  AND U9984 ( .A(\SUBBYTES[0].a/w2855 ), .B(\SUBBYTES[0].a/w2851 ), .Z(
        \SUBBYTES[0].a/w2892 ) );
  AND U9985 ( .A(\SUBBYTES[0].a/w2856 ), .B(\SUBBYTES[0].a/w2852 ), .Z(
        \SUBBYTES[0].a/w2890 ) );
  ANDN U9986 ( .A(\SUBBYTES[0].a/w2982 ), .B(n3252), .Z(\SUBBYTES[0].a/w2889 )
         );
  XNOR U9987 ( .A(\w1[0][17] ), .B(\w1[0][23] ), .Z(n3252) );
  XOR U9988 ( .A(g_input[17]), .B(e_input[17]), .Z(\w1[0][17] ) );
  AND U9989 ( .A(\w1[0][16] ), .B(\SUBBYTES[0].a/w2857 ), .Z(
        \SUBBYTES[0].a/w2885 ) );
  XOR U9990 ( .A(g_input[16]), .B(e_input[16]), .Z(\w1[0][16] ) );
  AND U9991 ( .A(\SUBBYTES[0].a/w2858 ), .B(\SUBBYTES[0].a/w2854 ), .Z(
        \SUBBYTES[0].a/w2883 ) );
  AND U9992 ( .A(\SUBBYTES[0].a/w2943 ), .B(\SUBBYTES[0].a/w2975 ), .Z(
        \SUBBYTES[0].a/w2882 ) );
  ANDN U9993 ( .A(\w1[0][120] ), .B(n3262), .Z(\SUBBYTES[0].a/w288 ) );
  ANDN U9994 ( .A(\SUBBYTES[0].a/w2964 ), .B(n3257), .Z(\SUBBYTES[0].a/w2877 )
         );
  XNOR U9995 ( .A(\w1[0][20] ), .B(\w1[0][23] ), .Z(n3257) );
  ANDN U9996 ( .A(\SUBBYTES[0].a/w2965 ), .B(n3258), .Z(\SUBBYTES[0].a/w2875 )
         );
  XNOR U9997 ( .A(\w1[0][18] ), .B(\w1[0][23] ), .Z(n3258) );
  XOR U9998 ( .A(g_input[23]), .B(e_input[23]), .Z(\w1[0][23] ) );
  IV U9999 ( .A(n3263), .Z(\w1[0][18] ) );
  ANDN U10000 ( .A(\SUBBYTES[0].a/w2967 ), .B(n3259), .Z(\SUBBYTES[0].a/w2874 ) );
  XOR U10001 ( .A(n3263), .B(\w1[0][20] ), .Z(n3259) );
  XOR U10002 ( .A(g_input[20]), .B(e_input[20]), .Z(\w1[0][20] ) );
  XNOR U10003 ( .A(g_input[18]), .B(e_input[18]), .Z(n3263) );
  AND U10004 ( .A(n3264), .B(\SUBBYTES[0].a/w163 ), .Z(\SUBBYTES[0].a/w286 )
         );
  AND U10005 ( .A(\SUBBYTES[0].a/w284 ), .B(n3265), .Z(\SUBBYTES[0].a/w285 )
         );
  XOR U10006 ( .A(\SUBBYTES[0].a/w228 ), .B(\SUBBYTES[0].a/n9 ), .Z(n3265) );
  AND U10007 ( .A(\SUBBYTES[0].a/w271 ), .B(\SUBBYTES[0].a/w273 ), .Z(
        \SUBBYTES[0].a/w280 ) );
  AND U10008 ( .A(\SUBBYTES[0].a/w272 ), .B(\SUBBYTES[0].a/w274 ), .Z(
        \SUBBYTES[0].a/w278 ) );
  AND U10009 ( .A(n3266), .B(\SUBBYTES[0].a/w2644 ), .Z(\SUBBYTES[0].a/w2779 )
         );
  AND U10010 ( .A(n3267), .B(\SUBBYTES[0].a/w2645 ), .Z(\SUBBYTES[0].a/w2777 )
         );
  AND U10011 ( .A(\SUBBYTES[0].a/w2775 ), .B(n3268), .Z(\SUBBYTES[0].a/w2776 )
         );
  ANDN U10012 ( .A(\w1[0][24] ), .B(n3269), .Z(\SUBBYTES[0].a/w2772 ) );
  AND U10013 ( .A(n3270), .B(\SUBBYTES[0].a/w2647 ), .Z(\SUBBYTES[0].a/w2770 )
         );
  AND U10014 ( .A(\SUBBYTES[0].a/w275 ), .B(\SUBBYTES[0].a/w276 ), .Z(
        \SUBBYTES[0].a/w277 ) );
  AND U10015 ( .A(\SUBBYTES[0].a/w2768 ), .B(n3271), .Z(\SUBBYTES[0].a/w2769 )
         );
  XOR U10016 ( .A(\SUBBYTES[0].a/w2712 ), .B(\SUBBYTES[0].a/n129 ), .Z(n3271)
         );
  AND U10017 ( .A(\SUBBYTES[0].a/w2755 ), .B(\SUBBYTES[0].a/w2757 ), .Z(
        \SUBBYTES[0].a/w2764 ) );
  AND U10018 ( .A(\SUBBYTES[0].a/w2756 ), .B(\SUBBYTES[0].a/w2758 ), .Z(
        \SUBBYTES[0].a/w2762 ) );
  AND U10019 ( .A(\SUBBYTES[0].a/w2759 ), .B(\SUBBYTES[0].a/w2760 ), .Z(
        \SUBBYTES[0].a/w2761 ) );
  AND U10020 ( .A(\SUBBYTES[0].a/w2648 ), .B(n3266), .Z(\SUBBYTES[0].a/w2747 )
         );
  XOR U10021 ( .A(\SUBBYTES[0].a/w2716 ), .B(n1165), .Z(n3266) );
  AND U10022 ( .A(\SUBBYTES[0].a/w2649 ), .B(n3267), .Z(\SUBBYTES[0].a/w2745 )
         );
  XOR U10023 ( .A(\SUBBYTES[0].a/n130 ), .B(\SUBBYTES[0].a/w2716 ), .Z(n3267)
         );
  ANDN U10024 ( .A(n3268), .B(n3272), .Z(\SUBBYTES[0].a/w2744 ) );
  XOR U10025 ( .A(n1165), .B(\SUBBYTES[0].a/n130 ), .Z(n3268) );
  ANDN U10026 ( .A(\SUBBYTES[0].a/w2650 ), .B(n3269), .Z(\SUBBYTES[0].a/w2740 ) );
  XNOR U10027 ( .A(\SUBBYTES[0].a/w2709 ), .B(\SUBBYTES[0].a/w2712 ), .Z(n3269) );
  AND U10028 ( .A(\SUBBYTES[0].a/w2651 ), .B(n3270), .Z(\SUBBYTES[0].a/w2738 )
         );
  XNOR U10029 ( .A(n3273), .B(\SUBBYTES[0].a/w2709 ), .Z(n3270) );
  AND U10030 ( .A(\SUBBYTES[0].a/w2736 ), .B(n3274), .Z(\SUBBYTES[0].a/w2737 )
         );
  XOR U10031 ( .A(n3275), .B(n3273), .Z(n3274) );
  IV U10032 ( .A(\SUBBYTES[0].a/n129 ), .Z(n3273) );
  ANDN U10033 ( .A(\SUBBYTES[0].a/w2755 ), .B(n3276), .Z(\SUBBYTES[0].a/w2732 ) );
  ANDN U10034 ( .A(\SUBBYTES[0].a/w2756 ), .B(n3277), .Z(\SUBBYTES[0].a/w2730 ) );
  ANDN U10035 ( .A(\SUBBYTES[0].a/w2759 ), .B(n3278), .Z(\SUBBYTES[0].a/w2729 ) );
  AND U10036 ( .A(\SUBBYTES[0].a/w2715 ), .B(\SUBBYTES[0].a/w2714 ), .Z(
        \SUBBYTES[0].a/w2716 ) );
  IV U10037 ( .A(n3275), .Z(\SUBBYTES[0].a/w2712 ) );
  NAND U10038 ( .A(\SUBBYTES[0].a/w2691 ), .B(\SUBBYTES[0].a/w2706 ), .Z(n3275) );
  AND U10039 ( .A(\SUBBYTES[0].a/w2708 ), .B(\SUBBYTES[0].a/w2714 ), .Z(
        \SUBBYTES[0].a/w2709 ) );
  AND U10040 ( .A(\SUBBYTES[0].a/w2693 ), .B(\SUBBYTES[0].a/w2691 ), .Z(
        \SUBBYTES[0].a/w2703 ) );
  AND U10041 ( .A(\SUBBYTES[0].a/w2694 ), .B(\SUBBYTES[0].a/w2692 ), .Z(
        \SUBBYTES[0].a/w2701 ) );
  AND U10042 ( .A(\SUBBYTES[0].a/w2708 ), .B(\SUBBYTES[0].a/w2715 ), .Z(
        \SUBBYTES[0].a/w2700 ) );
  AND U10043 ( .A(\SUBBYTES[0].a/w2648 ), .B(\SUBBYTES[0].a/w2644 ), .Z(
        \SUBBYTES[0].a/w2685 ) );
  AND U10044 ( .A(\SUBBYTES[0].a/w2649 ), .B(\SUBBYTES[0].a/w2645 ), .Z(
        \SUBBYTES[0].a/w2683 ) );
  ANDN U10045 ( .A(\SUBBYTES[0].a/w2775 ), .B(n3272), .Z(\SUBBYTES[0].a/w2682 ) );
  XNOR U10046 ( .A(\w1[0][25] ), .B(\w1[0][31] ), .Z(n3272) );
  XOR U10047 ( .A(g_input[25]), .B(e_input[25]), .Z(\w1[0][25] ) );
  AND U10048 ( .A(\w1[0][24] ), .B(\SUBBYTES[0].a/w2650 ), .Z(
        \SUBBYTES[0].a/w2678 ) );
  XOR U10049 ( .A(g_input[24]), .B(e_input[24]), .Z(\w1[0][24] ) );
  AND U10050 ( .A(\SUBBYTES[0].a/w2651 ), .B(\SUBBYTES[0].a/w2647 ), .Z(
        \SUBBYTES[0].a/w2676 ) );
  AND U10051 ( .A(\SUBBYTES[0].a/w2736 ), .B(\SUBBYTES[0].a/w2768 ), .Z(
        \SUBBYTES[0].a/w2675 ) );
  ANDN U10052 ( .A(\SUBBYTES[0].a/w2757 ), .B(n3276), .Z(\SUBBYTES[0].a/w2670 ) );
  XNOR U10053 ( .A(\w1[0][28] ), .B(\w1[0][31] ), .Z(n3276) );
  ANDN U10054 ( .A(\SUBBYTES[0].a/w2758 ), .B(n3277), .Z(\SUBBYTES[0].a/w2668 ) );
  XNOR U10055 ( .A(\w1[0][26] ), .B(\w1[0][31] ), .Z(n3277) );
  XOR U10056 ( .A(g_input[31]), .B(e_input[31]), .Z(\w1[0][31] ) );
  IV U10057 ( .A(n3279), .Z(\w1[0][26] ) );
  ANDN U10058 ( .A(\SUBBYTES[0].a/w2760 ), .B(n3278), .Z(\SUBBYTES[0].a/w2667 ) );
  XOR U10059 ( .A(n3279), .B(\w1[0][28] ), .Z(n3278) );
  XOR U10060 ( .A(g_input[28]), .B(e_input[28]), .Z(\w1[0][28] ) );
  XNOR U10061 ( .A(g_input[26]), .B(e_input[26]), .Z(n3279) );
  AND U10062 ( .A(\SUBBYTES[0].a/w164 ), .B(n3253), .Z(\SUBBYTES[0].a/w263 )
         );
  XOR U10063 ( .A(\SUBBYTES[0].a/w232 ), .B(n1153), .Z(n3253) );
  AND U10064 ( .A(\SUBBYTES[0].a/w165 ), .B(n3260), .Z(\SUBBYTES[0].a/w261 )
         );
  XOR U10065 ( .A(\SUBBYTES[0].a/n10 ), .B(\SUBBYTES[0].a/w232 ), .Z(n3260) );
  ANDN U10066 ( .A(n3261), .B(n3280), .Z(\SUBBYTES[0].a/w260 ) );
  XOR U10067 ( .A(n1153), .B(\SUBBYTES[0].a/n10 ), .Z(n3261) );
  AND U10068 ( .A(n3281), .B(\SUBBYTES[0].a/w2437 ), .Z(\SUBBYTES[0].a/w2572 )
         );
  AND U10069 ( .A(n3282), .B(\SUBBYTES[0].a/w2438 ), .Z(\SUBBYTES[0].a/w2570 )
         );
  AND U10070 ( .A(\SUBBYTES[0].a/w2568 ), .B(n3283), .Z(\SUBBYTES[0].a/w2569 )
         );
  ANDN U10071 ( .A(\w1[0][32] ), .B(n3284), .Z(\SUBBYTES[0].a/w2565 ) );
  AND U10072 ( .A(n3285), .B(\SUBBYTES[0].a/w2440 ), .Z(\SUBBYTES[0].a/w2563 )
         );
  AND U10073 ( .A(\SUBBYTES[0].a/w2561 ), .B(n3286), .Z(\SUBBYTES[0].a/w2562 )
         );
  XOR U10074 ( .A(\SUBBYTES[0].a/w2505 ), .B(\SUBBYTES[0].a/n119 ), .Z(n3286)
         );
  ANDN U10075 ( .A(\SUBBYTES[0].a/w166 ), .B(n3262), .Z(\SUBBYTES[0].a/w256 )
         );
  XNOR U10076 ( .A(\SUBBYTES[0].a/w225 ), .B(\SUBBYTES[0].a/w228 ), .Z(n3262)
         );
  AND U10077 ( .A(\SUBBYTES[0].a/w2548 ), .B(\SUBBYTES[0].a/w2550 ), .Z(
        \SUBBYTES[0].a/w2557 ) );
  AND U10078 ( .A(\SUBBYTES[0].a/w2549 ), .B(\SUBBYTES[0].a/w2551 ), .Z(
        \SUBBYTES[0].a/w2555 ) );
  AND U10079 ( .A(\SUBBYTES[0].a/w2552 ), .B(\SUBBYTES[0].a/w2553 ), .Z(
        \SUBBYTES[0].a/w2554 ) );
  AND U10080 ( .A(\SUBBYTES[0].a/w2441 ), .B(n3281), .Z(\SUBBYTES[0].a/w2540 )
         );
  XOR U10081 ( .A(\SUBBYTES[0].a/w2509 ), .B(n1164), .Z(n3281) );
  AND U10082 ( .A(\SUBBYTES[0].a/w167 ), .B(n3264), .Z(\SUBBYTES[0].a/w254 )
         );
  XNOR U10083 ( .A(n3287), .B(\SUBBYTES[0].a/w225 ), .Z(n3264) );
  AND U10084 ( .A(\SUBBYTES[0].a/w2442 ), .B(n3282), .Z(\SUBBYTES[0].a/w2538 )
         );
  XOR U10085 ( .A(\SUBBYTES[0].a/n120 ), .B(\SUBBYTES[0].a/w2509 ), .Z(n3282)
         );
  ANDN U10086 ( .A(n3283), .B(n3288), .Z(\SUBBYTES[0].a/w2537 ) );
  XOR U10087 ( .A(n1164), .B(\SUBBYTES[0].a/n120 ), .Z(n3283) );
  ANDN U10088 ( .A(\SUBBYTES[0].a/w2443 ), .B(n3284), .Z(\SUBBYTES[0].a/w2533 ) );
  XNOR U10089 ( .A(\SUBBYTES[0].a/w2502 ), .B(\SUBBYTES[0].a/w2505 ), .Z(n3284) );
  AND U10090 ( .A(\SUBBYTES[0].a/w2444 ), .B(n3285), .Z(\SUBBYTES[0].a/w2531 )
         );
  XNOR U10091 ( .A(n3289), .B(\SUBBYTES[0].a/w2502 ), .Z(n3285) );
  AND U10092 ( .A(\SUBBYTES[0].a/w2529 ), .B(n3290), .Z(\SUBBYTES[0].a/w2530 )
         );
  XOR U10093 ( .A(n3291), .B(n3289), .Z(n3290) );
  IV U10094 ( .A(\SUBBYTES[0].a/n119 ), .Z(n3289) );
  AND U10095 ( .A(\SUBBYTES[0].a/w252 ), .B(n3292), .Z(\SUBBYTES[0].a/w253 )
         );
  XOR U10096 ( .A(n3293), .B(n3287), .Z(n3292) );
  IV U10097 ( .A(\SUBBYTES[0].a/n9 ), .Z(n3287) );
  ANDN U10098 ( .A(\SUBBYTES[0].a/w2548 ), .B(n3294), .Z(\SUBBYTES[0].a/w2525 ) );
  ANDN U10099 ( .A(\SUBBYTES[0].a/w2549 ), .B(n3295), .Z(\SUBBYTES[0].a/w2523 ) );
  ANDN U10100 ( .A(\SUBBYTES[0].a/w2552 ), .B(n3296), .Z(\SUBBYTES[0].a/w2522 ) );
  AND U10101 ( .A(\SUBBYTES[0].a/w2508 ), .B(\SUBBYTES[0].a/w2507 ), .Z(
        \SUBBYTES[0].a/w2509 ) );
  IV U10102 ( .A(n3291), .Z(\SUBBYTES[0].a/w2505 ) );
  NAND U10103 ( .A(\SUBBYTES[0].a/w2484 ), .B(\SUBBYTES[0].a/w2499 ), .Z(n3291) );
  AND U10104 ( .A(\SUBBYTES[0].a/w2501 ), .B(\SUBBYTES[0].a/w2507 ), .Z(
        \SUBBYTES[0].a/w2502 ) );
  AND U10105 ( .A(\SUBBYTES[0].a/w2486 ), .B(\SUBBYTES[0].a/w2484 ), .Z(
        \SUBBYTES[0].a/w2496 ) );
  AND U10106 ( .A(\SUBBYTES[0].a/w2487 ), .B(\SUBBYTES[0].a/w2485 ), .Z(
        \SUBBYTES[0].a/w2494 ) );
  AND U10107 ( .A(\SUBBYTES[0].a/w2501 ), .B(\SUBBYTES[0].a/w2508 ), .Z(
        \SUBBYTES[0].a/w2493 ) );
  ANDN U10108 ( .A(\SUBBYTES[0].a/w271 ), .B(n3297), .Z(\SUBBYTES[0].a/w248 )
         );
  AND U10109 ( .A(\SUBBYTES[0].a/w2441 ), .B(\SUBBYTES[0].a/w2437 ), .Z(
        \SUBBYTES[0].a/w2478 ) );
  AND U10110 ( .A(\SUBBYTES[0].a/w2442 ), .B(\SUBBYTES[0].a/w2438 ), .Z(
        \SUBBYTES[0].a/w2476 ) );
  ANDN U10111 ( .A(\SUBBYTES[0].a/w2568 ), .B(n3288), .Z(\SUBBYTES[0].a/w2475 ) );
  XNOR U10112 ( .A(\w1[0][33] ), .B(\w1[0][39] ), .Z(n3288) );
  XOR U10113 ( .A(g_input[33]), .B(e_input[33]), .Z(\w1[0][33] ) );
  AND U10114 ( .A(\w1[0][32] ), .B(\SUBBYTES[0].a/w2443 ), .Z(
        \SUBBYTES[0].a/w2471 ) );
  XOR U10115 ( .A(g_input[32]), .B(e_input[32]), .Z(\w1[0][32] ) );
  AND U10116 ( .A(\SUBBYTES[0].a/w2444 ), .B(\SUBBYTES[0].a/w2440 ), .Z(
        \SUBBYTES[0].a/w2469 ) );
  AND U10117 ( .A(\SUBBYTES[0].a/w2529 ), .B(\SUBBYTES[0].a/w2561 ), .Z(
        \SUBBYTES[0].a/w2468 ) );
  ANDN U10118 ( .A(\SUBBYTES[0].a/w2550 ), .B(n3294), .Z(\SUBBYTES[0].a/w2463 ) );
  XNOR U10119 ( .A(\w1[0][36] ), .B(\w1[0][39] ), .Z(n3294) );
  ANDN U10120 ( .A(\SUBBYTES[0].a/w2551 ), .B(n3295), .Z(\SUBBYTES[0].a/w2461 ) );
  XNOR U10121 ( .A(\w1[0][34] ), .B(\w1[0][39] ), .Z(n3295) );
  XOR U10122 ( .A(g_input[39]), .B(e_input[39]), .Z(\w1[0][39] ) );
  IV U10123 ( .A(n3298), .Z(\w1[0][34] ) );
  ANDN U10124 ( .A(\SUBBYTES[0].a/w2553 ), .B(n3296), .Z(\SUBBYTES[0].a/w2460 ) );
  XOR U10125 ( .A(n3298), .B(\w1[0][36] ), .Z(n3296) );
  XOR U10126 ( .A(g_input[36]), .B(e_input[36]), .Z(\w1[0][36] ) );
  XNOR U10127 ( .A(g_input[34]), .B(e_input[34]), .Z(n3298) );
  ANDN U10128 ( .A(\SUBBYTES[0].a/w272 ), .B(n3299), .Z(\SUBBYTES[0].a/w246 )
         );
  ANDN U10129 ( .A(\SUBBYTES[0].a/w275 ), .B(n3300), .Z(\SUBBYTES[0].a/w245 )
         );
  AND U10130 ( .A(n3301), .B(\SUBBYTES[0].a/w2230 ), .Z(\SUBBYTES[0].a/w2365 )
         );
  AND U10131 ( .A(n3302), .B(\SUBBYTES[0].a/w2231 ), .Z(\SUBBYTES[0].a/w2363 )
         );
  AND U10132 ( .A(\SUBBYTES[0].a/w2361 ), .B(n3303), .Z(\SUBBYTES[0].a/w2362 )
         );
  ANDN U10133 ( .A(\w1[0][40] ), .B(n3304), .Z(\SUBBYTES[0].a/w2358 ) );
  AND U10134 ( .A(n3305), .B(\SUBBYTES[0].a/w2233 ), .Z(\SUBBYTES[0].a/w2356 )
         );
  AND U10135 ( .A(\SUBBYTES[0].a/w2354 ), .B(n3306), .Z(\SUBBYTES[0].a/w2355 )
         );
  XOR U10136 ( .A(\SUBBYTES[0].a/w2298 ), .B(\SUBBYTES[0].a/n109 ), .Z(n3306)
         );
  AND U10137 ( .A(\SUBBYTES[0].a/w2341 ), .B(\SUBBYTES[0].a/w2343 ), .Z(
        \SUBBYTES[0].a/w2350 ) );
  AND U10138 ( .A(\SUBBYTES[0].a/w2342 ), .B(\SUBBYTES[0].a/w2344 ), .Z(
        \SUBBYTES[0].a/w2348 ) );
  AND U10139 ( .A(\SUBBYTES[0].a/w2345 ), .B(\SUBBYTES[0].a/w2346 ), .Z(
        \SUBBYTES[0].a/w2347 ) );
  AND U10140 ( .A(\SUBBYTES[0].a/w2234 ), .B(n3301), .Z(\SUBBYTES[0].a/w2333 )
         );
  XOR U10141 ( .A(\SUBBYTES[0].a/w2302 ), .B(n1163), .Z(n3301) );
  AND U10142 ( .A(\SUBBYTES[0].a/w2235 ), .B(n3302), .Z(\SUBBYTES[0].a/w2331 )
         );
  XOR U10143 ( .A(\SUBBYTES[0].a/n110 ), .B(\SUBBYTES[0].a/w2302 ), .Z(n3302)
         );
  ANDN U10144 ( .A(n3303), .B(n3307), .Z(\SUBBYTES[0].a/w2330 ) );
  XOR U10145 ( .A(n1163), .B(\SUBBYTES[0].a/n110 ), .Z(n3303) );
  ANDN U10146 ( .A(\SUBBYTES[0].a/w2236 ), .B(n3304), .Z(\SUBBYTES[0].a/w2326 ) );
  XNOR U10147 ( .A(\SUBBYTES[0].a/w2295 ), .B(\SUBBYTES[0].a/w2298 ), .Z(n3304) );
  AND U10148 ( .A(\SUBBYTES[0].a/w2237 ), .B(n3305), .Z(\SUBBYTES[0].a/w2324 )
         );
  XNOR U10149 ( .A(n3308), .B(\SUBBYTES[0].a/w2295 ), .Z(n3305) );
  AND U10150 ( .A(\SUBBYTES[0].a/w2322 ), .B(n3309), .Z(\SUBBYTES[0].a/w2323 )
         );
  XOR U10151 ( .A(n3310), .B(n3308), .Z(n3309) );
  IV U10152 ( .A(\SUBBYTES[0].a/n109 ), .Z(n3308) );
  AND U10153 ( .A(\SUBBYTES[0].a/w231 ), .B(\SUBBYTES[0].a/w230 ), .Z(
        \SUBBYTES[0].a/w232 ) );
  ANDN U10154 ( .A(\SUBBYTES[0].a/w2341 ), .B(n3311), .Z(\SUBBYTES[0].a/w2318 ) );
  ANDN U10155 ( .A(\SUBBYTES[0].a/w2342 ), .B(n3312), .Z(\SUBBYTES[0].a/w2316 ) );
  ANDN U10156 ( .A(\SUBBYTES[0].a/w2345 ), .B(n3313), .Z(\SUBBYTES[0].a/w2315 ) );
  AND U10157 ( .A(\SUBBYTES[0].a/w2301 ), .B(\SUBBYTES[0].a/w2300 ), .Z(
        \SUBBYTES[0].a/w2302 ) );
  IV U10158 ( .A(n3310), .Z(\SUBBYTES[0].a/w2298 ) );
  NAND U10159 ( .A(\SUBBYTES[0].a/w2277 ), .B(\SUBBYTES[0].a/w2292 ), .Z(n3310) );
  AND U10160 ( .A(\SUBBYTES[0].a/w2294 ), .B(\SUBBYTES[0].a/w2300 ), .Z(
        \SUBBYTES[0].a/w2295 ) );
  AND U10161 ( .A(\SUBBYTES[0].a/w2279 ), .B(\SUBBYTES[0].a/w2277 ), .Z(
        \SUBBYTES[0].a/w2289 ) );
  AND U10162 ( .A(\SUBBYTES[0].a/w2280 ), .B(\SUBBYTES[0].a/w2278 ), .Z(
        \SUBBYTES[0].a/w2287 ) );
  AND U10163 ( .A(\SUBBYTES[0].a/w2294 ), .B(\SUBBYTES[0].a/w2301 ), .Z(
        \SUBBYTES[0].a/w2286 ) );
  IV U10164 ( .A(n3293), .Z(\SUBBYTES[0].a/w228 ) );
  NAND U10165 ( .A(\SUBBYTES[0].a/w207 ), .B(\SUBBYTES[0].a/w222 ), .Z(n3293)
         );
  AND U10166 ( .A(\SUBBYTES[0].a/w2234 ), .B(\SUBBYTES[0].a/w2230 ), .Z(
        \SUBBYTES[0].a/w2271 ) );
  AND U10167 ( .A(\SUBBYTES[0].a/w2235 ), .B(\SUBBYTES[0].a/w2231 ), .Z(
        \SUBBYTES[0].a/w2269 ) );
  ANDN U10168 ( .A(\SUBBYTES[0].a/w2361 ), .B(n3307), .Z(\SUBBYTES[0].a/w2268 ) );
  XNOR U10169 ( .A(\w1[0][41] ), .B(\w1[0][47] ), .Z(n3307) );
  XOR U10170 ( .A(g_input[41]), .B(e_input[41]), .Z(\w1[0][41] ) );
  AND U10171 ( .A(\w1[0][40] ), .B(\SUBBYTES[0].a/w2236 ), .Z(
        \SUBBYTES[0].a/w2264 ) );
  XOR U10172 ( .A(g_input[40]), .B(e_input[40]), .Z(\w1[0][40] ) );
  AND U10173 ( .A(\SUBBYTES[0].a/w2237 ), .B(\SUBBYTES[0].a/w2233 ), .Z(
        \SUBBYTES[0].a/w2262 ) );
  AND U10174 ( .A(\SUBBYTES[0].a/w2322 ), .B(\SUBBYTES[0].a/w2354 ), .Z(
        \SUBBYTES[0].a/w2261 ) );
  ANDN U10175 ( .A(\SUBBYTES[0].a/w2343 ), .B(n3311), .Z(\SUBBYTES[0].a/w2256 ) );
  XNOR U10176 ( .A(\w1[0][44] ), .B(\w1[0][47] ), .Z(n3311) );
  ANDN U10177 ( .A(\SUBBYTES[0].a/w2344 ), .B(n3312), .Z(\SUBBYTES[0].a/w2254 ) );
  XNOR U10178 ( .A(\w1[0][42] ), .B(\w1[0][47] ), .Z(n3312) );
  XOR U10179 ( .A(g_input[47]), .B(e_input[47]), .Z(\w1[0][47] ) );
  IV U10180 ( .A(n3314), .Z(\w1[0][42] ) );
  ANDN U10181 ( .A(\SUBBYTES[0].a/w2346 ), .B(n3313), .Z(\SUBBYTES[0].a/w2253 ) );
  XOR U10182 ( .A(n3314), .B(\w1[0][44] ), .Z(n3313) );
  XOR U10183 ( .A(g_input[44]), .B(e_input[44]), .Z(\w1[0][44] ) );
  XNOR U10184 ( .A(g_input[42]), .B(e_input[42]), .Z(n3314) );
  AND U10185 ( .A(\SUBBYTES[0].a/w224 ), .B(\SUBBYTES[0].a/w230 ), .Z(
        \SUBBYTES[0].a/w225 ) );
  AND U10186 ( .A(\SUBBYTES[0].a/w209 ), .B(\SUBBYTES[0].a/w207 ), .Z(
        \SUBBYTES[0].a/w219 ) );
  AND U10187 ( .A(\SUBBYTES[0].a/w210 ), .B(\SUBBYTES[0].a/w208 ), .Z(
        \SUBBYTES[0].a/w217 ) );
  AND U10188 ( .A(\SUBBYTES[0].a/w224 ), .B(\SUBBYTES[0].a/w231 ), .Z(
        \SUBBYTES[0].a/w216 ) );
  AND U10189 ( .A(n3315), .B(\SUBBYTES[0].a/w2023 ), .Z(\SUBBYTES[0].a/w2158 )
         );
  AND U10190 ( .A(n3316), .B(\SUBBYTES[0].a/w2024 ), .Z(\SUBBYTES[0].a/w2156 )
         );
  AND U10191 ( .A(\SUBBYTES[0].a/w2154 ), .B(n3317), .Z(\SUBBYTES[0].a/w2155 )
         );
  ANDN U10192 ( .A(\w1[0][48] ), .B(n3318), .Z(\SUBBYTES[0].a/w2151 ) );
  AND U10193 ( .A(n3319), .B(\SUBBYTES[0].a/w2026 ), .Z(\SUBBYTES[0].a/w2149 )
         );
  AND U10194 ( .A(\SUBBYTES[0].a/w2147 ), .B(n3320), .Z(\SUBBYTES[0].a/w2148 )
         );
  XOR U10195 ( .A(\SUBBYTES[0].a/w2091 ), .B(\SUBBYTES[0].a/n99 ), .Z(n3320)
         );
  AND U10196 ( .A(\SUBBYTES[0].a/w2134 ), .B(\SUBBYTES[0].a/w2136 ), .Z(
        \SUBBYTES[0].a/w2143 ) );
  AND U10197 ( .A(\SUBBYTES[0].a/w2135 ), .B(\SUBBYTES[0].a/w2137 ), .Z(
        \SUBBYTES[0].a/w2141 ) );
  AND U10198 ( .A(\SUBBYTES[0].a/w2138 ), .B(\SUBBYTES[0].a/w2139 ), .Z(
        \SUBBYTES[0].a/w2140 ) );
  AND U10199 ( .A(\SUBBYTES[0].a/w2027 ), .B(n3315), .Z(\SUBBYTES[0].a/w2126 )
         );
  XOR U10200 ( .A(\SUBBYTES[0].a/w2095 ), .B(n1162), .Z(n3315) );
  AND U10201 ( .A(\SUBBYTES[0].a/w2028 ), .B(n3316), .Z(\SUBBYTES[0].a/w2124 )
         );
  XOR U10202 ( .A(\SUBBYTES[0].a/n100 ), .B(\SUBBYTES[0].a/w2095 ), .Z(n3316)
         );
  ANDN U10203 ( .A(n3317), .B(n3321), .Z(\SUBBYTES[0].a/w2123 ) );
  XOR U10204 ( .A(n1162), .B(\SUBBYTES[0].a/n100 ), .Z(n3317) );
  ANDN U10205 ( .A(\SUBBYTES[0].a/w2029 ), .B(n3318), .Z(\SUBBYTES[0].a/w2119 ) );
  XNOR U10206 ( .A(\SUBBYTES[0].a/w2088 ), .B(\SUBBYTES[0].a/w2091 ), .Z(n3318) );
  AND U10207 ( .A(\SUBBYTES[0].a/w2030 ), .B(n3319), .Z(\SUBBYTES[0].a/w2117 )
         );
  XNOR U10208 ( .A(n3322), .B(\SUBBYTES[0].a/w2088 ), .Z(n3319) );
  AND U10209 ( .A(\SUBBYTES[0].a/w2115 ), .B(n3323), .Z(\SUBBYTES[0].a/w2116 )
         );
  XOR U10210 ( .A(n3324), .B(n3322), .Z(n3323) );
  IV U10211 ( .A(\SUBBYTES[0].a/n99 ), .Z(n3322) );
  ANDN U10212 ( .A(\SUBBYTES[0].a/w2134 ), .B(n3325), .Z(\SUBBYTES[0].a/w2111 ) );
  ANDN U10213 ( .A(\SUBBYTES[0].a/w2135 ), .B(n3326), .Z(\SUBBYTES[0].a/w2109 ) );
  ANDN U10214 ( .A(\SUBBYTES[0].a/w2138 ), .B(n3327), .Z(\SUBBYTES[0].a/w2108 ) );
  AND U10215 ( .A(\SUBBYTES[0].a/w2094 ), .B(\SUBBYTES[0].a/w2093 ), .Z(
        \SUBBYTES[0].a/w2095 ) );
  IV U10216 ( .A(n3324), .Z(\SUBBYTES[0].a/w2091 ) );
  NAND U10217 ( .A(\SUBBYTES[0].a/w2070 ), .B(\SUBBYTES[0].a/w2085 ), .Z(n3324) );
  AND U10218 ( .A(\SUBBYTES[0].a/w2087 ), .B(\SUBBYTES[0].a/w2093 ), .Z(
        \SUBBYTES[0].a/w2088 ) );
  AND U10219 ( .A(\SUBBYTES[0].a/w2072 ), .B(\SUBBYTES[0].a/w2070 ), .Z(
        \SUBBYTES[0].a/w2082 ) );
  AND U10220 ( .A(\SUBBYTES[0].a/w2073 ), .B(\SUBBYTES[0].a/w2071 ), .Z(
        \SUBBYTES[0].a/w2080 ) );
  AND U10221 ( .A(\SUBBYTES[0].a/w2087 ), .B(\SUBBYTES[0].a/w2094 ), .Z(
        \SUBBYTES[0].a/w2079 ) );
  AND U10222 ( .A(\SUBBYTES[0].a/w2027 ), .B(\SUBBYTES[0].a/w2023 ), .Z(
        \SUBBYTES[0].a/w2064 ) );
  AND U10223 ( .A(\SUBBYTES[0].a/w2028 ), .B(\SUBBYTES[0].a/w2024 ), .Z(
        \SUBBYTES[0].a/w2062 ) );
  ANDN U10224 ( .A(\SUBBYTES[0].a/w2154 ), .B(n3321), .Z(\SUBBYTES[0].a/w2061 ) );
  XNOR U10225 ( .A(\w1[0][49] ), .B(\w1[0][55] ), .Z(n3321) );
  XOR U10226 ( .A(g_input[49]), .B(e_input[49]), .Z(\w1[0][49] ) );
  AND U10227 ( .A(\w1[0][48] ), .B(\SUBBYTES[0].a/w2029 ), .Z(
        \SUBBYTES[0].a/w2057 ) );
  XOR U10228 ( .A(g_input[48]), .B(e_input[48]), .Z(\w1[0][48] ) );
  AND U10229 ( .A(\SUBBYTES[0].a/w2030 ), .B(\SUBBYTES[0].a/w2026 ), .Z(
        \SUBBYTES[0].a/w2055 ) );
  AND U10230 ( .A(\SUBBYTES[0].a/w2115 ), .B(\SUBBYTES[0].a/w2147 ), .Z(
        \SUBBYTES[0].a/w2054 ) );
  ANDN U10231 ( .A(\SUBBYTES[0].a/w2136 ), .B(n3325), .Z(\SUBBYTES[0].a/w2049 ) );
  XNOR U10232 ( .A(\w1[0][52] ), .B(\w1[0][55] ), .Z(n3325) );
  ANDN U10233 ( .A(\SUBBYTES[0].a/w2137 ), .B(n3326), .Z(\SUBBYTES[0].a/w2047 ) );
  XNOR U10234 ( .A(\w1[0][50] ), .B(\w1[0][55] ), .Z(n3326) );
  XOR U10235 ( .A(g_input[55]), .B(e_input[55]), .Z(\w1[0][55] ) );
  IV U10236 ( .A(n3328), .Z(\w1[0][50] ) );
  ANDN U10237 ( .A(\SUBBYTES[0].a/w2139 ), .B(n3327), .Z(\SUBBYTES[0].a/w2046 ) );
  XOR U10238 ( .A(n3328), .B(\w1[0][52] ), .Z(n3327) );
  XOR U10239 ( .A(g_input[52]), .B(e_input[52]), .Z(\w1[0][52] ) );
  XNOR U10240 ( .A(g_input[50]), .B(e_input[50]), .Z(n3328) );
  AND U10241 ( .A(\SUBBYTES[0].a/w164 ), .B(\SUBBYTES[0].a/w160 ), .Z(
        \SUBBYTES[0].a/w201 ) );
  AND U10242 ( .A(\SUBBYTES[0].a/w165 ), .B(\SUBBYTES[0].a/w161 ), .Z(
        \SUBBYTES[0].a/w199 ) );
  ANDN U10243 ( .A(\SUBBYTES[0].a/w291 ), .B(n3280), .Z(\SUBBYTES[0].a/w198 )
         );
  XNOR U10244 ( .A(\w1[0][121] ), .B(\w1[0][127] ), .Z(n3280) );
  XOR U10245 ( .A(g_input[121]), .B(e_input[121]), .Z(\w1[0][121] ) );
  AND U10246 ( .A(n3329), .B(\SUBBYTES[0].a/w1816 ), .Z(\SUBBYTES[0].a/w1951 )
         );
  AND U10247 ( .A(n3330), .B(\SUBBYTES[0].a/w1817 ), .Z(\SUBBYTES[0].a/w1949 )
         );
  AND U10248 ( .A(\SUBBYTES[0].a/w1947 ), .B(n3331), .Z(\SUBBYTES[0].a/w1948 )
         );
  ANDN U10249 ( .A(\w1[0][56] ), .B(n3332), .Z(\SUBBYTES[0].a/w1944 ) );
  AND U10250 ( .A(n3333), .B(\SUBBYTES[0].a/w1819 ), .Z(\SUBBYTES[0].a/w1942 )
         );
  AND U10251 ( .A(\SUBBYTES[0].a/w1940 ), .B(n3334), .Z(\SUBBYTES[0].a/w1941 )
         );
  XOR U10252 ( .A(\SUBBYTES[0].a/w1884 ), .B(\SUBBYTES[0].a/n89 ), .Z(n3334)
         );
  AND U10253 ( .A(\w1[0][120] ), .B(\SUBBYTES[0].a/w166 ), .Z(
        \SUBBYTES[0].a/w194 ) );
  XOR U10254 ( .A(g_input[120]), .B(e_input[120]), .Z(\w1[0][120] ) );
  AND U10255 ( .A(\SUBBYTES[0].a/w1927 ), .B(\SUBBYTES[0].a/w1929 ), .Z(
        \SUBBYTES[0].a/w1936 ) );
  AND U10256 ( .A(\SUBBYTES[0].a/w1928 ), .B(\SUBBYTES[0].a/w1930 ), .Z(
        \SUBBYTES[0].a/w1934 ) );
  AND U10257 ( .A(\SUBBYTES[0].a/w1931 ), .B(\SUBBYTES[0].a/w1932 ), .Z(
        \SUBBYTES[0].a/w1933 ) );
  AND U10258 ( .A(\SUBBYTES[0].a/w167 ), .B(\SUBBYTES[0].a/w163 ), .Z(
        \SUBBYTES[0].a/w192 ) );
  AND U10259 ( .A(\SUBBYTES[0].a/w1820 ), .B(n3329), .Z(\SUBBYTES[0].a/w1919 )
         );
  XOR U10260 ( .A(\SUBBYTES[0].a/w1888 ), .B(n1161), .Z(n3329) );
  AND U10261 ( .A(\SUBBYTES[0].a/w1821 ), .B(n3330), .Z(\SUBBYTES[0].a/w1917 )
         );
  XOR U10262 ( .A(\SUBBYTES[0].a/n90 ), .B(\SUBBYTES[0].a/w1888 ), .Z(n3330)
         );
  ANDN U10263 ( .A(n3331), .B(n3335), .Z(\SUBBYTES[0].a/w1916 ) );
  XOR U10264 ( .A(n1161), .B(\SUBBYTES[0].a/n90 ), .Z(n3331) );
  ANDN U10265 ( .A(\SUBBYTES[0].a/w1822 ), .B(n3332), .Z(\SUBBYTES[0].a/w1912 ) );
  XNOR U10266 ( .A(\SUBBYTES[0].a/w1881 ), .B(\SUBBYTES[0].a/w1884 ), .Z(n3332) );
  AND U10267 ( .A(\SUBBYTES[0].a/w1823 ), .B(n3333), .Z(\SUBBYTES[0].a/w1910 )
         );
  XNOR U10268 ( .A(n3336), .B(\SUBBYTES[0].a/w1881 ), .Z(n3333) );
  AND U10269 ( .A(\SUBBYTES[0].a/w252 ), .B(\SUBBYTES[0].a/w284 ), .Z(
        \SUBBYTES[0].a/w191 ) );
  AND U10270 ( .A(\SUBBYTES[0].a/w1908 ), .B(n3337), .Z(\SUBBYTES[0].a/w1909 )
         );
  XOR U10271 ( .A(n3338), .B(n3336), .Z(n3337) );
  IV U10272 ( .A(\SUBBYTES[0].a/n89 ), .Z(n3336) );
  ANDN U10273 ( .A(\SUBBYTES[0].a/w1927 ), .B(n3339), .Z(\SUBBYTES[0].a/w1904 ) );
  ANDN U10274 ( .A(\SUBBYTES[0].a/w1928 ), .B(n3340), .Z(\SUBBYTES[0].a/w1902 ) );
  ANDN U10275 ( .A(\SUBBYTES[0].a/w1931 ), .B(n3341), .Z(\SUBBYTES[0].a/w1901 ) );
  AND U10276 ( .A(\SUBBYTES[0].a/w1887 ), .B(\SUBBYTES[0].a/w1886 ), .Z(
        \SUBBYTES[0].a/w1888 ) );
  IV U10277 ( .A(n3338), .Z(\SUBBYTES[0].a/w1884 ) );
  NAND U10278 ( .A(\SUBBYTES[0].a/w1863 ), .B(\SUBBYTES[0].a/w1878 ), .Z(n3338) );
  AND U10279 ( .A(\SUBBYTES[0].a/w1880 ), .B(\SUBBYTES[0].a/w1886 ), .Z(
        \SUBBYTES[0].a/w1881 ) );
  AND U10280 ( .A(\SUBBYTES[0].a/w1865 ), .B(\SUBBYTES[0].a/w1863 ), .Z(
        \SUBBYTES[0].a/w1875 ) );
  AND U10281 ( .A(\SUBBYTES[0].a/w1866 ), .B(\SUBBYTES[0].a/w1864 ), .Z(
        \SUBBYTES[0].a/w1873 ) );
  AND U10282 ( .A(\SUBBYTES[0].a/w1880 ), .B(\SUBBYTES[0].a/w1887 ), .Z(
        \SUBBYTES[0].a/w1872 ) );
  ANDN U10283 ( .A(\SUBBYTES[0].a/w273 ), .B(n3297), .Z(\SUBBYTES[0].a/w186 )
         );
  XNOR U10284 ( .A(\w1[0][124] ), .B(\w1[0][127] ), .Z(n3297) );
  AND U10285 ( .A(\SUBBYTES[0].a/w1820 ), .B(\SUBBYTES[0].a/w1816 ), .Z(
        \SUBBYTES[0].a/w1857 ) );
  AND U10286 ( .A(\SUBBYTES[0].a/w1821 ), .B(\SUBBYTES[0].a/w1817 ), .Z(
        \SUBBYTES[0].a/w1855 ) );
  ANDN U10287 ( .A(\SUBBYTES[0].a/w1947 ), .B(n3335), .Z(\SUBBYTES[0].a/w1854 ) );
  XNOR U10288 ( .A(\w1[0][57] ), .B(\w1[0][63] ), .Z(n3335) );
  XOR U10289 ( .A(g_input[57]), .B(e_input[57]), .Z(\w1[0][57] ) );
  AND U10290 ( .A(\w1[0][56] ), .B(\SUBBYTES[0].a/w1822 ), .Z(
        \SUBBYTES[0].a/w1850 ) );
  XOR U10291 ( .A(g_input[56]), .B(e_input[56]), .Z(\w1[0][56] ) );
  AND U10292 ( .A(\SUBBYTES[0].a/w1823 ), .B(\SUBBYTES[0].a/w1819 ), .Z(
        \SUBBYTES[0].a/w1848 ) );
  AND U10293 ( .A(\SUBBYTES[0].a/w1908 ), .B(\SUBBYTES[0].a/w1940 ), .Z(
        \SUBBYTES[0].a/w1847 ) );
  ANDN U10294 ( .A(\SUBBYTES[0].a/w1929 ), .B(n3339), .Z(\SUBBYTES[0].a/w1842 ) );
  XNOR U10295 ( .A(\w1[0][60] ), .B(\w1[0][63] ), .Z(n3339) );
  ANDN U10296 ( .A(\SUBBYTES[0].a/w1930 ), .B(n3340), .Z(\SUBBYTES[0].a/w1840 ) );
  XNOR U10297 ( .A(\w1[0][58] ), .B(\w1[0][63] ), .Z(n3340) );
  XOR U10298 ( .A(g_input[63]), .B(e_input[63]), .Z(\w1[0][63] ) );
  IV U10299 ( .A(n3342), .Z(\w1[0][58] ) );
  ANDN U10300 ( .A(\SUBBYTES[0].a/w274 ), .B(n3299), .Z(\SUBBYTES[0].a/w184 )
         );
  XNOR U10301 ( .A(\w1[0][122] ), .B(\w1[0][127] ), .Z(n3299) );
  XOR U10302 ( .A(g_input[127]), .B(e_input[127]), .Z(\w1[0][127] ) );
  IV U10303 ( .A(n3343), .Z(\w1[0][122] ) );
  ANDN U10304 ( .A(\SUBBYTES[0].a/w1932 ), .B(n3341), .Z(\SUBBYTES[0].a/w1839 ) );
  XOR U10305 ( .A(n3342), .B(\w1[0][60] ), .Z(n3341) );
  XOR U10306 ( .A(g_input[60]), .B(e_input[60]), .Z(\w1[0][60] ) );
  XNOR U10307 ( .A(g_input[58]), .B(e_input[58]), .Z(n3342) );
  ANDN U10308 ( .A(\SUBBYTES[0].a/w276 ), .B(n3300), .Z(\SUBBYTES[0].a/w183 )
         );
  XOR U10309 ( .A(n3343), .B(\w1[0][124] ), .Z(n3300) );
  XOR U10310 ( .A(g_input[124]), .B(e_input[124]), .Z(\w1[0][124] ) );
  XNOR U10311 ( .A(g_input[122]), .B(e_input[122]), .Z(n3343) );
  AND U10312 ( .A(n3344), .B(\SUBBYTES[0].a/w1609 ), .Z(\SUBBYTES[0].a/w1744 )
         );
  AND U10313 ( .A(n3345), .B(\SUBBYTES[0].a/w1610 ), .Z(\SUBBYTES[0].a/w1742 )
         );
  AND U10314 ( .A(\SUBBYTES[0].a/w1740 ), .B(n3346), .Z(\SUBBYTES[0].a/w1741 )
         );
  ANDN U10315 ( .A(\w1[0][64] ), .B(n3347), .Z(\SUBBYTES[0].a/w1737 ) );
  AND U10316 ( .A(n3348), .B(\SUBBYTES[0].a/w1612 ), .Z(\SUBBYTES[0].a/w1735 )
         );
  AND U10317 ( .A(\SUBBYTES[0].a/w1733 ), .B(n3349), .Z(\SUBBYTES[0].a/w1734 )
         );
  XOR U10318 ( .A(\SUBBYTES[0].a/w1677 ), .B(\SUBBYTES[0].a/n79 ), .Z(n3349)
         );
  AND U10319 ( .A(\SUBBYTES[0].a/w1720 ), .B(\SUBBYTES[0].a/w1722 ), .Z(
        \SUBBYTES[0].a/w1729 ) );
  AND U10320 ( .A(\SUBBYTES[0].a/w1721 ), .B(\SUBBYTES[0].a/w1723 ), .Z(
        \SUBBYTES[0].a/w1727 ) );
  AND U10321 ( .A(\SUBBYTES[0].a/w1724 ), .B(\SUBBYTES[0].a/w1725 ), .Z(
        \SUBBYTES[0].a/w1726 ) );
  AND U10322 ( .A(\SUBBYTES[0].a/w1613 ), .B(n3344), .Z(\SUBBYTES[0].a/w1712 )
         );
  XOR U10323 ( .A(\SUBBYTES[0].a/w1681 ), .B(n1160), .Z(n3344) );
  AND U10324 ( .A(\SUBBYTES[0].a/w1614 ), .B(n3345), .Z(\SUBBYTES[0].a/w1710 )
         );
  XOR U10325 ( .A(\SUBBYTES[0].a/n80 ), .B(\SUBBYTES[0].a/w1681 ), .Z(n3345)
         );
  ANDN U10326 ( .A(n3346), .B(n3350), .Z(\SUBBYTES[0].a/w1709 ) );
  XOR U10327 ( .A(n1160), .B(\SUBBYTES[0].a/n80 ), .Z(n3346) );
  ANDN U10328 ( .A(\SUBBYTES[0].a/w1615 ), .B(n3347), .Z(\SUBBYTES[0].a/w1705 ) );
  XNOR U10329 ( .A(\SUBBYTES[0].a/w1674 ), .B(\SUBBYTES[0].a/w1677 ), .Z(n3347) );
  AND U10330 ( .A(\SUBBYTES[0].a/w1616 ), .B(n3348), .Z(\SUBBYTES[0].a/w1703 )
         );
  XNOR U10331 ( .A(n3351), .B(\SUBBYTES[0].a/w1674 ), .Z(n3348) );
  AND U10332 ( .A(\SUBBYTES[0].a/w1701 ), .B(n3352), .Z(\SUBBYTES[0].a/w1702 )
         );
  XOR U10333 ( .A(n3353), .B(n3351), .Z(n3352) );
  IV U10334 ( .A(\SUBBYTES[0].a/n79 ), .Z(n3351) );
  ANDN U10335 ( .A(\SUBBYTES[0].a/w1720 ), .B(n3354), .Z(\SUBBYTES[0].a/w1697 ) );
  ANDN U10336 ( .A(\SUBBYTES[0].a/w1721 ), .B(n3355), .Z(\SUBBYTES[0].a/w1695 ) );
  ANDN U10337 ( .A(\SUBBYTES[0].a/w1724 ), .B(n3356), .Z(\SUBBYTES[0].a/w1694 ) );
  AND U10338 ( .A(\SUBBYTES[0].a/w1680 ), .B(\SUBBYTES[0].a/w1679 ), .Z(
        \SUBBYTES[0].a/w1681 ) );
  IV U10339 ( .A(n3353), .Z(\SUBBYTES[0].a/w1677 ) );
  NAND U10340 ( .A(\SUBBYTES[0].a/w1656 ), .B(\SUBBYTES[0].a/w1671 ), .Z(n3353) );
  AND U10341 ( .A(\SUBBYTES[0].a/w1673 ), .B(\SUBBYTES[0].a/w1679 ), .Z(
        \SUBBYTES[0].a/w1674 ) );
  AND U10342 ( .A(\SUBBYTES[0].a/w1658 ), .B(\SUBBYTES[0].a/w1656 ), .Z(
        \SUBBYTES[0].a/w1668 ) );
  AND U10343 ( .A(\SUBBYTES[0].a/w1659 ), .B(\SUBBYTES[0].a/w1657 ), .Z(
        \SUBBYTES[0].a/w1666 ) );
  AND U10344 ( .A(\SUBBYTES[0].a/w1673 ), .B(\SUBBYTES[0].a/w1680 ), .Z(
        \SUBBYTES[0].a/w1665 ) );
  AND U10345 ( .A(\SUBBYTES[0].a/w1613 ), .B(\SUBBYTES[0].a/w1609 ), .Z(
        \SUBBYTES[0].a/w1650 ) );
  AND U10346 ( .A(\SUBBYTES[0].a/w1614 ), .B(\SUBBYTES[0].a/w1610 ), .Z(
        \SUBBYTES[0].a/w1648 ) );
  ANDN U10347 ( .A(\SUBBYTES[0].a/w1740 ), .B(n3350), .Z(\SUBBYTES[0].a/w1647 ) );
  XNOR U10348 ( .A(\w1[0][65] ), .B(\w1[0][71] ), .Z(n3350) );
  XOR U10349 ( .A(g_input[65]), .B(e_input[65]), .Z(\w1[0][65] ) );
  AND U10350 ( .A(\w1[0][64] ), .B(\SUBBYTES[0].a/w1615 ), .Z(
        \SUBBYTES[0].a/w1643 ) );
  XOR U10351 ( .A(g_input[64]), .B(e_input[64]), .Z(\w1[0][64] ) );
  AND U10352 ( .A(\SUBBYTES[0].a/w1616 ), .B(\SUBBYTES[0].a/w1612 ), .Z(
        \SUBBYTES[0].a/w1641 ) );
  AND U10353 ( .A(\SUBBYTES[0].a/w1701 ), .B(\SUBBYTES[0].a/w1733 ), .Z(
        \SUBBYTES[0].a/w1640 ) );
  ANDN U10354 ( .A(\SUBBYTES[0].a/w1722 ), .B(n3354), .Z(\SUBBYTES[0].a/w1635 ) );
  XNOR U10355 ( .A(\w1[0][68] ), .B(\w1[0][71] ), .Z(n3354) );
  ANDN U10356 ( .A(\SUBBYTES[0].a/w1723 ), .B(n3355), .Z(\SUBBYTES[0].a/w1633 ) );
  XNOR U10357 ( .A(\w1[0][66] ), .B(\w1[0][71] ), .Z(n3355) );
  XOR U10358 ( .A(g_input[71]), .B(e_input[71]), .Z(\w1[0][71] ) );
  IV U10359 ( .A(n3357), .Z(\w1[0][66] ) );
  ANDN U10360 ( .A(\SUBBYTES[0].a/w1725 ), .B(n3356), .Z(\SUBBYTES[0].a/w1632 ) );
  XOR U10361 ( .A(n3357), .B(\w1[0][68] ), .Z(n3356) );
  XOR U10362 ( .A(g_input[68]), .B(e_input[68]), .Z(\w1[0][68] ) );
  XNOR U10363 ( .A(g_input[66]), .B(e_input[66]), .Z(n3357) );
  AND U10364 ( .A(n3358), .B(\SUBBYTES[0].a/w1402 ), .Z(\SUBBYTES[0].a/w1537 )
         );
  AND U10365 ( .A(n3359), .B(\SUBBYTES[0].a/w1403 ), .Z(\SUBBYTES[0].a/w1535 )
         );
  AND U10366 ( .A(\SUBBYTES[0].a/w1533 ), .B(n3360), .Z(\SUBBYTES[0].a/w1534 )
         );
  ANDN U10367 ( .A(\w1[0][72] ), .B(n3361), .Z(\SUBBYTES[0].a/w1530 ) );
  AND U10368 ( .A(n3362), .B(\SUBBYTES[0].a/w1405 ), .Z(\SUBBYTES[0].a/w1528 )
         );
  AND U10369 ( .A(\SUBBYTES[0].a/w1526 ), .B(n3363), .Z(\SUBBYTES[0].a/w1527 )
         );
  XOR U10370 ( .A(\SUBBYTES[0].a/w1470 ), .B(\SUBBYTES[0].a/n69 ), .Z(n3363)
         );
  AND U10371 ( .A(\SUBBYTES[0].a/w1513 ), .B(\SUBBYTES[0].a/w1515 ), .Z(
        \SUBBYTES[0].a/w1522 ) );
  AND U10372 ( .A(\SUBBYTES[0].a/w1514 ), .B(\SUBBYTES[0].a/w1516 ), .Z(
        \SUBBYTES[0].a/w1520 ) );
  AND U10373 ( .A(\SUBBYTES[0].a/w1517 ), .B(\SUBBYTES[0].a/w1518 ), .Z(
        \SUBBYTES[0].a/w1519 ) );
  AND U10374 ( .A(\SUBBYTES[0].a/w1406 ), .B(n3358), .Z(\SUBBYTES[0].a/w1505 )
         );
  XOR U10375 ( .A(\SUBBYTES[0].a/w1474 ), .B(n1159), .Z(n3358) );
  AND U10376 ( .A(\SUBBYTES[0].a/w1407 ), .B(n3359), .Z(\SUBBYTES[0].a/w1503 )
         );
  XOR U10377 ( .A(\SUBBYTES[0].a/n70 ), .B(\SUBBYTES[0].a/w1474 ), .Z(n3359)
         );
  ANDN U10378 ( .A(n3360), .B(n3364), .Z(\SUBBYTES[0].a/w1502 ) );
  XOR U10379 ( .A(n1159), .B(\SUBBYTES[0].a/n70 ), .Z(n3360) );
  ANDN U10380 ( .A(\SUBBYTES[0].a/w1408 ), .B(n3361), .Z(\SUBBYTES[0].a/w1498 ) );
  XNOR U10381 ( .A(\SUBBYTES[0].a/w1467 ), .B(\SUBBYTES[0].a/w1470 ), .Z(n3361) );
  AND U10382 ( .A(\SUBBYTES[0].a/w1409 ), .B(n3362), .Z(\SUBBYTES[0].a/w1496 )
         );
  XNOR U10383 ( .A(n3365), .B(\SUBBYTES[0].a/w1467 ), .Z(n3362) );
  AND U10384 ( .A(\SUBBYTES[0].a/w1494 ), .B(n3366), .Z(\SUBBYTES[0].a/w1495 )
         );
  XOR U10385 ( .A(n3367), .B(n3365), .Z(n3366) );
  IV U10386 ( .A(\SUBBYTES[0].a/n69 ), .Z(n3365) );
  ANDN U10387 ( .A(\SUBBYTES[0].a/w1513 ), .B(n3368), .Z(\SUBBYTES[0].a/w1490 ) );
  ANDN U10388 ( .A(\SUBBYTES[0].a/w1514 ), .B(n3369), .Z(\SUBBYTES[0].a/w1488 ) );
  ANDN U10389 ( .A(\SUBBYTES[0].a/w1517 ), .B(n3370), .Z(\SUBBYTES[0].a/w1487 ) );
  AND U10390 ( .A(\SUBBYTES[0].a/w1473 ), .B(\SUBBYTES[0].a/w1472 ), .Z(
        \SUBBYTES[0].a/w1474 ) );
  IV U10391 ( .A(n3367), .Z(\SUBBYTES[0].a/w1470 ) );
  NAND U10392 ( .A(\SUBBYTES[0].a/w1449 ), .B(\SUBBYTES[0].a/w1464 ), .Z(n3367) );
  AND U10393 ( .A(\SUBBYTES[0].a/w1466 ), .B(\SUBBYTES[0].a/w1472 ), .Z(
        \SUBBYTES[0].a/w1467 ) );
  AND U10394 ( .A(\SUBBYTES[0].a/w1451 ), .B(\SUBBYTES[0].a/w1449 ), .Z(
        \SUBBYTES[0].a/w1461 ) );
  AND U10395 ( .A(\SUBBYTES[0].a/w1452 ), .B(\SUBBYTES[0].a/w1450 ), .Z(
        \SUBBYTES[0].a/w1459 ) );
  AND U10396 ( .A(\SUBBYTES[0].a/w1466 ), .B(\SUBBYTES[0].a/w1473 ), .Z(
        \SUBBYTES[0].a/w1458 ) );
  AND U10397 ( .A(\SUBBYTES[0].a/w1406 ), .B(\SUBBYTES[0].a/w1402 ), .Z(
        \SUBBYTES[0].a/w1443 ) );
  AND U10398 ( .A(\SUBBYTES[0].a/w1407 ), .B(\SUBBYTES[0].a/w1403 ), .Z(
        \SUBBYTES[0].a/w1441 ) );
  ANDN U10399 ( .A(\SUBBYTES[0].a/w1533 ), .B(n3364), .Z(\SUBBYTES[0].a/w1440 ) );
  XNOR U10400 ( .A(\w1[0][73] ), .B(\w1[0][79] ), .Z(n3364) );
  XOR U10401 ( .A(g_input[73]), .B(e_input[73]), .Z(\w1[0][73] ) );
  AND U10402 ( .A(\w1[0][72] ), .B(\SUBBYTES[0].a/w1408 ), .Z(
        \SUBBYTES[0].a/w1436 ) );
  XOR U10403 ( .A(g_input[72]), .B(e_input[72]), .Z(\w1[0][72] ) );
  AND U10404 ( .A(\SUBBYTES[0].a/w1409 ), .B(\SUBBYTES[0].a/w1405 ), .Z(
        \SUBBYTES[0].a/w1434 ) );
  AND U10405 ( .A(\SUBBYTES[0].a/w1494 ), .B(\SUBBYTES[0].a/w1526 ), .Z(
        \SUBBYTES[0].a/w1433 ) );
  ANDN U10406 ( .A(\SUBBYTES[0].a/w1515 ), .B(n3368), .Z(\SUBBYTES[0].a/w1428 ) );
  XNOR U10407 ( .A(\w1[0][76] ), .B(\w1[0][79] ), .Z(n3368) );
  ANDN U10408 ( .A(\SUBBYTES[0].a/w1516 ), .B(n3369), .Z(\SUBBYTES[0].a/w1426 ) );
  XNOR U10409 ( .A(\w1[0][74] ), .B(\w1[0][79] ), .Z(n3369) );
  XOR U10410 ( .A(g_input[79]), .B(e_input[79]), .Z(\w1[0][79] ) );
  IV U10411 ( .A(n3371), .Z(\w1[0][74] ) );
  ANDN U10412 ( .A(\SUBBYTES[0].a/w1518 ), .B(n3370), .Z(\SUBBYTES[0].a/w1425 ) );
  XOR U10413 ( .A(n3371), .B(\w1[0][76] ), .Z(n3370) );
  XOR U10414 ( .A(g_input[76]), .B(e_input[76]), .Z(\w1[0][76] ) );
  XNOR U10415 ( .A(g_input[74]), .B(e_input[74]), .Z(n3371) );
  AND U10416 ( .A(n3372), .B(\SUBBYTES[0].a/w1195 ), .Z(\SUBBYTES[0].a/w1330 )
         );
  AND U10417 ( .A(n3373), .B(\SUBBYTES[0].a/w1196 ), .Z(\SUBBYTES[0].a/w1328 )
         );
  AND U10418 ( .A(\SUBBYTES[0].a/w1326 ), .B(n3374), .Z(\SUBBYTES[0].a/w1327 )
         );
  ANDN U10419 ( .A(\w1[0][80] ), .B(n3375), .Z(\SUBBYTES[0].a/w1323 ) );
  AND U10420 ( .A(n3376), .B(\SUBBYTES[0].a/w1198 ), .Z(\SUBBYTES[0].a/w1321 )
         );
  AND U10421 ( .A(\SUBBYTES[0].a/w1319 ), .B(n3377), .Z(\SUBBYTES[0].a/w1320 )
         );
  XOR U10422 ( .A(\SUBBYTES[0].a/w1263 ), .B(\SUBBYTES[0].a/n59 ), .Z(n3377)
         );
  AND U10423 ( .A(\SUBBYTES[0].a/w1306 ), .B(\SUBBYTES[0].a/w1308 ), .Z(
        \SUBBYTES[0].a/w1315 ) );
  AND U10424 ( .A(\SUBBYTES[0].a/w1307 ), .B(\SUBBYTES[0].a/w1309 ), .Z(
        \SUBBYTES[0].a/w1313 ) );
  AND U10425 ( .A(\SUBBYTES[0].a/w1310 ), .B(\SUBBYTES[0].a/w1311 ), .Z(
        \SUBBYTES[0].a/w1312 ) );
  AND U10426 ( .A(\SUBBYTES[0].a/w1199 ), .B(n3372), .Z(\SUBBYTES[0].a/w1298 )
         );
  XOR U10427 ( .A(\SUBBYTES[0].a/w1267 ), .B(n1158), .Z(n3372) );
  AND U10428 ( .A(\SUBBYTES[0].a/w1200 ), .B(n3373), .Z(\SUBBYTES[0].a/w1296 )
         );
  XOR U10429 ( .A(\SUBBYTES[0].a/n60 ), .B(\SUBBYTES[0].a/w1267 ), .Z(n3373)
         );
  ANDN U10430 ( .A(n3374), .B(n3378), .Z(\SUBBYTES[0].a/w1295 ) );
  XOR U10431 ( .A(n1158), .B(\SUBBYTES[0].a/n60 ), .Z(n3374) );
  ANDN U10432 ( .A(\SUBBYTES[0].a/w1201 ), .B(n3375), .Z(\SUBBYTES[0].a/w1291 ) );
  XNOR U10433 ( .A(\SUBBYTES[0].a/w1260 ), .B(\SUBBYTES[0].a/w1263 ), .Z(n3375) );
  AND U10434 ( .A(\SUBBYTES[0].a/w1202 ), .B(n3376), .Z(\SUBBYTES[0].a/w1289 )
         );
  XNOR U10435 ( .A(n3379), .B(\SUBBYTES[0].a/w1260 ), .Z(n3376) );
  AND U10436 ( .A(\SUBBYTES[0].a/w1287 ), .B(n3380), .Z(\SUBBYTES[0].a/w1288 )
         );
  XOR U10437 ( .A(n3381), .B(n3379), .Z(n3380) );
  IV U10438 ( .A(\SUBBYTES[0].a/n59 ), .Z(n3379) );
  ANDN U10439 ( .A(\SUBBYTES[0].a/w1306 ), .B(n3382), .Z(\SUBBYTES[0].a/w1283 ) );
  ANDN U10440 ( .A(\SUBBYTES[0].a/w1307 ), .B(n3383), .Z(\SUBBYTES[0].a/w1281 ) );
  ANDN U10441 ( .A(\SUBBYTES[0].a/w1310 ), .B(n3384), .Z(\SUBBYTES[0].a/w1280 ) );
  AND U10442 ( .A(\SUBBYTES[0].a/w1266 ), .B(\SUBBYTES[0].a/w1265 ), .Z(
        \SUBBYTES[0].a/w1267 ) );
  IV U10443 ( .A(n3381), .Z(\SUBBYTES[0].a/w1263 ) );
  NAND U10444 ( .A(\SUBBYTES[0].a/w1242 ), .B(\SUBBYTES[0].a/w1257 ), .Z(n3381) );
  AND U10445 ( .A(\SUBBYTES[0].a/w1259 ), .B(\SUBBYTES[0].a/w1265 ), .Z(
        \SUBBYTES[0].a/w1260 ) );
  AND U10446 ( .A(\SUBBYTES[0].a/w1244 ), .B(\SUBBYTES[0].a/w1242 ), .Z(
        \SUBBYTES[0].a/w1254 ) );
  AND U10447 ( .A(\SUBBYTES[0].a/w1245 ), .B(\SUBBYTES[0].a/w1243 ), .Z(
        \SUBBYTES[0].a/w1252 ) );
  AND U10448 ( .A(\SUBBYTES[0].a/w1259 ), .B(\SUBBYTES[0].a/w1266 ), .Z(
        \SUBBYTES[0].a/w1251 ) );
  AND U10449 ( .A(\SUBBYTES[0].a/w1199 ), .B(\SUBBYTES[0].a/w1195 ), .Z(
        \SUBBYTES[0].a/w1236 ) );
  AND U10450 ( .A(\SUBBYTES[0].a/w1200 ), .B(\SUBBYTES[0].a/w1196 ), .Z(
        \SUBBYTES[0].a/w1234 ) );
  ANDN U10451 ( .A(\SUBBYTES[0].a/w1326 ), .B(n3378), .Z(\SUBBYTES[0].a/w1233 ) );
  XNOR U10452 ( .A(\w1[0][81] ), .B(\w1[0][87] ), .Z(n3378) );
  XOR U10453 ( .A(g_input[81]), .B(e_input[81]), .Z(\w1[0][81] ) );
  AND U10454 ( .A(\w1[0][80] ), .B(\SUBBYTES[0].a/w1201 ), .Z(
        \SUBBYTES[0].a/w1229 ) );
  XOR U10455 ( .A(g_input[80]), .B(e_input[80]), .Z(\w1[0][80] ) );
  AND U10456 ( .A(\SUBBYTES[0].a/w1202 ), .B(\SUBBYTES[0].a/w1198 ), .Z(
        \SUBBYTES[0].a/w1227 ) );
  AND U10457 ( .A(\SUBBYTES[0].a/w1287 ), .B(\SUBBYTES[0].a/w1319 ), .Z(
        \SUBBYTES[0].a/w1226 ) );
  ANDN U10458 ( .A(\SUBBYTES[0].a/w1308 ), .B(n3382), .Z(\SUBBYTES[0].a/w1221 ) );
  XNOR U10459 ( .A(\w1[0][84] ), .B(\w1[0][87] ), .Z(n3382) );
  ANDN U10460 ( .A(\SUBBYTES[0].a/w1309 ), .B(n3383), .Z(\SUBBYTES[0].a/w1219 ) );
  XNOR U10461 ( .A(\w1[0][82] ), .B(\w1[0][87] ), .Z(n3383) );
  XOR U10462 ( .A(g_input[87]), .B(e_input[87]), .Z(\w1[0][87] ) );
  IV U10463 ( .A(n3385), .Z(\w1[0][82] ) );
  ANDN U10464 ( .A(\SUBBYTES[0].a/w1311 ), .B(n3384), .Z(\SUBBYTES[0].a/w1218 ) );
  XOR U10465 ( .A(n3385), .B(\w1[0][84] ), .Z(n3384) );
  XOR U10466 ( .A(g_input[84]), .B(e_input[84]), .Z(\w1[0][84] ) );
  XNOR U10467 ( .A(g_input[82]), .B(e_input[82]), .Z(n3385) );
  AND U10468 ( .A(n3386), .B(\SUBBYTES[0].a/w988 ), .Z(\SUBBYTES[0].a/w1123 )
         );
  AND U10469 ( .A(n3387), .B(\SUBBYTES[0].a/w989 ), .Z(\SUBBYTES[0].a/w1121 )
         );
  AND U10470 ( .A(\SUBBYTES[0].a/w1119 ), .B(n3388), .Z(\SUBBYTES[0].a/w1120 )
         );
  ANDN U10471 ( .A(\w1[0][88] ), .B(n3389), .Z(\SUBBYTES[0].a/w1116 ) );
  AND U10472 ( .A(n3390), .B(\SUBBYTES[0].a/w991 ), .Z(\SUBBYTES[0].a/w1114 )
         );
  AND U10473 ( .A(\SUBBYTES[0].a/w1112 ), .B(n3391), .Z(\SUBBYTES[0].a/w1113 )
         );
  XOR U10474 ( .A(\SUBBYTES[0].a/w1056 ), .B(\SUBBYTES[0].a/n49 ), .Z(n3391)
         );
  AND U10475 ( .A(\SUBBYTES[0].a/w1099 ), .B(\SUBBYTES[0].a/w1101 ), .Z(
        \SUBBYTES[0].a/w1108 ) );
  AND U10476 ( .A(\SUBBYTES[0].a/w1100 ), .B(\SUBBYTES[0].a/w1102 ), .Z(
        \SUBBYTES[0].a/w1106 ) );
  AND U10477 ( .A(\SUBBYTES[0].a/w1103 ), .B(\SUBBYTES[0].a/w1104 ), .Z(
        \SUBBYTES[0].a/w1105 ) );
  AND U10478 ( .A(\SUBBYTES[0].a/w992 ), .B(n3386), .Z(\SUBBYTES[0].a/w1091 )
         );
  XOR U10479 ( .A(\SUBBYTES[0].a/w1060 ), .B(n1157), .Z(n3386) );
  AND U10480 ( .A(\SUBBYTES[0].a/w993 ), .B(n3387), .Z(\SUBBYTES[0].a/w1089 )
         );
  XOR U10481 ( .A(\SUBBYTES[0].a/n50 ), .B(\SUBBYTES[0].a/w1060 ), .Z(n3387)
         );
  ANDN U10482 ( .A(n3388), .B(n3392), .Z(\SUBBYTES[0].a/w1088 ) );
  XOR U10483 ( .A(n1157), .B(\SUBBYTES[0].a/n50 ), .Z(n3388) );
  ANDN U10484 ( .A(\SUBBYTES[0].a/w994 ), .B(n3389), .Z(\SUBBYTES[0].a/w1084 )
         );
  XNOR U10485 ( .A(\SUBBYTES[0].a/w1053 ), .B(\SUBBYTES[0].a/w1056 ), .Z(n3389) );
  AND U10486 ( .A(\SUBBYTES[0].a/w995 ), .B(n3390), .Z(\SUBBYTES[0].a/w1082 )
         );
  XNOR U10487 ( .A(n3393), .B(\SUBBYTES[0].a/w1053 ), .Z(n3390) );
  AND U10488 ( .A(\SUBBYTES[0].a/w1080 ), .B(n3394), .Z(\SUBBYTES[0].a/w1081 )
         );
  XOR U10489 ( .A(n3395), .B(n3393), .Z(n3394) );
  IV U10490 ( .A(\SUBBYTES[0].a/n49 ), .Z(n3393) );
  ANDN U10491 ( .A(\SUBBYTES[0].a/w1099 ), .B(n3396), .Z(\SUBBYTES[0].a/w1076 ) );
  ANDN U10492 ( .A(\SUBBYTES[0].a/w1100 ), .B(n3397), .Z(\SUBBYTES[0].a/w1074 ) );
  ANDN U10493 ( .A(\SUBBYTES[0].a/w1103 ), .B(n3398), .Z(\SUBBYTES[0].a/w1073 ) );
  AND U10494 ( .A(\SUBBYTES[0].a/w1059 ), .B(\SUBBYTES[0].a/w1058 ), .Z(
        \SUBBYTES[0].a/w1060 ) );
  IV U10495 ( .A(n3395), .Z(\SUBBYTES[0].a/w1056 ) );
  NAND U10496 ( .A(\SUBBYTES[0].a/w1035 ), .B(\SUBBYTES[0].a/w1050 ), .Z(n3395) );
  AND U10497 ( .A(\SUBBYTES[0].a/w1052 ), .B(\SUBBYTES[0].a/w1058 ), .Z(
        \SUBBYTES[0].a/w1053 ) );
  AND U10498 ( .A(\SUBBYTES[0].a/w1037 ), .B(\SUBBYTES[0].a/w1035 ), .Z(
        \SUBBYTES[0].a/w1047 ) );
  AND U10499 ( .A(\SUBBYTES[0].a/w1038 ), .B(\SUBBYTES[0].a/w1036 ), .Z(
        \SUBBYTES[0].a/w1045 ) );
  AND U10500 ( .A(\SUBBYTES[0].a/w1052 ), .B(\SUBBYTES[0].a/w1059 ), .Z(
        \SUBBYTES[0].a/w1044 ) );
  AND U10501 ( .A(\SUBBYTES[0].a/w992 ), .B(\SUBBYTES[0].a/w988 ), .Z(
        \SUBBYTES[0].a/w1029 ) );
  AND U10502 ( .A(\SUBBYTES[0].a/w993 ), .B(\SUBBYTES[0].a/w989 ), .Z(
        \SUBBYTES[0].a/w1027 ) );
  ANDN U10503 ( .A(\SUBBYTES[0].a/w1119 ), .B(n3392), .Z(\SUBBYTES[0].a/w1026 ) );
  XNOR U10504 ( .A(\w1[0][89] ), .B(\w1[0][95] ), .Z(n3392) );
  XOR U10505 ( .A(g_input[89]), .B(e_input[89]), .Z(\w1[0][89] ) );
  AND U10506 ( .A(\w1[0][88] ), .B(\SUBBYTES[0].a/w994 ), .Z(
        \SUBBYTES[0].a/w1022 ) );
  XOR U10507 ( .A(g_input[88]), .B(e_input[88]), .Z(\w1[0][88] ) );
  AND U10508 ( .A(\SUBBYTES[0].a/w995 ), .B(\SUBBYTES[0].a/w991 ), .Z(
        \SUBBYTES[0].a/w1020 ) );
  AND U10509 ( .A(\SUBBYTES[0].a/w1080 ), .B(\SUBBYTES[0].a/w1112 ), .Z(
        \SUBBYTES[0].a/w1019 ) );
  ANDN U10510 ( .A(\SUBBYTES[0].a/w1101 ), .B(n3396), .Z(\SUBBYTES[0].a/w1014 ) );
  XNOR U10511 ( .A(\w1[0][92] ), .B(\w1[0][95] ), .Z(n3396) );
  ANDN U10512 ( .A(\SUBBYTES[0].a/w1102 ), .B(n3397), .Z(\SUBBYTES[0].a/w1012 ) );
  XNOR U10513 ( .A(\w1[0][90] ), .B(\w1[0][95] ), .Z(n3397) );
  XOR U10514 ( .A(g_input[95]), .B(e_input[95]), .Z(\w1[0][95] ) );
  IV U10515 ( .A(n3399), .Z(\w1[0][90] ) );
  ANDN U10516 ( .A(\SUBBYTES[0].a/w1104 ), .B(n3398), .Z(\SUBBYTES[0].a/w1011 ) );
  XOR U10517 ( .A(n3399), .B(\w1[0][92] ), .Z(n3398) );
  XOR U10518 ( .A(g_input[92]), .B(e_input[92]), .Z(\w1[0][92] ) );
  XNOR U10519 ( .A(g_input[90]), .B(e_input[90]), .Z(n3399) );
  AND U10520 ( .A(\SUBBYTES[0].a/w2084 ), .B(\SUBBYTES[0].a/w2071 ), .Z(
        \SUBBYTES[0].a/n99 ) );
  AND U10521 ( .A(\SUBBYTES[0].a/w1877 ), .B(\SUBBYTES[0].a/w1866 ), .Z(
        \SUBBYTES[0].a/n90 ) );
  AND U10522 ( .A(\SUBBYTES[0].a/w221 ), .B(\SUBBYTES[0].a/w208 ), .Z(
        \SUBBYTES[0].a/n9 ) );
  AND U10523 ( .A(\SUBBYTES[0].a/w1877 ), .B(\SUBBYTES[0].a/w1864 ), .Z(
        \SUBBYTES[0].a/n89 ) );
  AND U10524 ( .A(\SUBBYTES[0].a/w1670 ), .B(\SUBBYTES[0].a/w1659 ), .Z(
        \SUBBYTES[0].a/n80 ) );
  AND U10525 ( .A(\SUBBYTES[0].a/w1670 ), .B(\SUBBYTES[0].a/w1657 ), .Z(
        \SUBBYTES[0].a/n79 ) );
  AND U10526 ( .A(\SUBBYTES[0].a/w1463 ), .B(\SUBBYTES[0].a/w1452 ), .Z(
        \SUBBYTES[0].a/n70 ) );
  AND U10527 ( .A(\SUBBYTES[0].a/w1463 ), .B(\SUBBYTES[0].a/w1450 ), .Z(
        \SUBBYTES[0].a/n69 ) );
  AND U10528 ( .A(\SUBBYTES[0].a/w1256 ), .B(\SUBBYTES[0].a/w1245 ), .Z(
        \SUBBYTES[0].a/n60 ) );
  AND U10529 ( .A(\SUBBYTES[0].a/w1256 ), .B(\SUBBYTES[0].a/w1243 ), .Z(
        \SUBBYTES[0].a/n59 ) );
  AND U10530 ( .A(\SUBBYTES[0].a/w1049 ), .B(\SUBBYTES[0].a/w1038 ), .Z(
        \SUBBYTES[0].a/n50 ) );
  AND U10531 ( .A(\SUBBYTES[0].a/w1049 ), .B(\SUBBYTES[0].a/w1036 ), .Z(
        \SUBBYTES[0].a/n49 ) );
  AND U10532 ( .A(\SUBBYTES[0].a/w842 ), .B(\SUBBYTES[0].a/w831 ), .Z(
        \SUBBYTES[0].a/n40 ) );
  AND U10533 ( .A(\SUBBYTES[0].a/w842 ), .B(\SUBBYTES[0].a/w829 ), .Z(
        \SUBBYTES[0].a/n39 ) );
  AND U10534 ( .A(\SUBBYTES[0].a/w635 ), .B(\SUBBYTES[0].a/w624 ), .Z(
        \SUBBYTES[0].a/n30 ) );
  AND U10535 ( .A(\SUBBYTES[0].a/w635 ), .B(\SUBBYTES[0].a/w622 ), .Z(
        \SUBBYTES[0].a/n29 ) );
  AND U10536 ( .A(\SUBBYTES[0].a/w428 ), .B(\SUBBYTES[0].a/w417 ), .Z(
        \SUBBYTES[0].a/n20 ) );
  AND U10537 ( .A(\SUBBYTES[0].a/w428 ), .B(\SUBBYTES[0].a/w415 ), .Z(
        \SUBBYTES[0].a/n19 ) );
  AND U10538 ( .A(\SUBBYTES[0].a/w3326 ), .B(\SUBBYTES[0].a/w3315 ), .Z(
        \SUBBYTES[0].a/n160 ) );
  AND U10539 ( .A(\SUBBYTES[0].a/w3326 ), .B(\SUBBYTES[0].a/w3313 ), .Z(
        \SUBBYTES[0].a/n159 ) );
  AND U10540 ( .A(\SUBBYTES[0].a/w3119 ), .B(\SUBBYTES[0].a/w3108 ), .Z(
        \SUBBYTES[0].a/n150 ) );
  AND U10541 ( .A(\SUBBYTES[0].a/w3119 ), .B(\SUBBYTES[0].a/w3106 ), .Z(
        \SUBBYTES[0].a/n149 ) );
  AND U10542 ( .A(\SUBBYTES[0].a/w2912 ), .B(\SUBBYTES[0].a/w2901 ), .Z(
        \SUBBYTES[0].a/n140 ) );
  AND U10543 ( .A(\SUBBYTES[0].a/w2912 ), .B(\SUBBYTES[0].a/w2899 ), .Z(
        \SUBBYTES[0].a/n139 ) );
  AND U10544 ( .A(\SUBBYTES[0].a/w2705 ), .B(\SUBBYTES[0].a/w2694 ), .Z(
        \SUBBYTES[0].a/n130 ) );
  AND U10545 ( .A(\SUBBYTES[0].a/w2705 ), .B(\SUBBYTES[0].a/w2692 ), .Z(
        \SUBBYTES[0].a/n129 ) );
  AND U10546 ( .A(\SUBBYTES[0].a/w2498 ), .B(\SUBBYTES[0].a/w2487 ), .Z(
        \SUBBYTES[0].a/n120 ) );
  AND U10547 ( .A(\SUBBYTES[0].a/w2498 ), .B(\SUBBYTES[0].a/w2485 ), .Z(
        \SUBBYTES[0].a/n119 ) );
  AND U10548 ( .A(\SUBBYTES[0].a/w2291 ), .B(\SUBBYTES[0].a/w2280 ), .Z(
        \SUBBYTES[0].a/n110 ) );
  AND U10549 ( .A(\SUBBYTES[0].a/w2291 ), .B(\SUBBYTES[0].a/w2278 ), .Z(
        \SUBBYTES[0].a/n109 ) );
  AND U10550 ( .A(\SUBBYTES[0].a/w2084 ), .B(\SUBBYTES[0].a/w2073 ), .Z(
        \SUBBYTES[0].a/n100 ) );
  AND U10551 ( .A(\SUBBYTES[0].a/w221 ), .B(\SUBBYTES[0].a/w210 ), .Z(
        \SUBBYTES[0].a/n10 ) );
endmodule

