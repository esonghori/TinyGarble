
module FA_256 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;


  AND U1 ( .A(A), .B(B), .Z(CO) );
  XOR U2 ( .A(B), .B(A), .Z(S) );
endmodule


module FA_511 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_510 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_509 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_508 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_507 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_506 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_505 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_504 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_503 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_502 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_501 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_500 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_499 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_498 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_497 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_496 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_495 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_494 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_493 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_492 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_491 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_490 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_489 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_488 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_487 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_486 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_485 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_484 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_483 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_482 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_481 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_480 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_479 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_478 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_477 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_476 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_475 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_474 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_473 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_472 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_471 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_470 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_469 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_468 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_467 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_466 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_465 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_464 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_463 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_462 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_461 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_460 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_459 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_458 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_457 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_456 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_455 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_454 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_453 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_452 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_451 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_450 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_449 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_448 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_447 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_446 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_445 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_444 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_443 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_442 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_441 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_440 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_439 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_438 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_437 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_436 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_435 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_434 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_433 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_432 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_431 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_430 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_429 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_428 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_427 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_426 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_425 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_424 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_423 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_422 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_421 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_420 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_419 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_418 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_417 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_416 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_415 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_414 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_413 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_412 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_411 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_410 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_409 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_408 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_407 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_406 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_405 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_404 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_403 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_402 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_401 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_400 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_399 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_398 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_397 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_396 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_395 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_394 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_393 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_392 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_391 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_390 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_389 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_388 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_387 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_386 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_385 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_384 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_383 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_382 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_381 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_380 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_379 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_378 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_377 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_376 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_375 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_374 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_373 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_372 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_371 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_370 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_369 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_368 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_367 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_366 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_365 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_364 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_363 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_362 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_361 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_360 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_359 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_358 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_357 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_356 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_355 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_354 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_353 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_352 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_351 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_350 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_349 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_348 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_347 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_346 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_345 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_344 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_343 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_342 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_341 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_340 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_339 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_338 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_337 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_336 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_335 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_334 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_333 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_332 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_331 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_330 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_329 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_328 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_327 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_326 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_325 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_324 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_323 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_322 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_321 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_320 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_319 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_318 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_317 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_316 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_315 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_314 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_313 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_312 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_311 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_310 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_309 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_308 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_307 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_306 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_305 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_304 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_303 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_302 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_301 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_300 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_299 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_298 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_297 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_296 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_295 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_294 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_293 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_292 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_291 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_290 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_289 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1, n2, n3;

  XNOR U1 ( .A(n1), .B(n2), .Z(S) );
  XOR U2 ( .A(CI), .B(n3), .Z(CO) );
  ANDN U3 ( .B(n2), .A(n1), .Z(n3) );
  XNOR U4 ( .A(A), .B(CI), .Z(n1) );
  XOR U5 ( .A(B), .B(CI), .Z(n2) );
endmodule


module FA_288 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_287 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_286 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_285 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_284 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_283 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_282 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_281 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_280 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_279 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_278 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_277 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_276 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_275 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_274 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_273 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_272 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_271 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_270 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_269 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_268 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_267 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_266 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_265 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_264 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_263 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_262 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_261 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_260 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_259 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  ANDN U2 ( .B(CI), .A(n1), .Z(CO) );
  XOR U3 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_258 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   n1;

  XOR U1 ( .A(CI), .B(n1), .Z(S) );
  XOR U2 ( .A(B), .B(CI), .Z(n1) );
endmodule


module FA_257 ( A, B, CI, S, CO );
  input A, B, CI;
  output S, CO;
  wire   B;
  assign S = B;

endmodule


module ADD_N256_1 ( A, B, CI, S, CO );
  input [255:0] A;
  input [255:0] B;
  output [255:0] S;
  input CI;
  output CO;

  wire   [255:1] C;

  FA_256 \FAINST[0].FA_  ( .A(A[0]), .B(B[0]), .CI(1'b0), .S(S[0]), .CO(C[1])
         );
  FA_511 \FAINST[1].FA_  ( .A(A[1]), .B(B[1]), .CI(C[1]), .S(S[1]), .CO(C[2])
         );
  FA_510 \FAINST[2].FA_  ( .A(A[2]), .B(B[2]), .CI(C[2]), .S(S[2]), .CO(C[3])
         );
  FA_509 \FAINST[3].FA_  ( .A(A[3]), .B(B[3]), .CI(C[3]), .S(S[3]), .CO(C[4])
         );
  FA_508 \FAINST[4].FA_  ( .A(A[4]), .B(B[4]), .CI(C[4]), .S(S[4]), .CO(C[5])
         );
  FA_507 \FAINST[5].FA_  ( .A(A[5]), .B(B[5]), .CI(C[5]), .S(S[5]), .CO(C[6])
         );
  FA_506 \FAINST[6].FA_  ( .A(A[6]), .B(B[6]), .CI(C[6]), .S(S[6]), .CO(C[7])
         );
  FA_505 \FAINST[7].FA_  ( .A(A[7]), .B(B[7]), .CI(C[7]), .S(S[7]), .CO(C[8])
         );
  FA_504 \FAINST[8].FA_  ( .A(A[8]), .B(B[8]), .CI(C[8]), .S(S[8]), .CO(C[9])
         );
  FA_503 \FAINST[9].FA_  ( .A(A[9]), .B(B[9]), .CI(C[9]), .S(S[9]), .CO(C[10])
         );
  FA_502 \FAINST[10].FA_  ( .A(A[10]), .B(B[10]), .CI(C[10]), .S(S[10]), .CO(
        C[11]) );
  FA_501 \FAINST[11].FA_  ( .A(A[11]), .B(B[11]), .CI(C[11]), .S(S[11]), .CO(
        C[12]) );
  FA_500 \FAINST[12].FA_  ( .A(A[12]), .B(B[12]), .CI(C[12]), .S(S[12]), .CO(
        C[13]) );
  FA_499 \FAINST[13].FA_  ( .A(A[13]), .B(B[13]), .CI(C[13]), .S(S[13]), .CO(
        C[14]) );
  FA_498 \FAINST[14].FA_  ( .A(A[14]), .B(B[14]), .CI(C[14]), .S(S[14]), .CO(
        C[15]) );
  FA_497 \FAINST[15].FA_  ( .A(A[15]), .B(B[15]), .CI(C[15]), .S(S[15]), .CO(
        C[16]) );
  FA_496 \FAINST[16].FA_  ( .A(A[16]), .B(B[16]), .CI(C[16]), .S(S[16]), .CO(
        C[17]) );
  FA_495 \FAINST[17].FA_  ( .A(A[17]), .B(B[17]), .CI(C[17]), .S(S[17]), .CO(
        C[18]) );
  FA_494 \FAINST[18].FA_  ( .A(A[18]), .B(B[18]), .CI(C[18]), .S(S[18]), .CO(
        C[19]) );
  FA_493 \FAINST[19].FA_  ( .A(A[19]), .B(B[19]), .CI(C[19]), .S(S[19]), .CO(
        C[20]) );
  FA_492 \FAINST[20].FA_  ( .A(A[20]), .B(B[20]), .CI(C[20]), .S(S[20]), .CO(
        C[21]) );
  FA_491 \FAINST[21].FA_  ( .A(A[21]), .B(B[21]), .CI(C[21]), .S(S[21]), .CO(
        C[22]) );
  FA_490 \FAINST[22].FA_  ( .A(A[22]), .B(B[22]), .CI(C[22]), .S(S[22]), .CO(
        C[23]) );
  FA_489 \FAINST[23].FA_  ( .A(A[23]), .B(B[23]), .CI(C[23]), .S(S[23]), .CO(
        C[24]) );
  FA_488 \FAINST[24].FA_  ( .A(A[24]), .B(B[24]), .CI(C[24]), .S(S[24]), .CO(
        C[25]) );
  FA_487 \FAINST[25].FA_  ( .A(A[25]), .B(B[25]), .CI(C[25]), .S(S[25]), .CO(
        C[26]) );
  FA_486 \FAINST[26].FA_  ( .A(A[26]), .B(B[26]), .CI(C[26]), .S(S[26]), .CO(
        C[27]) );
  FA_485 \FAINST[27].FA_  ( .A(A[27]), .B(B[27]), .CI(C[27]), .S(S[27]), .CO(
        C[28]) );
  FA_484 \FAINST[28].FA_  ( .A(A[28]), .B(B[28]), .CI(C[28]), .S(S[28]), .CO(
        C[29]) );
  FA_483 \FAINST[29].FA_  ( .A(A[29]), .B(B[29]), .CI(C[29]), .S(S[29]), .CO(
        C[30]) );
  FA_482 \FAINST[30].FA_  ( .A(A[30]), .B(B[30]), .CI(C[30]), .S(S[30]), .CO(
        C[31]) );
  FA_481 \FAINST[31].FA_  ( .A(A[31]), .B(B[31]), .CI(C[31]), .S(S[31]), .CO(
        C[32]) );
  FA_480 \FAINST[32].FA_  ( .A(A[32]), .B(B[32]), .CI(C[32]), .S(S[32]), .CO(
        C[33]) );
  FA_479 \FAINST[33].FA_  ( .A(A[33]), .B(B[33]), .CI(C[33]), .S(S[33]), .CO(
        C[34]) );
  FA_478 \FAINST[34].FA_  ( .A(A[34]), .B(B[34]), .CI(C[34]), .S(S[34]), .CO(
        C[35]) );
  FA_477 \FAINST[35].FA_  ( .A(A[35]), .B(B[35]), .CI(C[35]), .S(S[35]), .CO(
        C[36]) );
  FA_476 \FAINST[36].FA_  ( .A(A[36]), .B(B[36]), .CI(C[36]), .S(S[36]), .CO(
        C[37]) );
  FA_475 \FAINST[37].FA_  ( .A(A[37]), .B(B[37]), .CI(C[37]), .S(S[37]), .CO(
        C[38]) );
  FA_474 \FAINST[38].FA_  ( .A(A[38]), .B(B[38]), .CI(C[38]), .S(S[38]), .CO(
        C[39]) );
  FA_473 \FAINST[39].FA_  ( .A(A[39]), .B(B[39]), .CI(C[39]), .S(S[39]), .CO(
        C[40]) );
  FA_472 \FAINST[40].FA_  ( .A(A[40]), .B(B[40]), .CI(C[40]), .S(S[40]), .CO(
        C[41]) );
  FA_471 \FAINST[41].FA_  ( .A(A[41]), .B(B[41]), .CI(C[41]), .S(S[41]), .CO(
        C[42]) );
  FA_470 \FAINST[42].FA_  ( .A(A[42]), .B(B[42]), .CI(C[42]), .S(S[42]), .CO(
        C[43]) );
  FA_469 \FAINST[43].FA_  ( .A(A[43]), .B(B[43]), .CI(C[43]), .S(S[43]), .CO(
        C[44]) );
  FA_468 \FAINST[44].FA_  ( .A(A[44]), .B(B[44]), .CI(C[44]), .S(S[44]), .CO(
        C[45]) );
  FA_467 \FAINST[45].FA_  ( .A(A[45]), .B(B[45]), .CI(C[45]), .S(S[45]), .CO(
        C[46]) );
  FA_466 \FAINST[46].FA_  ( .A(A[46]), .B(B[46]), .CI(C[46]), .S(S[46]), .CO(
        C[47]) );
  FA_465 \FAINST[47].FA_  ( .A(A[47]), .B(B[47]), .CI(C[47]), .S(S[47]), .CO(
        C[48]) );
  FA_464 \FAINST[48].FA_  ( .A(A[48]), .B(B[48]), .CI(C[48]), .S(S[48]), .CO(
        C[49]) );
  FA_463 \FAINST[49].FA_  ( .A(A[49]), .B(B[49]), .CI(C[49]), .S(S[49]), .CO(
        C[50]) );
  FA_462 \FAINST[50].FA_  ( .A(A[50]), .B(B[50]), .CI(C[50]), .S(S[50]), .CO(
        C[51]) );
  FA_461 \FAINST[51].FA_  ( .A(A[51]), .B(B[51]), .CI(C[51]), .S(S[51]), .CO(
        C[52]) );
  FA_460 \FAINST[52].FA_  ( .A(A[52]), .B(B[52]), .CI(C[52]), .S(S[52]), .CO(
        C[53]) );
  FA_459 \FAINST[53].FA_  ( .A(A[53]), .B(B[53]), .CI(C[53]), .S(S[53]), .CO(
        C[54]) );
  FA_458 \FAINST[54].FA_  ( .A(A[54]), .B(B[54]), .CI(C[54]), .S(S[54]), .CO(
        C[55]) );
  FA_457 \FAINST[55].FA_  ( .A(A[55]), .B(B[55]), .CI(C[55]), .S(S[55]), .CO(
        C[56]) );
  FA_456 \FAINST[56].FA_  ( .A(A[56]), .B(B[56]), .CI(C[56]), .S(S[56]), .CO(
        C[57]) );
  FA_455 \FAINST[57].FA_  ( .A(A[57]), .B(B[57]), .CI(C[57]), .S(S[57]), .CO(
        C[58]) );
  FA_454 \FAINST[58].FA_  ( .A(A[58]), .B(B[58]), .CI(C[58]), .S(S[58]), .CO(
        C[59]) );
  FA_453 \FAINST[59].FA_  ( .A(A[59]), .B(B[59]), .CI(C[59]), .S(S[59]), .CO(
        C[60]) );
  FA_452 \FAINST[60].FA_  ( .A(A[60]), .B(B[60]), .CI(C[60]), .S(S[60]), .CO(
        C[61]) );
  FA_451 \FAINST[61].FA_  ( .A(A[61]), .B(B[61]), .CI(C[61]), .S(S[61]), .CO(
        C[62]) );
  FA_450 \FAINST[62].FA_  ( .A(A[62]), .B(B[62]), .CI(C[62]), .S(S[62]), .CO(
        C[63]) );
  FA_449 \FAINST[63].FA_  ( .A(A[63]), .B(B[63]), .CI(C[63]), .S(S[63]), .CO(
        C[64]) );
  FA_448 \FAINST[64].FA_  ( .A(A[64]), .B(B[64]), .CI(C[64]), .S(S[64]), .CO(
        C[65]) );
  FA_447 \FAINST[65].FA_  ( .A(A[65]), .B(B[65]), .CI(C[65]), .S(S[65]), .CO(
        C[66]) );
  FA_446 \FAINST[66].FA_  ( .A(A[66]), .B(B[66]), .CI(C[66]), .S(S[66]), .CO(
        C[67]) );
  FA_445 \FAINST[67].FA_  ( .A(A[67]), .B(B[67]), .CI(C[67]), .S(S[67]), .CO(
        C[68]) );
  FA_444 \FAINST[68].FA_  ( .A(A[68]), .B(B[68]), .CI(C[68]), .S(S[68]), .CO(
        C[69]) );
  FA_443 \FAINST[69].FA_  ( .A(A[69]), .B(B[69]), .CI(C[69]), .S(S[69]), .CO(
        C[70]) );
  FA_442 \FAINST[70].FA_  ( .A(A[70]), .B(B[70]), .CI(C[70]), .S(S[70]), .CO(
        C[71]) );
  FA_441 \FAINST[71].FA_  ( .A(A[71]), .B(B[71]), .CI(C[71]), .S(S[71]), .CO(
        C[72]) );
  FA_440 \FAINST[72].FA_  ( .A(A[72]), .B(B[72]), .CI(C[72]), .S(S[72]), .CO(
        C[73]) );
  FA_439 \FAINST[73].FA_  ( .A(A[73]), .B(B[73]), .CI(C[73]), .S(S[73]), .CO(
        C[74]) );
  FA_438 \FAINST[74].FA_  ( .A(A[74]), .B(B[74]), .CI(C[74]), .S(S[74]), .CO(
        C[75]) );
  FA_437 \FAINST[75].FA_  ( .A(A[75]), .B(B[75]), .CI(C[75]), .S(S[75]), .CO(
        C[76]) );
  FA_436 \FAINST[76].FA_  ( .A(A[76]), .B(B[76]), .CI(C[76]), .S(S[76]), .CO(
        C[77]) );
  FA_435 \FAINST[77].FA_  ( .A(A[77]), .B(B[77]), .CI(C[77]), .S(S[77]), .CO(
        C[78]) );
  FA_434 \FAINST[78].FA_  ( .A(A[78]), .B(B[78]), .CI(C[78]), .S(S[78]), .CO(
        C[79]) );
  FA_433 \FAINST[79].FA_  ( .A(A[79]), .B(B[79]), .CI(C[79]), .S(S[79]), .CO(
        C[80]) );
  FA_432 \FAINST[80].FA_  ( .A(A[80]), .B(B[80]), .CI(C[80]), .S(S[80]), .CO(
        C[81]) );
  FA_431 \FAINST[81].FA_  ( .A(A[81]), .B(B[81]), .CI(C[81]), .S(S[81]), .CO(
        C[82]) );
  FA_430 \FAINST[82].FA_  ( .A(A[82]), .B(B[82]), .CI(C[82]), .S(S[82]), .CO(
        C[83]) );
  FA_429 \FAINST[83].FA_  ( .A(A[83]), .B(B[83]), .CI(C[83]), .S(S[83]), .CO(
        C[84]) );
  FA_428 \FAINST[84].FA_  ( .A(A[84]), .B(B[84]), .CI(C[84]), .S(S[84]), .CO(
        C[85]) );
  FA_427 \FAINST[85].FA_  ( .A(A[85]), .B(B[85]), .CI(C[85]), .S(S[85]), .CO(
        C[86]) );
  FA_426 \FAINST[86].FA_  ( .A(A[86]), .B(B[86]), .CI(C[86]), .S(S[86]), .CO(
        C[87]) );
  FA_425 \FAINST[87].FA_  ( .A(A[87]), .B(B[87]), .CI(C[87]), .S(S[87]), .CO(
        C[88]) );
  FA_424 \FAINST[88].FA_  ( .A(A[88]), .B(B[88]), .CI(C[88]), .S(S[88]), .CO(
        C[89]) );
  FA_423 \FAINST[89].FA_  ( .A(A[89]), .B(B[89]), .CI(C[89]), .S(S[89]), .CO(
        C[90]) );
  FA_422 \FAINST[90].FA_  ( .A(A[90]), .B(B[90]), .CI(C[90]), .S(S[90]), .CO(
        C[91]) );
  FA_421 \FAINST[91].FA_  ( .A(A[91]), .B(B[91]), .CI(C[91]), .S(S[91]), .CO(
        C[92]) );
  FA_420 \FAINST[92].FA_  ( .A(A[92]), .B(B[92]), .CI(C[92]), .S(S[92]), .CO(
        C[93]) );
  FA_419 \FAINST[93].FA_  ( .A(A[93]), .B(B[93]), .CI(C[93]), .S(S[93]), .CO(
        C[94]) );
  FA_418 \FAINST[94].FA_  ( .A(A[94]), .B(B[94]), .CI(C[94]), .S(S[94]), .CO(
        C[95]) );
  FA_417 \FAINST[95].FA_  ( .A(A[95]), .B(B[95]), .CI(C[95]), .S(S[95]), .CO(
        C[96]) );
  FA_416 \FAINST[96].FA_  ( .A(A[96]), .B(B[96]), .CI(C[96]), .S(S[96]), .CO(
        C[97]) );
  FA_415 \FAINST[97].FA_  ( .A(A[97]), .B(B[97]), .CI(C[97]), .S(S[97]), .CO(
        C[98]) );
  FA_414 \FAINST[98].FA_  ( .A(A[98]), .B(B[98]), .CI(C[98]), .S(S[98]), .CO(
        C[99]) );
  FA_413 \FAINST[99].FA_  ( .A(A[99]), .B(B[99]), .CI(C[99]), .S(S[99]), .CO(
        C[100]) );
  FA_412 \FAINST[100].FA_  ( .A(A[100]), .B(B[100]), .CI(C[100]), .S(S[100]), 
        .CO(C[101]) );
  FA_411 \FAINST[101].FA_  ( .A(A[101]), .B(B[101]), .CI(C[101]), .S(S[101]), 
        .CO(C[102]) );
  FA_410 \FAINST[102].FA_  ( .A(A[102]), .B(B[102]), .CI(C[102]), .S(S[102]), 
        .CO(C[103]) );
  FA_409 \FAINST[103].FA_  ( .A(A[103]), .B(B[103]), .CI(C[103]), .S(S[103]), 
        .CO(C[104]) );
  FA_408 \FAINST[104].FA_  ( .A(A[104]), .B(B[104]), .CI(C[104]), .S(S[104]), 
        .CO(C[105]) );
  FA_407 \FAINST[105].FA_  ( .A(A[105]), .B(B[105]), .CI(C[105]), .S(S[105]), 
        .CO(C[106]) );
  FA_406 \FAINST[106].FA_  ( .A(A[106]), .B(B[106]), .CI(C[106]), .S(S[106]), 
        .CO(C[107]) );
  FA_405 \FAINST[107].FA_  ( .A(A[107]), .B(B[107]), .CI(C[107]), .S(S[107]), 
        .CO(C[108]) );
  FA_404 \FAINST[108].FA_  ( .A(A[108]), .B(B[108]), .CI(C[108]), .S(S[108]), 
        .CO(C[109]) );
  FA_403 \FAINST[109].FA_  ( .A(A[109]), .B(B[109]), .CI(C[109]), .S(S[109]), 
        .CO(C[110]) );
  FA_402 \FAINST[110].FA_  ( .A(A[110]), .B(B[110]), .CI(C[110]), .S(S[110]), 
        .CO(C[111]) );
  FA_401 \FAINST[111].FA_  ( .A(A[111]), .B(B[111]), .CI(C[111]), .S(S[111]), 
        .CO(C[112]) );
  FA_400 \FAINST[112].FA_  ( .A(A[112]), .B(B[112]), .CI(C[112]), .S(S[112]), 
        .CO(C[113]) );
  FA_399 \FAINST[113].FA_  ( .A(A[113]), .B(B[113]), .CI(C[113]), .S(S[113]), 
        .CO(C[114]) );
  FA_398 \FAINST[114].FA_  ( .A(A[114]), .B(B[114]), .CI(C[114]), .S(S[114]), 
        .CO(C[115]) );
  FA_397 \FAINST[115].FA_  ( .A(A[115]), .B(B[115]), .CI(C[115]), .S(S[115]), 
        .CO(C[116]) );
  FA_396 \FAINST[116].FA_  ( .A(A[116]), .B(B[116]), .CI(C[116]), .S(S[116]), 
        .CO(C[117]) );
  FA_395 \FAINST[117].FA_  ( .A(A[117]), .B(B[117]), .CI(C[117]), .S(S[117]), 
        .CO(C[118]) );
  FA_394 \FAINST[118].FA_  ( .A(A[118]), .B(B[118]), .CI(C[118]), .S(S[118]), 
        .CO(C[119]) );
  FA_393 \FAINST[119].FA_  ( .A(A[119]), .B(B[119]), .CI(C[119]), .S(S[119]), 
        .CO(C[120]) );
  FA_392 \FAINST[120].FA_  ( .A(A[120]), .B(B[120]), .CI(C[120]), .S(S[120]), 
        .CO(C[121]) );
  FA_391 \FAINST[121].FA_  ( .A(A[121]), .B(B[121]), .CI(C[121]), .S(S[121]), 
        .CO(C[122]) );
  FA_390 \FAINST[122].FA_  ( .A(A[122]), .B(B[122]), .CI(C[122]), .S(S[122]), 
        .CO(C[123]) );
  FA_389 \FAINST[123].FA_  ( .A(A[123]), .B(B[123]), .CI(C[123]), .S(S[123]), 
        .CO(C[124]) );
  FA_388 \FAINST[124].FA_  ( .A(A[124]), .B(B[124]), .CI(C[124]), .S(S[124]), 
        .CO(C[125]) );
  FA_387 \FAINST[125].FA_  ( .A(A[125]), .B(B[125]), .CI(C[125]), .S(S[125]), 
        .CO(C[126]) );
  FA_386 \FAINST[126].FA_  ( .A(A[126]), .B(B[126]), .CI(C[126]), .S(S[126]), 
        .CO(C[127]) );
  FA_385 \FAINST[127].FA_  ( .A(A[127]), .B(B[127]), .CI(C[127]), .S(S[127]), 
        .CO(C[128]) );
  FA_384 \FAINST[128].FA_  ( .A(A[128]), .B(B[128]), .CI(C[128]), .S(S[128]), 
        .CO(C[129]) );
  FA_383 \FAINST[129].FA_  ( .A(A[129]), .B(B[129]), .CI(C[129]), .S(S[129]), 
        .CO(C[130]) );
  FA_382 \FAINST[130].FA_  ( .A(A[130]), .B(B[130]), .CI(C[130]), .S(S[130]), 
        .CO(C[131]) );
  FA_381 \FAINST[131].FA_  ( .A(A[131]), .B(B[131]), .CI(C[131]), .S(S[131]), 
        .CO(C[132]) );
  FA_380 \FAINST[132].FA_  ( .A(A[132]), .B(B[132]), .CI(C[132]), .S(S[132]), 
        .CO(C[133]) );
  FA_379 \FAINST[133].FA_  ( .A(A[133]), .B(B[133]), .CI(C[133]), .S(S[133]), 
        .CO(C[134]) );
  FA_378 \FAINST[134].FA_  ( .A(A[134]), .B(B[134]), .CI(C[134]), .S(S[134]), 
        .CO(C[135]) );
  FA_377 \FAINST[135].FA_  ( .A(A[135]), .B(B[135]), .CI(C[135]), .S(S[135]), 
        .CO(C[136]) );
  FA_376 \FAINST[136].FA_  ( .A(A[136]), .B(B[136]), .CI(C[136]), .S(S[136]), 
        .CO(C[137]) );
  FA_375 \FAINST[137].FA_  ( .A(A[137]), .B(B[137]), .CI(C[137]), .S(S[137]), 
        .CO(C[138]) );
  FA_374 \FAINST[138].FA_  ( .A(A[138]), .B(B[138]), .CI(C[138]), .S(S[138]), 
        .CO(C[139]) );
  FA_373 \FAINST[139].FA_  ( .A(A[139]), .B(B[139]), .CI(C[139]), .S(S[139]), 
        .CO(C[140]) );
  FA_372 \FAINST[140].FA_  ( .A(A[140]), .B(B[140]), .CI(C[140]), .S(S[140]), 
        .CO(C[141]) );
  FA_371 \FAINST[141].FA_  ( .A(A[141]), .B(B[141]), .CI(C[141]), .S(S[141]), 
        .CO(C[142]) );
  FA_370 \FAINST[142].FA_  ( .A(A[142]), .B(B[142]), .CI(C[142]), .S(S[142]), 
        .CO(C[143]) );
  FA_369 \FAINST[143].FA_  ( .A(A[143]), .B(B[143]), .CI(C[143]), .S(S[143]), 
        .CO(C[144]) );
  FA_368 \FAINST[144].FA_  ( .A(A[144]), .B(B[144]), .CI(C[144]), .S(S[144]), 
        .CO(C[145]) );
  FA_367 \FAINST[145].FA_  ( .A(A[145]), .B(B[145]), .CI(C[145]), .S(S[145]), 
        .CO(C[146]) );
  FA_366 \FAINST[146].FA_  ( .A(A[146]), .B(B[146]), .CI(C[146]), .S(S[146]), 
        .CO(C[147]) );
  FA_365 \FAINST[147].FA_  ( .A(A[147]), .B(B[147]), .CI(C[147]), .S(S[147]), 
        .CO(C[148]) );
  FA_364 \FAINST[148].FA_  ( .A(A[148]), .B(B[148]), .CI(C[148]), .S(S[148]), 
        .CO(C[149]) );
  FA_363 \FAINST[149].FA_  ( .A(A[149]), .B(B[149]), .CI(C[149]), .S(S[149]), 
        .CO(C[150]) );
  FA_362 \FAINST[150].FA_  ( .A(A[150]), .B(B[150]), .CI(C[150]), .S(S[150]), 
        .CO(C[151]) );
  FA_361 \FAINST[151].FA_  ( .A(A[151]), .B(B[151]), .CI(C[151]), .S(S[151]), 
        .CO(C[152]) );
  FA_360 \FAINST[152].FA_  ( .A(A[152]), .B(B[152]), .CI(C[152]), .S(S[152]), 
        .CO(C[153]) );
  FA_359 \FAINST[153].FA_  ( .A(A[153]), .B(B[153]), .CI(C[153]), .S(S[153]), 
        .CO(C[154]) );
  FA_358 \FAINST[154].FA_  ( .A(A[154]), .B(B[154]), .CI(C[154]), .S(S[154]), 
        .CO(C[155]) );
  FA_357 \FAINST[155].FA_  ( .A(A[155]), .B(B[155]), .CI(C[155]), .S(S[155]), 
        .CO(C[156]) );
  FA_356 \FAINST[156].FA_  ( .A(A[156]), .B(B[156]), .CI(C[156]), .S(S[156]), 
        .CO(C[157]) );
  FA_355 \FAINST[157].FA_  ( .A(A[157]), .B(B[157]), .CI(C[157]), .S(S[157]), 
        .CO(C[158]) );
  FA_354 \FAINST[158].FA_  ( .A(A[158]), .B(B[158]), .CI(C[158]), .S(S[158]), 
        .CO(C[159]) );
  FA_353 \FAINST[159].FA_  ( .A(A[159]), .B(B[159]), .CI(C[159]), .S(S[159]), 
        .CO(C[160]) );
  FA_352 \FAINST[160].FA_  ( .A(A[160]), .B(B[160]), .CI(C[160]), .S(S[160]), 
        .CO(C[161]) );
  FA_351 \FAINST[161].FA_  ( .A(A[161]), .B(B[161]), .CI(C[161]), .S(S[161]), 
        .CO(C[162]) );
  FA_350 \FAINST[162].FA_  ( .A(A[162]), .B(B[162]), .CI(C[162]), .S(S[162]), 
        .CO(C[163]) );
  FA_349 \FAINST[163].FA_  ( .A(A[163]), .B(B[163]), .CI(C[163]), .S(S[163]), 
        .CO(C[164]) );
  FA_348 \FAINST[164].FA_  ( .A(A[164]), .B(B[164]), .CI(C[164]), .S(S[164]), 
        .CO(C[165]) );
  FA_347 \FAINST[165].FA_  ( .A(A[165]), .B(B[165]), .CI(C[165]), .S(S[165]), 
        .CO(C[166]) );
  FA_346 \FAINST[166].FA_  ( .A(A[166]), .B(B[166]), .CI(C[166]), .S(S[166]), 
        .CO(C[167]) );
  FA_345 \FAINST[167].FA_  ( .A(A[167]), .B(B[167]), .CI(C[167]), .S(S[167]), 
        .CO(C[168]) );
  FA_344 \FAINST[168].FA_  ( .A(A[168]), .B(B[168]), .CI(C[168]), .S(S[168]), 
        .CO(C[169]) );
  FA_343 \FAINST[169].FA_  ( .A(A[169]), .B(B[169]), .CI(C[169]), .S(S[169]), 
        .CO(C[170]) );
  FA_342 \FAINST[170].FA_  ( .A(A[170]), .B(B[170]), .CI(C[170]), .S(S[170]), 
        .CO(C[171]) );
  FA_341 \FAINST[171].FA_  ( .A(A[171]), .B(B[171]), .CI(C[171]), .S(S[171]), 
        .CO(C[172]) );
  FA_340 \FAINST[172].FA_  ( .A(A[172]), .B(B[172]), .CI(C[172]), .S(S[172]), 
        .CO(C[173]) );
  FA_339 \FAINST[173].FA_  ( .A(A[173]), .B(B[173]), .CI(C[173]), .S(S[173]), 
        .CO(C[174]) );
  FA_338 \FAINST[174].FA_  ( .A(A[174]), .B(B[174]), .CI(C[174]), .S(S[174]), 
        .CO(C[175]) );
  FA_337 \FAINST[175].FA_  ( .A(A[175]), .B(B[175]), .CI(C[175]), .S(S[175]), 
        .CO(C[176]) );
  FA_336 \FAINST[176].FA_  ( .A(A[176]), .B(B[176]), .CI(C[176]), .S(S[176]), 
        .CO(C[177]) );
  FA_335 \FAINST[177].FA_  ( .A(A[177]), .B(B[177]), .CI(C[177]), .S(S[177]), 
        .CO(C[178]) );
  FA_334 \FAINST[178].FA_  ( .A(A[178]), .B(B[178]), .CI(C[178]), .S(S[178]), 
        .CO(C[179]) );
  FA_333 \FAINST[179].FA_  ( .A(A[179]), .B(B[179]), .CI(C[179]), .S(S[179]), 
        .CO(C[180]) );
  FA_332 \FAINST[180].FA_  ( .A(A[180]), .B(B[180]), .CI(C[180]), .S(S[180]), 
        .CO(C[181]) );
  FA_331 \FAINST[181].FA_  ( .A(A[181]), .B(B[181]), .CI(C[181]), .S(S[181]), 
        .CO(C[182]) );
  FA_330 \FAINST[182].FA_  ( .A(A[182]), .B(B[182]), .CI(C[182]), .S(S[182]), 
        .CO(C[183]) );
  FA_329 \FAINST[183].FA_  ( .A(A[183]), .B(B[183]), .CI(C[183]), .S(S[183]), 
        .CO(C[184]) );
  FA_328 \FAINST[184].FA_  ( .A(A[184]), .B(B[184]), .CI(C[184]), .S(S[184]), 
        .CO(C[185]) );
  FA_327 \FAINST[185].FA_  ( .A(A[185]), .B(B[185]), .CI(C[185]), .S(S[185]), 
        .CO(C[186]) );
  FA_326 \FAINST[186].FA_  ( .A(A[186]), .B(B[186]), .CI(C[186]), .S(S[186]), 
        .CO(C[187]) );
  FA_325 \FAINST[187].FA_  ( .A(A[187]), .B(B[187]), .CI(C[187]), .S(S[187]), 
        .CO(C[188]) );
  FA_324 \FAINST[188].FA_  ( .A(A[188]), .B(B[188]), .CI(C[188]), .S(S[188]), 
        .CO(C[189]) );
  FA_323 \FAINST[189].FA_  ( .A(A[189]), .B(B[189]), .CI(C[189]), .S(S[189]), 
        .CO(C[190]) );
  FA_322 \FAINST[190].FA_  ( .A(A[190]), .B(B[190]), .CI(C[190]), .S(S[190]), 
        .CO(C[191]) );
  FA_321 \FAINST[191].FA_  ( .A(A[191]), .B(B[191]), .CI(C[191]), .S(S[191]), 
        .CO(C[192]) );
  FA_320 \FAINST[192].FA_  ( .A(A[192]), .B(B[192]), .CI(C[192]), .S(S[192]), 
        .CO(C[193]) );
  FA_319 \FAINST[193].FA_  ( .A(A[193]), .B(B[193]), .CI(C[193]), .S(S[193]), 
        .CO(C[194]) );
  FA_318 \FAINST[194].FA_  ( .A(A[194]), .B(B[194]), .CI(C[194]), .S(S[194]), 
        .CO(C[195]) );
  FA_317 \FAINST[195].FA_  ( .A(A[195]), .B(B[195]), .CI(C[195]), .S(S[195]), 
        .CO(C[196]) );
  FA_316 \FAINST[196].FA_  ( .A(A[196]), .B(B[196]), .CI(C[196]), .S(S[196]), 
        .CO(C[197]) );
  FA_315 \FAINST[197].FA_  ( .A(A[197]), .B(B[197]), .CI(C[197]), .S(S[197]), 
        .CO(C[198]) );
  FA_314 \FAINST[198].FA_  ( .A(A[198]), .B(B[198]), .CI(C[198]), .S(S[198]), 
        .CO(C[199]) );
  FA_313 \FAINST[199].FA_  ( .A(A[199]), .B(B[199]), .CI(C[199]), .S(S[199]), 
        .CO(C[200]) );
  FA_312 \FAINST[200].FA_  ( .A(A[200]), .B(B[200]), .CI(C[200]), .S(S[200]), 
        .CO(C[201]) );
  FA_311 \FAINST[201].FA_  ( .A(A[201]), .B(B[201]), .CI(C[201]), .S(S[201]), 
        .CO(C[202]) );
  FA_310 \FAINST[202].FA_  ( .A(A[202]), .B(B[202]), .CI(C[202]), .S(S[202]), 
        .CO(C[203]) );
  FA_309 \FAINST[203].FA_  ( .A(A[203]), .B(B[203]), .CI(C[203]), .S(S[203]), 
        .CO(C[204]) );
  FA_308 \FAINST[204].FA_  ( .A(A[204]), .B(B[204]), .CI(C[204]), .S(S[204]), 
        .CO(C[205]) );
  FA_307 \FAINST[205].FA_  ( .A(A[205]), .B(B[205]), .CI(C[205]), .S(S[205]), 
        .CO(C[206]) );
  FA_306 \FAINST[206].FA_  ( .A(A[206]), .B(B[206]), .CI(C[206]), .S(S[206]), 
        .CO(C[207]) );
  FA_305 \FAINST[207].FA_  ( .A(A[207]), .B(B[207]), .CI(C[207]), .S(S[207]), 
        .CO(C[208]) );
  FA_304 \FAINST[208].FA_  ( .A(A[208]), .B(B[208]), .CI(C[208]), .S(S[208]), 
        .CO(C[209]) );
  FA_303 \FAINST[209].FA_  ( .A(A[209]), .B(B[209]), .CI(C[209]), .S(S[209]), 
        .CO(C[210]) );
  FA_302 \FAINST[210].FA_  ( .A(A[210]), .B(B[210]), .CI(C[210]), .S(S[210]), 
        .CO(C[211]) );
  FA_301 \FAINST[211].FA_  ( .A(A[211]), .B(B[211]), .CI(C[211]), .S(S[211]), 
        .CO(C[212]) );
  FA_300 \FAINST[212].FA_  ( .A(A[212]), .B(B[212]), .CI(C[212]), .S(S[212]), 
        .CO(C[213]) );
  FA_299 \FAINST[213].FA_  ( .A(A[213]), .B(B[213]), .CI(C[213]), .S(S[213]), 
        .CO(C[214]) );
  FA_298 \FAINST[214].FA_  ( .A(A[214]), .B(B[214]), .CI(C[214]), .S(S[214]), 
        .CO(C[215]) );
  FA_297 \FAINST[215].FA_  ( .A(A[215]), .B(B[215]), .CI(C[215]), .S(S[215]), 
        .CO(C[216]) );
  FA_296 \FAINST[216].FA_  ( .A(A[216]), .B(B[216]), .CI(C[216]), .S(S[216]), 
        .CO(C[217]) );
  FA_295 \FAINST[217].FA_  ( .A(A[217]), .B(B[217]), .CI(C[217]), .S(S[217]), 
        .CO(C[218]) );
  FA_294 \FAINST[218].FA_  ( .A(A[218]), .B(B[218]), .CI(C[218]), .S(S[218]), 
        .CO(C[219]) );
  FA_293 \FAINST[219].FA_  ( .A(A[219]), .B(B[219]), .CI(C[219]), .S(S[219]), 
        .CO(C[220]) );
  FA_292 \FAINST[220].FA_  ( .A(A[220]), .B(B[220]), .CI(C[220]), .S(S[220]), 
        .CO(C[221]) );
  FA_291 \FAINST[221].FA_  ( .A(A[221]), .B(B[221]), .CI(C[221]), .S(S[221]), 
        .CO(C[222]) );
  FA_290 \FAINST[222].FA_  ( .A(A[222]), .B(B[222]), .CI(C[222]), .S(S[222]), 
        .CO(C[223]) );
  FA_289 \FAINST[223].FA_  ( .A(A[223]), .B(B[223]), .CI(C[223]), .S(S[223]), 
        .CO(C[224]) );
  FA_288 \FAINST[224].FA_  ( .A(1'b0), .B(B[224]), .CI(C[224]), .S(S[224]), 
        .CO(C[225]) );
  FA_287 \FAINST[225].FA_  ( .A(1'b0), .B(B[225]), .CI(C[225]), .S(S[225]), 
        .CO(C[226]) );
  FA_286 \FAINST[226].FA_  ( .A(1'b0), .B(B[226]), .CI(C[226]), .S(S[226]), 
        .CO(C[227]) );
  FA_285 \FAINST[227].FA_  ( .A(1'b0), .B(B[227]), .CI(C[227]), .S(S[227]), 
        .CO(C[228]) );
  FA_284 \FAINST[228].FA_  ( .A(1'b0), .B(B[228]), .CI(C[228]), .S(S[228]), 
        .CO(C[229]) );
  FA_283 \FAINST[229].FA_  ( .A(1'b0), .B(B[229]), .CI(C[229]), .S(S[229]), 
        .CO(C[230]) );
  FA_282 \FAINST[230].FA_  ( .A(1'b0), .B(B[230]), .CI(C[230]), .S(S[230]), 
        .CO(C[231]) );
  FA_281 \FAINST[231].FA_  ( .A(1'b0), .B(B[231]), .CI(C[231]), .S(S[231]), 
        .CO(C[232]) );
  FA_280 \FAINST[232].FA_  ( .A(1'b0), .B(B[232]), .CI(C[232]), .S(S[232]), 
        .CO(C[233]) );
  FA_279 \FAINST[233].FA_  ( .A(1'b0), .B(B[233]), .CI(C[233]), .S(S[233]), 
        .CO(C[234]) );
  FA_278 \FAINST[234].FA_  ( .A(1'b0), .B(B[234]), .CI(C[234]), .S(S[234]), 
        .CO(C[235]) );
  FA_277 \FAINST[235].FA_  ( .A(1'b0), .B(B[235]), .CI(C[235]), .S(S[235]), 
        .CO(C[236]) );
  FA_276 \FAINST[236].FA_  ( .A(1'b0), .B(B[236]), .CI(C[236]), .S(S[236]), 
        .CO(C[237]) );
  FA_275 \FAINST[237].FA_  ( .A(1'b0), .B(B[237]), .CI(C[237]), .S(S[237]), 
        .CO(C[238]) );
  FA_274 \FAINST[238].FA_  ( .A(1'b0), .B(B[238]), .CI(C[238]), .S(S[238]), 
        .CO(C[239]) );
  FA_273 \FAINST[239].FA_  ( .A(1'b0), .B(B[239]), .CI(C[239]), .S(S[239]), 
        .CO(C[240]) );
  FA_272 \FAINST[240].FA_  ( .A(1'b0), .B(B[240]), .CI(C[240]), .S(S[240]), 
        .CO(C[241]) );
  FA_271 \FAINST[241].FA_  ( .A(1'b0), .B(B[241]), .CI(C[241]), .S(S[241]), 
        .CO(C[242]) );
  FA_270 \FAINST[242].FA_  ( .A(1'b0), .B(B[242]), .CI(C[242]), .S(S[242]), 
        .CO(C[243]) );
  FA_269 \FAINST[243].FA_  ( .A(1'b0), .B(B[243]), .CI(C[243]), .S(S[243]), 
        .CO(C[244]) );
  FA_268 \FAINST[244].FA_  ( .A(1'b0), .B(B[244]), .CI(C[244]), .S(S[244]), 
        .CO(C[245]) );
  FA_267 \FAINST[245].FA_  ( .A(1'b0), .B(B[245]), .CI(C[245]), .S(S[245]), 
        .CO(C[246]) );
  FA_266 \FAINST[246].FA_  ( .A(1'b0), .B(B[246]), .CI(C[246]), .S(S[246]), 
        .CO(C[247]) );
  FA_265 \FAINST[247].FA_  ( .A(1'b0), .B(B[247]), .CI(C[247]), .S(S[247]), 
        .CO(C[248]) );
  FA_264 \FAINST[248].FA_  ( .A(1'b0), .B(B[248]), .CI(C[248]), .S(S[248]), 
        .CO(C[249]) );
  FA_263 \FAINST[249].FA_  ( .A(1'b0), .B(B[249]), .CI(C[249]), .S(S[249]), 
        .CO(C[250]) );
  FA_262 \FAINST[250].FA_  ( .A(1'b0), .B(B[250]), .CI(C[250]), .S(S[250]), 
        .CO(C[251]) );
  FA_261 \FAINST[251].FA_  ( .A(1'b0), .B(B[251]), .CI(C[251]), .S(S[251]), 
        .CO(C[252]) );
  FA_260 \FAINST[252].FA_  ( .A(1'b0), .B(B[252]), .CI(C[252]), .S(S[252]), 
        .CO(C[253]) );
  FA_259 \FAINST[253].FA_  ( .A(1'b0), .B(B[253]), .CI(C[253]), .S(S[253]), 
        .CO(C[254]) );
  FA_258 \FAINST[254].FA_  ( .A(1'b0), .B(B[254]), .CI(C[254]), .S(S[254]) );
  FA_257 \FAINST[255].FA_  ( .A(1'b0), .B(B[255]), .CI(1'b0), .S(S[255]) );
endmodule


module mult_N256_CC8_DW01_add_0 ( A, B, CI, SUM, CO );
  input [285:0] A;
  input [285:0] B;
  output [285:0] SUM;
  input CI;
  output CO;
  wire   \A[30] , \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] ,
         \A[23] , \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] ,
         \A[16] , \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] ,
         \A[8] , \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] ,
         \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272, n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281,
         n1282, n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291,
         n1292, n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301,
         n1302, n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311,
         n1312, n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321,
         n1322, n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331,
         n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341,
         n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351,
         n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361,
         n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371,
         n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381,
         n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391,
         n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441,
         n1442, n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451,
         n1452, n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461,
         n1462, n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471,
         n1472, n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481,
         n1482, n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491,
         n1492, n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501,
         n1502, n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511,
         n1512, n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521,
         n1522, n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531,
         n1532, n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541,
         n1542, n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551,
         n1552, n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561,
         n1562, n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571,
         n1572, n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581,
         n1582, n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591,
         n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601,
         n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611,
         n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621,
         n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631,
         n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641,
         n1642;
  assign SUM[30] = \A[30] ;
  assign \A[30]  = A[30];
  assign SUM[29] = \A[29] ;
  assign \A[29]  = A[29];
  assign SUM[28] = \A[28] ;
  assign \A[28]  = A[28];
  assign SUM[27] = \A[27] ;
  assign \A[27]  = A[27];
  assign SUM[26] = \A[26] ;
  assign \A[26]  = A[26];
  assign SUM[25] = \A[25] ;
  assign \A[25]  = A[25];
  assign SUM[24] = \A[24] ;
  assign \A[24]  = A[24];
  assign SUM[23] = \A[23] ;
  assign \A[23]  = A[23];
  assign SUM[22] = \A[22] ;
  assign \A[22]  = A[22];
  assign SUM[21] = \A[21] ;
  assign \A[21]  = A[21];
  assign SUM[20] = \A[20] ;
  assign \A[20]  = A[20];
  assign SUM[19] = \A[19] ;
  assign \A[19]  = A[19];
  assign SUM[18] = \A[18] ;
  assign \A[18]  = A[18];
  assign SUM[17] = \A[17] ;
  assign \A[17]  = A[17];
  assign SUM[16] = \A[16] ;
  assign \A[16]  = A[16];
  assign SUM[15] = \A[15] ;
  assign \A[15]  = A[15];
  assign SUM[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  NAND U2 ( .A(n15), .B(n18), .Z(n19) );
  XOR U3 ( .A(n1), .B(n2), .Z(SUM[99]) );
  NANDN U4 ( .A(n3), .B(n4), .Z(n2) );
  ANDN U5 ( .B(n5), .A(n6), .Z(n1) );
  NAND U6 ( .A(n7), .B(n8), .Z(n5) );
  XNOR U7 ( .A(n7), .B(n9), .Z(SUM[98]) );
  NANDN U8 ( .A(n6), .B(n8), .Z(n9) );
  NANDN U9 ( .A(n10), .B(n11), .Z(n7) );
  NAND U10 ( .A(n12), .B(n13), .Z(n11) );
  XNOR U11 ( .A(n12), .B(n14), .Z(SUM[97]) );
  NANDN U12 ( .A(n10), .B(n13), .Z(n14) );
  NAND U13 ( .A(n15), .B(n16), .Z(n12) );
  NANDN U14 ( .A(n17), .B(n18), .Z(n16) );
  XOR U15 ( .A(n17), .B(n19), .Z(SUM[96]) );
  XOR U16 ( .A(n20), .B(n21), .Z(SUM[95]) );
  OR U17 ( .A(n22), .B(n23), .Z(n21) );
  ANDN U18 ( .B(n24), .A(n25), .Z(n20) );
  NANDN U19 ( .A(n26), .B(n27), .Z(n24) );
  XNOR U20 ( .A(n27), .B(n28), .Z(SUM[94]) );
  OR U21 ( .A(n26), .B(n25), .Z(n28) );
  NANDN U22 ( .A(n29), .B(n30), .Z(n27) );
  NANDN U23 ( .A(n31), .B(n32), .Z(n30) );
  XNOR U24 ( .A(n32), .B(n33), .Z(SUM[93]) );
  OR U25 ( .A(n31), .B(n29), .Z(n33) );
  NANDN U26 ( .A(n34), .B(n35), .Z(n32) );
  NAND U27 ( .A(n36), .B(n37), .Z(n35) );
  XNOR U28 ( .A(n36), .B(n38), .Z(SUM[92]) );
  NANDN U29 ( .A(n34), .B(n37), .Z(n38) );
  NANDN U30 ( .A(n39), .B(n40), .Z(n36) );
  NANDN U31 ( .A(n41), .B(n42), .Z(n40) );
  XOR U32 ( .A(n43), .B(n44), .Z(SUM[91]) );
  NANDN U33 ( .A(n45), .B(n46), .Z(n44) );
  ANDN U34 ( .B(n47), .A(n48), .Z(n43) );
  NAND U35 ( .A(n49), .B(n50), .Z(n47) );
  XNOR U36 ( .A(n49), .B(n51), .Z(SUM[90]) );
  NANDN U37 ( .A(n48), .B(n50), .Z(n51) );
  NANDN U38 ( .A(n52), .B(n53), .Z(n49) );
  NAND U39 ( .A(n54), .B(n55), .Z(n53) );
  XNOR U40 ( .A(n54), .B(n56), .Z(SUM[89]) );
  NANDN U41 ( .A(n52), .B(n55), .Z(n56) );
  NANDN U42 ( .A(n57), .B(n58), .Z(n54) );
  NAND U43 ( .A(n42), .B(n59), .Z(n58) );
  XNOR U44 ( .A(n42), .B(n60), .Z(SUM[88]) );
  NANDN U45 ( .A(n57), .B(n59), .Z(n60) );
  NANDN U46 ( .A(n61), .B(n62), .Z(n42) );
  NANDN U47 ( .A(n63), .B(n64), .Z(n62) );
  XOR U48 ( .A(n65), .B(n66), .Z(SUM[87]) );
  NANDN U49 ( .A(n67), .B(n68), .Z(n66) );
  ANDN U50 ( .B(n69), .A(n70), .Z(n65) );
  NAND U51 ( .A(n71), .B(n72), .Z(n69) );
  XNOR U52 ( .A(n71), .B(n73), .Z(SUM[86]) );
  NANDN U53 ( .A(n70), .B(n72), .Z(n73) );
  NANDN U54 ( .A(n74), .B(n75), .Z(n71) );
  NAND U55 ( .A(n76), .B(n77), .Z(n75) );
  XNOR U56 ( .A(n76), .B(n78), .Z(SUM[85]) );
  NANDN U57 ( .A(n74), .B(n77), .Z(n78) );
  NANDN U58 ( .A(n79), .B(n80), .Z(n76) );
  NANDN U59 ( .A(n63), .B(n81), .Z(n80) );
  XOR U60 ( .A(n63), .B(n82), .Z(SUM[84]) );
  NANDN U61 ( .A(n79), .B(n81), .Z(n82) );
  ANDN U62 ( .B(n83), .A(n84), .Z(n63) );
  OR U63 ( .A(n85), .B(n86), .Z(n83) );
  XOR U64 ( .A(n87), .B(n88), .Z(SUM[83]) );
  NANDN U65 ( .A(n89), .B(n90), .Z(n88) );
  ANDN U66 ( .B(n91), .A(n92), .Z(n87) );
  NANDN U67 ( .A(n93), .B(n94), .Z(n91) );
  XNOR U68 ( .A(n94), .B(n95), .Z(SUM[82]) );
  OR U69 ( .A(n93), .B(n92), .Z(n95) );
  NANDN U70 ( .A(n96), .B(n97), .Z(n94) );
  NAND U71 ( .A(n98), .B(n99), .Z(n97) );
  XNOR U72 ( .A(n98), .B(n100), .Z(SUM[81]) );
  NANDN U73 ( .A(n96), .B(n99), .Z(n100) );
  NANDN U74 ( .A(n101), .B(n102), .Z(n98) );
  NANDN U75 ( .A(n86), .B(n103), .Z(n102) );
  XOR U76 ( .A(n86), .B(n104), .Z(SUM[80]) );
  NANDN U77 ( .A(n101), .B(n103), .Z(n104) );
  XOR U78 ( .A(n105), .B(n106), .Z(SUM[79]) );
  OR U79 ( .A(n107), .B(n108), .Z(n106) );
  ANDN U80 ( .B(n109), .A(n110), .Z(n105) );
  NANDN U81 ( .A(n111), .B(n112), .Z(n109) );
  XNOR U82 ( .A(n112), .B(n113), .Z(SUM[78]) );
  OR U83 ( .A(n111), .B(n110), .Z(n113) );
  NANDN U84 ( .A(n114), .B(n115), .Z(n112) );
  NANDN U85 ( .A(n116), .B(n117), .Z(n115) );
  XNOR U86 ( .A(n117), .B(n118), .Z(SUM[77]) );
  OR U87 ( .A(n116), .B(n114), .Z(n118) );
  NANDN U88 ( .A(n119), .B(n120), .Z(n117) );
  NAND U89 ( .A(n121), .B(n122), .Z(n120) );
  XNOR U90 ( .A(n121), .B(n123), .Z(SUM[76]) );
  NANDN U91 ( .A(n119), .B(n122), .Z(n123) );
  NANDN U92 ( .A(n124), .B(n125), .Z(n121) );
  NANDN U93 ( .A(n126), .B(n127), .Z(n125) );
  XOR U94 ( .A(n128), .B(n129), .Z(SUM[75]) );
  NANDN U95 ( .A(n130), .B(n131), .Z(n129) );
  ANDN U96 ( .B(n132), .A(n133), .Z(n128) );
  NAND U97 ( .A(n134), .B(n135), .Z(n132) );
  XNOR U98 ( .A(n134), .B(n136), .Z(SUM[74]) );
  NANDN U99 ( .A(n133), .B(n135), .Z(n136) );
  NANDN U100 ( .A(n137), .B(n138), .Z(n134) );
  NAND U101 ( .A(n139), .B(n140), .Z(n138) );
  XNOR U102 ( .A(n139), .B(n141), .Z(SUM[73]) );
  NANDN U103 ( .A(n137), .B(n140), .Z(n141) );
  NANDN U104 ( .A(n142), .B(n143), .Z(n139) );
  NAND U105 ( .A(n127), .B(n144), .Z(n143) );
  XNOR U106 ( .A(n127), .B(n145), .Z(SUM[72]) );
  NANDN U107 ( .A(n142), .B(n144), .Z(n145) );
  NANDN U108 ( .A(n146), .B(n147), .Z(n127) );
  NANDN U109 ( .A(n148), .B(n149), .Z(n147) );
  XOR U110 ( .A(n150), .B(n151), .Z(SUM[71]) );
  NANDN U111 ( .A(n152), .B(n153), .Z(n151) );
  ANDN U112 ( .B(n154), .A(n155), .Z(n150) );
  NAND U113 ( .A(n156), .B(n157), .Z(n154) );
  XNOR U114 ( .A(n156), .B(n158), .Z(SUM[70]) );
  NANDN U115 ( .A(n155), .B(n157), .Z(n158) );
  NANDN U116 ( .A(n159), .B(n160), .Z(n156) );
  NAND U117 ( .A(n161), .B(n162), .Z(n160) );
  XNOR U118 ( .A(n161), .B(n163), .Z(SUM[69]) );
  NANDN U119 ( .A(n159), .B(n162), .Z(n163) );
  NANDN U120 ( .A(n164), .B(n165), .Z(n161) );
  NANDN U121 ( .A(n148), .B(n166), .Z(n165) );
  XOR U122 ( .A(n148), .B(n167), .Z(SUM[68]) );
  NANDN U123 ( .A(n164), .B(n166), .Z(n167) );
  ANDN U124 ( .B(n168), .A(n169), .Z(n148) );
  OR U125 ( .A(n170), .B(n171), .Z(n168) );
  XOR U126 ( .A(n172), .B(n173), .Z(SUM[67]) );
  NANDN U127 ( .A(n174), .B(n175), .Z(n173) );
  ANDN U128 ( .B(n176), .A(n177), .Z(n172) );
  NANDN U129 ( .A(n178), .B(n179), .Z(n176) );
  XNOR U130 ( .A(n179), .B(n180), .Z(SUM[66]) );
  OR U131 ( .A(n178), .B(n177), .Z(n180) );
  NANDN U132 ( .A(n181), .B(n182), .Z(n179) );
  NAND U133 ( .A(n183), .B(n184), .Z(n182) );
  XNOR U134 ( .A(n183), .B(n185), .Z(SUM[65]) );
  NANDN U135 ( .A(n181), .B(n184), .Z(n185) );
  NANDN U136 ( .A(n186), .B(n187), .Z(n183) );
  NANDN U137 ( .A(n171), .B(n188), .Z(n187) );
  XOR U138 ( .A(n171), .B(n189), .Z(SUM[64]) );
  NANDN U139 ( .A(n186), .B(n188), .Z(n189) );
  XOR U140 ( .A(n190), .B(n191), .Z(SUM[63]) );
  OR U141 ( .A(n192), .B(n193), .Z(n191) );
  ANDN U142 ( .B(n194), .A(n195), .Z(n190) );
  NANDN U143 ( .A(n196), .B(n197), .Z(n194) );
  XNOR U144 ( .A(n197), .B(n198), .Z(SUM[62]) );
  OR U145 ( .A(n196), .B(n195), .Z(n198) );
  NANDN U146 ( .A(n199), .B(n200), .Z(n197) );
  NANDN U147 ( .A(n201), .B(n202), .Z(n200) );
  XNOR U148 ( .A(n202), .B(n203), .Z(SUM[61]) );
  OR U149 ( .A(n201), .B(n199), .Z(n203) );
  NANDN U150 ( .A(n204), .B(n205), .Z(n202) );
  NANDN U151 ( .A(n206), .B(n207), .Z(n205) );
  XNOR U152 ( .A(n207), .B(n208), .Z(SUM[60]) );
  OR U153 ( .A(n206), .B(n204), .Z(n208) );
  NANDN U154 ( .A(n209), .B(n210), .Z(n207) );
  NANDN U155 ( .A(n211), .B(n212), .Z(n210) );
  XOR U156 ( .A(n213), .B(n214), .Z(SUM[59]) );
  NANDN U157 ( .A(n215), .B(n216), .Z(n214) );
  ANDN U158 ( .B(n217), .A(n218), .Z(n213) );
  NAND U159 ( .A(n219), .B(n220), .Z(n217) );
  XNOR U160 ( .A(n219), .B(n221), .Z(SUM[58]) );
  NANDN U161 ( .A(n218), .B(n220), .Z(n221) );
  NANDN U162 ( .A(n222), .B(n223), .Z(n219) );
  NAND U163 ( .A(n224), .B(n225), .Z(n223) );
  XNOR U164 ( .A(n224), .B(n226), .Z(SUM[57]) );
  NANDN U165 ( .A(n222), .B(n225), .Z(n226) );
  NANDN U166 ( .A(n227), .B(n228), .Z(n224) );
  NAND U167 ( .A(n212), .B(n229), .Z(n228) );
  XNOR U168 ( .A(n212), .B(n230), .Z(SUM[56]) );
  NANDN U169 ( .A(n227), .B(n229), .Z(n230) );
  NANDN U170 ( .A(n231), .B(n232), .Z(n212) );
  OR U171 ( .A(n233), .B(n234), .Z(n232) );
  XOR U172 ( .A(n235), .B(n236), .Z(SUM[55]) );
  NANDN U173 ( .A(n237), .B(n238), .Z(n236) );
  ANDN U174 ( .B(n239), .A(n240), .Z(n235) );
  NAND U175 ( .A(n241), .B(n242), .Z(n239) );
  XNOR U176 ( .A(n241), .B(n243), .Z(SUM[54]) );
  NANDN U177 ( .A(n240), .B(n242), .Z(n243) );
  NANDN U178 ( .A(n244), .B(n245), .Z(n241) );
  NAND U179 ( .A(n246), .B(n247), .Z(n245) );
  XNOR U180 ( .A(n246), .B(n248), .Z(SUM[53]) );
  NANDN U181 ( .A(n244), .B(n247), .Z(n248) );
  NANDN U182 ( .A(n249), .B(n250), .Z(n246) );
  NANDN U183 ( .A(n234), .B(n251), .Z(n250) );
  XOR U184 ( .A(n234), .B(n252), .Z(SUM[52]) );
  NANDN U185 ( .A(n249), .B(n251), .Z(n252) );
  NOR U186 ( .A(n253), .B(n254), .Z(n234) );
  XOR U187 ( .A(n255), .B(n256), .Z(SUM[51]) );
  NANDN U188 ( .A(n257), .B(n258), .Z(n256) );
  ANDN U189 ( .B(n259), .A(n260), .Z(n255) );
  NAND U190 ( .A(n261), .B(n262), .Z(n259) );
  XNOR U191 ( .A(n261), .B(n263), .Z(SUM[50]) );
  NANDN U192 ( .A(n260), .B(n262), .Z(n263) );
  NANDN U193 ( .A(n264), .B(n265), .Z(n261) );
  NAND U194 ( .A(n266), .B(n267), .Z(n265) );
  XNOR U195 ( .A(n266), .B(n268), .Z(SUM[49]) );
  NANDN U196 ( .A(n264), .B(n267), .Z(n268) );
  NANDN U197 ( .A(n269), .B(n270), .Z(n266) );
  NANDN U198 ( .A(n271), .B(n272), .Z(n270) );
  XOR U199 ( .A(n271), .B(n273), .Z(SUM[48]) );
  NANDN U200 ( .A(n269), .B(n272), .Z(n273) );
  XOR U201 ( .A(n274), .B(n275), .Z(SUM[47]) );
  OR U202 ( .A(n276), .B(n277), .Z(n275) );
  ANDN U203 ( .B(n278), .A(n279), .Z(n274) );
  NANDN U204 ( .A(n280), .B(n281), .Z(n278) );
  XNOR U205 ( .A(n281), .B(n282), .Z(SUM[46]) );
  OR U206 ( .A(n280), .B(n279), .Z(n282) );
  NANDN U207 ( .A(n283), .B(n284), .Z(n281) );
  NANDN U208 ( .A(n285), .B(n286), .Z(n284) );
  XNOR U209 ( .A(n286), .B(n287), .Z(SUM[45]) );
  OR U210 ( .A(n285), .B(n283), .Z(n287) );
  NANDN U211 ( .A(n288), .B(n289), .Z(n286) );
  NAND U212 ( .A(n290), .B(n291), .Z(n289) );
  XNOR U213 ( .A(n290), .B(n292), .Z(SUM[44]) );
  NANDN U214 ( .A(n288), .B(n291), .Z(n292) );
  NANDN U215 ( .A(n293), .B(n294), .Z(n290) );
  NANDN U216 ( .A(n295), .B(n296), .Z(n294) );
  XOR U217 ( .A(n297), .B(n298), .Z(SUM[43]) );
  NANDN U218 ( .A(n299), .B(n300), .Z(n298) );
  ANDN U219 ( .B(n301), .A(n302), .Z(n297) );
  NAND U220 ( .A(n303), .B(n304), .Z(n301) );
  XNOR U221 ( .A(n303), .B(n305), .Z(SUM[42]) );
  NANDN U222 ( .A(n302), .B(n304), .Z(n305) );
  NANDN U223 ( .A(n306), .B(n307), .Z(n303) );
  NAND U224 ( .A(n308), .B(n309), .Z(n307) );
  XNOR U225 ( .A(n308), .B(n310), .Z(SUM[41]) );
  NANDN U226 ( .A(n306), .B(n309), .Z(n310) );
  NANDN U227 ( .A(n311), .B(n312), .Z(n308) );
  NAND U228 ( .A(n296), .B(n313), .Z(n312) );
  XNOR U229 ( .A(n296), .B(n314), .Z(SUM[40]) );
  NANDN U230 ( .A(n311), .B(n313), .Z(n314) );
  NANDN U231 ( .A(n315), .B(n316), .Z(n296) );
  NANDN U232 ( .A(n317), .B(n318), .Z(n316) );
  XOR U233 ( .A(n319), .B(n320), .Z(SUM[39]) );
  NANDN U234 ( .A(n321), .B(n322), .Z(n320) );
  ANDN U235 ( .B(n323), .A(n324), .Z(n319) );
  NAND U236 ( .A(n325), .B(n326), .Z(n323) );
  XNOR U237 ( .A(n325), .B(n327), .Z(SUM[38]) );
  NANDN U238 ( .A(n324), .B(n326), .Z(n327) );
  NANDN U239 ( .A(n328), .B(n329), .Z(n325) );
  NAND U240 ( .A(n330), .B(n331), .Z(n329) );
  XNOR U241 ( .A(n330), .B(n332), .Z(SUM[37]) );
  NANDN U242 ( .A(n328), .B(n331), .Z(n332) );
  NANDN U243 ( .A(n333), .B(n334), .Z(n330) );
  NANDN U244 ( .A(n317), .B(n335), .Z(n334) );
  XOR U245 ( .A(n317), .B(n336), .Z(SUM[36]) );
  NANDN U246 ( .A(n333), .B(n335), .Z(n336) );
  ANDN U247 ( .B(n337), .A(n338), .Z(n317) );
  NANDN U248 ( .A(n339), .B(n340), .Z(n337) );
  XOR U249 ( .A(n341), .B(n342), .Z(SUM[35]) );
  NANDN U250 ( .A(n343), .B(n344), .Z(n342) );
  ANDN U251 ( .B(n345), .A(n346), .Z(n341) );
  NANDN U252 ( .A(n347), .B(n348), .Z(n345) );
  XNOR U253 ( .A(n348), .B(n349), .Z(SUM[34]) );
  OR U254 ( .A(n347), .B(n346), .Z(n349) );
  NANDN U255 ( .A(n350), .B(n351), .Z(n348) );
  NAND U256 ( .A(n352), .B(n353), .Z(n351) );
  XNOR U257 ( .A(n352), .B(n354), .Z(SUM[33]) );
  NANDN U258 ( .A(n350), .B(n353), .Z(n354) );
  NANDN U259 ( .A(n355), .B(n356), .Z(n352) );
  NAND U260 ( .A(n357), .B(n340), .Z(n356) );
  XOR U261 ( .A(n340), .B(n358), .Z(SUM[32]) );
  ANDN U262 ( .B(n357), .A(n355), .Z(n358) );
  ANDN U263 ( .B(n359), .A(n340), .Z(SUM[31]) );
  OR U264 ( .A(A[31]), .B(B[31]), .Z(n359) );
  XOR U265 ( .A(n360), .B(n361), .Z(SUM[253]) );
  XNOR U266 ( .A(B[253]), .B(A[253]), .Z(n361) );
  ANDN U267 ( .B(n362), .A(n363), .Z(n360) );
  NAND U268 ( .A(n364), .B(n365), .Z(n362) );
  XNOR U269 ( .A(n364), .B(n366), .Z(SUM[252]) );
  NANDN U270 ( .A(n363), .B(n365), .Z(n366) );
  OR U271 ( .A(B[252]), .B(A[252]), .Z(n365) );
  AND U272 ( .A(B[252]), .B(A[252]), .Z(n363) );
  NANDN U273 ( .A(n367), .B(n368), .Z(n364) );
  NAND U274 ( .A(n369), .B(n370), .Z(n368) );
  XNOR U275 ( .A(n369), .B(n371), .Z(SUM[251]) );
  NANDN U276 ( .A(n367), .B(n370), .Z(n371) );
  OR U277 ( .A(B[251]), .B(A[251]), .Z(n370) );
  AND U278 ( .A(B[251]), .B(A[251]), .Z(n367) );
  NANDN U279 ( .A(n372), .B(n373), .Z(n369) );
  NAND U280 ( .A(n374), .B(n375), .Z(n373) );
  XNOR U281 ( .A(n374), .B(n376), .Z(SUM[250]) );
  NANDN U282 ( .A(n372), .B(n375), .Z(n376) );
  OR U283 ( .A(B[250]), .B(A[250]), .Z(n375) );
  AND U284 ( .A(B[250]), .B(A[250]), .Z(n372) );
  NANDN U285 ( .A(n377), .B(n378), .Z(n374) );
  NAND U286 ( .A(n379), .B(n380), .Z(n378) );
  XNOR U287 ( .A(n379), .B(n381), .Z(SUM[249]) );
  NANDN U288 ( .A(n377), .B(n380), .Z(n381) );
  OR U289 ( .A(B[249]), .B(A[249]), .Z(n380) );
  AND U290 ( .A(B[249]), .B(A[249]), .Z(n377) );
  NANDN U291 ( .A(n382), .B(n383), .Z(n379) );
  NAND U292 ( .A(n384), .B(n385), .Z(n383) );
  XNOR U293 ( .A(n384), .B(n386), .Z(SUM[248]) );
  NANDN U294 ( .A(n382), .B(n385), .Z(n386) );
  OR U295 ( .A(B[248]), .B(A[248]), .Z(n385) );
  AND U296 ( .A(B[248]), .B(A[248]), .Z(n382) );
  NANDN U297 ( .A(n387), .B(n388), .Z(n384) );
  NAND U298 ( .A(n389), .B(n390), .Z(n388) );
  XNOR U299 ( .A(n389), .B(n391), .Z(SUM[247]) );
  NANDN U300 ( .A(n387), .B(n390), .Z(n391) );
  OR U301 ( .A(B[247]), .B(A[247]), .Z(n390) );
  AND U302 ( .A(B[247]), .B(A[247]), .Z(n387) );
  NANDN U303 ( .A(n392), .B(n393), .Z(n389) );
  NAND U304 ( .A(n394), .B(n395), .Z(n393) );
  XNOR U305 ( .A(n394), .B(n396), .Z(SUM[246]) );
  NANDN U306 ( .A(n392), .B(n395), .Z(n396) );
  OR U307 ( .A(B[246]), .B(A[246]), .Z(n395) );
  AND U308 ( .A(B[246]), .B(A[246]), .Z(n392) );
  NANDN U309 ( .A(n397), .B(n398), .Z(n394) );
  NAND U310 ( .A(n399), .B(n400), .Z(n398) );
  XNOR U311 ( .A(n399), .B(n401), .Z(SUM[245]) );
  NANDN U312 ( .A(n397), .B(n400), .Z(n401) );
  OR U313 ( .A(B[245]), .B(A[245]), .Z(n400) );
  AND U314 ( .A(B[245]), .B(A[245]), .Z(n397) );
  NANDN U315 ( .A(n402), .B(n403), .Z(n399) );
  NAND U316 ( .A(n404), .B(n405), .Z(n403) );
  XNOR U317 ( .A(n404), .B(n406), .Z(SUM[244]) );
  NANDN U318 ( .A(n402), .B(n405), .Z(n406) );
  OR U319 ( .A(B[244]), .B(A[244]), .Z(n405) );
  AND U320 ( .A(B[244]), .B(A[244]), .Z(n402) );
  NANDN U321 ( .A(n407), .B(n408), .Z(n404) );
  NAND U322 ( .A(n409), .B(n410), .Z(n408) );
  XNOR U323 ( .A(n409), .B(n411), .Z(SUM[243]) );
  NANDN U324 ( .A(n407), .B(n410), .Z(n411) );
  OR U325 ( .A(B[243]), .B(A[243]), .Z(n410) );
  AND U326 ( .A(B[243]), .B(A[243]), .Z(n407) );
  NANDN U327 ( .A(n412), .B(n413), .Z(n409) );
  NAND U328 ( .A(n414), .B(n415), .Z(n413) );
  XNOR U329 ( .A(n414), .B(n416), .Z(SUM[242]) );
  NANDN U330 ( .A(n412), .B(n415), .Z(n416) );
  OR U331 ( .A(B[242]), .B(A[242]), .Z(n415) );
  AND U332 ( .A(B[242]), .B(A[242]), .Z(n412) );
  NANDN U333 ( .A(n417), .B(n418), .Z(n414) );
  NAND U334 ( .A(n419), .B(n420), .Z(n418) );
  XNOR U335 ( .A(n419), .B(n421), .Z(SUM[241]) );
  NANDN U336 ( .A(n417), .B(n420), .Z(n421) );
  OR U337 ( .A(B[241]), .B(A[241]), .Z(n420) );
  AND U338 ( .A(B[241]), .B(A[241]), .Z(n417) );
  NANDN U339 ( .A(n422), .B(n423), .Z(n419) );
  NAND U340 ( .A(n424), .B(n425), .Z(n423) );
  XNOR U341 ( .A(n424), .B(n426), .Z(SUM[240]) );
  NANDN U342 ( .A(n422), .B(n425), .Z(n426) );
  OR U343 ( .A(B[240]), .B(A[240]), .Z(n425) );
  AND U344 ( .A(B[240]), .B(A[240]), .Z(n422) );
  NANDN U345 ( .A(n427), .B(n428), .Z(n424) );
  NANDN U346 ( .A(n429), .B(n430), .Z(n428) );
  NANDN U347 ( .A(n431), .B(n432), .Z(n430) );
  NANDN U348 ( .A(n433), .B(n434), .Z(n432) );
  NANDN U349 ( .A(n435), .B(n436), .Z(n434) );
  NANDN U350 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U351 ( .A(n439), .B(n440), .Z(n438) );
  NANDN U352 ( .A(n441), .B(n442), .Z(n440) );
  NANDN U353 ( .A(n443), .B(n444), .Z(n442) );
  NANDN U354 ( .A(n445), .B(n446), .Z(n444) );
  NANDN U355 ( .A(n447), .B(n448), .Z(n446) );
  AND U356 ( .A(n449), .B(n450), .Z(n448) );
  NANDN U357 ( .A(n451), .B(n452), .Z(n450) );
  NANDN U358 ( .A(n451), .B(n453), .Z(n449) );
  XOR U359 ( .A(n454), .B(n455), .Z(SUM[239]) );
  OR U360 ( .A(n429), .B(n427), .Z(n455) );
  AND U361 ( .A(B[239]), .B(A[239]), .Z(n427) );
  NOR U362 ( .A(B[239]), .B(A[239]), .Z(n429) );
  ANDN U363 ( .B(n456), .A(n431), .Z(n454) );
  NANDN U364 ( .A(n433), .B(n457), .Z(n456) );
  XNOR U365 ( .A(n457), .B(n458), .Z(SUM[238]) );
  OR U366 ( .A(n433), .B(n431), .Z(n458) );
  AND U367 ( .A(B[238]), .B(A[238]), .Z(n431) );
  NOR U368 ( .A(B[238]), .B(A[238]), .Z(n433) );
  NANDN U369 ( .A(n435), .B(n459), .Z(n457) );
  NANDN U370 ( .A(n437), .B(n460), .Z(n459) );
  XNOR U371 ( .A(n460), .B(n461), .Z(SUM[237]) );
  OR U372 ( .A(n437), .B(n435), .Z(n461) );
  AND U373 ( .A(B[237]), .B(A[237]), .Z(n435) );
  NOR U374 ( .A(B[237]), .B(A[237]), .Z(n437) );
  NANDN U375 ( .A(n439), .B(n462), .Z(n460) );
  NANDN U376 ( .A(n441), .B(n463), .Z(n462) );
  XNOR U377 ( .A(n463), .B(n464), .Z(SUM[236]) );
  OR U378 ( .A(n441), .B(n439), .Z(n464) );
  AND U379 ( .A(B[236]), .B(A[236]), .Z(n439) );
  NOR U380 ( .A(B[236]), .B(A[236]), .Z(n441) );
  NANDN U381 ( .A(n443), .B(n465), .Z(n463) );
  NANDN U382 ( .A(n445), .B(n466), .Z(n465) );
  NAND U383 ( .A(n467), .B(n468), .Z(n445) );
  AND U384 ( .A(n469), .B(n470), .Z(n468) );
  AND U385 ( .A(n471), .B(n472), .Z(n467) );
  NANDN U386 ( .A(n473), .B(n474), .Z(n443) );
  NAND U387 ( .A(n475), .B(n472), .Z(n474) );
  NANDN U388 ( .A(n476), .B(n477), .Z(n475) );
  NAND U389 ( .A(n478), .B(n471), .Z(n477) );
  NANDN U390 ( .A(n479), .B(n480), .Z(n478) );
  NAND U391 ( .A(n470), .B(n481), .Z(n480) );
  XOR U392 ( .A(n482), .B(n483), .Z(SUM[235]) );
  NANDN U393 ( .A(n473), .B(n472), .Z(n483) );
  OR U394 ( .A(B[235]), .B(A[235]), .Z(n472) );
  AND U395 ( .A(B[235]), .B(A[235]), .Z(n473) );
  ANDN U396 ( .B(n484), .A(n476), .Z(n482) );
  NAND U397 ( .A(n485), .B(n471), .Z(n484) );
  XNOR U398 ( .A(n485), .B(n486), .Z(SUM[234]) );
  NANDN U399 ( .A(n476), .B(n471), .Z(n486) );
  OR U400 ( .A(B[234]), .B(A[234]), .Z(n471) );
  AND U401 ( .A(B[234]), .B(A[234]), .Z(n476) );
  NANDN U402 ( .A(n479), .B(n487), .Z(n485) );
  NAND U403 ( .A(n488), .B(n470), .Z(n487) );
  XNOR U404 ( .A(n488), .B(n489), .Z(SUM[233]) );
  NANDN U405 ( .A(n479), .B(n470), .Z(n489) );
  OR U406 ( .A(B[233]), .B(A[233]), .Z(n470) );
  AND U407 ( .A(B[233]), .B(A[233]), .Z(n479) );
  NANDN U408 ( .A(n481), .B(n490), .Z(n488) );
  NAND U409 ( .A(n466), .B(n469), .Z(n490) );
  XNOR U410 ( .A(n466), .B(n491), .Z(SUM[232]) );
  NANDN U411 ( .A(n481), .B(n469), .Z(n491) );
  OR U412 ( .A(B[232]), .B(A[232]), .Z(n469) );
  AND U413 ( .A(B[232]), .B(A[232]), .Z(n481) );
  NANDN U414 ( .A(n447), .B(n492), .Z(n466) );
  OR U415 ( .A(n451), .B(n493), .Z(n492) );
  NAND U416 ( .A(n494), .B(n495), .Z(n451) );
  AND U417 ( .A(n496), .B(n497), .Z(n495) );
  AND U418 ( .A(n498), .B(n499), .Z(n494) );
  NANDN U419 ( .A(n500), .B(n501), .Z(n447) );
  NAND U420 ( .A(n502), .B(n499), .Z(n501) );
  NANDN U421 ( .A(n503), .B(n504), .Z(n502) );
  NAND U422 ( .A(n505), .B(n498), .Z(n504) );
  NANDN U423 ( .A(n506), .B(n507), .Z(n505) );
  NAND U424 ( .A(n497), .B(n508), .Z(n507) );
  XOR U425 ( .A(n509), .B(n510), .Z(SUM[231]) );
  NANDN U426 ( .A(n500), .B(n499), .Z(n510) );
  OR U427 ( .A(B[231]), .B(A[231]), .Z(n499) );
  AND U428 ( .A(B[231]), .B(A[231]), .Z(n500) );
  ANDN U429 ( .B(n511), .A(n503), .Z(n509) );
  NAND U430 ( .A(n512), .B(n498), .Z(n511) );
  XNOR U431 ( .A(n512), .B(n513), .Z(SUM[230]) );
  NANDN U432 ( .A(n503), .B(n498), .Z(n513) );
  OR U433 ( .A(A[230]), .B(B[230]), .Z(n498) );
  AND U434 ( .A(A[230]), .B(B[230]), .Z(n503) );
  NANDN U435 ( .A(n506), .B(n514), .Z(n512) );
  NAND U436 ( .A(n515), .B(n497), .Z(n514) );
  XNOR U437 ( .A(n515), .B(n516), .Z(SUM[229]) );
  NANDN U438 ( .A(n506), .B(n497), .Z(n516) );
  OR U439 ( .A(A[229]), .B(B[229]), .Z(n497) );
  AND U440 ( .A(A[229]), .B(B[229]), .Z(n506) );
  NANDN U441 ( .A(n508), .B(n517), .Z(n515) );
  NANDN U442 ( .A(n493), .B(n496), .Z(n517) );
  XOR U443 ( .A(n493), .B(n518), .Z(SUM[228]) );
  NANDN U444 ( .A(n508), .B(n496), .Z(n518) );
  OR U445 ( .A(A[228]), .B(B[228]), .Z(n496) );
  AND U446 ( .A(A[228]), .B(B[228]), .Z(n508) );
  NOR U447 ( .A(n452), .B(n453), .Z(n493) );
  AND U448 ( .A(n519), .B(n520), .Z(n453) );
  AND U449 ( .A(n521), .B(n522), .Z(n520) );
  NOR U450 ( .A(n523), .B(n524), .Z(n522) );
  AND U451 ( .A(n525), .B(n526), .Z(n519) );
  NANDN U452 ( .A(n527), .B(n528), .Z(n452) );
  NAND U453 ( .A(n529), .B(n526), .Z(n528) );
  NANDN U454 ( .A(n530), .B(n531), .Z(n529) );
  NAND U455 ( .A(n532), .B(n525), .Z(n531) );
  NANDN U456 ( .A(n533), .B(n534), .Z(n532) );
  NAND U457 ( .A(n521), .B(n535), .Z(n534) );
  XOR U458 ( .A(n536), .B(n537), .Z(SUM[227]) );
  NANDN U459 ( .A(n527), .B(n526), .Z(n537) );
  OR U460 ( .A(B[227]), .B(A[227]), .Z(n526) );
  AND U461 ( .A(B[227]), .B(A[227]), .Z(n527) );
  ANDN U462 ( .B(n538), .A(n530), .Z(n536) );
  NAND U463 ( .A(n539), .B(n525), .Z(n538) );
  XNOR U464 ( .A(n539), .B(n540), .Z(SUM[226]) );
  NANDN U465 ( .A(n530), .B(n525), .Z(n540) );
  OR U466 ( .A(A[226]), .B(B[226]), .Z(n525) );
  AND U467 ( .A(A[226]), .B(B[226]), .Z(n530) );
  NANDN U468 ( .A(n533), .B(n541), .Z(n539) );
  NAND U469 ( .A(n542), .B(n521), .Z(n541) );
  XNOR U470 ( .A(n542), .B(n543), .Z(SUM[225]) );
  NANDN U471 ( .A(n533), .B(n521), .Z(n543) );
  OR U472 ( .A(A[225]), .B(B[225]), .Z(n521) );
  AND U473 ( .A(A[225]), .B(B[225]), .Z(n533) );
  NANDN U474 ( .A(n535), .B(n544), .Z(n542) );
  OR U475 ( .A(n523), .B(n524), .Z(n544) );
  XOR U476 ( .A(n523), .B(n545), .Z(SUM[224]) );
  OR U477 ( .A(n524), .B(n535), .Z(n545) );
  AND U478 ( .A(A[224]), .B(B[224]), .Z(n535) );
  NOR U479 ( .A(B[224]), .B(A[224]), .Z(n524) );
  ANDN U480 ( .B(n546), .A(n547), .Z(n523) );
  NANDN U481 ( .A(n548), .B(n549), .Z(n546) );
  NANDN U482 ( .A(n550), .B(n551), .Z(n549) );
  NANDN U483 ( .A(n552), .B(n553), .Z(n551) );
  NANDN U484 ( .A(n554), .B(n555), .Z(n553) );
  NANDN U485 ( .A(n556), .B(n557), .Z(n555) );
  NANDN U486 ( .A(n558), .B(n559), .Z(n557) );
  NANDN U487 ( .A(n560), .B(n561), .Z(n559) );
  NANDN U488 ( .A(n562), .B(n563), .Z(n561) );
  NANDN U489 ( .A(n564), .B(n565), .Z(n563) );
  NANDN U490 ( .A(n566), .B(n567), .Z(n565) );
  AND U491 ( .A(n568), .B(n569), .Z(n567) );
  NANDN U492 ( .A(n570), .B(n571), .Z(n569) );
  NANDN U493 ( .A(n570), .B(n572), .Z(n568) );
  XOR U494 ( .A(n573), .B(n574), .Z(SUM[223]) );
  OR U495 ( .A(n548), .B(n547), .Z(n574) );
  AND U496 ( .A(B[223]), .B(A[223]), .Z(n547) );
  NOR U497 ( .A(B[223]), .B(A[223]), .Z(n548) );
  ANDN U498 ( .B(n575), .A(n550), .Z(n573) );
  NANDN U499 ( .A(n552), .B(n576), .Z(n575) );
  XNOR U500 ( .A(n576), .B(n577), .Z(SUM[222]) );
  OR U501 ( .A(n552), .B(n550), .Z(n577) );
  AND U502 ( .A(B[222]), .B(A[222]), .Z(n550) );
  NOR U503 ( .A(B[222]), .B(A[222]), .Z(n552) );
  NANDN U504 ( .A(n554), .B(n578), .Z(n576) );
  NANDN U505 ( .A(n556), .B(n579), .Z(n578) );
  XNOR U506 ( .A(n579), .B(n580), .Z(SUM[221]) );
  OR U507 ( .A(n556), .B(n554), .Z(n580) );
  AND U508 ( .A(B[221]), .B(A[221]), .Z(n554) );
  NOR U509 ( .A(B[221]), .B(A[221]), .Z(n556) );
  NANDN U510 ( .A(n558), .B(n581), .Z(n579) );
  NANDN U511 ( .A(n560), .B(n582), .Z(n581) );
  XNOR U512 ( .A(n582), .B(n583), .Z(SUM[220]) );
  OR U513 ( .A(n560), .B(n558), .Z(n583) );
  AND U514 ( .A(B[220]), .B(A[220]), .Z(n558) );
  NOR U515 ( .A(B[220]), .B(A[220]), .Z(n560) );
  NANDN U516 ( .A(n562), .B(n584), .Z(n582) );
  NANDN U517 ( .A(n564), .B(n585), .Z(n584) );
  NAND U518 ( .A(n586), .B(n587), .Z(n564) );
  AND U519 ( .A(n588), .B(n589), .Z(n587) );
  AND U520 ( .A(n590), .B(n591), .Z(n586) );
  NANDN U521 ( .A(n592), .B(n593), .Z(n562) );
  NAND U522 ( .A(n594), .B(n591), .Z(n593) );
  NANDN U523 ( .A(n595), .B(n596), .Z(n594) );
  NAND U524 ( .A(n597), .B(n590), .Z(n596) );
  NANDN U525 ( .A(n598), .B(n599), .Z(n597) );
  NAND U526 ( .A(n589), .B(n600), .Z(n599) );
  XOR U527 ( .A(n601), .B(n602), .Z(SUM[219]) );
  NANDN U528 ( .A(n592), .B(n591), .Z(n602) );
  OR U529 ( .A(B[219]), .B(A[219]), .Z(n591) );
  AND U530 ( .A(B[219]), .B(A[219]), .Z(n592) );
  ANDN U531 ( .B(n603), .A(n595), .Z(n601) );
  NAND U532 ( .A(n604), .B(n590), .Z(n603) );
  XNOR U533 ( .A(n604), .B(n605), .Z(SUM[218]) );
  NANDN U534 ( .A(n595), .B(n590), .Z(n605) );
  OR U535 ( .A(B[218]), .B(A[218]), .Z(n590) );
  AND U536 ( .A(B[218]), .B(A[218]), .Z(n595) );
  NANDN U537 ( .A(n598), .B(n606), .Z(n604) );
  NAND U538 ( .A(n607), .B(n589), .Z(n606) );
  XNOR U539 ( .A(n607), .B(n608), .Z(SUM[217]) );
  NANDN U540 ( .A(n598), .B(n589), .Z(n608) );
  OR U541 ( .A(B[217]), .B(A[217]), .Z(n589) );
  AND U542 ( .A(B[217]), .B(A[217]), .Z(n598) );
  NANDN U543 ( .A(n600), .B(n609), .Z(n607) );
  NAND U544 ( .A(n585), .B(n588), .Z(n609) );
  XNOR U545 ( .A(n585), .B(n610), .Z(SUM[216]) );
  NANDN U546 ( .A(n600), .B(n588), .Z(n610) );
  OR U547 ( .A(B[216]), .B(A[216]), .Z(n588) );
  AND U548 ( .A(B[216]), .B(A[216]), .Z(n600) );
  NANDN U549 ( .A(n566), .B(n611), .Z(n585) );
  OR U550 ( .A(n570), .B(n612), .Z(n611) );
  NAND U551 ( .A(n613), .B(n614), .Z(n570) );
  AND U552 ( .A(n615), .B(n616), .Z(n614) );
  AND U553 ( .A(n617), .B(n618), .Z(n613) );
  NANDN U554 ( .A(n619), .B(n620), .Z(n566) );
  NAND U555 ( .A(n621), .B(n618), .Z(n620) );
  NANDN U556 ( .A(n622), .B(n623), .Z(n621) );
  NAND U557 ( .A(n624), .B(n617), .Z(n623) );
  NANDN U558 ( .A(n625), .B(n626), .Z(n624) );
  NAND U559 ( .A(n616), .B(n627), .Z(n626) );
  XOR U560 ( .A(n628), .B(n629), .Z(SUM[215]) );
  NANDN U561 ( .A(n619), .B(n618), .Z(n629) );
  OR U562 ( .A(B[215]), .B(A[215]), .Z(n618) );
  AND U563 ( .A(B[215]), .B(A[215]), .Z(n619) );
  ANDN U564 ( .B(n630), .A(n622), .Z(n628) );
  NAND U565 ( .A(n631), .B(n617), .Z(n630) );
  XNOR U566 ( .A(n631), .B(n632), .Z(SUM[214]) );
  NANDN U567 ( .A(n622), .B(n617), .Z(n632) );
  OR U568 ( .A(A[214]), .B(B[214]), .Z(n617) );
  AND U569 ( .A(A[214]), .B(B[214]), .Z(n622) );
  NANDN U570 ( .A(n625), .B(n633), .Z(n631) );
  NAND U571 ( .A(n634), .B(n616), .Z(n633) );
  XNOR U572 ( .A(n634), .B(n635), .Z(SUM[213]) );
  NANDN U573 ( .A(n625), .B(n616), .Z(n635) );
  OR U574 ( .A(A[213]), .B(B[213]), .Z(n616) );
  AND U575 ( .A(A[213]), .B(B[213]), .Z(n625) );
  NANDN U576 ( .A(n627), .B(n636), .Z(n634) );
  NANDN U577 ( .A(n612), .B(n615), .Z(n636) );
  XOR U578 ( .A(n612), .B(n637), .Z(SUM[212]) );
  NANDN U579 ( .A(n627), .B(n615), .Z(n637) );
  OR U580 ( .A(A[212]), .B(B[212]), .Z(n615) );
  AND U581 ( .A(A[212]), .B(B[212]), .Z(n627) );
  NOR U582 ( .A(n571), .B(n572), .Z(n612) );
  AND U583 ( .A(n638), .B(n639), .Z(n572) );
  AND U584 ( .A(n640), .B(n641), .Z(n639) );
  NOR U585 ( .A(n642), .B(n643), .Z(n641) );
  AND U586 ( .A(n644), .B(n645), .Z(n638) );
  NANDN U587 ( .A(n646), .B(n647), .Z(n571) );
  NAND U588 ( .A(n648), .B(n645), .Z(n647) );
  NANDN U589 ( .A(n649), .B(n650), .Z(n648) );
  NAND U590 ( .A(n651), .B(n644), .Z(n650) );
  NANDN U591 ( .A(n652), .B(n653), .Z(n651) );
  NAND U592 ( .A(n640), .B(n654), .Z(n653) );
  XOR U593 ( .A(n655), .B(n656), .Z(SUM[211]) );
  NANDN U594 ( .A(n646), .B(n645), .Z(n656) );
  OR U595 ( .A(B[211]), .B(A[211]), .Z(n645) );
  AND U596 ( .A(B[211]), .B(A[211]), .Z(n646) );
  ANDN U597 ( .B(n657), .A(n649), .Z(n655) );
  NAND U598 ( .A(n658), .B(n644), .Z(n657) );
  XNOR U599 ( .A(n658), .B(n659), .Z(SUM[210]) );
  NANDN U600 ( .A(n649), .B(n644), .Z(n659) );
  OR U601 ( .A(A[210]), .B(B[210]), .Z(n644) );
  AND U602 ( .A(A[210]), .B(B[210]), .Z(n649) );
  NANDN U603 ( .A(n652), .B(n660), .Z(n658) );
  NAND U604 ( .A(n661), .B(n640), .Z(n660) );
  XNOR U605 ( .A(n661), .B(n662), .Z(SUM[209]) );
  NANDN U606 ( .A(n652), .B(n640), .Z(n662) );
  OR U607 ( .A(A[209]), .B(B[209]), .Z(n640) );
  AND U608 ( .A(A[209]), .B(B[209]), .Z(n652) );
  NANDN U609 ( .A(n654), .B(n663), .Z(n661) );
  OR U610 ( .A(n642), .B(n643), .Z(n663) );
  XOR U611 ( .A(n642), .B(n664), .Z(SUM[208]) );
  OR U612 ( .A(n643), .B(n654), .Z(n664) );
  AND U613 ( .A(A[208]), .B(B[208]), .Z(n654) );
  NOR U614 ( .A(B[208]), .B(A[208]), .Z(n643) );
  ANDN U615 ( .B(n665), .A(n666), .Z(n642) );
  NANDN U616 ( .A(n667), .B(n668), .Z(n665) );
  NANDN U617 ( .A(n669), .B(n670), .Z(n668) );
  NANDN U618 ( .A(n671), .B(n672), .Z(n670) );
  NANDN U619 ( .A(n673), .B(n674), .Z(n672) );
  NANDN U620 ( .A(n675), .B(n676), .Z(n674) );
  NANDN U621 ( .A(n677), .B(n678), .Z(n676) );
  NANDN U622 ( .A(n679), .B(n680), .Z(n678) );
  NANDN U623 ( .A(n681), .B(n682), .Z(n680) );
  NANDN U624 ( .A(n683), .B(n684), .Z(n682) );
  NANDN U625 ( .A(n685), .B(n686), .Z(n684) );
  AND U626 ( .A(n687), .B(n688), .Z(n686) );
  NANDN U627 ( .A(n689), .B(n690), .Z(n688) );
  NANDN U628 ( .A(n689), .B(n691), .Z(n687) );
  XOR U629 ( .A(n692), .B(n693), .Z(SUM[207]) );
  OR U630 ( .A(n667), .B(n666), .Z(n693) );
  AND U631 ( .A(B[207]), .B(A[207]), .Z(n666) );
  NOR U632 ( .A(B[207]), .B(A[207]), .Z(n667) );
  ANDN U633 ( .B(n694), .A(n669), .Z(n692) );
  NANDN U634 ( .A(n671), .B(n695), .Z(n694) );
  XNOR U635 ( .A(n695), .B(n696), .Z(SUM[206]) );
  OR U636 ( .A(n671), .B(n669), .Z(n696) );
  AND U637 ( .A(B[206]), .B(A[206]), .Z(n669) );
  NOR U638 ( .A(B[206]), .B(A[206]), .Z(n671) );
  NANDN U639 ( .A(n673), .B(n697), .Z(n695) );
  NANDN U640 ( .A(n675), .B(n698), .Z(n697) );
  XNOR U641 ( .A(n698), .B(n699), .Z(SUM[205]) );
  OR U642 ( .A(n675), .B(n673), .Z(n699) );
  AND U643 ( .A(B[205]), .B(A[205]), .Z(n673) );
  NOR U644 ( .A(B[205]), .B(A[205]), .Z(n675) );
  NANDN U645 ( .A(n677), .B(n700), .Z(n698) );
  NANDN U646 ( .A(n679), .B(n701), .Z(n700) );
  XNOR U647 ( .A(n701), .B(n702), .Z(SUM[204]) );
  OR U648 ( .A(n679), .B(n677), .Z(n702) );
  AND U649 ( .A(B[204]), .B(A[204]), .Z(n677) );
  NOR U650 ( .A(B[204]), .B(A[204]), .Z(n679) );
  NANDN U651 ( .A(n681), .B(n703), .Z(n701) );
  NANDN U652 ( .A(n683), .B(n704), .Z(n703) );
  NAND U653 ( .A(n705), .B(n706), .Z(n683) );
  AND U654 ( .A(n707), .B(n708), .Z(n706) );
  AND U655 ( .A(n709), .B(n710), .Z(n705) );
  NANDN U656 ( .A(n711), .B(n712), .Z(n681) );
  NAND U657 ( .A(n713), .B(n710), .Z(n712) );
  NANDN U658 ( .A(n714), .B(n715), .Z(n713) );
  NAND U659 ( .A(n716), .B(n709), .Z(n715) );
  NANDN U660 ( .A(n717), .B(n718), .Z(n716) );
  NAND U661 ( .A(n708), .B(n719), .Z(n718) );
  XOR U662 ( .A(n720), .B(n721), .Z(SUM[203]) );
  NANDN U663 ( .A(n711), .B(n710), .Z(n721) );
  OR U664 ( .A(B[203]), .B(A[203]), .Z(n710) );
  AND U665 ( .A(B[203]), .B(A[203]), .Z(n711) );
  ANDN U666 ( .B(n722), .A(n714), .Z(n720) );
  NAND U667 ( .A(n723), .B(n709), .Z(n722) );
  XNOR U668 ( .A(n723), .B(n724), .Z(SUM[202]) );
  NANDN U669 ( .A(n714), .B(n709), .Z(n724) );
  OR U670 ( .A(B[202]), .B(A[202]), .Z(n709) );
  AND U671 ( .A(B[202]), .B(A[202]), .Z(n714) );
  NANDN U672 ( .A(n717), .B(n725), .Z(n723) );
  NAND U673 ( .A(n726), .B(n708), .Z(n725) );
  XNOR U674 ( .A(n726), .B(n727), .Z(SUM[201]) );
  NANDN U675 ( .A(n717), .B(n708), .Z(n727) );
  OR U676 ( .A(B[201]), .B(A[201]), .Z(n708) );
  AND U677 ( .A(B[201]), .B(A[201]), .Z(n717) );
  NANDN U678 ( .A(n719), .B(n728), .Z(n726) );
  NAND U679 ( .A(n704), .B(n707), .Z(n728) );
  XNOR U680 ( .A(n704), .B(n729), .Z(SUM[200]) );
  NANDN U681 ( .A(n719), .B(n707), .Z(n729) );
  OR U682 ( .A(B[200]), .B(A[200]), .Z(n707) );
  AND U683 ( .A(B[200]), .B(A[200]), .Z(n719) );
  NANDN U684 ( .A(n685), .B(n730), .Z(n704) );
  OR U685 ( .A(n689), .B(n731), .Z(n730) );
  NAND U686 ( .A(n732), .B(n733), .Z(n689) );
  AND U687 ( .A(n734), .B(n735), .Z(n733) );
  AND U688 ( .A(n736), .B(n737), .Z(n732) );
  NANDN U689 ( .A(n738), .B(n739), .Z(n685) );
  NAND U690 ( .A(n740), .B(n737), .Z(n739) );
  NANDN U691 ( .A(n741), .B(n742), .Z(n740) );
  NAND U692 ( .A(n743), .B(n736), .Z(n742) );
  NANDN U693 ( .A(n744), .B(n745), .Z(n743) );
  NAND U694 ( .A(n735), .B(n746), .Z(n745) );
  XOR U695 ( .A(n747), .B(n748), .Z(SUM[199]) );
  NANDN U696 ( .A(n738), .B(n737), .Z(n748) );
  OR U697 ( .A(B[199]), .B(A[199]), .Z(n737) );
  AND U698 ( .A(B[199]), .B(A[199]), .Z(n738) );
  ANDN U699 ( .B(n749), .A(n741), .Z(n747) );
  NAND U700 ( .A(n750), .B(n736), .Z(n749) );
  XNOR U701 ( .A(n750), .B(n751), .Z(SUM[198]) );
  NANDN U702 ( .A(n741), .B(n736), .Z(n751) );
  OR U703 ( .A(A[198]), .B(B[198]), .Z(n736) );
  AND U704 ( .A(A[198]), .B(B[198]), .Z(n741) );
  NANDN U705 ( .A(n744), .B(n752), .Z(n750) );
  NAND U706 ( .A(n753), .B(n735), .Z(n752) );
  XNOR U707 ( .A(n753), .B(n754), .Z(SUM[197]) );
  NANDN U708 ( .A(n744), .B(n735), .Z(n754) );
  OR U709 ( .A(A[197]), .B(B[197]), .Z(n735) );
  AND U710 ( .A(A[197]), .B(B[197]), .Z(n744) );
  NANDN U711 ( .A(n746), .B(n755), .Z(n753) );
  NANDN U712 ( .A(n731), .B(n734), .Z(n755) );
  XOR U713 ( .A(n731), .B(n756), .Z(SUM[196]) );
  NANDN U714 ( .A(n746), .B(n734), .Z(n756) );
  OR U715 ( .A(A[196]), .B(B[196]), .Z(n734) );
  AND U716 ( .A(A[196]), .B(B[196]), .Z(n746) );
  NOR U717 ( .A(n690), .B(n691), .Z(n731) );
  AND U718 ( .A(n757), .B(n758), .Z(n691) );
  AND U719 ( .A(n759), .B(n760), .Z(n758) );
  NOR U720 ( .A(n761), .B(n762), .Z(n760) );
  AND U721 ( .A(n763), .B(n764), .Z(n757) );
  NANDN U722 ( .A(n765), .B(n766), .Z(n690) );
  NAND U723 ( .A(n767), .B(n764), .Z(n766) );
  NANDN U724 ( .A(n768), .B(n769), .Z(n767) );
  NAND U725 ( .A(n770), .B(n763), .Z(n769) );
  NANDN U726 ( .A(n771), .B(n772), .Z(n770) );
  NAND U727 ( .A(n759), .B(n773), .Z(n772) );
  XOR U728 ( .A(n774), .B(n775), .Z(SUM[195]) );
  NANDN U729 ( .A(n765), .B(n764), .Z(n775) );
  OR U730 ( .A(B[195]), .B(A[195]), .Z(n764) );
  AND U731 ( .A(B[195]), .B(A[195]), .Z(n765) );
  ANDN U732 ( .B(n776), .A(n768), .Z(n774) );
  NAND U733 ( .A(n777), .B(n763), .Z(n776) );
  XNOR U734 ( .A(n777), .B(n778), .Z(SUM[194]) );
  NANDN U735 ( .A(n768), .B(n763), .Z(n778) );
  OR U736 ( .A(A[194]), .B(B[194]), .Z(n763) );
  AND U737 ( .A(A[194]), .B(B[194]), .Z(n768) );
  NANDN U738 ( .A(n771), .B(n779), .Z(n777) );
  NAND U739 ( .A(n780), .B(n759), .Z(n779) );
  XNOR U740 ( .A(n780), .B(n781), .Z(SUM[193]) );
  NANDN U741 ( .A(n771), .B(n759), .Z(n781) );
  OR U742 ( .A(A[193]), .B(B[193]), .Z(n759) );
  AND U743 ( .A(A[193]), .B(B[193]), .Z(n771) );
  NANDN U744 ( .A(n773), .B(n782), .Z(n780) );
  OR U745 ( .A(n761), .B(n762), .Z(n782) );
  XOR U746 ( .A(n761), .B(n783), .Z(SUM[192]) );
  OR U747 ( .A(n762), .B(n773), .Z(n783) );
  AND U748 ( .A(A[192]), .B(B[192]), .Z(n773) );
  NOR U749 ( .A(B[192]), .B(A[192]), .Z(n762) );
  ANDN U750 ( .B(n784), .A(n785), .Z(n761) );
  NANDN U751 ( .A(n786), .B(n787), .Z(n784) );
  NANDN U752 ( .A(n788), .B(n789), .Z(n787) );
  NANDN U753 ( .A(n790), .B(n791), .Z(n789) );
  NANDN U754 ( .A(n792), .B(n793), .Z(n791) );
  NANDN U755 ( .A(n794), .B(n795), .Z(n793) );
  NAND U756 ( .A(n796), .B(n797), .Z(n795) );
  NAND U757 ( .A(n798), .B(n799), .Z(n797) );
  AND U758 ( .A(n800), .B(n801), .Z(n799) );
  ANDN U759 ( .B(n802), .A(n803), .Z(n801) );
  NOR U760 ( .A(n804), .B(n805), .Z(n798) );
  ANDN U761 ( .B(n806), .A(n807), .Z(n796) );
  NAND U762 ( .A(n808), .B(n802), .Z(n806) );
  NANDN U763 ( .A(n809), .B(n810), .Z(n808) );
  NANDN U764 ( .A(n805), .B(n811), .Z(n810) );
  NANDN U765 ( .A(n812), .B(n813), .Z(n811) );
  NAND U766 ( .A(n814), .B(n800), .Z(n813) );
  XOR U767 ( .A(n815), .B(n816), .Z(SUM[191]) );
  OR U768 ( .A(n786), .B(n785), .Z(n816) );
  AND U769 ( .A(B[191]), .B(A[191]), .Z(n785) );
  NOR U770 ( .A(B[191]), .B(A[191]), .Z(n786) );
  ANDN U771 ( .B(n817), .A(n788), .Z(n815) );
  NANDN U772 ( .A(n790), .B(n818), .Z(n817) );
  XNOR U773 ( .A(n818), .B(n819), .Z(SUM[190]) );
  OR U774 ( .A(n790), .B(n788), .Z(n819) );
  AND U775 ( .A(B[190]), .B(A[190]), .Z(n788) );
  NOR U776 ( .A(B[190]), .B(A[190]), .Z(n790) );
  NANDN U777 ( .A(n792), .B(n820), .Z(n818) );
  NANDN U778 ( .A(n794), .B(n821), .Z(n820) );
  XNOR U779 ( .A(n821), .B(n822), .Z(SUM[189]) );
  OR U780 ( .A(n794), .B(n792), .Z(n822) );
  AND U781 ( .A(B[189]), .B(A[189]), .Z(n792) );
  NOR U782 ( .A(B[189]), .B(A[189]), .Z(n794) );
  NANDN U783 ( .A(n807), .B(n823), .Z(n821) );
  NAND U784 ( .A(n824), .B(n802), .Z(n823) );
  XNOR U785 ( .A(n824), .B(n825), .Z(SUM[188]) );
  NANDN U786 ( .A(n807), .B(n802), .Z(n825) );
  OR U787 ( .A(A[188]), .B(B[188]), .Z(n802) );
  AND U788 ( .A(B[188]), .B(A[188]), .Z(n807) );
  NANDN U789 ( .A(n809), .B(n826), .Z(n824) );
  NANDN U790 ( .A(n805), .B(n827), .Z(n826) );
  NAND U791 ( .A(n828), .B(n829), .Z(n805) );
  AND U792 ( .A(n830), .B(n831), .Z(n829) );
  AND U793 ( .A(n832), .B(n833), .Z(n828) );
  NANDN U794 ( .A(n834), .B(n835), .Z(n809) );
  NAND U795 ( .A(n836), .B(n833), .Z(n835) );
  NANDN U796 ( .A(n837), .B(n838), .Z(n836) );
  NAND U797 ( .A(n839), .B(n832), .Z(n838) );
  NANDN U798 ( .A(n840), .B(n841), .Z(n839) );
  NAND U799 ( .A(n831), .B(n842), .Z(n841) );
  XOR U800 ( .A(n843), .B(n844), .Z(SUM[187]) );
  NANDN U801 ( .A(n834), .B(n833), .Z(n844) );
  OR U802 ( .A(B[187]), .B(A[187]), .Z(n833) );
  AND U803 ( .A(B[187]), .B(A[187]), .Z(n834) );
  ANDN U804 ( .B(n845), .A(n837), .Z(n843) );
  NAND U805 ( .A(n846), .B(n832), .Z(n845) );
  XNOR U806 ( .A(n846), .B(n847), .Z(SUM[186]) );
  NANDN U807 ( .A(n837), .B(n832), .Z(n847) );
  OR U808 ( .A(B[186]), .B(A[186]), .Z(n832) );
  AND U809 ( .A(B[186]), .B(A[186]), .Z(n837) );
  NANDN U810 ( .A(n840), .B(n848), .Z(n846) );
  NAND U811 ( .A(n849), .B(n831), .Z(n848) );
  XNOR U812 ( .A(n849), .B(n850), .Z(SUM[185]) );
  NANDN U813 ( .A(n840), .B(n831), .Z(n850) );
  OR U814 ( .A(B[185]), .B(A[185]), .Z(n831) );
  AND U815 ( .A(B[185]), .B(A[185]), .Z(n840) );
  NANDN U816 ( .A(n842), .B(n851), .Z(n849) );
  NAND U817 ( .A(n827), .B(n830), .Z(n851) );
  XNOR U818 ( .A(n827), .B(n852), .Z(SUM[184]) );
  NANDN U819 ( .A(n842), .B(n830), .Z(n852) );
  OR U820 ( .A(B[184]), .B(A[184]), .Z(n830) );
  AND U821 ( .A(B[184]), .B(A[184]), .Z(n842) );
  NANDN U822 ( .A(n812), .B(n853), .Z(n827) );
  NANDN U823 ( .A(n854), .B(n800), .Z(n853) );
  AND U824 ( .A(n855), .B(n856), .Z(n800) );
  AND U825 ( .A(n857), .B(n858), .Z(n856) );
  AND U826 ( .A(n859), .B(n860), .Z(n855) );
  NANDN U827 ( .A(n861), .B(n862), .Z(n812) );
  NAND U828 ( .A(n863), .B(n860), .Z(n862) );
  NANDN U829 ( .A(n864), .B(n865), .Z(n863) );
  NAND U830 ( .A(n866), .B(n859), .Z(n865) );
  NANDN U831 ( .A(n867), .B(n868), .Z(n866) );
  NAND U832 ( .A(n858), .B(n869), .Z(n868) );
  XOR U833 ( .A(n870), .B(n871), .Z(SUM[183]) );
  NANDN U834 ( .A(n861), .B(n860), .Z(n871) );
  OR U835 ( .A(B[183]), .B(A[183]), .Z(n860) );
  AND U836 ( .A(B[183]), .B(A[183]), .Z(n861) );
  ANDN U837 ( .B(n872), .A(n864), .Z(n870) );
  NAND U838 ( .A(n873), .B(n859), .Z(n872) );
  XNOR U839 ( .A(n873), .B(n874), .Z(SUM[182]) );
  NANDN U840 ( .A(n864), .B(n859), .Z(n874) );
  OR U841 ( .A(B[182]), .B(A[182]), .Z(n859) );
  AND U842 ( .A(B[182]), .B(A[182]), .Z(n864) );
  NANDN U843 ( .A(n867), .B(n875), .Z(n873) );
  NAND U844 ( .A(n876), .B(n858), .Z(n875) );
  XNOR U845 ( .A(n876), .B(n877), .Z(SUM[181]) );
  NANDN U846 ( .A(n867), .B(n858), .Z(n877) );
  OR U847 ( .A(B[181]), .B(A[181]), .Z(n858) );
  AND U848 ( .A(B[181]), .B(A[181]), .Z(n867) );
  NANDN U849 ( .A(n869), .B(n878), .Z(n876) );
  NANDN U850 ( .A(n854), .B(n857), .Z(n878) );
  XOR U851 ( .A(n854), .B(n879), .Z(SUM[180]) );
  NANDN U852 ( .A(n869), .B(n857), .Z(n879) );
  OR U853 ( .A(B[180]), .B(A[180]), .Z(n857) );
  AND U854 ( .A(B[180]), .B(A[180]), .Z(n869) );
  ANDN U855 ( .B(n880), .A(n814), .Z(n854) );
  NANDN U856 ( .A(n881), .B(n882), .Z(n814) );
  NAND U857 ( .A(n883), .B(n884), .Z(n882) );
  NANDN U858 ( .A(n885), .B(n886), .Z(n883) );
  NANDN U859 ( .A(n887), .B(n888), .Z(n886) );
  NANDN U860 ( .A(n889), .B(n890), .Z(n888) );
  NAND U861 ( .A(n891), .B(n892), .Z(n890) );
  OR U862 ( .A(n804), .B(n803), .Z(n880) );
  NAND U863 ( .A(n893), .B(n894), .Z(n804) );
  AND U864 ( .A(n895), .B(n891), .Z(n894) );
  ANDN U865 ( .B(n884), .A(n887), .Z(n893) );
  XOR U866 ( .A(n896), .B(n897), .Z(SUM[179]) );
  NANDN U867 ( .A(n881), .B(n884), .Z(n897) );
  OR U868 ( .A(B[179]), .B(A[179]), .Z(n884) );
  AND U869 ( .A(B[179]), .B(A[179]), .Z(n881) );
  ANDN U870 ( .B(n898), .A(n885), .Z(n896) );
  NANDN U871 ( .A(n887), .B(n899), .Z(n898) );
  XNOR U872 ( .A(n899), .B(n900), .Z(SUM[178]) );
  OR U873 ( .A(n887), .B(n885), .Z(n900) );
  AND U874 ( .A(B[178]), .B(A[178]), .Z(n885) );
  NOR U875 ( .A(B[178]), .B(A[178]), .Z(n887) );
  NANDN U876 ( .A(n889), .B(n901), .Z(n899) );
  NAND U877 ( .A(n902), .B(n891), .Z(n901) );
  XNOR U878 ( .A(n902), .B(n903), .Z(SUM[177]) );
  NANDN U879 ( .A(n889), .B(n891), .Z(n903) );
  OR U880 ( .A(B[177]), .B(A[177]), .Z(n891) );
  AND U881 ( .A(B[177]), .B(A[177]), .Z(n889) );
  NANDN U882 ( .A(n892), .B(n904), .Z(n902) );
  NANDN U883 ( .A(n803), .B(n895), .Z(n904) );
  XOR U884 ( .A(n803), .B(n905), .Z(SUM[176]) );
  NANDN U885 ( .A(n892), .B(n895), .Z(n905) );
  OR U886 ( .A(B[176]), .B(A[176]), .Z(n895) );
  AND U887 ( .A(A[176]), .B(B[176]), .Z(n892) );
  ANDN U888 ( .B(n906), .A(n907), .Z(n803) );
  NANDN U889 ( .A(n908), .B(n909), .Z(n906) );
  NANDN U890 ( .A(n910), .B(n911), .Z(n909) );
  NANDN U891 ( .A(n912), .B(n913), .Z(n911) );
  NANDN U892 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U893 ( .A(n916), .B(n917), .Z(n915) );
  NAND U894 ( .A(n918), .B(n919), .Z(n917) );
  NAND U895 ( .A(n920), .B(n921), .Z(n919) );
  AND U896 ( .A(n922), .B(n923), .Z(n921) );
  ANDN U897 ( .B(n924), .A(n925), .Z(n923) );
  NOR U898 ( .A(n926), .B(n927), .Z(n920) );
  ANDN U899 ( .B(n928), .A(n929), .Z(n918) );
  NAND U900 ( .A(n930), .B(n924), .Z(n928) );
  NANDN U901 ( .A(n931), .B(n932), .Z(n930) );
  NANDN U902 ( .A(n927), .B(n933), .Z(n932) );
  NANDN U903 ( .A(n934), .B(n935), .Z(n933) );
  NAND U904 ( .A(n936), .B(n922), .Z(n935) );
  XOR U905 ( .A(n937), .B(n938), .Z(SUM[175]) );
  OR U906 ( .A(n908), .B(n907), .Z(n938) );
  AND U907 ( .A(B[175]), .B(A[175]), .Z(n907) );
  NOR U908 ( .A(B[175]), .B(A[175]), .Z(n908) );
  ANDN U909 ( .B(n939), .A(n910), .Z(n937) );
  NANDN U910 ( .A(n912), .B(n940), .Z(n939) );
  XNOR U911 ( .A(n940), .B(n941), .Z(SUM[174]) );
  OR U912 ( .A(n912), .B(n910), .Z(n941) );
  AND U913 ( .A(B[174]), .B(A[174]), .Z(n910) );
  NOR U914 ( .A(B[174]), .B(A[174]), .Z(n912) );
  NANDN U915 ( .A(n914), .B(n942), .Z(n940) );
  NANDN U916 ( .A(n916), .B(n943), .Z(n942) );
  XNOR U917 ( .A(n943), .B(n944), .Z(SUM[173]) );
  OR U918 ( .A(n916), .B(n914), .Z(n944) );
  AND U919 ( .A(B[173]), .B(A[173]), .Z(n914) );
  NOR U920 ( .A(B[173]), .B(A[173]), .Z(n916) );
  NANDN U921 ( .A(n929), .B(n945), .Z(n943) );
  NAND U922 ( .A(n946), .B(n924), .Z(n945) );
  XNOR U923 ( .A(n946), .B(n947), .Z(SUM[172]) );
  NANDN U924 ( .A(n929), .B(n924), .Z(n947) );
  OR U925 ( .A(A[172]), .B(B[172]), .Z(n924) );
  AND U926 ( .A(B[172]), .B(A[172]), .Z(n929) );
  NANDN U927 ( .A(n931), .B(n948), .Z(n946) );
  NANDN U928 ( .A(n927), .B(n949), .Z(n948) );
  NAND U929 ( .A(n950), .B(n951), .Z(n927) );
  AND U930 ( .A(n952), .B(n953), .Z(n951) );
  AND U931 ( .A(n954), .B(n955), .Z(n950) );
  NANDN U932 ( .A(n956), .B(n957), .Z(n931) );
  NAND U933 ( .A(n958), .B(n955), .Z(n957) );
  NANDN U934 ( .A(n959), .B(n960), .Z(n958) );
  NAND U935 ( .A(n961), .B(n954), .Z(n960) );
  NANDN U936 ( .A(n962), .B(n963), .Z(n961) );
  NAND U937 ( .A(n953), .B(n964), .Z(n963) );
  XOR U938 ( .A(n965), .B(n966), .Z(SUM[171]) );
  NANDN U939 ( .A(n956), .B(n955), .Z(n966) );
  OR U940 ( .A(B[171]), .B(A[171]), .Z(n955) );
  AND U941 ( .A(B[171]), .B(A[171]), .Z(n956) );
  ANDN U942 ( .B(n967), .A(n959), .Z(n965) );
  NAND U943 ( .A(n968), .B(n954), .Z(n967) );
  XNOR U944 ( .A(n968), .B(n969), .Z(SUM[170]) );
  NANDN U945 ( .A(n959), .B(n954), .Z(n969) );
  OR U946 ( .A(B[170]), .B(A[170]), .Z(n954) );
  AND U947 ( .A(B[170]), .B(A[170]), .Z(n959) );
  NANDN U948 ( .A(n962), .B(n970), .Z(n968) );
  NAND U949 ( .A(n971), .B(n953), .Z(n970) );
  XNOR U950 ( .A(n971), .B(n972), .Z(SUM[169]) );
  NANDN U951 ( .A(n962), .B(n953), .Z(n972) );
  OR U952 ( .A(B[169]), .B(A[169]), .Z(n953) );
  AND U953 ( .A(B[169]), .B(A[169]), .Z(n962) );
  NANDN U954 ( .A(n964), .B(n973), .Z(n971) );
  NAND U955 ( .A(n949), .B(n952), .Z(n973) );
  XNOR U956 ( .A(n949), .B(n974), .Z(SUM[168]) );
  NANDN U957 ( .A(n964), .B(n952), .Z(n974) );
  OR U958 ( .A(B[168]), .B(A[168]), .Z(n952) );
  AND U959 ( .A(B[168]), .B(A[168]), .Z(n964) );
  NANDN U960 ( .A(n934), .B(n975), .Z(n949) );
  NANDN U961 ( .A(n976), .B(n922), .Z(n975) );
  AND U962 ( .A(n977), .B(n978), .Z(n922) );
  AND U963 ( .A(n979), .B(n980), .Z(n978) );
  AND U964 ( .A(n981), .B(n982), .Z(n977) );
  NANDN U965 ( .A(n983), .B(n984), .Z(n934) );
  NAND U966 ( .A(n985), .B(n982), .Z(n984) );
  NANDN U967 ( .A(n986), .B(n987), .Z(n985) );
  NAND U968 ( .A(n988), .B(n981), .Z(n987) );
  NANDN U969 ( .A(n989), .B(n990), .Z(n988) );
  NAND U970 ( .A(n980), .B(n991), .Z(n990) );
  XOR U971 ( .A(n992), .B(n993), .Z(SUM[167]) );
  NANDN U972 ( .A(n983), .B(n982), .Z(n993) );
  OR U973 ( .A(B[167]), .B(A[167]), .Z(n982) );
  AND U974 ( .A(B[167]), .B(A[167]), .Z(n983) );
  ANDN U975 ( .B(n994), .A(n986), .Z(n992) );
  NAND U976 ( .A(n995), .B(n981), .Z(n994) );
  XNOR U977 ( .A(n995), .B(n996), .Z(SUM[166]) );
  NANDN U978 ( .A(n986), .B(n981), .Z(n996) );
  OR U979 ( .A(B[166]), .B(A[166]), .Z(n981) );
  AND U980 ( .A(B[166]), .B(A[166]), .Z(n986) );
  NANDN U981 ( .A(n989), .B(n997), .Z(n995) );
  NAND U982 ( .A(n998), .B(n980), .Z(n997) );
  XNOR U983 ( .A(n998), .B(n999), .Z(SUM[165]) );
  NANDN U984 ( .A(n989), .B(n980), .Z(n999) );
  OR U985 ( .A(B[165]), .B(A[165]), .Z(n980) );
  AND U986 ( .A(B[165]), .B(A[165]), .Z(n989) );
  NANDN U987 ( .A(n991), .B(n1000), .Z(n998) );
  NANDN U988 ( .A(n976), .B(n979), .Z(n1000) );
  XOR U989 ( .A(n976), .B(n1001), .Z(SUM[164]) );
  NANDN U990 ( .A(n991), .B(n979), .Z(n1001) );
  OR U991 ( .A(B[164]), .B(A[164]), .Z(n979) );
  AND U992 ( .A(B[164]), .B(A[164]), .Z(n991) );
  ANDN U993 ( .B(n1002), .A(n936), .Z(n976) );
  NANDN U994 ( .A(n1003), .B(n1004), .Z(n936) );
  NAND U995 ( .A(n1005), .B(n1006), .Z(n1004) );
  NANDN U996 ( .A(n1007), .B(n1008), .Z(n1005) );
  NANDN U997 ( .A(n1009), .B(n1010), .Z(n1008) );
  NANDN U998 ( .A(n1011), .B(n1012), .Z(n1010) );
  NAND U999 ( .A(n1013), .B(n1014), .Z(n1012) );
  OR U1000 ( .A(n926), .B(n925), .Z(n1002) );
  NAND U1001 ( .A(n1015), .B(n1016), .Z(n926) );
  AND U1002 ( .A(n1017), .B(n1013), .Z(n1016) );
  ANDN U1003 ( .B(n1006), .A(n1009), .Z(n1015) );
  XOR U1004 ( .A(n1018), .B(n1019), .Z(SUM[163]) );
  NANDN U1005 ( .A(n1003), .B(n1006), .Z(n1019) );
  OR U1006 ( .A(B[163]), .B(A[163]), .Z(n1006) );
  AND U1007 ( .A(B[163]), .B(A[163]), .Z(n1003) );
  ANDN U1008 ( .B(n1020), .A(n1007), .Z(n1018) );
  NANDN U1009 ( .A(n1009), .B(n1021), .Z(n1020) );
  XNOR U1010 ( .A(n1021), .B(n1022), .Z(SUM[162]) );
  OR U1011 ( .A(n1009), .B(n1007), .Z(n1022) );
  AND U1012 ( .A(B[162]), .B(A[162]), .Z(n1007) );
  NOR U1013 ( .A(B[162]), .B(A[162]), .Z(n1009) );
  NANDN U1014 ( .A(n1011), .B(n1023), .Z(n1021) );
  NAND U1015 ( .A(n1024), .B(n1013), .Z(n1023) );
  XNOR U1016 ( .A(n1024), .B(n1025), .Z(SUM[161]) );
  NANDN U1017 ( .A(n1011), .B(n1013), .Z(n1025) );
  OR U1018 ( .A(B[161]), .B(A[161]), .Z(n1013) );
  AND U1019 ( .A(B[161]), .B(A[161]), .Z(n1011) );
  NANDN U1020 ( .A(n1014), .B(n1026), .Z(n1024) );
  NANDN U1021 ( .A(n925), .B(n1017), .Z(n1026) );
  XOR U1022 ( .A(n925), .B(n1027), .Z(SUM[160]) );
  NANDN U1023 ( .A(n1014), .B(n1017), .Z(n1027) );
  OR U1024 ( .A(B[160]), .B(A[160]), .Z(n1017) );
  AND U1025 ( .A(A[160]), .B(B[160]), .Z(n1014) );
  ANDN U1026 ( .B(n1028), .A(n1029), .Z(n925) );
  NANDN U1027 ( .A(n1030), .B(n1031), .Z(n1028) );
  NANDN U1028 ( .A(n1032), .B(n1033), .Z(n1031) );
  NANDN U1029 ( .A(n1034), .B(n1035), .Z(n1033) );
  NANDN U1030 ( .A(n1036), .B(n1037), .Z(n1035) );
  NANDN U1031 ( .A(n1038), .B(n1039), .Z(n1037) );
  NAND U1032 ( .A(n1040), .B(n1041), .Z(n1039) );
  NAND U1033 ( .A(n1042), .B(n1043), .Z(n1041) );
  AND U1034 ( .A(n1044), .B(n1045), .Z(n1043) );
  ANDN U1035 ( .B(n1046), .A(n1047), .Z(n1045) );
  NOR U1036 ( .A(n1048), .B(n1049), .Z(n1042) );
  ANDN U1037 ( .B(n1050), .A(n1051), .Z(n1040) );
  NAND U1038 ( .A(n1052), .B(n1046), .Z(n1050) );
  NANDN U1039 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U1040 ( .A(n1049), .B(n1055), .Z(n1054) );
  NANDN U1041 ( .A(n1056), .B(n1057), .Z(n1055) );
  NAND U1042 ( .A(n1058), .B(n1044), .Z(n1057) );
  XOR U1043 ( .A(n1059), .B(n1060), .Z(SUM[159]) );
  OR U1044 ( .A(n1030), .B(n1029), .Z(n1060) );
  AND U1045 ( .A(B[159]), .B(A[159]), .Z(n1029) );
  NOR U1046 ( .A(B[159]), .B(A[159]), .Z(n1030) );
  ANDN U1047 ( .B(n1061), .A(n1032), .Z(n1059) );
  NANDN U1048 ( .A(n1034), .B(n1062), .Z(n1061) );
  XNOR U1049 ( .A(n1062), .B(n1063), .Z(SUM[158]) );
  OR U1050 ( .A(n1034), .B(n1032), .Z(n1063) );
  AND U1051 ( .A(B[158]), .B(A[158]), .Z(n1032) );
  NOR U1052 ( .A(B[158]), .B(A[158]), .Z(n1034) );
  NANDN U1053 ( .A(n1036), .B(n1064), .Z(n1062) );
  NANDN U1054 ( .A(n1038), .B(n1065), .Z(n1064) );
  XNOR U1055 ( .A(n1065), .B(n1066), .Z(SUM[157]) );
  OR U1056 ( .A(n1038), .B(n1036), .Z(n1066) );
  AND U1057 ( .A(B[157]), .B(A[157]), .Z(n1036) );
  NOR U1058 ( .A(B[157]), .B(A[157]), .Z(n1038) );
  NANDN U1059 ( .A(n1051), .B(n1067), .Z(n1065) );
  NAND U1060 ( .A(n1068), .B(n1046), .Z(n1067) );
  XNOR U1061 ( .A(n1068), .B(n1069), .Z(SUM[156]) );
  NANDN U1062 ( .A(n1051), .B(n1046), .Z(n1069) );
  OR U1063 ( .A(A[156]), .B(B[156]), .Z(n1046) );
  AND U1064 ( .A(B[156]), .B(A[156]), .Z(n1051) );
  NANDN U1065 ( .A(n1053), .B(n1070), .Z(n1068) );
  NANDN U1066 ( .A(n1049), .B(n1071), .Z(n1070) );
  NAND U1067 ( .A(n1072), .B(n1073), .Z(n1049) );
  AND U1068 ( .A(n1074), .B(n1075), .Z(n1073) );
  AND U1069 ( .A(n1076), .B(n1077), .Z(n1072) );
  NANDN U1070 ( .A(n1078), .B(n1079), .Z(n1053) );
  NAND U1071 ( .A(n1080), .B(n1077), .Z(n1079) );
  NANDN U1072 ( .A(n1081), .B(n1082), .Z(n1080) );
  NAND U1073 ( .A(n1083), .B(n1076), .Z(n1082) );
  NANDN U1074 ( .A(n1084), .B(n1085), .Z(n1083) );
  NAND U1075 ( .A(n1075), .B(n1086), .Z(n1085) );
  XOR U1076 ( .A(n1087), .B(n1088), .Z(SUM[155]) );
  NANDN U1077 ( .A(n1078), .B(n1077), .Z(n1088) );
  OR U1078 ( .A(B[155]), .B(A[155]), .Z(n1077) );
  AND U1079 ( .A(B[155]), .B(A[155]), .Z(n1078) );
  ANDN U1080 ( .B(n1089), .A(n1081), .Z(n1087) );
  NAND U1081 ( .A(n1090), .B(n1076), .Z(n1089) );
  XNOR U1082 ( .A(n1090), .B(n1091), .Z(SUM[154]) );
  NANDN U1083 ( .A(n1081), .B(n1076), .Z(n1091) );
  OR U1084 ( .A(B[154]), .B(A[154]), .Z(n1076) );
  AND U1085 ( .A(B[154]), .B(A[154]), .Z(n1081) );
  NANDN U1086 ( .A(n1084), .B(n1092), .Z(n1090) );
  NAND U1087 ( .A(n1093), .B(n1075), .Z(n1092) );
  XNOR U1088 ( .A(n1093), .B(n1094), .Z(SUM[153]) );
  NANDN U1089 ( .A(n1084), .B(n1075), .Z(n1094) );
  OR U1090 ( .A(B[153]), .B(A[153]), .Z(n1075) );
  AND U1091 ( .A(B[153]), .B(A[153]), .Z(n1084) );
  NANDN U1092 ( .A(n1086), .B(n1095), .Z(n1093) );
  NAND U1093 ( .A(n1071), .B(n1074), .Z(n1095) );
  XNOR U1094 ( .A(n1071), .B(n1096), .Z(SUM[152]) );
  NANDN U1095 ( .A(n1086), .B(n1074), .Z(n1096) );
  OR U1096 ( .A(B[152]), .B(A[152]), .Z(n1074) );
  AND U1097 ( .A(B[152]), .B(A[152]), .Z(n1086) );
  NANDN U1098 ( .A(n1056), .B(n1097), .Z(n1071) );
  NANDN U1099 ( .A(n1098), .B(n1044), .Z(n1097) );
  AND U1100 ( .A(n1099), .B(n1100), .Z(n1044) );
  AND U1101 ( .A(n1101), .B(n1102), .Z(n1100) );
  AND U1102 ( .A(n1103), .B(n1104), .Z(n1099) );
  NANDN U1103 ( .A(n1105), .B(n1106), .Z(n1056) );
  NAND U1104 ( .A(n1107), .B(n1104), .Z(n1106) );
  NANDN U1105 ( .A(n1108), .B(n1109), .Z(n1107) );
  NAND U1106 ( .A(n1110), .B(n1103), .Z(n1109) );
  NANDN U1107 ( .A(n1111), .B(n1112), .Z(n1110) );
  NAND U1108 ( .A(n1102), .B(n1113), .Z(n1112) );
  XOR U1109 ( .A(n1114), .B(n1115), .Z(SUM[151]) );
  NANDN U1110 ( .A(n1105), .B(n1104), .Z(n1115) );
  OR U1111 ( .A(B[151]), .B(A[151]), .Z(n1104) );
  AND U1112 ( .A(B[151]), .B(A[151]), .Z(n1105) );
  ANDN U1113 ( .B(n1116), .A(n1108), .Z(n1114) );
  NAND U1114 ( .A(n1117), .B(n1103), .Z(n1116) );
  XNOR U1115 ( .A(n1117), .B(n1118), .Z(SUM[150]) );
  NANDN U1116 ( .A(n1108), .B(n1103), .Z(n1118) );
  OR U1117 ( .A(B[150]), .B(A[150]), .Z(n1103) );
  AND U1118 ( .A(B[150]), .B(A[150]), .Z(n1108) );
  NANDN U1119 ( .A(n1111), .B(n1119), .Z(n1117) );
  NAND U1120 ( .A(n1120), .B(n1102), .Z(n1119) );
  XNOR U1121 ( .A(n1120), .B(n1121), .Z(SUM[149]) );
  NANDN U1122 ( .A(n1111), .B(n1102), .Z(n1121) );
  OR U1123 ( .A(B[149]), .B(A[149]), .Z(n1102) );
  AND U1124 ( .A(B[149]), .B(A[149]), .Z(n1111) );
  NANDN U1125 ( .A(n1113), .B(n1122), .Z(n1120) );
  NANDN U1126 ( .A(n1098), .B(n1101), .Z(n1122) );
  XOR U1127 ( .A(n1098), .B(n1123), .Z(SUM[148]) );
  NANDN U1128 ( .A(n1113), .B(n1101), .Z(n1123) );
  OR U1129 ( .A(B[148]), .B(A[148]), .Z(n1101) );
  AND U1130 ( .A(B[148]), .B(A[148]), .Z(n1113) );
  ANDN U1131 ( .B(n1124), .A(n1058), .Z(n1098) );
  NANDN U1132 ( .A(n1125), .B(n1126), .Z(n1058) );
  NAND U1133 ( .A(n1127), .B(n1128), .Z(n1126) );
  NANDN U1134 ( .A(n1129), .B(n1130), .Z(n1127) );
  NANDN U1135 ( .A(n1131), .B(n1132), .Z(n1130) );
  NANDN U1136 ( .A(n1133), .B(n1134), .Z(n1132) );
  NAND U1137 ( .A(n1135), .B(n1136), .Z(n1134) );
  OR U1138 ( .A(n1048), .B(n1047), .Z(n1124) );
  NAND U1139 ( .A(n1137), .B(n1138), .Z(n1048) );
  AND U1140 ( .A(n1139), .B(n1135), .Z(n1138) );
  ANDN U1141 ( .B(n1128), .A(n1131), .Z(n1137) );
  XOR U1142 ( .A(n1140), .B(n1141), .Z(SUM[147]) );
  NANDN U1143 ( .A(n1125), .B(n1128), .Z(n1141) );
  OR U1144 ( .A(B[147]), .B(A[147]), .Z(n1128) );
  AND U1145 ( .A(B[147]), .B(A[147]), .Z(n1125) );
  ANDN U1146 ( .B(n1142), .A(n1129), .Z(n1140) );
  NANDN U1147 ( .A(n1131), .B(n1143), .Z(n1142) );
  XNOR U1148 ( .A(n1143), .B(n1144), .Z(SUM[146]) );
  OR U1149 ( .A(n1131), .B(n1129), .Z(n1144) );
  AND U1150 ( .A(B[146]), .B(A[146]), .Z(n1129) );
  NOR U1151 ( .A(B[146]), .B(A[146]), .Z(n1131) );
  NANDN U1152 ( .A(n1133), .B(n1145), .Z(n1143) );
  NAND U1153 ( .A(n1146), .B(n1135), .Z(n1145) );
  XNOR U1154 ( .A(n1146), .B(n1147), .Z(SUM[145]) );
  NANDN U1155 ( .A(n1133), .B(n1135), .Z(n1147) );
  OR U1156 ( .A(B[145]), .B(A[145]), .Z(n1135) );
  AND U1157 ( .A(B[145]), .B(A[145]), .Z(n1133) );
  NANDN U1158 ( .A(n1136), .B(n1148), .Z(n1146) );
  NANDN U1159 ( .A(n1047), .B(n1139), .Z(n1148) );
  XOR U1160 ( .A(n1047), .B(n1149), .Z(SUM[144]) );
  NANDN U1161 ( .A(n1136), .B(n1139), .Z(n1149) );
  OR U1162 ( .A(B[144]), .B(A[144]), .Z(n1139) );
  AND U1163 ( .A(A[144]), .B(B[144]), .Z(n1136) );
  ANDN U1164 ( .B(n1150), .A(n1151), .Z(n1047) );
  NANDN U1165 ( .A(n1152), .B(n1153), .Z(n1150) );
  NANDN U1166 ( .A(n1154), .B(n1155), .Z(n1153) );
  NANDN U1167 ( .A(n1156), .B(n1157), .Z(n1155) );
  NANDN U1168 ( .A(n1158), .B(n1159), .Z(n1157) );
  NANDN U1169 ( .A(n1160), .B(n1161), .Z(n1159) );
  NAND U1170 ( .A(n1162), .B(n1163), .Z(n1161) );
  NAND U1171 ( .A(n1164), .B(n1165), .Z(n1163) );
  AND U1172 ( .A(n1166), .B(n1167), .Z(n1165) );
  ANDN U1173 ( .B(n1168), .A(n1169), .Z(n1167) );
  NOR U1174 ( .A(n1170), .B(n1171), .Z(n1164) );
  ANDN U1175 ( .B(n1172), .A(n1173), .Z(n1162) );
  NAND U1176 ( .A(n1174), .B(n1168), .Z(n1172) );
  NANDN U1177 ( .A(n1175), .B(n1176), .Z(n1174) );
  NANDN U1178 ( .A(n1171), .B(n1177), .Z(n1176) );
  NANDN U1179 ( .A(n1178), .B(n1179), .Z(n1177) );
  NAND U1180 ( .A(n1180), .B(n1166), .Z(n1179) );
  XOR U1181 ( .A(n1181), .B(n1182), .Z(SUM[143]) );
  OR U1182 ( .A(n1152), .B(n1151), .Z(n1182) );
  AND U1183 ( .A(B[143]), .B(A[143]), .Z(n1151) );
  NOR U1184 ( .A(B[143]), .B(A[143]), .Z(n1152) );
  ANDN U1185 ( .B(n1183), .A(n1154), .Z(n1181) );
  NANDN U1186 ( .A(n1156), .B(n1184), .Z(n1183) );
  XNOR U1187 ( .A(n1184), .B(n1185), .Z(SUM[142]) );
  OR U1188 ( .A(n1156), .B(n1154), .Z(n1185) );
  AND U1189 ( .A(B[142]), .B(A[142]), .Z(n1154) );
  NOR U1190 ( .A(B[142]), .B(A[142]), .Z(n1156) );
  NANDN U1191 ( .A(n1158), .B(n1186), .Z(n1184) );
  NANDN U1192 ( .A(n1160), .B(n1187), .Z(n1186) );
  XNOR U1193 ( .A(n1187), .B(n1188), .Z(SUM[141]) );
  OR U1194 ( .A(n1160), .B(n1158), .Z(n1188) );
  AND U1195 ( .A(B[141]), .B(A[141]), .Z(n1158) );
  NOR U1196 ( .A(B[141]), .B(A[141]), .Z(n1160) );
  NANDN U1197 ( .A(n1173), .B(n1189), .Z(n1187) );
  NAND U1198 ( .A(n1190), .B(n1168), .Z(n1189) );
  XNOR U1199 ( .A(n1190), .B(n1191), .Z(SUM[140]) );
  NANDN U1200 ( .A(n1173), .B(n1168), .Z(n1191) );
  OR U1201 ( .A(A[140]), .B(B[140]), .Z(n1168) );
  AND U1202 ( .A(B[140]), .B(A[140]), .Z(n1173) );
  NANDN U1203 ( .A(n1175), .B(n1192), .Z(n1190) );
  NANDN U1204 ( .A(n1171), .B(n1193), .Z(n1192) );
  NAND U1205 ( .A(n1194), .B(n1195), .Z(n1171) );
  AND U1206 ( .A(n1196), .B(n1197), .Z(n1195) );
  AND U1207 ( .A(n1198), .B(n1199), .Z(n1194) );
  NANDN U1208 ( .A(n1200), .B(n1201), .Z(n1175) );
  NAND U1209 ( .A(n1202), .B(n1199), .Z(n1201) );
  NANDN U1210 ( .A(n1203), .B(n1204), .Z(n1202) );
  NAND U1211 ( .A(n1205), .B(n1198), .Z(n1204) );
  NANDN U1212 ( .A(n1206), .B(n1207), .Z(n1205) );
  NAND U1213 ( .A(n1197), .B(n1208), .Z(n1207) );
  XOR U1214 ( .A(n1209), .B(n1210), .Z(SUM[139]) );
  NANDN U1215 ( .A(n1200), .B(n1199), .Z(n1210) );
  OR U1216 ( .A(B[139]), .B(A[139]), .Z(n1199) );
  AND U1217 ( .A(B[139]), .B(A[139]), .Z(n1200) );
  ANDN U1218 ( .B(n1211), .A(n1203), .Z(n1209) );
  NAND U1219 ( .A(n1212), .B(n1198), .Z(n1211) );
  XNOR U1220 ( .A(n1212), .B(n1213), .Z(SUM[138]) );
  NANDN U1221 ( .A(n1203), .B(n1198), .Z(n1213) );
  OR U1222 ( .A(B[138]), .B(A[138]), .Z(n1198) );
  AND U1223 ( .A(B[138]), .B(A[138]), .Z(n1203) );
  NANDN U1224 ( .A(n1206), .B(n1214), .Z(n1212) );
  NAND U1225 ( .A(n1215), .B(n1197), .Z(n1214) );
  XNOR U1226 ( .A(n1215), .B(n1216), .Z(SUM[137]) );
  NANDN U1227 ( .A(n1206), .B(n1197), .Z(n1216) );
  OR U1228 ( .A(B[137]), .B(A[137]), .Z(n1197) );
  AND U1229 ( .A(B[137]), .B(A[137]), .Z(n1206) );
  NANDN U1230 ( .A(n1208), .B(n1217), .Z(n1215) );
  NAND U1231 ( .A(n1193), .B(n1196), .Z(n1217) );
  XNOR U1232 ( .A(n1193), .B(n1218), .Z(SUM[136]) );
  NANDN U1233 ( .A(n1208), .B(n1196), .Z(n1218) );
  OR U1234 ( .A(B[136]), .B(A[136]), .Z(n1196) );
  AND U1235 ( .A(B[136]), .B(A[136]), .Z(n1208) );
  NANDN U1236 ( .A(n1178), .B(n1219), .Z(n1193) );
  NANDN U1237 ( .A(n1220), .B(n1166), .Z(n1219) );
  AND U1238 ( .A(n1221), .B(n1222), .Z(n1166) );
  AND U1239 ( .A(n1223), .B(n1224), .Z(n1222) );
  AND U1240 ( .A(n1225), .B(n1226), .Z(n1221) );
  NANDN U1241 ( .A(n1227), .B(n1228), .Z(n1178) );
  NAND U1242 ( .A(n1229), .B(n1226), .Z(n1228) );
  NANDN U1243 ( .A(n1230), .B(n1231), .Z(n1229) );
  NAND U1244 ( .A(n1232), .B(n1225), .Z(n1231) );
  NANDN U1245 ( .A(n1233), .B(n1234), .Z(n1232) );
  NAND U1246 ( .A(n1224), .B(n1235), .Z(n1234) );
  XOR U1247 ( .A(n1236), .B(n1237), .Z(SUM[135]) );
  NANDN U1248 ( .A(n1227), .B(n1226), .Z(n1237) );
  OR U1249 ( .A(B[135]), .B(A[135]), .Z(n1226) );
  AND U1250 ( .A(B[135]), .B(A[135]), .Z(n1227) );
  ANDN U1251 ( .B(n1238), .A(n1230), .Z(n1236) );
  NAND U1252 ( .A(n1239), .B(n1225), .Z(n1238) );
  XNOR U1253 ( .A(n1239), .B(n1240), .Z(SUM[134]) );
  NANDN U1254 ( .A(n1230), .B(n1225), .Z(n1240) );
  OR U1255 ( .A(B[134]), .B(A[134]), .Z(n1225) );
  AND U1256 ( .A(B[134]), .B(A[134]), .Z(n1230) );
  NANDN U1257 ( .A(n1233), .B(n1241), .Z(n1239) );
  NAND U1258 ( .A(n1242), .B(n1224), .Z(n1241) );
  XNOR U1259 ( .A(n1242), .B(n1243), .Z(SUM[133]) );
  NANDN U1260 ( .A(n1233), .B(n1224), .Z(n1243) );
  OR U1261 ( .A(B[133]), .B(A[133]), .Z(n1224) );
  AND U1262 ( .A(B[133]), .B(A[133]), .Z(n1233) );
  NANDN U1263 ( .A(n1235), .B(n1244), .Z(n1242) );
  NANDN U1264 ( .A(n1220), .B(n1223), .Z(n1244) );
  XOR U1265 ( .A(n1220), .B(n1245), .Z(SUM[132]) );
  NANDN U1266 ( .A(n1235), .B(n1223), .Z(n1245) );
  OR U1267 ( .A(B[132]), .B(A[132]), .Z(n1223) );
  AND U1268 ( .A(B[132]), .B(A[132]), .Z(n1235) );
  ANDN U1269 ( .B(n1246), .A(n1180), .Z(n1220) );
  NANDN U1270 ( .A(n1247), .B(n1248), .Z(n1180) );
  NAND U1271 ( .A(n1249), .B(n1250), .Z(n1248) );
  NANDN U1272 ( .A(n1251), .B(n1252), .Z(n1249) );
  NANDN U1273 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1274 ( .A(n1255), .B(n1256), .Z(n1254) );
  NAND U1275 ( .A(n1257), .B(n1258), .Z(n1256) );
  OR U1276 ( .A(n1170), .B(n1169), .Z(n1246) );
  NAND U1277 ( .A(n1259), .B(n1260), .Z(n1170) );
  AND U1278 ( .A(n1261), .B(n1257), .Z(n1260) );
  ANDN U1279 ( .B(n1250), .A(n1253), .Z(n1259) );
  XOR U1280 ( .A(n1262), .B(n1263), .Z(SUM[131]) );
  NANDN U1281 ( .A(n1247), .B(n1250), .Z(n1263) );
  OR U1282 ( .A(B[131]), .B(A[131]), .Z(n1250) );
  AND U1283 ( .A(B[131]), .B(A[131]), .Z(n1247) );
  ANDN U1284 ( .B(n1264), .A(n1251), .Z(n1262) );
  NANDN U1285 ( .A(n1253), .B(n1265), .Z(n1264) );
  XNOR U1286 ( .A(n1265), .B(n1266), .Z(SUM[130]) );
  OR U1287 ( .A(n1253), .B(n1251), .Z(n1266) );
  AND U1288 ( .A(B[130]), .B(A[130]), .Z(n1251) );
  NOR U1289 ( .A(B[130]), .B(A[130]), .Z(n1253) );
  NANDN U1290 ( .A(n1255), .B(n1267), .Z(n1265) );
  NAND U1291 ( .A(n1268), .B(n1257), .Z(n1267) );
  XNOR U1292 ( .A(n1268), .B(n1269), .Z(SUM[129]) );
  NANDN U1293 ( .A(n1255), .B(n1257), .Z(n1269) );
  OR U1294 ( .A(B[129]), .B(A[129]), .Z(n1257) );
  AND U1295 ( .A(B[129]), .B(A[129]), .Z(n1255) );
  NANDN U1296 ( .A(n1258), .B(n1270), .Z(n1268) );
  NANDN U1297 ( .A(n1169), .B(n1261), .Z(n1270) );
  XOR U1298 ( .A(n1169), .B(n1271), .Z(SUM[128]) );
  NANDN U1299 ( .A(n1258), .B(n1261), .Z(n1271) );
  OR U1300 ( .A(B[128]), .B(A[128]), .Z(n1261) );
  AND U1301 ( .A(A[128]), .B(B[128]), .Z(n1258) );
  ANDN U1302 ( .B(n1272), .A(n1273), .Z(n1169) );
  NANDN U1303 ( .A(n1274), .B(n1275), .Z(n1272) );
  NANDN U1304 ( .A(n1276), .B(n1277), .Z(n1275) );
  NANDN U1305 ( .A(n1278), .B(n1279), .Z(n1277) );
  NANDN U1306 ( .A(n1280), .B(n1281), .Z(n1279) );
  NANDN U1307 ( .A(n1282), .B(n1283), .Z(n1281) );
  NAND U1308 ( .A(n1284), .B(n1285), .Z(n1283) );
  NAND U1309 ( .A(n1286), .B(n1287), .Z(n1285) );
  AND U1310 ( .A(n1288), .B(n1289), .Z(n1287) );
  ANDN U1311 ( .B(n1290), .A(n1291), .Z(n1289) );
  NOR U1312 ( .A(n1292), .B(n1293), .Z(n1286) );
  ANDN U1313 ( .B(n1294), .A(n1295), .Z(n1284) );
  NAND U1314 ( .A(n1296), .B(n1290), .Z(n1294) );
  NANDN U1315 ( .A(n1297), .B(n1298), .Z(n1296) );
  NANDN U1316 ( .A(n1293), .B(n1299), .Z(n1298) );
  NANDN U1317 ( .A(n1300), .B(n1301), .Z(n1299) );
  NAND U1318 ( .A(n1302), .B(n1288), .Z(n1301) );
  XOR U1319 ( .A(n1303), .B(n1304), .Z(SUM[127]) );
  OR U1320 ( .A(n1274), .B(n1273), .Z(n1304) );
  AND U1321 ( .A(B[127]), .B(A[127]), .Z(n1273) );
  NOR U1322 ( .A(B[127]), .B(A[127]), .Z(n1274) );
  ANDN U1323 ( .B(n1305), .A(n1276), .Z(n1303) );
  NANDN U1324 ( .A(n1278), .B(n1306), .Z(n1305) );
  XNOR U1325 ( .A(n1306), .B(n1307), .Z(SUM[126]) );
  OR U1326 ( .A(n1278), .B(n1276), .Z(n1307) );
  AND U1327 ( .A(B[126]), .B(A[126]), .Z(n1276) );
  NOR U1328 ( .A(B[126]), .B(A[126]), .Z(n1278) );
  NANDN U1329 ( .A(n1280), .B(n1308), .Z(n1306) );
  NANDN U1330 ( .A(n1282), .B(n1309), .Z(n1308) );
  XNOR U1331 ( .A(n1309), .B(n1310), .Z(SUM[125]) );
  OR U1332 ( .A(n1282), .B(n1280), .Z(n1310) );
  AND U1333 ( .A(B[125]), .B(A[125]), .Z(n1280) );
  NOR U1334 ( .A(B[125]), .B(A[125]), .Z(n1282) );
  NANDN U1335 ( .A(n1295), .B(n1311), .Z(n1309) );
  NAND U1336 ( .A(n1312), .B(n1290), .Z(n1311) );
  XNOR U1337 ( .A(n1312), .B(n1313), .Z(SUM[124]) );
  NANDN U1338 ( .A(n1295), .B(n1290), .Z(n1313) );
  OR U1339 ( .A(A[124]), .B(B[124]), .Z(n1290) );
  AND U1340 ( .A(B[124]), .B(A[124]), .Z(n1295) );
  NANDN U1341 ( .A(n1297), .B(n1314), .Z(n1312) );
  NANDN U1342 ( .A(n1293), .B(n1315), .Z(n1314) );
  NAND U1343 ( .A(n1316), .B(n1317), .Z(n1293) );
  AND U1344 ( .A(n1318), .B(n1319), .Z(n1317) );
  AND U1345 ( .A(n1320), .B(n1321), .Z(n1316) );
  NANDN U1346 ( .A(n1322), .B(n1323), .Z(n1297) );
  NAND U1347 ( .A(n1324), .B(n1321), .Z(n1323) );
  NANDN U1348 ( .A(n1325), .B(n1326), .Z(n1324) );
  NAND U1349 ( .A(n1327), .B(n1320), .Z(n1326) );
  NANDN U1350 ( .A(n1328), .B(n1329), .Z(n1327) );
  NAND U1351 ( .A(n1319), .B(n1330), .Z(n1329) );
  XOR U1352 ( .A(n1331), .B(n1332), .Z(SUM[123]) );
  NANDN U1353 ( .A(n1322), .B(n1321), .Z(n1332) );
  OR U1354 ( .A(B[123]), .B(A[123]), .Z(n1321) );
  AND U1355 ( .A(B[123]), .B(A[123]), .Z(n1322) );
  ANDN U1356 ( .B(n1333), .A(n1325), .Z(n1331) );
  NAND U1357 ( .A(n1334), .B(n1320), .Z(n1333) );
  XNOR U1358 ( .A(n1334), .B(n1335), .Z(SUM[122]) );
  NANDN U1359 ( .A(n1325), .B(n1320), .Z(n1335) );
  OR U1360 ( .A(B[122]), .B(A[122]), .Z(n1320) );
  AND U1361 ( .A(B[122]), .B(A[122]), .Z(n1325) );
  NANDN U1362 ( .A(n1328), .B(n1336), .Z(n1334) );
  NAND U1363 ( .A(n1337), .B(n1319), .Z(n1336) );
  XNOR U1364 ( .A(n1337), .B(n1338), .Z(SUM[121]) );
  NANDN U1365 ( .A(n1328), .B(n1319), .Z(n1338) );
  OR U1366 ( .A(B[121]), .B(A[121]), .Z(n1319) );
  AND U1367 ( .A(B[121]), .B(A[121]), .Z(n1328) );
  NANDN U1368 ( .A(n1330), .B(n1339), .Z(n1337) );
  NAND U1369 ( .A(n1315), .B(n1318), .Z(n1339) );
  XNOR U1370 ( .A(n1315), .B(n1340), .Z(SUM[120]) );
  NANDN U1371 ( .A(n1330), .B(n1318), .Z(n1340) );
  OR U1372 ( .A(B[120]), .B(A[120]), .Z(n1318) );
  AND U1373 ( .A(B[120]), .B(A[120]), .Z(n1330) );
  NANDN U1374 ( .A(n1300), .B(n1341), .Z(n1315) );
  NANDN U1375 ( .A(n1342), .B(n1288), .Z(n1341) );
  AND U1376 ( .A(n1343), .B(n1344), .Z(n1288) );
  AND U1377 ( .A(n1345), .B(n1346), .Z(n1344) );
  AND U1378 ( .A(n1347), .B(n1348), .Z(n1343) );
  NANDN U1379 ( .A(n1349), .B(n1350), .Z(n1300) );
  NAND U1380 ( .A(n1351), .B(n1348), .Z(n1350) );
  NANDN U1381 ( .A(n1352), .B(n1353), .Z(n1351) );
  NAND U1382 ( .A(n1354), .B(n1347), .Z(n1353) );
  NANDN U1383 ( .A(n1355), .B(n1356), .Z(n1354) );
  NAND U1384 ( .A(n1346), .B(n1357), .Z(n1356) );
  XOR U1385 ( .A(n1358), .B(n1359), .Z(SUM[119]) );
  NANDN U1386 ( .A(n1349), .B(n1348), .Z(n1359) );
  OR U1387 ( .A(B[119]), .B(A[119]), .Z(n1348) );
  AND U1388 ( .A(B[119]), .B(A[119]), .Z(n1349) );
  ANDN U1389 ( .B(n1360), .A(n1352), .Z(n1358) );
  NAND U1390 ( .A(n1361), .B(n1347), .Z(n1360) );
  XNOR U1391 ( .A(n1361), .B(n1362), .Z(SUM[118]) );
  NANDN U1392 ( .A(n1352), .B(n1347), .Z(n1362) );
  OR U1393 ( .A(B[118]), .B(A[118]), .Z(n1347) );
  AND U1394 ( .A(B[118]), .B(A[118]), .Z(n1352) );
  NANDN U1395 ( .A(n1355), .B(n1363), .Z(n1361) );
  NAND U1396 ( .A(n1364), .B(n1346), .Z(n1363) );
  XNOR U1397 ( .A(n1364), .B(n1365), .Z(SUM[117]) );
  NANDN U1398 ( .A(n1355), .B(n1346), .Z(n1365) );
  OR U1399 ( .A(B[117]), .B(A[117]), .Z(n1346) );
  AND U1400 ( .A(B[117]), .B(A[117]), .Z(n1355) );
  NANDN U1401 ( .A(n1357), .B(n1366), .Z(n1364) );
  NANDN U1402 ( .A(n1342), .B(n1345), .Z(n1366) );
  XOR U1403 ( .A(n1342), .B(n1367), .Z(SUM[116]) );
  NANDN U1404 ( .A(n1357), .B(n1345), .Z(n1367) );
  OR U1405 ( .A(B[116]), .B(A[116]), .Z(n1345) );
  AND U1406 ( .A(B[116]), .B(A[116]), .Z(n1357) );
  ANDN U1407 ( .B(n1368), .A(n1302), .Z(n1342) );
  NANDN U1408 ( .A(n1369), .B(n1370), .Z(n1302) );
  NAND U1409 ( .A(n1371), .B(n1372), .Z(n1370) );
  NANDN U1410 ( .A(n1373), .B(n1374), .Z(n1371) );
  NANDN U1411 ( .A(n1375), .B(n1376), .Z(n1374) );
  NANDN U1412 ( .A(n1377), .B(n1378), .Z(n1376) );
  NAND U1413 ( .A(n1379), .B(n1380), .Z(n1378) );
  OR U1414 ( .A(n1292), .B(n1291), .Z(n1368) );
  NAND U1415 ( .A(n1381), .B(n1382), .Z(n1292) );
  AND U1416 ( .A(n1383), .B(n1379), .Z(n1382) );
  ANDN U1417 ( .B(n1372), .A(n1375), .Z(n1381) );
  XOR U1418 ( .A(n1384), .B(n1385), .Z(SUM[115]) );
  NANDN U1419 ( .A(n1369), .B(n1372), .Z(n1385) );
  OR U1420 ( .A(B[115]), .B(A[115]), .Z(n1372) );
  AND U1421 ( .A(B[115]), .B(A[115]), .Z(n1369) );
  ANDN U1422 ( .B(n1386), .A(n1373), .Z(n1384) );
  NANDN U1423 ( .A(n1375), .B(n1387), .Z(n1386) );
  XNOR U1424 ( .A(n1387), .B(n1388), .Z(SUM[114]) );
  OR U1425 ( .A(n1375), .B(n1373), .Z(n1388) );
  AND U1426 ( .A(B[114]), .B(A[114]), .Z(n1373) );
  NOR U1427 ( .A(B[114]), .B(A[114]), .Z(n1375) );
  NANDN U1428 ( .A(n1377), .B(n1389), .Z(n1387) );
  NAND U1429 ( .A(n1390), .B(n1379), .Z(n1389) );
  XNOR U1430 ( .A(n1390), .B(n1391), .Z(SUM[113]) );
  NANDN U1431 ( .A(n1377), .B(n1379), .Z(n1391) );
  OR U1432 ( .A(B[113]), .B(A[113]), .Z(n1379) );
  AND U1433 ( .A(B[113]), .B(A[113]), .Z(n1377) );
  NANDN U1434 ( .A(n1380), .B(n1392), .Z(n1390) );
  NANDN U1435 ( .A(n1291), .B(n1383), .Z(n1392) );
  XOR U1436 ( .A(n1291), .B(n1393), .Z(SUM[112]) );
  NANDN U1437 ( .A(n1380), .B(n1383), .Z(n1393) );
  OR U1438 ( .A(B[112]), .B(A[112]), .Z(n1383) );
  AND U1439 ( .A(A[112]), .B(B[112]), .Z(n1380) );
  ANDN U1440 ( .B(n1394), .A(n1395), .Z(n1291) );
  NANDN U1441 ( .A(n1396), .B(n1397), .Z(n1394) );
  NANDN U1442 ( .A(n1398), .B(n1399), .Z(n1397) );
  NANDN U1443 ( .A(n1400), .B(n1401), .Z(n1399) );
  NANDN U1444 ( .A(n1402), .B(n1403), .Z(n1401) );
  NANDN U1445 ( .A(n1404), .B(n1405), .Z(n1403) );
  NAND U1446 ( .A(n1406), .B(n1407), .Z(n1405) );
  NAND U1447 ( .A(n1408), .B(n1409), .Z(n1407) );
  AND U1448 ( .A(n1410), .B(n1411), .Z(n1409) );
  ANDN U1449 ( .B(n1412), .A(n17), .Z(n1411) );
  NOR U1450 ( .A(n1413), .B(n1414), .Z(n1408) );
  ANDN U1451 ( .B(n1415), .A(n1416), .Z(n1406) );
  NAND U1452 ( .A(n1417), .B(n1412), .Z(n1415) );
  NANDN U1453 ( .A(n1418), .B(n1419), .Z(n1417) );
  NANDN U1454 ( .A(n1414), .B(n1420), .Z(n1419) );
  NANDN U1455 ( .A(n1421), .B(n1422), .Z(n1420) );
  NAND U1456 ( .A(n1423), .B(n1410), .Z(n1422) );
  XOR U1457 ( .A(n1424), .B(n1425), .Z(SUM[111]) );
  OR U1458 ( .A(n1396), .B(n1395), .Z(n1425) );
  AND U1459 ( .A(B[111]), .B(A[111]), .Z(n1395) );
  NOR U1460 ( .A(B[111]), .B(A[111]), .Z(n1396) );
  ANDN U1461 ( .B(n1426), .A(n1398), .Z(n1424) );
  NANDN U1462 ( .A(n1400), .B(n1427), .Z(n1426) );
  XNOR U1463 ( .A(n1427), .B(n1428), .Z(SUM[110]) );
  OR U1464 ( .A(n1400), .B(n1398), .Z(n1428) );
  AND U1465 ( .A(B[110]), .B(A[110]), .Z(n1398) );
  NOR U1466 ( .A(B[110]), .B(A[110]), .Z(n1400) );
  NANDN U1467 ( .A(n1402), .B(n1429), .Z(n1427) );
  NANDN U1468 ( .A(n1404), .B(n1430), .Z(n1429) );
  XNOR U1469 ( .A(n1430), .B(n1431), .Z(SUM[109]) );
  OR U1470 ( .A(n1404), .B(n1402), .Z(n1431) );
  AND U1471 ( .A(B[109]), .B(A[109]), .Z(n1402) );
  NOR U1472 ( .A(B[109]), .B(A[109]), .Z(n1404) );
  NANDN U1473 ( .A(n1416), .B(n1432), .Z(n1430) );
  NAND U1474 ( .A(n1433), .B(n1412), .Z(n1432) );
  XNOR U1475 ( .A(n1433), .B(n1434), .Z(SUM[108]) );
  NANDN U1476 ( .A(n1416), .B(n1412), .Z(n1434) );
  OR U1477 ( .A(A[108]), .B(B[108]), .Z(n1412) );
  AND U1478 ( .A(B[108]), .B(A[108]), .Z(n1416) );
  NANDN U1479 ( .A(n1418), .B(n1435), .Z(n1433) );
  NANDN U1480 ( .A(n1414), .B(n1436), .Z(n1435) );
  NAND U1481 ( .A(n1437), .B(n1438), .Z(n1414) );
  AND U1482 ( .A(n1439), .B(n1440), .Z(n1438) );
  AND U1483 ( .A(n1441), .B(n1442), .Z(n1437) );
  NANDN U1484 ( .A(n1443), .B(n1444), .Z(n1418) );
  NAND U1485 ( .A(n1445), .B(n1442), .Z(n1444) );
  NANDN U1486 ( .A(n1446), .B(n1447), .Z(n1445) );
  NAND U1487 ( .A(n1448), .B(n1441), .Z(n1447) );
  NANDN U1488 ( .A(n1449), .B(n1450), .Z(n1448) );
  NAND U1489 ( .A(n1440), .B(n1451), .Z(n1450) );
  XOR U1490 ( .A(n1452), .B(n1453), .Z(SUM[107]) );
  NANDN U1491 ( .A(n1443), .B(n1442), .Z(n1453) );
  OR U1492 ( .A(B[107]), .B(A[107]), .Z(n1442) );
  AND U1493 ( .A(B[107]), .B(A[107]), .Z(n1443) );
  ANDN U1494 ( .B(n1454), .A(n1446), .Z(n1452) );
  NAND U1495 ( .A(n1455), .B(n1441), .Z(n1454) );
  XNOR U1496 ( .A(n1455), .B(n1456), .Z(SUM[106]) );
  NANDN U1497 ( .A(n1446), .B(n1441), .Z(n1456) );
  OR U1498 ( .A(B[106]), .B(A[106]), .Z(n1441) );
  AND U1499 ( .A(B[106]), .B(A[106]), .Z(n1446) );
  NANDN U1500 ( .A(n1449), .B(n1457), .Z(n1455) );
  NAND U1501 ( .A(n1458), .B(n1440), .Z(n1457) );
  XNOR U1502 ( .A(n1458), .B(n1459), .Z(SUM[105]) );
  NANDN U1503 ( .A(n1449), .B(n1440), .Z(n1459) );
  OR U1504 ( .A(B[105]), .B(A[105]), .Z(n1440) );
  AND U1505 ( .A(B[105]), .B(A[105]), .Z(n1449) );
  NANDN U1506 ( .A(n1451), .B(n1460), .Z(n1458) );
  NAND U1507 ( .A(n1436), .B(n1439), .Z(n1460) );
  XNOR U1508 ( .A(n1436), .B(n1461), .Z(SUM[104]) );
  NANDN U1509 ( .A(n1451), .B(n1439), .Z(n1461) );
  OR U1510 ( .A(B[104]), .B(A[104]), .Z(n1439) );
  AND U1511 ( .A(B[104]), .B(A[104]), .Z(n1451) );
  NANDN U1512 ( .A(n1421), .B(n1462), .Z(n1436) );
  NANDN U1513 ( .A(n1463), .B(n1410), .Z(n1462) );
  AND U1514 ( .A(n1464), .B(n1465), .Z(n1410) );
  AND U1515 ( .A(n1466), .B(n1467), .Z(n1465) );
  AND U1516 ( .A(n1468), .B(n1469), .Z(n1464) );
  NANDN U1517 ( .A(n1470), .B(n1471), .Z(n1421) );
  NAND U1518 ( .A(n1472), .B(n1469), .Z(n1471) );
  NANDN U1519 ( .A(n1473), .B(n1474), .Z(n1472) );
  NAND U1520 ( .A(n1475), .B(n1468), .Z(n1474) );
  NANDN U1521 ( .A(n1476), .B(n1477), .Z(n1475) );
  NAND U1522 ( .A(n1467), .B(n1478), .Z(n1477) );
  XOR U1523 ( .A(n1479), .B(n1480), .Z(SUM[103]) );
  NANDN U1524 ( .A(n1470), .B(n1469), .Z(n1480) );
  OR U1525 ( .A(B[103]), .B(A[103]), .Z(n1469) );
  AND U1526 ( .A(B[103]), .B(A[103]), .Z(n1470) );
  ANDN U1527 ( .B(n1481), .A(n1473), .Z(n1479) );
  NAND U1528 ( .A(n1482), .B(n1468), .Z(n1481) );
  XNOR U1529 ( .A(n1482), .B(n1483), .Z(SUM[102]) );
  NANDN U1530 ( .A(n1473), .B(n1468), .Z(n1483) );
  OR U1531 ( .A(B[102]), .B(A[102]), .Z(n1468) );
  AND U1532 ( .A(B[102]), .B(A[102]), .Z(n1473) );
  NANDN U1533 ( .A(n1476), .B(n1484), .Z(n1482) );
  NAND U1534 ( .A(n1485), .B(n1467), .Z(n1484) );
  XNOR U1535 ( .A(n1485), .B(n1486), .Z(SUM[101]) );
  NANDN U1536 ( .A(n1476), .B(n1467), .Z(n1486) );
  OR U1537 ( .A(B[101]), .B(A[101]), .Z(n1467) );
  AND U1538 ( .A(B[101]), .B(A[101]), .Z(n1476) );
  NANDN U1539 ( .A(n1478), .B(n1487), .Z(n1485) );
  NANDN U1540 ( .A(n1463), .B(n1466), .Z(n1487) );
  XOR U1541 ( .A(n1463), .B(n1488), .Z(SUM[100]) );
  NANDN U1542 ( .A(n1478), .B(n1466), .Z(n1488) );
  OR U1543 ( .A(B[100]), .B(A[100]), .Z(n1466) );
  AND U1544 ( .A(B[100]), .B(A[100]), .Z(n1478) );
  ANDN U1545 ( .B(n1489), .A(n1423), .Z(n1463) );
  NANDN U1546 ( .A(n3), .B(n1490), .Z(n1423) );
  NAND U1547 ( .A(n1491), .B(n4), .Z(n1490) );
  NANDN U1548 ( .A(n6), .B(n1492), .Z(n1491) );
  NAND U1549 ( .A(n1493), .B(n8), .Z(n1492) );
  NANDN U1550 ( .A(n10), .B(n1494), .Z(n1493) );
  NANDN U1551 ( .A(n15), .B(n13), .Z(n1494) );
  NAND U1552 ( .A(B[96]), .B(A[96]), .Z(n15) );
  AND U1553 ( .A(B[97]), .B(A[97]), .Z(n10) );
  AND U1554 ( .A(A[98]), .B(B[98]), .Z(n6) );
  AND U1555 ( .A(B[99]), .B(A[99]), .Z(n3) );
  OR U1556 ( .A(n1413), .B(n17), .Z(n1489) );
  ANDN U1557 ( .B(n1495), .A(n23), .Z(n17) );
  AND U1558 ( .A(B[95]), .B(A[95]), .Z(n23) );
  NANDN U1559 ( .A(n22), .B(n1496), .Z(n1495) );
  NANDN U1560 ( .A(n25), .B(n1497), .Z(n1496) );
  NANDN U1561 ( .A(n26), .B(n1498), .Z(n1497) );
  NANDN U1562 ( .A(n29), .B(n1499), .Z(n1498) );
  NANDN U1563 ( .A(n31), .B(n1500), .Z(n1499) );
  NAND U1564 ( .A(n1501), .B(n1502), .Z(n1500) );
  NAND U1565 ( .A(n1503), .B(n1504), .Z(n1502) );
  AND U1566 ( .A(n64), .B(n1505), .Z(n1504) );
  ANDN U1567 ( .B(n37), .A(n86), .Z(n1505) );
  ANDN U1568 ( .B(n1506), .A(n108), .Z(n86) );
  AND U1569 ( .A(B[79]), .B(A[79]), .Z(n108) );
  NANDN U1570 ( .A(n107), .B(n1507), .Z(n1506) );
  NANDN U1571 ( .A(n110), .B(n1508), .Z(n1507) );
  NANDN U1572 ( .A(n111), .B(n1509), .Z(n1508) );
  NANDN U1573 ( .A(n114), .B(n1510), .Z(n1509) );
  NANDN U1574 ( .A(n116), .B(n1511), .Z(n1510) );
  NAND U1575 ( .A(n1512), .B(n1513), .Z(n1511) );
  NAND U1576 ( .A(n1514), .B(n1515), .Z(n1513) );
  AND U1577 ( .A(n149), .B(n1516), .Z(n1515) );
  ANDN U1578 ( .B(n122), .A(n171), .Z(n1516) );
  ANDN U1579 ( .B(n1517), .A(n193), .Z(n171) );
  AND U1580 ( .A(B[63]), .B(A[63]), .Z(n193) );
  NANDN U1581 ( .A(n192), .B(n1518), .Z(n1517) );
  NANDN U1582 ( .A(n195), .B(n1519), .Z(n1518) );
  NANDN U1583 ( .A(n196), .B(n1520), .Z(n1519) );
  NANDN U1584 ( .A(n199), .B(n1521), .Z(n1520) );
  NANDN U1585 ( .A(n201), .B(n1522), .Z(n1521) );
  NANDN U1586 ( .A(n204), .B(n1523), .Z(n1522) );
  NANDN U1587 ( .A(n206), .B(n1524), .Z(n1523) );
  NANDN U1588 ( .A(n209), .B(n1525), .Z(n1524) );
  NANDN U1589 ( .A(n211), .B(n1526), .Z(n1525) );
  NANDN U1590 ( .A(n231), .B(n1527), .Z(n1526) );
  AND U1591 ( .A(n1528), .B(n1529), .Z(n1527) );
  NANDN U1592 ( .A(n233), .B(n253), .Z(n1529) );
  NANDN U1593 ( .A(n257), .B(n1530), .Z(n253) );
  NAND U1594 ( .A(n1531), .B(n258), .Z(n1530) );
  NANDN U1595 ( .A(n260), .B(n1532), .Z(n1531) );
  NAND U1596 ( .A(n1533), .B(n262), .Z(n1532) );
  NANDN U1597 ( .A(n264), .B(n1534), .Z(n1533) );
  NAND U1598 ( .A(n267), .B(n269), .Z(n1534) );
  AND U1599 ( .A(A[48]), .B(B[48]), .Z(n269) );
  AND U1600 ( .A(A[49]), .B(B[49]), .Z(n264) );
  AND U1601 ( .A(A[50]), .B(B[50]), .Z(n260) );
  AND U1602 ( .A(B[51]), .B(A[51]), .Z(n257) );
  NANDN U1603 ( .A(n233), .B(n254), .Z(n1528) );
  AND U1604 ( .A(n1535), .B(n1536), .Z(n254) );
  AND U1605 ( .A(n262), .B(n1537), .Z(n1536) );
  AND U1606 ( .A(n272), .B(n267), .Z(n1537) );
  OR U1607 ( .A(A[49]), .B(B[49]), .Z(n267) );
  OR U1608 ( .A(A[48]), .B(B[48]), .Z(n272) );
  OR U1609 ( .A(A[50]), .B(B[50]), .Z(n262) );
  ANDN U1610 ( .B(n258), .A(n271), .Z(n1535) );
  ANDN U1611 ( .B(n1538), .A(n277), .Z(n271) );
  AND U1612 ( .A(B[47]), .B(A[47]), .Z(n277) );
  NANDN U1613 ( .A(n276), .B(n1539), .Z(n1538) );
  NANDN U1614 ( .A(n279), .B(n1540), .Z(n1539) );
  NANDN U1615 ( .A(n280), .B(n1541), .Z(n1540) );
  NANDN U1616 ( .A(n283), .B(n1542), .Z(n1541) );
  NANDN U1617 ( .A(n285), .B(n1543), .Z(n1542) );
  NAND U1618 ( .A(n1544), .B(n1545), .Z(n1543) );
  NAND U1619 ( .A(n1546), .B(n1547), .Z(n1545) );
  ANDN U1620 ( .B(n1548), .A(n295), .Z(n1547) );
  AND U1621 ( .A(n291), .B(n318), .Z(n1548) );
  ANDN U1622 ( .B(n340), .A(n339), .Z(n1546) );
  NAND U1623 ( .A(n1549), .B(n1550), .Z(n339) );
  AND U1624 ( .A(n357), .B(n353), .Z(n1550) );
  OR U1625 ( .A(B[32]), .B(A[32]), .Z(n357) );
  ANDN U1626 ( .B(n344), .A(n347), .Z(n1549) );
  AND U1627 ( .A(A[31]), .B(B[31]), .Z(n340) );
  ANDN U1628 ( .B(n1551), .A(n288), .Z(n1544) );
  AND U1629 ( .A(B[44]), .B(A[44]), .Z(n288) );
  NAND U1630 ( .A(n1552), .B(n291), .Z(n1551) );
  OR U1631 ( .A(A[44]), .B(B[44]), .Z(n291) );
  NANDN U1632 ( .A(n293), .B(n1553), .Z(n1552) );
  NANDN U1633 ( .A(n295), .B(n1554), .Z(n1553) );
  NANDN U1634 ( .A(n315), .B(n1555), .Z(n1554) );
  NAND U1635 ( .A(n338), .B(n318), .Z(n1555) );
  AND U1636 ( .A(n1556), .B(n1557), .Z(n318) );
  AND U1637 ( .A(n335), .B(n331), .Z(n1557) );
  OR U1638 ( .A(B[36]), .B(A[36]), .Z(n335) );
  AND U1639 ( .A(n326), .B(n322), .Z(n1556) );
  NANDN U1640 ( .A(n343), .B(n1558), .Z(n338) );
  NAND U1641 ( .A(n1559), .B(n344), .Z(n1558) );
  OR U1642 ( .A(B[35]), .B(A[35]), .Z(n344) );
  NANDN U1643 ( .A(n346), .B(n1560), .Z(n1559) );
  NANDN U1644 ( .A(n347), .B(n1561), .Z(n1560) );
  NANDN U1645 ( .A(n350), .B(n1562), .Z(n1561) );
  NAND U1646 ( .A(n353), .B(n355), .Z(n1562) );
  AND U1647 ( .A(A[32]), .B(B[32]), .Z(n355) );
  OR U1648 ( .A(B[33]), .B(A[33]), .Z(n353) );
  AND U1649 ( .A(B[33]), .B(A[33]), .Z(n350) );
  NOR U1650 ( .A(B[34]), .B(A[34]), .Z(n347) );
  AND U1651 ( .A(B[34]), .B(A[34]), .Z(n346) );
  AND U1652 ( .A(B[35]), .B(A[35]), .Z(n343) );
  NANDN U1653 ( .A(n321), .B(n1563), .Z(n315) );
  NAND U1654 ( .A(n1564), .B(n322), .Z(n1563) );
  OR U1655 ( .A(B[39]), .B(A[39]), .Z(n322) );
  NANDN U1656 ( .A(n324), .B(n1565), .Z(n1564) );
  NAND U1657 ( .A(n1566), .B(n326), .Z(n1565) );
  OR U1658 ( .A(B[38]), .B(A[38]), .Z(n326) );
  NANDN U1659 ( .A(n328), .B(n1567), .Z(n1566) );
  NAND U1660 ( .A(n331), .B(n333), .Z(n1567) );
  AND U1661 ( .A(B[36]), .B(A[36]), .Z(n333) );
  OR U1662 ( .A(B[37]), .B(A[37]), .Z(n331) );
  AND U1663 ( .A(B[37]), .B(A[37]), .Z(n328) );
  AND U1664 ( .A(B[38]), .B(A[38]), .Z(n324) );
  AND U1665 ( .A(B[39]), .B(A[39]), .Z(n321) );
  NAND U1666 ( .A(n1568), .B(n1569), .Z(n295) );
  AND U1667 ( .A(n313), .B(n309), .Z(n1569) );
  OR U1668 ( .A(B[40]), .B(A[40]), .Z(n313) );
  AND U1669 ( .A(n304), .B(n300), .Z(n1568) );
  NANDN U1670 ( .A(n299), .B(n1570), .Z(n293) );
  NAND U1671 ( .A(n1571), .B(n300), .Z(n1570) );
  OR U1672 ( .A(B[43]), .B(A[43]), .Z(n300) );
  NANDN U1673 ( .A(n302), .B(n1572), .Z(n1571) );
  NAND U1674 ( .A(n1573), .B(n304), .Z(n1572) );
  OR U1675 ( .A(B[42]), .B(A[42]), .Z(n304) );
  NANDN U1676 ( .A(n306), .B(n1574), .Z(n1573) );
  NAND U1677 ( .A(n309), .B(n311), .Z(n1574) );
  AND U1678 ( .A(B[40]), .B(A[40]), .Z(n311) );
  OR U1679 ( .A(B[41]), .B(A[41]), .Z(n309) );
  AND U1680 ( .A(B[41]), .B(A[41]), .Z(n306) );
  AND U1681 ( .A(B[42]), .B(A[42]), .Z(n302) );
  AND U1682 ( .A(B[43]), .B(A[43]), .Z(n299) );
  NOR U1683 ( .A(B[45]), .B(A[45]), .Z(n285) );
  AND U1684 ( .A(B[45]), .B(A[45]), .Z(n283) );
  NOR U1685 ( .A(B[46]), .B(A[46]), .Z(n280) );
  AND U1686 ( .A(B[46]), .B(A[46]), .Z(n279) );
  NOR U1687 ( .A(B[47]), .B(A[47]), .Z(n276) );
  OR U1688 ( .A(B[51]), .B(A[51]), .Z(n258) );
  NAND U1689 ( .A(n1575), .B(n1576), .Z(n233) );
  AND U1690 ( .A(n251), .B(n247), .Z(n1576) );
  OR U1691 ( .A(A[52]), .B(B[52]), .Z(n251) );
  AND U1692 ( .A(n242), .B(n238), .Z(n1575) );
  NANDN U1693 ( .A(n237), .B(n1577), .Z(n231) );
  NAND U1694 ( .A(n1578), .B(n238), .Z(n1577) );
  OR U1695 ( .A(B[55]), .B(A[55]), .Z(n238) );
  NANDN U1696 ( .A(n240), .B(n1579), .Z(n1578) );
  NAND U1697 ( .A(n1580), .B(n242), .Z(n1579) );
  OR U1698 ( .A(A[54]), .B(B[54]), .Z(n242) );
  NANDN U1699 ( .A(n244), .B(n1581), .Z(n1580) );
  NAND U1700 ( .A(n247), .B(n249), .Z(n1581) );
  AND U1701 ( .A(A[52]), .B(B[52]), .Z(n249) );
  OR U1702 ( .A(A[53]), .B(B[53]), .Z(n247) );
  AND U1703 ( .A(A[53]), .B(B[53]), .Z(n244) );
  AND U1704 ( .A(A[54]), .B(B[54]), .Z(n240) );
  AND U1705 ( .A(B[55]), .B(A[55]), .Z(n237) );
  NAND U1706 ( .A(n1582), .B(n1583), .Z(n211) );
  AND U1707 ( .A(n229), .B(n225), .Z(n1583) );
  OR U1708 ( .A(B[56]), .B(A[56]), .Z(n229) );
  AND U1709 ( .A(n220), .B(n216), .Z(n1582) );
  NANDN U1710 ( .A(n215), .B(n1584), .Z(n209) );
  NAND U1711 ( .A(n1585), .B(n216), .Z(n1584) );
  OR U1712 ( .A(B[59]), .B(A[59]), .Z(n216) );
  NANDN U1713 ( .A(n218), .B(n1586), .Z(n1585) );
  NAND U1714 ( .A(n1587), .B(n220), .Z(n1586) );
  OR U1715 ( .A(B[58]), .B(A[58]), .Z(n220) );
  NANDN U1716 ( .A(n222), .B(n1588), .Z(n1587) );
  NAND U1717 ( .A(n225), .B(n227), .Z(n1588) );
  AND U1718 ( .A(B[56]), .B(A[56]), .Z(n227) );
  OR U1719 ( .A(B[57]), .B(A[57]), .Z(n225) );
  AND U1720 ( .A(B[57]), .B(A[57]), .Z(n222) );
  AND U1721 ( .A(B[58]), .B(A[58]), .Z(n218) );
  AND U1722 ( .A(B[59]), .B(A[59]), .Z(n215) );
  NOR U1723 ( .A(B[60]), .B(A[60]), .Z(n206) );
  AND U1724 ( .A(B[60]), .B(A[60]), .Z(n204) );
  NOR U1725 ( .A(B[61]), .B(A[61]), .Z(n201) );
  AND U1726 ( .A(B[61]), .B(A[61]), .Z(n199) );
  NOR U1727 ( .A(B[62]), .B(A[62]), .Z(n196) );
  AND U1728 ( .A(B[62]), .B(A[62]), .Z(n195) );
  NOR U1729 ( .A(B[63]), .B(A[63]), .Z(n192) );
  NOR U1730 ( .A(n170), .B(n126), .Z(n1514) );
  NAND U1731 ( .A(n1589), .B(n1590), .Z(n170) );
  AND U1732 ( .A(n188), .B(n184), .Z(n1590) );
  OR U1733 ( .A(B[64]), .B(A[64]), .Z(n188) );
  ANDN U1734 ( .B(n175), .A(n178), .Z(n1589) );
  ANDN U1735 ( .B(n1591), .A(n119), .Z(n1512) );
  AND U1736 ( .A(B[76]), .B(A[76]), .Z(n119) );
  NAND U1737 ( .A(n1592), .B(n122), .Z(n1591) );
  OR U1738 ( .A(A[76]), .B(B[76]), .Z(n122) );
  NANDN U1739 ( .A(n124), .B(n1593), .Z(n1592) );
  NANDN U1740 ( .A(n126), .B(n1594), .Z(n1593) );
  NANDN U1741 ( .A(n146), .B(n1595), .Z(n1594) );
  NAND U1742 ( .A(n169), .B(n149), .Z(n1595) );
  AND U1743 ( .A(n1596), .B(n1597), .Z(n149) );
  AND U1744 ( .A(n166), .B(n162), .Z(n1597) );
  OR U1745 ( .A(B[68]), .B(A[68]), .Z(n166) );
  AND U1746 ( .A(n157), .B(n153), .Z(n1596) );
  NANDN U1747 ( .A(n174), .B(n1598), .Z(n169) );
  NAND U1748 ( .A(n1599), .B(n175), .Z(n1598) );
  OR U1749 ( .A(B[67]), .B(A[67]), .Z(n175) );
  NANDN U1750 ( .A(n177), .B(n1600), .Z(n1599) );
  NANDN U1751 ( .A(n178), .B(n1601), .Z(n1600) );
  NANDN U1752 ( .A(n181), .B(n1602), .Z(n1601) );
  NAND U1753 ( .A(n184), .B(n186), .Z(n1602) );
  AND U1754 ( .A(A[64]), .B(B[64]), .Z(n186) );
  OR U1755 ( .A(B[65]), .B(A[65]), .Z(n184) );
  AND U1756 ( .A(B[65]), .B(A[65]), .Z(n181) );
  NOR U1757 ( .A(B[66]), .B(A[66]), .Z(n178) );
  AND U1758 ( .A(B[66]), .B(A[66]), .Z(n177) );
  AND U1759 ( .A(B[67]), .B(A[67]), .Z(n174) );
  NANDN U1760 ( .A(n152), .B(n1603), .Z(n146) );
  NAND U1761 ( .A(n1604), .B(n153), .Z(n1603) );
  OR U1762 ( .A(B[71]), .B(A[71]), .Z(n153) );
  NANDN U1763 ( .A(n155), .B(n1605), .Z(n1604) );
  NAND U1764 ( .A(n1606), .B(n157), .Z(n1605) );
  OR U1765 ( .A(B[70]), .B(A[70]), .Z(n157) );
  NANDN U1766 ( .A(n159), .B(n1607), .Z(n1606) );
  NAND U1767 ( .A(n162), .B(n164), .Z(n1607) );
  AND U1768 ( .A(B[68]), .B(A[68]), .Z(n164) );
  OR U1769 ( .A(B[69]), .B(A[69]), .Z(n162) );
  AND U1770 ( .A(B[69]), .B(A[69]), .Z(n159) );
  AND U1771 ( .A(B[70]), .B(A[70]), .Z(n155) );
  AND U1772 ( .A(B[71]), .B(A[71]), .Z(n152) );
  NAND U1773 ( .A(n1608), .B(n1609), .Z(n126) );
  AND U1774 ( .A(n144), .B(n140), .Z(n1609) );
  OR U1775 ( .A(B[72]), .B(A[72]), .Z(n144) );
  AND U1776 ( .A(n135), .B(n131), .Z(n1608) );
  NANDN U1777 ( .A(n130), .B(n1610), .Z(n124) );
  NAND U1778 ( .A(n1611), .B(n131), .Z(n1610) );
  OR U1779 ( .A(B[75]), .B(A[75]), .Z(n131) );
  NANDN U1780 ( .A(n133), .B(n1612), .Z(n1611) );
  NAND U1781 ( .A(n1613), .B(n135), .Z(n1612) );
  OR U1782 ( .A(B[74]), .B(A[74]), .Z(n135) );
  NANDN U1783 ( .A(n137), .B(n1614), .Z(n1613) );
  NAND U1784 ( .A(n140), .B(n142), .Z(n1614) );
  AND U1785 ( .A(B[72]), .B(A[72]), .Z(n142) );
  OR U1786 ( .A(B[73]), .B(A[73]), .Z(n140) );
  AND U1787 ( .A(B[73]), .B(A[73]), .Z(n137) );
  AND U1788 ( .A(B[74]), .B(A[74]), .Z(n133) );
  AND U1789 ( .A(B[75]), .B(A[75]), .Z(n130) );
  NOR U1790 ( .A(B[77]), .B(A[77]), .Z(n116) );
  AND U1791 ( .A(B[77]), .B(A[77]), .Z(n114) );
  NOR U1792 ( .A(B[78]), .B(A[78]), .Z(n111) );
  AND U1793 ( .A(B[78]), .B(A[78]), .Z(n110) );
  NOR U1794 ( .A(B[79]), .B(A[79]), .Z(n107) );
  NOR U1795 ( .A(n85), .B(n41), .Z(n1503) );
  NAND U1796 ( .A(n1615), .B(n1616), .Z(n85) );
  AND U1797 ( .A(n103), .B(n99), .Z(n1616) );
  OR U1798 ( .A(B[80]), .B(A[80]), .Z(n103) );
  ANDN U1799 ( .B(n90), .A(n93), .Z(n1615) );
  ANDN U1800 ( .B(n1617), .A(n34), .Z(n1501) );
  AND U1801 ( .A(B[92]), .B(A[92]), .Z(n34) );
  NAND U1802 ( .A(n1618), .B(n37), .Z(n1617) );
  OR U1803 ( .A(A[92]), .B(B[92]), .Z(n37) );
  NANDN U1804 ( .A(n39), .B(n1619), .Z(n1618) );
  NANDN U1805 ( .A(n41), .B(n1620), .Z(n1619) );
  NANDN U1806 ( .A(n61), .B(n1621), .Z(n1620) );
  NAND U1807 ( .A(n84), .B(n64), .Z(n1621) );
  AND U1808 ( .A(n1622), .B(n1623), .Z(n64) );
  AND U1809 ( .A(n81), .B(n77), .Z(n1623) );
  OR U1810 ( .A(B[84]), .B(A[84]), .Z(n81) );
  AND U1811 ( .A(n72), .B(n68), .Z(n1622) );
  NANDN U1812 ( .A(n89), .B(n1624), .Z(n84) );
  NAND U1813 ( .A(n1625), .B(n90), .Z(n1624) );
  OR U1814 ( .A(B[83]), .B(A[83]), .Z(n90) );
  NANDN U1815 ( .A(n92), .B(n1626), .Z(n1625) );
  NANDN U1816 ( .A(n93), .B(n1627), .Z(n1626) );
  NANDN U1817 ( .A(n96), .B(n1628), .Z(n1627) );
  NAND U1818 ( .A(n99), .B(n101), .Z(n1628) );
  AND U1819 ( .A(A[80]), .B(B[80]), .Z(n101) );
  OR U1820 ( .A(B[81]), .B(A[81]), .Z(n99) );
  AND U1821 ( .A(B[81]), .B(A[81]), .Z(n96) );
  NOR U1822 ( .A(B[82]), .B(A[82]), .Z(n93) );
  AND U1823 ( .A(B[82]), .B(A[82]), .Z(n92) );
  AND U1824 ( .A(B[83]), .B(A[83]), .Z(n89) );
  NANDN U1825 ( .A(n67), .B(n1629), .Z(n61) );
  NAND U1826 ( .A(n1630), .B(n68), .Z(n1629) );
  OR U1827 ( .A(B[87]), .B(A[87]), .Z(n68) );
  NANDN U1828 ( .A(n70), .B(n1631), .Z(n1630) );
  NAND U1829 ( .A(n1632), .B(n72), .Z(n1631) );
  OR U1830 ( .A(B[86]), .B(A[86]), .Z(n72) );
  NANDN U1831 ( .A(n74), .B(n1633), .Z(n1632) );
  NAND U1832 ( .A(n77), .B(n79), .Z(n1633) );
  AND U1833 ( .A(B[84]), .B(A[84]), .Z(n79) );
  OR U1834 ( .A(B[85]), .B(A[85]), .Z(n77) );
  AND U1835 ( .A(B[85]), .B(A[85]), .Z(n74) );
  AND U1836 ( .A(B[86]), .B(A[86]), .Z(n70) );
  AND U1837 ( .A(B[87]), .B(A[87]), .Z(n67) );
  NAND U1838 ( .A(n1634), .B(n1635), .Z(n41) );
  AND U1839 ( .A(n59), .B(n55), .Z(n1635) );
  OR U1840 ( .A(B[88]), .B(A[88]), .Z(n59) );
  AND U1841 ( .A(n50), .B(n46), .Z(n1634) );
  NANDN U1842 ( .A(n45), .B(n1636), .Z(n39) );
  NAND U1843 ( .A(n1637), .B(n46), .Z(n1636) );
  OR U1844 ( .A(B[91]), .B(A[91]), .Z(n46) );
  NANDN U1845 ( .A(n48), .B(n1638), .Z(n1637) );
  NAND U1846 ( .A(n1639), .B(n50), .Z(n1638) );
  OR U1847 ( .A(B[90]), .B(A[90]), .Z(n50) );
  NANDN U1848 ( .A(n52), .B(n1640), .Z(n1639) );
  NAND U1849 ( .A(n55), .B(n57), .Z(n1640) );
  AND U1850 ( .A(B[88]), .B(A[88]), .Z(n57) );
  OR U1851 ( .A(B[89]), .B(A[89]), .Z(n55) );
  AND U1852 ( .A(B[89]), .B(A[89]), .Z(n52) );
  AND U1853 ( .A(B[90]), .B(A[90]), .Z(n48) );
  AND U1854 ( .A(B[91]), .B(A[91]), .Z(n45) );
  NOR U1855 ( .A(B[93]), .B(A[93]), .Z(n31) );
  AND U1856 ( .A(B[93]), .B(A[93]), .Z(n29) );
  NOR U1857 ( .A(B[94]), .B(A[94]), .Z(n26) );
  AND U1858 ( .A(B[94]), .B(A[94]), .Z(n25) );
  NOR U1859 ( .A(B[95]), .B(A[95]), .Z(n22) );
  NAND U1860 ( .A(n1641), .B(n1642), .Z(n1413) );
  AND U1861 ( .A(n13), .B(n8), .Z(n1642) );
  OR U1862 ( .A(B[98]), .B(A[98]), .Z(n8) );
  OR U1863 ( .A(B[97]), .B(A[97]), .Z(n13) );
  AND U1864 ( .A(n4), .B(n18), .Z(n1641) );
  OR U1865 ( .A(B[96]), .B(A[96]), .Z(n18) );
  OR U1866 ( .A(B[99]), .B(A[99]), .Z(n4) );
endmodule


module mult_N256_CC8_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [255:0] B;
  output [287:0] PRODUCT;
  input TC;
  wire   \A1[284] , \A1[283] , \A1[282] , \A1[281] , \A1[280] , \A1[279] ,
         \A1[278] , \A1[277] , \A1[276] , \A1[275] , \A1[274] , \A1[273] ,
         \A1[272] , \A1[271] , \A1[270] , \A1[269] , \A1[268] , \A1[267] ,
         \A1[266] , \A1[265] , \A1[264] , \A1[263] , \A1[262] , \A1[261] ,
         \A1[260] , \A1[259] , \A1[258] , \A1[257] , \A1[256] , \A1[255] ,
         \A1[254] , \A1[253] , \A1[252] , \A1[251] , \A1[250] , \A1[249] ,
         \A1[248] , \A1[247] , \A1[246] , \A1[245] , \A1[244] , \A1[243] ,
         \A1[242] , \A1[241] , \A1[240] , \A1[239] , \A1[238] , \A1[237] ,
         \A1[236] , \A1[235] , \A1[234] , \A1[233] , \A1[232] , \A1[231] ,
         \A1[230] , \A1[229] , \A1[228] , \A1[227] , \A1[226] , \A1[225] ,
         \A1[224] , \A1[223] , \A1[222] , \A1[221] , \A1[220] , \A1[219] ,
         \A1[218] , \A1[217] , \A1[216] , \A1[215] , \A1[214] , \A1[213] ,
         \A1[212] , \A1[211] , \A1[210] , \A1[209] , \A1[208] , \A1[207] ,
         \A1[206] , \A1[205] , \A1[204] , \A1[203] , \A1[202] , \A1[201] ,
         \A1[200] , \A1[199] , \A1[198] , \A1[197] , \A1[196] , \A1[195] ,
         \A1[194] , \A1[193] , \A1[192] , \A1[191] , \A1[190] , \A1[189] ,
         \A1[188] , \A1[187] , \A1[186] , \A1[185] , \A1[184] , \A1[183] ,
         \A1[182] , \A1[181] , \A1[180] , \A1[179] , \A1[178] , \A1[177] ,
         \A1[176] , \A1[175] , \A1[174] , \A1[173] , \A1[172] , \A1[171] ,
         \A1[170] , \A1[169] , \A1[168] , \A1[167] , \A1[166] , \A1[165] ,
         \A1[164] , \A1[163] , \A1[162] , \A1[161] , \A1[160] , \A1[159] ,
         \A1[158] , \A1[157] , \A1[156] , \A1[155] , \A1[154] , \A1[153] ,
         \A1[152] , \A1[151] , \A1[150] , \A1[149] , \A1[148] , \A1[147] ,
         \A1[146] , \A1[145] , \A1[144] , \A1[143] , \A1[142] , \A1[141] ,
         \A1[140] , \A1[139] , \A1[138] , \A1[137] , \A1[136] , \A1[135] ,
         \A1[134] , \A1[133] , \A1[132] , \A1[131] , \A1[130] , \A1[129] ,
         \A1[128] , \A1[127] , \A1[126] , \A1[125] , \A1[124] , \A1[123] ,
         \A1[122] , \A1[121] , \A1[120] , \A1[119] , \A1[118] , \A1[117] ,
         \A1[116] , \A1[115] , \A1[114] , \A1[113] , \A1[112] , \A1[111] ,
         \A1[110] , \A1[109] , \A1[108] , \A1[107] , \A1[106] , \A1[105] ,
         \A1[104] , \A1[103] , \A1[102] , \A1[101] , \A1[100] , \A1[99] ,
         \A1[98] , \A1[97] , \A1[96] , \A1[95] , \A1[94] , \A1[93] , \A1[92] ,
         \A1[91] , \A1[90] , \A1[89] , \A1[88] , \A1[87] , \A1[86] , \A1[85] ,
         \A1[84] , \A1[83] , \A1[82] , \A1[81] , \A1[80] , \A1[79] , \A1[78] ,
         \A1[77] , \A1[76] , \A1[75] , \A1[74] , \A1[73] , \A1[72] , \A1[71] ,
         \A1[70] , \A1[69] , \A1[68] , \A1[67] , \A1[66] , \A1[65] , \A1[64] ,
         \A1[63] , \A1[62] , \A1[61] , \A1[60] , \A1[59] , \A1[58] , \A1[57] ,
         \A1[56] , \A1[55] , \A1[54] , \A1[53] , \A1[52] , \A1[51] , \A1[50] ,
         \A1[49] , \A1[48] , \A1[47] , \A1[46] , \A1[45] , \A1[44] , \A1[43] ,
         \A1[42] , \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] ,
         \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] ,
         \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] ,
         \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] ,
         \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] ,
         \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] ,
         \A1[0] , \A2[285] , \A2[284] , \A2[283] , \A2[282] , \A2[281] ,
         \A2[280] , \A2[279] , \A2[278] , \A2[277] , \A2[276] , \A2[275] ,
         \A2[274] , \A2[273] , \A2[272] , \A2[271] , \A2[270] , \A2[269] ,
         \A2[268] , \A2[267] , \A2[266] , \A2[265] , \A2[264] , \A2[263] ,
         \A2[262] , \A2[261] , \A2[260] , \A2[259] , \A2[258] , \A2[257] ,
         \A2[256] , \A2[255] , \A2[254] , \A2[253] , \A2[252] , \A2[251] ,
         \A2[250] , \A2[249] , \A2[248] , \A2[247] , \A2[246] , \A2[245] ,
         \A2[244] , \A2[243] , \A2[242] , \A2[241] , \A2[240] , \A2[239] ,
         \A2[238] , \A2[237] , \A2[236] , \A2[235] , \A2[234] , \A2[233] ,
         \A2[232] , \A2[231] , \A2[230] , \A2[229] , \A2[228] , \A2[227] ,
         \A2[226] , \A2[225] , \A2[224] , \A2[223] , \A2[222] , \A2[221] ,
         \A2[220] , \A2[219] , \A2[218] , \A2[217] , \A2[216] , \A2[215] ,
         \A2[214] , \A2[213] , \A2[212] , \A2[211] , \A2[210] , \A2[209] ,
         \A2[208] , \A2[207] , \A2[206] , \A2[205] , \A2[204] , \A2[203] ,
         \A2[202] , \A2[201] , \A2[200] , \A2[199] , \A2[198] , \A2[197] ,
         \A2[196] , \A2[195] , \A2[194] , \A2[193] , \A2[192] , \A2[191] ,
         \A2[190] , \A2[189] , \A2[188] , \A2[187] , \A2[186] , \A2[185] ,
         \A2[184] , \A2[183] , \A2[182] , \A2[181] , \A2[180] , \A2[179] ,
         \A2[178] , \A2[177] , \A2[176] , \A2[175] , \A2[174] , \A2[173] ,
         \A2[172] , \A2[171] , \A2[170] , \A2[169] , \A2[168] , \A2[167] ,
         \A2[166] , \A2[165] , \A2[164] , \A2[163] , \A2[162] , \A2[161] ,
         \A2[160] , \A2[159] , \A2[158] , \A2[157] , \A2[156] , \A2[155] ,
         \A2[154] , \A2[153] , \A2[152] , \A2[151] , \A2[150] , \A2[149] ,
         \A2[148] , \A2[147] , \A2[146] , \A2[145] , \A2[144] , \A2[143] ,
         \A2[142] , \A2[141] , \A2[140] , \A2[139] , \A2[138] , \A2[137] ,
         \A2[136] , \A2[135] , \A2[134] , \A2[133] , \A2[132] , \A2[131] ,
         \A2[130] , \A2[129] , \A2[128] , \A2[127] , \A2[126] , \A2[125] ,
         \A2[124] , \A2[123] , \A2[122] , \A2[121] , \A2[120] , \A2[119] ,
         \A2[118] , \A2[117] , \A2[116] , \A2[115] , \A2[114] , \A2[113] ,
         \A2[112] , \A2[111] , \A2[110] , \A2[109] , \A2[108] , \A2[107] ,
         \A2[106] , \A2[105] , \A2[104] , \A2[103] , \A2[102] , \A2[101] ,
         \A2[100] , \A2[99] , \A2[98] , \A2[97] , \A2[96] , \A2[95] , \A2[94] ,
         \A2[93] , \A2[92] , \A2[91] , \A2[90] , \A2[89] , \A2[88] , \A2[87] ,
         \A2[86] , \A2[85] , \A2[84] , \A2[83] , \A2[82] , \A2[81] , \A2[80] ,
         \A2[79] , \A2[78] , \A2[77] , \A2[76] , \A2[75] , \A2[74] , \A2[73] ,
         \A2[72] , \A2[71] , \A2[70] , \A2[69] , \A2[68] , \A2[67] , \A2[66] ,
         \A2[65] , \A2[64] , \A2[63] , \A2[62] , \A2[61] , \A2[60] , \A2[59] ,
         \A2[58] , \A2[57] , \A2[56] , \A2[55] , \A2[54] , \A2[53] , \A2[52] ,
         \A2[51] , \A2[50] , \A2[49] , \A2[48] , \A2[47] , \A2[46] , \A2[45] ,
         \A2[44] , \A2[43] , \A2[42] , \A2[41] , \A2[40] , \A2[39] , \A2[38] ,
         \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] , \A2[32] , \A2[31] ,
         n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043,
         n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053,
         n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063,
         n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073,
         n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083,
         n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093,
         n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103,
         n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113,
         n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122, n1123,
         n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132, n1133,
         n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142, n1143,
         n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152, n1153,
         n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162, n1163,
         n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172, n1173,
         n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182, n1183,
         n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192, n1193,
         n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202, n1203,
         n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212, n1213,
         n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222, n1223,
         n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232, n1233,
         n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242, n1243,
         n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252, n1253,
         n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262, n1263,
         n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272, n1273,
         n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282, n1283,
         n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292, n1293,
         n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302, n1303,
         n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312, n1313,
         n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322, n1323,
         n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332, n1333,
         n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342, n1343,
         n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352, n1353,
         n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362, n1363,
         n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372, n1373,
         n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382, n1383,
         n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392, n1393,
         n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402, n1403,
         n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412, n1413,
         n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422, n1423,
         n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432, n1433,
         n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442, n1443,
         n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452, n1453,
         n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462, n1463,
         n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472, n1473,
         n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482, n1483,
         n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492, n1493,
         n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502, n1503,
         n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512, n1513,
         n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522, n1523,
         n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532, n1533,
         n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542, n1543,
         n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552, n1553,
         n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562, n1563,
         n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572, n1573,
         n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582, n1583,
         n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592, n1593,
         n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602, n1603,
         n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612, n1613,
         n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622, n1623,
         n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632, n1633,
         n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642, n1643,
         n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652, n1653,
         n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662, n1663,
         n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672, n1673,
         n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682, n1683,
         n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692, n1693,
         n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702, n1703,
         n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712, n1713,
         n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722, n1723,
         n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732, n1733,
         n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742, n1743,
         n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752, n1753,
         n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762, n1763,
         n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772, n1773,
         n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782, n1783,
         n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792, n1793,
         n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802, n1803,
         n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812, n1813,
         n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822, n1823,
         n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832, n1833,
         n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842, n1843,
         n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852, n1853,
         n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862, n1863,
         n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872, n1873,
         n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882, n1883,
         n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892, n1893,
         n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902, n1903,
         n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912, n1913,
         n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922, n1923,
         n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932, n1933,
         n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942, n1943,
         n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952, n1953,
         n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962, n1963,
         n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972, n1973,
         n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982, n1983,
         n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992, n1993,
         n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002, n2003,
         n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012, n2013,
         n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022, n2023,
         n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032, n2033,
         n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042, n2043,
         n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052, n2053,
         n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062, n2063,
         n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072, n2073,
         n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082, n2083,
         n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092, n2093,
         n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102, n2103,
         n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112, n2113,
         n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122, n2123,
         n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132, n2133,
         n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142, n2143,
         n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152, n2153,
         n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162, n2163,
         n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172, n2173,
         n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182, n2183,
         n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192, n2193,
         n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202, n2203,
         n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212, n2213,
         n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222, n2223,
         n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232, n2233,
         n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242, n2243,
         n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252, n2253,
         n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262, n2263,
         n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272, n2273,
         n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282, n2283,
         n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292, n2293,
         n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302, n2303,
         n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312, n2313,
         n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322, n2323,
         n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332, n2333,
         n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342, n2343,
         n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352, n2353,
         n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362, n2363,
         n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372, n2373,
         n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382, n2383,
         n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392, n2393,
         n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402, n2403,
         n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412, n2413,
         n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422, n2423,
         n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432, n2433,
         n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442, n2443,
         n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452, n2453,
         n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462, n2463,
         n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472, n2473,
         n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482, n2483,
         n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492, n2493,
         n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502, n2503,
         n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512, n2513,
         n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522, n2523,
         n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532, n2533,
         n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542, n2543,
         n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552, n2553,
         n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562, n2563,
         n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572, n2573,
         n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582, n2583,
         n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592, n2593,
         n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602, n2603,
         n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612, n2613,
         n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622, n2623,
         n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632, n2633,
         n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642, n2643,
         n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652, n2653,
         n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662, n2663,
         n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672, n2673,
         n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682, n2683,
         n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692, n2693,
         n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702, n2703,
         n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712, n2713,
         n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722, n2723,
         n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732, n2733,
         n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742, n2743,
         n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752, n2753,
         n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762, n2763,
         n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772, n2773,
         n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782, n2783,
         n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792, n2793,
         n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802, n2803,
         n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812, n2813,
         n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822, n2823,
         n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832, n2833,
         n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842, n2843,
         n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852, n2853,
         n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862, n2863,
         n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872, n2873,
         n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882, n2883,
         n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892, n2893,
         n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902, n2903,
         n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912, n2913,
         n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922, n2923,
         n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932, n2933,
         n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942, n2943,
         n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952, n2953,
         n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962, n2963,
         n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972, n2973,
         n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982, n2983,
         n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992, n2993,
         n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002, n3003,
         n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012, n3013,
         n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022, n3023,
         n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032, n3033,
         n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042, n3043,
         n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052, n3053,
         n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062, n3063,
         n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072, n3073,
         n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082, n3083,
         n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092, n3093,
         n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102, n3103,
         n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112, n3113,
         n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122, n3123,
         n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132, n3133,
         n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142, n3143,
         n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152, n3153,
         n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162, n3163,
         n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172, n3173,
         n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182, n3183,
         n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192, n3193,
         n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202, n3203,
         n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212, n3213,
         n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222, n3223,
         n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232, n3233,
         n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242, n3243,
         n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252, n3253,
         n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262, n3263,
         n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272, n3273,
         n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282, n3283,
         n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292, n3293,
         n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302, n3303,
         n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312, n3313,
         n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322, n3323,
         n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332, n3333,
         n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342, n3343,
         n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352, n3353,
         n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362, n3363,
         n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372, n3373,
         n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382, n3383,
         n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392, n3393,
         n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402, n3403,
         n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412, n3413,
         n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422, n3423,
         n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432, n3433,
         n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442, n3443,
         n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452, n3453,
         n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462, n3463,
         n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472, n3473,
         n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482, n3483,
         n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492, n3493,
         n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502, n3503,
         n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512, n3513,
         n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522, n3523,
         n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532, n3533,
         n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542, n3543,
         n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552, n3553,
         n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562, n3563,
         n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572, n3573,
         n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582, n3583,
         n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592, n3593,
         n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602, n3603,
         n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612, n3613,
         n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622, n3623,
         n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632, n3633,
         n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642, n3643,
         n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652, n3653,
         n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662, n3663,
         n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672, n3673,
         n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682, n3683,
         n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692, n3693,
         n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702, n3703,
         n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712, n3713,
         n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722, n3723,
         n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732, n3733,
         n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742, n3743,
         n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752, n3753,
         n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762, n3763,
         n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772, n3773,
         n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782, n3783,
         n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792, n3793,
         n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802, n3803,
         n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812, n3813,
         n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822, n3823,
         n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832, n3833,
         n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842, n3843,
         n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852, n3853,
         n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862, n3863,
         n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872, n3873,
         n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882, n3883,
         n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892, n3893,
         n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902, n3903,
         n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912, n3913,
         n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922, n3923,
         n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932, n3933,
         n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942, n3943,
         n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952, n3953,
         n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962, n3963,
         n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972, n3973,
         n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982, n3983,
         n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992, n3993,
         n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002, n4003,
         n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012, n4013,
         n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022, n4023,
         n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032, n4033,
         n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042, n4043,
         n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052, n4053,
         n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062, n4063,
         n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072, n4073,
         n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082, n4083,
         n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092, n4093,
         n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102, n4103,
         n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112, n4113,
         n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122, n4123,
         n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132, n4133,
         n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142, n4143,
         n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152, n4153,
         n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162, n4163,
         n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172, n4173,
         n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182, n4183,
         n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192, n4193,
         n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202, n4203,
         n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212, n4213,
         n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222, n4223,
         n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232, n4233,
         n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242, n4243,
         n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252, n4253,
         n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262, n4263,
         n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272, n4273,
         n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282, n4283,
         n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292, n4293,
         n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302, n4303,
         n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312, n4313,
         n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322, n4323,
         n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332, n4333,
         n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342, n4343,
         n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352, n4353,
         n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362, n4363,
         n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372, n4373,
         n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382, n4383,
         n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392, n4393,
         n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402, n4403,
         n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412, n4413,
         n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422, n4423,
         n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432, n4433,
         n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442, n4443,
         n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452, n4453,
         n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462, n4463,
         n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472, n4473,
         n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482, n4483,
         n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492, n4493,
         n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502, n4503,
         n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512, n4513,
         n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522, n4523,
         n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532, n4533,
         n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542, n4543,
         n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552, n4553,
         n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562, n4563,
         n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572, n4573,
         n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582, n4583,
         n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592, n4593,
         n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602, n4603,
         n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612, n4613,
         n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622, n4623,
         n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632, n4633,
         n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642, n4643,
         n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652, n4653,
         n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662, n4663,
         n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672, n4673,
         n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682, n4683,
         n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692, n4693,
         n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702, n4703,
         n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712, n4713,
         n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722, n4723,
         n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732, n4733,
         n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742, n4743,
         n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752, n4753,
         n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762, n4763,
         n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772, n4773,
         n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782, n4783,
         n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792, n4793,
         n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802, n4803,
         n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812, n4813,
         n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822, n4823,
         n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832, n4833,
         n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842, n4843,
         n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852, n4853,
         n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862, n4863,
         n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872, n4873,
         n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882, n4883,
         n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892, n4893,
         n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902, n4903,
         n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912, n4913,
         n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922, n4923,
         n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932, n4933,
         n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942, n4943,
         n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952, n4953,
         n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962, n4963,
         n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972, n4973,
         n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982, n4983,
         n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992, n4993,
         n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002, n5003,
         n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012, n5013,
         n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022, n5023,
         n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032, n5033,
         n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042, n5043,
         n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052, n5053,
         n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062, n5063,
         n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072, n5073,
         n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082, n5083,
         n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092, n5093,
         n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102, n5103,
         n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112, n5113,
         n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122, n5123,
         n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132, n5133,
         n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142, n5143,
         n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152, n5153,
         n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162, n5163,
         n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172, n5173,
         n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182, n5183,
         n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192, n5193,
         n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202, n5203,
         n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212, n5213,
         n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222, n5223,
         n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232, n5233,
         n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242, n5243,
         n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252, n5253,
         n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262, n5263,
         n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272, n5273,
         n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282, n5283,
         n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292, n5293,
         n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302, n5303,
         n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312, n5313,
         n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322, n5323,
         n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332, n5333,
         n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342, n5343,
         n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352, n5353,
         n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362, n5363,
         n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372, n5373,
         n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382, n5383,
         n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392, n5393,
         n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402, n5403,
         n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412, n5413,
         n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422, n5423,
         n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432, n5433,
         n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442, n5443,
         n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452, n5453,
         n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462, n5463,
         n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472, n5473,
         n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482, n5483,
         n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492, n5493,
         n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502, n5503,
         n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512, n5513,
         n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522, n5523,
         n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532, n5533,
         n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542, n5543,
         n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552, n5553,
         n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562, n5563,
         n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572, n5573,
         n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582, n5583,
         n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592, n5593,
         n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602, n5603,
         n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612, n5613,
         n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622, n5623,
         n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632, n5633,
         n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642, n5643,
         n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652, n5653,
         n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662, n5663,
         n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672, n5673,
         n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682, n5683,
         n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692, n5693,
         n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702, n5703,
         n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712, n5713,
         n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722, n5723,
         n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732, n5733,
         n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742, n5743,
         n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752, n5753,
         n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762, n5763,
         n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772, n5773,
         n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782, n5783,
         n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792, n5793,
         n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802, n5803,
         n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812, n5813,
         n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822, n5823,
         n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832, n5833,
         n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842, n5843,
         n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852, n5853,
         n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862, n5863,
         n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872, n5873,
         n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882, n5883,
         n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892, n5893,
         n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902, n5903,
         n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912, n5913,
         n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922, n5923,
         n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932, n5933,
         n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942, n5943,
         n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952, n5953,
         n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962, n5963,
         n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972, n5973,
         n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982, n5983,
         n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992, n5993,
         n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002, n6003,
         n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012, n6013,
         n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022, n6023,
         n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032, n6033,
         n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042, n6043,
         n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052, n6053,
         n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062, n6063,
         n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072, n6073,
         n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082, n6083,
         n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092, n6093,
         n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102, n6103,
         n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112, n6113,
         n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122, n6123,
         n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132, n6133,
         n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142, n6143,
         n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152, n6153,
         n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162, n6163,
         n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172, n6173,
         n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182, n6183,
         n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192, n6193,
         n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202, n6203,
         n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212, n6213,
         n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222, n6223,
         n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232, n6233,
         n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242, n6243,
         n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252, n6253,
         n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262, n6263,
         n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272, n6273,
         n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282, n6283,
         n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292, n6293,
         n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302, n6303,
         n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312, n6313,
         n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322, n6323,
         n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332, n6333,
         n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342, n6343,
         n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352, n6353,
         n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362, n6363,
         n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372, n6373,
         n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382, n6383,
         n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392, n6393,
         n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402, n6403,
         n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412, n6413,
         n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422, n6423,
         n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432, n6433,
         n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442, n6443,
         n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452, n6453,
         n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462, n6463,
         n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472, n6473,
         n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482, n6483,
         n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492, n6493,
         n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502, n6503,
         n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512, n6513,
         n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522, n6523,
         n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532, n6533,
         n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542, n6543,
         n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552, n6553,
         n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562, n6563,
         n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572, n6573,
         n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582, n6583,
         n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592, n6593,
         n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602, n6603,
         n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612, n6613,
         n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622, n6623,
         n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632, n6633,
         n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642, n6643,
         n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652, n6653,
         n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662, n6663,
         n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672, n6673,
         n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682, n6683,
         n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692, n6693,
         n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702, n6703,
         n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712, n6713,
         n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722, n6723,
         n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732, n6733,
         n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742, n6743,
         n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752, n6753,
         n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762, n6763,
         n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772, n6773,
         n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782, n6783,
         n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792, n6793,
         n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802, n6803,
         n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812, n6813,
         n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822, n6823,
         n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832, n6833,
         n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842, n6843,
         n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852, n6853,
         n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862, n6863,
         n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872, n6873,
         n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882, n6883,
         n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892, n6893,
         n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902, n6903,
         n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912, n6913,
         n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922, n6923,
         n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932, n6933,
         n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942, n6943,
         n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952, n6953,
         n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962, n6963,
         n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972, n6973,
         n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982, n6983,
         n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992, n6993,
         n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002, n7003,
         n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012, n7013,
         n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022, n7023,
         n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032, n7033,
         n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042, n7043,
         n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052, n7053,
         n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062, n7063,
         n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072, n7073,
         n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082, n7083,
         n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092, n7093,
         n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102, n7103,
         n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112, n7113,
         n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122, n7123,
         n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132, n7133,
         n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142, n7143,
         n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152, n7153,
         n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162, n7163,
         n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172, n7173,
         n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182, n7183,
         n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192, n7193,
         n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202, n7203,
         n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212, n7213,
         n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222, n7223,
         n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232, n7233,
         n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242, n7243,
         n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252, n7253,
         n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262, n7263,
         n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272, n7273,
         n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282, n7283,
         n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292, n7293,
         n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302, n7303,
         n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312, n7313,
         n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322, n7323,
         n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332, n7333,
         n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342, n7343,
         n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352, n7353,
         n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362, n7363,
         n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372, n7373,
         n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382, n7383,
         n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392, n7393,
         n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402, n7403,
         n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412, n7413,
         n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422, n7423,
         n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432, n7433,
         n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442, n7443,
         n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452, n7453,
         n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462, n7463,
         n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472, n7473,
         n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482, n7483,
         n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492, n7493,
         n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502, n7503,
         n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512, n7513,
         n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522, n7523,
         n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532, n7533,
         n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542, n7543,
         n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552, n7553,
         n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562, n7563,
         n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572, n7573,
         n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582, n7583,
         n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592, n7593,
         n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602, n7603,
         n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612, n7613,
         n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622, n7623,
         n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632, n7633,
         n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642, n7643,
         n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652, n7653,
         n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662, n7663,
         n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672, n7673,
         n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682, n7683,
         n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692, n7693,
         n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702, n7703,
         n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712, n7713,
         n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722, n7723,
         n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732, n7733,
         n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742, n7743,
         n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752, n7753,
         n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762, n7763,
         n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772, n7773,
         n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782, n7783,
         n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792, n7793,
         n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802, n7803,
         n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812, n7813,
         n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822, n7823,
         n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832, n7833,
         n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842, n7843,
         n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852, n7853,
         n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862, n7863,
         n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872, n7873,
         n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882, n7883,
         n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892, n7893,
         n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902, n7903,
         n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912, n7913,
         n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922, n7923,
         n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932, n7933,
         n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942, n7943,
         n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952, n7953,
         n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962, n7963,
         n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972, n7973,
         n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982, n7983,
         n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992, n7993,
         n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002, n8003,
         n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012, n8013,
         n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022, n8023,
         n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032, n8033,
         n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042, n8043,
         n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052, n8053,
         n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062, n8063,
         n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072, n8073,
         n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082, n8083,
         n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092, n8093,
         n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102, n8103,
         n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112, n8113,
         n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122, n8123,
         n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132, n8133,
         n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142, n8143,
         n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152, n8153,
         n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162, n8163,
         n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172, n8173,
         n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182, n8183,
         n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192, n8193,
         n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202, n8203,
         n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212, n8213,
         n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222, n8223,
         n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232, n8233,
         n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242, n8243,
         n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252, n8253,
         n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262, n8263,
         n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272, n8273,
         n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282, n8283,
         n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292, n8293,
         n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302, n8303,
         n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312, n8313,
         n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322, n8323,
         n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332, n8333,
         n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342, n8343,
         n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352, n8353,
         n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362, n8363,
         n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372, n8373,
         n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382, n8383,
         n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392, n8393,
         n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402, n8403,
         n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412, n8413,
         n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422, n8423,
         n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432, n8433,
         n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442, n8443,
         n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452, n8453,
         n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462, n8463,
         n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472, n8473,
         n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482, n8483,
         n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492, n8493,
         n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502, n8503,
         n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512, n8513,
         n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522, n8523,
         n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532, n8533,
         n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542, n8543,
         n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552, n8553,
         n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562, n8563,
         n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572, n8573,
         n8574, n8575, n8576, n8577, n8578, n8579, n8580, n8581, n8582, n8583,
         n8584, n8585, n8586, n8587, n8588, n8589, n8590, n8591, n8592, n8593,
         n8594, n8595, n8596, n8597, n8598, n8599, n8600, n8601, n8602, n8603,
         n8604, n8605, n8606, n8607, n8608, n8609, n8610, n8611, n8612, n8613,
         n8614, n8615, n8616, n8617, n8618, n8619, n8620, n8621, n8622, n8623,
         n8624, n8625, n8626, n8627, n8628, n8629, n8630, n8631, n8632, n8633,
         n8634, n8635, n8636, n8637, n8638, n8639, n8640, n8641, n8642, n8643,
         n8644, n8645, n8646, n8647, n8648, n8649, n8650, n8651, n8652, n8653,
         n8654, n8655, n8656, n8657, n8658, n8659, n8660, n8661, n8662, n8663,
         n8664, n8665, n8666, n8667, n8668, n8669, n8670, n8671, n8672, n8673,
         n8674, n8675, n8676, n8677, n8678, n8679, n8680, n8681, n8682, n8683,
         n8684, n8685, n8686, n8687, n8688, n8689, n8690, n8691, n8692, n8693,
         n8694, n8695, n8696, n8697, n8698, n8699, n8700, n8701, n8702, n8703,
         n8704, n8705, n8706, n8707, n8708, n8709, n8710, n8711, n8712, n8713,
         n8714, n8715, n8716, n8717, n8718, n8719, n8720, n8721, n8722, n8723,
         n8724, n8725, n8726, n8727, n8728, n8729, n8730, n8731, n8732, n8733,
         n8734, n8735, n8736, n8737, n8738, n8739, n8740, n8741, n8742, n8743,
         n8744, n8745, n8746, n8747, n8748, n8749, n8750, n8751, n8752, n8753,
         n8754, n8755, n8756, n8757, n8758, n8759, n8760, n8761, n8762, n8763,
         n8764, n8765, n8766, n8767, n8768, n8769, n8770, n8771, n8772, n8773,
         n8774, n8775, n8776, n8777, n8778, n8779, n8780, n8781, n8782, n8783,
         n8784, n8785, n8786, n8787, n8788, n8789, n8790, n8791, n8792, n8793,
         n8794, n8795, n8796, n8797, n8798, n8799, n8800, n8801, n8802, n8803,
         n8804, n8805, n8806, n8807, n8808, n8809, n8810, n8811, n8812, n8813,
         n8814, n8815, n8816, n8817, n8818, n8819, n8820, n8821, n8822, n8823,
         n8824, n8825, n8826, n8827, n8828, n8829, n8830, n8831, n8832, n8833,
         n8834, n8835, n8836, n8837, n8838, n8839, n8840, n8841, n8842, n8843,
         n8844, n8845, n8846, n8847, n8848, n8849, n8850, n8851, n8852, n8853,
         n8854, n8855, n8856, n8857, n8858, n8859, n8860, n8861, n8862, n8863,
         n8864, n8865, n8866, n8867, n8868, n8869, n8870, n8871, n8872, n8873,
         n8874, n8875, n8876, n8877, n8878, n8879, n8880, n8881, n8882, n8883,
         n8884, n8885, n8886, n8887, n8888, n8889, n8890, n8891, n8892, n8893,
         n8894, n8895, n8896, n8897, n8898, n8899, n8900, n8901, n8902, n8903,
         n8904, n8905, n8906, n8907, n8908, n8909, n8910, n8911, n8912, n8913,
         n8914, n8915, n8916, n8917, n8918, n8919, n8920, n8921, n8922, n8923,
         n8924, n8925, n8926, n8927, n8928, n8929, n8930, n8931, n8932, n8933,
         n8934, n8935, n8936, n8937, n8938, n8939, n8940, n8941, n8942, n8943,
         n8944, n8945, n8946, n8947, n8948, n8949, n8950, n8951, n8952, n8953,
         n8954, n8955, n8956, n8957, n8958, n8959, n8960, n8961, n8962, n8963,
         n8964, n8965, n8966, n8967, n8968, n8969, n8970, n8971, n8972, n8973,
         n8974, n8975, n8976, n8977, n8978, n8979, n8980, n8981, n8982, n8983,
         n8984, n8985, n8986, n8987, n8988, n8989, n8990, n8991, n8992, n8993,
         n8994, n8995, n8996, n8997, n8998, n8999, n9000, n9001, n9002, n9003,
         n9004, n9005, n9006, n9007, n9008, n9009, n9010, n9011, n9012, n9013,
         n9014, n9015, n9016, n9017, n9018, n9019, n9020, n9021, n9022, n9023,
         n9024, n9025, n9026, n9027, n9028, n9029, n9030, n9031, n9032, n9033,
         n9034, n9035, n9036, n9037, n9038, n9039, n9040, n9041, n9042, n9043,
         n9044, n9045, n9046, n9047, n9048, n9049, n9050, n9051, n9052, n9053,
         n9054, n9055, n9056, n9057, n9058, n9059, n9060, n9061, n9062, n9063,
         n9064, n9065, n9066, n9067, n9068, n9069, n9070, n9071, n9072, n9073,
         n9074, n9075, n9076, n9077, n9078, n9079, n9080, n9081, n9082, n9083,
         n9084, n9085, n9086, n9087, n9088, n9089, n9090, n9091, n9092, n9093,
         n9094, n9095, n9096, n9097, n9098, n9099, n9100, n9101, n9102, n9103,
         n9104, n9105, n9106, n9107, n9108, n9109, n9110, n9111, n9112, n9113,
         n9114, n9115, n9116, n9117, n9118, n9119, n9120, n9121, n9122, n9123,
         n9124, n9125, n9126, n9127, n9128, n9129, n9130, n9131, n9132, n9133,
         n9134, n9135, n9136, n9137, n9138, n9139, n9140, n9141, n9142, n9143,
         n9144, n9145, n9146, n9147, n9148, n9149, n9150, n9151, n9152, n9153,
         n9154, n9155, n9156, n9157, n9158, n9159, n9160, n9161, n9162, n9163,
         n9164, n9165, n9166, n9167, n9168, n9169, n9170, n9171, n9172, n9173,
         n9174, n9175, n9176, n9177, n9178, n9179, n9180, n9181, n9182, n9183,
         n9184, n9185, n9186, n9187, n9188, n9189, n9190, n9191, n9192, n9193,
         n9194, n9195, n9196, n9197, n9198, n9199, n9200, n9201, n9202, n9203,
         n9204, n9205, n9206, n9207, n9208, n9209, n9210, n9211, n9212, n9213,
         n9214, n9215, n9216, n9217, n9218, n9219, n9220, n9221, n9222, n9223,
         n9224, n9225, n9226, n9227, n9228, n9229, n9230, n9231, n9232, n9233,
         n9234, n9235, n9236, n9237, n9238, n9239, n9240, n9241, n9242, n9243,
         n9244, n9245, n9246, n9247, n9248, n9249, n9250, n9251, n9252, n9253,
         n9254, n9255, n9256, n9257, n9258, n9259, n9260, n9261, n9262, n9263,
         n9264, n9265, n9266, n9267, n9268, n9269, n9270, n9271, n9272, n9273,
         n9274, n9275, n9276, n9277, n9278, n9279, n9280, n9281, n9282, n9283,
         n9284, n9285, n9286, n9287, n9288, n9289, n9290, n9291, n9292, n9293,
         n9294, n9295, n9296, n9297, n9298, n9299, n9300, n9301, n9302, n9303,
         n9304, n9305, n9306, n9307, n9308, n9309, n9310, n9311, n9312, n9313,
         n9314, n9315, n9316, n9317, n9318, n9319, n9320, n9321, n9322, n9323,
         n9324, n9325, n9326, n9327, n9328, n9329, n9330, n9331, n9332, n9333,
         n9334, n9335, n9336, n9337, n9338, n9339, n9340, n9341, n9342, n9343,
         n9344, n9345, n9346, n9347, n9348, n9349, n9350, n9351, n9352, n9353,
         n9354, n9355, n9356, n9357, n9358, n9359, n9360, n9361, n9362, n9363,
         n9364, n9365, n9366, n9367, n9368, n9369, n9370, n9371, n9372, n9373,
         n9374, n9375, n9376, n9377, n9378, n9379, n9380, n9381, n9382, n9383,
         n9384, n9385, n9386, n9387, n9388, n9389, n9390, n9391, n9392, n9393,
         n9394, n9395, n9396, n9397, n9398, n9399, n9400, n9401, n9402, n9403,
         n9404, n9405, n9406, n9407, n9408, n9409, n9410, n9411, n9412, n9413,
         n9414, n9415, n9416, n9417, n9418, n9419, n9420, n9421, n9422, n9423,
         n9424, n9425, n9426, n9427, n9428, n9429, n9430, n9431, n9432, n9433,
         n9434, n9435, n9436, n9437, n9438, n9439, n9440, n9441, n9442, n9443,
         n9444, n9445, n9446, n9447, n9448, n9449, n9450, n9451, n9452, n9453,
         n9454, n9455, n9456, n9457, n9458, n9459, n9460, n9461, n9462, n9463,
         n9464, n9465, n9466, n9467, n9468, n9469, n9470, n9471, n9472, n9473,
         n9474, n9475, n9476, n9477, n9478, n9479, n9480, n9481, n9482, n9483,
         n9484, n9485, n9486, n9487, n9488, n9489, n9490, n9491, n9492, n9493,
         n9494, n9495, n9496, n9497, n9498, n9499, n9500, n9501, n9502, n9503,
         n9504, n9505, n9506, n9507, n9508, n9509, n9510, n9511, n9512, n9513,
         n9514, n9515, n9516, n9517, n9518, n9519, n9520, n9521, n9522, n9523,
         n9524, n9525, n9526, n9527, n9528, n9529, n9530, n9531, n9532, n9533,
         n9534, n9535, n9536, n9537, n9538, n9539, n9540, n9541, n9542, n9543,
         n9544, n9545, n9546, n9547, n9548, n9549, n9550, n9551, n9552, n9553,
         n9554, n9555, n9556, n9557, n9558, n9559, n9560, n9561, n9562, n9563,
         n9564, n9565, n9566, n9567, n9568, n9569, n9570, n9571, n9572, n9573,
         n9574, n9575, n9576, n9577, n9578, n9579, n9580, n9581, n9582, n9583,
         n9584, n9585, n9586, n9587, n9588, n9589, n9590, n9591, n9592, n9593,
         n9594, n9595, n9596, n9597, n9598, n9599, n9600, n9601, n9602, n9603,
         n9604, n9605, n9606, n9607, n9608, n9609, n9610, n9611, n9612, n9613,
         n9614, n9615, n9616, n9617, n9618, n9619, n9620, n9621, n9622, n9623,
         n9624, n9625, n9626, n9627, n9628, n9629, n9630, n9631, n9632, n9633,
         n9634, n9635, n9636, n9637, n9638, n9639, n9640, n9641, n9642, n9643,
         n9644, n9645, n9646, n9647, n9648, n9649, n9650, n9651, n9652, n9653,
         n9654, n9655, n9656, n9657, n9658, n9659, n9660, n9661, n9662, n9663,
         n9664, n9665, n9666, n9667, n9668, n9669, n9670, n9671, n9672, n9673,
         n9674, n9675, n9676, n9677, n9678, n9679, n9680, n9681, n9682, n9683,
         n9684, n9685, n9686, n9687, n9688, n9689, n9690, n9691, n9692, n9693,
         n9694, n9695, n9696, n9697, n9698, n9699, n9700, n9701, n9702, n9703,
         n9704, n9705, n9706, n9707, n9708, n9709, n9710, n9711, n9712, n9713,
         n9714, n9715, n9716, n9717, n9718, n9719, n9720, n9721, n9722, n9723,
         n9724, n9725, n9726, n9727, n9728, n9729, n9730, n9731, n9732, n9733,
         n9734, n9735, n9736, n9737, n9738, n9739, n9740, n9741, n9742, n9743,
         n9744, n9745, n9746, n9747, n9748, n9749, n9750, n9751, n9752, n9753,
         n9754, n9755, n9756, n9757, n9758, n9759, n9760, n9761, n9762, n9763,
         n9764, n9765, n9766, n9767, n9768, n9769, n9770, n9771, n9772, n9773,
         n9774, n9775, n9776, n9777, n9778, n9779, n9780, n9781, n9782, n9783,
         n9784, n9785, n9786, n9787, n9788, n9789, n9790, n9791, n9792, n9793,
         n9794, n9795, n9796, n9797, n9798, n9799, n9800, n9801, n9802, n9803,
         n9804, n9805, n9806, n9807, n9808, n9809, n9810, n9811, n9812, n9813,
         n9814, n9815, n9816, n9817, n9818, n9819, n9820, n9821, n9822, n9823,
         n9824, n9825, n9826, n9827, n9828, n9829, n9830, n9831, n9832, n9833,
         n9834, n9835, n9836, n9837, n9838, n9839, n9840, n9841, n9842, n9843,
         n9844, n9845, n9846, n9847, n9848, n9849, n9850, n9851, n9852, n9853,
         n9854, n9855, n9856, n9857, n9858, n9859, n9860, n9861, n9862, n9863,
         n9864, n9865, n9866, n9867, n9868, n9869, n9870, n9871, n9872, n9873,
         n9874, n9875, n9876, n9877, n9878, n9879, n9880, n9881, n9882, n9883,
         n9884, n9885, n9886, n9887, n9888, n9889, n9890, n9891, n9892, n9893,
         n9894, n9895, n9896, n9897, n9898, n9899, n9900, n9901, n9902, n9903,
         n9904, n9905, n9906, n9907, n9908, n9909, n9910, n9911, n9912, n9913,
         n9914, n9915, n9916, n9917, n9918, n9919, n9920, n9921, n9922, n9923,
         n9924, n9925, n9926, n9927, n9928, n9929, n9930, n9931, n9932, n9933,
         n9934, n9935, n9936, n9937, n9938, n9939, n9940, n9941, n9942, n9943,
         n9944, n9945, n9946, n9947, n9948, n9949, n9950, n9951, n9952, n9953,
         n9954, n9955, n9956, n9957, n9958, n9959, n9960, n9961, n9962, n9963,
         n9964, n9965, n9966, n9967, n9968, n9969, n9970, n9971, n9972, n9973,
         n9974, n9975, n9976, n9977, n9978, n9979, n9980, n9981, n9982, n9983,
         n9984, n9985, n9986, n9987, n9988, n9989, n9990, n9991, n9992, n9993,
         n9994, n9995, n9996, n9997, n9998, n9999, n10000, n10001, n10002,
         n10003, n10004, n10005, n10006, n10007, n10008, n10009, n10010,
         n10011, n10012, n10013, n10014, n10015, n10016, n10017, n10018,
         n10019, n10020, n10021, n10022, n10023, n10024, n10025, n10026,
         n10027, n10028, n10029, n10030, n10031, n10032, n10033, n10034,
         n10035, n10036, n10037, n10038, n10039, n10040, n10041, n10042,
         n10043, n10044, n10045, n10046, n10047, n10048, n10049, n10050,
         n10051, n10052, n10053, n10054, n10055, n10056, n10057, n10058,
         n10059, n10060, n10061, n10062, n10063, n10064, n10065, n10066,
         n10067, n10068, n10069, n10070, n10071, n10072, n10073, n10074,
         n10075, n10076, n10077, n10078, n10079, n10080, n10081, n10082,
         n10083, n10084, n10085, n10086, n10087, n10088, n10089, n10090,
         n10091, n10092, n10093, n10094, n10095, n10096, n10097, n10098,
         n10099, n10100, n10101, n10102, n10103, n10104, n10105, n10106,
         n10107, n10108, n10109, n10110, n10111, n10112, n10113, n10114,
         n10115, n10116, n10117, n10118, n10119, n10120, n10121, n10122,
         n10123, n10124, n10125, n10126, n10127, n10128, n10129, n10130,
         n10131, n10132, n10133, n10134, n10135, n10136, n10137, n10138,
         n10139, n10140, n10141, n10142, n10143, n10144, n10145, n10146,
         n10147, n10148, n10149, n10150, n10151, n10152, n10153, n10154,
         n10155, n10156, n10157, n10158, n10159, n10160, n10161, n10162,
         n10163, n10164, n10165, n10166, n10167, n10168, n10169, n10170,
         n10171, n10172, n10173, n10174, n10175, n10176, n10177, n10178,
         n10179, n10180, n10181, n10182, n10183, n10184, n10185, n10186,
         n10187, n10188, n10189, n10190, n10191, n10192, n10193, n10194,
         n10195, n10196, n10197, n10198, n10199, n10200, n10201, n10202,
         n10203, n10204, n10205, n10206, n10207, n10208, n10209, n10210,
         n10211, n10212, n10213, n10214, n10215, n10216, n10217, n10218,
         n10219, n10220, n10221, n10222, n10223, n10224, n10225, n10226,
         n10227, n10228, n10229, n10230, n10231, n10232, n10233, n10234,
         n10235, n10236, n10237, n10238, n10239, n10240, n10241, n10242,
         n10243, n10244, n10245, n10246, n10247, n10248, n10249, n10250,
         n10251, n10252, n10253, n10254, n10255, n10256, n10257, n10258,
         n10259, n10260, n10261, n10262, n10263, n10264, n10265, n10266,
         n10267, n10268, n10269, n10270, n10271, n10272, n10273, n10274,
         n10275, n10276, n10277, n10278, n10279, n10280, n10281, n10282,
         n10283, n10284, n10285, n10286, n10287, n10288, n10289, n10290,
         n10291, n10292, n10293, n10294, n10295, n10296, n10297, n10298,
         n10299, n10300, n10301, n10302, n10303, n10304, n10305, n10306,
         n10307, n10308, n10309, n10310, n10311, n10312, n10313, n10314,
         n10315, n10316, n10317, n10318, n10319, n10320, n10321, n10322,
         n10323, n10324, n10325, n10326, n10327, n10328, n10329, n10330,
         n10331, n10332, n10333, n10334, n10335, n10336, n10337, n10338,
         n10339, n10340, n10341, n10342, n10343, n10344, n10345, n10346,
         n10347, n10348, n10349, n10350, n10351, n10352, n10353, n10354,
         n10355, n10356, n10357, n10358, n10359, n10360, n10361, n10362,
         n10363, n10364, n10365, n10366, n10367, n10368, n10369, n10370,
         n10371, n10372, n10373, n10374, n10375, n10376, n10377, n10378,
         n10379, n10380, n10381, n10382, n10383, n10384, n10385, n10386,
         n10387, n10388, n10389, n10390, n10391, n10392, n10393, n10394,
         n10395, n10396, n10397, n10398, n10399, n10400, n10401, n10402,
         n10403, n10404, n10405, n10406, n10407, n10408, n10409, n10410,
         n10411, n10412, n10413, n10414, n10415, n10416, n10417, n10418,
         n10419, n10420, n10421, n10422, n10423, n10424, n10425, n10426,
         n10427, n10428, n10429, n10430, n10431, n10432, n10433, n10434,
         n10435, n10436, n10437, n10438, n10439, n10440, n10441, n10442,
         n10443, n10444, n10445, n10446, n10447, n10448, n10449, n10450,
         n10451, n10452, n10453, n10454, n10455, n10456, n10457, n10458,
         n10459, n10460, n10461, n10462, n10463, n10464, n10465, n10466,
         n10467, n10468, n10469, n10470, n10471, n10472, n10473, n10474,
         n10475, n10476, n10477, n10478, n10479, n10480, n10481, n10482,
         n10483, n10484, n10485, n10486, n10487, n10488, n10489, n10490,
         n10491, n10492, n10493, n10494, n10495, n10496, n10497, n10498,
         n10499, n10500, n10501, n10502, n10503, n10504, n10505, n10506,
         n10507, n10508, n10509, n10510, n10511, n10512, n10513, n10514,
         n10515, n10516, n10517, n10518, n10519, n10520, n10521, n10522,
         n10523, n10524, n10525, n10526, n10527, n10528, n10529, n10530,
         n10531, n10532, n10533, n10534, n10535, n10536, n10537, n10538,
         n10539, n10540, n10541, n10542, n10543, n10544, n10545, n10546,
         n10547, n10548, n10549, n10550, n10551, n10552, n10553, n10554,
         n10555, n10556, n10557, n10558, n10559, n10560, n10561, n10562,
         n10563, n10564, n10565, n10566, n10567, n10568, n10569, n10570,
         n10571, n10572, n10573, n10574, n10575, n10576, n10577, n10578,
         n10579, n10580, n10581, n10582, n10583, n10584, n10585, n10586,
         n10587, n10588, n10589, n10590, n10591, n10592, n10593, n10594,
         n10595, n10596, n10597, n10598, n10599, n10600, n10601, n10602,
         n10603, n10604, n10605, n10606, n10607, n10608, n10609, n10610,
         n10611, n10612, n10613, n10614, n10615, n10616, n10617, n10618,
         n10619, n10620, n10621, n10622, n10623, n10624, n10625, n10626,
         n10627, n10628, n10629, n10630, n10631, n10632, n10633, n10634,
         n10635, n10636, n10637, n10638, n10639, n10640, n10641, n10642,
         n10643, n10644, n10645, n10646, n10647, n10648, n10649, n10650,
         n10651, n10652, n10653, n10654, n10655, n10656, n10657, n10658,
         n10659, n10660, n10661, n10662, n10663, n10664, n10665, n10666,
         n10667, n10668, n10669, n10670, n10671, n10672, n10673, n10674,
         n10675, n10676, n10677, n10678, n10679, n10680, n10681, n10682,
         n10683, n10684, n10685, n10686, n10687, n10688, n10689, n10690,
         n10691, n10692, n10693, n10694, n10695, n10696, n10697, n10698,
         n10699, n10700, n10701, n10702, n10703, n10704, n10705, n10706,
         n10707, n10708, n10709, n10710, n10711, n10712, n10713, n10714,
         n10715, n10716, n10717, n10718, n10719, n10720, n10721, n10722,
         n10723, n10724, n10725, n10726, n10727, n10728, n10729, n10730,
         n10731, n10732, n10733, n10734, n10735, n10736, n10737, n10738,
         n10739, n10740, n10741, n10742, n10743, n10744, n10745, n10746,
         n10747, n10748, n10749, n10750, n10751, n10752, n10753, n10754,
         n10755, n10756, n10757, n10758, n10759, n10760, n10761, n10762,
         n10763, n10764, n10765, n10766, n10767, n10768, n10769, n10770,
         n10771, n10772, n10773, n10774, n10775, n10776, n10777, n10778,
         n10779, n10780, n10781, n10782, n10783, n10784, n10785, n10786,
         n10787, n10788, n10789, n10790, n10791, n10792, n10793, n10794,
         n10795, n10796, n10797, n10798, n10799, n10800, n10801, n10802,
         n10803, n10804, n10805, n10806, n10807, n10808, n10809, n10810,
         n10811, n10812, n10813, n10814, n10815, n10816, n10817, n10818,
         n10819, n10820, n10821, n10822, n10823, n10824, n10825, n10826,
         n10827, n10828, n10829, n10830, n10831, n10832, n10833, n10834,
         n10835, n10836, n10837, n10838, n10839, n10840, n10841, n10842,
         n10843, n10844, n10845, n10846, n10847, n10848, n10849, n10850,
         n10851, n10852, n10853, n10854, n10855, n10856, n10857, n10858,
         n10859, n10860, n10861, n10862, n10863, n10864, n10865, n10866,
         n10867, n10868, n10869, n10870, n10871, n10872, n10873, n10874,
         n10875, n10876, n10877, n10878, n10879, n10880, n10881, n10882,
         n10883, n10884, n10885, n10886, n10887, n10888, n10889, n10890,
         n10891, n10892, n10893, n10894, n10895, n10896, n10897, n10898,
         n10899, n10900, n10901, n10902, n10903, n10904, n10905, n10906,
         n10907, n10908, n10909, n10910, n10911, n10912, n10913, n10914,
         n10915, n10916, n10917, n10918, n10919, n10920, n10921, n10922,
         n10923, n10924, n10925, n10926, n10927, n10928, n10929, n10930,
         n10931, n10932, n10933, n10934, n10935, n10936, n10937, n10938,
         n10939, n10940, n10941, n10942, n10943, n10944, n10945, n10946,
         n10947, n10948, n10949, n10950, n10951, n10952, n10953, n10954,
         n10955, n10956, n10957, n10958, n10959, n10960, n10961, n10962,
         n10963, n10964, n10965, n10966, n10967, n10968, n10969, n10970,
         n10971, n10972, n10973, n10974, n10975, n10976, n10977, n10978,
         n10979, n10980, n10981, n10982, n10983, n10984, n10985, n10986,
         n10987, n10988, n10989, n10990, n10991, n10992, n10993, n10994,
         n10995, n10996, n10997, n10998, n10999, n11000, n11001, n11002,
         n11003, n11004, n11005, n11006, n11007, n11008, n11009, n11010,
         n11011, n11012, n11013, n11014, n11015, n11016, n11017, n11018,
         n11019, n11020, n11021, n11022, n11023, n11024, n11025, n11026,
         n11027, n11028, n11029, n11030, n11031, n11032, n11033, n11034,
         n11035, n11036, n11037, n11038, n11039, n11040, n11041, n11042,
         n11043, n11044, n11045, n11046, n11047, n11048, n11049, n11050,
         n11051, n11052, n11053, n11054, n11055, n11056, n11057, n11058,
         n11059, n11060, n11061, n11062, n11063, n11064, n11065, n11066,
         n11067, n11068, n11069, n11070, n11071, n11072, n11073, n11074,
         n11075, n11076, n11077, n11078, n11079, n11080, n11081, n11082,
         n11083, n11084, n11085, n11086, n11087, n11088, n11089, n11090,
         n11091, n11092, n11093, n11094, n11095, n11096, n11097, n11098,
         n11099, n11100, n11101, n11102, n11103, n11104, n11105, n11106,
         n11107, n11108, n11109, n11110, n11111, n11112, n11113, n11114,
         n11115, n11116, n11117, n11118, n11119, n11120, n11121, n11122,
         n11123, n11124, n11125, n11126, n11127, n11128, n11129, n11130,
         n11131, n11132, n11133, n11134, n11135, n11136, n11137, n11138,
         n11139, n11140, n11141, n11142, n11143, n11144, n11145, n11146,
         n11147, n11148, n11149, n11150, n11151, n11152, n11153, n11154,
         n11155, n11156, n11157, n11158, n11159, n11160, n11161, n11162,
         n11163, n11164, n11165, n11166, n11167, n11168, n11169, n11170,
         n11171, n11172, n11173, n11174, n11175, n11176, n11177, n11178,
         n11179, n11180, n11181, n11182, n11183, n11184, n11185, n11186,
         n11187, n11188, n11189, n11190, n11191, n11192, n11193, n11194,
         n11195, n11196, n11197, n11198, n11199, n11200, n11201, n11202,
         n11203, n11204, n11205, n11206, n11207, n11208, n11209, n11210,
         n11211, n11212, n11213, n11214, n11215, n11216, n11217, n11218,
         n11219, n11220, n11221, n11222, n11223, n11224, n11225, n11226,
         n11227, n11228, n11229, n11230, n11231, n11232, n11233, n11234,
         n11235, n11236, n11237, n11238, n11239, n11240, n11241, n11242,
         n11243, n11244, n11245, n11246, n11247, n11248, n11249, n11250,
         n11251, n11252, n11253, n11254, n11255, n11256, n11257, n11258,
         n11259, n11260, n11261, n11262, n11263, n11264, n11265, n11266,
         n11267, n11268, n11269, n11270, n11271, n11272, n11273, n11274,
         n11275, n11276, n11277, n11278, n11279, n11280, n11281, n11282,
         n11283, n11284, n11285, n11286, n11287, n11288, n11289, n11290,
         n11291, n11292, n11293, n11294, n11295, n11296, n11297, n11298,
         n11299, n11300, n11301, n11302, n11303, n11304, n11305, n11306,
         n11307, n11308, n11309, n11310, n11311, n11312, n11313, n11314,
         n11315, n11316, n11317, n11318, n11319, n11320, n11321, n11322,
         n11323, n11324, n11325, n11326, n11327, n11328, n11329, n11330,
         n11331, n11332, n11333, n11334, n11335, n11336, n11337, n11338,
         n11339, n11340, n11341, n11342, n11343, n11344, n11345, n11346,
         n11347, n11348, n11349, n11350, n11351, n11352, n11353, n11354,
         n11355, n11356, n11357, n11358, n11359, n11360, n11361, n11362,
         n11363, n11364, n11365, n11366, n11367, n11368, n11369, n11370,
         n11371, n11372, n11373, n11374, n11375, n11376, n11377, n11378,
         n11379, n11380, n11381, n11382, n11383, n11384, n11385, n11386,
         n11387, n11388, n11389, n11390, n11391, n11392, n11393, n11394,
         n11395, n11396, n11397, n11398, n11399, n11400, n11401, n11402,
         n11403, n11404, n11405, n11406, n11407, n11408, n11409, n11410,
         n11411, n11412, n11413, n11414, n11415, n11416, n11417, n11418,
         n11419, n11420, n11421, n11422, n11423, n11424, n11425, n11426,
         n11427, n11428, n11429, n11430, n11431, n11432, n11433, n11434,
         n11435, n11436, n11437, n11438, n11439, n11440, n11441, n11442,
         n11443, n11444, n11445, n11446, n11447, n11448, n11449, n11450,
         n11451, n11452, n11453, n11454, n11455, n11456, n11457, n11458,
         n11459, n11460, n11461, n11462, n11463, n11464, n11465, n11466,
         n11467, n11468, n11469, n11470, n11471, n11472, n11473, n11474,
         n11475, n11476, n11477, n11478, n11479, n11480, n11481, n11482,
         n11483, n11484, n11485, n11486, n11487, n11488, n11489, n11490,
         n11491, n11492, n11493, n11494, n11495, n11496, n11497, n11498,
         n11499, n11500, n11501, n11502, n11503, n11504, n11505, n11506,
         n11507, n11508, n11509, n11510, n11511, n11512, n11513, n11514,
         n11515, n11516, n11517, n11518, n11519, n11520, n11521, n11522,
         n11523, n11524, n11525, n11526, n11527, n11528, n11529, n11530,
         n11531, n11532, n11533, n11534, n11535, n11536, n11537, n11538,
         n11539, n11540, n11541, n11542, n11543, n11544, n11545, n11546,
         n11547, n11548, n11549, n11550, n11551, n11552, n11553, n11554,
         n11555, n11556, n11557, n11558, n11559, n11560, n11561, n11562,
         n11563, n11564, n11565, n11566, n11567, n11568, n11569, n11570,
         n11571, n11572, n11573, n11574, n11575, n11576, n11577, n11578,
         n11579, n11580, n11581, n11582, n11583, n11584, n11585, n11586,
         n11587, n11588, n11589, n11590, n11591, n11592, n11593, n11594,
         n11595, n11596, n11597, n11598, n11599, n11600, n11601, n11602,
         n11603, n11604, n11605, n11606, n11607, n11608, n11609, n11610,
         n11611, n11612, n11613, n11614, n11615, n11616, n11617, n11618,
         n11619, n11620, n11621, n11622, n11623, n11624, n11625, n11626,
         n11627, n11628, n11629, n11630, n11631, n11632, n11633, n11634,
         n11635, n11636, n11637, n11638, n11639, n11640, n11641, n11642,
         n11643, n11644, n11645, n11646, n11647, n11648, n11649, n11650,
         n11651, n11652, n11653, n11654, n11655, n11656, n11657, n11658,
         n11659, n11660, n11661, n11662, n11663, n11664, n11665, n11666,
         n11667, n11668, n11669, n11670, n11671, n11672, n11673, n11674,
         n11675, n11676, n11677, n11678, n11679, n11680, n11681, n11682,
         n11683, n11684, n11685, n11686, n11687, n11688, n11689, n11690,
         n11691, n11692, n11693, n11694, n11695, n11696, n11697, n11698,
         n11699, n11700, n11701, n11702, n11703, n11704, n11705, n11706,
         n11707, n11708, n11709, n11710, n11711, n11712, n11713, n11714,
         n11715, n11716, n11717, n11718, n11719, n11720, n11721, n11722,
         n11723, n11724, n11725, n11726, n11727, n11728, n11729, n11730,
         n11731, n11732, n11733, n11734, n11735, n11736, n11737, n11738,
         n11739, n11740, n11741, n11742, n11743, n11744, n11745, n11746,
         n11747, n11748, n11749, n11750, n11751, n11752, n11753, n11754,
         n11755, n11756, n11757, n11758, n11759, n11760, n11761, n11762,
         n11763, n11764, n11765, n11766, n11767, n11768, n11769, n11770,
         n11771, n11772, n11773, n11774, n11775, n11776, n11777, n11778,
         n11779, n11780, n11781, n11782, n11783, n11784, n11785, n11786,
         n11787, n11788, n11789, n11790, n11791, n11792, n11793, n11794,
         n11795, n11796, n11797, n11798, n11799, n11800, n11801, n11802,
         n11803, n11804, n11805, n11806, n11807, n11808, n11809, n11810,
         n11811, n11812, n11813, n11814, n11815, n11816, n11817, n11818,
         n11819, n11820, n11821, n11822, n11823, n11824, n11825, n11826,
         n11827, n11828, n11829, n11830, n11831, n11832, n11833, n11834,
         n11835, n11836, n11837, n11838, n11839, n11840, n11841, n11842,
         n11843, n11844, n11845, n11846, n11847, n11848, n11849, n11850,
         n11851, n11852, n11853, n11854, n11855, n11856, n11857, n11858,
         n11859, n11860, n11861, n11862, n11863, n11864, n11865, n11866,
         n11867, n11868, n11869, n11870, n11871, n11872, n11873, n11874,
         n11875, n11876, n11877, n11878, n11879, n11880, n11881, n11882,
         n11883, n11884, n11885, n11886, n11887, n11888, n11889, n11890,
         n11891, n11892, n11893, n11894, n11895, n11896, n11897, n11898,
         n11899, n11900, n11901, n11902, n11903, n11904, n11905, n11906,
         n11907, n11908, n11909, n11910, n11911, n11912, n11913, n11914,
         n11915, n11916, n11917, n11918, n11919, n11920, n11921, n11922,
         n11923, n11924, n11925, n11926, n11927, n11928, n11929, n11930,
         n11931, n11932, n11933, n11934, n11935, n11936, n11937, n11938,
         n11939, n11940, n11941, n11942, n11943, n11944, n11945, n11946,
         n11947, n11948, n11949, n11950, n11951, n11952, n11953, n11954,
         n11955, n11956, n11957, n11958, n11959, n11960, n11961, n11962,
         n11963, n11964, n11965, n11966, n11967, n11968, n11969, n11970,
         n11971, n11972, n11973, n11974, n11975, n11976, n11977, n11978,
         n11979, n11980, n11981, n11982, n11983, n11984, n11985, n11986,
         n11987, n11988, n11989, n11990, n11991, n11992, n11993, n11994,
         n11995, n11996, n11997, n11998, n11999, n12000, n12001, n12002,
         n12003, n12004, n12005, n12006, n12007, n12008, n12009, n12010,
         n12011, n12012, n12013, n12014, n12015, n12016, n12017, n12018,
         n12019, n12020, n12021, n12022, n12023, n12024, n12025, n12026,
         n12027, n12028, n12029, n12030, n12031, n12032, n12033, n12034,
         n12035, n12036, n12037, n12038, n12039, n12040, n12041, n12042,
         n12043, n12044, n12045, n12046, n12047, n12048, n12049, n12050,
         n12051, n12052, n12053, n12054, n12055, n12056, n12057, n12058,
         n12059, n12060, n12061, n12062, n12063, n12064, n12065, n12066,
         n12067, n12068, n12069, n12070, n12071, n12072, n12073, n12074,
         n12075, n12076, n12077, n12078, n12079, n12080, n12081, n12082,
         n12083, n12084, n12085, n12086, n12087, n12088, n12089, n12090,
         n12091, n12092, n12093, n12094, n12095, n12096, n12097, n12098,
         n12099, n12100, n12101, n12102, n12103, n12104, n12105, n12106,
         n12107, n12108, n12109, n12110, n12111, n12112, n12113, n12114,
         n12115, n12116, n12117, n12118, n12119, n12120, n12121, n12122,
         n12123, n12124, n12125, n12126, n12127, n12128, n12129, n12130,
         n12131, n12132, n12133, n12134, n12135, n12136, n12137, n12138,
         n12139, n12140, n12141, n12142, n12143, n12144, n12145, n12146,
         n12147, n12148, n12149, n12150, n12151, n12152, n12153, n12154,
         n12155, n12156, n12157, n12158, n12159, n12160, n12161, n12162,
         n12163, n12164, n12165, n12166, n12167, n12168, n12169, n12170,
         n12171, n12172, n12173, n12174, n12175, n12176, n12177, n12178,
         n12179, n12180, n12181, n12182, n12183, n12184, n12185, n12186,
         n12187, n12188, n12189, n12190, n12191, n12192, n12193, n12194,
         n12195, n12196, n12197, n12198, n12199, n12200, n12201, n12202,
         n12203, n12204, n12205, n12206, n12207, n12208, n12209, n12210,
         n12211, n12212, n12213, n12214, n12215, n12216, n12217, n12218,
         n12219, n12220, n12221, n12222, n12223, n12224, n12225, n12226,
         n12227, n12228, n12229, n12230, n12231, n12232, n12233, n12234,
         n12235, n12236, n12237, n12238, n12239, n12240, n12241, n12242,
         n12243, n12244, n12245, n12246, n12247, n12248, n12249, n12250,
         n12251, n12252, n12253, n12254, n12255, n12256, n12257, n12258,
         n12259, n12260, n12261, n12262, n12263, n12264, n12265, n12266,
         n12267, n12268, n12269, n12270, n12271, n12272, n12273, n12274,
         n12275, n12276, n12277, n12278, n12279, n12280, n12281, n12282,
         n12283, n12284, n12285, n12286, n12287, n12288, n12289, n12290,
         n12291, n12292, n12293, n12294, n12295, n12296, n12297, n12298,
         n12299, n12300, n12301, n12302, n12303, n12304, n12305, n12306,
         n12307, n12308, n12309, n12310, n12311, n12312, n12313, n12314,
         n12315, n12316, n12317, n12318, n12319, n12320, n12321, n12322,
         n12323, n12324, n12325, n12326, n12327, n12328, n12329, n12330,
         n12331, n12332, n12333, n12334, n12335, n12336, n12337, n12338,
         n12339, n12340, n12341, n12342, n12343, n12344, n12345, n12346,
         n12347, n12348, n12349, n12350, n12351, n12352, n12353, n12354,
         n12355, n12356, n12357, n12358, n12359, n12360, n12361, n12362,
         n12363, n12364, n12365, n12366, n12367, n12368, n12369, n12370,
         n12371, n12372, n12373, n12374, n12375, n12376, n12377, n12378,
         n12379, n12380, n12381, n12382, n12383, n12384, n12385, n12386,
         n12387, n12388, n12389, n12390, n12391, n12392, n12393, n12394,
         n12395, n12396, n12397, n12398, n12399, n12400, n12401, n12402,
         n12403, n12404, n12405, n12406, n12407, n12408, n12409, n12410,
         n12411, n12412, n12413, n12414, n12415, n12416, n12417, n12418,
         n12419, n12420, n12421, n12422, n12423, n12424, n12425, n12426,
         n12427, n12428, n12429, n12430, n12431, n12432, n12433, n12434,
         n12435, n12436, n12437, n12438, n12439, n12440, n12441, n12442,
         n12443, n12444, n12445, n12446, n12447, n12448, n12449, n12450,
         n12451, n12452, n12453, n12454, n12455, n12456, n12457, n12458,
         n12459, n12460, n12461, n12462, n12463, n12464, n12465, n12466,
         n12467, n12468, n12469, n12470, n12471, n12472, n12473, n12474,
         n12475, n12476, n12477, n12478, n12479, n12480, n12481, n12482,
         n12483, n12484, n12485, n12486, n12487, n12488, n12489, n12490,
         n12491, n12492, n12493, n12494, n12495, n12496, n12497, n12498,
         n12499, n12500, n12501, n12502, n12503, n12504, n12505, n12506,
         n12507, n12508, n12509, n12510, n12511, n12512, n12513, n12514,
         n12515, n12516, n12517, n12518, n12519, n12520, n12521, n12522,
         n12523, n12524, n12525, n12526, n12527, n12528, n12529, n12530,
         n12531, n12532, n12533, n12534, n12535, n12536, n12537, n12538,
         n12539, n12540, n12541, n12542, n12543, n12544, n12545, n12546,
         n12547, n12548, n12549, n12550, n12551, n12552, n12553, n12554,
         n12555, n12556, n12557, n12558, n12559, n12560, n12561, n12562,
         n12563, n12564, n12565, n12566, n12567, n12568, n12569, n12570,
         n12571, n12572, n12573, n12574, n12575, n12576, n12577, n12578,
         n12579, n12580, n12581, n12582, n12583, n12584, n12585, n12586,
         n12587, n12588, n12589, n12590, n12591, n12592, n12593, n12594,
         n12595, n12596, n12597, n12598, n12599, n12600, n12601, n12602,
         n12603, n12604, n12605, n12606, n12607, n12608, n12609, n12610,
         n12611, n12612, n12613, n12614, n12615, n12616, n12617, n12618,
         n12619, n12620, n12621, n12622, n12623, n12624, n12625, n12626,
         n12627, n12628, n12629, n12630, n12631, n12632, n12633, n12634,
         n12635, n12636, n12637, n12638, n12639, n12640, n12641, n12642,
         n12643, n12644, n12645, n12646, n12647, n12648, n12649, n12650,
         n12651, n12652, n12653, n12654, n12655, n12656, n12657, n12658,
         n12659, n12660, n12661, n12662, n12663, n12664, n12665, n12666,
         n12667, n12668, n12669, n12670, n12671, n12672, n12673, n12674,
         n12675, n12676, n12677, n12678, n12679, n12680, n12681, n12682,
         n12683, n12684, n12685, n12686, n12687, n12688, n12689, n12690,
         n12691, n12692, n12693, n12694, n12695, n12696, n12697, n12698,
         n12699, n12700, n12701, n12702, n12703, n12704, n12705, n12706,
         n12707, n12708, n12709, n12710, n12711, n12712, n12713, n12714,
         n12715, n12716, n12717, n12718, n12719, n12720, n12721, n12722,
         n12723, n12724, n12725, n12726, n12727, n12728, n12729, n12730,
         n12731, n12732, n12733, n12734, n12735, n12736, n12737, n12738,
         n12739, n12740, n12741, n12742, n12743, n12744, n12745, n12746,
         n12747, n12748, n12749, n12750, n12751, n12752, n12753, n12754,
         n12755, n12756, n12757, n12758, n12759, n12760, n12761, n12762,
         n12763, n12764, n12765, n12766, n12767, n12768, n12769, n12770,
         n12771, n12772, n12773, n12774, n12775, n12776, n12777, n12778,
         n12779, n12780, n12781, n12782, n12783, n12784, n12785, n12786,
         n12787, n12788, n12789, n12790, n12791, n12792, n12793, n12794,
         n12795, n12796, n12797, n12798, n12799, n12800, n12801, n12802,
         n12803, n12804, n12805, n12806, n12807, n12808, n12809, n12810,
         n12811, n12812, n12813, n12814, n12815, n12816, n12817, n12818,
         n12819, n12820, n12821, n12822, n12823, n12824, n12825, n12826,
         n12827, n12828, n12829, n12830, n12831, n12832, n12833, n12834,
         n12835, n12836, n12837, n12838, n12839, n12840, n12841, n12842,
         n12843, n12844, n12845, n12846, n12847, n12848, n12849, n12850,
         n12851, n12852, n12853, n12854, n12855, n12856, n12857, n12858,
         n12859, n12860, n12861, n12862, n12863, n12864, n12865, n12866,
         n12867, n12868, n12869, n12870, n12871, n12872, n12873, n12874,
         n12875, n12876, n12877, n12878, n12879, n12880, n12881, n12882,
         n12883, n12884, n12885, n12886, n12887, n12888, n12889, n12890,
         n12891, n12892, n12893, n12894, n12895, n12896, n12897, n12898,
         n12899, n12900, n12901, n12902, n12903, n12904, n12905, n12906,
         n12907, n12908, n12909, n12910, n12911, n12912, n12913, n12914,
         n12915, n12916, n12917, n12918, n12919, n12920, n12921, n12922,
         n12923, n12924, n12925, n12926, n12927, n12928, n12929, n12930,
         n12931, n12932, n12933, n12934, n12935, n12936, n12937, n12938,
         n12939, n12940, n12941, n12942, n12943, n12944, n12945, n12946,
         n12947, n12948, n12949, n12950, n12951, n12952, n12953, n12954,
         n12955, n12956, n12957, n12958, n12959, n12960, n12961, n12962,
         n12963, n12964, n12965, n12966, n12967, n12968, n12969, n12970,
         n12971, n12972, n12973, n12974, n12975, n12976, n12977, n12978,
         n12979, n12980, n12981, n12982, n12983, n12984, n12985, n12986,
         n12987, n12988, n12989, n12990, n12991, n12992, n12993, n12994,
         n12995, n12996, n12997, n12998, n12999, n13000, n13001, n13002,
         n13003, n13004, n13005, n13006, n13007, n13008, n13009, n13010,
         n13011, n13012, n13013, n13014, n13015, n13016, n13017, n13018,
         n13019, n13020, n13021, n13022, n13023, n13024, n13025, n13026,
         n13027, n13028, n13029, n13030, n13031, n13032, n13033, n13034,
         n13035, n13036, n13037, n13038, n13039, n13040, n13041, n13042,
         n13043, n13044, n13045, n13046, n13047, n13048, n13049, n13050,
         n13051, n13052, n13053, n13054, n13055, n13056, n13057, n13058,
         n13059, n13060, n13061, n13062, n13063, n13064, n13065, n13066,
         n13067, n13068, n13069, n13070, n13071, n13072, n13073, n13074,
         n13075, n13076, n13077, n13078, n13079, n13080, n13081, n13082,
         n13083, n13084, n13085, n13086, n13087, n13088, n13089, n13090,
         n13091, n13092, n13093, n13094, n13095, n13096, n13097, n13098,
         n13099, n13100, n13101, n13102, n13103, n13104, n13105, n13106,
         n13107, n13108, n13109, n13110, n13111, n13112, n13113, n13114,
         n13115, n13116, n13117, n13118, n13119, n13120, n13121, n13122,
         n13123, n13124, n13125, n13126, n13127, n13128, n13129, n13130,
         n13131, n13132, n13133, n13134, n13135, n13136, n13137, n13138,
         n13139, n13140, n13141, n13142, n13143, n13144, n13145, n13146,
         n13147, n13148, n13149, n13150, n13151, n13152, n13153, n13154,
         n13155, n13156, n13157, n13158, n13159, n13160, n13161, n13162,
         n13163, n13164, n13165, n13166, n13167, n13168, n13169, n13170,
         n13171, n13172, n13173, n13174, n13175, n13176, n13177, n13178,
         n13179, n13180, n13181, n13182, n13183, n13184, n13185, n13186,
         n13187, n13188, n13189, n13190, n13191, n13192, n13193, n13194,
         n13195, n13196, n13197, n13198, n13199, n13200, n13201, n13202,
         n13203, n13204, n13205, n13206, n13207, n13208, n13209, n13210,
         n13211, n13212, n13213, n13214, n13215, n13216, n13217, n13218,
         n13219, n13220, n13221, n13222, n13223, n13224, n13225, n13226,
         n13227, n13228, n13229, n13230, n13231, n13232, n13233, n13234,
         n13235, n13236, n13237, n13238, n13239, n13240, n13241, n13242,
         n13243, n13244, n13245, n13246, n13247, n13248, n13249, n13250,
         n13251, n13252, n13253, n13254, n13255, n13256, n13257, n13258,
         n13259, n13260, n13261, n13262, n13263, n13264, n13265, n13266,
         n13267, n13268, n13269, n13270, n13271, n13272, n13273, n13274,
         n13275, n13276, n13277, n13278, n13279, n13280, n13281, n13282,
         n13283, n13284, n13285, n13286, n13287, n13288, n13289, n13290,
         n13291, n13292, n13293, n13294, n13295, n13296, n13297, n13298,
         n13299, n13300, n13301, n13302, n13303, n13304, n13305, n13306,
         n13307, n13308, n13309, n13310, n13311, n13312, n13313, n13314,
         n13315, n13316, n13317, n13318, n13319, n13320, n13321, n13322,
         n13323, n13324, n13325, n13326, n13327, n13328, n13329, n13330,
         n13331, n13332, n13333, n13334, n13335, n13336, n13337, n13338,
         n13339, n13340, n13341, n13342, n13343, n13344, n13345, n13346,
         n13347, n13348, n13349, n13350, n13351, n13352, n13353, n13354,
         n13355, n13356, n13357, n13358, n13359, n13360, n13361, n13362,
         n13363, n13364, n13365, n13366, n13367, n13368, n13369, n13370,
         n13371, n13372, n13373, n13374, n13375, n13376, n13377, n13378,
         n13379, n13380, n13381, n13382, n13383, n13384, n13385, n13386,
         n13387, n13388, n13389, n13390, n13391, n13392, n13393, n13394,
         n13395, n13396, n13397, n13398, n13399, n13400, n13401, n13402,
         n13403, n13404, n13405, n13406, n13407, n13408, n13409, n13410,
         n13411, n13412, n13413, n13414, n13415, n13416, n13417, n13418,
         n13419, n13420, n13421, n13422, n13423, n13424, n13425, n13426,
         n13427, n13428, n13429, n13430, n13431, n13432, n13433, n13434,
         n13435, n13436, n13437, n13438, n13439, n13440, n13441, n13442,
         n13443, n13444, n13445, n13446, n13447, n13448, n13449, n13450,
         n13451, n13452, n13453, n13454, n13455, n13456, n13457, n13458,
         n13459, n13460, n13461, n13462, n13463, n13464, n13465, n13466,
         n13467, n13468, n13469, n13470, n13471, n13472, n13473, n13474,
         n13475, n13476, n13477, n13478, n13479, n13480, n13481, n13482,
         n13483, n13484, n13485, n13486, n13487, n13488, n13489, n13490,
         n13491, n13492, n13493, n13494, n13495, n13496, n13497, n13498,
         n13499, n13500, n13501, n13502, n13503, n13504, n13505, n13506,
         n13507, n13508, n13509, n13510, n13511, n13512, n13513, n13514,
         n13515, n13516, n13517, n13518, n13519, n13520, n13521, n13522,
         n13523, n13524, n13525, n13526, n13527, n13528, n13529, n13530,
         n13531, n13532, n13533, n13534, n13535, n13536, n13537, n13538,
         n13539, n13540, n13541, n13542, n13543, n13544, n13545, n13546,
         n13547, n13548, n13549, n13550, n13551, n13552, n13553, n13554,
         n13555, n13556, n13557, n13558, n13559, n13560, n13561, n13562,
         n13563, n13564, n13565, n13566, n13567, n13568, n13569, n13570,
         n13571, n13572, n13573, n13574, n13575, n13576, n13577, n13578,
         n13579, n13580, n13581, n13582, n13583, n13584, n13585, n13586,
         n13587, n13588, n13589, n13590, n13591, n13592, n13593, n13594,
         n13595, n13596, n13597, n13598, n13599, n13600, n13601, n13602,
         n13603, n13604, n13605, n13606, n13607, n13608, n13609, n13610,
         n13611, n13612, n13613, n13614, n13615, n13616, n13617, n13618,
         n13619, n13620, n13621, n13622, n13623, n13624, n13625, n13626,
         n13627, n13628, n13629, n13630, n13631, n13632, n13633, n13634,
         n13635, n13636, n13637, n13638, n13639, n13640, n13641, n13642,
         n13643, n13644, n13645, n13646, n13647, n13648, n13649, n13650,
         n13651, n13652, n13653, n13654, n13655, n13656, n13657, n13658,
         n13659, n13660, n13661, n13662, n13663, n13664, n13665, n13666,
         n13667, n13668, n13669, n13670, n13671, n13672, n13673, n13674,
         n13675, n13676, n13677, n13678, n13679, n13680, n13681, n13682,
         n13683, n13684, n13685, n13686, n13687, n13688, n13689, n13690,
         n13691, n13692, n13693, n13694, n13695, n13696, n13697, n13698,
         n13699, n13700, n13701, n13702, n13703, n13704, n13705, n13706,
         n13707, n13708, n13709, n13710, n13711, n13712, n13713, n13714,
         n13715, n13716, n13717, n13718, n13719, n13720, n13721, n13722,
         n13723, n13724, n13725, n13726, n13727, n13728, n13729, n13730,
         n13731, n13732, n13733, n13734, n13735, n13736, n13737, n13738,
         n13739, n13740, n13741, n13742, n13743, n13744, n13745, n13746,
         n13747, n13748, n13749, n13750, n13751, n13752, n13753, n13754,
         n13755, n13756, n13757, n13758, n13759, n13760, n13761, n13762,
         n13763, n13764, n13765, n13766, n13767, n13768, n13769, n13770,
         n13771, n13772, n13773, n13774, n13775, n13776, n13777, n13778,
         n13779, n13780, n13781, n13782, n13783, n13784, n13785, n13786,
         n13787, n13788, n13789, n13790, n13791, n13792, n13793, n13794,
         n13795, n13796, n13797, n13798, n13799, n13800, n13801, n13802,
         n13803, n13804, n13805, n13806, n13807, n13808, n13809, n13810,
         n13811, n13812, n13813, n13814, n13815, n13816, n13817, n13818,
         n13819, n13820, n13821, n13822, n13823, n13824, n13825, n13826,
         n13827, n13828, n13829, n13830, n13831, n13832, n13833, n13834,
         n13835, n13836, n13837, n13838, n13839, n13840, n13841, n13842,
         n13843, n13844, n13845, n13846, n13847, n13848, n13849, n13850,
         n13851, n13852, n13853, n13854, n13855, n13856, n13857, n13858,
         n13859, n13860, n13861, n13862, n13863, n13864, n13865, n13866,
         n13867, n13868, n13869, n13870, n13871, n13872, n13873, n13874,
         n13875, n13876, n13877, n13878, n13879, n13880, n13881, n13882,
         n13883, n13884, n13885, n13886, n13887, n13888, n13889, n13890,
         n13891, n13892, n13893, n13894, n13895, n13896, n13897, n13898,
         n13899, n13900, n13901, n13902, n13903, n13904, n13905, n13906,
         n13907, n13908, n13909, n13910, n13911, n13912, n13913, n13914,
         n13915, n13916, n13917, n13918, n13919, n13920, n13921, n13922,
         n13923, n13924, n13925, n13926, n13927, n13928, n13929, n13930,
         n13931, n13932, n13933, n13934, n13935, n13936, n13937, n13938,
         n13939, n13940, n13941, n13942, n13943, n13944, n13945, n13946,
         n13947, n13948, n13949, n13950, n13951, n13952, n13953, n13954,
         n13955, n13956, n13957, n13958, n13959, n13960, n13961, n13962,
         n13963, n13964, n13965, n13966, n13967, n13968, n13969, n13970,
         n13971, n13972, n13973, n13974, n13975, n13976, n13977, n13978,
         n13979, n13980, n13981, n13982, n13983, n13984, n13985, n13986,
         n13987, n13988, n13989, n13990, n13991, n13992, n13993, n13994,
         n13995, n13996, n13997, n13998, n13999, n14000, n14001, n14002,
         n14003, n14004, n14005, n14006, n14007, n14008, n14009, n14010,
         n14011, n14012, n14013, n14014, n14015, n14016, n14017, n14018,
         n14019, n14020, n14021, n14022, n14023, n14024, n14025, n14026,
         n14027, n14028, n14029, n14030, n14031, n14032, n14033, n14034,
         n14035, n14036, n14037, n14038, n14039, n14040, n14041, n14042,
         n14043, n14044, n14045, n14046, n14047, n14048, n14049, n14050,
         n14051, n14052, n14053, n14054, n14055, n14056, n14057, n14058,
         n14059, n14060, n14061, n14062, n14063, n14064, n14065, n14066,
         n14067, n14068, n14069, n14070, n14071, n14072, n14073, n14074,
         n14075, n14076, n14077, n14078, n14079, n14080, n14081, n14082,
         n14083, n14084, n14085, n14086, n14087, n14088, n14089, n14090,
         n14091, n14092, n14093, n14094, n14095, n14096, n14097, n14098,
         n14099, n14100, n14101, n14102, n14103, n14104, n14105, n14106,
         n14107, n14108, n14109, n14110, n14111, n14112, n14113, n14114,
         n14115, n14116, n14117, n14118, n14119, n14120, n14121, n14122,
         n14123, n14124, n14125, n14126, n14127, n14128, n14129, n14130,
         n14131, n14132, n14133, n14134, n14135, n14136, n14137, n14138,
         n14139, n14140, n14141, n14142, n14143, n14144, n14145, n14146,
         n14147, n14148, n14149, n14150, n14151, n14152, n14153, n14154,
         n14155, n14156, n14157, n14158, n14159, n14160, n14161, n14162,
         n14163, n14164, n14165, n14166, n14167, n14168, n14169, n14170,
         n14171, n14172, n14173, n14174, n14175, n14176, n14177, n14178,
         n14179, n14180, n14181, n14182, n14183, n14184, n14185, n14186,
         n14187, n14188, n14189, n14190, n14191, n14192, n14193, n14194,
         n14195, n14196, n14197, n14198, n14199, n14200, n14201, n14202,
         n14203, n14204, n14205, n14206, n14207, n14208, n14209, n14210,
         n14211, n14212, n14213, n14214, n14215, n14216, n14217, n14218,
         n14219, n14220, n14221, n14222, n14223, n14224, n14225, n14226,
         n14227, n14228, n14229, n14230, n14231, n14232, n14233, n14234,
         n14235, n14236, n14237, n14238, n14239, n14240, n14241, n14242,
         n14243, n14244, n14245, n14246, n14247, n14248, n14249, n14250,
         n14251, n14252, n14253, n14254, n14255, n14256, n14257, n14258,
         n14259, n14260, n14261, n14262, n14263, n14264, n14265, n14266,
         n14267, n14268, n14269, n14270, n14271, n14272, n14273, n14274,
         n14275, n14276, n14277, n14278, n14279, n14280, n14281, n14282,
         n14283, n14284, n14285, n14286, n14287, n14288, n14289, n14290,
         n14291, n14292, n14293, n14294, n14295, n14296, n14297, n14298,
         n14299, n14300, n14301, n14302, n14303, n14304, n14305, n14306,
         n14307, n14308, n14309, n14310, n14311, n14312, n14313, n14314,
         n14315, n14316, n14317, n14318, n14319, n14320, n14321, n14322,
         n14323, n14324, n14325, n14326, n14327, n14328, n14329, n14330,
         n14331, n14332, n14333, n14334, n14335, n14336, n14337, n14338,
         n14339, n14340, n14341, n14342, n14343, n14344, n14345, n14346,
         n14347, n14348, n14349, n14350, n14351, n14352, n14353, n14354,
         n14355, n14356, n14357, n14358, n14359, n14360, n14361, n14362,
         n14363, n14364, n14365, n14366, n14367, n14368, n14369, n14370,
         n14371, n14372, n14373, n14374, n14375, n14376, n14377, n14378,
         n14379, n14380, n14381, n14382, n14383, n14384, n14385, n14386,
         n14387, n14388, n14389, n14390, n14391, n14392, n14393, n14394,
         n14395, n14396, n14397, n14398, n14399, n14400, n14401, n14402,
         n14403, n14404, n14405, n14406, n14407, n14408, n14409, n14410,
         n14411, n14412, n14413, n14414, n14415, n14416, n14417, n14418,
         n14419, n14420, n14421, n14422, n14423, n14424, n14425, n14426,
         n14427, n14428, n14429, n14430, n14431, n14432, n14433, n14434,
         n14435, n14436, n14437, n14438, n14439, n14440, n14441, n14442,
         n14443, n14444, n14445, n14446, n14447, n14448, n14449, n14450,
         n14451, n14452, n14453, n14454, n14455, n14456, n14457, n14458,
         n14459, n14460, n14461, n14462, n14463, n14464, n14465, n14466,
         n14467, n14468, n14469, n14470, n14471, n14472, n14473, n14474,
         n14475, n14476, n14477, n14478, n14479, n14480, n14481, n14482,
         n14483, n14484, n14485, n14486, n14487, n14488, n14489, n14490,
         n14491, n14492, n14493, n14494, n14495, n14496, n14497, n14498,
         n14499, n14500, n14501, n14502, n14503, n14504, n14505, n14506,
         n14507, n14508, n14509, n14510, n14511, n14512, n14513, n14514,
         n14515, n14516, n14517, n14518, n14519, n14520, n14521, n14522,
         n14523, n14524, n14525, n14526, n14527, n14528, n14529, n14530,
         n14531, n14532, n14533, n14534, n14535, n14536, n14537, n14538,
         n14539, n14540, n14541, n14542, n14543, n14544, n14545, n14546,
         n14547, n14548, n14549, n14550, n14551, n14552, n14553, n14554,
         n14555, n14556, n14557, n14558, n14559, n14560, n14561, n14562,
         n14563, n14564, n14565, n14566, n14567, n14568, n14569, n14570,
         n14571, n14572, n14573, n14574, n14575, n14576, n14577, n14578,
         n14579, n14580, n14581, n14582, n14583, n14584, n14585, n14586,
         n14587, n14588, n14589, n14590, n14591, n14592, n14593, n14594,
         n14595, n14596, n14597, n14598, n14599, n14600, n14601, n14602,
         n14603, n14604, n14605, n14606, n14607, n14608, n14609, n14610,
         n14611, n14612, n14613, n14614, n14615, n14616, n14617, n14618,
         n14619, n14620, n14621, n14622, n14623, n14624, n14625, n14626,
         n14627, n14628, n14629, n14630, n14631, n14632, n14633, n14634,
         n14635, n14636, n14637, n14638, n14639, n14640, n14641, n14642,
         n14643, n14644, n14645, n14646, n14647, n14648, n14649, n14650,
         n14651, n14652, n14653, n14654, n14655, n14656, n14657, n14658,
         n14659, n14660, n14661, n14662, n14663, n14664, n14665, n14666,
         n14667, n14668, n14669, n14670, n14671, n14672, n14673, n14674,
         n14675, n14676, n14677, n14678, n14679, n14680, n14681, n14682,
         n14683, n14684, n14685, n14686, n14687, n14688, n14689, n14690,
         n14691, n14692, n14693, n14694, n14695, n14696, n14697, n14698,
         n14699, n14700, n14701, n14702, n14703, n14704, n14705, n14706,
         n14707, n14708, n14709, n14710, n14711, n14712, n14713, n14714,
         n14715, n14716, n14717, n14718, n14719, n14720, n14721, n14722,
         n14723, n14724, n14725, n14726, n14727, n14728, n14729, n14730,
         n14731, n14732, n14733, n14734, n14735, n14736, n14737, n14738,
         n14739, n14740, n14741, n14742, n14743, n14744, n14745, n14746,
         n14747, n14748, n14749, n14750, n14751, n14752, n14753, n14754,
         n14755, n14756, n14757, n14758, n14759, n14760, n14761, n14762,
         n14763, n14764, n14765, n14766, n14767, n14768, n14769, n14770,
         n14771, n14772, n14773, n14774, n14775, n14776, n14777, n14778,
         n14779, n14780, n14781, n14782, n14783, n14784, n14785, n14786,
         n14787, n14788, n14789, n14790, n14791, n14792, n14793, n14794,
         n14795, n14796, n14797, n14798, n14799, n14800, n14801, n14802,
         n14803, n14804, n14805, n14806, n14807, n14808, n14809, n14810,
         n14811, n14812, n14813, n14814, n14815, n14816, n14817, n14818,
         n14819, n14820, n14821, n14822, n14823, n14824, n14825, n14826,
         n14827, n14828, n14829, n14830, n14831, n14832, n14833, n14834,
         n14835, n14836, n14837, n14838, n14839, n14840, n14841, n14842,
         n14843, n14844, n14845, n14846, n14847, n14848, n14849, n14850,
         n14851, n14852, n14853, n14854, n14855, n14856, n14857, n14858,
         n14859, n14860, n14861, n14862, n14863, n14864, n14865, n14866,
         n14867, n14868, n14869, n14870, n14871, n14872, n14873, n14874,
         n14875, n14876, n14877, n14878, n14879, n14880, n14881, n14882,
         n14883, n14884, n14885, n14886, n14887, n14888, n14889, n14890,
         n14891, n14892, n14893, n14894, n14895, n14896, n14897, n14898,
         n14899, n14900, n14901, n14902, n14903, n14904, n14905, n14906,
         n14907, n14908, n14909, n14910, n14911, n14912, n14913, n14914,
         n14915, n14916, n14917, n14918, n14919, n14920, n14921, n14922,
         n14923, n14924, n14925, n14926, n14927, n14928, n14929, n14930,
         n14931, n14932, n14933, n14934, n14935, n14936, n14937, n14938,
         n14939, n14940, n14941, n14942, n14943, n14944, n14945, n14946,
         n14947, n14948, n14949, n14950, n14951, n14952, n14953, n14954,
         n14955, n14956, n14957, n14958, n14959, n14960, n14961, n14962,
         n14963, n14964, n14965, n14966, n14967, n14968, n14969, n14970,
         n14971, n14972, n14973, n14974, n14975, n14976, n14977, n14978,
         n14979, n14980, n14981, n14982, n14983, n14984, n14985, n14986,
         n14987, n14988, n14989, n14990, n14991, n14992, n14993, n14994,
         n14995, n14996, n14997, n14998, n14999, n15000, n15001, n15002,
         n15003, n15004, n15005, n15006, n15007, n15008, n15009, n15010,
         n15011, n15012, n15013, n15014, n15015, n15016, n15017, n15018,
         n15019, n15020, n15021, n15022, n15023, n15024, n15025, n15026,
         n15027, n15028, n15029, n15030, n15031, n15032, n15033, n15034,
         n15035, n15036, n15037, n15038, n15039, n15040, n15041, n15042,
         n15043, n15044, n15045, n15046, n15047, n15048, n15049, n15050,
         n15051, n15052, n15053, n15054, n15055, n15056, n15057, n15058,
         n15059, n15060, n15061, n15062, n15063, n15064, n15065, n15066,
         n15067, n15068, n15069, n15070, n15071, n15072, n15073, n15074,
         n15075, n15076, n15077, n15078, n15079, n15080, n15081, n15082,
         n15083, n15084, n15085, n15086, n15087, n15088, n15089, n15090,
         n15091, n15092, n15093, n15094, n15095, n15096, n15097, n15098,
         n15099, n15100, n15101, n15102, n15103, n15104, n15105, n15106,
         n15107, n15108, n15109, n15110, n15111, n15112, n15113, n15114,
         n15115, n15116, n15117, n15118, n15119, n15120, n15121, n15122,
         n15123, n15124, n15125, n15126, n15127, n15128, n15129, n15130,
         n15131, n15132, n15133, n15134, n15135, n15136, n15137, n15138,
         n15139, n15140, n15141, n15142, n15143, n15144, n15145, n15146,
         n15147, n15148, n15149, n15150, n15151, n15152, n15153, n15154,
         n15155, n15156, n15157, n15158, n15159, n15160, n15161, n15162,
         n15163, n15164, n15165, n15166, n15167, n15168, n15169, n15170,
         n15171, n15172, n15173, n15174, n15175, n15176, n15177, n15178,
         n15179, n15180, n15181, n15182, n15183, n15184, n15185, n15186,
         n15187, n15188, n15189, n15190, n15191, n15192, n15193, n15194,
         n15195, n15196, n15197, n15198, n15199, n15200, n15201, n15202,
         n15203, n15204, n15205, n15206, n15207, n15208, n15209, n15210,
         n15211, n15212, n15213, n15214, n15215, n15216, n15217, n15218,
         n15219, n15220, n15221, n15222, n15223, n15224, n15225, n15226,
         n15227, n15228, n15229, n15230, n15231, n15232, n15233, n15234,
         n15235, n15236, n15237, n15238, n15239, n15240, n15241, n15242,
         n15243, n15244, n15245, n15246, n15247, n15248, n15249, n15250,
         n15251, n15252, n15253, n15254, n15255, n15256, n15257, n15258,
         n15259, n15260, n15261, n15262, n15263, n15264, n15265, n15266,
         n15267, n15268, n15269, n15270, n15271, n15272, n15273, n15274,
         n15275, n15276, n15277, n15278, n15279, n15280, n15281, n15282,
         n15283, n15284, n15285, n15286, n15287, n15288, n15289, n15290,
         n15291, n15292, n15293, n15294, n15295, n15296, n15297, n15298,
         n15299, n15300, n15301, n15302, n15303, n15304, n15305, n15306,
         n15307, n15308, n15309, n15310, n15311, n15312, n15313, n15314,
         n15315, n15316, n15317, n15318, n15319, n15320, n15321, n15322,
         n15323, n15324, n15325, n15326, n15327, n15328, n15329, n15330,
         n15331, n15332, n15333, n15334, n15335, n15336, n15337, n15338,
         n15339, n15340, n15341, n15342, n15343, n15344, n15345, n15346,
         n15347, n15348, n15349, n15350, n15351, n15352, n15353, n15354,
         n15355, n15356, n15357, n15358, n15359, n15360, n15361, n15362,
         n15363, n15364, n15365, n15366, n15367, n15368, n15369, n15370,
         n15371, n15372, n15373, n15374, n15375, n15376, n15377, n15378,
         n15379, n15380, n15381, n15382, n15383, n15384, n15385, n15386,
         n15387, n15388, n15389, n15390, n15391, n15392, n15393, n15394,
         n15395, n15396, n15397, n15398, n15399, n15400, n15401, n15402,
         n15403, n15404, n15405, n15406, n15407, n15408, n15409, n15410,
         n15411, n15412, n15413, n15414, n15415, n15416, n15417, n15418,
         n15419, n15420, n15421, n15422, n15423, n15424, n15425, n15426,
         n15427, n15428, n15429, n15430, n15431, n15432, n15433, n15434,
         n15435, n15436, n15437, n15438, n15439, n15440, n15441, n15442,
         n15443, n15444, n15445, n15446, n15447, n15448, n15449, n15450,
         n15451, n15452, n15453, n15454, n15455, n15456, n15457, n15458,
         n15459, n15460, n15461, n15462, n15463, n15464, n15465, n15466,
         n15467, n15468, n15469, n15470, n15471, n15472, n15473, n15474,
         n15475, n15476, n15477, n15478, n15479, n15480, n15481, n15482,
         n15483, n15484, n15485, n15486, n15487, n15488, n15489, n15490,
         n15491, n15492, n15493, n15494, n15495, n15496, n15497, n15498,
         n15499, n15500, n15501, n15502, n15503, n15504, n15505, n15506,
         n15507, n15508, n15509, n15510, n15511, n15512, n15513, n15514,
         n15515, n15516, n15517, n15518, n15519, n15520, n15521, n15522,
         n15523, n15524, n15525, n15526, n15527, n15528, n15529, n15530,
         n15531, n15532, n15533, n15534, n15535, n15536, n15537, n15538,
         n15539, n15540, n15541, n15542, n15543, n15544, n15545, n15546,
         n15547, n15548, n15549, n15550, n15551, n15552, n15553, n15554,
         n15555, n15556, n15557, n15558, n15559, n15560, n15561, n15562,
         n15563, n15564, n15565, n15566, n15567, n15568, n15569, n15570,
         n15571, n15572, n15573, n15574, n15575, n15576, n15577, n15578,
         n15579, n15580, n15581, n15582, n15583, n15584, n15585, n15586,
         n15587, n15588, n15589, n15590, n15591, n15592, n15593, n15594,
         n15595, n15596, n15597, n15598, n15599, n15600, n15601, n15602,
         n15603, n15604, n15605, n15606, n15607, n15608, n15609, n15610,
         n15611, n15612, n15613, n15614, n15615, n15616, n15617, n15618,
         n15619, n15620, n15621, n15622, n15623, n15624, n15625, n15626,
         n15627, n15628, n15629, n15630, n15631, n15632, n15633, n15634,
         n15635, n15636, n15637, n15638, n15639, n15640, n15641, n15642,
         n15643, n15644, n15645, n15646, n15647, n15648, n15649, n15650,
         n15651, n15652, n15653, n15654, n15655, n15656, n15657, n15658,
         n15659, n15660, n15661, n15662, n15663, n15664, n15665, n15666,
         n15667, n15668, n15669, n15670, n15671, n15672, n15673, n15674,
         n15675, n15676, n15677, n15678, n15679, n15680, n15681, n15682,
         n15683, n15684, n15685, n15686, n15687, n15688, n15689, n15690,
         n15691, n15692, n15693, n15694, n15695, n15696, n15697, n15698,
         n15699, n15700, n15701, n15702, n15703, n15704, n15705, n15706,
         n15707, n15708, n15709, n15710, n15711, n15712, n15713, n15714,
         n15715, n15716, n15717, n15718, n15719, n15720, n15721, n15722,
         n15723, n15724, n15725, n15726, n15727, n15728, n15729, n15730,
         n15731, n15732, n15733, n15734, n15735, n15736, n15737, n15738,
         n15739, n15740, n15741, n15742, n15743, n15744, n15745, n15746,
         n15747, n15748, n15749, n15750, n15751, n15752, n15753, n15754,
         n15755, n15756, n15757, n15758, n15759, n15760, n15761, n15762,
         n15763, n15764, n15765, n15766, n15767, n15768, n15769, n15770,
         n15771, n15772, n15773, n15774, n15775, n15776, n15777, n15778,
         n15779, n15780, n15781, n15782, n15783, n15784, n15785, n15786,
         n15787, n15788, n15789, n15790, n15791, n15792, n15793, n15794,
         n15795, n15796, n15797, n15798, n15799, n15800, n15801, n15802,
         n15803, n15804, n15805, n15806, n15807, n15808, n15809, n15810,
         n15811, n15812, n15813, n15814, n15815, n15816, n15817, n15818,
         n15819, n15820, n15821, n15822, n15823, n15824, n15825, n15826,
         n15827, n15828, n15829, n15830, n15831, n15832, n15833, n15834,
         n15835, n15836, n15837, n15838, n15839, n15840, n15841, n15842,
         n15843, n15844, n15845, n15846, n15847, n15848, n15849, n15850,
         n15851, n15852, n15853, n15854, n15855, n15856, n15857, n15858,
         n15859, n15860, n15861, n15862, n15863, n15864, n15865, n15866,
         n15867, n15868, n15869, n15870, n15871, n15872, n15873, n15874,
         n15875, n15876, n15877, n15878, n15879, n15880, n15881, n15882,
         n15883, n15884, n15885, n15886, n15887, n15888, n15889, n15890,
         n15891, n15892, n15893, n15894, n15895, n15896, n15897, n15898,
         n15899, n15900, n15901, n15902, n15903, n15904, n15905, n15906,
         n15907, n15908, n15909, n15910, n15911, n15912, n15913, n15914,
         n15915, n15916, n15917, n15918, n15919, n15920, n15921, n15922,
         n15923, n15924, n15925, n15926, n15927, n15928, n15929, n15930,
         n15931, n15932, n15933, n15934, n15935, n15936, n15937, n15938,
         n15939, n15940, n15941, n15942, n15943, n15944, n15945, n15946,
         n15947, n15948, n15949, n15950, n15951, n15952, n15953, n15954,
         n15955, n15956, n15957, n15958, n15959, n15960, n15961, n15962,
         n15963, n15964, n15965, n15966, n15967, n15968, n15969, n15970,
         n15971, n15972, n15973, n15974, n15975, n15976, n15977, n15978,
         n15979, n15980, n15981, n15982, n15983, n15984, n15985, n15986,
         n15987, n15988, n15989, n15990, n15991, n15992, n15993, n15994,
         n15995, n15996, n15997, n15998, n15999, n16000, n16001, n16002,
         n16003, n16004, n16005, n16006, n16007, n16008, n16009, n16010,
         n16011, n16012, n16013, n16014, n16015, n16016, n16017, n16018,
         n16019, n16020, n16021, n16022, n16023, n16024, n16025, n16026,
         n16027, n16028, n16029, n16030, n16031, n16032, n16033, n16034,
         n16035, n16036, n16037, n16038, n16039, n16040, n16041, n16042,
         n16043, n16044, n16045, n16046, n16047, n16048, n16049, n16050,
         n16051, n16052, n16053, n16054, n16055, n16056, n16057, n16058,
         n16059, n16060, n16061, n16062, n16063, n16064, n16065, n16066,
         n16067, n16068, n16069, n16070, n16071, n16072, n16073, n16074,
         n16075, n16076, n16077, n16078, n16079, n16080, n16081, n16082,
         n16083, n16084, n16085, n16086, n16087, n16088, n16089, n16090,
         n16091, n16092, n16093, n16094, n16095, n16096, n16097, n16098,
         n16099, n16100, n16101, n16102, n16103, n16104, n16105, n16106,
         n16107, n16108, n16109, n16110, n16111, n16112, n16113, n16114,
         n16115, n16116, n16117, n16118, n16119, n16120, n16121, n16122,
         n16123, n16124, n16125, n16126, n16127, n16128, n16129, n16130,
         n16131, n16132, n16133, n16134, n16135, n16136, n16137, n16138,
         n16139, n16140, n16141, n16142, n16143, n16144, n16145, n16146,
         n16147, n16148, n16149, n16150, n16151, n16152, n16153, n16154,
         n16155, n16156, n16157, n16158, n16159, n16160, n16161, n16162,
         n16163, n16164, n16165, n16166, n16167, n16168, n16169, n16170,
         n16171, n16172, n16173, n16174, n16175, n16176, n16177, n16178,
         n16179, n16180, n16181, n16182, n16183, n16184, n16185, n16186,
         n16187, n16188, n16189, n16190, n16191, n16192, n16193, n16194,
         n16195, n16196, n16197, n16198, n16199, n16200, n16201, n16202,
         n16203, n16204, n16205, n16206, n16207, n16208, n16209, n16210,
         n16211, n16212, n16213, n16214, n16215, n16216, n16217, n16218,
         n16219, n16220, n16221, n16222, n16223, n16224, n16225, n16226,
         n16227, n16228, n16229, n16230, n16231, n16232, n16233, n16234,
         n16235, n16236, n16237, n16238, n16239, n16240, n16241, n16242,
         n16243, n16244, n16245, n16246, n16247, n16248, n16249, n16250,
         n16251, n16252, n16253, n16254, n16255, n16256, n16257, n16258,
         n16259, n16260, n16261, n16262, n16263, n16264, n16265, n16266,
         n16267, n16268, n16269, n16270, n16271, n16272, n16273, n16274,
         n16275, n16276, n16277, n16278, n16279, n16280, n16281, n16282,
         n16283, n16284, n16285, n16286, n16287, n16288, n16289, n16290,
         n16291, n16292, n16293, n16294, n16295, n16296, n16297, n16298,
         n16299, n16300, n16301, n16302, n16303, n16304, n16305, n16306,
         n16307, n16308, n16309, n16310, n16311, n16312, n16313, n16314,
         n16315, n16316, n16317, n16318, n16319, n16320, n16321, n16322,
         n16323, n16324, n16325, n16326, n16327, n16328, n16329, n16330,
         n16331, n16332, n16333, n16334, n16335, n16336, n16337, n16338,
         n16339, n16340, n16341, n16342, n16343, n16344, n16345, n16346,
         n16347, n16348, n16349, n16350, n16351, n16352, n16353, n16354,
         n16355, n16356, n16357, n16358, n16359, n16360, n16361, n16362,
         n16363, n16364, n16365, n16366, n16367, n16368, n16369, n16370,
         n16371, n16372, n16373, n16374, n16375, n16376, n16377, n16378,
         n16379, n16380, n16381, n16382, n16383, n16384, n16385, n16386,
         n16387, n16388, n16389, n16390, n16391, n16392, n16393, n16394,
         n16395, n16396, n16397, n16398, n16399, n16400, n16401, n16402,
         n16403, n16404, n16405, n16406, n16407, n16408, n16409, n16410,
         n16411, n16412, n16413, n16414, n16415, n16416, n16417, n16418,
         n16419, n16420, n16421, n16422, n16423, n16424, n16425, n16426,
         n16427, n16428, n16429, n16430, n16431, n16432, n16433, n16434,
         n16435, n16436, n16437, n16438, n16439, n16440, n16441, n16442,
         n16443, n16444, n16445, n16446, n16447, n16448, n16449, n16450,
         n16451, n16452, n16453, n16454, n16455, n16456, n16457, n16458,
         n16459, n16460, n16461, n16462, n16463, n16464, n16465, n16466,
         n16467, n16468, n16469, n16470, n16471, n16472, n16473, n16474,
         n16475, n16476, n16477, n16478, n16479, n16480, n16481, n16482,
         n16483, n16484, n16485, n16486, n16487, n16488, n16489, n16490,
         n16491, n16492, n16493, n16494, n16495, n16496, n16497, n16498,
         n16499, n16500, n16501, n16502, n16503, n16504, n16505, n16506,
         n16507, n16508, n16509, n16510, n16511, n16512, n16513, n16514,
         n16515, n16516, n16517, n16518, n16519, n16520, n16521, n16522,
         n16523, n16524, n16525, n16526, n16527, n16528, n16529, n16530,
         n16531, n16532, n16533, n16534, n16535, n16536, n16537, n16538,
         n16539, n16540, n16541, n16542, n16543, n16544, n16545, n16546,
         n16547, n16548, n16549, n16550, n16551, n16552, n16553, n16554,
         n16555, n16556, n16557, n16558, n16559, n16560, n16561, n16562,
         n16563, n16564, n16565, n16566, n16567, n16568, n16569, n16570,
         n16571, n16572, n16573, n16574, n16575, n16576, n16577, n16578,
         n16579, n16580, n16581, n16582, n16583, n16584, n16585, n16586,
         n16587, n16588, n16589, n16590, n16591, n16592, n16593, n16594,
         n16595, n16596, n16597, n16598, n16599, n16600, n16601, n16602,
         n16603, n16604, n16605, n16606, n16607, n16608, n16609, n16610,
         n16611, n16612, n16613, n16614, n16615, n16616, n16617, n16618,
         n16619, n16620, n16621, n16622, n16623, n16624, n16625, n16626,
         n16627, n16628, n16629, n16630, n16631, n16632, n16633, n16634,
         n16635, n16636, n16637, n16638, n16639, n16640, n16641, n16642,
         n16643, n16644, n16645, n16646, n16647, n16648, n16649, n16650,
         n16651, n16652, n16653, n16654, n16655, n16656, n16657, n16658,
         n16659, n16660, n16661, n16662, n16663, n16664, n16665, n16666,
         n16667, n16668, n16669, n16670, n16671, n16672, n16673, n16674,
         n16675, n16676, n16677, n16678, n16679, n16680, n16681, n16682,
         n16683, n16684, n16685, n16686, n16687, n16688, n16689, n16690,
         n16691, n16692, n16693, n16694, n16695, n16696, n16697, n16698,
         n16699, n16700, n16701, n16702, n16703, n16704, n16705, n16706,
         n16707, n16708, n16709, n16710, n16711, n16712, n16713, n16714,
         n16715, n16716, n16717, n16718, n16719, n16720, n16721, n16722,
         n16723, n16724, n16725, n16726, n16727, n16728, n16729, n16730,
         n16731, n16732, n16733, n16734, n16735, n16736, n16737, n16738,
         n16739, n16740, n16741, n16742, n16743, n16744, n16745, n16746,
         n16747, n16748, n16749, n16750, n16751, n16752, n16753, n16754,
         n16755, n16756, n16757, n16758, n16759, n16760, n16761, n16762,
         n16763, n16764, n16765, n16766, n16767, n16768, n16769, n16770,
         n16771, n16772, n16773, n16774, n16775, n16776, n16777, n16778,
         n16779, n16780, n16781, n16782, n16783, n16784, n16785, n16786,
         n16787, n16788, n16789, n16790, n16791, n16792, n16793, n16794,
         n16795, n16796, n16797, n16798, n16799, n16800, n16801, n16802,
         n16803, n16804, n16805, n16806, n16807, n16808, n16809, n16810,
         n16811, n16812, n16813, n16814, n16815, n16816, n16817, n16818,
         n16819, n16820, n16821, n16822, n16823, n16824, n16825, n16826,
         n16827, n16828, n16829, n16830, n16831, n16832, n16833, n16834,
         n16835, n16836, n16837, n16838, n16839, n16840, n16841, n16842,
         n16843, n16844, n16845, n16846, n16847, n16848, n16849, n16850,
         n16851, n16852, n16853, n16854, n16855, n16856, n16857, n16858,
         n16859, n16860, n16861, n16862, n16863, n16864, n16865, n16866,
         n16867, n16868, n16869, n16870, n16871, n16872, n16873, n16874,
         n16875, n16876, n16877, n16878, n16879, n16880, n16881, n16882,
         n16883, n16884, n16885, n16886, n16887, n16888, n16889, n16890,
         n16891, n16892, n16893, n16894, n16895, n16896, n16897, n16898,
         n16899, n16900, n16901, n16902, n16903, n16904, n16905, n16906,
         n16907, n16908, n16909, n16910, n16911, n16912, n16913, n16914,
         n16915, n16916, n16917, n16918, n16919, n16920, n16921, n16922,
         n16923, n16924, n16925, n16926, n16927, n16928, n16929, n16930,
         n16931, n16932, n16933, n16934, n16935, n16936, n16937, n16938,
         n16939, n16940, n16941, n16942, n16943, n16944, n16945, n16946,
         n16947, n16948, n16949, n16950, n16951, n16952, n16953, n16954,
         n16955, n16956, n16957, n16958, n16959, n16960, n16961, n16962,
         n16963, n16964, n16965, n16966, n16967, n16968, n16969, n16970,
         n16971, n16972, n16973, n16974, n16975, n16976, n16977, n16978,
         n16979, n16980, n16981, n16982, n16983, n16984, n16985, n16986,
         n16987, n16988, n16989, n16990, n16991, n16992, n16993, n16994,
         n16995, n16996, n16997, n16998, n16999, n17000, n17001, n17002,
         n17003, n17004, n17005, n17006, n17007, n17008, n17009, n17010,
         n17011, n17012, n17013, n17014, n17015, n17016, n17017, n17018,
         n17019, n17020, n17021, n17022, n17023, n17024, n17025, n17026,
         n17027, n17028, n17029, n17030, n17031, n17032, n17033, n17034,
         n17035, n17036, n17037, n17038, n17039, n17040, n17041, n17042,
         n17043, n17044, n17045, n17046, n17047, n17048, n17049, n17050,
         n17051, n17052, n17053, n17054, n17055, n17056, n17057, n17058,
         n17059, n17060, n17061, n17062, n17063, n17064, n17065, n17066,
         n17067, n17068, n17069, n17070, n17071, n17072, n17073, n17074,
         n17075, n17076, n17077, n17078, n17079, n17080, n17081, n17082,
         n17083, n17084, n17085, n17086, n17087, n17088, n17089, n17090,
         n17091, n17092, n17093, n17094, n17095, n17096, n17097, n17098,
         n17099, n17100, n17101, n17102, n17103, n17104, n17105, n17106,
         n17107, n17108, n17109, n17110, n17111, n17112, n17113, n17114,
         n17115, n17116, n17117, n17118, n17119, n17120, n17121, n17122,
         n17123, n17124, n17125, n17126, n17127, n17128, n17129, n17130,
         n17131, n17132, n17133, n17134, n17135, n17136, n17137, n17138,
         n17139, n17140, n17141, n17142, n17143, n17144, n17145, n17146,
         n17147, n17148, n17149, n17150, n17151, n17152, n17153, n17154,
         n17155, n17156, n17157, n17158, n17159, n17160, n17161, n17162,
         n17163, n17164, n17165, n17166, n17167, n17168, n17169, n17170,
         n17171, n17172, n17173, n17174, n17175, n17176, n17177, n17178,
         n17179, n17180, n17181, n17182, n17183, n17184, n17185, n17186,
         n17187, n17188, n17189, n17190, n17191, n17192, n17193, n17194,
         n17195, n17196, n17197, n17198, n17199, n17200, n17201, n17202,
         n17203, n17204, n17205, n17206, n17207, n17208, n17209, n17210,
         n17211, n17212, n17213, n17214, n17215, n17216, n17217, n17218,
         n17219, n17220, n17221, n17222, n17223, n17224, n17225, n17226,
         n17227, n17228, n17229, n17230, n17231, n17232, n17233, n17234,
         n17235, n17236, n17237, n17238, n17239, n17240, n17241, n17242,
         n17243, n17244, n17245, n17246, n17247, n17248, n17249, n17250,
         n17251, n17252, n17253, n17254, n17255, n17256, n17257, n17258,
         n17259, n17260, n17261, n17262, n17263, n17264, n17265, n17266,
         n17267, n17268, n17269, n17270, n17271, n17272, n17273, n17274,
         n17275, n17276, n17277, n17278, n17279, n17280, n17281, n17282,
         n17283, n17284, n17285, n17286, n17287, n17288, n17289, n17290,
         n17291, n17292, n17293, n17294, n17295, n17296, n17297, n17298,
         n17299, n17300, n17301, n17302, n17303, n17304, n17305, n17306,
         n17307, n17308, n17309, n17310, n17311, n17312, n17313, n17314,
         n17315, n17316, n17317, n17318, n17319, n17320, n17321, n17322,
         n17323, n17324, n17325, n17326, n17327, n17328, n17329, n17330,
         n17331, n17332, n17333, n17334, n17335, n17336, n17337, n17338,
         n17339, n17340, n17341, n17342, n17343, n17344, n17345, n17346,
         n17347, n17348, n17349, n17350, n17351, n17352, n17353, n17354,
         n17355, n17356, n17357, n17358, n17359, n17360, n17361, n17362,
         n17363, n17364, n17365, n17366, n17367, n17368, n17369, n17370,
         n17371, n17372, n17373, n17374, n17375, n17376, n17377, n17378,
         n17379, n17380, n17381, n17382, n17383, n17384, n17385, n17386,
         n17387, n17388, n17389, n17390, n17391, n17392, n17393, n17394,
         n17395, n17396, n17397, n17398, n17399, n17400, n17401, n17402,
         n17403, n17404, n17405, n17406, n17407, n17408, n17409, n17410,
         n17411, n17412, n17413, n17414, n17415, n17416, n17417, n17418,
         n17419, n17420, n17421, n17422, n17423, n17424, n17425, n17426,
         n17427, n17428, n17429, n17430, n17431, n17432, n17433, n17434,
         n17435, n17436, n17437, n17438, n17439, n17440, n17441, n17442,
         n17443, n17444, n17445, n17446, n17447, n17448, n17449, n17450,
         n17451, n17452, n17453, n17454, n17455, n17456, n17457, n17458,
         n17459, n17460, n17461, n17462, n17463, n17464, n17465, n17466,
         n17467, n17468, n17469, n17470, n17471, n17472, n17473, n17474,
         n17475, n17476, n17477, n17478, n17479, n17480, n17481, n17482,
         n17483, n17484, n17485, n17486, n17487, n17488, n17489, n17490,
         n17491, n17492, n17493, n17494, n17495, n17496, n17497, n17498,
         n17499, n17500, n17501, n17502, n17503, n17504, n17505, n17506,
         n17507, n17508, n17509, n17510, n17511, n17512, n17513, n17514,
         n17515, n17516, n17517, n17518, n17519, n17520, n17521, n17522,
         n17523, n17524, n17525, n17526, n17527, n17528, n17529, n17530,
         n17531, n17532, n17533, n17534, n17535, n17536, n17537, n17538,
         n17539, n17540, n17541, n17542, n17543, n17544, n17545, n17546,
         n17547, n17548, n17549, n17550, n17551, n17552, n17553, n17554,
         n17555, n17556, n17557, n17558, n17559, n17560, n17561, n17562,
         n17563, n17564, n17565, n17566, n17567, n17568, n17569, n17570,
         n17571, n17572, n17573, n17574, n17575, n17576, n17577, n17578,
         n17579, n17580, n17581, n17582, n17583, n17584, n17585, n17586,
         n17587, n17588, n17589, n17590, n17591, n17592, n17593, n17594,
         n17595, n17596, n17597, n17598, n17599, n17600, n17601, n17602,
         n17603, n17604, n17605, n17606, n17607, n17608, n17609, n17610,
         n17611, n17612, n17613, n17614, n17615, n17616, n17617, n17618,
         n17619, n17620, n17621, n17622, n17623, n17624, n17625, n17626,
         n17627, n17628, n17629, n17630, n17631, n17632, n17633, n17634,
         n17635, n17636, n17637, n17638, n17639, n17640, n17641, n17642,
         n17643, n17644, n17645, n17646, n17647, n17648, n17649, n17650,
         n17651, n17652, n17653, n17654, n17655, n17656, n17657, n17658,
         n17659, n17660, n17661, n17662, n17663, n17664, n17665, n17666,
         n17667, n17668, n17669, n17670, n17671, n17672, n17673, n17674,
         n17675, n17676, n17677, n17678, n17679, n17680, n17681, n17682,
         n17683, n17684, n17685, n17686, n17687, n17688, n17689, n17690,
         n17691, n17692, n17693, n17694, n17695, n17696, n17697, n17698,
         n17699, n17700, n17701, n17702, n17703, n17704, n17705, n17706,
         n17707, n17708, n17709, n17710, n17711, n17712, n17713, n17714,
         n17715, n17716, n17717, n17718, n17719, n17720, n17721, n17722,
         n17723, n17724, n17725, n17726, n17727, n17728, n17729, n17730,
         n17731, n17732, n17733, n17734, n17735, n17736, n17737, n17738,
         n17739, n17740, n17741, n17742, n17743, n17744, n17745, n17746,
         n17747, n17748, n17749, n17750, n17751, n17752, n17753, n17754,
         n17755, n17756, n17757, n17758, n17759, n17760, n17761, n17762,
         n17763, n17764, n17765, n17766, n17767, n17768, n17769, n17770,
         n17771, n17772, n17773, n17774, n17775, n17776, n17777, n17778,
         n17779, n17780, n17781, n17782, n17783, n17784, n17785, n17786,
         n17787, n17788, n17789, n17790, n17791, n17792, n17793, n17794,
         n17795, n17796, n17797, n17798, n17799, n17800, n17801, n17802,
         n17803, n17804, n17805, n17806, n17807, n17808, n17809, n17810,
         n17811, n17812, n17813, n17814, n17815, n17816, n17817, n17818,
         n17819, n17820, n17821, n17822, n17823, n17824, n17825, n17826,
         n17827, n17828, n17829, n17830, n17831, n17832, n17833, n17834,
         n17835, n17836, n17837, n17838, n17839, n17840, n17841, n17842,
         n17843, n17844, n17845, n17846, n17847, n17848, n17849, n17850,
         n17851, n17852, n17853, n17854, n17855, n17856, n17857, n17858,
         n17859, n17860, n17861, n17862, n17863, n17864, n17865, n17866,
         n17867, n17868, n17869, n17870, n17871, n17872, n17873, n17874,
         n17875, n17876, n17877, n17878, n17879, n17880, n17881, n17882,
         n17883, n17884, n17885, n17886, n17887, n17888, n17889, n17890,
         n17891, n17892, n17893, n17894, n17895, n17896, n17897, n17898,
         n17899, n17900, n17901, n17902, n17903, n17904, n17905, n17906,
         n17907, n17908, n17909, n17910, n17911, n17912, n17913, n17914,
         n17915, n17916, n17917, n17918, n17919, n17920, n17921, n17922,
         n17923, n17924, n17925, n17926, n17927, n17928, n17929, n17930,
         n17931, n17932, n17933, n17934, n17935, n17936, n17937, n17938,
         n17939, n17940, n17941, n17942, n17943, n17944, n17945, n17946,
         n17947, n17948, n17949, n17950, n17951, n17952, n17953, n17954,
         n17955, n17956, n17957, n17958, n17959, n17960, n17961, n17962,
         n17963, n17964, n17965, n17966, n17967, n17968, n17969, n17970,
         n17971, n17972, n17973, n17974, n17975, n17976, n17977, n17978,
         n17979, n17980, n17981, n17982, n17983, n17984, n17985, n17986,
         n17987, n17988, n17989, n17990, n17991, n17992, n17993, n17994,
         n17995, n17996, n17997, n17998, n17999, n18000, n18001, n18002,
         n18003, n18004, n18005, n18006, n18007, n18008, n18009, n18010,
         n18011, n18012, n18013, n18014, n18015, n18016, n18017, n18018,
         n18019, n18020, n18021, n18022, n18023, n18024, n18025, n18026,
         n18027, n18028, n18029, n18030, n18031, n18032, n18033, n18034,
         n18035, n18036, n18037, n18038, n18039, n18040, n18041, n18042,
         n18043, n18044, n18045, n18046, n18047, n18048, n18049, n18050,
         n18051, n18052, n18053, n18054, n18055, n18056, n18057, n18058,
         n18059, n18060, n18061, n18062, n18063, n18064, n18065, n18066,
         n18067, n18068, n18069, n18070, n18071, n18072, n18073, n18074,
         n18075, n18076, n18077, n18078, n18079, n18080, n18081, n18082,
         n18083, n18084, n18085, n18086, n18087, n18088, n18089, n18090,
         n18091, n18092, n18093, n18094, n18095, n18096, n18097, n18098,
         n18099, n18100, n18101, n18102, n18103, n18104, n18105, n18106,
         n18107, n18108, n18109, n18110, n18111, n18112, n18113, n18114,
         n18115, n18116, n18117, n18118, n18119, n18120, n18121, n18122,
         n18123, n18124, n18125, n18126, n18127, n18128, n18129, n18130,
         n18131, n18132, n18133, n18134, n18135, n18136, n18137, n18138,
         n18139, n18140, n18141, n18142, n18143, n18144, n18145, n18146,
         n18147, n18148, n18149, n18150, n18151, n18152, n18153, n18154,
         n18155, n18156, n18157, n18158, n18159, n18160, n18161, n18162,
         n18163, n18164, n18165, n18166, n18167, n18168, n18169, n18170,
         n18171, n18172, n18173, n18174, n18175, n18176, n18177, n18178,
         n18179, n18180, n18181, n18182, n18183, n18184, n18185, n18186,
         n18187, n18188, n18189, n18190, n18191, n18192, n18193, n18194,
         n18195, n18196, n18197, n18198, n18199, n18200, n18201, n18202,
         n18203, n18204, n18205, n18206, n18207, n18208, n18209, n18210,
         n18211, n18212, n18213, n18214, n18215, n18216, n18217, n18218,
         n18219, n18220, n18221, n18222, n18223, n18224, n18225, n18226,
         n18227, n18228, n18229, n18230, n18231, n18232, n18233, n18234,
         n18235, n18236, n18237, n18238, n18239, n18240, n18241, n18242,
         n18243, n18244, n18245, n18246, n18247, n18248, n18249, n18250,
         n18251, n18252, n18253, n18254, n18255, n18256, n18257, n18258,
         n18259, n18260, n18261, n18262, n18263, n18264, n18265, n18266,
         n18267, n18268, n18269, n18270, n18271, n18272, n18273, n18274,
         n18275, n18276, n18277, n18278, n18279, n18280, n18281, n18282,
         n18283, n18284, n18285, n18286, n18287, n18288, n18289, n18290,
         n18291, n18292, n18293, n18294, n18295, n18296, n18297, n18298,
         n18299, n18300, n18301, n18302, n18303, n18304, n18305, n18306,
         n18307, n18308, n18309, n18310, n18311, n18312, n18313, n18314,
         n18315, n18316, n18317, n18318, n18319, n18320, n18321, n18322,
         n18323, n18324, n18325, n18326, n18327, n18328, n18329, n18330,
         n18331, n18332, n18333, n18334, n18335, n18336, n18337, n18338,
         n18339, n18340, n18341, n18342, n18343, n18344, n18345, n18346,
         n18347, n18348, n18349, n18350, n18351, n18352, n18353, n18354,
         n18355, n18356, n18357, n18358, n18359, n18360, n18361, n18362,
         n18363, n18364, n18365, n18366, n18367, n18368, n18369, n18370,
         n18371, n18372, n18373, n18374, n18375, n18376, n18377, n18378,
         n18379, n18380, n18381, n18382, n18383, n18384, n18385, n18386,
         n18387, n18388, n18389, n18390, n18391, n18392, n18393, n18394,
         n18395, n18396, n18397, n18398, n18399, n18400, n18401, n18402,
         n18403, n18404, n18405, n18406, n18407, n18408, n18409, n18410,
         n18411, n18412, n18413, n18414, n18415, n18416, n18417, n18418,
         n18419, n18420, n18421, n18422, n18423, n18424, n18425, n18426,
         n18427, n18428, n18429, n18430, n18431, n18432, n18433, n18434,
         n18435, n18436, n18437, n18438, n18439, n18440, n18441, n18442,
         n18443, n18444, n18445, n18446, n18447, n18448, n18449, n18450,
         n18451, n18452, n18453, n18454, n18455, n18456, n18457, n18458,
         n18459, n18460, n18461, n18462, n18463, n18464, n18465, n18466,
         n18467, n18468, n18469, n18470, n18471, n18472, n18473, n18474,
         n18475, n18476, n18477, n18478, n18479, n18480, n18481, n18482,
         n18483, n18484, n18485, n18486, n18487, n18488, n18489, n18490,
         n18491, n18492, n18493, n18494, n18495, n18496, n18497, n18498,
         n18499, n18500, n18501, n18502, n18503, n18504, n18505, n18506,
         n18507, n18508, n18509, n18510, n18511, n18512, n18513, n18514,
         n18515, n18516, n18517, n18518, n18519, n18520, n18521, n18522,
         n18523, n18524, n18525, n18526, n18527, n18528, n18529, n18530,
         n18531, n18532, n18533, n18534, n18535, n18536, n18537, n18538,
         n18539, n18540, n18541, n18542, n18543, n18544, n18545, n18546,
         n18547, n18548, n18549, n18550, n18551, n18552, n18553, n18554,
         n18555, n18556, n18557, n18558, n18559, n18560, n18561, n18562,
         n18563, n18564, n18565, n18566, n18567, n18568, n18569, n18570,
         n18571, n18572, n18573, n18574, n18575, n18576, n18577, n18578,
         n18579, n18580, n18581, n18582, n18583, n18584, n18585, n18586,
         n18587, n18588, n18589, n18590, n18591, n18592, n18593, n18594,
         n18595, n18596, n18597, n18598, n18599, n18600, n18601, n18602,
         n18603, n18604, n18605, n18606, n18607, n18608, n18609, n18610,
         n18611, n18612, n18613, n18614, n18615, n18616, n18617, n18618,
         n18619, n18620, n18621, n18622, n18623, n18624, n18625, n18626,
         n18627, n18628, n18629, n18630, n18631, n18632, n18633, n18634,
         n18635, n18636, n18637, n18638, n18639, n18640, n18641, n18642,
         n18643, n18644, n18645, n18646, n18647, n18648, n18649, n18650,
         n18651, n18652, n18653, n18654, n18655, n18656, n18657, n18658,
         n18659, n18660, n18661, n18662, n18663, n18664, n18665, n18666,
         n18667, n18668, n18669, n18670, n18671, n18672, n18673, n18674,
         n18675, n18676, n18677, n18678, n18679, n18680, n18681, n18682,
         n18683, n18684, n18685, n18686, n18687, n18688, n18689, n18690,
         n18691, n18692, n18693, n18694, n18695, n18696, n18697, n18698,
         n18699, n18700, n18701, n18702, n18703, n18704, n18705, n18706,
         n18707, n18708, n18709, n18710, n18711, n18712, n18713, n18714,
         n18715, n18716, n18717, n18718, n18719, n18720, n18721, n18722,
         n18723, n18724, n18725, n18726, n18727, n18728, n18729, n18730,
         n18731, n18732, n18733, n18734, n18735, n18736, n18737, n18738,
         n18739, n18740, n18741, n18742, n18743, n18744, n18745, n18746,
         n18747, n18748, n18749, n18750, n18751, n18752, n18753, n18754,
         n18755, n18756, n18757, n18758, n18759, n18760, n18761, n18762,
         n18763, n18764, n18765, n18766, n18767, n18768, n18769, n18770,
         n18771, n18772, n18773, n18774, n18775, n18776, n18777, n18778,
         n18779, n18780, n18781, n18782, n18783, n18784, n18785, n18786,
         n18787, n18788, n18789, n18790, n18791, n18792, n18793, n18794,
         n18795, n18796, n18797, n18798, n18799, n18800, n18801, n18802,
         n18803, n18804, n18805, n18806, n18807, n18808, n18809, n18810,
         n18811, n18812, n18813, n18814, n18815, n18816, n18817, n18818,
         n18819, n18820, n18821, n18822, n18823, n18824, n18825, n18826,
         n18827, n18828, n18829, n18830, n18831, n18832, n18833, n18834,
         n18835, n18836, n18837, n18838, n18839, n18840, n18841, n18842,
         n18843, n18844, n18845, n18846, n18847, n18848, n18849, n18850,
         n18851, n18852, n18853, n18854, n18855, n18856, n18857, n18858,
         n18859, n18860, n18861, n18862, n18863, n18864, n18865, n18866,
         n18867, n18868, n18869, n18870, n18871, n18872, n18873, n18874,
         n18875, n18876, n18877, n18878, n18879, n18880, n18881, n18882,
         n18883, n18884, n18885, n18886, n18887, n18888, n18889, n18890,
         n18891, n18892, n18893, n18894, n18895, n18896, n18897, n18898,
         n18899, n18900, n18901, n18902, n18903, n18904, n18905, n18906,
         n18907, n18908, n18909, n18910, n18911, n18912, n18913, n18914,
         n18915, n18916, n18917, n18918, n18919, n18920, n18921, n18922,
         n18923, n18924, n18925, n18926, n18927, n18928, n18929, n18930,
         n18931, n18932, n18933, n18934, n18935, n18936, n18937, n18938,
         n18939, n18940, n18941, n18942, n18943, n18944, n18945, n18946,
         n18947, n18948, n18949, n18950, n18951, n18952, n18953, n18954,
         n18955, n18956, n18957, n18958, n18959, n18960, n18961, n18962,
         n18963, n18964, n18965, n18966, n18967, n18968, n18969, n18970,
         n18971, n18972, n18973, n18974, n18975, n18976, n18977, n18978,
         n18979, n18980, n18981, n18982, n18983, n18984, n18985, n18986,
         n18987, n18988, n18989, n18990, n18991, n18992, n18993, n18994,
         n18995, n18996, n18997, n18998, n18999, n19000, n19001, n19002,
         n19003, n19004, n19005, n19006, n19007, n19008, n19009, n19010,
         n19011, n19012, n19013, n19014, n19015, n19016, n19017, n19018,
         n19019, n19020, n19021, n19022, n19023, n19024, n19025, n19026,
         n19027, n19028, n19029, n19030, n19031, n19032, n19033, n19034,
         n19035, n19036, n19037, n19038, n19039, n19040, n19041, n19042,
         n19043, n19044, n19045, n19046, n19047, n19048, n19049, n19050,
         n19051, n19052, n19053, n19054, n19055, n19056, n19057, n19058,
         n19059, n19060, n19061, n19062, n19063, n19064, n19065, n19066,
         n19067, n19068, n19069, n19070, n19071, n19072, n19073, n19074,
         n19075, n19076, n19077, n19078, n19079, n19080, n19081, n19082,
         n19083, n19084, n19085, n19086, n19087, n19088, n19089, n19090,
         n19091, n19092, n19093, n19094, n19095, n19096, n19097, n19098,
         n19099, n19100, n19101, n19102, n19103, n19104, n19105, n19106,
         n19107, n19108, n19109, n19110, n19111, n19112, n19113, n19114,
         n19115, n19116, n19117, n19118, n19119, n19120, n19121, n19122,
         n19123, n19124, n19125, n19126, n19127, n19128, n19129, n19130,
         n19131, n19132, n19133, n19134, n19135, n19136, n19137, n19138,
         n19139, n19140, n19141, n19142, n19143, n19144, n19145, n19146,
         n19147, n19148, n19149, n19150, n19151, n19152, n19153, n19154,
         n19155, n19156, n19157, n19158, n19159, n19160, n19161, n19162,
         n19163, n19164, n19165, n19166, n19167, n19168, n19169, n19170,
         n19171, n19172, n19173, n19174, n19175, n19176, n19177, n19178,
         n19179, n19180, n19181, n19182, n19183, n19184, n19185, n19186,
         n19187, n19188, n19189, n19190, n19191, n19192, n19193, n19194,
         n19195, n19196, n19197, n19198, n19199, n19200, n19201, n19202,
         n19203, n19204, n19205, n19206, n19207, n19208, n19209, n19210,
         n19211, n19212, n19213, n19214, n19215, n19216, n19217, n19218,
         n19219, n19220, n19221, n19222, n19223, n19224, n19225, n19226,
         n19227, n19228, n19229, n19230, n19231, n19232, n19233, n19234,
         n19235, n19236, n19237, n19238, n19239, n19240, n19241, n19242,
         n19243, n19244, n19245, n19246, n19247, n19248, n19249, n19250,
         n19251, n19252, n19253, n19254, n19255, n19256, n19257, n19258,
         n19259, n19260, n19261, n19262, n19263, n19264, n19265, n19266,
         n19267, n19268, n19269, n19270, n19271, n19272, n19273, n19274,
         n19275, n19276, n19277, n19278, n19279, n19280, n19281, n19282,
         n19283, n19284, n19285, n19286, n19287, n19288, n19289, n19290,
         n19291, n19292, n19293, n19294, n19295, n19296, n19297, n19298,
         n19299, n19300, n19301, n19302, n19303, n19304, n19305, n19306,
         n19307, n19308, n19309, n19310, n19311, n19312, n19313, n19314,
         n19315, n19316, n19317, n19318, n19319, n19320, n19321, n19322,
         n19323, n19324, n19325, n19326, n19327, n19328, n19329, n19330,
         n19331, n19332, n19333, n19334, n19335, n19336, n19337, n19338,
         n19339, n19340, n19341, n19342, n19343, n19344, n19345, n19346,
         n19347, n19348, n19349, n19350, n19351, n19352, n19353, n19354,
         n19355, n19356, n19357, n19358, n19359, n19360, n19361, n19362,
         n19363, n19364, n19365, n19366, n19367, n19368, n19369, n19370,
         n19371, n19372, n19373, n19374, n19375, n19376, n19377, n19378,
         n19379, n19380, n19381, n19382, n19383, n19384, n19385, n19386,
         n19387, n19388, n19389, n19390, n19391, n19392, n19393, n19394,
         n19395, n19396, n19397, n19398, n19399, n19400, n19401, n19402,
         n19403, n19404, n19405, n19406, n19407, n19408, n19409, n19410,
         n19411, n19412, n19413, n19414, n19415, n19416, n19417, n19418,
         n19419, n19420, n19421, n19422, n19423, n19424, n19425, n19426,
         n19427, n19428, n19429, n19430, n19431, n19432, n19433, n19434,
         n19435, n19436, n19437, n19438, n19439, n19440, n19441, n19442,
         n19443, n19444, n19445, n19446, n19447, n19448, n19449, n19450,
         n19451, n19452, n19453, n19454, n19455, n19456, n19457, n19458,
         n19459, n19460, n19461, n19462, n19463, n19464, n19465, n19466,
         n19467, n19468, n19469, n19470, n19471, n19472, n19473, n19474,
         n19475, n19476, n19477, n19478, n19479, n19480, n19481, n19482,
         n19483, n19484, n19485, n19486, n19487, n19488, n19489, n19490,
         n19491, n19492, n19493, n19494, n19495, n19496, n19497, n19498,
         n19499, n19500, n19501, n19502, n19503, n19504, n19505, n19506,
         n19507, n19508, n19509, n19510, n19511, n19512, n19513, n19514,
         n19515, n19516, n19517, n19518, n19519, n19520, n19521, n19522,
         n19523, n19524, n19525, n19526, n19527, n19528, n19529, n19530,
         n19531, n19532, n19533, n19534, n19535, n19536, n19537, n19538,
         n19539, n19540, n19541, n19542, n19543, n19544, n19545, n19546,
         n19547, n19548, n19549, n19550, n19551, n19552, n19553, n19554,
         n19555, n19556, n19557, n19558, n19559, n19560, n19561, n19562,
         n19563, n19564, n19565, n19566, n19567, n19568, n19569, n19570,
         n19571, n19572, n19573, n19574, n19575, n19576, n19577, n19578,
         n19579, n19580, n19581, n19582, n19583, n19584, n19585, n19586,
         n19587, n19588, n19589, n19590, n19591, n19592, n19593, n19594,
         n19595, n19596, n19597, n19598, n19599, n19600, n19601, n19602,
         n19603, n19604, n19605, n19606, n19607, n19608, n19609, n19610,
         n19611, n19612, n19613, n19614, n19615, n19616, n19617, n19618,
         n19619, n19620, n19621, n19622, n19623, n19624, n19625, n19626,
         n19627, n19628, n19629, n19630, n19631, n19632, n19633, n19634,
         n19635, n19636, n19637, n19638, n19639, n19640, n19641, n19642,
         n19643, n19644, n19645, n19646, n19647, n19648, n19649, n19650,
         n19651, n19652, n19653, n19654, n19655, n19656, n19657, n19658,
         n19659, n19660, n19661, n19662, n19663, n19664, n19665, n19666,
         n19667, n19668, n19669, n19670, n19671, n19672, n19673, n19674,
         n19675, n19676, n19677, n19678, n19679, n19680, n19681, n19682,
         n19683, n19684, n19685, n19686, n19687, n19688, n19689, n19690,
         n19691, n19692, n19693, n19694, n19695, n19696, n19697, n19698,
         n19699, n19700, n19701, n19702, n19703, n19704, n19705, n19706,
         n19707, n19708, n19709, n19710, n19711, n19712, n19713, n19714,
         n19715, n19716, n19717, n19718, n19719, n19720, n19721, n19722,
         n19723, n19724, n19725, n19726, n19727, n19728, n19729, n19730,
         n19731, n19732, n19733, n19734, n19735, n19736, n19737, n19738,
         n19739, n19740, n19741, n19742, n19743, n19744, n19745, n19746,
         n19747, n19748, n19749, n19750, n19751, n19752, n19753, n19754,
         n19755, n19756, n19757, n19758, n19759, n19760, n19761, n19762,
         n19763, n19764, n19765, n19766, n19767, n19768, n19769, n19770,
         n19771, n19772, n19773, n19774, n19775, n19776, n19777, n19778,
         n19779, n19780, n19781, n19782, n19783, n19784, n19785, n19786,
         n19787, n19788, n19789, n19790, n19791, n19792, n19793, n19794,
         n19795, n19796, n19797, n19798, n19799, n19800, n19801, n19802,
         n19803, n19804, n19805, n19806, n19807, n19808, n19809, n19810,
         n19811, n19812, n19813, n19814, n19815, n19816, n19817, n19818,
         n19819, n19820, n19821, n19822, n19823, n19824, n19825, n19826,
         n19827, n19828, n19829, n19830, n19831, n19832, n19833, n19834,
         n19835, n19836, n19837, n19838, n19839, n19840, n19841, n19842,
         n19843, n19844, n19845, n19846, n19847, n19848, n19849, n19850,
         n19851, n19852, n19853, n19854, n19855, n19856, n19857, n19858,
         n19859, n19860, n19861, n19862, n19863, n19864, n19865, n19866,
         n19867, n19868, n19869, n19870, n19871, n19872, n19873, n19874,
         n19875, n19876, n19877, n19878, n19879, n19880, n19881, n19882,
         n19883, n19884, n19885, n19886, n19887, n19888, n19889, n19890,
         n19891, n19892, n19893, n19894, n19895, n19896, n19897, n19898,
         n19899, n19900, n19901, n19902, n19903, n19904, n19905, n19906,
         n19907, n19908, n19909, n19910, n19911, n19912, n19913, n19914,
         n19915, n19916, n19917, n19918, n19919, n19920, n19921, n19922,
         n19923, n19924, n19925, n19926, n19927, n19928, n19929, n19930,
         n19931, n19932, n19933, n19934, n19935, n19936, n19937, n19938,
         n19939, n19940, n19941, n19942, n19943, n19944, n19945, n19946,
         n19947, n19948, n19949, n19950, n19951, n19952, n19953, n19954,
         n19955, n19956, n19957, n19958, n19959, n19960, n19961, n19962,
         n19963, n19964, n19965, n19966, n19967, n19968, n19969, n19970,
         n19971, n19972, n19973, n19974, n19975, n19976, n19977, n19978,
         n19979, n19980, n19981, n19982, n19983, n19984, n19985, n19986,
         n19987, n19988, n19989, n19990, n19991, n19992, n19993, n19994,
         n19995, n19996, n19997, n19998, n19999, n20000, n20001, n20002,
         n20003, n20004, n20005, n20006, n20007, n20008, n20009, n20010,
         n20011, n20012, n20013, n20014, n20015, n20016, n20017, n20018,
         n20019, n20020, n20021, n20022, n20023, n20024, n20025, n20026,
         n20027, n20028, n20029, n20030, n20031, n20032, n20033, n20034,
         n20035, n20036, n20037, n20038, n20039, n20040, n20041, n20042,
         n20043, n20044, n20045, n20046, n20047, n20048, n20049, n20050,
         n20051, n20052, n20053, n20054, n20055, n20056, n20057, n20058,
         n20059, n20060, n20061, n20062, n20063, n20064, n20065, n20066,
         n20067, n20068, n20069, n20070, n20071, n20072, n20073, n20074,
         n20075, n20076, n20077, n20078, n20079, n20080, n20081, n20082,
         n20083, n20084, n20085, n20086, n20087, n20088, n20089, n20090,
         n20091, n20092, n20093, n20094, n20095, n20096, n20097, n20098,
         n20099, n20100, n20101, n20102, n20103, n20104, n20105, n20106,
         n20107, n20108, n20109, n20110, n20111, n20112, n20113, n20114,
         n20115, n20116, n20117, n20118, n20119, n20120, n20121, n20122,
         n20123, n20124, n20125, n20126, n20127, n20128, n20129, n20130,
         n20131, n20132, n20133, n20134, n20135, n20136, n20137, n20138,
         n20139, n20140, n20141, n20142, n20143, n20144, n20145, n20146,
         n20147, n20148, n20149, n20150, n20151, n20152, n20153, n20154,
         n20155, n20156, n20157, n20158, n20159, n20160, n20161, n20162,
         n20163, n20164, n20165, n20166, n20167, n20168, n20169, n20170,
         n20171, n20172, n20173, n20174, n20175, n20176, n20177, n20178,
         n20179, n20180, n20181, n20182, n20183, n20184, n20185, n20186,
         n20187, n20188, n20189, n20190, n20191, n20192, n20193, n20194,
         n20195, n20196, n20197, n20198, n20199, n20200, n20201, n20202,
         n20203, n20204, n20205, n20206, n20207, n20208, n20209, n20210,
         n20211, n20212, n20213, n20214, n20215, n20216, n20217, n20218,
         n20219, n20220, n20221, n20222, n20223, n20224, n20225, n20226,
         n20227, n20228, n20229, n20230, n20231, n20232, n20233, n20234,
         n20235, n20236, n20237, n20238, n20239, n20240, n20241, n20242,
         n20243, n20244, n20245, n20246, n20247, n20248, n20249, n20250,
         n20251, n20252, n20253, n20254, n20255, n20256, n20257, n20258,
         n20259, n20260, n20261, n20262, n20263, n20264, n20265, n20266,
         n20267, n20268, n20269, n20270, n20271, n20272, n20273, n20274,
         n20275, n20276, n20277, n20278, n20279, n20280, n20281, n20282,
         n20283, n20284, n20285, n20286, n20287, n20288, n20289, n20290,
         n20291, n20292, n20293, n20294, n20295, n20296, n20297, n20298,
         n20299, n20300, n20301, n20302, n20303, n20304, n20305, n20306,
         n20307, n20308, n20309, n20310, n20311, n20312, n20313, n20314,
         n20315, n20316, n20317, n20318, n20319, n20320, n20321, n20322,
         n20323, n20324, n20325, n20326, n20327, n20328, n20329, n20330,
         n20331, n20332, n20333, n20334, n20335, n20336, n20337, n20338,
         n20339, n20340, n20341, n20342, n20343, n20344, n20345, n20346,
         n20347, n20348, n20349, n20350, n20351, n20352, n20353, n20354,
         n20355, n20356, n20357, n20358, n20359, n20360, n20361, n20362,
         n20363, n20364, n20365, n20366, n20367, n20368, n20369, n20370,
         n20371, n20372, n20373, n20374, n20375, n20376, n20377, n20378,
         n20379, n20380, n20381, n20382, n20383, n20384, n20385, n20386,
         n20387, n20388, n20389, n20390, n20391, n20392, n20393, n20394,
         n20395, n20396, n20397, n20398, n20399, n20400, n20401, n20402,
         n20403, n20404, n20405, n20406, n20407, n20408, n20409, n20410,
         n20411, n20412, n20413, n20414, n20415, n20416, n20417, n20418,
         n20419, n20420, n20421, n20422, n20423, n20424, n20425, n20426,
         n20427, n20428, n20429, n20430, n20431, n20432, n20433, n20434,
         n20435, n20436, n20437, n20438, n20439, n20440, n20441, n20442,
         n20443, n20444, n20445, n20446, n20447, n20448, n20449, n20450,
         n20451, n20452, n20453, n20454, n20455, n20456, n20457, n20458,
         n20459, n20460, n20461, n20462, n20463, n20464, n20465, n20466,
         n20467, n20468, n20469, n20470, n20471, n20472, n20473, n20474,
         n20475, n20476, n20477, n20478, n20479, n20480, n20481, n20482,
         n20483, n20484, n20485, n20486, n20487, n20488, n20489, n20490,
         n20491, n20492, n20493, n20494, n20495, n20496, n20497, n20498,
         n20499, n20500, n20501, n20502, n20503, n20504, n20505, n20506,
         n20507, n20508, n20509, n20510, n20511, n20512, n20513, n20514,
         n20515, n20516, n20517, n20518, n20519, n20520, n20521, n20522,
         n20523, n20524, n20525, n20526, n20527, n20528, n20529, n20530,
         n20531, n20532, n20533, n20534, n20535, n20536, n20537, n20538,
         n20539, n20540, n20541, n20542, n20543, n20544, n20545, n20546,
         n20547, n20548, n20549, n20550, n20551, n20552, n20553, n20554,
         n20555, n20556, n20557, n20558, n20559, n20560, n20561, n20562,
         n20563, n20564, n20565, n20566, n20567, n20568, n20569, n20570,
         n20571, n20572, n20573, n20574, n20575, n20576, n20577, n20578,
         n20579, n20580, n20581, n20582, n20583, n20584, n20585, n20586,
         n20587, n20588, n20589, n20590, n20591, n20592, n20593, n20594,
         n20595, n20596, n20597, n20598, n20599, n20600, n20601, n20602,
         n20603, n20604, n20605, n20606, n20607, n20608, n20609, n20610,
         n20611, n20612, n20613, n20614, n20615, n20616, n20617, n20618,
         n20619, n20620, n20621, n20622, n20623, n20624, n20625, n20626,
         n20627, n20628, n20629, n20630, n20631, n20632, n20633, n20634,
         n20635, n20636, n20637, n20638, n20639, n20640, n20641, n20642,
         n20643, n20644, n20645, n20646, n20647, n20648, n20649, n20650,
         n20651, n20652, n20653, n20654, n20655, n20656, n20657, n20658,
         n20659, n20660, n20661, n20662, n20663, n20664, n20665, n20666,
         n20667, n20668, n20669, n20670, n20671, n20672, n20673, n20674,
         n20675, n20676, n20677, n20678, n20679, n20680, n20681, n20682,
         n20683, n20684, n20685, n20686, n20687, n20688, n20689, n20690,
         n20691, n20692, n20693, n20694, n20695, n20696, n20697, n20698,
         n20699, n20700, n20701, n20702, n20703, n20704, n20705, n20706,
         n20707, n20708, n20709, n20710, n20711, n20712, n20713, n20714,
         n20715, n20716, n20717, n20718, n20719, n20720, n20721, n20722,
         n20723, n20724, n20725, n20726, n20727, n20728, n20729, n20730,
         n20731, n20732, n20733, n20734, n20735, n20736, n20737, n20738,
         n20739, n20740, n20741, n20742, n20743, n20744, n20745, n20746,
         n20747, n20748, n20749, n20750, n20751, n20752, n20753, n20754,
         n20755, n20756, n20757, n20758, n20759, n20760, n20761, n20762,
         n20763, n20764, n20765, n20766, n20767, n20768, n20769, n20770,
         n20771, n20772, n20773, n20774, n20775, n20776, n20777, n20778,
         n20779, n20780, n20781, n20782, n20783, n20784, n20785, n20786,
         n20787, n20788, n20789, n20790, n20791, n20792, n20793, n20794,
         n20795, n20796, n20797, n20798, n20799, n20800, n20801, n20802,
         n20803, n20804, n20805, n20806, n20807, n20808, n20809, n20810,
         n20811, n20812, n20813, n20814, n20815, n20816, n20817, n20818,
         n20819, n20820, n20821, n20822, n20823, n20824, n20825, n20826,
         n20827, n20828, n20829, n20830, n20831, n20832, n20833, n20834,
         n20835, n20836, n20837, n20838, n20839, n20840, n20841, n20842,
         n20843, n20844, n20845, n20846, n20847, n20848, n20849, n20850,
         n20851, n20852, n20853, n20854, n20855, n20856, n20857, n20858,
         n20859, n20860, n20861, n20862, n20863, n20864, n20865, n20866,
         n20867, n20868, n20869, n20870, n20871, n20872, n20873, n20874,
         n20875, n20876, n20877, n20878, n20879, n20880, n20881, n20882,
         n20883, n20884, n20885, n20886, n20887, n20888, n20889, n20890,
         n20891, n20892, n20893, n20894, n20895, n20896, n20897, n20898,
         n20899, n20900, n20901, n20902, n20903, n20904, n20905, n20906,
         n20907, n20908, n20909, n20910, n20911, n20912, n20913, n20914,
         n20915, n20916, n20917, n20918, n20919, n20920, n20921, n20922,
         n20923, n20924, n20925, n20926, n20927, n20928, n20929, n20930,
         n20931, n20932, n20933, n20934, n20935, n20936, n20937, n20938,
         n20939, n20940, n20941, n20942, n20943, n20944, n20945, n20946,
         n20947, n20948, n20949, n20950, n20951, n20952, n20953, n20954,
         n20955, n20956, n20957, n20958, n20959, n20960, n20961, n20962,
         n20963, n20964, n20965, n20966, n20967, n20968, n20969, n20970,
         n20971, n20972, n20973, n20974, n20975, n20976, n20977, n20978,
         n20979, n20980, n20981, n20982, n20983, n20984, n20985, n20986,
         n20987, n20988, n20989, n20990, n20991, n20992, n20993, n20994,
         n20995, n20996, n20997, n20998, n20999, n21000, n21001, n21002,
         n21003, n21004, n21005, n21006, n21007, n21008, n21009, n21010,
         n21011, n21012, n21013, n21014, n21015, n21016, n21017, n21018,
         n21019, n21020, n21021, n21022, n21023, n21024, n21025, n21026,
         n21027, n21028, n21029, n21030, n21031, n21032, n21033, n21034,
         n21035, n21036, n21037, n21038, n21039, n21040, n21041, n21042,
         n21043, n21044, n21045, n21046, n21047, n21048, n21049, n21050,
         n21051, n21052, n21053, n21054, n21055, n21056, n21057, n21058,
         n21059, n21060, n21061, n21062, n21063, n21064, n21065, n21066,
         n21067, n21068, n21069, n21070, n21071, n21072, n21073, n21074,
         n21075, n21076, n21077, n21078, n21079, n21080, n21081, n21082,
         n21083, n21084, n21085, n21086, n21087, n21088, n21089, n21090,
         n21091, n21092, n21093, n21094, n21095, n21096, n21097, n21098,
         n21099, n21100, n21101, n21102, n21103, n21104, n21105, n21106,
         n21107, n21108, n21109, n21110, n21111, n21112, n21113, n21114,
         n21115, n21116, n21117, n21118, n21119, n21120, n21121, n21122,
         n21123, n21124, n21125, n21126, n21127, n21128, n21129, n21130,
         n21131, n21132, n21133, n21134, n21135, n21136, n21137, n21138,
         n21139, n21140, n21141, n21142, n21143, n21144, n21145, n21146,
         n21147, n21148, n21149, n21150, n21151, n21152, n21153, n21154,
         n21155, n21156, n21157, n21158, n21159, n21160, n21161, n21162,
         n21163, n21164, n21165, n21166, n21167, n21168, n21169, n21170,
         n21171, n21172, n21173, n21174, n21175, n21176, n21177, n21178,
         n21179, n21180, n21181, n21182, n21183, n21184, n21185, n21186,
         n21187, n21188, n21189, n21190, n21191, n21192, n21193, n21194,
         n21195, n21196, n21197, n21198, n21199, n21200, n21201, n21202,
         n21203, n21204, n21205, n21206, n21207, n21208, n21209, n21210,
         n21211, n21212, n21213, n21214, n21215, n21216, n21217, n21218,
         n21219, n21220, n21221, n21222, n21223, n21224, n21225, n21226,
         n21227, n21228, n21229, n21230, n21231, n21232, n21233, n21234,
         n21235, n21236, n21237, n21238, n21239, n21240, n21241, n21242,
         n21243, n21244, n21245, n21246, n21247, n21248, n21249, n21250,
         n21251, n21252, n21253, n21254, n21255, n21256, n21257, n21258,
         n21259, n21260, n21261, n21262, n21263, n21264, n21265, n21266,
         n21267, n21268, n21269, n21270, n21271, n21272, n21273, n21274,
         n21275, n21276, n21277, n21278, n21279, n21280, n21281, n21282,
         n21283, n21284, n21285, n21286, n21287, n21288, n21289, n21290,
         n21291, n21292, n21293, n21294, n21295, n21296, n21297, n21298,
         n21299, n21300, n21301, n21302, n21303, n21304, n21305, n21306,
         n21307, n21308, n21309, n21310, n21311, n21312, n21313, n21314,
         n21315, n21316, n21317, n21318, n21319, n21320, n21321, n21322,
         n21323, n21324, n21325, n21326, n21327, n21328, n21329, n21330,
         n21331, n21332, n21333, n21334, n21335, n21336, n21337, n21338,
         n21339, n21340, n21341, n21342, n21343, n21344, n21345, n21346,
         n21347, n21348, n21349, n21350, n21351, n21352, n21353, n21354,
         n21355, n21356, n21357, n21358, n21359, n21360, n21361, n21362,
         n21363, n21364, n21365, n21366, n21367, n21368, n21369, n21370,
         n21371, n21372, n21373, n21374, n21375, n21376, n21377, n21378,
         n21379, n21380, n21381, n21382, n21383, n21384, n21385, n21386,
         n21387, n21388, n21389, n21390, n21391, n21392, n21393, n21394,
         n21395, n21396, n21397, n21398, n21399, n21400, n21401, n21402,
         n21403, n21404, n21405, n21406, n21407, n21408, n21409, n21410,
         n21411, n21412, n21413, n21414, n21415, n21416, n21417, n21418,
         n21419, n21420, n21421, n21422, n21423, n21424, n21425, n21426,
         n21427, n21428, n21429, n21430, n21431, n21432, n21433, n21434,
         n21435, n21436, n21437, n21438, n21439, n21440, n21441, n21442,
         n21443, n21444, n21445, n21446, n21447, n21448, n21449, n21450,
         n21451, n21452, n21453, n21454, n21455, n21456, n21457, n21458,
         n21459, n21460, n21461, n21462, n21463, n21464, n21465, n21466,
         n21467, n21468, n21469, n21470, n21471, n21472, n21473, n21474,
         n21475, n21476, n21477, n21478, n21479, n21480, n21481, n21482,
         n21483, n21484, n21485, n21486, n21487, n21488, n21489, n21490,
         n21491, n21492, n21493, n21494, n21495, n21496, n21497, n21498,
         n21499, n21500, n21501, n21502, n21503, n21504, n21505, n21506,
         n21507, n21508, n21509, n21510, n21511, n21512, n21513, n21514,
         n21515, n21516, n21517, n21518, n21519, n21520, n21521, n21522,
         n21523, n21524, n21525, n21526, n21527, n21528, n21529, n21530,
         n21531, n21532, n21533, n21534, n21535, n21536, n21537, n21538,
         n21539, n21540, n21541, n21542, n21543, n21544, n21545, n21546,
         n21547, n21548, n21549, n21550, n21551, n21552, n21553, n21554,
         n21555, n21556, n21557, n21558, n21559, n21560, n21561, n21562,
         n21563, n21564, n21565, n21566, n21567, n21568, n21569, n21570,
         n21571, n21572, n21573, n21574, n21575, n21576, n21577, n21578,
         n21579, n21580, n21581, n21582, n21583, n21584, n21585, n21586,
         n21587, n21588, n21589, n21590, n21591, n21592, n21593, n21594,
         n21595, n21596, n21597, n21598, n21599, n21600, n21601, n21602,
         n21603, n21604, n21605, n21606, n21607, n21608, n21609, n21610,
         n21611, n21612, n21613, n21614, n21615, n21616, n21617, n21618,
         n21619, n21620, n21621, n21622, n21623, n21624, n21625, n21626,
         n21627, n21628, n21629, n21630, n21631, n21632, n21633, n21634,
         n21635, n21636, n21637, n21638, n21639, n21640, n21641, n21642,
         n21643, n21644, n21645, n21646, n21647, n21648, n21649, n21650,
         n21651, n21652, n21653, n21654, n21655, n21656, n21657, n21658,
         n21659, n21660, n21661, n21662, n21663, n21664, n21665, n21666,
         n21667, n21668, n21669, n21670, n21671, n21672, n21673, n21674,
         n21675, n21676, n21677, n21678, n21679, n21680, n21681, n21682,
         n21683, n21684, n21685, n21686, n21687, n21688, n21689, n21690,
         n21691, n21692, n21693, n21694, n21695, n21696, n21697, n21698,
         n21699, n21700, n21701, n21702, n21703, n21704, n21705, n21706,
         n21707, n21708, n21709, n21710, n21711, n21712, n21713, n21714,
         n21715, n21716, n21717, n21718, n21719, n21720, n21721, n21722,
         n21723, n21724, n21725, n21726, n21727, n21728, n21729, n21730,
         n21731, n21732, n21733, n21734, n21735, n21736, n21737, n21738,
         n21739, n21740, n21741, n21742, n21743, n21744, n21745, n21746,
         n21747, n21748, n21749, n21750, n21751, n21752, n21753, n21754,
         n21755, n21756, n21757, n21758, n21759, n21760, n21761, n21762,
         n21763, n21764, n21765, n21766, n21767, n21768, n21769, n21770,
         n21771, n21772, n21773, n21774, n21775, n21776, n21777, n21778,
         n21779, n21780, n21781, n21782, n21783, n21784, n21785, n21786,
         n21787, n21788, n21789, n21790, n21791, n21792, n21793, n21794,
         n21795, n21796, n21797, n21798, n21799, n21800, n21801, n21802,
         n21803, n21804, n21805, n21806, n21807, n21808, n21809, n21810,
         n21811, n21812, n21813, n21814, n21815, n21816, n21817, n21818,
         n21819, n21820, n21821, n21822, n21823, n21824, n21825, n21826,
         n21827, n21828, n21829, n21830, n21831, n21832, n21833, n21834,
         n21835, n21836, n21837, n21838, n21839, n21840, n21841, n21842,
         n21843, n21844, n21845, n21846, n21847, n21848, n21849, n21850,
         n21851, n21852, n21853, n21854, n21855, n21856, n21857, n21858,
         n21859, n21860, n21861, n21862, n21863, n21864, n21865, n21866,
         n21867, n21868, n21869, n21870, n21871, n21872, n21873, n21874,
         n21875, n21876, n21877, n21878, n21879, n21880, n21881, n21882,
         n21883, n21884, n21885, n21886, n21887, n21888, n21889, n21890,
         n21891, n21892, n21893, n21894, n21895, n21896, n21897, n21898,
         n21899, n21900, n21901, n21902, n21903, n21904, n21905, n21906,
         n21907, n21908, n21909, n21910, n21911, n21912, n21913, n21914,
         n21915, n21916, n21917, n21918, n21919, n21920, n21921, n21922,
         n21923, n21924, n21925, n21926, n21927, n21928, n21929, n21930,
         n21931, n21932, n21933, n21934, n21935, n21936, n21937, n21938,
         n21939, n21940, n21941, n21942, n21943, n21944, n21945, n21946,
         n21947, n21948, n21949, n21950, n21951, n21952, n21953, n21954,
         n21955, n21956, n21957, n21958, n21959, n21960, n21961, n21962,
         n21963, n21964, n21965, n21966, n21967, n21968, n21969, n21970,
         n21971, n21972, n21973, n21974, n21975, n21976, n21977, n21978,
         n21979, n21980, n21981, n21982, n21983, n21984, n21985, n21986,
         n21987, n21988, n21989, n21990, n21991, n21992, n21993, n21994,
         n21995, n21996, n21997, n21998, n21999, n22000, n22001, n22002,
         n22003, n22004, n22005, n22006, n22007, n22008, n22009, n22010,
         n22011, n22012, n22013, n22014, n22015, n22016, n22017, n22018,
         n22019, n22020, n22021, n22022, n22023, n22024, n22025, n22026,
         n22027, n22028, n22029, n22030, n22031, n22032, n22033, n22034,
         n22035, n22036, n22037, n22038, n22039, n22040, n22041, n22042,
         n22043, n22044, n22045, n22046, n22047, n22048, n22049, n22050,
         n22051, n22052, n22053, n22054, n22055, n22056, n22057, n22058,
         n22059, n22060, n22061, n22062, n22063, n22064, n22065, n22066,
         n22067, n22068, n22069, n22070, n22071, n22072, n22073, n22074,
         n22075, n22076, n22077, n22078, n22079, n22080, n22081, n22082,
         n22083, n22084, n22085, n22086, n22087, n22088, n22089, n22090,
         n22091, n22092, n22093, n22094, n22095, n22096, n22097, n22098,
         n22099, n22100, n22101, n22102, n22103, n22104, n22105, n22106,
         n22107, n22108, n22109, n22110, n22111, n22112, n22113, n22114,
         n22115, n22116, n22117, n22118, n22119, n22120, n22121, n22122,
         n22123, n22124, n22125, n22126, n22127, n22128, n22129, n22130,
         n22131, n22132, n22133, n22134, n22135, n22136, n22137, n22138,
         n22139, n22140, n22141, n22142, n22143, n22144, n22145, n22146,
         n22147, n22148, n22149, n22150, n22151, n22152, n22153, n22154,
         n22155, n22156, n22157, n22158, n22159, n22160, n22161, n22162,
         n22163, n22164, n22165, n22166, n22167, n22168, n22169, n22170,
         n22171, n22172, n22173, n22174, n22175, n22176, n22177, n22178,
         n22179, n22180, n22181, n22182, n22183, n22184, n22185, n22186,
         n22187, n22188, n22189, n22190, n22191, n22192, n22193, n22194,
         n22195, n22196, n22197, n22198, n22199, n22200, n22201, n22202,
         n22203, n22204, n22205, n22206, n22207, n22208, n22209, n22210,
         n22211, n22212, n22213, n22214, n22215, n22216, n22217, n22218,
         n22219, n22220, n22221, n22222, n22223, n22224, n22225, n22226,
         n22227, n22228, n22229, n22230, n22231, n22232, n22233, n22234,
         n22235, n22236, n22237, n22238, n22239, n22240, n22241, n22242,
         n22243, n22244, n22245, n22246, n22247, n22248, n22249, n22250,
         n22251, n22252, n22253, n22254, n22255, n22256, n22257, n22258,
         n22259, n22260, n22261, n22262, n22263, n22264, n22265, n22266,
         n22267, n22268, n22269, n22270, n22271, n22272, n22273, n22274,
         n22275, n22276, n22277, n22278, n22279, n22280, n22281, n22282,
         n22283, n22284, n22285, n22286, n22287, n22288, n22289, n22290,
         n22291, n22292, n22293, n22294, n22295, n22296, n22297, n22298,
         n22299, n22300, n22301, n22302, n22303, n22304, n22305, n22306,
         n22307, n22308, n22309, n22310, n22311, n22312, n22313, n22314,
         n22315, n22316, n22317, n22318, n22319, n22320, n22321, n22322,
         n22323, n22324, n22325, n22326, n22327, n22328, n22329, n22330,
         n22331, n22332, n22333, n22334, n22335, n22336, n22337, n22338,
         n22339, n22340, n22341, n22342, n22343, n22344, n22345, n22346,
         n22347, n22348, n22349, n22350, n22351, n22352, n22353, n22354,
         n22355, n22356, n22357, n22358, n22359, n22360, n22361, n22362,
         n22363, n22364, n22365, n22366, n22367, n22368, n22369, n22370,
         n22371, n22372, n22373, n22374, n22375, n22376, n22377, n22378,
         n22379, n22380, n22381, n22382, n22383, n22384, n22385, n22386,
         n22387, n22388, n22389, n22390, n22391, n22392, n22393, n22394,
         n22395, n22396, n22397, n22398, n22399, n22400, n22401, n22402,
         n22403, n22404, n22405, n22406, n22407, n22408, n22409, n22410,
         n22411, n22412, n22413, n22414, n22415, n22416, n22417, n22418,
         n22419, n22420, n22421, n22422, n22423, n22424, n22425, n22426,
         n22427, n22428, n22429, n22430, n22431, n22432, n22433, n22434,
         n22435, n22436, n22437, n22438, n22439, n22440, n22441, n22442,
         n22443, n22444, n22445, n22446, n22447, n22448, n22449, n22450,
         n22451, n22452, n22453, n22454, n22455, n22456, n22457, n22458,
         n22459, n22460, n22461, n22462, n22463, n22464, n22465, n22466,
         n22467, n22468, n22469, n22470, n22471, n22472, n22473, n22474,
         n22475, n22476, n22477, n22478, n22479, n22480, n22481, n22482,
         n22483, n22484, n22485, n22486, n22487, n22488, n22489, n22490,
         n22491, n22492, n22493, n22494, n22495, n22496, n22497, n22498,
         n22499, n22500, n22501, n22502, n22503, n22504, n22505, n22506,
         n22507, n22508, n22509, n22510, n22511, n22512, n22513, n22514,
         n22515, n22516, n22517, n22518, n22519, n22520, n22521, n22522,
         n22523, n22524, n22525, n22526, n22527, n22528, n22529, n22530,
         n22531, n22532, n22533, n22534, n22535, n22536, n22537, n22538,
         n22539, n22540, n22541, n22542, n22543, n22544, n22545, n22546,
         n22547, n22548, n22549, n22550, n22551, n22552, n22553, n22554,
         n22555, n22556, n22557, n22558, n22559, n22560, n22561, n22562,
         n22563, n22564, n22565, n22566, n22567, n22568, n22569, n22570,
         n22571, n22572, n22573, n22574, n22575, n22576, n22577, n22578,
         n22579, n22580, n22581, n22582, n22583, n22584, n22585, n22586,
         n22587, n22588, n22589, n22590, n22591, n22592, n22593, n22594,
         n22595, n22596, n22597, n22598, n22599, n22600, n22601, n22602,
         n22603, n22604, n22605, n22606, n22607, n22608, n22609, n22610,
         n22611, n22612, n22613, n22614, n22615, n22616, n22617, n22618,
         n22619, n22620, n22621, n22622, n22623, n22624, n22625, n22626,
         n22627, n22628, n22629, n22630, n22631, n22632, n22633, n22634,
         n22635, n22636, n22637, n22638, n22639, n22640, n22641, n22642,
         n22643, n22644, n22645, n22646, n22647, n22648, n22649, n22650,
         n22651, n22652, n22653, n22654, n22655, n22656, n22657, n22658,
         n22659, n22660, n22661, n22662, n22663, n22664, n22665, n22666,
         n22667, n22668, n22669, n22670, n22671, n22672, n22673, n22674,
         n22675, n22676, n22677, n22678, n22679, n22680, n22681, n22682,
         n22683, n22684, n22685, n22686, n22687, n22688, n22689, n22690,
         n22691, n22692, n22693, n22694, n22695, n22696, n22697, n22698,
         n22699, n22700, n22701, n22702, n22703, n22704, n22705, n22706,
         n22707, n22708, n22709, n22710, n22711, n22712, n22713, n22714,
         n22715, n22716, n22717, n22718, n22719, n22720, n22721, n22722,
         n22723, n22724, n22725, n22726, n22727, n22728, n22729, n22730,
         n22731, n22732, n22733, n22734, n22735, n22736, n22737, n22738,
         n22739, n22740, n22741, n22742, n22743, n22744, n22745, n22746,
         n22747, n22748, n22749, n22750, n22751, n22752, n22753, n22754,
         n22755, n22756, n22757, n22758, n22759, n22760, n22761, n22762,
         n22763, n22764, n22765, n22766, n22767, n22768, n22769, n22770,
         n22771, n22772, n22773, n22774, n22775, n22776, n22777, n22778,
         n22779, n22780, n22781, n22782, n22783, n22784, n22785, n22786,
         n22787, n22788, n22789, n22790, n22791, n22792, n22793, n22794,
         n22795, n22796, n22797, n22798, n22799, n22800, n22801, n22802,
         n22803, n22804, n22805, n22806, n22807, n22808, n22809, n22810,
         n22811, n22812, n22813, n22814, n22815, n22816, n22817, n22818,
         n22819, n22820, n22821, n22822, n22823, n22824, n22825, n22826,
         n22827, n22828, n22829, n22830, n22831, n22832, n22833, n22834,
         n22835, n22836, n22837, n22838, n22839, n22840, n22841, n22842,
         n22843, n22844, n22845, n22846, n22847, n22848, n22849, n22850,
         n22851, n22852, n22853, n22854, n22855, n22856, n22857, n22858,
         n22859, n22860, n22861, n22862, n22863, n22864, n22865, n22866,
         n22867, n22868, n22869, n22870, n22871, n22872, n22873, n22874,
         n22875, n22876, n22877, n22878, n22879, n22880, n22881, n22882,
         n22883, n22884, n22885, n22886, n22887, n22888, n22889, n22890,
         n22891, n22892, n22893, n22894, n22895, n22896, n22897, n22898,
         n22899, n22900, n22901, n22902, n22903, n22904, n22905, n22906,
         n22907, n22908, n22909, n22910, n22911, n22912, n22913, n22914,
         n22915, n22916, n22917, n22918, n22919, n22920, n22921, n22922,
         n22923, n22924, n22925, n22926, n22927, n22928, n22929, n22930,
         n22931, n22932, n22933, n22934, n22935, n22936, n22937, n22938,
         n22939, n22940, n22941, n22942, n22943, n22944, n22945, n22946,
         n22947, n22948, n22949, n22950, n22951, n22952, n22953, n22954,
         n22955, n22956, n22957, n22958, n22959, n22960, n22961, n22962,
         n22963, n22964, n22965, n22966, n22967, n22968, n22969, n22970,
         n22971, n22972, n22973, n22974, n22975, n22976, n22977, n22978,
         n22979, n22980, n22981, n22982, n22983, n22984, n22985, n22986,
         n22987, n22988, n22989, n22990, n22991, n22992, n22993, n22994,
         n22995, n22996, n22997, n22998, n22999, n23000, n23001, n23002,
         n23003, n23004, n23005, n23006, n23007, n23008, n23009, n23010,
         n23011, n23012, n23013, n23014, n23015, n23016, n23017, n23018,
         n23019, n23020, n23021, n23022, n23023, n23024, n23025, n23026,
         n23027, n23028, n23029, n23030, n23031, n23032, n23033, n23034,
         n23035, n23036, n23037, n23038, n23039, n23040, n23041, n23042,
         n23043, n23044, n23045, n23046, n23047, n23048, n23049, n23050,
         n23051, n23052, n23053, n23054, n23055, n23056, n23057, n23058,
         n23059, n23060, n23061, n23062, n23063, n23064, n23065, n23066,
         n23067, n23068, n23069, n23070, n23071, n23072, n23073, n23074,
         n23075, n23076, n23077, n23078, n23079, n23080, n23081, n23082,
         n23083, n23084, n23085, n23086, n23087, n23088, n23089, n23090,
         n23091, n23092, n23093, n23094, n23095, n23096, n23097, n23098,
         n23099, n23100, n23101, n23102, n23103, n23104, n23105, n23106,
         n23107, n23108, n23109, n23110, n23111, n23112, n23113, n23114,
         n23115, n23116, n23117, n23118, n23119, n23120, n23121, n23122,
         n23123, n23124, n23125, n23126, n23127, n23128, n23129, n23130,
         n23131, n23132, n23133, n23134, n23135, n23136, n23137, n23138,
         n23139, n23140, n23141, n23142, n23143, n23144, n23145, n23146,
         n23147, n23148, n23149, n23150, n23151, n23152, n23153, n23154,
         n23155, n23156, n23157, n23158, n23159, n23160, n23161, n23162,
         n23163, n23164, n23165, n23166, n23167, n23168, n23169, n23170,
         n23171, n23172, n23173, n23174, n23175, n23176, n23177, n23178,
         n23179, n23180, n23181, n23182, n23183, n23184, n23185, n23186,
         n23187, n23188, n23189, n23190, n23191, n23192, n23193, n23194,
         n23195, n23196, n23197, n23198, n23199, n23200, n23201, n23202,
         n23203, n23204, n23205, n23206, n23207, n23208, n23209, n23210,
         n23211, n23212, n23213, n23214, n23215, n23216, n23217, n23218,
         n23219, n23220, n23221, n23222, n23223, n23224, n23225, n23226,
         n23227, n23228, n23229, n23230, n23231, n23232, n23233, n23234,
         n23235, n23236, n23237, n23238, n23239, n23240, n23241, n23242,
         n23243, n23244, n23245, n23246, n23247, n23248, n23249, n23250,
         n23251, n23252, n23253, n23254, n23255, n23256, n23257, n23258,
         n23259, n23260, n23261, n23262, n23263, n23264, n23265, n23266,
         n23267, n23268, n23269, n23270, n23271, n23272, n23273, n23274,
         n23275, n23276, n23277, n23278, n23279, n23280, n23281, n23282,
         n23283, n23284, n23285, n23286, n23287, n23288, n23289, n23290,
         n23291, n23292, n23293, n23294, n23295, n23296, n23297, n23298,
         n23299, n23300, n23301, n23302, n23303, n23304, n23305, n23306,
         n23307, n23308, n23309, n23310, n23311, n23312, n23313, n23314,
         n23315, n23316, n23317, n23318, n23319, n23320, n23321, n23322,
         n23323, n23324, n23325, n23326, n23327, n23328, n23329, n23330,
         n23331, n23332, n23333, n23334, n23335, n23336, n23337, n23338,
         n23339, n23340, n23341, n23342, n23343, n23344, n23345, n23346,
         n23347, n23348, n23349, n23350, n23351, n23352, n23353, n23354,
         n23355, n23356, n23357, n23358, n23359, n23360, n23361, n23362,
         n23363, n23364, n23365, n23366, n23367, n23368, n23369, n23370,
         n23371, n23372, n23373, n23374, n23375, n23376, n23377, n23378,
         n23379, n23380, n23381, n23382, n23383, n23384, n23385, n23386,
         n23387, n23388, n23389, n23390, n23391, n23392, n23393, n23394,
         n23395, n23396, n23397, n23398, n23399, n23400, n23401, n23402,
         n23403, n23404, n23405, n23406, n23407, n23408, n23409, n23410,
         n23411, n23412, n23413, n23414, n23415, n23416, n23417, n23418,
         n23419, n23420, n23421, n23422, n23423, n23424, n23425, n23426,
         n23427, n23428, n23429, n23430, n23431, n23432, n23433, n23434,
         n23435, n23436, n23437, n23438, n23439, n23440, n23441, n23442,
         n23443, n23444, n23445, n23446, n23447, n23448, n23449, n23450,
         n23451, n23452, n23453, n23454, n23455, n23456, n23457, n23458,
         n23459, n23460, n23461, n23462, n23463, n23464, n23465, n23466,
         n23467, n23468, n23469, n23470, n23471, n23472, n23473, n23474,
         n23475, n23476, n23477, n23478, n23479, n23480, n23481, n23482,
         n23483, n23484, n23485, n23486, n23487, n23488, n23489, n23490,
         n23491, n23492, n23493, n23494, n23495, n23496, n23497, n23498,
         n23499, n23500, n23501, n23502, n23503, n23504, n23505, n23506,
         n23507, n23508, n23509, n23510, n23511, n23512, n23513, n23514,
         n23515, n23516, n23517, n23518, n23519, n23520, n23521, n23522,
         n23523, n23524, n23525, n23526, n23527, n23528, n23529, n23530,
         n23531, n23532, n23533, n23534, n23535, n23536, n23537, n23538,
         n23539, n23540, n23541, n23542, n23543, n23544, n23545, n23546,
         n23547, n23548, n23549, n23550, n23551, n23552, n23553, n23554,
         n23555, n23556, n23557, n23558, n23559, n23560, n23561, n23562,
         n23563, n23564, n23565, n23566, n23567, n23568, n23569, n23570,
         n23571, n23572, n23573, n23574, n23575, n23576, n23577, n23578,
         n23579, n23580, n23581, n23582, n23583, n23584, n23585, n23586,
         n23587, n23588, n23589, n23590, n23591, n23592, n23593, n23594,
         n23595, n23596, n23597, n23598, n23599, n23600, n23601, n23602,
         n23603, n23604, n23605, n23606, n23607, n23608, n23609, n23610,
         n23611, n23612, n23613, n23614, n23615, n23616, n23617, n23618,
         n23619, n23620, n23621, n23622, n23623, n23624, n23625, n23626,
         n23627, n23628, n23629, n23630, n23631, n23632, n23633, n23634,
         n23635, n23636, n23637, n23638, n23639, n23640, n23641, n23642,
         n23643, n23644, n23645, n23646, n23647, n23648, n23649, n23650,
         n23651, n23652, n23653, n23654, n23655, n23656, n23657, n23658,
         n23659, n23660, n23661, n23662, n23663, n23664, n23665, n23666,
         n23667, n23668, n23669, n23670, n23671, n23672, n23673, n23674,
         n23675, n23676, n23677, n23678, n23679, n23680, n23681, n23682,
         n23683, n23684, n23685, n23686, n23687, n23688, n23689, n23690,
         n23691, n23692, n23693, n23694, n23695, n23696, n23697, n23698,
         n23699, n23700, n23701, n23702, n23703, n23704, n23705, n23706,
         n23707, n23708, n23709, n23710, n23711, n23712, n23713, n23714,
         n23715, n23716, n23717, n23718, n23719, n23720, n23721, n23722,
         n23723, n23724, n23725, n23726, n23727, n23728, n23729, n23730,
         n23731, n23732, n23733, n23734, n23735, n23736, n23737, n23738,
         n23739, n23740, n23741, n23742, n23743, n23744, n23745, n23746,
         n23747, n23748, n23749, n23750, n23751, n23752, n23753, n23754,
         n23755, n23756, n23757, n23758, n23759, n23760, n23761, n23762,
         n23763, n23764, n23765, n23766, n23767, n23768, n23769, n23770,
         n23771, n23772, n23773, n23774, n23775, n23776, n23777, n23778,
         n23779, n23780, n23781, n23782, n23783, n23784, n23785, n23786,
         n23787, n23788, n23789, n23790, n23791, n23792, n23793, n23794,
         n23795, n23796, n23797, n23798, n23799, n23800, n23801, n23802,
         n23803, n23804, n23805, n23806, n23807, n23808, n23809, n23810,
         n23811, n23812, n23813, n23814, n23815, n23816, n23817, n23818,
         n23819, n23820, n23821, n23822, n23823, n23824, n23825, n23826,
         n23827, n23828, n23829, n23830, n23831, n23832, n23833, n23834,
         n23835, n23836, n23837, n23838, n23839, n23840, n23841, n23842,
         n23843, n23844, n23845, n23846, n23847, n23848, n23849, n23850,
         n23851, n23852, n23853, n23854, n23855, n23856, n23857, n23858,
         n23859, n23860, n23861, n23862, n23863, n23864, n23865, n23866,
         n23867, n23868, n23869, n23870, n23871, n23872, n23873, n23874,
         n23875, n23876, n23877, n23878, n23879, n23880, n23881, n23882,
         n23883, n23884, n23885, n23886, n23887, n23888, n23889, n23890,
         n23891, n23892, n23893, n23894, n23895, n23896, n23897, n23898,
         n23899, n23900, n23901, n23902, n23903, n23904, n23905, n23906,
         n23907, n23908, n23909, n23910, n23911, n23912, n23913, n23914,
         n23915, n23916, n23917, n23918, n23919, n23920, n23921, n23922,
         n23923, n23924, n23925, n23926, n23927, n23928, n23929, n23930,
         n23931, n23932, n23933, n23934, n23935, n23936, n23937, n23938,
         n23939, n23940, n23941, n23942, n23943, n23944, n23945, n23946,
         n23947, n23948, n23949, n23950, n23951, n23952, n23953, n23954,
         n23955, n23956, n23957, n23958, n23959, n23960, n23961, n23962,
         n23963, n23964, n23965, n23966, n23967, n23968, n23969, n23970,
         n23971, n23972, n23973, n23974, n23975, n23976, n23977, n23978,
         n23979, n23980, n23981, n23982, n23983, n23984, n23985, n23986,
         n23987, n23988, n23989, n23990, n23991, n23992, n23993, n23994,
         n23995, n23996, n23997, n23998, n23999, n24000, n24001, n24002,
         n24003, n24004, n24005, n24006, n24007, n24008, n24009, n24010,
         n24011, n24012, n24013, n24014, n24015, n24016, n24017, n24018,
         n24019, n24020, n24021, n24022, n24023, n24024, n24025, n24026,
         n24027, n24028, n24029, n24030, n24031, n24032, n24033, n24034,
         n24035, n24036, n24037, n24038, n24039, n24040, n24041, n24042,
         n24043, n24044, n24045, n24046, n24047, n24048, n24049, n24050,
         n24051, n24052, n24053, n24054, n24055, n24056, n24057, n24058,
         n24059, n24060, n24061, n24062, n24063, n24064, n24065, n24066,
         n24067, n24068, n24069, n24070, n24071, n24072, n24073, n24074,
         n24075, n24076, n24077, n24078, n24079, n24080, n24081, n24082,
         n24083, n24084, n24085, n24086, n24087, n24088, n24089, n24090,
         n24091, n24092, n24093, n24094, n24095, n24096, n24097, n24098,
         n24099, n24100, n24101, n24102, n24103, n24104, n24105, n24106,
         n24107, n24108, n24109, n24110, n24111, n24112, n24113, n24114,
         n24115, n24116, n24117, n24118, n24119, n24120, n24121, n24122,
         n24123, n24124, n24125, n24126, n24127, n24128, n24129, n24130,
         n24131, n24132, n24133, n24134, n24135, n24136, n24137, n24138,
         n24139, n24140, n24141, n24142, n24143, n24144, n24145, n24146,
         n24147, n24148, n24149, n24150, n24151, n24152, n24153, n24154,
         n24155, n24156, n24157, n24158, n24159, n24160, n24161, n24162,
         n24163, n24164, n24165, n24166, n24167, n24168, n24169, n24170,
         n24171, n24172, n24173, n24174, n24175, n24176, n24177, n24178,
         n24179, n24180, n24181, n24182, n24183, n24184, n24185, n24186,
         n24187, n24188, n24189, n24190, n24191, n24192, n24193, n24194,
         n24195, n24196, n24197, n24198, n24199, n24200, n24201, n24202,
         n24203, n24204, n24205, n24206, n24207, n24208, n24209, n24210,
         n24211, n24212, n24213, n24214, n24215, n24216, n24217, n24218,
         n24219, n24220, n24221, n24222, n24223, n24224, n24225, n24226,
         n24227, n24228, n24229, n24230, n24231, n24232, n24233, n24234,
         n24235, n24236, n24237, n24238, n24239, n24240, n24241, n24242,
         n24243, n24244, n24245, n24246, n24247, n24248, n24249, n24250,
         n24251, n24252, n24253, n24254, n24255, n24256, n24257, n24258,
         n24259, n24260, n24261, n24262, n24263, n24264, n24265, n24266,
         n24267, n24268, n24269, n24270, n24271, n24272, n24273, n24274,
         n24275, n24276, n24277, n24278, n24279, n24280, n24281, n24282,
         n24283, n24284, n24285, n24286, n24287, n24288, n24289, n24290,
         n24291, n24292, n24293, n24294, n24295, n24296, n24297, n24298,
         n24299, n24300, n24301, n24302, n24303, n24304, n24305, n24306,
         n24307, n24308, n24309, n24310, n24311, n24312, n24313, n24314,
         n24315, n24316, n24317, n24318, n24319, n24320, n24321, n24322,
         n24323, n24324, n24325, n24326, n24327, n24328, n24329, n24330,
         n24331, n24332, n24333, n24334, n24335, n24336, n24337, n24338,
         n24339, n24340, n24341, n24342, n24343, n24344, n24345, n24346,
         n24347, n24348, n24349, n24350, n24351, n24352, n24353, n24354,
         n24355, n24356, n24357, n24358, n24359, n24360, n24361, n24362,
         n24363, n24364, n24365, n24366, n24367, n24368, n24369, n24370,
         n24371, n24372, n24373, n24374, n24375, n24376, n24377, n24378,
         n24379, n24380, n24381, n24382, n24383, n24384, n24385, n24386,
         n24387, n24388, n24389, n24390, n24391, n24392, n24393, n24394,
         n24395, n24396, n24397, n24398, n24399, n24400, n24401, n24402,
         n24403, n24404, n24405, n24406, n24407, n24408, n24409, n24410,
         n24411, n24412, n24413, n24414, n24415, n24416, n24417, n24418,
         n24419, n24420, n24421, n24422, n24423, n24424, n24425, n24426,
         n24427, n24428, n24429, n24430, n24431, n24432, n24433, n24434,
         n24435, n24436, n24437, n24438, n24439, n24440, n24441, n24442,
         n24443, n24444, n24445, n24446, n24447, n24448, n24449, n24450,
         n24451, n24452, n24453, n24454, n24455, n24456, n24457, n24458,
         n24459, n24460, n24461, n24462, n24463, n24464, n24465, n24466,
         n24467, n24468, n24469, n24470, n24471, n24472, n24473, n24474,
         n24475, n24476, n24477, n24478, n24479, n24480, n24481, n24482,
         n24483, n24484, n24485, n24486, n24487, n24488, n24489, n24490,
         n24491, n24492, n24493, n24494, n24495, n24496, n24497, n24498,
         n24499, n24500, n24501, n24502, n24503, n24504, n24505, n24506,
         n24507, n24508, n24509, n24510, n24511, n24512, n24513, n24514,
         n24515, n24516, n24517, n24518, n24519, n24520, n24521, n24522,
         n24523, n24524, n24525, n24526, n24527, n24528, n24529, n24530,
         n24531, n24532, n24533, n24534, n24535, n24536, n24537, n24538,
         n24539, n24540, n24541, n24542, n24543, n24544, n24545, n24546,
         n24547, n24548, n24549, n24550, n24551, n24552, n24553, n24554,
         n24555, n24556, n24557, n24558, n24559, n24560, n24561, n24562,
         n24563, n24564, n24565, n24566, n24567, n24568, n24569, n24570,
         n24571, n24572, n24573, n24574, n24575, n24576, n24577, n24578,
         n24579, n24580, n24581, n24582, n24583, n24584, n24585, n24586,
         n24587, n24588, n24589, n24590, n24591, n24592, n24593, n24594,
         n24595, n24596, n24597, n24598, n24599, n24600, n24601, n24602,
         n24603, n24604, n24605, n24606, n24607, n24608, n24609, n24610,
         n24611, n24612, n24613, n24614, n24615, n24616, n24617, n24618,
         n24619, n24620, n24621, n24622, n24623, n24624, n24625, n24626,
         n24627, n24628, n24629, n24630, n24631, n24632, n24633, n24634,
         n24635, n24636, n24637, n24638, n24639, n24640, n24641, n24642,
         n24643, n24644, n24645, n24646, n24647, n24648, n24649, n24650,
         n24651, n24652, n24653, n24654, n24655, n24656, n24657, n24658,
         n24659, n24660, n24661, n24662, n24663, n24664, n24665, n24666,
         n24667, n24668, n24669, n24670, n24671, n24672, n24673, n24674,
         n24675, n24676, n24677, n24678, n24679, n24680, n24681, n24682,
         n24683, n24684, n24685, n24686, n24687, n24688, n24689, n24690,
         n24691, n24692, n24693, n24694, n24695, n24696, n24697, n24698,
         n24699, n24700, n24701, n24702, n24703, n24704, n24705, n24706,
         n24707, n24708, n24709, n24710, n24711, n24712, n24713, n24714,
         n24715, n24716, n24717, n24718, n24719, n24720, n24721, n24722,
         n24723, n24724, n24725, n24726, n24727, n24728, n24729, n24730,
         n24731, n24732, n24733, n24734, n24735, n24736, n24737, n24738,
         n24739, n24740, n24741, n24742, n24743, n24744, n24745, n24746,
         n24747, n24748, n24749, n24750, n24751, n24752, n24753, n24754,
         n24755, n24756, n24757, n24758, n24759, n24760, n24761, n24762,
         n24763, n24764, n24765, n24766, n24767, n24768, n24769, n24770,
         n24771, n24772, n24773, n24774, n24775, n24776, n24777, n24778,
         n24779, n24780, n24781, n24782, n24783, n24784, n24785, n24786,
         n24787, n24788, n24789, n24790, n24791, n24792, n24793, n24794,
         n24795, n24796, n24797, n24798, n24799, n24800, n24801, n24802,
         n24803, n24804, n24805, n24806, n24807, n24808, n24809, n24810,
         n24811, n24812, n24813, n24814, n24815, n24816, n24817, n24818,
         n24819, n24820, n24821, n24822, n24823, n24824, n24825, n24826,
         n24827, n24828, n24829, n24830, n24831, n24832, n24833, n24834,
         n24835, n24836, n24837, n24838, n24839, n24840, n24841, n24842,
         n24843, n24844, n24845, n24846, n24847, n24848, n24849, n24850,
         n24851, n24852, n24853, n24854, n24855, n24856, n24857, n24858,
         n24859, n24860, n24861, n24862, n24863, n24864, n24865, n24866,
         n24867, n24868, n24869, n24870, n24871, n24872, n24873, n24874,
         n24875, n24876, n24877, n24878, n24879, n24880, n24881, n24882,
         n24883, n24884, n24885, n24886, n24887, n24888, n24889, n24890,
         n24891, n24892, n24893, n24894, n24895, n24896, n24897, n24898,
         n24899, n24900, n24901, n24902, n24903, n24904, n24905, n24906,
         n24907, n24908, n24909, n24910, n24911, n24912, n24913, n24914,
         n24915, n24916, n24917, n24918, n24919, n24920, n24921, n24922,
         n24923, n24924, n24925, n24926, n24927, n24928, n24929, n24930,
         n24931, n24932, n24933, n24934, n24935, n24936, n24937, n24938,
         n24939, n24940, n24941, n24942, n24943, n24944, n24945, n24946,
         n24947, n24948, n24949, n24950, n24951, n24952, n24953, n24954,
         n24955, n24956, n24957, n24958, n24959, n24960, n24961, n24962,
         n24963, n24964, n24965, n24966, n24967, n24968, n24969, n24970,
         n24971, n24972, n24973, n24974, n24975, n24976, n24977, n24978,
         n24979, n24980, n24981, n24982, n24983, n24984, n24985, n24986,
         n24987, n24988, n24989, n24990, n24991, n24992, n24993, n24994,
         n24995, n24996, n24997, n24998, n24999, n25000, n25001, n25002,
         n25003, n25004, n25005, n25006, n25007, n25008, n25009, n25010,
         n25011, n25012, n25013, n25014, n25015, n25016, n25017, n25018,
         n25019, n25020, n25021, n25022, n25023, n25024, n25025, n25026,
         n25027, n25028, n25029, n25030, n25031, n25032, n25033, n25034,
         n25035, n25036, n25037, n25038, n25039, n25040, n25041, n25042,
         n25043, n25044, n25045, n25046, n25047, n25048, n25049, n25050,
         n25051, n25052, n25053, n25054, n25055, n25056, n25057, n25058,
         n25059, n25060, n25061, n25062, n25063, n25064, n25065, n25066,
         n25067, n25068, n25069, n25070, n25071, n25072, n25073, n25074,
         n25075, n25076, n25077, n25078, n25079, n25080, n25081, n25082,
         n25083, n25084, n25085, n25086, n25087, n25088, n25089, n25090,
         n25091, n25092, n25093, n25094, n25095, n25096, n25097, n25098,
         n25099, n25100, n25101, n25102, n25103, n25104, n25105, n25106,
         n25107, n25108, n25109, n25110, n25111, n25112, n25113, n25114,
         n25115, n25116, n25117, n25118, n25119, n25120, n25121, n25122,
         n25123, n25124, n25125, n25126, n25127, n25128, n25129, n25130,
         n25131, n25132, n25133, n25134, n25135, n25136, n25137, n25138,
         n25139, n25140, n25141, n25142, n25143, n25144, n25145, n25146,
         n25147, n25148, n25149, n25150, n25151, n25152, n25153, n25154,
         n25155, n25156, n25157, n25158, n25159, n25160, n25161, n25162,
         n25163, n25164, n25165, n25166, n25167, n25168, n25169, n25170,
         n25171, n25172, n25173, n25174, n25175, n25176, n25177, n25178,
         n25179, n25180, n25181, n25182, n25183, n25184, n25185, n25186,
         n25187, n25188, n25189, n25190, n25191, n25192, n25193, n25194,
         n25195, n25196, n25197, n25198, n25199, n25200, n25201, n25202,
         n25203, n25204, n25205, n25206, n25207, n25208, n25209, n25210,
         n25211, n25212, n25213, n25214, n25215, n25216, n25217, n25218,
         n25219, n25220, n25221, n25222, n25223, n25224, n25225, n25226,
         n25227, n25228, n25229, n25230, n25231, n25232, n25233, n25234,
         n25235, n25236, n25237, n25238, n25239, n25240, n25241, n25242,
         n25243, n25244, n25245, n25246, n25247, n25248, n25249, n25250,
         n25251, n25252, n25253, n25254, n25255, n25256, n25257, n25258,
         n25259, n25260, n25261, n25262, n25263, n25264, n25265, n25266,
         n25267, n25268, n25269, n25270, n25271, n25272, n25273, n25274,
         n25275, n25276, n25277, n25278, n25279, n25280, n25281, n25282,
         n25283, n25284, n25285, n25286, n25287, n25288, n25289, n25290,
         n25291, n25292, n25293, n25294, n25295, n25296, n25297, n25298,
         n25299, n25300, n25301, n25302, n25303, n25304, n25305, n25306,
         n25307, n25308, n25309, n25310, n25311, n25312, n25313, n25314,
         n25315, n25316, n25317, n25318, n25319, n25320, n25321, n25322,
         n25323, n25324, n25325, n25326, n25327, n25328, n25329, n25330,
         n25331, n25332, n25333, n25334, n25335, n25336, n25337, n25338,
         n25339, n25340, n25341, n25342, n25343, n25344, n25345, n25346,
         n25347, n25348, n25349, n25350, n25351, n25352, n25353, n25354,
         n25355, n25356, n25357, n25358, n25359, n25360, n25361, n25362,
         n25363, n25364, n25365, n25366, n25367, n25368, n25369, n25370,
         n25371, n25372, n25373, n25374, n25375, n25376, n25377, n25378,
         n25379, n25380, n25381, n25382, n25383, n25384, n25385, n25386,
         n25387, n25388, n25389, n25390, n25391, n25392, n25393, n25394,
         n25395, n25396, n25397, n25398, n25399, n25400, n25401, n25402,
         n25403, n25404, n25405, n25406, n25407, n25408, n25409, n25410,
         n25411, n25412, n25413, n25414, n25415, n25416, n25417, n25418,
         n25419, n25420, n25421, n25422, n25423, n25424, n25425, n25426,
         n25427, n25428, n25429, n25430, n25431, n25432, n25433, n25434,
         n25435, n25436, n25437, n25438, n25439, n25440, n25441, n25442,
         n25443, n25444, n25445, n25446, n25447, n25448, n25449, n25450,
         n25451, n25452, n25453, n25454, n25455, n25456, n25457, n25458,
         n25459, n25460, n25461, n25462, n25463, n25464, n25465, n25466,
         n25467, n25468, n25469, n25470, n25471, n25472, n25473, n25474,
         n25475, n25476, n25477, n25478, n25479, n25480, n25481, n25482,
         n25483, n25484, n25485, n25486, n25487, n25488, n25489, n25490,
         n25491, n25492, n25493, n25494, n25495, n25496, n25497, n25498,
         n25499, n25500, n25501, n25502, n25503, n25504, n25505, n25506,
         n25507, n25508, n25509, n25510, n25511, n25512, n25513, n25514,
         n25515, n25516, n25517, n25518, n25519, n25520, n25521, n25522,
         n25523, n25524, n25525, n25526, n25527, n25528, n25529, n25530,
         n25531, n25532, n25533, n25534, n25535, n25536, n25537, n25538,
         n25539, n25540, n25541, n25542, n25543, n25544, n25545, n25546,
         n25547, n25548, n25549, n25550, n25551, n25552, n25553, n25554,
         n25555, n25556, n25557, n25558, n25559, n25560, n25561, n25562,
         n25563, n25564, n25565, n25566, n25567, n25568, n25569, n25570,
         n25571, n25572, n25573, n25574, n25575, n25576, n25577, n25578,
         n25579, n25580, n25581, n25582, n25583, n25584, n25585, n25586,
         n25587, n25588, n25589, n25590, n25591, n25592, n25593, n25594,
         n25595, n25596, n25597, n25598, n25599, n25600, n25601, n25602,
         n25603, n25604, n25605, n25606, n25607, n25608, n25609, n25610,
         n25611, n25612, n25613, n25614, n25615, n25616, n25617, n25618,
         n25619, n25620, n25621, n25622, n25623, n25624, n25625, n25626,
         n25627, n25628, n25629, n25630, n25631, n25632, n25633, n25634,
         n25635, n25636, n25637, n25638, n25639, n25640, n25641, n25642,
         n25643, n25644, n25645, n25646, n25647, n25648, n25649, n25650,
         n25651, n25652, n25653, n25654, n25655, n25656, n25657, n25658,
         n25659, n25660, n25661, n25662, n25663, n25664, n25665, n25666,
         n25667, n25668, n25669, n25670, n25671, n25672, n25673, n25674,
         n25675, n25676, n25677, n25678, n25679, n25680, n25681, n25682,
         n25683, n25684, n25685, n25686, n25687, n25688, n25689, n25690,
         n25691, n25692, n25693, n25694, n25695, n25696, n25697, n25698,
         n25699, n25700, n25701, n25702, n25703, n25704, n25705, n25706,
         n25707, n25708, n25709, n25710, n25711, n25712, n25713, n25714,
         n25715, n25716, n25717, n25718, n25719, n25720, n25721, n25722,
         n25723, n25724, n25725, n25726, n25727, n25728, n25729, n25730,
         n25731, n25732, n25733, n25734, n25735, n25736, n25737, n25738,
         n25739, n25740, n25741, n25742, n25743, n25744, n25745, n25746,
         n25747, n25748, n25749, n25750, n25751, n25752, n25753, n25754,
         n25755, n25756, n25757, n25758, n25759, n25760, n25761, n25762,
         n25763, n25764, n25765, n25766, n25767, n25768, n25769, n25770,
         n25771, n25772, n25773, n25774, n25775, n25776, n25777, n25778,
         n25779, n25780, n25781, n25782, n25783, n25784, n25785, n25786,
         n25787, n25788, n25789, n25790, n25791, n25792, n25793, n25794,
         n25795, n25796, n25797, n25798, n25799, n25800, n25801, n25802,
         n25803, n25804, n25805, n25806, n25807, n25808, n25809, n25810,
         n25811, n25812, n25813, n25814, n25815, n25816, n25817, n25818,
         n25819, n25820, n25821, n25822, n25823, n25824, n25825, n25826,
         n25827, n25828, n25829, n25830, n25831, n25832, n25833, n25834,
         n25835, n25836, n25837, n25838, n25839, n25840, n25841, n25842,
         n25843, n25844, n25845, n25846, n25847, n25848, n25849, n25850,
         n25851, n25852, n25853, n25854, n25855, n25856, n25857, n25858,
         n25859, n25860, n25861, n25862, n25863, n25864, n25865, n25866,
         n25867, n25868, n25869, n25870, n25871, n25872, n25873, n25874,
         n25875, n25876, n25877, n25878, n25879, n25880, n25881, n25882,
         n25883, n25884, n25885, n25886, n25887, n25888, n25889, n25890,
         n25891, n25892, n25893, n25894, n25895, n25896, n25897, n25898,
         n25899, n25900, n25901, n25902, n25903, n25904, n25905, n25906,
         n25907, n25908, n25909, n25910, n25911, n25912, n25913, n25914,
         n25915, n25916, n25917, n25918, n25919, n25920, n25921, n25922,
         n25923, n25924, n25925, n25926, n25927, n25928, n25929, n25930,
         n25931, n25932, n25933, n25934, n25935, n25936, n25937, n25938,
         n25939, n25940, n25941, n25942, n25943, n25944, n25945, n25946,
         n25947, n25948, n25949, n25950, n25951, n25952, n25953, n25954,
         n25955, n25956, n25957, n25958, n25959, n25960, n25961, n25962,
         n25963, n25964, n25965, n25966, n25967, n25968, n25969, n25970,
         n25971, n25972, n25973, n25974, n25975, n25976, n25977, n25978,
         n25979, n25980, n25981, n25982, n25983, n25984, n25985, n25986,
         n25987, n25988, n25989, n25990, n25991, n25992, n25993, n25994,
         n25995, n25996, n25997, n25998, n25999, n26000, n26001, n26002,
         n26003, n26004, n26005, n26006, n26007, n26008, n26009, n26010,
         n26011, n26012, n26013, n26014, n26015, n26016, n26017, n26018,
         n26019, n26020, n26021, n26022, n26023, n26024, n26025, n26026,
         n26027, n26028, n26029, n26030, n26031, n26032, n26033, n26034,
         n26035, n26036, n26037, n26038, n26039, n26040, n26041, n26042,
         n26043, n26044, n26045, n26046, n26047, n26048, n26049, n26050,
         n26051, n26052, n26053, n26054, n26055, n26056, n26057, n26058,
         n26059, n26060, n26061, n26062, n26063, n26064, n26065, n26066,
         n26067, n26068, n26069, n26070, n26071, n26072, n26073, n26074,
         n26075, n26076, n26077, n26078, n26079, n26080, n26081, n26082,
         n26083, n26084, n26085, n26086, n26087, n26088, n26089, n26090,
         n26091, n26092, n26093, n26094, n26095, n26096, n26097, n26098,
         n26099, n26100, n26101, n26102, n26103, n26104, n26105, n26106,
         n26107, n26108, n26109, n26110, n26111, n26112, n26113, n26114,
         n26115, n26116, n26117, n26118, n26119, n26120, n26121, n26122,
         n26123, n26124, n26125, n26126, n26127, n26128, n26129, n26130,
         n26131, n26132, n26133, n26134, n26135, n26136, n26137, n26138,
         n26139, n26140, n26141, n26142, n26143, n26144, n26145, n26146,
         n26147, n26148, n26149, n26150, n26151, n26152, n26153, n26154,
         n26155, n26156, n26157, n26158, n26159, n26160, n26161, n26162,
         n26163, n26164, n26165, n26166, n26167, n26168, n26169, n26170,
         n26171, n26172, n26173, n26174, n26175, n26176, n26177, n26178,
         n26179, n26180, n26181, n26182, n26183, n26184, n26185, n26186,
         n26187, n26188, n26189, n26190, n26191, n26192, n26193, n26194,
         n26195, n26196, n26197, n26198, n26199, n26200, n26201, n26202,
         n26203, n26204, n26205, n26206, n26207, n26208, n26209, n26210,
         n26211, n26212, n26213, n26214, n26215, n26216, n26217, n26218,
         n26219, n26220, n26221, n26222, n26223, n26224, n26225, n26226,
         n26227, n26228, n26229, n26230, n26231, n26232, n26233, n26234,
         n26235, n26236, n26237, n26238, n26239, n26240, n26241, n26242,
         n26243, n26244, n26245, n26246, n26247, n26248, n26249, n26250,
         n26251, n26252, n26253, n26254, n26255, n26256, n26257, n26258,
         n26259, n26260, n26261, n26262, n26263, n26264, n26265, n26266,
         n26267, n26268, n26269, n26270, n26271, n26272, n26273, n26274,
         n26275, n26276, n26277, n26278, n26279, n26280, n26281, n26282,
         n26283, n26284, n26285, n26286, n26287, n26288, n26289, n26290,
         n26291, n26292, n26293, n26294, n26295, n26296, n26297, n26298,
         n26299, n26300, n26301, n26302, n26303, n26304, n26305, n26306,
         n26307, n26308, n26309, n26310, n26311, n26312, n26313, n26314,
         n26315, n26316, n26317, n26318, n26319, n26320, n26321, n26322,
         n26323, n26324, n26325, n26326, n26327, n26328, n26329, n26330,
         n26331, n26332, n26333, n26334, n26335, n26336, n26337, n26338,
         n26339, n26340, n26341, n26342, n26343, n26344, n26345, n26346,
         n26347, n26348, n26349, n26350, n26351, n26352, n26353, n26354,
         n26355, n26356, n26357, n26358, n26359, n26360, n26361, n26362,
         n26363, n26364, n26365, n26366, n26367, n26368, n26369, n26370,
         n26371, n26372, n26373, n26374, n26375, n26376, n26377, n26378,
         n26379, n26380, n26381, n26382, n26383, n26384, n26385, n26386,
         n26387, n26388, n26389, n26390, n26391, n26392, n26393, n26394,
         n26395, n26396, n26397, n26398, n26399, n26400, n26401, n26402,
         n26403, n26404, n26405, n26406, n26407, n26408, n26409, n26410,
         n26411, n26412, n26413, n26414, n26415, n26416, n26417, n26418,
         n26419, n26420, n26421, n26422, n26423, n26424, n26425, n26426,
         n26427, n26428, n26429, n26430, n26431, n26432, n26433, n26434,
         n26435, n26436, n26437, n26438, n26439, n26440, n26441, n26442,
         n26443, n26444, n26445, n26446, n26447, n26448, n26449, n26450,
         n26451, n26452, n26453, n26454, n26455, n26456, n26457, n26458,
         n26459, n26460, n26461, n26462, n26463, n26464, n26465, n26466,
         n26467, n26468, n26469, n26470, n26471, n26472, n26473, n26474,
         n26475, n26476, n26477, n26478, n26479, n26480, n26481, n26482,
         n26483, n26484, n26485, n26486, n26487, n26488, n26489, n26490,
         n26491, n26492, n26493, n26494, n26495, n26496, n26497, n26498,
         n26499, n26500, n26501, n26502, n26503, n26504, n26505, n26506,
         n26507, n26508, n26509, n26510, n26511, n26512, n26513, n26514,
         n26515, n26516, n26517, n26518, n26519, n26520, n26521, n26522,
         n26523, n26524, n26525, n26526, n26527, n26528, n26529, n26530,
         n26531, n26532, n26533, n26534, n26535, n26536, n26537, n26538,
         n26539, n26540, n26541, n26542, n26543, n26544, n26545, n26546,
         n26547, n26548, n26549, n26550, n26551, n26552, n26553, n26554,
         n26555, n26556, n26557, n26558, n26559, n26560, n26561, n26562,
         n26563, n26564, n26565, n26566, n26567, n26568, n26569, n26570,
         n26571, n26572, n26573, n26574, n26575, n26576, n26577, n26578,
         n26579, n26580, n26581, n26582, n26583, n26584, n26585, n26586,
         n26587, n26588, n26589, n26590, n26591, n26592, n26593, n26594,
         n26595, n26596, n26597, n26598, n26599, n26600, n26601, n26602,
         n26603, n26604, n26605, n26606, n26607, n26608, n26609, n26610,
         n26611, n26612, n26613, n26614, n26615, n26616, n26617, n26618,
         n26619, n26620, n26621, n26622, n26623, n26624, n26625, n26626,
         n26627, n26628, n26629, n26630, n26631, n26632, n26633, n26634,
         n26635, n26636, n26637, n26638, n26639, n26640, n26641, n26642,
         n26643, n26644, n26645, n26646, n26647, n26648, n26649, n26650,
         n26651, n26652, n26653, n26654, n26655, n26656, n26657, n26658,
         n26659, n26660, n26661, n26662, n26663, n26664, n26665, n26666,
         n26667, n26668, n26669, n26670, n26671, n26672, n26673, n26674,
         n26675, n26676, n26677, n26678, n26679, n26680, n26681, n26682,
         n26683, n26684, n26685, n26686, n26687, n26688, n26689, n26690,
         n26691, n26692, n26693, n26694, n26695, n26696, n26697, n26698,
         n26699, n26700, n26701, n26702, n26703, n26704, n26705, n26706,
         n26707, n26708, n26709, n26710, n26711, n26712, n26713, n26714,
         n26715, n26716, n26717, n26718, n26719, n26720, n26721, n26722,
         n26723, n26724, n26725, n26726, n26727, n26728, n26729, n26730,
         n26731, n26732, n26733, n26734, n26735, n26736, n26737, n26738,
         n26739, n26740, n26741, n26742, n26743, n26744, n26745, n26746,
         n26747, n26748, n26749, n26750, n26751, n26752, n26753, n26754,
         n26755, n26756, n26757, n26758, n26759, n26760, n26761, n26762,
         n26763, n26764, n26765, n26766, n26767, n26768, n26769, n26770,
         n26771, n26772, n26773, n26774, n26775, n26776, n26777, n26778,
         n26779, n26780, n26781, n26782, n26783, n26784, n26785, n26786,
         n26787, n26788, n26789, n26790, n26791, n26792, n26793, n26794,
         n26795, n26796, n26797, n26798, n26799, n26800, n26801, n26802,
         n26803, n26804, n26805, n26806, n26807, n26808, n26809, n26810,
         n26811, n26812, n26813, n26814, n26815, n26816, n26817, n26818,
         n26819, n26820, n26821, n26822, n26823, n26824, n26825, n26826,
         n26827, n26828, n26829, n26830, n26831, n26832, n26833, n26834,
         n26835, n26836, n26837, n26838, n26839, n26840, n26841, n26842,
         n26843, n26844, n26845, n26846, n26847, n26848, n26849, n26850,
         n26851, n26852, n26853, n26854, n26855, n26856, n26857, n26858,
         n26859, n26860, n26861, n26862, n26863, n26864, n26865, n26866,
         n26867, n26868, n26869, n26870, n26871, n26872, n26873, n26874,
         n26875, n26876, n26877, n26878, n26879, n26880, n26881, n26882,
         n26883, n26884, n26885, n26886, n26887, n26888, n26889, n26890,
         n26891, n26892, n26893, n26894, n26895, n26896, n26897, n26898,
         n26899, n26900, n26901, n26902, n26903, n26904, n26905, n26906,
         n26907, n26908, n26909, n26910, n26911, n26912, n26913, n26914,
         n26915, n26916, n26917, n26918, n26919, n26920, n26921, n26922,
         n26923, n26924, n26925, n26926, n26927, n26928, n26929, n26930,
         n26931, n26932, n26933, n26934, n26935, n26936, n26937, n26938,
         n26939, n26940, n26941, n26942, n26943, n26944, n26945, n26946,
         n26947, n26948, n26949, n26950, n26951, n26952, n26953, n26954,
         n26955, n26956, n26957, n26958, n26959, n26960, n26961, n26962,
         n26963, n26964, n26965, n26966, n26967, n26968, n26969, n26970,
         n26971, n26972, n26973, n26974, n26975, n26976, n26977, n26978,
         n26979, n26980, n26981, n26982, n26983, n26984, n26985, n26986,
         n26987, n26988, n26989, n26990, n26991, n26992, n26993, n26994,
         n26995, n26996, n26997, n26998, n26999, n27000, n27001, n27002,
         n27003, n27004, n27005, n27006, n27007, n27008, n27009, n27010,
         n27011, n27012, n27013, n27014, n27015, n27016, n27017, n27018,
         n27019, n27020, n27021, n27022, n27023, n27024, n27025, n27026,
         n27027, n27028, n27029, n27030, n27031, n27032, n27033, n27034,
         n27035, n27036, n27037, n27038, n27039, n27040, n27041, n27042,
         n27043, n27044, n27045, n27046, n27047, n27048, n27049, n27050,
         n27051, n27052, n27053, n27054, n27055, n27056, n27057, n27058,
         n27059, n27060, n27061, n27062, n27063, n27064, n27065, n27066,
         n27067, n27068, n27069, n27070, n27071, n27072, n27073, n27074,
         n27075, n27076, n27077, n27078, n27079, n27080, n27081, n27082,
         n27083, n27084, n27085, n27086, n27087, n27088, n27089, n27090,
         n27091, n27092, n27093, n27094, n27095, n27096, n27097, n27098,
         n27099, n27100, n27101, n27102, n27103, n27104, n27105, n27106,
         n27107, n27108, n27109, n27110, n27111, n27112, n27113, n27114,
         n27115, n27116, n27117, n27118, n27119, n27120, n27121, n27122,
         n27123, n27124, n27125, n27126, n27127, n27128, n27129, n27130,
         n27131, n27132, n27133, n27134, n27135, n27136, n27137, n27138,
         n27139, n27140, n27141, n27142, n27143, n27144, n27145, n27146,
         n27147, n27148, n27149, n27150, n27151, n27152, n27153, n27154,
         n27155, n27156, n27157, n27158, n27159, n27160, n27161, n27162,
         n27163, n27164, n27165, n27166, n27167, n27168, n27169, n27170,
         n27171, n27172, n27173, n27174, n27175, n27176, n27177, n27178,
         n27179, n27180, n27181, n27182, n27183, n27184, n27185, n27186,
         n27187, n27188, n27189, n27190, n27191, n27192, n27193, n27194,
         n27195, n27196, n27197, n27198, n27199, n27200, n27201, n27202,
         n27203, n27204, n27205, n27206, n27207, n27208, n27209, n27210,
         n27211, n27212, n27213, n27214, n27215, n27216, n27217, n27218,
         n27219, n27220, n27221, n27222, n27223, n27224, n27225, n27226,
         n27227, n27228, n27229, n27230, n27231, n27232, n27233, n27234,
         n27235, n27236, n27237, n27238, n27239, n27240, n27241, n27242,
         n27243, n27244, n27245, n27246, n27247, n27248, n27249, n27250,
         n27251, n27252, n27253, n27254, n27255, n27256, n27257, n27258,
         n27259, n27260, n27261, n27262, n27263, n27264, n27265, n27266,
         n27267, n27268, n27269, n27270, n27271, n27272, n27273, n27274,
         n27275, n27276, n27277, n27278, n27279, n27280, n27281, n27282,
         n27283, n27284, n27285, n27286, n27287, n27288, n27289, n27290,
         n27291, n27292, n27293, n27294, n27295, n27296, n27297, n27298,
         n27299, n27300, n27301, n27302, n27303, n27304, n27305, n27306,
         n27307, n27308, n27309, n27310, n27311, n27312, n27313, n27314,
         n27315, n27316, n27317, n27318, n27319, n27320, n27321, n27322,
         n27323, n27324, n27325, n27326, n27327, n27328, n27329, n27330,
         n27331, n27332, n27333, n27334, n27335, n27336, n27337, n27338,
         n27339, n27340, n27341, n27342, n27343, n27344, n27345, n27346,
         n27347, n27348, n27349, n27350, n27351, n27352, n27353, n27354,
         n27355, n27356, n27357, n27358, n27359, n27360, n27361, n27362,
         n27363, n27364, n27365, n27366, n27367, n27368, n27369, n27370,
         n27371, n27372, n27373, n27374, n27375, n27376, n27377, n27378,
         n27379, n27380, n27381, n27382, n27383, n27384, n27385, n27386,
         n27387, n27388, n27389, n27390, n27391, n27392, n27393, n27394,
         n27395, n27396, n27397, n27398, n27399, n27400, n27401, n27402,
         n27403, n27404, n27405, n27406, n27407, n27408, n27409, n27410,
         n27411, n27412, n27413, n27414, n27415, n27416, n27417, n27418,
         n27419, n27420, n27421, n27422, n27423, n27424, n27425, n27426,
         n27427, n27428, n27429, n27430, n27431, n27432, n27433, n27434,
         n27435, n27436, n27437, n27438, n27439, n27440, n27441, n27442,
         n27443, n27444, n27445, n27446, n27447, n27448, n27449, n27450,
         n27451, n27452, n27453, n27454, n27455, n27456, n27457, n27458,
         n27459, n27460, n27461, n27462, n27463, n27464, n27465, n27466,
         n27467, n27468, n27469, n27470, n27471, n27472, n27473, n27474,
         n27475, n27476, n27477, n27478, n27479, n27480, n27481, n27482,
         n27483, n27484, n27485, n27486, n27487, n27488, n27489, n27490,
         n27491, n27492, n27493, n27494, n27495, n27496, n27497, n27498,
         n27499, n27500, n27501, n27502, n27503, n27504, n27505, n27506,
         n27507, n27508, n27509, n27510, n27511, n27512, n27513, n27514,
         n27515, n27516, n27517, n27518, n27519, n27520, n27521, n27522,
         n27523, n27524, n27525, n27526, n27527, n27528, n27529, n27530,
         n27531, n27532, n27533, n27534, n27535, n27536, n27537, n27538,
         n27539, n27540, n27541, n27542, n27543, n27544, n27545, n27546,
         n27547, n27548, n27549, n27550, n27551, n27552, n27553, n27554,
         n27555, n27556, n27557, n27558, n27559, n27560, n27561, n27562,
         n27563, n27564, n27565, n27566, n27567, n27568, n27569, n27570,
         n27571, n27572, n27573, n27574, n27575, n27576, n27577, n27578,
         n27579, n27580, n27581, n27582, n27583, n27584, n27585, n27586,
         n27587, n27588, n27589, n27590, n27591, n27592, n27593, n27594,
         n27595, n27596, n27597, n27598, n27599, n27600, n27601, n27602,
         n27603, n27604, n27605, n27606, n27607, n27608, n27609, n27610,
         n27611, n27612, n27613, n27614, n27615, n27616, n27617, n27618,
         n27619, n27620, n27621, n27622, n27623, n27624, n27625, n27626,
         n27627, n27628, n27629, n27630, n27631, n27632, n27633, n27634,
         n27635, n27636, n27637, n27638, n27639, n27640, n27641, n27642,
         n27643, n27644, n27645, n27646, n27647, n27648, n27649, n27650,
         n27651, n27652, n27653, n27654, n27655, n27656, n27657, n27658,
         n27659, n27660, n27661, n27662, n27663, n27664, n27665, n27666,
         n27667, n27668, n27669, n27670, n27671, n27672, n27673, n27674,
         n27675, n27676, n27677, n27678, n27679, n27680, n27681, n27682,
         n27683, n27684, n27685, n27686, n27687, n27688, n27689, n27690,
         n27691, n27692, n27693, n27694, n27695, n27696, n27697, n27698,
         n27699, n27700, n27701, n27702, n27703, n27704, n27705, n27706,
         n27707, n27708, n27709, n27710, n27711, n27712, n27713, n27714,
         n27715, n27716, n27717, n27718, n27719, n27720, n27721, n27722,
         n27723, n27724, n27725, n27726, n27727, n27728, n27729, n27730,
         n27731, n27732, n27733, n27734, n27735, n27736, n27737, n27738,
         n27739, n27740, n27741, n27742, n27743, n27744, n27745, n27746,
         n27747, n27748, n27749, n27750, n27751, n27752, n27753, n27754,
         n27755, n27756, n27757, n27758, n27759, n27760, n27761, n27762,
         n27763, n27764, n27765, n27766, n27767, n27768, n27769, n27770,
         n27771, n27772, n27773, n27774, n27775, n27776, n27777, n27778,
         n27779, n27780, n27781, n27782, n27783, n27784, n27785, n27786,
         n27787, n27788, n27789, n27790, n27791, n27792, n27793, n27794,
         n27795, n27796, n27797, n27798, n27799, n27800, n27801, n27802,
         n27803, n27804, n27805, n27806, n27807, n27808, n27809, n27810,
         n27811, n27812, n27813, n27814, n27815, n27816, n27817, n27818,
         n27819, n27820, n27821, n27822, n27823, n27824, n27825, n27826,
         n27827, n27828, n27829, n27830, n27831, n27832, n27833, n27834,
         n27835, n27836, n27837, n27838, n27839, n27840, n27841, n27842,
         n27843, n27844, n27845, n27846, n27847, n27848, n27849, n27850,
         n27851, n27852, n27853, n27854, n27855, n27856, n27857, n27858,
         n27859, n27860, n27861, n27862, n27863, n27864, n27865, n27866,
         n27867, n27868, n27869, n27870, n27871, n27872, n27873, n27874,
         n27875, n27876, n27877, n27878, n27879, n27880, n27881, n27882,
         n27883, n27884, n27885, n27886, n27887, n27888, n27889, n27890,
         n27891, n27892, n27893, n27894, n27895, n27896, n27897, n27898,
         n27899, n27900, n27901, n27902, n27903, n27904, n27905, n27906,
         n27907, n27908, n27909, n27910, n27911, n27912, n27913, n27914,
         n27915, n27916, n27917, n27918, n27919, n27920, n27921, n27922,
         n27923, n27924, n27925, n27926, n27927, n27928, n27929, n27930,
         n27931, n27932, n27933, n27934, n27935, n27936, n27937, n27938,
         n27939, n27940, n27941, n27942, n27943, n27944, n27945, n27946,
         n27947, n27948, n27949, n27950, n27951, n27952, n27953, n27954,
         n27955, n27956, n27957, n27958, n27959, n27960, n27961, n27962,
         n27963, n27964, n27965, n27966, n27967, n27968, n27969, n27970,
         n27971, n27972, n27973, n27974, n27975, n27976, n27977, n27978,
         n27979, n27980, n27981, n27982, n27983, n27984, n27985, n27986,
         n27987, n27988, n27989, n27990, n27991, n27992, n27993, n27994,
         n27995, n27996, n27997, n27998, n27999, n28000, n28001, n28002,
         n28003, n28004, n28005, n28006, n28007, n28008, n28009, n28010,
         n28011, n28012, n28013, n28014, n28015, n28016, n28017, n28018,
         n28019, n28020, n28021, n28022, n28023, n28024, n28025, n28026,
         n28027, n28028, n28029, n28030, n28031, n28032, n28033, n28034,
         n28035, n28036, n28037, n28038, n28039, n28040, n28041, n28042,
         n28043, n28044, n28045, n28046, n28047, n28048, n28049, n28050,
         n28051, n28052, n28053, n28054, n28055, n28056, n28057, n28058,
         n28059, n28060, n28061, n28062, n28063, n28064, n28065, n28066,
         n28067, n28068, n28069, n28070, n28071, n28072, n28073, n28074,
         n28075, n28076, n28077, n28078, n28079, n28080, n28081, n28082,
         n28083, n28084, n28085, n28086, n28087, n28088, n28089, n28090,
         n28091, n28092, n28093, n28094, n28095, n28096, n28097, n28098,
         n28099, n28100, n28101, n28102, n28103, n28104, n28105, n28106,
         n28107, n28108, n28109, n28110, n28111, n28112, n28113, n28114,
         n28115, n28116, n28117, n28118, n28119, n28120, n28121, n28122,
         n28123, n28124, n28125, n28126, n28127, n28128, n28129, n28130,
         n28131, n28132, n28133, n28134, n28135, n28136, n28137, n28138,
         n28139, n28140, n28141, n28142, n28143, n28144, n28145, n28146,
         n28147, n28148, n28149, n28150, n28151, n28152, n28153, n28154,
         n28155, n28156, n28157, n28158, n28159, n28160, n28161, n28162,
         n28163, n28164, n28165, n28166, n28167, n28168, n28169, n28170,
         n28171, n28172, n28173, n28174, n28175, n28176, n28177, n28178,
         n28179, n28180, n28181, n28182, n28183, n28184, n28185, n28186,
         n28187, n28188, n28189, n28190, n28191, n28192, n28193, n28194,
         n28195, n28196, n28197, n28198, n28199, n28200, n28201, n28202,
         n28203, n28204, n28205, n28206, n28207, n28208, n28209, n28210,
         n28211, n28212, n28213, n28214, n28215, n28216, n28217, n28218,
         n28219, n28220, n28221, n28222, n28223, n28224, n28225, n28226,
         n28227, n28228, n28229, n28230, n28231, n28232, n28233, n28234,
         n28235, n28236, n28237, n28238, n28239, n28240, n28241, n28242,
         n28243, n28244, n28245, n28246, n28247, n28248, n28249, n28250,
         n28251, n28252, n28253, n28254, n28255, n28256, n28257, n28258,
         n28259, n28260, n28261, n28262, n28263, n28264, n28265, n28266,
         n28267, n28268, n28269, n28270, n28271, n28272, n28273, n28274,
         n28275, n28276, n28277, n28278, n28279, n28280, n28281, n28282,
         n28283, n28284, n28285, n28286, n28287, n28288, n28289, n28290,
         n28291, n28292, n28293, n28294, n28295, n28296, n28297, n28298,
         n28299, n28300, n28301, n28302, n28303, n28304, n28305, n28306,
         n28307, n28308, n28309, n28310, n28311, n28312, n28313, n28314,
         n28315, n28316, n28317, n28318, n28319, n28320, n28321, n28322,
         n28323, n28324, n28325, n28326, n28327, n28328, n28329, n28330,
         n28331, n28332, n28333, n28334, n28335, n28336, n28337, n28338,
         n28339, n28340, n28341, n28342, n28343, n28344, n28345, n28346,
         n28347, n28348, n28349, n28350, n28351, n28352, n28353, n28354,
         n28355, n28356, n28357, n28358, n28359, n28360, n28361, n28362,
         n28363, n28364, n28365, n28366, n28367, n28368, n28369, n28370,
         n28371, n28372, n28373, n28374, n28375, n28376, n28377, n28378,
         n28379, n28380, n28381, n28382, n28383, n28384, n28385, n28386,
         n28387, n28388, n28389, n28390, n28391, n28392, n28393, n28394,
         n28395, n28396, n28397, n28398, n28399, n28400, n28401, n28402,
         n28403, n28404, n28405, n28406, n28407, n28408, n28409, n28410,
         n28411, n28412, n28413, n28414, n28415, n28416, n28417, n28418,
         n28419, n28420, n28421, n28422, n28423, n28424, n28425, n28426,
         n28427, n28428, n28429, n28430, n28431, n28432, n28433, n28434,
         n28435, n28436, n28437, n28438, n28439, n28440, n28441, n28442,
         n28443, n28444, n28445, n28446, n28447, n28448, n28449, n28450,
         n28451, n28452, n28453, n28454, n28455, n28456, n28457, n28458,
         n28459, n28460, n28461, n28462, n28463, n28464, n28465, n28466,
         n28467, n28468, n28469, n28470, n28471, n28472, n28473, n28474,
         n28475, n28476, n28477, n28478, n28479, n28480, n28481, n28482,
         n28483, n28484, n28485, n28486, n28487, n28488, n28489, n28490,
         n28491, n28492, n28493, n28494, n28495, n28496, n28497, n28498,
         n28499, n28500, n28501, n28502, n28503, n28504, n28505, n28506,
         n28507, n28508, n28509, n28510, n28511, n28512, n28513, n28514,
         n28515, n28516, n28517, n28518, n28519, n28520, n28521, n28522,
         n28523, n28524, n28525, n28526, n28527, n28528, n28529, n28530,
         n28531, n28532, n28533, n28534, n28535, n28536, n28537, n28538,
         n28539, n28540, n28541, n28542, n28543, n28544, n28545, n28546,
         n28547, n28548, n28549, n28550, n28551, n28552, n28553, n28554,
         n28555, n28556, n28557, n28558, n28559, n28560, n28561, n28562,
         n28563, n28564, n28565, n28566, n28567, n28568, n28569, n28570,
         n28571, n28572, n28573, n28574, n28575, n28576, n28577, n28578,
         n28579, n28580, n28581, n28582, n28583, n28584, n28585, n28586,
         n28587, n28588, n28589, n28590, n28591, n28592, n28593, n28594,
         n28595, n28596, n28597, n28598, n28599, n28600, n28601, n28602,
         n28603, n28604, n28605, n28606, n28607, n28608, n28609, n28610,
         n28611, n28612, n28613, n28614, n28615, n28616, n28617, n28618,
         n28619, n28620, n28621, n28622, n28623, n28624, n28625, n28626,
         n28627, n28628, n28629, n28630, n28631, n28632, n28633, n28634,
         n28635, n28636, n28637, n28638, n28639, n28640, n28641, n28642,
         n28643, n28644, n28645, n28646, n28647, n28648, n28649, n28650,
         n28651, n28652, n28653, n28654, n28655, n28656, n28657, n28658,
         n28659, n28660, n28661, n28662, n28663, n28664, n28665, n28666,
         n28667, n28668, n28669, n28670, n28671, n28672, n28673, n28674,
         n28675, n28676, n28677, n28678, n28679, n28680, n28681, n28682,
         n28683, n28684, n28685, n28686, n28687, n28688, n28689, n28690,
         n28691, n28692, n28693, n28694, n28695, n28696, n28697, n28698,
         n28699, n28700, n28701, n28702, n28703, n28704, n28705, n28706,
         n28707, n28708, n28709, n28710, n28711, n28712, n28713, n28714,
         n28715, n28716, n28717, n28718, n28719, n28720, n28721, n28722,
         n28723, n28724, n28725, n28726, n28727, n28728, n28729, n28730,
         n28731, n28732, n28733, n28734, n28735, n28736, n28737, n28738,
         n28739, n28740, n28741, n28742, n28743, n28744, n28745, n28746,
         n28747, n28748, n28749, n28750, n28751, n28752, n28753, n28754,
         n28755, n28756, n28757, n28758, n28759, n28760, n28761, n28762,
         n28763, n28764, n28765, n28766, n28767, n28768, n28769, n28770,
         n28771, n28772, n28773, n28774, n28775, n28776, n28777, n28778,
         n28779, n28780, n28781, n28782, n28783, n28784, n28785, n28786,
         n28787, n28788, n28789, n28790, n28791, n28792, n28793, n28794,
         n28795, n28796, n28797, n28798, n28799, n28800, n28801, n28802,
         n28803, n28804, n28805, n28806, n28807, n28808, n28809, n28810,
         n28811, n28812, n28813, n28814, n28815, n28816, n28817, n28818,
         n28819, n28820, n28821, n28822, n28823, n28824, n28825, n28826,
         n28827, n28828, n28829, n28830, n28831, n28832, n28833, n28834,
         n28835, n28836, n28837, n28838, n28839, n28840, n28841, n28842,
         n28843, n28844, n28845, n28846, n28847, n28848, n28849, n28850,
         n28851, n28852, n28853, n28854, n28855, n28856, n28857, n28858,
         n28859, n28860, n28861, n28862, n28863, n28864, n28865, n28866,
         n28867, n28868, n28869, n28870, n28871, n28872, n28873, n28874,
         n28875, n28876, n28877, n28878, n28879, n28880, n28881, n28882,
         n28883, n28884, n28885, n28886, n28887, n28888, n28889, n28890,
         n28891, n28892, n28893, n28894, n28895, n28896, n28897, n28898,
         n28899, n28900, n28901, n28902, n28903, n28904, n28905, n28906,
         n28907, n28908, n28909, n28910, n28911, n28912, n28913, n28914,
         n28915, n28916, n28917, n28918, n28919, n28920, n28921, n28922,
         n28923, n28924, n28925, n28926, n28927, n28928, n28929, n28930,
         n28931, n28932, n28933, n28934, n28935, n28936, n28937, n28938,
         n28939, n28940, n28941, n28942, n28943, n28944, n28945, n28946,
         n28947, n28948, n28949, n28950, n28951, n28952, n28953, n28954,
         n28955, n28956, n28957, n28958, n28959, n28960, n28961, n28962,
         n28963, n28964, n28965, n28966, n28967, n28968, n28969, n28970,
         n28971, n28972, n28973, n28974, n28975, n28976, n28977, n28978,
         n28979, n28980, n28981, n28982, n28983, n28984, n28985, n28986,
         n28987, n28988, n28989, n28990, n28991, n28992, n28993, n28994,
         n28995, n28996, n28997, n28998, n28999, n29000, n29001, n29002,
         n29003, n29004, n29005, n29006, n29007, n29008, n29009, n29010,
         n29011, n29012, n29013, n29014, n29015, n29016, n29017, n29018,
         n29019, n29020, n29021, n29022, n29023, n29024, n29025, n29026,
         n29027, n29028, n29029, n29030, n29031, n29032, n29033, n29034,
         n29035, n29036, n29037, n29038, n29039, n29040, n29041, n29042,
         n29043, n29044, n29045, n29046, n29047, n29048, n29049, n29050,
         n29051, n29052, n29053, n29054, n29055, n29056, n29057, n29058,
         n29059, n29060, n29061, n29062, n29063, n29064, n29065, n29066,
         n29067, n29068, n29069, n29070, n29071, n29072, n29073, n29074,
         n29075, n29076, n29077, n29078, n29079, n29080, n29081, n29082,
         n29083, n29084, n29085, n29086, n29087, n29088, n29089, n29090,
         n29091, n29092, n29093, n29094, n29095, n29096, n29097, n29098,
         n29099, n29100, n29101, n29102, n29103, n29104, n29105, n29106,
         n29107, n29108, n29109, n29110, n29111, n29112, n29113, n29114,
         n29115, n29116, n29117, n29118, n29119, n29120, n29121, n29122,
         n29123, n29124, n29125, n29126, n29127, n29128, n29129, n29130,
         n29131, n29132, n29133, n29134, n29135, n29136, n29137, n29138,
         n29139, n29140, n29141, n29142, n29143, n29144, n29145, n29146,
         n29147, n29148, n29149, n29150, n29151, n29152, n29153, n29154,
         n29155, n29156, n29157, n29158, n29159, n29160, n29161, n29162,
         n29163, n29164, n29165, n29166, n29167, n29168, n29169, n29170,
         n29171, n29172, n29173, n29174, n29175, n29176, n29177, n29178,
         n29179, n29180, n29181, n29182, n29183, n29184, n29185, n29186,
         n29187, n29188, n29189, n29190, n29191, n29192, n29193, n29194,
         n29195, n29196, n29197, n29198, n29199, n29200, n29201, n29202,
         n29203, n29204, n29205, n29206, n29207, n29208, n29209, n29210,
         n29211, n29212, n29213, n29214, n29215, n29216, n29217, n29218,
         n29219, n29220, n29221, n29222, n29223, n29224, n29225, n29226,
         n29227, n29228, n29229, n29230, n29231, n29232, n29233, n29234,
         n29235, n29236, n29237, n29238, n29239, n29240, n29241, n29242,
         n29243, n29244, n29245, n29246, n29247, n29248, n29249, n29250,
         n29251, n29252, n29253, n29254, n29255, n29256, n29257, n29258,
         n29259, n29260, n29261, n29262, n29263, n29264, n29265, n29266,
         n29267, n29268, n29269, n29270, n29271, n29272, n29273, n29274,
         n29275, n29276, n29277, n29278, n29279, n29280, n29281, n29282,
         n29283, n29284, n29285, n29286, n29287, n29288, n29289, n29290,
         n29291, n29292, n29293, n29294, n29295, n29296, n29297, n29298,
         n29299, n29300, n29301, n29302, n29303, n29304, n29305, n29306,
         n29307, n29308, n29309, n29310, n29311, n29312, n29313, n29314,
         n29315, n29316, n29317, n29318, n29319, n29320, n29321, n29322,
         n29323, n29324, n29325, n29326, n29327, n29328, n29329, n29330,
         n29331, n29332, n29333, n29334, n29335, n29336, n29337, n29338,
         n29339, n29340, n29341, n29342, n29343, n29344, n29345, n29346,
         n29347, n29348, n29349, n29350, n29351, n29352, n29353, n29354,
         n29355, n29356, n29357, n29358, n29359, n29360, n29361, n29362,
         n29363, n29364, n29365, n29366, n29367, n29368, n29369, n29370,
         n29371, n29372, n29373, n29374, n29375, n29376, n29377, n29378,
         n29379, n29380, n29381, n29382, n29383, n29384, n29385, n29386,
         n29387, n29388, n29389, n29390, n29391, n29392, n29393, n29394,
         n29395, n29396, n29397, n29398, n29399, n29400, n29401, n29402,
         n29403, n29404, n29405, n29406, n29407, n29408, n29409, n29410,
         n29411, n29412, n29413, n29414, n29415, n29416, n29417, n29418,
         n29419, n29420, n29421, n29422, n29423, n29424, n29425, n29426,
         n29427, n29428, n29429, n29430, n29431, n29432, n29433, n29434,
         n29435, n29436, n29437, n29438, n29439, n29440, n29441, n29442,
         n29443, n29444, n29445, n29446, n29447, n29448, n29449, n29450,
         n29451, n29452, n29453, n29454, n29455, n29456, n29457, n29458,
         n29459, n29460, n29461, n29462, n29463, n29464, n29465, n29466,
         n29467, n29468, n29469, n29470, n29471, n29472, n29473, n29474,
         n29475, n29476, n29477, n29478, n29479, n29480, n29481, n29482,
         n29483, n29484, n29485, n29486, n29487, n29488, n29489, n29490,
         n29491, n29492, n29493, n29494, n29495, n29496, n29497, n29498,
         n29499, n29500, n29501, n29502, n29503, n29504, n29505, n29506,
         n29507, n29508, n29509, n29510, n29511, n29512, n29513, n29514,
         n29515, n29516, n29517, n29518, n29519, n29520, n29521, n29522,
         n29523, n29524, n29525, n29526, n29527, n29528, n29529, n29530,
         n29531, n29532, n29533, n29534, n29535, n29536, n29537, n29538,
         n29539, n29540, n29541, n29542, n29543, n29544, n29545, n29546,
         n29547, n29548, n29549, n29550, n29551, n29552, n29553, n29554,
         n29555, n29556, n29557, n29558, n29559, n29560, n29561, n29562,
         n29563, n29564, n29565, n29566, n29567, n29568, n29569, n29570,
         n29571, n29572, n29573, n29574, n29575, n29576, n29577, n29578,
         n29579, n29580, n29581, n29582, n29583, n29584, n29585, n29586,
         n29587, n29588, n29589, n29590, n29591, n29592, n29593, n29594,
         n29595, n29596, n29597, n29598, n29599, n29600, n29601, n29602,
         n29603, n29604, n29605, n29606, n29607, n29608, n29609, n29610,
         n29611, n29612, n29613, n29614, n29615, n29616, n29617, n29618,
         n29619, n29620, n29621, n29622, n29623, n29624, n29625, n29626,
         n29627, n29628, n29629, n29630, n29631, n29632, n29633, n29634,
         n29635, n29636, n29637, n29638, n29639, n29640, n29641, n29642,
         n29643, n29644, n29645, n29646, n29647, n29648, n29649, n29650,
         n29651, n29652, n29653, n29654, n29655, n29656, n29657, n29658,
         n29659, n29660, n29661, n29662, n29663, n29664, n29665, n29666,
         n29667, n29668, n29669, n29670, n29671, n29672, n29673, n29674,
         n29675, n29676, n29677, n29678, n29679, n29680, n29681, n29682,
         n29683, n29684, n29685, n29686, n29687, n29688, n29689, n29690,
         n29691, n29692, n29693, n29694, n29695, n29696, n29697, n29698,
         n29699, n29700, n29701, n29702, n29703, n29704, n29705, n29706,
         n29707, n29708, n29709, n29710, n29711, n29712, n29713, n29714,
         n29715, n29716, n29717, n29718, n29719, n29720, n29721, n29722,
         n29723, n29724, n29725, n29726, n29727, n29728, n29729, n29730,
         n29731, n29732, n29733, n29734, n29735, n29736, n29737, n29738,
         n29739, n29740, n29741, n29742, n29743, n29744, n29745, n29746,
         n29747, n29748, n29749, n29750, n29751, n29752, n29753, n29754,
         n29755, n29756, n29757, n29758, n29759, n29760, n29761, n29762,
         n29763, n29764, n29765, n29766, n29767, n29768, n29769, n29770,
         n29771, n29772, n29773, n29774, n29775, n29776, n29777, n29778,
         n29779, n29780, n29781, n29782, n29783, n29784, n29785, n29786,
         n29787, n29788, n29789, n29790, n29791, n29792, n29793, n29794,
         n29795, n29796, n29797, n29798, n29799, n29800, n29801, n29802,
         n29803, n29804, n29805, n29806, n29807, n29808, n29809, n29810,
         n29811, n29812, n29813, n29814, n29815, n29816, n29817, n29818,
         n29819, n29820, n29821, n29822, n29823, n29824, n29825, n29826,
         n29827, n29828, n29829, n29830, n29831, n29832, n29833, n29834,
         n29835, n29836, n29837, n29838, n29839, n29840, n29841, n29842,
         n29843, n29844, n29845, n29846, n29847, n29848, n29849, n29850,
         n29851, n29852, n29853, n29854, n29855, n29856, n29857, n29858,
         n29859, n29860, n29861, n29862, n29863, n29864, n29865, n29866,
         n29867, n29868, n29869, n29870, n29871, n29872, n29873, n29874,
         n29875, n29876, n29877, n29878, n29879, n29880, n29881, n29882,
         n29883, n29884, n29885, n29886, n29887, n29888, n29889, n29890,
         n29891, n29892, n29893, n29894, n29895, n29896, n29897, n29898,
         n29899, n29900, n29901, n29902, n29903, n29904, n29905, n29906,
         n29907, n29908, n29909, n29910, n29911, n29912, n29913, n29914,
         n29915, n29916, n29917, n29918, n29919, n29920, n29921, n29922,
         n29923, n29924, n29925, n29926, n29927, n29928, n29929, n29930,
         n29931, n29932, n29933, n29934, n29935, n29936, n29937, n29938,
         n29939, n29940, n29941, n29942, n29943, n29944, n29945, n29946,
         n29947, n29948, n29949, n29950, n29951, n29952, n29953, n29954,
         n29955, n29956, n29957, n29958, n29959, n29960, n29961, n29962,
         n29963, n29964, n29965, n29966, n29967, n29968, n29969, n29970,
         n29971, n29972, n29973, n29974, n29975, n29976, n29977, n29978,
         n29979, n29980, n29981, n29982, n29983, n29984, n29985, n29986,
         n29987, n29988, n29989, n29990, n29991, n29992, n29993, n29994,
         n29995, n29996, n29997, n29998, n29999, n30000, n30001, n30002,
         n30003, n30004, n30005, n30006, n30007, n30008, n30009, n30010,
         n30011, n30012, n30013, n30014, n30015, n30016, n30017, n30018,
         n30019, n30020, n30021, n30022, n30023, n30024, n30025, n30026,
         n30027, n30028, n30029, n30030, n30031, n30032, n30033, n30034,
         n30035, n30036, n30037, n30038, n30039, n30040, n30041, n30042,
         n30043, n30044, n30045, n30046, n30047, n30048, n30049, n30050,
         n30051, n30052, n30053, n30054, n30055, n30056, n30057, n30058,
         n30059, n30060, n30061, n30062, n30063, n30064, n30065, n30066,
         n30067, n30068, n30069, n30070, n30071, n30072, n30073, n30074,
         n30075, n30076, n30077, n30078, n30079, n30080, n30081, n30082,
         n30083, n30084, n30085, n30086, n30087, n30088, n30089, n30090,
         n30091, n30092, n30093, n30094, n30095, n30096, n30097, n30098,
         n30099, n30100, n30101, n30102, n30103, n30104, n30105, n30106,
         n30107, n30108, n30109, n30110, n30111, n30112, n30113, n30114,
         n30115, n30116, n30117, n30118, n30119, n30120, n30121, n30122,
         n30123, n30124, n30125, n30126, n30127, n30128, n30129, n30130,
         n30131, n30132, n30133, n30134, n30135, n30136, n30137, n30138,
         n30139, n30140, n30141, n30142, n30143, n30144, n30145, n30146,
         n30147, n30148, n30149, n30150, n30151, n30152, n30153, n30154,
         n30155, n30156, n30157, n30158, n30159, n30160, n30161, n30162,
         n30163, n30164, n30165, n30166, n30167, n30168, n30169, n30170,
         n30171, n30172, n30173, n30174, n30175, n30176, n30177, n30178,
         n30179, n30180, n30181, n30182, n30183, n30184, n30185, n30186,
         n30187, n30188, n30189, n30190, n30191, n30192, n30193, n30194,
         n30195, n30196, n30197, n30198, n30199, n30200, n30201, n30202,
         n30203, n30204, n30205, n30206, n30207, n30208, n30209, n30210,
         n30211, n30212, n30213, n30214, n30215, n30216, n30217, n30218,
         n30219, n30220, n30221, n30222, n30223, n30224, n30225, n30226,
         n30227, n30228, n30229, n30230, n30231, n30232, n30233, n30234,
         n30235, n30236, n30237, n30238, n30239, n30240, n30241, n30242,
         n30243, n30244, n30245, n30246, n30247, n30248, n30249, n30250,
         n30251, n30252, n30253, n30254, n30255, n30256, n30257, n30258,
         n30259, n30260, n30261, n30262, n30263, n30264, n30265, n30266,
         n30267, n30268, n30269, n30270, n30271, n30272, n30273, n30274,
         n30275, n30276, n30277, n30278, n30279, n30280, n30281, n30282,
         n30283, n30284, n30285, n30286, n30287, n30288, n30289, n30290,
         n30291, n30292, n30293, n30294, n30295, n30296, n30297, n30298,
         n30299, n30300, n30301, n30302, n30303, n30304, n30305, n30306,
         n30307, n30308, n30309, n30310, n30311, n30312, n30313, n30314,
         n30315, n30316, n30317, n30318, n30319, n30320, n30321, n30322,
         n30323, n30324, n30325, n30326, n30327, n30328, n30329, n30330,
         n30331, n30332, n30333, n30334, n30335, n30336, n30337, n30338,
         n30339, n30340, n30341, n30342, n30343, n30344, n30345, n30346,
         n30347, n30348, n30349, n30350, n30351, n30352, n30353, n30354,
         n30355, n30356, n30357, n30358, n30359, n30360, n30361, n30362,
         n30363, n30364, n30365, n30366, n30367, n30368, n30369, n30370,
         n30371, n30372, n30373, n30374, n30375, n30376, n30377, n30378,
         n30379, n30380, n30381, n30382, n30383, n30384, n30385, n30386,
         n30387, n30388, n30389, n30390, n30391, n30392, n30393, n30394,
         n30395, n30396, n30397, n30398, n30399, n30400, n30401, n30402,
         n30403, n30404, n30405, n30406, n30407, n30408, n30409, n30410,
         n30411, n30412, n30413, n30414, n30415, n30416, n30417, n30418,
         n30419, n30420, n30421, n30422, n30423, n30424, n30425, n30426,
         n30427, n30428, n30429, n30430, n30431, n30432, n30433, n30434,
         n30435, n30436, n30437, n30438, n30439, n30440, n30441, n30442,
         n30443, n30444, n30445, n30446, n30447, n30448, n30449, n30450,
         n30451, n30452, n30453, n30454, n30455, n30456, n30457, n30458,
         n30459, n30460, n30461, n30462, n30463, n30464, n30465, n30466,
         n30467, n30468, n30469, n30470, n30471, n30472, n30473, n30474,
         n30475, n30476, n30477, n30478, n30479, n30480, n30481, n30482,
         n30483, n30484, n30485, n30486, n30487, n30488, n30489, n30490,
         n30491, n30492, n30493, n30494, n30495, n30496, n30497, n30498,
         n30499, n30500, n30501, n30502, n30503, n30504, n30505, n30506,
         n30507, n30508, n30509, n30510, n30511, n30512, n30513, n30514,
         n30515, n30516, n30517, n30518, n30519, n30520, n30521, n30522,
         n30523, n30524, n30525, n30526, n30527, n30528, n30529, n30530,
         n30531, n30532, n30533, n30534, n30535, n30536, n30537, n30538,
         n30539, n30540, n30541, n30542, n30543, n30544, n30545, n30546,
         n30547, n30548, n30549, n30550, n30551, n30552, n30553, n30554,
         n30555, n30556, n30557, n30558, n30559, n30560, n30561, n30562,
         n30563, n30564, n30565, n30566, n30567, n30568, n30569, n30570,
         n30571, n30572, n30573, n30574, n30575, n30576, n30577, n30578,
         n30579, n30580, n30581, n30582, n30583, n30584, n30585, n30586,
         n30587, n30588, n30589, n30590, n30591, n30592, n30593, n30594,
         n30595, n30596, n30597, n30598, n30599, n30600, n30601, n30602,
         n30603, n30604, n30605, n30606, n30607, n30608, n30609, n30610,
         n30611, n30612, n30613, n30614, n30615, n30616, n30617, n30618,
         n30619, n30620, n30621, n30622, n30623, n30624, n30625, n30626,
         n30627, n30628, n30629, n30630, n30631, n30632, n30633, n30634,
         n30635, n30636, n30637, n30638, n30639, n30640, n30641, n30642,
         n30643, n30644, n30645, n30646, n30647, n30648, n30649, n30650,
         n30651, n30652, n30653, n30654, n30655, n30656, n30657, n30658,
         n30659, n30660, n30661, n30662, n30663, n30664, n30665, n30666,
         n30667, n30668, n30669, n30670, n30671, n30672, n30673, n30674,
         n30675, n30676, n30677, n30678, n30679, n30680, n30681, n30682,
         n30683, n30684, n30685, n30686, n30687, n30688, n30689, n30690,
         n30691, n30692, n30693, n30694, n30695, n30696, n30697, n30698,
         n30699, n30700, n30701, n30702, n30703, n30704, n30705, n30706,
         n30707, n30708, n30709, n30710, n30711, n30712, n30713, n30714,
         n30715, n30716, n30717, n30718, n30719, n30720, n30721, n30722,
         n30723, n30724, n30725, n30726, n30727, n30728, n30729, n30730,
         n30731, n30732, n30733, n30734, n30735, n30736, n30737, n30738,
         n30739, n30740, n30741, n30742, n30743, n30744, n30745, n30746,
         n30747, n30748, n30749, n30750, n30751, n30752, n30753, n30754,
         n30755, n30756, n30757, n30758, n30759, n30760, n30761, n30762,
         n30763, n30764, n30765, n30766, n30767, n30768, n30769, n30770,
         n30771, n30772, n30773, n30774, n30775, n30776, n30777, n30778,
         n30779, n30780, n30781, n30782, n30783, n30784, n30785, n30786,
         n30787, n30788, n30789, n30790, n30791, n30792, n30793, n30794,
         n30795, n30796, n30797, n30798, n30799, n30800, n30801, n30802,
         n30803, n30804, n30805, n30806, n30807, n30808, n30809, n30810,
         n30811, n30812, n30813, n30814, n30815, n30816, n30817, n30818,
         n30819, n30820, n30821, n30822, n30823, n30824, n30825, n30826,
         n30827, n30828, n30829, n30830, n30831, n30832, n30833, n30834,
         n30835, n30836, n30837, n30838, n30839, n30840, n30841, n30842,
         n30843, n30844, n30845, n30846, n30847, n30848, n30849, n30850,
         n30851, n30852, n30853, n30854, n30855, n30856, n30857, n30858,
         n30859, n30860, n30861, n30862, n30863, n30864, n30865, n30866,
         n30867, n30868, n30869, n30870, n30871, n30872, n30873, n30874,
         n30875, n30876, n30877, n30878, n30879, n30880, n30881, n30882,
         n30883, n30884, n30885, n30886, n30887, n30888, n30889, n30890,
         n30891, n30892, n30893, n30894, n30895, n30896, n30897, n30898,
         n30899, n30900, n30901, n30902, n30903, n30904, n30905, n30906,
         n30907, n30908, n30909, n30910, n30911, n30912, n30913, n30914,
         n30915, n30916, n30917, n30918, n30919, n30920, n30921, n30922,
         n30923, n30924, n30925, n30926, n30927, n30928, n30929, n30930,
         n30931, n30932, n30933, n30934, n30935, n30936, n30937, n30938,
         n30939, n30940, n30941, n30942, n30943, n30944, n30945, n30946,
         n30947, n30948, n30949, n30950, n30951, n30952, n30953, n30954,
         n30955, n30956, n30957, n30958, n30959, n30960, n30961, n30962,
         n30963, n30964, n30965, n30966, n30967, n30968, n30969, n30970,
         n30971, n30972, n30973, n30974, n30975, n30976, n30977, n30978,
         n30979, n30980, n30981, n30982, n30983, n30984, n30985, n30986,
         n30987, n30988, n30989, n30990, n30991, n30992, n30993, n30994,
         n30995, n30996, n30997, n30998, n30999, n31000, n31001, n31002,
         n31003, n31004, n31005, n31006, n31007, n31008, n31009, n31010,
         n31011, n31012, n31013, n31014, n31015, n31016, n31017, n31018,
         n31019, n31020, n31021, n31022, n31023, n31024, n31025, n31026,
         n31027, n31028, n31029, n31030, n31031, n31032, n31033, n31034,
         n31035, n31036, n31037, n31038, n31039, n31040, n31041, n31042,
         n31043, n31044, n31045, n31046, n31047, n31048, n31049, n31050,
         n31051, n31052, n31053, n31054, n31055, n31056, n31057, n31058,
         n31059, n31060, n31061, n31062, n31063, n31064, n31065, n31066,
         n31067, n31068, n31069, n31070, n31071, n31072, n31073, n31074,
         n31075, n31076, n31077, n31078, n31079, n31080, n31081, n31082,
         n31083, n31084, n31085, n31086, n31087, n31088, n31089, n31090,
         n31091, n31092, n31093, n31094, n31095, n31096, n31097, n31098,
         n31099, n31100, n31101, n31102, n31103, n31104, n31105, n31106,
         n31107, n31108, n31109, n31110, n31111, n31112, n31113, n31114,
         n31115, n31116, n31117, n31118, n31119, n31120, n31121, n31122,
         n31123, n31124, n31125, n31126, n31127, n31128, n31129, n31130,
         n31131, n31132, n31133, n31134, n31135, n31136, n31137, n31138,
         n31139, n31140, n31141, n31142, n31143, n31144, n31145, n31146,
         n31147, n31148, n31149, n31150, n31151, n31152, n31153, n31154,
         n31155, n31156, n31157, n31158, n31159, n31160, n31161, n31162,
         n31163, n31164, n31165, n31166, n31167, n31168, n31169, n31170,
         n31171, n31172, n31173, n31174, n31175, n31176, n31177, n31178,
         n31179, n31180, n31181, n31182, n31183, n31184, n31185, n31186,
         n31187, n31188, n31189, n31190, n31191, n31192, n31193, n31194,
         n31195, n31196, n31197, n31198, n31199, n31200, n31201, n31202,
         n31203, n31204, n31205, n31206, n31207, n31208, n31209, n31210,
         n31211, n31212, n31213, n31214, n31215, n31216, n31217, n31218,
         n31219, n31220, n31221, n31222, n31223, n31224, n31225, n31226,
         n31227, n31228, n31229, n31230, n31231, n31232, n31233, n31234,
         n31235, n31236, n31237, n31238, n31239, n31240, n31241, n31242,
         n31243, n31244, n31245, n31246, n31247, n31248, n31249, n31250,
         n31251, n31252, n31253, n31254, n31255, n31256, n31257, n31258,
         n31259, n31260, n31261, n31262, n31263, n31264, n31265, n31266,
         n31267, n31268, n31269, n31270, n31271, n31272, n31273, n31274,
         n31275, n31276, n31277, n31278, n31279, n31280, n31281, n31282,
         n31283, n31284, n31285, n31286, n31287, n31288, n31289, n31290,
         n31291, n31292, n31293, n31294, n31295, n31296, n31297, n31298,
         n31299, n31300, n31301, n31302, n31303, n31304, n31305, n31306,
         n31307, n31308, n31309, n31310, n31311, n31312, n31313, n31314,
         n31315, n31316, n31317, n31318, n31319, n31320, n31321, n31322,
         n31323, n31324, n31325, n31326, n31327, n31328, n31329, n31330,
         n31331, n31332, n31333, n31334, n31335, n31336, n31337, n31338,
         n31339, n31340, n31341, n31342, n31343, n31344, n31345, n31346,
         n31347, n31348, n31349, n31350, n31351, n31352, n31353, n31354,
         n31355, n31356, n31357, n31358, n31359, n31360, n31361, n31362,
         n31363, n31364, n31365, n31366, n31367, n31368, n31369, n31370,
         n31371, n31372, n31373, n31374, n31375, n31376, n31377, n31378,
         n31379, n31380, n31381, n31382, n31383, n31384, n31385, n31386,
         n31387, n31388, n31389, n31390, n31391, n31392, n31393, n31394,
         n31395, n31396, n31397, n31398, n31399, n31400, n31401, n31402,
         n31403, n31404, n31405, n31406, n31407, n31408, n31409, n31410,
         n31411, n31412, n31413, n31414, n31415, n31416, n31417, n31418,
         n31419, n31420, n31421, n31422, n31423, n31424, n31425, n31426,
         n31427, n31428, n31429, n31430, n31431, n31432, n31433, n31434,
         n31435, n31436, n31437, n31438, n31439, n31440, n31441, n31442,
         n31443, n31444, n31445, n31446, n31447, n31448, n31449, n31450,
         n31451, n31452, n31453, n31454, n31455, n31456, n31457, n31458,
         n31459, n31460, n31461, n31462, n31463, n31464, n31465, n31466,
         n31467, n31468, n31469, n31470, n31471, n31472, n31473, n31474,
         n31475, n31476, n31477, n31478, n31479, n31480, n31481, n31482,
         n31483, n31484, n31485, n31486, n31487, n31488, n31489, n31490,
         n31491, n31492, n31493, n31494, n31495, n31496, n31497, n31498,
         n31499, n31500, n31501, n31502, n31503, n31504, n31505, n31506,
         n31507, n31508, n31509, n31510, n31511, n31512, n31513, n31514,
         n31515, n31516, n31517, n31518, n31519, n31520, n31521, n31522,
         n31523, n31524, n31525, n31526, n31527, n31528, n31529, n31530,
         n31531, n31532, n31533, n31534, n31535, n31536, n31537, n31538,
         n31539, n31540, n31541, n31542, n31543, n31544, n31545, n31546,
         n31547, n31548, n31549, n31550, n31551, n31552, n31553, n31554,
         n31555, n31556, n31557, n31558, n31559, n31560, n31561, n31562,
         n31563, n31564, n31565, n31566, n31567, n31568, n31569, n31570,
         n31571, n31572, n31573, n31574, n31575, n31576, n31577, n31578,
         n31579, n31580, n31581, n31582, n31583, n31584, n31585, n31586,
         n31587, n31588, n31589, n31590, n31591, n31592, n31593, n31594,
         n31595, n31596, n31597, n31598, n31599, n31600, n31601, n31602,
         n31603, n31604, n31605, n31606, n31607, n31608, n31609, n31610,
         n31611, n31612, n31613, n31614, n31615, n31616, n31617, n31618,
         n31619, n31620, n31621, n31622, n31623, n31624, n31625, n31626,
         n31627, n31628, n31629, n31630, n31631, n31632, n31633, n31634,
         n31635, n31636, n31637, n31638, n31639, n31640, n31641, n31642,
         n31643, n31644, n31645, n31646, n31647, n31648, n31649, n31650,
         n31651, n31652, n31653, n31654, n31655, n31656, n31657, n31658,
         n31659, n31660, n31661, n31662, n31663, n31664, n31665, n31666,
         n31667, n31668, n31669, n31670, n31671, n31672, n31673, n31674,
         n31675, n31676, n31677, n31678, n31679, n31680, n31681, n31682,
         n31683, n31684, n31685, n31686, n31687, n31688, n31689, n31690,
         n31691, n31692, n31693, n31694, n31695, n31696, n31697, n31698,
         n31699, n31700, n31701, n31702, n31703, n31704, n31705, n31706,
         n31707, n31708, n31709, n31710, n31711, n31712, n31713, n31714,
         n31715, n31716, n31717, n31718, n31719, n31720, n31721, n31722,
         n31723, n31724, n31725, n31726, n31727, n31728, n31729, n31730,
         n31731, n31732, n31733, n31734, n31735, n31736, n31737, n31738,
         n31739, n31740, n31741, n31742, n31743, n31744, n31745, n31746,
         n31747, n31748, n31749, n31750, n31751, n31752, n31753, n31754,
         n31755, n31756, n31757, n31758, n31759, n31760, n31761, n31762,
         n31763, n31764, n31765, n31766, n31767, n31768, n31769, n31770,
         n31771, n31772, n31773, n31774, n31775, n31776, n31777, n31778,
         n31779, n31780, n31781, n31782, n31783, n31784, n31785, n31786,
         n31787, n31788, n31789, n31790, n31791, n31792, n31793, n31794,
         n31795, n31796, n31797, n31798, n31799, n31800, n31801, n31802,
         n31803, n31804, n31805, n31806, n31807, n31808, n31809, n31810,
         n31811, n31812, n31813, n31814, n31815, n31816, n31817, n31818,
         n31819, n31820, n31821, n31822, n31823, n31824, n31825, n31826,
         n31827, n31828, n31829, n31830, n31831, n31832, n31833, n31834,
         n31835, n31836, n31837, n31838, n31839, n31840, n31841, n31842,
         n31843, n31844, n31845, n31846, n31847, n31848, n31849, n31850,
         n31851, n31852, n31853, n31854, n31855, n31856, n31857, n31858,
         n31859, n31860, n31861, n31862, n31863, n31864, n31865, n31866,
         n31867, n31868, n31869, n31870, n31871, n31872, n31873, n31874,
         n31875, n31876, n31877, n31878, n31879, n31880, n31881, n31882,
         n31883, n31884, n31885, n31886, n31887, n31888, n31889, n31890,
         n31891, n31892, n31893, n31894, n31895, n31896, n31897, n31898,
         n31899, n31900, n31901, n31902, n31903, n31904, n31905, n31906,
         n31907, n31908, n31909, n31910, n31911, n31912, n31913, n31914,
         n31915, n31916, n31917, n31918, n31919, n31920, n31921, n31922,
         n31923, n31924, n31925, n31926, n31927, n31928, n31929, n31930,
         n31931, n31932, n31933, n31934, n31935, n31936, n31937, n31938,
         n31939, n31940, n31941, n31942, n31943, n31944, n31945, n31946,
         n31947, n31948, n31949, n31950, n31951, n31952, n31953, n31954,
         n31955, n31956, n31957, n31958, n31959, n31960, n31961, n31962,
         n31963, n31964, n31965, n31966, n31967, n31968, n31969, n31970,
         n31971, n31972, n31973, n31974, n31975, n31976, n31977, n31978,
         n31979, n31980, n31981, n31982, n31983, n31984, n31985, n31986,
         n31987, n31988, n31989, n31990, n31991, n31992, n31993, n31994,
         n31995, n31996, n31997, n31998, n31999, n32000, n32001, n32002,
         n32003, n32004, n32005, n32006, n32007, n32008, n32009, n32010,
         n32011, n32012, n32013, n32014, n32015, n32016, n32017, n32018,
         n32019, n32020, n32021, n32022, n32023, n32024, n32025, n32026,
         n32027, n32028, n32029, n32030, n32031, n32032, n32033, n32034,
         n32035, n32036, n32037, n32038, n32039, n32040, n32041, n32042,
         n32043, n32044, n32045, n32046, n32047, n32048, n32049, n32050,
         n32051, n32052, n32053, n32054, n32055, n32056, n32057, n32058,
         n32059, n32060, n32061, n32062, n32063, n32064, n32065, n32066,
         n32067, n32068, n32069, n32070, n32071, n32072, n32073, n32074,
         n32075, n32076, n32077, n32078, n32079, n32080, n32081, n32082,
         n32083, n32084, n32085, n32086, n32087, n32088, n32089, n32090,
         n32091, n32092, n32093, n32094, n32095, n32096, n32097, n32098,
         n32099, n32100, n32101, n32102, n32103, n32104, n32105, n32106,
         n32107, n32108, n32109, n32110, n32111, n32112, n32113, n32114,
         n32115, n32116, n32117, n32118, n32119, n32120, n32121, n32122,
         n32123, n32124, n32125, n32126, n32127, n32128, n32129, n32130,
         n32131, n32132, n32133, n32134, n32135, n32136, n32137, n32138,
         n32139, n32140, n32141, n32142, n32143, n32144, n32145, n32146,
         n32147, n32148, n32149, n32150, n32151, n32152, n32153, n32154,
         n32155, n32156, n32157, n32158, n32159, n32160, n32161, n32162,
         n32163, n32164, n32165, n32166, n32167, n32168, n32169, n32170,
         n32171, n32172, n32173, n32174, n32175, n32176, n32177, n32178,
         n32179, n32180, n32181, n32182, n32183, n32184, n32185, n32186,
         n32187, n32188, n32189, n32190, n32191, n32192, n32193, n32194,
         n32195, n32196, n32197, n32198, n32199, n32200, n32201, n32202,
         n32203, n32204, n32205, n32206, n32207, n32208, n32209, n32210,
         n32211, n32212, n32213, n32214, n32215, n32216, n32217, n32218,
         n32219, n32220, n32221, n32222, n32223, n32224, n32225, n32226,
         n32227, n32228, n32229, n32230, n32231, n32232, n32233, n32234,
         n32235, n32236, n32237, n32238, n32239, n32240, n32241, n32242,
         n32243, n32244, n32245, n32246, n32247, n32248, n32249, n32250,
         n32251, n32252, n32253, n32254, n32255, n32256, n32257, n32258,
         n32259, n32260, n32261, n32262, n32263, n32264, n32265, n32266,
         n32267, n32268, n32269, n32270, n32271, n32272, n32273, n32274,
         n32275, n32276, n32277, n32278, n32279, n32280, n32281, n32282,
         n32283, n32284, n32285, n32286, n32287, n32288, n32289, n32290,
         n32291, n32292, n32293, n32294, n32295, n32296, n32297, n32298,
         n32299, n32300, n32301, n32302, n32303, n32304, n32305, n32306,
         n32307, n32308, n32309, n32310, n32311, n32312, n32313, n32314,
         n32315, n32316, n32317, n32318, n32319, n32320, n32321, n32322,
         n32323, n32324, n32325, n32326, n32327, n32328, n32329, n32330,
         n32331, n32332, n32333, n32334, n32335, n32336, n32337, n32338,
         n32339, n32340, n32341, n32342, n32343, n32344, n32345, n32346,
         n32347, n32348, n32349, n32350, n32351, n32352, n32353, n32354,
         n32355, n32356, n32357, n32358, n32359, n32360, n32361, n32362,
         n32363, n32364, n32365, n32366, n32367, n32368, n32369, n32370,
         n32371, n32372, n32373, n32374, n32375, n32376, n32377, n32378,
         n32379, n32380, n32381, n32382, n32383, n32384, n32385, n32386,
         n32387, n32388, n32389, n32390, n32391, n32392, n32393, n32394,
         n32395, n32396, n32397, n32398, n32399, n32400, n32401, n32402,
         n32403, n32404, n32405, n32406, n32407, n32408, n32409, n32410,
         n32411, n32412, n32413, n32414, n32415, n32416, n32417, n32418,
         n32419, n32420, n32421, n32422, n32423, n32424, n32425, n32426,
         n32427, n32428, n32429, n32430, n32431, n32432, n32433, n32434,
         n32435, n32436, n32437, n32438, n32439, n32440, n32441, n32442,
         n32443, n32444, n32445, n32446, n32447, n32448, n32449, n32450,
         n32451, n32452, n32453, n32454, n32455, n32456, n32457, n32458,
         n32459, n32460, n32461, n32462, n32463, n32464, n32465, n32466,
         n32467, n32468, n32469, n32470, n32471, n32472, n32473, n32474,
         n32475, n32476, n32477, n32478, n32479, n32480, n32481, n32482,
         n32483, n32484, n32485, n32486, n32487, n32488, n32489, n32490,
         n32491, n32492, n32493, n32494, n32495, n32496, n32497, n32498,
         n32499, n32500, n32501, n32502, n32503, n32504, n32505, n32506,
         n32507, n32508, n32509, n32510, n32511, n32512, n32513, n32514,
         n32515, n32516, n32517, n32518, n32519, n32520, n32521, n32522,
         n32523, n32524, n32525, n32526, n32527, n32528, n32529, n32530,
         n32531, n32532, n32533, n32534, n32535, n32536, n32537, n32538,
         n32539, n32540, n32541, n32542, n32543, n32544, n32545, n32546,
         n32547, n32548, n32549, n32550, n32551, n32552, n32553, n32554,
         n32555, n32556, n32557, n32558, n32559, n32560, n32561, n32562,
         n32563, n32564, n32565, n32566, n32567, n32568, n32569, n32570,
         n32571, n32572, n32573, n32574, n32575, n32576, n32577, n32578,
         n32579, n32580, n32581, n32582, n32583, n32584, n32585, n32586,
         n32587, n32588, n32589, n32590, n32591, n32592, n32593, n32594,
         n32595, n32596, n32597, n32598, n32599, n32600, n32601, n32602,
         n32603, n32604, n32605, n32606, n32607, n32608, n32609, n32610,
         n32611, n32612, n32613, n32614, n32615, n32616, n32617, n32618,
         n32619, n32620, n32621, n32622, n32623, n32624, n32625, n32626,
         n32627, n32628, n32629, n32630, n32631, n32632, n32633, n32634,
         n32635, n32636, n32637, n32638, n32639, n32640, n32641, n32642,
         n32643, n32644, n32645, n32646, n32647, n32648, n32649, n32650,
         n32651, n32652, n32653, n32654, n32655, n32656, n32657, n32658,
         n32659, n32660, n32661, n32662, n32663, n32664, n32665, n32666,
         n32667, n32668, n32669, n32670, n32671, n32672, n32673, n32674,
         n32675, n32676, n32677, n32678, n32679, n32680, n32681, n32682,
         n32683, n32684, n32685, n32686, n32687, n32688, n32689, n32690,
         n32691, n32692, n32693, n32694, n32695, n32696, n32697, n32698,
         n32699, n32700, n32701, n32702, n32703, n32704, n32705, n32706,
         n32707, n32708, n32709, n32710, n32711, n32712, n32713, n32714,
         n32715, n32716, n32717, n32718, n32719, n32720, n32721, n32722,
         n32723, n32724, n32725, n32726, n32727, n32728, n32729, n32730,
         n32731, n32732, n32733, n32734, n32735, n32736, n32737, n32738,
         n32739, n32740, n32741, n32742, n32743, n32744, n32745, n32746,
         n32747, n32748, n32749, n32750, n32751, n32752, n32753, n32754,
         n32755, n32756, n32757, n32758, n32759, n32760, n32761, n32762,
         n32763, n32764, n32765, n32766, n32767, n32768, n32769, n32770,
         n32771, n32772, n32773, n32774, n32775, n32776, n32777, n32778,
         n32779, n32780, n32781, n32782, n32783, n32784, n32785, n32786,
         n32787, n32788, n32789, n32790, n32791, n32792, n32793, n32794,
         n32795, n32796, n32797, n32798, n32799, n32800, n32801, n32802,
         n32803, n32804, n32805, n32806, n32807, n32808, n32809, n32810,
         n32811, n32812, n32813, n32814, n32815, n32816, n32817, n32818,
         n32819, n32820, n32821, n32822, n32823, n32824, n32825, n32826,
         n32827, n32828, n32829, n32830, n32831, n32832, n32833, n32834,
         n32835, n32836, n32837, n32838, n32839, n32840, n32841, n32842,
         n32843, n32844, n32845, n32846, n32847, n32848, n32849, n32850,
         n32851, n32852, n32853, n32854, n32855, n32856, n32857, n32858,
         n32859, n32860, n32861, n32862, n32863, n32864, n32865, n32866,
         n32867, n32868, n32869, n32870, n32871, n32872, n32873, n32874,
         n32875, n32876, n32877, n32878, n32879, n32880, n32881, n32882,
         n32883, n32884, n32885, n32886, n32887, n32888, n32889, n32890,
         n32891, n32892, n32893, n32894, n32895, n32896, n32897, n32898,
         n32899, n32900, n32901, n32902, n32903, n32904, n32905, n32906,
         n32907, n32908, n32909, n32910, n32911, n32912, n32913, n32914,
         n32915, n32916, n32917, n32918, n32919, n32920, n32921, n32922,
         n32923, n32924, n32925, n32926, n32927, n32928, n32929, n32930,
         n32931, n32932, n32933, n32934, n32935, n32936, n32937, n32938,
         n32939, n32940, n32941, n32942, n32943, n32944, n32945, n32946,
         n32947, n32948, n32949, n32950, n32951, n32952, n32953, n32954,
         n32955, n32956, n32957, n32958, n32959, n32960, n32961, n32962,
         n32963, n32964, n32965, n32966, n32967, n32968, n32969, n32970,
         n32971, n32972, n32973, n32974, n32975, n32976, n32977, n32978,
         n32979, n32980, n32981, n32982, n32983, n32984, n32985, n32986,
         n32987, n32988, n32989, n32990, n32991, n32992, n32993, n32994,
         n32995, n32996, n32997, n32998, n32999, n33000, n33001, n33002,
         n33003, n33004, n33005, n33006, n33007, n33008, n33009, n33010,
         n33011, n33012, n33013, n33014, n33015, n33016, n33017, n33018,
         n33019, n33020, n33021, n33022, n33023, n33024, n33025, n33026,
         n33027, n33028, n33029, n33030, n33031, n33032, n33033, n33034,
         n33035, n33036, n33037, n33038, n33039, n33040, n33041, n33042,
         n33043, n33044, n33045, n33046, n33047, n33048, n33049, n33050,
         n33051, n33052, n33053, n33054, n33055, n33056, n33057, n33058,
         n33059, n33060, n33061, n33062, n33063, n33064, n33065, n33066,
         n33067, n33068, n33069, n33070, n33071, n33072, n33073, n33074,
         n33075, n33076, n33077, n33078, n33079, n33080, n33081, n33082,
         n33083, n33084, n33085, n33086, n33087, n33088, n33089, n33090,
         n33091, n33092, n33093, n33094, n33095, n33096, n33097, n33098,
         n33099, n33100, n33101, n33102, n33103, n33104, n33105, n33106,
         n33107, n33108, n33109, n33110, n33111, n33112, n33113, n33114,
         n33115, n33116, n33117, n33118, n33119, n33120, n33121, n33122,
         n33123, n33124, n33125, n33126, n33127, n33128, n33129, n33130,
         n33131, n33132, n33133, n33134, n33135, n33136, n33137, n33138,
         n33139, n33140, n33141, n33142, n33143, n33144, n33145, n33146,
         n33147, n33148, n33149, n33150, n33151, n33152, n33153, n33154,
         n33155, n33156, n33157, n33158, n33159, n33160, n33161, n33162,
         n33163, n33164, n33165, n33166, n33167, n33168, n33169, n33170,
         n33171, n33172, n33173, n33174, n33175, n33176, n33177, n33178,
         n33179, n33180, n33181, n33182, n33183, n33184, n33185, n33186,
         n33187, n33188, n33189, n33190, n33191, n33192, n33193, n33194,
         n33195, n33196, n33197, n33198, n33199, n33200, n33201, n33202,
         n33203, n33204, n33205, n33206, n33207, n33208, n33209, n33210,
         n33211, n33212, n33213, n33214, n33215, n33216, n33217, n33218,
         n33219, n33220, n33221, n33222, n33223, n33224, n33225, n33226,
         n33227, n33228, n33229, n33230, n33231, n33232, n33233, n33234,
         n33235, n33236, n33237, n33238, n33239, n33240, n33241, n33242,
         n33243, n33244, n33245, n33246, n33247, n33248, n33249, n33250,
         n33251, n33252, n33253, n33254, n33255, n33256, n33257, n33258,
         n33259, n33260, n33261, n33262, n33263, n33264, n33265, n33266,
         n33267, n33268, n33269, n33270, n33271, n33272, n33273, n33274,
         n33275, n33276, n33277, n33278, n33279, n33280, n33281, n33282,
         n33283, n33284, n33285, n33286, n33287, n33288, n33289, n33290,
         n33291, n33292, n33293, n33294, n33295, n33296, n33297, n33298,
         n33299, n33300, n33301, n33302, n33303, n33304, n33305, n33306,
         n33307, n33308, n33309, n33310, n33311, n33312, n33313, n33314,
         n33315, n33316, n33317, n33318, n33319, n33320, n33321, n33322,
         n33323, n33324, n33325, n33326, n33327, n33328, n33329, n33330,
         n33331, n33332, n33333, n33334, n33335, n33336, n33337, n33338,
         n33339, n33340, n33341, n33342, n33343, n33344, n33345, n33346,
         n33347, n33348, n33349, n33350, n33351, n33352, n33353, n33354,
         n33355, n33356, n33357, n33358, n33359, n33360, n33361, n33362,
         n33363, n33364, n33365, n33366, n33367, n33368, n33369, n33370,
         n33371, n33372, n33373, n33374, n33375, n33376, n33377, n33378,
         n33379, n33380, n33381, n33382, n33383, n33384, n33385, n33386,
         n33387, n33388, n33389, n33390, n33391, n33392, n33393, n33394,
         n33395, n33396, n33397, n33398, n33399, n33400, n33401, n33402,
         n33403, n33404, n33405, n33406, n33407, n33408, n33409, n33410,
         n33411, n33412, n33413, n33414, n33415, n33416, n33417, n33418,
         n33419, n33420, n33421, n33422, n33423, n33424, n33425, n33426,
         n33427, n33428, n33429, n33430, n33431, n33432, n33433, n33434,
         n33435, n33436, n33437, n33438, n33439, n33440, n33441, n33442,
         n33443, n33444, n33445, n33446, n33447, n33448, n33449, n33450,
         n33451, n33452, n33453, n33454, n33455, n33456, n33457, n33458,
         n33459, n33460, n33461, n33462, n33463, n33464, n33465, n33466,
         n33467, n33468, n33469, n33470, n33471, n33472, n33473, n33474,
         n33475, n33476, n33477, n33478, n33479, n33480, n33481, n33482,
         n33483, n33484, n33485, n33486, n33487, n33488, n33489, n33490,
         n33491, n33492, n33493, n33494, n33495, n33496, n33497, n33498,
         n33499, n33500, n33501, n33502, n33503, n33504, n33505, n33506,
         n33507, n33508, n33509, n33510, n33511, n33512, n33513, n33514,
         n33515, n33516, n33517, n33518, n33519, n33520, n33521, n33522,
         n33523, n33524, n33525, n33526, n33527, n33528, n33529, n33530,
         n33531, n33532, n33533, n33534, n33535, n33536, n33537, n33538,
         n33539, n33540, n33541, n33542, n33543, n33544, n33545, n33546,
         n33547, n33548, n33549, n33550, n33551, n33552, n33553, n33554,
         n33555, n33556, n33557, n33558, n33559, n33560, n33561, n33562,
         n33563, n33564, n33565, n33566, n33567, n33568, n33569, n33570,
         n33571, n33572, n33573, n33574, n33575, n33576, n33577, n33578,
         n33579, n33580, n33581, n33582, n33583, n33584, n33585, n33586,
         n33587, n33588, n33589, n33590, n33591, n33592, n33593, n33594,
         n33595, n33596, n33597, n33598, n33599, n33600, n33601, n33602,
         n33603, n33604, n33605, n33606, n33607, n33608, n33609, n33610,
         n33611, n33612, n33613, n33614, n33615, n33616, n33617, n33618,
         n33619, n33620, n33621, n33622, n33623, n33624, n33625, n33626,
         n33627, n33628, n33629, n33630, n33631, n33632, n33633, n33634,
         n33635, n33636, n33637, n33638, n33639, n33640, n33641, n33642,
         n33643, n33644, n33645, n33646, n33647, n33648, n33649, n33650,
         n33651, n33652, n33653, n33654, n33655, n33656, n33657, n33658,
         n33659, n33660, n33661, n33662, n33663, n33664, n33665, n33666,
         n33667, n33668, n33669, n33670, n33671, n33672, n33673, n33674,
         n33675, n33676, n33677, n33678, n33679, n33680, n33681, n33682,
         n33683, n33684, n33685, n33686, n33687, n33688, n33689, n33690,
         n33691, n33692, n33693, n33694, n33695, n33696, n33697, n33698,
         n33699, n33700, n33701, n33702, n33703, n33704, n33705, n33706,
         n33707, n33708, n33709, n33710, n33711, n33712, n33713, n33714,
         n33715, n33716, n33717, n33718, n33719, n33720, n33721, n33722,
         n33723, n33724, n33725, n33726, n33727, n33728, n33729, n33730,
         n33731, n33732, n33733, n33734, n33735, n33736, n33737, n33738,
         n33739, n33740, n33741, n33742, n33743, n33744, n33745, n33746,
         n33747, n33748, n33749, n33750, n33751, n33752, n33753, n33754,
         n33755, n33756, n33757, n33758, n33759, n33760, n33761, n33762,
         n33763, n33764, n33765, n33766, n33767, n33768, n33769, n33770,
         n33771, n33772, n33773, n33774, n33775, n33776, n33777, n33778,
         n33779, n33780, n33781, n33782, n33783, n33784, n33785, n33786,
         n33787, n33788, n33789, n33790, n33791, n33792, n33793, n33794,
         n33795, n33796, n33797, n33798, n33799, n33800, n33801, n33802,
         n33803, n33804, n33805, n33806, n33807, n33808, n33809, n33810,
         n33811, n33812, n33813, n33814, n33815, n33816, n33817, n33818,
         n33819, n33820, n33821, n33822, n33823, n33824, n33825, n33826,
         n33827, n33828, n33829, n33830, n33831, n33832, n33833, n33834,
         n33835, n33836, n33837, n33838, n33839, n33840, n33841, n33842,
         n33843, n33844, n33845, n33846, n33847, n33848, n33849, n33850,
         n33851, n33852, n33853, n33854, n33855, n33856, n33857, n33858,
         n33859, n33860, n33861, n33862, n33863, n33864, n33865, n33866,
         n33867, n33868, n33869, n33870, n33871, n33872, n33873, n33874,
         n33875, n33876, n33877, n33878, n33879, n33880, n33881, n33882,
         n33883, n33884, n33885, n33886, n33887, n33888, n33889, n33890,
         n33891, n33892, n33893, n33894, n33895, n33896, n33897, n33898,
         n33899, n33900, n33901, n33902, n33903, n33904, n33905, n33906,
         n33907, n33908, n33909, n33910, n33911, n33912, n33913, n33914,
         n33915, n33916, n33917, n33918, n33919, n33920, n33921, n33922,
         n33923, n33924, n33925, n33926, n33927, n33928, n33929, n33930,
         n33931, n33932, n33933, n33934, n33935, n33936, n33937, n33938,
         n33939, n33940, n33941, n33942, n33943, n33944, n33945, n33946,
         n33947, n33948, n33949, n33950, n33951, n33952, n33953, n33954,
         n33955, n33956, n33957, n33958, n33959, n33960, n33961, n33962,
         n33963, n33964, n33965, n33966, n33967, n33968, n33969, n33970,
         n33971, n33972, n33973, n33974, n33975, n33976, n33977, n33978,
         n33979, n33980, n33981, n33982, n33983, n33984, n33985, n33986,
         n33987, n33988, n33989, n33990, n33991, n33992, n33993, n33994,
         n33995, n33996, n33997, n33998, n33999, n34000, n34001, n34002,
         n34003, n34004, n34005, n34006, n34007, n34008, n34009, n34010,
         n34011, n34012, n34013, n34014, n34015, n34016, n34017, n34018,
         n34019, n34020, n34021, n34022, n34023, n34024, n34025, n34026,
         n34027, n34028, n34029, n34030, n34031, n34032, n34033, n34034,
         n34035, n34036, n34037, n34038, n34039, n34040, n34041, n34042,
         n34043, n34044, n34045, n34046, n34047, n34048, n34049, n34050,
         n34051, n34052, n34053, n34054, n34055, n34056, n34057, n34058,
         n34059, n34060, n34061, n34062, n34063, n34064, n34065, n34066,
         n34067, n34068, n34069, n34070, n34071, n34072, n34073, n34074,
         n34075, n34076, n34077, n34078, n34079, n34080, n34081, n34082,
         n34083, n34084, n34085, n34086, n34087, n34088, n34089, n34090,
         n34091, n34092, n34093, n34094, n34095, n34096, n34097, n34098,
         n34099, n34100, n34101, n34102, n34103, n34104, n34105, n34106,
         n34107, n34108, n34109, n34110, n34111, n34112, n34113, n34114,
         n34115, n34116, n34117, n34118, n34119, n34120, n34121, n34122,
         n34123, n34124, n34125, n34126, n34127, n34128, n34129, n34130,
         n34131, n34132, n34133, n34134, n34135, n34136, n34137, n34138,
         n34139, n34140, n34141, n34142, n34143, n34144, n34145, n34146,
         n34147, n34148, n34149, n34150, n34151, n34152, n34153, n34154,
         n34155, n34156, n34157, n34158, n34159, n34160, n34161, n34162,
         n34163, n34164, n34165, n34166, n34167, n34168, n34169, n34170,
         n34171, n34172, n34173, n34174, n34175, n34176, n34177, n34178,
         n34179, n34180, n34181, n34182, n34183, n34184, n34185, n34186,
         n34187, n34188, n34189, n34190, n34191, n34192, n34193, n34194,
         n34195, n34196, n34197, n34198, n34199, n34200, n34201, n34202,
         n34203, n34204, n34205, n34206, n34207, n34208, n34209, n34210,
         n34211, n34212, n34213, n34214, n34215, n34216, n34217, n34218,
         n34219, n34220, n34221, n34222, n34223, n34224, n34225, n34226,
         n34227, n34228, n34229, n34230, n34231, n34232, n34233, n34234,
         n34235, n34236, n34237, n34238, n34239, n34240, n34241, n34242,
         n34243, n34244, n34245, n34246, n34247, n34248, n34249, n34250,
         n34251, n34252, n34253, n34254, n34255, n34256, n34257, n34258,
         n34259, n34260, n34261, n34262, n34263, n34264, n34265, n34266,
         n34267, n34268, n34269, n34270, n34271, n34272, n34273, n34274,
         n34275, n34276, n34277, n34278, n34279, n34280, n34281, n34282,
         n34283, n34284, n34285, n34286, n34287, n34288, n34289, n34290,
         n34291, n34292, n34293, n34294, n34295, n34296, n34297, n34298,
         n34299, n34300, n34301, n34302, n34303, n34304, n34305, n34306,
         n34307, n34308, n34309, n34310, n34311, n34312, n34313, n34314,
         n34315, n34316, n34317, n34318, n34319, n34320, n34321, n34322,
         n34323, n34324, n34325, n34326, n34327, n34328, n34329, n34330,
         n34331, n34332, n34333, n34334, n34335, n34336, n34337, n34338,
         n34339, n34340, n34341, n34342, n34343, n34344, n34345, n34346,
         n34347, n34348, n34349, n34350, n34351, n34352, n34353, n34354,
         n34355, n34356, n34357, n34358, n34359, n34360, n34361, n34362,
         n34363, n34364, n34365, n34366, n34367, n34368, n34369, n34370,
         n34371, n34372, n34373, n34374, n34375, n34376, n34377, n34378,
         n34379, n34380, n34381, n34382, n34383, n34384, n34385, n34386,
         n34387, n34388, n34389, n34390, n34391, n34392, n34393, n34394,
         n34395, n34396, n34397, n34398, n34399, n34400, n34401, n34402,
         n34403, n34404, n34405, n34406, n34407, n34408, n34409, n34410,
         n34411, n34412, n34413, n34414, n34415, n34416, n34417, n34418,
         n34419, n34420, n34421, n34422, n34423, n34424, n34425, n34426,
         n34427, n34428, n34429, n34430, n34431, n34432, n34433, n34434,
         n34435, n34436, n34437, n34438, n34439, n34440, n34441, n34442,
         n34443, n34444, n34445, n34446, n34447, n34448, n34449, n34450,
         n34451, n34452, n34453, n34454, n34455, n34456, n34457, n34458,
         n34459, n34460, n34461, n34462, n34463, n34464, n34465, n34466,
         n34467, n34468, n34469, n34470, n34471, n34472, n34473, n34474,
         n34475, n34476, n34477, n34478, n34479, n34480, n34481, n34482,
         n34483, n34484, n34485, n34486, n34487, n34488, n34489, n34490,
         n34491, n34492, n34493, n34494, n34495, n34496, n34497, n34498,
         n34499, n34500, n34501, n34502, n34503, n34504, n34505, n34506,
         n34507, n34508, n34509, n34510, n34511, n34512, n34513, n34514,
         n34515, n34516, n34517, n34518, n34519, n34520, n34521, n34522,
         n34523, n34524, n34525, n34526, n34527, n34528, n34529, n34530,
         n34531, n34532, n34533, n34534, n34535, n34536, n34537, n34538,
         n34539, n34540, n34541, n34542, n34543, n34544, n34545, n34546,
         n34547, n34548, n34549, n34550, n34551, n34552, n34553, n34554,
         n34555, n34556, n34557, n34558, n34559, n34560, n34561, n34562,
         n34563, n34564, n34565, n34566, n34567, n34568, n34569, n34570,
         n34571, n34572, n34573, n34574, n34575, n34576, n34577, n34578,
         n34579, n34580, n34581, n34582, n34583, n34584, n34585, n34586,
         n34587, n34588, n34589, n34590, n34591, n34592, n34593, n34594,
         n34595, n34596, n34597, n34598, n34599, n34600, n34601, n34602,
         n34603, n34604, n34605, n34606, n34607, n34608, n34609, n34610,
         n34611, n34612, n34613, n34614, n34615, n34616, n34617, n34618,
         n34619, n34620, n34621, n34622, n34623, n34624, n34625, n34626,
         n34627, n34628, n34629, n34630, n34631, n34632, n34633, n34634,
         n34635, n34636, n34637, n34638, n34639, n34640, n34641, n34642,
         n34643, n34644, n34645, n34646, n34647, n34648, n34649, n34650,
         n34651, n34652, n34653, n34654, n34655, n34656, n34657, n34658,
         n34659, n34660, n34661, n34662, n34663, n34664, n34665, n34666,
         n34667, n34668, n34669, n34670, n34671, n34672, n34673, n34674,
         n34675, n34676, n34677, n34678, n34679, n34680, n34681, n34682,
         n34683, n34684, n34685, n34686, n34687, n34688, n34689, n34690,
         n34691, n34692, n34693, n34694, n34695, n34696, n34697, n34698,
         n34699, n34700, n34701, n34702, n34703, n34704, n34705, n34706,
         n34707, n34708, n34709, n34710, n34711, n34712, n34713, n34714,
         n34715, n34716, n34717, n34718, n34719, n34720, n34721, n34722,
         n34723, n34724, n34725, n34726, n34727, n34728, n34729, n34730,
         n34731, n34732, n34733, n34734, n34735, n34736, n34737, n34738,
         n34739, n34740, n34741, n34742, n34743, n34744, n34745, n34746,
         n34747, n34748, n34749, n34750, n34751, n34752, n34753, n34754,
         n34755, n34756, n34757, n34758, n34759, n34760, n34761, n34762,
         n34763, n34764, n34765, n34766, n34767, n34768, n34769, n34770,
         n34771, n34772, n34773, n34774, n34775, n34776, n34777, n34778,
         n34779, n34780, n34781, n34782, n34783, n34784, n34785, n34786,
         n34787, n34788, n34789, n34790, n34791, n34792, n34793, n34794,
         n34795, n34796, n34797, n34798, n34799, n34800, n34801, n34802,
         n34803, n34804, n34805, n34806, n34807, n34808, n34809, n34810,
         n34811, n34812, n34813, n34814, n34815, n34816, n34817, n34818,
         n34819, n34820, n34821, n34822, n34823, n34824, n34825, n34826,
         n34827, n34828, n34829, n34830, n34831, n34832, n34833, n34834,
         n34835, n34836, n34837, n34838, n34839, n34840, n34841, n34842,
         n34843, n34844, n34845, n34846, n34847, n34848, n34849, n34850,
         n34851, n34852, n34853, n34854, n34855, n34856, n34857, n34858,
         n34859, n34860, n34861, n34862, n34863, n34864, n34865, n34866,
         n34867, n34868, n34869, n34870, n34871, n34872, n34873, n34874,
         n34875, n34876, n34877, n34878, n34879, n34880, n34881, n34882,
         n34883, n34884, n34885, n34886, n34887, n34888, n34889, n34890,
         n34891, n34892, n34893, n34894, n34895, n34896, n34897, n34898,
         n34899, n34900, n34901, n34902, n34903, n34904, n34905, n34906,
         n34907, n34908, n34909, n34910, n34911, n34912, n34913, n34914,
         n34915, n34916, n34917, n34918, n34919, n34920, n34921, n34922,
         n34923, n34924, n34925, n34926, n34927, n34928, n34929, n34930,
         n34931, n34932, n34933, n34934, n34935, n34936, n34937, n34938,
         n34939, n34940, n34941, n34942, n34943, n34944, n34945, n34946,
         n34947, n34948, n34949, n34950, n34951, n34952, n34953, n34954,
         n34955, n34956, n34957, n34958, n34959, n34960, n34961, n34962,
         n34963, n34964, n34965, n34966, n34967, n34968, n34969, n34970,
         n34971, n34972, n34973, n34974, n34975, n34976, n34977, n34978,
         n34979, n34980, n34981, n34982, n34983, n34984, n34985, n34986,
         n34987, n34988, n34989, n34990, n34991, n34992, n34993, n34994,
         n34995, n34996, n34997, n34998, n34999, n35000, n35001, n35002,
         n35003, n35004, n35005, n35006, n35007, n35008, n35009, n35010,
         n35011, n35012, n35013, n35014, n35015, n35016, n35017, n35018,
         n35019, n35020, n35021, n35022, n35023, n35024, n35025, n35026,
         n35027, n35028, n35029, n35030, n35031, n35032, n35033, n35034,
         n35035, n35036, n35037, n35038, n35039, n35040, n35041, n35042,
         n35043, n35044, n35045, n35046, n35047, n35048, n35049, n35050,
         n35051, n35052, n35053, n35054, n35055, n35056, n35057, n35058,
         n35059, n35060, n35061, n35062, n35063, n35064, n35065, n35066,
         n35067, n35068, n35069, n35070, n35071, n35072, n35073, n35074,
         n35075, n35076, n35077, n35078, n35079, n35080, n35081, n35082,
         n35083, n35084, n35085, n35086, n35087, n35088, n35089, n35090,
         n35091, n35092, n35093, n35094, n35095, n35096, n35097, n35098,
         n35099, n35100, n35101, n35102, n35103, n35104, n35105, n35106,
         n35107, n35108, n35109, n35110, n35111, n35112, n35113, n35114,
         n35115, n35116, n35117, n35118, n35119, n35120, n35121, n35122,
         n35123, n35124, n35125, n35126, n35127, n35128, n35129, n35130,
         n35131, n35132, n35133, n35134, n35135, n35136, n35137, n35138,
         n35139, n35140, n35141, n35142, n35143, n35144, n35145, n35146,
         n35147, n35148, n35149, n35150, n35151, n35152, n35153, n35154,
         n35155, n35156, n35157, n35158, n35159, n35160, n35161, n35162,
         n35163, n35164, n35165, n35166, n35167, n35168, n35169, n35170,
         n35171, n35172, n35173, n35174, n35175, n35176, n35177, n35178,
         n35179, n35180, n35181, n35182, n35183, n35184, n35185, n35186,
         n35187, n35188, n35189, n35190, n35191, n35192, n35193, n35194,
         n35195, n35196, n35197, n35198, n35199, n35200, n35201, n35202,
         n35203, n35204, n35205, n35206, n35207, n35208, n35209, n35210,
         n35211, n35212, n35213, n35214, n35215, n35216, n35217, n35218,
         n35219, n35220, n35221, n35222, n35223, n35224, n35225, n35226,
         n35227, n35228, n35229, n35230, n35231, n35232, n35233, n35234,
         n35235, n35236, n35237, n35238, n35239, n35240, n35241, n35242,
         n35243, n35244, n35245, n35246, n35247, n35248, n35249, n35250,
         n35251, n35252, n35253, n35254, n35255, n35256, n35257, n35258,
         n35259, n35260, n35261, n35262, n35263, n35264, n35265, n35266,
         n35267, n35268, n35269, n35270, n35271, n35272, n35273, n35274,
         n35275, n35276, n35277, n35278, n35279, n35280, n35281, n35282,
         n35283, n35284, n35285, n35286, n35287, n35288, n35289, n35290,
         n35291, n35292, n35293, n35294, n35295, n35296, n35297, n35298,
         n35299, n35300, n35301, n35302, n35303, n35304, n35305, n35306,
         n35307, n35308, n35309, n35310, n35311, n35312, n35313, n35314,
         n35315, n35316, n35317, n35318, n35319, n35320, n35321, n35322,
         n35323, n35324, n35325, n35326, n35327, n35328, n35329, n35330,
         n35331, n35332, n35333, n35334, n35335, n35336, n35337, n35338,
         n35339, n35340, n35341, n35342, n35343, n35344, n35345, n35346,
         n35347, n35348, n35349, n35350, n35351, n35352, n35353, n35354,
         n35355, n35356, n35357, n35358, n35359, n35360, n35361, n35362,
         n35363, n35364, n35365, n35366, n35367, n35368, n35369, n35370,
         n35371, n35372, n35373, n35374, n35375, n35376, n35377, n35378,
         n35379, n35380, n35381, n35382, n35383, n35384, n35385, n35386,
         n35387, n35388, n35389, n35390, n35391, n35392, n35393, n35394,
         n35395, n35396, n35397, n35398, n35399, n35400, n35401, n35402,
         n35403, n35404, n35405, n35406, n35407, n35408, n35409, n35410,
         n35411, n35412, n35413, n35414, n35415, n35416, n35417, n35418,
         n35419, n35420, n35421, n35422, n35423, n35424, n35425, n35426,
         n35427, n35428, n35429, n35430, n35431, n35432, n35433, n35434,
         n35435, n35436, n35437, n35438, n35439, n35440, n35441, n35442,
         n35443, n35444, n35445, n35446, n35447, n35448, n35449, n35450,
         n35451, n35452, n35453, n35454, n35455, n35456, n35457, n35458,
         n35459, n35460, n35461, n35462, n35463, n35464, n35465, n35466,
         n35467, n35468, n35469, n35470, n35471, n35472, n35473, n35474,
         n35475, n35476, n35477, n35478, n35479, n35480, n35481, n35482,
         n35483, n35484, n35485, n35486, n35487, n35488, n35489, n35490,
         n35491, n35492, n35493, n35494, n35495, n35496, n35497, n35498,
         n35499, n35500, n35501, n35502, n35503, n35504, n35505, n35506,
         n35507, n35508, n35509, n35510, n35511, n35512, n35513, n35514,
         n35515, n35516, n35517, n35518, n35519, n35520, n35521, n35522,
         n35523, n35524, n35525, n35526, n35527, n35528, n35529, n35530,
         n35531, n35532, n35533, n35534, n35535, n35536, n35537, n35538,
         n35539, n35540, n35541, n35542, n35543, n35544, n35545, n35546,
         n35547, n35548, n35549, n35550, n35551, n35552, n35553, n35554,
         n35555, n35556, n35557, n35558, n35559, n35560, n35561, n35562,
         n35563, n35564, n35565, n35566, n35567, n35568, n35569, n35570,
         n35571, n35572, n35573, n35574, n35575, n35576, n35577, n35578,
         n35579, n35580, n35581, n35582, n35583, n35584, n35585, n35586,
         n35587, n35588, n35589, n35590, n35591, n35592, n35593, n35594,
         n35595, n35596, n35597, n35598, n35599, n35600, n35601, n35602,
         n35603, n35604, n35605, n35606, n35607, n35608, n35609, n35610,
         n35611, n35612, n35613, n35614, n35615, n35616, n35617, n35618,
         n35619, n35620, n35621, n35622, n35623, n35624, n35625, n35626,
         n35627, n35628, n35629, n35630, n35631, n35632, n35633, n35634,
         n35635, n35636, n35637, n35638, n35639, n35640, n35641, n35642,
         n35643, n35644, n35645, n35646, n35647, n35648, n35649, n35650,
         n35651, n35652, n35653, n35654, n35655, n35656, n35657, n35658,
         n35659, n35660, n35661, n35662, n35663, n35664, n35665, n35666,
         n35667, n35668, n35669, n35670, n35671, n35672, n35673, n35674,
         n35675, n35676, n35677, n35678, n35679, n35680, n35681, n35682,
         n35683, n35684, n35685, n35686, n35687, n35688, n35689, n35690,
         n35691, n35692, n35693, n35694, n35695, n35696, n35697, n35698,
         n35699, n35700, n35701, n35702, n35703, n35704, n35705, n35706,
         n35707, n35708, n35709, n35710, n35711, n35712, n35713, n35714,
         n35715, n35716, n35717, n35718, n35719, n35720, n35721, n35722,
         n35723, n35724, n35725, n35726, n35727, n35728, n35729, n35730,
         n35731, n35732, n35733, n35734, n35735, n35736, n35737, n35738,
         n35739, n35740, n35741, n35742, n35743, n35744, n35745, n35746,
         n35747, n35748, n35749, n35750, n35751, n35752, n35753, n35754,
         n35755, n35756, n35757, n35758, n35759, n35760, n35761, n35762,
         n35763, n35764, n35765, n35766, n35767, n35768, n35769, n35770,
         n35771, n35772, n35773, n35774, n35775, n35776, n35777, n35778,
         n35779, n35780, n35781, n35782, n35783, n35784, n35785, n35786,
         n35787, n35788, n35789, n35790, n35791, n35792, n35793, n35794,
         n35795, n35796, n35797, n35798, n35799, n35800, n35801, n35802,
         n35803, n35804, n35805, n35806, n35807, n35808, n35809, n35810,
         n35811, n35812, n35813, n35814, n35815, n35816, n35817, n35818,
         n35819, n35820, n35821, n35822, n35823, n35824, n35825, n35826,
         n35827, n35828, n35829, n35830, n35831, n35832, n35833, n35834,
         n35835, n35836, n35837, n35838, n35839, n35840, n35841, n35842,
         n35843, n35844, n35845, n35846, n35847, n35848, n35849, n35850,
         n35851, n35852, n35853, n35854, n35855, n35856, n35857, n35858,
         n35859, n35860, n35861, n35862, n35863, n35864, n35865, n35866,
         n35867, n35868, n35869, n35870, n35871, n35872, n35873, n35874,
         n35875, n35876, n35877, n35878, n35879, n35880, n35881, n35882,
         n35883, n35884, n35885, n35886, n35887, n35888, n35889, n35890,
         n35891, n35892, n35893, n35894, n35895, n35896, n35897, n35898,
         n35899, n35900, n35901, n35902, n35903, n35904, n35905, n35906,
         n35907, n35908, n35909, n35910, n35911, n35912, n35913, n35914,
         n35915, n35916, n35917, n35918, n35919, n35920, n35921, n35922,
         n35923, n35924, n35925, n35926, n35927, n35928, n35929, n35930,
         n35931, n35932, n35933, n35934, n35935, n35936, n35937, n35938,
         n35939, n35940, n35941, n35942, n35943, n35944, n35945, n35946,
         n35947, n35948, n35949, n35950, n35951, n35952, n35953, n35954,
         n35955, n35956, n35957, n35958, n35959, n35960, n35961, n35962,
         n35963, n35964, n35965, n35966, n35967, n35968, n35969, n35970,
         n35971, n35972, n35973, n35974, n35975, n35976, n35977, n35978,
         n35979, n35980, n35981, n35982, n35983, n35984, n35985, n35986,
         n35987, n35988, n35989, n35990, n35991, n35992, n35993, n35994,
         n35995, n35996, n35997, n35998, n35999, n36000, n36001, n36002,
         n36003, n36004, n36005, n36006, n36007, n36008, n36009, n36010,
         n36011, n36012, n36013, n36014, n36015, n36016, n36017, n36018,
         n36019, n36020, n36021, n36022, n36023, n36024, n36025, n36026,
         n36027, n36028, n36029, n36030, n36031, n36032, n36033, n36034,
         n36035, n36036, n36037, n36038, n36039, n36040, n36041, n36042,
         n36043, n36044, n36045, n36046, n36047, n36048, n36049, n36050,
         n36051, n36052, n36053, n36054, n36055, n36056, n36057, n36058,
         n36059, n36060, n36061, n36062, n36063, n36064, n36065, n36066,
         n36067, n36068, n36069, n36070, n36071, n36072, n36073, n36074,
         n36075, n36076, n36077, n36078, n36079, n36080, n36081, n36082,
         n36083, n36084, n36085, n36086, n36087, n36088, n36089, n36090,
         n36091, n36092, n36093, n36094, n36095, n36096, n36097, n36098,
         n36099, n36100, n36101, n36102, n36103, n36104, n36105, n36106,
         n36107, n36108, n36109, n36110, n36111, n36112, n36113, n36114,
         n36115, n36116, n36117, n36118, n36119, n36120, n36121, n36122,
         n36123, n36124, n36125, n36126, n36127, n36128, n36129, n36130,
         n36131, n36132, n36133, n36134, n36135, n36136, n36137, n36138,
         n36139, n36140, n36141, n36142, n36143, n36144, n36145, n36146,
         n36147, n36148, n36149, n36150, n36151, n36152, n36153, n36154,
         n36155, n36156, n36157, n36158, n36159, n36160, n36161, n36162,
         n36163, n36164, n36165, n36166, n36167, n36168, n36169, n36170,
         n36171, n36172, n36173, n36174, n36175, n36176, n36177, n36178,
         n36179, n36180, n36181, n36182, n36183, n36184, n36185, n36186,
         n36187, n36188, n36189, n36190, n36191, n36192, n36193, n36194,
         n36195, n36196, n36197, n36198, n36199, n36200, n36201, n36202,
         n36203, n36204, n36205, n36206, n36207, n36208, n36209, n36210,
         n36211, n36212, n36213, n36214, n36215, n36216, n36217, n36218,
         n36219, n36220, n36221, n36222, n36223, n36224, n36225, n36226,
         n36227, n36228, n36229, n36230, n36231, n36232, n36233, n36234,
         n36235, n36236, n36237, n36238, n36239, n36240, n36241, n36242,
         n36243, n36244, n36245, n36246, n36247, n36248, n36249, n36250,
         n36251, n36252, n36253, n36254, n36255, n36256, n36257, n36258,
         n36259, n36260, n36261, n36262, n36263, n36264, n36265, n36266,
         n36267, n36268, n36269, n36270, n36271, n36272, n36273, n36274,
         n36275, n36276, n36277, n36278, n36279, n36280, n36281, n36282,
         n36283, n36284, n36285, n36286, n36287, n36288, n36289, n36290,
         n36291, n36292, n36293, n36294, n36295, n36296, n36297, n36298,
         n36299, n36300, n36301, n36302, n36303, n36304, n36305, n36306,
         n36307, n36308, n36309, n36310, n36311, n36312, n36313, n36314,
         n36315, n36316, n36317, n36318, n36319, n36320, n36321, n36322,
         n36323, n36324, n36325, n36326, n36327, n36328, n36329, n36330,
         n36331, n36332, n36333, n36334, n36335, n36336, n36337, n36338,
         n36339, n36340, n36341, n36342, n36343, n36344, n36345, n36346,
         n36347, n36348, n36349, n36350, n36351, n36352, n36353, n36354,
         n36355, n36356, n36357, n36358, n36359, n36360, n36361, n36362,
         n36363, n36364, n36365, n36366, n36367, n36368, n36369, n36370,
         n36371, n36372, n36373, n36374, n36375, n36376, n36377, n36378,
         n36379, n36380, n36381, n36382, n36383, n36384, n36385, n36386,
         n36387, n36388, n36389, n36390, n36391, n36392, n36393, n36394,
         n36395, n36396, n36397, n36398, n36399, n36400, n36401, n36402,
         n36403, n36404, n36405, n36406, n36407, n36408, n36409, n36410,
         n36411, n36412, n36413, n36414, n36415, n36416, n36417, n36418,
         n36419, n36420, n36421, n36422, n36423, n36424, n36425, n36426,
         n36427, n36428, n36429, n36430, n36431, n36432, n36433, n36434,
         n36435, n36436, n36437, n36438, n36439, n36440, n36441, n36442,
         n36443, n36444, n36445, n36446, n36447, n36448, n36449, n36450,
         n36451, n36452, n36453, n36454, n36455, n36456, n36457, n36458,
         n36459, n36460, n36461, n36462, n36463, n36464, n36465, n36466,
         n36467, n36468, n36469, n36470, n36471, n36472, n36473, n36474,
         n36475, n36476, n36477, n36478, n36479, n36480, n36481, n36482,
         n36483, n36484, n36485, n36486, n36487, n36488, n36489, n36490,
         n36491, n36492, n36493, n36494, n36495, n36496, n36497, n36498,
         n36499, n36500, n36501, n36502, n36503, n36504, n36505, n36506,
         n36507, n36508, n36509, n36510, n36511, n36512, n36513, n36514,
         n36515, n36516, n36517, n36518, n36519, n36520, n36521, n36522,
         n36523, n36524, n36525, n36526, n36527, n36528, n36529, n36530,
         n36531, n36532, n36533, n36534, n36535, n36536, n36537, n36538,
         n36539, n36540, n36541, n36542, n36543, n36544, n36545, n36546,
         n36547, n36548, n36549, n36550, n36551, n36552, n36553, n36554,
         n36555, n36556, n36557, n36558, n36559, n36560, n36561, n36562,
         n36563, n36564, n36565, n36566, n36567, n36568, n36569, n36570,
         n36571, n36572, n36573, n36574, n36575, n36576, n36577, n36578,
         n36579, n36580, n36581, n36582, n36583, n36584, n36585, n36586,
         n36587, n36588, n36589, n36590, n36591, n36592, n36593, n36594,
         n36595, n36596, n36597, n36598, n36599, n36600, n36601, n36602,
         n36603, n36604, n36605, n36606, n36607, n36608, n36609, n36610,
         n36611, n36612, n36613, n36614, n36615, n36616, n36617, n36618,
         n36619, n36620, n36621, n36622, n36623, n36624, n36625, n36626,
         n36627, n36628, n36629, n36630, n36631, n36632, n36633, n36634,
         n36635, n36636, n36637, n36638, n36639, n36640, n36641, n36642,
         n36643, n36644, n36645, n36646, n36647, n36648, n36649, n36650,
         n36651, n36652, n36653, n36654, n36655, n36656, n36657, n36658,
         n36659, n36660, n36661, n36662, n36663, n36664, n36665, n36666,
         n36667, n36668, n36669, n36670, n36671, n36672, n36673, n36674,
         n36675, n36676, n36677, n36678, n36679, n36680, n36681, n36682,
         n36683, n36684, n36685, n36686, n36687, n36688, n36689, n36690,
         n36691, n36692, n36693, n36694, n36695, n36696, n36697, n36698,
         n36699, n36700, n36701, n36702, n36703, n36704, n36705, n36706,
         n36707, n36708, n36709, n36710, n36711, n36712, n36713, n36714,
         n36715, n36716, n36717, n36718, n36719, n36720, n36721, n36722,
         n36723, n36724, n36725, n36726, n36727, n36728, n36729, n36730,
         n36731, n36732, n36733, n36734, n36735, n36736, n36737, n36738,
         n36739, n36740, n36741, n36742, n36743, n36744, n36745, n36746,
         n36747, n36748, n36749, n36750, n36751, n36752, n36753, n36754,
         n36755, n36756, n36757, n36758, n36759, n36760, n36761, n36762,
         n36763, n36764, n36765, n36766, n36767, n36768, n36769, n36770,
         n36771, n36772, n36773, n36774, n36775, n36776, n36777, n36778,
         n36779, n36780, n36781, n36782, n36783, n36784, n36785, n36786,
         n36787, n36788, n36789, n36790, n36791, n36792, n36793, n36794,
         n36795, n36796, n36797, n36798, n36799, n36800, n36801, n36802,
         n36803, n36804, n36805, n36806, n36807, n36808, n36809, n36810,
         n36811, n36812, n36813, n36814, n36815, n36816, n36817, n36818,
         n36819, n36820, n36821, n36822, n36823, n36824, n36825, n36826,
         n36827, n36828, n36829, n36830, n36831, n36832, n36833, n36834,
         n36835, n36836, n36837, n36838, n36839, n36840, n36841, n36842,
         n36843, n36844, n36845, n36846, n36847, n36848, n36849, n36850,
         n36851, n36852, n36853, n36854, n36855, n36856, n36857, n36858,
         n36859, n36860, n36861, n36862, n36863, n36864, n36865, n36866,
         n36867, n36868, n36869, n36870, n36871, n36872, n36873, n36874,
         n36875, n36876, n36877, n36878, n36879, n36880, n36881, n36882,
         n36883, n36884, n36885, n36886, n36887, n36888, n36889, n36890,
         n36891, n36892, n36893, n36894, n36895, n36896, n36897, n36898,
         n36899, n36900, n36901, n36902, n36903, n36904, n36905, n36906,
         n36907, n36908, n36909, n36910, n36911, n36912, n36913, n36914,
         n36915, n36916, n36917, n36918, n36919, n36920, n36921, n36922,
         n36923, n36924, n36925, n36926, n36927, n36928, n36929, n36930,
         n36931, n36932, n36933, n36934, n36935, n36936, n36937, n36938,
         n36939, n36940, n36941, n36942, n36943, n36944, n36945, n36946,
         n36947, n36948, n36949, n36950, n36951, n36952, n36953, n36954,
         n36955, n36956, n36957, n36958, n36959, n36960, n36961, n36962,
         n36963, n36964, n36965, n36966, n36967, n36968, n36969, n36970,
         n36971, n36972, n36973, n36974, n36975, n36976, n36977, n36978,
         n36979, n36980, n36981, n36982, n36983, n36984, n36985, n36986,
         n36987, n36988, n36989, n36990, n36991, n36992, n36993, n36994,
         n36995, n36996, n36997, n36998, n36999, n37000, n37001, n37002,
         n37003, n37004, n37005, n37006, n37007, n37008, n37009, n37010,
         n37011, n37012, n37013, n37014, n37015, n37016, n37017, n37018,
         n37019, n37020, n37021, n37022, n37023, n37024, n37025, n37026,
         n37027, n37028, n37029, n37030, n37031, n37032, n37033, n37034,
         n37035, n37036, n37037, n37038, n37039, n37040, n37041, n37042,
         n37043, n37044, n37045, n37046, n37047, n37048, n37049, n37050,
         n37051, n37052, n37053, n37054, n37055, n37056, n37057, n37058,
         n37059, n37060, n37061, n37062, n37063, n37064, n37065, n37066,
         n37067, n37068, n37069, n37070, n37071, n37072, n37073, n37074,
         n37075, n37076, n37077, n37078, n37079, n37080, n37081, n37082,
         n37083, n37084, n37085, n37086, n37087, n37088, n37089, n37090,
         n37091, n37092, n37093, n37094, n37095, n37096, n37097, n37098,
         n37099, n37100, n37101, n37102, n37103, n37104, n37105, n37106,
         n37107, n37108, n37109, n37110, n37111, n37112, n37113, n37114,
         n37115, n37116, n37117, n37118, n37119, n37120, n37121, n37122,
         n37123, n37124, n37125, n37126, n37127, n37128, n37129, n37130,
         n37131, n37132, n37133, n37134, n37135, n37136, n37137, n37138,
         n37139, n37140, n37141, n37142, n37143, n37144, n37145, n37146,
         n37147, n37148, n37149, n37150, n37151, n37152, n37153, n37154,
         n37155, n37156, n37157, n37158, n37159, n37160, n37161, n37162,
         n37163, n37164, n37165, n37166, n37167, n37168, n37169, n37170,
         n37171, n37172, n37173, n37174, n37175, n37176, n37177, n37178,
         n37179, n37180, n37181, n37182, n37183, n37184, n37185, n37186,
         n37187, n37188, n37189, n37190, n37191, n37192, n37193, n37194,
         n37195, n37196, n37197, n37198, n37199, n37200, n37201, n37202,
         n37203, n37204, n37205, n37206, n37207, n37208, n37209, n37210,
         n37211, n37212, n37213, n37214, n37215, n37216, n37217, n37218,
         n37219, n37220, n37221, n37222, n37223, n37224, n37225, n37226,
         n37227, n37228, n37229, n37230, n37231, n37232, n37233, n37234,
         n37235, n37236, n37237, n37238, n37239, n37240, n37241, n37242,
         n37243, n37244, n37245, n37246, n37247, n37248, n37249, n37250,
         n37251, n37252, n37253, n37254, n37255, n37256, n37257, n37258,
         n37259, n37260, n37261, n37262, n37263, n37264, n37265, n37266,
         n37267, n37268, n37269, n37270, n37271, n37272, n37273, n37274,
         n37275, n37276, n37277, n37278, n37279, n37280, n37281, n37282,
         n37283, n37284, n37285, n37286, n37287, n37288, n37289, n37290,
         n37291, n37292, n37293, n37294, n37295, n37296, n37297, n37298,
         n37299, n37300, n37301, n37302, n37303, n37304, n37305, n37306,
         n37307, n37308, n37309, n37310, n37311, n37312, n37313, n37314,
         n37315, n37316, n37317, n37318, n37319, n37320, n37321, n37322,
         n37323, n37324, n37325, n37326, n37327, n37328, n37329, n37330,
         n37331, n37332, n37333, n37334, n37335, n37336, n37337, n37338,
         n37339, n37340, n37341, n37342, n37343, n37344, n37345, n37346,
         n37347, n37348, n37349, n37350, n37351, n37352, n37353, n37354,
         n37355, n37356, n37357, n37358, n37359, n37360, n37361, n37362,
         n37363, n37364, n37365, n37366, n37367, n37368, n37369, n37370,
         n37371, n37372, n37373, n37374, n37375, n37376, n37377, n37378,
         n37379, n37380, n37381, n37382, n37383, n37384, n37385, n37386,
         n37387, n37388, n37389, n37390, n37391, n37392, n37393, n37394,
         n37395, n37396, n37397, n37398, n37399, n37400, n37401, n37402,
         n37403, n37404, n37405, n37406, n37407, n37408, n37409, n37410,
         n37411, n37412, n37413, n37414, n37415, n37416, n37417, n37418,
         n37419, n37420, n37421, n37422, n37423, n37424, n37425, n37426,
         n37427, n37428, n37429, n37430, n37431, n37432, n37433, n37434,
         n37435, n37436, n37437, n37438, n37439, n37440, n37441, n37442,
         n37443, n37444, n37445, n37446, n37447, n37448, n37449, n37450,
         n37451, n37452, n37453, n37454, n37455, n37456, n37457, n37458,
         n37459, n37460, n37461, n37462, n37463, n37464, n37465, n37466,
         n37467, n37468, n37469, n37470, n37471, n37472, n37473, n37474,
         n37475, n37476, n37477, n37478, n37479, n37480, n37481, n37482,
         n37483, n37484, n37485, n37486, n37487, n37488, n37489, n37490,
         n37491, n37492, n37493, n37494, n37495, n37496, n37497, n37498,
         n37499, n37500, n37501, n37502, n37503, n37504, n37505, n37506,
         n37507, n37508, n37509, n37510, n37511, n37512, n37513, n37514,
         n37515, n37516, n37517, n37518, n37519, n37520, n37521, n37522,
         n37523, n37524, n37525, n37526, n37527, n37528, n37529, n37530,
         n37531, n37532, n37533, n37534, n37535, n37536, n37537, n37538,
         n37539, n37540, n37541, n37542, n37543, n37544, n37545, n37546,
         n37547, n37548, n37549, n37550, n37551, n37552, n37553, n37554,
         n37555, n37556, n37557, n37558, n37559, n37560, n37561, n37562,
         n37563, n37564, n37565, n37566, n37567, n37568, n37569, n37570,
         n37571, n37572, n37573, n37574, n37575, n37576, n37577, n37578,
         n37579, n37580, n37581, n37582, n37583, n37584, n37585, n37586,
         n37587, n37588, n37589, n37590, n37591, n37592, n37593, n37594,
         n37595, n37596, n37597, n37598, n37599, n37600, n37601, n37602,
         n37603, n37604, n37605, n37606, n37607, n37608, n37609, n37610,
         n37611, n37612, n37613, n37614, n37615, n37616, n37617, n37618,
         n37619, n37620, n37621, n37622, n37623, n37624, n37625, n37626,
         n37627, n37628, n37629, n37630, n37631, n37632, n37633, n37634,
         n37635, n37636, n37637, n37638, n37639, n37640, n37641, n37642,
         n37643, n37644, n37645, n37646, n37647, n37648, n37649, n37650,
         n37651, n37652, n37653, n37654, n37655, n37656, n37657, n37658,
         n37659, n37660, n37661, n37662, n37663, n37664, n37665, n37666,
         n37667, n37668, n37669, n37670, n37671, n37672, n37673, n37674,
         n37675, n37676, n37677, n37678, n37679, n37680, n37681, n37682,
         n37683, n37684, n37685, n37686, n37687, n37688, n37689, n37690,
         n37691, n37692, n37693, n37694, n37695, n37696, n37697, n37698,
         n37699, n37700, n37701, n37702, n37703, n37704, n37705, n37706,
         n37707, n37708, n37709, n37710, n37711, n37712, n37713, n37714,
         n37715, n37716, n37717, n37718, n37719, n37720, n37721, n37722,
         n37723, n37724, n37725, n37726, n37727, n37728, n37729, n37730,
         n37731, n37732, n37733, n37734, n37735, n37736, n37737, n37738,
         n37739, n37740, n37741, n37742, n37743, n37744, n37745, n37746,
         n37747, n37748, n37749, n37750, n37751, n37752, n37753, n37754,
         n37755, n37756, n37757, n37758, n37759, n37760, n37761, n37762,
         n37763, n37764, n37765, n37766, n37767, n37768, n37769, n37770,
         n37771, n37772, n37773, n37774, n37775, n37776, n37777, n37778,
         n37779, n37780, n37781, n37782, n37783, n37784, n37785, n37786,
         n37787, n37788, n37789, n37790, n37791, n37792, n37793, n37794,
         n37795, n37796, n37797, n37798, n37799, n37800, n37801, n37802,
         n37803, n37804, n37805, n37806, n37807, n37808, n37809, n37810,
         n37811, n37812, n37813, n37814, n37815, n37816, n37817, n37818,
         n37819, n37820, n37821, n37822, n37823, n37824, n37825, n37826,
         n37827, n37828, n37829, n37830, n37831, n37832, n37833, n37834,
         n37835, n37836, n37837, n37838, n37839, n37840, n37841, n37842,
         n37843, n37844, n37845, n37846, n37847, n37848, n37849, n37850,
         n37851, n37852, n37853, n37854, n37855, n37856, n37857, n37858,
         n37859, n37860, n37861, n37862, n37863, n37864, n37865, n37866,
         n37867, n37868, n37869, n37870, n37871, n37872, n37873, n37874,
         n37875, n37876, n37877, n37878, n37879, n37880, n37881, n37882,
         n37883, n37884, n37885, n37886, n37887, n37888, n37889, n37890,
         n37891, n37892, n37893, n37894, n37895, n37896, n37897, n37898,
         n37899, n37900, n37901, n37902, n37903, n37904, n37905, n37906,
         n37907, n37908, n37909, n37910, n37911, n37912, n37913, n37914,
         n37915, n37916, n37917, n37918, n37919, n37920, n37921, n37922,
         n37923, n37924, n37925, n37926, n37927, n37928, n37929, n37930,
         n37931, n37932, n37933, n37934, n37935, n37936, n37937, n37938,
         n37939, n37940, n37941, n37942, n37943, n37944, n37945, n37946,
         n37947, n37948, n37949, n37950, n37951, n37952, n37953, n37954,
         n37955, n37956, n37957, n37958, n37959, n37960, n37961, n37962,
         n37963, n37964, n37965, n37966, n37967, n37968, n37969, n37970,
         n37971, n37972, n37973, n37974, n37975, n37976, n37977, n37978,
         n37979, n37980, n37981, n37982, n37983, n37984, n37985, n37986,
         n37987, n37988, n37989, n37990, n37991, n37992, n37993, n37994,
         n37995, n37996, n37997, n37998, n37999, n38000, n38001, n38002,
         n38003, n38004, n38005, n38006, n38007, n38008, n38009, n38010,
         n38011, n38012, n38013, n38014, n38015, n38016, n38017, n38018,
         n38019, n38020, n38021, n38022, n38023, n38024, n38025, n38026,
         n38027, n38028, n38029, n38030, n38031, n38032, n38033, n38034,
         n38035, n38036, n38037, n38038, n38039, n38040, n38041, n38042,
         n38043, n38044, n38045, n38046, n38047, n38048, n38049, n38050,
         n38051, n38052, n38053, n38054, n38055, n38056, n38057, n38058,
         n38059, n38060, n38061, n38062, n38063, n38064, n38065, n38066,
         n38067, n38068, n38069, n38070, n38071, n38072, n38073, n38074,
         n38075, n38076, n38077, n38078, n38079, n38080, n38081, n38082,
         n38083, n38084, n38085, n38086, n38087, n38088, n38089, n38090,
         n38091, n38092, n38093, n38094, n38095, n38096, n38097, n38098,
         n38099, n38100, n38101, n38102, n38103, n38104, n38105, n38106,
         n38107, n38108, n38109, n38110, n38111, n38112, n38113, n38114,
         n38115, n38116, n38117, n38118, n38119, n38120, n38121, n38122,
         n38123, n38124, n38125, n38126, n38127, n38128, n38129, n38130,
         n38131, n38132, n38133, n38134, n38135, n38136, n38137, n38138,
         n38139, n38140, n38141, n38142, n38143, n38144, n38145, n38146,
         n38147, n38148, n38149, n38150, n38151, n38152, n38153, n38154,
         n38155, n38156, n38157, n38158, n38159, n38160, n38161, n38162,
         n38163, n38164, n38165, n38166, n38167, n38168, n38169, n38170,
         n38171, n38172, n38173, n38174, n38175, n38176, n38177, n38178,
         n38179, n38180, n38181, n38182, n38183, n38184, n38185, n38186,
         n38187, n38188, n38189, n38190, n38191, n38192, n38193, n38194,
         n38195, n38196, n38197, n38198, n38199, n38200, n38201, n38202,
         n38203, n38204, n38205, n38206, n38207, n38208, n38209, n38210,
         n38211, n38212, n38213, n38214, n38215, n38216, n38217, n38218,
         n38219, n38220, n38221, n38222, n38223, n38224, n38225, n38226,
         n38227, n38228, n38229, n38230, n38231, n38232, n38233, n38234,
         n38235, n38236, n38237, n38238, n38239, n38240, n38241, n38242,
         n38243, n38244, n38245, n38246, n38247, n38248, n38249, n38250,
         n38251, n38252, n38253, n38254, n38255, n38256, n38257, n38258,
         n38259, n38260, n38261, n38262, n38263, n38264, n38265, n38266,
         n38267, n38268, n38269, n38270, n38271, n38272, n38273, n38274,
         n38275, n38276, n38277, n38278, n38279, n38280, n38281, n38282,
         n38283, n38284, n38285, n38286, n38287, n38288, n38289, n38290,
         n38291, n38292, n38293, n38294, n38295, n38296, n38297, n38298,
         n38299, n38300, n38301, n38302, n38303, n38304, n38305, n38306,
         n38307, n38308, n38309, n38310, n38311, n38312, n38313, n38314,
         n38315, n38316, n38317, n38318, n38319, n38320, n38321, n38322,
         n38323, n38324, n38325, n38326, n38327, n38328, n38329, n38330,
         n38331, n38332, n38333, n38334, n38335, n38336, n38337, n38338,
         n38339, n38340, n38341, n38342, n38343, n38344, n38345, n38346,
         n38347, n38348, n38349, n38350, n38351, n38352, n38353, n38354,
         n38355, n38356, n38357, n38358, n38359, n38360, n38361, n38362,
         n38363, n38364, n38365, n38366, n38367, n38368, n38369, n38370,
         n38371, n38372, n38373, n38374, n38375, n38376, n38377, n38378,
         n38379, n38380, n38381, n38382, n38383, n38384, n38385, n38386,
         n38387, n38388, n38389, n38390, n38391, n38392, n38393, n38394,
         n38395, n38396, n38397, n38398, n38399, n38400, n38401, n38402,
         n38403, n38404, n38405, n38406, n38407, n38408, n38409, n38410,
         n38411, n38412, n38413, n38414, n38415, n38416, n38417, n38418,
         n38419, n38420, n38421, n38422, n38423, n38424, n38425, n38426,
         n38427, n38428, n38429, n38430, n38431, n38432, n38433, n38434,
         n38435, n38436, n38437, n38438, n38439, n38440, n38441, n38442,
         n38443, n38444, n38445, n38446, n38447, n38448, n38449, n38450,
         n38451, n38452, n38453, n38454, n38455, n38456, n38457, n38458,
         n38459, n38460, n38461, n38462, n38463, n38464, n38465, n38466,
         n38467, n38468, n38469, n38470, n38471, n38472, n38473, n38474,
         n38475, n38476, n38477, n38478, n38479, n38480, n38481, n38482,
         n38483, n38484, n38485, n38486, n38487, n38488, n38489, n38490,
         n38491, n38492, n38493, n38494, n38495, n38496, n38497, n38498,
         n38499, n38500, n38501, n38502, n38503, n38504, n38505, n38506,
         n38507, n38508, n38509, n38510, n38511, n38512, n38513, n38514,
         n38515, n38516, n38517, n38518, n38519, n38520, n38521, n38522,
         n38523, n38524, n38525, n38526, n38527, n38528, n38529, n38530,
         n38531, n38532, n38533, n38534, n38535, n38536, n38537, n38538,
         n38539, n38540, n38541, n38542, n38543, n38544, n38545, n38546,
         n38547, n38548, n38549, n38550, n38551, n38552, n38553, n38554,
         n38555, n38556, n38557, n38558, n38559, n38560, n38561, n38562,
         n38563, n38564, n38565, n38566, n38567, n38568, n38569, n38570,
         n38571, n38572, n38573, n38574, n38575, n38576, n38577, n38578,
         n38579, n38580, n38581, n38582, n38583, n38584, n38585, n38586,
         n38587, n38588, n38589, n38590, n38591, n38592, n38593, n38594,
         n38595, n38596, n38597, n38598, n38599, n38600, n38601, n38602,
         n38603, n38604, n38605, n38606, n38607, n38608, n38609, n38610,
         n38611, n38612, n38613, n38614, n38615, n38616, n38617, n38618,
         n38619, n38620, n38621, n38622, n38623, n38624, n38625, n38626,
         n38627, n38628, n38629, n38630, n38631, n38632, n38633, n38634,
         n38635, n38636, n38637, n38638, n38639, n38640, n38641, n38642,
         n38643, n38644, n38645, n38646, n38647, n38648, n38649, n38650,
         n38651, n38652, n38653, n38654, n38655, n38656, n38657, n38658,
         n38659, n38660, n38661, n38662, n38663, n38664, n38665, n38666,
         n38667, n38668, n38669, n38670, n38671, n38672, n38673, n38674,
         n38675, n38676, n38677, n38678, n38679, n38680, n38681, n38682,
         n38683, n38684, n38685, n38686, n38687, n38688, n38689, n38690,
         n38691, n38692, n38693, n38694, n38695, n38696, n38697, n38698,
         n38699, n38700, n38701, n38702, n38703, n38704, n38705, n38706,
         n38707, n38708, n38709, n38710, n38711, n38712, n38713, n38714,
         n38715, n38716, n38717, n38718, n38719, n38720, n38721, n38722,
         n38723, n38724, n38725, n38726, n38727, n38728, n38729, n38730,
         n38731, n38732, n38733, n38734, n38735, n38736, n38737, n38738,
         n38739, n38740, n38741, n38742, n38743, n38744, n38745, n38746,
         n38747, n38748, n38749, n38750, n38751, n38752, n38753, n38754,
         n38755, n38756, n38757, n38758, n38759, n38760, n38761, n38762,
         n38763, n38764, n38765, n38766, n38767, n38768, n38769, n38770,
         n38771, n38772, n38773, n38774, n38775, n38776, n38777, n38778,
         n38779, n38780, n38781, n38782, n38783, n38784, n38785, n38786,
         n38787, n38788, n38789, n38790, n38791, n38792, n38793, n38794,
         n38795, n38796, n38797, n38798, n38799, n38800, n38801, n38802,
         n38803, n38804, n38805, n38806, n38807, n38808, n38809, n38810,
         n38811, n38812, n38813, n38814, n38815, n38816, n38817, n38818,
         n38819, n38820, n38821, n38822, n38823, n38824, n38825, n38826,
         n38827, n38828, n38829, n38830, n38831, n38832, n38833, n38834,
         n38835, n38836, n38837, n38838, n38839, n38840, n38841, n38842,
         n38843, n38844, n38845, n38846, n38847, n38848, n38849, n38850,
         n38851, n38852, n38853, n38854, n38855, n38856, n38857, n38858,
         n38859, n38860, n38861, n38862, n38863, n38864, n38865, n38866,
         n38867, n38868, n38869, n38870, n38871, n38872, n38873, n38874,
         n38875, n38876, n38877, n38878, n38879, n38880, n38881, n38882,
         n38883, n38884, n38885, n38886, n38887, n38888, n38889, n38890,
         n38891, n38892, n38893, n38894, n38895, n38896, n38897, n38898,
         n38899, n38900, n38901, n38902, n38903, n38904, n38905, n38906,
         n38907, n38908, n38909, n38910, n38911, n38912, n38913, n38914,
         n38915, n38916, n38917, n38918, n38919, n38920, n38921, n38922,
         n38923, n38924, n38925, n38926, n38927, n38928, n38929, n38930,
         n38931, n38932, n38933, n38934, n38935, n38936, n38937, n38938,
         n38939, n38940, n38941, n38942, n38943, n38944, n38945, n38946,
         n38947, n38948, n38949, n38950, n38951, n38952, n38953, n38954,
         n38955, n38956, n38957, n38958, n38959, n38960, n38961, n38962,
         n38963, n38964, n38965, n38966, n38967, n38968, n38969, n38970,
         n38971, n38972, n38973, n38974, n38975, n38976, n38977, n38978,
         n38979, n38980, n38981, n38982, n38983, n38984, n38985, n38986,
         n38987, n38988, n38989, n38990, n38991, n38992, n38993, n38994,
         n38995, n38996, n38997, n38998, n38999, n39000, n39001, n39002,
         n39003, n39004, n39005, n39006, n39007, n39008, n39009, n39010,
         n39011, n39012, n39013, n39014, n39015, n39016, n39017, n39018,
         n39019, n39020, n39021, n39022, n39023, n39024, n39025, n39026,
         n39027, n39028, n39029, n39030, n39031, n39032, n39033, n39034,
         n39035, n39036, n39037, n39038, n39039, n39040, n39041, n39042,
         n39043, n39044, n39045, n39046, n39047, n39048, n39049, n39050,
         n39051, n39052, n39053, n39054, n39055, n39056, n39057, n39058,
         n39059, n39060, n39061, n39062, n39063, n39064, n39065, n39066,
         n39067, n39068, n39069, n39070, n39071, n39072, n39073, n39074,
         n39075, n39076, n39077, n39078, n39079, n39080, n39081, n39082,
         n39083, n39084, n39085, n39086, n39087, n39088, n39089, n39090,
         n39091, n39092, n39093, n39094, n39095, n39096, n39097, n39098,
         n39099, n39100, n39101, n39102, n39103, n39104, n39105, n39106,
         n39107, n39108, n39109, n39110, n39111, n39112, n39113, n39114,
         n39115, n39116, n39117, n39118, n39119, n39120, n39121, n39122,
         n39123, n39124, n39125, n39126, n39127, n39128, n39129, n39130,
         n39131, n39132, n39133, n39134, n39135, n39136, n39137, n39138,
         n39139, n39140, n39141, n39142, n39143, n39144, n39145, n39146,
         n39147, n39148, n39149, n39150, n39151, n39152, n39153, n39154,
         n39155, n39156, n39157, n39158, n39159, n39160, n39161, n39162,
         n39163, n39164, n39165, n39166, n39167, n39168, n39169, n39170,
         n39171, n39172, n39173, n39174, n39175, n39176, n39177, n39178,
         n39179, n39180, n39181, n39182, n39183, n39184, n39185, n39186,
         n39187, n39188, n39189, n39190, n39191, n39192, n39193, n39194,
         n39195, n39196, n39197, n39198, n39199, n39200, n39201, n39202,
         n39203, n39204, n39205, n39206, n39207, n39208, n39209, n39210,
         n39211, n39212, n39213, n39214, n39215, n39216, n39217, n39218,
         n39219, n39220, n39221, n39222, n39223, n39224, n39225, n39226,
         n39227, n39228, n39229, n39230, n39231, n39232, n39233, n39234,
         n39235, n39236, n39237, n39238, n39239, n39240, n39241, n39242,
         n39243, n39244, n39245, n39246, n39247, n39248, n39249, n39250,
         n39251, n39252, n39253, n39254, n39255, n39256, n39257, n39258,
         n39259, n39260, n39261, n39262, n39263, n39264, n39265, n39266,
         n39267, n39268, n39269, n39270, n39271, n39272, n39273, n39274,
         n39275, n39276, n39277, n39278, n39279, n39280, n39281, n39282,
         n39283, n39284, n39285, n39286, n39287, n39288, n39289, n39290,
         n39291, n39292, n39293, n39294, n39295, n39296, n39297, n39298,
         n39299, n39300, n39301, n39302, n39303, n39304, n39305, n39306,
         n39307, n39308, n39309, n39310, n39311, n39312, n39313, n39314,
         n39315, n39316, n39317, n39318, n39319, n39320, n39321, n39322,
         n39323, n39324, n39325, n39326, n39327, n39328, n39329, n39330,
         n39331, n39332, n39333, n39334, n39335, n39336, n39337, n39338,
         n39339, n39340, n39341, n39342, n39343, n39344, n39345, n39346,
         n39347, n39348, n39349, n39350, n39351, n39352, n39353, n39354,
         n39355, n39356, n39357, n39358, n39359, n39360, n39361, n39362,
         n39363, n39364, n39365, n39366, n39367, n39368, n39369, n39370,
         n39371, n39372, n39373, n39374, n39375, n39376, n39377, n39378,
         n39379, n39380, n39381, n39382, n39383, n39384, n39385, n39386,
         n39387, n39388, n39389, n39390, n39391, n39392, n39393, n39394,
         n39395, n39396, n39397, n39398, n39399, n39400, n39401, n39402,
         n39403, n39404, n39405, n39406, n39407, n39408, n39409, n39410,
         n39411, n39412, n39413, n39414, n39415, n39416, n39417, n39418,
         n39419, n39420, n39421, n39422, n39423, n39424, n39425, n39426,
         n39427, n39428, n39429, n39430, n39431, n39432, n39433, n39434,
         n39435, n39436, n39437, n39438, n39439, n39440, n39441, n39442,
         n39443, n39444, n39445, n39446, n39447, n39448, n39449, n39450,
         n39451, n39452, n39453, n39454, n39455, n39456, n39457, n39458,
         n39459, n39460, n39461, n39462, n39463, n39464, n39465, n39466,
         n39467, n39468, n39469, n39470, n39471, n39472, n39473, n39474,
         n39475, n39476, n39477, n39478, n39479, n39480, n39481, n39482,
         n39483, n39484, n39485, n39486, n39487, n39488, n39489, n39490,
         n39491, n39492, n39493, n39494, n39495, n39496, n39497, n39498,
         n39499, n39500, n39501, n39502, n39503, n39504, n39505, n39506,
         n39507, n39508, n39509, n39510, n39511, n39512, n39513, n39514,
         n39515, n39516, n39517, n39518, n39519, n39520, n39521, n39522,
         n39523, n39524, n39525, n39526, n39527, n39528, n39529, n39530,
         n39531, n39532, n39533, n39534, n39535, n39536, n39537, n39538,
         n39539, n39540, n39541, n39542, n39543, n39544, n39545, n39546,
         n39547, n39548, n39549, n39550, n39551, n39552, n39553, n39554,
         n39555, n39556, n39557, n39558, n39559, n39560, n39561, n39562,
         n39563, n39564, n39565, n39566, n39567, n39568, n39569, n39570,
         n39571, n39572, n39573, n39574, n39575, n39576, n39577, n39578,
         n39579, n39580, n39581, n39582, n39583, n39584, n39585, n39586,
         n39587, n39588, n39589, n39590, n39591, n39592, n39593, n39594,
         n39595, n39596, n39597, n39598, n39599, n39600, n39601, n39602,
         n39603, n39604, n39605, n39606, n39607, n39608, n39609, n39610,
         n39611, n39612, n39613, n39614, n39615, n39616, n39617, n39618,
         n39619, n39620, n39621, n39622, n39623, n39624, n39625, n39626,
         n39627, n39628, n39629, n39630, n39631, n39632, n39633, n39634,
         n39635, n39636, n39637, n39638, n39639, n39640, n39641, n39642,
         n39643, n39644, n39645, n39646, n39647, n39648, n39649, n39650,
         n39651, n39652, n39653, n39654, n39655, n39656, n39657, n39658,
         n39659, n39660, n39661, n39662, n39663, n39664, n39665, n39666,
         n39667, n39668, n39669, n39670, n39671, n39672, n39673, n39674,
         n39675, n39676, n39677, n39678, n39679, n39680, n39681, n39682,
         n39683, n39684, n39685, n39686, n39687, n39688, n39689, n39690,
         n39691, n39692, n39693, n39694, n39695, n39696, n39697, n39698,
         n39699, n39700, n39701, n39702, n39703, n39704, n39705, n39706,
         n39707, n39708, n39709, n39710, n39711, n39712, n39713, n39714,
         n39715, n39716, n39717, n39718, n39719, n39720, n39721, n39722,
         n39723, n39724, n39725, n39726, n39727, n39728, n39729, n39730,
         n39731, n39732, n39733, n39734, n39735, n39736, n39737, n39738,
         n39739, n39740, n39741, n39742, n39743, n39744, n39745, n39746,
         n39747, n39748, n39749, n39750, n39751, n39752, n39753, n39754,
         n39755, n39756, n39757, n39758, n39759, n39760, n39761, n39762,
         n39763, n39764, n39765, n39766, n39767, n39768, n39769, n39770,
         n39771, n39772, n39773, n39774, n39775, n39776, n39777, n39778,
         n39779, n39780, n39781, n39782, n39783, n39784, n39785, n39786,
         n39787, n39788, n39789, n39790, n39791, n39792, n39793, n39794,
         n39795, n39796, n39797, n39798, n39799, n39800, n39801, n39802,
         n39803, n39804, n39805, n39806, n39807, n39808, n39809, n39810,
         n39811, n39812, n39813, n39814, n39815, n39816, n39817, n39818,
         n39819, n39820, n39821, n39822, n39823, n39824, n39825, n39826,
         n39827, n39828, n39829, n39830, n39831, n39832, n39833, n39834,
         n39835, n39836, n39837, n39838, n39839, n39840, n39841, n39842,
         n39843, n39844, n39845, n39846, n39847, n39848, n39849, n39850,
         n39851, n39852, n39853, n39854, n39855, n39856, n39857, n39858,
         n39859, n39860, n39861, n39862, n39863, n39864, n39865, n39866,
         n39867, n39868, n39869, n39870, n39871, n39872, n39873, n39874,
         n39875, n39876, n39877, n39878, n39879, n39880, n39881, n39882,
         n39883, n39884, n39885, n39886, n39887, n39888, n39889, n39890,
         n39891, n39892, n39893, n39894, n39895, n39896, n39897, n39898,
         n39899, n39900, n39901, n39902, n39903, n39904, n39905, n39906,
         n39907, n39908, n39909, n39910, n39911, n39912, n39913, n39914,
         n39915, n39916, n39917, n39918, n39919, n39920, n39921, n39922,
         n39923, n39924, n39925, n39926, n39927, n39928, n39929, n39930,
         n39931, n39932, n39933, n39934, n39935, n39936, n39937, n39938,
         n39939, n39940, n39941, n39942, n39943, n39944, n39945, n39946,
         n39947, n39948, n39949, n39950, n39951, n39952, n39953, n39954,
         n39955, n39956, n39957, n39958, n39959, n39960, n39961, n39962,
         n39963, n39964, n39965, n39966, n39967, n39968, n39969, n39970,
         n39971, n39972, n39973, n39974, n39975, n39976, n39977, n39978,
         n39979, n39980, n39981, n39982, n39983, n39984, n39985, n39986,
         n39987, n39988, n39989, n39990, n39991, n39992, n39993, n39994,
         n39995, n39996, n39997, n39998, n39999, n40000, n40001, n40002,
         n40003, n40004, n40005, n40006, n40007, n40008, n40009, n40010,
         n40011, n40012, n40013, n40014, n40015, n40016, n40017, n40018,
         n40019, n40020, n40021, n40022, n40023, n40024, n40025, n40026,
         n40027, n40028, n40029, n40030, n40031, n40032, n40033, n40034,
         n40035, n40036, n40037, n40038, n40039, n40040, n40041, n40042,
         n40043, n40044, n40045, n40046, n40047, n40048, n40049, n40050,
         n40051, n40052, n40053, n40054, n40055, n40056, n40057, n40058,
         n40059, n40060, n40061, n40062, n40063, n40064, n40065, n40066,
         n40067, n40068, n40069, n40070, n40071, n40072, n40073, n40074,
         n40075, n40076, n40077, n40078, n40079, n40080, n40081, n40082,
         n40083, n40084, n40085, n40086, n40087, n40088, n40089, n40090,
         n40091, n40092, n40093, n40094, n40095, n40096, n40097, n40098,
         n40099, n40100, n40101, n40102, n40103, n40104, n40105, n40106,
         n40107, n40108, n40109, n40110, n40111, n40112, n40113, n40114,
         n40115, n40116, n40117, n40118, n40119, n40120, n40121, n40122,
         n40123, n40124, n40125, n40126, n40127, n40128, n40129, n40130,
         n40131, n40132, n40133, n40134, n40135, n40136, n40137, n40138,
         n40139, n40140, n40141, n40142, n40143, n40144, n40145, n40146,
         n40147, n40148, n40149, n40150, n40151, n40152, n40153, n40154,
         n40155, n40156, n40157, n40158, n40159, n40160, n40161, n40162,
         n40163, n40164, n40165, n40166, n40167, n40168, n40169, n40170,
         n40171, n40172, n40173, n40174, n40175, n40176, n40177, n40178,
         n40179, n40180, n40181, n40182, n40183, n40184, n40185, n40186,
         n40187, n40188, n40189, n40190, n40191, n40192, n40193, n40194,
         n40195, n40196, n40197, n40198, n40199, n40200, n40201, n40202,
         n40203, n40204, n40205, n40206, n40207, n40208, n40209, n40210,
         n40211, n40212, n40213, n40214, n40215, n40216, n40217, n40218,
         n40219, n40220, n40221, n40222, n40223, n40224, n40225, n40226,
         n40227, n40228, n40229, n40230, n40231, n40232, n40233, n40234,
         n40235, n40236, n40237, n40238, n40239, n40240, n40241, n40242,
         n40243, n40244, n40245, n40246, n40247, n40248, n40249, n40250,
         n40251, n40252, n40253, n40254, n40255, n40256, n40257, n40258,
         n40259, n40260, n40261, n40262, n40263, n40264, n40265, n40266,
         n40267, n40268, n40269, n40270, n40271, n40272, n40273, n40274,
         n40275, n40276, n40277, n40278, n40279, n40280, n40281, n40282,
         n40283, n40284, n40285, n40286, n40287, n40288, n40289, n40290,
         n40291, n40292, n40293, n40294, n40295, n40296, n40297, n40298,
         n40299, n40300, n40301, n40302, n40303, n40304, n40305, n40306,
         n40307, n40308, n40309, n40310, n40311, n40312, n40313, n40314,
         n40315, n40316, n40317, n40318, n40319, n40320, n40321, n40322,
         n40323, n40324, n40325, n40326, n40327, n40328, n40329, n40330,
         n40331, n40332, n40333, n40334, n40335, n40336, n40337, n40338,
         n40339, n40340, n40341, n40342, n40343, n40344, n40345, n40346,
         n40347, n40348, n40349, n40350, n40351, n40352, n40353, n40354,
         n40355, n40356, n40357, n40358, n40359, n40360, n40361, n40362,
         n40363, n40364, n40365, n40366, n40367, n40368, n40369, n40370,
         n40371, n40372, n40373, n40374, n40375, n40376, n40377, n40378,
         n40379, n40380, n40381, n40382, n40383, n40384, n40385, n40386,
         n40387, n40388, n40389, n40390, n40391, n40392, n40393, n40394,
         n40395, n40396, n40397, n40398, n40399, n40400, n40401, n40402,
         n40403, n40404, n40405, n40406, n40407, n40408, n40409, n40410,
         n40411, n40412, n40413, n40414, n40415, n40416, n40417, n40418,
         n40419, n40420, n40421, n40422, n40423, n40424, n40425, n40426,
         n40427, n40428, n40429, n40430, n40431, n40432, n40433, n40434,
         n40435, n40436, n40437, n40438, n40439, n40440, n40441, n40442,
         n40443, n40444, n40445, n40446, n40447, n40448, n40449, n40450,
         n40451, n40452, n40453, n40454, n40455, n40456, n40457, n40458,
         n40459, n40460, n40461, n40462, n40463, n40464, n40465, n40466,
         n40467, n40468, n40469, n40470, n40471, n40472, n40473, n40474,
         n40475, n40476, n40477, n40478, n40479, n40480, n40481, n40482,
         n40483, n40484, n40485, n40486, n40487, n40488, n40489, n40490,
         n40491, n40492, n40493, n40494, n40495, n40496, n40497, n40498,
         n40499, n40500, n40501, n40502, n40503, n40504, n40505, n40506,
         n40507, n40508, n40509, n40510, n40511, n40512, n40513, n40514,
         n40515, n40516, n40517, n40518, n40519, n40520, n40521, n40522,
         n40523, n40524, n40525, n40526, n40527, n40528, n40529, n40530,
         n40531, n40532, n40533, n40534, n40535, n40536, n40537, n40538,
         n40539, n40540, n40541, n40542, n40543, n40544, n40545, n40546,
         n40547, n40548, n40549, n40550, n40551, n40552, n40553, n40554,
         n40555, n40556, n40557, n40558, n40559, n40560, n40561, n40562,
         n40563, n40564, n40565, n40566, n40567, n40568, n40569, n40570,
         n40571, n40572, n40573, n40574, n40575, n40576, n40577, n40578,
         n40579, n40580, n40581, n40582, n40583, n40584, n40585, n40586,
         n40587, n40588, n40589, n40590, n40591, n40592, n40593, n40594,
         n40595, n40596, n40597, n40598, n40599, n40600, n40601, n40602,
         n40603, n40604, n40605, n40606, n40607, n40608, n40609, n40610,
         n40611, n40612, n40613, n40614, n40615, n40616, n40617, n40618,
         n40619, n40620, n40621, n40622, n40623, n40624, n40625, n40626,
         n40627, n40628, n40629, n40630, n40631, n40632, n40633, n40634,
         n40635, n40636, n40637, n40638, n40639, n40640, n40641, n40642,
         n40643, n40644, n40645, n40646, n40647, n40648, n40649, n40650,
         n40651, n40652, n40653, n40654, n40655, n40656, n40657, n40658,
         n40659, n40660, n40661, n40662, n40663, n40664, n40665, n40666,
         n40667, n40668, n40669, n40670, n40671, n40672, n40673, n40674,
         n40675, n40676, n40677, n40678, n40679, n40680, n40681, n40682,
         n40683, n40684, n40685, n40686, n40687, n40688, n40689, n40690,
         n40691, n40692, n40693, n40694, n40695, n40696, n40697, n40698,
         n40699, n40700, n40701, n40702, n40703, n40704, n40705, n40706,
         n40707, n40708, n40709, n40710, n40711, n40712, n40713, n40714,
         n40715, n40716, n40717, n40718, n40719, n40720, n40721, n40722,
         n40723, n40724, n40725, n40726, n40727, n40728, n40729, n40730,
         n40731, n40732, n40733, n40734, n40735, n40736, n40737, n40738,
         n40739, n40740, n40741, n40742, n40743, n40744, n40745, n40746,
         n40747, n40748, n40749, n40750, n40751, n40752, n40753, n40754,
         n40755, n40756, n40757, n40758, n40759, n40760, n40761, n40762,
         n40763, n40764, n40765, n40766, n40767, n40768, n40769, n40770,
         n40771, n40772, n40773, n40774, n40775, n40776, n40777, n40778,
         n40779, n40780, n40781, n40782, n40783, n40784, n40785, n40786,
         n40787, n40788, n40789, n40790, n40791, n40792, n40793, n40794,
         n40795, n40796, n40797, n40798, n40799, n40800, n40801, n40802,
         n40803, n40804, n40805, n40806, n40807, n40808, n40809, n40810,
         n40811, n40812, n40813, n40814, n40815, n40816, n40817, n40818,
         n40819, n40820, n40821, n40822, n40823, n40824, n40825, n40826,
         n40827, n40828, n40829, n40830, n40831, n40832, n40833, n40834,
         n40835, n40836, n40837, n40838, n40839, n40840, n40841, n40842,
         n40843, n40844, n40845, n40846, n40847, n40848, n40849, n40850,
         n40851, n40852, n40853, n40854, n40855, n40856, n40857, n40858,
         n40859, n40860, n40861, n40862, n40863, n40864, n40865, n40866,
         n40867, n40868, n40869, n40870, n40871, n40872, n40873, n40874,
         n40875, n40876, n40877, n40878, n40879, n40880, n40881, n40882,
         n40883, n40884, n40885, n40886, n40887, n40888, n40889, n40890,
         n40891, n40892, n40893, n40894, n40895, n40896, n40897, n40898,
         n40899, n40900, n40901, n40902, n40903, n40904, n40905, n40906,
         n40907, n40908, n40909, n40910, n40911, n40912, n40913, n40914,
         n40915, n40916, n40917, n40918, n40919, n40920, n40921, n40922,
         n40923, n40924, n40925, n40926, n40927, n40928, n40929, n40930,
         n40931, n40932, n40933, n40934, n40935, n40936, n40937, n40938,
         n40939, n40940, n40941, n40942, n40943, n40944, n40945, n40946,
         n40947, n40948, n40949, n40950, n40951, n40952, n40953, n40954,
         n40955, n40956, n40957, n40958, n40959, n40960, n40961, n40962,
         n40963, n40964, n40965, n40966, n40967, n40968, n40969, n40970,
         n40971, n40972, n40973, n40974, n40975, n40976, n40977, n40978,
         n40979, n40980, n40981, n40982, n40983, n40984, n40985, n40986,
         n40987, n40988, n40989, n40990, n40991, n40992, n40993, n40994,
         n40995, n40996, n40997, n40998, n40999, n41000, n41001, n41002,
         n41003, n41004, n41005, n41006, n41007, n41008, n41009, n41010,
         n41011, n41012, n41013, n41014, n41015, n41016, n41017, n41018,
         n41019, n41020, n41021, n41022, n41023, n41024, n41025, n41026,
         n41027, n41028, n41029, n41030, n41031, n41032, n41033, n41034,
         n41035, n41036, n41037, n41038, n41039, n41040, n41041, n41042,
         n41043, n41044, n41045, n41046, n41047, n41048, n41049, n41050,
         n41051, n41052, n41053, n41054, n41055, n41056, n41057, n41058,
         n41059, n41060, n41061, n41062, n41063, n41064, n41065, n41066,
         n41067, n41068, n41069, n41070, n41071, n41072, n41073, n41074,
         n41075, n41076, n41077, n41078, n41079, n41080, n41081, n41082,
         n41083, n41084, n41085, n41086, n41087, n41088, n41089, n41090,
         n41091, n41092, n41093, n41094, n41095, n41096, n41097, n41098,
         n41099, n41100, n41101, n41102, n41103, n41104, n41105, n41106,
         n41107, n41108, n41109, n41110, n41111, n41112, n41113, n41114,
         n41115, n41116, n41117, n41118, n41119, n41120, n41121, n41122,
         n41123, n41124, n41125, n41126, n41127, n41128, n41129, n41130,
         n41131, n41132, n41133, n41134, n41135, n41136, n41137, n41138,
         n41139, n41140, n41141, n41142, n41143, n41144, n41145, n41146,
         n41147, n41148, n41149, n41150, n41151, n41152, n41153, n41154,
         n41155, n41156, n41157, n41158, n41159, n41160, n41161, n41162,
         n41163, n41164, n41165, n41166, n41167, n41168, n41169, n41170,
         n41171, n41172, n41173, n41174, n41175, n41176, n41177, n41178,
         n41179, n41180, n41181, n41182, n41183, n41184, n41185, n41186,
         n41187, n41188, n41189, n41190, n41191, n41192, n41193, n41194,
         n41195, n41196, n41197, n41198, n41199, n41200, n41201, n41202,
         n41203, n41204, n41205, n41206, n41207, n41208, n41209, n41210,
         n41211, n41212, n41213, n41214, n41215, n41216, n41217, n41218,
         n41219, n41220, n41221, n41222, n41223, n41224, n41225, n41226,
         n41227, n41228, n41229, n41230, n41231, n41232, n41233, n41234,
         n41235, n41236, n41237, n41238, n41239, n41240, n41241, n41242,
         n41243, n41244, n41245, n41246, n41247, n41248, n41249, n41250,
         n41251, n41252, n41253, n41254, n41255, n41256, n41257, n41258,
         n41259, n41260, n41261, n41262, n41263, n41264, n41265, n41266,
         n41267, n41268, n41269, n41270, n41271, n41272, n41273, n41274,
         n41275, n41276, n41277, n41278, n41279, n41280, n41281, n41282,
         n41283, n41284, n41285, n41286, n41287, n41288, n41289, n41290,
         n41291, n41292, n41293, n41294, n41295, n41296, n41297, n41298,
         n41299, n41300, n41301, n41302, n41303, n41304, n41305, n41306,
         n41307, n41308, n41309, n41310, n41311, n41312, n41313, n41314,
         n41315, n41316, n41317, n41318, n41319, n41320, n41321, n41322,
         n41323, n41324, n41325, n41326, n41327, n41328, n41329, n41330,
         n41331, n41332, n41333, n41334, n41335, n41336, n41337, n41338,
         n41339, n41340, n41341, n41342, n41343, n41344, n41345, n41346,
         n41347, n41348, n41349, n41350, n41351, n41352, n41353, n41354,
         n41355, n41356, n41357, n41358, n41359, n41360, n41361, n41362,
         n41363, n41364, n41365, n41366, n41367, n41368, n41369, n41370,
         n41371, n41372, n41373, n41374, n41375, n41376, n41377, n41378,
         n41379, n41380, n41381, n41382, n41383, n41384, n41385, n41386,
         n41387, n41388, n41389, n41390, n41391, n41392, n41393, n41394,
         n41395, n41396, n41397, n41398, n41399, n41400, n41401, n41402,
         n41403, n41404, n41405, n41406, n41407, n41408, n41409, n41410,
         n41411, n41412, n41413, n41414, n41415, n41416, n41417, n41418,
         n41419, n41420, n41421, n41422, n41423, n41424, n41425, n41426,
         n41427, n41428, n41429, n41430, n41431, n41432, n41433, n41434,
         n41435, n41436, n41437, n41438, n41439, n41440, n41441, n41442,
         n41443, n41444, n41445, n41446, n41447, n41448, n41449, n41450,
         n41451, n41452, n41453, n41454, n41455, n41456, n41457, n41458,
         n41459, n41460, n41461, n41462, n41463, n41464, n41465, n41466,
         n41467, n41468, n41469, n41470, n41471, n41472, n41473, n41474,
         n41475, n41476, n41477, n41478, n41479, n41480, n41481, n41482,
         n41483, n41484, n41485, n41486, n41487, n41488, n41489, n41490,
         n41491, n41492, n41493, n41494, n41495, n41496, n41497, n41498,
         n41499, n41500, n41501, n41502, n41503, n41504, n41505, n41506,
         n41507, n41508, n41509, n41510, n41511, n41512, n41513, n41514,
         n41515, n41516, n41517, n41518, n41519, n41520, n41521, n41522,
         n41523, n41524, n41525, n41526, n41527, n41528, n41529, n41530,
         n41531, n41532, n41533, n41534, n41535, n41536, n41537, n41538,
         n41539, n41540, n41541, n41542, n41543, n41544, n41545, n41546,
         n41547, n41548, n41549, n41550, n41551, n41552, n41553, n41554,
         n41555, n41556, n41557, n41558, n41559, n41560, n41561, n41562,
         n41563, n41564, n41565, n41566, n41567, n41568, n41569, n41570,
         n41571, n41572, n41573, n41574, n41575, n41576, n41577, n41578,
         n41579, n41580, n41581, n41582, n41583, n41584, n41585, n41586,
         n41587, n41588, n41589, n41590, n41591, n41592, n41593, n41594,
         n41595, n41596, n41597, n41598, n41599, n41600, n41601, n41602,
         n41603, n41604, n41605, n41606, n41607, n41608, n41609, n41610,
         n41611, n41612, n41613, n41614, n41615, n41616, n41617, n41618,
         n41619, n41620, n41621, n41622, n41623, n41624, n41625, n41626,
         n41627, n41628, n41629, n41630, n41631, n41632, n41633, n41634,
         n41635, n41636, n41637, n41638, n41639, n41640, n41641, n41642,
         n41643, n41644, n41645, n41646, n41647, n41648, n41649, n41650,
         n41651, n41652, n41653, n41654, n41655, n41656, n41657, n41658,
         n41659, n41660, n41661, n41662, n41663, n41664, n41665, n41666,
         n41667, n41668, n41669, n41670, n41671, n41672, n41673, n41674,
         n41675, n41676, n41677, n41678, n41679, n41680, n41681, n41682,
         n41683, n41684, n41685, n41686, n41687, n41688, n41689, n41690,
         n41691, n41692, n41693, n41694, n41695, n41696, n41697, n41698,
         n41699, n41700, n41701, n41702, n41703, n41704, n41705, n41706,
         n41707, n41708, n41709, n41710, n41711, n41712, n41713, n41714,
         n41715, n41716, n41717, n41718, n41719, n41720, n41721, n41722,
         n41723, n41724, n41725, n41726, n41727, n41728, n41729, n41730,
         n41731, n41732, n41733, n41734, n41735, n41736, n41737, n41738,
         n41739, n41740, n41741, n41742, n41743, n41744, n41745, n41746,
         n41747, n41748, n41749, n41750, n41751, n41752, n41753, n41754,
         n41755, n41756, n41757, n41758, n41759, n41760, n41761, n41762,
         n41763, n41764, n41765, n41766, n41767, n41768, n41769, n41770,
         n41771, n41772, n41773, n41774, n41775, n41776, n41777, n41778,
         n41779, n41780, n41781, n41782, n41783, n41784, n41785, n41786,
         n41787, n41788, n41789, n41790, n41791, n41792, n41793, n41794,
         n41795, n41796, n41797, n41798, n41799, n41800, n41801, n41802,
         n41803, n41804, n41805, n41806, n41807, n41808, n41809, n41810,
         n41811, n41812, n41813, n41814, n41815, n41816, n41817, n41818,
         n41819, n41820, n41821, n41822, n41823, n41824, n41825, n41826,
         n41827, n41828, n41829, n41830, n41831, n41832, n41833, n41834,
         n41835, n41836, n41837, n41838, n41839, n41840, n41841, n41842,
         n41843, n41844, n41845, n41846, n41847, n41848, n41849, n41850,
         n41851, n41852, n41853, n41854, n41855, n41856, n41857, n41858,
         n41859, n41860, n41861, n41862, n41863, n41864, n41865, n41866,
         n41867, n41868, n41869, n41870, n41871, n41872, n41873, n41874,
         n41875, n41876, n41877, n41878, n41879, n41880, n41881, n41882,
         n41883, n41884, n41885, n41886, n41887, n41888, n41889, n41890,
         n41891, n41892, n41893, n41894, n41895, n41896, n41897, n41898,
         n41899, n41900, n41901, n41902, n41903, n41904, n41905, n41906,
         n41907, n41908, n41909, n41910, n41911, n41912, n41913, n41914,
         n41915, n41916, n41917, n41918, n41919, n41920, n41921, n41922,
         n41923, n41924, n41925, n41926, n41927, n41928, n41929, n41930,
         n41931, n41932, n41933, n41934, n41935, n41936, n41937, n41938,
         n41939, n41940, n41941, n41942, n41943, n41944, n41945, n41946,
         n41947, n41948, n41949, n41950, n41951, n41952, n41953, n41954,
         n41955, n41956, n41957, n41958, n41959, n41960, n41961, n41962,
         n41963, n41964, n41965, n41966, n41967, n41968, n41969, n41970,
         n41971, n41972, n41973, n41974, n41975, n41976, n41977, n41978,
         n41979, n41980, n41981, n41982, n41983, n41984, n41985, n41986,
         n41987, n41988, n41989, n41990, n41991, n41992, n41993, n41994,
         n41995, n41996, n41997, n41998, n41999, n42000, n42001, n42002,
         n42003, n42004, n42005, n42006, n42007, n42008, n42009, n42010,
         n42011, n42012, n42013, n42014, n42015, n42016, n42017, n42018,
         n42019, n42020, n42021, n42022, n42023, n42024, n42025, n42026,
         n42027, n42028, n42029, n42030, n42031, n42032, n42033, n42034,
         n42035, n42036, n42037, n42038, n42039, n42040, n42041, n42042,
         n42043, n42044, n42045, n42046, n42047, n42048, n42049, n42050,
         n42051, n42052, n42053, n42054, n42055, n42056, n42057, n42058,
         n42059, n42060, n42061, n42062, n42063, n42064, n42065, n42066,
         n42067, n42068, n42069, n42070, n42071, n42072, n42073, n42074,
         n42075, n42076, n42077, n42078, n42079, n42080, n42081, n42082,
         n42083, n42084, n42085, n42086, n42087, n42088, n42089, n42090,
         n42091, n42092, n42093, n42094, n42095, n42096, n42097, n42098,
         n42099, n42100, n42101, n42102, n42103, n42104, n42105, n42106,
         n42107, n42108, n42109, n42110, n42111, n42112, n42113, n42114,
         n42115, n42116, n42117, n42118, n42119, n42120, n42121, n42122,
         n42123, n42124, n42125, n42126, n42127, n42128, n42129, n42130,
         n42131, n42132, n42133, n42134, n42135, n42136, n42137, n42138,
         n42139, n42140, n42141, n42142, n42143, n42144, n42145, n42146,
         n42147, n42148, n42149, n42150, n42151, n42152, n42153, n42154,
         n42155, n42156, n42157, n42158, n42159, n42160, n42161, n42162,
         n42163, n42164, n42165, n42166, n42167, n42168, n42169, n42170,
         n42171, n42172, n42173, n42174, n42175, n42176, n42177, n42178,
         n42179, n42180, n42181, n42182, n42183, n42184, n42185, n42186,
         n42187, n42188, n42189, n42190, n42191, n42192, n42193, n42194,
         n42195, n42196, n42197, n42198, n42199, n42200, n42201, n42202,
         n42203, n42204, n42205, n42206, n42207, n42208, n42209, n42210,
         n42211, n42212, n42213, n42214, n42215, n42216, n42217, n42218,
         n42219, n42220, n42221, n42222, n42223, n42224, n42225, n42226,
         n42227, n42228, n42229, n42230, n42231, n42232, n42233, n42234,
         n42235, n42236, n42237, n42238, n42239, n42240, n42241, n42242,
         n42243, n42244, n42245, n42246, n42247, n42248, n42249, n42250,
         n42251, n42252, n42253, n42254, n42255, n42256, n42257, n42258,
         n42259, n42260, n42261, n42262, n42263, n42264, n42265, n42266,
         n42267, n42268, n42269, n42270, n42271, n42272, n42273, n42274,
         n42275, n42276, n42277, n42278, n42279, n42280, n42281, n42282,
         n42283, n42284, n42285, n42286, n42287, n42288, n42289, n42290,
         n42291, n42292, n42293, n42294, n42295, n42296, n42297, n42298,
         n42299, n42300, n42301, n42302, n42303, n42304, n42305, n42306,
         n42307, n42308, n42309, n42310, n42311, n42312, n42313, n42314,
         n42315, n42316, n42317, n42318, n42319, n42320, n42321, n42322,
         n42323, n42324, n42325, n42326, n42327, n42328, n42329, n42330,
         n42331, n42332, n42333, n42334, n42335, n42336, n42337, n42338,
         n42339, n42340, n42341, n42342, n42343, n42344, n42345, n42346,
         n42347, n42348, n42349, n42350, n42351, n42352, n42353, n42354,
         n42355, n42356, n42357, n42358, n42359, n42360, n42361, n42362,
         n42363, n42364, n42365, n42366, n42367, n42368, n42369, n42370,
         n42371, n42372, n42373, n42374, n42375, n42376, n42377, n42378,
         n42379, n42380, n42381, n42382, n42383, n42384, n42385, n42386,
         n42387, n42388, n42389, n42390, n42391, n42392, n42393, n42394,
         n42395, n42396, n42397, n42398, n42399, n42400, n42401, n42402,
         n42403, n42404, n42405, n42406, n42407, n42408, n42409, n42410,
         n42411, n42412, n42413, n42414, n42415, n42416, n42417, n42418,
         n42419, n42420, n42421, n42422, n42423, n42424, n42425, n42426,
         n42427, n42428, n42429, n42430, n42431, n42432, n42433, n42434,
         n42435, n42436, n42437, n42438, n42439, n42440, n42441, n42442,
         n42443, n42444, n42445, n42446, n42447, n42448, n42449, n42450,
         n42451, n42452, n42453, n42454, n42455, n42456, n42457, n42458,
         n42459, n42460, n42461, n42462, n42463, n42464, n42465, n42466,
         n42467, n42468, n42469, n42470, n42471, n42472, n42473, n42474,
         n42475, n42476, n42477, n42478, n42479, n42480, n42481, n42482,
         n42483, n42484, n42485, n42486, n42487, n42488, n42489, n42490,
         n42491, n42492, n42493, n42494, n42495, n42496, n42497, n42498,
         n42499, n42500, n42501, n42502, n42503, n42504, n42505, n42506,
         n42507, n42508, n42509, n42510, n42511, n42512, n42513, n42514,
         n42515, n42516, n42517, n42518, n42519, n42520, n42521, n42522,
         n42523, n42524, n42525, n42526, n42527, n42528, n42529, n42530,
         n42531, n42532, n42533, n42534, n42535, n42536, n42537, n42538,
         n42539, n42540, n42541, n42542, n42543, n42544, n42545, n42546,
         n42547, n42548, n42549, n42550, n42551, n42552, n42553, n42554,
         n42555, n42556, n42557, n42558, n42559, n42560, n42561, n42562,
         n42563, n42564, n42565, n42566, n42567, n42568, n42569, n42570,
         n42571, n42572, n42573, n42574, n42575, n42576, n42577, n42578,
         n42579, n42580, n42581, n42582, n42583, n42584, n42585, n42586,
         n42587, n42588, n42589, n42590, n42591, n42592, n42593, n42594,
         n42595, n42596, n42597, n42598, n42599, n42600, n42601, n42602,
         n42603, n42604, n42605, n42606, n42607, n42608, n42609, n42610,
         n42611, n42612, n42613, n42614, n42615, n42616, n42617, n42618,
         n42619, n42620, n42621, n42622, n42623, n42624, n42625, n42626,
         n42627, n42628, n42629, n42630, n42631, n42632, n42633, n42634,
         n42635, n42636, n42637, n42638, n42639, n42640, n42641, n42642,
         n42643, n42644, n42645, n42646, n42647, n42648, n42649, n42650,
         n42651, n42652, n42653, n42654, n42655, n42656, n42657, n42658,
         n42659, n42660, n42661, n42662, n42663, n42664, n42665, n42666,
         n42667, n42668, n42669, n42670, n42671, n42672, n42673, n42674,
         n42675, n42676, n42677, n42678, n42679, n42680, n42681, n42682,
         n42683, n42684, n42685, n42686, n42687, n42688, n42689, n42690,
         n42691, n42692, n42693, n42694, n42695, n42696, n42697, n42698,
         n42699, n42700, n42701, n42702, n42703, n42704, n42705, n42706,
         n42707, n42708, n42709, n42710, n42711, n42712, n42713, n42714,
         n42715, n42716, n42717, n42718, n42719, n42720, n42721, n42722,
         n42723, n42724, n42725, n42726, n42727, n42728, n42729, n42730,
         n42731, n42732, n42733, n42734, n42735, n42736, n42737, n42738,
         n42739, n42740, n42741, n42742, n42743, n42744, n42745, n42746,
         n42747, n42748, n42749, n42750, n42751, n42752, n42753, n42754,
         n42755, n42756, n42757, n42758, n42759, n42760, n42761, n42762,
         n42763, n42764, n42765, n42766, n42767, n42768, n42769, n42770,
         n42771, n42772, n42773, n42774, n42775, n42776, n42777, n42778,
         n42779, n42780, n42781, n42782, n42783, n42784, n42785, n42786,
         n42787, n42788, n42789, n42790, n42791, n42792, n42793, n42794,
         n42795, n42796, n42797, n42798, n42799, n42800, n42801, n42802,
         n42803, n42804, n42805, n42806, n42807, n42808, n42809, n42810,
         n42811, n42812, n42813, n42814, n42815, n42816, n42817, n42818,
         n42819, n42820, n42821, n42822, n42823, n42824, n42825, n42826,
         n42827, n42828, n42829, n42830, n42831, n42832, n42833, n42834,
         n42835, n42836, n42837, n42838, n42839, n42840, n42841, n42842,
         n42843, n42844, n42845, n42846, n42847, n42848, n42849, n42850,
         n42851, n42852, n42853, n42854, n42855, n42856, n42857, n42858,
         n42859, n42860, n42861, n42862, n42863, n42864, n42865, n42866,
         n42867, n42868, n42869, n42870, n42871, n42872, n42873, n42874,
         n42875, n42876, n42877, n42878, n42879, n42880, n42881, n42882,
         n42883, n42884, n42885, n42886, n42887, n42888, n42889, n42890,
         n42891, n42892, n42893, n42894, n42895, n42896, n42897, n42898,
         n42899, n42900, n42901, n42902, n42903, n42904, n42905, n42906,
         n42907, n42908, n42909, n42910, n42911, n42912, n42913, n42914,
         n42915, n42916, n42917, n42918, n42919, n42920, n42921, n42922,
         n42923, n42924, n42925, n42926, n42927, n42928, n42929, n42930,
         n42931, n42932, n42933, n42934, n42935, n42936, n42937, n42938,
         n42939, n42940, n42941, n42942, n42943, n42944, n42945, n42946,
         n42947, n42948, n42949, n42950, n42951, n42952, n42953, n42954,
         n42955, n42956, n42957, n42958, n42959, n42960, n42961, n42962,
         n42963, n42964, n42965, n42966, n42967, n42968, n42969, n42970,
         n42971, n42972, n42973, n42974, n42975, n42976, n42977, n42978,
         n42979, n42980, n42981, n42982, n42983, n42984, n42985, n42986,
         n42987, n42988, n42989, n42990, n42991, n42992, n42993, n42994,
         n42995, n42996, n42997, n42998, n42999, n43000, n43001, n43002,
         n43003, n43004, n43005, n43006, n43007, n43008, n43009, n43010,
         n43011, n43012, n43013, n43014, n43015, n43016, n43017, n43018,
         n43019, n43020, n43021, n43022, n43023, n43024, n43025, n43026,
         n43027, n43028, n43029, n43030, n43031, n43032, n43033, n43034,
         n43035, n43036, n43037, n43038, n43039, n43040, n43041, n43042,
         n43043, n43044, n43045, n43046, n43047, n43048, n43049, n43050,
         n43051, n43052, n43053, n43054, n43055, n43056, n43057, n43058,
         n43059, n43060, n43061, n43062, n43063, n43064, n43065, n43066,
         n43067, n43068, n43069, n43070, n43071, n43072, n43073, n43074,
         n43075, n43076, n43077, n43078, n43079, n43080, n43081, n43082,
         n43083, n43084, n43085, n43086, n43087, n43088, n43089, n43090,
         n43091, n43092, n43093, n43094, n43095, n43096, n43097, n43098,
         n43099, n43100, n43101, n43102, n43103, n43104, n43105, n43106,
         n43107, n43108, n43109, n43110, n43111, n43112, n43113, n43114,
         n43115, n43116, n43117, n43118, n43119, n43120, n43121, n43122,
         n43123, n43124, n43125, n43126, n43127, n43128, n43129, n43130,
         n43131, n43132, n43133, n43134, n43135, n43136, n43137, n43138,
         n43139, n43140, n43141, n43142, n43143, n43144, n43145, n43146,
         n43147, n43148, n43149, n43150, n43151, n43152, n43153, n43154,
         n43155, n43156, n43157, n43158, n43159, n43160, n43161, n43162,
         n43163, n43164, n43165, n43166, n43167, n43168, n43169, n43170,
         n43171, n43172, n43173, n43174, n43175, n43176, n43177, n43178,
         n43179, n43180, n43181, n43182, n43183, n43184, n43185, n43186,
         n43187, n43188, n43189, n43190, n43191, n43192, n43193, n43194,
         n43195, n43196, n43197, n43198, n43199, n43200, n43201, n43202,
         n43203, n43204, n43205, n43206, n43207, n43208, n43209, n43210,
         n43211, n43212, n43213, n43214, n43215, n43216, n43217, n43218,
         n43219, n43220, n43221, n43222, n43223, n43224, n43225, n43226,
         n43227, n43228, n43229, n43230, n43231, n43232, n43233, n43234,
         n43235, n43236, n43237, n43238, n43239, n43240, n43241, n43242,
         n43243, n43244, n43245, n43246, n43247, n43248, n43249, n43250,
         n43251, n43252, n43253, n43254, n43255, n43256, n43257, n43258,
         n43259, n43260, n43261, n43262, n43263, n43264, n43265, n43266,
         n43267, n43268, n43269, n43270, n43271, n43272, n43273, n43274,
         n43275, n43276, n43277, n43278, n43279, n43280, n43281, n43282,
         n43283, n43284, n43285, n43286, n43287, n43288, n43289, n43290,
         n43291, n43292, n43293, n43294, n43295, n43296, n43297, n43298,
         n43299, n43300, n43301, n43302, n43303, n43304, n43305, n43306,
         n43307, n43308, n43309, n43310, n43311, n43312, n43313, n43314,
         n43315, n43316, n43317, n43318, n43319, n43320, n43321, n43322,
         n43323, n43324, n43325, n43326, n43327, n43328, n43329, n43330,
         n43331, n43332, n43333, n43334, n43335, n43336, n43337, n43338,
         n43339, n43340, n43341, n43342, n43343, n43344, n43345, n43346,
         n43347, n43348, n43349, n43350, n43351, n43352, n43353, n43354,
         n43355, n43356, n43357, n43358, n43359, n43360, n43361, n43362,
         n43363, n43364, n43365, n43366, n43367, n43368, n43369, n43370,
         n43371, n43372, n43373, n43374, n43375, n43376, n43377, n43378,
         n43379, n43380, n43381, n43382, n43383, n43384, n43385, n43386,
         n43387, n43388, n43389, n43390, n43391, n43392, n43393, n43394,
         n43395, n43396, n43397, n43398, n43399, n43400, n43401, n43402,
         n43403, n43404, n43405, n43406, n43407, n43408, n43409, n43410,
         n43411, n43412, n43413, n43414, n43415, n43416, n43417, n43418,
         n43419, n43420, n43421, n43422, n43423, n43424, n43425, n43426,
         n43427, n43428, n43429, n43430, n43431, n43432, n43433, n43434,
         n43435, n43436, n43437, n43438, n43439, n43440, n43441, n43442,
         n43443, n43444, n43445, n43446, n43447, n43448, n43449, n43450,
         n43451, n43452, n43453, n43454, n43455, n43456, n43457, n43458,
         n43459, n43460, n43461, n43462, n43463, n43464, n43465, n43466,
         n43467, n43468, n43469, n43470, n43471, n43472, n43473, n43474,
         n43475, n43476, n43477, n43478, n43479, n43480, n43481, n43482,
         n43483, n43484, n43485, n43486, n43487, n43488, n43489, n43490,
         n43491, n43492, n43493, n43494, n43495, n43496, n43497, n43498,
         n43499, n43500, n43501, n43502, n43503, n43504, n43505, n43506,
         n43507, n43508, n43509, n43510, n43511, n43512, n43513, n43514,
         n43515, n43516, n43517, n43518, n43519, n43520, n43521, n43522,
         n43523, n43524, n43525, n43526, n43527, n43528, n43529, n43530,
         n43531, n43532, n43533, n43534, n43535, n43536, n43537, n43538,
         n43539, n43540, n43541, n43542, n43543, n43544, n43545, n43546,
         n43547, n43548, n43549, n43550, n43551, n43552, n43553, n43554,
         n43555, n43556, n43557, n43558, n43559, n43560, n43561, n43562,
         n43563, n43564, n43565, n43566, n43567, n43568, n43569, n43570,
         n43571, n43572, n43573, n43574, n43575, n43576, n43577, n43578,
         n43579, n43580, n43581, n43582, n43583, n43584, n43585, n43586,
         n43587, n43588, n43589, n43590, n43591, n43592, n43593, n43594,
         n43595, n43596, n43597, n43598, n43599, n43600, n43601, n43602,
         n43603, n43604, n43605, n43606, n43607, n43608, n43609, n43610,
         n43611, n43612, n43613, n43614, n43615, n43616, n43617, n43618,
         n43619, n43620, n43621, n43622, n43623, n43624, n43625, n43626,
         n43627, n43628, n43629, n43630, n43631, n43632, n43633, n43634,
         n43635, n43636, n43637, n43638, n43639, n43640, n43641, n43642,
         n43643, n43644, n43645, n43646, n43647, n43648, n43649, n43650,
         n43651, n43652, n43653, n43654, n43655, n43656, n43657, n43658,
         n43659, n43660, n43661, n43662, n43663, n43664, n43665, n43666,
         n43667, n43668, n43669, n43670, n43671, n43672, n43673, n43674,
         n43675, n43676, n43677, n43678, n43679, n43680, n43681, n43682,
         n43683, n43684, n43685, n43686, n43687, n43688, n43689, n43690,
         n43691, n43692, n43693, n43694, n43695, n43696, n43697, n43698,
         n43699, n43700, n43701, n43702, n43703, n43704, n43705, n43706,
         n43707, n43708, n43709, n43710, n43711, n43712, n43713, n43714,
         n43715, n43716, n43717, n43718, n43719, n43720, n43721, n43722,
         n43723, n43724, n43725, n43726, n43727, n43728, n43729, n43730,
         n43731, n43732, n43733, n43734, n43735, n43736, n43737, n43738,
         n43739, n43740, n43741, n43742, n43743, n43744, n43745, n43746,
         n43747, n43748, n43749, n43750, n43751, n43752, n43753, n43754,
         n43755, n43756, n43757, n43758, n43759, n43760, n43761, n43762,
         n43763, n43764, n43765, n43766, n43767, n43768, n43769, n43770,
         n43771, n43772, n43773, n43774, n43775, n43776, n43777, n43778,
         n43779, n43780, n43781, n43782, n43783, n43784, n43785, n43786,
         n43787, n43788, n43789, n43790, n43791, n43792, n43793, n43794,
         n43795, n43796, n43797, n43798, n43799, n43800, n43801, n43802,
         n43803, n43804, n43805, n43806, n43807, n43808, n43809, n43810,
         n43811, n43812, n43813, n43814, n43815, n43816, n43817, n43818,
         n43819, n43820, n43821, n43822, n43823, n43824, n43825, n43826,
         n43827, n43828, n43829, n43830, n43831, n43832, n43833, n43834,
         n43835, n43836, n43837, n43838, n43839, n43840, n43841, n43842,
         n43843, n43844, n43845, n43846, n43847, n43848, n43849, n43850,
         n43851, n43852, n43853, n43854, n43855, n43856, n43857, n43858,
         n43859, n43860, n43861, n43862, n43863, n43864, n43865, n43866,
         n43867, n43868, n43869, n43870, n43871, n43872, n43873, n43874,
         n43875, n43876, n43877, n43878, n43879, n43880, n43881, n43882,
         n43883, n43884, n43885, n43886, n43887, n43888, n43889, n43890,
         n43891, n43892, n43893, n43894, n43895, n43896, n43897, n43898,
         n43899, n43900, n43901, n43902, n43903, n43904, n43905, n43906,
         n43907, n43908, n43909, n43910, n43911, n43912, n43913, n43914,
         n43915, n43916, n43917, n43918, n43919, n43920, n43921, n43922,
         n43923, n43924, n43925, n43926, n43927, n43928, n43929, n43930,
         n43931, n43932, n43933, n43934, n43935, n43936, n43937, n43938,
         n43939, n43940, n43941, n43942, n43943, n43944, n43945, n43946,
         n43947, n43948, n43949, n43950, n43951, n43952, n43953, n43954,
         n43955, n43956, n43957, n43958, n43959, n43960, n43961, n43962,
         n43963, n43964, n43965, n43966, n43967, n43968, n43969, n43970,
         n43971, n43972, n43973, n43974, n43975, n43976, n43977, n43978,
         n43979, n43980, n43981, n43982, n43983, n43984, n43985, n43986,
         n43987, n43988, n43989, n43990, n43991, n43992, n43993, n43994,
         n43995, n43996, n43997, n43998, n43999, n44000, n44001, n44002,
         n44003, n44004, n44005, n44006, n44007, n44008, n44009, n44010,
         n44011, n44012, n44013, n44014, n44015, n44016, n44017, n44018,
         n44019, n44020, n44021, n44022, n44023, n44024, n44025, n44026,
         n44027, n44028, n44029, n44030, n44031, n44032, n44033, n44034,
         n44035, n44036, n44037, n44038, n44039, n44040, n44041, n44042,
         n44043, n44044, n44045, n44046, n44047, n44048, n44049, n44050,
         n44051, n44052, n44053, n44054, n44055, n44056, n44057, n44058,
         n44059, n44060, n44061, n44062, n44063, n44064, n44065, n44066,
         n44067, n44068, n44069, n44070, n44071, n44072, n44073, n44074,
         n44075, n44076, n44077, n44078, n44079, n44080, n44081, n44082,
         n44083, n44084, n44085, n44086, n44087, n44088, n44089, n44090,
         n44091, n44092, n44093, n44094, n44095, n44096, n44097, n44098,
         n44099, n44100, n44101, n44102, n44103, n44104, n44105, n44106,
         n44107, n44108, n44109, n44110, n44111, n44112, n44113, n44114,
         n44115, n44116, n44117, n44118, n44119, n44120, n44121, n44122,
         n44123, n44124, n44125, n44126, n44127, n44128, n44129, n44130,
         n44131, n44132, n44133, n44134, n44135, n44136, n44137, n44138,
         n44139, n44140, n44141, n44142, n44143, n44144, n44145, n44146,
         n44147, n44148, n44149, n44150, n44151, n44152, n44153, n44154,
         n44155, n44156, n44157, n44158, n44159, n44160, n44161, n44162,
         n44163, n44164, n44165, n44166, n44167, n44168, n44169, n44170,
         n44171, n44172, n44173, n44174, n44175, n44176, n44177, n44178,
         n44179, n44180, n44181, n44182, n44183, n44184, n44185, n44186,
         n44187, n44188, n44189, n44190, n44191, n44192, n44193, n44194,
         n44195, n44196, n44197, n44198, n44199, n44200, n44201, n44202,
         n44203, n44204, n44205, n44206, n44207, n44208, n44209, n44210,
         n44211, n44212, n44213, n44214, n44215, n44216, n44217, n44218,
         n44219, n44220, n44221, n44222, n44223, n44224, n44225, n44226,
         n44227, n44228, n44229, n44230, n44231, n44232, n44233, n44234,
         n44235, n44236, n44237, n44238, n44239, n44240, n44241, n44242,
         n44243, n44244, n44245, n44246, n44247, n44248, n44249, n44250,
         n44251, n44252, n44253, n44254, n44255, n44256, n44257, n44258,
         n44259, n44260, n44261, n44262, n44263, n44264, n44265, n44266,
         n44267, n44268, n44269, n44270, n44271, n44272, n44273, n44274,
         n44275, n44276, n44277, n44278, n44279, n44280, n44281, n44282,
         n44283, n44284, n44285, n44286, n44287, n44288, n44289, n44290,
         n44291, n44292, n44293, n44294, n44295, n44296, n44297, n44298,
         n44299, n44300, n44301, n44302, n44303, n44304, n44305, n44306,
         n44307, n44308, n44309, n44310, n44311, n44312, n44313, n44314,
         n44315, n44316, n44317, n44318, n44319, n44320, n44321, n44322,
         n44323, n44324, n44325, n44326, n44327, n44328, n44329, n44330,
         n44331, n44332, n44333, n44334, n44335, n44336, n44337, n44338,
         n44339, n44340, n44341, n44342, n44343, n44344, n44345, n44346,
         n44347, n44348, n44349, n44350, n44351, n44352, n44353, n44354,
         n44355, n44356, n44357, n44358, n44359, n44360, n44361, n44362,
         n44363, n44364, n44365, n44366, n44367, n44368, n44369, n44370,
         n44371, n44372, n44373, n44374, n44375, n44376, n44377, n44378,
         n44379, n44380, n44381, n44382, n44383, n44384, n44385, n44386,
         n44387, n44388, n44389, n44390, n44391, n44392, n44393, n44394,
         n44395, n44396, n44397, n44398, n44399, n44400, n44401, n44402,
         n44403, n44404, n44405, n44406, n44407, n44408, n44409, n44410,
         n44411, n44412, n44413, n44414, n44415, n44416, n44417, n44418,
         n44419, n44420, n44421, n44422, n44423, n44424, n44425, n44426,
         n44427, n44428, n44429, n44430, n44431, n44432, n44433, n44434,
         n44435, n44436, n44437, n44438, n44439, n44440, n44441, n44442,
         n44443, n44444, n44445, n44446, n44447, n44448, n44449, n44450,
         n44451, n44452, n44453, n44454, n44455, n44456, n44457, n44458,
         n44459, n44460, n44461, n44462, n44463, n44464, n44465, n44466,
         n44467, n44468, n44469, n44470, n44471, n44472, n44473, n44474,
         n44475, n44476, n44477, n44478, n44479, n44480, n44481, n44482,
         n44483, n44484, n44485, n44486, n44487, n44488, n44489, n44490,
         n44491, n44492, n44493, n44494, n44495, n44496, n44497, n44498,
         n44499, n44500, n44501, n44502, n44503, n44504, n44505, n44506,
         n44507, n44508, n44509, n44510, n44511, n44512, n44513, n44514,
         n44515, n44516, n44517, n44518, n44519, n44520, n44521, n44522,
         n44523, n44524, n44525, n44526, n44527, n44528, n44529, n44530,
         n44531, n44532, n44533, n44534, n44535, n44536, n44537, n44538,
         n44539, n44540, n44541, n44542, n44543, n44544, n44545, n44546,
         n44547, n44548, n44549, n44550, n44551, n44552, n44553, n44554,
         n44555, n44556, n44557, n44558, n44559, n44560, n44561, n44562,
         n44563, n44564, n44565, n44566, n44567, n44568, n44569, n44570,
         n44571, n44572, n44573, n44574, n44575, n44576, n44577, n44578,
         n44579, n44580, n44581, n44582, n44583, n44584, n44585, n44586,
         n44587, n44588, n44589, n44590, n44591, n44592, n44593, n44594,
         n44595, n44596, n44597, n44598, n44599, n44600, n44601, n44602,
         n44603, n44604, n44605, n44606, n44607, n44608, n44609, n44610,
         n44611, n44612, n44613, n44614, n44615, n44616, n44617, n44618,
         n44619, n44620, n44621, n44622, n44623, n44624, n44625, n44626,
         n44627, n44628, n44629, n44630, n44631, n44632, n44633, n44634,
         n44635, n44636, n44637, n44638, n44639, n44640, n44641, n44642,
         n44643, n44644, n44645, n44646, n44647, n44648, n44649, n44650,
         n44651, n44652, n44653, n44654, n44655, n44656, n44657, n44658,
         n44659, n44660, n44661, n44662, n44663, n44664, n44665, n44666,
         n44667, n44668, n44669, n44670, n44671, n44672, n44673, n44674,
         n44675, n44676, n44677, n44678, n44679, n44680, n44681, n44682,
         n44683, n44684, n44685, n44686, n44687, n44688, n44689, n44690,
         n44691, n44692, n44693, n44694, n44695, n44696, n44697, n44698,
         n44699, n44700, n44701, n44702, n44703, n44704, n44705, n44706,
         n44707, n44708, n44709, n44710, n44711, n44712, n44713, n44714,
         n44715, n44716, n44717, n44718, n44719, n44720, n44721, n44722,
         n44723, n44724, n44725, n44726, n44727, n44728, n44729, n44730,
         n44731, n44732, n44733, n44734, n44735, n44736, n44737, n44738,
         n44739, n44740, n44741, n44742, n44743, n44744, n44745, n44746,
         n44747, n44748, n44749, n44750, n44751, n44752, n44753, n44754,
         n44755, n44756, n44757, n44758, n44759, n44760, n44761, n44762,
         n44763, n44764, n44765, n44766, n44767, n44768, n44769, n44770,
         n44771, n44772, n44773, n44774, n44775, n44776, n44777, n44778,
         n44779, n44780, n44781, n44782, n44783, n44784, n44785, n44786,
         n44787, n44788, n44789, n44790, n44791, n44792, n44793, n44794,
         n44795, n44796, n44797, n44798, n44799, n44800, n44801, n44802,
         n44803, n44804, n44805, n44806, n44807, n44808, n44809, n44810,
         n44811, n44812, n44813, n44814, n44815, n44816, n44817, n44818,
         n44819, n44820, n44821, n44822, n44823, n44824, n44825, n44826,
         n44827, n44828, n44829, n44830, n44831, n44832, n44833, n44834,
         n44835, n44836, n44837, n44838, n44839, n44840, n44841, n44842,
         n44843, n44844, n44845, n44846, n44847, n44848, n44849, n44850,
         n44851, n44852, n44853, n44854, n44855, n44856, n44857, n44858,
         n44859, n44860, n44861, n44862, n44863, n44864, n44865, n44866,
         n44867, n44868, n44869, n44870, n44871, n44872, n44873, n44874,
         n44875, n44876, n44877, n44878, n44879, n44880, n44881, n44882,
         n44883, n44884, n44885, n44886, n44887, n44888, n44889, n44890,
         n44891, n44892, n44893, n44894, n44895, n44896, n44897, n44898,
         n44899, n44900, n44901, n44902, n44903, n44904, n44905, n44906,
         n44907, n44908, n44909, n44910, n44911, n44912, n44913, n44914,
         n44915, n44916, n44917, n44918, n44919, n44920, n44921, n44922,
         n44923, n44924, n44925, n44926, n44927, n44928, n44929, n44930,
         n44931, n44932, n44933, n44934, n44935, n44936, n44937, n44938,
         n44939, n44940, n44941, n44942, n44943, n44944, n44945, n44946,
         n44947, n44948, n44949, n44950, n44951, n44952, n44953, n44954,
         n44955, n44956, n44957, n44958, n44959, n44960, n44961, n44962,
         n44963, n44964, n44965, n44966, n44967, n44968, n44969, n44970,
         n44971, n44972, n44973, n44974, n44975, n44976, n44977, n44978,
         n44979, n44980, n44981, n44982, n44983, n44984, n44985, n44986,
         n44987, n44988, n44989, n44990, n44991, n44992, n44993, n44994,
         n44995, n44996, n44997, n44998, n44999, n45000, n45001, n45002,
         n45003, n45004, n45005, n45006, n45007, n45008, n45009, n45010,
         n45011, n45012, n45013, n45014, n45015, n45016, n45017, n45018,
         n45019, n45020, n45021, n45022, n45023, n45024, n45025, n45026,
         n45027, n45028, n45029, n45030, n45031, n45032, n45033, n45034,
         n45035, n45036, n45037, n45038, n45039, n45040, n45041, n45042,
         n45043, n45044, n45045, n45046, n45047, n45048, n45049, n45050,
         n45051, n45052, n45053, n45054, n45055, n45056, n45057, n45058,
         n45059, n45060, n45061, n45062, n45063, n45064, n45065, n45066,
         n45067, n45068, n45069, n45070, n45071, n45072, n45073, n45074,
         n45075, n45076, n45077, n45078, n45079, n45080, n45081, n45082,
         n45083, n45084, n45085, n45086, n45087, n45088, n45089, n45090,
         n45091, n45092, n45093, n45094, n45095, n45096, n45097, n45098,
         n45099, n45100, n45101, n45102, n45103, n45104, n45105, n45106,
         n45107, n45108, n45109, n45110, n45111, n45112, n45113, n45114,
         n45115, n45116, n45117, n45118, n45119, n45120, n45121, n45122,
         n45123, n45124, n45125, n45126, n45127, n45128, n45129, n45130,
         n45131, n45132, n45133, n45134, n45135, n45136, n45137, n45138,
         n45139, n45140, n45141, n45142, n45143, n45144, n45145, n45146,
         n45147, n45148, n45149, n45150, n45151, n45152, n45153, n45154,
         n45155, n45156, n45157, n45158, n45159, n45160, n45161, n45162,
         n45163, n45164, n45165, n45166, n45167, n45168, n45169, n45170,
         n45171, n45172, n45173, n45174, n45175, n45176, n45177, n45178,
         n45179, n45180, n45181, n45182, n45183, n45184, n45185, n45186,
         n45187, n45188, n45189, n45190, n45191, n45192, n45193, n45194,
         n45195, n45196, n45197, n45198, n45199, n45200, n45201, n45202,
         n45203, n45204, n45205, n45206, n45207, n45208, n45209, n45210,
         n45211, n45212, n45213, n45214, n45215, n45216, n45217, n45218,
         n45219, n45220, n45221, n45222, n45223, n45224, n45225, n45226,
         n45227, n45228, n45229, n45230, n45231, n45232, n45233, n45234,
         n45235, n45236, n45237, n45238, n45239, n45240, n45241, n45242,
         n45243, n45244, n45245, n45246, n45247, n45248, n45249, n45250,
         n45251, n45252, n45253, n45254, n45255, n45256, n45257, n45258,
         n45259, n45260, n45261, n45262, n45263, n45264, n45265, n45266,
         n45267, n45268, n45269, n45270, n45271, n45272, n45273, n45274,
         n45275, n45276, n45277, n45278, n45279, n45280, n45281, n45282,
         n45283, n45284, n45285, n45286, n45287, n45288, n45289, n45290,
         n45291, n45292, n45293, n45294, n45295, n45296, n45297, n45298,
         n45299, n45300, n45301, n45302, n45303, n45304, n45305, n45306,
         n45307, n45308, n45309, n45310, n45311, n45312, n45313, n45314,
         n45315, n45316, n45317, n45318, n45319, n45320, n45321, n45322,
         n45323, n45324, n45325, n45326, n45327, n45328, n45329, n45330,
         n45331, n45332, n45333, n45334, n45335, n45336, n45337, n45338,
         n45339, n45340, n45341, n45342, n45343, n45344, n45345, n45346,
         n45347, n45348, n45349, n45350, n45351, n45352, n45353, n45354,
         n45355, n45356, n45357, n45358, n45359, n45360, n45361, n45362,
         n45363, n45364, n45365, n45366, n45367, n45368, n45369, n45370,
         n45371, n45372, n45373, n45374, n45375, n45376, n45377, n45378,
         n45379, n45380, n45381, n45382, n45383, n45384, n45385, n45386,
         n45387, n45388, n45389, n45390, n45391, n45392, n45393, n45394,
         n45395, n45396, n45397, n45398, n45399, n45400, n45401, n45402,
         n45403, n45404, n45405, n45406, n45407, n45408, n45409, n45410,
         n45411, n45412, n45413, n45414, n45415, n45416, n45417, n45418,
         n45419, n45420, n45421, n45422, n45423, n45424, n45425, n45426,
         n45427, n45428, n45429, n45430, n45431, n45432, n45433, n45434,
         n45435, n45436, n45437, n45438, n45439, n45440, n45441, n45442,
         n45443, n45444, n45445, n45446, n45447, n45448, n45449, n45450,
         n45451, n45452, n45453, n45454, n45455, n45456, n45457, n45458,
         n45459, n45460, n45461, n45462, n45463, n45464, n45465, n45466,
         n45467, n45468, n45469, n45470, n45471, n45472, n45473, n45474,
         n45475, n45476, n45477, n45478, n45479, n45480, n45481, n45482,
         n45483, n45484, n45485, n45486, n45487, n45488, n45489, n45490,
         n45491, n45492, n45493, n45494, n45495, n45496, n45497, n45498,
         n45499, n45500, n45501, n45502, n45503, n45504, n45505, n45506,
         n45507, n45508, n45509, n45510, n45511, n45512, n45513, n45514,
         n45515, n45516, n45517, n45518, n45519, n45520, n45521, n45522,
         n45523, n45524, n45525, n45526, n45527, n45528, n45529, n45530,
         n45531, n45532, n45533, n45534, n45535, n45536, n45537, n45538,
         n45539, n45540, n45541, n45542, n45543, n45544, n45545, n45546,
         n45547, n45548, n45549, n45550, n45551, n45552, n45553, n45554,
         n45555, n45556, n45557, n45558, n45559, n45560, n45561, n45562,
         n45563, n45564, n45565, n45566, n45567, n45568, n45569, n45570,
         n45571, n45572, n45573, n45574, n45575, n45576, n45577, n45578,
         n45579, n45580, n45581, n45582, n45583, n45584, n45585, n45586,
         n45587, n45588, n45589, n45590, n45591, n45592, n45593, n45594,
         n45595, n45596, n45597, n45598, n45599, n45600, n45601, n45602,
         n45603, n45604, n45605, n45606, n45607, n45608, n45609, n45610,
         n45611, n45612, n45613, n45614, n45615, n45616, n45617, n45618,
         n45619, n45620, n45621, n45622, n45623, n45624, n45625, n45626,
         n45627, n45628, n45629, n45630, n45631, n45632, n45633, n45634,
         n45635, n45636, n45637, n45638, n45639, n45640, n45641, n45642,
         n45643, n45644, n45645, n45646, n45647, n45648, n45649, n45650,
         n45651, n45652, n45653, n45654, n45655, n45656, n45657, n45658,
         n45659, n45660, n45661, n45662, n45663, n45664, n45665, n45666,
         n45667, n45668, n45669, n45670, n45671, n45672, n45673, n45674,
         n45675, n45676, n45677, n45678, n45679, n45680, n45681, n45682,
         n45683, n45684, n45685, n45686, n45687, n45688, n45689, n45690,
         n45691, n45692, n45693, n45694, n45695, n45696, n45697, n45698,
         n45699, n45700, n45701, n45702, n45703, n45704, n45705, n45706,
         n45707, n45708, n45709, n45710, n45711, n45712, n45713, n45714,
         n45715, n45716, n45717, n45718, n45719, n45720, n45721, n45722,
         n45723, n45724, n45725, n45726, n45727, n45728, n45729, n45730,
         n45731, n45732, n45733, n45734, n45735, n45736, n45737, n45738,
         n45739, n45740, n45741, n45742, n45743, n45744, n45745, n45746,
         n45747, n45748, n45749, n45750, n45751, n45752, n45753, n45754,
         n45755, n45756, n45757, n45758, n45759, n45760, n45761, n45762,
         n45763, n45764, n45765, n45766, n45767, n45768, n45769, n45770,
         n45771, n45772, n45773, n45774, n45775, n45776, n45777, n45778,
         n45779, n45780, n45781, n45782, n45783, n45784, n45785, n45786,
         n45787, n45788, n45789, n45790, n45791, n45792, n45793, n45794,
         n45795, n45796, n45797, n45798, n45799, n45800, n45801, n45802,
         n45803, n45804, n45805, n45806, n45807, n45808, n45809, n45810,
         n45811, n45812, n45813, n45814, n45815, n45816, n45817, n45818,
         n45819, n45820, n45821, n45822, n45823, n45824, n45825, n45826,
         n45827, n45828, n45829, n45830, n45831, n45832, n45833, n45834,
         n45835, n45836, n45837, n45838, n45839, n45840, n45841, n45842,
         n45843, n45844, n45845, n45846, n45847, n45848, n45849, n45850,
         n45851, n45852, n45853, n45854, n45855, n45856, n45857, n45858,
         n45859, n45860, n45861, n45862, n45863, n45864, n45865, n45866,
         n45867, n45868, n45869, n45870, n45871, n45872, n45873, n45874,
         n45875, n45876, n45877, n45878, n45879, n45880, n45881, n45882,
         n45883, n45884, n45885, n45886, n45887, n45888, n45889, n45890,
         n45891, n45892, n45893, n45894, n45895, n45896, n45897, n45898,
         n45899, n45900, n45901, n45902, n45903, n45904, n45905, n45906,
         n45907, n45908, n45909, n45910, n45911, n45912, n45913, n45914,
         n45915, n45916, n45917, n45918, n45919, n45920, n45921, n45922,
         n45923, n45924, n45925, n45926, n45927, n45928, n45929, n45930,
         n45931, n45932, n45933, n45934, n45935, n45936, n45937, n45938,
         n45939, n45940, n45941, n45942, n45943, n45944, n45945, n45946,
         n45947, n45948, n45949, n45950, n45951, n45952, n45953, n45954,
         n45955, n45956, n45957, n45958, n45959, n45960, n45961, n45962,
         n45963, n45964, n45965, n45966, n45967, n45968, n45969, n45970,
         n45971, n45972, n45973, n45974, n45975, n45976, n45977, n45978,
         n45979, n45980, n45981, n45982, n45983, n45984, n45985, n45986,
         n45987, n45988, n45989, n45990, n45991, n45992, n45993, n45994,
         n45995, n45996, n45997, n45998, n45999, n46000, n46001, n46002,
         n46003, n46004, n46005, n46006, n46007, n46008, n46009, n46010,
         n46011, n46012, n46013, n46014, n46015, n46016, n46017, n46018,
         n46019, n46020, n46021, n46022, n46023, n46024, n46025, n46026,
         n46027, n46028, n46029, n46030, n46031, n46032, n46033, n46034,
         n46035, n46036, n46037, n46038, n46039, n46040, n46041, n46042,
         n46043, n46044, n46045, n46046, n46047, n46048, n46049, n46050,
         n46051, n46052, n46053, n46054, n46055, n46056, n46057, n46058,
         n46059, n46060, n46061, n46062, n46063, n46064, n46065, n46066,
         n46067, n46068, n46069, n46070, n46071, n46072, n46073, n46074,
         n46075, n46076, n46077, n46078, n46079, n46080, n46081, n46082,
         n46083, n46084, n46085, n46086, n46087, n46088, n46089, n46090,
         n46091, n46092, n46093, n46094, n46095, n46096, n46097, n46098,
         n46099, n46100, n46101, n46102, n46103, n46104, n46105, n46106,
         n46107, n46108, n46109, n46110, n46111, n46112, n46113, n46114,
         n46115, n46116, n46117, n46118, n46119, n46120, n46121, n46122,
         n46123, n46124, n46125, n46126, n46127, n46128, n46129, n46130,
         n46131, n46132, n46133, n46134, n46135, n46136, n46137, n46138,
         n46139, n46140, n46141, n46142, n46143, n46144, n46145, n46146,
         n46147, n46148, n46149, n46150, n46151, n46152, n46153, n46154,
         n46155, n46156, n46157, n46158, n46159, n46160, n46161, n46162,
         n46163, n46164, n46165, n46166, n46167, n46168, n46169, n46170,
         n46171, n46172, n46173, n46174, n46175, n46176, n46177, n46178,
         n46179, n46180, n46181, n46182, n46183, n46184, n46185, n46186,
         n46187, n46188, n46189, n46190, n46191, n46192, n46193, n46194,
         n46195, n46196, n46197, n46198, n46199, n46200, n46201, n46202,
         n46203, n46204, n46205, n46206, n46207, n46208, n46209, n46210,
         n46211, n46212, n46213, n46214, n46215, n46216, n46217, n46218,
         n46219, n46220, n46221, n46222, n46223, n46224, n46225, n46226,
         n46227, n46228, n46229, n46230, n46231, n46232, n46233, n46234,
         n46235, n46236, n46237, n46238, n46239, n46240, n46241, n46242,
         n46243, n46244, n46245, n46246, n46247, n46248, n46249, n46250,
         n46251, n46252, n46253, n46254, n46255, n46256, n46257, n46258,
         n46259, n46260, n46261, n46262, n46263, n46264, n46265, n46266,
         n46267, n46268, n46269, n46270, n46271, n46272, n46273, n46274,
         n46275, n46276, n46277, n46278, n46279, n46280, n46281, n46282,
         n46283, n46284, n46285, n46286, n46287, n46288, n46289, n46290,
         n46291, n46292, n46293, n46294, n46295, n46296, n46297, n46298,
         n46299, n46300, n46301, n46302, n46303, n46304, n46305, n46306,
         n46307, n46308, n46309, n46310, n46311, n46312, n46313, n46314,
         n46315, n46316, n46317, n46318, n46319, n46320, n46321, n46322,
         n46323, n46324, n46325, n46326, n46327, n46328, n46329, n46330,
         n46331, n46332, n46333, n46334, n46335, n46336, n46337, n46338,
         n46339, n46340, n46341, n46342, n46343, n46344, n46345, n46346,
         n46347, n46348, n46349, n46350, n46351, n46352, n46353, n46354,
         n46355, n46356, n46357, n46358, n46359, n46360, n46361, n46362,
         n46363, n46364, n46365, n46366, n46367, n46368, n46369, n46370,
         n46371, n46372, n46373, n46374, n46375, n46376, n46377, n46378,
         n46379, n46380, n46381, n46382, n46383, n46384, n46385, n46386,
         n46387, n46388, n46389, n46390, n46391, n46392, n46393, n46394,
         n46395, n46396, n46397, n46398, n46399, n46400, n46401, n46402,
         n46403, n46404, n46405, n46406, n46407, n46408, n46409, n46410,
         n46411, n46412, n46413, n46414, n46415, n46416, n46417, n46418,
         n46419, n46420, n46421, n46422, n46423, n46424, n46425, n46426,
         n46427, n46428, n46429, n46430, n46431, n46432, n46433, n46434,
         n46435, n46436, n46437, n46438, n46439, n46440, n46441, n46442,
         n46443, n46444, n46445, n46446, n46447, n46448, n46449, n46450,
         n46451, n46452, n46453, n46454, n46455, n46456, n46457, n46458,
         n46459, n46460, n46461, n46462, n46463, n46464, n46465, n46466,
         n46467, n46468, n46469, n46470, n46471, n46472, n46473, n46474,
         n46475, n46476, n46477, n46478, n46479, n46480, n46481, n46482,
         n46483, n46484, n46485, n46486, n46487, n46488, n46489, n46490,
         n46491, n46492, n46493, n46494, n46495, n46496, n46497, n46498,
         n46499, n46500, n46501, n46502, n46503, n46504, n46505, n46506,
         n46507, n46508, n46509, n46510, n46511, n46512, n46513, n46514,
         n46515, n46516, n46517, n46518, n46519, n46520, n46521, n46522,
         n46523, n46524, n46525, n46526, n46527, n46528, n46529, n46530,
         n46531, n46532, n46533, n46534, n46535, n46536, n46537, n46538,
         n46539, n46540, n46541, n46542, n46543, n46544, n46545, n46546,
         n46547, n46548, n46549, n46550, n46551, n46552, n46553, n46554,
         n46555, n46556, n46557, n46558, n46559, n46560, n46561, n46562,
         n46563, n46564, n46565, n46566, n46567, n46568, n46569, n46570,
         n46571, n46572, n46573, n46574, n46575, n46576, n46577, n46578,
         n46579, n46580, n46581, n46582, n46583, n46584, n46585, n46586,
         n46587, n46588, n46589, n46590, n46591, n46592, n46593, n46594,
         n46595, n46596, n46597, n46598, n46599, n46600, n46601, n46602,
         n46603, n46604, n46605, n46606, n46607, n46608, n46609, n46610,
         n46611, n46612, n46613, n46614, n46615, n46616, n46617, n46618,
         n46619, n46620, n46621, n46622, n46623, n46624, n46625, n46626,
         n46627, n46628, n46629, n46630, n46631, n46632, n46633, n46634,
         n46635, n46636, n46637, n46638, n46639, n46640, n46641, n46642,
         n46643, n46644, n46645, n46646, n46647, n46648, n46649, n46650,
         n46651, n46652, n46653, n46654, n46655, n46656, n46657, n46658,
         n46659, n46660, n46661, n46662, n46663, n46664, n46665, n46666,
         n46667, n46668, n46669, n46670, n46671, n46672, n46673, n46674,
         n46675, n46676, n46677, n46678, n46679, n46680, n46681, n46682,
         n46683, n46684, n46685, n46686, n46687, n46688, n46689, n46690,
         n46691, n46692, n46693, n46694, n46695, n46696, n46697, n46698,
         n46699, n46700, n46701, n46702, n46703, n46704, n46705, n46706,
         n46707, n46708, n46709, n46710, n46711, n46712, n46713, n46714,
         n46715, n46716, n46717, n46718, n46719, n46720, n46721, n46722,
         n46723, n46724, n46725, n46726, n46727, n46728, n46729, n46730,
         n46731, n46732, n46733, n46734, n46735, n46736, n46737, n46738,
         n46739, n46740, n46741, n46742, n46743, n46744, n46745, n46746,
         n46747, n46748, n46749, n46750, n46751, n46752, n46753, n46754,
         n46755, n46756, n46757, n46758, n46759, n46760, n46761, n46762,
         n46763, n46764, n46765, n46766, n46767, n46768, n46769, n46770,
         n46771, n46772, n46773, n46774, n46775, n46776, n46777, n46778,
         n46779, n46780, n46781, n46782, n46783, n46784, n46785, n46786,
         n46787, n46788, n46789, n46790, n46791, n46792, n46793, n46794,
         n46795, n46796, n46797, n46798, n46799, n46800, n46801, n46802,
         n46803, n46804, n46805, n46806, n46807, n46808, n46809, n46810,
         n46811, n46812, n46813, n46814, n46815, n46816, n46817, n46818,
         n46819, n46820, n46821, n46822, n46823, n46824, n46825, n46826,
         n46827, n46828, n46829, n46830, n46831, n46832, n46833, n46834,
         n46835, n46836, n46837, n46838, n46839, n46840, n46841, n46842,
         n46843, n46844, n46845, n46846, n46847, n46848, n46849, n46850,
         n46851, n46852, n46853, n46854, n46855, n46856, n46857, n46858,
         n46859, n46860, n46861, n46862, n46863, n46864, n46865, n46866,
         n46867, n46868, n46869, n46870, n46871, n46872, n46873, n46874,
         n46875, n46876, n46877, n46878, n46879, n46880, n46881, n46882,
         n46883, n46884, n46885, n46886, n46887, n46888, n46889, n46890,
         n46891, n46892, n46893, n46894, n46895, n46896, n46897, n46898,
         n46899, n46900, n46901, n46902, n46903, n46904, n46905, n46906,
         n46907, n46908, n46909, n46910, n46911, n46912, n46913, n46914,
         n46915, n46916, n46917, n46918, n46919, n46920, n46921, n46922,
         n46923, n46924, n46925, n46926, n46927, n46928, n46929, n46930,
         n46931, n46932, n46933, n46934, n46935, n46936, n46937, n46938,
         n46939, n46940, n46941, n46942, n46943, n46944, n46945, n46946,
         n46947, n46948, n46949, n46950, n46951, n46952, n46953, n46954,
         n46955, n46956, n46957, n46958, n46959, n46960, n46961, n46962,
         n46963, n46964, n46965, n46966, n46967, n46968, n46969, n46970,
         n46971, n46972, n46973, n46974, n46975, n46976, n46977, n46978,
         n46979, n46980, n46981, n46982, n46983, n46984, n46985, n46986,
         n46987, n46988, n46989, n46990, n46991, n46992, n46993, n46994,
         n46995, n46996, n46997, n46998, n46999, n47000, n47001, n47002,
         n47003, n47004, n47005, n47006, n47007, n47008, n47009, n47010,
         n47011, n47012, n47013, n47014, n47015, n47016, n47017, n47018,
         n47019, n47020, n47021, n47022, n47023, n47024, n47025, n47026,
         n47027, n47028, n47029, n47030, n47031, n47032, n47033, n47034,
         n47035, n47036, n47037, n47038, n47039, n47040, n47041, n47042,
         n47043, n47044, n47045, n47046, n47047, n47048, n47049, n47050,
         n47051, n47052, n47053, n47054, n47055, n47056, n47057, n47058,
         n47059, n47060, n47061, n47062, n47063, n47064, n47065, n47066,
         n47067, n47068, n47069, n47070, n47071, n47072, n47073, n47074,
         n47075, n47076, n47077, n47078, n47079, n47080, n47081, n47082,
         n47083, n47084, n47085, n47086, n47087, n47088, n47089, n47090,
         n47091, n47092, n47093, n47094, n47095, n47096, n47097, n47098,
         n47099, n47100, n47101, n47102, n47103, n47104, n47105, n47106,
         n47107, n47108, n47109, n47110, n47111, n47112, n47113, n47114,
         n47115, n47116, n47117, n47118, n47119, n47120, n47121, n47122,
         n47123, n47124, n47125, n47126, n47127, n47128, n47129, n47130,
         n47131, n47132, n47133, n47134, n47135, n47136, n47137, n47138,
         n47139, n47140, n47141, n47142, n47143, n47144, n47145, n47146,
         n47147, n47148, n47149, n47150, n47151, n47152, n47153, n47154,
         n47155, n47156, n47157, n47158, n47159, n47160, n47161, n47162,
         n47163, n47164, n47165, n47166, n47167, n47168, n47169, n47170,
         n47171, n47172, n47173, n47174, n47175, n47176, n47177, n47178,
         n47179, n47180, n47181, n47182, n47183, n47184, n47185, n47186,
         n47187, n47188, n47189, n47190, n47191, n47192, n47193, n47194,
         n47195, n47196, n47197, n47198, n47199, n47200, n47201, n47202,
         n47203, n47204, n47205, n47206, n47207, n47208, n47209, n47210,
         n47211, n47212, n47213, n47214, n47215, n47216, n47217, n47218,
         n47219, n47220, n47221, n47222, n47223, n47224, n47225, n47226,
         n47227, n47228, n47229, n47230, n47231, n47232, n47233, n47234,
         n47235, n47236, n47237, n47238, n47239, n47240, n47241, n47242,
         n47243, n47244, n47245, n47246, n47247, n47248, n47249, n47250,
         n47251, n47252, n47253, n47254, n47255, n47256, n47257, n47258,
         n47259, n47260, n47261, n47262, n47263, n47264, n47265, n47266,
         n47267, n47268, n47269, n47270, n47271, n47272, n47273, n47274,
         n47275, n47276, n47277, n47278, n47279, n47280, n47281, n47282,
         n47283, n47284, n47285, n47286, n47287, n47288, n47289, n47290,
         n47291, n47292, n47293, n47294, n47295, n47296, n47297, n47298,
         n47299, n47300, n47301, n47302, n47303, n47304, n47305, n47306,
         n47307, n47308, n47309, n47310, n47311, n47312, n47313, n47314,
         n47315, n47316, n47317, n47318, n47319, n47320, n47321, n47322,
         n47323, n47324, n47325, n47326, n47327, n47328, n47329, n47330,
         n47331, n47332, n47333, n47334, n47335, n47336, n47337, n47338,
         n47339, n47340, n47341, n47342, n47343, n47344, n47345, n47346,
         n47347, n47348, n47349, n47350, n47351, n47352, n47353, n47354,
         n47355, n47356, n47357, n47358, n47359, n47360, n47361, n47362,
         n47363, n47364, n47365, n47366, n47367, n47368, n47369, n47370,
         n47371, n47372, n47373, n47374, n47375, n47376, n47377, n47378,
         n47379, n47380, n47381, n47382, n47383, n47384, n47385, n47386,
         n47387, n47388, n47389, n47390, n47391, n47392, n47393, n47394,
         n47395, n47396, n47397, n47398, n47399, n47400, n47401, n47402,
         n47403, n47404, n47405, n47406, n47407, n47408, n47409, n47410,
         n47411, n47412, n47413, n47414, n47415, n47416, n47417, n47418,
         n47419, n47420, n47421, n47422, n47423, n47424, n47425, n47426,
         n47427, n47428, n47429, n47430, n47431, n47432, n47433, n47434,
         n47435, n47436, n47437, n47438, n47439, n47440, n47441, n47442,
         n47443, n47444, n47445, n47446, n47447, n47448, n47449, n47450,
         n47451, n47452, n47453, n47454, n47455, n47456, n47457, n47458,
         n47459, n47460, n47461, n47462, n47463, n47464, n47465, n47466,
         n47467, n47468, n47469, n47470, n47471, n47472, n47473, n47474,
         n47475, n47476, n47477, n47478, n47479, n47480, n47481, n47482,
         n47483, n47484, n47485, n47486, n47487, n47488, n47489, n47490,
         n47491, n47492, n47493, n47494, n47495, n47496, n47497, n47498,
         n47499, n47500, n47501, n47502, n47503, n47504, n47505, n47506,
         n47507, n47508, n47509, n47510, n47511, n47512, n47513, n47514,
         n47515, n47516, n47517, n47518, n47519, n47520, n47521, n47522,
         n47523, n47524, n47525, n47526, n47527, n47528, n47529, n47530,
         n47531, n47532, n47533, n47534, n47535, n47536, n47537, n47538,
         n47539, n47540, n47541, n47542, n47543, n47544, n47545, n47546,
         n47547, n47548, n47549, n47550, n47551, n47552, n47553, n47554,
         n47555, n47556, n47557, n47558, n47559, n47560, n47561, n47562,
         n47563, n47564, n47565, n47566, n47567, n47568, n47569, n47570,
         n47571, n47572, n47573, n47574, n47575, n47576, n47577, n47578,
         n47579, n47580, n47581, n47582, n47583, n47584, n47585, n47586,
         n47587, n47588, n47589, n47590, n47591, n47592, n47593, n47594,
         n47595, n47596, n47597, n47598, n47599, n47600, n47601, n47602,
         n47603, n47604, n47605, n47606, n47607, n47608, n47609, n47610,
         n47611, n47612, n47613, n47614, n47615, n47616, n47617, n47618,
         n47619, n47620, n47621, n47622, n47623, n47624, n47625, n47626,
         n47627, n47628, n47629, n47630, n47631, n47632, n47633, n47634,
         n47635, n47636, n47637, n47638, n47639, n47640, n47641, n47642,
         n47643, n47644, n47645, n47646, n47647, n47648, n47649, n47650,
         n47651, n47652, n47653, n47654, n47655, n47656, n47657, n47658,
         n47659, n47660, n47661, n47662, n47663, n47664, n47665, n47666,
         n47667, n47668, n47669, n47670, n47671, n47672, n47673, n47674,
         n47675, n47676, n47677, n47678, n47679, n47680, n47681, n47682,
         n47683, n47684, n47685, n47686, n47687, n47688, n47689, n47690,
         n47691, n47692, n47693, n47694, n47695, n47696, n47697, n47698,
         n47699, n47700, n47701, n47702, n47703, n47704, n47705, n47706,
         n47707, n47708, n47709, n47710, n47711, n47712, n47713, n47714,
         n47715, n47716, n47717, n47718, n47719, n47720, n47721, n47722,
         n47723, n47724, n47725, n47726, n47727, n47728, n47729, n47730,
         n47731, n47732, n47733, n47734, n47735, n47736, n47737, n47738,
         n47739, n47740, n47741, n47742, n47743, n47744, n47745, n47746,
         n47747, n47748, n47749, n47750, n47751, n47752, n47753, n47754,
         n47755, n47756, n47757, n47758, n47759, n47760, n47761, n47762,
         n47763, n47764, n47765, n47766, n47767, n47768, n47769, n47770,
         n47771, n47772, n47773, n47774, n47775, n47776, n47777, n47778,
         n47779, n47780, n47781, n47782, n47783, n47784, n47785, n47786,
         n47787, n47788, n47789, n47790, n47791, n47792, n47793, n47794,
         n47795, n47796, n47797, n47798, n47799, n47800, n47801, n47802,
         n47803, n47804, n47805, n47806, n47807, n47808, n47809, n47810,
         n47811, n47812, n47813, n47814, n47815, n47816, n47817, n47818,
         n47819, n47820, n47821, n47822, n47823, n47824, n47825, n47826,
         n47827, n47828, n47829, n47830, n47831, n47832, n47833, n47834,
         n47835, n47836, n47837, n47838, n47839, n47840, n47841, n47842,
         n47843, n47844, n47845, n47846, n47847, n47848, n47849, n47850,
         n47851, n47852, n47853, n47854, n47855, n47856, n47857, n47858,
         n47859, n47860, n47861, n47862, n47863, n47864, n47865, n47866,
         n47867, n47868, n47869, n47870, n47871, n47872, n47873, n47874,
         n47875, n47876, n47877, n47878, n47879, n47880, n47881, n47882,
         n47883, n47884, n47885, n47886, n47887, n47888, n47889, n47890,
         n47891, n47892, n47893, n47894, n47895, n47896, n47897, n47898,
         n47899, n47900, n47901, n47902, n47903, n47904, n47905, n47906,
         n47907, n47908, n47909, n47910, n47911, n47912, n47913, n47914,
         n47915, n47916, n47917, n47918, n47919, n47920, n47921, n47922,
         n47923, n47924, n47925, n47926, n47927, n47928, n47929, n47930,
         n47931, n47932, n47933, n47934, n47935, n47936, n47937, n47938,
         n47939, n47940, n47941, n47942, n47943, n47944, n47945, n47946,
         n47947, n47948, n47949, n47950, n47951, n47952, n47953, n47954,
         n47955, n47956, n47957, n47958, n47959, n47960, n47961, n47962,
         n47963, n47964, n47965, n47966, n47967, n47968, n47969, n47970,
         n47971, n47972, n47973, n47974, n47975, n47976, n47977, n47978,
         n47979, n47980, n47981, n47982, n47983, n47984, n47985, n47986,
         n47987, n47988, n47989, n47990, n47991, n47992, n47993, n47994,
         n47995, n47996, n47997, n47998, n47999, n48000, n48001, n48002,
         n48003, n48004, n48005, n48006, n48007, n48008, n48009, n48010,
         n48011, n48012, n48013, n48014, n48015, n48016, n48017, n48018,
         n48019, n48020, n48021, n48022, n48023, n48024, n48025, n48026,
         n48027, n48028, n48029, n48030, n48031, n48032, n48033, n48034,
         n48035, n48036, n48037, n48038, n48039, n48040, n48041, n48042,
         n48043, n48044, n48045, n48046, n48047, n48048, n48049, n48050,
         n48051, n48052, n48053, n48054, n48055, n48056, n48057, n48058,
         n48059, n48060, n48061, n48062, n48063, n48064, n48065, n48066,
         n48067, n48068, n48069, n48070, n48071, n48072, n48073, n48074,
         n48075, n48076, n48077, n48078, n48079, n48080, n48081, n48082,
         n48083, n48084, n48085, n48086, n48087, n48088, n48089, n48090,
         n48091, n48092, n48093, n48094, n48095, n48096, n48097, n48098,
         n48099, n48100, n48101, n48102, n48103, n48104, n48105, n48106,
         n48107, n48108, n48109, n48110, n48111, n48112, n48113, n48114,
         n48115, n48116, n48117, n48118, n48119, n48120, n48121, n48122,
         n48123, n48124, n48125, n48126, n48127, n48128, n48129, n48130,
         n48131, n48132, n48133, n48134, n48135, n48136, n48137, n48138,
         n48139, n48140, n48141, n48142, n48143, n48144, n48145, n48146,
         n48147, n48148, n48149, n48150, n48151, n48152, n48153, n48154,
         n48155, n48156, n48157, n48158, n48159, n48160, n48161, n48162,
         n48163, n48164, n48165, n48166, n48167, n48168, n48169, n48170,
         n48171, n48172, n48173, n48174, n48175, n48176, n48177, n48178,
         n48179, n48180, n48181, n48182, n48183, n48184, n48185, n48186,
         n48187, n48188, n48189, n48190, n48191, n48192, n48193, n48194,
         n48195, n48196, n48197, n48198, n48199, n48200, n48201, n48202,
         n48203, n48204, n48205, n48206, n48207, n48208, n48209, n48210,
         n48211, n48212, n48213, n48214, n48215, n48216, n48217, n48218,
         n48219, n48220, n48221, n48222, n48223, n48224, n48225, n48226,
         n48227, n48228, n48229, n48230, n48231, n48232, n48233, n48234,
         n48235, n48236, n48237, n48238, n48239, n48240, n48241, n48242,
         n48243, n48244, n48245, n48246, n48247, n48248, n48249, n48250,
         n48251, n48252, n48253, n48254, n48255, n48256, n48257, n48258,
         n48259, n48260, n48261, n48262, n48263, n48264, n48265, n48266,
         n48267, n48268, n48269, n48270, n48271, n48272, n48273, n48274,
         n48275, n48276, n48277, n48278, n48279, n48280, n48281, n48282,
         n48283, n48284, n48285, n48286, n48287, n48288, n48289, n48290,
         n48291, n48292, n48293, n48294, n48295, n48296, n48297, n48298,
         n48299, n48300, n48301, n48302, n48303, n48304, n48305, n48306,
         n48307, n48308, n48309, n48310, n48311, n48312, n48313, n48314,
         n48315, n48316, n48317, n48318, n48319, n48320, n48321, n48322,
         n48323, n48324, n48325, n48326, n48327, n48328, n48329, n48330,
         n48331, n48332, n48333, n48334, n48335, n48336, n48337, n48338,
         n48339, n48340, n48341, n48342, n48343, n48344, n48345, n48346,
         n48347, n48348, n48349, n48350, n48351, n48352, n48353, n48354,
         n48355, n48356, n48357, n48358, n48359, n48360, n48361, n48362,
         n48363, n48364, n48365, n48366, n48367, n48368, n48369, n48370,
         n48371, n48372, n48373, n48374, n48375, n48376, n48377, n48378,
         n48379, n48380, n48381, n48382, n48383, n48384, n48385, n48386,
         n48387, n48388, n48389, n48390, n48391, n48392, n48393, n48394,
         n48395, n48396, n48397, n48398, n48399, n48400, n48401, n48402,
         n48403, n48404, n48405, n48406, n48407, n48408, n48409, n48410,
         n48411, n48412, n48413, n48414, n48415, n48416, n48417, n48418,
         n48419, n48420, n48421, n48422, n48423, n48424, n48425, n48426,
         n48427, n48428, n48429, n48430, n48431, n48432, n48433, n48434,
         n48435, n48436, n48437, n48438, n48439, n48440, n48441, n48442,
         n48443, n48444, n48445, n48446, n48447, n48448, n48449, n48450,
         n48451, n48452, n48453, n48454, n48455, n48456, n48457, n48458,
         n48459, n48460, n48461, n48462, n48463, n48464, n48465, n48466,
         n48467, n48468, n48469, n48470, n48471, n48472, n48473, n48474,
         n48475, n48476, n48477, n48478, n48479, n48480, n48481, n48482,
         n48483, n48484, n48485, n48486, n48487, n48488, n48489, n48490,
         n48491, n48492, n48493, n48494, n48495, n48496, n48497, n48498,
         n48499, n48500, n48501, n48502, n48503, n48504, n48505, n48506,
         n48507, n48508, n48509, n48510, n48511, n48512, n48513, n48514,
         n48515, n48516, n48517, n48518, n48519, n48520, n48521, n48522,
         n48523, n48524, n48525, n48526, n48527, n48528, n48529, n48530,
         n48531, n48532, n48533, n48534, n48535, n48536, n48537, n48538,
         n48539, n48540, n48541, n48542, n48543, n48544, n48545, n48546,
         n48547, n48548, n48549, n48550, n48551, n48552, n48553, n48554,
         n48555, n48556, n48557, n48558, n48559, n48560, n48561, n48562,
         n48563, n48564, n48565, n48566, n48567, n48568, n48569, n48570,
         n48571, n48572, n48573, n48574, n48575, n48576, n48577, n48578,
         n48579, n48580, n48581, n48582, n48583, n48584, n48585, n48586,
         n48587, n48588, n48589, n48590, n48591, n48592, n48593, n48594,
         n48595, n48596, n48597, n48598, n48599, n48600, n48601, n48602,
         n48603, n48604, n48605, n48606, n48607, n48608, n48609, n48610,
         n48611, n48612, n48613, n48614, n48615, n48616, n48617, n48618,
         n48619, n48620, n48621, n48622, n48623, n48624, n48625, n48626,
         n48627, n48628, n48629, n48630, n48631, n48632, n48633, n48634,
         n48635, n48636, n48637, n48638, n48639, n48640, n48641, n48642,
         n48643, n48644, n48645, n48646, n48647, n48648, n48649, n48650,
         n48651, n48652, n48653, n48654, n48655, n48656, n48657, n48658,
         n48659, n48660, n48661, n48662, n48663, n48664, n48665, n48666,
         n48667, n48668, n48669, n48670, n48671, n48672, n48673, n48674,
         n48675, n48676, n48677, n48678, n48679, n48680, n48681, n48682,
         n48683, n48684, n48685, n48686, n48687, n48688, n48689, n48690,
         n48691, n48692, n48693, n48694, n48695, n48696, n48697, n48698,
         n48699, n48700, n48701, n48702, n48703, n48704, n48705, n48706,
         n48707, n48708, n48709, n48710, n48711, n48712, n48713, n48714,
         n48715, n48716, n48717, n48718, n48719, n48720, n48721, n48722,
         n48723, n48724, n48725, n48726, n48727, n48728, n48729, n48730,
         n48731, n48732, n48733, n48734, n48735, n48736, n48737, n48738,
         n48739, n48740, n48741, n48742, n48743, n48744, n48745, n48746,
         n48747, n48748, n48749, n48750, n48751, n48752, n48753, n48754,
         n48755, n48756, n48757, n48758, n48759, n48760, n48761, n48762,
         n48763, n48764, n48765, n48766, n48767, n48768, n48769, n48770,
         n48771, n48772, n48773, n48774, n48775, n48776, n48777, n48778,
         n48779, n48780, n48781, n48782, n48783, n48784, n48785, n48786,
         n48787, n48788, n48789, n48790, n48791, n48792, n48793, n48794,
         n48795, n48796, n48797, n48798, n48799, n48800, n48801, n48802,
         n48803, n48804, n48805, n48806, n48807, n48808, n48809, n48810,
         n48811, n48812, n48813, n48814, n48815, n48816, n48817, n48818,
         n48819, n48820, n48821, n48822, n48823, n48824, n48825, n48826,
         n48827, n48828, n48829, n48830, n48831, n48832, n48833, n48834,
         n48835, n48836, n48837, n48838, n48839, n48840, n48841, n48842,
         n48843, n48844, n48845, n48846, n48847, n48848, n48849, n48850,
         n48851, n48852, n48853, n48854, n48855, n48856, n48857, n48858,
         n48859, n48860, n48861, n48862, n48863, n48864, n48865, n48866,
         n48867, n48868, n48869, n48870, n48871, n48872, n48873, n48874,
         n48875, n48876, n48877, n48878, n48879, n48880, n48881, n48882,
         n48883, n48884, n48885, n48886, n48887, n48888, n48889, n48890,
         n48891, n48892, n48893, n48894, n48895, n48896, n48897, n48898,
         n48899, n48900, n48901, n48902, n48903, n48904, n48905, n48906,
         n48907, n48908, n48909, n48910, n48911, n48912, n48913, n48914,
         n48915, n48916, n48917, n48918, n48919, n48920, n48921, n48922,
         n48923, n48924, n48925, n48926, n48927, n48928, n48929, n48930,
         n48931, n48932, n48933, n48934, n48935, n48936, n48937, n48938,
         n48939, n48940, n48941, n48942, n48943, n48944, n48945, n48946,
         n48947, n48948, n48949, n48950, n48951, n48952, n48953, n48954,
         n48955, n48956, n48957, n48958, n48959, n48960, n48961, n48962,
         n48963, n48964, n48965, n48966, n48967, n48968, n48969, n48970,
         n48971, n48972, n48973, n48974, n48975, n48976, n48977, n48978,
         n48979, n48980, n48981, n48982, n48983, n48984, n48985, n48986,
         n48987, n48988, n48989, n48990, n48991, n48992, n48993, n48994,
         n48995, n48996, n48997, n48998, n48999, n49000, n49001, n49002,
         n49003, n49004, n49005, n49006, n49007, n49008, n49009, n49010,
         n49011, n49012, n49013, n49014, n49015, n49016, n49017, n49018,
         n49019, n49020, n49021, n49022, n49023, n49024, n49025, n49026,
         n49027, n49028, n49029, n49030, n49031, n49032, n49033, n49034,
         n49035, n49036, n49037, n49038, n49039, n49040, n49041, n49042,
         n49043, n49044, n49045, n49046, n49047, n49048, n49049, n49050,
         n49051, n49052, n49053, n49054, n49055, n49056, n49057, n49058,
         n49059, n49060, n49061, n49062, n49063, n49064, n49065, n49066,
         n49067, n49068, n49069, n49070, n49071, n49072, n49073, n49074,
         n49075, n49076, n49077, n49078, n49079, n49080, n49081, n49082,
         n49083, n49084, n49085, n49086, n49087, n49088, n49089, n49090,
         n49091, n49092, n49093, n49094, n49095, n49096, n49097, n49098,
         n49099, n49100, n49101, n49102, n49103, n49104, n49105, n49106,
         n49107, n49108, n49109, n49110, n49111, n49112, n49113, n49114,
         n49115, n49116, n49117, n49118, n49119, n49120, n49121, n49122,
         n49123, n49124, n49125, n49126, n49127, n49128, n49129, n49130,
         n49131, n49132, n49133, n49134, n49135, n49136, n49137, n49138,
         n49139, n49140, n49141, n49142, n49143, n49144, n49145, n49146,
         n49147, n49148, n49149, n49150, n49151, n49152, n49153, n49154,
         n49155, n49156, n49157, n49158, n49159, n49160, n49161, n49162,
         n49163, n49164, n49165, n49166, n49167, n49168, n49169, n49170,
         n49171, n49172, n49173, n49174, n49175, n49176, n49177, n49178,
         n49179, n49180, n49181, n49182, n49183, n49184, n49185, n49186,
         n49187, n49188, n49189, n49190, n49191, n49192, n49193, n49194,
         n49195, n49196, n49197, n49198, n49199, n49200, n49201, n49202,
         n49203, n49204, n49205, n49206, n49207, n49208, n49209, n49210,
         n49211, n49212, n49213, n49214, n49215, n49216, n49217, n49218,
         n49219, n49220, n49221, n49222, n49223, n49224, n49225, n49226,
         n49227, n49228, n49229, n49230, n49231, n49232, n49233, n49234,
         n49235, n49236, n49237, n49238, n49239, n49240, n49241, n49242,
         n49243, n49244, n49245, n49246, n49247, n49248, n49249, n49250,
         n49251, n49252, n49253, n49254, n49255, n49256, n49257, n49258,
         n49259, n49260, n49261, n49262, n49263, n49264, n49265, n49266,
         n49267, n49268, n49269, n49270, n49271, n49272, n49273, n49274,
         n49275, n49276, n49277, n49278, n49279, n49280, n49281, n49282,
         n49283, n49284, n49285, n49286, n49287, n49288, n49289, n49290,
         n49291, n49292, n49293, n49294, n49295, n49296, n49297, n49298,
         n49299, n49300, n49301, n49302, n49303, n49304, n49305, n49306,
         n49307, n49308, n49309, n49310, n49311, n49312, n49313, n49314,
         n49315, n49316, n49317, n49318, n49319, n49320, n49321, n49322,
         n49323, n49324, n49325, n49326, n49327, n49328, n49329, n49330,
         n49331, n49332, n49333, n49334, n49335, n49336, n49337, n49338,
         n49339, n49340, n49341, n49342, n49343, n49344, n49345, n49346,
         n49347, n49348, n49349, n49350, n49351, n49352, n49353, n49354,
         n49355, n49356, n49357, n49358, n49359, n49360, n49361, n49362,
         n49363, n49364, n49365, n49366, n49367, n49368, n49369, n49370,
         n49371, n49372, n49373, n49374, n49375, n49376, n49377, n49378,
         n49379, n49380, n49381, n49382, n49383, n49384, n49385, n49386,
         n49387, n49388, n49389, n49390, n49391, n49392, n49393, n49394,
         n49395, n49396, n49397, n49398, n49399, n49400, n49401, n49402,
         n49403, n49404, n49405, n49406, n49407, n49408, n49409, n49410,
         n49411, n49412, n49413, n49414, n49415, n49416, n49417, n49418,
         n49419, n49420, n49421, n49422, n49423, n49424, n49425, n49426,
         n49427, n49428, n49429, n49430, n49431, n49432, n49433, n49434,
         n49435, n49436, n49437, n49438, n49439, n49440, n49441, n49442,
         n49443, n49444, n49445, n49446, n49447, n49448, n49449, n49450,
         n49451, n49452, n49453, n49454, n49455, n49456, n49457, n49458,
         n49459, n49460, n49461, n49462, n49463, n49464, n49465, n49466,
         n49467, n49468, n49469, n49470, n49471, n49472, n49473, n49474,
         n49475, n49476, n49477, n49478, n49479, n49480, n49481, n49482,
         n49483, n49484, n49485, n49486, n49487, n49488, n49489, n49490,
         n49491, n49492, n49493, n49494, n49495, n49496, n49497, n49498,
         n49499, n49500, n49501, n49502, n49503, n49504, n49505, n49506,
         n49507, n49508, n49509, n49510, n49511, n49512, n49513, n49514,
         n49515, n49516, n49517, n49518, n49519, n49520, n49521, n49522,
         n49523, n49524, n49525, n49526, n49527, n49528, n49529, n49530,
         n49531, n49532, n49533, n49534, n49535, n49536, n49537, n49538,
         n49539, n49540, n49541, n49542, n49543, n49544, n49545, n49546,
         n49547, n49548, n49549, n49550, n49551, n49552, n49553, n49554,
         n49555, n49556, n49557, n49558, n49559, n49560, n49561, n49562,
         n49563, n49564, n49565, n49566, n49567, n49568, n49569, n49570,
         n49571, n49572, n49573, n49574, n49575, n49576, n49577, n49578,
         n49579, n49580, n49581, n49582, n49583, n49584, n49585, n49586,
         n49587, n49588, n49589, n49590, n49591, n49592, n49593, n49594,
         n49595, n49596, n49597, n49598, n49599, n49600, n49601, n49602,
         n49603, n49604, n49605, n49606, n49607, n49608, n49609, n49610,
         n49611, n49612, n49613, n49614, n49615, n49616, n49617, n49618,
         n49619, n49620, n49621, n49622, n49623, n49624, n49625, n49626,
         n49627, n49628, n49629, n49630, n49631, n49632, n49633, n49634,
         n49635, n49636, n49637, n49638, n49639, n49640, n49641, n49642,
         n49643, n49644, n49645, n49646, n49647, n49648, n49649, n49650,
         n49651, n49652, n49653, n49654, n49655, n49656, n49657, n49658,
         n49659, n49660, n49661, n49662, n49663, n49664, n49665, n49666,
         n49667, n49668, n49669, n49670, n49671, n49672, n49673, n49674,
         n49675, n49676, n49677, n49678, n49679, n49680, n49681, n49682,
         n49683, n49684, n49685, n49686, n49687, n49688, n49689, n49690,
         n49691, n49692, n49693, n49694, n49695, n49696, n49697, n49698,
         n49699, n49700, n49701, n49702, n49703, n49704, n49705, n49706,
         n49707, n49708, n49709, n49710, n49711, n49712, n49713, n49714,
         n49715, n49716, n49717, n49718, n49719, n49720, n49721, n49722,
         n49723, n49724, n49725, n49726, n49727, n49728, n49729, n49730,
         n49731, n49732, n49733, n49734, n49735, n49736, n49737, n49738,
         n49739, n49740, n49741, n49742, n49743, n49744, n49745, n49746,
         n49747, n49748, n49749, n49750, n49751, n49752, n49753, n49754,
         n49755, n49756, n49757, n49758, n49759, n49760, n49761, n49762,
         n49763, n49764, n49765, n49766, n49767, n49768, n49769, n49770,
         n49771, n49772, n49773, n49774, n49775, n49776, n49777, n49778,
         n49779, n49780, n49781, n49782, n49783, n49784, n49785, n49786,
         n49787, n49788, n49789, n49790, n49791, n49792, n49793, n49794,
         n49795, n49796, n49797, n49798, n49799, n49800, n49801, n49802,
         n49803, n49804, n49805, n49806, n49807, n49808, n49809, n49810,
         n49811, n49812, n49813, n49814, n49815, n49816, n49817, n49818,
         n49819, n49820, n49821, n49822, n49823, n49824, n49825, n49826,
         n49827, n49828, n49829, n49830, n49831, n49832, n49833, n49834,
         n49835, n49836, n49837, n49838, n49839, n49840, n49841, n49842,
         n49843, n49844, n49845, n49846, n49847, n49848, n49849, n49850,
         n49851, n49852, n49853, n49854, n49855, n49856, n49857, n49858,
         n49859, n49860, n49861, n49862, n49863, n49864, n49865, n49866,
         n49867, n49868, n49869, n49870, n49871, n49872, n49873, n49874,
         n49875, n49876, n49877, n49878, n49879, n49880, n49881, n49882,
         n49883, n49884, n49885, n49886, n49887, n49888, n49889, n49890,
         n49891, n49892, n49893, n49894, n49895, n49896, n49897, n49898,
         n49899, n49900, n49901, n49902, n49903, n49904, n49905, n49906,
         n49907, n49908, n49909, n49910, n49911, n49912, n49913, n49914,
         n49915, n49916, n49917, n49918, n49919, n49920, n49921, n49922,
         n49923, n49924, n49925, n49926, n49927, n49928, n49929, n49930,
         n49931, n49932, n49933, n49934, n49935, n49936, n49937, n49938,
         n49939, n49940, n49941, n49942, n49943, n49944, n49945, n49946,
         n49947, n49948, n49949, n49950, n49951, n49952, n49953, n49954,
         n49955, n49956, n49957, n49958, n49959, n49960, n49961, n49962,
         n49963, n49964, n49965, n49966, n49967, n49968, n49969, n49970,
         n49971, n49972, n49973, n49974, n49975, n49976, n49977, n49978,
         n49979, n49980, n49981, n49982, n49983, n49984, n49985, n49986,
         n49987, n49988, n49989, n49990, n49991, n49992, n49993, n49994,
         n49995, n49996, n49997, n49998, n49999, n50000, n50001, n50002,
         n50003, n50004, n50005, n50006, n50007, n50008, n50009, n50010,
         n50011, n50012, n50013, n50014, n50015, n50016, n50017, n50018,
         n50019, n50020, n50021, n50022, n50023, n50024, n50025, n50026,
         n50027, n50028, n50029, n50030, n50031, n50032, n50033, n50034,
         n50035, n50036, n50037, n50038, n50039, n50040, n50041, n50042,
         n50043, n50044, n50045, n50046, n50047, n50048, n50049, n50050,
         n50051, n50052, n50053, n50054, n50055, n50056, n50057, n50058,
         n50059, n50060, n50061, n50062, n50063, n50064, n50065, n50066,
         n50067, n50068, n50069, n50070, n50071, n50072, n50073, n50074,
         n50075, n50076, n50077, n50078, n50079, n50080, n50081, n50082,
         n50083, n50084, n50085, n50086, n50087, n50088, n50089, n50090,
         n50091, n50092, n50093, n50094, n50095, n50096, n50097, n50098,
         n50099, n50100, n50101, n50102, n50103, n50104, n50105, n50106,
         n50107, n50108, n50109, n50110, n50111, n50112, n50113, n50114,
         n50115, n50116, n50117, n50118, n50119, n50120, n50121, n50122,
         n50123, n50124, n50125, n50126, n50127, n50128, n50129, n50130,
         n50131, n50132, n50133, n50134, n50135, n50136, n50137, n50138,
         n50139, n50140, n50141, n50142, n50143, n50144, n50145, n50146,
         n50147, n50148, n50149, n50150, n50151, n50152, n50153, n50154,
         n50155, n50156, n50157, n50158, n50159, n50160, n50161, n50162,
         n50163, n50164, n50165, n50166, n50167, n50168, n50169, n50170,
         n50171, n50172, n50173, n50174, n50175, n50176, n50177, n50178,
         n50179, n50180, n50181, n50182, n50183, n50184, n50185, n50186,
         n50187, n50188, n50189, n50190, n50191, n50192, n50193, n50194,
         n50195, n50196, n50197, n50198, n50199, n50200, n50201, n50202,
         n50203, n50204, n50205, n50206, n50207, n50208, n50209, n50210,
         n50211, n50212, n50213, n50214, n50215, n50216, n50217, n50218,
         n50219, n50220, n50221, n50222, n50223, n50224, n50225, n50226,
         n50227, n50228, n50229, n50230, n50231, n50232, n50233, n50234,
         n50235, n50236, n50237, n50238, n50239, n50240, n50241, n50242,
         n50243, n50244, n50245, n50246, n50247, n50248, n50249, n50250,
         n50251, n50252, n50253, n50254, n50255, n50256, n50257, n50258,
         n50259, n50260, n50261, n50262, n50263, n50264, n50265, n50266,
         n50267, n50268, n50269, n50270, n50271, n50272, n50273, n50274,
         n50275, n50276, n50277, n50278, n50279, n50280, n50281, n50282,
         n50283, n50284, n50285, n50286, n50287, n50288, n50289, n50290,
         n50291, n50292, n50293, n50294, n50295, n50296, n50297, n50298,
         n50299, n50300, n50301, n50302, n50303, n50304, n50305, n50306,
         n50307, n50308, n50309, n50310, n50311, n50312, n50313, n50314,
         n50315, n50316, n50317, n50318, n50319, n50320, n50321, n50322,
         n50323, n50324, n50325, n50326, n50327, n50328, n50329, n50330,
         n50331, n50332, n50333, n50334, n50335, n50336, n50337, n50338,
         n50339, n50340, n50341, n50342, n50343, n50344, n50345, n50346,
         n50347, n50348, n50349, n50350, n50351, n50352, n50353, n50354,
         n50355, n50356, n50357, n50358, n50359, n50360, n50361, n50362,
         n50363, n50364, n50365, n50366, n50367, n50368, n50369, n50370,
         n50371, n50372, n50373, n50374, n50375, n50376, n50377, n50378,
         n50379, n50380, n50381, n50382, n50383, n50384, n50385, n50386,
         n50387, n50388, n50389, n50390, n50391, n50392, n50393, n50394,
         n50395, n50396, n50397, n50398, n50399, n50400, n50401, n50402,
         n50403, n50404, n50405, n50406, n50407, n50408, n50409, n50410,
         n50411, n50412, n50413, n50414, n50415, n50416, n50417, n50418,
         n50419, n50420, n50421, n50422, n50423, n50424, n50425, n50426,
         n50427, n50428, n50429, n50430, n50431, n50432, n50433, n50434,
         n50435, n50436, n50437, n50438, n50439, n50440, n50441, n50442,
         n50443, n50444, n50445, n50446, n50447, n50448, n50449, n50450,
         n50451, n50452, n50453, n50454, n50455, n50456, n50457, n50458,
         n50459, n50460, n50461, n50462, n50463, n50464, n50465, n50466,
         n50467, n50468, n50469, n50470, n50471, n50472, n50473, n50474,
         n50475, n50476, n50477, n50478, n50479, n50480, n50481, n50482,
         n50483, n50484, n50485, n50486, n50487, n50488, n50489, n50490,
         n50491, n50492, n50493, n50494, n50495, n50496, n50497, n50498,
         n50499, n50500, n50501, n50502, n50503, n50504, n50505, n50506,
         n50507, n50508, n50509, n50510, n50511, n50512, n50513, n50514,
         n50515, n50516, n50517, n50518, n50519, n50520, n50521, n50522,
         n50523, n50524, n50525, n50526, n50527, n50528, n50529, n50530,
         n50531, n50532, n50533, n50534, n50535, n50536, n50537, n50538,
         n50539, n50540, n50541, n50542, n50543, n50544, n50545, n50546,
         n50547, n50548, n50549, n50550, n50551, n50552, n50553, n50554,
         n50555, n50556, n50557, n50558, n50559, n50560, n50561, n50562,
         n50563, n50564, n50565, n50566, n50567, n50568, n50569, n50570,
         n50571, n50572, n50573, n50574, n50575, n50576, n50577, n50578,
         n50579, n50580, n50581, n50582, n50583, n50584, n50585, n50586,
         n50587, n50588, n50589, n50590, n50591, n50592, n50593, n50594,
         n50595, n50596, n50597, n50598, n50599, n50600, n50601, n50602,
         n50603, n50604, n50605, n50606, n50607, n50608, n50609, n50610,
         n50611, n50612, n50613, n50614, n50615, n50616, n50617, n50618,
         n50619, n50620, n50621, n50622, n50623, n50624, n50625, n50626,
         n50627, n50628, n50629, n50630, n50631, n50632, n50633, n50634,
         n50635, n50636, n50637, n50638, n50639, n50640, n50641, n50642,
         n50643, n50644, n50645, n50646, n50647, n50648, n50649, n50650,
         n50651, n50652, n50653, n50654, n50655, n50656, n50657, n50658,
         n50659, n50660, n50661, n50662, n50663, n50664, n50665, n50666,
         n50667, n50668, n50669, n50670, n50671, n50672, n50673, n50674,
         n50675, n50676, n50677, n50678, n50679, n50680, n50681, n50682,
         n50683, n50684, n50685, n50686, n50687, n50688, n50689, n50690,
         n50691, n50692, n50693, n50694, n50695, n50696, n50697, n50698,
         n50699, n50700, n50701, n50702, n50703, n50704, n50705, n50706,
         n50707, n50708, n50709, n50710, n50711, n50712, n50713, n50714,
         n50715, n50716, n50717, n50718, n50719, n50720, n50721, n50722,
         n50723, n50724, n50725, n50726, n50727, n50728, n50729, n50730,
         n50731, n50732, n50733, n50734, n50735, n50736, n50737, n50738,
         n50739, n50740, n50741, n50742, n50743, n50744, n50745, n50746,
         n50747, n50748, n50749, n50750, n50751, n50752, n50753, n50754,
         n50755, n50756, n50757, n50758, n50759, n50760, n50761, n50762,
         n50763, n50764, n50765, n50766, n50767, n50768, n50769, n50770,
         n50771, n50772, n50773, n50774, n50775, n50776, n50777, n50778,
         n50779, n50780, n50781, n50782, n50783, n50784, n50785, n50786,
         n50787, n50788, n50789, n50790, n50791, n50792, n50793, n50794,
         n50795, n50796, n50797, n50798, n50799, n50800, n50801, n50802,
         n50803, n50804, n50805, n50806, n50807, n50808, n50809, n50810,
         n50811, n50812, n50813, n50814, n50815, n50816, n50817, n50818,
         n50819, n50820, n50821, n50822, n50823, n50824, n50825, n50826,
         n50827, n50828, n50829, n50830, n50831, n50832, n50833, n50834,
         n50835, n50836, n50837, n50838, n50839, n50840, n50841, n50842,
         n50843, n50844, n50845, n50846, n50847, n50848, n50849, n50850,
         n50851, n50852, n50853, n50854, n50855, n50856, n50857, n50858,
         n50859, n50860, n50861, n50862, n50863, n50864, n50865, n50866,
         n50867, n50868, n50869, n50870, n50871, n50872, n50873, n50874,
         n50875, n50876, n50877, n50878, n50879, n50880, n50881, n50882,
         n50883, n50884, n50885, n50886, n50887, n50888, n50889, n50890,
         n50891, n50892, n50893, n50894, n50895, n50896, n50897, n50898,
         n50899, n50900, n50901, n50902, n50903, n50904, n50905, n50906,
         n50907, n50908, n50909, n50910, n50911, n50912, n50913, n50914,
         n50915, n50916, n50917, n50918, n50919, n50920, n50921, n50922,
         n50923, n50924, n50925, n50926, n50927, n50928, n50929, n50930,
         n50931, n50932, n50933, n50934, n50935, n50936, n50937, n50938,
         n50939, n50940, n50941, n50942, n50943, n50944, n50945, n50946,
         n50947, n50948, n50949, n50950, n50951, n50952, n50953, n50954,
         n50955, n50956, n50957, n50958, n50959, n50960, n50961, n50962,
         n50963, n50964, n50965, n50966, n50967, n50968, n50969, n50970,
         n50971, n50972, n50973, n50974, n50975, n50976, n50977, n50978,
         n50979, n50980, n50981, n50982, n50983, n50984, n50985, n50986,
         n50987, n50988, n50989, n50990, n50991, n50992, n50993, n50994,
         n50995, n50996, n50997, n50998, n50999, n51000, n51001, n51002,
         n51003, n51004, n51005, n51006, n51007, n51008, n51009, n51010,
         n51011, n51012, n51013, n51014, n51015, n51016, n51017, n51018,
         n51019, n51020, n51021, n51022, n51023, n51024, n51025, n51026,
         n51027, n51028, n51029, n51030, n51031, n51032, n51033, n51034,
         n51035, n51036, n51037, n51038, n51039, n51040, n51041, n51042,
         n51043, n51044, n51045, n51046, n51047, n51048, n51049, n51050,
         n51051, n51052, n51053, n51054, n51055, n51056, n51057, n51058,
         n51059, n51060, n51061, n51062, n51063, n51064, n51065, n51066,
         n51067, n51068, n51069, n51070, n51071, n51072, n51073, n51074,
         n51075, n51076, n51077, n51078, n51079, n51080, n51081, n51082,
         n51083, n51084, n51085, n51086, n51087, n51088, n51089, n51090,
         n51091, n51092, n51093, n51094, n51095, n51096, n51097, n51098,
         n51099, n51100, n51101, n51102, n51103, n51104, n51105, n51106,
         n51107, n51108, n51109, n51110, n51111, n51112, n51113, n51114,
         n51115, n51116, n51117, n51118, n51119, n51120, n51121, n51122,
         n51123, n51124, n51125, n51126, n51127, n51128, n51129, n51130,
         n51131, n51132, n51133, n51134, n51135, n51136, n51137, n51138,
         n51139, n51140, n51141, n51142, n51143, n51144, n51145, n51146,
         n51147, n51148, n51149, n51150, n51151, n51152, n51153, n51154,
         n51155, n51156, n51157, n51158, n51159, n51160, n51161, n51162,
         n51163, n51164, n51165, n51166, n51167, n51168, n51169, n51170,
         n51171, n51172, n51173, n51174, n51175, n51176, n51177, n51178,
         n51179, n51180, n51181, n51182, n51183, n51184, n51185, n51186,
         n51187, n51188, n51189, n51190, n51191, n51192, n51193, n51194,
         n51195, n51196, n51197, n51198, n51199, n51200, n51201, n51202,
         n51203, n51204, n51205, n51206, n51207, n51208, n51209, n51210,
         n51211, n51212, n51213, n51214, n51215, n51216, n51217, n51218,
         n51219, n51220, n51221, n51222, n51223, n51224, n51225, n51226,
         n51227, n51228, n51229, n51230, n51231, n51232, n51233, n51234,
         n51235, n51236, n51237, n51238, n51239, n51240, n51241, n51242,
         n51243, n51244, n51245, n51246, n51247, n51248, n51249, n51250,
         n51251, n51252, n51253, n51254, n51255, n51256, n51257, n51258,
         n51259, n51260, n51261, n51262, n51263, n51264, n51265, n51266,
         n51267, n51268, n51269, n51270, n51271, n51272, n51273, n51274,
         n51275, n51276, n51277, n51278, n51279, n51280, n51281, n51282,
         n51283, n51284, n51285, n51286, n51287, n51288, n51289, n51290,
         n51291, n51292, n51293, n51294, n51295, n51296, n51297, n51298,
         n51299, n51300, n51301, n51302, n51303, n51304, n51305, n51306,
         n51307, n51308, n51309, n51310, n51311, n51312, n51313, n51314,
         n51315, n51316, n51317, n51318, n51319, n51320, n51321, n51322,
         n51323, n51324, n51325, n51326, n51327, n51328, n51329, n51330,
         n51331, n51332, n51333, n51334, n51335, n51336, n51337, n51338,
         n51339, n51340, n51341, n51342, n51343, n51344, n51345, n51346,
         n51347, n51348, n51349, n51350, n51351, n51352, n51353, n51354,
         n51355, n51356, n51357, n51358, n51359, n51360, n51361, n51362,
         n51363, n51364, n51365, n51366, n51367, n51368, n51369, n51370,
         n51371, n51372, n51373, n51374, n51375, n51376, n51377, n51378,
         n51379, n51380, n51381, n51382, n51383, n51384, n51385, n51386,
         n51387, n51388, n51389, n51390, n51391, n51392, n51393, n51394,
         n51395, n51396, n51397, n51398, n51399, n51400, n51401, n51402,
         n51403, n51404, n51405, n51406, n51407, n51408, n51409, n51410,
         n51411, n51412, n51413, n51414, n51415, n51416, n51417, n51418,
         n51419, n51420, n51421, n51422, n51423, n51424, n51425, n51426,
         n51427, n51428, n51429, n51430, n51431, n51432, n51433, n51434,
         n51435, n51436, n51437, n51438, n51439, n51440, n51441, n51442,
         n51443, n51444, n51445, n51446, n51447, n51448, n51449, n51450,
         n51451, n51452, n51453, n51454, n51455, n51456, n51457, n51458,
         n51459, n51460, n51461, n51462, n51463, n51464, n51465, n51466,
         n51467, n51468, n51469, n51470, n51471, n51472, n51473, n51474,
         n51475, n51476, n51477, n51478, n51479, n51480, n51481, n51482,
         n51483, n51484, n51485, n51486, n51487, n51488, n51489, n51490,
         n51491, n51492, n51493, n51494, n51495, n51496, n51497, n51498,
         n51499, n51500, n51501, n51502, n51503, n51504, n51505, n51506,
         n51507, n51508, n51509, n51510, n51511, n51512, n51513, n51514,
         n51515, n51516, n51517, n51518, n51519, n51520, n51521, n51522,
         n51523, n51524, n51525, n51526, n51527, n51528, n51529, n51530,
         n51531, n51532, n51533, n51534, n51535, n51536, n51537, n51538,
         n51539, n51540, n51541, n51542, n51543, n51544, n51545, n51546,
         n51547, n51548, n51549, n51550, n51551, n51552, n51553, n51554,
         n51555, n51556, n51557, n51558, n51559, n51560, n51561, n51562,
         n51563, n51564, n51565, n51566, n51567, n51568, n51569, n51570,
         n51571, n51572, n51573, n51574, n51575, n51576, n51577, n51578,
         n51579, n51580, n51581, n51582, n51583, n51584, n51585, n51586,
         n51587, n51588, n51589, n51590, n51591, n51592, n51593, n51594,
         n51595, n51596, n51597, n51598, n51599, n51600, n51601, n51602,
         n51603, n51604, n51605, n51606, n51607, n51608, n51609, n51610,
         n51611, n51612, n51613, n51614, n51615, n51616, n51617, n51618,
         n51619, n51620, n51621, n51622, n51623, n51624, n51625, n51626,
         n51627, n51628, n51629, n51630, n51631, n51632, n51633, n51634,
         n51635, n51636, n51637, n51638, n51639, n51640, n51641, n51642,
         n51643, n51644, n51645, n51646, n51647, n51648, n51649, n51650,
         n51651, n51652, n51653, n51654, n51655, n51656, n51657, n51658,
         n51659, n51660, n51661, n51662, n51663, n51664, n51665, n51666,
         n51667, n51668, n51669, n51670, n51671, n51672, n51673, n51674,
         n51675, n51676, n51677, n51678, n51679, n51680, n51681, n51682,
         n51683, n51684, n51685, n51686, n51687, n51688, n51689, n51690,
         n51691, n51692, n51693, n51694, n51695, n51696, n51697, n51698,
         n51699, n51700, n51701, n51702, n51703, n51704, n51705, n51706,
         n51707, n51708, n51709, n51710, n51711, n51712, n51713, n51714,
         n51715, n51716, n51717, n51718, n51719, n51720, n51721, n51722,
         n51723, n51724, n51725, n51726, n51727, n51728, n51729, n51730,
         n51731, n51732, n51733, n51734, n51735, n51736, n51737, n51738,
         n51739, n51740, n51741, n51742, n51743, n51744, n51745, n51746,
         n51747, n51748, n51749, n51750, n51751, n51752, n51753, n51754,
         n51755, n51756, n51757, n51758, n51759, n51760, n51761, n51762,
         n51763, n51764, n51765, n51766, n51767, n51768, n51769, n51770,
         n51771, n51772, n51773, n51774, n51775, n51776, n51777, n51778,
         n51779, n51780, n51781, n51782, n51783, n51784, n51785, n51786,
         n51787, n51788, n51789, n51790, n51791, n51792, n51793, n51794,
         n51795, n51796, n51797, n51798, n51799, n51800, n51801, n51802,
         n51803, n51804, n51805, n51806, n51807, n51808, n51809, n51810,
         n51811, n51812, n51813, n51814, n51815, n51816, n51817, n51818,
         n51819, n51820, n51821, n51822, n51823, n51824, n51825, n51826,
         n51827, n51828, n51829, n51830, n51831, n51832, n51833, n51834,
         n51835, n51836, n51837, n51838, n51839, n51840, n51841, n51842,
         n51843, n51844, n51845, n51846, n51847, n51848, n51849, n51850,
         n51851, n51852, n51853, n51854, n51855, n51856, n51857, n51858,
         n51859, n51860, n51861, n51862, n51863, n51864, n51865, n51866,
         n51867, n51868, n51869, n51870, n51871, n51872, n51873, n51874,
         n51875, n51876, n51877, n51878, n51879, n51880, n51881, n51882,
         n51883, n51884, n51885, n51886, n51887, n51888, n51889, n51890,
         n51891, n51892, n51893, n51894, n51895, n51896, n51897, n51898,
         n51899, n51900, n51901, n51902, n51903, n51904, n51905, n51906,
         n51907, n51908, n51909, n51910, n51911, n51912, n51913, n51914,
         n51915, n51916, n51917, n51918, n51919, n51920, n51921, n51922,
         n51923, n51924, n51925, n51926, n51927, n51928, n51929, n51930,
         n51931, n51932, n51933, n51934, n51935, n51936, n51937, n51938,
         n51939, n51940, n51941, n51942, n51943, n51944, n51945, n51946,
         n51947, n51948, n51949, n51950, n51951, n51952, n51953, n51954,
         n51955, n51956, n51957, n51958, n51959, n51960, n51961, n51962,
         n51963, n51964, n51965, n51966, n51967, n51968, n51969, n51970,
         n51971, n51972, n51973, n51974, n51975, n51976, n51977, n51978,
         n51979, n51980, n51981, n51982, n51983, n51984, n51985, n51986,
         n51987, n51988, n51989, n51990, n51991, n51992, n51993, n51994,
         n51995, n51996, n51997, n51998, n51999, n52000, n52001, n52002,
         n52003, n52004, n52005, n52006, n52007, n52008, n52009, n52010,
         n52011, n52012, n52013, n52014, n52015, n52016, n52017, n52018,
         n52019, n52020, n52021, n52022, n52023, n52024, n52025, n52026,
         n52027, n52028, n52029, n52030, n52031, n52032, n52033, n52034,
         n52035, n52036, n52037, n52038, n52039, n52040, n52041, n52042,
         n52043, n52044, n52045, n52046, n52047, n52048, n52049, n52050,
         n52051, n52052, n52053, n52054, n52055, n52056, n52057, n52058,
         n52059, n52060, n52061, n52062, n52063, n52064, n52065, n52066,
         n52067, n52068, n52069, n52070, n52071, n52072, n52073, n52074,
         n52075, n52076, n52077, n52078, n52079, n52080, n52081, n52082,
         n52083, n52084, n52085, n52086, n52087, n52088, n52089, n52090,
         n52091, n52092, n52093, n52094, n52095, n52096, n52097, n52098,
         n52099, n52100, n52101, n52102, n52103, n52104, n52105, n52106,
         n52107, n52108, n52109, n52110, n52111, n52112, n52113, n52114,
         n52115, n52116, n52117, n52118, n52119, n52120, n52121, n52122,
         n52123, n52124, n52125, n52126, n52127, n52128, n52129, n52130,
         n52131, n52132, n52133, n52134, n52135, n52136, n52137, n52138,
         n52139, n52140, n52141, n52142, n52143, n52144, n52145, n52146,
         n52147, n52148, n52149, n52150, n52151, n52152, n52153, n52154,
         n52155, n52156, n52157, n52158, n52159, n52160, n52161, n52162,
         n52163, n52164, n52165, n52166, n52167, n52168, n52169, n52170,
         n52171, n52172, n52173, n52174, n52175, n52176, n52177, n52178,
         n52179, n52180, n52181, n52182, n52183, n52184, n52185, n52186,
         n52187, n52188, n52189, n52190, n52191, n52192, n52193, n52194,
         n52195, n52196, n52197, n52198, n52199, n52200, n52201, n52202,
         n52203, n52204, n52205, n52206, n52207, n52208, n52209, n52210,
         n52211, n52212, n52213, n52214, n52215, n52216, n52217, n52218,
         n52219, n52220, n52221, n52222, n52223, n52224, n52225, n52226,
         n52227, n52228, n52229, n52230, n52231, n52232, n52233, n52234,
         n52235, n52236, n52237, n52238, n52239, n52240, n52241, n52242,
         n52243, n52244, n52245, n52246, n52247, n52248, n52249, n52250,
         n52251, n52252, n52253, n52254, n52255, n52256, n52257, n52258,
         n52259, n52260, n52261, n52262, n52263, n52264, n52265, n52266,
         n52267, n52268, n52269, n52270, n52271, n52272, n52273, n52274,
         n52275, n52276, n52277, n52278, n52279, n52280, n52281, n52282,
         n52283, n52284, n52285, n52286, n52287, n52288, n52289, n52290,
         n52291, n52292, n52293, n52294, n52295, n52296, n52297, n52298,
         n52299, n52300, n52301, n52302, n52303, n52304, n52305, n52306,
         n52307, n52308, n52309, n52310, n52311, n52312, n52313, n52314,
         n52315, n52316, n52317, n52318, n52319, n52320, n52321, n52322,
         n52323, n52324, n52325, n52326, n52327, n52328, n52329, n52330,
         n52331, n52332, n52333, n52334, n52335, n52336, n52337, n52338,
         n52339, n52340, n52341, n52342, n52343, n52344, n52345, n52346,
         n52347, n52348, n52349, n52350, n52351, n52352, n52353, n52354,
         n52355, n52356, n52357, n52358, n52359, n52360, n52361, n52362,
         n52363, n52364, n52365, n52366, n52367, n52368, n52369, n52370,
         n52371, n52372, n52373, n52374, n52375, n52376, n52377, n52378,
         n52379, n52380, n52381, n52382, n52383, n52384, n52385, n52386,
         n52387, n52388, n52389, n52390, n52391, n52392, n52393, n52394,
         n52395, n52396, n52397, n52398, n52399, n52400, n52401, n52402,
         n52403, n52404, n52405, n52406, n52407, n52408, n52409, n52410,
         n52411, n52412, n52413, n52414, n52415, n52416, n52417, n52418,
         n52419, n52420, n52421, n52422, n52423, n52424, n52425, n52426,
         n52427, n52428, n52429, n52430, n52431, n52432, n52433, n52434,
         n52435, n52436, n52437, n52438, n52439, n52440, n52441, n52442,
         n52443, n52444, n52445, n52446, n52447, n52448, n52449, n52450,
         n52451, n52452, n52453, n52454, n52455, n52456, n52457, n52458,
         n52459, n52460, n52461, n52462, n52463, n52464, n52465, n52466,
         n52467, n52468, n52469, n52470, n52471, n52472, n52473, n52474,
         n52475, n52476, n52477, n52478, n52479, n52480, n52481, n52482,
         n52483, n52484, n52485, n52486, n52487, n52488, n52489, n52490,
         n52491, n52492, n52493, n52494, n52495, n52496, n52497, n52498,
         n52499, n52500, n52501, n52502, n52503, n52504, n52505, n52506,
         n52507, n52508, n52509, n52510, n52511, n52512, n52513, n52514,
         n52515, n52516, n52517, n52518, n52519, n52520, n52521, n52522,
         n52523, n52524, n52525, n52526, n52527, n52528, n52529, n52530,
         n52531, n52532, n52533, n52534, n52535, n52536, n52537, n52538,
         n52539, n52540, n52541, n52542, n52543, n52544, n52545, n52546,
         n52547, n52548, n52549, n52550, n52551, n52552, n52553, n52554,
         n52555, n52556, n52557, n52558, n52559, n52560, n52561, n52562,
         n52563, n52564, n52565, n52566, n52567, n52568, n52569, n52570,
         n52571, n52572, n52573, n52574, n52575, n52576, n52577, n52578,
         n52579, n52580, n52581, n52582, n52583, n52584, n52585, n52586,
         n52587, n52588, n52589, n52590, n52591, n52592, n52593, n52594,
         n52595, n52596, n52597, n52598, n52599, n52600, n52601, n52602,
         n52603, n52604, n52605, n52606, n52607, n52608, n52609, n52610,
         n52611, n52612, n52613, n52614, n52615, n52616, n52617, n52618,
         n52619, n52620, n52621, n52622, n52623, n52624, n52625, n52626,
         n52627, n52628, n52629, n52630, n52631, n52632, n52633, n52634,
         n52635, n52636, n52637, n52638, n52639, n52640, n52641, n52642,
         n52643, n52644, n52645, n52646, n52647, n52648, n52649, n52650,
         n52651, n52652, n52653, n52654, n52655, n52656, n52657, n52658,
         n52659, n52660, n52661, n52662, n52663, n52664, n52665, n52666,
         n52667, n52668, n52669, n52670, n52671, n52672, n52673, n52674,
         n52675, n52676, n52677, n52678, n52679, n52680, n52681, n52682,
         n52683, n52684, n52685, n52686, n52687, n52688, n52689, n52690,
         n52691, n52692, n52693, n52694, n52695, n52696, n52697, n52698,
         n52699, n52700, n52701, n52702, n52703, n52704, n52705, n52706,
         n52707, n52708, n52709, n52710, n52711, n52712, n52713, n52714,
         n52715, n52716, n52717, n52718, n52719, n52720, n52721, n52722,
         n52723, n52724, n52725, n52726, n52727, n52728, n52729, n52730,
         n52731, n52732, n52733, n52734, n52735, n52736, n52737, n52738,
         n52739, n52740, n52741, n52742, n52743, n52744, n52745, n52746,
         n52747, n52748, n52749, n52750, n52751, n52752, n52753, n52754,
         n52755, n52756, n52757, n52758, n52759, n52760, n52761, n52762,
         n52763, n52764, n52765, n52766, n52767, n52768, n52769, n52770,
         n52771, n52772, n52773, n52774, n52775, n52776, n52777, n52778,
         n52779, n52780, n52781, n52782, n52783, n52784, n52785, n52786,
         n52787, n52788, n52789, n52790, n52791, n52792, n52793, n52794,
         n52795, n52796, n52797, n52798, n52799, n52800, n52801, n52802,
         n52803, n52804, n52805, n52806, n52807, n52808, n52809, n52810,
         n52811, n52812, n52813, n52814, n52815, n52816, n52817, n52818,
         n52819, n52820, n52821, n52822, n52823, n52824, n52825, n52826,
         n52827, n52828, n52829, n52830, n52831, n52832, n52833, n52834,
         n52835, n52836, n52837, n52838, n52839, n52840, n52841, n52842,
         n52843, n52844, n52845, n52846, n52847, n52848, n52849, n52850,
         n52851, n52852, n52853, n52854, n52855, n52856, n52857, n52858,
         n52859, n52860, n52861, n52862, n52863, n52864, n52865, n52866,
         n52867, n52868, n52869, n52870, n52871, n52872, n52873, n52874,
         n52875, n52876, n52877, n52878, n52879, n52880, n52881, n52882,
         n52883, n52884, n52885, n52886, n52887, n52888, n52889, n52890,
         n52891, n52892, n52893, n52894, n52895, n52896, n52897, n52898,
         n52899, n52900, n52901, n52902, n52903, n52904, n52905, n52906,
         n52907, n52908, n52909, n52910, n52911, n52912, n52913, n52914,
         n52915, n52916, n52917, n52918, n52919, n52920, n52921, n52922,
         n52923, n52924, n52925, n52926, n52927, n52928, n52929, n52930,
         n52931, n52932, n52933, n52934, n52935, n52936, n52937, n52938,
         n52939, n52940, n52941, n52942, n52943, n52944, n52945, n52946,
         n52947, n52948, n52949, n52950, n52951, n52952, n52953, n52954,
         n52955, n52956, n52957, n52958, n52959, n52960, n52961, n52962,
         n52963, n52964, n52965, n52966, n52967, n52968, n52969, n52970,
         n52971, n52972, n52973, n52974, n52975, n52976, n52977, n52978,
         n52979, n52980, n52981, n52982, n52983, n52984, n52985, n52986,
         n52987, n52988, n52989, n52990, n52991, n52992, n52993, n52994,
         n52995, n52996, n52997, n52998, n52999, n53000, n53001, n53002,
         n53003, n53004, n53005, n53006, n53007, n53008, n53009, n53010,
         n53011, n53012, n53013, n53014, n53015, n53016, n53017, n53018,
         n53019, n53020, n53021, n53022, n53023, n53024, n53025, n53026,
         n53027, n53028, n53029, n53030, n53031, n53032, n53033, n53034,
         n53035, n53036, n53037, n53038, n53039, n53040, n53041, n53042,
         n53043, n53044, n53045, n53046, n53047, n53048, n53049, n53050,
         n53051, n53052, n53053, n53054, n53055, n53056, n53057, n53058,
         n53059, n53060, n53061, n53062, n53063, n53064, n53065, n53066,
         n53067, n53068, n53069, n53070, n53071, n53072, n53073, n53074,
         n53075, n53076, n53077, n53078, n53079, n53080, n53081, n53082,
         n53083, n53084, n53085, n53086, n53087, n53088, n53089, n53090,
         n53091, n53092, n53093, n53094, n53095, n53096, n53097, n53098,
         n53099, n53100, n53101, n53102, n53103, n53104, n53105, n53106,
         n53107, n53108, n53109, n53110, n53111, n53112, n53113, n53114,
         n53115, n53116, n53117, n53118, n53119, n53120, n53121, n53122,
         n53123, n53124, n53125, n53126, n53127, n53128, n53129, n53130,
         n53131, n53132, n53133, n53134, n53135, n53136, n53137, n53138,
         n53139, n53140, n53141, n53142, n53143, n53144, n53145, n53146,
         n53147, n53148, n53149, n53150, n53151, n53152, n53153, n53154,
         n53155, n53156, n53157, n53158, n53159, n53160, n53161, n53162,
         n53163, n53164, n53165, n53166, n53167, n53168, n53169, n53170,
         n53171, n53172, n53173, n53174, n53175, n53176, n53177, n53178,
         n53179, n53180, n53181, n53182, n53183, n53184, n53185, n53186,
         n53187, n53188, n53189, n53190, n53191, n53192, n53193, n53194,
         n53195, n53196, n53197, n53198, n53199, n53200, n53201, n53202,
         n53203, n53204, n53205, n53206, n53207, n53208, n53209, n53210,
         n53211, n53212, n53213, n53214, n53215, n53216, n53217, n53218,
         n53219, n53220, n53221, n53222, n53223, n53224, n53225, n53226,
         n53227, n53228, n53229, n53230, n53231, n53232, n53233, n53234,
         n53235, n53236, n53237, n53238, n53239, n53240, n53241, n53242,
         n53243, n53244, n53245, n53246, n53247, n53248, n53249, n53250,
         n53251, n53252, n53253, n53254, n53255, n53256, n53257, n53258,
         n53259, n53260, n53261, n53262, n53263, n53264, n53265, n53266,
         n53267, n53268, n53269, n53270, n53271, n53272, n53273, n53274,
         n53275, n53276, n53277, n53278, n53279, n53280, n53281, n53282,
         n53283, n53284, n53285, n53286, n53287, n53288, n53289, n53290,
         n53291, n53292, n53293, n53294, n53295, n53296, n53297, n53298,
         n53299, n53300, n53301, n53302, n53303, n53304, n53305, n53306,
         n53307, n53308, n53309, n53310, n53311, n53312, n53313, n53314,
         n53315, n53316, n53317, n53318, n53319, n53320, n53321, n53322,
         n53323, n53324, n53325, n53326, n53327, n53328, n53329, n53330,
         n53331, n53332, n53333, n53334, n53335, n53336, n53337, n53338,
         n53339, n53340, n53341, n53342, n53343, n53344, n53345, n53346,
         n53347, n53348, n53349, n53350, n53351, n53352, n53353, n53354,
         n53355, n53356, n53357, n53358, n53359, n53360, n53361, n53362,
         n53363, n53364, n53365, n53366, n53367, n53368, n53369, n53370,
         n53371, n53372, n53373, n53374, n53375, n53376, n53377, n53378,
         n53379, n53380, n53381, n53382, n53383, n53384, n53385, n53386,
         n53387, n53388, n53389, n53390, n53391, n53392, n53393, n53394,
         n53395, n53396, n53397, n53398, n53399, n53400, n53401, n53402,
         n53403, n53404, n53405, n53406, n53407, n53408, n53409, n53410,
         n53411, n53412, n53413, n53414, n53415, n53416, n53417, n53418,
         n53419, n53420, n53421, n53422, n53423, n53424, n53425, n53426,
         n53427, n53428, n53429, n53430, n53431, n53432, n53433, n53434,
         n53435, n53436, n53437, n53438, n53439, n53440, n53441, n53442,
         n53443, n53444, n53445, n53446, n53447, n53448, n53449, n53450,
         n53451, n53452, n53453, n53454, n53455, n53456, n53457, n53458,
         n53459, n53460, n53461, n53462, n53463, n53464, n53465, n53466,
         n53467, n53468, n53469, n53470, n53471, n53472, n53473, n53474,
         n53475, n53476, n53477, n53478, n53479, n53480, n53481, n53482,
         n53483, n53484, n53485, n53486, n53487, n53488, n53489, n53490,
         n53491, n53492, n53493, n53494, n53495, n53496, n53497, n53498,
         n53499, n53500, n53501, n53502, n53503, n53504, n53505, n53506,
         n53507, n53508, n53509, n53510, n53511, n53512, n53513, n53514,
         n53515, n53516, n53517, n53518, n53519, n53520, n53521, n53522,
         n53523, n53524, n53525, n53526, n53527, n53528, n53529, n53530,
         n53531, n53532, n53533, n53534, n53535, n53536, n53537, n53538,
         n53539, n53540, n53541, n53542, n53543, n53544, n53545, n53546,
         n53547, n53548, n53549, n53550, n53551, n53552, n53553, n53554,
         n53555, n53556, n53557, n53558, n53559, n53560, n53561, n53562,
         n53563, n53564, n53565, n53566, n53567, n53568, n53569, n53570,
         n53571, n53572, n53573, n53574, n53575, n53576, n53577, n53578,
         n53579, n53580, n53581, n53582, n53583, n53584, n53585, n53586,
         n53587, n53588, n53589, n53590, n53591, n53592, n53593, n53594,
         n53595, n53596, n53597, n53598, n53599, n53600, n53601, n53602,
         n53603, n53604, n53605, n53606, n53607, n53608, n53609, n53610,
         n53611, n53612, n53613, n53614, n53615, n53616, n53617, n53618,
         n53619, n53620, n53621, n53622, n53623, n53624, n53625, n53626,
         n53627, n53628, n53629, n53630, n53631, n53632, n53633, n53634,
         n53635, n53636, n53637, n53638, n53639, n53640, n53641, n53642,
         n53643, n53644, n53645, n53646, n53647, n53648, n53649, n53650,
         n53651, n53652, n53653, n53654, n53655, n53656, n53657, n53658,
         n53659, n53660, n53661, n53662, n53663, n53664, n53665, n53666,
         n53667, n53668, n53669, n53670, n53671, n53672, n53673, n53674,
         n53675, n53676, n53677, n53678, n53679, n53680, n53681, n53682,
         n53683, n53684, n53685, n53686, n53687, n53688, n53689, n53690,
         n53691, n53692, n53693, n53694, n53695, n53696, n53697, n53698,
         n53699, n53700, n53701, n53702, n53703, n53704, n53705, n53706,
         n53707, n53708, n53709, n53710, n53711, n53712, n53713, n53714,
         n53715, n53716, n53717, n53718, n53719, n53720, n53721, n53722,
         n53723, n53724, n53725, n53726, n53727, n53728, n53729, n53730,
         n53731, n53732, n53733, n53734, n53735, n53736, n53737, n53738,
         n53739, n53740, n53741, n53742, n53743, n53744, n53745, n53746,
         n53747, n53748, n53749, n53750, n53751, n53752, n53753, n53754,
         n53755, n53756, n53757, n53758, n53759, n53760, n53761, n53762,
         n53763, n53764, n53765, n53766, n53767, n53768, n53769, n53770,
         n53771, n53772, n53773, n53774, n53775, n53776, n53777, n53778,
         n53779, n53780, n53781, n53782, n53783, n53784, n53785, n53786,
         n53787, n53788, n53789, n53790, n53791, n53792, n53793, n53794,
         n53795, n53796, n53797, n53798, n53799, n53800, n53801, n53802,
         n53803, n53804, n53805, n53806, n53807, n53808, n53809, n53810,
         n53811, n53812, n53813, n53814, n53815, n53816, n53817, n53818,
         n53819, n53820, n53821, n53822, n53823, n53824, n53825, n53826,
         n53827, n53828, n53829, n53830, n53831, n53832, n53833, n53834,
         n53835, n53836, n53837, n53838, n53839, n53840, n53841, n53842,
         n53843, n53844, n53845, n53846, n53847, n53848, n53849, n53850,
         n53851, n53852, n53853, n53854, n53855, n53856, n53857, n53858,
         n53859, n53860, n53861, n53862, n53863, n53864, n53865, n53866,
         n53867, n53868, n53869, n53870, n53871, n53872, n53873, n53874,
         n53875, n53876, n53877, n53878, n53879, n53880, n53881, n53882,
         n53883, n53884, n53885, n53886, n53887, n53888, n53889, n53890,
         n53891, n53892, n53893, n53894, n53895, n53896, n53897, n53898,
         n53899, n53900, n53901, n53902, n53903, n53904, n53905, n53906,
         n53907, n53908, n53909, n53910, n53911, n53912, n53913, n53914,
         n53915, n53916, n53917, n53918, n53919, n53920, n53921, n53922,
         n53923, n53924, n53925, n53926, n53927, n53928, n53929, n53930,
         n53931, n53932, n53933, n53934, n53935, n53936, n53937, n53938,
         n53939, n53940, n53941, n53942, n53943, n53944, n53945, n53946,
         n53947, n53948, n53949, n53950, n53951, n53952, n53953, n53954,
         n53955, n53956, n53957, n53958, n53959, n53960, n53961, n53962,
         n53963, n53964, n53965, n53966, n53967, n53968, n53969, n53970,
         n53971, n53972, n53973, n53974, n53975, n53976, n53977, n53978,
         n53979, n53980, n53981, n53982, n53983, n53984, n53985, n53986,
         n53987, n53988, n53989, n53990, n53991, n53992, n53993, n53994,
         n53995, n53996, n53997, n53998, n53999, n54000, n54001, n54002,
         n54003, n54004, n54005, n54006, n54007, n54008, n54009, n54010,
         n54011, n54012, n54013, n54014, n54015, n54016, n54017, n54018,
         n54019, n54020, n54021, n54022, n54023, n54024, n54025, n54026,
         n54027, n54028, n54029, n54030, n54031, n54032, n54033, n54034,
         n54035, n54036, n54037, n54038, n54039, n54040, n54041, n54042,
         n54043, n54044, n54045, n54046, n54047, n54048, n54049, n54050,
         n54051, n54052, n54053, n54054, n54055, n54056, n54057, n54058,
         n54059, n54060, n54061, n54062, n54063, n54064, n54065, n54066,
         n54067, n54068, n54069, n54070, n54071, n54072, n54073, n54074,
         n54075, n54076, n54077, n54078, n54079, n54080, n54081, n54082,
         n54083, n54084, n54085, n54086, n54087, n54088, n54089, n54090,
         n54091, n54092, n54093, n54094, n54095, n54096, n54097, n54098,
         n54099, n54100, n54101, n54102, n54103, n54104, n54105, n54106,
         n54107, n54108, n54109, n54110, n54111, n54112, n54113, n54114,
         n54115, n54116, n54117, n54118, n54119, n54120, n54121, n54122,
         n54123, n54124, n54125, n54126, n54127, n54128, n54129, n54130,
         n54131, n54132, n54133, n54134, n54135, n54136, n54137, n54138,
         n54139, n54140, n54141, n54142, n54143, n54144, n54145, n54146,
         n54147, n54148, n54149, n54150, n54151, n54152, n54153, n54154,
         n54155, n54156, n54157, n54158, n54159, n54160, n54161, n54162,
         n54163, n54164, n54165, n54166, n54167, n54168, n54169, n54170,
         n54171, n54172, n54173, n54174, n54175, n54176, n54177, n54178,
         n54179, n54180, n54181, n54182, n54183, n54184, n54185, n54186,
         n54187, n54188, n54189, n54190, n54191, n54192, n54193, n54194,
         n54195, n54196, n54197, n54198, n54199, n54200, n54201, n54202,
         n54203, n54204, n54205, n54206, n54207, n54208, n54209, n54210,
         n54211, n54212, n54213, n54214, n54215, n54216, n54217, n54218,
         n54219, n54220, n54221, n54222, n54223, n54224, n54225, n54226,
         n54227, n54228, n54229, n54230, n54231, n54232, n54233, n54234,
         n54235, n54236, n54237, n54238, n54239, n54240, n54241, n54242,
         n54243, n54244, n54245, n54246, n54247, n54248, n54249, n54250,
         n54251, n54252, n54253, n54254, n54255, n54256, n54257, n54258,
         n54259, n54260, n54261, n54262, n54263, n54264, n54265, n54266,
         n54267, n54268, n54269, n54270, n54271, n54272, n54273, n54274,
         n54275, n54276, n54277, n54278, n54279, n54280, n54281, n54282,
         n54283, n54284, n54285, n54286, n54287, n54288, n54289, n54290,
         n54291, n54292, n54293, n54294, n54295, n54296, n54297, n54298,
         n54299, n54300, n54301, n54302, n54303, n54304, n54305, n54306,
         n54307, n54308, n54309, n54310, n54311, n54312, n54313, n54314,
         n54315, n54316, n54317, n54318, n54319, n54320, n54321, n54322,
         n54323, n54324, n54325, n54326, n54327, n54328, n54329, n54330,
         n54331, n54332, n54333, n54334, n54335, n54336, n54337, n54338,
         n54339, n54340, n54341, n54342, n54343, n54344, n54345, n54346,
         n54347, n54348, n54349, n54350, n54351, n54352, n54353, n54354,
         n54355, n54356, n54357, n54358, n54359, n54360, n54361, n54362,
         n54363, n54364, n54365, n54366, n54367, n54368, n54369, n54370,
         n54371, n54372, n54373, n54374, n54375, n54376, n54377, n54378,
         n54379, n54380, n54381, n54382, n54383, n54384, n54385, n54386,
         n54387, n54388, n54389, n54390, n54391, n54392, n54393, n54394,
         n54395, n54396, n54397, n54398, n54399, n54400, n54401, n54402,
         n54403, n54404, n54405, n54406, n54407, n54408, n54409, n54410,
         n54411, n54412, n54413, n54414, n54415, n54416, n54417, n54418,
         n54419, n54420, n54421, n54422, n54423, n54424, n54425, n54426,
         n54427, n54428, n54429, n54430, n54431, n54432, n54433, n54434,
         n54435, n54436, n54437, n54438, n54439, n54440, n54441, n54442,
         n54443, n54444, n54445, n54446, n54447, n54448, n54449, n54450,
         n54451, n54452, n54453, n54454, n54455, n54456, n54457, n54458,
         n54459, n54460, n54461, n54462, n54463, n54464, n54465, n54466,
         n54467, n54468, n54469, n54470, n54471, n54472, n54473, n54474,
         n54475, n54476, n54477, n54478, n54479, n54480, n54481, n54482,
         n54483, n54484, n54485, n54486, n54487, n54488, n54489, n54490,
         n54491, n54492, n54493, n54494, n54495, n54496, n54497, n54498,
         n54499, n54500, n54501, n54502, n54503, n54504, n54505, n54506,
         n54507, n54508, n54509, n54510, n54511, n54512, n54513, n54514,
         n54515, n54516, n54517, n54518, n54519, n54520, n54521, n54522,
         n54523, n54524, n54525, n54526, n54527, n54528, n54529, n54530,
         n54531, n54532, n54533, n54534, n54535, n54536, n54537, n54538,
         n54539, n54540, n54541, n54542, n54543, n54544, n54545, n54546,
         n54547, n54548, n54549, n54550, n54551, n54552, n54553, n54554,
         n54555, n54556, n54557, n54558, n54559, n54560, n54561, n54562,
         n54563, n54564, n54565, n54566, n54567, n54568, n54569, n54570,
         n54571, n54572, n54573, n54574, n54575, n54576, n54577, n54578,
         n54579, n54580, n54581, n54582, n54583, n54584, n54585, n54586,
         n54587, n54588, n54589, n54590, n54591, n54592, n54593, n54594,
         n54595, n54596, n54597, n54598, n54599, n54600, n54601, n54602,
         n54603, n54604, n54605, n54606, n54607, n54608, n54609, n54610,
         n54611, n54612, n54613, n54614, n54615, n54616, n54617, n54618,
         n54619, n54620, n54621, n54622, n54623, n54624, n54625, n54626,
         n54627, n54628, n54629, n54630, n54631, n54632, n54633, n54634,
         n54635, n54636, n54637, n54638, n54639, n54640, n54641, n54642,
         n54643, n54644, n54645, n54646, n54647, n54648, n54649, n54650,
         n54651, n54652, n54653, n54654, n54655, n54656, n54657, n54658,
         n54659, n54660, n54661, n54662, n54663, n54664, n54665, n54666,
         n54667, n54668, n54669, n54670, n54671, n54672, n54673, n54674,
         n54675, n54676, n54677, n54678, n54679, n54680, n54681, n54682,
         n54683, n54684, n54685, n54686, n54687, n54688, n54689, n54690,
         n54691, n54692, n54693, n54694, n54695, n54696, n54697, n54698,
         n54699, n54700, n54701, n54702, n54703, n54704, n54705, n54706,
         n54707, n54708, n54709, n54710, n54711, n54712, n54713, n54714,
         n54715, n54716, n54717, n54718, n54719, n54720, n54721, n54722,
         n54723, n54724, n54725, n54726, n54727, n54728, n54729, n54730,
         n54731, n54732, n54733, n54734, n54735, n54736, n54737, n54738,
         n54739, n54740, n54741, n54742, n54743, n54744, n54745, n54746,
         n54747, n54748, n54749, n54750, n54751, n54752, n54753, n54754,
         n54755, n54756, n54757, n54758, n54759, n54760, n54761, n54762,
         n54763, n54764, n54765, n54766, n54767, n54768, n54769, n54770,
         n54771, n54772, n54773, n54774, n54775, n54776, n54777, n54778,
         n54779, n54780, n54781, n54782, n54783, n54784, n54785, n54786,
         n54787, n54788, n54789, n54790, n54791, n54792, n54793, n54794,
         n54795, n54796, n54797, n54798, n54799, n54800, n54801, n54802,
         n54803, n54804, n54805, n54806, n54807, n54808, n54809, n54810,
         n54811, n54812, n54813, n54814, n54815, n54816, n54817, n54818,
         n54819, n54820, n54821, n54822, n54823, n54824, n54825, n54826,
         n54827, n54828, n54829, n54830, n54831, n54832, n54833, n54834,
         n54835, n54836, n54837, n54838, n54839, n54840, n54841, n54842,
         n54843, n54844, n54845, n54846, n54847, n54848, n54849, n54850,
         n54851, n54852, n54853, n54854, n54855, n54856, n54857, n54858,
         n54859, n54860, n54861, n54862, n54863, n54864, n54865, n54866,
         n54867, n54868, n54869, n54870, n54871, n54872, n54873, n54874,
         n54875, n54876, n54877, n54878, n54879, n54880, n54881, n54882,
         n54883, n54884, n54885, n54886, n54887, n54888, n54889, n54890,
         n54891, n54892, n54893, n54894, n54895, n54896, n54897, n54898,
         n54899, n54900, n54901, n54902, n54903, n54904, n54905;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31;

  mult_N256_CC8_DW01_add_0 FS_1 ( .A({1'b0, \A1[284] , \A1[283] , \A1[282] , 
        \A1[281] , \A1[280] , \A1[279] , \A1[278] , \A1[277] , \A1[276] , 
        \A1[275] , \A1[274] , \A1[273] , \A1[272] , \A1[271] , \A1[270] , 
        \A1[269] , \A1[268] , \A1[267] , \A1[266] , \A1[265] , \A1[264] , 
        \A1[263] , \A1[262] , \A1[261] , \A1[260] , \A1[259] , \A1[258] , 
        \A1[257] , \A1[256] , \A1[255] , \A1[254] , \A1[253] , \A1[252] , 
        \A1[251] , \A1[250] , \A1[249] , \A1[248] , \A1[247] , \A1[246] , 
        \A1[245] , \A1[244] , \A1[243] , \A1[242] , \A1[241] , \A1[240] , 
        \A1[239] , \A1[238] , \A1[237] , \A1[236] , \A1[235] , \A1[234] , 
        \A1[233] , \A1[232] , \A1[231] , \A1[230] , \A1[229] , \A1[228] , 
        \A1[227] , \A1[226] , \A1[225] , \A1[224] , \A1[223] , \A1[222] , 
        \A1[221] , \A1[220] , \A1[219] , \A1[218] , \A1[217] , \A1[216] , 
        \A1[215] , \A1[214] , \A1[213] , \A1[212] , \A1[211] , \A1[210] , 
        \A1[209] , \A1[208] , \A1[207] , \A1[206] , \A1[205] , \A1[204] , 
        \A1[203] , \A1[202] , \A1[201] , \A1[200] , \A1[199] , \A1[198] , 
        \A1[197] , \A1[196] , \A1[195] , \A1[194] , \A1[193] , \A1[192] , 
        \A1[191] , \A1[190] , \A1[189] , \A1[188] , \A1[187] , \A1[186] , 
        \A1[185] , \A1[184] , \A1[183] , \A1[182] , \A1[181] , \A1[180] , 
        \A1[179] , \A1[178] , \A1[177] , \A1[176] , \A1[175] , \A1[174] , 
        \A1[173] , \A1[172] , \A1[171] , \A1[170] , \A1[169] , \A1[168] , 
        \A1[167] , \A1[166] , \A1[165] , \A1[164] , \A1[163] , \A1[162] , 
        \A1[161] , \A1[160] , \A1[159] , \A1[158] , \A1[157] , \A1[156] , 
        \A1[155] , \A1[154] , \A1[153] , \A1[152] , \A1[151] , \A1[150] , 
        \A1[149] , \A1[148] , \A1[147] , \A1[146] , \A1[145] , \A1[144] , 
        \A1[143] , \A1[142] , \A1[141] , \A1[140] , \A1[139] , \A1[138] , 
        \A1[137] , \A1[136] , \A1[135] , \A1[134] , \A1[133] , \A1[132] , 
        \A1[131] , \A1[130] , \A1[129] , \A1[128] , \A1[127] , \A1[126] , 
        \A1[125] , \A1[124] , \A1[123] , \A1[122] , \A1[121] , \A1[120] , 
        \A1[119] , \A1[118] , \A1[117] , \A1[116] , \A1[115] , \A1[114] , 
        \A1[113] , \A1[112] , \A1[111] , \A1[110] , \A1[109] , \A1[108] , 
        \A1[107] , \A1[106] , \A1[105] , \A1[104] , \A1[103] , \A1[102] , 
        \A1[101] , \A1[100] , \A1[99] , \A1[98] , \A1[97] , \A1[96] , \A1[95] , 
        \A1[94] , \A1[93] , \A1[92] , \A1[91] , \A1[90] , \A1[89] , \A1[88] , 
        \A1[87] , \A1[86] , \A1[85] , \A1[84] , \A1[83] , \A1[82] , \A1[81] , 
        \A1[80] , \A1[79] , \A1[78] , \A1[77] , \A1[76] , \A1[75] , \A1[74] , 
        \A1[73] , \A1[72] , \A1[71] , \A1[70] , \A1[69] , \A1[68] , \A1[67] , 
        \A1[66] , \A1[65] , \A1[64] , \A1[63] , \A1[62] , \A1[61] , \A1[60] , 
        \A1[59] , \A1[58] , \A1[57] , \A1[56] , \A1[55] , \A1[54] , \A1[53] , 
        \A1[52] , \A1[51] , \A1[50] , \A1[49] , \A1[48] , \A1[47] , \A1[46] , 
        \A1[45] , \A1[44] , \A1[43] , \A1[42] , \A1[41] , \A1[40] , \A1[39] , 
        \A1[38] , \A1[37] , \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , 
        \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] , \A1[26] , \A1[25] , 
        \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , 
        \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , 
        \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , 
        \A1[3] , \A1[2] , \A1[1] , \A1[0] }), .B({\A2[285] , \A2[284] , 
        \A2[283] , \A2[282] , \A2[281] , \A2[280] , \A2[279] , \A2[278] , 
        \A2[277] , \A2[276] , \A2[275] , \A2[274] , \A2[273] , \A2[272] , 
        \A2[271] , \A2[270] , \A2[269] , \A2[268] , \A2[267] , \A2[266] , 
        \A2[265] , \A2[264] , \A2[263] , \A2[262] , \A2[261] , \A2[260] , 
        \A2[259] , \A2[258] , \A2[257] , \A2[256] , \A2[255] , \A2[254] , 
        \A2[253] , \A2[252] , \A2[251] , \A2[250] , \A2[249] , \A2[248] , 
        \A2[247] , \A2[246] , \A2[245] , \A2[244] , \A2[243] , \A2[242] , 
        \A2[241] , \A2[240] , \A2[239] , \A2[238] , \A2[237] , \A2[236] , 
        \A2[235] , \A2[234] , \A2[233] , \A2[232] , \A2[231] , \A2[230] , 
        \A2[229] , \A2[228] , \A2[227] , \A2[226] , \A2[225] , \A2[224] , 
        \A2[223] , \A2[222] , \A2[221] , \A2[220] , \A2[219] , \A2[218] , 
        \A2[217] , \A2[216] , \A2[215] , \A2[214] , \A2[213] , \A2[212] , 
        \A2[211] , \A2[210] , \A2[209] , \A2[208] , \A2[207] , \A2[206] , 
        \A2[205] , \A2[204] , \A2[203] , \A2[202] , \A2[201] , \A2[200] , 
        \A2[199] , \A2[198] , \A2[197] , \A2[196] , \A2[195] , \A2[194] , 
        \A2[193] , \A2[192] , \A2[191] , \A2[190] , \A2[189] , \A2[188] , 
        \A2[187] , \A2[186] , \A2[185] , \A2[184] , \A2[183] , \A2[182] , 
        \A2[181] , \A2[180] , \A2[179] , \A2[178] , \A2[177] , \A2[176] , 
        \A2[175] , \A2[174] , \A2[173] , \A2[172] , \A2[171] , \A2[170] , 
        \A2[169] , \A2[168] , \A2[167] , \A2[166] , \A2[165] , \A2[164] , 
        \A2[163] , \A2[162] , \A2[161] , \A2[160] , \A2[159] , \A2[158] , 
        \A2[157] , \A2[156] , \A2[155] , \A2[154] , \A2[153] , \A2[152] , 
        \A2[151] , \A2[150] , \A2[149] , \A2[148] , \A2[147] , \A2[146] , 
        \A2[145] , \A2[144] , \A2[143] , \A2[142] , \A2[141] , \A2[140] , 
        \A2[139] , \A2[138] , \A2[137] , \A2[136] , \A2[135] , \A2[134] , 
        \A2[133] , \A2[132] , \A2[131] , \A2[130] , \A2[129] , \A2[128] , 
        \A2[127] , \A2[126] , \A2[125] , \A2[124] , \A2[123] , \A2[122] , 
        \A2[121] , \A2[120] , \A2[119] , \A2[118] , \A2[117] , \A2[116] , 
        \A2[115] , \A2[114] , \A2[113] , \A2[112] , \A2[111] , \A2[110] , 
        \A2[109] , \A2[108] , \A2[107] , \A2[106] , \A2[105] , \A2[104] , 
        \A2[103] , \A2[102] , \A2[101] , \A2[100] , \A2[99] , \A2[98] , 
        \A2[97] , \A2[96] , \A2[95] , \A2[94] , \A2[93] , \A2[92] , \A2[91] , 
        \A2[90] , \A2[89] , \A2[88] , \A2[87] , \A2[86] , \A2[85] , \A2[84] , 
        \A2[83] , \A2[82] , \A2[81] , \A2[80] , \A2[79] , \A2[78] , \A2[77] , 
        \A2[76] , \A2[75] , \A2[74] , \A2[73] , \A2[72] , \A2[71] , \A2[70] , 
        \A2[69] , \A2[68] , \A2[67] , \A2[66] , \A2[65] , \A2[64] , \A2[63] , 
        \A2[62] , \A2[61] , \A2[60] , \A2[59] , \A2[58] , \A2[57] , \A2[56] , 
        \A2[55] , \A2[54] , \A2[53] , \A2[52] , \A2[51] , \A2[50] , \A2[49] , 
        \A2[48] , \A2[47] , \A2[46] , \A2[45] , \A2[44] , \A2[43] , \A2[42] , 
        \A2[41] , \A2[40] , \A2[39] , \A2[38] , \A2[37] , \A2[36] , \A2[35] , 
        \A2[34] , \A2[33] , \A2[32] , \A2[31] , 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .CI(1'b0), .SUM({SYNOPSYS_UNCONNECTED__0, 
        SYNOPSYS_UNCONNECTED__1, SYNOPSYS_UNCONNECTED__2, 
        SYNOPSYS_UNCONNECTED__3, SYNOPSYS_UNCONNECTED__4, 
        SYNOPSYS_UNCONNECTED__5, SYNOPSYS_UNCONNECTED__6, 
        SYNOPSYS_UNCONNECTED__7, SYNOPSYS_UNCONNECTED__8, 
        SYNOPSYS_UNCONNECTED__9, SYNOPSYS_UNCONNECTED__10, 
        SYNOPSYS_UNCONNECTED__11, SYNOPSYS_UNCONNECTED__12, 
        SYNOPSYS_UNCONNECTED__13, SYNOPSYS_UNCONNECTED__14, 
        SYNOPSYS_UNCONNECTED__15, SYNOPSYS_UNCONNECTED__16, 
        SYNOPSYS_UNCONNECTED__17, SYNOPSYS_UNCONNECTED__18, 
        SYNOPSYS_UNCONNECTED__19, SYNOPSYS_UNCONNECTED__20, 
        SYNOPSYS_UNCONNECTED__21, SYNOPSYS_UNCONNECTED__22, 
        SYNOPSYS_UNCONNECTED__23, SYNOPSYS_UNCONNECTED__24, 
        SYNOPSYS_UNCONNECTED__25, SYNOPSYS_UNCONNECTED__26, 
        SYNOPSYS_UNCONNECTED__27, SYNOPSYS_UNCONNECTED__28, 
        SYNOPSYS_UNCONNECTED__29, SYNOPSYS_UNCONNECTED__30, 
        SYNOPSYS_UNCONNECTED__31, PRODUCT[255:2]}) );
  OR U2 ( .A(n54875), .B(n54872), .Z(n54884) );
  NANDN U3 ( .A(n3296), .B(n3295), .Z(n3291) );
  OR U4 ( .A(n52215), .B(n52213), .Z(n52323) );
  NANDN U5 ( .A(n2744), .B(n2743), .Z(n2739) );
  NANDN U6 ( .A(n2255), .B(n2254), .Z(n2250) );
  OR U7 ( .A(n52167), .B(n52165), .Z(n52305) );
  NANDN U8 ( .A(n1826), .B(n1825), .Z(n1821) );
  NANDN U9 ( .A(n1463), .B(n1462), .Z(n1458) );
  OR U10 ( .A(n52119), .B(n52117), .Z(n52287) );
  NANDN U11 ( .A(n1163), .B(n1162), .Z(n1158) );
  NANDN U12 ( .A(n922), .B(n921), .Z(n917) );
  OR U13 ( .A(n52071), .B(n52069), .Z(n52269) );
  NANDN U14 ( .A(n748), .B(n747), .Z(n743) );
  OR U15 ( .A(n52039), .B(n52037), .Z(n52257) );
  NANDN U16 ( .A(n637), .B(n636), .Z(n632) );
  OR U17 ( .A(n49418), .B(n49415), .Z(n49469) );
  OR U18 ( .A(n24375), .B(n24374), .Z(n24370) );
  OR U19 ( .A(n24952), .B(n24951), .Z(n24947) );
  OR U20 ( .A(n25378), .B(n25377), .Z(n25373) );
  OR U21 ( .A(n25804), .B(n25803), .Z(n25799) );
  OR U22 ( .A(n26230), .B(n26229), .Z(n26225) );
  OR U23 ( .A(n26656), .B(n26655), .Z(n26651) );
  OR U24 ( .A(n27226), .B(n27225), .Z(n27221) );
  OR U25 ( .A(n27652), .B(n27651), .Z(n27647) );
  OR U26 ( .A(n28078), .B(n28077), .Z(n28073) );
  OR U27 ( .A(n28504), .B(n28503), .Z(n28499) );
  OR U28 ( .A(n28930), .B(n28929), .Z(n28925) );
  OR U29 ( .A(n29497), .B(n29496), .Z(n29492) );
  OR U30 ( .A(n29923), .B(n29922), .Z(n29918) );
  OR U31 ( .A(n30349), .B(n30348), .Z(n30344) );
  OR U32 ( .A(n30775), .B(n30774), .Z(n30770) );
  OR U33 ( .A(n31201), .B(n31200), .Z(n31196) );
  OR U34 ( .A(n31757), .B(n31756), .Z(n31752) );
  OR U35 ( .A(n32183), .B(n32182), .Z(n32178) );
  OR U36 ( .A(n32609), .B(n32608), .Z(n32604) );
  OR U37 ( .A(n33035), .B(n33034), .Z(n33030) );
  OR U38 ( .A(n33461), .B(n33460), .Z(n33456) );
  OR U39 ( .A(n34010), .B(n34009), .Z(n34005) );
  OR U40 ( .A(n34436), .B(n34435), .Z(n34431) );
  OR U41 ( .A(n34862), .B(n34861), .Z(n34857) );
  OR U42 ( .A(n35288), .B(n35287), .Z(n35283) );
  OR U43 ( .A(n35714), .B(n35713), .Z(n35709) );
  OR U44 ( .A(n36256), .B(n36255), .Z(n36251) );
  OR U45 ( .A(n36682), .B(n36681), .Z(n36677) );
  OR U46 ( .A(n37108), .B(n37107), .Z(n37103) );
  OR U47 ( .A(n37534), .B(n37533), .Z(n37529) );
  OR U48 ( .A(n37960), .B(n37959), .Z(n37955) );
  OR U49 ( .A(n38495), .B(n38494), .Z(n38490) );
  OR U50 ( .A(n38921), .B(n38920), .Z(n38916) );
  OR U51 ( .A(n39347), .B(n39346), .Z(n39342) );
  OR U52 ( .A(n39773), .B(n39772), .Z(n39768) );
  OR U53 ( .A(n40199), .B(n40198), .Z(n40194) );
  OR U54 ( .A(n40727), .B(n40726), .Z(n40722) );
  OR U55 ( .A(n41153), .B(n41152), .Z(n41148) );
  OR U56 ( .A(n41579), .B(n41578), .Z(n41574) );
  OR U57 ( .A(n42005), .B(n42004), .Z(n42000) );
  OR U58 ( .A(n42431), .B(n42430), .Z(n42426) );
  OR U59 ( .A(n42952), .B(n42951), .Z(n42947) );
  OR U60 ( .A(n43378), .B(n43377), .Z(n43373) );
  OR U61 ( .A(n43804), .B(n43803), .Z(n43799) );
  OR U62 ( .A(n44230), .B(n44229), .Z(n44225) );
  OR U63 ( .A(n44656), .B(n44655), .Z(n44651) );
  OR U64 ( .A(n45170), .B(n45169), .Z(n45165) );
  OR U65 ( .A(n45596), .B(n45595), .Z(n45591) );
  OR U66 ( .A(n46022), .B(n46021), .Z(n46017) );
  OR U67 ( .A(n46448), .B(n46447), .Z(n46443) );
  OR U68 ( .A(n46874), .B(n46873), .Z(n46869) );
  OR U69 ( .A(n47381), .B(n47380), .Z(n47376) );
  OR U70 ( .A(n47807), .B(n47806), .Z(n47802) );
  OR U71 ( .A(n48233), .B(n48232), .Z(n48228) );
  OR U72 ( .A(n48659), .B(n48658), .Z(n48654) );
  OR U73 ( .A(n49085), .B(n49084), .Z(n49080) );
  OR U74 ( .A(n49904), .B(n49903), .Z(n49899) );
  OR U75 ( .A(n50330), .B(n50329), .Z(n50325) );
  OR U76 ( .A(n50756), .B(n50755), .Z(n50751) );
  OR U77 ( .A(n51182), .B(n51181), .Z(n51177) );
  OR U78 ( .A(n51608), .B(n51607), .Z(n51603) );
  OR U79 ( .A(n54893), .B(n54890), .Z(n54895) );
  OR U80 ( .A(n54850), .B(n54847), .Z(n54866) );
  OR U81 ( .A(n54779), .B(n54776), .Z(n54809) );
  OR U82 ( .A(n54680), .B(n54677), .Z(n54724) );
  OR U83 ( .A(n54553), .B(n54550), .Z(n54611) );
  OR U84 ( .A(n54398), .B(n54395), .Z(n54470) );
  OR U85 ( .A(n54215), .B(n54212), .Z(n54301) );
  OR U86 ( .A(n54004), .B(n54001), .Z(n54104) );
  OR U87 ( .A(n53765), .B(n53762), .Z(n53879) );
  OR U88 ( .A(n53498), .B(n53495), .Z(n53626) );
  OR U89 ( .A(n53203), .B(n53200), .Z(n53345) );
  OR U90 ( .A(n52880), .B(n52877), .Z(n53036) );
  OR U91 ( .A(n52529), .B(n52526), .Z(n52699) );
  OR U92 ( .A(n4555), .B(n4554), .Z(n4550) );
  OR U93 ( .A(n4981), .B(n4980), .Z(n4976) );
  OR U94 ( .A(n5407), .B(n5406), .Z(n5402) );
  OR U95 ( .A(n5833), .B(n5832), .Z(n5828) );
  OR U96 ( .A(n6262), .B(n6261), .Z(n6257) );
  OR U97 ( .A(n6688), .B(n6687), .Z(n6683) );
  OR U98 ( .A(n7114), .B(n7113), .Z(n7109) );
  OR U99 ( .A(n7540), .B(n7539), .Z(n7535) );
  OR U100 ( .A(n7966), .B(n7965), .Z(n7961) );
  OR U101 ( .A(n8396), .B(n8395), .Z(n8391) );
  OR U102 ( .A(n8822), .B(n8821), .Z(n8817) );
  OR U103 ( .A(n9248), .B(n9247), .Z(n9243) );
  OR U104 ( .A(n9674), .B(n9673), .Z(n9669) );
  OR U105 ( .A(n10100), .B(n10099), .Z(n10095) );
  OR U106 ( .A(n10529), .B(n10528), .Z(n10524) );
  OR U107 ( .A(n10955), .B(n10954), .Z(n10950) );
  OR U108 ( .A(n11381), .B(n11380), .Z(n11376) );
  OR U109 ( .A(n11807), .B(n11806), .Z(n11802) );
  NANDN U110 ( .A(n3699), .B(n3698), .Z(n3694) );
  OR U111 ( .A(n12233), .B(n12232), .Z(n12228) );
  OR U112 ( .A(n23949), .B(n23948), .Z(n23944) );
  OR U113 ( .A(n52231), .B(n52229), .Z(n52329) );
  NAND U114 ( .A(B[255]), .B(n16854), .Z(n16641) );
  OR U115 ( .A(n12663), .B(n12662), .Z(n12658) );
  OR U116 ( .A(n23523), .B(n23522), .Z(n23518) );
  OR U117 ( .A(n17064), .B(n17063), .Z(n17059) );
  OR U118 ( .A(n23097), .B(n23096), .Z(n23092) );
  OR U119 ( .A(n22671), .B(n22670), .Z(n22666) );
  OR U120 ( .A(n17490), .B(n17489), .Z(n17485) );
  OR U121 ( .A(n22087), .B(n22086), .Z(n22082) );
  OR U122 ( .A(n21661), .B(n21660), .Z(n21656) );
  OR U123 ( .A(n18088), .B(n18087), .Z(n18083) );
  OR U124 ( .A(n21235), .B(n21234), .Z(n21230) );
  OR U125 ( .A(n20809), .B(n20808), .Z(n20804) );
  OR U126 ( .A(n18514), .B(n18513), .Z(n18509) );
  OR U127 ( .A(n20383), .B(n20382), .Z(n20378) );
  OR U128 ( .A(n19792), .B(n19791), .Z(n19787) );
  OR U129 ( .A(n18940), .B(n18939), .Z(n18935) );
  OR U130 ( .A(n19366), .B(n19365), .Z(n19361) );
  NANDN U131 ( .A(n3105), .B(n3104), .Z(n3100) );
  OR U132 ( .A(n13157), .B(n13156), .Z(n13152) );
  OR U133 ( .A(n15672), .B(n15671), .Z(n15667) );
  NANDN U134 ( .A(n2574), .B(n2573), .Z(n2569) );
  OR U135 ( .A(n52183), .B(n52181), .Z(n52311) );
  OR U136 ( .A(n20176), .B(n20175), .Z(n20171) );
  NANDN U137 ( .A(n2103), .B(n2102), .Z(n2098) );
  OR U138 ( .A(n24745), .B(n24744), .Z(n24740) );
  OR U139 ( .A(n29290), .B(n29289), .Z(n29285) );
  NANDN U140 ( .A(n1698), .B(n1697), .Z(n1693) );
  OR U141 ( .A(n52135), .B(n52133), .Z(n52293) );
  OR U142 ( .A(n33803), .B(n33802), .Z(n33798) );
  NANDN U143 ( .A(n1356), .B(n1355), .Z(n1351) );
  OR U144 ( .A(n38288), .B(n38287), .Z(n38283) );
  OR U145 ( .A(n42745), .B(n42744), .Z(n42740) );
  NANDN U146 ( .A(n1077), .B(n1076), .Z(n1072) );
  OR U147 ( .A(n52087), .B(n52085), .Z(n52275) );
  OR U148 ( .A(n47174), .B(n47173), .Z(n47169) );
  NANDN U149 ( .A(n857), .B(n856), .Z(n852) );
  OR U150 ( .A(n49673), .B(n49670), .Z(n49682) );
  OR U151 ( .A(n49616), .B(n49613), .Z(n49639) );
  NANDN U152 ( .A(n704), .B(n703), .Z(n699) );
  NANDN U153 ( .A(n51843), .B(n51842), .Z(n51838) );
  OR U154 ( .A(n49531), .B(n49528), .Z(n49568) );
  OR U155 ( .A(n614), .B(n617), .Z(n52030) );
  NANDN U156 ( .A(n613), .B(n612), .Z(n608) );
  OR U157 ( .A(n49361), .B(n49359), .Z(n49404) );
  OR U158 ( .A(n49331), .B(n49329), .Z(n49392) );
  OR U159 ( .A(n24588), .B(n24587), .Z(n24583) );
  OR U160 ( .A(n25165), .B(n25164), .Z(n25160) );
  OR U161 ( .A(n25591), .B(n25590), .Z(n25586) );
  OR U162 ( .A(n26017), .B(n26016), .Z(n26012) );
  OR U163 ( .A(n26443), .B(n26442), .Z(n26438) );
  OR U164 ( .A(n26869), .B(n26868), .Z(n26864) );
  OR U165 ( .A(n27439), .B(n27438), .Z(n27434) );
  OR U166 ( .A(n27865), .B(n27864), .Z(n27860) );
  OR U167 ( .A(n28291), .B(n28290), .Z(n28286) );
  OR U168 ( .A(n28717), .B(n28716), .Z(n28712) );
  OR U169 ( .A(n29143), .B(n29142), .Z(n29138) );
  OR U170 ( .A(n29710), .B(n29709), .Z(n29705) );
  OR U171 ( .A(n30136), .B(n30135), .Z(n30131) );
  OR U172 ( .A(n30562), .B(n30561), .Z(n30557) );
  OR U173 ( .A(n30988), .B(n30987), .Z(n30983) );
  OR U174 ( .A(n31414), .B(n31413), .Z(n31409) );
  OR U175 ( .A(n31970), .B(n31969), .Z(n31965) );
  OR U176 ( .A(n32396), .B(n32395), .Z(n32391) );
  OR U177 ( .A(n32822), .B(n32821), .Z(n32817) );
  OR U178 ( .A(n33248), .B(n33247), .Z(n33243) );
  OR U179 ( .A(n33674), .B(n33673), .Z(n33669) );
  OR U180 ( .A(n34223), .B(n34222), .Z(n34218) );
  OR U181 ( .A(n34649), .B(n34648), .Z(n34644) );
  OR U182 ( .A(n35075), .B(n35074), .Z(n35070) );
  OR U183 ( .A(n35501), .B(n35500), .Z(n35496) );
  OR U184 ( .A(n35927), .B(n35926), .Z(n35922) );
  OR U185 ( .A(n36469), .B(n36468), .Z(n36464) );
  OR U186 ( .A(n36895), .B(n36894), .Z(n36890) );
  OR U187 ( .A(n37321), .B(n37320), .Z(n37316) );
  OR U188 ( .A(n37747), .B(n37746), .Z(n37742) );
  OR U189 ( .A(n38173), .B(n38172), .Z(n38168) );
  OR U190 ( .A(n38708), .B(n38707), .Z(n38703) );
  OR U191 ( .A(n39134), .B(n39133), .Z(n39129) );
  OR U192 ( .A(n39560), .B(n39559), .Z(n39555) );
  OR U193 ( .A(n39986), .B(n39985), .Z(n39981) );
  OR U194 ( .A(n40412), .B(n40411), .Z(n40407) );
  OR U195 ( .A(n40940), .B(n40939), .Z(n40935) );
  OR U196 ( .A(n41366), .B(n41365), .Z(n41361) );
  OR U197 ( .A(n41792), .B(n41791), .Z(n41787) );
  OR U198 ( .A(n42218), .B(n42217), .Z(n42213) );
  OR U199 ( .A(n42644), .B(n42643), .Z(n42639) );
  OR U200 ( .A(n43165), .B(n43164), .Z(n43160) );
  OR U201 ( .A(n43591), .B(n43590), .Z(n43586) );
  OR U202 ( .A(n44017), .B(n44016), .Z(n44012) );
  OR U203 ( .A(n44443), .B(n44442), .Z(n44438) );
  OR U204 ( .A(n44869), .B(n44868), .Z(n44864) );
  OR U205 ( .A(n45383), .B(n45382), .Z(n45378) );
  OR U206 ( .A(n45809), .B(n45808), .Z(n45804) );
  OR U207 ( .A(n46235), .B(n46234), .Z(n46230) );
  OR U208 ( .A(n46661), .B(n46660), .Z(n46656) );
  OR U209 ( .A(n47087), .B(n47086), .Z(n47082) );
  OR U210 ( .A(n47594), .B(n47593), .Z(n47589) );
  OR U211 ( .A(n48020), .B(n48019), .Z(n48015) );
  OR U212 ( .A(n48446), .B(n48445), .Z(n48441) );
  OR U213 ( .A(n48872), .B(n48871), .Z(n48867) );
  OR U214 ( .A(n49298), .B(n49297), .Z(n49293) );
  OR U215 ( .A(n50117), .B(n50116), .Z(n50112) );
  OR U216 ( .A(n50543), .B(n50542), .Z(n50538) );
  OR U217 ( .A(n50969), .B(n50968), .Z(n50964) );
  OR U218 ( .A(n51395), .B(n51394), .Z(n51390) );
  OR U219 ( .A(n51821), .B(n51820), .Z(n51816) );
  NANDN U220 ( .A(n3912), .B(n3915), .Z(n52245) );
  OR U221 ( .A(n54818), .B(n54815), .Z(n54841) );
  OR U222 ( .A(n54733), .B(n54730), .Z(n54770) );
  OR U223 ( .A(n54620), .B(n54617), .Z(n54671) );
  OR U224 ( .A(n54479), .B(n54476), .Z(n54544) );
  OR U225 ( .A(n54310), .B(n54307), .Z(n54389) );
  OR U226 ( .A(n54113), .B(n54110), .Z(n54206) );
  OR U227 ( .A(n53888), .B(n53885), .Z(n53995) );
  OR U228 ( .A(n53635), .B(n53632), .Z(n53756) );
  OR U229 ( .A(n53354), .B(n53351), .Z(n53489) );
  OR U230 ( .A(n53045), .B(n53042), .Z(n53194) );
  OR U231 ( .A(n52708), .B(n52705), .Z(n52871) );
  OR U232 ( .A(n52343), .B(n52340), .Z(n52520) );
  OR U233 ( .A(n4128), .B(n4127), .Z(n4123) );
  OR U234 ( .A(n4342), .B(n4341), .Z(n4337) );
  OR U235 ( .A(n4768), .B(n4767), .Z(n4763) );
  OR U236 ( .A(n5194), .B(n5193), .Z(n5189) );
  OR U237 ( .A(n5620), .B(n5619), .Z(n5615) );
  OR U238 ( .A(n6046), .B(n6045), .Z(n6041) );
  OR U239 ( .A(n6475), .B(n6474), .Z(n6470) );
  OR U240 ( .A(n6901), .B(n6900), .Z(n6896) );
  OR U241 ( .A(n7327), .B(n7326), .Z(n7322) );
  OR U242 ( .A(n7753), .B(n7752), .Z(n7748) );
  OR U243 ( .A(n8179), .B(n8178), .Z(n8174) );
  OR U244 ( .A(n8609), .B(n8608), .Z(n8604) );
  OR U245 ( .A(n9035), .B(n9034), .Z(n9030) );
  OR U246 ( .A(n9461), .B(n9460), .Z(n9456) );
  OR U247 ( .A(n9887), .B(n9886), .Z(n9882) );
  OR U248 ( .A(n10313), .B(n10312), .Z(n10308) );
  OR U249 ( .A(n10742), .B(n10741), .Z(n10737) );
  OR U250 ( .A(n11168), .B(n11167), .Z(n11163) );
  OR U251 ( .A(n11594), .B(n11593), .Z(n11589) );
  OR U252 ( .A(n12020), .B(n12019), .Z(n12015) );
  OR U253 ( .A(n24162), .B(n24161), .Z(n24157) );
  NANDN U254 ( .A(n52011), .B(n52010), .Z(n52006) );
  NANDN U255 ( .A(n3494), .B(n3493), .Z(n3489) );
  OR U256 ( .A(n12446), .B(n12445), .Z(n12441) );
  OR U257 ( .A(n23736), .B(n23735), .Z(n23731) );
  OR U258 ( .A(n16852), .B(n16851), .Z(n16847) );
  OR U259 ( .A(n23310), .B(n23309), .Z(n23305) );
  OR U260 ( .A(n17277), .B(n17276), .Z(n17272) );
  OR U261 ( .A(n22884), .B(n22883), .Z(n22879) );
  OR U262 ( .A(n22300), .B(n22299), .Z(n22295) );
  OR U263 ( .A(n17703), .B(n17702), .Z(n17698) );
  OR U264 ( .A(n21874), .B(n21873), .Z(n21869) );
  OR U265 ( .A(n21448), .B(n21447), .Z(n21443) );
  OR U266 ( .A(n18301), .B(n18300), .Z(n18296) );
  OR U267 ( .A(n21022), .B(n21021), .Z(n21017) );
  OR U268 ( .A(n20596), .B(n20595), .Z(n20591) );
  OR U269 ( .A(n18727), .B(n18726), .Z(n18722) );
  OR U270 ( .A(n20005), .B(n20004), .Z(n20000) );
  OR U271 ( .A(n19579), .B(n19578), .Z(n19574) );
  OR U272 ( .A(n19153), .B(n19152), .Z(n19148) );
  OR U273 ( .A(n12863), .B(n12862), .Z(n12858) );
  NANDN U274 ( .A(n51997), .B(n51996), .Z(n51992) );
  NANDN U275 ( .A(n16436), .B(n16433), .Z(n16432) );
  NANDN U276 ( .A(n2921), .B(n2920), .Z(n2916) );
  OR U277 ( .A(n14068), .B(n14067), .Z(n14063) );
  NANDN U278 ( .A(n51983), .B(n51982), .Z(n51978) );
  OR U279 ( .A(n52199), .B(n52197), .Z(n52317) );
  OR U280 ( .A(n17881), .B(n17880), .Z(n17876) );
  NANDN U281 ( .A(n51969), .B(n51968), .Z(n51964) );
  NANDN U282 ( .A(n2411), .B(n2410), .Z(n2406) );
  OR U283 ( .A(n22464), .B(n22463), .Z(n22459) );
  NANDN U284 ( .A(n51955), .B(n51954), .Z(n51950) );
  NANDN U285 ( .A(n1961), .B(n1960), .Z(n1956) );
  OR U286 ( .A(n27019), .B(n27018), .Z(n27014) );
  NANDN U287 ( .A(n51941), .B(n51940), .Z(n51936) );
  OR U288 ( .A(n52151), .B(n52149), .Z(n52299) );
  OR U289 ( .A(n31550), .B(n31549), .Z(n31545) );
  NANDN U290 ( .A(n51927), .B(n51926), .Z(n51922) );
  NANDN U291 ( .A(n1577), .B(n1576), .Z(n1572) );
  OR U292 ( .A(n36049), .B(n36048), .Z(n36044) );
  NANDN U293 ( .A(n51913), .B(n51912), .Z(n51908) );
  NANDN U294 ( .A(n1256), .B(n1255), .Z(n1251) );
  OR U295 ( .A(n40520), .B(n40519), .Z(n40515) );
  NANDN U296 ( .A(n51899), .B(n51898), .Z(n51894) );
  OR U297 ( .A(n52103), .B(n52101), .Z(n52281) );
  OR U298 ( .A(n44963), .B(n44962), .Z(n44958) );
  NANDN U299 ( .A(n51885), .B(n51884), .Z(n51880) );
  NANDN U300 ( .A(n994), .B(n993), .Z(n989) );
  OR U301 ( .A(n49691), .B(n49688), .Z(n49693) );
  NANDN U302 ( .A(n51871), .B(n51870), .Z(n51866) );
  NANDN U303 ( .A(n799), .B(n798), .Z(n794) );
  OR U304 ( .A(n49648), .B(n49645), .Z(n49664) );
  NANDN U305 ( .A(n51857), .B(n51856), .Z(n51852) );
  OR U306 ( .A(n52055), .B(n52053), .Z(n52263) );
  OR U307 ( .A(n49577), .B(n49574), .Z(n49607) );
  NANDN U308 ( .A(n667), .B(n666), .Z(n662) );
  OR U309 ( .A(n49478), .B(n49475), .Z(n49522) );
  OR U310 ( .A(n51624), .B(n51625), .Z(n51623) );
  NANDN U311 ( .A(n606), .B(n605), .Z(n601) );
  OR U312 ( .A(n49382), .B(n49379), .Z(n49408) );
  OR U313 ( .A(n49346), .B(n49344), .Z(n49398) );
  OR U314 ( .A(n49316), .B(n49314), .Z(n49386) );
  OR U315 ( .A(n12886), .B(n12887), .Z(n12885) );
  OR U316 ( .A(n12933), .B(n12934), .Z(n12932) );
  OR U317 ( .A(n13201), .B(n13202), .Z(n13200) );
  OR U318 ( .A(n13304), .B(n13305), .Z(n13303) );
  OR U319 ( .A(n13435), .B(n13436), .Z(n13434) );
  OR U320 ( .A(n13594), .B(n13595), .Z(n13593) );
  OR U321 ( .A(n13781), .B(n13782), .Z(n13780) );
  OR U322 ( .A(n14182), .B(n14183), .Z(n14181) );
  OR U323 ( .A(n14425), .B(n14426), .Z(n14424) );
  OR U324 ( .A(n14696), .B(n14697), .Z(n14695) );
  OR U325 ( .A(n14995), .B(n14996), .Z(n14994) );
  OR U326 ( .A(n15322), .B(n15323), .Z(n15321) );
  OR U327 ( .A(n15856), .B(n15857), .Z(n15855) );
  OR U328 ( .A(n16239), .B(n16240), .Z(n16238) );
  IV U329 ( .A(n16638), .Z(n3) );
  IV U330 ( .A(B[100]), .Z(n4) );
  IV U331 ( .A(n51829), .Z(n5) );
  IV U332 ( .A(B[99]), .Z(n6) );
  IV U333 ( .A(n52036), .Z(n7) );
  IV U334 ( .A(n52044), .Z(n8) );
  IV U335 ( .A(B[97]), .Z(n9) );
  IV U336 ( .A(n52052), .Z(n10) );
  IV U337 ( .A(B[96]), .Z(n11) );
  IV U338 ( .A(n52060), .Z(n12) );
  IV U339 ( .A(B[95]), .Z(n13) );
  IV U340 ( .A(n52068), .Z(n14) );
  IV U341 ( .A(B[94]), .Z(n15) );
  IV U342 ( .A(n52076), .Z(n16) );
  IV U343 ( .A(B[93]), .Z(n17) );
  IV U344 ( .A(n52084), .Z(n18) );
  IV U345 ( .A(B[92]), .Z(n19) );
  IV U346 ( .A(n52092), .Z(n20) );
  IV U347 ( .A(B[91]), .Z(n21) );
  IV U348 ( .A(n52100), .Z(n22) );
  IV U349 ( .A(B[90]), .Z(n23) );
  IV U350 ( .A(n52108), .Z(n24) );
  IV U351 ( .A(B[89]), .Z(n25) );
  IV U352 ( .A(n52116), .Z(n26) );
  IV U353 ( .A(B[88]), .Z(n27) );
  IV U354 ( .A(n52124), .Z(n28) );
  IV U355 ( .A(B[87]), .Z(n29) );
  IV U356 ( .A(n52132), .Z(n30) );
  IV U357 ( .A(B[86]), .Z(n31) );
  IV U358 ( .A(n52140), .Z(n32) );
  IV U359 ( .A(B[85]), .Z(n33) );
  IV U360 ( .A(n52148), .Z(n34) );
  IV U361 ( .A(n52156), .Z(n35) );
  IV U362 ( .A(n52164), .Z(n36) );
  IV U363 ( .A(n52172), .Z(n37) );
  IV U364 ( .A(n52180), .Z(n38) );
  IV U365 ( .A(n52188), .Z(n39) );
  IV U366 ( .A(n52196), .Z(n40) );
  IV U367 ( .A(n52204), .Z(n41) );
  IV U368 ( .A(n52212), .Z(n42) );
  IV U369 ( .A(n52220), .Z(n43) );
  IV U370 ( .A(n52228), .Z(n44) );
  IV U371 ( .A(n52236), .Z(n45) );
  IV U372 ( .A(n52336), .Z(n46) );
  IV U373 ( .A(n52244), .Z(n47) );
  IV U374 ( .A(n3904), .Z(n48) );
  IV U375 ( .A(n49313), .Z(n49) );
  IV U376 ( .A(n49328), .Z(n50) );
  IV U377 ( .A(n49343), .Z(n51) );
  IV U378 ( .A(n49358), .Z(n52) );
  IV U379 ( .A(n49378), .Z(n53) );
  IV U380 ( .A(A[31]), .Z(n54) );
  IV U381 ( .A(A[30]), .Z(n55) );
  IV U382 ( .A(A[29]), .Z(n56) );
  IV U383 ( .A(A[28]), .Z(n57) );
  IV U384 ( .A(A[27]), .Z(n58) );
  IV U385 ( .A(A[26]), .Z(n59) );
  IV U386 ( .A(A[25]), .Z(n60) );
  IV U387 ( .A(A[24]), .Z(n61) );
  IV U388 ( .A(A[23]), .Z(n62) );
  IV U389 ( .A(A[22]), .Z(n63) );
  IV U390 ( .A(A[21]), .Z(n64) );
  IV U391 ( .A(A[20]), .Z(n65) );
  IV U392 ( .A(A[19]), .Z(n66) );
  IV U393 ( .A(A[18]), .Z(n67) );
  IV U394 ( .A(A[17]), .Z(n68) );
  IV U395 ( .A(A[16]), .Z(n69) );
  IV U396 ( .A(A[15]), .Z(n70) );
  IV U397 ( .A(A[14]), .Z(n71) );
  IV U398 ( .A(A[13]), .Z(n72) );
  IV U399 ( .A(A[12]), .Z(n73) );
  IV U400 ( .A(A[11]), .Z(n74) );
  IV U401 ( .A(A[10]), .Z(n75) );
  IV U402 ( .A(A[9]), .Z(n76) );
  IV U403 ( .A(A[8]), .Z(n77) );
  IV U404 ( .A(A[7]), .Z(n78) );
  IV U405 ( .A(A[6]), .Z(n79) );
  IV U406 ( .A(A[5]), .Z(n80) );
  IV U407 ( .A(A[4]), .Z(n81) );
  IV U408 ( .A(A[3]), .Z(n82) );
  XNOR U409 ( .A(n84), .B(n85), .Z(PRODUCT[1]) );
  AND U410 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
  AND U411 ( .A(n86), .B(n87), .Z(\A2[99] ) );
  AND U412 ( .A(n88), .B(n89), .Z(\A2[98] ) );
  AND U413 ( .A(n90), .B(n91), .Z(\A2[97] ) );
  AND U414 ( .A(n92), .B(n93), .Z(\A2[96] ) );
  AND U415 ( .A(n94), .B(n95), .Z(\A2[95] ) );
  AND U416 ( .A(n96), .B(n97), .Z(\A2[94] ) );
  AND U417 ( .A(n98), .B(n99), .Z(\A2[93] ) );
  AND U418 ( .A(n100), .B(n101), .Z(\A2[92] ) );
  AND U419 ( .A(n102), .B(n103), .Z(\A2[91] ) );
  AND U420 ( .A(n104), .B(n105), .Z(\A2[90] ) );
  AND U421 ( .A(n106), .B(n107), .Z(\A2[89] ) );
  AND U422 ( .A(n108), .B(n109), .Z(\A2[88] ) );
  AND U423 ( .A(n110), .B(n111), .Z(\A2[87] ) );
  AND U424 ( .A(n112), .B(n113), .Z(\A2[86] ) );
  AND U425 ( .A(n114), .B(n115), .Z(\A2[85] ) );
  AND U426 ( .A(n116), .B(n117), .Z(\A2[84] ) );
  AND U427 ( .A(n118), .B(n119), .Z(\A2[83] ) );
  AND U428 ( .A(n120), .B(n121), .Z(\A2[82] ) );
  AND U429 ( .A(n122), .B(n123), .Z(\A2[81] ) );
  AND U430 ( .A(n124), .B(n125), .Z(\A2[80] ) );
  AND U431 ( .A(n126), .B(n127), .Z(\A2[79] ) );
  AND U432 ( .A(n128), .B(n129), .Z(\A2[78] ) );
  AND U433 ( .A(n130), .B(n131), .Z(\A2[77] ) );
  AND U434 ( .A(n132), .B(n133), .Z(\A2[76] ) );
  AND U435 ( .A(n134), .B(n135), .Z(\A2[75] ) );
  AND U436 ( .A(n136), .B(n137), .Z(\A2[74] ) );
  AND U437 ( .A(n138), .B(n139), .Z(\A2[73] ) );
  AND U438 ( .A(n140), .B(n141), .Z(\A2[72] ) );
  AND U439 ( .A(n142), .B(n143), .Z(\A2[71] ) );
  AND U440 ( .A(n144), .B(n145), .Z(\A2[70] ) );
  AND U441 ( .A(n146), .B(n147), .Z(\A2[69] ) );
  AND U442 ( .A(n148), .B(n149), .Z(\A2[68] ) );
  AND U443 ( .A(n150), .B(n151), .Z(\A2[67] ) );
  AND U444 ( .A(n152), .B(n153), .Z(\A2[66] ) );
  AND U445 ( .A(n154), .B(n155), .Z(\A2[65] ) );
  AND U446 ( .A(n156), .B(n157), .Z(\A2[64] ) );
  AND U447 ( .A(n158), .B(n159), .Z(\A2[63] ) );
  AND U448 ( .A(n160), .B(n161), .Z(\A2[62] ) );
  AND U449 ( .A(n162), .B(n163), .Z(\A2[61] ) );
  AND U450 ( .A(n164), .B(n165), .Z(\A2[60] ) );
  AND U451 ( .A(n166), .B(n167), .Z(\A2[59] ) );
  AND U452 ( .A(n168), .B(n169), .Z(\A2[58] ) );
  AND U453 ( .A(n170), .B(n171), .Z(\A2[57] ) );
  AND U454 ( .A(n172), .B(n173), .Z(\A2[56] ) );
  AND U455 ( .A(n174), .B(n175), .Z(\A2[55] ) );
  AND U456 ( .A(n176), .B(n177), .Z(\A2[54] ) );
  AND U457 ( .A(n178), .B(n179), .Z(\A2[53] ) );
  AND U458 ( .A(n180), .B(n181), .Z(\A2[52] ) );
  AND U459 ( .A(n182), .B(n183), .Z(\A2[51] ) );
  AND U460 ( .A(n184), .B(n185), .Z(\A2[50] ) );
  AND U461 ( .A(n186), .B(n187), .Z(\A2[49] ) );
  AND U462 ( .A(n188), .B(n189), .Z(\A2[48] ) );
  AND U463 ( .A(n190), .B(n191), .Z(\A2[47] ) );
  AND U464 ( .A(n192), .B(n193), .Z(\A2[46] ) );
  AND U465 ( .A(n194), .B(n195), .Z(\A2[45] ) );
  AND U466 ( .A(n196), .B(n197), .Z(\A2[44] ) );
  AND U467 ( .A(n198), .B(n199), .Z(\A2[43] ) );
  AND U468 ( .A(n200), .B(n201), .Z(\A2[42] ) );
  AND U469 ( .A(n202), .B(n203), .Z(\A2[41] ) );
  AND U470 ( .A(n204), .B(n205), .Z(\A2[40] ) );
  AND U471 ( .A(n206), .B(n207), .Z(\A2[39] ) );
  AND U472 ( .A(n208), .B(n209), .Z(\A2[38] ) );
  AND U473 ( .A(n210), .B(n211), .Z(\A2[37] ) );
  AND U474 ( .A(n212), .B(n213), .Z(\A2[36] ) );
  AND U475 ( .A(n214), .B(n215), .Z(\A2[35] ) );
  AND U476 ( .A(n216), .B(n217), .Z(\A2[34] ) );
  AND U477 ( .A(n218), .B(n219), .Z(\A2[33] ) );
  AND U478 ( .A(n220), .B(n221), .Z(\A2[32] ) );
  AND U479 ( .A(n222), .B(n223), .Z(\A2[31] ) );
  AND U480 ( .A(n224), .B(A[31]), .Z(\A2[285] ) );
  AND U481 ( .A(n225), .B(n226), .Z(\A2[284] ) );
  AND U482 ( .A(n227), .B(n228), .Z(\A2[283] ) );
  AND U483 ( .A(n229), .B(n230), .Z(\A2[282] ) );
  AND U484 ( .A(n231), .B(n232), .Z(\A2[281] ) );
  AND U485 ( .A(n233), .B(n234), .Z(\A2[280] ) );
  AND U486 ( .A(n235), .B(n236), .Z(\A2[279] ) );
  AND U487 ( .A(n237), .B(n238), .Z(\A2[278] ) );
  AND U488 ( .A(n239), .B(n240), .Z(\A2[277] ) );
  AND U489 ( .A(n241), .B(n242), .Z(\A2[276] ) );
  AND U490 ( .A(n243), .B(n244), .Z(\A2[275] ) );
  AND U491 ( .A(n245), .B(n246), .Z(\A2[274] ) );
  AND U492 ( .A(n247), .B(n248), .Z(\A2[273] ) );
  AND U493 ( .A(n249), .B(n250), .Z(\A2[272] ) );
  AND U494 ( .A(n251), .B(n252), .Z(\A2[271] ) );
  AND U495 ( .A(n253), .B(n254), .Z(\A2[270] ) );
  AND U496 ( .A(n255), .B(n256), .Z(\A2[269] ) );
  AND U497 ( .A(n257), .B(n258), .Z(\A2[268] ) );
  AND U498 ( .A(n259), .B(n260), .Z(\A2[267] ) );
  AND U499 ( .A(n261), .B(n262), .Z(\A2[266] ) );
  AND U500 ( .A(n263), .B(n264), .Z(\A2[265] ) );
  AND U501 ( .A(n265), .B(n266), .Z(\A2[264] ) );
  AND U502 ( .A(n267), .B(n268), .Z(\A2[263] ) );
  AND U503 ( .A(n269), .B(n270), .Z(\A2[262] ) );
  AND U504 ( .A(n271), .B(n272), .Z(\A2[261] ) );
  AND U505 ( .A(n273), .B(n274), .Z(\A2[260] ) );
  AND U506 ( .A(n275), .B(n276), .Z(\A2[259] ) );
  AND U507 ( .A(n277), .B(n278), .Z(\A2[258] ) );
  AND U508 ( .A(n279), .B(n280), .Z(\A2[257] ) );
  AND U509 ( .A(n281), .B(n282), .Z(\A2[256] ) );
  AND U510 ( .A(n283), .B(n284), .Z(\A2[255] ) );
  AND U511 ( .A(n285), .B(n286), .Z(\A2[254] ) );
  AND U512 ( .A(n287), .B(n288), .Z(\A2[253] ) );
  AND U513 ( .A(n289), .B(n290), .Z(\A2[252] ) );
  AND U514 ( .A(n291), .B(n292), .Z(\A2[251] ) );
  AND U515 ( .A(n293), .B(n294), .Z(\A2[250] ) );
  AND U516 ( .A(n295), .B(n296), .Z(\A2[249] ) );
  AND U517 ( .A(n297), .B(n298), .Z(\A2[248] ) );
  AND U518 ( .A(n299), .B(n300), .Z(\A2[247] ) );
  AND U519 ( .A(n301), .B(n302), .Z(\A2[246] ) );
  AND U520 ( .A(n303), .B(n304), .Z(\A2[245] ) );
  AND U521 ( .A(n305), .B(n306), .Z(\A2[244] ) );
  AND U522 ( .A(n307), .B(n308), .Z(\A2[243] ) );
  AND U523 ( .A(n309), .B(n310), .Z(\A2[242] ) );
  AND U524 ( .A(n311), .B(n312), .Z(\A2[241] ) );
  AND U525 ( .A(n313), .B(n314), .Z(\A2[240] ) );
  AND U526 ( .A(n315), .B(n316), .Z(\A2[239] ) );
  AND U527 ( .A(n317), .B(n318), .Z(\A2[238] ) );
  AND U528 ( .A(n319), .B(n320), .Z(\A2[237] ) );
  AND U529 ( .A(n321), .B(n322), .Z(\A2[236] ) );
  AND U530 ( .A(n323), .B(n324), .Z(\A2[235] ) );
  AND U531 ( .A(n325), .B(n326), .Z(\A2[234] ) );
  AND U532 ( .A(n327), .B(n328), .Z(\A2[233] ) );
  AND U533 ( .A(n329), .B(n330), .Z(\A2[232] ) );
  AND U534 ( .A(n331), .B(n332), .Z(\A2[231] ) );
  AND U535 ( .A(n333), .B(n334), .Z(\A2[230] ) );
  AND U536 ( .A(n335), .B(n336), .Z(\A2[229] ) );
  AND U537 ( .A(n337), .B(n338), .Z(\A2[228] ) );
  AND U538 ( .A(n339), .B(n340), .Z(\A2[227] ) );
  AND U539 ( .A(n341), .B(n342), .Z(\A2[226] ) );
  AND U540 ( .A(n343), .B(n344), .Z(\A2[225] ) );
  AND U541 ( .A(n345), .B(n346), .Z(\A2[224] ) );
  AND U542 ( .A(n347), .B(n348), .Z(\A2[223] ) );
  AND U543 ( .A(n349), .B(n350), .Z(\A2[222] ) );
  AND U544 ( .A(n351), .B(n352), .Z(\A2[221] ) );
  AND U545 ( .A(n353), .B(n354), .Z(\A2[220] ) );
  AND U546 ( .A(n355), .B(n356), .Z(\A2[219] ) );
  AND U547 ( .A(n357), .B(n358), .Z(\A2[218] ) );
  AND U548 ( .A(n359), .B(n360), .Z(\A2[217] ) );
  AND U549 ( .A(n361), .B(n362), .Z(\A2[216] ) );
  AND U550 ( .A(n363), .B(n364), .Z(\A2[215] ) );
  AND U551 ( .A(n365), .B(n366), .Z(\A2[214] ) );
  AND U552 ( .A(n367), .B(n368), .Z(\A2[213] ) );
  AND U553 ( .A(n369), .B(n370), .Z(\A2[212] ) );
  AND U554 ( .A(n371), .B(n372), .Z(\A2[211] ) );
  AND U555 ( .A(n373), .B(n374), .Z(\A2[210] ) );
  AND U556 ( .A(n375), .B(n376), .Z(\A2[209] ) );
  AND U557 ( .A(n377), .B(n378), .Z(\A2[208] ) );
  AND U558 ( .A(n379), .B(n380), .Z(\A2[207] ) );
  AND U559 ( .A(n381), .B(n382), .Z(\A2[206] ) );
  AND U560 ( .A(n383), .B(n384), .Z(\A2[205] ) );
  AND U561 ( .A(n385), .B(n386), .Z(\A2[204] ) );
  AND U562 ( .A(n387), .B(n388), .Z(\A2[203] ) );
  AND U563 ( .A(n389), .B(n390), .Z(\A2[202] ) );
  AND U564 ( .A(n391), .B(n392), .Z(\A2[201] ) );
  AND U565 ( .A(n393), .B(n394), .Z(\A2[200] ) );
  AND U566 ( .A(n395), .B(n396), .Z(\A2[199] ) );
  AND U567 ( .A(n397), .B(n398), .Z(\A2[198] ) );
  AND U568 ( .A(n399), .B(n400), .Z(\A2[197] ) );
  AND U569 ( .A(n401), .B(n402), .Z(\A2[196] ) );
  AND U570 ( .A(n403), .B(n404), .Z(\A2[195] ) );
  AND U571 ( .A(n405), .B(n406), .Z(\A2[194] ) );
  AND U572 ( .A(n407), .B(n408), .Z(\A2[193] ) );
  AND U573 ( .A(n409), .B(n410), .Z(\A2[192] ) );
  AND U574 ( .A(n411), .B(n412), .Z(\A2[191] ) );
  AND U575 ( .A(n413), .B(n414), .Z(\A2[190] ) );
  AND U576 ( .A(n415), .B(n416), .Z(\A2[189] ) );
  AND U577 ( .A(n417), .B(n418), .Z(\A2[188] ) );
  AND U578 ( .A(n419), .B(n420), .Z(\A2[187] ) );
  AND U579 ( .A(n421), .B(n422), .Z(\A2[186] ) );
  AND U580 ( .A(n423), .B(n424), .Z(\A2[185] ) );
  AND U581 ( .A(n425), .B(n426), .Z(\A2[184] ) );
  AND U582 ( .A(n427), .B(n428), .Z(\A2[183] ) );
  AND U583 ( .A(n429), .B(n430), .Z(\A2[182] ) );
  AND U584 ( .A(n431), .B(n432), .Z(\A2[181] ) );
  AND U585 ( .A(n433), .B(n434), .Z(\A2[180] ) );
  AND U586 ( .A(n435), .B(n436), .Z(\A2[179] ) );
  AND U587 ( .A(n437), .B(n438), .Z(\A2[178] ) );
  AND U588 ( .A(n439), .B(n440), .Z(\A2[177] ) );
  AND U589 ( .A(n441), .B(n442), .Z(\A2[176] ) );
  AND U590 ( .A(n443), .B(n444), .Z(\A2[175] ) );
  AND U591 ( .A(n445), .B(n446), .Z(\A2[174] ) );
  AND U592 ( .A(n447), .B(n448), .Z(\A2[173] ) );
  AND U593 ( .A(n449), .B(n450), .Z(\A2[172] ) );
  AND U594 ( .A(n451), .B(n452), .Z(\A2[171] ) );
  AND U595 ( .A(n453), .B(n454), .Z(\A2[170] ) );
  AND U596 ( .A(n455), .B(n456), .Z(\A2[169] ) );
  AND U597 ( .A(n457), .B(n458), .Z(\A2[168] ) );
  AND U598 ( .A(n459), .B(n460), .Z(\A2[167] ) );
  AND U599 ( .A(n461), .B(n462), .Z(\A2[166] ) );
  AND U600 ( .A(n463), .B(n464), .Z(\A2[165] ) );
  AND U601 ( .A(n465), .B(n466), .Z(\A2[164] ) );
  AND U602 ( .A(n467), .B(n468), .Z(\A2[163] ) );
  AND U603 ( .A(n469), .B(n470), .Z(\A2[162] ) );
  AND U604 ( .A(n471), .B(n472), .Z(\A2[161] ) );
  AND U605 ( .A(n473), .B(n474), .Z(\A2[160] ) );
  AND U606 ( .A(n475), .B(n476), .Z(\A2[159] ) );
  AND U607 ( .A(n477), .B(n478), .Z(\A2[158] ) );
  AND U608 ( .A(n479), .B(n480), .Z(\A2[157] ) );
  AND U609 ( .A(n481), .B(n482), .Z(\A2[156] ) );
  AND U610 ( .A(n483), .B(n484), .Z(\A2[155] ) );
  AND U611 ( .A(n485), .B(n486), .Z(\A2[154] ) );
  AND U612 ( .A(n487), .B(n488), .Z(\A2[153] ) );
  AND U613 ( .A(n489), .B(n490), .Z(\A2[152] ) );
  AND U614 ( .A(n491), .B(n492), .Z(\A2[151] ) );
  AND U615 ( .A(n493), .B(n494), .Z(\A2[150] ) );
  AND U616 ( .A(n495), .B(n496), .Z(\A2[149] ) );
  AND U617 ( .A(n497), .B(n498), .Z(\A2[148] ) );
  AND U618 ( .A(n499), .B(n500), .Z(\A2[147] ) );
  AND U619 ( .A(n501), .B(n502), .Z(\A2[146] ) );
  AND U620 ( .A(n503), .B(n504), .Z(\A2[145] ) );
  AND U621 ( .A(n505), .B(n506), .Z(\A2[144] ) );
  AND U622 ( .A(n507), .B(n508), .Z(\A2[143] ) );
  AND U623 ( .A(n509), .B(n510), .Z(\A2[142] ) );
  AND U624 ( .A(n511), .B(n512), .Z(\A2[141] ) );
  AND U625 ( .A(n513), .B(n514), .Z(\A2[140] ) );
  AND U626 ( .A(n515), .B(n516), .Z(\A2[139] ) );
  AND U627 ( .A(n517), .B(n518), .Z(\A2[138] ) );
  AND U628 ( .A(n519), .B(n520), .Z(\A2[137] ) );
  AND U629 ( .A(n521), .B(n522), .Z(\A2[136] ) );
  AND U630 ( .A(n523), .B(n524), .Z(\A2[135] ) );
  AND U631 ( .A(n525), .B(n526), .Z(\A2[134] ) );
  AND U632 ( .A(n527), .B(n528), .Z(\A2[133] ) );
  AND U633 ( .A(n529), .B(n530), .Z(\A2[132] ) );
  AND U634 ( .A(n531), .B(n532), .Z(\A2[131] ) );
  AND U635 ( .A(n533), .B(n534), .Z(\A2[130] ) );
  AND U636 ( .A(n535), .B(n536), .Z(\A2[129] ) );
  AND U637 ( .A(n537), .B(n538), .Z(\A2[128] ) );
  AND U638 ( .A(n539), .B(n540), .Z(\A2[127] ) );
  AND U639 ( .A(n541), .B(n542), .Z(\A2[126] ) );
  AND U640 ( .A(n543), .B(n544), .Z(\A2[125] ) );
  AND U641 ( .A(n545), .B(n546), .Z(\A2[124] ) );
  AND U642 ( .A(n547), .B(n548), .Z(\A2[123] ) );
  AND U643 ( .A(n549), .B(n550), .Z(\A2[122] ) );
  AND U644 ( .A(n551), .B(n552), .Z(\A2[121] ) );
  AND U645 ( .A(n553), .B(n554), .Z(\A2[120] ) );
  AND U646 ( .A(n555), .B(n556), .Z(\A2[119] ) );
  AND U647 ( .A(n557), .B(n558), .Z(\A2[118] ) );
  AND U648 ( .A(n559), .B(n560), .Z(\A2[117] ) );
  AND U649 ( .A(n561), .B(n562), .Z(\A2[116] ) );
  AND U650 ( .A(n563), .B(n564), .Z(\A2[115] ) );
  AND U651 ( .A(n565), .B(n566), .Z(\A2[114] ) );
  AND U652 ( .A(n567), .B(n568), .Z(\A2[113] ) );
  AND U653 ( .A(n569), .B(n570), .Z(\A2[112] ) );
  AND U654 ( .A(n571), .B(n572), .Z(\A2[111] ) );
  AND U655 ( .A(n573), .B(n574), .Z(\A2[110] ) );
  AND U656 ( .A(n575), .B(n576), .Z(\A2[109] ) );
  AND U657 ( .A(n577), .B(n578), .Z(\A2[108] ) );
  AND U658 ( .A(n579), .B(n580), .Z(\A2[107] ) );
  AND U659 ( .A(n581), .B(n582), .Z(\A2[106] ) );
  AND U660 ( .A(n583), .B(n584), .Z(\A2[105] ) );
  AND U661 ( .A(n585), .B(n586), .Z(\A2[104] ) );
  AND U662 ( .A(n587), .B(n588), .Z(\A2[103] ) );
  AND U663 ( .A(n589), .B(n590), .Z(\A2[102] ) );
  AND U664 ( .A(n591), .B(n592), .Z(\A2[101] ) );
  AND U665 ( .A(n593), .B(n594), .Z(\A2[100] ) );
  XOR U666 ( .A(n595), .B(n596), .Z(\A1[9] ) );
  XNOR U667 ( .A(n597), .B(n49), .Z(n596) );
  XOR U668 ( .A(n594), .B(n593), .Z(\A1[99] ) );
  XOR U669 ( .A(n598), .B(n599), .Z(n593) );
  XNOR U670 ( .A(n600), .B(n5), .Z(n599) );
  NAND U671 ( .A(n601), .B(n602), .Z(n594) );
  NANDN U672 ( .A(n603), .B(n604), .Z(n602) );
  NANDN U673 ( .A(n605), .B(n606), .Z(n604) );
  XOR U674 ( .A(n87), .B(n86), .Z(\A1[98] ) );
  XNOR U675 ( .A(n603), .B(n607), .Z(n86) );
  XNOR U676 ( .A(n605), .B(n606), .Z(n607) );
  AND U677 ( .A(n608), .B(n609), .Z(n606) );
  NAND U678 ( .A(n610), .B(n611), .Z(n609) );
  NANDN U679 ( .A(n612), .B(n613), .Z(n610) );
  ANDN U680 ( .B(B[69]), .A(n54), .Z(n605) );
  XOR U681 ( .A(n614), .B(n615), .Z(n603) );
  XOR U682 ( .A(n616), .B(n617), .Z(n615) );
  NAND U683 ( .A(n618), .B(n619), .Z(n87) );
  NANDN U684 ( .A(n620), .B(n621), .Z(n619) );
  OR U685 ( .A(n622), .B(n623), .Z(n621) );
  NAND U686 ( .A(n623), .B(n622), .Z(n618) );
  XOR U687 ( .A(n89), .B(n88), .Z(\A1[97] ) );
  XOR U688 ( .A(n623), .B(n624), .Z(n88) );
  XNOR U689 ( .A(n622), .B(n620), .Z(n624) );
  AND U690 ( .A(n625), .B(n626), .Z(n620) );
  NANDN U691 ( .A(n627), .B(n628), .Z(n626) );
  NANDN U692 ( .A(n629), .B(n630), .Z(n628) );
  NANDN U693 ( .A(n630), .B(n629), .Z(n625) );
  ANDN U694 ( .B(B[68]), .A(n54), .Z(n622) );
  XOR U695 ( .A(n611), .B(n631), .Z(n623) );
  XNOR U696 ( .A(n612), .B(n613), .Z(n631) );
  AND U697 ( .A(n632), .B(n633), .Z(n613) );
  NANDN U698 ( .A(n634), .B(n635), .Z(n633) );
  NANDN U699 ( .A(n636), .B(n637), .Z(n635) );
  ANDN U700 ( .B(B[69]), .A(n55), .Z(n612) );
  XOR U701 ( .A(n638), .B(n639), .Z(n611) );
  XNOR U702 ( .A(n640), .B(n7), .Z(n639) );
  NAND U703 ( .A(n641), .B(n642), .Z(n89) );
  NANDN U704 ( .A(n643), .B(n644), .Z(n642) );
  OR U705 ( .A(n645), .B(n646), .Z(n644) );
  NAND U706 ( .A(n646), .B(n645), .Z(n641) );
  XOR U707 ( .A(n91), .B(n90), .Z(\A1[96] ) );
  XOR U708 ( .A(n646), .B(n647), .Z(n90) );
  XNOR U709 ( .A(n645), .B(n643), .Z(n647) );
  AND U710 ( .A(n648), .B(n649), .Z(n643) );
  NANDN U711 ( .A(n650), .B(n651), .Z(n649) );
  NANDN U712 ( .A(n652), .B(n653), .Z(n651) );
  NANDN U713 ( .A(n653), .B(n652), .Z(n648) );
  ANDN U714 ( .B(B[67]), .A(n54), .Z(n645) );
  XNOR U715 ( .A(n630), .B(n654), .Z(n646) );
  XNOR U716 ( .A(n629), .B(n627), .Z(n654) );
  AND U717 ( .A(n655), .B(n656), .Z(n627) );
  NANDN U718 ( .A(n657), .B(n658), .Z(n656) );
  OR U719 ( .A(n659), .B(n660), .Z(n658) );
  NAND U720 ( .A(n660), .B(n659), .Z(n655) );
  ANDN U721 ( .B(B[68]), .A(n55), .Z(n629) );
  XOR U722 ( .A(n634), .B(n661), .Z(n630) );
  XNOR U723 ( .A(n636), .B(n637), .Z(n661) );
  AND U724 ( .A(n662), .B(n663), .Z(n637) );
  NAND U725 ( .A(n664), .B(n665), .Z(n663) );
  NANDN U726 ( .A(n666), .B(n667), .Z(n664) );
  ANDN U727 ( .B(B[69]), .A(n56), .Z(n636) );
  XNOR U728 ( .A(n668), .B(n669), .Z(n634) );
  XNOR U729 ( .A(n670), .B(n8), .Z(n669) );
  NAND U730 ( .A(n671), .B(n672), .Z(n91) );
  NANDN U731 ( .A(n673), .B(n674), .Z(n672) );
  OR U732 ( .A(n675), .B(n676), .Z(n674) );
  NAND U733 ( .A(n676), .B(n675), .Z(n671) );
  XOR U734 ( .A(n93), .B(n92), .Z(\A1[95] ) );
  XOR U735 ( .A(n676), .B(n677), .Z(n92) );
  XNOR U736 ( .A(n675), .B(n673), .Z(n677) );
  AND U737 ( .A(n678), .B(n679), .Z(n673) );
  NANDN U738 ( .A(n680), .B(n681), .Z(n679) );
  NANDN U739 ( .A(n682), .B(n683), .Z(n681) );
  NANDN U740 ( .A(n683), .B(n682), .Z(n678) );
  ANDN U741 ( .B(B[66]), .A(n54), .Z(n675) );
  XNOR U742 ( .A(n653), .B(n684), .Z(n676) );
  XNOR U743 ( .A(n652), .B(n650), .Z(n684) );
  AND U744 ( .A(n685), .B(n686), .Z(n650) );
  NANDN U745 ( .A(n687), .B(n688), .Z(n686) );
  OR U746 ( .A(n689), .B(n690), .Z(n688) );
  NAND U747 ( .A(n690), .B(n689), .Z(n685) );
  ANDN U748 ( .B(B[67]), .A(n55), .Z(n652) );
  XNOR U749 ( .A(n660), .B(n691), .Z(n653) );
  XNOR U750 ( .A(n659), .B(n657), .Z(n691) );
  AND U751 ( .A(n692), .B(n693), .Z(n657) );
  NANDN U752 ( .A(n694), .B(n695), .Z(n693) );
  NANDN U753 ( .A(n696), .B(n697), .Z(n695) );
  NANDN U754 ( .A(n697), .B(n696), .Z(n692) );
  ANDN U755 ( .B(B[68]), .A(n56), .Z(n659) );
  XOR U756 ( .A(n665), .B(n698), .Z(n660) );
  XNOR U757 ( .A(n666), .B(n667), .Z(n698) );
  AND U758 ( .A(n699), .B(n700), .Z(n667) );
  NANDN U759 ( .A(n701), .B(n702), .Z(n700) );
  NANDN U760 ( .A(n703), .B(n704), .Z(n702) );
  ANDN U761 ( .B(B[69]), .A(n57), .Z(n666) );
  XOR U762 ( .A(n705), .B(n706), .Z(n665) );
  XNOR U763 ( .A(n707), .B(n10), .Z(n706) );
  NAND U764 ( .A(n708), .B(n709), .Z(n93) );
  NANDN U765 ( .A(n710), .B(n711), .Z(n709) );
  OR U766 ( .A(n712), .B(n713), .Z(n711) );
  NAND U767 ( .A(n713), .B(n712), .Z(n708) );
  XOR U768 ( .A(n95), .B(n94), .Z(\A1[94] ) );
  XOR U769 ( .A(n713), .B(n714), .Z(n94) );
  XNOR U770 ( .A(n712), .B(n710), .Z(n714) );
  AND U771 ( .A(n715), .B(n716), .Z(n710) );
  NANDN U772 ( .A(n717), .B(n718), .Z(n716) );
  NANDN U773 ( .A(n719), .B(n720), .Z(n718) );
  NANDN U774 ( .A(n720), .B(n719), .Z(n715) );
  ANDN U775 ( .B(B[65]), .A(n54), .Z(n712) );
  XNOR U776 ( .A(n683), .B(n721), .Z(n713) );
  XNOR U777 ( .A(n682), .B(n680), .Z(n721) );
  AND U778 ( .A(n722), .B(n723), .Z(n680) );
  NANDN U779 ( .A(n724), .B(n725), .Z(n723) );
  OR U780 ( .A(n726), .B(n727), .Z(n725) );
  NAND U781 ( .A(n727), .B(n726), .Z(n722) );
  ANDN U782 ( .B(B[66]), .A(n55), .Z(n682) );
  XNOR U783 ( .A(n690), .B(n728), .Z(n683) );
  XNOR U784 ( .A(n689), .B(n687), .Z(n728) );
  AND U785 ( .A(n729), .B(n730), .Z(n687) );
  NANDN U786 ( .A(n731), .B(n732), .Z(n730) );
  NANDN U787 ( .A(n733), .B(n734), .Z(n732) );
  NANDN U788 ( .A(n734), .B(n733), .Z(n729) );
  ANDN U789 ( .B(B[67]), .A(n56), .Z(n689) );
  XNOR U790 ( .A(n697), .B(n735), .Z(n690) );
  XNOR U791 ( .A(n696), .B(n694), .Z(n735) );
  AND U792 ( .A(n736), .B(n737), .Z(n694) );
  NANDN U793 ( .A(n738), .B(n739), .Z(n737) );
  OR U794 ( .A(n740), .B(n741), .Z(n739) );
  NAND U795 ( .A(n741), .B(n740), .Z(n736) );
  ANDN U796 ( .B(B[68]), .A(n57), .Z(n696) );
  XOR U797 ( .A(n701), .B(n742), .Z(n697) );
  XNOR U798 ( .A(n703), .B(n704), .Z(n742) );
  AND U799 ( .A(n743), .B(n744), .Z(n704) );
  NAND U800 ( .A(n745), .B(n746), .Z(n744) );
  NANDN U801 ( .A(n747), .B(n748), .Z(n745) );
  ANDN U802 ( .B(B[69]), .A(n58), .Z(n703) );
  XNOR U803 ( .A(n749), .B(n750), .Z(n701) );
  XNOR U804 ( .A(n751), .B(n12), .Z(n750) );
  NAND U805 ( .A(n752), .B(n753), .Z(n95) );
  NANDN U806 ( .A(n754), .B(n755), .Z(n753) );
  OR U807 ( .A(n756), .B(n757), .Z(n755) );
  NAND U808 ( .A(n757), .B(n756), .Z(n752) );
  XOR U809 ( .A(n97), .B(n96), .Z(\A1[93] ) );
  XOR U810 ( .A(n757), .B(n758), .Z(n96) );
  XNOR U811 ( .A(n756), .B(n754), .Z(n758) );
  AND U812 ( .A(n759), .B(n760), .Z(n754) );
  NANDN U813 ( .A(n761), .B(n762), .Z(n760) );
  NANDN U814 ( .A(n763), .B(n764), .Z(n762) );
  NANDN U815 ( .A(n764), .B(n763), .Z(n759) );
  ANDN U816 ( .B(B[64]), .A(n54), .Z(n756) );
  XNOR U817 ( .A(n720), .B(n765), .Z(n757) );
  XNOR U818 ( .A(n719), .B(n717), .Z(n765) );
  AND U819 ( .A(n766), .B(n767), .Z(n717) );
  NANDN U820 ( .A(n768), .B(n769), .Z(n767) );
  OR U821 ( .A(n770), .B(n771), .Z(n769) );
  NAND U822 ( .A(n771), .B(n770), .Z(n766) );
  ANDN U823 ( .B(B[65]), .A(n55), .Z(n719) );
  XNOR U824 ( .A(n727), .B(n772), .Z(n720) );
  XNOR U825 ( .A(n726), .B(n724), .Z(n772) );
  AND U826 ( .A(n773), .B(n774), .Z(n724) );
  NANDN U827 ( .A(n775), .B(n776), .Z(n774) );
  NANDN U828 ( .A(n777), .B(n778), .Z(n776) );
  NANDN U829 ( .A(n778), .B(n777), .Z(n773) );
  ANDN U830 ( .B(B[66]), .A(n56), .Z(n726) );
  XNOR U831 ( .A(n734), .B(n779), .Z(n727) );
  XNOR U832 ( .A(n733), .B(n731), .Z(n779) );
  AND U833 ( .A(n780), .B(n781), .Z(n731) );
  NANDN U834 ( .A(n782), .B(n783), .Z(n781) );
  OR U835 ( .A(n784), .B(n785), .Z(n783) );
  NAND U836 ( .A(n785), .B(n784), .Z(n780) );
  ANDN U837 ( .B(B[67]), .A(n57), .Z(n733) );
  XNOR U838 ( .A(n741), .B(n786), .Z(n734) );
  XNOR U839 ( .A(n740), .B(n738), .Z(n786) );
  AND U840 ( .A(n787), .B(n788), .Z(n738) );
  NANDN U841 ( .A(n789), .B(n790), .Z(n788) );
  NANDN U842 ( .A(n791), .B(n792), .Z(n790) );
  NANDN U843 ( .A(n792), .B(n791), .Z(n787) );
  ANDN U844 ( .B(B[68]), .A(n58), .Z(n740) );
  XOR U845 ( .A(n746), .B(n793), .Z(n741) );
  XNOR U846 ( .A(n747), .B(n748), .Z(n793) );
  AND U847 ( .A(n794), .B(n795), .Z(n748) );
  NANDN U848 ( .A(n796), .B(n797), .Z(n795) );
  NANDN U849 ( .A(n798), .B(n799), .Z(n797) );
  ANDN U850 ( .B(B[69]), .A(n59), .Z(n747) );
  XOR U851 ( .A(n800), .B(n801), .Z(n746) );
  XNOR U852 ( .A(n802), .B(n14), .Z(n801) );
  NAND U853 ( .A(n803), .B(n804), .Z(n97) );
  NANDN U854 ( .A(n805), .B(n806), .Z(n804) );
  OR U855 ( .A(n807), .B(n808), .Z(n806) );
  NAND U856 ( .A(n808), .B(n807), .Z(n803) );
  XOR U857 ( .A(n99), .B(n98), .Z(\A1[92] ) );
  XOR U858 ( .A(n808), .B(n809), .Z(n98) );
  XNOR U859 ( .A(n807), .B(n805), .Z(n809) );
  AND U860 ( .A(n810), .B(n811), .Z(n805) );
  NANDN U861 ( .A(n812), .B(n813), .Z(n811) );
  NANDN U862 ( .A(n814), .B(n815), .Z(n813) );
  NANDN U863 ( .A(n815), .B(n814), .Z(n810) );
  ANDN U864 ( .B(B[63]), .A(n54), .Z(n807) );
  XNOR U865 ( .A(n764), .B(n816), .Z(n808) );
  XNOR U866 ( .A(n763), .B(n761), .Z(n816) );
  AND U867 ( .A(n817), .B(n818), .Z(n761) );
  NANDN U868 ( .A(n819), .B(n820), .Z(n818) );
  OR U869 ( .A(n821), .B(n822), .Z(n820) );
  NAND U870 ( .A(n822), .B(n821), .Z(n817) );
  ANDN U871 ( .B(B[64]), .A(n55), .Z(n763) );
  XNOR U872 ( .A(n771), .B(n823), .Z(n764) );
  XNOR U873 ( .A(n770), .B(n768), .Z(n823) );
  AND U874 ( .A(n824), .B(n825), .Z(n768) );
  NANDN U875 ( .A(n826), .B(n827), .Z(n825) );
  NANDN U876 ( .A(n828), .B(n829), .Z(n827) );
  NANDN U877 ( .A(n829), .B(n828), .Z(n824) );
  ANDN U878 ( .B(B[65]), .A(n56), .Z(n770) );
  XNOR U879 ( .A(n778), .B(n830), .Z(n771) );
  XNOR U880 ( .A(n777), .B(n775), .Z(n830) );
  AND U881 ( .A(n831), .B(n832), .Z(n775) );
  NANDN U882 ( .A(n833), .B(n834), .Z(n832) );
  OR U883 ( .A(n835), .B(n836), .Z(n834) );
  NAND U884 ( .A(n836), .B(n835), .Z(n831) );
  ANDN U885 ( .B(B[66]), .A(n57), .Z(n777) );
  XNOR U886 ( .A(n785), .B(n837), .Z(n778) );
  XNOR U887 ( .A(n784), .B(n782), .Z(n837) );
  AND U888 ( .A(n838), .B(n839), .Z(n782) );
  NANDN U889 ( .A(n840), .B(n841), .Z(n839) );
  NANDN U890 ( .A(n842), .B(n843), .Z(n841) );
  NANDN U891 ( .A(n843), .B(n842), .Z(n838) );
  ANDN U892 ( .B(B[67]), .A(n58), .Z(n784) );
  XNOR U893 ( .A(n792), .B(n844), .Z(n785) );
  XNOR U894 ( .A(n791), .B(n789), .Z(n844) );
  AND U895 ( .A(n845), .B(n846), .Z(n789) );
  NANDN U896 ( .A(n847), .B(n848), .Z(n846) );
  OR U897 ( .A(n849), .B(n850), .Z(n848) );
  NAND U898 ( .A(n850), .B(n849), .Z(n845) );
  ANDN U899 ( .B(B[68]), .A(n59), .Z(n791) );
  XOR U900 ( .A(n796), .B(n851), .Z(n792) );
  XNOR U901 ( .A(n798), .B(n799), .Z(n851) );
  AND U902 ( .A(n852), .B(n853), .Z(n799) );
  NAND U903 ( .A(n854), .B(n855), .Z(n853) );
  NANDN U904 ( .A(n856), .B(n857), .Z(n854) );
  ANDN U905 ( .B(B[69]), .A(n60), .Z(n798) );
  XNOR U906 ( .A(n858), .B(n859), .Z(n796) );
  XNOR U907 ( .A(n860), .B(n16), .Z(n859) );
  NAND U908 ( .A(n861), .B(n862), .Z(n99) );
  NANDN U909 ( .A(n863), .B(n864), .Z(n862) );
  OR U910 ( .A(n865), .B(n866), .Z(n864) );
  NAND U911 ( .A(n866), .B(n865), .Z(n861) );
  XOR U912 ( .A(n101), .B(n100), .Z(\A1[91] ) );
  XOR U913 ( .A(n866), .B(n867), .Z(n100) );
  XNOR U914 ( .A(n865), .B(n863), .Z(n867) );
  AND U915 ( .A(n868), .B(n869), .Z(n863) );
  NANDN U916 ( .A(n870), .B(n871), .Z(n869) );
  NANDN U917 ( .A(n872), .B(n873), .Z(n871) );
  NANDN U918 ( .A(n873), .B(n872), .Z(n868) );
  ANDN U919 ( .B(B[62]), .A(n54), .Z(n865) );
  XNOR U920 ( .A(n815), .B(n874), .Z(n866) );
  XNOR U921 ( .A(n814), .B(n812), .Z(n874) );
  AND U922 ( .A(n875), .B(n876), .Z(n812) );
  NANDN U923 ( .A(n877), .B(n878), .Z(n876) );
  OR U924 ( .A(n879), .B(n880), .Z(n878) );
  NAND U925 ( .A(n880), .B(n879), .Z(n875) );
  ANDN U926 ( .B(B[63]), .A(n55), .Z(n814) );
  XNOR U927 ( .A(n822), .B(n881), .Z(n815) );
  XNOR U928 ( .A(n821), .B(n819), .Z(n881) );
  AND U929 ( .A(n882), .B(n883), .Z(n819) );
  NANDN U930 ( .A(n884), .B(n885), .Z(n883) );
  NANDN U931 ( .A(n886), .B(n887), .Z(n885) );
  NANDN U932 ( .A(n887), .B(n886), .Z(n882) );
  ANDN U933 ( .B(B[64]), .A(n56), .Z(n821) );
  XNOR U934 ( .A(n829), .B(n888), .Z(n822) );
  XNOR U935 ( .A(n828), .B(n826), .Z(n888) );
  AND U936 ( .A(n889), .B(n890), .Z(n826) );
  NANDN U937 ( .A(n891), .B(n892), .Z(n890) );
  OR U938 ( .A(n893), .B(n894), .Z(n892) );
  NAND U939 ( .A(n894), .B(n893), .Z(n889) );
  ANDN U940 ( .B(B[65]), .A(n57), .Z(n828) );
  XNOR U941 ( .A(n836), .B(n895), .Z(n829) );
  XNOR U942 ( .A(n835), .B(n833), .Z(n895) );
  AND U943 ( .A(n896), .B(n897), .Z(n833) );
  NANDN U944 ( .A(n898), .B(n899), .Z(n897) );
  NANDN U945 ( .A(n900), .B(n901), .Z(n899) );
  NANDN U946 ( .A(n901), .B(n900), .Z(n896) );
  ANDN U947 ( .B(B[66]), .A(n58), .Z(n835) );
  XNOR U948 ( .A(n843), .B(n902), .Z(n836) );
  XNOR U949 ( .A(n842), .B(n840), .Z(n902) );
  AND U950 ( .A(n903), .B(n904), .Z(n840) );
  NANDN U951 ( .A(n905), .B(n906), .Z(n904) );
  OR U952 ( .A(n907), .B(n908), .Z(n906) );
  NAND U953 ( .A(n908), .B(n907), .Z(n903) );
  ANDN U954 ( .B(B[67]), .A(n59), .Z(n842) );
  XNOR U955 ( .A(n850), .B(n909), .Z(n843) );
  XNOR U956 ( .A(n849), .B(n847), .Z(n909) );
  AND U957 ( .A(n910), .B(n911), .Z(n847) );
  NANDN U958 ( .A(n912), .B(n913), .Z(n911) );
  NANDN U959 ( .A(n914), .B(n915), .Z(n913) );
  NANDN U960 ( .A(n915), .B(n914), .Z(n910) );
  ANDN U961 ( .B(B[68]), .A(n60), .Z(n849) );
  XOR U962 ( .A(n855), .B(n916), .Z(n850) );
  XNOR U963 ( .A(n856), .B(n857), .Z(n916) );
  AND U964 ( .A(n917), .B(n918), .Z(n857) );
  NANDN U965 ( .A(n919), .B(n920), .Z(n918) );
  NANDN U966 ( .A(n921), .B(n922), .Z(n920) );
  ANDN U967 ( .B(B[69]), .A(n61), .Z(n856) );
  XOR U968 ( .A(n923), .B(n924), .Z(n855) );
  XNOR U969 ( .A(n925), .B(n18), .Z(n924) );
  NAND U970 ( .A(n926), .B(n927), .Z(n101) );
  NANDN U971 ( .A(n928), .B(n929), .Z(n927) );
  OR U972 ( .A(n930), .B(n931), .Z(n929) );
  NAND U973 ( .A(n931), .B(n930), .Z(n926) );
  XOR U974 ( .A(n103), .B(n102), .Z(\A1[90] ) );
  XOR U975 ( .A(n931), .B(n932), .Z(n102) );
  XNOR U976 ( .A(n930), .B(n928), .Z(n932) );
  AND U977 ( .A(n933), .B(n934), .Z(n928) );
  NANDN U978 ( .A(n935), .B(n936), .Z(n934) );
  NANDN U979 ( .A(n937), .B(n938), .Z(n936) );
  NANDN U980 ( .A(n938), .B(n937), .Z(n933) );
  ANDN U981 ( .B(B[61]), .A(n54), .Z(n930) );
  XNOR U982 ( .A(n873), .B(n939), .Z(n931) );
  XNOR U983 ( .A(n872), .B(n870), .Z(n939) );
  AND U984 ( .A(n940), .B(n941), .Z(n870) );
  NANDN U985 ( .A(n942), .B(n943), .Z(n941) );
  OR U986 ( .A(n944), .B(n945), .Z(n943) );
  NAND U987 ( .A(n945), .B(n944), .Z(n940) );
  ANDN U988 ( .B(B[62]), .A(n55), .Z(n872) );
  XNOR U989 ( .A(n880), .B(n946), .Z(n873) );
  XNOR U990 ( .A(n879), .B(n877), .Z(n946) );
  AND U991 ( .A(n947), .B(n948), .Z(n877) );
  NANDN U992 ( .A(n949), .B(n950), .Z(n948) );
  NANDN U993 ( .A(n951), .B(n952), .Z(n950) );
  NANDN U994 ( .A(n952), .B(n951), .Z(n947) );
  ANDN U995 ( .B(B[63]), .A(n56), .Z(n879) );
  XNOR U996 ( .A(n887), .B(n953), .Z(n880) );
  XNOR U997 ( .A(n886), .B(n884), .Z(n953) );
  AND U998 ( .A(n954), .B(n955), .Z(n884) );
  NANDN U999 ( .A(n956), .B(n957), .Z(n955) );
  OR U1000 ( .A(n958), .B(n959), .Z(n957) );
  NAND U1001 ( .A(n959), .B(n958), .Z(n954) );
  ANDN U1002 ( .B(B[64]), .A(n57), .Z(n886) );
  XNOR U1003 ( .A(n894), .B(n960), .Z(n887) );
  XNOR U1004 ( .A(n893), .B(n891), .Z(n960) );
  AND U1005 ( .A(n961), .B(n962), .Z(n891) );
  NANDN U1006 ( .A(n963), .B(n964), .Z(n962) );
  NANDN U1007 ( .A(n965), .B(n966), .Z(n964) );
  NANDN U1008 ( .A(n966), .B(n965), .Z(n961) );
  ANDN U1009 ( .B(B[65]), .A(n58), .Z(n893) );
  XNOR U1010 ( .A(n901), .B(n967), .Z(n894) );
  XNOR U1011 ( .A(n900), .B(n898), .Z(n967) );
  AND U1012 ( .A(n968), .B(n969), .Z(n898) );
  NANDN U1013 ( .A(n970), .B(n971), .Z(n969) );
  OR U1014 ( .A(n972), .B(n973), .Z(n971) );
  NAND U1015 ( .A(n973), .B(n972), .Z(n968) );
  ANDN U1016 ( .B(B[66]), .A(n59), .Z(n900) );
  XNOR U1017 ( .A(n908), .B(n974), .Z(n901) );
  XNOR U1018 ( .A(n907), .B(n905), .Z(n974) );
  AND U1019 ( .A(n975), .B(n976), .Z(n905) );
  NANDN U1020 ( .A(n977), .B(n978), .Z(n976) );
  NANDN U1021 ( .A(n979), .B(n980), .Z(n978) );
  NANDN U1022 ( .A(n980), .B(n979), .Z(n975) );
  ANDN U1023 ( .B(B[67]), .A(n60), .Z(n907) );
  XNOR U1024 ( .A(n915), .B(n981), .Z(n908) );
  XNOR U1025 ( .A(n914), .B(n912), .Z(n981) );
  AND U1026 ( .A(n982), .B(n983), .Z(n912) );
  NANDN U1027 ( .A(n984), .B(n985), .Z(n983) );
  OR U1028 ( .A(n986), .B(n987), .Z(n985) );
  NAND U1029 ( .A(n987), .B(n986), .Z(n982) );
  ANDN U1030 ( .B(B[68]), .A(n61), .Z(n914) );
  XOR U1031 ( .A(n919), .B(n988), .Z(n915) );
  XNOR U1032 ( .A(n921), .B(n922), .Z(n988) );
  AND U1033 ( .A(n989), .B(n990), .Z(n922) );
  NAND U1034 ( .A(n991), .B(n992), .Z(n990) );
  NANDN U1035 ( .A(n993), .B(n994), .Z(n991) );
  ANDN U1036 ( .B(B[69]), .A(n62), .Z(n921) );
  XNOR U1037 ( .A(n995), .B(n996), .Z(n919) );
  XNOR U1038 ( .A(n997), .B(n20), .Z(n996) );
  NAND U1039 ( .A(n998), .B(n999), .Z(n103) );
  NANDN U1040 ( .A(n1000), .B(n1001), .Z(n999) );
  OR U1041 ( .A(n1002), .B(n1003), .Z(n1001) );
  NAND U1042 ( .A(n1003), .B(n1002), .Z(n998) );
  XNOR U1043 ( .A(n1004), .B(n1005), .Z(\A1[8] ) );
  XNOR U1044 ( .A(n1006), .B(n1007), .Z(n1005) );
  XOR U1045 ( .A(n105), .B(n104), .Z(\A1[89] ) );
  XOR U1046 ( .A(n1003), .B(n1008), .Z(n104) );
  XNOR U1047 ( .A(n1002), .B(n1000), .Z(n1008) );
  AND U1048 ( .A(n1009), .B(n1010), .Z(n1000) );
  NANDN U1049 ( .A(n1011), .B(n1012), .Z(n1010) );
  NANDN U1050 ( .A(n1013), .B(n1014), .Z(n1012) );
  NANDN U1051 ( .A(n1014), .B(n1013), .Z(n1009) );
  ANDN U1052 ( .B(B[60]), .A(n54), .Z(n1002) );
  XNOR U1053 ( .A(n938), .B(n1015), .Z(n1003) );
  XNOR U1054 ( .A(n937), .B(n935), .Z(n1015) );
  AND U1055 ( .A(n1016), .B(n1017), .Z(n935) );
  NANDN U1056 ( .A(n1018), .B(n1019), .Z(n1017) );
  OR U1057 ( .A(n1020), .B(n1021), .Z(n1019) );
  NAND U1058 ( .A(n1021), .B(n1020), .Z(n1016) );
  ANDN U1059 ( .B(B[61]), .A(n55), .Z(n937) );
  XNOR U1060 ( .A(n945), .B(n1022), .Z(n938) );
  XNOR U1061 ( .A(n944), .B(n942), .Z(n1022) );
  AND U1062 ( .A(n1023), .B(n1024), .Z(n942) );
  NANDN U1063 ( .A(n1025), .B(n1026), .Z(n1024) );
  NANDN U1064 ( .A(n1027), .B(n1028), .Z(n1026) );
  NANDN U1065 ( .A(n1028), .B(n1027), .Z(n1023) );
  ANDN U1066 ( .B(B[62]), .A(n56), .Z(n944) );
  XNOR U1067 ( .A(n952), .B(n1029), .Z(n945) );
  XNOR U1068 ( .A(n951), .B(n949), .Z(n1029) );
  AND U1069 ( .A(n1030), .B(n1031), .Z(n949) );
  NANDN U1070 ( .A(n1032), .B(n1033), .Z(n1031) );
  OR U1071 ( .A(n1034), .B(n1035), .Z(n1033) );
  NAND U1072 ( .A(n1035), .B(n1034), .Z(n1030) );
  ANDN U1073 ( .B(B[63]), .A(n57), .Z(n951) );
  XNOR U1074 ( .A(n959), .B(n1036), .Z(n952) );
  XNOR U1075 ( .A(n958), .B(n956), .Z(n1036) );
  AND U1076 ( .A(n1037), .B(n1038), .Z(n956) );
  NANDN U1077 ( .A(n1039), .B(n1040), .Z(n1038) );
  NANDN U1078 ( .A(n1041), .B(n1042), .Z(n1040) );
  NANDN U1079 ( .A(n1042), .B(n1041), .Z(n1037) );
  ANDN U1080 ( .B(B[64]), .A(n58), .Z(n958) );
  XNOR U1081 ( .A(n966), .B(n1043), .Z(n959) );
  XNOR U1082 ( .A(n965), .B(n963), .Z(n1043) );
  AND U1083 ( .A(n1044), .B(n1045), .Z(n963) );
  NANDN U1084 ( .A(n1046), .B(n1047), .Z(n1045) );
  OR U1085 ( .A(n1048), .B(n1049), .Z(n1047) );
  NAND U1086 ( .A(n1049), .B(n1048), .Z(n1044) );
  ANDN U1087 ( .B(B[65]), .A(n59), .Z(n965) );
  XNOR U1088 ( .A(n973), .B(n1050), .Z(n966) );
  XNOR U1089 ( .A(n972), .B(n970), .Z(n1050) );
  AND U1090 ( .A(n1051), .B(n1052), .Z(n970) );
  NANDN U1091 ( .A(n1053), .B(n1054), .Z(n1052) );
  NANDN U1092 ( .A(n1055), .B(n1056), .Z(n1054) );
  NANDN U1093 ( .A(n1056), .B(n1055), .Z(n1051) );
  ANDN U1094 ( .B(B[66]), .A(n60), .Z(n972) );
  XNOR U1095 ( .A(n980), .B(n1057), .Z(n973) );
  XNOR U1096 ( .A(n979), .B(n977), .Z(n1057) );
  AND U1097 ( .A(n1058), .B(n1059), .Z(n977) );
  NANDN U1098 ( .A(n1060), .B(n1061), .Z(n1059) );
  OR U1099 ( .A(n1062), .B(n1063), .Z(n1061) );
  NAND U1100 ( .A(n1063), .B(n1062), .Z(n1058) );
  ANDN U1101 ( .B(B[67]), .A(n61), .Z(n979) );
  XNOR U1102 ( .A(n987), .B(n1064), .Z(n980) );
  XNOR U1103 ( .A(n986), .B(n984), .Z(n1064) );
  AND U1104 ( .A(n1065), .B(n1066), .Z(n984) );
  NANDN U1105 ( .A(n1067), .B(n1068), .Z(n1066) );
  NANDN U1106 ( .A(n1069), .B(n1070), .Z(n1068) );
  NANDN U1107 ( .A(n1070), .B(n1069), .Z(n1065) );
  ANDN U1108 ( .B(B[68]), .A(n62), .Z(n986) );
  XOR U1109 ( .A(n992), .B(n1071), .Z(n987) );
  XNOR U1110 ( .A(n993), .B(n994), .Z(n1071) );
  AND U1111 ( .A(n1072), .B(n1073), .Z(n994) );
  NANDN U1112 ( .A(n1074), .B(n1075), .Z(n1073) );
  NANDN U1113 ( .A(n1076), .B(n1077), .Z(n1075) );
  ANDN U1114 ( .B(B[69]), .A(n63), .Z(n993) );
  XOR U1115 ( .A(n1078), .B(n1079), .Z(n992) );
  XNOR U1116 ( .A(n1080), .B(n22), .Z(n1079) );
  NAND U1117 ( .A(n1081), .B(n1082), .Z(n105) );
  NANDN U1118 ( .A(n1083), .B(n1084), .Z(n1082) );
  OR U1119 ( .A(n1085), .B(n1086), .Z(n1084) );
  NAND U1120 ( .A(n1086), .B(n1085), .Z(n1081) );
  XOR U1121 ( .A(n107), .B(n106), .Z(\A1[88] ) );
  XOR U1122 ( .A(n1086), .B(n1087), .Z(n106) );
  XNOR U1123 ( .A(n1085), .B(n1083), .Z(n1087) );
  AND U1124 ( .A(n1088), .B(n1089), .Z(n1083) );
  NANDN U1125 ( .A(n1090), .B(n1091), .Z(n1089) );
  NANDN U1126 ( .A(n1092), .B(n1093), .Z(n1091) );
  NANDN U1127 ( .A(n1093), .B(n1092), .Z(n1088) );
  ANDN U1128 ( .B(B[59]), .A(n54), .Z(n1085) );
  XNOR U1129 ( .A(n1014), .B(n1094), .Z(n1086) );
  XNOR U1130 ( .A(n1013), .B(n1011), .Z(n1094) );
  AND U1131 ( .A(n1095), .B(n1096), .Z(n1011) );
  NANDN U1132 ( .A(n1097), .B(n1098), .Z(n1096) );
  OR U1133 ( .A(n1099), .B(n1100), .Z(n1098) );
  NAND U1134 ( .A(n1100), .B(n1099), .Z(n1095) );
  ANDN U1135 ( .B(B[60]), .A(n55), .Z(n1013) );
  XNOR U1136 ( .A(n1021), .B(n1101), .Z(n1014) );
  XNOR U1137 ( .A(n1020), .B(n1018), .Z(n1101) );
  AND U1138 ( .A(n1102), .B(n1103), .Z(n1018) );
  NANDN U1139 ( .A(n1104), .B(n1105), .Z(n1103) );
  NANDN U1140 ( .A(n1106), .B(n1107), .Z(n1105) );
  NANDN U1141 ( .A(n1107), .B(n1106), .Z(n1102) );
  ANDN U1142 ( .B(B[61]), .A(n56), .Z(n1020) );
  XNOR U1143 ( .A(n1028), .B(n1108), .Z(n1021) );
  XNOR U1144 ( .A(n1027), .B(n1025), .Z(n1108) );
  AND U1145 ( .A(n1109), .B(n1110), .Z(n1025) );
  NANDN U1146 ( .A(n1111), .B(n1112), .Z(n1110) );
  OR U1147 ( .A(n1113), .B(n1114), .Z(n1112) );
  NAND U1148 ( .A(n1114), .B(n1113), .Z(n1109) );
  ANDN U1149 ( .B(B[62]), .A(n57), .Z(n1027) );
  XNOR U1150 ( .A(n1035), .B(n1115), .Z(n1028) );
  XNOR U1151 ( .A(n1034), .B(n1032), .Z(n1115) );
  AND U1152 ( .A(n1116), .B(n1117), .Z(n1032) );
  NANDN U1153 ( .A(n1118), .B(n1119), .Z(n1117) );
  NANDN U1154 ( .A(n1120), .B(n1121), .Z(n1119) );
  NANDN U1155 ( .A(n1121), .B(n1120), .Z(n1116) );
  ANDN U1156 ( .B(B[63]), .A(n58), .Z(n1034) );
  XNOR U1157 ( .A(n1042), .B(n1122), .Z(n1035) );
  XNOR U1158 ( .A(n1041), .B(n1039), .Z(n1122) );
  AND U1159 ( .A(n1123), .B(n1124), .Z(n1039) );
  NANDN U1160 ( .A(n1125), .B(n1126), .Z(n1124) );
  OR U1161 ( .A(n1127), .B(n1128), .Z(n1126) );
  NAND U1162 ( .A(n1128), .B(n1127), .Z(n1123) );
  ANDN U1163 ( .B(B[64]), .A(n59), .Z(n1041) );
  XNOR U1164 ( .A(n1049), .B(n1129), .Z(n1042) );
  XNOR U1165 ( .A(n1048), .B(n1046), .Z(n1129) );
  AND U1166 ( .A(n1130), .B(n1131), .Z(n1046) );
  NANDN U1167 ( .A(n1132), .B(n1133), .Z(n1131) );
  NANDN U1168 ( .A(n1134), .B(n1135), .Z(n1133) );
  NANDN U1169 ( .A(n1135), .B(n1134), .Z(n1130) );
  ANDN U1170 ( .B(B[65]), .A(n60), .Z(n1048) );
  XNOR U1171 ( .A(n1056), .B(n1136), .Z(n1049) );
  XNOR U1172 ( .A(n1055), .B(n1053), .Z(n1136) );
  AND U1173 ( .A(n1137), .B(n1138), .Z(n1053) );
  NANDN U1174 ( .A(n1139), .B(n1140), .Z(n1138) );
  OR U1175 ( .A(n1141), .B(n1142), .Z(n1140) );
  NAND U1176 ( .A(n1142), .B(n1141), .Z(n1137) );
  ANDN U1177 ( .B(B[66]), .A(n61), .Z(n1055) );
  XNOR U1178 ( .A(n1063), .B(n1143), .Z(n1056) );
  XNOR U1179 ( .A(n1062), .B(n1060), .Z(n1143) );
  AND U1180 ( .A(n1144), .B(n1145), .Z(n1060) );
  NANDN U1181 ( .A(n1146), .B(n1147), .Z(n1145) );
  NANDN U1182 ( .A(n1148), .B(n1149), .Z(n1147) );
  NANDN U1183 ( .A(n1149), .B(n1148), .Z(n1144) );
  ANDN U1184 ( .B(B[67]), .A(n62), .Z(n1062) );
  XNOR U1185 ( .A(n1070), .B(n1150), .Z(n1063) );
  XNOR U1186 ( .A(n1069), .B(n1067), .Z(n1150) );
  AND U1187 ( .A(n1151), .B(n1152), .Z(n1067) );
  NANDN U1188 ( .A(n1153), .B(n1154), .Z(n1152) );
  OR U1189 ( .A(n1155), .B(n1156), .Z(n1154) );
  NAND U1190 ( .A(n1156), .B(n1155), .Z(n1151) );
  ANDN U1191 ( .B(B[68]), .A(n63), .Z(n1069) );
  XOR U1192 ( .A(n1074), .B(n1157), .Z(n1070) );
  XNOR U1193 ( .A(n1076), .B(n1077), .Z(n1157) );
  AND U1194 ( .A(n1158), .B(n1159), .Z(n1077) );
  NAND U1195 ( .A(n1160), .B(n1161), .Z(n1159) );
  NANDN U1196 ( .A(n1162), .B(n1163), .Z(n1160) );
  ANDN U1197 ( .B(B[69]), .A(n64), .Z(n1076) );
  XNOR U1198 ( .A(n1164), .B(n1165), .Z(n1074) );
  XNOR U1199 ( .A(n1166), .B(n24), .Z(n1165) );
  NAND U1200 ( .A(n1167), .B(n1168), .Z(n107) );
  NANDN U1201 ( .A(n1169), .B(n1170), .Z(n1168) );
  OR U1202 ( .A(n1171), .B(n1172), .Z(n1170) );
  NAND U1203 ( .A(n1172), .B(n1171), .Z(n1167) );
  XOR U1204 ( .A(n109), .B(n108), .Z(\A1[87] ) );
  XOR U1205 ( .A(n1172), .B(n1173), .Z(n108) );
  XNOR U1206 ( .A(n1171), .B(n1169), .Z(n1173) );
  AND U1207 ( .A(n1174), .B(n1175), .Z(n1169) );
  NANDN U1208 ( .A(n1176), .B(n1177), .Z(n1175) );
  NANDN U1209 ( .A(n1178), .B(n1179), .Z(n1177) );
  NANDN U1210 ( .A(n1179), .B(n1178), .Z(n1174) );
  ANDN U1211 ( .B(B[58]), .A(n54), .Z(n1171) );
  XNOR U1212 ( .A(n1093), .B(n1180), .Z(n1172) );
  XNOR U1213 ( .A(n1092), .B(n1090), .Z(n1180) );
  AND U1214 ( .A(n1181), .B(n1182), .Z(n1090) );
  NANDN U1215 ( .A(n1183), .B(n1184), .Z(n1182) );
  OR U1216 ( .A(n1185), .B(n1186), .Z(n1184) );
  NAND U1217 ( .A(n1186), .B(n1185), .Z(n1181) );
  ANDN U1218 ( .B(B[59]), .A(n55), .Z(n1092) );
  XNOR U1219 ( .A(n1100), .B(n1187), .Z(n1093) );
  XNOR U1220 ( .A(n1099), .B(n1097), .Z(n1187) );
  AND U1221 ( .A(n1188), .B(n1189), .Z(n1097) );
  NANDN U1222 ( .A(n1190), .B(n1191), .Z(n1189) );
  NANDN U1223 ( .A(n1192), .B(n1193), .Z(n1191) );
  NANDN U1224 ( .A(n1193), .B(n1192), .Z(n1188) );
  ANDN U1225 ( .B(B[60]), .A(n56), .Z(n1099) );
  XNOR U1226 ( .A(n1107), .B(n1194), .Z(n1100) );
  XNOR U1227 ( .A(n1106), .B(n1104), .Z(n1194) );
  AND U1228 ( .A(n1195), .B(n1196), .Z(n1104) );
  NANDN U1229 ( .A(n1197), .B(n1198), .Z(n1196) );
  OR U1230 ( .A(n1199), .B(n1200), .Z(n1198) );
  NAND U1231 ( .A(n1200), .B(n1199), .Z(n1195) );
  ANDN U1232 ( .B(B[61]), .A(n57), .Z(n1106) );
  XNOR U1233 ( .A(n1114), .B(n1201), .Z(n1107) );
  XNOR U1234 ( .A(n1113), .B(n1111), .Z(n1201) );
  AND U1235 ( .A(n1202), .B(n1203), .Z(n1111) );
  NANDN U1236 ( .A(n1204), .B(n1205), .Z(n1203) );
  NANDN U1237 ( .A(n1206), .B(n1207), .Z(n1205) );
  NANDN U1238 ( .A(n1207), .B(n1206), .Z(n1202) );
  ANDN U1239 ( .B(B[62]), .A(n58), .Z(n1113) );
  XNOR U1240 ( .A(n1121), .B(n1208), .Z(n1114) );
  XNOR U1241 ( .A(n1120), .B(n1118), .Z(n1208) );
  AND U1242 ( .A(n1209), .B(n1210), .Z(n1118) );
  NANDN U1243 ( .A(n1211), .B(n1212), .Z(n1210) );
  OR U1244 ( .A(n1213), .B(n1214), .Z(n1212) );
  NAND U1245 ( .A(n1214), .B(n1213), .Z(n1209) );
  ANDN U1246 ( .B(B[63]), .A(n59), .Z(n1120) );
  XNOR U1247 ( .A(n1128), .B(n1215), .Z(n1121) );
  XNOR U1248 ( .A(n1127), .B(n1125), .Z(n1215) );
  AND U1249 ( .A(n1216), .B(n1217), .Z(n1125) );
  NANDN U1250 ( .A(n1218), .B(n1219), .Z(n1217) );
  NANDN U1251 ( .A(n1220), .B(n1221), .Z(n1219) );
  NANDN U1252 ( .A(n1221), .B(n1220), .Z(n1216) );
  ANDN U1253 ( .B(B[64]), .A(n60), .Z(n1127) );
  XNOR U1254 ( .A(n1135), .B(n1222), .Z(n1128) );
  XNOR U1255 ( .A(n1134), .B(n1132), .Z(n1222) );
  AND U1256 ( .A(n1223), .B(n1224), .Z(n1132) );
  NANDN U1257 ( .A(n1225), .B(n1226), .Z(n1224) );
  OR U1258 ( .A(n1227), .B(n1228), .Z(n1226) );
  NAND U1259 ( .A(n1228), .B(n1227), .Z(n1223) );
  ANDN U1260 ( .B(B[65]), .A(n61), .Z(n1134) );
  XNOR U1261 ( .A(n1142), .B(n1229), .Z(n1135) );
  XNOR U1262 ( .A(n1141), .B(n1139), .Z(n1229) );
  AND U1263 ( .A(n1230), .B(n1231), .Z(n1139) );
  NANDN U1264 ( .A(n1232), .B(n1233), .Z(n1231) );
  NANDN U1265 ( .A(n1234), .B(n1235), .Z(n1233) );
  NANDN U1266 ( .A(n1235), .B(n1234), .Z(n1230) );
  ANDN U1267 ( .B(B[66]), .A(n62), .Z(n1141) );
  XNOR U1268 ( .A(n1149), .B(n1236), .Z(n1142) );
  XNOR U1269 ( .A(n1148), .B(n1146), .Z(n1236) );
  AND U1270 ( .A(n1237), .B(n1238), .Z(n1146) );
  NANDN U1271 ( .A(n1239), .B(n1240), .Z(n1238) );
  OR U1272 ( .A(n1241), .B(n1242), .Z(n1240) );
  NAND U1273 ( .A(n1242), .B(n1241), .Z(n1237) );
  ANDN U1274 ( .B(B[67]), .A(n63), .Z(n1148) );
  XNOR U1275 ( .A(n1156), .B(n1243), .Z(n1149) );
  XNOR U1276 ( .A(n1155), .B(n1153), .Z(n1243) );
  AND U1277 ( .A(n1244), .B(n1245), .Z(n1153) );
  NANDN U1278 ( .A(n1246), .B(n1247), .Z(n1245) );
  NANDN U1279 ( .A(n1248), .B(n1249), .Z(n1247) );
  NANDN U1280 ( .A(n1249), .B(n1248), .Z(n1244) );
  ANDN U1281 ( .B(B[68]), .A(n64), .Z(n1155) );
  XOR U1282 ( .A(n1161), .B(n1250), .Z(n1156) );
  XNOR U1283 ( .A(n1162), .B(n1163), .Z(n1250) );
  AND U1284 ( .A(n1251), .B(n1252), .Z(n1163) );
  NANDN U1285 ( .A(n1253), .B(n1254), .Z(n1252) );
  NANDN U1286 ( .A(n1255), .B(n1256), .Z(n1254) );
  ANDN U1287 ( .B(B[69]), .A(n65), .Z(n1162) );
  XOR U1288 ( .A(n1257), .B(n1258), .Z(n1161) );
  XNOR U1289 ( .A(n1259), .B(n26), .Z(n1258) );
  NAND U1290 ( .A(n1260), .B(n1261), .Z(n109) );
  NANDN U1291 ( .A(n1262), .B(n1263), .Z(n1261) );
  OR U1292 ( .A(n1264), .B(n1265), .Z(n1263) );
  NAND U1293 ( .A(n1265), .B(n1264), .Z(n1260) );
  XOR U1294 ( .A(n111), .B(n110), .Z(\A1[86] ) );
  XOR U1295 ( .A(n1265), .B(n1266), .Z(n110) );
  XNOR U1296 ( .A(n1264), .B(n1262), .Z(n1266) );
  AND U1297 ( .A(n1267), .B(n1268), .Z(n1262) );
  NANDN U1298 ( .A(n1269), .B(n1270), .Z(n1268) );
  NANDN U1299 ( .A(n1271), .B(n1272), .Z(n1270) );
  NANDN U1300 ( .A(n1272), .B(n1271), .Z(n1267) );
  ANDN U1301 ( .B(B[57]), .A(n54), .Z(n1264) );
  XNOR U1302 ( .A(n1179), .B(n1273), .Z(n1265) );
  XNOR U1303 ( .A(n1178), .B(n1176), .Z(n1273) );
  AND U1304 ( .A(n1274), .B(n1275), .Z(n1176) );
  NANDN U1305 ( .A(n1276), .B(n1277), .Z(n1275) );
  OR U1306 ( .A(n1278), .B(n1279), .Z(n1277) );
  NAND U1307 ( .A(n1279), .B(n1278), .Z(n1274) );
  ANDN U1308 ( .B(B[58]), .A(n55), .Z(n1178) );
  XNOR U1309 ( .A(n1186), .B(n1280), .Z(n1179) );
  XNOR U1310 ( .A(n1185), .B(n1183), .Z(n1280) );
  AND U1311 ( .A(n1281), .B(n1282), .Z(n1183) );
  NANDN U1312 ( .A(n1283), .B(n1284), .Z(n1282) );
  NANDN U1313 ( .A(n1285), .B(n1286), .Z(n1284) );
  NANDN U1314 ( .A(n1286), .B(n1285), .Z(n1281) );
  ANDN U1315 ( .B(B[59]), .A(n56), .Z(n1185) );
  XNOR U1316 ( .A(n1193), .B(n1287), .Z(n1186) );
  XNOR U1317 ( .A(n1192), .B(n1190), .Z(n1287) );
  AND U1318 ( .A(n1288), .B(n1289), .Z(n1190) );
  NANDN U1319 ( .A(n1290), .B(n1291), .Z(n1289) );
  OR U1320 ( .A(n1292), .B(n1293), .Z(n1291) );
  NAND U1321 ( .A(n1293), .B(n1292), .Z(n1288) );
  ANDN U1322 ( .B(B[60]), .A(n57), .Z(n1192) );
  XNOR U1323 ( .A(n1200), .B(n1294), .Z(n1193) );
  XNOR U1324 ( .A(n1199), .B(n1197), .Z(n1294) );
  AND U1325 ( .A(n1295), .B(n1296), .Z(n1197) );
  NANDN U1326 ( .A(n1297), .B(n1298), .Z(n1296) );
  NANDN U1327 ( .A(n1299), .B(n1300), .Z(n1298) );
  NANDN U1328 ( .A(n1300), .B(n1299), .Z(n1295) );
  ANDN U1329 ( .B(B[61]), .A(n58), .Z(n1199) );
  XNOR U1330 ( .A(n1207), .B(n1301), .Z(n1200) );
  XNOR U1331 ( .A(n1206), .B(n1204), .Z(n1301) );
  AND U1332 ( .A(n1302), .B(n1303), .Z(n1204) );
  NANDN U1333 ( .A(n1304), .B(n1305), .Z(n1303) );
  OR U1334 ( .A(n1306), .B(n1307), .Z(n1305) );
  NAND U1335 ( .A(n1307), .B(n1306), .Z(n1302) );
  ANDN U1336 ( .B(B[62]), .A(n59), .Z(n1206) );
  XNOR U1337 ( .A(n1214), .B(n1308), .Z(n1207) );
  XNOR U1338 ( .A(n1213), .B(n1211), .Z(n1308) );
  AND U1339 ( .A(n1309), .B(n1310), .Z(n1211) );
  NANDN U1340 ( .A(n1311), .B(n1312), .Z(n1310) );
  NANDN U1341 ( .A(n1313), .B(n1314), .Z(n1312) );
  NANDN U1342 ( .A(n1314), .B(n1313), .Z(n1309) );
  ANDN U1343 ( .B(B[63]), .A(n60), .Z(n1213) );
  XNOR U1344 ( .A(n1221), .B(n1315), .Z(n1214) );
  XNOR U1345 ( .A(n1220), .B(n1218), .Z(n1315) );
  AND U1346 ( .A(n1316), .B(n1317), .Z(n1218) );
  NANDN U1347 ( .A(n1318), .B(n1319), .Z(n1317) );
  OR U1348 ( .A(n1320), .B(n1321), .Z(n1319) );
  NAND U1349 ( .A(n1321), .B(n1320), .Z(n1316) );
  ANDN U1350 ( .B(B[64]), .A(n61), .Z(n1220) );
  XNOR U1351 ( .A(n1228), .B(n1322), .Z(n1221) );
  XNOR U1352 ( .A(n1227), .B(n1225), .Z(n1322) );
  AND U1353 ( .A(n1323), .B(n1324), .Z(n1225) );
  NANDN U1354 ( .A(n1325), .B(n1326), .Z(n1324) );
  NANDN U1355 ( .A(n1327), .B(n1328), .Z(n1326) );
  NANDN U1356 ( .A(n1328), .B(n1327), .Z(n1323) );
  ANDN U1357 ( .B(B[65]), .A(n62), .Z(n1227) );
  XNOR U1358 ( .A(n1235), .B(n1329), .Z(n1228) );
  XNOR U1359 ( .A(n1234), .B(n1232), .Z(n1329) );
  AND U1360 ( .A(n1330), .B(n1331), .Z(n1232) );
  NANDN U1361 ( .A(n1332), .B(n1333), .Z(n1331) );
  OR U1362 ( .A(n1334), .B(n1335), .Z(n1333) );
  NAND U1363 ( .A(n1335), .B(n1334), .Z(n1330) );
  ANDN U1364 ( .B(B[66]), .A(n63), .Z(n1234) );
  XNOR U1365 ( .A(n1242), .B(n1336), .Z(n1235) );
  XNOR U1366 ( .A(n1241), .B(n1239), .Z(n1336) );
  AND U1367 ( .A(n1337), .B(n1338), .Z(n1239) );
  NANDN U1368 ( .A(n1339), .B(n1340), .Z(n1338) );
  NANDN U1369 ( .A(n1341), .B(n1342), .Z(n1340) );
  NANDN U1370 ( .A(n1342), .B(n1341), .Z(n1337) );
  ANDN U1371 ( .B(B[67]), .A(n64), .Z(n1241) );
  XNOR U1372 ( .A(n1249), .B(n1343), .Z(n1242) );
  XNOR U1373 ( .A(n1248), .B(n1246), .Z(n1343) );
  AND U1374 ( .A(n1344), .B(n1345), .Z(n1246) );
  NANDN U1375 ( .A(n1346), .B(n1347), .Z(n1345) );
  OR U1376 ( .A(n1348), .B(n1349), .Z(n1347) );
  NAND U1377 ( .A(n1349), .B(n1348), .Z(n1344) );
  ANDN U1378 ( .B(B[68]), .A(n65), .Z(n1248) );
  XOR U1379 ( .A(n1253), .B(n1350), .Z(n1249) );
  XNOR U1380 ( .A(n1255), .B(n1256), .Z(n1350) );
  AND U1381 ( .A(n1351), .B(n1352), .Z(n1256) );
  NAND U1382 ( .A(n1353), .B(n1354), .Z(n1352) );
  NANDN U1383 ( .A(n1355), .B(n1356), .Z(n1353) );
  ANDN U1384 ( .B(B[69]), .A(n66), .Z(n1255) );
  XNOR U1385 ( .A(n1357), .B(n1358), .Z(n1253) );
  XNOR U1386 ( .A(n1359), .B(n28), .Z(n1358) );
  NAND U1387 ( .A(n1360), .B(n1361), .Z(n111) );
  NANDN U1388 ( .A(n1362), .B(n1363), .Z(n1361) );
  OR U1389 ( .A(n1364), .B(n1365), .Z(n1363) );
  NAND U1390 ( .A(n1365), .B(n1364), .Z(n1360) );
  XOR U1391 ( .A(n113), .B(n112), .Z(\A1[85] ) );
  XOR U1392 ( .A(n1365), .B(n1366), .Z(n112) );
  XNOR U1393 ( .A(n1364), .B(n1362), .Z(n1366) );
  AND U1394 ( .A(n1367), .B(n1368), .Z(n1362) );
  NANDN U1395 ( .A(n1369), .B(n1370), .Z(n1368) );
  NANDN U1396 ( .A(n1371), .B(n1372), .Z(n1370) );
  NANDN U1397 ( .A(n1372), .B(n1371), .Z(n1367) );
  ANDN U1398 ( .B(B[56]), .A(n54), .Z(n1364) );
  XNOR U1399 ( .A(n1272), .B(n1373), .Z(n1365) );
  XNOR U1400 ( .A(n1271), .B(n1269), .Z(n1373) );
  AND U1401 ( .A(n1374), .B(n1375), .Z(n1269) );
  NANDN U1402 ( .A(n1376), .B(n1377), .Z(n1375) );
  OR U1403 ( .A(n1378), .B(n1379), .Z(n1377) );
  NAND U1404 ( .A(n1379), .B(n1378), .Z(n1374) );
  ANDN U1405 ( .B(B[57]), .A(n55), .Z(n1271) );
  XNOR U1406 ( .A(n1279), .B(n1380), .Z(n1272) );
  XNOR U1407 ( .A(n1278), .B(n1276), .Z(n1380) );
  AND U1408 ( .A(n1381), .B(n1382), .Z(n1276) );
  NANDN U1409 ( .A(n1383), .B(n1384), .Z(n1382) );
  NANDN U1410 ( .A(n1385), .B(n1386), .Z(n1384) );
  NANDN U1411 ( .A(n1386), .B(n1385), .Z(n1381) );
  ANDN U1412 ( .B(B[58]), .A(n56), .Z(n1278) );
  XNOR U1413 ( .A(n1286), .B(n1387), .Z(n1279) );
  XNOR U1414 ( .A(n1285), .B(n1283), .Z(n1387) );
  AND U1415 ( .A(n1388), .B(n1389), .Z(n1283) );
  NANDN U1416 ( .A(n1390), .B(n1391), .Z(n1389) );
  OR U1417 ( .A(n1392), .B(n1393), .Z(n1391) );
  NAND U1418 ( .A(n1393), .B(n1392), .Z(n1388) );
  ANDN U1419 ( .B(B[59]), .A(n57), .Z(n1285) );
  XNOR U1420 ( .A(n1293), .B(n1394), .Z(n1286) );
  XNOR U1421 ( .A(n1292), .B(n1290), .Z(n1394) );
  AND U1422 ( .A(n1395), .B(n1396), .Z(n1290) );
  NANDN U1423 ( .A(n1397), .B(n1398), .Z(n1396) );
  NANDN U1424 ( .A(n1399), .B(n1400), .Z(n1398) );
  NANDN U1425 ( .A(n1400), .B(n1399), .Z(n1395) );
  ANDN U1426 ( .B(B[60]), .A(n58), .Z(n1292) );
  XNOR U1427 ( .A(n1300), .B(n1401), .Z(n1293) );
  XNOR U1428 ( .A(n1299), .B(n1297), .Z(n1401) );
  AND U1429 ( .A(n1402), .B(n1403), .Z(n1297) );
  NANDN U1430 ( .A(n1404), .B(n1405), .Z(n1403) );
  OR U1431 ( .A(n1406), .B(n1407), .Z(n1405) );
  NAND U1432 ( .A(n1407), .B(n1406), .Z(n1402) );
  ANDN U1433 ( .B(B[61]), .A(n59), .Z(n1299) );
  XNOR U1434 ( .A(n1307), .B(n1408), .Z(n1300) );
  XNOR U1435 ( .A(n1306), .B(n1304), .Z(n1408) );
  AND U1436 ( .A(n1409), .B(n1410), .Z(n1304) );
  NANDN U1437 ( .A(n1411), .B(n1412), .Z(n1410) );
  NANDN U1438 ( .A(n1413), .B(n1414), .Z(n1412) );
  NANDN U1439 ( .A(n1414), .B(n1413), .Z(n1409) );
  ANDN U1440 ( .B(B[62]), .A(n60), .Z(n1306) );
  XNOR U1441 ( .A(n1314), .B(n1415), .Z(n1307) );
  XNOR U1442 ( .A(n1313), .B(n1311), .Z(n1415) );
  AND U1443 ( .A(n1416), .B(n1417), .Z(n1311) );
  NANDN U1444 ( .A(n1418), .B(n1419), .Z(n1417) );
  OR U1445 ( .A(n1420), .B(n1421), .Z(n1419) );
  NAND U1446 ( .A(n1421), .B(n1420), .Z(n1416) );
  ANDN U1447 ( .B(B[63]), .A(n61), .Z(n1313) );
  XNOR U1448 ( .A(n1321), .B(n1422), .Z(n1314) );
  XNOR U1449 ( .A(n1320), .B(n1318), .Z(n1422) );
  AND U1450 ( .A(n1423), .B(n1424), .Z(n1318) );
  NANDN U1451 ( .A(n1425), .B(n1426), .Z(n1424) );
  NANDN U1452 ( .A(n1427), .B(n1428), .Z(n1426) );
  NANDN U1453 ( .A(n1428), .B(n1427), .Z(n1423) );
  ANDN U1454 ( .B(B[64]), .A(n62), .Z(n1320) );
  XNOR U1455 ( .A(n1328), .B(n1429), .Z(n1321) );
  XNOR U1456 ( .A(n1327), .B(n1325), .Z(n1429) );
  AND U1457 ( .A(n1430), .B(n1431), .Z(n1325) );
  NANDN U1458 ( .A(n1432), .B(n1433), .Z(n1431) );
  OR U1459 ( .A(n1434), .B(n1435), .Z(n1433) );
  NAND U1460 ( .A(n1435), .B(n1434), .Z(n1430) );
  ANDN U1461 ( .B(B[65]), .A(n63), .Z(n1327) );
  XNOR U1462 ( .A(n1335), .B(n1436), .Z(n1328) );
  XNOR U1463 ( .A(n1334), .B(n1332), .Z(n1436) );
  AND U1464 ( .A(n1437), .B(n1438), .Z(n1332) );
  NANDN U1465 ( .A(n1439), .B(n1440), .Z(n1438) );
  NANDN U1466 ( .A(n1441), .B(n1442), .Z(n1440) );
  NANDN U1467 ( .A(n1442), .B(n1441), .Z(n1437) );
  ANDN U1468 ( .B(B[66]), .A(n64), .Z(n1334) );
  XNOR U1469 ( .A(n1342), .B(n1443), .Z(n1335) );
  XNOR U1470 ( .A(n1341), .B(n1339), .Z(n1443) );
  AND U1471 ( .A(n1444), .B(n1445), .Z(n1339) );
  NANDN U1472 ( .A(n1446), .B(n1447), .Z(n1445) );
  OR U1473 ( .A(n1448), .B(n1449), .Z(n1447) );
  NAND U1474 ( .A(n1449), .B(n1448), .Z(n1444) );
  ANDN U1475 ( .B(B[67]), .A(n65), .Z(n1341) );
  XNOR U1476 ( .A(n1349), .B(n1450), .Z(n1342) );
  XNOR U1477 ( .A(n1348), .B(n1346), .Z(n1450) );
  AND U1478 ( .A(n1451), .B(n1452), .Z(n1346) );
  NANDN U1479 ( .A(n1453), .B(n1454), .Z(n1452) );
  NANDN U1480 ( .A(n1455), .B(n1456), .Z(n1454) );
  NANDN U1481 ( .A(n1456), .B(n1455), .Z(n1451) );
  ANDN U1482 ( .B(B[68]), .A(n66), .Z(n1348) );
  XOR U1483 ( .A(n1354), .B(n1457), .Z(n1349) );
  XNOR U1484 ( .A(n1355), .B(n1356), .Z(n1457) );
  AND U1485 ( .A(n1458), .B(n1459), .Z(n1356) );
  NANDN U1486 ( .A(n1460), .B(n1461), .Z(n1459) );
  NANDN U1487 ( .A(n1462), .B(n1463), .Z(n1461) );
  ANDN U1488 ( .B(B[69]), .A(n67), .Z(n1355) );
  XOR U1489 ( .A(n1464), .B(n1465), .Z(n1354) );
  XNOR U1490 ( .A(n1466), .B(n30), .Z(n1465) );
  NAND U1491 ( .A(n1467), .B(n1468), .Z(n113) );
  NANDN U1492 ( .A(n1469), .B(n1470), .Z(n1468) );
  OR U1493 ( .A(n1471), .B(n1472), .Z(n1470) );
  NAND U1494 ( .A(n1472), .B(n1471), .Z(n1467) );
  XOR U1495 ( .A(n115), .B(n114), .Z(\A1[84] ) );
  XOR U1496 ( .A(n1472), .B(n1473), .Z(n114) );
  XNOR U1497 ( .A(n1471), .B(n1469), .Z(n1473) );
  AND U1498 ( .A(n1474), .B(n1475), .Z(n1469) );
  NANDN U1499 ( .A(n1476), .B(n1477), .Z(n1475) );
  NANDN U1500 ( .A(n1478), .B(n1479), .Z(n1477) );
  NANDN U1501 ( .A(n1479), .B(n1478), .Z(n1474) );
  ANDN U1502 ( .B(B[55]), .A(n54), .Z(n1471) );
  XNOR U1503 ( .A(n1372), .B(n1480), .Z(n1472) );
  XNOR U1504 ( .A(n1371), .B(n1369), .Z(n1480) );
  AND U1505 ( .A(n1481), .B(n1482), .Z(n1369) );
  NANDN U1506 ( .A(n1483), .B(n1484), .Z(n1482) );
  OR U1507 ( .A(n1485), .B(n1486), .Z(n1484) );
  NAND U1508 ( .A(n1486), .B(n1485), .Z(n1481) );
  ANDN U1509 ( .B(B[56]), .A(n55), .Z(n1371) );
  XNOR U1510 ( .A(n1379), .B(n1487), .Z(n1372) );
  XNOR U1511 ( .A(n1378), .B(n1376), .Z(n1487) );
  AND U1512 ( .A(n1488), .B(n1489), .Z(n1376) );
  NANDN U1513 ( .A(n1490), .B(n1491), .Z(n1489) );
  NANDN U1514 ( .A(n1492), .B(n1493), .Z(n1491) );
  NANDN U1515 ( .A(n1493), .B(n1492), .Z(n1488) );
  ANDN U1516 ( .B(B[57]), .A(n56), .Z(n1378) );
  XNOR U1517 ( .A(n1386), .B(n1494), .Z(n1379) );
  XNOR U1518 ( .A(n1385), .B(n1383), .Z(n1494) );
  AND U1519 ( .A(n1495), .B(n1496), .Z(n1383) );
  NANDN U1520 ( .A(n1497), .B(n1498), .Z(n1496) );
  OR U1521 ( .A(n1499), .B(n1500), .Z(n1498) );
  NAND U1522 ( .A(n1500), .B(n1499), .Z(n1495) );
  ANDN U1523 ( .B(B[58]), .A(n57), .Z(n1385) );
  XNOR U1524 ( .A(n1393), .B(n1501), .Z(n1386) );
  XNOR U1525 ( .A(n1392), .B(n1390), .Z(n1501) );
  AND U1526 ( .A(n1502), .B(n1503), .Z(n1390) );
  NANDN U1527 ( .A(n1504), .B(n1505), .Z(n1503) );
  NANDN U1528 ( .A(n1506), .B(n1507), .Z(n1505) );
  NANDN U1529 ( .A(n1507), .B(n1506), .Z(n1502) );
  ANDN U1530 ( .B(B[59]), .A(n58), .Z(n1392) );
  XNOR U1531 ( .A(n1400), .B(n1508), .Z(n1393) );
  XNOR U1532 ( .A(n1399), .B(n1397), .Z(n1508) );
  AND U1533 ( .A(n1509), .B(n1510), .Z(n1397) );
  NANDN U1534 ( .A(n1511), .B(n1512), .Z(n1510) );
  OR U1535 ( .A(n1513), .B(n1514), .Z(n1512) );
  NAND U1536 ( .A(n1514), .B(n1513), .Z(n1509) );
  ANDN U1537 ( .B(B[60]), .A(n59), .Z(n1399) );
  XNOR U1538 ( .A(n1407), .B(n1515), .Z(n1400) );
  XNOR U1539 ( .A(n1406), .B(n1404), .Z(n1515) );
  AND U1540 ( .A(n1516), .B(n1517), .Z(n1404) );
  NANDN U1541 ( .A(n1518), .B(n1519), .Z(n1517) );
  NANDN U1542 ( .A(n1520), .B(n1521), .Z(n1519) );
  NANDN U1543 ( .A(n1521), .B(n1520), .Z(n1516) );
  ANDN U1544 ( .B(B[61]), .A(n60), .Z(n1406) );
  XNOR U1545 ( .A(n1414), .B(n1522), .Z(n1407) );
  XNOR U1546 ( .A(n1413), .B(n1411), .Z(n1522) );
  AND U1547 ( .A(n1523), .B(n1524), .Z(n1411) );
  NANDN U1548 ( .A(n1525), .B(n1526), .Z(n1524) );
  OR U1549 ( .A(n1527), .B(n1528), .Z(n1526) );
  NAND U1550 ( .A(n1528), .B(n1527), .Z(n1523) );
  ANDN U1551 ( .B(B[62]), .A(n61), .Z(n1413) );
  XNOR U1552 ( .A(n1421), .B(n1529), .Z(n1414) );
  XNOR U1553 ( .A(n1420), .B(n1418), .Z(n1529) );
  AND U1554 ( .A(n1530), .B(n1531), .Z(n1418) );
  NANDN U1555 ( .A(n1532), .B(n1533), .Z(n1531) );
  NANDN U1556 ( .A(n1534), .B(n1535), .Z(n1533) );
  NANDN U1557 ( .A(n1535), .B(n1534), .Z(n1530) );
  ANDN U1558 ( .B(B[63]), .A(n62), .Z(n1420) );
  XNOR U1559 ( .A(n1428), .B(n1536), .Z(n1421) );
  XNOR U1560 ( .A(n1427), .B(n1425), .Z(n1536) );
  AND U1561 ( .A(n1537), .B(n1538), .Z(n1425) );
  NANDN U1562 ( .A(n1539), .B(n1540), .Z(n1538) );
  OR U1563 ( .A(n1541), .B(n1542), .Z(n1540) );
  NAND U1564 ( .A(n1542), .B(n1541), .Z(n1537) );
  ANDN U1565 ( .B(B[64]), .A(n63), .Z(n1427) );
  XNOR U1566 ( .A(n1435), .B(n1543), .Z(n1428) );
  XNOR U1567 ( .A(n1434), .B(n1432), .Z(n1543) );
  AND U1568 ( .A(n1544), .B(n1545), .Z(n1432) );
  NANDN U1569 ( .A(n1546), .B(n1547), .Z(n1545) );
  NANDN U1570 ( .A(n1548), .B(n1549), .Z(n1547) );
  NANDN U1571 ( .A(n1549), .B(n1548), .Z(n1544) );
  ANDN U1572 ( .B(B[65]), .A(n64), .Z(n1434) );
  XNOR U1573 ( .A(n1442), .B(n1550), .Z(n1435) );
  XNOR U1574 ( .A(n1441), .B(n1439), .Z(n1550) );
  AND U1575 ( .A(n1551), .B(n1552), .Z(n1439) );
  NANDN U1576 ( .A(n1553), .B(n1554), .Z(n1552) );
  OR U1577 ( .A(n1555), .B(n1556), .Z(n1554) );
  NAND U1578 ( .A(n1556), .B(n1555), .Z(n1551) );
  ANDN U1579 ( .B(B[66]), .A(n65), .Z(n1441) );
  XNOR U1580 ( .A(n1449), .B(n1557), .Z(n1442) );
  XNOR U1581 ( .A(n1448), .B(n1446), .Z(n1557) );
  AND U1582 ( .A(n1558), .B(n1559), .Z(n1446) );
  NANDN U1583 ( .A(n1560), .B(n1561), .Z(n1559) );
  NANDN U1584 ( .A(n1562), .B(n1563), .Z(n1561) );
  NANDN U1585 ( .A(n1563), .B(n1562), .Z(n1558) );
  ANDN U1586 ( .B(B[67]), .A(n66), .Z(n1448) );
  XNOR U1587 ( .A(n1456), .B(n1564), .Z(n1449) );
  XNOR U1588 ( .A(n1455), .B(n1453), .Z(n1564) );
  AND U1589 ( .A(n1565), .B(n1566), .Z(n1453) );
  NANDN U1590 ( .A(n1567), .B(n1568), .Z(n1566) );
  OR U1591 ( .A(n1569), .B(n1570), .Z(n1568) );
  NAND U1592 ( .A(n1570), .B(n1569), .Z(n1565) );
  ANDN U1593 ( .B(B[68]), .A(n67), .Z(n1455) );
  XOR U1594 ( .A(n1460), .B(n1571), .Z(n1456) );
  XNOR U1595 ( .A(n1462), .B(n1463), .Z(n1571) );
  AND U1596 ( .A(n1572), .B(n1573), .Z(n1463) );
  NAND U1597 ( .A(n1574), .B(n1575), .Z(n1573) );
  NANDN U1598 ( .A(n1576), .B(n1577), .Z(n1574) );
  ANDN U1599 ( .B(B[69]), .A(n68), .Z(n1462) );
  XNOR U1600 ( .A(n1578), .B(n1579), .Z(n1460) );
  XNOR U1601 ( .A(n1580), .B(n32), .Z(n1579) );
  NAND U1602 ( .A(n1581), .B(n1582), .Z(n115) );
  NANDN U1603 ( .A(n1583), .B(n1584), .Z(n1582) );
  OR U1604 ( .A(n1585), .B(n1586), .Z(n1584) );
  NAND U1605 ( .A(n1586), .B(n1585), .Z(n1581) );
  XOR U1606 ( .A(n117), .B(n116), .Z(\A1[83] ) );
  XOR U1607 ( .A(n1586), .B(n1587), .Z(n116) );
  XNOR U1608 ( .A(n1585), .B(n1583), .Z(n1587) );
  AND U1609 ( .A(n1588), .B(n1589), .Z(n1583) );
  NANDN U1610 ( .A(n1590), .B(n1591), .Z(n1589) );
  NANDN U1611 ( .A(n1592), .B(n1593), .Z(n1591) );
  NANDN U1612 ( .A(n1593), .B(n1592), .Z(n1588) );
  ANDN U1613 ( .B(B[54]), .A(n54), .Z(n1585) );
  XNOR U1614 ( .A(n1479), .B(n1594), .Z(n1586) );
  XNOR U1615 ( .A(n1478), .B(n1476), .Z(n1594) );
  AND U1616 ( .A(n1595), .B(n1596), .Z(n1476) );
  NANDN U1617 ( .A(n1597), .B(n1598), .Z(n1596) );
  OR U1618 ( .A(n1599), .B(n1600), .Z(n1598) );
  NAND U1619 ( .A(n1600), .B(n1599), .Z(n1595) );
  ANDN U1620 ( .B(B[55]), .A(n55), .Z(n1478) );
  XNOR U1621 ( .A(n1486), .B(n1601), .Z(n1479) );
  XNOR U1622 ( .A(n1485), .B(n1483), .Z(n1601) );
  AND U1623 ( .A(n1602), .B(n1603), .Z(n1483) );
  NANDN U1624 ( .A(n1604), .B(n1605), .Z(n1603) );
  NANDN U1625 ( .A(n1606), .B(n1607), .Z(n1605) );
  NANDN U1626 ( .A(n1607), .B(n1606), .Z(n1602) );
  ANDN U1627 ( .B(B[56]), .A(n56), .Z(n1485) );
  XNOR U1628 ( .A(n1493), .B(n1608), .Z(n1486) );
  XNOR U1629 ( .A(n1492), .B(n1490), .Z(n1608) );
  AND U1630 ( .A(n1609), .B(n1610), .Z(n1490) );
  NANDN U1631 ( .A(n1611), .B(n1612), .Z(n1610) );
  OR U1632 ( .A(n1613), .B(n1614), .Z(n1612) );
  NAND U1633 ( .A(n1614), .B(n1613), .Z(n1609) );
  ANDN U1634 ( .B(B[57]), .A(n57), .Z(n1492) );
  XNOR U1635 ( .A(n1500), .B(n1615), .Z(n1493) );
  XNOR U1636 ( .A(n1499), .B(n1497), .Z(n1615) );
  AND U1637 ( .A(n1616), .B(n1617), .Z(n1497) );
  NANDN U1638 ( .A(n1618), .B(n1619), .Z(n1617) );
  NANDN U1639 ( .A(n1620), .B(n1621), .Z(n1619) );
  NANDN U1640 ( .A(n1621), .B(n1620), .Z(n1616) );
  ANDN U1641 ( .B(B[58]), .A(n58), .Z(n1499) );
  XNOR U1642 ( .A(n1507), .B(n1622), .Z(n1500) );
  XNOR U1643 ( .A(n1506), .B(n1504), .Z(n1622) );
  AND U1644 ( .A(n1623), .B(n1624), .Z(n1504) );
  NANDN U1645 ( .A(n1625), .B(n1626), .Z(n1624) );
  OR U1646 ( .A(n1627), .B(n1628), .Z(n1626) );
  NAND U1647 ( .A(n1628), .B(n1627), .Z(n1623) );
  ANDN U1648 ( .B(B[59]), .A(n59), .Z(n1506) );
  XNOR U1649 ( .A(n1514), .B(n1629), .Z(n1507) );
  XNOR U1650 ( .A(n1513), .B(n1511), .Z(n1629) );
  AND U1651 ( .A(n1630), .B(n1631), .Z(n1511) );
  NANDN U1652 ( .A(n1632), .B(n1633), .Z(n1631) );
  NANDN U1653 ( .A(n1634), .B(n1635), .Z(n1633) );
  NANDN U1654 ( .A(n1635), .B(n1634), .Z(n1630) );
  ANDN U1655 ( .B(B[60]), .A(n60), .Z(n1513) );
  XNOR U1656 ( .A(n1521), .B(n1636), .Z(n1514) );
  XNOR U1657 ( .A(n1520), .B(n1518), .Z(n1636) );
  AND U1658 ( .A(n1637), .B(n1638), .Z(n1518) );
  NANDN U1659 ( .A(n1639), .B(n1640), .Z(n1638) );
  OR U1660 ( .A(n1641), .B(n1642), .Z(n1640) );
  NAND U1661 ( .A(n1642), .B(n1641), .Z(n1637) );
  ANDN U1662 ( .B(B[61]), .A(n61), .Z(n1520) );
  XNOR U1663 ( .A(n1528), .B(n1643), .Z(n1521) );
  XNOR U1664 ( .A(n1527), .B(n1525), .Z(n1643) );
  AND U1665 ( .A(n1644), .B(n1645), .Z(n1525) );
  NANDN U1666 ( .A(n1646), .B(n1647), .Z(n1645) );
  NANDN U1667 ( .A(n1648), .B(n1649), .Z(n1647) );
  NANDN U1668 ( .A(n1649), .B(n1648), .Z(n1644) );
  ANDN U1669 ( .B(B[62]), .A(n62), .Z(n1527) );
  XNOR U1670 ( .A(n1535), .B(n1650), .Z(n1528) );
  XNOR U1671 ( .A(n1534), .B(n1532), .Z(n1650) );
  AND U1672 ( .A(n1651), .B(n1652), .Z(n1532) );
  NANDN U1673 ( .A(n1653), .B(n1654), .Z(n1652) );
  OR U1674 ( .A(n1655), .B(n1656), .Z(n1654) );
  NAND U1675 ( .A(n1656), .B(n1655), .Z(n1651) );
  ANDN U1676 ( .B(B[63]), .A(n63), .Z(n1534) );
  XNOR U1677 ( .A(n1542), .B(n1657), .Z(n1535) );
  XNOR U1678 ( .A(n1541), .B(n1539), .Z(n1657) );
  AND U1679 ( .A(n1658), .B(n1659), .Z(n1539) );
  NANDN U1680 ( .A(n1660), .B(n1661), .Z(n1659) );
  NANDN U1681 ( .A(n1662), .B(n1663), .Z(n1661) );
  NANDN U1682 ( .A(n1663), .B(n1662), .Z(n1658) );
  ANDN U1683 ( .B(B[64]), .A(n64), .Z(n1541) );
  XNOR U1684 ( .A(n1549), .B(n1664), .Z(n1542) );
  XNOR U1685 ( .A(n1548), .B(n1546), .Z(n1664) );
  AND U1686 ( .A(n1665), .B(n1666), .Z(n1546) );
  NANDN U1687 ( .A(n1667), .B(n1668), .Z(n1666) );
  OR U1688 ( .A(n1669), .B(n1670), .Z(n1668) );
  NAND U1689 ( .A(n1670), .B(n1669), .Z(n1665) );
  ANDN U1690 ( .B(B[65]), .A(n65), .Z(n1548) );
  XNOR U1691 ( .A(n1556), .B(n1671), .Z(n1549) );
  XNOR U1692 ( .A(n1555), .B(n1553), .Z(n1671) );
  AND U1693 ( .A(n1672), .B(n1673), .Z(n1553) );
  NANDN U1694 ( .A(n1674), .B(n1675), .Z(n1673) );
  NANDN U1695 ( .A(n1676), .B(n1677), .Z(n1675) );
  NANDN U1696 ( .A(n1677), .B(n1676), .Z(n1672) );
  ANDN U1697 ( .B(B[66]), .A(n66), .Z(n1555) );
  XNOR U1698 ( .A(n1563), .B(n1678), .Z(n1556) );
  XNOR U1699 ( .A(n1562), .B(n1560), .Z(n1678) );
  AND U1700 ( .A(n1679), .B(n1680), .Z(n1560) );
  NANDN U1701 ( .A(n1681), .B(n1682), .Z(n1680) );
  OR U1702 ( .A(n1683), .B(n1684), .Z(n1682) );
  NAND U1703 ( .A(n1684), .B(n1683), .Z(n1679) );
  ANDN U1704 ( .B(B[67]), .A(n67), .Z(n1562) );
  XNOR U1705 ( .A(n1570), .B(n1685), .Z(n1563) );
  XNOR U1706 ( .A(n1569), .B(n1567), .Z(n1685) );
  AND U1707 ( .A(n1686), .B(n1687), .Z(n1567) );
  NANDN U1708 ( .A(n1688), .B(n1689), .Z(n1687) );
  NANDN U1709 ( .A(n1690), .B(n1691), .Z(n1689) );
  NANDN U1710 ( .A(n1691), .B(n1690), .Z(n1686) );
  ANDN U1711 ( .B(B[68]), .A(n68), .Z(n1569) );
  XOR U1712 ( .A(n1575), .B(n1692), .Z(n1570) );
  XNOR U1713 ( .A(n1576), .B(n1577), .Z(n1692) );
  AND U1714 ( .A(n1693), .B(n1694), .Z(n1577) );
  NANDN U1715 ( .A(n1695), .B(n1696), .Z(n1694) );
  NANDN U1716 ( .A(n1697), .B(n1698), .Z(n1696) );
  ANDN U1717 ( .B(B[69]), .A(n69), .Z(n1576) );
  XOR U1718 ( .A(n1699), .B(n1700), .Z(n1575) );
  XNOR U1719 ( .A(n1701), .B(n34), .Z(n1700) );
  NAND U1720 ( .A(n1702), .B(n1703), .Z(n117) );
  NANDN U1721 ( .A(n1704), .B(n1705), .Z(n1703) );
  OR U1722 ( .A(n1706), .B(n1707), .Z(n1705) );
  NAND U1723 ( .A(n1707), .B(n1706), .Z(n1702) );
  XOR U1724 ( .A(n119), .B(n118), .Z(\A1[82] ) );
  XOR U1725 ( .A(n1707), .B(n1708), .Z(n118) );
  XNOR U1726 ( .A(n1706), .B(n1704), .Z(n1708) );
  AND U1727 ( .A(n1709), .B(n1710), .Z(n1704) );
  NANDN U1728 ( .A(n1711), .B(n1712), .Z(n1710) );
  NANDN U1729 ( .A(n1713), .B(n1714), .Z(n1712) );
  NANDN U1730 ( .A(n1714), .B(n1713), .Z(n1709) );
  ANDN U1731 ( .B(B[53]), .A(n54), .Z(n1706) );
  XNOR U1732 ( .A(n1593), .B(n1715), .Z(n1707) );
  XNOR U1733 ( .A(n1592), .B(n1590), .Z(n1715) );
  AND U1734 ( .A(n1716), .B(n1717), .Z(n1590) );
  NANDN U1735 ( .A(n1718), .B(n1719), .Z(n1717) );
  OR U1736 ( .A(n1720), .B(n1721), .Z(n1719) );
  NAND U1737 ( .A(n1721), .B(n1720), .Z(n1716) );
  ANDN U1738 ( .B(B[54]), .A(n55), .Z(n1592) );
  XNOR U1739 ( .A(n1600), .B(n1722), .Z(n1593) );
  XNOR U1740 ( .A(n1599), .B(n1597), .Z(n1722) );
  AND U1741 ( .A(n1723), .B(n1724), .Z(n1597) );
  NANDN U1742 ( .A(n1725), .B(n1726), .Z(n1724) );
  NANDN U1743 ( .A(n1727), .B(n1728), .Z(n1726) );
  NANDN U1744 ( .A(n1728), .B(n1727), .Z(n1723) );
  ANDN U1745 ( .B(B[55]), .A(n56), .Z(n1599) );
  XNOR U1746 ( .A(n1607), .B(n1729), .Z(n1600) );
  XNOR U1747 ( .A(n1606), .B(n1604), .Z(n1729) );
  AND U1748 ( .A(n1730), .B(n1731), .Z(n1604) );
  NANDN U1749 ( .A(n1732), .B(n1733), .Z(n1731) );
  OR U1750 ( .A(n1734), .B(n1735), .Z(n1733) );
  NAND U1751 ( .A(n1735), .B(n1734), .Z(n1730) );
  ANDN U1752 ( .B(B[56]), .A(n57), .Z(n1606) );
  XNOR U1753 ( .A(n1614), .B(n1736), .Z(n1607) );
  XNOR U1754 ( .A(n1613), .B(n1611), .Z(n1736) );
  AND U1755 ( .A(n1737), .B(n1738), .Z(n1611) );
  NANDN U1756 ( .A(n1739), .B(n1740), .Z(n1738) );
  NANDN U1757 ( .A(n1741), .B(n1742), .Z(n1740) );
  NANDN U1758 ( .A(n1742), .B(n1741), .Z(n1737) );
  ANDN U1759 ( .B(B[57]), .A(n58), .Z(n1613) );
  XNOR U1760 ( .A(n1621), .B(n1743), .Z(n1614) );
  XNOR U1761 ( .A(n1620), .B(n1618), .Z(n1743) );
  AND U1762 ( .A(n1744), .B(n1745), .Z(n1618) );
  NANDN U1763 ( .A(n1746), .B(n1747), .Z(n1745) );
  OR U1764 ( .A(n1748), .B(n1749), .Z(n1747) );
  NAND U1765 ( .A(n1749), .B(n1748), .Z(n1744) );
  ANDN U1766 ( .B(B[58]), .A(n59), .Z(n1620) );
  XNOR U1767 ( .A(n1628), .B(n1750), .Z(n1621) );
  XNOR U1768 ( .A(n1627), .B(n1625), .Z(n1750) );
  AND U1769 ( .A(n1751), .B(n1752), .Z(n1625) );
  NANDN U1770 ( .A(n1753), .B(n1754), .Z(n1752) );
  NANDN U1771 ( .A(n1755), .B(n1756), .Z(n1754) );
  NANDN U1772 ( .A(n1756), .B(n1755), .Z(n1751) );
  ANDN U1773 ( .B(B[59]), .A(n60), .Z(n1627) );
  XNOR U1774 ( .A(n1635), .B(n1757), .Z(n1628) );
  XNOR U1775 ( .A(n1634), .B(n1632), .Z(n1757) );
  AND U1776 ( .A(n1758), .B(n1759), .Z(n1632) );
  NANDN U1777 ( .A(n1760), .B(n1761), .Z(n1759) );
  OR U1778 ( .A(n1762), .B(n1763), .Z(n1761) );
  NAND U1779 ( .A(n1763), .B(n1762), .Z(n1758) );
  ANDN U1780 ( .B(B[60]), .A(n61), .Z(n1634) );
  XNOR U1781 ( .A(n1642), .B(n1764), .Z(n1635) );
  XNOR U1782 ( .A(n1641), .B(n1639), .Z(n1764) );
  AND U1783 ( .A(n1765), .B(n1766), .Z(n1639) );
  NANDN U1784 ( .A(n1767), .B(n1768), .Z(n1766) );
  NANDN U1785 ( .A(n1769), .B(n1770), .Z(n1768) );
  NANDN U1786 ( .A(n1770), .B(n1769), .Z(n1765) );
  ANDN U1787 ( .B(B[61]), .A(n62), .Z(n1641) );
  XNOR U1788 ( .A(n1649), .B(n1771), .Z(n1642) );
  XNOR U1789 ( .A(n1648), .B(n1646), .Z(n1771) );
  AND U1790 ( .A(n1772), .B(n1773), .Z(n1646) );
  NANDN U1791 ( .A(n1774), .B(n1775), .Z(n1773) );
  OR U1792 ( .A(n1776), .B(n1777), .Z(n1775) );
  NAND U1793 ( .A(n1777), .B(n1776), .Z(n1772) );
  ANDN U1794 ( .B(B[62]), .A(n63), .Z(n1648) );
  XNOR U1795 ( .A(n1656), .B(n1778), .Z(n1649) );
  XNOR U1796 ( .A(n1655), .B(n1653), .Z(n1778) );
  AND U1797 ( .A(n1779), .B(n1780), .Z(n1653) );
  NANDN U1798 ( .A(n1781), .B(n1782), .Z(n1780) );
  NANDN U1799 ( .A(n1783), .B(n1784), .Z(n1782) );
  NANDN U1800 ( .A(n1784), .B(n1783), .Z(n1779) );
  ANDN U1801 ( .B(B[63]), .A(n64), .Z(n1655) );
  XNOR U1802 ( .A(n1663), .B(n1785), .Z(n1656) );
  XNOR U1803 ( .A(n1662), .B(n1660), .Z(n1785) );
  AND U1804 ( .A(n1786), .B(n1787), .Z(n1660) );
  NANDN U1805 ( .A(n1788), .B(n1789), .Z(n1787) );
  OR U1806 ( .A(n1790), .B(n1791), .Z(n1789) );
  NAND U1807 ( .A(n1791), .B(n1790), .Z(n1786) );
  ANDN U1808 ( .B(B[64]), .A(n65), .Z(n1662) );
  XNOR U1809 ( .A(n1670), .B(n1792), .Z(n1663) );
  XNOR U1810 ( .A(n1669), .B(n1667), .Z(n1792) );
  AND U1811 ( .A(n1793), .B(n1794), .Z(n1667) );
  NANDN U1812 ( .A(n1795), .B(n1796), .Z(n1794) );
  NANDN U1813 ( .A(n1797), .B(n1798), .Z(n1796) );
  NANDN U1814 ( .A(n1798), .B(n1797), .Z(n1793) );
  ANDN U1815 ( .B(B[65]), .A(n66), .Z(n1669) );
  XNOR U1816 ( .A(n1677), .B(n1799), .Z(n1670) );
  XNOR U1817 ( .A(n1676), .B(n1674), .Z(n1799) );
  AND U1818 ( .A(n1800), .B(n1801), .Z(n1674) );
  NANDN U1819 ( .A(n1802), .B(n1803), .Z(n1801) );
  OR U1820 ( .A(n1804), .B(n1805), .Z(n1803) );
  NAND U1821 ( .A(n1805), .B(n1804), .Z(n1800) );
  ANDN U1822 ( .B(B[66]), .A(n67), .Z(n1676) );
  XNOR U1823 ( .A(n1684), .B(n1806), .Z(n1677) );
  XNOR U1824 ( .A(n1683), .B(n1681), .Z(n1806) );
  AND U1825 ( .A(n1807), .B(n1808), .Z(n1681) );
  NANDN U1826 ( .A(n1809), .B(n1810), .Z(n1808) );
  NANDN U1827 ( .A(n1811), .B(n1812), .Z(n1810) );
  NANDN U1828 ( .A(n1812), .B(n1811), .Z(n1807) );
  ANDN U1829 ( .B(B[67]), .A(n68), .Z(n1683) );
  XNOR U1830 ( .A(n1691), .B(n1813), .Z(n1684) );
  XNOR U1831 ( .A(n1690), .B(n1688), .Z(n1813) );
  AND U1832 ( .A(n1814), .B(n1815), .Z(n1688) );
  NANDN U1833 ( .A(n1816), .B(n1817), .Z(n1815) );
  OR U1834 ( .A(n1818), .B(n1819), .Z(n1817) );
  NAND U1835 ( .A(n1819), .B(n1818), .Z(n1814) );
  ANDN U1836 ( .B(B[68]), .A(n69), .Z(n1690) );
  XOR U1837 ( .A(n1695), .B(n1820), .Z(n1691) );
  XNOR U1838 ( .A(n1697), .B(n1698), .Z(n1820) );
  AND U1839 ( .A(n1821), .B(n1822), .Z(n1698) );
  NAND U1840 ( .A(n1823), .B(n1824), .Z(n1822) );
  NANDN U1841 ( .A(n1825), .B(n1826), .Z(n1823) );
  ANDN U1842 ( .B(B[69]), .A(n70), .Z(n1697) );
  XNOR U1843 ( .A(n1827), .B(n1828), .Z(n1695) );
  XNOR U1844 ( .A(n1829), .B(n35), .Z(n1828) );
  NAND U1845 ( .A(n1830), .B(n1831), .Z(n119) );
  NANDN U1846 ( .A(n1832), .B(n1833), .Z(n1831) );
  OR U1847 ( .A(n1834), .B(n1835), .Z(n1833) );
  NAND U1848 ( .A(n1835), .B(n1834), .Z(n1830) );
  XOR U1849 ( .A(n121), .B(n120), .Z(\A1[81] ) );
  XOR U1850 ( .A(n1835), .B(n1836), .Z(n120) );
  XNOR U1851 ( .A(n1834), .B(n1832), .Z(n1836) );
  AND U1852 ( .A(n1837), .B(n1838), .Z(n1832) );
  NANDN U1853 ( .A(n1839), .B(n1840), .Z(n1838) );
  NANDN U1854 ( .A(n1841), .B(n1842), .Z(n1840) );
  NANDN U1855 ( .A(n1842), .B(n1841), .Z(n1837) );
  ANDN U1856 ( .B(B[52]), .A(n54), .Z(n1834) );
  XNOR U1857 ( .A(n1714), .B(n1843), .Z(n1835) );
  XNOR U1858 ( .A(n1713), .B(n1711), .Z(n1843) );
  AND U1859 ( .A(n1844), .B(n1845), .Z(n1711) );
  NANDN U1860 ( .A(n1846), .B(n1847), .Z(n1845) );
  OR U1861 ( .A(n1848), .B(n1849), .Z(n1847) );
  NAND U1862 ( .A(n1849), .B(n1848), .Z(n1844) );
  ANDN U1863 ( .B(B[53]), .A(n55), .Z(n1713) );
  XNOR U1864 ( .A(n1721), .B(n1850), .Z(n1714) );
  XNOR U1865 ( .A(n1720), .B(n1718), .Z(n1850) );
  AND U1866 ( .A(n1851), .B(n1852), .Z(n1718) );
  NANDN U1867 ( .A(n1853), .B(n1854), .Z(n1852) );
  NANDN U1868 ( .A(n1855), .B(n1856), .Z(n1854) );
  NANDN U1869 ( .A(n1856), .B(n1855), .Z(n1851) );
  ANDN U1870 ( .B(B[54]), .A(n56), .Z(n1720) );
  XNOR U1871 ( .A(n1728), .B(n1857), .Z(n1721) );
  XNOR U1872 ( .A(n1727), .B(n1725), .Z(n1857) );
  AND U1873 ( .A(n1858), .B(n1859), .Z(n1725) );
  NANDN U1874 ( .A(n1860), .B(n1861), .Z(n1859) );
  OR U1875 ( .A(n1862), .B(n1863), .Z(n1861) );
  NAND U1876 ( .A(n1863), .B(n1862), .Z(n1858) );
  ANDN U1877 ( .B(B[55]), .A(n57), .Z(n1727) );
  XNOR U1878 ( .A(n1735), .B(n1864), .Z(n1728) );
  XNOR U1879 ( .A(n1734), .B(n1732), .Z(n1864) );
  AND U1880 ( .A(n1865), .B(n1866), .Z(n1732) );
  NANDN U1881 ( .A(n1867), .B(n1868), .Z(n1866) );
  NANDN U1882 ( .A(n1869), .B(n1870), .Z(n1868) );
  NANDN U1883 ( .A(n1870), .B(n1869), .Z(n1865) );
  ANDN U1884 ( .B(B[56]), .A(n58), .Z(n1734) );
  XNOR U1885 ( .A(n1742), .B(n1871), .Z(n1735) );
  XNOR U1886 ( .A(n1741), .B(n1739), .Z(n1871) );
  AND U1887 ( .A(n1872), .B(n1873), .Z(n1739) );
  NANDN U1888 ( .A(n1874), .B(n1875), .Z(n1873) );
  OR U1889 ( .A(n1876), .B(n1877), .Z(n1875) );
  NAND U1890 ( .A(n1877), .B(n1876), .Z(n1872) );
  ANDN U1891 ( .B(B[57]), .A(n59), .Z(n1741) );
  XNOR U1892 ( .A(n1749), .B(n1878), .Z(n1742) );
  XNOR U1893 ( .A(n1748), .B(n1746), .Z(n1878) );
  AND U1894 ( .A(n1879), .B(n1880), .Z(n1746) );
  NANDN U1895 ( .A(n1881), .B(n1882), .Z(n1880) );
  NANDN U1896 ( .A(n1883), .B(n1884), .Z(n1882) );
  NANDN U1897 ( .A(n1884), .B(n1883), .Z(n1879) );
  ANDN U1898 ( .B(B[58]), .A(n60), .Z(n1748) );
  XNOR U1899 ( .A(n1756), .B(n1885), .Z(n1749) );
  XNOR U1900 ( .A(n1755), .B(n1753), .Z(n1885) );
  AND U1901 ( .A(n1886), .B(n1887), .Z(n1753) );
  NANDN U1902 ( .A(n1888), .B(n1889), .Z(n1887) );
  OR U1903 ( .A(n1890), .B(n1891), .Z(n1889) );
  NAND U1904 ( .A(n1891), .B(n1890), .Z(n1886) );
  ANDN U1905 ( .B(B[59]), .A(n61), .Z(n1755) );
  XNOR U1906 ( .A(n1763), .B(n1892), .Z(n1756) );
  XNOR U1907 ( .A(n1762), .B(n1760), .Z(n1892) );
  AND U1908 ( .A(n1893), .B(n1894), .Z(n1760) );
  NANDN U1909 ( .A(n1895), .B(n1896), .Z(n1894) );
  NANDN U1910 ( .A(n1897), .B(n1898), .Z(n1896) );
  NANDN U1911 ( .A(n1898), .B(n1897), .Z(n1893) );
  ANDN U1912 ( .B(B[60]), .A(n62), .Z(n1762) );
  XNOR U1913 ( .A(n1770), .B(n1899), .Z(n1763) );
  XNOR U1914 ( .A(n1769), .B(n1767), .Z(n1899) );
  AND U1915 ( .A(n1900), .B(n1901), .Z(n1767) );
  NANDN U1916 ( .A(n1902), .B(n1903), .Z(n1901) );
  OR U1917 ( .A(n1904), .B(n1905), .Z(n1903) );
  NAND U1918 ( .A(n1905), .B(n1904), .Z(n1900) );
  ANDN U1919 ( .B(B[61]), .A(n63), .Z(n1769) );
  XNOR U1920 ( .A(n1777), .B(n1906), .Z(n1770) );
  XNOR U1921 ( .A(n1776), .B(n1774), .Z(n1906) );
  AND U1922 ( .A(n1907), .B(n1908), .Z(n1774) );
  NANDN U1923 ( .A(n1909), .B(n1910), .Z(n1908) );
  NANDN U1924 ( .A(n1911), .B(n1912), .Z(n1910) );
  NANDN U1925 ( .A(n1912), .B(n1911), .Z(n1907) );
  ANDN U1926 ( .B(B[62]), .A(n64), .Z(n1776) );
  XNOR U1927 ( .A(n1784), .B(n1913), .Z(n1777) );
  XNOR U1928 ( .A(n1783), .B(n1781), .Z(n1913) );
  AND U1929 ( .A(n1914), .B(n1915), .Z(n1781) );
  NANDN U1930 ( .A(n1916), .B(n1917), .Z(n1915) );
  OR U1931 ( .A(n1918), .B(n1919), .Z(n1917) );
  NAND U1932 ( .A(n1919), .B(n1918), .Z(n1914) );
  ANDN U1933 ( .B(B[63]), .A(n65), .Z(n1783) );
  XNOR U1934 ( .A(n1791), .B(n1920), .Z(n1784) );
  XNOR U1935 ( .A(n1790), .B(n1788), .Z(n1920) );
  AND U1936 ( .A(n1921), .B(n1922), .Z(n1788) );
  NANDN U1937 ( .A(n1923), .B(n1924), .Z(n1922) );
  NANDN U1938 ( .A(n1925), .B(n1926), .Z(n1924) );
  NANDN U1939 ( .A(n1926), .B(n1925), .Z(n1921) );
  ANDN U1940 ( .B(B[64]), .A(n66), .Z(n1790) );
  XNOR U1941 ( .A(n1798), .B(n1927), .Z(n1791) );
  XNOR U1942 ( .A(n1797), .B(n1795), .Z(n1927) );
  AND U1943 ( .A(n1928), .B(n1929), .Z(n1795) );
  NANDN U1944 ( .A(n1930), .B(n1931), .Z(n1929) );
  OR U1945 ( .A(n1932), .B(n1933), .Z(n1931) );
  NAND U1946 ( .A(n1933), .B(n1932), .Z(n1928) );
  ANDN U1947 ( .B(B[65]), .A(n67), .Z(n1797) );
  XNOR U1948 ( .A(n1805), .B(n1934), .Z(n1798) );
  XNOR U1949 ( .A(n1804), .B(n1802), .Z(n1934) );
  AND U1950 ( .A(n1935), .B(n1936), .Z(n1802) );
  NANDN U1951 ( .A(n1937), .B(n1938), .Z(n1936) );
  NANDN U1952 ( .A(n1939), .B(n1940), .Z(n1938) );
  NANDN U1953 ( .A(n1940), .B(n1939), .Z(n1935) );
  ANDN U1954 ( .B(B[66]), .A(n68), .Z(n1804) );
  XNOR U1955 ( .A(n1812), .B(n1941), .Z(n1805) );
  XNOR U1956 ( .A(n1811), .B(n1809), .Z(n1941) );
  AND U1957 ( .A(n1942), .B(n1943), .Z(n1809) );
  NANDN U1958 ( .A(n1944), .B(n1945), .Z(n1943) );
  OR U1959 ( .A(n1946), .B(n1947), .Z(n1945) );
  NAND U1960 ( .A(n1947), .B(n1946), .Z(n1942) );
  ANDN U1961 ( .B(B[67]), .A(n69), .Z(n1811) );
  XNOR U1962 ( .A(n1819), .B(n1948), .Z(n1812) );
  XNOR U1963 ( .A(n1818), .B(n1816), .Z(n1948) );
  AND U1964 ( .A(n1949), .B(n1950), .Z(n1816) );
  NANDN U1965 ( .A(n1951), .B(n1952), .Z(n1950) );
  NANDN U1966 ( .A(n1953), .B(n1954), .Z(n1952) );
  NANDN U1967 ( .A(n1954), .B(n1953), .Z(n1949) );
  ANDN U1968 ( .B(B[68]), .A(n70), .Z(n1818) );
  XOR U1969 ( .A(n1824), .B(n1955), .Z(n1819) );
  XNOR U1970 ( .A(n1825), .B(n1826), .Z(n1955) );
  AND U1971 ( .A(n1956), .B(n1957), .Z(n1826) );
  NANDN U1972 ( .A(n1958), .B(n1959), .Z(n1957) );
  NANDN U1973 ( .A(n1960), .B(n1961), .Z(n1959) );
  ANDN U1974 ( .B(B[69]), .A(n71), .Z(n1825) );
  XOR U1975 ( .A(n1962), .B(n1963), .Z(n1824) );
  XNOR U1976 ( .A(n1964), .B(n36), .Z(n1963) );
  NAND U1977 ( .A(n1965), .B(n1966), .Z(n121) );
  NANDN U1978 ( .A(n1967), .B(n1968), .Z(n1966) );
  OR U1979 ( .A(n1969), .B(n1970), .Z(n1968) );
  NAND U1980 ( .A(n1970), .B(n1969), .Z(n1965) );
  XOR U1981 ( .A(n123), .B(n122), .Z(\A1[80] ) );
  XOR U1982 ( .A(n1970), .B(n1971), .Z(n122) );
  XNOR U1983 ( .A(n1969), .B(n1967), .Z(n1971) );
  AND U1984 ( .A(n1972), .B(n1973), .Z(n1967) );
  NANDN U1985 ( .A(n1974), .B(n1975), .Z(n1973) );
  NANDN U1986 ( .A(n1976), .B(n1977), .Z(n1975) );
  NANDN U1987 ( .A(n1977), .B(n1976), .Z(n1972) );
  ANDN U1988 ( .B(B[51]), .A(n54), .Z(n1969) );
  XNOR U1989 ( .A(n1842), .B(n1978), .Z(n1970) );
  XNOR U1990 ( .A(n1841), .B(n1839), .Z(n1978) );
  AND U1991 ( .A(n1979), .B(n1980), .Z(n1839) );
  NANDN U1992 ( .A(n1981), .B(n1982), .Z(n1980) );
  OR U1993 ( .A(n1983), .B(n1984), .Z(n1982) );
  NAND U1994 ( .A(n1984), .B(n1983), .Z(n1979) );
  ANDN U1995 ( .B(B[52]), .A(n55), .Z(n1841) );
  XNOR U1996 ( .A(n1849), .B(n1985), .Z(n1842) );
  XNOR U1997 ( .A(n1848), .B(n1846), .Z(n1985) );
  AND U1998 ( .A(n1986), .B(n1987), .Z(n1846) );
  NANDN U1999 ( .A(n1988), .B(n1989), .Z(n1987) );
  NANDN U2000 ( .A(n1990), .B(n1991), .Z(n1989) );
  NANDN U2001 ( .A(n1991), .B(n1990), .Z(n1986) );
  ANDN U2002 ( .B(B[53]), .A(n56), .Z(n1848) );
  XNOR U2003 ( .A(n1856), .B(n1992), .Z(n1849) );
  XNOR U2004 ( .A(n1855), .B(n1853), .Z(n1992) );
  AND U2005 ( .A(n1993), .B(n1994), .Z(n1853) );
  NANDN U2006 ( .A(n1995), .B(n1996), .Z(n1994) );
  OR U2007 ( .A(n1997), .B(n1998), .Z(n1996) );
  NAND U2008 ( .A(n1998), .B(n1997), .Z(n1993) );
  ANDN U2009 ( .B(B[54]), .A(n57), .Z(n1855) );
  XNOR U2010 ( .A(n1863), .B(n1999), .Z(n1856) );
  XNOR U2011 ( .A(n1862), .B(n1860), .Z(n1999) );
  AND U2012 ( .A(n2000), .B(n2001), .Z(n1860) );
  NANDN U2013 ( .A(n2002), .B(n2003), .Z(n2001) );
  NANDN U2014 ( .A(n2004), .B(n2005), .Z(n2003) );
  NANDN U2015 ( .A(n2005), .B(n2004), .Z(n2000) );
  ANDN U2016 ( .B(B[55]), .A(n58), .Z(n1862) );
  XNOR U2017 ( .A(n1870), .B(n2006), .Z(n1863) );
  XNOR U2018 ( .A(n1869), .B(n1867), .Z(n2006) );
  AND U2019 ( .A(n2007), .B(n2008), .Z(n1867) );
  NANDN U2020 ( .A(n2009), .B(n2010), .Z(n2008) );
  OR U2021 ( .A(n2011), .B(n2012), .Z(n2010) );
  NAND U2022 ( .A(n2012), .B(n2011), .Z(n2007) );
  ANDN U2023 ( .B(B[56]), .A(n59), .Z(n1869) );
  XNOR U2024 ( .A(n1877), .B(n2013), .Z(n1870) );
  XNOR U2025 ( .A(n1876), .B(n1874), .Z(n2013) );
  AND U2026 ( .A(n2014), .B(n2015), .Z(n1874) );
  NANDN U2027 ( .A(n2016), .B(n2017), .Z(n2015) );
  NANDN U2028 ( .A(n2018), .B(n2019), .Z(n2017) );
  NANDN U2029 ( .A(n2019), .B(n2018), .Z(n2014) );
  ANDN U2030 ( .B(B[57]), .A(n60), .Z(n1876) );
  XNOR U2031 ( .A(n1884), .B(n2020), .Z(n1877) );
  XNOR U2032 ( .A(n1883), .B(n1881), .Z(n2020) );
  AND U2033 ( .A(n2021), .B(n2022), .Z(n1881) );
  NANDN U2034 ( .A(n2023), .B(n2024), .Z(n2022) );
  OR U2035 ( .A(n2025), .B(n2026), .Z(n2024) );
  NAND U2036 ( .A(n2026), .B(n2025), .Z(n2021) );
  ANDN U2037 ( .B(B[58]), .A(n61), .Z(n1883) );
  XNOR U2038 ( .A(n1891), .B(n2027), .Z(n1884) );
  XNOR U2039 ( .A(n1890), .B(n1888), .Z(n2027) );
  AND U2040 ( .A(n2028), .B(n2029), .Z(n1888) );
  NANDN U2041 ( .A(n2030), .B(n2031), .Z(n2029) );
  NANDN U2042 ( .A(n2032), .B(n2033), .Z(n2031) );
  NANDN U2043 ( .A(n2033), .B(n2032), .Z(n2028) );
  ANDN U2044 ( .B(B[59]), .A(n62), .Z(n1890) );
  XNOR U2045 ( .A(n1898), .B(n2034), .Z(n1891) );
  XNOR U2046 ( .A(n1897), .B(n1895), .Z(n2034) );
  AND U2047 ( .A(n2035), .B(n2036), .Z(n1895) );
  NANDN U2048 ( .A(n2037), .B(n2038), .Z(n2036) );
  OR U2049 ( .A(n2039), .B(n2040), .Z(n2038) );
  NAND U2050 ( .A(n2040), .B(n2039), .Z(n2035) );
  ANDN U2051 ( .B(B[60]), .A(n63), .Z(n1897) );
  XNOR U2052 ( .A(n1905), .B(n2041), .Z(n1898) );
  XNOR U2053 ( .A(n1904), .B(n1902), .Z(n2041) );
  AND U2054 ( .A(n2042), .B(n2043), .Z(n1902) );
  NANDN U2055 ( .A(n2044), .B(n2045), .Z(n2043) );
  NANDN U2056 ( .A(n2046), .B(n2047), .Z(n2045) );
  NANDN U2057 ( .A(n2047), .B(n2046), .Z(n2042) );
  ANDN U2058 ( .B(B[61]), .A(n64), .Z(n1904) );
  XNOR U2059 ( .A(n1912), .B(n2048), .Z(n1905) );
  XNOR U2060 ( .A(n1911), .B(n1909), .Z(n2048) );
  AND U2061 ( .A(n2049), .B(n2050), .Z(n1909) );
  NANDN U2062 ( .A(n2051), .B(n2052), .Z(n2050) );
  OR U2063 ( .A(n2053), .B(n2054), .Z(n2052) );
  NAND U2064 ( .A(n2054), .B(n2053), .Z(n2049) );
  ANDN U2065 ( .B(B[62]), .A(n65), .Z(n1911) );
  XNOR U2066 ( .A(n1919), .B(n2055), .Z(n1912) );
  XNOR U2067 ( .A(n1918), .B(n1916), .Z(n2055) );
  AND U2068 ( .A(n2056), .B(n2057), .Z(n1916) );
  NANDN U2069 ( .A(n2058), .B(n2059), .Z(n2057) );
  NANDN U2070 ( .A(n2060), .B(n2061), .Z(n2059) );
  NANDN U2071 ( .A(n2061), .B(n2060), .Z(n2056) );
  ANDN U2072 ( .B(B[63]), .A(n66), .Z(n1918) );
  XNOR U2073 ( .A(n1926), .B(n2062), .Z(n1919) );
  XNOR U2074 ( .A(n1925), .B(n1923), .Z(n2062) );
  AND U2075 ( .A(n2063), .B(n2064), .Z(n1923) );
  NANDN U2076 ( .A(n2065), .B(n2066), .Z(n2064) );
  OR U2077 ( .A(n2067), .B(n2068), .Z(n2066) );
  NAND U2078 ( .A(n2068), .B(n2067), .Z(n2063) );
  ANDN U2079 ( .B(B[64]), .A(n67), .Z(n1925) );
  XNOR U2080 ( .A(n1933), .B(n2069), .Z(n1926) );
  XNOR U2081 ( .A(n1932), .B(n1930), .Z(n2069) );
  AND U2082 ( .A(n2070), .B(n2071), .Z(n1930) );
  NANDN U2083 ( .A(n2072), .B(n2073), .Z(n2071) );
  NANDN U2084 ( .A(n2074), .B(n2075), .Z(n2073) );
  NANDN U2085 ( .A(n2075), .B(n2074), .Z(n2070) );
  ANDN U2086 ( .B(B[65]), .A(n68), .Z(n1932) );
  XNOR U2087 ( .A(n1940), .B(n2076), .Z(n1933) );
  XNOR U2088 ( .A(n1939), .B(n1937), .Z(n2076) );
  AND U2089 ( .A(n2077), .B(n2078), .Z(n1937) );
  NANDN U2090 ( .A(n2079), .B(n2080), .Z(n2078) );
  OR U2091 ( .A(n2081), .B(n2082), .Z(n2080) );
  NAND U2092 ( .A(n2082), .B(n2081), .Z(n2077) );
  ANDN U2093 ( .B(B[66]), .A(n69), .Z(n1939) );
  XNOR U2094 ( .A(n1947), .B(n2083), .Z(n1940) );
  XNOR U2095 ( .A(n1946), .B(n1944), .Z(n2083) );
  AND U2096 ( .A(n2084), .B(n2085), .Z(n1944) );
  NANDN U2097 ( .A(n2086), .B(n2087), .Z(n2085) );
  NANDN U2098 ( .A(n2088), .B(n2089), .Z(n2087) );
  NANDN U2099 ( .A(n2089), .B(n2088), .Z(n2084) );
  ANDN U2100 ( .B(B[67]), .A(n70), .Z(n1946) );
  XNOR U2101 ( .A(n1954), .B(n2090), .Z(n1947) );
  XNOR U2102 ( .A(n1953), .B(n1951), .Z(n2090) );
  AND U2103 ( .A(n2091), .B(n2092), .Z(n1951) );
  NANDN U2104 ( .A(n2093), .B(n2094), .Z(n2092) );
  OR U2105 ( .A(n2095), .B(n2096), .Z(n2094) );
  NAND U2106 ( .A(n2096), .B(n2095), .Z(n2091) );
  ANDN U2107 ( .B(B[68]), .A(n71), .Z(n1953) );
  XOR U2108 ( .A(n1958), .B(n2097), .Z(n1954) );
  XNOR U2109 ( .A(n1960), .B(n1961), .Z(n2097) );
  AND U2110 ( .A(n2098), .B(n2099), .Z(n1961) );
  NAND U2111 ( .A(n2100), .B(n2101), .Z(n2099) );
  NANDN U2112 ( .A(n2102), .B(n2103), .Z(n2100) );
  ANDN U2113 ( .B(B[69]), .A(n72), .Z(n1960) );
  XNOR U2114 ( .A(n2104), .B(n2105), .Z(n1958) );
  XNOR U2115 ( .A(n2106), .B(n37), .Z(n2105) );
  NAND U2116 ( .A(n2107), .B(n2108), .Z(n123) );
  NANDN U2117 ( .A(n2109), .B(n2110), .Z(n2108) );
  OR U2118 ( .A(n2111), .B(n2112), .Z(n2110) );
  NAND U2119 ( .A(n2112), .B(n2111), .Z(n2107) );
  XOR U2120 ( .A(n2113), .B(n2114), .Z(\A1[7] ) );
  XNOR U2121 ( .A(n2115), .B(n50), .Z(n2114) );
  XOR U2122 ( .A(n125), .B(n124), .Z(\A1[79] ) );
  XOR U2123 ( .A(n2112), .B(n2116), .Z(n124) );
  XNOR U2124 ( .A(n2111), .B(n2109), .Z(n2116) );
  AND U2125 ( .A(n2117), .B(n2118), .Z(n2109) );
  NANDN U2126 ( .A(n2119), .B(n2120), .Z(n2118) );
  NANDN U2127 ( .A(n2121), .B(n2122), .Z(n2120) );
  NANDN U2128 ( .A(n2122), .B(n2121), .Z(n2117) );
  ANDN U2129 ( .B(B[50]), .A(n54), .Z(n2111) );
  XNOR U2130 ( .A(n1977), .B(n2123), .Z(n2112) );
  XNOR U2131 ( .A(n1976), .B(n1974), .Z(n2123) );
  AND U2132 ( .A(n2124), .B(n2125), .Z(n1974) );
  NANDN U2133 ( .A(n2126), .B(n2127), .Z(n2125) );
  OR U2134 ( .A(n2128), .B(n2129), .Z(n2127) );
  NAND U2135 ( .A(n2129), .B(n2128), .Z(n2124) );
  ANDN U2136 ( .B(B[51]), .A(n55), .Z(n1976) );
  XNOR U2137 ( .A(n1984), .B(n2130), .Z(n1977) );
  XNOR U2138 ( .A(n1983), .B(n1981), .Z(n2130) );
  AND U2139 ( .A(n2131), .B(n2132), .Z(n1981) );
  NANDN U2140 ( .A(n2133), .B(n2134), .Z(n2132) );
  NANDN U2141 ( .A(n2135), .B(n2136), .Z(n2134) );
  NANDN U2142 ( .A(n2136), .B(n2135), .Z(n2131) );
  ANDN U2143 ( .B(B[52]), .A(n56), .Z(n1983) );
  XNOR U2144 ( .A(n1991), .B(n2137), .Z(n1984) );
  XNOR U2145 ( .A(n1990), .B(n1988), .Z(n2137) );
  AND U2146 ( .A(n2138), .B(n2139), .Z(n1988) );
  NANDN U2147 ( .A(n2140), .B(n2141), .Z(n2139) );
  OR U2148 ( .A(n2142), .B(n2143), .Z(n2141) );
  NAND U2149 ( .A(n2143), .B(n2142), .Z(n2138) );
  ANDN U2150 ( .B(B[53]), .A(n57), .Z(n1990) );
  XNOR U2151 ( .A(n1998), .B(n2144), .Z(n1991) );
  XNOR U2152 ( .A(n1997), .B(n1995), .Z(n2144) );
  AND U2153 ( .A(n2145), .B(n2146), .Z(n1995) );
  NANDN U2154 ( .A(n2147), .B(n2148), .Z(n2146) );
  NANDN U2155 ( .A(n2149), .B(n2150), .Z(n2148) );
  NANDN U2156 ( .A(n2150), .B(n2149), .Z(n2145) );
  ANDN U2157 ( .B(B[54]), .A(n58), .Z(n1997) );
  XNOR U2158 ( .A(n2005), .B(n2151), .Z(n1998) );
  XNOR U2159 ( .A(n2004), .B(n2002), .Z(n2151) );
  AND U2160 ( .A(n2152), .B(n2153), .Z(n2002) );
  NANDN U2161 ( .A(n2154), .B(n2155), .Z(n2153) );
  OR U2162 ( .A(n2156), .B(n2157), .Z(n2155) );
  NAND U2163 ( .A(n2157), .B(n2156), .Z(n2152) );
  ANDN U2164 ( .B(B[55]), .A(n59), .Z(n2004) );
  XNOR U2165 ( .A(n2012), .B(n2158), .Z(n2005) );
  XNOR U2166 ( .A(n2011), .B(n2009), .Z(n2158) );
  AND U2167 ( .A(n2159), .B(n2160), .Z(n2009) );
  NANDN U2168 ( .A(n2161), .B(n2162), .Z(n2160) );
  NANDN U2169 ( .A(n2163), .B(n2164), .Z(n2162) );
  NANDN U2170 ( .A(n2164), .B(n2163), .Z(n2159) );
  ANDN U2171 ( .B(B[56]), .A(n60), .Z(n2011) );
  XNOR U2172 ( .A(n2019), .B(n2165), .Z(n2012) );
  XNOR U2173 ( .A(n2018), .B(n2016), .Z(n2165) );
  AND U2174 ( .A(n2166), .B(n2167), .Z(n2016) );
  NANDN U2175 ( .A(n2168), .B(n2169), .Z(n2167) );
  OR U2176 ( .A(n2170), .B(n2171), .Z(n2169) );
  NAND U2177 ( .A(n2171), .B(n2170), .Z(n2166) );
  ANDN U2178 ( .B(B[57]), .A(n61), .Z(n2018) );
  XNOR U2179 ( .A(n2026), .B(n2172), .Z(n2019) );
  XNOR U2180 ( .A(n2025), .B(n2023), .Z(n2172) );
  AND U2181 ( .A(n2173), .B(n2174), .Z(n2023) );
  NANDN U2182 ( .A(n2175), .B(n2176), .Z(n2174) );
  NANDN U2183 ( .A(n2177), .B(n2178), .Z(n2176) );
  NANDN U2184 ( .A(n2178), .B(n2177), .Z(n2173) );
  ANDN U2185 ( .B(B[58]), .A(n62), .Z(n2025) );
  XNOR U2186 ( .A(n2033), .B(n2179), .Z(n2026) );
  XNOR U2187 ( .A(n2032), .B(n2030), .Z(n2179) );
  AND U2188 ( .A(n2180), .B(n2181), .Z(n2030) );
  NANDN U2189 ( .A(n2182), .B(n2183), .Z(n2181) );
  OR U2190 ( .A(n2184), .B(n2185), .Z(n2183) );
  NAND U2191 ( .A(n2185), .B(n2184), .Z(n2180) );
  ANDN U2192 ( .B(B[59]), .A(n63), .Z(n2032) );
  XNOR U2193 ( .A(n2040), .B(n2186), .Z(n2033) );
  XNOR U2194 ( .A(n2039), .B(n2037), .Z(n2186) );
  AND U2195 ( .A(n2187), .B(n2188), .Z(n2037) );
  NANDN U2196 ( .A(n2189), .B(n2190), .Z(n2188) );
  NANDN U2197 ( .A(n2191), .B(n2192), .Z(n2190) );
  NANDN U2198 ( .A(n2192), .B(n2191), .Z(n2187) );
  ANDN U2199 ( .B(B[60]), .A(n64), .Z(n2039) );
  XNOR U2200 ( .A(n2047), .B(n2193), .Z(n2040) );
  XNOR U2201 ( .A(n2046), .B(n2044), .Z(n2193) );
  AND U2202 ( .A(n2194), .B(n2195), .Z(n2044) );
  NANDN U2203 ( .A(n2196), .B(n2197), .Z(n2195) );
  OR U2204 ( .A(n2198), .B(n2199), .Z(n2197) );
  NAND U2205 ( .A(n2199), .B(n2198), .Z(n2194) );
  ANDN U2206 ( .B(B[61]), .A(n65), .Z(n2046) );
  XNOR U2207 ( .A(n2054), .B(n2200), .Z(n2047) );
  XNOR U2208 ( .A(n2053), .B(n2051), .Z(n2200) );
  AND U2209 ( .A(n2201), .B(n2202), .Z(n2051) );
  NANDN U2210 ( .A(n2203), .B(n2204), .Z(n2202) );
  NANDN U2211 ( .A(n2205), .B(n2206), .Z(n2204) );
  NANDN U2212 ( .A(n2206), .B(n2205), .Z(n2201) );
  ANDN U2213 ( .B(B[62]), .A(n66), .Z(n2053) );
  XNOR U2214 ( .A(n2061), .B(n2207), .Z(n2054) );
  XNOR U2215 ( .A(n2060), .B(n2058), .Z(n2207) );
  AND U2216 ( .A(n2208), .B(n2209), .Z(n2058) );
  NANDN U2217 ( .A(n2210), .B(n2211), .Z(n2209) );
  OR U2218 ( .A(n2212), .B(n2213), .Z(n2211) );
  NAND U2219 ( .A(n2213), .B(n2212), .Z(n2208) );
  ANDN U2220 ( .B(B[63]), .A(n67), .Z(n2060) );
  XNOR U2221 ( .A(n2068), .B(n2214), .Z(n2061) );
  XNOR U2222 ( .A(n2067), .B(n2065), .Z(n2214) );
  AND U2223 ( .A(n2215), .B(n2216), .Z(n2065) );
  NANDN U2224 ( .A(n2217), .B(n2218), .Z(n2216) );
  NANDN U2225 ( .A(n2219), .B(n2220), .Z(n2218) );
  NANDN U2226 ( .A(n2220), .B(n2219), .Z(n2215) );
  ANDN U2227 ( .B(B[64]), .A(n68), .Z(n2067) );
  XNOR U2228 ( .A(n2075), .B(n2221), .Z(n2068) );
  XNOR U2229 ( .A(n2074), .B(n2072), .Z(n2221) );
  AND U2230 ( .A(n2222), .B(n2223), .Z(n2072) );
  NANDN U2231 ( .A(n2224), .B(n2225), .Z(n2223) );
  OR U2232 ( .A(n2226), .B(n2227), .Z(n2225) );
  NAND U2233 ( .A(n2227), .B(n2226), .Z(n2222) );
  ANDN U2234 ( .B(B[65]), .A(n69), .Z(n2074) );
  XNOR U2235 ( .A(n2082), .B(n2228), .Z(n2075) );
  XNOR U2236 ( .A(n2081), .B(n2079), .Z(n2228) );
  AND U2237 ( .A(n2229), .B(n2230), .Z(n2079) );
  NANDN U2238 ( .A(n2231), .B(n2232), .Z(n2230) );
  NANDN U2239 ( .A(n2233), .B(n2234), .Z(n2232) );
  NANDN U2240 ( .A(n2234), .B(n2233), .Z(n2229) );
  ANDN U2241 ( .B(B[66]), .A(n70), .Z(n2081) );
  XNOR U2242 ( .A(n2089), .B(n2235), .Z(n2082) );
  XNOR U2243 ( .A(n2088), .B(n2086), .Z(n2235) );
  AND U2244 ( .A(n2236), .B(n2237), .Z(n2086) );
  NANDN U2245 ( .A(n2238), .B(n2239), .Z(n2237) );
  OR U2246 ( .A(n2240), .B(n2241), .Z(n2239) );
  NAND U2247 ( .A(n2241), .B(n2240), .Z(n2236) );
  ANDN U2248 ( .B(B[67]), .A(n71), .Z(n2088) );
  XNOR U2249 ( .A(n2096), .B(n2242), .Z(n2089) );
  XNOR U2250 ( .A(n2095), .B(n2093), .Z(n2242) );
  AND U2251 ( .A(n2243), .B(n2244), .Z(n2093) );
  NANDN U2252 ( .A(n2245), .B(n2246), .Z(n2244) );
  NANDN U2253 ( .A(n2247), .B(n2248), .Z(n2246) );
  NANDN U2254 ( .A(n2248), .B(n2247), .Z(n2243) );
  ANDN U2255 ( .B(B[68]), .A(n72), .Z(n2095) );
  XOR U2256 ( .A(n2101), .B(n2249), .Z(n2096) );
  XNOR U2257 ( .A(n2102), .B(n2103), .Z(n2249) );
  AND U2258 ( .A(n2250), .B(n2251), .Z(n2103) );
  NANDN U2259 ( .A(n2252), .B(n2253), .Z(n2251) );
  NANDN U2260 ( .A(n2254), .B(n2255), .Z(n2253) );
  ANDN U2261 ( .B(B[69]), .A(n73), .Z(n2102) );
  XOR U2262 ( .A(n2256), .B(n2257), .Z(n2101) );
  XNOR U2263 ( .A(n2258), .B(n38), .Z(n2257) );
  NAND U2264 ( .A(n2259), .B(n2260), .Z(n125) );
  NANDN U2265 ( .A(n2261), .B(n2262), .Z(n2260) );
  OR U2266 ( .A(n2263), .B(n2264), .Z(n2262) );
  NAND U2267 ( .A(n2264), .B(n2263), .Z(n2259) );
  XOR U2268 ( .A(n127), .B(n126), .Z(\A1[78] ) );
  XOR U2269 ( .A(n2264), .B(n2265), .Z(n126) );
  XNOR U2270 ( .A(n2263), .B(n2261), .Z(n2265) );
  AND U2271 ( .A(n2266), .B(n2267), .Z(n2261) );
  NANDN U2272 ( .A(n2268), .B(n2269), .Z(n2267) );
  NANDN U2273 ( .A(n2270), .B(n2271), .Z(n2269) );
  NANDN U2274 ( .A(n2271), .B(n2270), .Z(n2266) );
  ANDN U2275 ( .B(B[49]), .A(n54), .Z(n2263) );
  XNOR U2276 ( .A(n2122), .B(n2272), .Z(n2264) );
  XNOR U2277 ( .A(n2121), .B(n2119), .Z(n2272) );
  AND U2278 ( .A(n2273), .B(n2274), .Z(n2119) );
  NANDN U2279 ( .A(n2275), .B(n2276), .Z(n2274) );
  OR U2280 ( .A(n2277), .B(n2278), .Z(n2276) );
  NAND U2281 ( .A(n2278), .B(n2277), .Z(n2273) );
  ANDN U2282 ( .B(B[50]), .A(n55), .Z(n2121) );
  XNOR U2283 ( .A(n2129), .B(n2279), .Z(n2122) );
  XNOR U2284 ( .A(n2128), .B(n2126), .Z(n2279) );
  AND U2285 ( .A(n2280), .B(n2281), .Z(n2126) );
  NANDN U2286 ( .A(n2282), .B(n2283), .Z(n2281) );
  NANDN U2287 ( .A(n2284), .B(n2285), .Z(n2283) );
  NANDN U2288 ( .A(n2285), .B(n2284), .Z(n2280) );
  ANDN U2289 ( .B(B[51]), .A(n56), .Z(n2128) );
  XNOR U2290 ( .A(n2136), .B(n2286), .Z(n2129) );
  XNOR U2291 ( .A(n2135), .B(n2133), .Z(n2286) );
  AND U2292 ( .A(n2287), .B(n2288), .Z(n2133) );
  NANDN U2293 ( .A(n2289), .B(n2290), .Z(n2288) );
  OR U2294 ( .A(n2291), .B(n2292), .Z(n2290) );
  NAND U2295 ( .A(n2292), .B(n2291), .Z(n2287) );
  ANDN U2296 ( .B(B[52]), .A(n57), .Z(n2135) );
  XNOR U2297 ( .A(n2143), .B(n2293), .Z(n2136) );
  XNOR U2298 ( .A(n2142), .B(n2140), .Z(n2293) );
  AND U2299 ( .A(n2294), .B(n2295), .Z(n2140) );
  NANDN U2300 ( .A(n2296), .B(n2297), .Z(n2295) );
  NANDN U2301 ( .A(n2298), .B(n2299), .Z(n2297) );
  NANDN U2302 ( .A(n2299), .B(n2298), .Z(n2294) );
  ANDN U2303 ( .B(B[53]), .A(n58), .Z(n2142) );
  XNOR U2304 ( .A(n2150), .B(n2300), .Z(n2143) );
  XNOR U2305 ( .A(n2149), .B(n2147), .Z(n2300) );
  AND U2306 ( .A(n2301), .B(n2302), .Z(n2147) );
  NANDN U2307 ( .A(n2303), .B(n2304), .Z(n2302) );
  OR U2308 ( .A(n2305), .B(n2306), .Z(n2304) );
  NAND U2309 ( .A(n2306), .B(n2305), .Z(n2301) );
  ANDN U2310 ( .B(B[54]), .A(n59), .Z(n2149) );
  XNOR U2311 ( .A(n2157), .B(n2307), .Z(n2150) );
  XNOR U2312 ( .A(n2156), .B(n2154), .Z(n2307) );
  AND U2313 ( .A(n2308), .B(n2309), .Z(n2154) );
  NANDN U2314 ( .A(n2310), .B(n2311), .Z(n2309) );
  NANDN U2315 ( .A(n2312), .B(n2313), .Z(n2311) );
  NANDN U2316 ( .A(n2313), .B(n2312), .Z(n2308) );
  ANDN U2317 ( .B(B[55]), .A(n60), .Z(n2156) );
  XNOR U2318 ( .A(n2164), .B(n2314), .Z(n2157) );
  XNOR U2319 ( .A(n2163), .B(n2161), .Z(n2314) );
  AND U2320 ( .A(n2315), .B(n2316), .Z(n2161) );
  NANDN U2321 ( .A(n2317), .B(n2318), .Z(n2316) );
  OR U2322 ( .A(n2319), .B(n2320), .Z(n2318) );
  NAND U2323 ( .A(n2320), .B(n2319), .Z(n2315) );
  ANDN U2324 ( .B(B[56]), .A(n61), .Z(n2163) );
  XNOR U2325 ( .A(n2171), .B(n2321), .Z(n2164) );
  XNOR U2326 ( .A(n2170), .B(n2168), .Z(n2321) );
  AND U2327 ( .A(n2322), .B(n2323), .Z(n2168) );
  NANDN U2328 ( .A(n2324), .B(n2325), .Z(n2323) );
  NANDN U2329 ( .A(n2326), .B(n2327), .Z(n2325) );
  NANDN U2330 ( .A(n2327), .B(n2326), .Z(n2322) );
  ANDN U2331 ( .B(B[57]), .A(n62), .Z(n2170) );
  XNOR U2332 ( .A(n2178), .B(n2328), .Z(n2171) );
  XNOR U2333 ( .A(n2177), .B(n2175), .Z(n2328) );
  AND U2334 ( .A(n2329), .B(n2330), .Z(n2175) );
  NANDN U2335 ( .A(n2331), .B(n2332), .Z(n2330) );
  OR U2336 ( .A(n2333), .B(n2334), .Z(n2332) );
  NAND U2337 ( .A(n2334), .B(n2333), .Z(n2329) );
  ANDN U2338 ( .B(B[58]), .A(n63), .Z(n2177) );
  XNOR U2339 ( .A(n2185), .B(n2335), .Z(n2178) );
  XNOR U2340 ( .A(n2184), .B(n2182), .Z(n2335) );
  AND U2341 ( .A(n2336), .B(n2337), .Z(n2182) );
  NANDN U2342 ( .A(n2338), .B(n2339), .Z(n2337) );
  NANDN U2343 ( .A(n2340), .B(n2341), .Z(n2339) );
  NANDN U2344 ( .A(n2341), .B(n2340), .Z(n2336) );
  ANDN U2345 ( .B(B[59]), .A(n64), .Z(n2184) );
  XNOR U2346 ( .A(n2192), .B(n2342), .Z(n2185) );
  XNOR U2347 ( .A(n2191), .B(n2189), .Z(n2342) );
  AND U2348 ( .A(n2343), .B(n2344), .Z(n2189) );
  NANDN U2349 ( .A(n2345), .B(n2346), .Z(n2344) );
  OR U2350 ( .A(n2347), .B(n2348), .Z(n2346) );
  NAND U2351 ( .A(n2348), .B(n2347), .Z(n2343) );
  ANDN U2352 ( .B(B[60]), .A(n65), .Z(n2191) );
  XNOR U2353 ( .A(n2199), .B(n2349), .Z(n2192) );
  XNOR U2354 ( .A(n2198), .B(n2196), .Z(n2349) );
  AND U2355 ( .A(n2350), .B(n2351), .Z(n2196) );
  NANDN U2356 ( .A(n2352), .B(n2353), .Z(n2351) );
  NANDN U2357 ( .A(n2354), .B(n2355), .Z(n2353) );
  NANDN U2358 ( .A(n2355), .B(n2354), .Z(n2350) );
  ANDN U2359 ( .B(B[61]), .A(n66), .Z(n2198) );
  XNOR U2360 ( .A(n2206), .B(n2356), .Z(n2199) );
  XNOR U2361 ( .A(n2205), .B(n2203), .Z(n2356) );
  AND U2362 ( .A(n2357), .B(n2358), .Z(n2203) );
  NANDN U2363 ( .A(n2359), .B(n2360), .Z(n2358) );
  OR U2364 ( .A(n2361), .B(n2362), .Z(n2360) );
  NAND U2365 ( .A(n2362), .B(n2361), .Z(n2357) );
  ANDN U2366 ( .B(B[62]), .A(n67), .Z(n2205) );
  XNOR U2367 ( .A(n2213), .B(n2363), .Z(n2206) );
  XNOR U2368 ( .A(n2212), .B(n2210), .Z(n2363) );
  AND U2369 ( .A(n2364), .B(n2365), .Z(n2210) );
  NANDN U2370 ( .A(n2366), .B(n2367), .Z(n2365) );
  NANDN U2371 ( .A(n2368), .B(n2369), .Z(n2367) );
  NANDN U2372 ( .A(n2369), .B(n2368), .Z(n2364) );
  ANDN U2373 ( .B(B[63]), .A(n68), .Z(n2212) );
  XNOR U2374 ( .A(n2220), .B(n2370), .Z(n2213) );
  XNOR U2375 ( .A(n2219), .B(n2217), .Z(n2370) );
  AND U2376 ( .A(n2371), .B(n2372), .Z(n2217) );
  NANDN U2377 ( .A(n2373), .B(n2374), .Z(n2372) );
  OR U2378 ( .A(n2375), .B(n2376), .Z(n2374) );
  NAND U2379 ( .A(n2376), .B(n2375), .Z(n2371) );
  ANDN U2380 ( .B(B[64]), .A(n69), .Z(n2219) );
  XNOR U2381 ( .A(n2227), .B(n2377), .Z(n2220) );
  XNOR U2382 ( .A(n2226), .B(n2224), .Z(n2377) );
  AND U2383 ( .A(n2378), .B(n2379), .Z(n2224) );
  NANDN U2384 ( .A(n2380), .B(n2381), .Z(n2379) );
  NANDN U2385 ( .A(n2382), .B(n2383), .Z(n2381) );
  NANDN U2386 ( .A(n2383), .B(n2382), .Z(n2378) );
  ANDN U2387 ( .B(B[65]), .A(n70), .Z(n2226) );
  XNOR U2388 ( .A(n2234), .B(n2384), .Z(n2227) );
  XNOR U2389 ( .A(n2233), .B(n2231), .Z(n2384) );
  AND U2390 ( .A(n2385), .B(n2386), .Z(n2231) );
  NANDN U2391 ( .A(n2387), .B(n2388), .Z(n2386) );
  OR U2392 ( .A(n2389), .B(n2390), .Z(n2388) );
  NAND U2393 ( .A(n2390), .B(n2389), .Z(n2385) );
  ANDN U2394 ( .B(B[66]), .A(n71), .Z(n2233) );
  XNOR U2395 ( .A(n2241), .B(n2391), .Z(n2234) );
  XNOR U2396 ( .A(n2240), .B(n2238), .Z(n2391) );
  AND U2397 ( .A(n2392), .B(n2393), .Z(n2238) );
  NANDN U2398 ( .A(n2394), .B(n2395), .Z(n2393) );
  NANDN U2399 ( .A(n2396), .B(n2397), .Z(n2395) );
  NANDN U2400 ( .A(n2397), .B(n2396), .Z(n2392) );
  ANDN U2401 ( .B(B[67]), .A(n72), .Z(n2240) );
  XNOR U2402 ( .A(n2248), .B(n2398), .Z(n2241) );
  XNOR U2403 ( .A(n2247), .B(n2245), .Z(n2398) );
  AND U2404 ( .A(n2399), .B(n2400), .Z(n2245) );
  NANDN U2405 ( .A(n2401), .B(n2402), .Z(n2400) );
  OR U2406 ( .A(n2403), .B(n2404), .Z(n2402) );
  NAND U2407 ( .A(n2404), .B(n2403), .Z(n2399) );
  ANDN U2408 ( .B(B[68]), .A(n73), .Z(n2247) );
  XOR U2409 ( .A(n2252), .B(n2405), .Z(n2248) );
  XNOR U2410 ( .A(n2254), .B(n2255), .Z(n2405) );
  AND U2411 ( .A(n2406), .B(n2407), .Z(n2255) );
  NAND U2412 ( .A(n2408), .B(n2409), .Z(n2407) );
  NANDN U2413 ( .A(n2410), .B(n2411), .Z(n2408) );
  ANDN U2414 ( .B(B[69]), .A(n74), .Z(n2254) );
  XNOR U2415 ( .A(n2412), .B(n2413), .Z(n2252) );
  XNOR U2416 ( .A(n2414), .B(n39), .Z(n2413) );
  NAND U2417 ( .A(n2415), .B(n2416), .Z(n127) );
  NANDN U2418 ( .A(n2417), .B(n2418), .Z(n2416) );
  OR U2419 ( .A(n2419), .B(n2420), .Z(n2418) );
  NAND U2420 ( .A(n2420), .B(n2419), .Z(n2415) );
  XOR U2421 ( .A(n129), .B(n128), .Z(\A1[77] ) );
  XOR U2422 ( .A(n2420), .B(n2421), .Z(n128) );
  XNOR U2423 ( .A(n2419), .B(n2417), .Z(n2421) );
  AND U2424 ( .A(n2422), .B(n2423), .Z(n2417) );
  NANDN U2425 ( .A(n2424), .B(n2425), .Z(n2423) );
  NANDN U2426 ( .A(n2426), .B(n2427), .Z(n2425) );
  NANDN U2427 ( .A(n2427), .B(n2426), .Z(n2422) );
  ANDN U2428 ( .B(B[48]), .A(n54), .Z(n2419) );
  XNOR U2429 ( .A(n2271), .B(n2428), .Z(n2420) );
  XNOR U2430 ( .A(n2270), .B(n2268), .Z(n2428) );
  AND U2431 ( .A(n2429), .B(n2430), .Z(n2268) );
  NANDN U2432 ( .A(n2431), .B(n2432), .Z(n2430) );
  OR U2433 ( .A(n2433), .B(n2434), .Z(n2432) );
  NAND U2434 ( .A(n2434), .B(n2433), .Z(n2429) );
  ANDN U2435 ( .B(B[49]), .A(n55), .Z(n2270) );
  XNOR U2436 ( .A(n2278), .B(n2435), .Z(n2271) );
  XNOR U2437 ( .A(n2277), .B(n2275), .Z(n2435) );
  AND U2438 ( .A(n2436), .B(n2437), .Z(n2275) );
  NANDN U2439 ( .A(n2438), .B(n2439), .Z(n2437) );
  NANDN U2440 ( .A(n2440), .B(n2441), .Z(n2439) );
  NANDN U2441 ( .A(n2441), .B(n2440), .Z(n2436) );
  ANDN U2442 ( .B(B[50]), .A(n56), .Z(n2277) );
  XNOR U2443 ( .A(n2285), .B(n2442), .Z(n2278) );
  XNOR U2444 ( .A(n2284), .B(n2282), .Z(n2442) );
  AND U2445 ( .A(n2443), .B(n2444), .Z(n2282) );
  NANDN U2446 ( .A(n2445), .B(n2446), .Z(n2444) );
  OR U2447 ( .A(n2447), .B(n2448), .Z(n2446) );
  NAND U2448 ( .A(n2448), .B(n2447), .Z(n2443) );
  ANDN U2449 ( .B(B[51]), .A(n57), .Z(n2284) );
  XNOR U2450 ( .A(n2292), .B(n2449), .Z(n2285) );
  XNOR U2451 ( .A(n2291), .B(n2289), .Z(n2449) );
  AND U2452 ( .A(n2450), .B(n2451), .Z(n2289) );
  NANDN U2453 ( .A(n2452), .B(n2453), .Z(n2451) );
  NANDN U2454 ( .A(n2454), .B(n2455), .Z(n2453) );
  NANDN U2455 ( .A(n2455), .B(n2454), .Z(n2450) );
  ANDN U2456 ( .B(B[52]), .A(n58), .Z(n2291) );
  XNOR U2457 ( .A(n2299), .B(n2456), .Z(n2292) );
  XNOR U2458 ( .A(n2298), .B(n2296), .Z(n2456) );
  AND U2459 ( .A(n2457), .B(n2458), .Z(n2296) );
  NANDN U2460 ( .A(n2459), .B(n2460), .Z(n2458) );
  OR U2461 ( .A(n2461), .B(n2462), .Z(n2460) );
  NAND U2462 ( .A(n2462), .B(n2461), .Z(n2457) );
  ANDN U2463 ( .B(B[53]), .A(n59), .Z(n2298) );
  XNOR U2464 ( .A(n2306), .B(n2463), .Z(n2299) );
  XNOR U2465 ( .A(n2305), .B(n2303), .Z(n2463) );
  AND U2466 ( .A(n2464), .B(n2465), .Z(n2303) );
  NANDN U2467 ( .A(n2466), .B(n2467), .Z(n2465) );
  NANDN U2468 ( .A(n2468), .B(n2469), .Z(n2467) );
  NANDN U2469 ( .A(n2469), .B(n2468), .Z(n2464) );
  ANDN U2470 ( .B(B[54]), .A(n60), .Z(n2305) );
  XNOR U2471 ( .A(n2313), .B(n2470), .Z(n2306) );
  XNOR U2472 ( .A(n2312), .B(n2310), .Z(n2470) );
  AND U2473 ( .A(n2471), .B(n2472), .Z(n2310) );
  NANDN U2474 ( .A(n2473), .B(n2474), .Z(n2472) );
  OR U2475 ( .A(n2475), .B(n2476), .Z(n2474) );
  NAND U2476 ( .A(n2476), .B(n2475), .Z(n2471) );
  ANDN U2477 ( .B(B[55]), .A(n61), .Z(n2312) );
  XNOR U2478 ( .A(n2320), .B(n2477), .Z(n2313) );
  XNOR U2479 ( .A(n2319), .B(n2317), .Z(n2477) );
  AND U2480 ( .A(n2478), .B(n2479), .Z(n2317) );
  NANDN U2481 ( .A(n2480), .B(n2481), .Z(n2479) );
  NANDN U2482 ( .A(n2482), .B(n2483), .Z(n2481) );
  NANDN U2483 ( .A(n2483), .B(n2482), .Z(n2478) );
  ANDN U2484 ( .B(B[56]), .A(n62), .Z(n2319) );
  XNOR U2485 ( .A(n2327), .B(n2484), .Z(n2320) );
  XNOR U2486 ( .A(n2326), .B(n2324), .Z(n2484) );
  AND U2487 ( .A(n2485), .B(n2486), .Z(n2324) );
  NANDN U2488 ( .A(n2487), .B(n2488), .Z(n2486) );
  OR U2489 ( .A(n2489), .B(n2490), .Z(n2488) );
  NAND U2490 ( .A(n2490), .B(n2489), .Z(n2485) );
  ANDN U2491 ( .B(B[57]), .A(n63), .Z(n2326) );
  XNOR U2492 ( .A(n2334), .B(n2491), .Z(n2327) );
  XNOR U2493 ( .A(n2333), .B(n2331), .Z(n2491) );
  AND U2494 ( .A(n2492), .B(n2493), .Z(n2331) );
  NANDN U2495 ( .A(n2494), .B(n2495), .Z(n2493) );
  NANDN U2496 ( .A(n2496), .B(n2497), .Z(n2495) );
  NANDN U2497 ( .A(n2497), .B(n2496), .Z(n2492) );
  ANDN U2498 ( .B(B[58]), .A(n64), .Z(n2333) );
  XNOR U2499 ( .A(n2341), .B(n2498), .Z(n2334) );
  XNOR U2500 ( .A(n2340), .B(n2338), .Z(n2498) );
  AND U2501 ( .A(n2499), .B(n2500), .Z(n2338) );
  NANDN U2502 ( .A(n2501), .B(n2502), .Z(n2500) );
  OR U2503 ( .A(n2503), .B(n2504), .Z(n2502) );
  NAND U2504 ( .A(n2504), .B(n2503), .Z(n2499) );
  ANDN U2505 ( .B(B[59]), .A(n65), .Z(n2340) );
  XNOR U2506 ( .A(n2348), .B(n2505), .Z(n2341) );
  XNOR U2507 ( .A(n2347), .B(n2345), .Z(n2505) );
  AND U2508 ( .A(n2506), .B(n2507), .Z(n2345) );
  NANDN U2509 ( .A(n2508), .B(n2509), .Z(n2507) );
  NANDN U2510 ( .A(n2510), .B(n2511), .Z(n2509) );
  NANDN U2511 ( .A(n2511), .B(n2510), .Z(n2506) );
  ANDN U2512 ( .B(B[60]), .A(n66), .Z(n2347) );
  XNOR U2513 ( .A(n2355), .B(n2512), .Z(n2348) );
  XNOR U2514 ( .A(n2354), .B(n2352), .Z(n2512) );
  AND U2515 ( .A(n2513), .B(n2514), .Z(n2352) );
  NANDN U2516 ( .A(n2515), .B(n2516), .Z(n2514) );
  OR U2517 ( .A(n2517), .B(n2518), .Z(n2516) );
  NAND U2518 ( .A(n2518), .B(n2517), .Z(n2513) );
  ANDN U2519 ( .B(B[61]), .A(n67), .Z(n2354) );
  XNOR U2520 ( .A(n2362), .B(n2519), .Z(n2355) );
  XNOR U2521 ( .A(n2361), .B(n2359), .Z(n2519) );
  AND U2522 ( .A(n2520), .B(n2521), .Z(n2359) );
  NANDN U2523 ( .A(n2522), .B(n2523), .Z(n2521) );
  NANDN U2524 ( .A(n2524), .B(n2525), .Z(n2523) );
  NANDN U2525 ( .A(n2525), .B(n2524), .Z(n2520) );
  ANDN U2526 ( .B(B[62]), .A(n68), .Z(n2361) );
  XNOR U2527 ( .A(n2369), .B(n2526), .Z(n2362) );
  XNOR U2528 ( .A(n2368), .B(n2366), .Z(n2526) );
  AND U2529 ( .A(n2527), .B(n2528), .Z(n2366) );
  NANDN U2530 ( .A(n2529), .B(n2530), .Z(n2528) );
  OR U2531 ( .A(n2531), .B(n2532), .Z(n2530) );
  NAND U2532 ( .A(n2532), .B(n2531), .Z(n2527) );
  ANDN U2533 ( .B(B[63]), .A(n69), .Z(n2368) );
  XNOR U2534 ( .A(n2376), .B(n2533), .Z(n2369) );
  XNOR U2535 ( .A(n2375), .B(n2373), .Z(n2533) );
  AND U2536 ( .A(n2534), .B(n2535), .Z(n2373) );
  NANDN U2537 ( .A(n2536), .B(n2537), .Z(n2535) );
  NANDN U2538 ( .A(n2538), .B(n2539), .Z(n2537) );
  NANDN U2539 ( .A(n2539), .B(n2538), .Z(n2534) );
  ANDN U2540 ( .B(B[64]), .A(n70), .Z(n2375) );
  XNOR U2541 ( .A(n2383), .B(n2540), .Z(n2376) );
  XNOR U2542 ( .A(n2382), .B(n2380), .Z(n2540) );
  AND U2543 ( .A(n2541), .B(n2542), .Z(n2380) );
  NANDN U2544 ( .A(n2543), .B(n2544), .Z(n2542) );
  OR U2545 ( .A(n2545), .B(n2546), .Z(n2544) );
  NAND U2546 ( .A(n2546), .B(n2545), .Z(n2541) );
  ANDN U2547 ( .B(B[65]), .A(n71), .Z(n2382) );
  XNOR U2548 ( .A(n2390), .B(n2547), .Z(n2383) );
  XNOR U2549 ( .A(n2389), .B(n2387), .Z(n2547) );
  AND U2550 ( .A(n2548), .B(n2549), .Z(n2387) );
  NANDN U2551 ( .A(n2550), .B(n2551), .Z(n2549) );
  NANDN U2552 ( .A(n2552), .B(n2553), .Z(n2551) );
  NANDN U2553 ( .A(n2553), .B(n2552), .Z(n2548) );
  ANDN U2554 ( .B(B[66]), .A(n72), .Z(n2389) );
  XNOR U2555 ( .A(n2397), .B(n2554), .Z(n2390) );
  XNOR U2556 ( .A(n2396), .B(n2394), .Z(n2554) );
  AND U2557 ( .A(n2555), .B(n2556), .Z(n2394) );
  NANDN U2558 ( .A(n2557), .B(n2558), .Z(n2556) );
  OR U2559 ( .A(n2559), .B(n2560), .Z(n2558) );
  NAND U2560 ( .A(n2560), .B(n2559), .Z(n2555) );
  ANDN U2561 ( .B(B[67]), .A(n73), .Z(n2396) );
  XNOR U2562 ( .A(n2404), .B(n2561), .Z(n2397) );
  XNOR U2563 ( .A(n2403), .B(n2401), .Z(n2561) );
  AND U2564 ( .A(n2562), .B(n2563), .Z(n2401) );
  NANDN U2565 ( .A(n2564), .B(n2565), .Z(n2563) );
  NANDN U2566 ( .A(n2566), .B(n2567), .Z(n2565) );
  NANDN U2567 ( .A(n2567), .B(n2566), .Z(n2562) );
  ANDN U2568 ( .B(B[68]), .A(n74), .Z(n2403) );
  XOR U2569 ( .A(n2409), .B(n2568), .Z(n2404) );
  XNOR U2570 ( .A(n2410), .B(n2411), .Z(n2568) );
  AND U2571 ( .A(n2569), .B(n2570), .Z(n2411) );
  NANDN U2572 ( .A(n2571), .B(n2572), .Z(n2570) );
  NANDN U2573 ( .A(n2573), .B(n2574), .Z(n2572) );
  ANDN U2574 ( .B(B[69]), .A(n75), .Z(n2410) );
  XOR U2575 ( .A(n2575), .B(n2576), .Z(n2409) );
  XNOR U2576 ( .A(n2577), .B(n40), .Z(n2576) );
  NAND U2577 ( .A(n2578), .B(n2579), .Z(n129) );
  NANDN U2578 ( .A(n2580), .B(n2581), .Z(n2579) );
  OR U2579 ( .A(n2582), .B(n2583), .Z(n2581) );
  NAND U2580 ( .A(n2583), .B(n2582), .Z(n2578) );
  XOR U2581 ( .A(n131), .B(n130), .Z(\A1[76] ) );
  XOR U2582 ( .A(n2583), .B(n2584), .Z(n130) );
  XNOR U2583 ( .A(n2582), .B(n2580), .Z(n2584) );
  AND U2584 ( .A(n2585), .B(n2586), .Z(n2580) );
  NANDN U2585 ( .A(n2587), .B(n2588), .Z(n2586) );
  NANDN U2586 ( .A(n2589), .B(n2590), .Z(n2588) );
  NANDN U2587 ( .A(n2590), .B(n2589), .Z(n2585) );
  ANDN U2588 ( .B(B[47]), .A(n54), .Z(n2582) );
  XNOR U2589 ( .A(n2427), .B(n2591), .Z(n2583) );
  XNOR U2590 ( .A(n2426), .B(n2424), .Z(n2591) );
  AND U2591 ( .A(n2592), .B(n2593), .Z(n2424) );
  NANDN U2592 ( .A(n2594), .B(n2595), .Z(n2593) );
  OR U2593 ( .A(n2596), .B(n2597), .Z(n2595) );
  NAND U2594 ( .A(n2597), .B(n2596), .Z(n2592) );
  ANDN U2595 ( .B(B[48]), .A(n55), .Z(n2426) );
  XNOR U2596 ( .A(n2434), .B(n2598), .Z(n2427) );
  XNOR U2597 ( .A(n2433), .B(n2431), .Z(n2598) );
  AND U2598 ( .A(n2599), .B(n2600), .Z(n2431) );
  NANDN U2599 ( .A(n2601), .B(n2602), .Z(n2600) );
  NANDN U2600 ( .A(n2603), .B(n2604), .Z(n2602) );
  NANDN U2601 ( .A(n2604), .B(n2603), .Z(n2599) );
  ANDN U2602 ( .B(B[49]), .A(n56), .Z(n2433) );
  XNOR U2603 ( .A(n2441), .B(n2605), .Z(n2434) );
  XNOR U2604 ( .A(n2440), .B(n2438), .Z(n2605) );
  AND U2605 ( .A(n2606), .B(n2607), .Z(n2438) );
  NANDN U2606 ( .A(n2608), .B(n2609), .Z(n2607) );
  OR U2607 ( .A(n2610), .B(n2611), .Z(n2609) );
  NAND U2608 ( .A(n2611), .B(n2610), .Z(n2606) );
  ANDN U2609 ( .B(B[50]), .A(n57), .Z(n2440) );
  XNOR U2610 ( .A(n2448), .B(n2612), .Z(n2441) );
  XNOR U2611 ( .A(n2447), .B(n2445), .Z(n2612) );
  AND U2612 ( .A(n2613), .B(n2614), .Z(n2445) );
  NANDN U2613 ( .A(n2615), .B(n2616), .Z(n2614) );
  NANDN U2614 ( .A(n2617), .B(n2618), .Z(n2616) );
  NANDN U2615 ( .A(n2618), .B(n2617), .Z(n2613) );
  ANDN U2616 ( .B(B[51]), .A(n58), .Z(n2447) );
  XNOR U2617 ( .A(n2455), .B(n2619), .Z(n2448) );
  XNOR U2618 ( .A(n2454), .B(n2452), .Z(n2619) );
  AND U2619 ( .A(n2620), .B(n2621), .Z(n2452) );
  NANDN U2620 ( .A(n2622), .B(n2623), .Z(n2621) );
  OR U2621 ( .A(n2624), .B(n2625), .Z(n2623) );
  NAND U2622 ( .A(n2625), .B(n2624), .Z(n2620) );
  ANDN U2623 ( .B(B[52]), .A(n59), .Z(n2454) );
  XNOR U2624 ( .A(n2462), .B(n2626), .Z(n2455) );
  XNOR U2625 ( .A(n2461), .B(n2459), .Z(n2626) );
  AND U2626 ( .A(n2627), .B(n2628), .Z(n2459) );
  NANDN U2627 ( .A(n2629), .B(n2630), .Z(n2628) );
  NANDN U2628 ( .A(n2631), .B(n2632), .Z(n2630) );
  NANDN U2629 ( .A(n2632), .B(n2631), .Z(n2627) );
  ANDN U2630 ( .B(B[53]), .A(n60), .Z(n2461) );
  XNOR U2631 ( .A(n2469), .B(n2633), .Z(n2462) );
  XNOR U2632 ( .A(n2468), .B(n2466), .Z(n2633) );
  AND U2633 ( .A(n2634), .B(n2635), .Z(n2466) );
  NANDN U2634 ( .A(n2636), .B(n2637), .Z(n2635) );
  OR U2635 ( .A(n2638), .B(n2639), .Z(n2637) );
  NAND U2636 ( .A(n2639), .B(n2638), .Z(n2634) );
  ANDN U2637 ( .B(B[54]), .A(n61), .Z(n2468) );
  XNOR U2638 ( .A(n2476), .B(n2640), .Z(n2469) );
  XNOR U2639 ( .A(n2475), .B(n2473), .Z(n2640) );
  AND U2640 ( .A(n2641), .B(n2642), .Z(n2473) );
  NANDN U2641 ( .A(n2643), .B(n2644), .Z(n2642) );
  NANDN U2642 ( .A(n2645), .B(n2646), .Z(n2644) );
  NANDN U2643 ( .A(n2646), .B(n2645), .Z(n2641) );
  ANDN U2644 ( .B(B[55]), .A(n62), .Z(n2475) );
  XNOR U2645 ( .A(n2483), .B(n2647), .Z(n2476) );
  XNOR U2646 ( .A(n2482), .B(n2480), .Z(n2647) );
  AND U2647 ( .A(n2648), .B(n2649), .Z(n2480) );
  NANDN U2648 ( .A(n2650), .B(n2651), .Z(n2649) );
  OR U2649 ( .A(n2652), .B(n2653), .Z(n2651) );
  NAND U2650 ( .A(n2653), .B(n2652), .Z(n2648) );
  ANDN U2651 ( .B(B[56]), .A(n63), .Z(n2482) );
  XNOR U2652 ( .A(n2490), .B(n2654), .Z(n2483) );
  XNOR U2653 ( .A(n2489), .B(n2487), .Z(n2654) );
  AND U2654 ( .A(n2655), .B(n2656), .Z(n2487) );
  NANDN U2655 ( .A(n2657), .B(n2658), .Z(n2656) );
  NANDN U2656 ( .A(n2659), .B(n2660), .Z(n2658) );
  NANDN U2657 ( .A(n2660), .B(n2659), .Z(n2655) );
  ANDN U2658 ( .B(B[57]), .A(n64), .Z(n2489) );
  XNOR U2659 ( .A(n2497), .B(n2661), .Z(n2490) );
  XNOR U2660 ( .A(n2496), .B(n2494), .Z(n2661) );
  AND U2661 ( .A(n2662), .B(n2663), .Z(n2494) );
  NANDN U2662 ( .A(n2664), .B(n2665), .Z(n2663) );
  OR U2663 ( .A(n2666), .B(n2667), .Z(n2665) );
  NAND U2664 ( .A(n2667), .B(n2666), .Z(n2662) );
  ANDN U2665 ( .B(B[58]), .A(n65), .Z(n2496) );
  XNOR U2666 ( .A(n2504), .B(n2668), .Z(n2497) );
  XNOR U2667 ( .A(n2503), .B(n2501), .Z(n2668) );
  AND U2668 ( .A(n2669), .B(n2670), .Z(n2501) );
  NANDN U2669 ( .A(n2671), .B(n2672), .Z(n2670) );
  NANDN U2670 ( .A(n2673), .B(n2674), .Z(n2672) );
  NANDN U2671 ( .A(n2674), .B(n2673), .Z(n2669) );
  ANDN U2672 ( .B(B[59]), .A(n66), .Z(n2503) );
  XNOR U2673 ( .A(n2511), .B(n2675), .Z(n2504) );
  XNOR U2674 ( .A(n2510), .B(n2508), .Z(n2675) );
  AND U2675 ( .A(n2676), .B(n2677), .Z(n2508) );
  NANDN U2676 ( .A(n2678), .B(n2679), .Z(n2677) );
  OR U2677 ( .A(n2680), .B(n2681), .Z(n2679) );
  NAND U2678 ( .A(n2681), .B(n2680), .Z(n2676) );
  ANDN U2679 ( .B(B[60]), .A(n67), .Z(n2510) );
  XNOR U2680 ( .A(n2518), .B(n2682), .Z(n2511) );
  XNOR U2681 ( .A(n2517), .B(n2515), .Z(n2682) );
  AND U2682 ( .A(n2683), .B(n2684), .Z(n2515) );
  NANDN U2683 ( .A(n2685), .B(n2686), .Z(n2684) );
  NANDN U2684 ( .A(n2687), .B(n2688), .Z(n2686) );
  NANDN U2685 ( .A(n2688), .B(n2687), .Z(n2683) );
  ANDN U2686 ( .B(B[61]), .A(n68), .Z(n2517) );
  XNOR U2687 ( .A(n2525), .B(n2689), .Z(n2518) );
  XNOR U2688 ( .A(n2524), .B(n2522), .Z(n2689) );
  AND U2689 ( .A(n2690), .B(n2691), .Z(n2522) );
  NANDN U2690 ( .A(n2692), .B(n2693), .Z(n2691) );
  OR U2691 ( .A(n2694), .B(n2695), .Z(n2693) );
  NAND U2692 ( .A(n2695), .B(n2694), .Z(n2690) );
  ANDN U2693 ( .B(B[62]), .A(n69), .Z(n2524) );
  XNOR U2694 ( .A(n2532), .B(n2696), .Z(n2525) );
  XNOR U2695 ( .A(n2531), .B(n2529), .Z(n2696) );
  AND U2696 ( .A(n2697), .B(n2698), .Z(n2529) );
  NANDN U2697 ( .A(n2699), .B(n2700), .Z(n2698) );
  NANDN U2698 ( .A(n2701), .B(n2702), .Z(n2700) );
  NANDN U2699 ( .A(n2702), .B(n2701), .Z(n2697) );
  ANDN U2700 ( .B(B[63]), .A(n70), .Z(n2531) );
  XNOR U2701 ( .A(n2539), .B(n2703), .Z(n2532) );
  XNOR U2702 ( .A(n2538), .B(n2536), .Z(n2703) );
  AND U2703 ( .A(n2704), .B(n2705), .Z(n2536) );
  NANDN U2704 ( .A(n2706), .B(n2707), .Z(n2705) );
  OR U2705 ( .A(n2708), .B(n2709), .Z(n2707) );
  NAND U2706 ( .A(n2709), .B(n2708), .Z(n2704) );
  ANDN U2707 ( .B(B[64]), .A(n71), .Z(n2538) );
  XNOR U2708 ( .A(n2546), .B(n2710), .Z(n2539) );
  XNOR U2709 ( .A(n2545), .B(n2543), .Z(n2710) );
  AND U2710 ( .A(n2711), .B(n2712), .Z(n2543) );
  NANDN U2711 ( .A(n2713), .B(n2714), .Z(n2712) );
  NANDN U2712 ( .A(n2715), .B(n2716), .Z(n2714) );
  NANDN U2713 ( .A(n2716), .B(n2715), .Z(n2711) );
  ANDN U2714 ( .B(B[65]), .A(n72), .Z(n2545) );
  XNOR U2715 ( .A(n2553), .B(n2717), .Z(n2546) );
  XNOR U2716 ( .A(n2552), .B(n2550), .Z(n2717) );
  AND U2717 ( .A(n2718), .B(n2719), .Z(n2550) );
  NANDN U2718 ( .A(n2720), .B(n2721), .Z(n2719) );
  OR U2719 ( .A(n2722), .B(n2723), .Z(n2721) );
  NAND U2720 ( .A(n2723), .B(n2722), .Z(n2718) );
  ANDN U2721 ( .B(B[66]), .A(n73), .Z(n2552) );
  XNOR U2722 ( .A(n2560), .B(n2724), .Z(n2553) );
  XNOR U2723 ( .A(n2559), .B(n2557), .Z(n2724) );
  AND U2724 ( .A(n2725), .B(n2726), .Z(n2557) );
  NANDN U2725 ( .A(n2727), .B(n2728), .Z(n2726) );
  NANDN U2726 ( .A(n2729), .B(n2730), .Z(n2728) );
  NANDN U2727 ( .A(n2730), .B(n2729), .Z(n2725) );
  ANDN U2728 ( .B(B[67]), .A(n74), .Z(n2559) );
  XNOR U2729 ( .A(n2567), .B(n2731), .Z(n2560) );
  XNOR U2730 ( .A(n2566), .B(n2564), .Z(n2731) );
  AND U2731 ( .A(n2732), .B(n2733), .Z(n2564) );
  NANDN U2732 ( .A(n2734), .B(n2735), .Z(n2733) );
  OR U2733 ( .A(n2736), .B(n2737), .Z(n2735) );
  NAND U2734 ( .A(n2737), .B(n2736), .Z(n2732) );
  ANDN U2735 ( .B(B[68]), .A(n75), .Z(n2566) );
  XOR U2736 ( .A(n2571), .B(n2738), .Z(n2567) );
  XNOR U2737 ( .A(n2573), .B(n2574), .Z(n2738) );
  AND U2738 ( .A(n2739), .B(n2740), .Z(n2574) );
  NAND U2739 ( .A(n2741), .B(n2742), .Z(n2740) );
  NANDN U2740 ( .A(n2743), .B(n2744), .Z(n2741) );
  ANDN U2741 ( .B(B[69]), .A(n76), .Z(n2573) );
  XNOR U2742 ( .A(n2745), .B(n2746), .Z(n2571) );
  XNOR U2743 ( .A(n2747), .B(n41), .Z(n2746) );
  NAND U2744 ( .A(n2748), .B(n2749), .Z(n131) );
  NANDN U2745 ( .A(n2750), .B(n2751), .Z(n2749) );
  OR U2746 ( .A(n2752), .B(n2753), .Z(n2751) );
  NAND U2747 ( .A(n2753), .B(n2752), .Z(n2748) );
  XOR U2748 ( .A(n133), .B(n132), .Z(\A1[75] ) );
  XOR U2749 ( .A(n2753), .B(n2754), .Z(n132) );
  XNOR U2750 ( .A(n2752), .B(n2750), .Z(n2754) );
  AND U2751 ( .A(n2755), .B(n2756), .Z(n2750) );
  NANDN U2752 ( .A(n2757), .B(n2758), .Z(n2756) );
  NANDN U2753 ( .A(n2759), .B(n2760), .Z(n2758) );
  NANDN U2754 ( .A(n2760), .B(n2759), .Z(n2755) );
  ANDN U2755 ( .B(B[46]), .A(n54), .Z(n2752) );
  XNOR U2756 ( .A(n2590), .B(n2761), .Z(n2753) );
  XNOR U2757 ( .A(n2589), .B(n2587), .Z(n2761) );
  AND U2758 ( .A(n2762), .B(n2763), .Z(n2587) );
  NANDN U2759 ( .A(n2764), .B(n2765), .Z(n2763) );
  OR U2760 ( .A(n2766), .B(n2767), .Z(n2765) );
  NAND U2761 ( .A(n2767), .B(n2766), .Z(n2762) );
  ANDN U2762 ( .B(B[47]), .A(n55), .Z(n2589) );
  XNOR U2763 ( .A(n2597), .B(n2768), .Z(n2590) );
  XNOR U2764 ( .A(n2596), .B(n2594), .Z(n2768) );
  AND U2765 ( .A(n2769), .B(n2770), .Z(n2594) );
  NANDN U2766 ( .A(n2771), .B(n2772), .Z(n2770) );
  NANDN U2767 ( .A(n2773), .B(n2774), .Z(n2772) );
  NANDN U2768 ( .A(n2774), .B(n2773), .Z(n2769) );
  ANDN U2769 ( .B(B[48]), .A(n56), .Z(n2596) );
  XNOR U2770 ( .A(n2604), .B(n2775), .Z(n2597) );
  XNOR U2771 ( .A(n2603), .B(n2601), .Z(n2775) );
  AND U2772 ( .A(n2776), .B(n2777), .Z(n2601) );
  NANDN U2773 ( .A(n2778), .B(n2779), .Z(n2777) );
  OR U2774 ( .A(n2780), .B(n2781), .Z(n2779) );
  NAND U2775 ( .A(n2781), .B(n2780), .Z(n2776) );
  ANDN U2776 ( .B(B[49]), .A(n57), .Z(n2603) );
  XNOR U2777 ( .A(n2611), .B(n2782), .Z(n2604) );
  XNOR U2778 ( .A(n2610), .B(n2608), .Z(n2782) );
  AND U2779 ( .A(n2783), .B(n2784), .Z(n2608) );
  NANDN U2780 ( .A(n2785), .B(n2786), .Z(n2784) );
  NANDN U2781 ( .A(n2787), .B(n2788), .Z(n2786) );
  NANDN U2782 ( .A(n2788), .B(n2787), .Z(n2783) );
  ANDN U2783 ( .B(B[50]), .A(n58), .Z(n2610) );
  XNOR U2784 ( .A(n2618), .B(n2789), .Z(n2611) );
  XNOR U2785 ( .A(n2617), .B(n2615), .Z(n2789) );
  AND U2786 ( .A(n2790), .B(n2791), .Z(n2615) );
  NANDN U2787 ( .A(n2792), .B(n2793), .Z(n2791) );
  OR U2788 ( .A(n2794), .B(n2795), .Z(n2793) );
  NAND U2789 ( .A(n2795), .B(n2794), .Z(n2790) );
  ANDN U2790 ( .B(B[51]), .A(n59), .Z(n2617) );
  XNOR U2791 ( .A(n2625), .B(n2796), .Z(n2618) );
  XNOR U2792 ( .A(n2624), .B(n2622), .Z(n2796) );
  AND U2793 ( .A(n2797), .B(n2798), .Z(n2622) );
  NANDN U2794 ( .A(n2799), .B(n2800), .Z(n2798) );
  NANDN U2795 ( .A(n2801), .B(n2802), .Z(n2800) );
  NANDN U2796 ( .A(n2802), .B(n2801), .Z(n2797) );
  ANDN U2797 ( .B(B[52]), .A(n60), .Z(n2624) );
  XNOR U2798 ( .A(n2632), .B(n2803), .Z(n2625) );
  XNOR U2799 ( .A(n2631), .B(n2629), .Z(n2803) );
  AND U2800 ( .A(n2804), .B(n2805), .Z(n2629) );
  NANDN U2801 ( .A(n2806), .B(n2807), .Z(n2805) );
  OR U2802 ( .A(n2808), .B(n2809), .Z(n2807) );
  NAND U2803 ( .A(n2809), .B(n2808), .Z(n2804) );
  ANDN U2804 ( .B(B[53]), .A(n61), .Z(n2631) );
  XNOR U2805 ( .A(n2639), .B(n2810), .Z(n2632) );
  XNOR U2806 ( .A(n2638), .B(n2636), .Z(n2810) );
  AND U2807 ( .A(n2811), .B(n2812), .Z(n2636) );
  NANDN U2808 ( .A(n2813), .B(n2814), .Z(n2812) );
  NANDN U2809 ( .A(n2815), .B(n2816), .Z(n2814) );
  NANDN U2810 ( .A(n2816), .B(n2815), .Z(n2811) );
  ANDN U2811 ( .B(B[54]), .A(n62), .Z(n2638) );
  XNOR U2812 ( .A(n2646), .B(n2817), .Z(n2639) );
  XNOR U2813 ( .A(n2645), .B(n2643), .Z(n2817) );
  AND U2814 ( .A(n2818), .B(n2819), .Z(n2643) );
  NANDN U2815 ( .A(n2820), .B(n2821), .Z(n2819) );
  OR U2816 ( .A(n2822), .B(n2823), .Z(n2821) );
  NAND U2817 ( .A(n2823), .B(n2822), .Z(n2818) );
  ANDN U2818 ( .B(B[55]), .A(n63), .Z(n2645) );
  XNOR U2819 ( .A(n2653), .B(n2824), .Z(n2646) );
  XNOR U2820 ( .A(n2652), .B(n2650), .Z(n2824) );
  AND U2821 ( .A(n2825), .B(n2826), .Z(n2650) );
  NANDN U2822 ( .A(n2827), .B(n2828), .Z(n2826) );
  NANDN U2823 ( .A(n2829), .B(n2830), .Z(n2828) );
  NANDN U2824 ( .A(n2830), .B(n2829), .Z(n2825) );
  ANDN U2825 ( .B(B[56]), .A(n64), .Z(n2652) );
  XNOR U2826 ( .A(n2660), .B(n2831), .Z(n2653) );
  XNOR U2827 ( .A(n2659), .B(n2657), .Z(n2831) );
  AND U2828 ( .A(n2832), .B(n2833), .Z(n2657) );
  NANDN U2829 ( .A(n2834), .B(n2835), .Z(n2833) );
  OR U2830 ( .A(n2836), .B(n2837), .Z(n2835) );
  NAND U2831 ( .A(n2837), .B(n2836), .Z(n2832) );
  ANDN U2832 ( .B(B[57]), .A(n65), .Z(n2659) );
  XNOR U2833 ( .A(n2667), .B(n2838), .Z(n2660) );
  XNOR U2834 ( .A(n2666), .B(n2664), .Z(n2838) );
  AND U2835 ( .A(n2839), .B(n2840), .Z(n2664) );
  NANDN U2836 ( .A(n2841), .B(n2842), .Z(n2840) );
  NANDN U2837 ( .A(n2843), .B(n2844), .Z(n2842) );
  NANDN U2838 ( .A(n2844), .B(n2843), .Z(n2839) );
  ANDN U2839 ( .B(B[58]), .A(n66), .Z(n2666) );
  XNOR U2840 ( .A(n2674), .B(n2845), .Z(n2667) );
  XNOR U2841 ( .A(n2673), .B(n2671), .Z(n2845) );
  AND U2842 ( .A(n2846), .B(n2847), .Z(n2671) );
  NANDN U2843 ( .A(n2848), .B(n2849), .Z(n2847) );
  OR U2844 ( .A(n2850), .B(n2851), .Z(n2849) );
  NAND U2845 ( .A(n2851), .B(n2850), .Z(n2846) );
  ANDN U2846 ( .B(B[59]), .A(n67), .Z(n2673) );
  XNOR U2847 ( .A(n2681), .B(n2852), .Z(n2674) );
  XNOR U2848 ( .A(n2680), .B(n2678), .Z(n2852) );
  AND U2849 ( .A(n2853), .B(n2854), .Z(n2678) );
  NANDN U2850 ( .A(n2855), .B(n2856), .Z(n2854) );
  NANDN U2851 ( .A(n2857), .B(n2858), .Z(n2856) );
  NANDN U2852 ( .A(n2858), .B(n2857), .Z(n2853) );
  ANDN U2853 ( .B(B[60]), .A(n68), .Z(n2680) );
  XNOR U2854 ( .A(n2688), .B(n2859), .Z(n2681) );
  XNOR U2855 ( .A(n2687), .B(n2685), .Z(n2859) );
  AND U2856 ( .A(n2860), .B(n2861), .Z(n2685) );
  NANDN U2857 ( .A(n2862), .B(n2863), .Z(n2861) );
  OR U2858 ( .A(n2864), .B(n2865), .Z(n2863) );
  NAND U2859 ( .A(n2865), .B(n2864), .Z(n2860) );
  ANDN U2860 ( .B(B[61]), .A(n69), .Z(n2687) );
  XNOR U2861 ( .A(n2695), .B(n2866), .Z(n2688) );
  XNOR U2862 ( .A(n2694), .B(n2692), .Z(n2866) );
  AND U2863 ( .A(n2867), .B(n2868), .Z(n2692) );
  NANDN U2864 ( .A(n2869), .B(n2870), .Z(n2868) );
  NANDN U2865 ( .A(n2871), .B(n2872), .Z(n2870) );
  NANDN U2866 ( .A(n2872), .B(n2871), .Z(n2867) );
  ANDN U2867 ( .B(B[62]), .A(n70), .Z(n2694) );
  XNOR U2868 ( .A(n2702), .B(n2873), .Z(n2695) );
  XNOR U2869 ( .A(n2701), .B(n2699), .Z(n2873) );
  AND U2870 ( .A(n2874), .B(n2875), .Z(n2699) );
  NANDN U2871 ( .A(n2876), .B(n2877), .Z(n2875) );
  OR U2872 ( .A(n2878), .B(n2879), .Z(n2877) );
  NAND U2873 ( .A(n2879), .B(n2878), .Z(n2874) );
  ANDN U2874 ( .B(B[63]), .A(n71), .Z(n2701) );
  XNOR U2875 ( .A(n2709), .B(n2880), .Z(n2702) );
  XNOR U2876 ( .A(n2708), .B(n2706), .Z(n2880) );
  AND U2877 ( .A(n2881), .B(n2882), .Z(n2706) );
  NANDN U2878 ( .A(n2883), .B(n2884), .Z(n2882) );
  NANDN U2879 ( .A(n2885), .B(n2886), .Z(n2884) );
  NANDN U2880 ( .A(n2886), .B(n2885), .Z(n2881) );
  ANDN U2881 ( .B(B[64]), .A(n72), .Z(n2708) );
  XNOR U2882 ( .A(n2716), .B(n2887), .Z(n2709) );
  XNOR U2883 ( .A(n2715), .B(n2713), .Z(n2887) );
  AND U2884 ( .A(n2888), .B(n2889), .Z(n2713) );
  NANDN U2885 ( .A(n2890), .B(n2891), .Z(n2889) );
  OR U2886 ( .A(n2892), .B(n2893), .Z(n2891) );
  NAND U2887 ( .A(n2893), .B(n2892), .Z(n2888) );
  ANDN U2888 ( .B(B[65]), .A(n73), .Z(n2715) );
  XNOR U2889 ( .A(n2723), .B(n2894), .Z(n2716) );
  XNOR U2890 ( .A(n2722), .B(n2720), .Z(n2894) );
  AND U2891 ( .A(n2895), .B(n2896), .Z(n2720) );
  NANDN U2892 ( .A(n2897), .B(n2898), .Z(n2896) );
  NANDN U2893 ( .A(n2899), .B(n2900), .Z(n2898) );
  NANDN U2894 ( .A(n2900), .B(n2899), .Z(n2895) );
  ANDN U2895 ( .B(B[66]), .A(n74), .Z(n2722) );
  XNOR U2896 ( .A(n2730), .B(n2901), .Z(n2723) );
  XNOR U2897 ( .A(n2729), .B(n2727), .Z(n2901) );
  AND U2898 ( .A(n2902), .B(n2903), .Z(n2727) );
  NANDN U2899 ( .A(n2904), .B(n2905), .Z(n2903) );
  OR U2900 ( .A(n2906), .B(n2907), .Z(n2905) );
  NAND U2901 ( .A(n2907), .B(n2906), .Z(n2902) );
  ANDN U2902 ( .B(B[67]), .A(n75), .Z(n2729) );
  XNOR U2903 ( .A(n2737), .B(n2908), .Z(n2730) );
  XNOR U2904 ( .A(n2736), .B(n2734), .Z(n2908) );
  AND U2905 ( .A(n2909), .B(n2910), .Z(n2734) );
  NANDN U2906 ( .A(n2911), .B(n2912), .Z(n2910) );
  NANDN U2907 ( .A(n2913), .B(n2914), .Z(n2912) );
  NANDN U2908 ( .A(n2914), .B(n2913), .Z(n2909) );
  ANDN U2909 ( .B(B[68]), .A(n76), .Z(n2736) );
  XOR U2910 ( .A(n2742), .B(n2915), .Z(n2737) );
  XNOR U2911 ( .A(n2743), .B(n2744), .Z(n2915) );
  AND U2912 ( .A(n2916), .B(n2917), .Z(n2744) );
  NANDN U2913 ( .A(n2918), .B(n2919), .Z(n2917) );
  NANDN U2914 ( .A(n2920), .B(n2921), .Z(n2919) );
  ANDN U2915 ( .B(B[69]), .A(n77), .Z(n2743) );
  XOR U2916 ( .A(n2922), .B(n2923), .Z(n2742) );
  XNOR U2917 ( .A(n2924), .B(n42), .Z(n2923) );
  NAND U2918 ( .A(n2925), .B(n2926), .Z(n133) );
  NANDN U2919 ( .A(n2927), .B(n2928), .Z(n2926) );
  OR U2920 ( .A(n2929), .B(n2930), .Z(n2928) );
  NAND U2921 ( .A(n2930), .B(n2929), .Z(n2925) );
  XOR U2922 ( .A(n135), .B(n134), .Z(\A1[74] ) );
  XOR U2923 ( .A(n2930), .B(n2931), .Z(n134) );
  XNOR U2924 ( .A(n2929), .B(n2927), .Z(n2931) );
  AND U2925 ( .A(n2932), .B(n2933), .Z(n2927) );
  NANDN U2926 ( .A(n2934), .B(n2935), .Z(n2933) );
  NANDN U2927 ( .A(n2936), .B(n2937), .Z(n2935) );
  NANDN U2928 ( .A(n2937), .B(n2936), .Z(n2932) );
  ANDN U2929 ( .B(B[45]), .A(n54), .Z(n2929) );
  XNOR U2930 ( .A(n2760), .B(n2938), .Z(n2930) );
  XNOR U2931 ( .A(n2759), .B(n2757), .Z(n2938) );
  AND U2932 ( .A(n2939), .B(n2940), .Z(n2757) );
  NANDN U2933 ( .A(n2941), .B(n2942), .Z(n2940) );
  OR U2934 ( .A(n2943), .B(n2944), .Z(n2942) );
  NAND U2935 ( .A(n2944), .B(n2943), .Z(n2939) );
  ANDN U2936 ( .B(B[46]), .A(n55), .Z(n2759) );
  XNOR U2937 ( .A(n2767), .B(n2945), .Z(n2760) );
  XNOR U2938 ( .A(n2766), .B(n2764), .Z(n2945) );
  AND U2939 ( .A(n2946), .B(n2947), .Z(n2764) );
  NANDN U2940 ( .A(n2948), .B(n2949), .Z(n2947) );
  NANDN U2941 ( .A(n2950), .B(n2951), .Z(n2949) );
  NANDN U2942 ( .A(n2951), .B(n2950), .Z(n2946) );
  ANDN U2943 ( .B(B[47]), .A(n56), .Z(n2766) );
  XNOR U2944 ( .A(n2774), .B(n2952), .Z(n2767) );
  XNOR U2945 ( .A(n2773), .B(n2771), .Z(n2952) );
  AND U2946 ( .A(n2953), .B(n2954), .Z(n2771) );
  NANDN U2947 ( .A(n2955), .B(n2956), .Z(n2954) );
  OR U2948 ( .A(n2957), .B(n2958), .Z(n2956) );
  NAND U2949 ( .A(n2958), .B(n2957), .Z(n2953) );
  ANDN U2950 ( .B(B[48]), .A(n57), .Z(n2773) );
  XNOR U2951 ( .A(n2781), .B(n2959), .Z(n2774) );
  XNOR U2952 ( .A(n2780), .B(n2778), .Z(n2959) );
  AND U2953 ( .A(n2960), .B(n2961), .Z(n2778) );
  NANDN U2954 ( .A(n2962), .B(n2963), .Z(n2961) );
  NANDN U2955 ( .A(n2964), .B(n2965), .Z(n2963) );
  NANDN U2956 ( .A(n2965), .B(n2964), .Z(n2960) );
  ANDN U2957 ( .B(B[49]), .A(n58), .Z(n2780) );
  XNOR U2958 ( .A(n2788), .B(n2966), .Z(n2781) );
  XNOR U2959 ( .A(n2787), .B(n2785), .Z(n2966) );
  AND U2960 ( .A(n2967), .B(n2968), .Z(n2785) );
  NANDN U2961 ( .A(n2969), .B(n2970), .Z(n2968) );
  OR U2962 ( .A(n2971), .B(n2972), .Z(n2970) );
  NAND U2963 ( .A(n2972), .B(n2971), .Z(n2967) );
  ANDN U2964 ( .B(B[50]), .A(n59), .Z(n2787) );
  XNOR U2965 ( .A(n2795), .B(n2973), .Z(n2788) );
  XNOR U2966 ( .A(n2794), .B(n2792), .Z(n2973) );
  AND U2967 ( .A(n2974), .B(n2975), .Z(n2792) );
  NANDN U2968 ( .A(n2976), .B(n2977), .Z(n2975) );
  NANDN U2969 ( .A(n2978), .B(n2979), .Z(n2977) );
  NANDN U2970 ( .A(n2979), .B(n2978), .Z(n2974) );
  ANDN U2971 ( .B(B[51]), .A(n60), .Z(n2794) );
  XNOR U2972 ( .A(n2802), .B(n2980), .Z(n2795) );
  XNOR U2973 ( .A(n2801), .B(n2799), .Z(n2980) );
  AND U2974 ( .A(n2981), .B(n2982), .Z(n2799) );
  NANDN U2975 ( .A(n2983), .B(n2984), .Z(n2982) );
  OR U2976 ( .A(n2985), .B(n2986), .Z(n2984) );
  NAND U2977 ( .A(n2986), .B(n2985), .Z(n2981) );
  ANDN U2978 ( .B(B[52]), .A(n61), .Z(n2801) );
  XNOR U2979 ( .A(n2809), .B(n2987), .Z(n2802) );
  XNOR U2980 ( .A(n2808), .B(n2806), .Z(n2987) );
  AND U2981 ( .A(n2988), .B(n2989), .Z(n2806) );
  NANDN U2982 ( .A(n2990), .B(n2991), .Z(n2989) );
  NANDN U2983 ( .A(n2992), .B(n2993), .Z(n2991) );
  NANDN U2984 ( .A(n2993), .B(n2992), .Z(n2988) );
  ANDN U2985 ( .B(B[53]), .A(n62), .Z(n2808) );
  XNOR U2986 ( .A(n2816), .B(n2994), .Z(n2809) );
  XNOR U2987 ( .A(n2815), .B(n2813), .Z(n2994) );
  AND U2988 ( .A(n2995), .B(n2996), .Z(n2813) );
  NANDN U2989 ( .A(n2997), .B(n2998), .Z(n2996) );
  OR U2990 ( .A(n2999), .B(n3000), .Z(n2998) );
  NAND U2991 ( .A(n3000), .B(n2999), .Z(n2995) );
  ANDN U2992 ( .B(B[54]), .A(n63), .Z(n2815) );
  XNOR U2993 ( .A(n2823), .B(n3001), .Z(n2816) );
  XNOR U2994 ( .A(n2822), .B(n2820), .Z(n3001) );
  AND U2995 ( .A(n3002), .B(n3003), .Z(n2820) );
  NANDN U2996 ( .A(n3004), .B(n3005), .Z(n3003) );
  NANDN U2997 ( .A(n3006), .B(n3007), .Z(n3005) );
  NANDN U2998 ( .A(n3007), .B(n3006), .Z(n3002) );
  ANDN U2999 ( .B(B[55]), .A(n64), .Z(n2822) );
  XNOR U3000 ( .A(n2830), .B(n3008), .Z(n2823) );
  XNOR U3001 ( .A(n2829), .B(n2827), .Z(n3008) );
  AND U3002 ( .A(n3009), .B(n3010), .Z(n2827) );
  NANDN U3003 ( .A(n3011), .B(n3012), .Z(n3010) );
  OR U3004 ( .A(n3013), .B(n3014), .Z(n3012) );
  NAND U3005 ( .A(n3014), .B(n3013), .Z(n3009) );
  ANDN U3006 ( .B(B[56]), .A(n65), .Z(n2829) );
  XNOR U3007 ( .A(n2837), .B(n3015), .Z(n2830) );
  XNOR U3008 ( .A(n2836), .B(n2834), .Z(n3015) );
  AND U3009 ( .A(n3016), .B(n3017), .Z(n2834) );
  NANDN U3010 ( .A(n3018), .B(n3019), .Z(n3017) );
  NANDN U3011 ( .A(n3020), .B(n3021), .Z(n3019) );
  NANDN U3012 ( .A(n3021), .B(n3020), .Z(n3016) );
  ANDN U3013 ( .B(B[57]), .A(n66), .Z(n2836) );
  XNOR U3014 ( .A(n2844), .B(n3022), .Z(n2837) );
  XNOR U3015 ( .A(n2843), .B(n2841), .Z(n3022) );
  AND U3016 ( .A(n3023), .B(n3024), .Z(n2841) );
  NANDN U3017 ( .A(n3025), .B(n3026), .Z(n3024) );
  OR U3018 ( .A(n3027), .B(n3028), .Z(n3026) );
  NAND U3019 ( .A(n3028), .B(n3027), .Z(n3023) );
  ANDN U3020 ( .B(B[58]), .A(n67), .Z(n2843) );
  XNOR U3021 ( .A(n2851), .B(n3029), .Z(n2844) );
  XNOR U3022 ( .A(n2850), .B(n2848), .Z(n3029) );
  AND U3023 ( .A(n3030), .B(n3031), .Z(n2848) );
  NANDN U3024 ( .A(n3032), .B(n3033), .Z(n3031) );
  NANDN U3025 ( .A(n3034), .B(n3035), .Z(n3033) );
  NANDN U3026 ( .A(n3035), .B(n3034), .Z(n3030) );
  ANDN U3027 ( .B(B[59]), .A(n68), .Z(n2850) );
  XNOR U3028 ( .A(n2858), .B(n3036), .Z(n2851) );
  XNOR U3029 ( .A(n2857), .B(n2855), .Z(n3036) );
  AND U3030 ( .A(n3037), .B(n3038), .Z(n2855) );
  NANDN U3031 ( .A(n3039), .B(n3040), .Z(n3038) );
  OR U3032 ( .A(n3041), .B(n3042), .Z(n3040) );
  NAND U3033 ( .A(n3042), .B(n3041), .Z(n3037) );
  ANDN U3034 ( .B(B[60]), .A(n69), .Z(n2857) );
  XNOR U3035 ( .A(n2865), .B(n3043), .Z(n2858) );
  XNOR U3036 ( .A(n2864), .B(n2862), .Z(n3043) );
  AND U3037 ( .A(n3044), .B(n3045), .Z(n2862) );
  NANDN U3038 ( .A(n3046), .B(n3047), .Z(n3045) );
  NANDN U3039 ( .A(n3048), .B(n3049), .Z(n3047) );
  NANDN U3040 ( .A(n3049), .B(n3048), .Z(n3044) );
  ANDN U3041 ( .B(B[61]), .A(n70), .Z(n2864) );
  XNOR U3042 ( .A(n2872), .B(n3050), .Z(n2865) );
  XNOR U3043 ( .A(n2871), .B(n2869), .Z(n3050) );
  AND U3044 ( .A(n3051), .B(n3052), .Z(n2869) );
  NANDN U3045 ( .A(n3053), .B(n3054), .Z(n3052) );
  OR U3046 ( .A(n3055), .B(n3056), .Z(n3054) );
  NAND U3047 ( .A(n3056), .B(n3055), .Z(n3051) );
  ANDN U3048 ( .B(B[62]), .A(n71), .Z(n2871) );
  XNOR U3049 ( .A(n2879), .B(n3057), .Z(n2872) );
  XNOR U3050 ( .A(n2878), .B(n2876), .Z(n3057) );
  AND U3051 ( .A(n3058), .B(n3059), .Z(n2876) );
  NANDN U3052 ( .A(n3060), .B(n3061), .Z(n3059) );
  NANDN U3053 ( .A(n3062), .B(n3063), .Z(n3061) );
  NANDN U3054 ( .A(n3063), .B(n3062), .Z(n3058) );
  ANDN U3055 ( .B(B[63]), .A(n72), .Z(n2878) );
  XNOR U3056 ( .A(n2886), .B(n3064), .Z(n2879) );
  XNOR U3057 ( .A(n2885), .B(n2883), .Z(n3064) );
  AND U3058 ( .A(n3065), .B(n3066), .Z(n2883) );
  NANDN U3059 ( .A(n3067), .B(n3068), .Z(n3066) );
  OR U3060 ( .A(n3069), .B(n3070), .Z(n3068) );
  NAND U3061 ( .A(n3070), .B(n3069), .Z(n3065) );
  ANDN U3062 ( .B(B[64]), .A(n73), .Z(n2885) );
  XNOR U3063 ( .A(n2893), .B(n3071), .Z(n2886) );
  XNOR U3064 ( .A(n2892), .B(n2890), .Z(n3071) );
  AND U3065 ( .A(n3072), .B(n3073), .Z(n2890) );
  NANDN U3066 ( .A(n3074), .B(n3075), .Z(n3073) );
  NANDN U3067 ( .A(n3076), .B(n3077), .Z(n3075) );
  NANDN U3068 ( .A(n3077), .B(n3076), .Z(n3072) );
  ANDN U3069 ( .B(B[65]), .A(n74), .Z(n2892) );
  XNOR U3070 ( .A(n2900), .B(n3078), .Z(n2893) );
  XNOR U3071 ( .A(n2899), .B(n2897), .Z(n3078) );
  AND U3072 ( .A(n3079), .B(n3080), .Z(n2897) );
  NANDN U3073 ( .A(n3081), .B(n3082), .Z(n3080) );
  OR U3074 ( .A(n3083), .B(n3084), .Z(n3082) );
  NAND U3075 ( .A(n3084), .B(n3083), .Z(n3079) );
  ANDN U3076 ( .B(B[66]), .A(n75), .Z(n2899) );
  XNOR U3077 ( .A(n2907), .B(n3085), .Z(n2900) );
  XNOR U3078 ( .A(n2906), .B(n2904), .Z(n3085) );
  AND U3079 ( .A(n3086), .B(n3087), .Z(n2904) );
  NANDN U3080 ( .A(n3088), .B(n3089), .Z(n3087) );
  NANDN U3081 ( .A(n3090), .B(n3091), .Z(n3089) );
  NANDN U3082 ( .A(n3091), .B(n3090), .Z(n3086) );
  ANDN U3083 ( .B(B[67]), .A(n76), .Z(n2906) );
  XNOR U3084 ( .A(n2914), .B(n3092), .Z(n2907) );
  XNOR U3085 ( .A(n2913), .B(n2911), .Z(n3092) );
  AND U3086 ( .A(n3093), .B(n3094), .Z(n2911) );
  NANDN U3087 ( .A(n3095), .B(n3096), .Z(n3094) );
  OR U3088 ( .A(n3097), .B(n3098), .Z(n3096) );
  NAND U3089 ( .A(n3098), .B(n3097), .Z(n3093) );
  ANDN U3090 ( .B(B[68]), .A(n77), .Z(n2913) );
  XOR U3091 ( .A(n2918), .B(n3099), .Z(n2914) );
  XNOR U3092 ( .A(n2920), .B(n2921), .Z(n3099) );
  AND U3093 ( .A(n3100), .B(n3101), .Z(n2921) );
  NAND U3094 ( .A(n3102), .B(n3103), .Z(n3101) );
  NANDN U3095 ( .A(n3104), .B(n3105), .Z(n3102) );
  ANDN U3096 ( .B(B[69]), .A(n78), .Z(n2920) );
  XNOR U3097 ( .A(n3106), .B(n3107), .Z(n2918) );
  XNOR U3098 ( .A(n3108), .B(n43), .Z(n3107) );
  NAND U3099 ( .A(n3109), .B(n3110), .Z(n135) );
  NANDN U3100 ( .A(n3111), .B(n3112), .Z(n3110) );
  OR U3101 ( .A(n3113), .B(n3114), .Z(n3112) );
  NAND U3102 ( .A(n3114), .B(n3113), .Z(n3109) );
  XOR U3103 ( .A(n137), .B(n136), .Z(\A1[73] ) );
  XOR U3104 ( .A(n3114), .B(n3115), .Z(n136) );
  XNOR U3105 ( .A(n3113), .B(n3111), .Z(n3115) );
  AND U3106 ( .A(n3116), .B(n3117), .Z(n3111) );
  NANDN U3107 ( .A(n3118), .B(n3119), .Z(n3117) );
  NANDN U3108 ( .A(n3120), .B(n3121), .Z(n3119) );
  NANDN U3109 ( .A(n3121), .B(n3120), .Z(n3116) );
  ANDN U3110 ( .B(B[44]), .A(n54), .Z(n3113) );
  XNOR U3111 ( .A(n2937), .B(n3122), .Z(n3114) );
  XNOR U3112 ( .A(n2936), .B(n2934), .Z(n3122) );
  AND U3113 ( .A(n3123), .B(n3124), .Z(n2934) );
  NANDN U3114 ( .A(n3125), .B(n3126), .Z(n3124) );
  OR U3115 ( .A(n3127), .B(n3128), .Z(n3126) );
  NAND U3116 ( .A(n3128), .B(n3127), .Z(n3123) );
  ANDN U3117 ( .B(B[45]), .A(n55), .Z(n2936) );
  XNOR U3118 ( .A(n2944), .B(n3129), .Z(n2937) );
  XNOR U3119 ( .A(n2943), .B(n2941), .Z(n3129) );
  AND U3120 ( .A(n3130), .B(n3131), .Z(n2941) );
  NANDN U3121 ( .A(n3132), .B(n3133), .Z(n3131) );
  NANDN U3122 ( .A(n3134), .B(n3135), .Z(n3133) );
  NANDN U3123 ( .A(n3135), .B(n3134), .Z(n3130) );
  ANDN U3124 ( .B(B[46]), .A(n56), .Z(n2943) );
  XNOR U3125 ( .A(n2951), .B(n3136), .Z(n2944) );
  XNOR U3126 ( .A(n2950), .B(n2948), .Z(n3136) );
  AND U3127 ( .A(n3137), .B(n3138), .Z(n2948) );
  NANDN U3128 ( .A(n3139), .B(n3140), .Z(n3138) );
  OR U3129 ( .A(n3141), .B(n3142), .Z(n3140) );
  NAND U3130 ( .A(n3142), .B(n3141), .Z(n3137) );
  ANDN U3131 ( .B(B[47]), .A(n57), .Z(n2950) );
  XNOR U3132 ( .A(n2958), .B(n3143), .Z(n2951) );
  XNOR U3133 ( .A(n2957), .B(n2955), .Z(n3143) );
  AND U3134 ( .A(n3144), .B(n3145), .Z(n2955) );
  NANDN U3135 ( .A(n3146), .B(n3147), .Z(n3145) );
  NANDN U3136 ( .A(n3148), .B(n3149), .Z(n3147) );
  NANDN U3137 ( .A(n3149), .B(n3148), .Z(n3144) );
  ANDN U3138 ( .B(B[48]), .A(n58), .Z(n2957) );
  XNOR U3139 ( .A(n2965), .B(n3150), .Z(n2958) );
  XNOR U3140 ( .A(n2964), .B(n2962), .Z(n3150) );
  AND U3141 ( .A(n3151), .B(n3152), .Z(n2962) );
  NANDN U3142 ( .A(n3153), .B(n3154), .Z(n3152) );
  OR U3143 ( .A(n3155), .B(n3156), .Z(n3154) );
  NAND U3144 ( .A(n3156), .B(n3155), .Z(n3151) );
  ANDN U3145 ( .B(B[49]), .A(n59), .Z(n2964) );
  XNOR U3146 ( .A(n2972), .B(n3157), .Z(n2965) );
  XNOR U3147 ( .A(n2971), .B(n2969), .Z(n3157) );
  AND U3148 ( .A(n3158), .B(n3159), .Z(n2969) );
  NANDN U3149 ( .A(n3160), .B(n3161), .Z(n3159) );
  NANDN U3150 ( .A(n3162), .B(n3163), .Z(n3161) );
  NANDN U3151 ( .A(n3163), .B(n3162), .Z(n3158) );
  ANDN U3152 ( .B(B[50]), .A(n60), .Z(n2971) );
  XNOR U3153 ( .A(n2979), .B(n3164), .Z(n2972) );
  XNOR U3154 ( .A(n2978), .B(n2976), .Z(n3164) );
  AND U3155 ( .A(n3165), .B(n3166), .Z(n2976) );
  NANDN U3156 ( .A(n3167), .B(n3168), .Z(n3166) );
  OR U3157 ( .A(n3169), .B(n3170), .Z(n3168) );
  NAND U3158 ( .A(n3170), .B(n3169), .Z(n3165) );
  ANDN U3159 ( .B(B[51]), .A(n61), .Z(n2978) );
  XNOR U3160 ( .A(n2986), .B(n3171), .Z(n2979) );
  XNOR U3161 ( .A(n2985), .B(n2983), .Z(n3171) );
  AND U3162 ( .A(n3172), .B(n3173), .Z(n2983) );
  NANDN U3163 ( .A(n3174), .B(n3175), .Z(n3173) );
  NANDN U3164 ( .A(n3176), .B(n3177), .Z(n3175) );
  NANDN U3165 ( .A(n3177), .B(n3176), .Z(n3172) );
  ANDN U3166 ( .B(B[52]), .A(n62), .Z(n2985) );
  XNOR U3167 ( .A(n2993), .B(n3178), .Z(n2986) );
  XNOR U3168 ( .A(n2992), .B(n2990), .Z(n3178) );
  AND U3169 ( .A(n3179), .B(n3180), .Z(n2990) );
  NANDN U3170 ( .A(n3181), .B(n3182), .Z(n3180) );
  OR U3171 ( .A(n3183), .B(n3184), .Z(n3182) );
  NAND U3172 ( .A(n3184), .B(n3183), .Z(n3179) );
  ANDN U3173 ( .B(B[53]), .A(n63), .Z(n2992) );
  XNOR U3174 ( .A(n3000), .B(n3185), .Z(n2993) );
  XNOR U3175 ( .A(n2999), .B(n2997), .Z(n3185) );
  AND U3176 ( .A(n3186), .B(n3187), .Z(n2997) );
  NANDN U3177 ( .A(n3188), .B(n3189), .Z(n3187) );
  NANDN U3178 ( .A(n3190), .B(n3191), .Z(n3189) );
  NANDN U3179 ( .A(n3191), .B(n3190), .Z(n3186) );
  ANDN U3180 ( .B(B[54]), .A(n64), .Z(n2999) );
  XNOR U3181 ( .A(n3007), .B(n3192), .Z(n3000) );
  XNOR U3182 ( .A(n3006), .B(n3004), .Z(n3192) );
  AND U3183 ( .A(n3193), .B(n3194), .Z(n3004) );
  NANDN U3184 ( .A(n3195), .B(n3196), .Z(n3194) );
  OR U3185 ( .A(n3197), .B(n3198), .Z(n3196) );
  NAND U3186 ( .A(n3198), .B(n3197), .Z(n3193) );
  ANDN U3187 ( .B(B[55]), .A(n65), .Z(n3006) );
  XNOR U3188 ( .A(n3014), .B(n3199), .Z(n3007) );
  XNOR U3189 ( .A(n3013), .B(n3011), .Z(n3199) );
  AND U3190 ( .A(n3200), .B(n3201), .Z(n3011) );
  NANDN U3191 ( .A(n3202), .B(n3203), .Z(n3201) );
  NANDN U3192 ( .A(n3204), .B(n3205), .Z(n3203) );
  NANDN U3193 ( .A(n3205), .B(n3204), .Z(n3200) );
  ANDN U3194 ( .B(B[56]), .A(n66), .Z(n3013) );
  XNOR U3195 ( .A(n3021), .B(n3206), .Z(n3014) );
  XNOR U3196 ( .A(n3020), .B(n3018), .Z(n3206) );
  AND U3197 ( .A(n3207), .B(n3208), .Z(n3018) );
  NANDN U3198 ( .A(n3209), .B(n3210), .Z(n3208) );
  OR U3199 ( .A(n3211), .B(n3212), .Z(n3210) );
  NAND U3200 ( .A(n3212), .B(n3211), .Z(n3207) );
  ANDN U3201 ( .B(B[57]), .A(n67), .Z(n3020) );
  XNOR U3202 ( .A(n3028), .B(n3213), .Z(n3021) );
  XNOR U3203 ( .A(n3027), .B(n3025), .Z(n3213) );
  AND U3204 ( .A(n3214), .B(n3215), .Z(n3025) );
  NANDN U3205 ( .A(n3216), .B(n3217), .Z(n3215) );
  NANDN U3206 ( .A(n3218), .B(n3219), .Z(n3217) );
  NANDN U3207 ( .A(n3219), .B(n3218), .Z(n3214) );
  ANDN U3208 ( .B(B[58]), .A(n68), .Z(n3027) );
  XNOR U3209 ( .A(n3035), .B(n3220), .Z(n3028) );
  XNOR U3210 ( .A(n3034), .B(n3032), .Z(n3220) );
  AND U3211 ( .A(n3221), .B(n3222), .Z(n3032) );
  NANDN U3212 ( .A(n3223), .B(n3224), .Z(n3222) );
  OR U3213 ( .A(n3225), .B(n3226), .Z(n3224) );
  NAND U3214 ( .A(n3226), .B(n3225), .Z(n3221) );
  ANDN U3215 ( .B(B[59]), .A(n69), .Z(n3034) );
  XNOR U3216 ( .A(n3042), .B(n3227), .Z(n3035) );
  XNOR U3217 ( .A(n3041), .B(n3039), .Z(n3227) );
  AND U3218 ( .A(n3228), .B(n3229), .Z(n3039) );
  NANDN U3219 ( .A(n3230), .B(n3231), .Z(n3229) );
  NANDN U3220 ( .A(n3232), .B(n3233), .Z(n3231) );
  NANDN U3221 ( .A(n3233), .B(n3232), .Z(n3228) );
  ANDN U3222 ( .B(B[60]), .A(n70), .Z(n3041) );
  XNOR U3223 ( .A(n3049), .B(n3234), .Z(n3042) );
  XNOR U3224 ( .A(n3048), .B(n3046), .Z(n3234) );
  AND U3225 ( .A(n3235), .B(n3236), .Z(n3046) );
  NANDN U3226 ( .A(n3237), .B(n3238), .Z(n3236) );
  OR U3227 ( .A(n3239), .B(n3240), .Z(n3238) );
  NAND U3228 ( .A(n3240), .B(n3239), .Z(n3235) );
  ANDN U3229 ( .B(B[61]), .A(n71), .Z(n3048) );
  XNOR U3230 ( .A(n3056), .B(n3241), .Z(n3049) );
  XNOR U3231 ( .A(n3055), .B(n3053), .Z(n3241) );
  AND U3232 ( .A(n3242), .B(n3243), .Z(n3053) );
  NANDN U3233 ( .A(n3244), .B(n3245), .Z(n3243) );
  NANDN U3234 ( .A(n3246), .B(n3247), .Z(n3245) );
  NANDN U3235 ( .A(n3247), .B(n3246), .Z(n3242) );
  ANDN U3236 ( .B(B[62]), .A(n72), .Z(n3055) );
  XNOR U3237 ( .A(n3063), .B(n3248), .Z(n3056) );
  XNOR U3238 ( .A(n3062), .B(n3060), .Z(n3248) );
  AND U3239 ( .A(n3249), .B(n3250), .Z(n3060) );
  NANDN U3240 ( .A(n3251), .B(n3252), .Z(n3250) );
  OR U3241 ( .A(n3253), .B(n3254), .Z(n3252) );
  NAND U3242 ( .A(n3254), .B(n3253), .Z(n3249) );
  ANDN U3243 ( .B(B[63]), .A(n73), .Z(n3062) );
  XNOR U3244 ( .A(n3070), .B(n3255), .Z(n3063) );
  XNOR U3245 ( .A(n3069), .B(n3067), .Z(n3255) );
  AND U3246 ( .A(n3256), .B(n3257), .Z(n3067) );
  NANDN U3247 ( .A(n3258), .B(n3259), .Z(n3257) );
  NANDN U3248 ( .A(n3260), .B(n3261), .Z(n3259) );
  NANDN U3249 ( .A(n3261), .B(n3260), .Z(n3256) );
  ANDN U3250 ( .B(B[64]), .A(n74), .Z(n3069) );
  XNOR U3251 ( .A(n3077), .B(n3262), .Z(n3070) );
  XNOR U3252 ( .A(n3076), .B(n3074), .Z(n3262) );
  AND U3253 ( .A(n3263), .B(n3264), .Z(n3074) );
  NANDN U3254 ( .A(n3265), .B(n3266), .Z(n3264) );
  OR U3255 ( .A(n3267), .B(n3268), .Z(n3266) );
  NAND U3256 ( .A(n3268), .B(n3267), .Z(n3263) );
  ANDN U3257 ( .B(B[65]), .A(n75), .Z(n3076) );
  XNOR U3258 ( .A(n3084), .B(n3269), .Z(n3077) );
  XNOR U3259 ( .A(n3083), .B(n3081), .Z(n3269) );
  AND U3260 ( .A(n3270), .B(n3271), .Z(n3081) );
  NANDN U3261 ( .A(n3272), .B(n3273), .Z(n3271) );
  NANDN U3262 ( .A(n3274), .B(n3275), .Z(n3273) );
  NANDN U3263 ( .A(n3275), .B(n3274), .Z(n3270) );
  ANDN U3264 ( .B(B[66]), .A(n76), .Z(n3083) );
  XNOR U3265 ( .A(n3091), .B(n3276), .Z(n3084) );
  XNOR U3266 ( .A(n3090), .B(n3088), .Z(n3276) );
  AND U3267 ( .A(n3277), .B(n3278), .Z(n3088) );
  NANDN U3268 ( .A(n3279), .B(n3280), .Z(n3278) );
  OR U3269 ( .A(n3281), .B(n3282), .Z(n3280) );
  NAND U3270 ( .A(n3282), .B(n3281), .Z(n3277) );
  ANDN U3271 ( .B(B[67]), .A(n77), .Z(n3090) );
  XNOR U3272 ( .A(n3098), .B(n3283), .Z(n3091) );
  XNOR U3273 ( .A(n3097), .B(n3095), .Z(n3283) );
  AND U3274 ( .A(n3284), .B(n3285), .Z(n3095) );
  NANDN U3275 ( .A(n3286), .B(n3287), .Z(n3285) );
  NANDN U3276 ( .A(n3288), .B(n3289), .Z(n3287) );
  NANDN U3277 ( .A(n3289), .B(n3288), .Z(n3284) );
  ANDN U3278 ( .B(B[68]), .A(n78), .Z(n3097) );
  XOR U3279 ( .A(n3103), .B(n3290), .Z(n3098) );
  XNOR U3280 ( .A(n3104), .B(n3105), .Z(n3290) );
  AND U3281 ( .A(n3291), .B(n3292), .Z(n3105) );
  NANDN U3282 ( .A(n3293), .B(n3294), .Z(n3292) );
  NANDN U3283 ( .A(n3295), .B(n3296), .Z(n3294) );
  ANDN U3284 ( .B(B[69]), .A(n79), .Z(n3104) );
  XOR U3285 ( .A(n3297), .B(n3298), .Z(n3103) );
  XNOR U3286 ( .A(n3299), .B(n44), .Z(n3298) );
  NAND U3287 ( .A(n3300), .B(n3301), .Z(n137) );
  NANDN U3288 ( .A(n3302), .B(n3303), .Z(n3301) );
  OR U3289 ( .A(n3304), .B(n3305), .Z(n3303) );
  NAND U3290 ( .A(n3305), .B(n3304), .Z(n3300) );
  XOR U3291 ( .A(n139), .B(n138), .Z(\A1[72] ) );
  XOR U3292 ( .A(n3305), .B(n3306), .Z(n138) );
  XNOR U3293 ( .A(n3304), .B(n3302), .Z(n3306) );
  AND U3294 ( .A(n3307), .B(n3308), .Z(n3302) );
  NANDN U3295 ( .A(n3309), .B(n3310), .Z(n3308) );
  NANDN U3296 ( .A(n3311), .B(n3312), .Z(n3310) );
  NANDN U3297 ( .A(n3312), .B(n3311), .Z(n3307) );
  ANDN U3298 ( .B(B[43]), .A(n54), .Z(n3304) );
  XNOR U3299 ( .A(n3121), .B(n3313), .Z(n3305) );
  XNOR U3300 ( .A(n3120), .B(n3118), .Z(n3313) );
  AND U3301 ( .A(n3314), .B(n3315), .Z(n3118) );
  NANDN U3302 ( .A(n3316), .B(n3317), .Z(n3315) );
  OR U3303 ( .A(n3318), .B(n3319), .Z(n3317) );
  NAND U3304 ( .A(n3319), .B(n3318), .Z(n3314) );
  ANDN U3305 ( .B(B[44]), .A(n55), .Z(n3120) );
  XNOR U3306 ( .A(n3128), .B(n3320), .Z(n3121) );
  XNOR U3307 ( .A(n3127), .B(n3125), .Z(n3320) );
  AND U3308 ( .A(n3321), .B(n3322), .Z(n3125) );
  NANDN U3309 ( .A(n3323), .B(n3324), .Z(n3322) );
  NANDN U3310 ( .A(n3325), .B(n3326), .Z(n3324) );
  NANDN U3311 ( .A(n3326), .B(n3325), .Z(n3321) );
  ANDN U3312 ( .B(B[45]), .A(n56), .Z(n3127) );
  XNOR U3313 ( .A(n3135), .B(n3327), .Z(n3128) );
  XNOR U3314 ( .A(n3134), .B(n3132), .Z(n3327) );
  AND U3315 ( .A(n3328), .B(n3329), .Z(n3132) );
  NANDN U3316 ( .A(n3330), .B(n3331), .Z(n3329) );
  OR U3317 ( .A(n3332), .B(n3333), .Z(n3331) );
  NAND U3318 ( .A(n3333), .B(n3332), .Z(n3328) );
  ANDN U3319 ( .B(B[46]), .A(n57), .Z(n3134) );
  XNOR U3320 ( .A(n3142), .B(n3334), .Z(n3135) );
  XNOR U3321 ( .A(n3141), .B(n3139), .Z(n3334) );
  AND U3322 ( .A(n3335), .B(n3336), .Z(n3139) );
  NANDN U3323 ( .A(n3337), .B(n3338), .Z(n3336) );
  NANDN U3324 ( .A(n3339), .B(n3340), .Z(n3338) );
  NANDN U3325 ( .A(n3340), .B(n3339), .Z(n3335) );
  ANDN U3326 ( .B(B[47]), .A(n58), .Z(n3141) );
  XNOR U3327 ( .A(n3149), .B(n3341), .Z(n3142) );
  XNOR U3328 ( .A(n3148), .B(n3146), .Z(n3341) );
  AND U3329 ( .A(n3342), .B(n3343), .Z(n3146) );
  NANDN U3330 ( .A(n3344), .B(n3345), .Z(n3343) );
  OR U3331 ( .A(n3346), .B(n3347), .Z(n3345) );
  NAND U3332 ( .A(n3347), .B(n3346), .Z(n3342) );
  ANDN U3333 ( .B(B[48]), .A(n59), .Z(n3148) );
  XNOR U3334 ( .A(n3156), .B(n3348), .Z(n3149) );
  XNOR U3335 ( .A(n3155), .B(n3153), .Z(n3348) );
  AND U3336 ( .A(n3349), .B(n3350), .Z(n3153) );
  NANDN U3337 ( .A(n3351), .B(n3352), .Z(n3350) );
  NANDN U3338 ( .A(n3353), .B(n3354), .Z(n3352) );
  NANDN U3339 ( .A(n3354), .B(n3353), .Z(n3349) );
  ANDN U3340 ( .B(B[49]), .A(n60), .Z(n3155) );
  XNOR U3341 ( .A(n3163), .B(n3355), .Z(n3156) );
  XNOR U3342 ( .A(n3162), .B(n3160), .Z(n3355) );
  AND U3343 ( .A(n3356), .B(n3357), .Z(n3160) );
  NANDN U3344 ( .A(n3358), .B(n3359), .Z(n3357) );
  OR U3345 ( .A(n3360), .B(n3361), .Z(n3359) );
  NAND U3346 ( .A(n3361), .B(n3360), .Z(n3356) );
  ANDN U3347 ( .B(B[50]), .A(n61), .Z(n3162) );
  XNOR U3348 ( .A(n3170), .B(n3362), .Z(n3163) );
  XNOR U3349 ( .A(n3169), .B(n3167), .Z(n3362) );
  AND U3350 ( .A(n3363), .B(n3364), .Z(n3167) );
  NANDN U3351 ( .A(n3365), .B(n3366), .Z(n3364) );
  NANDN U3352 ( .A(n3367), .B(n3368), .Z(n3366) );
  NANDN U3353 ( .A(n3368), .B(n3367), .Z(n3363) );
  ANDN U3354 ( .B(B[51]), .A(n62), .Z(n3169) );
  XNOR U3355 ( .A(n3177), .B(n3369), .Z(n3170) );
  XNOR U3356 ( .A(n3176), .B(n3174), .Z(n3369) );
  AND U3357 ( .A(n3370), .B(n3371), .Z(n3174) );
  NANDN U3358 ( .A(n3372), .B(n3373), .Z(n3371) );
  OR U3359 ( .A(n3374), .B(n3375), .Z(n3373) );
  NAND U3360 ( .A(n3375), .B(n3374), .Z(n3370) );
  ANDN U3361 ( .B(B[52]), .A(n63), .Z(n3176) );
  XNOR U3362 ( .A(n3184), .B(n3376), .Z(n3177) );
  XNOR U3363 ( .A(n3183), .B(n3181), .Z(n3376) );
  AND U3364 ( .A(n3377), .B(n3378), .Z(n3181) );
  NANDN U3365 ( .A(n3379), .B(n3380), .Z(n3378) );
  NANDN U3366 ( .A(n3381), .B(n3382), .Z(n3380) );
  NANDN U3367 ( .A(n3382), .B(n3381), .Z(n3377) );
  ANDN U3368 ( .B(B[53]), .A(n64), .Z(n3183) );
  XNOR U3369 ( .A(n3191), .B(n3383), .Z(n3184) );
  XNOR U3370 ( .A(n3190), .B(n3188), .Z(n3383) );
  AND U3371 ( .A(n3384), .B(n3385), .Z(n3188) );
  NANDN U3372 ( .A(n3386), .B(n3387), .Z(n3385) );
  OR U3373 ( .A(n3388), .B(n3389), .Z(n3387) );
  NAND U3374 ( .A(n3389), .B(n3388), .Z(n3384) );
  ANDN U3375 ( .B(B[54]), .A(n65), .Z(n3190) );
  XNOR U3376 ( .A(n3198), .B(n3390), .Z(n3191) );
  XNOR U3377 ( .A(n3197), .B(n3195), .Z(n3390) );
  AND U3378 ( .A(n3391), .B(n3392), .Z(n3195) );
  NANDN U3379 ( .A(n3393), .B(n3394), .Z(n3392) );
  NANDN U3380 ( .A(n3395), .B(n3396), .Z(n3394) );
  NANDN U3381 ( .A(n3396), .B(n3395), .Z(n3391) );
  ANDN U3382 ( .B(B[55]), .A(n66), .Z(n3197) );
  XNOR U3383 ( .A(n3205), .B(n3397), .Z(n3198) );
  XNOR U3384 ( .A(n3204), .B(n3202), .Z(n3397) );
  AND U3385 ( .A(n3398), .B(n3399), .Z(n3202) );
  NANDN U3386 ( .A(n3400), .B(n3401), .Z(n3399) );
  OR U3387 ( .A(n3402), .B(n3403), .Z(n3401) );
  NAND U3388 ( .A(n3403), .B(n3402), .Z(n3398) );
  ANDN U3389 ( .B(B[56]), .A(n67), .Z(n3204) );
  XNOR U3390 ( .A(n3212), .B(n3404), .Z(n3205) );
  XNOR U3391 ( .A(n3211), .B(n3209), .Z(n3404) );
  AND U3392 ( .A(n3405), .B(n3406), .Z(n3209) );
  NANDN U3393 ( .A(n3407), .B(n3408), .Z(n3406) );
  NANDN U3394 ( .A(n3409), .B(n3410), .Z(n3408) );
  NANDN U3395 ( .A(n3410), .B(n3409), .Z(n3405) );
  ANDN U3396 ( .B(B[57]), .A(n68), .Z(n3211) );
  XNOR U3397 ( .A(n3219), .B(n3411), .Z(n3212) );
  XNOR U3398 ( .A(n3218), .B(n3216), .Z(n3411) );
  AND U3399 ( .A(n3412), .B(n3413), .Z(n3216) );
  NANDN U3400 ( .A(n3414), .B(n3415), .Z(n3413) );
  OR U3401 ( .A(n3416), .B(n3417), .Z(n3415) );
  NAND U3402 ( .A(n3417), .B(n3416), .Z(n3412) );
  ANDN U3403 ( .B(B[58]), .A(n69), .Z(n3218) );
  XNOR U3404 ( .A(n3226), .B(n3418), .Z(n3219) );
  XNOR U3405 ( .A(n3225), .B(n3223), .Z(n3418) );
  AND U3406 ( .A(n3419), .B(n3420), .Z(n3223) );
  NANDN U3407 ( .A(n3421), .B(n3422), .Z(n3420) );
  NANDN U3408 ( .A(n3423), .B(n3424), .Z(n3422) );
  NANDN U3409 ( .A(n3424), .B(n3423), .Z(n3419) );
  ANDN U3410 ( .B(B[59]), .A(n70), .Z(n3225) );
  XNOR U3411 ( .A(n3233), .B(n3425), .Z(n3226) );
  XNOR U3412 ( .A(n3232), .B(n3230), .Z(n3425) );
  AND U3413 ( .A(n3426), .B(n3427), .Z(n3230) );
  NANDN U3414 ( .A(n3428), .B(n3429), .Z(n3427) );
  OR U3415 ( .A(n3430), .B(n3431), .Z(n3429) );
  NAND U3416 ( .A(n3431), .B(n3430), .Z(n3426) );
  ANDN U3417 ( .B(B[60]), .A(n71), .Z(n3232) );
  XNOR U3418 ( .A(n3240), .B(n3432), .Z(n3233) );
  XNOR U3419 ( .A(n3239), .B(n3237), .Z(n3432) );
  AND U3420 ( .A(n3433), .B(n3434), .Z(n3237) );
  NANDN U3421 ( .A(n3435), .B(n3436), .Z(n3434) );
  NANDN U3422 ( .A(n3437), .B(n3438), .Z(n3436) );
  NANDN U3423 ( .A(n3438), .B(n3437), .Z(n3433) );
  ANDN U3424 ( .B(B[61]), .A(n72), .Z(n3239) );
  XNOR U3425 ( .A(n3247), .B(n3439), .Z(n3240) );
  XNOR U3426 ( .A(n3246), .B(n3244), .Z(n3439) );
  AND U3427 ( .A(n3440), .B(n3441), .Z(n3244) );
  NANDN U3428 ( .A(n3442), .B(n3443), .Z(n3441) );
  OR U3429 ( .A(n3444), .B(n3445), .Z(n3443) );
  NAND U3430 ( .A(n3445), .B(n3444), .Z(n3440) );
  ANDN U3431 ( .B(B[62]), .A(n73), .Z(n3246) );
  XNOR U3432 ( .A(n3254), .B(n3446), .Z(n3247) );
  XNOR U3433 ( .A(n3253), .B(n3251), .Z(n3446) );
  AND U3434 ( .A(n3447), .B(n3448), .Z(n3251) );
  NANDN U3435 ( .A(n3449), .B(n3450), .Z(n3448) );
  NANDN U3436 ( .A(n3451), .B(n3452), .Z(n3450) );
  NANDN U3437 ( .A(n3452), .B(n3451), .Z(n3447) );
  ANDN U3438 ( .B(B[63]), .A(n74), .Z(n3253) );
  XNOR U3439 ( .A(n3261), .B(n3453), .Z(n3254) );
  XNOR U3440 ( .A(n3260), .B(n3258), .Z(n3453) );
  AND U3441 ( .A(n3454), .B(n3455), .Z(n3258) );
  NANDN U3442 ( .A(n3456), .B(n3457), .Z(n3455) );
  OR U3443 ( .A(n3458), .B(n3459), .Z(n3457) );
  NAND U3444 ( .A(n3459), .B(n3458), .Z(n3454) );
  ANDN U3445 ( .B(B[64]), .A(n75), .Z(n3260) );
  XNOR U3446 ( .A(n3268), .B(n3460), .Z(n3261) );
  XNOR U3447 ( .A(n3267), .B(n3265), .Z(n3460) );
  AND U3448 ( .A(n3461), .B(n3462), .Z(n3265) );
  NANDN U3449 ( .A(n3463), .B(n3464), .Z(n3462) );
  NANDN U3450 ( .A(n3465), .B(n3466), .Z(n3464) );
  NANDN U3451 ( .A(n3466), .B(n3465), .Z(n3461) );
  ANDN U3452 ( .B(B[65]), .A(n76), .Z(n3267) );
  XNOR U3453 ( .A(n3275), .B(n3467), .Z(n3268) );
  XNOR U3454 ( .A(n3274), .B(n3272), .Z(n3467) );
  AND U3455 ( .A(n3468), .B(n3469), .Z(n3272) );
  NANDN U3456 ( .A(n3470), .B(n3471), .Z(n3469) );
  OR U3457 ( .A(n3472), .B(n3473), .Z(n3471) );
  NAND U3458 ( .A(n3473), .B(n3472), .Z(n3468) );
  ANDN U3459 ( .B(B[66]), .A(n77), .Z(n3274) );
  XNOR U3460 ( .A(n3282), .B(n3474), .Z(n3275) );
  XNOR U3461 ( .A(n3281), .B(n3279), .Z(n3474) );
  AND U3462 ( .A(n3475), .B(n3476), .Z(n3279) );
  NANDN U3463 ( .A(n3477), .B(n3478), .Z(n3476) );
  NANDN U3464 ( .A(n3479), .B(n3480), .Z(n3478) );
  NANDN U3465 ( .A(n3480), .B(n3479), .Z(n3475) );
  ANDN U3466 ( .B(B[67]), .A(n78), .Z(n3281) );
  XNOR U3467 ( .A(n3289), .B(n3481), .Z(n3282) );
  XNOR U3468 ( .A(n3288), .B(n3286), .Z(n3481) );
  AND U3469 ( .A(n3482), .B(n3483), .Z(n3286) );
  NANDN U3470 ( .A(n3484), .B(n3485), .Z(n3483) );
  OR U3471 ( .A(n3486), .B(n3487), .Z(n3485) );
  NAND U3472 ( .A(n3487), .B(n3486), .Z(n3482) );
  ANDN U3473 ( .B(B[68]), .A(n79), .Z(n3288) );
  XOR U3474 ( .A(n3293), .B(n3488), .Z(n3289) );
  XNOR U3475 ( .A(n3295), .B(n3296), .Z(n3488) );
  AND U3476 ( .A(n3489), .B(n3490), .Z(n3296) );
  NAND U3477 ( .A(n3491), .B(n3492), .Z(n3490) );
  NANDN U3478 ( .A(n3493), .B(n3494), .Z(n3491) );
  ANDN U3479 ( .B(B[69]), .A(n80), .Z(n3295) );
  XNOR U3480 ( .A(n3495), .B(n3496), .Z(n3293) );
  XNOR U3481 ( .A(n3497), .B(n45), .Z(n3496) );
  NAND U3482 ( .A(n3498), .B(n3499), .Z(n139) );
  NANDN U3483 ( .A(n3500), .B(n3501), .Z(n3499) );
  OR U3484 ( .A(n3502), .B(n3503), .Z(n3501) );
  NAND U3485 ( .A(n3503), .B(n3502), .Z(n3498) );
  XOR U3486 ( .A(n141), .B(n140), .Z(\A1[71] ) );
  XOR U3487 ( .A(n3503), .B(n3504), .Z(n140) );
  XNOR U3488 ( .A(n3502), .B(n3500), .Z(n3504) );
  AND U3489 ( .A(n3505), .B(n3506), .Z(n3500) );
  NANDN U3490 ( .A(n3507), .B(n3508), .Z(n3506) );
  NANDN U3491 ( .A(n3509), .B(n3510), .Z(n3508) );
  NANDN U3492 ( .A(n3510), .B(n3509), .Z(n3505) );
  ANDN U3493 ( .B(B[42]), .A(n54), .Z(n3502) );
  XNOR U3494 ( .A(n3312), .B(n3511), .Z(n3503) );
  XNOR U3495 ( .A(n3311), .B(n3309), .Z(n3511) );
  AND U3496 ( .A(n3512), .B(n3513), .Z(n3309) );
  NANDN U3497 ( .A(n3514), .B(n3515), .Z(n3513) );
  OR U3498 ( .A(n3516), .B(n3517), .Z(n3515) );
  NAND U3499 ( .A(n3517), .B(n3516), .Z(n3512) );
  ANDN U3500 ( .B(B[43]), .A(n55), .Z(n3311) );
  XNOR U3501 ( .A(n3319), .B(n3518), .Z(n3312) );
  XNOR U3502 ( .A(n3318), .B(n3316), .Z(n3518) );
  AND U3503 ( .A(n3519), .B(n3520), .Z(n3316) );
  NANDN U3504 ( .A(n3521), .B(n3522), .Z(n3520) );
  NANDN U3505 ( .A(n3523), .B(n3524), .Z(n3522) );
  NANDN U3506 ( .A(n3524), .B(n3523), .Z(n3519) );
  ANDN U3507 ( .B(B[44]), .A(n56), .Z(n3318) );
  XNOR U3508 ( .A(n3326), .B(n3525), .Z(n3319) );
  XNOR U3509 ( .A(n3325), .B(n3323), .Z(n3525) );
  AND U3510 ( .A(n3526), .B(n3527), .Z(n3323) );
  NANDN U3511 ( .A(n3528), .B(n3529), .Z(n3527) );
  OR U3512 ( .A(n3530), .B(n3531), .Z(n3529) );
  NAND U3513 ( .A(n3531), .B(n3530), .Z(n3526) );
  ANDN U3514 ( .B(B[45]), .A(n57), .Z(n3325) );
  XNOR U3515 ( .A(n3333), .B(n3532), .Z(n3326) );
  XNOR U3516 ( .A(n3332), .B(n3330), .Z(n3532) );
  AND U3517 ( .A(n3533), .B(n3534), .Z(n3330) );
  NANDN U3518 ( .A(n3535), .B(n3536), .Z(n3534) );
  NANDN U3519 ( .A(n3537), .B(n3538), .Z(n3536) );
  NANDN U3520 ( .A(n3538), .B(n3537), .Z(n3533) );
  ANDN U3521 ( .B(B[46]), .A(n58), .Z(n3332) );
  XNOR U3522 ( .A(n3340), .B(n3539), .Z(n3333) );
  XNOR U3523 ( .A(n3339), .B(n3337), .Z(n3539) );
  AND U3524 ( .A(n3540), .B(n3541), .Z(n3337) );
  NANDN U3525 ( .A(n3542), .B(n3543), .Z(n3541) );
  OR U3526 ( .A(n3544), .B(n3545), .Z(n3543) );
  NAND U3527 ( .A(n3545), .B(n3544), .Z(n3540) );
  ANDN U3528 ( .B(B[47]), .A(n59), .Z(n3339) );
  XNOR U3529 ( .A(n3347), .B(n3546), .Z(n3340) );
  XNOR U3530 ( .A(n3346), .B(n3344), .Z(n3546) );
  AND U3531 ( .A(n3547), .B(n3548), .Z(n3344) );
  NANDN U3532 ( .A(n3549), .B(n3550), .Z(n3548) );
  NANDN U3533 ( .A(n3551), .B(n3552), .Z(n3550) );
  NANDN U3534 ( .A(n3552), .B(n3551), .Z(n3547) );
  ANDN U3535 ( .B(B[48]), .A(n60), .Z(n3346) );
  XNOR U3536 ( .A(n3354), .B(n3553), .Z(n3347) );
  XNOR U3537 ( .A(n3353), .B(n3351), .Z(n3553) );
  AND U3538 ( .A(n3554), .B(n3555), .Z(n3351) );
  NANDN U3539 ( .A(n3556), .B(n3557), .Z(n3555) );
  OR U3540 ( .A(n3558), .B(n3559), .Z(n3557) );
  NAND U3541 ( .A(n3559), .B(n3558), .Z(n3554) );
  ANDN U3542 ( .B(B[49]), .A(n61), .Z(n3353) );
  XNOR U3543 ( .A(n3361), .B(n3560), .Z(n3354) );
  XNOR U3544 ( .A(n3360), .B(n3358), .Z(n3560) );
  AND U3545 ( .A(n3561), .B(n3562), .Z(n3358) );
  NANDN U3546 ( .A(n3563), .B(n3564), .Z(n3562) );
  NANDN U3547 ( .A(n3565), .B(n3566), .Z(n3564) );
  NANDN U3548 ( .A(n3566), .B(n3565), .Z(n3561) );
  ANDN U3549 ( .B(B[50]), .A(n62), .Z(n3360) );
  XNOR U3550 ( .A(n3368), .B(n3567), .Z(n3361) );
  XNOR U3551 ( .A(n3367), .B(n3365), .Z(n3567) );
  AND U3552 ( .A(n3568), .B(n3569), .Z(n3365) );
  NANDN U3553 ( .A(n3570), .B(n3571), .Z(n3569) );
  OR U3554 ( .A(n3572), .B(n3573), .Z(n3571) );
  NAND U3555 ( .A(n3573), .B(n3572), .Z(n3568) );
  ANDN U3556 ( .B(B[51]), .A(n63), .Z(n3367) );
  XNOR U3557 ( .A(n3375), .B(n3574), .Z(n3368) );
  XNOR U3558 ( .A(n3374), .B(n3372), .Z(n3574) );
  AND U3559 ( .A(n3575), .B(n3576), .Z(n3372) );
  NANDN U3560 ( .A(n3577), .B(n3578), .Z(n3576) );
  NANDN U3561 ( .A(n3579), .B(n3580), .Z(n3578) );
  NANDN U3562 ( .A(n3580), .B(n3579), .Z(n3575) );
  ANDN U3563 ( .B(B[52]), .A(n64), .Z(n3374) );
  XNOR U3564 ( .A(n3382), .B(n3581), .Z(n3375) );
  XNOR U3565 ( .A(n3381), .B(n3379), .Z(n3581) );
  AND U3566 ( .A(n3582), .B(n3583), .Z(n3379) );
  NANDN U3567 ( .A(n3584), .B(n3585), .Z(n3583) );
  OR U3568 ( .A(n3586), .B(n3587), .Z(n3585) );
  NAND U3569 ( .A(n3587), .B(n3586), .Z(n3582) );
  ANDN U3570 ( .B(B[53]), .A(n65), .Z(n3381) );
  XNOR U3571 ( .A(n3389), .B(n3588), .Z(n3382) );
  XNOR U3572 ( .A(n3388), .B(n3386), .Z(n3588) );
  AND U3573 ( .A(n3589), .B(n3590), .Z(n3386) );
  NANDN U3574 ( .A(n3591), .B(n3592), .Z(n3590) );
  NANDN U3575 ( .A(n3593), .B(n3594), .Z(n3592) );
  NANDN U3576 ( .A(n3594), .B(n3593), .Z(n3589) );
  ANDN U3577 ( .B(B[54]), .A(n66), .Z(n3388) );
  XNOR U3578 ( .A(n3396), .B(n3595), .Z(n3389) );
  XNOR U3579 ( .A(n3395), .B(n3393), .Z(n3595) );
  AND U3580 ( .A(n3596), .B(n3597), .Z(n3393) );
  NANDN U3581 ( .A(n3598), .B(n3599), .Z(n3597) );
  OR U3582 ( .A(n3600), .B(n3601), .Z(n3599) );
  NAND U3583 ( .A(n3601), .B(n3600), .Z(n3596) );
  ANDN U3584 ( .B(B[55]), .A(n67), .Z(n3395) );
  XNOR U3585 ( .A(n3403), .B(n3602), .Z(n3396) );
  XNOR U3586 ( .A(n3402), .B(n3400), .Z(n3602) );
  AND U3587 ( .A(n3603), .B(n3604), .Z(n3400) );
  NANDN U3588 ( .A(n3605), .B(n3606), .Z(n3604) );
  NANDN U3589 ( .A(n3607), .B(n3608), .Z(n3606) );
  NANDN U3590 ( .A(n3608), .B(n3607), .Z(n3603) );
  ANDN U3591 ( .B(B[56]), .A(n68), .Z(n3402) );
  XNOR U3592 ( .A(n3410), .B(n3609), .Z(n3403) );
  XNOR U3593 ( .A(n3409), .B(n3407), .Z(n3609) );
  AND U3594 ( .A(n3610), .B(n3611), .Z(n3407) );
  NANDN U3595 ( .A(n3612), .B(n3613), .Z(n3611) );
  OR U3596 ( .A(n3614), .B(n3615), .Z(n3613) );
  NAND U3597 ( .A(n3615), .B(n3614), .Z(n3610) );
  ANDN U3598 ( .B(B[57]), .A(n69), .Z(n3409) );
  XNOR U3599 ( .A(n3417), .B(n3616), .Z(n3410) );
  XNOR U3600 ( .A(n3416), .B(n3414), .Z(n3616) );
  AND U3601 ( .A(n3617), .B(n3618), .Z(n3414) );
  NANDN U3602 ( .A(n3619), .B(n3620), .Z(n3618) );
  NANDN U3603 ( .A(n3621), .B(n3622), .Z(n3620) );
  NANDN U3604 ( .A(n3622), .B(n3621), .Z(n3617) );
  ANDN U3605 ( .B(B[58]), .A(n70), .Z(n3416) );
  XNOR U3606 ( .A(n3424), .B(n3623), .Z(n3417) );
  XNOR U3607 ( .A(n3423), .B(n3421), .Z(n3623) );
  AND U3608 ( .A(n3624), .B(n3625), .Z(n3421) );
  NANDN U3609 ( .A(n3626), .B(n3627), .Z(n3625) );
  OR U3610 ( .A(n3628), .B(n3629), .Z(n3627) );
  NAND U3611 ( .A(n3629), .B(n3628), .Z(n3624) );
  ANDN U3612 ( .B(B[59]), .A(n71), .Z(n3423) );
  XNOR U3613 ( .A(n3431), .B(n3630), .Z(n3424) );
  XNOR U3614 ( .A(n3430), .B(n3428), .Z(n3630) );
  AND U3615 ( .A(n3631), .B(n3632), .Z(n3428) );
  NANDN U3616 ( .A(n3633), .B(n3634), .Z(n3632) );
  NANDN U3617 ( .A(n3635), .B(n3636), .Z(n3634) );
  NANDN U3618 ( .A(n3636), .B(n3635), .Z(n3631) );
  ANDN U3619 ( .B(B[60]), .A(n72), .Z(n3430) );
  XNOR U3620 ( .A(n3438), .B(n3637), .Z(n3431) );
  XNOR U3621 ( .A(n3437), .B(n3435), .Z(n3637) );
  AND U3622 ( .A(n3638), .B(n3639), .Z(n3435) );
  NANDN U3623 ( .A(n3640), .B(n3641), .Z(n3639) );
  OR U3624 ( .A(n3642), .B(n3643), .Z(n3641) );
  NAND U3625 ( .A(n3643), .B(n3642), .Z(n3638) );
  ANDN U3626 ( .B(B[61]), .A(n73), .Z(n3437) );
  XNOR U3627 ( .A(n3445), .B(n3644), .Z(n3438) );
  XNOR U3628 ( .A(n3444), .B(n3442), .Z(n3644) );
  AND U3629 ( .A(n3645), .B(n3646), .Z(n3442) );
  NANDN U3630 ( .A(n3647), .B(n3648), .Z(n3646) );
  NANDN U3631 ( .A(n3649), .B(n3650), .Z(n3648) );
  NANDN U3632 ( .A(n3650), .B(n3649), .Z(n3645) );
  ANDN U3633 ( .B(B[62]), .A(n74), .Z(n3444) );
  XNOR U3634 ( .A(n3452), .B(n3651), .Z(n3445) );
  XNOR U3635 ( .A(n3451), .B(n3449), .Z(n3651) );
  AND U3636 ( .A(n3652), .B(n3653), .Z(n3449) );
  NANDN U3637 ( .A(n3654), .B(n3655), .Z(n3653) );
  OR U3638 ( .A(n3656), .B(n3657), .Z(n3655) );
  NAND U3639 ( .A(n3657), .B(n3656), .Z(n3652) );
  ANDN U3640 ( .B(B[63]), .A(n75), .Z(n3451) );
  XNOR U3641 ( .A(n3459), .B(n3658), .Z(n3452) );
  XNOR U3642 ( .A(n3458), .B(n3456), .Z(n3658) );
  AND U3643 ( .A(n3659), .B(n3660), .Z(n3456) );
  NANDN U3644 ( .A(n3661), .B(n3662), .Z(n3660) );
  NANDN U3645 ( .A(n3663), .B(n3664), .Z(n3662) );
  NANDN U3646 ( .A(n3664), .B(n3663), .Z(n3659) );
  ANDN U3647 ( .B(B[64]), .A(n76), .Z(n3458) );
  XNOR U3648 ( .A(n3466), .B(n3665), .Z(n3459) );
  XNOR U3649 ( .A(n3465), .B(n3463), .Z(n3665) );
  AND U3650 ( .A(n3666), .B(n3667), .Z(n3463) );
  NANDN U3651 ( .A(n3668), .B(n3669), .Z(n3667) );
  OR U3652 ( .A(n3670), .B(n3671), .Z(n3669) );
  NAND U3653 ( .A(n3671), .B(n3670), .Z(n3666) );
  ANDN U3654 ( .B(B[65]), .A(n77), .Z(n3465) );
  XNOR U3655 ( .A(n3473), .B(n3672), .Z(n3466) );
  XNOR U3656 ( .A(n3472), .B(n3470), .Z(n3672) );
  AND U3657 ( .A(n3673), .B(n3674), .Z(n3470) );
  NANDN U3658 ( .A(n3675), .B(n3676), .Z(n3674) );
  NANDN U3659 ( .A(n3677), .B(n3678), .Z(n3676) );
  NANDN U3660 ( .A(n3678), .B(n3677), .Z(n3673) );
  ANDN U3661 ( .B(B[66]), .A(n78), .Z(n3472) );
  XNOR U3662 ( .A(n3480), .B(n3679), .Z(n3473) );
  XNOR U3663 ( .A(n3479), .B(n3477), .Z(n3679) );
  AND U3664 ( .A(n3680), .B(n3681), .Z(n3477) );
  NANDN U3665 ( .A(n3682), .B(n3683), .Z(n3681) );
  OR U3666 ( .A(n3684), .B(n3685), .Z(n3683) );
  NAND U3667 ( .A(n3685), .B(n3684), .Z(n3680) );
  ANDN U3668 ( .B(B[67]), .A(n79), .Z(n3479) );
  XNOR U3669 ( .A(n3487), .B(n3686), .Z(n3480) );
  XNOR U3670 ( .A(n3486), .B(n3484), .Z(n3686) );
  AND U3671 ( .A(n3687), .B(n3688), .Z(n3484) );
  NANDN U3672 ( .A(n3689), .B(n3690), .Z(n3688) );
  NANDN U3673 ( .A(n3691), .B(n3692), .Z(n3690) );
  NANDN U3674 ( .A(n3692), .B(n3691), .Z(n3687) );
  ANDN U3675 ( .B(B[68]), .A(n80), .Z(n3486) );
  XOR U3676 ( .A(n3492), .B(n3693), .Z(n3487) );
  XNOR U3677 ( .A(n3493), .B(n3494), .Z(n3693) );
  AND U3678 ( .A(n3694), .B(n3695), .Z(n3494) );
  NANDN U3679 ( .A(n3696), .B(n3697), .Z(n3695) );
  NANDN U3680 ( .A(n3698), .B(n3699), .Z(n3697) );
  ANDN U3681 ( .B(B[69]), .A(n81), .Z(n3493) );
  XNOR U3682 ( .A(n3700), .B(n3701), .Z(n3492) );
  XNOR U3683 ( .A(n3702), .B(n47), .Z(n3701) );
  NAND U3684 ( .A(n3703), .B(n3704), .Z(n141) );
  NANDN U3685 ( .A(n3705), .B(n3706), .Z(n3704) );
  OR U3686 ( .A(n3707), .B(n3708), .Z(n3706) );
  NAND U3687 ( .A(n3708), .B(n3707), .Z(n3703) );
  XOR U3688 ( .A(n143), .B(n142), .Z(\A1[70] ) );
  XOR U3689 ( .A(n3708), .B(n3709), .Z(n142) );
  XNOR U3690 ( .A(n3707), .B(n3705), .Z(n3709) );
  AND U3691 ( .A(n3710), .B(n3711), .Z(n3705) );
  NANDN U3692 ( .A(n3712), .B(n3713), .Z(n3711) );
  NANDN U3693 ( .A(n3714), .B(n3715), .Z(n3713) );
  NANDN U3694 ( .A(n3715), .B(n3714), .Z(n3710) );
  ANDN U3695 ( .B(B[41]), .A(n54), .Z(n3707) );
  XNOR U3696 ( .A(n3510), .B(n3716), .Z(n3708) );
  XNOR U3697 ( .A(n3509), .B(n3507), .Z(n3716) );
  AND U3698 ( .A(n3717), .B(n3718), .Z(n3507) );
  NANDN U3699 ( .A(n3719), .B(n3720), .Z(n3718) );
  OR U3700 ( .A(n3721), .B(n3722), .Z(n3720) );
  NAND U3701 ( .A(n3722), .B(n3721), .Z(n3717) );
  ANDN U3702 ( .B(B[42]), .A(n55), .Z(n3509) );
  XNOR U3703 ( .A(n3517), .B(n3723), .Z(n3510) );
  XNOR U3704 ( .A(n3516), .B(n3514), .Z(n3723) );
  AND U3705 ( .A(n3724), .B(n3725), .Z(n3514) );
  NANDN U3706 ( .A(n3726), .B(n3727), .Z(n3725) );
  NANDN U3707 ( .A(n3728), .B(n3729), .Z(n3727) );
  NANDN U3708 ( .A(n3729), .B(n3728), .Z(n3724) );
  ANDN U3709 ( .B(B[43]), .A(n56), .Z(n3516) );
  XNOR U3710 ( .A(n3524), .B(n3730), .Z(n3517) );
  XNOR U3711 ( .A(n3523), .B(n3521), .Z(n3730) );
  AND U3712 ( .A(n3731), .B(n3732), .Z(n3521) );
  NANDN U3713 ( .A(n3733), .B(n3734), .Z(n3732) );
  OR U3714 ( .A(n3735), .B(n3736), .Z(n3734) );
  NAND U3715 ( .A(n3736), .B(n3735), .Z(n3731) );
  ANDN U3716 ( .B(B[44]), .A(n57), .Z(n3523) );
  XNOR U3717 ( .A(n3531), .B(n3737), .Z(n3524) );
  XNOR U3718 ( .A(n3530), .B(n3528), .Z(n3737) );
  AND U3719 ( .A(n3738), .B(n3739), .Z(n3528) );
  NANDN U3720 ( .A(n3740), .B(n3741), .Z(n3739) );
  NANDN U3721 ( .A(n3742), .B(n3743), .Z(n3741) );
  NANDN U3722 ( .A(n3743), .B(n3742), .Z(n3738) );
  ANDN U3723 ( .B(B[45]), .A(n58), .Z(n3530) );
  XNOR U3724 ( .A(n3538), .B(n3744), .Z(n3531) );
  XNOR U3725 ( .A(n3537), .B(n3535), .Z(n3744) );
  AND U3726 ( .A(n3745), .B(n3746), .Z(n3535) );
  NANDN U3727 ( .A(n3747), .B(n3748), .Z(n3746) );
  OR U3728 ( .A(n3749), .B(n3750), .Z(n3748) );
  NAND U3729 ( .A(n3750), .B(n3749), .Z(n3745) );
  ANDN U3730 ( .B(B[46]), .A(n59), .Z(n3537) );
  XNOR U3731 ( .A(n3545), .B(n3751), .Z(n3538) );
  XNOR U3732 ( .A(n3544), .B(n3542), .Z(n3751) );
  AND U3733 ( .A(n3752), .B(n3753), .Z(n3542) );
  NANDN U3734 ( .A(n3754), .B(n3755), .Z(n3753) );
  NANDN U3735 ( .A(n3756), .B(n3757), .Z(n3755) );
  NANDN U3736 ( .A(n3757), .B(n3756), .Z(n3752) );
  ANDN U3737 ( .B(B[47]), .A(n60), .Z(n3544) );
  XNOR U3738 ( .A(n3552), .B(n3758), .Z(n3545) );
  XNOR U3739 ( .A(n3551), .B(n3549), .Z(n3758) );
  AND U3740 ( .A(n3759), .B(n3760), .Z(n3549) );
  NANDN U3741 ( .A(n3761), .B(n3762), .Z(n3760) );
  OR U3742 ( .A(n3763), .B(n3764), .Z(n3762) );
  NAND U3743 ( .A(n3764), .B(n3763), .Z(n3759) );
  ANDN U3744 ( .B(B[48]), .A(n61), .Z(n3551) );
  XNOR U3745 ( .A(n3559), .B(n3765), .Z(n3552) );
  XNOR U3746 ( .A(n3558), .B(n3556), .Z(n3765) );
  AND U3747 ( .A(n3766), .B(n3767), .Z(n3556) );
  NANDN U3748 ( .A(n3768), .B(n3769), .Z(n3767) );
  NANDN U3749 ( .A(n3770), .B(n3771), .Z(n3769) );
  NANDN U3750 ( .A(n3771), .B(n3770), .Z(n3766) );
  ANDN U3751 ( .B(B[49]), .A(n62), .Z(n3558) );
  XNOR U3752 ( .A(n3566), .B(n3772), .Z(n3559) );
  XNOR U3753 ( .A(n3565), .B(n3563), .Z(n3772) );
  AND U3754 ( .A(n3773), .B(n3774), .Z(n3563) );
  NANDN U3755 ( .A(n3775), .B(n3776), .Z(n3774) );
  OR U3756 ( .A(n3777), .B(n3778), .Z(n3776) );
  NAND U3757 ( .A(n3778), .B(n3777), .Z(n3773) );
  ANDN U3758 ( .B(B[50]), .A(n63), .Z(n3565) );
  XNOR U3759 ( .A(n3573), .B(n3779), .Z(n3566) );
  XNOR U3760 ( .A(n3572), .B(n3570), .Z(n3779) );
  AND U3761 ( .A(n3780), .B(n3781), .Z(n3570) );
  NANDN U3762 ( .A(n3782), .B(n3783), .Z(n3781) );
  NANDN U3763 ( .A(n3784), .B(n3785), .Z(n3783) );
  NANDN U3764 ( .A(n3785), .B(n3784), .Z(n3780) );
  ANDN U3765 ( .B(B[51]), .A(n64), .Z(n3572) );
  XNOR U3766 ( .A(n3580), .B(n3786), .Z(n3573) );
  XNOR U3767 ( .A(n3579), .B(n3577), .Z(n3786) );
  AND U3768 ( .A(n3787), .B(n3788), .Z(n3577) );
  NANDN U3769 ( .A(n3789), .B(n3790), .Z(n3788) );
  OR U3770 ( .A(n3791), .B(n3792), .Z(n3790) );
  NAND U3771 ( .A(n3792), .B(n3791), .Z(n3787) );
  ANDN U3772 ( .B(B[52]), .A(n65), .Z(n3579) );
  XNOR U3773 ( .A(n3587), .B(n3793), .Z(n3580) );
  XNOR U3774 ( .A(n3586), .B(n3584), .Z(n3793) );
  AND U3775 ( .A(n3794), .B(n3795), .Z(n3584) );
  NANDN U3776 ( .A(n3796), .B(n3797), .Z(n3795) );
  NANDN U3777 ( .A(n3798), .B(n3799), .Z(n3797) );
  NANDN U3778 ( .A(n3799), .B(n3798), .Z(n3794) );
  ANDN U3779 ( .B(B[53]), .A(n66), .Z(n3586) );
  XNOR U3780 ( .A(n3594), .B(n3800), .Z(n3587) );
  XNOR U3781 ( .A(n3593), .B(n3591), .Z(n3800) );
  AND U3782 ( .A(n3801), .B(n3802), .Z(n3591) );
  NANDN U3783 ( .A(n3803), .B(n3804), .Z(n3802) );
  OR U3784 ( .A(n3805), .B(n3806), .Z(n3804) );
  NAND U3785 ( .A(n3806), .B(n3805), .Z(n3801) );
  ANDN U3786 ( .B(B[54]), .A(n67), .Z(n3593) );
  XNOR U3787 ( .A(n3601), .B(n3807), .Z(n3594) );
  XNOR U3788 ( .A(n3600), .B(n3598), .Z(n3807) );
  AND U3789 ( .A(n3808), .B(n3809), .Z(n3598) );
  NANDN U3790 ( .A(n3810), .B(n3811), .Z(n3809) );
  NANDN U3791 ( .A(n3812), .B(n3813), .Z(n3811) );
  NANDN U3792 ( .A(n3813), .B(n3812), .Z(n3808) );
  ANDN U3793 ( .B(B[55]), .A(n68), .Z(n3600) );
  XNOR U3794 ( .A(n3608), .B(n3814), .Z(n3601) );
  XNOR U3795 ( .A(n3607), .B(n3605), .Z(n3814) );
  AND U3796 ( .A(n3815), .B(n3816), .Z(n3605) );
  NANDN U3797 ( .A(n3817), .B(n3818), .Z(n3816) );
  OR U3798 ( .A(n3819), .B(n3820), .Z(n3818) );
  NAND U3799 ( .A(n3820), .B(n3819), .Z(n3815) );
  ANDN U3800 ( .B(B[56]), .A(n69), .Z(n3607) );
  XNOR U3801 ( .A(n3615), .B(n3821), .Z(n3608) );
  XNOR U3802 ( .A(n3614), .B(n3612), .Z(n3821) );
  AND U3803 ( .A(n3822), .B(n3823), .Z(n3612) );
  NANDN U3804 ( .A(n3824), .B(n3825), .Z(n3823) );
  NANDN U3805 ( .A(n3826), .B(n3827), .Z(n3825) );
  NANDN U3806 ( .A(n3827), .B(n3826), .Z(n3822) );
  ANDN U3807 ( .B(B[57]), .A(n70), .Z(n3614) );
  XNOR U3808 ( .A(n3622), .B(n3828), .Z(n3615) );
  XNOR U3809 ( .A(n3621), .B(n3619), .Z(n3828) );
  AND U3810 ( .A(n3829), .B(n3830), .Z(n3619) );
  NANDN U3811 ( .A(n3831), .B(n3832), .Z(n3830) );
  OR U3812 ( .A(n3833), .B(n3834), .Z(n3832) );
  NAND U3813 ( .A(n3834), .B(n3833), .Z(n3829) );
  ANDN U3814 ( .B(B[58]), .A(n71), .Z(n3621) );
  XNOR U3815 ( .A(n3629), .B(n3835), .Z(n3622) );
  XNOR U3816 ( .A(n3628), .B(n3626), .Z(n3835) );
  AND U3817 ( .A(n3836), .B(n3837), .Z(n3626) );
  NANDN U3818 ( .A(n3838), .B(n3839), .Z(n3837) );
  NANDN U3819 ( .A(n3840), .B(n3841), .Z(n3839) );
  NANDN U3820 ( .A(n3841), .B(n3840), .Z(n3836) );
  ANDN U3821 ( .B(B[59]), .A(n72), .Z(n3628) );
  XNOR U3822 ( .A(n3636), .B(n3842), .Z(n3629) );
  XNOR U3823 ( .A(n3635), .B(n3633), .Z(n3842) );
  AND U3824 ( .A(n3843), .B(n3844), .Z(n3633) );
  NANDN U3825 ( .A(n3845), .B(n3846), .Z(n3844) );
  OR U3826 ( .A(n3847), .B(n3848), .Z(n3846) );
  NAND U3827 ( .A(n3848), .B(n3847), .Z(n3843) );
  ANDN U3828 ( .B(B[60]), .A(n73), .Z(n3635) );
  XNOR U3829 ( .A(n3643), .B(n3849), .Z(n3636) );
  XNOR U3830 ( .A(n3642), .B(n3640), .Z(n3849) );
  AND U3831 ( .A(n3850), .B(n3851), .Z(n3640) );
  NANDN U3832 ( .A(n3852), .B(n3853), .Z(n3851) );
  NANDN U3833 ( .A(n3854), .B(n3855), .Z(n3853) );
  NANDN U3834 ( .A(n3855), .B(n3854), .Z(n3850) );
  ANDN U3835 ( .B(B[61]), .A(n74), .Z(n3642) );
  XNOR U3836 ( .A(n3650), .B(n3856), .Z(n3643) );
  XNOR U3837 ( .A(n3649), .B(n3647), .Z(n3856) );
  AND U3838 ( .A(n3857), .B(n3858), .Z(n3647) );
  NANDN U3839 ( .A(n3859), .B(n3860), .Z(n3858) );
  OR U3840 ( .A(n3861), .B(n3862), .Z(n3860) );
  NAND U3841 ( .A(n3862), .B(n3861), .Z(n3857) );
  ANDN U3842 ( .B(B[62]), .A(n75), .Z(n3649) );
  XNOR U3843 ( .A(n3657), .B(n3863), .Z(n3650) );
  XNOR U3844 ( .A(n3656), .B(n3654), .Z(n3863) );
  AND U3845 ( .A(n3864), .B(n3865), .Z(n3654) );
  NANDN U3846 ( .A(n3866), .B(n3867), .Z(n3865) );
  NANDN U3847 ( .A(n3868), .B(n3869), .Z(n3867) );
  NANDN U3848 ( .A(n3869), .B(n3868), .Z(n3864) );
  ANDN U3849 ( .B(B[63]), .A(n76), .Z(n3656) );
  XNOR U3850 ( .A(n3664), .B(n3870), .Z(n3657) );
  XNOR U3851 ( .A(n3663), .B(n3661), .Z(n3870) );
  AND U3852 ( .A(n3871), .B(n3872), .Z(n3661) );
  NANDN U3853 ( .A(n3873), .B(n3874), .Z(n3872) );
  OR U3854 ( .A(n3875), .B(n3876), .Z(n3874) );
  NAND U3855 ( .A(n3876), .B(n3875), .Z(n3871) );
  ANDN U3856 ( .B(B[64]), .A(n77), .Z(n3663) );
  XNOR U3857 ( .A(n3671), .B(n3877), .Z(n3664) );
  XNOR U3858 ( .A(n3670), .B(n3668), .Z(n3877) );
  AND U3859 ( .A(n3878), .B(n3879), .Z(n3668) );
  NANDN U3860 ( .A(n3880), .B(n3881), .Z(n3879) );
  NANDN U3861 ( .A(n3882), .B(n3883), .Z(n3881) );
  NANDN U3862 ( .A(n3883), .B(n3882), .Z(n3878) );
  ANDN U3863 ( .B(B[65]), .A(n78), .Z(n3670) );
  XNOR U3864 ( .A(n3678), .B(n3884), .Z(n3671) );
  XNOR U3865 ( .A(n3677), .B(n3675), .Z(n3884) );
  AND U3866 ( .A(n3885), .B(n3886), .Z(n3675) );
  NANDN U3867 ( .A(n3887), .B(n3888), .Z(n3886) );
  OR U3868 ( .A(n3889), .B(n3890), .Z(n3888) );
  NAND U3869 ( .A(n3890), .B(n3889), .Z(n3885) );
  ANDN U3870 ( .B(B[66]), .A(n79), .Z(n3677) );
  XNOR U3871 ( .A(n3685), .B(n3891), .Z(n3678) );
  XNOR U3872 ( .A(n3684), .B(n3682), .Z(n3891) );
  AND U3873 ( .A(n3892), .B(n3893), .Z(n3682) );
  NANDN U3874 ( .A(n3894), .B(n3895), .Z(n3893) );
  NANDN U3875 ( .A(n3896), .B(n3897), .Z(n3895) );
  NANDN U3876 ( .A(n3897), .B(n3896), .Z(n3892) );
  ANDN U3877 ( .B(B[67]), .A(n80), .Z(n3684) );
  XNOR U3878 ( .A(n3692), .B(n3898), .Z(n3685) );
  XNOR U3879 ( .A(n3691), .B(n3689), .Z(n3898) );
  AND U3880 ( .A(n3899), .B(n3900), .Z(n3689) );
  NANDN U3881 ( .A(n3901), .B(n3902), .Z(n3900) );
  NANDN U3882 ( .A(n3903), .B(n3904), .Z(n3902) );
  NAND U3883 ( .A(n48), .B(n3903), .Z(n3899) );
  ANDN U3884 ( .B(B[68]), .A(n81), .Z(n3691) );
  XOR U3885 ( .A(n3696), .B(n3905), .Z(n3692) );
  XNOR U3886 ( .A(n3698), .B(n3699), .Z(n3905) );
  AND U3887 ( .A(n3906), .B(n3907), .Z(n3699) );
  NANDN U3888 ( .A(n3908), .B(n3909), .Z(n3907) );
  NANDN U3889 ( .A(n3910), .B(n3911), .Z(n3909) );
  NANDN U3890 ( .A(n3911), .B(n3910), .Z(n3906) );
  ANDN U3891 ( .B(B[69]), .A(n82), .Z(n3698) );
  XNOR U3892 ( .A(n3912), .B(n3913), .Z(n3696) );
  XOR U3893 ( .A(n3914), .B(n3915), .Z(n3913) );
  NAND U3894 ( .A(n3916), .B(n3917), .Z(n143) );
  NANDN U3895 ( .A(n3918), .B(n3919), .Z(n3917) );
  OR U3896 ( .A(n3920), .B(n3921), .Z(n3919) );
  NAND U3897 ( .A(n3921), .B(n3920), .Z(n3916) );
  XNOR U3898 ( .A(n3922), .B(n3923), .Z(\A1[6] ) );
  XNOR U3899 ( .A(n3924), .B(n3925), .Z(n3923) );
  XOR U3900 ( .A(n145), .B(n144), .Z(\A1[69] ) );
  XOR U3901 ( .A(n3921), .B(n3926), .Z(n144) );
  XNOR U3902 ( .A(n3920), .B(n3918), .Z(n3926) );
  AND U3903 ( .A(n3927), .B(n3928), .Z(n3918) );
  NANDN U3904 ( .A(n3929), .B(n3930), .Z(n3928) );
  NANDN U3905 ( .A(n3931), .B(n3932), .Z(n3930) );
  NANDN U3906 ( .A(n3932), .B(n3931), .Z(n3927) );
  ANDN U3907 ( .B(B[40]), .A(n54), .Z(n3920) );
  XNOR U3908 ( .A(n3715), .B(n3933), .Z(n3921) );
  XNOR U3909 ( .A(n3714), .B(n3712), .Z(n3933) );
  AND U3910 ( .A(n3934), .B(n3935), .Z(n3712) );
  NANDN U3911 ( .A(n3936), .B(n3937), .Z(n3935) );
  OR U3912 ( .A(n3938), .B(n3939), .Z(n3937) );
  NAND U3913 ( .A(n3939), .B(n3938), .Z(n3934) );
  ANDN U3914 ( .B(B[41]), .A(n55), .Z(n3714) );
  XNOR U3915 ( .A(n3722), .B(n3940), .Z(n3715) );
  XNOR U3916 ( .A(n3721), .B(n3719), .Z(n3940) );
  AND U3917 ( .A(n3941), .B(n3942), .Z(n3719) );
  NANDN U3918 ( .A(n3943), .B(n3944), .Z(n3942) );
  NANDN U3919 ( .A(n3945), .B(n3946), .Z(n3944) );
  NANDN U3920 ( .A(n3946), .B(n3945), .Z(n3941) );
  ANDN U3921 ( .B(B[42]), .A(n56), .Z(n3721) );
  XNOR U3922 ( .A(n3729), .B(n3947), .Z(n3722) );
  XNOR U3923 ( .A(n3728), .B(n3726), .Z(n3947) );
  AND U3924 ( .A(n3948), .B(n3949), .Z(n3726) );
  NANDN U3925 ( .A(n3950), .B(n3951), .Z(n3949) );
  OR U3926 ( .A(n3952), .B(n3953), .Z(n3951) );
  NAND U3927 ( .A(n3953), .B(n3952), .Z(n3948) );
  ANDN U3928 ( .B(B[43]), .A(n57), .Z(n3728) );
  XNOR U3929 ( .A(n3736), .B(n3954), .Z(n3729) );
  XNOR U3930 ( .A(n3735), .B(n3733), .Z(n3954) );
  AND U3931 ( .A(n3955), .B(n3956), .Z(n3733) );
  NANDN U3932 ( .A(n3957), .B(n3958), .Z(n3956) );
  NANDN U3933 ( .A(n3959), .B(n3960), .Z(n3958) );
  NANDN U3934 ( .A(n3960), .B(n3959), .Z(n3955) );
  ANDN U3935 ( .B(B[44]), .A(n58), .Z(n3735) );
  XNOR U3936 ( .A(n3743), .B(n3961), .Z(n3736) );
  XNOR U3937 ( .A(n3742), .B(n3740), .Z(n3961) );
  AND U3938 ( .A(n3962), .B(n3963), .Z(n3740) );
  NANDN U3939 ( .A(n3964), .B(n3965), .Z(n3963) );
  OR U3940 ( .A(n3966), .B(n3967), .Z(n3965) );
  NAND U3941 ( .A(n3967), .B(n3966), .Z(n3962) );
  ANDN U3942 ( .B(B[45]), .A(n59), .Z(n3742) );
  XNOR U3943 ( .A(n3750), .B(n3968), .Z(n3743) );
  XNOR U3944 ( .A(n3749), .B(n3747), .Z(n3968) );
  AND U3945 ( .A(n3969), .B(n3970), .Z(n3747) );
  NANDN U3946 ( .A(n3971), .B(n3972), .Z(n3970) );
  NANDN U3947 ( .A(n3973), .B(n3974), .Z(n3972) );
  NANDN U3948 ( .A(n3974), .B(n3973), .Z(n3969) );
  ANDN U3949 ( .B(B[46]), .A(n60), .Z(n3749) );
  XNOR U3950 ( .A(n3757), .B(n3975), .Z(n3750) );
  XNOR U3951 ( .A(n3756), .B(n3754), .Z(n3975) );
  AND U3952 ( .A(n3976), .B(n3977), .Z(n3754) );
  NANDN U3953 ( .A(n3978), .B(n3979), .Z(n3977) );
  OR U3954 ( .A(n3980), .B(n3981), .Z(n3979) );
  NAND U3955 ( .A(n3981), .B(n3980), .Z(n3976) );
  ANDN U3956 ( .B(B[47]), .A(n61), .Z(n3756) );
  XNOR U3957 ( .A(n3764), .B(n3982), .Z(n3757) );
  XNOR U3958 ( .A(n3763), .B(n3761), .Z(n3982) );
  AND U3959 ( .A(n3983), .B(n3984), .Z(n3761) );
  NANDN U3960 ( .A(n3985), .B(n3986), .Z(n3984) );
  NANDN U3961 ( .A(n3987), .B(n3988), .Z(n3986) );
  NANDN U3962 ( .A(n3988), .B(n3987), .Z(n3983) );
  ANDN U3963 ( .B(B[48]), .A(n62), .Z(n3763) );
  XNOR U3964 ( .A(n3771), .B(n3989), .Z(n3764) );
  XNOR U3965 ( .A(n3770), .B(n3768), .Z(n3989) );
  AND U3966 ( .A(n3990), .B(n3991), .Z(n3768) );
  NANDN U3967 ( .A(n3992), .B(n3993), .Z(n3991) );
  OR U3968 ( .A(n3994), .B(n3995), .Z(n3993) );
  NAND U3969 ( .A(n3995), .B(n3994), .Z(n3990) );
  ANDN U3970 ( .B(B[49]), .A(n63), .Z(n3770) );
  XNOR U3971 ( .A(n3778), .B(n3996), .Z(n3771) );
  XNOR U3972 ( .A(n3777), .B(n3775), .Z(n3996) );
  AND U3973 ( .A(n3997), .B(n3998), .Z(n3775) );
  NANDN U3974 ( .A(n3999), .B(n4000), .Z(n3998) );
  NANDN U3975 ( .A(n4001), .B(n4002), .Z(n4000) );
  NANDN U3976 ( .A(n4002), .B(n4001), .Z(n3997) );
  ANDN U3977 ( .B(B[50]), .A(n64), .Z(n3777) );
  XNOR U3978 ( .A(n3785), .B(n4003), .Z(n3778) );
  XNOR U3979 ( .A(n3784), .B(n3782), .Z(n4003) );
  AND U3980 ( .A(n4004), .B(n4005), .Z(n3782) );
  NANDN U3981 ( .A(n4006), .B(n4007), .Z(n4005) );
  OR U3982 ( .A(n4008), .B(n4009), .Z(n4007) );
  NAND U3983 ( .A(n4009), .B(n4008), .Z(n4004) );
  ANDN U3984 ( .B(B[51]), .A(n65), .Z(n3784) );
  XNOR U3985 ( .A(n3792), .B(n4010), .Z(n3785) );
  XNOR U3986 ( .A(n3791), .B(n3789), .Z(n4010) );
  AND U3987 ( .A(n4011), .B(n4012), .Z(n3789) );
  NANDN U3988 ( .A(n4013), .B(n4014), .Z(n4012) );
  NANDN U3989 ( .A(n4015), .B(n4016), .Z(n4014) );
  NANDN U3990 ( .A(n4016), .B(n4015), .Z(n4011) );
  ANDN U3991 ( .B(B[52]), .A(n66), .Z(n3791) );
  XNOR U3992 ( .A(n3799), .B(n4017), .Z(n3792) );
  XNOR U3993 ( .A(n3798), .B(n3796), .Z(n4017) );
  AND U3994 ( .A(n4018), .B(n4019), .Z(n3796) );
  NANDN U3995 ( .A(n4020), .B(n4021), .Z(n4019) );
  OR U3996 ( .A(n4022), .B(n4023), .Z(n4021) );
  NAND U3997 ( .A(n4023), .B(n4022), .Z(n4018) );
  ANDN U3998 ( .B(B[53]), .A(n67), .Z(n3798) );
  XNOR U3999 ( .A(n3806), .B(n4024), .Z(n3799) );
  XNOR U4000 ( .A(n3805), .B(n3803), .Z(n4024) );
  AND U4001 ( .A(n4025), .B(n4026), .Z(n3803) );
  NANDN U4002 ( .A(n4027), .B(n4028), .Z(n4026) );
  NANDN U4003 ( .A(n4029), .B(n4030), .Z(n4028) );
  NANDN U4004 ( .A(n4030), .B(n4029), .Z(n4025) );
  ANDN U4005 ( .B(B[54]), .A(n68), .Z(n3805) );
  XNOR U4006 ( .A(n3813), .B(n4031), .Z(n3806) );
  XNOR U4007 ( .A(n3812), .B(n3810), .Z(n4031) );
  AND U4008 ( .A(n4032), .B(n4033), .Z(n3810) );
  NANDN U4009 ( .A(n4034), .B(n4035), .Z(n4033) );
  OR U4010 ( .A(n4036), .B(n4037), .Z(n4035) );
  NAND U4011 ( .A(n4037), .B(n4036), .Z(n4032) );
  ANDN U4012 ( .B(B[55]), .A(n69), .Z(n3812) );
  XNOR U4013 ( .A(n3820), .B(n4038), .Z(n3813) );
  XNOR U4014 ( .A(n3819), .B(n3817), .Z(n4038) );
  AND U4015 ( .A(n4039), .B(n4040), .Z(n3817) );
  NANDN U4016 ( .A(n4041), .B(n4042), .Z(n4040) );
  NANDN U4017 ( .A(n4043), .B(n4044), .Z(n4042) );
  NANDN U4018 ( .A(n4044), .B(n4043), .Z(n4039) );
  ANDN U4019 ( .B(B[56]), .A(n70), .Z(n3819) );
  XNOR U4020 ( .A(n3827), .B(n4045), .Z(n3820) );
  XNOR U4021 ( .A(n3826), .B(n3824), .Z(n4045) );
  AND U4022 ( .A(n4046), .B(n4047), .Z(n3824) );
  NANDN U4023 ( .A(n4048), .B(n4049), .Z(n4047) );
  OR U4024 ( .A(n4050), .B(n4051), .Z(n4049) );
  NAND U4025 ( .A(n4051), .B(n4050), .Z(n4046) );
  ANDN U4026 ( .B(B[57]), .A(n71), .Z(n3826) );
  XNOR U4027 ( .A(n3834), .B(n4052), .Z(n3827) );
  XNOR U4028 ( .A(n3833), .B(n3831), .Z(n4052) );
  AND U4029 ( .A(n4053), .B(n4054), .Z(n3831) );
  NANDN U4030 ( .A(n4055), .B(n4056), .Z(n4054) );
  NANDN U4031 ( .A(n4057), .B(n4058), .Z(n4056) );
  NANDN U4032 ( .A(n4058), .B(n4057), .Z(n4053) );
  ANDN U4033 ( .B(B[58]), .A(n72), .Z(n3833) );
  XNOR U4034 ( .A(n3841), .B(n4059), .Z(n3834) );
  XNOR U4035 ( .A(n3840), .B(n3838), .Z(n4059) );
  AND U4036 ( .A(n4060), .B(n4061), .Z(n3838) );
  NANDN U4037 ( .A(n4062), .B(n4063), .Z(n4061) );
  OR U4038 ( .A(n4064), .B(n4065), .Z(n4063) );
  NAND U4039 ( .A(n4065), .B(n4064), .Z(n4060) );
  ANDN U4040 ( .B(B[59]), .A(n73), .Z(n3840) );
  XNOR U4041 ( .A(n3848), .B(n4066), .Z(n3841) );
  XNOR U4042 ( .A(n3847), .B(n3845), .Z(n4066) );
  AND U4043 ( .A(n4067), .B(n4068), .Z(n3845) );
  NANDN U4044 ( .A(n4069), .B(n4070), .Z(n4068) );
  NANDN U4045 ( .A(n4071), .B(n4072), .Z(n4070) );
  NANDN U4046 ( .A(n4072), .B(n4071), .Z(n4067) );
  ANDN U4047 ( .B(B[60]), .A(n74), .Z(n3847) );
  XNOR U4048 ( .A(n3855), .B(n4073), .Z(n3848) );
  XNOR U4049 ( .A(n3854), .B(n3852), .Z(n4073) );
  AND U4050 ( .A(n4074), .B(n4075), .Z(n3852) );
  NANDN U4051 ( .A(n4076), .B(n4077), .Z(n4075) );
  OR U4052 ( .A(n4078), .B(n4079), .Z(n4077) );
  NAND U4053 ( .A(n4079), .B(n4078), .Z(n4074) );
  ANDN U4054 ( .B(B[61]), .A(n75), .Z(n3854) );
  XNOR U4055 ( .A(n3862), .B(n4080), .Z(n3855) );
  XNOR U4056 ( .A(n3861), .B(n3859), .Z(n4080) );
  AND U4057 ( .A(n4081), .B(n4082), .Z(n3859) );
  NANDN U4058 ( .A(n4083), .B(n4084), .Z(n4082) );
  NANDN U4059 ( .A(n4085), .B(n4086), .Z(n4084) );
  NANDN U4060 ( .A(n4086), .B(n4085), .Z(n4081) );
  ANDN U4061 ( .B(B[62]), .A(n76), .Z(n3861) );
  XNOR U4062 ( .A(n3869), .B(n4087), .Z(n3862) );
  XNOR U4063 ( .A(n3868), .B(n3866), .Z(n4087) );
  AND U4064 ( .A(n4088), .B(n4089), .Z(n3866) );
  NANDN U4065 ( .A(n4090), .B(n4091), .Z(n4089) );
  OR U4066 ( .A(n4092), .B(n4093), .Z(n4091) );
  NAND U4067 ( .A(n4093), .B(n4092), .Z(n4088) );
  ANDN U4068 ( .B(B[63]), .A(n77), .Z(n3868) );
  XNOR U4069 ( .A(n3876), .B(n4094), .Z(n3869) );
  XNOR U4070 ( .A(n3875), .B(n3873), .Z(n4094) );
  AND U4071 ( .A(n4095), .B(n4096), .Z(n3873) );
  NANDN U4072 ( .A(n4097), .B(n4098), .Z(n4096) );
  NANDN U4073 ( .A(n4099), .B(n4100), .Z(n4098) );
  NANDN U4074 ( .A(n4100), .B(n4099), .Z(n4095) );
  ANDN U4075 ( .B(B[64]), .A(n78), .Z(n3875) );
  XNOR U4076 ( .A(n3883), .B(n4101), .Z(n3876) );
  XNOR U4077 ( .A(n3882), .B(n3880), .Z(n4101) );
  AND U4078 ( .A(n4102), .B(n4103), .Z(n3880) );
  NANDN U4079 ( .A(n4104), .B(n4105), .Z(n4103) );
  OR U4080 ( .A(n4106), .B(n4107), .Z(n4105) );
  NAND U4081 ( .A(n4107), .B(n4106), .Z(n4102) );
  ANDN U4082 ( .B(B[65]), .A(n79), .Z(n3882) );
  XNOR U4083 ( .A(n3890), .B(n4108), .Z(n3883) );
  XNOR U4084 ( .A(n3889), .B(n3887), .Z(n4108) );
  AND U4085 ( .A(n4109), .B(n4110), .Z(n3887) );
  NANDN U4086 ( .A(n4111), .B(n4112), .Z(n4110) );
  NANDN U4087 ( .A(n4113), .B(n4114), .Z(n4112) );
  NANDN U4088 ( .A(n4114), .B(n4113), .Z(n4109) );
  ANDN U4089 ( .B(B[66]), .A(n80), .Z(n3889) );
  XNOR U4090 ( .A(n3897), .B(n4115), .Z(n3890) );
  XNOR U4091 ( .A(n3896), .B(n3894), .Z(n4115) );
  AND U4092 ( .A(n4116), .B(n4117), .Z(n3894) );
  NANDN U4093 ( .A(n4118), .B(n4119), .Z(n4117) );
  OR U4094 ( .A(n4120), .B(n4121), .Z(n4119) );
  NAND U4095 ( .A(n4121), .B(n4120), .Z(n4116) );
  ANDN U4096 ( .B(B[67]), .A(n81), .Z(n3896) );
  XNOR U4097 ( .A(n48), .B(n4122), .Z(n3897) );
  XNOR U4098 ( .A(n3903), .B(n3901), .Z(n4122) );
  AND U4099 ( .A(n4123), .B(n4124), .Z(n3901) );
  NANDN U4100 ( .A(n4125), .B(n4126), .Z(n4124) );
  NAND U4101 ( .A(n4127), .B(n4128), .Z(n4126) );
  ANDN U4102 ( .B(B[68]), .A(n82), .Z(n3903) );
  XNOR U4103 ( .A(n3908), .B(n4129), .Z(n3904) );
  XOR U4104 ( .A(n3910), .B(n3911), .Z(n4129) );
  NAND U4105 ( .A(B[69]), .B(A[2]), .Z(n3911) );
  ANDN U4106 ( .B(n4130), .A(n4131), .Z(n3910) );
  AND U4107 ( .A(A[0]), .B(B[70]), .Z(n4130) );
  XNOR U4108 ( .A(n4132), .B(n4133), .Z(n3908) );
  NAND U4109 ( .A(B[71]), .B(A[0]), .Z(n4133) );
  NAND U4110 ( .A(n4134), .B(n4135), .Z(n145) );
  NANDN U4111 ( .A(n4136), .B(n4137), .Z(n4135) );
  OR U4112 ( .A(n4138), .B(n4139), .Z(n4137) );
  NAND U4113 ( .A(n4139), .B(n4138), .Z(n4134) );
  XOR U4114 ( .A(n147), .B(n146), .Z(\A1[68] ) );
  XOR U4115 ( .A(n4139), .B(n4140), .Z(n146) );
  XNOR U4116 ( .A(n4138), .B(n4136), .Z(n4140) );
  AND U4117 ( .A(n4141), .B(n4142), .Z(n4136) );
  NANDN U4118 ( .A(n4143), .B(n4144), .Z(n4142) );
  NANDN U4119 ( .A(n4145), .B(n4146), .Z(n4144) );
  NANDN U4120 ( .A(n4146), .B(n4145), .Z(n4141) );
  ANDN U4121 ( .B(B[39]), .A(n54), .Z(n4138) );
  XNOR U4122 ( .A(n3932), .B(n4147), .Z(n4139) );
  XNOR U4123 ( .A(n3931), .B(n3929), .Z(n4147) );
  AND U4124 ( .A(n4148), .B(n4149), .Z(n3929) );
  NANDN U4125 ( .A(n4150), .B(n4151), .Z(n4149) );
  OR U4126 ( .A(n4152), .B(n4153), .Z(n4151) );
  NAND U4127 ( .A(n4153), .B(n4152), .Z(n4148) );
  ANDN U4128 ( .B(B[40]), .A(n55), .Z(n3931) );
  XNOR U4129 ( .A(n3939), .B(n4154), .Z(n3932) );
  XNOR U4130 ( .A(n3938), .B(n3936), .Z(n4154) );
  AND U4131 ( .A(n4155), .B(n4156), .Z(n3936) );
  NANDN U4132 ( .A(n4157), .B(n4158), .Z(n4156) );
  NANDN U4133 ( .A(n4159), .B(n4160), .Z(n4158) );
  NANDN U4134 ( .A(n4160), .B(n4159), .Z(n4155) );
  ANDN U4135 ( .B(B[41]), .A(n56), .Z(n3938) );
  XNOR U4136 ( .A(n3946), .B(n4161), .Z(n3939) );
  XNOR U4137 ( .A(n3945), .B(n3943), .Z(n4161) );
  AND U4138 ( .A(n4162), .B(n4163), .Z(n3943) );
  NANDN U4139 ( .A(n4164), .B(n4165), .Z(n4163) );
  OR U4140 ( .A(n4166), .B(n4167), .Z(n4165) );
  NAND U4141 ( .A(n4167), .B(n4166), .Z(n4162) );
  ANDN U4142 ( .B(B[42]), .A(n57), .Z(n3945) );
  XNOR U4143 ( .A(n3953), .B(n4168), .Z(n3946) );
  XNOR U4144 ( .A(n3952), .B(n3950), .Z(n4168) );
  AND U4145 ( .A(n4169), .B(n4170), .Z(n3950) );
  NANDN U4146 ( .A(n4171), .B(n4172), .Z(n4170) );
  NANDN U4147 ( .A(n4173), .B(n4174), .Z(n4172) );
  NANDN U4148 ( .A(n4174), .B(n4173), .Z(n4169) );
  ANDN U4149 ( .B(B[43]), .A(n58), .Z(n3952) );
  XNOR U4150 ( .A(n3960), .B(n4175), .Z(n3953) );
  XNOR U4151 ( .A(n3959), .B(n3957), .Z(n4175) );
  AND U4152 ( .A(n4176), .B(n4177), .Z(n3957) );
  NANDN U4153 ( .A(n4178), .B(n4179), .Z(n4177) );
  OR U4154 ( .A(n4180), .B(n4181), .Z(n4179) );
  NAND U4155 ( .A(n4181), .B(n4180), .Z(n4176) );
  ANDN U4156 ( .B(B[44]), .A(n59), .Z(n3959) );
  XNOR U4157 ( .A(n3967), .B(n4182), .Z(n3960) );
  XNOR U4158 ( .A(n3966), .B(n3964), .Z(n4182) );
  AND U4159 ( .A(n4183), .B(n4184), .Z(n3964) );
  NANDN U4160 ( .A(n4185), .B(n4186), .Z(n4184) );
  NANDN U4161 ( .A(n4187), .B(n4188), .Z(n4186) );
  NANDN U4162 ( .A(n4188), .B(n4187), .Z(n4183) );
  ANDN U4163 ( .B(B[45]), .A(n60), .Z(n3966) );
  XNOR U4164 ( .A(n3974), .B(n4189), .Z(n3967) );
  XNOR U4165 ( .A(n3973), .B(n3971), .Z(n4189) );
  AND U4166 ( .A(n4190), .B(n4191), .Z(n3971) );
  NANDN U4167 ( .A(n4192), .B(n4193), .Z(n4191) );
  OR U4168 ( .A(n4194), .B(n4195), .Z(n4193) );
  NAND U4169 ( .A(n4195), .B(n4194), .Z(n4190) );
  ANDN U4170 ( .B(B[46]), .A(n61), .Z(n3973) );
  XNOR U4171 ( .A(n3981), .B(n4196), .Z(n3974) );
  XNOR U4172 ( .A(n3980), .B(n3978), .Z(n4196) );
  AND U4173 ( .A(n4197), .B(n4198), .Z(n3978) );
  NANDN U4174 ( .A(n4199), .B(n4200), .Z(n4198) );
  NANDN U4175 ( .A(n4201), .B(n4202), .Z(n4200) );
  NANDN U4176 ( .A(n4202), .B(n4201), .Z(n4197) );
  ANDN U4177 ( .B(B[47]), .A(n62), .Z(n3980) );
  XNOR U4178 ( .A(n3988), .B(n4203), .Z(n3981) );
  XNOR U4179 ( .A(n3987), .B(n3985), .Z(n4203) );
  AND U4180 ( .A(n4204), .B(n4205), .Z(n3985) );
  NANDN U4181 ( .A(n4206), .B(n4207), .Z(n4205) );
  OR U4182 ( .A(n4208), .B(n4209), .Z(n4207) );
  NAND U4183 ( .A(n4209), .B(n4208), .Z(n4204) );
  ANDN U4184 ( .B(B[48]), .A(n63), .Z(n3987) );
  XNOR U4185 ( .A(n3995), .B(n4210), .Z(n3988) );
  XNOR U4186 ( .A(n3994), .B(n3992), .Z(n4210) );
  AND U4187 ( .A(n4211), .B(n4212), .Z(n3992) );
  NANDN U4188 ( .A(n4213), .B(n4214), .Z(n4212) );
  NANDN U4189 ( .A(n4215), .B(n4216), .Z(n4214) );
  NANDN U4190 ( .A(n4216), .B(n4215), .Z(n4211) );
  ANDN U4191 ( .B(B[49]), .A(n64), .Z(n3994) );
  XNOR U4192 ( .A(n4002), .B(n4217), .Z(n3995) );
  XNOR U4193 ( .A(n4001), .B(n3999), .Z(n4217) );
  AND U4194 ( .A(n4218), .B(n4219), .Z(n3999) );
  NANDN U4195 ( .A(n4220), .B(n4221), .Z(n4219) );
  OR U4196 ( .A(n4222), .B(n4223), .Z(n4221) );
  NAND U4197 ( .A(n4223), .B(n4222), .Z(n4218) );
  ANDN U4198 ( .B(B[50]), .A(n65), .Z(n4001) );
  XNOR U4199 ( .A(n4009), .B(n4224), .Z(n4002) );
  XNOR U4200 ( .A(n4008), .B(n4006), .Z(n4224) );
  AND U4201 ( .A(n4225), .B(n4226), .Z(n4006) );
  NANDN U4202 ( .A(n4227), .B(n4228), .Z(n4226) );
  NANDN U4203 ( .A(n4229), .B(n4230), .Z(n4228) );
  NANDN U4204 ( .A(n4230), .B(n4229), .Z(n4225) );
  ANDN U4205 ( .B(B[51]), .A(n66), .Z(n4008) );
  XNOR U4206 ( .A(n4016), .B(n4231), .Z(n4009) );
  XNOR U4207 ( .A(n4015), .B(n4013), .Z(n4231) );
  AND U4208 ( .A(n4232), .B(n4233), .Z(n4013) );
  NANDN U4209 ( .A(n4234), .B(n4235), .Z(n4233) );
  OR U4210 ( .A(n4236), .B(n4237), .Z(n4235) );
  NAND U4211 ( .A(n4237), .B(n4236), .Z(n4232) );
  ANDN U4212 ( .B(B[52]), .A(n67), .Z(n4015) );
  XNOR U4213 ( .A(n4023), .B(n4238), .Z(n4016) );
  XNOR U4214 ( .A(n4022), .B(n4020), .Z(n4238) );
  AND U4215 ( .A(n4239), .B(n4240), .Z(n4020) );
  NANDN U4216 ( .A(n4241), .B(n4242), .Z(n4240) );
  NANDN U4217 ( .A(n4243), .B(n4244), .Z(n4242) );
  NANDN U4218 ( .A(n4244), .B(n4243), .Z(n4239) );
  ANDN U4219 ( .B(B[53]), .A(n68), .Z(n4022) );
  XNOR U4220 ( .A(n4030), .B(n4245), .Z(n4023) );
  XNOR U4221 ( .A(n4029), .B(n4027), .Z(n4245) );
  AND U4222 ( .A(n4246), .B(n4247), .Z(n4027) );
  NANDN U4223 ( .A(n4248), .B(n4249), .Z(n4247) );
  OR U4224 ( .A(n4250), .B(n4251), .Z(n4249) );
  NAND U4225 ( .A(n4251), .B(n4250), .Z(n4246) );
  ANDN U4226 ( .B(B[54]), .A(n69), .Z(n4029) );
  XNOR U4227 ( .A(n4037), .B(n4252), .Z(n4030) );
  XNOR U4228 ( .A(n4036), .B(n4034), .Z(n4252) );
  AND U4229 ( .A(n4253), .B(n4254), .Z(n4034) );
  NANDN U4230 ( .A(n4255), .B(n4256), .Z(n4254) );
  NANDN U4231 ( .A(n4257), .B(n4258), .Z(n4256) );
  NANDN U4232 ( .A(n4258), .B(n4257), .Z(n4253) );
  ANDN U4233 ( .B(B[55]), .A(n70), .Z(n4036) );
  XNOR U4234 ( .A(n4044), .B(n4259), .Z(n4037) );
  XNOR U4235 ( .A(n4043), .B(n4041), .Z(n4259) );
  AND U4236 ( .A(n4260), .B(n4261), .Z(n4041) );
  NANDN U4237 ( .A(n4262), .B(n4263), .Z(n4261) );
  OR U4238 ( .A(n4264), .B(n4265), .Z(n4263) );
  NAND U4239 ( .A(n4265), .B(n4264), .Z(n4260) );
  ANDN U4240 ( .B(B[56]), .A(n71), .Z(n4043) );
  XNOR U4241 ( .A(n4051), .B(n4266), .Z(n4044) );
  XNOR U4242 ( .A(n4050), .B(n4048), .Z(n4266) );
  AND U4243 ( .A(n4267), .B(n4268), .Z(n4048) );
  NANDN U4244 ( .A(n4269), .B(n4270), .Z(n4268) );
  NANDN U4245 ( .A(n4271), .B(n4272), .Z(n4270) );
  NANDN U4246 ( .A(n4272), .B(n4271), .Z(n4267) );
  ANDN U4247 ( .B(B[57]), .A(n72), .Z(n4050) );
  XNOR U4248 ( .A(n4058), .B(n4273), .Z(n4051) );
  XNOR U4249 ( .A(n4057), .B(n4055), .Z(n4273) );
  AND U4250 ( .A(n4274), .B(n4275), .Z(n4055) );
  NANDN U4251 ( .A(n4276), .B(n4277), .Z(n4275) );
  OR U4252 ( .A(n4278), .B(n4279), .Z(n4277) );
  NAND U4253 ( .A(n4279), .B(n4278), .Z(n4274) );
  ANDN U4254 ( .B(B[58]), .A(n73), .Z(n4057) );
  XNOR U4255 ( .A(n4065), .B(n4280), .Z(n4058) );
  XNOR U4256 ( .A(n4064), .B(n4062), .Z(n4280) );
  AND U4257 ( .A(n4281), .B(n4282), .Z(n4062) );
  NANDN U4258 ( .A(n4283), .B(n4284), .Z(n4282) );
  NANDN U4259 ( .A(n4285), .B(n4286), .Z(n4284) );
  NANDN U4260 ( .A(n4286), .B(n4285), .Z(n4281) );
  ANDN U4261 ( .B(B[59]), .A(n74), .Z(n4064) );
  XNOR U4262 ( .A(n4072), .B(n4287), .Z(n4065) );
  XNOR U4263 ( .A(n4071), .B(n4069), .Z(n4287) );
  AND U4264 ( .A(n4288), .B(n4289), .Z(n4069) );
  NANDN U4265 ( .A(n4290), .B(n4291), .Z(n4289) );
  OR U4266 ( .A(n4292), .B(n4293), .Z(n4291) );
  NAND U4267 ( .A(n4293), .B(n4292), .Z(n4288) );
  ANDN U4268 ( .B(B[60]), .A(n75), .Z(n4071) );
  XNOR U4269 ( .A(n4079), .B(n4294), .Z(n4072) );
  XNOR U4270 ( .A(n4078), .B(n4076), .Z(n4294) );
  AND U4271 ( .A(n4295), .B(n4296), .Z(n4076) );
  NANDN U4272 ( .A(n4297), .B(n4298), .Z(n4296) );
  NANDN U4273 ( .A(n4299), .B(n4300), .Z(n4298) );
  NANDN U4274 ( .A(n4300), .B(n4299), .Z(n4295) );
  ANDN U4275 ( .B(B[61]), .A(n76), .Z(n4078) );
  XNOR U4276 ( .A(n4086), .B(n4301), .Z(n4079) );
  XNOR U4277 ( .A(n4085), .B(n4083), .Z(n4301) );
  AND U4278 ( .A(n4302), .B(n4303), .Z(n4083) );
  NANDN U4279 ( .A(n4304), .B(n4305), .Z(n4303) );
  OR U4280 ( .A(n4306), .B(n4307), .Z(n4305) );
  NAND U4281 ( .A(n4307), .B(n4306), .Z(n4302) );
  ANDN U4282 ( .B(B[62]), .A(n77), .Z(n4085) );
  XNOR U4283 ( .A(n4093), .B(n4308), .Z(n4086) );
  XNOR U4284 ( .A(n4092), .B(n4090), .Z(n4308) );
  AND U4285 ( .A(n4309), .B(n4310), .Z(n4090) );
  NANDN U4286 ( .A(n4311), .B(n4312), .Z(n4310) );
  NANDN U4287 ( .A(n4313), .B(n4314), .Z(n4312) );
  NANDN U4288 ( .A(n4314), .B(n4313), .Z(n4309) );
  ANDN U4289 ( .B(B[63]), .A(n78), .Z(n4092) );
  XNOR U4290 ( .A(n4100), .B(n4315), .Z(n4093) );
  XNOR U4291 ( .A(n4099), .B(n4097), .Z(n4315) );
  AND U4292 ( .A(n4316), .B(n4317), .Z(n4097) );
  NANDN U4293 ( .A(n4318), .B(n4319), .Z(n4317) );
  OR U4294 ( .A(n4320), .B(n4321), .Z(n4319) );
  NAND U4295 ( .A(n4321), .B(n4320), .Z(n4316) );
  ANDN U4296 ( .B(B[64]), .A(n79), .Z(n4099) );
  XNOR U4297 ( .A(n4107), .B(n4322), .Z(n4100) );
  XNOR U4298 ( .A(n4106), .B(n4104), .Z(n4322) );
  AND U4299 ( .A(n4323), .B(n4324), .Z(n4104) );
  NANDN U4300 ( .A(n4325), .B(n4326), .Z(n4324) );
  NANDN U4301 ( .A(n4327), .B(n4328), .Z(n4326) );
  NANDN U4302 ( .A(n4328), .B(n4327), .Z(n4323) );
  ANDN U4303 ( .B(B[65]), .A(n80), .Z(n4106) );
  XNOR U4304 ( .A(n4114), .B(n4329), .Z(n4107) );
  XNOR U4305 ( .A(n4113), .B(n4111), .Z(n4329) );
  AND U4306 ( .A(n4330), .B(n4331), .Z(n4111) );
  NANDN U4307 ( .A(n4332), .B(n4333), .Z(n4331) );
  OR U4308 ( .A(n4334), .B(n4335), .Z(n4333) );
  NAND U4309 ( .A(n4335), .B(n4334), .Z(n4330) );
  ANDN U4310 ( .B(B[66]), .A(n81), .Z(n4113) );
  XNOR U4311 ( .A(n4121), .B(n4336), .Z(n4114) );
  XNOR U4312 ( .A(n4120), .B(n4118), .Z(n4336) );
  AND U4313 ( .A(n4337), .B(n4338), .Z(n4118) );
  NANDN U4314 ( .A(n4339), .B(n4340), .Z(n4338) );
  NAND U4315 ( .A(n4341), .B(n4342), .Z(n4340) );
  ANDN U4316 ( .B(B[67]), .A(n82), .Z(n4120) );
  XOR U4317 ( .A(n4127), .B(n4343), .Z(n4121) );
  XNOR U4318 ( .A(n4125), .B(n4128), .Z(n4343) );
  NAND U4319 ( .A(B[68]), .B(A[2]), .Z(n4128) );
  NAND U4320 ( .A(B[69]), .B(n4344), .Z(n4125) );
  ANDN U4321 ( .B(A[0]), .A(n4345), .Z(n4344) );
  XNOR U4322 ( .A(n4131), .B(n4346), .Z(n4127) );
  NAND U4323 ( .A(A[0]), .B(B[70]), .Z(n4346) );
  NAND U4324 ( .A(B[69]), .B(A[1]), .Z(n4131) );
  NAND U4325 ( .A(n4347), .B(n4348), .Z(n147) );
  NANDN U4326 ( .A(n4349), .B(n4350), .Z(n4348) );
  OR U4327 ( .A(n4351), .B(n4352), .Z(n4350) );
  NAND U4328 ( .A(n4352), .B(n4351), .Z(n4347) );
  XOR U4329 ( .A(n149), .B(n148), .Z(\A1[67] ) );
  XOR U4330 ( .A(n4352), .B(n4353), .Z(n148) );
  XNOR U4331 ( .A(n4351), .B(n4349), .Z(n4353) );
  AND U4332 ( .A(n4354), .B(n4355), .Z(n4349) );
  NANDN U4333 ( .A(n4356), .B(n4357), .Z(n4355) );
  NANDN U4334 ( .A(n4358), .B(n4359), .Z(n4357) );
  NANDN U4335 ( .A(n4359), .B(n4358), .Z(n4354) );
  ANDN U4336 ( .B(B[38]), .A(n54), .Z(n4351) );
  XNOR U4337 ( .A(n4146), .B(n4360), .Z(n4352) );
  XNOR U4338 ( .A(n4145), .B(n4143), .Z(n4360) );
  AND U4339 ( .A(n4361), .B(n4362), .Z(n4143) );
  NANDN U4340 ( .A(n4363), .B(n4364), .Z(n4362) );
  OR U4341 ( .A(n4365), .B(n4366), .Z(n4364) );
  NAND U4342 ( .A(n4366), .B(n4365), .Z(n4361) );
  ANDN U4343 ( .B(B[39]), .A(n55), .Z(n4145) );
  XNOR U4344 ( .A(n4153), .B(n4367), .Z(n4146) );
  XNOR U4345 ( .A(n4152), .B(n4150), .Z(n4367) );
  AND U4346 ( .A(n4368), .B(n4369), .Z(n4150) );
  NANDN U4347 ( .A(n4370), .B(n4371), .Z(n4369) );
  NANDN U4348 ( .A(n4372), .B(n4373), .Z(n4371) );
  NANDN U4349 ( .A(n4373), .B(n4372), .Z(n4368) );
  ANDN U4350 ( .B(B[40]), .A(n56), .Z(n4152) );
  XNOR U4351 ( .A(n4160), .B(n4374), .Z(n4153) );
  XNOR U4352 ( .A(n4159), .B(n4157), .Z(n4374) );
  AND U4353 ( .A(n4375), .B(n4376), .Z(n4157) );
  NANDN U4354 ( .A(n4377), .B(n4378), .Z(n4376) );
  OR U4355 ( .A(n4379), .B(n4380), .Z(n4378) );
  NAND U4356 ( .A(n4380), .B(n4379), .Z(n4375) );
  ANDN U4357 ( .B(B[41]), .A(n57), .Z(n4159) );
  XNOR U4358 ( .A(n4167), .B(n4381), .Z(n4160) );
  XNOR U4359 ( .A(n4166), .B(n4164), .Z(n4381) );
  AND U4360 ( .A(n4382), .B(n4383), .Z(n4164) );
  NANDN U4361 ( .A(n4384), .B(n4385), .Z(n4383) );
  NANDN U4362 ( .A(n4386), .B(n4387), .Z(n4385) );
  NANDN U4363 ( .A(n4387), .B(n4386), .Z(n4382) );
  ANDN U4364 ( .B(B[42]), .A(n58), .Z(n4166) );
  XNOR U4365 ( .A(n4174), .B(n4388), .Z(n4167) );
  XNOR U4366 ( .A(n4173), .B(n4171), .Z(n4388) );
  AND U4367 ( .A(n4389), .B(n4390), .Z(n4171) );
  NANDN U4368 ( .A(n4391), .B(n4392), .Z(n4390) );
  OR U4369 ( .A(n4393), .B(n4394), .Z(n4392) );
  NAND U4370 ( .A(n4394), .B(n4393), .Z(n4389) );
  ANDN U4371 ( .B(B[43]), .A(n59), .Z(n4173) );
  XNOR U4372 ( .A(n4181), .B(n4395), .Z(n4174) );
  XNOR U4373 ( .A(n4180), .B(n4178), .Z(n4395) );
  AND U4374 ( .A(n4396), .B(n4397), .Z(n4178) );
  NANDN U4375 ( .A(n4398), .B(n4399), .Z(n4397) );
  NANDN U4376 ( .A(n4400), .B(n4401), .Z(n4399) );
  NANDN U4377 ( .A(n4401), .B(n4400), .Z(n4396) );
  ANDN U4378 ( .B(B[44]), .A(n60), .Z(n4180) );
  XNOR U4379 ( .A(n4188), .B(n4402), .Z(n4181) );
  XNOR U4380 ( .A(n4187), .B(n4185), .Z(n4402) );
  AND U4381 ( .A(n4403), .B(n4404), .Z(n4185) );
  NANDN U4382 ( .A(n4405), .B(n4406), .Z(n4404) );
  OR U4383 ( .A(n4407), .B(n4408), .Z(n4406) );
  NAND U4384 ( .A(n4408), .B(n4407), .Z(n4403) );
  ANDN U4385 ( .B(B[45]), .A(n61), .Z(n4187) );
  XNOR U4386 ( .A(n4195), .B(n4409), .Z(n4188) );
  XNOR U4387 ( .A(n4194), .B(n4192), .Z(n4409) );
  AND U4388 ( .A(n4410), .B(n4411), .Z(n4192) );
  NANDN U4389 ( .A(n4412), .B(n4413), .Z(n4411) );
  NANDN U4390 ( .A(n4414), .B(n4415), .Z(n4413) );
  NANDN U4391 ( .A(n4415), .B(n4414), .Z(n4410) );
  ANDN U4392 ( .B(B[46]), .A(n62), .Z(n4194) );
  XNOR U4393 ( .A(n4202), .B(n4416), .Z(n4195) );
  XNOR U4394 ( .A(n4201), .B(n4199), .Z(n4416) );
  AND U4395 ( .A(n4417), .B(n4418), .Z(n4199) );
  NANDN U4396 ( .A(n4419), .B(n4420), .Z(n4418) );
  OR U4397 ( .A(n4421), .B(n4422), .Z(n4420) );
  NAND U4398 ( .A(n4422), .B(n4421), .Z(n4417) );
  ANDN U4399 ( .B(B[47]), .A(n63), .Z(n4201) );
  XNOR U4400 ( .A(n4209), .B(n4423), .Z(n4202) );
  XNOR U4401 ( .A(n4208), .B(n4206), .Z(n4423) );
  AND U4402 ( .A(n4424), .B(n4425), .Z(n4206) );
  NANDN U4403 ( .A(n4426), .B(n4427), .Z(n4425) );
  NANDN U4404 ( .A(n4428), .B(n4429), .Z(n4427) );
  NANDN U4405 ( .A(n4429), .B(n4428), .Z(n4424) );
  ANDN U4406 ( .B(B[48]), .A(n64), .Z(n4208) );
  XNOR U4407 ( .A(n4216), .B(n4430), .Z(n4209) );
  XNOR U4408 ( .A(n4215), .B(n4213), .Z(n4430) );
  AND U4409 ( .A(n4431), .B(n4432), .Z(n4213) );
  NANDN U4410 ( .A(n4433), .B(n4434), .Z(n4432) );
  OR U4411 ( .A(n4435), .B(n4436), .Z(n4434) );
  NAND U4412 ( .A(n4436), .B(n4435), .Z(n4431) );
  ANDN U4413 ( .B(B[49]), .A(n65), .Z(n4215) );
  XNOR U4414 ( .A(n4223), .B(n4437), .Z(n4216) );
  XNOR U4415 ( .A(n4222), .B(n4220), .Z(n4437) );
  AND U4416 ( .A(n4438), .B(n4439), .Z(n4220) );
  NANDN U4417 ( .A(n4440), .B(n4441), .Z(n4439) );
  NANDN U4418 ( .A(n4442), .B(n4443), .Z(n4441) );
  NANDN U4419 ( .A(n4443), .B(n4442), .Z(n4438) );
  ANDN U4420 ( .B(B[50]), .A(n66), .Z(n4222) );
  XNOR U4421 ( .A(n4230), .B(n4444), .Z(n4223) );
  XNOR U4422 ( .A(n4229), .B(n4227), .Z(n4444) );
  AND U4423 ( .A(n4445), .B(n4446), .Z(n4227) );
  NANDN U4424 ( .A(n4447), .B(n4448), .Z(n4446) );
  OR U4425 ( .A(n4449), .B(n4450), .Z(n4448) );
  NAND U4426 ( .A(n4450), .B(n4449), .Z(n4445) );
  ANDN U4427 ( .B(B[51]), .A(n67), .Z(n4229) );
  XNOR U4428 ( .A(n4237), .B(n4451), .Z(n4230) );
  XNOR U4429 ( .A(n4236), .B(n4234), .Z(n4451) );
  AND U4430 ( .A(n4452), .B(n4453), .Z(n4234) );
  NANDN U4431 ( .A(n4454), .B(n4455), .Z(n4453) );
  NANDN U4432 ( .A(n4456), .B(n4457), .Z(n4455) );
  NANDN U4433 ( .A(n4457), .B(n4456), .Z(n4452) );
  ANDN U4434 ( .B(B[52]), .A(n68), .Z(n4236) );
  XNOR U4435 ( .A(n4244), .B(n4458), .Z(n4237) );
  XNOR U4436 ( .A(n4243), .B(n4241), .Z(n4458) );
  AND U4437 ( .A(n4459), .B(n4460), .Z(n4241) );
  NANDN U4438 ( .A(n4461), .B(n4462), .Z(n4460) );
  OR U4439 ( .A(n4463), .B(n4464), .Z(n4462) );
  NAND U4440 ( .A(n4464), .B(n4463), .Z(n4459) );
  ANDN U4441 ( .B(B[53]), .A(n69), .Z(n4243) );
  XNOR U4442 ( .A(n4251), .B(n4465), .Z(n4244) );
  XNOR U4443 ( .A(n4250), .B(n4248), .Z(n4465) );
  AND U4444 ( .A(n4466), .B(n4467), .Z(n4248) );
  NANDN U4445 ( .A(n4468), .B(n4469), .Z(n4467) );
  NANDN U4446 ( .A(n4470), .B(n4471), .Z(n4469) );
  NANDN U4447 ( .A(n4471), .B(n4470), .Z(n4466) );
  ANDN U4448 ( .B(B[54]), .A(n70), .Z(n4250) );
  XNOR U4449 ( .A(n4258), .B(n4472), .Z(n4251) );
  XNOR U4450 ( .A(n4257), .B(n4255), .Z(n4472) );
  AND U4451 ( .A(n4473), .B(n4474), .Z(n4255) );
  NANDN U4452 ( .A(n4475), .B(n4476), .Z(n4474) );
  OR U4453 ( .A(n4477), .B(n4478), .Z(n4476) );
  NAND U4454 ( .A(n4478), .B(n4477), .Z(n4473) );
  ANDN U4455 ( .B(B[55]), .A(n71), .Z(n4257) );
  XNOR U4456 ( .A(n4265), .B(n4479), .Z(n4258) );
  XNOR U4457 ( .A(n4264), .B(n4262), .Z(n4479) );
  AND U4458 ( .A(n4480), .B(n4481), .Z(n4262) );
  NANDN U4459 ( .A(n4482), .B(n4483), .Z(n4481) );
  NANDN U4460 ( .A(n4484), .B(n4485), .Z(n4483) );
  NANDN U4461 ( .A(n4485), .B(n4484), .Z(n4480) );
  ANDN U4462 ( .B(B[56]), .A(n72), .Z(n4264) );
  XNOR U4463 ( .A(n4272), .B(n4486), .Z(n4265) );
  XNOR U4464 ( .A(n4271), .B(n4269), .Z(n4486) );
  AND U4465 ( .A(n4487), .B(n4488), .Z(n4269) );
  NANDN U4466 ( .A(n4489), .B(n4490), .Z(n4488) );
  OR U4467 ( .A(n4491), .B(n4492), .Z(n4490) );
  NAND U4468 ( .A(n4492), .B(n4491), .Z(n4487) );
  ANDN U4469 ( .B(B[57]), .A(n73), .Z(n4271) );
  XNOR U4470 ( .A(n4279), .B(n4493), .Z(n4272) );
  XNOR U4471 ( .A(n4278), .B(n4276), .Z(n4493) );
  AND U4472 ( .A(n4494), .B(n4495), .Z(n4276) );
  NANDN U4473 ( .A(n4496), .B(n4497), .Z(n4495) );
  NANDN U4474 ( .A(n4498), .B(n4499), .Z(n4497) );
  NANDN U4475 ( .A(n4499), .B(n4498), .Z(n4494) );
  ANDN U4476 ( .B(B[58]), .A(n74), .Z(n4278) );
  XNOR U4477 ( .A(n4286), .B(n4500), .Z(n4279) );
  XNOR U4478 ( .A(n4285), .B(n4283), .Z(n4500) );
  AND U4479 ( .A(n4501), .B(n4502), .Z(n4283) );
  NANDN U4480 ( .A(n4503), .B(n4504), .Z(n4502) );
  OR U4481 ( .A(n4505), .B(n4506), .Z(n4504) );
  NAND U4482 ( .A(n4506), .B(n4505), .Z(n4501) );
  ANDN U4483 ( .B(B[59]), .A(n75), .Z(n4285) );
  XNOR U4484 ( .A(n4293), .B(n4507), .Z(n4286) );
  XNOR U4485 ( .A(n4292), .B(n4290), .Z(n4507) );
  AND U4486 ( .A(n4508), .B(n4509), .Z(n4290) );
  NANDN U4487 ( .A(n4510), .B(n4511), .Z(n4509) );
  NANDN U4488 ( .A(n4512), .B(n4513), .Z(n4511) );
  NANDN U4489 ( .A(n4513), .B(n4512), .Z(n4508) );
  ANDN U4490 ( .B(B[60]), .A(n76), .Z(n4292) );
  XNOR U4491 ( .A(n4300), .B(n4514), .Z(n4293) );
  XNOR U4492 ( .A(n4299), .B(n4297), .Z(n4514) );
  AND U4493 ( .A(n4515), .B(n4516), .Z(n4297) );
  NANDN U4494 ( .A(n4517), .B(n4518), .Z(n4516) );
  OR U4495 ( .A(n4519), .B(n4520), .Z(n4518) );
  NAND U4496 ( .A(n4520), .B(n4519), .Z(n4515) );
  ANDN U4497 ( .B(B[61]), .A(n77), .Z(n4299) );
  XNOR U4498 ( .A(n4307), .B(n4521), .Z(n4300) );
  XNOR U4499 ( .A(n4306), .B(n4304), .Z(n4521) );
  AND U4500 ( .A(n4522), .B(n4523), .Z(n4304) );
  NANDN U4501 ( .A(n4524), .B(n4525), .Z(n4523) );
  NANDN U4502 ( .A(n4526), .B(n4527), .Z(n4525) );
  NANDN U4503 ( .A(n4527), .B(n4526), .Z(n4522) );
  ANDN U4504 ( .B(B[62]), .A(n78), .Z(n4306) );
  XNOR U4505 ( .A(n4314), .B(n4528), .Z(n4307) );
  XNOR U4506 ( .A(n4313), .B(n4311), .Z(n4528) );
  AND U4507 ( .A(n4529), .B(n4530), .Z(n4311) );
  NANDN U4508 ( .A(n4531), .B(n4532), .Z(n4530) );
  OR U4509 ( .A(n4533), .B(n4534), .Z(n4532) );
  NAND U4510 ( .A(n4534), .B(n4533), .Z(n4529) );
  ANDN U4511 ( .B(B[63]), .A(n79), .Z(n4313) );
  XNOR U4512 ( .A(n4321), .B(n4535), .Z(n4314) );
  XNOR U4513 ( .A(n4320), .B(n4318), .Z(n4535) );
  AND U4514 ( .A(n4536), .B(n4537), .Z(n4318) );
  NANDN U4515 ( .A(n4538), .B(n4539), .Z(n4537) );
  NANDN U4516 ( .A(n4540), .B(n4541), .Z(n4539) );
  NANDN U4517 ( .A(n4541), .B(n4540), .Z(n4536) );
  ANDN U4518 ( .B(B[64]), .A(n80), .Z(n4320) );
  XNOR U4519 ( .A(n4328), .B(n4542), .Z(n4321) );
  XNOR U4520 ( .A(n4327), .B(n4325), .Z(n4542) );
  AND U4521 ( .A(n4543), .B(n4544), .Z(n4325) );
  NANDN U4522 ( .A(n4545), .B(n4546), .Z(n4544) );
  OR U4523 ( .A(n4547), .B(n4548), .Z(n4546) );
  NAND U4524 ( .A(n4548), .B(n4547), .Z(n4543) );
  ANDN U4525 ( .B(B[65]), .A(n81), .Z(n4327) );
  XNOR U4526 ( .A(n4335), .B(n4549), .Z(n4328) );
  XNOR U4527 ( .A(n4334), .B(n4332), .Z(n4549) );
  AND U4528 ( .A(n4550), .B(n4551), .Z(n4332) );
  NANDN U4529 ( .A(n4552), .B(n4553), .Z(n4551) );
  NAND U4530 ( .A(n4554), .B(n4555), .Z(n4553) );
  ANDN U4531 ( .B(B[66]), .A(n82), .Z(n4334) );
  XOR U4532 ( .A(n4341), .B(n4556), .Z(n4335) );
  XNOR U4533 ( .A(n4339), .B(n4342), .Z(n4556) );
  NAND U4534 ( .A(A[2]), .B(B[67]), .Z(n4342) );
  NANDN U4535 ( .A(n4557), .B(n4558), .Z(n4339) );
  AND U4536 ( .A(A[0]), .B(B[68]), .Z(n4558) );
  XNOR U4537 ( .A(n4345), .B(n4559), .Z(n4341) );
  NAND U4538 ( .A(B[69]), .B(A[0]), .Z(n4559) );
  NAND U4539 ( .A(B[68]), .B(A[1]), .Z(n4345) );
  NAND U4540 ( .A(n4560), .B(n4561), .Z(n149) );
  NANDN U4541 ( .A(n4562), .B(n4563), .Z(n4561) );
  OR U4542 ( .A(n4564), .B(n4565), .Z(n4563) );
  NAND U4543 ( .A(n4565), .B(n4564), .Z(n4560) );
  XOR U4544 ( .A(n151), .B(n150), .Z(\A1[66] ) );
  XOR U4545 ( .A(n4565), .B(n4566), .Z(n150) );
  XNOR U4546 ( .A(n4564), .B(n4562), .Z(n4566) );
  AND U4547 ( .A(n4567), .B(n4568), .Z(n4562) );
  NANDN U4548 ( .A(n4569), .B(n4570), .Z(n4568) );
  NANDN U4549 ( .A(n4571), .B(n4572), .Z(n4570) );
  NANDN U4550 ( .A(n4572), .B(n4571), .Z(n4567) );
  ANDN U4551 ( .B(B[37]), .A(n54), .Z(n4564) );
  XNOR U4552 ( .A(n4359), .B(n4573), .Z(n4565) );
  XNOR U4553 ( .A(n4358), .B(n4356), .Z(n4573) );
  AND U4554 ( .A(n4574), .B(n4575), .Z(n4356) );
  NANDN U4555 ( .A(n4576), .B(n4577), .Z(n4575) );
  OR U4556 ( .A(n4578), .B(n4579), .Z(n4577) );
  NAND U4557 ( .A(n4579), .B(n4578), .Z(n4574) );
  ANDN U4558 ( .B(B[38]), .A(n55), .Z(n4358) );
  XNOR U4559 ( .A(n4366), .B(n4580), .Z(n4359) );
  XNOR U4560 ( .A(n4365), .B(n4363), .Z(n4580) );
  AND U4561 ( .A(n4581), .B(n4582), .Z(n4363) );
  NANDN U4562 ( .A(n4583), .B(n4584), .Z(n4582) );
  NANDN U4563 ( .A(n4585), .B(n4586), .Z(n4584) );
  NANDN U4564 ( .A(n4586), .B(n4585), .Z(n4581) );
  ANDN U4565 ( .B(B[39]), .A(n56), .Z(n4365) );
  XNOR U4566 ( .A(n4373), .B(n4587), .Z(n4366) );
  XNOR U4567 ( .A(n4372), .B(n4370), .Z(n4587) );
  AND U4568 ( .A(n4588), .B(n4589), .Z(n4370) );
  NANDN U4569 ( .A(n4590), .B(n4591), .Z(n4589) );
  OR U4570 ( .A(n4592), .B(n4593), .Z(n4591) );
  NAND U4571 ( .A(n4593), .B(n4592), .Z(n4588) );
  ANDN U4572 ( .B(B[40]), .A(n57), .Z(n4372) );
  XNOR U4573 ( .A(n4380), .B(n4594), .Z(n4373) );
  XNOR U4574 ( .A(n4379), .B(n4377), .Z(n4594) );
  AND U4575 ( .A(n4595), .B(n4596), .Z(n4377) );
  NANDN U4576 ( .A(n4597), .B(n4598), .Z(n4596) );
  NANDN U4577 ( .A(n4599), .B(n4600), .Z(n4598) );
  NANDN U4578 ( .A(n4600), .B(n4599), .Z(n4595) );
  ANDN U4579 ( .B(B[41]), .A(n58), .Z(n4379) );
  XNOR U4580 ( .A(n4387), .B(n4601), .Z(n4380) );
  XNOR U4581 ( .A(n4386), .B(n4384), .Z(n4601) );
  AND U4582 ( .A(n4602), .B(n4603), .Z(n4384) );
  NANDN U4583 ( .A(n4604), .B(n4605), .Z(n4603) );
  OR U4584 ( .A(n4606), .B(n4607), .Z(n4605) );
  NAND U4585 ( .A(n4607), .B(n4606), .Z(n4602) );
  ANDN U4586 ( .B(B[42]), .A(n59), .Z(n4386) );
  XNOR U4587 ( .A(n4394), .B(n4608), .Z(n4387) );
  XNOR U4588 ( .A(n4393), .B(n4391), .Z(n4608) );
  AND U4589 ( .A(n4609), .B(n4610), .Z(n4391) );
  NANDN U4590 ( .A(n4611), .B(n4612), .Z(n4610) );
  NANDN U4591 ( .A(n4613), .B(n4614), .Z(n4612) );
  NANDN U4592 ( .A(n4614), .B(n4613), .Z(n4609) );
  ANDN U4593 ( .B(B[43]), .A(n60), .Z(n4393) );
  XNOR U4594 ( .A(n4401), .B(n4615), .Z(n4394) );
  XNOR U4595 ( .A(n4400), .B(n4398), .Z(n4615) );
  AND U4596 ( .A(n4616), .B(n4617), .Z(n4398) );
  NANDN U4597 ( .A(n4618), .B(n4619), .Z(n4617) );
  OR U4598 ( .A(n4620), .B(n4621), .Z(n4619) );
  NAND U4599 ( .A(n4621), .B(n4620), .Z(n4616) );
  ANDN U4600 ( .B(B[44]), .A(n61), .Z(n4400) );
  XNOR U4601 ( .A(n4408), .B(n4622), .Z(n4401) );
  XNOR U4602 ( .A(n4407), .B(n4405), .Z(n4622) );
  AND U4603 ( .A(n4623), .B(n4624), .Z(n4405) );
  NANDN U4604 ( .A(n4625), .B(n4626), .Z(n4624) );
  NANDN U4605 ( .A(n4627), .B(n4628), .Z(n4626) );
  NANDN U4606 ( .A(n4628), .B(n4627), .Z(n4623) );
  ANDN U4607 ( .B(B[45]), .A(n62), .Z(n4407) );
  XNOR U4608 ( .A(n4415), .B(n4629), .Z(n4408) );
  XNOR U4609 ( .A(n4414), .B(n4412), .Z(n4629) );
  AND U4610 ( .A(n4630), .B(n4631), .Z(n4412) );
  NANDN U4611 ( .A(n4632), .B(n4633), .Z(n4631) );
  OR U4612 ( .A(n4634), .B(n4635), .Z(n4633) );
  NAND U4613 ( .A(n4635), .B(n4634), .Z(n4630) );
  ANDN U4614 ( .B(B[46]), .A(n63), .Z(n4414) );
  XNOR U4615 ( .A(n4422), .B(n4636), .Z(n4415) );
  XNOR U4616 ( .A(n4421), .B(n4419), .Z(n4636) );
  AND U4617 ( .A(n4637), .B(n4638), .Z(n4419) );
  NANDN U4618 ( .A(n4639), .B(n4640), .Z(n4638) );
  NANDN U4619 ( .A(n4641), .B(n4642), .Z(n4640) );
  NANDN U4620 ( .A(n4642), .B(n4641), .Z(n4637) );
  ANDN U4621 ( .B(B[47]), .A(n64), .Z(n4421) );
  XNOR U4622 ( .A(n4429), .B(n4643), .Z(n4422) );
  XNOR U4623 ( .A(n4428), .B(n4426), .Z(n4643) );
  AND U4624 ( .A(n4644), .B(n4645), .Z(n4426) );
  NANDN U4625 ( .A(n4646), .B(n4647), .Z(n4645) );
  OR U4626 ( .A(n4648), .B(n4649), .Z(n4647) );
  NAND U4627 ( .A(n4649), .B(n4648), .Z(n4644) );
  ANDN U4628 ( .B(B[48]), .A(n65), .Z(n4428) );
  XNOR U4629 ( .A(n4436), .B(n4650), .Z(n4429) );
  XNOR U4630 ( .A(n4435), .B(n4433), .Z(n4650) );
  AND U4631 ( .A(n4651), .B(n4652), .Z(n4433) );
  NANDN U4632 ( .A(n4653), .B(n4654), .Z(n4652) );
  NANDN U4633 ( .A(n4655), .B(n4656), .Z(n4654) );
  NANDN U4634 ( .A(n4656), .B(n4655), .Z(n4651) );
  ANDN U4635 ( .B(B[49]), .A(n66), .Z(n4435) );
  XNOR U4636 ( .A(n4443), .B(n4657), .Z(n4436) );
  XNOR U4637 ( .A(n4442), .B(n4440), .Z(n4657) );
  AND U4638 ( .A(n4658), .B(n4659), .Z(n4440) );
  NANDN U4639 ( .A(n4660), .B(n4661), .Z(n4659) );
  OR U4640 ( .A(n4662), .B(n4663), .Z(n4661) );
  NAND U4641 ( .A(n4663), .B(n4662), .Z(n4658) );
  ANDN U4642 ( .B(B[50]), .A(n67), .Z(n4442) );
  XNOR U4643 ( .A(n4450), .B(n4664), .Z(n4443) );
  XNOR U4644 ( .A(n4449), .B(n4447), .Z(n4664) );
  AND U4645 ( .A(n4665), .B(n4666), .Z(n4447) );
  NANDN U4646 ( .A(n4667), .B(n4668), .Z(n4666) );
  NANDN U4647 ( .A(n4669), .B(n4670), .Z(n4668) );
  NANDN U4648 ( .A(n4670), .B(n4669), .Z(n4665) );
  ANDN U4649 ( .B(B[51]), .A(n68), .Z(n4449) );
  XNOR U4650 ( .A(n4457), .B(n4671), .Z(n4450) );
  XNOR U4651 ( .A(n4456), .B(n4454), .Z(n4671) );
  AND U4652 ( .A(n4672), .B(n4673), .Z(n4454) );
  NANDN U4653 ( .A(n4674), .B(n4675), .Z(n4673) );
  OR U4654 ( .A(n4676), .B(n4677), .Z(n4675) );
  NAND U4655 ( .A(n4677), .B(n4676), .Z(n4672) );
  ANDN U4656 ( .B(B[52]), .A(n69), .Z(n4456) );
  XNOR U4657 ( .A(n4464), .B(n4678), .Z(n4457) );
  XNOR U4658 ( .A(n4463), .B(n4461), .Z(n4678) );
  AND U4659 ( .A(n4679), .B(n4680), .Z(n4461) );
  NANDN U4660 ( .A(n4681), .B(n4682), .Z(n4680) );
  NANDN U4661 ( .A(n4683), .B(n4684), .Z(n4682) );
  NANDN U4662 ( .A(n4684), .B(n4683), .Z(n4679) );
  ANDN U4663 ( .B(B[53]), .A(n70), .Z(n4463) );
  XNOR U4664 ( .A(n4471), .B(n4685), .Z(n4464) );
  XNOR U4665 ( .A(n4470), .B(n4468), .Z(n4685) );
  AND U4666 ( .A(n4686), .B(n4687), .Z(n4468) );
  NANDN U4667 ( .A(n4688), .B(n4689), .Z(n4687) );
  OR U4668 ( .A(n4690), .B(n4691), .Z(n4689) );
  NAND U4669 ( .A(n4691), .B(n4690), .Z(n4686) );
  ANDN U4670 ( .B(B[54]), .A(n71), .Z(n4470) );
  XNOR U4671 ( .A(n4478), .B(n4692), .Z(n4471) );
  XNOR U4672 ( .A(n4477), .B(n4475), .Z(n4692) );
  AND U4673 ( .A(n4693), .B(n4694), .Z(n4475) );
  NANDN U4674 ( .A(n4695), .B(n4696), .Z(n4694) );
  NANDN U4675 ( .A(n4697), .B(n4698), .Z(n4696) );
  NANDN U4676 ( .A(n4698), .B(n4697), .Z(n4693) );
  ANDN U4677 ( .B(B[55]), .A(n72), .Z(n4477) );
  XNOR U4678 ( .A(n4485), .B(n4699), .Z(n4478) );
  XNOR U4679 ( .A(n4484), .B(n4482), .Z(n4699) );
  AND U4680 ( .A(n4700), .B(n4701), .Z(n4482) );
  NANDN U4681 ( .A(n4702), .B(n4703), .Z(n4701) );
  OR U4682 ( .A(n4704), .B(n4705), .Z(n4703) );
  NAND U4683 ( .A(n4705), .B(n4704), .Z(n4700) );
  ANDN U4684 ( .B(B[56]), .A(n73), .Z(n4484) );
  XNOR U4685 ( .A(n4492), .B(n4706), .Z(n4485) );
  XNOR U4686 ( .A(n4491), .B(n4489), .Z(n4706) );
  AND U4687 ( .A(n4707), .B(n4708), .Z(n4489) );
  NANDN U4688 ( .A(n4709), .B(n4710), .Z(n4708) );
  NANDN U4689 ( .A(n4711), .B(n4712), .Z(n4710) );
  NANDN U4690 ( .A(n4712), .B(n4711), .Z(n4707) );
  ANDN U4691 ( .B(B[57]), .A(n74), .Z(n4491) );
  XNOR U4692 ( .A(n4499), .B(n4713), .Z(n4492) );
  XNOR U4693 ( .A(n4498), .B(n4496), .Z(n4713) );
  AND U4694 ( .A(n4714), .B(n4715), .Z(n4496) );
  NANDN U4695 ( .A(n4716), .B(n4717), .Z(n4715) );
  OR U4696 ( .A(n4718), .B(n4719), .Z(n4717) );
  NAND U4697 ( .A(n4719), .B(n4718), .Z(n4714) );
  ANDN U4698 ( .B(B[58]), .A(n75), .Z(n4498) );
  XNOR U4699 ( .A(n4506), .B(n4720), .Z(n4499) );
  XNOR U4700 ( .A(n4505), .B(n4503), .Z(n4720) );
  AND U4701 ( .A(n4721), .B(n4722), .Z(n4503) );
  NANDN U4702 ( .A(n4723), .B(n4724), .Z(n4722) );
  NANDN U4703 ( .A(n4725), .B(n4726), .Z(n4724) );
  NANDN U4704 ( .A(n4726), .B(n4725), .Z(n4721) );
  ANDN U4705 ( .B(B[59]), .A(n76), .Z(n4505) );
  XNOR U4706 ( .A(n4513), .B(n4727), .Z(n4506) );
  XNOR U4707 ( .A(n4512), .B(n4510), .Z(n4727) );
  AND U4708 ( .A(n4728), .B(n4729), .Z(n4510) );
  NANDN U4709 ( .A(n4730), .B(n4731), .Z(n4729) );
  OR U4710 ( .A(n4732), .B(n4733), .Z(n4731) );
  NAND U4711 ( .A(n4733), .B(n4732), .Z(n4728) );
  ANDN U4712 ( .B(B[60]), .A(n77), .Z(n4512) );
  XNOR U4713 ( .A(n4520), .B(n4734), .Z(n4513) );
  XNOR U4714 ( .A(n4519), .B(n4517), .Z(n4734) );
  AND U4715 ( .A(n4735), .B(n4736), .Z(n4517) );
  NANDN U4716 ( .A(n4737), .B(n4738), .Z(n4736) );
  NANDN U4717 ( .A(n4739), .B(n4740), .Z(n4738) );
  NANDN U4718 ( .A(n4740), .B(n4739), .Z(n4735) );
  ANDN U4719 ( .B(B[61]), .A(n78), .Z(n4519) );
  XNOR U4720 ( .A(n4527), .B(n4741), .Z(n4520) );
  XNOR U4721 ( .A(n4526), .B(n4524), .Z(n4741) );
  AND U4722 ( .A(n4742), .B(n4743), .Z(n4524) );
  NANDN U4723 ( .A(n4744), .B(n4745), .Z(n4743) );
  OR U4724 ( .A(n4746), .B(n4747), .Z(n4745) );
  NAND U4725 ( .A(n4747), .B(n4746), .Z(n4742) );
  ANDN U4726 ( .B(B[62]), .A(n79), .Z(n4526) );
  XNOR U4727 ( .A(n4534), .B(n4748), .Z(n4527) );
  XNOR U4728 ( .A(n4533), .B(n4531), .Z(n4748) );
  AND U4729 ( .A(n4749), .B(n4750), .Z(n4531) );
  NANDN U4730 ( .A(n4751), .B(n4752), .Z(n4750) );
  NANDN U4731 ( .A(n4753), .B(n4754), .Z(n4752) );
  NANDN U4732 ( .A(n4754), .B(n4753), .Z(n4749) );
  ANDN U4733 ( .B(B[63]), .A(n80), .Z(n4533) );
  XNOR U4734 ( .A(n4541), .B(n4755), .Z(n4534) );
  XNOR U4735 ( .A(n4540), .B(n4538), .Z(n4755) );
  AND U4736 ( .A(n4756), .B(n4757), .Z(n4538) );
  NANDN U4737 ( .A(n4758), .B(n4759), .Z(n4757) );
  OR U4738 ( .A(n4760), .B(n4761), .Z(n4759) );
  NAND U4739 ( .A(n4761), .B(n4760), .Z(n4756) );
  ANDN U4740 ( .B(B[64]), .A(n81), .Z(n4540) );
  XNOR U4741 ( .A(n4548), .B(n4762), .Z(n4541) );
  XNOR U4742 ( .A(n4547), .B(n4545), .Z(n4762) );
  AND U4743 ( .A(n4763), .B(n4764), .Z(n4545) );
  NANDN U4744 ( .A(n4765), .B(n4766), .Z(n4764) );
  NAND U4745 ( .A(n4767), .B(n4768), .Z(n4766) );
  ANDN U4746 ( .B(B[65]), .A(n82), .Z(n4547) );
  XOR U4747 ( .A(n4554), .B(n4769), .Z(n4548) );
  XNOR U4748 ( .A(n4552), .B(n4555), .Z(n4769) );
  NAND U4749 ( .A(A[2]), .B(B[66]), .Z(n4555) );
  NANDN U4750 ( .A(n4770), .B(n4771), .Z(n4552) );
  AND U4751 ( .A(A[0]), .B(B[67]), .Z(n4771) );
  XNOR U4752 ( .A(n4557), .B(n4772), .Z(n4554) );
  NAND U4753 ( .A(A[0]), .B(B[68]), .Z(n4772) );
  NAND U4754 ( .A(B[67]), .B(A[1]), .Z(n4557) );
  NAND U4755 ( .A(n4773), .B(n4774), .Z(n151) );
  NANDN U4756 ( .A(n4775), .B(n4776), .Z(n4774) );
  OR U4757 ( .A(n4777), .B(n4778), .Z(n4776) );
  NAND U4758 ( .A(n4778), .B(n4777), .Z(n4773) );
  XOR U4759 ( .A(n153), .B(n152), .Z(\A1[65] ) );
  XOR U4760 ( .A(n4778), .B(n4779), .Z(n152) );
  XNOR U4761 ( .A(n4777), .B(n4775), .Z(n4779) );
  AND U4762 ( .A(n4780), .B(n4781), .Z(n4775) );
  NANDN U4763 ( .A(n4782), .B(n4783), .Z(n4781) );
  NANDN U4764 ( .A(n4784), .B(n4785), .Z(n4783) );
  NANDN U4765 ( .A(n4785), .B(n4784), .Z(n4780) );
  ANDN U4766 ( .B(B[36]), .A(n54), .Z(n4777) );
  XNOR U4767 ( .A(n4572), .B(n4786), .Z(n4778) );
  XNOR U4768 ( .A(n4571), .B(n4569), .Z(n4786) );
  AND U4769 ( .A(n4787), .B(n4788), .Z(n4569) );
  NANDN U4770 ( .A(n4789), .B(n4790), .Z(n4788) );
  OR U4771 ( .A(n4791), .B(n4792), .Z(n4790) );
  NAND U4772 ( .A(n4792), .B(n4791), .Z(n4787) );
  ANDN U4773 ( .B(B[37]), .A(n55), .Z(n4571) );
  XNOR U4774 ( .A(n4579), .B(n4793), .Z(n4572) );
  XNOR U4775 ( .A(n4578), .B(n4576), .Z(n4793) );
  AND U4776 ( .A(n4794), .B(n4795), .Z(n4576) );
  NANDN U4777 ( .A(n4796), .B(n4797), .Z(n4795) );
  NANDN U4778 ( .A(n4798), .B(n4799), .Z(n4797) );
  NANDN U4779 ( .A(n4799), .B(n4798), .Z(n4794) );
  ANDN U4780 ( .B(B[38]), .A(n56), .Z(n4578) );
  XNOR U4781 ( .A(n4586), .B(n4800), .Z(n4579) );
  XNOR U4782 ( .A(n4585), .B(n4583), .Z(n4800) );
  AND U4783 ( .A(n4801), .B(n4802), .Z(n4583) );
  NANDN U4784 ( .A(n4803), .B(n4804), .Z(n4802) );
  OR U4785 ( .A(n4805), .B(n4806), .Z(n4804) );
  NAND U4786 ( .A(n4806), .B(n4805), .Z(n4801) );
  ANDN U4787 ( .B(B[39]), .A(n57), .Z(n4585) );
  XNOR U4788 ( .A(n4593), .B(n4807), .Z(n4586) );
  XNOR U4789 ( .A(n4592), .B(n4590), .Z(n4807) );
  AND U4790 ( .A(n4808), .B(n4809), .Z(n4590) );
  NANDN U4791 ( .A(n4810), .B(n4811), .Z(n4809) );
  NANDN U4792 ( .A(n4812), .B(n4813), .Z(n4811) );
  NANDN U4793 ( .A(n4813), .B(n4812), .Z(n4808) );
  ANDN U4794 ( .B(B[40]), .A(n58), .Z(n4592) );
  XNOR U4795 ( .A(n4600), .B(n4814), .Z(n4593) );
  XNOR U4796 ( .A(n4599), .B(n4597), .Z(n4814) );
  AND U4797 ( .A(n4815), .B(n4816), .Z(n4597) );
  NANDN U4798 ( .A(n4817), .B(n4818), .Z(n4816) );
  OR U4799 ( .A(n4819), .B(n4820), .Z(n4818) );
  NAND U4800 ( .A(n4820), .B(n4819), .Z(n4815) );
  ANDN U4801 ( .B(B[41]), .A(n59), .Z(n4599) );
  XNOR U4802 ( .A(n4607), .B(n4821), .Z(n4600) );
  XNOR U4803 ( .A(n4606), .B(n4604), .Z(n4821) );
  AND U4804 ( .A(n4822), .B(n4823), .Z(n4604) );
  NANDN U4805 ( .A(n4824), .B(n4825), .Z(n4823) );
  NANDN U4806 ( .A(n4826), .B(n4827), .Z(n4825) );
  NANDN U4807 ( .A(n4827), .B(n4826), .Z(n4822) );
  ANDN U4808 ( .B(B[42]), .A(n60), .Z(n4606) );
  XNOR U4809 ( .A(n4614), .B(n4828), .Z(n4607) );
  XNOR U4810 ( .A(n4613), .B(n4611), .Z(n4828) );
  AND U4811 ( .A(n4829), .B(n4830), .Z(n4611) );
  NANDN U4812 ( .A(n4831), .B(n4832), .Z(n4830) );
  OR U4813 ( .A(n4833), .B(n4834), .Z(n4832) );
  NAND U4814 ( .A(n4834), .B(n4833), .Z(n4829) );
  ANDN U4815 ( .B(B[43]), .A(n61), .Z(n4613) );
  XNOR U4816 ( .A(n4621), .B(n4835), .Z(n4614) );
  XNOR U4817 ( .A(n4620), .B(n4618), .Z(n4835) );
  AND U4818 ( .A(n4836), .B(n4837), .Z(n4618) );
  NANDN U4819 ( .A(n4838), .B(n4839), .Z(n4837) );
  NANDN U4820 ( .A(n4840), .B(n4841), .Z(n4839) );
  NANDN U4821 ( .A(n4841), .B(n4840), .Z(n4836) );
  ANDN U4822 ( .B(B[44]), .A(n62), .Z(n4620) );
  XNOR U4823 ( .A(n4628), .B(n4842), .Z(n4621) );
  XNOR U4824 ( .A(n4627), .B(n4625), .Z(n4842) );
  AND U4825 ( .A(n4843), .B(n4844), .Z(n4625) );
  NANDN U4826 ( .A(n4845), .B(n4846), .Z(n4844) );
  OR U4827 ( .A(n4847), .B(n4848), .Z(n4846) );
  NAND U4828 ( .A(n4848), .B(n4847), .Z(n4843) );
  ANDN U4829 ( .B(B[45]), .A(n63), .Z(n4627) );
  XNOR U4830 ( .A(n4635), .B(n4849), .Z(n4628) );
  XNOR U4831 ( .A(n4634), .B(n4632), .Z(n4849) );
  AND U4832 ( .A(n4850), .B(n4851), .Z(n4632) );
  NANDN U4833 ( .A(n4852), .B(n4853), .Z(n4851) );
  NANDN U4834 ( .A(n4854), .B(n4855), .Z(n4853) );
  NANDN U4835 ( .A(n4855), .B(n4854), .Z(n4850) );
  ANDN U4836 ( .B(B[46]), .A(n64), .Z(n4634) );
  XNOR U4837 ( .A(n4642), .B(n4856), .Z(n4635) );
  XNOR U4838 ( .A(n4641), .B(n4639), .Z(n4856) );
  AND U4839 ( .A(n4857), .B(n4858), .Z(n4639) );
  NANDN U4840 ( .A(n4859), .B(n4860), .Z(n4858) );
  OR U4841 ( .A(n4861), .B(n4862), .Z(n4860) );
  NAND U4842 ( .A(n4862), .B(n4861), .Z(n4857) );
  ANDN U4843 ( .B(B[47]), .A(n65), .Z(n4641) );
  XNOR U4844 ( .A(n4649), .B(n4863), .Z(n4642) );
  XNOR U4845 ( .A(n4648), .B(n4646), .Z(n4863) );
  AND U4846 ( .A(n4864), .B(n4865), .Z(n4646) );
  NANDN U4847 ( .A(n4866), .B(n4867), .Z(n4865) );
  NANDN U4848 ( .A(n4868), .B(n4869), .Z(n4867) );
  NANDN U4849 ( .A(n4869), .B(n4868), .Z(n4864) );
  ANDN U4850 ( .B(B[48]), .A(n66), .Z(n4648) );
  XNOR U4851 ( .A(n4656), .B(n4870), .Z(n4649) );
  XNOR U4852 ( .A(n4655), .B(n4653), .Z(n4870) );
  AND U4853 ( .A(n4871), .B(n4872), .Z(n4653) );
  NANDN U4854 ( .A(n4873), .B(n4874), .Z(n4872) );
  OR U4855 ( .A(n4875), .B(n4876), .Z(n4874) );
  NAND U4856 ( .A(n4876), .B(n4875), .Z(n4871) );
  ANDN U4857 ( .B(B[49]), .A(n67), .Z(n4655) );
  XNOR U4858 ( .A(n4663), .B(n4877), .Z(n4656) );
  XNOR U4859 ( .A(n4662), .B(n4660), .Z(n4877) );
  AND U4860 ( .A(n4878), .B(n4879), .Z(n4660) );
  NANDN U4861 ( .A(n4880), .B(n4881), .Z(n4879) );
  NANDN U4862 ( .A(n4882), .B(n4883), .Z(n4881) );
  NANDN U4863 ( .A(n4883), .B(n4882), .Z(n4878) );
  ANDN U4864 ( .B(B[50]), .A(n68), .Z(n4662) );
  XNOR U4865 ( .A(n4670), .B(n4884), .Z(n4663) );
  XNOR U4866 ( .A(n4669), .B(n4667), .Z(n4884) );
  AND U4867 ( .A(n4885), .B(n4886), .Z(n4667) );
  NANDN U4868 ( .A(n4887), .B(n4888), .Z(n4886) );
  OR U4869 ( .A(n4889), .B(n4890), .Z(n4888) );
  NAND U4870 ( .A(n4890), .B(n4889), .Z(n4885) );
  ANDN U4871 ( .B(B[51]), .A(n69), .Z(n4669) );
  XNOR U4872 ( .A(n4677), .B(n4891), .Z(n4670) );
  XNOR U4873 ( .A(n4676), .B(n4674), .Z(n4891) );
  AND U4874 ( .A(n4892), .B(n4893), .Z(n4674) );
  NANDN U4875 ( .A(n4894), .B(n4895), .Z(n4893) );
  NANDN U4876 ( .A(n4896), .B(n4897), .Z(n4895) );
  NANDN U4877 ( .A(n4897), .B(n4896), .Z(n4892) );
  ANDN U4878 ( .B(B[52]), .A(n70), .Z(n4676) );
  XNOR U4879 ( .A(n4684), .B(n4898), .Z(n4677) );
  XNOR U4880 ( .A(n4683), .B(n4681), .Z(n4898) );
  AND U4881 ( .A(n4899), .B(n4900), .Z(n4681) );
  NANDN U4882 ( .A(n4901), .B(n4902), .Z(n4900) );
  OR U4883 ( .A(n4903), .B(n4904), .Z(n4902) );
  NAND U4884 ( .A(n4904), .B(n4903), .Z(n4899) );
  ANDN U4885 ( .B(B[53]), .A(n71), .Z(n4683) );
  XNOR U4886 ( .A(n4691), .B(n4905), .Z(n4684) );
  XNOR U4887 ( .A(n4690), .B(n4688), .Z(n4905) );
  AND U4888 ( .A(n4906), .B(n4907), .Z(n4688) );
  NANDN U4889 ( .A(n4908), .B(n4909), .Z(n4907) );
  NANDN U4890 ( .A(n4910), .B(n4911), .Z(n4909) );
  NANDN U4891 ( .A(n4911), .B(n4910), .Z(n4906) );
  ANDN U4892 ( .B(B[54]), .A(n72), .Z(n4690) );
  XNOR U4893 ( .A(n4698), .B(n4912), .Z(n4691) );
  XNOR U4894 ( .A(n4697), .B(n4695), .Z(n4912) );
  AND U4895 ( .A(n4913), .B(n4914), .Z(n4695) );
  NANDN U4896 ( .A(n4915), .B(n4916), .Z(n4914) );
  OR U4897 ( .A(n4917), .B(n4918), .Z(n4916) );
  NAND U4898 ( .A(n4918), .B(n4917), .Z(n4913) );
  ANDN U4899 ( .B(B[55]), .A(n73), .Z(n4697) );
  XNOR U4900 ( .A(n4705), .B(n4919), .Z(n4698) );
  XNOR U4901 ( .A(n4704), .B(n4702), .Z(n4919) );
  AND U4902 ( .A(n4920), .B(n4921), .Z(n4702) );
  NANDN U4903 ( .A(n4922), .B(n4923), .Z(n4921) );
  NANDN U4904 ( .A(n4924), .B(n4925), .Z(n4923) );
  NANDN U4905 ( .A(n4925), .B(n4924), .Z(n4920) );
  ANDN U4906 ( .B(B[56]), .A(n74), .Z(n4704) );
  XNOR U4907 ( .A(n4712), .B(n4926), .Z(n4705) );
  XNOR U4908 ( .A(n4711), .B(n4709), .Z(n4926) );
  AND U4909 ( .A(n4927), .B(n4928), .Z(n4709) );
  NANDN U4910 ( .A(n4929), .B(n4930), .Z(n4928) );
  OR U4911 ( .A(n4931), .B(n4932), .Z(n4930) );
  NAND U4912 ( .A(n4932), .B(n4931), .Z(n4927) );
  ANDN U4913 ( .B(B[57]), .A(n75), .Z(n4711) );
  XNOR U4914 ( .A(n4719), .B(n4933), .Z(n4712) );
  XNOR U4915 ( .A(n4718), .B(n4716), .Z(n4933) );
  AND U4916 ( .A(n4934), .B(n4935), .Z(n4716) );
  NANDN U4917 ( .A(n4936), .B(n4937), .Z(n4935) );
  NANDN U4918 ( .A(n4938), .B(n4939), .Z(n4937) );
  NANDN U4919 ( .A(n4939), .B(n4938), .Z(n4934) );
  ANDN U4920 ( .B(B[58]), .A(n76), .Z(n4718) );
  XNOR U4921 ( .A(n4726), .B(n4940), .Z(n4719) );
  XNOR U4922 ( .A(n4725), .B(n4723), .Z(n4940) );
  AND U4923 ( .A(n4941), .B(n4942), .Z(n4723) );
  NANDN U4924 ( .A(n4943), .B(n4944), .Z(n4942) );
  OR U4925 ( .A(n4945), .B(n4946), .Z(n4944) );
  NAND U4926 ( .A(n4946), .B(n4945), .Z(n4941) );
  ANDN U4927 ( .B(B[59]), .A(n77), .Z(n4725) );
  XNOR U4928 ( .A(n4733), .B(n4947), .Z(n4726) );
  XNOR U4929 ( .A(n4732), .B(n4730), .Z(n4947) );
  AND U4930 ( .A(n4948), .B(n4949), .Z(n4730) );
  NANDN U4931 ( .A(n4950), .B(n4951), .Z(n4949) );
  NANDN U4932 ( .A(n4952), .B(n4953), .Z(n4951) );
  NANDN U4933 ( .A(n4953), .B(n4952), .Z(n4948) );
  ANDN U4934 ( .B(B[60]), .A(n78), .Z(n4732) );
  XNOR U4935 ( .A(n4740), .B(n4954), .Z(n4733) );
  XNOR U4936 ( .A(n4739), .B(n4737), .Z(n4954) );
  AND U4937 ( .A(n4955), .B(n4956), .Z(n4737) );
  NANDN U4938 ( .A(n4957), .B(n4958), .Z(n4956) );
  OR U4939 ( .A(n4959), .B(n4960), .Z(n4958) );
  NAND U4940 ( .A(n4960), .B(n4959), .Z(n4955) );
  ANDN U4941 ( .B(B[61]), .A(n79), .Z(n4739) );
  XNOR U4942 ( .A(n4747), .B(n4961), .Z(n4740) );
  XNOR U4943 ( .A(n4746), .B(n4744), .Z(n4961) );
  AND U4944 ( .A(n4962), .B(n4963), .Z(n4744) );
  NANDN U4945 ( .A(n4964), .B(n4965), .Z(n4963) );
  NANDN U4946 ( .A(n4966), .B(n4967), .Z(n4965) );
  NANDN U4947 ( .A(n4967), .B(n4966), .Z(n4962) );
  ANDN U4948 ( .B(B[62]), .A(n80), .Z(n4746) );
  XNOR U4949 ( .A(n4754), .B(n4968), .Z(n4747) );
  XNOR U4950 ( .A(n4753), .B(n4751), .Z(n4968) );
  AND U4951 ( .A(n4969), .B(n4970), .Z(n4751) );
  NANDN U4952 ( .A(n4971), .B(n4972), .Z(n4970) );
  OR U4953 ( .A(n4973), .B(n4974), .Z(n4972) );
  NAND U4954 ( .A(n4974), .B(n4973), .Z(n4969) );
  ANDN U4955 ( .B(B[63]), .A(n81), .Z(n4753) );
  XNOR U4956 ( .A(n4761), .B(n4975), .Z(n4754) );
  XNOR U4957 ( .A(n4760), .B(n4758), .Z(n4975) );
  AND U4958 ( .A(n4976), .B(n4977), .Z(n4758) );
  NANDN U4959 ( .A(n4978), .B(n4979), .Z(n4977) );
  NAND U4960 ( .A(n4980), .B(n4981), .Z(n4979) );
  ANDN U4961 ( .B(B[64]), .A(n82), .Z(n4760) );
  XOR U4962 ( .A(n4767), .B(n4982), .Z(n4761) );
  XNOR U4963 ( .A(n4765), .B(n4768), .Z(n4982) );
  NAND U4964 ( .A(A[2]), .B(B[65]), .Z(n4768) );
  NANDN U4965 ( .A(n4983), .B(n4984), .Z(n4765) );
  AND U4966 ( .A(A[0]), .B(B[66]), .Z(n4984) );
  XNOR U4967 ( .A(n4770), .B(n4985), .Z(n4767) );
  NAND U4968 ( .A(A[0]), .B(B[67]), .Z(n4985) );
  NAND U4969 ( .A(B[66]), .B(A[1]), .Z(n4770) );
  NAND U4970 ( .A(n4986), .B(n4987), .Z(n153) );
  NANDN U4971 ( .A(n4988), .B(n4989), .Z(n4987) );
  OR U4972 ( .A(n4990), .B(n4991), .Z(n4989) );
  NAND U4973 ( .A(n4991), .B(n4990), .Z(n4986) );
  XOR U4974 ( .A(n155), .B(n154), .Z(\A1[64] ) );
  XOR U4975 ( .A(n4991), .B(n4992), .Z(n154) );
  XNOR U4976 ( .A(n4990), .B(n4988), .Z(n4992) );
  AND U4977 ( .A(n4993), .B(n4994), .Z(n4988) );
  NANDN U4978 ( .A(n4995), .B(n4996), .Z(n4994) );
  NANDN U4979 ( .A(n4997), .B(n4998), .Z(n4996) );
  NANDN U4980 ( .A(n4998), .B(n4997), .Z(n4993) );
  ANDN U4981 ( .B(B[35]), .A(n54), .Z(n4990) );
  XNOR U4982 ( .A(n4785), .B(n4999), .Z(n4991) );
  XNOR U4983 ( .A(n4784), .B(n4782), .Z(n4999) );
  AND U4984 ( .A(n5000), .B(n5001), .Z(n4782) );
  NANDN U4985 ( .A(n5002), .B(n5003), .Z(n5001) );
  OR U4986 ( .A(n5004), .B(n5005), .Z(n5003) );
  NAND U4987 ( .A(n5005), .B(n5004), .Z(n5000) );
  ANDN U4988 ( .B(B[36]), .A(n55), .Z(n4784) );
  XNOR U4989 ( .A(n4792), .B(n5006), .Z(n4785) );
  XNOR U4990 ( .A(n4791), .B(n4789), .Z(n5006) );
  AND U4991 ( .A(n5007), .B(n5008), .Z(n4789) );
  NANDN U4992 ( .A(n5009), .B(n5010), .Z(n5008) );
  NANDN U4993 ( .A(n5011), .B(n5012), .Z(n5010) );
  NANDN U4994 ( .A(n5012), .B(n5011), .Z(n5007) );
  ANDN U4995 ( .B(B[37]), .A(n56), .Z(n4791) );
  XNOR U4996 ( .A(n4799), .B(n5013), .Z(n4792) );
  XNOR U4997 ( .A(n4798), .B(n4796), .Z(n5013) );
  AND U4998 ( .A(n5014), .B(n5015), .Z(n4796) );
  NANDN U4999 ( .A(n5016), .B(n5017), .Z(n5015) );
  OR U5000 ( .A(n5018), .B(n5019), .Z(n5017) );
  NAND U5001 ( .A(n5019), .B(n5018), .Z(n5014) );
  ANDN U5002 ( .B(B[38]), .A(n57), .Z(n4798) );
  XNOR U5003 ( .A(n4806), .B(n5020), .Z(n4799) );
  XNOR U5004 ( .A(n4805), .B(n4803), .Z(n5020) );
  AND U5005 ( .A(n5021), .B(n5022), .Z(n4803) );
  NANDN U5006 ( .A(n5023), .B(n5024), .Z(n5022) );
  NANDN U5007 ( .A(n5025), .B(n5026), .Z(n5024) );
  NANDN U5008 ( .A(n5026), .B(n5025), .Z(n5021) );
  ANDN U5009 ( .B(B[39]), .A(n58), .Z(n4805) );
  XNOR U5010 ( .A(n4813), .B(n5027), .Z(n4806) );
  XNOR U5011 ( .A(n4812), .B(n4810), .Z(n5027) );
  AND U5012 ( .A(n5028), .B(n5029), .Z(n4810) );
  NANDN U5013 ( .A(n5030), .B(n5031), .Z(n5029) );
  OR U5014 ( .A(n5032), .B(n5033), .Z(n5031) );
  NAND U5015 ( .A(n5033), .B(n5032), .Z(n5028) );
  ANDN U5016 ( .B(B[40]), .A(n59), .Z(n4812) );
  XNOR U5017 ( .A(n4820), .B(n5034), .Z(n4813) );
  XNOR U5018 ( .A(n4819), .B(n4817), .Z(n5034) );
  AND U5019 ( .A(n5035), .B(n5036), .Z(n4817) );
  NANDN U5020 ( .A(n5037), .B(n5038), .Z(n5036) );
  NANDN U5021 ( .A(n5039), .B(n5040), .Z(n5038) );
  NANDN U5022 ( .A(n5040), .B(n5039), .Z(n5035) );
  ANDN U5023 ( .B(B[41]), .A(n60), .Z(n4819) );
  XNOR U5024 ( .A(n4827), .B(n5041), .Z(n4820) );
  XNOR U5025 ( .A(n4826), .B(n4824), .Z(n5041) );
  AND U5026 ( .A(n5042), .B(n5043), .Z(n4824) );
  NANDN U5027 ( .A(n5044), .B(n5045), .Z(n5043) );
  OR U5028 ( .A(n5046), .B(n5047), .Z(n5045) );
  NAND U5029 ( .A(n5047), .B(n5046), .Z(n5042) );
  ANDN U5030 ( .B(B[42]), .A(n61), .Z(n4826) );
  XNOR U5031 ( .A(n4834), .B(n5048), .Z(n4827) );
  XNOR U5032 ( .A(n4833), .B(n4831), .Z(n5048) );
  AND U5033 ( .A(n5049), .B(n5050), .Z(n4831) );
  NANDN U5034 ( .A(n5051), .B(n5052), .Z(n5050) );
  NANDN U5035 ( .A(n5053), .B(n5054), .Z(n5052) );
  NANDN U5036 ( .A(n5054), .B(n5053), .Z(n5049) );
  ANDN U5037 ( .B(B[43]), .A(n62), .Z(n4833) );
  XNOR U5038 ( .A(n4841), .B(n5055), .Z(n4834) );
  XNOR U5039 ( .A(n4840), .B(n4838), .Z(n5055) );
  AND U5040 ( .A(n5056), .B(n5057), .Z(n4838) );
  NANDN U5041 ( .A(n5058), .B(n5059), .Z(n5057) );
  OR U5042 ( .A(n5060), .B(n5061), .Z(n5059) );
  NAND U5043 ( .A(n5061), .B(n5060), .Z(n5056) );
  ANDN U5044 ( .B(B[44]), .A(n63), .Z(n4840) );
  XNOR U5045 ( .A(n4848), .B(n5062), .Z(n4841) );
  XNOR U5046 ( .A(n4847), .B(n4845), .Z(n5062) );
  AND U5047 ( .A(n5063), .B(n5064), .Z(n4845) );
  NANDN U5048 ( .A(n5065), .B(n5066), .Z(n5064) );
  NANDN U5049 ( .A(n5067), .B(n5068), .Z(n5066) );
  NANDN U5050 ( .A(n5068), .B(n5067), .Z(n5063) );
  ANDN U5051 ( .B(B[45]), .A(n64), .Z(n4847) );
  XNOR U5052 ( .A(n4855), .B(n5069), .Z(n4848) );
  XNOR U5053 ( .A(n4854), .B(n4852), .Z(n5069) );
  AND U5054 ( .A(n5070), .B(n5071), .Z(n4852) );
  NANDN U5055 ( .A(n5072), .B(n5073), .Z(n5071) );
  OR U5056 ( .A(n5074), .B(n5075), .Z(n5073) );
  NAND U5057 ( .A(n5075), .B(n5074), .Z(n5070) );
  ANDN U5058 ( .B(B[46]), .A(n65), .Z(n4854) );
  XNOR U5059 ( .A(n4862), .B(n5076), .Z(n4855) );
  XNOR U5060 ( .A(n4861), .B(n4859), .Z(n5076) );
  AND U5061 ( .A(n5077), .B(n5078), .Z(n4859) );
  NANDN U5062 ( .A(n5079), .B(n5080), .Z(n5078) );
  NANDN U5063 ( .A(n5081), .B(n5082), .Z(n5080) );
  NANDN U5064 ( .A(n5082), .B(n5081), .Z(n5077) );
  ANDN U5065 ( .B(B[47]), .A(n66), .Z(n4861) );
  XNOR U5066 ( .A(n4869), .B(n5083), .Z(n4862) );
  XNOR U5067 ( .A(n4868), .B(n4866), .Z(n5083) );
  AND U5068 ( .A(n5084), .B(n5085), .Z(n4866) );
  NANDN U5069 ( .A(n5086), .B(n5087), .Z(n5085) );
  OR U5070 ( .A(n5088), .B(n5089), .Z(n5087) );
  NAND U5071 ( .A(n5089), .B(n5088), .Z(n5084) );
  ANDN U5072 ( .B(B[48]), .A(n67), .Z(n4868) );
  XNOR U5073 ( .A(n4876), .B(n5090), .Z(n4869) );
  XNOR U5074 ( .A(n4875), .B(n4873), .Z(n5090) );
  AND U5075 ( .A(n5091), .B(n5092), .Z(n4873) );
  NANDN U5076 ( .A(n5093), .B(n5094), .Z(n5092) );
  NANDN U5077 ( .A(n5095), .B(n5096), .Z(n5094) );
  NANDN U5078 ( .A(n5096), .B(n5095), .Z(n5091) );
  ANDN U5079 ( .B(B[49]), .A(n68), .Z(n4875) );
  XNOR U5080 ( .A(n4883), .B(n5097), .Z(n4876) );
  XNOR U5081 ( .A(n4882), .B(n4880), .Z(n5097) );
  AND U5082 ( .A(n5098), .B(n5099), .Z(n4880) );
  NANDN U5083 ( .A(n5100), .B(n5101), .Z(n5099) );
  OR U5084 ( .A(n5102), .B(n5103), .Z(n5101) );
  NAND U5085 ( .A(n5103), .B(n5102), .Z(n5098) );
  ANDN U5086 ( .B(B[50]), .A(n69), .Z(n4882) );
  XNOR U5087 ( .A(n4890), .B(n5104), .Z(n4883) );
  XNOR U5088 ( .A(n4889), .B(n4887), .Z(n5104) );
  AND U5089 ( .A(n5105), .B(n5106), .Z(n4887) );
  NANDN U5090 ( .A(n5107), .B(n5108), .Z(n5106) );
  NANDN U5091 ( .A(n5109), .B(n5110), .Z(n5108) );
  NANDN U5092 ( .A(n5110), .B(n5109), .Z(n5105) );
  ANDN U5093 ( .B(B[51]), .A(n70), .Z(n4889) );
  XNOR U5094 ( .A(n4897), .B(n5111), .Z(n4890) );
  XNOR U5095 ( .A(n4896), .B(n4894), .Z(n5111) );
  AND U5096 ( .A(n5112), .B(n5113), .Z(n4894) );
  NANDN U5097 ( .A(n5114), .B(n5115), .Z(n5113) );
  OR U5098 ( .A(n5116), .B(n5117), .Z(n5115) );
  NAND U5099 ( .A(n5117), .B(n5116), .Z(n5112) );
  ANDN U5100 ( .B(B[52]), .A(n71), .Z(n4896) );
  XNOR U5101 ( .A(n4904), .B(n5118), .Z(n4897) );
  XNOR U5102 ( .A(n4903), .B(n4901), .Z(n5118) );
  AND U5103 ( .A(n5119), .B(n5120), .Z(n4901) );
  NANDN U5104 ( .A(n5121), .B(n5122), .Z(n5120) );
  NANDN U5105 ( .A(n5123), .B(n5124), .Z(n5122) );
  NANDN U5106 ( .A(n5124), .B(n5123), .Z(n5119) );
  ANDN U5107 ( .B(B[53]), .A(n72), .Z(n4903) );
  XNOR U5108 ( .A(n4911), .B(n5125), .Z(n4904) );
  XNOR U5109 ( .A(n4910), .B(n4908), .Z(n5125) );
  AND U5110 ( .A(n5126), .B(n5127), .Z(n4908) );
  NANDN U5111 ( .A(n5128), .B(n5129), .Z(n5127) );
  OR U5112 ( .A(n5130), .B(n5131), .Z(n5129) );
  NAND U5113 ( .A(n5131), .B(n5130), .Z(n5126) );
  ANDN U5114 ( .B(B[54]), .A(n73), .Z(n4910) );
  XNOR U5115 ( .A(n4918), .B(n5132), .Z(n4911) );
  XNOR U5116 ( .A(n4917), .B(n4915), .Z(n5132) );
  AND U5117 ( .A(n5133), .B(n5134), .Z(n4915) );
  NANDN U5118 ( .A(n5135), .B(n5136), .Z(n5134) );
  NANDN U5119 ( .A(n5137), .B(n5138), .Z(n5136) );
  NANDN U5120 ( .A(n5138), .B(n5137), .Z(n5133) );
  ANDN U5121 ( .B(B[55]), .A(n74), .Z(n4917) );
  XNOR U5122 ( .A(n4925), .B(n5139), .Z(n4918) );
  XNOR U5123 ( .A(n4924), .B(n4922), .Z(n5139) );
  AND U5124 ( .A(n5140), .B(n5141), .Z(n4922) );
  NANDN U5125 ( .A(n5142), .B(n5143), .Z(n5141) );
  OR U5126 ( .A(n5144), .B(n5145), .Z(n5143) );
  NAND U5127 ( .A(n5145), .B(n5144), .Z(n5140) );
  ANDN U5128 ( .B(B[56]), .A(n75), .Z(n4924) );
  XNOR U5129 ( .A(n4932), .B(n5146), .Z(n4925) );
  XNOR U5130 ( .A(n4931), .B(n4929), .Z(n5146) );
  AND U5131 ( .A(n5147), .B(n5148), .Z(n4929) );
  NANDN U5132 ( .A(n5149), .B(n5150), .Z(n5148) );
  NANDN U5133 ( .A(n5151), .B(n5152), .Z(n5150) );
  NANDN U5134 ( .A(n5152), .B(n5151), .Z(n5147) );
  ANDN U5135 ( .B(B[57]), .A(n76), .Z(n4931) );
  XNOR U5136 ( .A(n4939), .B(n5153), .Z(n4932) );
  XNOR U5137 ( .A(n4938), .B(n4936), .Z(n5153) );
  AND U5138 ( .A(n5154), .B(n5155), .Z(n4936) );
  NANDN U5139 ( .A(n5156), .B(n5157), .Z(n5155) );
  OR U5140 ( .A(n5158), .B(n5159), .Z(n5157) );
  NAND U5141 ( .A(n5159), .B(n5158), .Z(n5154) );
  ANDN U5142 ( .B(B[58]), .A(n77), .Z(n4938) );
  XNOR U5143 ( .A(n4946), .B(n5160), .Z(n4939) );
  XNOR U5144 ( .A(n4945), .B(n4943), .Z(n5160) );
  AND U5145 ( .A(n5161), .B(n5162), .Z(n4943) );
  NANDN U5146 ( .A(n5163), .B(n5164), .Z(n5162) );
  NANDN U5147 ( .A(n5165), .B(n5166), .Z(n5164) );
  NANDN U5148 ( .A(n5166), .B(n5165), .Z(n5161) );
  ANDN U5149 ( .B(B[59]), .A(n78), .Z(n4945) );
  XNOR U5150 ( .A(n4953), .B(n5167), .Z(n4946) );
  XNOR U5151 ( .A(n4952), .B(n4950), .Z(n5167) );
  AND U5152 ( .A(n5168), .B(n5169), .Z(n4950) );
  NANDN U5153 ( .A(n5170), .B(n5171), .Z(n5169) );
  OR U5154 ( .A(n5172), .B(n5173), .Z(n5171) );
  NAND U5155 ( .A(n5173), .B(n5172), .Z(n5168) );
  ANDN U5156 ( .B(B[60]), .A(n79), .Z(n4952) );
  XNOR U5157 ( .A(n4960), .B(n5174), .Z(n4953) );
  XNOR U5158 ( .A(n4959), .B(n4957), .Z(n5174) );
  AND U5159 ( .A(n5175), .B(n5176), .Z(n4957) );
  NANDN U5160 ( .A(n5177), .B(n5178), .Z(n5176) );
  NANDN U5161 ( .A(n5179), .B(n5180), .Z(n5178) );
  NANDN U5162 ( .A(n5180), .B(n5179), .Z(n5175) );
  ANDN U5163 ( .B(B[61]), .A(n80), .Z(n4959) );
  XNOR U5164 ( .A(n4967), .B(n5181), .Z(n4960) );
  XNOR U5165 ( .A(n4966), .B(n4964), .Z(n5181) );
  AND U5166 ( .A(n5182), .B(n5183), .Z(n4964) );
  NANDN U5167 ( .A(n5184), .B(n5185), .Z(n5183) );
  OR U5168 ( .A(n5186), .B(n5187), .Z(n5185) );
  NAND U5169 ( .A(n5187), .B(n5186), .Z(n5182) );
  ANDN U5170 ( .B(B[62]), .A(n81), .Z(n4966) );
  XNOR U5171 ( .A(n4974), .B(n5188), .Z(n4967) );
  XNOR U5172 ( .A(n4973), .B(n4971), .Z(n5188) );
  AND U5173 ( .A(n5189), .B(n5190), .Z(n4971) );
  NANDN U5174 ( .A(n5191), .B(n5192), .Z(n5190) );
  NAND U5175 ( .A(n5193), .B(n5194), .Z(n5192) );
  ANDN U5176 ( .B(B[63]), .A(n82), .Z(n4973) );
  XOR U5177 ( .A(n4980), .B(n5195), .Z(n4974) );
  XNOR U5178 ( .A(n4978), .B(n4981), .Z(n5195) );
  NAND U5179 ( .A(A[2]), .B(B[64]), .Z(n4981) );
  NANDN U5180 ( .A(n5196), .B(n5197), .Z(n4978) );
  AND U5181 ( .A(A[0]), .B(B[65]), .Z(n5197) );
  XNOR U5182 ( .A(n4983), .B(n5198), .Z(n4980) );
  NAND U5183 ( .A(A[0]), .B(B[66]), .Z(n5198) );
  NAND U5184 ( .A(B[65]), .B(A[1]), .Z(n4983) );
  NAND U5185 ( .A(n5199), .B(n5200), .Z(n155) );
  NANDN U5186 ( .A(n5201), .B(n5202), .Z(n5200) );
  OR U5187 ( .A(n5203), .B(n5204), .Z(n5202) );
  NAND U5188 ( .A(n5204), .B(n5203), .Z(n5199) );
  XOR U5189 ( .A(n157), .B(n156), .Z(\A1[63] ) );
  XOR U5190 ( .A(n5204), .B(n5205), .Z(n156) );
  XNOR U5191 ( .A(n5203), .B(n5201), .Z(n5205) );
  AND U5192 ( .A(n5206), .B(n5207), .Z(n5201) );
  NANDN U5193 ( .A(n5208), .B(n5209), .Z(n5207) );
  NANDN U5194 ( .A(n5210), .B(n5211), .Z(n5209) );
  NANDN U5195 ( .A(n5211), .B(n5210), .Z(n5206) );
  ANDN U5196 ( .B(B[34]), .A(n54), .Z(n5203) );
  XNOR U5197 ( .A(n4998), .B(n5212), .Z(n5204) );
  XNOR U5198 ( .A(n4997), .B(n4995), .Z(n5212) );
  AND U5199 ( .A(n5213), .B(n5214), .Z(n4995) );
  NANDN U5200 ( .A(n5215), .B(n5216), .Z(n5214) );
  OR U5201 ( .A(n5217), .B(n5218), .Z(n5216) );
  NAND U5202 ( .A(n5218), .B(n5217), .Z(n5213) );
  ANDN U5203 ( .B(B[35]), .A(n55), .Z(n4997) );
  XNOR U5204 ( .A(n5005), .B(n5219), .Z(n4998) );
  XNOR U5205 ( .A(n5004), .B(n5002), .Z(n5219) );
  AND U5206 ( .A(n5220), .B(n5221), .Z(n5002) );
  NANDN U5207 ( .A(n5222), .B(n5223), .Z(n5221) );
  NANDN U5208 ( .A(n5224), .B(n5225), .Z(n5223) );
  NANDN U5209 ( .A(n5225), .B(n5224), .Z(n5220) );
  ANDN U5210 ( .B(B[36]), .A(n56), .Z(n5004) );
  XNOR U5211 ( .A(n5012), .B(n5226), .Z(n5005) );
  XNOR U5212 ( .A(n5011), .B(n5009), .Z(n5226) );
  AND U5213 ( .A(n5227), .B(n5228), .Z(n5009) );
  NANDN U5214 ( .A(n5229), .B(n5230), .Z(n5228) );
  OR U5215 ( .A(n5231), .B(n5232), .Z(n5230) );
  NAND U5216 ( .A(n5232), .B(n5231), .Z(n5227) );
  ANDN U5217 ( .B(B[37]), .A(n57), .Z(n5011) );
  XNOR U5218 ( .A(n5019), .B(n5233), .Z(n5012) );
  XNOR U5219 ( .A(n5018), .B(n5016), .Z(n5233) );
  AND U5220 ( .A(n5234), .B(n5235), .Z(n5016) );
  NANDN U5221 ( .A(n5236), .B(n5237), .Z(n5235) );
  NANDN U5222 ( .A(n5238), .B(n5239), .Z(n5237) );
  NANDN U5223 ( .A(n5239), .B(n5238), .Z(n5234) );
  ANDN U5224 ( .B(B[38]), .A(n58), .Z(n5018) );
  XNOR U5225 ( .A(n5026), .B(n5240), .Z(n5019) );
  XNOR U5226 ( .A(n5025), .B(n5023), .Z(n5240) );
  AND U5227 ( .A(n5241), .B(n5242), .Z(n5023) );
  NANDN U5228 ( .A(n5243), .B(n5244), .Z(n5242) );
  OR U5229 ( .A(n5245), .B(n5246), .Z(n5244) );
  NAND U5230 ( .A(n5246), .B(n5245), .Z(n5241) );
  ANDN U5231 ( .B(B[39]), .A(n59), .Z(n5025) );
  XNOR U5232 ( .A(n5033), .B(n5247), .Z(n5026) );
  XNOR U5233 ( .A(n5032), .B(n5030), .Z(n5247) );
  AND U5234 ( .A(n5248), .B(n5249), .Z(n5030) );
  NANDN U5235 ( .A(n5250), .B(n5251), .Z(n5249) );
  NANDN U5236 ( .A(n5252), .B(n5253), .Z(n5251) );
  NANDN U5237 ( .A(n5253), .B(n5252), .Z(n5248) );
  ANDN U5238 ( .B(B[40]), .A(n60), .Z(n5032) );
  XNOR U5239 ( .A(n5040), .B(n5254), .Z(n5033) );
  XNOR U5240 ( .A(n5039), .B(n5037), .Z(n5254) );
  AND U5241 ( .A(n5255), .B(n5256), .Z(n5037) );
  NANDN U5242 ( .A(n5257), .B(n5258), .Z(n5256) );
  OR U5243 ( .A(n5259), .B(n5260), .Z(n5258) );
  NAND U5244 ( .A(n5260), .B(n5259), .Z(n5255) );
  ANDN U5245 ( .B(B[41]), .A(n61), .Z(n5039) );
  XNOR U5246 ( .A(n5047), .B(n5261), .Z(n5040) );
  XNOR U5247 ( .A(n5046), .B(n5044), .Z(n5261) );
  AND U5248 ( .A(n5262), .B(n5263), .Z(n5044) );
  NANDN U5249 ( .A(n5264), .B(n5265), .Z(n5263) );
  NANDN U5250 ( .A(n5266), .B(n5267), .Z(n5265) );
  NANDN U5251 ( .A(n5267), .B(n5266), .Z(n5262) );
  ANDN U5252 ( .B(B[42]), .A(n62), .Z(n5046) );
  XNOR U5253 ( .A(n5054), .B(n5268), .Z(n5047) );
  XNOR U5254 ( .A(n5053), .B(n5051), .Z(n5268) );
  AND U5255 ( .A(n5269), .B(n5270), .Z(n5051) );
  NANDN U5256 ( .A(n5271), .B(n5272), .Z(n5270) );
  OR U5257 ( .A(n5273), .B(n5274), .Z(n5272) );
  NAND U5258 ( .A(n5274), .B(n5273), .Z(n5269) );
  ANDN U5259 ( .B(B[43]), .A(n63), .Z(n5053) );
  XNOR U5260 ( .A(n5061), .B(n5275), .Z(n5054) );
  XNOR U5261 ( .A(n5060), .B(n5058), .Z(n5275) );
  AND U5262 ( .A(n5276), .B(n5277), .Z(n5058) );
  NANDN U5263 ( .A(n5278), .B(n5279), .Z(n5277) );
  NANDN U5264 ( .A(n5280), .B(n5281), .Z(n5279) );
  NANDN U5265 ( .A(n5281), .B(n5280), .Z(n5276) );
  ANDN U5266 ( .B(B[44]), .A(n64), .Z(n5060) );
  XNOR U5267 ( .A(n5068), .B(n5282), .Z(n5061) );
  XNOR U5268 ( .A(n5067), .B(n5065), .Z(n5282) );
  AND U5269 ( .A(n5283), .B(n5284), .Z(n5065) );
  NANDN U5270 ( .A(n5285), .B(n5286), .Z(n5284) );
  OR U5271 ( .A(n5287), .B(n5288), .Z(n5286) );
  NAND U5272 ( .A(n5288), .B(n5287), .Z(n5283) );
  ANDN U5273 ( .B(B[45]), .A(n65), .Z(n5067) );
  XNOR U5274 ( .A(n5075), .B(n5289), .Z(n5068) );
  XNOR U5275 ( .A(n5074), .B(n5072), .Z(n5289) );
  AND U5276 ( .A(n5290), .B(n5291), .Z(n5072) );
  NANDN U5277 ( .A(n5292), .B(n5293), .Z(n5291) );
  NANDN U5278 ( .A(n5294), .B(n5295), .Z(n5293) );
  NANDN U5279 ( .A(n5295), .B(n5294), .Z(n5290) );
  ANDN U5280 ( .B(B[46]), .A(n66), .Z(n5074) );
  XNOR U5281 ( .A(n5082), .B(n5296), .Z(n5075) );
  XNOR U5282 ( .A(n5081), .B(n5079), .Z(n5296) );
  AND U5283 ( .A(n5297), .B(n5298), .Z(n5079) );
  NANDN U5284 ( .A(n5299), .B(n5300), .Z(n5298) );
  OR U5285 ( .A(n5301), .B(n5302), .Z(n5300) );
  NAND U5286 ( .A(n5302), .B(n5301), .Z(n5297) );
  ANDN U5287 ( .B(B[47]), .A(n67), .Z(n5081) );
  XNOR U5288 ( .A(n5089), .B(n5303), .Z(n5082) );
  XNOR U5289 ( .A(n5088), .B(n5086), .Z(n5303) );
  AND U5290 ( .A(n5304), .B(n5305), .Z(n5086) );
  NANDN U5291 ( .A(n5306), .B(n5307), .Z(n5305) );
  NANDN U5292 ( .A(n5308), .B(n5309), .Z(n5307) );
  NANDN U5293 ( .A(n5309), .B(n5308), .Z(n5304) );
  ANDN U5294 ( .B(B[48]), .A(n68), .Z(n5088) );
  XNOR U5295 ( .A(n5096), .B(n5310), .Z(n5089) );
  XNOR U5296 ( .A(n5095), .B(n5093), .Z(n5310) );
  AND U5297 ( .A(n5311), .B(n5312), .Z(n5093) );
  NANDN U5298 ( .A(n5313), .B(n5314), .Z(n5312) );
  OR U5299 ( .A(n5315), .B(n5316), .Z(n5314) );
  NAND U5300 ( .A(n5316), .B(n5315), .Z(n5311) );
  ANDN U5301 ( .B(B[49]), .A(n69), .Z(n5095) );
  XNOR U5302 ( .A(n5103), .B(n5317), .Z(n5096) );
  XNOR U5303 ( .A(n5102), .B(n5100), .Z(n5317) );
  AND U5304 ( .A(n5318), .B(n5319), .Z(n5100) );
  NANDN U5305 ( .A(n5320), .B(n5321), .Z(n5319) );
  NANDN U5306 ( .A(n5322), .B(n5323), .Z(n5321) );
  NANDN U5307 ( .A(n5323), .B(n5322), .Z(n5318) );
  ANDN U5308 ( .B(B[50]), .A(n70), .Z(n5102) );
  XNOR U5309 ( .A(n5110), .B(n5324), .Z(n5103) );
  XNOR U5310 ( .A(n5109), .B(n5107), .Z(n5324) );
  AND U5311 ( .A(n5325), .B(n5326), .Z(n5107) );
  NANDN U5312 ( .A(n5327), .B(n5328), .Z(n5326) );
  OR U5313 ( .A(n5329), .B(n5330), .Z(n5328) );
  NAND U5314 ( .A(n5330), .B(n5329), .Z(n5325) );
  ANDN U5315 ( .B(B[51]), .A(n71), .Z(n5109) );
  XNOR U5316 ( .A(n5117), .B(n5331), .Z(n5110) );
  XNOR U5317 ( .A(n5116), .B(n5114), .Z(n5331) );
  AND U5318 ( .A(n5332), .B(n5333), .Z(n5114) );
  NANDN U5319 ( .A(n5334), .B(n5335), .Z(n5333) );
  NANDN U5320 ( .A(n5336), .B(n5337), .Z(n5335) );
  NANDN U5321 ( .A(n5337), .B(n5336), .Z(n5332) );
  ANDN U5322 ( .B(B[52]), .A(n72), .Z(n5116) );
  XNOR U5323 ( .A(n5124), .B(n5338), .Z(n5117) );
  XNOR U5324 ( .A(n5123), .B(n5121), .Z(n5338) );
  AND U5325 ( .A(n5339), .B(n5340), .Z(n5121) );
  NANDN U5326 ( .A(n5341), .B(n5342), .Z(n5340) );
  OR U5327 ( .A(n5343), .B(n5344), .Z(n5342) );
  NAND U5328 ( .A(n5344), .B(n5343), .Z(n5339) );
  ANDN U5329 ( .B(B[53]), .A(n73), .Z(n5123) );
  XNOR U5330 ( .A(n5131), .B(n5345), .Z(n5124) );
  XNOR U5331 ( .A(n5130), .B(n5128), .Z(n5345) );
  AND U5332 ( .A(n5346), .B(n5347), .Z(n5128) );
  NANDN U5333 ( .A(n5348), .B(n5349), .Z(n5347) );
  NANDN U5334 ( .A(n5350), .B(n5351), .Z(n5349) );
  NANDN U5335 ( .A(n5351), .B(n5350), .Z(n5346) );
  ANDN U5336 ( .B(B[54]), .A(n74), .Z(n5130) );
  XNOR U5337 ( .A(n5138), .B(n5352), .Z(n5131) );
  XNOR U5338 ( .A(n5137), .B(n5135), .Z(n5352) );
  AND U5339 ( .A(n5353), .B(n5354), .Z(n5135) );
  NANDN U5340 ( .A(n5355), .B(n5356), .Z(n5354) );
  OR U5341 ( .A(n5357), .B(n5358), .Z(n5356) );
  NAND U5342 ( .A(n5358), .B(n5357), .Z(n5353) );
  ANDN U5343 ( .B(B[55]), .A(n75), .Z(n5137) );
  XNOR U5344 ( .A(n5145), .B(n5359), .Z(n5138) );
  XNOR U5345 ( .A(n5144), .B(n5142), .Z(n5359) );
  AND U5346 ( .A(n5360), .B(n5361), .Z(n5142) );
  NANDN U5347 ( .A(n5362), .B(n5363), .Z(n5361) );
  NANDN U5348 ( .A(n5364), .B(n5365), .Z(n5363) );
  NANDN U5349 ( .A(n5365), .B(n5364), .Z(n5360) );
  ANDN U5350 ( .B(B[56]), .A(n76), .Z(n5144) );
  XNOR U5351 ( .A(n5152), .B(n5366), .Z(n5145) );
  XNOR U5352 ( .A(n5151), .B(n5149), .Z(n5366) );
  AND U5353 ( .A(n5367), .B(n5368), .Z(n5149) );
  NANDN U5354 ( .A(n5369), .B(n5370), .Z(n5368) );
  OR U5355 ( .A(n5371), .B(n5372), .Z(n5370) );
  NAND U5356 ( .A(n5372), .B(n5371), .Z(n5367) );
  ANDN U5357 ( .B(B[57]), .A(n77), .Z(n5151) );
  XNOR U5358 ( .A(n5159), .B(n5373), .Z(n5152) );
  XNOR U5359 ( .A(n5158), .B(n5156), .Z(n5373) );
  AND U5360 ( .A(n5374), .B(n5375), .Z(n5156) );
  NANDN U5361 ( .A(n5376), .B(n5377), .Z(n5375) );
  NANDN U5362 ( .A(n5378), .B(n5379), .Z(n5377) );
  NANDN U5363 ( .A(n5379), .B(n5378), .Z(n5374) );
  ANDN U5364 ( .B(B[58]), .A(n78), .Z(n5158) );
  XNOR U5365 ( .A(n5166), .B(n5380), .Z(n5159) );
  XNOR U5366 ( .A(n5165), .B(n5163), .Z(n5380) );
  AND U5367 ( .A(n5381), .B(n5382), .Z(n5163) );
  NANDN U5368 ( .A(n5383), .B(n5384), .Z(n5382) );
  OR U5369 ( .A(n5385), .B(n5386), .Z(n5384) );
  NAND U5370 ( .A(n5386), .B(n5385), .Z(n5381) );
  ANDN U5371 ( .B(B[59]), .A(n79), .Z(n5165) );
  XNOR U5372 ( .A(n5173), .B(n5387), .Z(n5166) );
  XNOR U5373 ( .A(n5172), .B(n5170), .Z(n5387) );
  AND U5374 ( .A(n5388), .B(n5389), .Z(n5170) );
  NANDN U5375 ( .A(n5390), .B(n5391), .Z(n5389) );
  NANDN U5376 ( .A(n5392), .B(n5393), .Z(n5391) );
  NANDN U5377 ( .A(n5393), .B(n5392), .Z(n5388) );
  ANDN U5378 ( .B(B[60]), .A(n80), .Z(n5172) );
  XNOR U5379 ( .A(n5180), .B(n5394), .Z(n5173) );
  XNOR U5380 ( .A(n5179), .B(n5177), .Z(n5394) );
  AND U5381 ( .A(n5395), .B(n5396), .Z(n5177) );
  NANDN U5382 ( .A(n5397), .B(n5398), .Z(n5396) );
  OR U5383 ( .A(n5399), .B(n5400), .Z(n5398) );
  NAND U5384 ( .A(n5400), .B(n5399), .Z(n5395) );
  ANDN U5385 ( .B(B[61]), .A(n81), .Z(n5179) );
  XNOR U5386 ( .A(n5187), .B(n5401), .Z(n5180) );
  XNOR U5387 ( .A(n5186), .B(n5184), .Z(n5401) );
  AND U5388 ( .A(n5402), .B(n5403), .Z(n5184) );
  NANDN U5389 ( .A(n5404), .B(n5405), .Z(n5403) );
  NAND U5390 ( .A(n5406), .B(n5407), .Z(n5405) );
  ANDN U5391 ( .B(B[62]), .A(n82), .Z(n5186) );
  XOR U5392 ( .A(n5193), .B(n5408), .Z(n5187) );
  XNOR U5393 ( .A(n5191), .B(n5194), .Z(n5408) );
  NAND U5394 ( .A(A[2]), .B(B[63]), .Z(n5194) );
  NANDN U5395 ( .A(n5409), .B(n5410), .Z(n5191) );
  AND U5396 ( .A(A[0]), .B(B[64]), .Z(n5410) );
  XNOR U5397 ( .A(n5196), .B(n5411), .Z(n5193) );
  NAND U5398 ( .A(A[0]), .B(B[65]), .Z(n5411) );
  NAND U5399 ( .A(B[64]), .B(A[1]), .Z(n5196) );
  NAND U5400 ( .A(n5412), .B(n5413), .Z(n157) );
  NANDN U5401 ( .A(n5414), .B(n5415), .Z(n5413) );
  OR U5402 ( .A(n5416), .B(n5417), .Z(n5415) );
  NAND U5403 ( .A(n5417), .B(n5416), .Z(n5412) );
  XOR U5404 ( .A(n159), .B(n158), .Z(\A1[62] ) );
  XOR U5405 ( .A(n5417), .B(n5418), .Z(n158) );
  XNOR U5406 ( .A(n5416), .B(n5414), .Z(n5418) );
  AND U5407 ( .A(n5419), .B(n5420), .Z(n5414) );
  NANDN U5408 ( .A(n5421), .B(n5422), .Z(n5420) );
  NANDN U5409 ( .A(n5423), .B(n5424), .Z(n5422) );
  NANDN U5410 ( .A(n5424), .B(n5423), .Z(n5419) );
  ANDN U5411 ( .B(B[33]), .A(n54), .Z(n5416) );
  XNOR U5412 ( .A(n5211), .B(n5425), .Z(n5417) );
  XNOR U5413 ( .A(n5210), .B(n5208), .Z(n5425) );
  AND U5414 ( .A(n5426), .B(n5427), .Z(n5208) );
  NANDN U5415 ( .A(n5428), .B(n5429), .Z(n5427) );
  OR U5416 ( .A(n5430), .B(n5431), .Z(n5429) );
  NAND U5417 ( .A(n5431), .B(n5430), .Z(n5426) );
  ANDN U5418 ( .B(B[34]), .A(n55), .Z(n5210) );
  XNOR U5419 ( .A(n5218), .B(n5432), .Z(n5211) );
  XNOR U5420 ( .A(n5217), .B(n5215), .Z(n5432) );
  AND U5421 ( .A(n5433), .B(n5434), .Z(n5215) );
  NANDN U5422 ( .A(n5435), .B(n5436), .Z(n5434) );
  NANDN U5423 ( .A(n5437), .B(n5438), .Z(n5436) );
  NANDN U5424 ( .A(n5438), .B(n5437), .Z(n5433) );
  ANDN U5425 ( .B(B[35]), .A(n56), .Z(n5217) );
  XNOR U5426 ( .A(n5225), .B(n5439), .Z(n5218) );
  XNOR U5427 ( .A(n5224), .B(n5222), .Z(n5439) );
  AND U5428 ( .A(n5440), .B(n5441), .Z(n5222) );
  NANDN U5429 ( .A(n5442), .B(n5443), .Z(n5441) );
  OR U5430 ( .A(n5444), .B(n5445), .Z(n5443) );
  NAND U5431 ( .A(n5445), .B(n5444), .Z(n5440) );
  ANDN U5432 ( .B(B[36]), .A(n57), .Z(n5224) );
  XNOR U5433 ( .A(n5232), .B(n5446), .Z(n5225) );
  XNOR U5434 ( .A(n5231), .B(n5229), .Z(n5446) );
  AND U5435 ( .A(n5447), .B(n5448), .Z(n5229) );
  NANDN U5436 ( .A(n5449), .B(n5450), .Z(n5448) );
  NANDN U5437 ( .A(n5451), .B(n5452), .Z(n5450) );
  NANDN U5438 ( .A(n5452), .B(n5451), .Z(n5447) );
  ANDN U5439 ( .B(B[37]), .A(n58), .Z(n5231) );
  XNOR U5440 ( .A(n5239), .B(n5453), .Z(n5232) );
  XNOR U5441 ( .A(n5238), .B(n5236), .Z(n5453) );
  AND U5442 ( .A(n5454), .B(n5455), .Z(n5236) );
  NANDN U5443 ( .A(n5456), .B(n5457), .Z(n5455) );
  OR U5444 ( .A(n5458), .B(n5459), .Z(n5457) );
  NAND U5445 ( .A(n5459), .B(n5458), .Z(n5454) );
  ANDN U5446 ( .B(B[38]), .A(n59), .Z(n5238) );
  XNOR U5447 ( .A(n5246), .B(n5460), .Z(n5239) );
  XNOR U5448 ( .A(n5245), .B(n5243), .Z(n5460) );
  AND U5449 ( .A(n5461), .B(n5462), .Z(n5243) );
  NANDN U5450 ( .A(n5463), .B(n5464), .Z(n5462) );
  NANDN U5451 ( .A(n5465), .B(n5466), .Z(n5464) );
  NANDN U5452 ( .A(n5466), .B(n5465), .Z(n5461) );
  ANDN U5453 ( .B(B[39]), .A(n60), .Z(n5245) );
  XNOR U5454 ( .A(n5253), .B(n5467), .Z(n5246) );
  XNOR U5455 ( .A(n5252), .B(n5250), .Z(n5467) );
  AND U5456 ( .A(n5468), .B(n5469), .Z(n5250) );
  NANDN U5457 ( .A(n5470), .B(n5471), .Z(n5469) );
  OR U5458 ( .A(n5472), .B(n5473), .Z(n5471) );
  NAND U5459 ( .A(n5473), .B(n5472), .Z(n5468) );
  ANDN U5460 ( .B(B[40]), .A(n61), .Z(n5252) );
  XNOR U5461 ( .A(n5260), .B(n5474), .Z(n5253) );
  XNOR U5462 ( .A(n5259), .B(n5257), .Z(n5474) );
  AND U5463 ( .A(n5475), .B(n5476), .Z(n5257) );
  NANDN U5464 ( .A(n5477), .B(n5478), .Z(n5476) );
  NANDN U5465 ( .A(n5479), .B(n5480), .Z(n5478) );
  NANDN U5466 ( .A(n5480), .B(n5479), .Z(n5475) );
  ANDN U5467 ( .B(B[41]), .A(n62), .Z(n5259) );
  XNOR U5468 ( .A(n5267), .B(n5481), .Z(n5260) );
  XNOR U5469 ( .A(n5266), .B(n5264), .Z(n5481) );
  AND U5470 ( .A(n5482), .B(n5483), .Z(n5264) );
  NANDN U5471 ( .A(n5484), .B(n5485), .Z(n5483) );
  OR U5472 ( .A(n5486), .B(n5487), .Z(n5485) );
  NAND U5473 ( .A(n5487), .B(n5486), .Z(n5482) );
  ANDN U5474 ( .B(B[42]), .A(n63), .Z(n5266) );
  XNOR U5475 ( .A(n5274), .B(n5488), .Z(n5267) );
  XNOR U5476 ( .A(n5273), .B(n5271), .Z(n5488) );
  AND U5477 ( .A(n5489), .B(n5490), .Z(n5271) );
  NANDN U5478 ( .A(n5491), .B(n5492), .Z(n5490) );
  NANDN U5479 ( .A(n5493), .B(n5494), .Z(n5492) );
  NANDN U5480 ( .A(n5494), .B(n5493), .Z(n5489) );
  ANDN U5481 ( .B(B[43]), .A(n64), .Z(n5273) );
  XNOR U5482 ( .A(n5281), .B(n5495), .Z(n5274) );
  XNOR U5483 ( .A(n5280), .B(n5278), .Z(n5495) );
  AND U5484 ( .A(n5496), .B(n5497), .Z(n5278) );
  NANDN U5485 ( .A(n5498), .B(n5499), .Z(n5497) );
  OR U5486 ( .A(n5500), .B(n5501), .Z(n5499) );
  NAND U5487 ( .A(n5501), .B(n5500), .Z(n5496) );
  ANDN U5488 ( .B(B[44]), .A(n65), .Z(n5280) );
  XNOR U5489 ( .A(n5288), .B(n5502), .Z(n5281) );
  XNOR U5490 ( .A(n5287), .B(n5285), .Z(n5502) );
  AND U5491 ( .A(n5503), .B(n5504), .Z(n5285) );
  NANDN U5492 ( .A(n5505), .B(n5506), .Z(n5504) );
  NANDN U5493 ( .A(n5507), .B(n5508), .Z(n5506) );
  NANDN U5494 ( .A(n5508), .B(n5507), .Z(n5503) );
  ANDN U5495 ( .B(B[45]), .A(n66), .Z(n5287) );
  XNOR U5496 ( .A(n5295), .B(n5509), .Z(n5288) );
  XNOR U5497 ( .A(n5294), .B(n5292), .Z(n5509) );
  AND U5498 ( .A(n5510), .B(n5511), .Z(n5292) );
  NANDN U5499 ( .A(n5512), .B(n5513), .Z(n5511) );
  OR U5500 ( .A(n5514), .B(n5515), .Z(n5513) );
  NAND U5501 ( .A(n5515), .B(n5514), .Z(n5510) );
  ANDN U5502 ( .B(B[46]), .A(n67), .Z(n5294) );
  XNOR U5503 ( .A(n5302), .B(n5516), .Z(n5295) );
  XNOR U5504 ( .A(n5301), .B(n5299), .Z(n5516) );
  AND U5505 ( .A(n5517), .B(n5518), .Z(n5299) );
  NANDN U5506 ( .A(n5519), .B(n5520), .Z(n5518) );
  NANDN U5507 ( .A(n5521), .B(n5522), .Z(n5520) );
  NANDN U5508 ( .A(n5522), .B(n5521), .Z(n5517) );
  ANDN U5509 ( .B(B[47]), .A(n68), .Z(n5301) );
  XNOR U5510 ( .A(n5309), .B(n5523), .Z(n5302) );
  XNOR U5511 ( .A(n5308), .B(n5306), .Z(n5523) );
  AND U5512 ( .A(n5524), .B(n5525), .Z(n5306) );
  NANDN U5513 ( .A(n5526), .B(n5527), .Z(n5525) );
  OR U5514 ( .A(n5528), .B(n5529), .Z(n5527) );
  NAND U5515 ( .A(n5529), .B(n5528), .Z(n5524) );
  ANDN U5516 ( .B(B[48]), .A(n69), .Z(n5308) );
  XNOR U5517 ( .A(n5316), .B(n5530), .Z(n5309) );
  XNOR U5518 ( .A(n5315), .B(n5313), .Z(n5530) );
  AND U5519 ( .A(n5531), .B(n5532), .Z(n5313) );
  NANDN U5520 ( .A(n5533), .B(n5534), .Z(n5532) );
  NANDN U5521 ( .A(n5535), .B(n5536), .Z(n5534) );
  NANDN U5522 ( .A(n5536), .B(n5535), .Z(n5531) );
  ANDN U5523 ( .B(B[49]), .A(n70), .Z(n5315) );
  XNOR U5524 ( .A(n5323), .B(n5537), .Z(n5316) );
  XNOR U5525 ( .A(n5322), .B(n5320), .Z(n5537) );
  AND U5526 ( .A(n5538), .B(n5539), .Z(n5320) );
  NANDN U5527 ( .A(n5540), .B(n5541), .Z(n5539) );
  OR U5528 ( .A(n5542), .B(n5543), .Z(n5541) );
  NAND U5529 ( .A(n5543), .B(n5542), .Z(n5538) );
  ANDN U5530 ( .B(B[50]), .A(n71), .Z(n5322) );
  XNOR U5531 ( .A(n5330), .B(n5544), .Z(n5323) );
  XNOR U5532 ( .A(n5329), .B(n5327), .Z(n5544) );
  AND U5533 ( .A(n5545), .B(n5546), .Z(n5327) );
  NANDN U5534 ( .A(n5547), .B(n5548), .Z(n5546) );
  NANDN U5535 ( .A(n5549), .B(n5550), .Z(n5548) );
  NANDN U5536 ( .A(n5550), .B(n5549), .Z(n5545) );
  ANDN U5537 ( .B(B[51]), .A(n72), .Z(n5329) );
  XNOR U5538 ( .A(n5337), .B(n5551), .Z(n5330) );
  XNOR U5539 ( .A(n5336), .B(n5334), .Z(n5551) );
  AND U5540 ( .A(n5552), .B(n5553), .Z(n5334) );
  NANDN U5541 ( .A(n5554), .B(n5555), .Z(n5553) );
  OR U5542 ( .A(n5556), .B(n5557), .Z(n5555) );
  NAND U5543 ( .A(n5557), .B(n5556), .Z(n5552) );
  ANDN U5544 ( .B(B[52]), .A(n73), .Z(n5336) );
  XNOR U5545 ( .A(n5344), .B(n5558), .Z(n5337) );
  XNOR U5546 ( .A(n5343), .B(n5341), .Z(n5558) );
  AND U5547 ( .A(n5559), .B(n5560), .Z(n5341) );
  NANDN U5548 ( .A(n5561), .B(n5562), .Z(n5560) );
  NANDN U5549 ( .A(n5563), .B(n5564), .Z(n5562) );
  NANDN U5550 ( .A(n5564), .B(n5563), .Z(n5559) );
  ANDN U5551 ( .B(B[53]), .A(n74), .Z(n5343) );
  XNOR U5552 ( .A(n5351), .B(n5565), .Z(n5344) );
  XNOR U5553 ( .A(n5350), .B(n5348), .Z(n5565) );
  AND U5554 ( .A(n5566), .B(n5567), .Z(n5348) );
  NANDN U5555 ( .A(n5568), .B(n5569), .Z(n5567) );
  OR U5556 ( .A(n5570), .B(n5571), .Z(n5569) );
  NAND U5557 ( .A(n5571), .B(n5570), .Z(n5566) );
  ANDN U5558 ( .B(B[54]), .A(n75), .Z(n5350) );
  XNOR U5559 ( .A(n5358), .B(n5572), .Z(n5351) );
  XNOR U5560 ( .A(n5357), .B(n5355), .Z(n5572) );
  AND U5561 ( .A(n5573), .B(n5574), .Z(n5355) );
  NANDN U5562 ( .A(n5575), .B(n5576), .Z(n5574) );
  NANDN U5563 ( .A(n5577), .B(n5578), .Z(n5576) );
  NANDN U5564 ( .A(n5578), .B(n5577), .Z(n5573) );
  ANDN U5565 ( .B(B[55]), .A(n76), .Z(n5357) );
  XNOR U5566 ( .A(n5365), .B(n5579), .Z(n5358) );
  XNOR U5567 ( .A(n5364), .B(n5362), .Z(n5579) );
  AND U5568 ( .A(n5580), .B(n5581), .Z(n5362) );
  NANDN U5569 ( .A(n5582), .B(n5583), .Z(n5581) );
  OR U5570 ( .A(n5584), .B(n5585), .Z(n5583) );
  NAND U5571 ( .A(n5585), .B(n5584), .Z(n5580) );
  ANDN U5572 ( .B(B[56]), .A(n77), .Z(n5364) );
  XNOR U5573 ( .A(n5372), .B(n5586), .Z(n5365) );
  XNOR U5574 ( .A(n5371), .B(n5369), .Z(n5586) );
  AND U5575 ( .A(n5587), .B(n5588), .Z(n5369) );
  NANDN U5576 ( .A(n5589), .B(n5590), .Z(n5588) );
  NANDN U5577 ( .A(n5591), .B(n5592), .Z(n5590) );
  NANDN U5578 ( .A(n5592), .B(n5591), .Z(n5587) );
  ANDN U5579 ( .B(B[57]), .A(n78), .Z(n5371) );
  XNOR U5580 ( .A(n5379), .B(n5593), .Z(n5372) );
  XNOR U5581 ( .A(n5378), .B(n5376), .Z(n5593) );
  AND U5582 ( .A(n5594), .B(n5595), .Z(n5376) );
  NANDN U5583 ( .A(n5596), .B(n5597), .Z(n5595) );
  OR U5584 ( .A(n5598), .B(n5599), .Z(n5597) );
  NAND U5585 ( .A(n5599), .B(n5598), .Z(n5594) );
  ANDN U5586 ( .B(B[58]), .A(n79), .Z(n5378) );
  XNOR U5587 ( .A(n5386), .B(n5600), .Z(n5379) );
  XNOR U5588 ( .A(n5385), .B(n5383), .Z(n5600) );
  AND U5589 ( .A(n5601), .B(n5602), .Z(n5383) );
  NANDN U5590 ( .A(n5603), .B(n5604), .Z(n5602) );
  NANDN U5591 ( .A(n5605), .B(n5606), .Z(n5604) );
  NANDN U5592 ( .A(n5606), .B(n5605), .Z(n5601) );
  ANDN U5593 ( .B(B[59]), .A(n80), .Z(n5385) );
  XNOR U5594 ( .A(n5393), .B(n5607), .Z(n5386) );
  XNOR U5595 ( .A(n5392), .B(n5390), .Z(n5607) );
  AND U5596 ( .A(n5608), .B(n5609), .Z(n5390) );
  NANDN U5597 ( .A(n5610), .B(n5611), .Z(n5609) );
  OR U5598 ( .A(n5612), .B(n5613), .Z(n5611) );
  NAND U5599 ( .A(n5613), .B(n5612), .Z(n5608) );
  ANDN U5600 ( .B(B[60]), .A(n81), .Z(n5392) );
  XNOR U5601 ( .A(n5400), .B(n5614), .Z(n5393) );
  XNOR U5602 ( .A(n5399), .B(n5397), .Z(n5614) );
  AND U5603 ( .A(n5615), .B(n5616), .Z(n5397) );
  NANDN U5604 ( .A(n5617), .B(n5618), .Z(n5616) );
  NAND U5605 ( .A(n5619), .B(n5620), .Z(n5618) );
  ANDN U5606 ( .B(B[61]), .A(n82), .Z(n5399) );
  XOR U5607 ( .A(n5406), .B(n5621), .Z(n5400) );
  XNOR U5608 ( .A(n5404), .B(n5407), .Z(n5621) );
  NAND U5609 ( .A(A[2]), .B(B[62]), .Z(n5407) );
  NANDN U5610 ( .A(n5622), .B(n5623), .Z(n5404) );
  AND U5611 ( .A(A[0]), .B(B[63]), .Z(n5623) );
  XNOR U5612 ( .A(n5409), .B(n5624), .Z(n5406) );
  NAND U5613 ( .A(A[0]), .B(B[64]), .Z(n5624) );
  NAND U5614 ( .A(B[63]), .B(A[1]), .Z(n5409) );
  NAND U5615 ( .A(n5625), .B(n5626), .Z(n159) );
  NANDN U5616 ( .A(n5627), .B(n5628), .Z(n5626) );
  OR U5617 ( .A(n5629), .B(n5630), .Z(n5628) );
  NAND U5618 ( .A(n5630), .B(n5629), .Z(n5625) );
  XOR U5619 ( .A(n161), .B(n160), .Z(\A1[61] ) );
  XOR U5620 ( .A(n5630), .B(n5631), .Z(n160) );
  XNOR U5621 ( .A(n5629), .B(n5627), .Z(n5631) );
  AND U5622 ( .A(n5632), .B(n5633), .Z(n5627) );
  NANDN U5623 ( .A(n5634), .B(n5635), .Z(n5633) );
  NANDN U5624 ( .A(n5636), .B(n5637), .Z(n5635) );
  NANDN U5625 ( .A(n5637), .B(n5636), .Z(n5632) );
  ANDN U5626 ( .B(B[32]), .A(n54), .Z(n5629) );
  XNOR U5627 ( .A(n5424), .B(n5638), .Z(n5630) );
  XNOR U5628 ( .A(n5423), .B(n5421), .Z(n5638) );
  AND U5629 ( .A(n5639), .B(n5640), .Z(n5421) );
  NANDN U5630 ( .A(n5641), .B(n5642), .Z(n5640) );
  OR U5631 ( .A(n5643), .B(n5644), .Z(n5642) );
  NAND U5632 ( .A(n5644), .B(n5643), .Z(n5639) );
  ANDN U5633 ( .B(B[33]), .A(n55), .Z(n5423) );
  XNOR U5634 ( .A(n5431), .B(n5645), .Z(n5424) );
  XNOR U5635 ( .A(n5430), .B(n5428), .Z(n5645) );
  AND U5636 ( .A(n5646), .B(n5647), .Z(n5428) );
  NANDN U5637 ( .A(n5648), .B(n5649), .Z(n5647) );
  NANDN U5638 ( .A(n5650), .B(n5651), .Z(n5649) );
  NANDN U5639 ( .A(n5651), .B(n5650), .Z(n5646) );
  ANDN U5640 ( .B(B[34]), .A(n56), .Z(n5430) );
  XNOR U5641 ( .A(n5438), .B(n5652), .Z(n5431) );
  XNOR U5642 ( .A(n5437), .B(n5435), .Z(n5652) );
  AND U5643 ( .A(n5653), .B(n5654), .Z(n5435) );
  NANDN U5644 ( .A(n5655), .B(n5656), .Z(n5654) );
  OR U5645 ( .A(n5657), .B(n5658), .Z(n5656) );
  NAND U5646 ( .A(n5658), .B(n5657), .Z(n5653) );
  ANDN U5647 ( .B(B[35]), .A(n57), .Z(n5437) );
  XNOR U5648 ( .A(n5445), .B(n5659), .Z(n5438) );
  XNOR U5649 ( .A(n5444), .B(n5442), .Z(n5659) );
  AND U5650 ( .A(n5660), .B(n5661), .Z(n5442) );
  NANDN U5651 ( .A(n5662), .B(n5663), .Z(n5661) );
  NANDN U5652 ( .A(n5664), .B(n5665), .Z(n5663) );
  NANDN U5653 ( .A(n5665), .B(n5664), .Z(n5660) );
  ANDN U5654 ( .B(B[36]), .A(n58), .Z(n5444) );
  XNOR U5655 ( .A(n5452), .B(n5666), .Z(n5445) );
  XNOR U5656 ( .A(n5451), .B(n5449), .Z(n5666) );
  AND U5657 ( .A(n5667), .B(n5668), .Z(n5449) );
  NANDN U5658 ( .A(n5669), .B(n5670), .Z(n5668) );
  OR U5659 ( .A(n5671), .B(n5672), .Z(n5670) );
  NAND U5660 ( .A(n5672), .B(n5671), .Z(n5667) );
  ANDN U5661 ( .B(B[37]), .A(n59), .Z(n5451) );
  XNOR U5662 ( .A(n5459), .B(n5673), .Z(n5452) );
  XNOR U5663 ( .A(n5458), .B(n5456), .Z(n5673) );
  AND U5664 ( .A(n5674), .B(n5675), .Z(n5456) );
  NANDN U5665 ( .A(n5676), .B(n5677), .Z(n5675) );
  NANDN U5666 ( .A(n5678), .B(n5679), .Z(n5677) );
  NANDN U5667 ( .A(n5679), .B(n5678), .Z(n5674) );
  ANDN U5668 ( .B(B[38]), .A(n60), .Z(n5458) );
  XNOR U5669 ( .A(n5466), .B(n5680), .Z(n5459) );
  XNOR U5670 ( .A(n5465), .B(n5463), .Z(n5680) );
  AND U5671 ( .A(n5681), .B(n5682), .Z(n5463) );
  NANDN U5672 ( .A(n5683), .B(n5684), .Z(n5682) );
  OR U5673 ( .A(n5685), .B(n5686), .Z(n5684) );
  NAND U5674 ( .A(n5686), .B(n5685), .Z(n5681) );
  ANDN U5675 ( .B(B[39]), .A(n61), .Z(n5465) );
  XNOR U5676 ( .A(n5473), .B(n5687), .Z(n5466) );
  XNOR U5677 ( .A(n5472), .B(n5470), .Z(n5687) );
  AND U5678 ( .A(n5688), .B(n5689), .Z(n5470) );
  NANDN U5679 ( .A(n5690), .B(n5691), .Z(n5689) );
  NANDN U5680 ( .A(n5692), .B(n5693), .Z(n5691) );
  NANDN U5681 ( .A(n5693), .B(n5692), .Z(n5688) );
  ANDN U5682 ( .B(B[40]), .A(n62), .Z(n5472) );
  XNOR U5683 ( .A(n5480), .B(n5694), .Z(n5473) );
  XNOR U5684 ( .A(n5479), .B(n5477), .Z(n5694) );
  AND U5685 ( .A(n5695), .B(n5696), .Z(n5477) );
  NANDN U5686 ( .A(n5697), .B(n5698), .Z(n5696) );
  OR U5687 ( .A(n5699), .B(n5700), .Z(n5698) );
  NAND U5688 ( .A(n5700), .B(n5699), .Z(n5695) );
  ANDN U5689 ( .B(B[41]), .A(n63), .Z(n5479) );
  XNOR U5690 ( .A(n5487), .B(n5701), .Z(n5480) );
  XNOR U5691 ( .A(n5486), .B(n5484), .Z(n5701) );
  AND U5692 ( .A(n5702), .B(n5703), .Z(n5484) );
  NANDN U5693 ( .A(n5704), .B(n5705), .Z(n5703) );
  NANDN U5694 ( .A(n5706), .B(n5707), .Z(n5705) );
  NANDN U5695 ( .A(n5707), .B(n5706), .Z(n5702) );
  ANDN U5696 ( .B(B[42]), .A(n64), .Z(n5486) );
  XNOR U5697 ( .A(n5494), .B(n5708), .Z(n5487) );
  XNOR U5698 ( .A(n5493), .B(n5491), .Z(n5708) );
  AND U5699 ( .A(n5709), .B(n5710), .Z(n5491) );
  NANDN U5700 ( .A(n5711), .B(n5712), .Z(n5710) );
  OR U5701 ( .A(n5713), .B(n5714), .Z(n5712) );
  NAND U5702 ( .A(n5714), .B(n5713), .Z(n5709) );
  ANDN U5703 ( .B(B[43]), .A(n65), .Z(n5493) );
  XNOR U5704 ( .A(n5501), .B(n5715), .Z(n5494) );
  XNOR U5705 ( .A(n5500), .B(n5498), .Z(n5715) );
  AND U5706 ( .A(n5716), .B(n5717), .Z(n5498) );
  NANDN U5707 ( .A(n5718), .B(n5719), .Z(n5717) );
  NANDN U5708 ( .A(n5720), .B(n5721), .Z(n5719) );
  NANDN U5709 ( .A(n5721), .B(n5720), .Z(n5716) );
  ANDN U5710 ( .B(B[44]), .A(n66), .Z(n5500) );
  XNOR U5711 ( .A(n5508), .B(n5722), .Z(n5501) );
  XNOR U5712 ( .A(n5507), .B(n5505), .Z(n5722) );
  AND U5713 ( .A(n5723), .B(n5724), .Z(n5505) );
  NANDN U5714 ( .A(n5725), .B(n5726), .Z(n5724) );
  OR U5715 ( .A(n5727), .B(n5728), .Z(n5726) );
  NAND U5716 ( .A(n5728), .B(n5727), .Z(n5723) );
  ANDN U5717 ( .B(B[45]), .A(n67), .Z(n5507) );
  XNOR U5718 ( .A(n5515), .B(n5729), .Z(n5508) );
  XNOR U5719 ( .A(n5514), .B(n5512), .Z(n5729) );
  AND U5720 ( .A(n5730), .B(n5731), .Z(n5512) );
  NANDN U5721 ( .A(n5732), .B(n5733), .Z(n5731) );
  NANDN U5722 ( .A(n5734), .B(n5735), .Z(n5733) );
  NANDN U5723 ( .A(n5735), .B(n5734), .Z(n5730) );
  ANDN U5724 ( .B(B[46]), .A(n68), .Z(n5514) );
  XNOR U5725 ( .A(n5522), .B(n5736), .Z(n5515) );
  XNOR U5726 ( .A(n5521), .B(n5519), .Z(n5736) );
  AND U5727 ( .A(n5737), .B(n5738), .Z(n5519) );
  NANDN U5728 ( .A(n5739), .B(n5740), .Z(n5738) );
  OR U5729 ( .A(n5741), .B(n5742), .Z(n5740) );
  NAND U5730 ( .A(n5742), .B(n5741), .Z(n5737) );
  ANDN U5731 ( .B(B[47]), .A(n69), .Z(n5521) );
  XNOR U5732 ( .A(n5529), .B(n5743), .Z(n5522) );
  XNOR U5733 ( .A(n5528), .B(n5526), .Z(n5743) );
  AND U5734 ( .A(n5744), .B(n5745), .Z(n5526) );
  NANDN U5735 ( .A(n5746), .B(n5747), .Z(n5745) );
  NANDN U5736 ( .A(n5748), .B(n5749), .Z(n5747) );
  NANDN U5737 ( .A(n5749), .B(n5748), .Z(n5744) );
  ANDN U5738 ( .B(B[48]), .A(n70), .Z(n5528) );
  XNOR U5739 ( .A(n5536), .B(n5750), .Z(n5529) );
  XNOR U5740 ( .A(n5535), .B(n5533), .Z(n5750) );
  AND U5741 ( .A(n5751), .B(n5752), .Z(n5533) );
  NANDN U5742 ( .A(n5753), .B(n5754), .Z(n5752) );
  OR U5743 ( .A(n5755), .B(n5756), .Z(n5754) );
  NAND U5744 ( .A(n5756), .B(n5755), .Z(n5751) );
  ANDN U5745 ( .B(B[49]), .A(n71), .Z(n5535) );
  XNOR U5746 ( .A(n5543), .B(n5757), .Z(n5536) );
  XNOR U5747 ( .A(n5542), .B(n5540), .Z(n5757) );
  AND U5748 ( .A(n5758), .B(n5759), .Z(n5540) );
  NANDN U5749 ( .A(n5760), .B(n5761), .Z(n5759) );
  NANDN U5750 ( .A(n5762), .B(n5763), .Z(n5761) );
  NANDN U5751 ( .A(n5763), .B(n5762), .Z(n5758) );
  ANDN U5752 ( .B(B[50]), .A(n72), .Z(n5542) );
  XNOR U5753 ( .A(n5550), .B(n5764), .Z(n5543) );
  XNOR U5754 ( .A(n5549), .B(n5547), .Z(n5764) );
  AND U5755 ( .A(n5765), .B(n5766), .Z(n5547) );
  NANDN U5756 ( .A(n5767), .B(n5768), .Z(n5766) );
  OR U5757 ( .A(n5769), .B(n5770), .Z(n5768) );
  NAND U5758 ( .A(n5770), .B(n5769), .Z(n5765) );
  ANDN U5759 ( .B(B[51]), .A(n73), .Z(n5549) );
  XNOR U5760 ( .A(n5557), .B(n5771), .Z(n5550) );
  XNOR U5761 ( .A(n5556), .B(n5554), .Z(n5771) );
  AND U5762 ( .A(n5772), .B(n5773), .Z(n5554) );
  NANDN U5763 ( .A(n5774), .B(n5775), .Z(n5773) );
  NANDN U5764 ( .A(n5776), .B(n5777), .Z(n5775) );
  NANDN U5765 ( .A(n5777), .B(n5776), .Z(n5772) );
  ANDN U5766 ( .B(B[52]), .A(n74), .Z(n5556) );
  XNOR U5767 ( .A(n5564), .B(n5778), .Z(n5557) );
  XNOR U5768 ( .A(n5563), .B(n5561), .Z(n5778) );
  AND U5769 ( .A(n5779), .B(n5780), .Z(n5561) );
  NANDN U5770 ( .A(n5781), .B(n5782), .Z(n5780) );
  OR U5771 ( .A(n5783), .B(n5784), .Z(n5782) );
  NAND U5772 ( .A(n5784), .B(n5783), .Z(n5779) );
  ANDN U5773 ( .B(B[53]), .A(n75), .Z(n5563) );
  XNOR U5774 ( .A(n5571), .B(n5785), .Z(n5564) );
  XNOR U5775 ( .A(n5570), .B(n5568), .Z(n5785) );
  AND U5776 ( .A(n5786), .B(n5787), .Z(n5568) );
  NANDN U5777 ( .A(n5788), .B(n5789), .Z(n5787) );
  NANDN U5778 ( .A(n5790), .B(n5791), .Z(n5789) );
  NANDN U5779 ( .A(n5791), .B(n5790), .Z(n5786) );
  ANDN U5780 ( .B(B[54]), .A(n76), .Z(n5570) );
  XNOR U5781 ( .A(n5578), .B(n5792), .Z(n5571) );
  XNOR U5782 ( .A(n5577), .B(n5575), .Z(n5792) );
  AND U5783 ( .A(n5793), .B(n5794), .Z(n5575) );
  NANDN U5784 ( .A(n5795), .B(n5796), .Z(n5794) );
  OR U5785 ( .A(n5797), .B(n5798), .Z(n5796) );
  NAND U5786 ( .A(n5798), .B(n5797), .Z(n5793) );
  ANDN U5787 ( .B(B[55]), .A(n77), .Z(n5577) );
  XNOR U5788 ( .A(n5585), .B(n5799), .Z(n5578) );
  XNOR U5789 ( .A(n5584), .B(n5582), .Z(n5799) );
  AND U5790 ( .A(n5800), .B(n5801), .Z(n5582) );
  NANDN U5791 ( .A(n5802), .B(n5803), .Z(n5801) );
  NANDN U5792 ( .A(n5804), .B(n5805), .Z(n5803) );
  NANDN U5793 ( .A(n5805), .B(n5804), .Z(n5800) );
  ANDN U5794 ( .B(B[56]), .A(n78), .Z(n5584) );
  XNOR U5795 ( .A(n5592), .B(n5806), .Z(n5585) );
  XNOR U5796 ( .A(n5591), .B(n5589), .Z(n5806) );
  AND U5797 ( .A(n5807), .B(n5808), .Z(n5589) );
  NANDN U5798 ( .A(n5809), .B(n5810), .Z(n5808) );
  OR U5799 ( .A(n5811), .B(n5812), .Z(n5810) );
  NAND U5800 ( .A(n5812), .B(n5811), .Z(n5807) );
  ANDN U5801 ( .B(B[57]), .A(n79), .Z(n5591) );
  XNOR U5802 ( .A(n5599), .B(n5813), .Z(n5592) );
  XNOR U5803 ( .A(n5598), .B(n5596), .Z(n5813) );
  AND U5804 ( .A(n5814), .B(n5815), .Z(n5596) );
  NANDN U5805 ( .A(n5816), .B(n5817), .Z(n5815) );
  NANDN U5806 ( .A(n5818), .B(n5819), .Z(n5817) );
  NANDN U5807 ( .A(n5819), .B(n5818), .Z(n5814) );
  ANDN U5808 ( .B(B[58]), .A(n80), .Z(n5598) );
  XNOR U5809 ( .A(n5606), .B(n5820), .Z(n5599) );
  XNOR U5810 ( .A(n5605), .B(n5603), .Z(n5820) );
  AND U5811 ( .A(n5821), .B(n5822), .Z(n5603) );
  NANDN U5812 ( .A(n5823), .B(n5824), .Z(n5822) );
  OR U5813 ( .A(n5825), .B(n5826), .Z(n5824) );
  NAND U5814 ( .A(n5826), .B(n5825), .Z(n5821) );
  ANDN U5815 ( .B(B[59]), .A(n81), .Z(n5605) );
  XNOR U5816 ( .A(n5613), .B(n5827), .Z(n5606) );
  XNOR U5817 ( .A(n5612), .B(n5610), .Z(n5827) );
  AND U5818 ( .A(n5828), .B(n5829), .Z(n5610) );
  NANDN U5819 ( .A(n5830), .B(n5831), .Z(n5829) );
  NAND U5820 ( .A(n5832), .B(n5833), .Z(n5831) );
  ANDN U5821 ( .B(B[60]), .A(n82), .Z(n5612) );
  XOR U5822 ( .A(n5619), .B(n5834), .Z(n5613) );
  XNOR U5823 ( .A(n5617), .B(n5620), .Z(n5834) );
  NAND U5824 ( .A(A[2]), .B(B[61]), .Z(n5620) );
  NANDN U5825 ( .A(n5835), .B(n5836), .Z(n5617) );
  AND U5826 ( .A(A[0]), .B(B[62]), .Z(n5836) );
  XNOR U5827 ( .A(n5622), .B(n5837), .Z(n5619) );
  NAND U5828 ( .A(A[0]), .B(B[63]), .Z(n5837) );
  NAND U5829 ( .A(B[62]), .B(A[1]), .Z(n5622) );
  NAND U5830 ( .A(n5838), .B(n5839), .Z(n161) );
  NANDN U5831 ( .A(n5840), .B(n5841), .Z(n5839) );
  OR U5832 ( .A(n5842), .B(n5843), .Z(n5841) );
  NAND U5833 ( .A(n5843), .B(n5842), .Z(n5838) );
  XOR U5834 ( .A(n163), .B(n162), .Z(\A1[60] ) );
  XOR U5835 ( .A(n5843), .B(n5844), .Z(n162) );
  XNOR U5836 ( .A(n5842), .B(n5840), .Z(n5844) );
  AND U5837 ( .A(n5845), .B(n5846), .Z(n5840) );
  NANDN U5838 ( .A(n5847), .B(n5848), .Z(n5846) );
  NANDN U5839 ( .A(n5849), .B(n5850), .Z(n5848) );
  NANDN U5840 ( .A(n5850), .B(n5849), .Z(n5845) );
  ANDN U5841 ( .B(B[31]), .A(n54), .Z(n5842) );
  XNOR U5842 ( .A(n5637), .B(n5851), .Z(n5843) );
  XNOR U5843 ( .A(n5636), .B(n5634), .Z(n5851) );
  AND U5844 ( .A(n5852), .B(n5853), .Z(n5634) );
  NANDN U5845 ( .A(n5854), .B(n5855), .Z(n5853) );
  OR U5846 ( .A(n5856), .B(n5857), .Z(n5855) );
  NAND U5847 ( .A(n5857), .B(n5856), .Z(n5852) );
  ANDN U5848 ( .B(B[32]), .A(n55), .Z(n5636) );
  XNOR U5849 ( .A(n5644), .B(n5858), .Z(n5637) );
  XNOR U5850 ( .A(n5643), .B(n5641), .Z(n5858) );
  AND U5851 ( .A(n5859), .B(n5860), .Z(n5641) );
  NANDN U5852 ( .A(n5861), .B(n5862), .Z(n5860) );
  NANDN U5853 ( .A(n5863), .B(n5864), .Z(n5862) );
  NANDN U5854 ( .A(n5864), .B(n5863), .Z(n5859) );
  ANDN U5855 ( .B(B[33]), .A(n56), .Z(n5643) );
  XNOR U5856 ( .A(n5651), .B(n5865), .Z(n5644) );
  XNOR U5857 ( .A(n5650), .B(n5648), .Z(n5865) );
  AND U5858 ( .A(n5866), .B(n5867), .Z(n5648) );
  NANDN U5859 ( .A(n5868), .B(n5869), .Z(n5867) );
  OR U5860 ( .A(n5870), .B(n5871), .Z(n5869) );
  NAND U5861 ( .A(n5871), .B(n5870), .Z(n5866) );
  ANDN U5862 ( .B(B[34]), .A(n57), .Z(n5650) );
  XNOR U5863 ( .A(n5658), .B(n5872), .Z(n5651) );
  XNOR U5864 ( .A(n5657), .B(n5655), .Z(n5872) );
  AND U5865 ( .A(n5873), .B(n5874), .Z(n5655) );
  NANDN U5866 ( .A(n5875), .B(n5876), .Z(n5874) );
  NANDN U5867 ( .A(n5877), .B(n5878), .Z(n5876) );
  NANDN U5868 ( .A(n5878), .B(n5877), .Z(n5873) );
  ANDN U5869 ( .B(B[35]), .A(n58), .Z(n5657) );
  XNOR U5870 ( .A(n5665), .B(n5879), .Z(n5658) );
  XNOR U5871 ( .A(n5664), .B(n5662), .Z(n5879) );
  AND U5872 ( .A(n5880), .B(n5881), .Z(n5662) );
  NANDN U5873 ( .A(n5882), .B(n5883), .Z(n5881) );
  OR U5874 ( .A(n5884), .B(n5885), .Z(n5883) );
  NAND U5875 ( .A(n5885), .B(n5884), .Z(n5880) );
  ANDN U5876 ( .B(B[36]), .A(n59), .Z(n5664) );
  XNOR U5877 ( .A(n5672), .B(n5886), .Z(n5665) );
  XNOR U5878 ( .A(n5671), .B(n5669), .Z(n5886) );
  AND U5879 ( .A(n5887), .B(n5888), .Z(n5669) );
  NANDN U5880 ( .A(n5889), .B(n5890), .Z(n5888) );
  NANDN U5881 ( .A(n5891), .B(n5892), .Z(n5890) );
  NANDN U5882 ( .A(n5892), .B(n5891), .Z(n5887) );
  ANDN U5883 ( .B(B[37]), .A(n60), .Z(n5671) );
  XNOR U5884 ( .A(n5679), .B(n5893), .Z(n5672) );
  XNOR U5885 ( .A(n5678), .B(n5676), .Z(n5893) );
  AND U5886 ( .A(n5894), .B(n5895), .Z(n5676) );
  NANDN U5887 ( .A(n5896), .B(n5897), .Z(n5895) );
  OR U5888 ( .A(n5898), .B(n5899), .Z(n5897) );
  NAND U5889 ( .A(n5899), .B(n5898), .Z(n5894) );
  ANDN U5890 ( .B(B[38]), .A(n61), .Z(n5678) );
  XNOR U5891 ( .A(n5686), .B(n5900), .Z(n5679) );
  XNOR U5892 ( .A(n5685), .B(n5683), .Z(n5900) );
  AND U5893 ( .A(n5901), .B(n5902), .Z(n5683) );
  NANDN U5894 ( .A(n5903), .B(n5904), .Z(n5902) );
  NANDN U5895 ( .A(n5905), .B(n5906), .Z(n5904) );
  NANDN U5896 ( .A(n5906), .B(n5905), .Z(n5901) );
  ANDN U5897 ( .B(B[39]), .A(n62), .Z(n5685) );
  XNOR U5898 ( .A(n5693), .B(n5907), .Z(n5686) );
  XNOR U5899 ( .A(n5692), .B(n5690), .Z(n5907) );
  AND U5900 ( .A(n5908), .B(n5909), .Z(n5690) );
  NANDN U5901 ( .A(n5910), .B(n5911), .Z(n5909) );
  OR U5902 ( .A(n5912), .B(n5913), .Z(n5911) );
  NAND U5903 ( .A(n5913), .B(n5912), .Z(n5908) );
  ANDN U5904 ( .B(B[40]), .A(n63), .Z(n5692) );
  XNOR U5905 ( .A(n5700), .B(n5914), .Z(n5693) );
  XNOR U5906 ( .A(n5699), .B(n5697), .Z(n5914) );
  AND U5907 ( .A(n5915), .B(n5916), .Z(n5697) );
  NANDN U5908 ( .A(n5917), .B(n5918), .Z(n5916) );
  NANDN U5909 ( .A(n5919), .B(n5920), .Z(n5918) );
  NANDN U5910 ( .A(n5920), .B(n5919), .Z(n5915) );
  ANDN U5911 ( .B(B[41]), .A(n64), .Z(n5699) );
  XNOR U5912 ( .A(n5707), .B(n5921), .Z(n5700) );
  XNOR U5913 ( .A(n5706), .B(n5704), .Z(n5921) );
  AND U5914 ( .A(n5922), .B(n5923), .Z(n5704) );
  NANDN U5915 ( .A(n5924), .B(n5925), .Z(n5923) );
  OR U5916 ( .A(n5926), .B(n5927), .Z(n5925) );
  NAND U5917 ( .A(n5927), .B(n5926), .Z(n5922) );
  ANDN U5918 ( .B(B[42]), .A(n65), .Z(n5706) );
  XNOR U5919 ( .A(n5714), .B(n5928), .Z(n5707) );
  XNOR U5920 ( .A(n5713), .B(n5711), .Z(n5928) );
  AND U5921 ( .A(n5929), .B(n5930), .Z(n5711) );
  NANDN U5922 ( .A(n5931), .B(n5932), .Z(n5930) );
  NANDN U5923 ( .A(n5933), .B(n5934), .Z(n5932) );
  NANDN U5924 ( .A(n5934), .B(n5933), .Z(n5929) );
  ANDN U5925 ( .B(B[43]), .A(n66), .Z(n5713) );
  XNOR U5926 ( .A(n5721), .B(n5935), .Z(n5714) );
  XNOR U5927 ( .A(n5720), .B(n5718), .Z(n5935) );
  AND U5928 ( .A(n5936), .B(n5937), .Z(n5718) );
  NANDN U5929 ( .A(n5938), .B(n5939), .Z(n5937) );
  OR U5930 ( .A(n5940), .B(n5941), .Z(n5939) );
  NAND U5931 ( .A(n5941), .B(n5940), .Z(n5936) );
  ANDN U5932 ( .B(B[44]), .A(n67), .Z(n5720) );
  XNOR U5933 ( .A(n5728), .B(n5942), .Z(n5721) );
  XNOR U5934 ( .A(n5727), .B(n5725), .Z(n5942) );
  AND U5935 ( .A(n5943), .B(n5944), .Z(n5725) );
  NANDN U5936 ( .A(n5945), .B(n5946), .Z(n5944) );
  NANDN U5937 ( .A(n5947), .B(n5948), .Z(n5946) );
  NANDN U5938 ( .A(n5948), .B(n5947), .Z(n5943) );
  ANDN U5939 ( .B(B[45]), .A(n68), .Z(n5727) );
  XNOR U5940 ( .A(n5735), .B(n5949), .Z(n5728) );
  XNOR U5941 ( .A(n5734), .B(n5732), .Z(n5949) );
  AND U5942 ( .A(n5950), .B(n5951), .Z(n5732) );
  NANDN U5943 ( .A(n5952), .B(n5953), .Z(n5951) );
  OR U5944 ( .A(n5954), .B(n5955), .Z(n5953) );
  NAND U5945 ( .A(n5955), .B(n5954), .Z(n5950) );
  ANDN U5946 ( .B(B[46]), .A(n69), .Z(n5734) );
  XNOR U5947 ( .A(n5742), .B(n5956), .Z(n5735) );
  XNOR U5948 ( .A(n5741), .B(n5739), .Z(n5956) );
  AND U5949 ( .A(n5957), .B(n5958), .Z(n5739) );
  NANDN U5950 ( .A(n5959), .B(n5960), .Z(n5958) );
  NANDN U5951 ( .A(n5961), .B(n5962), .Z(n5960) );
  NANDN U5952 ( .A(n5962), .B(n5961), .Z(n5957) );
  ANDN U5953 ( .B(B[47]), .A(n70), .Z(n5741) );
  XNOR U5954 ( .A(n5749), .B(n5963), .Z(n5742) );
  XNOR U5955 ( .A(n5748), .B(n5746), .Z(n5963) );
  AND U5956 ( .A(n5964), .B(n5965), .Z(n5746) );
  NANDN U5957 ( .A(n5966), .B(n5967), .Z(n5965) );
  OR U5958 ( .A(n5968), .B(n5969), .Z(n5967) );
  NAND U5959 ( .A(n5969), .B(n5968), .Z(n5964) );
  ANDN U5960 ( .B(B[48]), .A(n71), .Z(n5748) );
  XNOR U5961 ( .A(n5756), .B(n5970), .Z(n5749) );
  XNOR U5962 ( .A(n5755), .B(n5753), .Z(n5970) );
  AND U5963 ( .A(n5971), .B(n5972), .Z(n5753) );
  NANDN U5964 ( .A(n5973), .B(n5974), .Z(n5972) );
  NANDN U5965 ( .A(n5975), .B(n5976), .Z(n5974) );
  NANDN U5966 ( .A(n5976), .B(n5975), .Z(n5971) );
  ANDN U5967 ( .B(B[49]), .A(n72), .Z(n5755) );
  XNOR U5968 ( .A(n5763), .B(n5977), .Z(n5756) );
  XNOR U5969 ( .A(n5762), .B(n5760), .Z(n5977) );
  AND U5970 ( .A(n5978), .B(n5979), .Z(n5760) );
  NANDN U5971 ( .A(n5980), .B(n5981), .Z(n5979) );
  OR U5972 ( .A(n5982), .B(n5983), .Z(n5981) );
  NAND U5973 ( .A(n5983), .B(n5982), .Z(n5978) );
  ANDN U5974 ( .B(B[50]), .A(n73), .Z(n5762) );
  XNOR U5975 ( .A(n5770), .B(n5984), .Z(n5763) );
  XNOR U5976 ( .A(n5769), .B(n5767), .Z(n5984) );
  AND U5977 ( .A(n5985), .B(n5986), .Z(n5767) );
  NANDN U5978 ( .A(n5987), .B(n5988), .Z(n5986) );
  NANDN U5979 ( .A(n5989), .B(n5990), .Z(n5988) );
  NANDN U5980 ( .A(n5990), .B(n5989), .Z(n5985) );
  ANDN U5981 ( .B(B[51]), .A(n74), .Z(n5769) );
  XNOR U5982 ( .A(n5777), .B(n5991), .Z(n5770) );
  XNOR U5983 ( .A(n5776), .B(n5774), .Z(n5991) );
  AND U5984 ( .A(n5992), .B(n5993), .Z(n5774) );
  NANDN U5985 ( .A(n5994), .B(n5995), .Z(n5993) );
  OR U5986 ( .A(n5996), .B(n5997), .Z(n5995) );
  NAND U5987 ( .A(n5997), .B(n5996), .Z(n5992) );
  ANDN U5988 ( .B(B[52]), .A(n75), .Z(n5776) );
  XNOR U5989 ( .A(n5784), .B(n5998), .Z(n5777) );
  XNOR U5990 ( .A(n5783), .B(n5781), .Z(n5998) );
  AND U5991 ( .A(n5999), .B(n6000), .Z(n5781) );
  NANDN U5992 ( .A(n6001), .B(n6002), .Z(n6000) );
  NANDN U5993 ( .A(n6003), .B(n6004), .Z(n6002) );
  NANDN U5994 ( .A(n6004), .B(n6003), .Z(n5999) );
  ANDN U5995 ( .B(B[53]), .A(n76), .Z(n5783) );
  XNOR U5996 ( .A(n5791), .B(n6005), .Z(n5784) );
  XNOR U5997 ( .A(n5790), .B(n5788), .Z(n6005) );
  AND U5998 ( .A(n6006), .B(n6007), .Z(n5788) );
  NANDN U5999 ( .A(n6008), .B(n6009), .Z(n6007) );
  OR U6000 ( .A(n6010), .B(n6011), .Z(n6009) );
  NAND U6001 ( .A(n6011), .B(n6010), .Z(n6006) );
  ANDN U6002 ( .B(B[54]), .A(n77), .Z(n5790) );
  XNOR U6003 ( .A(n5798), .B(n6012), .Z(n5791) );
  XNOR U6004 ( .A(n5797), .B(n5795), .Z(n6012) );
  AND U6005 ( .A(n6013), .B(n6014), .Z(n5795) );
  NANDN U6006 ( .A(n6015), .B(n6016), .Z(n6014) );
  NANDN U6007 ( .A(n6017), .B(n6018), .Z(n6016) );
  NANDN U6008 ( .A(n6018), .B(n6017), .Z(n6013) );
  ANDN U6009 ( .B(B[55]), .A(n78), .Z(n5797) );
  XNOR U6010 ( .A(n5805), .B(n6019), .Z(n5798) );
  XNOR U6011 ( .A(n5804), .B(n5802), .Z(n6019) );
  AND U6012 ( .A(n6020), .B(n6021), .Z(n5802) );
  NANDN U6013 ( .A(n6022), .B(n6023), .Z(n6021) );
  OR U6014 ( .A(n6024), .B(n6025), .Z(n6023) );
  NAND U6015 ( .A(n6025), .B(n6024), .Z(n6020) );
  ANDN U6016 ( .B(B[56]), .A(n79), .Z(n5804) );
  XNOR U6017 ( .A(n5812), .B(n6026), .Z(n5805) );
  XNOR U6018 ( .A(n5811), .B(n5809), .Z(n6026) );
  AND U6019 ( .A(n6027), .B(n6028), .Z(n5809) );
  NANDN U6020 ( .A(n6029), .B(n6030), .Z(n6028) );
  NANDN U6021 ( .A(n6031), .B(n6032), .Z(n6030) );
  NANDN U6022 ( .A(n6032), .B(n6031), .Z(n6027) );
  ANDN U6023 ( .B(B[57]), .A(n80), .Z(n5811) );
  XNOR U6024 ( .A(n5819), .B(n6033), .Z(n5812) );
  XNOR U6025 ( .A(n5818), .B(n5816), .Z(n6033) );
  AND U6026 ( .A(n6034), .B(n6035), .Z(n5816) );
  NANDN U6027 ( .A(n6036), .B(n6037), .Z(n6035) );
  OR U6028 ( .A(n6038), .B(n6039), .Z(n6037) );
  NAND U6029 ( .A(n6039), .B(n6038), .Z(n6034) );
  ANDN U6030 ( .B(B[58]), .A(n81), .Z(n5818) );
  XNOR U6031 ( .A(n5826), .B(n6040), .Z(n5819) );
  XNOR U6032 ( .A(n5825), .B(n5823), .Z(n6040) );
  AND U6033 ( .A(n6041), .B(n6042), .Z(n5823) );
  NANDN U6034 ( .A(n6043), .B(n6044), .Z(n6042) );
  NAND U6035 ( .A(n6045), .B(n6046), .Z(n6044) );
  ANDN U6036 ( .B(B[59]), .A(n82), .Z(n5825) );
  XOR U6037 ( .A(n5832), .B(n6047), .Z(n5826) );
  XNOR U6038 ( .A(n5830), .B(n5833), .Z(n6047) );
  NAND U6039 ( .A(A[2]), .B(B[60]), .Z(n5833) );
  NANDN U6040 ( .A(n6048), .B(n6049), .Z(n5830) );
  AND U6041 ( .A(A[0]), .B(B[61]), .Z(n6049) );
  XNOR U6042 ( .A(n5835), .B(n6050), .Z(n5832) );
  NAND U6043 ( .A(A[0]), .B(B[62]), .Z(n6050) );
  NAND U6044 ( .A(B[61]), .B(A[1]), .Z(n5835) );
  NAND U6045 ( .A(n6051), .B(n6052), .Z(n163) );
  NANDN U6046 ( .A(n6053), .B(n6054), .Z(n6052) );
  OR U6047 ( .A(n6055), .B(n6056), .Z(n6054) );
  NAND U6048 ( .A(n6056), .B(n6055), .Z(n6051) );
  XOR U6049 ( .A(n6057), .B(n6058), .Z(\A1[5] ) );
  XNOR U6050 ( .A(n6059), .B(n51), .Z(n6058) );
  XOR U6051 ( .A(n165), .B(n164), .Z(\A1[59] ) );
  XOR U6052 ( .A(n6056), .B(n6060), .Z(n164) );
  XNOR U6053 ( .A(n6055), .B(n6053), .Z(n6060) );
  AND U6054 ( .A(n6061), .B(n6062), .Z(n6053) );
  NANDN U6055 ( .A(n6063), .B(n6064), .Z(n6062) );
  NANDN U6056 ( .A(n6065), .B(n6066), .Z(n6064) );
  NANDN U6057 ( .A(n6066), .B(n6065), .Z(n6061) );
  ANDN U6058 ( .B(B[30]), .A(n54), .Z(n6055) );
  XNOR U6059 ( .A(n5850), .B(n6067), .Z(n6056) );
  XNOR U6060 ( .A(n5849), .B(n5847), .Z(n6067) );
  AND U6061 ( .A(n6068), .B(n6069), .Z(n5847) );
  NANDN U6062 ( .A(n6070), .B(n6071), .Z(n6069) );
  OR U6063 ( .A(n6072), .B(n6073), .Z(n6071) );
  NAND U6064 ( .A(n6073), .B(n6072), .Z(n6068) );
  ANDN U6065 ( .B(B[31]), .A(n55), .Z(n5849) );
  XNOR U6066 ( .A(n5857), .B(n6074), .Z(n5850) );
  XNOR U6067 ( .A(n5856), .B(n5854), .Z(n6074) );
  AND U6068 ( .A(n6075), .B(n6076), .Z(n5854) );
  NANDN U6069 ( .A(n6077), .B(n6078), .Z(n6076) );
  NANDN U6070 ( .A(n6079), .B(n6080), .Z(n6078) );
  NANDN U6071 ( .A(n6080), .B(n6079), .Z(n6075) );
  ANDN U6072 ( .B(B[32]), .A(n56), .Z(n5856) );
  XNOR U6073 ( .A(n5864), .B(n6081), .Z(n5857) );
  XNOR U6074 ( .A(n5863), .B(n5861), .Z(n6081) );
  AND U6075 ( .A(n6082), .B(n6083), .Z(n5861) );
  NANDN U6076 ( .A(n6084), .B(n6085), .Z(n6083) );
  OR U6077 ( .A(n6086), .B(n6087), .Z(n6085) );
  NAND U6078 ( .A(n6087), .B(n6086), .Z(n6082) );
  ANDN U6079 ( .B(B[33]), .A(n57), .Z(n5863) );
  XNOR U6080 ( .A(n5871), .B(n6088), .Z(n5864) );
  XNOR U6081 ( .A(n5870), .B(n5868), .Z(n6088) );
  AND U6082 ( .A(n6089), .B(n6090), .Z(n5868) );
  NANDN U6083 ( .A(n6091), .B(n6092), .Z(n6090) );
  NANDN U6084 ( .A(n6093), .B(n6094), .Z(n6092) );
  NANDN U6085 ( .A(n6094), .B(n6093), .Z(n6089) );
  ANDN U6086 ( .B(B[34]), .A(n58), .Z(n5870) );
  XNOR U6087 ( .A(n5878), .B(n6095), .Z(n5871) );
  XNOR U6088 ( .A(n5877), .B(n5875), .Z(n6095) );
  AND U6089 ( .A(n6096), .B(n6097), .Z(n5875) );
  NANDN U6090 ( .A(n6098), .B(n6099), .Z(n6097) );
  OR U6091 ( .A(n6100), .B(n6101), .Z(n6099) );
  NAND U6092 ( .A(n6101), .B(n6100), .Z(n6096) );
  ANDN U6093 ( .B(B[35]), .A(n59), .Z(n5877) );
  XNOR U6094 ( .A(n5885), .B(n6102), .Z(n5878) );
  XNOR U6095 ( .A(n5884), .B(n5882), .Z(n6102) );
  AND U6096 ( .A(n6103), .B(n6104), .Z(n5882) );
  NANDN U6097 ( .A(n6105), .B(n6106), .Z(n6104) );
  NANDN U6098 ( .A(n6107), .B(n6108), .Z(n6106) );
  NANDN U6099 ( .A(n6108), .B(n6107), .Z(n6103) );
  ANDN U6100 ( .B(B[36]), .A(n60), .Z(n5884) );
  XNOR U6101 ( .A(n5892), .B(n6109), .Z(n5885) );
  XNOR U6102 ( .A(n5891), .B(n5889), .Z(n6109) );
  AND U6103 ( .A(n6110), .B(n6111), .Z(n5889) );
  NANDN U6104 ( .A(n6112), .B(n6113), .Z(n6111) );
  OR U6105 ( .A(n6114), .B(n6115), .Z(n6113) );
  NAND U6106 ( .A(n6115), .B(n6114), .Z(n6110) );
  ANDN U6107 ( .B(B[37]), .A(n61), .Z(n5891) );
  XNOR U6108 ( .A(n5899), .B(n6116), .Z(n5892) );
  XNOR U6109 ( .A(n5898), .B(n5896), .Z(n6116) );
  AND U6110 ( .A(n6117), .B(n6118), .Z(n5896) );
  NANDN U6111 ( .A(n6119), .B(n6120), .Z(n6118) );
  NANDN U6112 ( .A(n6121), .B(n6122), .Z(n6120) );
  NANDN U6113 ( .A(n6122), .B(n6121), .Z(n6117) );
  ANDN U6114 ( .B(B[38]), .A(n62), .Z(n5898) );
  XNOR U6115 ( .A(n5906), .B(n6123), .Z(n5899) );
  XNOR U6116 ( .A(n5905), .B(n5903), .Z(n6123) );
  AND U6117 ( .A(n6124), .B(n6125), .Z(n5903) );
  NANDN U6118 ( .A(n6126), .B(n6127), .Z(n6125) );
  OR U6119 ( .A(n6128), .B(n6129), .Z(n6127) );
  NAND U6120 ( .A(n6129), .B(n6128), .Z(n6124) );
  ANDN U6121 ( .B(B[39]), .A(n63), .Z(n5905) );
  XNOR U6122 ( .A(n5913), .B(n6130), .Z(n5906) );
  XNOR U6123 ( .A(n5912), .B(n5910), .Z(n6130) );
  AND U6124 ( .A(n6131), .B(n6132), .Z(n5910) );
  NANDN U6125 ( .A(n6133), .B(n6134), .Z(n6132) );
  NANDN U6126 ( .A(n6135), .B(n6136), .Z(n6134) );
  NANDN U6127 ( .A(n6136), .B(n6135), .Z(n6131) );
  ANDN U6128 ( .B(B[40]), .A(n64), .Z(n5912) );
  XNOR U6129 ( .A(n5920), .B(n6137), .Z(n5913) );
  XNOR U6130 ( .A(n5919), .B(n5917), .Z(n6137) );
  AND U6131 ( .A(n6138), .B(n6139), .Z(n5917) );
  NANDN U6132 ( .A(n6140), .B(n6141), .Z(n6139) );
  OR U6133 ( .A(n6142), .B(n6143), .Z(n6141) );
  NAND U6134 ( .A(n6143), .B(n6142), .Z(n6138) );
  ANDN U6135 ( .B(B[41]), .A(n65), .Z(n5919) );
  XNOR U6136 ( .A(n5927), .B(n6144), .Z(n5920) );
  XNOR U6137 ( .A(n5926), .B(n5924), .Z(n6144) );
  AND U6138 ( .A(n6145), .B(n6146), .Z(n5924) );
  NANDN U6139 ( .A(n6147), .B(n6148), .Z(n6146) );
  NANDN U6140 ( .A(n6149), .B(n6150), .Z(n6148) );
  NANDN U6141 ( .A(n6150), .B(n6149), .Z(n6145) );
  ANDN U6142 ( .B(B[42]), .A(n66), .Z(n5926) );
  XNOR U6143 ( .A(n5934), .B(n6151), .Z(n5927) );
  XNOR U6144 ( .A(n5933), .B(n5931), .Z(n6151) );
  AND U6145 ( .A(n6152), .B(n6153), .Z(n5931) );
  NANDN U6146 ( .A(n6154), .B(n6155), .Z(n6153) );
  OR U6147 ( .A(n6156), .B(n6157), .Z(n6155) );
  NAND U6148 ( .A(n6157), .B(n6156), .Z(n6152) );
  ANDN U6149 ( .B(B[43]), .A(n67), .Z(n5933) );
  XNOR U6150 ( .A(n5941), .B(n6158), .Z(n5934) );
  XNOR U6151 ( .A(n5940), .B(n5938), .Z(n6158) );
  AND U6152 ( .A(n6159), .B(n6160), .Z(n5938) );
  NANDN U6153 ( .A(n6161), .B(n6162), .Z(n6160) );
  NANDN U6154 ( .A(n6163), .B(n6164), .Z(n6162) );
  NANDN U6155 ( .A(n6164), .B(n6163), .Z(n6159) );
  ANDN U6156 ( .B(B[44]), .A(n68), .Z(n5940) );
  XNOR U6157 ( .A(n5948), .B(n6165), .Z(n5941) );
  XNOR U6158 ( .A(n5947), .B(n5945), .Z(n6165) );
  AND U6159 ( .A(n6166), .B(n6167), .Z(n5945) );
  NANDN U6160 ( .A(n6168), .B(n6169), .Z(n6167) );
  OR U6161 ( .A(n6170), .B(n6171), .Z(n6169) );
  NAND U6162 ( .A(n6171), .B(n6170), .Z(n6166) );
  ANDN U6163 ( .B(B[45]), .A(n69), .Z(n5947) );
  XNOR U6164 ( .A(n5955), .B(n6172), .Z(n5948) );
  XNOR U6165 ( .A(n5954), .B(n5952), .Z(n6172) );
  AND U6166 ( .A(n6173), .B(n6174), .Z(n5952) );
  NANDN U6167 ( .A(n6175), .B(n6176), .Z(n6174) );
  NANDN U6168 ( .A(n6177), .B(n6178), .Z(n6176) );
  NANDN U6169 ( .A(n6178), .B(n6177), .Z(n6173) );
  ANDN U6170 ( .B(B[46]), .A(n70), .Z(n5954) );
  XNOR U6171 ( .A(n5962), .B(n6179), .Z(n5955) );
  XNOR U6172 ( .A(n5961), .B(n5959), .Z(n6179) );
  AND U6173 ( .A(n6180), .B(n6181), .Z(n5959) );
  NANDN U6174 ( .A(n6182), .B(n6183), .Z(n6181) );
  OR U6175 ( .A(n6184), .B(n6185), .Z(n6183) );
  NAND U6176 ( .A(n6185), .B(n6184), .Z(n6180) );
  ANDN U6177 ( .B(B[47]), .A(n71), .Z(n5961) );
  XNOR U6178 ( .A(n5969), .B(n6186), .Z(n5962) );
  XNOR U6179 ( .A(n5968), .B(n5966), .Z(n6186) );
  AND U6180 ( .A(n6187), .B(n6188), .Z(n5966) );
  NANDN U6181 ( .A(n6189), .B(n6190), .Z(n6188) );
  NANDN U6182 ( .A(n6191), .B(n6192), .Z(n6190) );
  NANDN U6183 ( .A(n6192), .B(n6191), .Z(n6187) );
  ANDN U6184 ( .B(B[48]), .A(n72), .Z(n5968) );
  XNOR U6185 ( .A(n5976), .B(n6193), .Z(n5969) );
  XNOR U6186 ( .A(n5975), .B(n5973), .Z(n6193) );
  AND U6187 ( .A(n6194), .B(n6195), .Z(n5973) );
  NANDN U6188 ( .A(n6196), .B(n6197), .Z(n6195) );
  OR U6189 ( .A(n6198), .B(n6199), .Z(n6197) );
  NAND U6190 ( .A(n6199), .B(n6198), .Z(n6194) );
  ANDN U6191 ( .B(B[49]), .A(n73), .Z(n5975) );
  XNOR U6192 ( .A(n5983), .B(n6200), .Z(n5976) );
  XNOR U6193 ( .A(n5982), .B(n5980), .Z(n6200) );
  AND U6194 ( .A(n6201), .B(n6202), .Z(n5980) );
  NANDN U6195 ( .A(n6203), .B(n6204), .Z(n6202) );
  NANDN U6196 ( .A(n6205), .B(n6206), .Z(n6204) );
  NANDN U6197 ( .A(n6206), .B(n6205), .Z(n6201) );
  ANDN U6198 ( .B(B[50]), .A(n74), .Z(n5982) );
  XNOR U6199 ( .A(n5990), .B(n6207), .Z(n5983) );
  XNOR U6200 ( .A(n5989), .B(n5987), .Z(n6207) );
  AND U6201 ( .A(n6208), .B(n6209), .Z(n5987) );
  NANDN U6202 ( .A(n6210), .B(n6211), .Z(n6209) );
  OR U6203 ( .A(n6212), .B(n6213), .Z(n6211) );
  NAND U6204 ( .A(n6213), .B(n6212), .Z(n6208) );
  ANDN U6205 ( .B(B[51]), .A(n75), .Z(n5989) );
  XNOR U6206 ( .A(n5997), .B(n6214), .Z(n5990) );
  XNOR U6207 ( .A(n5996), .B(n5994), .Z(n6214) );
  AND U6208 ( .A(n6215), .B(n6216), .Z(n5994) );
  NANDN U6209 ( .A(n6217), .B(n6218), .Z(n6216) );
  NANDN U6210 ( .A(n6219), .B(n6220), .Z(n6218) );
  NANDN U6211 ( .A(n6220), .B(n6219), .Z(n6215) );
  ANDN U6212 ( .B(B[52]), .A(n76), .Z(n5996) );
  XNOR U6213 ( .A(n6004), .B(n6221), .Z(n5997) );
  XNOR U6214 ( .A(n6003), .B(n6001), .Z(n6221) );
  AND U6215 ( .A(n6222), .B(n6223), .Z(n6001) );
  NANDN U6216 ( .A(n6224), .B(n6225), .Z(n6223) );
  OR U6217 ( .A(n6226), .B(n6227), .Z(n6225) );
  NAND U6218 ( .A(n6227), .B(n6226), .Z(n6222) );
  ANDN U6219 ( .B(B[53]), .A(n77), .Z(n6003) );
  XNOR U6220 ( .A(n6011), .B(n6228), .Z(n6004) );
  XNOR U6221 ( .A(n6010), .B(n6008), .Z(n6228) );
  AND U6222 ( .A(n6229), .B(n6230), .Z(n6008) );
  NANDN U6223 ( .A(n6231), .B(n6232), .Z(n6230) );
  NANDN U6224 ( .A(n6233), .B(n6234), .Z(n6232) );
  NANDN U6225 ( .A(n6234), .B(n6233), .Z(n6229) );
  ANDN U6226 ( .B(B[54]), .A(n78), .Z(n6010) );
  XNOR U6227 ( .A(n6018), .B(n6235), .Z(n6011) );
  XNOR U6228 ( .A(n6017), .B(n6015), .Z(n6235) );
  AND U6229 ( .A(n6236), .B(n6237), .Z(n6015) );
  NANDN U6230 ( .A(n6238), .B(n6239), .Z(n6237) );
  OR U6231 ( .A(n6240), .B(n6241), .Z(n6239) );
  NAND U6232 ( .A(n6241), .B(n6240), .Z(n6236) );
  ANDN U6233 ( .B(B[55]), .A(n79), .Z(n6017) );
  XNOR U6234 ( .A(n6025), .B(n6242), .Z(n6018) );
  XNOR U6235 ( .A(n6024), .B(n6022), .Z(n6242) );
  AND U6236 ( .A(n6243), .B(n6244), .Z(n6022) );
  NANDN U6237 ( .A(n6245), .B(n6246), .Z(n6244) );
  NANDN U6238 ( .A(n6247), .B(n6248), .Z(n6246) );
  NANDN U6239 ( .A(n6248), .B(n6247), .Z(n6243) );
  ANDN U6240 ( .B(B[56]), .A(n80), .Z(n6024) );
  XNOR U6241 ( .A(n6032), .B(n6249), .Z(n6025) );
  XNOR U6242 ( .A(n6031), .B(n6029), .Z(n6249) );
  AND U6243 ( .A(n6250), .B(n6251), .Z(n6029) );
  NANDN U6244 ( .A(n6252), .B(n6253), .Z(n6251) );
  OR U6245 ( .A(n6254), .B(n6255), .Z(n6253) );
  NAND U6246 ( .A(n6255), .B(n6254), .Z(n6250) );
  ANDN U6247 ( .B(B[57]), .A(n81), .Z(n6031) );
  XNOR U6248 ( .A(n6039), .B(n6256), .Z(n6032) );
  XNOR U6249 ( .A(n6038), .B(n6036), .Z(n6256) );
  AND U6250 ( .A(n6257), .B(n6258), .Z(n6036) );
  NANDN U6251 ( .A(n6259), .B(n6260), .Z(n6258) );
  NAND U6252 ( .A(n6261), .B(n6262), .Z(n6260) );
  ANDN U6253 ( .B(B[58]), .A(n82), .Z(n6038) );
  XOR U6254 ( .A(n6045), .B(n6263), .Z(n6039) );
  XNOR U6255 ( .A(n6043), .B(n6046), .Z(n6263) );
  NAND U6256 ( .A(A[2]), .B(B[59]), .Z(n6046) );
  NANDN U6257 ( .A(n6264), .B(n6265), .Z(n6043) );
  AND U6258 ( .A(A[0]), .B(B[60]), .Z(n6265) );
  XNOR U6259 ( .A(n6048), .B(n6266), .Z(n6045) );
  NAND U6260 ( .A(A[0]), .B(B[61]), .Z(n6266) );
  NAND U6261 ( .A(B[60]), .B(A[1]), .Z(n6048) );
  NAND U6262 ( .A(n6267), .B(n6268), .Z(n165) );
  NANDN U6263 ( .A(n6269), .B(n6270), .Z(n6268) );
  OR U6264 ( .A(n6271), .B(n6272), .Z(n6270) );
  NAND U6265 ( .A(n6272), .B(n6271), .Z(n6267) );
  XOR U6266 ( .A(n167), .B(n166), .Z(\A1[58] ) );
  XOR U6267 ( .A(n6272), .B(n6273), .Z(n166) );
  XNOR U6268 ( .A(n6271), .B(n6269), .Z(n6273) );
  AND U6269 ( .A(n6274), .B(n6275), .Z(n6269) );
  NANDN U6270 ( .A(n6276), .B(n6277), .Z(n6275) );
  NANDN U6271 ( .A(n6278), .B(n6279), .Z(n6277) );
  NANDN U6272 ( .A(n6279), .B(n6278), .Z(n6274) );
  ANDN U6273 ( .B(B[29]), .A(n54), .Z(n6271) );
  XNOR U6274 ( .A(n6066), .B(n6280), .Z(n6272) );
  XNOR U6275 ( .A(n6065), .B(n6063), .Z(n6280) );
  AND U6276 ( .A(n6281), .B(n6282), .Z(n6063) );
  NANDN U6277 ( .A(n6283), .B(n6284), .Z(n6282) );
  OR U6278 ( .A(n6285), .B(n6286), .Z(n6284) );
  NAND U6279 ( .A(n6286), .B(n6285), .Z(n6281) );
  ANDN U6280 ( .B(B[30]), .A(n55), .Z(n6065) );
  XNOR U6281 ( .A(n6073), .B(n6287), .Z(n6066) );
  XNOR U6282 ( .A(n6072), .B(n6070), .Z(n6287) );
  AND U6283 ( .A(n6288), .B(n6289), .Z(n6070) );
  NANDN U6284 ( .A(n6290), .B(n6291), .Z(n6289) );
  NANDN U6285 ( .A(n6292), .B(n6293), .Z(n6291) );
  NANDN U6286 ( .A(n6293), .B(n6292), .Z(n6288) );
  ANDN U6287 ( .B(B[31]), .A(n56), .Z(n6072) );
  XNOR U6288 ( .A(n6080), .B(n6294), .Z(n6073) );
  XNOR U6289 ( .A(n6079), .B(n6077), .Z(n6294) );
  AND U6290 ( .A(n6295), .B(n6296), .Z(n6077) );
  NANDN U6291 ( .A(n6297), .B(n6298), .Z(n6296) );
  OR U6292 ( .A(n6299), .B(n6300), .Z(n6298) );
  NAND U6293 ( .A(n6300), .B(n6299), .Z(n6295) );
  ANDN U6294 ( .B(B[32]), .A(n57), .Z(n6079) );
  XNOR U6295 ( .A(n6087), .B(n6301), .Z(n6080) );
  XNOR U6296 ( .A(n6086), .B(n6084), .Z(n6301) );
  AND U6297 ( .A(n6302), .B(n6303), .Z(n6084) );
  NANDN U6298 ( .A(n6304), .B(n6305), .Z(n6303) );
  NANDN U6299 ( .A(n6306), .B(n6307), .Z(n6305) );
  NANDN U6300 ( .A(n6307), .B(n6306), .Z(n6302) );
  ANDN U6301 ( .B(B[33]), .A(n58), .Z(n6086) );
  XNOR U6302 ( .A(n6094), .B(n6308), .Z(n6087) );
  XNOR U6303 ( .A(n6093), .B(n6091), .Z(n6308) );
  AND U6304 ( .A(n6309), .B(n6310), .Z(n6091) );
  NANDN U6305 ( .A(n6311), .B(n6312), .Z(n6310) );
  OR U6306 ( .A(n6313), .B(n6314), .Z(n6312) );
  NAND U6307 ( .A(n6314), .B(n6313), .Z(n6309) );
  ANDN U6308 ( .B(B[34]), .A(n59), .Z(n6093) );
  XNOR U6309 ( .A(n6101), .B(n6315), .Z(n6094) );
  XNOR U6310 ( .A(n6100), .B(n6098), .Z(n6315) );
  AND U6311 ( .A(n6316), .B(n6317), .Z(n6098) );
  NANDN U6312 ( .A(n6318), .B(n6319), .Z(n6317) );
  NANDN U6313 ( .A(n6320), .B(n6321), .Z(n6319) );
  NANDN U6314 ( .A(n6321), .B(n6320), .Z(n6316) );
  ANDN U6315 ( .B(B[35]), .A(n60), .Z(n6100) );
  XNOR U6316 ( .A(n6108), .B(n6322), .Z(n6101) );
  XNOR U6317 ( .A(n6107), .B(n6105), .Z(n6322) );
  AND U6318 ( .A(n6323), .B(n6324), .Z(n6105) );
  NANDN U6319 ( .A(n6325), .B(n6326), .Z(n6324) );
  OR U6320 ( .A(n6327), .B(n6328), .Z(n6326) );
  NAND U6321 ( .A(n6328), .B(n6327), .Z(n6323) );
  ANDN U6322 ( .B(B[36]), .A(n61), .Z(n6107) );
  XNOR U6323 ( .A(n6115), .B(n6329), .Z(n6108) );
  XNOR U6324 ( .A(n6114), .B(n6112), .Z(n6329) );
  AND U6325 ( .A(n6330), .B(n6331), .Z(n6112) );
  NANDN U6326 ( .A(n6332), .B(n6333), .Z(n6331) );
  NANDN U6327 ( .A(n6334), .B(n6335), .Z(n6333) );
  NANDN U6328 ( .A(n6335), .B(n6334), .Z(n6330) );
  ANDN U6329 ( .B(B[37]), .A(n62), .Z(n6114) );
  XNOR U6330 ( .A(n6122), .B(n6336), .Z(n6115) );
  XNOR U6331 ( .A(n6121), .B(n6119), .Z(n6336) );
  AND U6332 ( .A(n6337), .B(n6338), .Z(n6119) );
  NANDN U6333 ( .A(n6339), .B(n6340), .Z(n6338) );
  OR U6334 ( .A(n6341), .B(n6342), .Z(n6340) );
  NAND U6335 ( .A(n6342), .B(n6341), .Z(n6337) );
  ANDN U6336 ( .B(B[38]), .A(n63), .Z(n6121) );
  XNOR U6337 ( .A(n6129), .B(n6343), .Z(n6122) );
  XNOR U6338 ( .A(n6128), .B(n6126), .Z(n6343) );
  AND U6339 ( .A(n6344), .B(n6345), .Z(n6126) );
  NANDN U6340 ( .A(n6346), .B(n6347), .Z(n6345) );
  NANDN U6341 ( .A(n6348), .B(n6349), .Z(n6347) );
  NANDN U6342 ( .A(n6349), .B(n6348), .Z(n6344) );
  ANDN U6343 ( .B(B[39]), .A(n64), .Z(n6128) );
  XNOR U6344 ( .A(n6136), .B(n6350), .Z(n6129) );
  XNOR U6345 ( .A(n6135), .B(n6133), .Z(n6350) );
  AND U6346 ( .A(n6351), .B(n6352), .Z(n6133) );
  NANDN U6347 ( .A(n6353), .B(n6354), .Z(n6352) );
  OR U6348 ( .A(n6355), .B(n6356), .Z(n6354) );
  NAND U6349 ( .A(n6356), .B(n6355), .Z(n6351) );
  ANDN U6350 ( .B(B[40]), .A(n65), .Z(n6135) );
  XNOR U6351 ( .A(n6143), .B(n6357), .Z(n6136) );
  XNOR U6352 ( .A(n6142), .B(n6140), .Z(n6357) );
  AND U6353 ( .A(n6358), .B(n6359), .Z(n6140) );
  NANDN U6354 ( .A(n6360), .B(n6361), .Z(n6359) );
  NANDN U6355 ( .A(n6362), .B(n6363), .Z(n6361) );
  NANDN U6356 ( .A(n6363), .B(n6362), .Z(n6358) );
  ANDN U6357 ( .B(B[41]), .A(n66), .Z(n6142) );
  XNOR U6358 ( .A(n6150), .B(n6364), .Z(n6143) );
  XNOR U6359 ( .A(n6149), .B(n6147), .Z(n6364) );
  AND U6360 ( .A(n6365), .B(n6366), .Z(n6147) );
  NANDN U6361 ( .A(n6367), .B(n6368), .Z(n6366) );
  OR U6362 ( .A(n6369), .B(n6370), .Z(n6368) );
  NAND U6363 ( .A(n6370), .B(n6369), .Z(n6365) );
  ANDN U6364 ( .B(B[42]), .A(n67), .Z(n6149) );
  XNOR U6365 ( .A(n6157), .B(n6371), .Z(n6150) );
  XNOR U6366 ( .A(n6156), .B(n6154), .Z(n6371) );
  AND U6367 ( .A(n6372), .B(n6373), .Z(n6154) );
  NANDN U6368 ( .A(n6374), .B(n6375), .Z(n6373) );
  NANDN U6369 ( .A(n6376), .B(n6377), .Z(n6375) );
  NANDN U6370 ( .A(n6377), .B(n6376), .Z(n6372) );
  ANDN U6371 ( .B(B[43]), .A(n68), .Z(n6156) );
  XNOR U6372 ( .A(n6164), .B(n6378), .Z(n6157) );
  XNOR U6373 ( .A(n6163), .B(n6161), .Z(n6378) );
  AND U6374 ( .A(n6379), .B(n6380), .Z(n6161) );
  NANDN U6375 ( .A(n6381), .B(n6382), .Z(n6380) );
  OR U6376 ( .A(n6383), .B(n6384), .Z(n6382) );
  NAND U6377 ( .A(n6384), .B(n6383), .Z(n6379) );
  ANDN U6378 ( .B(B[44]), .A(n69), .Z(n6163) );
  XNOR U6379 ( .A(n6171), .B(n6385), .Z(n6164) );
  XNOR U6380 ( .A(n6170), .B(n6168), .Z(n6385) );
  AND U6381 ( .A(n6386), .B(n6387), .Z(n6168) );
  NANDN U6382 ( .A(n6388), .B(n6389), .Z(n6387) );
  NANDN U6383 ( .A(n6390), .B(n6391), .Z(n6389) );
  NANDN U6384 ( .A(n6391), .B(n6390), .Z(n6386) );
  ANDN U6385 ( .B(B[45]), .A(n70), .Z(n6170) );
  XNOR U6386 ( .A(n6178), .B(n6392), .Z(n6171) );
  XNOR U6387 ( .A(n6177), .B(n6175), .Z(n6392) );
  AND U6388 ( .A(n6393), .B(n6394), .Z(n6175) );
  NANDN U6389 ( .A(n6395), .B(n6396), .Z(n6394) );
  OR U6390 ( .A(n6397), .B(n6398), .Z(n6396) );
  NAND U6391 ( .A(n6398), .B(n6397), .Z(n6393) );
  ANDN U6392 ( .B(B[46]), .A(n71), .Z(n6177) );
  XNOR U6393 ( .A(n6185), .B(n6399), .Z(n6178) );
  XNOR U6394 ( .A(n6184), .B(n6182), .Z(n6399) );
  AND U6395 ( .A(n6400), .B(n6401), .Z(n6182) );
  NANDN U6396 ( .A(n6402), .B(n6403), .Z(n6401) );
  NANDN U6397 ( .A(n6404), .B(n6405), .Z(n6403) );
  NANDN U6398 ( .A(n6405), .B(n6404), .Z(n6400) );
  ANDN U6399 ( .B(B[47]), .A(n72), .Z(n6184) );
  XNOR U6400 ( .A(n6192), .B(n6406), .Z(n6185) );
  XNOR U6401 ( .A(n6191), .B(n6189), .Z(n6406) );
  AND U6402 ( .A(n6407), .B(n6408), .Z(n6189) );
  NANDN U6403 ( .A(n6409), .B(n6410), .Z(n6408) );
  OR U6404 ( .A(n6411), .B(n6412), .Z(n6410) );
  NAND U6405 ( .A(n6412), .B(n6411), .Z(n6407) );
  ANDN U6406 ( .B(B[48]), .A(n73), .Z(n6191) );
  XNOR U6407 ( .A(n6199), .B(n6413), .Z(n6192) );
  XNOR U6408 ( .A(n6198), .B(n6196), .Z(n6413) );
  AND U6409 ( .A(n6414), .B(n6415), .Z(n6196) );
  NANDN U6410 ( .A(n6416), .B(n6417), .Z(n6415) );
  NANDN U6411 ( .A(n6418), .B(n6419), .Z(n6417) );
  NANDN U6412 ( .A(n6419), .B(n6418), .Z(n6414) );
  ANDN U6413 ( .B(B[49]), .A(n74), .Z(n6198) );
  XNOR U6414 ( .A(n6206), .B(n6420), .Z(n6199) );
  XNOR U6415 ( .A(n6205), .B(n6203), .Z(n6420) );
  AND U6416 ( .A(n6421), .B(n6422), .Z(n6203) );
  NANDN U6417 ( .A(n6423), .B(n6424), .Z(n6422) );
  OR U6418 ( .A(n6425), .B(n6426), .Z(n6424) );
  NAND U6419 ( .A(n6426), .B(n6425), .Z(n6421) );
  ANDN U6420 ( .B(B[50]), .A(n75), .Z(n6205) );
  XNOR U6421 ( .A(n6213), .B(n6427), .Z(n6206) );
  XNOR U6422 ( .A(n6212), .B(n6210), .Z(n6427) );
  AND U6423 ( .A(n6428), .B(n6429), .Z(n6210) );
  NANDN U6424 ( .A(n6430), .B(n6431), .Z(n6429) );
  NANDN U6425 ( .A(n6432), .B(n6433), .Z(n6431) );
  NANDN U6426 ( .A(n6433), .B(n6432), .Z(n6428) );
  ANDN U6427 ( .B(B[51]), .A(n76), .Z(n6212) );
  XNOR U6428 ( .A(n6220), .B(n6434), .Z(n6213) );
  XNOR U6429 ( .A(n6219), .B(n6217), .Z(n6434) );
  AND U6430 ( .A(n6435), .B(n6436), .Z(n6217) );
  NANDN U6431 ( .A(n6437), .B(n6438), .Z(n6436) );
  OR U6432 ( .A(n6439), .B(n6440), .Z(n6438) );
  NAND U6433 ( .A(n6440), .B(n6439), .Z(n6435) );
  ANDN U6434 ( .B(B[52]), .A(n77), .Z(n6219) );
  XNOR U6435 ( .A(n6227), .B(n6441), .Z(n6220) );
  XNOR U6436 ( .A(n6226), .B(n6224), .Z(n6441) );
  AND U6437 ( .A(n6442), .B(n6443), .Z(n6224) );
  NANDN U6438 ( .A(n6444), .B(n6445), .Z(n6443) );
  NANDN U6439 ( .A(n6446), .B(n6447), .Z(n6445) );
  NANDN U6440 ( .A(n6447), .B(n6446), .Z(n6442) );
  ANDN U6441 ( .B(B[53]), .A(n78), .Z(n6226) );
  XNOR U6442 ( .A(n6234), .B(n6448), .Z(n6227) );
  XNOR U6443 ( .A(n6233), .B(n6231), .Z(n6448) );
  AND U6444 ( .A(n6449), .B(n6450), .Z(n6231) );
  NANDN U6445 ( .A(n6451), .B(n6452), .Z(n6450) );
  OR U6446 ( .A(n6453), .B(n6454), .Z(n6452) );
  NAND U6447 ( .A(n6454), .B(n6453), .Z(n6449) );
  ANDN U6448 ( .B(B[54]), .A(n79), .Z(n6233) );
  XNOR U6449 ( .A(n6241), .B(n6455), .Z(n6234) );
  XNOR U6450 ( .A(n6240), .B(n6238), .Z(n6455) );
  AND U6451 ( .A(n6456), .B(n6457), .Z(n6238) );
  NANDN U6452 ( .A(n6458), .B(n6459), .Z(n6457) );
  NANDN U6453 ( .A(n6460), .B(n6461), .Z(n6459) );
  NANDN U6454 ( .A(n6461), .B(n6460), .Z(n6456) );
  ANDN U6455 ( .B(B[55]), .A(n80), .Z(n6240) );
  XNOR U6456 ( .A(n6248), .B(n6462), .Z(n6241) );
  XNOR U6457 ( .A(n6247), .B(n6245), .Z(n6462) );
  AND U6458 ( .A(n6463), .B(n6464), .Z(n6245) );
  NANDN U6459 ( .A(n6465), .B(n6466), .Z(n6464) );
  OR U6460 ( .A(n6467), .B(n6468), .Z(n6466) );
  NAND U6461 ( .A(n6468), .B(n6467), .Z(n6463) );
  ANDN U6462 ( .B(B[56]), .A(n81), .Z(n6247) );
  XNOR U6463 ( .A(n6255), .B(n6469), .Z(n6248) );
  XNOR U6464 ( .A(n6254), .B(n6252), .Z(n6469) );
  AND U6465 ( .A(n6470), .B(n6471), .Z(n6252) );
  NANDN U6466 ( .A(n6472), .B(n6473), .Z(n6471) );
  NAND U6467 ( .A(n6474), .B(n6475), .Z(n6473) );
  ANDN U6468 ( .B(B[57]), .A(n82), .Z(n6254) );
  XOR U6469 ( .A(n6261), .B(n6476), .Z(n6255) );
  XNOR U6470 ( .A(n6259), .B(n6262), .Z(n6476) );
  NAND U6471 ( .A(A[2]), .B(B[58]), .Z(n6262) );
  NANDN U6472 ( .A(n6477), .B(n6478), .Z(n6259) );
  AND U6473 ( .A(A[0]), .B(B[59]), .Z(n6478) );
  XNOR U6474 ( .A(n6264), .B(n6479), .Z(n6261) );
  NAND U6475 ( .A(A[0]), .B(B[60]), .Z(n6479) );
  NAND U6476 ( .A(B[59]), .B(A[1]), .Z(n6264) );
  NAND U6477 ( .A(n6480), .B(n6481), .Z(n167) );
  NANDN U6478 ( .A(n6482), .B(n6483), .Z(n6481) );
  OR U6479 ( .A(n6484), .B(n6485), .Z(n6483) );
  NAND U6480 ( .A(n6485), .B(n6484), .Z(n6480) );
  XOR U6481 ( .A(n169), .B(n168), .Z(\A1[57] ) );
  XOR U6482 ( .A(n6485), .B(n6486), .Z(n168) );
  XNOR U6483 ( .A(n6484), .B(n6482), .Z(n6486) );
  AND U6484 ( .A(n6487), .B(n6488), .Z(n6482) );
  NANDN U6485 ( .A(n6489), .B(n6490), .Z(n6488) );
  NANDN U6486 ( .A(n6491), .B(n6492), .Z(n6490) );
  NANDN U6487 ( .A(n6492), .B(n6491), .Z(n6487) );
  ANDN U6488 ( .B(B[28]), .A(n54), .Z(n6484) );
  XNOR U6489 ( .A(n6279), .B(n6493), .Z(n6485) );
  XNOR U6490 ( .A(n6278), .B(n6276), .Z(n6493) );
  AND U6491 ( .A(n6494), .B(n6495), .Z(n6276) );
  NANDN U6492 ( .A(n6496), .B(n6497), .Z(n6495) );
  OR U6493 ( .A(n6498), .B(n6499), .Z(n6497) );
  NAND U6494 ( .A(n6499), .B(n6498), .Z(n6494) );
  ANDN U6495 ( .B(B[29]), .A(n55), .Z(n6278) );
  XNOR U6496 ( .A(n6286), .B(n6500), .Z(n6279) );
  XNOR U6497 ( .A(n6285), .B(n6283), .Z(n6500) );
  AND U6498 ( .A(n6501), .B(n6502), .Z(n6283) );
  NANDN U6499 ( .A(n6503), .B(n6504), .Z(n6502) );
  NANDN U6500 ( .A(n6505), .B(n6506), .Z(n6504) );
  NANDN U6501 ( .A(n6506), .B(n6505), .Z(n6501) );
  ANDN U6502 ( .B(B[30]), .A(n56), .Z(n6285) );
  XNOR U6503 ( .A(n6293), .B(n6507), .Z(n6286) );
  XNOR U6504 ( .A(n6292), .B(n6290), .Z(n6507) );
  AND U6505 ( .A(n6508), .B(n6509), .Z(n6290) );
  NANDN U6506 ( .A(n6510), .B(n6511), .Z(n6509) );
  OR U6507 ( .A(n6512), .B(n6513), .Z(n6511) );
  NAND U6508 ( .A(n6513), .B(n6512), .Z(n6508) );
  ANDN U6509 ( .B(B[31]), .A(n57), .Z(n6292) );
  XNOR U6510 ( .A(n6300), .B(n6514), .Z(n6293) );
  XNOR U6511 ( .A(n6299), .B(n6297), .Z(n6514) );
  AND U6512 ( .A(n6515), .B(n6516), .Z(n6297) );
  NANDN U6513 ( .A(n6517), .B(n6518), .Z(n6516) );
  NANDN U6514 ( .A(n6519), .B(n6520), .Z(n6518) );
  NANDN U6515 ( .A(n6520), .B(n6519), .Z(n6515) );
  ANDN U6516 ( .B(B[32]), .A(n58), .Z(n6299) );
  XNOR U6517 ( .A(n6307), .B(n6521), .Z(n6300) );
  XNOR U6518 ( .A(n6306), .B(n6304), .Z(n6521) );
  AND U6519 ( .A(n6522), .B(n6523), .Z(n6304) );
  NANDN U6520 ( .A(n6524), .B(n6525), .Z(n6523) );
  OR U6521 ( .A(n6526), .B(n6527), .Z(n6525) );
  NAND U6522 ( .A(n6527), .B(n6526), .Z(n6522) );
  ANDN U6523 ( .B(B[33]), .A(n59), .Z(n6306) );
  XNOR U6524 ( .A(n6314), .B(n6528), .Z(n6307) );
  XNOR U6525 ( .A(n6313), .B(n6311), .Z(n6528) );
  AND U6526 ( .A(n6529), .B(n6530), .Z(n6311) );
  NANDN U6527 ( .A(n6531), .B(n6532), .Z(n6530) );
  NANDN U6528 ( .A(n6533), .B(n6534), .Z(n6532) );
  NANDN U6529 ( .A(n6534), .B(n6533), .Z(n6529) );
  ANDN U6530 ( .B(B[34]), .A(n60), .Z(n6313) );
  XNOR U6531 ( .A(n6321), .B(n6535), .Z(n6314) );
  XNOR U6532 ( .A(n6320), .B(n6318), .Z(n6535) );
  AND U6533 ( .A(n6536), .B(n6537), .Z(n6318) );
  NANDN U6534 ( .A(n6538), .B(n6539), .Z(n6537) );
  OR U6535 ( .A(n6540), .B(n6541), .Z(n6539) );
  NAND U6536 ( .A(n6541), .B(n6540), .Z(n6536) );
  ANDN U6537 ( .B(B[35]), .A(n61), .Z(n6320) );
  XNOR U6538 ( .A(n6328), .B(n6542), .Z(n6321) );
  XNOR U6539 ( .A(n6327), .B(n6325), .Z(n6542) );
  AND U6540 ( .A(n6543), .B(n6544), .Z(n6325) );
  NANDN U6541 ( .A(n6545), .B(n6546), .Z(n6544) );
  NANDN U6542 ( .A(n6547), .B(n6548), .Z(n6546) );
  NANDN U6543 ( .A(n6548), .B(n6547), .Z(n6543) );
  ANDN U6544 ( .B(B[36]), .A(n62), .Z(n6327) );
  XNOR U6545 ( .A(n6335), .B(n6549), .Z(n6328) );
  XNOR U6546 ( .A(n6334), .B(n6332), .Z(n6549) );
  AND U6547 ( .A(n6550), .B(n6551), .Z(n6332) );
  NANDN U6548 ( .A(n6552), .B(n6553), .Z(n6551) );
  OR U6549 ( .A(n6554), .B(n6555), .Z(n6553) );
  NAND U6550 ( .A(n6555), .B(n6554), .Z(n6550) );
  ANDN U6551 ( .B(B[37]), .A(n63), .Z(n6334) );
  XNOR U6552 ( .A(n6342), .B(n6556), .Z(n6335) );
  XNOR U6553 ( .A(n6341), .B(n6339), .Z(n6556) );
  AND U6554 ( .A(n6557), .B(n6558), .Z(n6339) );
  NANDN U6555 ( .A(n6559), .B(n6560), .Z(n6558) );
  NANDN U6556 ( .A(n6561), .B(n6562), .Z(n6560) );
  NANDN U6557 ( .A(n6562), .B(n6561), .Z(n6557) );
  ANDN U6558 ( .B(B[38]), .A(n64), .Z(n6341) );
  XNOR U6559 ( .A(n6349), .B(n6563), .Z(n6342) );
  XNOR U6560 ( .A(n6348), .B(n6346), .Z(n6563) );
  AND U6561 ( .A(n6564), .B(n6565), .Z(n6346) );
  NANDN U6562 ( .A(n6566), .B(n6567), .Z(n6565) );
  OR U6563 ( .A(n6568), .B(n6569), .Z(n6567) );
  NAND U6564 ( .A(n6569), .B(n6568), .Z(n6564) );
  ANDN U6565 ( .B(B[39]), .A(n65), .Z(n6348) );
  XNOR U6566 ( .A(n6356), .B(n6570), .Z(n6349) );
  XNOR U6567 ( .A(n6355), .B(n6353), .Z(n6570) );
  AND U6568 ( .A(n6571), .B(n6572), .Z(n6353) );
  NANDN U6569 ( .A(n6573), .B(n6574), .Z(n6572) );
  NANDN U6570 ( .A(n6575), .B(n6576), .Z(n6574) );
  NANDN U6571 ( .A(n6576), .B(n6575), .Z(n6571) );
  ANDN U6572 ( .B(B[40]), .A(n66), .Z(n6355) );
  XNOR U6573 ( .A(n6363), .B(n6577), .Z(n6356) );
  XNOR U6574 ( .A(n6362), .B(n6360), .Z(n6577) );
  AND U6575 ( .A(n6578), .B(n6579), .Z(n6360) );
  NANDN U6576 ( .A(n6580), .B(n6581), .Z(n6579) );
  OR U6577 ( .A(n6582), .B(n6583), .Z(n6581) );
  NAND U6578 ( .A(n6583), .B(n6582), .Z(n6578) );
  ANDN U6579 ( .B(B[41]), .A(n67), .Z(n6362) );
  XNOR U6580 ( .A(n6370), .B(n6584), .Z(n6363) );
  XNOR U6581 ( .A(n6369), .B(n6367), .Z(n6584) );
  AND U6582 ( .A(n6585), .B(n6586), .Z(n6367) );
  NANDN U6583 ( .A(n6587), .B(n6588), .Z(n6586) );
  NANDN U6584 ( .A(n6589), .B(n6590), .Z(n6588) );
  NANDN U6585 ( .A(n6590), .B(n6589), .Z(n6585) );
  ANDN U6586 ( .B(B[42]), .A(n68), .Z(n6369) );
  XNOR U6587 ( .A(n6377), .B(n6591), .Z(n6370) );
  XNOR U6588 ( .A(n6376), .B(n6374), .Z(n6591) );
  AND U6589 ( .A(n6592), .B(n6593), .Z(n6374) );
  NANDN U6590 ( .A(n6594), .B(n6595), .Z(n6593) );
  OR U6591 ( .A(n6596), .B(n6597), .Z(n6595) );
  NAND U6592 ( .A(n6597), .B(n6596), .Z(n6592) );
  ANDN U6593 ( .B(B[43]), .A(n69), .Z(n6376) );
  XNOR U6594 ( .A(n6384), .B(n6598), .Z(n6377) );
  XNOR U6595 ( .A(n6383), .B(n6381), .Z(n6598) );
  AND U6596 ( .A(n6599), .B(n6600), .Z(n6381) );
  NANDN U6597 ( .A(n6601), .B(n6602), .Z(n6600) );
  NANDN U6598 ( .A(n6603), .B(n6604), .Z(n6602) );
  NANDN U6599 ( .A(n6604), .B(n6603), .Z(n6599) );
  ANDN U6600 ( .B(B[44]), .A(n70), .Z(n6383) );
  XNOR U6601 ( .A(n6391), .B(n6605), .Z(n6384) );
  XNOR U6602 ( .A(n6390), .B(n6388), .Z(n6605) );
  AND U6603 ( .A(n6606), .B(n6607), .Z(n6388) );
  NANDN U6604 ( .A(n6608), .B(n6609), .Z(n6607) );
  OR U6605 ( .A(n6610), .B(n6611), .Z(n6609) );
  NAND U6606 ( .A(n6611), .B(n6610), .Z(n6606) );
  ANDN U6607 ( .B(B[45]), .A(n71), .Z(n6390) );
  XNOR U6608 ( .A(n6398), .B(n6612), .Z(n6391) );
  XNOR U6609 ( .A(n6397), .B(n6395), .Z(n6612) );
  AND U6610 ( .A(n6613), .B(n6614), .Z(n6395) );
  NANDN U6611 ( .A(n6615), .B(n6616), .Z(n6614) );
  NANDN U6612 ( .A(n6617), .B(n6618), .Z(n6616) );
  NANDN U6613 ( .A(n6618), .B(n6617), .Z(n6613) );
  ANDN U6614 ( .B(B[46]), .A(n72), .Z(n6397) );
  XNOR U6615 ( .A(n6405), .B(n6619), .Z(n6398) );
  XNOR U6616 ( .A(n6404), .B(n6402), .Z(n6619) );
  AND U6617 ( .A(n6620), .B(n6621), .Z(n6402) );
  NANDN U6618 ( .A(n6622), .B(n6623), .Z(n6621) );
  OR U6619 ( .A(n6624), .B(n6625), .Z(n6623) );
  NAND U6620 ( .A(n6625), .B(n6624), .Z(n6620) );
  ANDN U6621 ( .B(B[47]), .A(n73), .Z(n6404) );
  XNOR U6622 ( .A(n6412), .B(n6626), .Z(n6405) );
  XNOR U6623 ( .A(n6411), .B(n6409), .Z(n6626) );
  AND U6624 ( .A(n6627), .B(n6628), .Z(n6409) );
  NANDN U6625 ( .A(n6629), .B(n6630), .Z(n6628) );
  NANDN U6626 ( .A(n6631), .B(n6632), .Z(n6630) );
  NANDN U6627 ( .A(n6632), .B(n6631), .Z(n6627) );
  ANDN U6628 ( .B(B[48]), .A(n74), .Z(n6411) );
  XNOR U6629 ( .A(n6419), .B(n6633), .Z(n6412) );
  XNOR U6630 ( .A(n6418), .B(n6416), .Z(n6633) );
  AND U6631 ( .A(n6634), .B(n6635), .Z(n6416) );
  NANDN U6632 ( .A(n6636), .B(n6637), .Z(n6635) );
  OR U6633 ( .A(n6638), .B(n6639), .Z(n6637) );
  NAND U6634 ( .A(n6639), .B(n6638), .Z(n6634) );
  ANDN U6635 ( .B(B[49]), .A(n75), .Z(n6418) );
  XNOR U6636 ( .A(n6426), .B(n6640), .Z(n6419) );
  XNOR U6637 ( .A(n6425), .B(n6423), .Z(n6640) );
  AND U6638 ( .A(n6641), .B(n6642), .Z(n6423) );
  NANDN U6639 ( .A(n6643), .B(n6644), .Z(n6642) );
  NANDN U6640 ( .A(n6645), .B(n6646), .Z(n6644) );
  NANDN U6641 ( .A(n6646), .B(n6645), .Z(n6641) );
  ANDN U6642 ( .B(B[50]), .A(n76), .Z(n6425) );
  XNOR U6643 ( .A(n6433), .B(n6647), .Z(n6426) );
  XNOR U6644 ( .A(n6432), .B(n6430), .Z(n6647) );
  AND U6645 ( .A(n6648), .B(n6649), .Z(n6430) );
  NANDN U6646 ( .A(n6650), .B(n6651), .Z(n6649) );
  OR U6647 ( .A(n6652), .B(n6653), .Z(n6651) );
  NAND U6648 ( .A(n6653), .B(n6652), .Z(n6648) );
  ANDN U6649 ( .B(B[51]), .A(n77), .Z(n6432) );
  XNOR U6650 ( .A(n6440), .B(n6654), .Z(n6433) );
  XNOR U6651 ( .A(n6439), .B(n6437), .Z(n6654) );
  AND U6652 ( .A(n6655), .B(n6656), .Z(n6437) );
  NANDN U6653 ( .A(n6657), .B(n6658), .Z(n6656) );
  NANDN U6654 ( .A(n6659), .B(n6660), .Z(n6658) );
  NANDN U6655 ( .A(n6660), .B(n6659), .Z(n6655) );
  ANDN U6656 ( .B(B[52]), .A(n78), .Z(n6439) );
  XNOR U6657 ( .A(n6447), .B(n6661), .Z(n6440) );
  XNOR U6658 ( .A(n6446), .B(n6444), .Z(n6661) );
  AND U6659 ( .A(n6662), .B(n6663), .Z(n6444) );
  NANDN U6660 ( .A(n6664), .B(n6665), .Z(n6663) );
  OR U6661 ( .A(n6666), .B(n6667), .Z(n6665) );
  NAND U6662 ( .A(n6667), .B(n6666), .Z(n6662) );
  ANDN U6663 ( .B(B[53]), .A(n79), .Z(n6446) );
  XNOR U6664 ( .A(n6454), .B(n6668), .Z(n6447) );
  XNOR U6665 ( .A(n6453), .B(n6451), .Z(n6668) );
  AND U6666 ( .A(n6669), .B(n6670), .Z(n6451) );
  NANDN U6667 ( .A(n6671), .B(n6672), .Z(n6670) );
  NANDN U6668 ( .A(n6673), .B(n6674), .Z(n6672) );
  NANDN U6669 ( .A(n6674), .B(n6673), .Z(n6669) );
  ANDN U6670 ( .B(B[54]), .A(n80), .Z(n6453) );
  XNOR U6671 ( .A(n6461), .B(n6675), .Z(n6454) );
  XNOR U6672 ( .A(n6460), .B(n6458), .Z(n6675) );
  AND U6673 ( .A(n6676), .B(n6677), .Z(n6458) );
  NANDN U6674 ( .A(n6678), .B(n6679), .Z(n6677) );
  OR U6675 ( .A(n6680), .B(n6681), .Z(n6679) );
  NAND U6676 ( .A(n6681), .B(n6680), .Z(n6676) );
  ANDN U6677 ( .B(B[55]), .A(n81), .Z(n6460) );
  XNOR U6678 ( .A(n6468), .B(n6682), .Z(n6461) );
  XNOR U6679 ( .A(n6467), .B(n6465), .Z(n6682) );
  AND U6680 ( .A(n6683), .B(n6684), .Z(n6465) );
  NANDN U6681 ( .A(n6685), .B(n6686), .Z(n6684) );
  NAND U6682 ( .A(n6687), .B(n6688), .Z(n6686) );
  ANDN U6683 ( .B(B[56]), .A(n82), .Z(n6467) );
  XOR U6684 ( .A(n6474), .B(n6689), .Z(n6468) );
  XNOR U6685 ( .A(n6472), .B(n6475), .Z(n6689) );
  NAND U6686 ( .A(A[2]), .B(B[57]), .Z(n6475) );
  NANDN U6687 ( .A(n6690), .B(n6691), .Z(n6472) );
  AND U6688 ( .A(A[0]), .B(B[58]), .Z(n6691) );
  XNOR U6689 ( .A(n6477), .B(n6692), .Z(n6474) );
  NAND U6690 ( .A(A[0]), .B(B[59]), .Z(n6692) );
  NAND U6691 ( .A(B[58]), .B(A[1]), .Z(n6477) );
  NAND U6692 ( .A(n6693), .B(n6694), .Z(n169) );
  NANDN U6693 ( .A(n6695), .B(n6696), .Z(n6694) );
  OR U6694 ( .A(n6697), .B(n6698), .Z(n6696) );
  NAND U6695 ( .A(n6698), .B(n6697), .Z(n6693) );
  XOR U6696 ( .A(n171), .B(n170), .Z(\A1[56] ) );
  XOR U6697 ( .A(n6698), .B(n6699), .Z(n170) );
  XNOR U6698 ( .A(n6697), .B(n6695), .Z(n6699) );
  AND U6699 ( .A(n6700), .B(n6701), .Z(n6695) );
  NANDN U6700 ( .A(n6702), .B(n6703), .Z(n6701) );
  NANDN U6701 ( .A(n6704), .B(n6705), .Z(n6703) );
  NANDN U6702 ( .A(n6705), .B(n6704), .Z(n6700) );
  ANDN U6703 ( .B(B[27]), .A(n54), .Z(n6697) );
  XNOR U6704 ( .A(n6492), .B(n6706), .Z(n6698) );
  XNOR U6705 ( .A(n6491), .B(n6489), .Z(n6706) );
  AND U6706 ( .A(n6707), .B(n6708), .Z(n6489) );
  NANDN U6707 ( .A(n6709), .B(n6710), .Z(n6708) );
  OR U6708 ( .A(n6711), .B(n6712), .Z(n6710) );
  NAND U6709 ( .A(n6712), .B(n6711), .Z(n6707) );
  ANDN U6710 ( .B(B[28]), .A(n55), .Z(n6491) );
  XNOR U6711 ( .A(n6499), .B(n6713), .Z(n6492) );
  XNOR U6712 ( .A(n6498), .B(n6496), .Z(n6713) );
  AND U6713 ( .A(n6714), .B(n6715), .Z(n6496) );
  NANDN U6714 ( .A(n6716), .B(n6717), .Z(n6715) );
  NANDN U6715 ( .A(n6718), .B(n6719), .Z(n6717) );
  NANDN U6716 ( .A(n6719), .B(n6718), .Z(n6714) );
  ANDN U6717 ( .B(B[29]), .A(n56), .Z(n6498) );
  XNOR U6718 ( .A(n6506), .B(n6720), .Z(n6499) );
  XNOR U6719 ( .A(n6505), .B(n6503), .Z(n6720) );
  AND U6720 ( .A(n6721), .B(n6722), .Z(n6503) );
  NANDN U6721 ( .A(n6723), .B(n6724), .Z(n6722) );
  OR U6722 ( .A(n6725), .B(n6726), .Z(n6724) );
  NAND U6723 ( .A(n6726), .B(n6725), .Z(n6721) );
  ANDN U6724 ( .B(B[30]), .A(n57), .Z(n6505) );
  XNOR U6725 ( .A(n6513), .B(n6727), .Z(n6506) );
  XNOR U6726 ( .A(n6512), .B(n6510), .Z(n6727) );
  AND U6727 ( .A(n6728), .B(n6729), .Z(n6510) );
  NANDN U6728 ( .A(n6730), .B(n6731), .Z(n6729) );
  NANDN U6729 ( .A(n6732), .B(n6733), .Z(n6731) );
  NANDN U6730 ( .A(n6733), .B(n6732), .Z(n6728) );
  ANDN U6731 ( .B(B[31]), .A(n58), .Z(n6512) );
  XNOR U6732 ( .A(n6520), .B(n6734), .Z(n6513) );
  XNOR U6733 ( .A(n6519), .B(n6517), .Z(n6734) );
  AND U6734 ( .A(n6735), .B(n6736), .Z(n6517) );
  NANDN U6735 ( .A(n6737), .B(n6738), .Z(n6736) );
  OR U6736 ( .A(n6739), .B(n6740), .Z(n6738) );
  NAND U6737 ( .A(n6740), .B(n6739), .Z(n6735) );
  ANDN U6738 ( .B(B[32]), .A(n59), .Z(n6519) );
  XNOR U6739 ( .A(n6527), .B(n6741), .Z(n6520) );
  XNOR U6740 ( .A(n6526), .B(n6524), .Z(n6741) );
  AND U6741 ( .A(n6742), .B(n6743), .Z(n6524) );
  NANDN U6742 ( .A(n6744), .B(n6745), .Z(n6743) );
  NANDN U6743 ( .A(n6746), .B(n6747), .Z(n6745) );
  NANDN U6744 ( .A(n6747), .B(n6746), .Z(n6742) );
  ANDN U6745 ( .B(B[33]), .A(n60), .Z(n6526) );
  XNOR U6746 ( .A(n6534), .B(n6748), .Z(n6527) );
  XNOR U6747 ( .A(n6533), .B(n6531), .Z(n6748) );
  AND U6748 ( .A(n6749), .B(n6750), .Z(n6531) );
  NANDN U6749 ( .A(n6751), .B(n6752), .Z(n6750) );
  OR U6750 ( .A(n6753), .B(n6754), .Z(n6752) );
  NAND U6751 ( .A(n6754), .B(n6753), .Z(n6749) );
  ANDN U6752 ( .B(B[34]), .A(n61), .Z(n6533) );
  XNOR U6753 ( .A(n6541), .B(n6755), .Z(n6534) );
  XNOR U6754 ( .A(n6540), .B(n6538), .Z(n6755) );
  AND U6755 ( .A(n6756), .B(n6757), .Z(n6538) );
  NANDN U6756 ( .A(n6758), .B(n6759), .Z(n6757) );
  NANDN U6757 ( .A(n6760), .B(n6761), .Z(n6759) );
  NANDN U6758 ( .A(n6761), .B(n6760), .Z(n6756) );
  ANDN U6759 ( .B(B[35]), .A(n62), .Z(n6540) );
  XNOR U6760 ( .A(n6548), .B(n6762), .Z(n6541) );
  XNOR U6761 ( .A(n6547), .B(n6545), .Z(n6762) );
  AND U6762 ( .A(n6763), .B(n6764), .Z(n6545) );
  NANDN U6763 ( .A(n6765), .B(n6766), .Z(n6764) );
  OR U6764 ( .A(n6767), .B(n6768), .Z(n6766) );
  NAND U6765 ( .A(n6768), .B(n6767), .Z(n6763) );
  ANDN U6766 ( .B(B[36]), .A(n63), .Z(n6547) );
  XNOR U6767 ( .A(n6555), .B(n6769), .Z(n6548) );
  XNOR U6768 ( .A(n6554), .B(n6552), .Z(n6769) );
  AND U6769 ( .A(n6770), .B(n6771), .Z(n6552) );
  NANDN U6770 ( .A(n6772), .B(n6773), .Z(n6771) );
  NANDN U6771 ( .A(n6774), .B(n6775), .Z(n6773) );
  NANDN U6772 ( .A(n6775), .B(n6774), .Z(n6770) );
  ANDN U6773 ( .B(B[37]), .A(n64), .Z(n6554) );
  XNOR U6774 ( .A(n6562), .B(n6776), .Z(n6555) );
  XNOR U6775 ( .A(n6561), .B(n6559), .Z(n6776) );
  AND U6776 ( .A(n6777), .B(n6778), .Z(n6559) );
  NANDN U6777 ( .A(n6779), .B(n6780), .Z(n6778) );
  OR U6778 ( .A(n6781), .B(n6782), .Z(n6780) );
  NAND U6779 ( .A(n6782), .B(n6781), .Z(n6777) );
  ANDN U6780 ( .B(B[38]), .A(n65), .Z(n6561) );
  XNOR U6781 ( .A(n6569), .B(n6783), .Z(n6562) );
  XNOR U6782 ( .A(n6568), .B(n6566), .Z(n6783) );
  AND U6783 ( .A(n6784), .B(n6785), .Z(n6566) );
  NANDN U6784 ( .A(n6786), .B(n6787), .Z(n6785) );
  NANDN U6785 ( .A(n6788), .B(n6789), .Z(n6787) );
  NANDN U6786 ( .A(n6789), .B(n6788), .Z(n6784) );
  ANDN U6787 ( .B(B[39]), .A(n66), .Z(n6568) );
  XNOR U6788 ( .A(n6576), .B(n6790), .Z(n6569) );
  XNOR U6789 ( .A(n6575), .B(n6573), .Z(n6790) );
  AND U6790 ( .A(n6791), .B(n6792), .Z(n6573) );
  NANDN U6791 ( .A(n6793), .B(n6794), .Z(n6792) );
  OR U6792 ( .A(n6795), .B(n6796), .Z(n6794) );
  NAND U6793 ( .A(n6796), .B(n6795), .Z(n6791) );
  ANDN U6794 ( .B(B[40]), .A(n67), .Z(n6575) );
  XNOR U6795 ( .A(n6583), .B(n6797), .Z(n6576) );
  XNOR U6796 ( .A(n6582), .B(n6580), .Z(n6797) );
  AND U6797 ( .A(n6798), .B(n6799), .Z(n6580) );
  NANDN U6798 ( .A(n6800), .B(n6801), .Z(n6799) );
  NANDN U6799 ( .A(n6802), .B(n6803), .Z(n6801) );
  NANDN U6800 ( .A(n6803), .B(n6802), .Z(n6798) );
  ANDN U6801 ( .B(B[41]), .A(n68), .Z(n6582) );
  XNOR U6802 ( .A(n6590), .B(n6804), .Z(n6583) );
  XNOR U6803 ( .A(n6589), .B(n6587), .Z(n6804) );
  AND U6804 ( .A(n6805), .B(n6806), .Z(n6587) );
  NANDN U6805 ( .A(n6807), .B(n6808), .Z(n6806) );
  OR U6806 ( .A(n6809), .B(n6810), .Z(n6808) );
  NAND U6807 ( .A(n6810), .B(n6809), .Z(n6805) );
  ANDN U6808 ( .B(B[42]), .A(n69), .Z(n6589) );
  XNOR U6809 ( .A(n6597), .B(n6811), .Z(n6590) );
  XNOR U6810 ( .A(n6596), .B(n6594), .Z(n6811) );
  AND U6811 ( .A(n6812), .B(n6813), .Z(n6594) );
  NANDN U6812 ( .A(n6814), .B(n6815), .Z(n6813) );
  NANDN U6813 ( .A(n6816), .B(n6817), .Z(n6815) );
  NANDN U6814 ( .A(n6817), .B(n6816), .Z(n6812) );
  ANDN U6815 ( .B(B[43]), .A(n70), .Z(n6596) );
  XNOR U6816 ( .A(n6604), .B(n6818), .Z(n6597) );
  XNOR U6817 ( .A(n6603), .B(n6601), .Z(n6818) );
  AND U6818 ( .A(n6819), .B(n6820), .Z(n6601) );
  NANDN U6819 ( .A(n6821), .B(n6822), .Z(n6820) );
  OR U6820 ( .A(n6823), .B(n6824), .Z(n6822) );
  NAND U6821 ( .A(n6824), .B(n6823), .Z(n6819) );
  ANDN U6822 ( .B(B[44]), .A(n71), .Z(n6603) );
  XNOR U6823 ( .A(n6611), .B(n6825), .Z(n6604) );
  XNOR U6824 ( .A(n6610), .B(n6608), .Z(n6825) );
  AND U6825 ( .A(n6826), .B(n6827), .Z(n6608) );
  NANDN U6826 ( .A(n6828), .B(n6829), .Z(n6827) );
  NANDN U6827 ( .A(n6830), .B(n6831), .Z(n6829) );
  NANDN U6828 ( .A(n6831), .B(n6830), .Z(n6826) );
  ANDN U6829 ( .B(B[45]), .A(n72), .Z(n6610) );
  XNOR U6830 ( .A(n6618), .B(n6832), .Z(n6611) );
  XNOR U6831 ( .A(n6617), .B(n6615), .Z(n6832) );
  AND U6832 ( .A(n6833), .B(n6834), .Z(n6615) );
  NANDN U6833 ( .A(n6835), .B(n6836), .Z(n6834) );
  OR U6834 ( .A(n6837), .B(n6838), .Z(n6836) );
  NAND U6835 ( .A(n6838), .B(n6837), .Z(n6833) );
  ANDN U6836 ( .B(B[46]), .A(n73), .Z(n6617) );
  XNOR U6837 ( .A(n6625), .B(n6839), .Z(n6618) );
  XNOR U6838 ( .A(n6624), .B(n6622), .Z(n6839) );
  AND U6839 ( .A(n6840), .B(n6841), .Z(n6622) );
  NANDN U6840 ( .A(n6842), .B(n6843), .Z(n6841) );
  NANDN U6841 ( .A(n6844), .B(n6845), .Z(n6843) );
  NANDN U6842 ( .A(n6845), .B(n6844), .Z(n6840) );
  ANDN U6843 ( .B(B[47]), .A(n74), .Z(n6624) );
  XNOR U6844 ( .A(n6632), .B(n6846), .Z(n6625) );
  XNOR U6845 ( .A(n6631), .B(n6629), .Z(n6846) );
  AND U6846 ( .A(n6847), .B(n6848), .Z(n6629) );
  NANDN U6847 ( .A(n6849), .B(n6850), .Z(n6848) );
  OR U6848 ( .A(n6851), .B(n6852), .Z(n6850) );
  NAND U6849 ( .A(n6852), .B(n6851), .Z(n6847) );
  ANDN U6850 ( .B(B[48]), .A(n75), .Z(n6631) );
  XNOR U6851 ( .A(n6639), .B(n6853), .Z(n6632) );
  XNOR U6852 ( .A(n6638), .B(n6636), .Z(n6853) );
  AND U6853 ( .A(n6854), .B(n6855), .Z(n6636) );
  NANDN U6854 ( .A(n6856), .B(n6857), .Z(n6855) );
  NANDN U6855 ( .A(n6858), .B(n6859), .Z(n6857) );
  NANDN U6856 ( .A(n6859), .B(n6858), .Z(n6854) );
  ANDN U6857 ( .B(B[49]), .A(n76), .Z(n6638) );
  XNOR U6858 ( .A(n6646), .B(n6860), .Z(n6639) );
  XNOR U6859 ( .A(n6645), .B(n6643), .Z(n6860) );
  AND U6860 ( .A(n6861), .B(n6862), .Z(n6643) );
  NANDN U6861 ( .A(n6863), .B(n6864), .Z(n6862) );
  OR U6862 ( .A(n6865), .B(n6866), .Z(n6864) );
  NAND U6863 ( .A(n6866), .B(n6865), .Z(n6861) );
  ANDN U6864 ( .B(B[50]), .A(n77), .Z(n6645) );
  XNOR U6865 ( .A(n6653), .B(n6867), .Z(n6646) );
  XNOR U6866 ( .A(n6652), .B(n6650), .Z(n6867) );
  AND U6867 ( .A(n6868), .B(n6869), .Z(n6650) );
  NANDN U6868 ( .A(n6870), .B(n6871), .Z(n6869) );
  NANDN U6869 ( .A(n6872), .B(n6873), .Z(n6871) );
  NANDN U6870 ( .A(n6873), .B(n6872), .Z(n6868) );
  ANDN U6871 ( .B(B[51]), .A(n78), .Z(n6652) );
  XNOR U6872 ( .A(n6660), .B(n6874), .Z(n6653) );
  XNOR U6873 ( .A(n6659), .B(n6657), .Z(n6874) );
  AND U6874 ( .A(n6875), .B(n6876), .Z(n6657) );
  NANDN U6875 ( .A(n6877), .B(n6878), .Z(n6876) );
  OR U6876 ( .A(n6879), .B(n6880), .Z(n6878) );
  NAND U6877 ( .A(n6880), .B(n6879), .Z(n6875) );
  ANDN U6878 ( .B(B[52]), .A(n79), .Z(n6659) );
  XNOR U6879 ( .A(n6667), .B(n6881), .Z(n6660) );
  XNOR U6880 ( .A(n6666), .B(n6664), .Z(n6881) );
  AND U6881 ( .A(n6882), .B(n6883), .Z(n6664) );
  NANDN U6882 ( .A(n6884), .B(n6885), .Z(n6883) );
  NANDN U6883 ( .A(n6886), .B(n6887), .Z(n6885) );
  NANDN U6884 ( .A(n6887), .B(n6886), .Z(n6882) );
  ANDN U6885 ( .B(B[53]), .A(n80), .Z(n6666) );
  XNOR U6886 ( .A(n6674), .B(n6888), .Z(n6667) );
  XNOR U6887 ( .A(n6673), .B(n6671), .Z(n6888) );
  AND U6888 ( .A(n6889), .B(n6890), .Z(n6671) );
  NANDN U6889 ( .A(n6891), .B(n6892), .Z(n6890) );
  OR U6890 ( .A(n6893), .B(n6894), .Z(n6892) );
  NAND U6891 ( .A(n6894), .B(n6893), .Z(n6889) );
  ANDN U6892 ( .B(B[54]), .A(n81), .Z(n6673) );
  XNOR U6893 ( .A(n6681), .B(n6895), .Z(n6674) );
  XNOR U6894 ( .A(n6680), .B(n6678), .Z(n6895) );
  AND U6895 ( .A(n6896), .B(n6897), .Z(n6678) );
  NANDN U6896 ( .A(n6898), .B(n6899), .Z(n6897) );
  NAND U6897 ( .A(n6900), .B(n6901), .Z(n6899) );
  ANDN U6898 ( .B(B[55]), .A(n82), .Z(n6680) );
  XOR U6899 ( .A(n6687), .B(n6902), .Z(n6681) );
  XNOR U6900 ( .A(n6685), .B(n6688), .Z(n6902) );
  NAND U6901 ( .A(A[2]), .B(B[56]), .Z(n6688) );
  NANDN U6902 ( .A(n6903), .B(n6904), .Z(n6685) );
  AND U6903 ( .A(A[0]), .B(B[57]), .Z(n6904) );
  XNOR U6904 ( .A(n6690), .B(n6905), .Z(n6687) );
  NAND U6905 ( .A(A[0]), .B(B[58]), .Z(n6905) );
  NAND U6906 ( .A(B[57]), .B(A[1]), .Z(n6690) );
  NAND U6907 ( .A(n6906), .B(n6907), .Z(n171) );
  NANDN U6908 ( .A(n6908), .B(n6909), .Z(n6907) );
  OR U6909 ( .A(n6910), .B(n6911), .Z(n6909) );
  NAND U6910 ( .A(n6911), .B(n6910), .Z(n6906) );
  XOR U6911 ( .A(n173), .B(n172), .Z(\A1[55] ) );
  XOR U6912 ( .A(n6911), .B(n6912), .Z(n172) );
  XNOR U6913 ( .A(n6910), .B(n6908), .Z(n6912) );
  AND U6914 ( .A(n6913), .B(n6914), .Z(n6908) );
  NANDN U6915 ( .A(n6915), .B(n6916), .Z(n6914) );
  NANDN U6916 ( .A(n6917), .B(n6918), .Z(n6916) );
  NANDN U6917 ( .A(n6918), .B(n6917), .Z(n6913) );
  ANDN U6918 ( .B(B[26]), .A(n54), .Z(n6910) );
  XNOR U6919 ( .A(n6705), .B(n6919), .Z(n6911) );
  XNOR U6920 ( .A(n6704), .B(n6702), .Z(n6919) );
  AND U6921 ( .A(n6920), .B(n6921), .Z(n6702) );
  NANDN U6922 ( .A(n6922), .B(n6923), .Z(n6921) );
  OR U6923 ( .A(n6924), .B(n6925), .Z(n6923) );
  NAND U6924 ( .A(n6925), .B(n6924), .Z(n6920) );
  ANDN U6925 ( .B(B[27]), .A(n55), .Z(n6704) );
  XNOR U6926 ( .A(n6712), .B(n6926), .Z(n6705) );
  XNOR U6927 ( .A(n6711), .B(n6709), .Z(n6926) );
  AND U6928 ( .A(n6927), .B(n6928), .Z(n6709) );
  NANDN U6929 ( .A(n6929), .B(n6930), .Z(n6928) );
  NANDN U6930 ( .A(n6931), .B(n6932), .Z(n6930) );
  NANDN U6931 ( .A(n6932), .B(n6931), .Z(n6927) );
  ANDN U6932 ( .B(B[28]), .A(n56), .Z(n6711) );
  XNOR U6933 ( .A(n6719), .B(n6933), .Z(n6712) );
  XNOR U6934 ( .A(n6718), .B(n6716), .Z(n6933) );
  AND U6935 ( .A(n6934), .B(n6935), .Z(n6716) );
  NANDN U6936 ( .A(n6936), .B(n6937), .Z(n6935) );
  OR U6937 ( .A(n6938), .B(n6939), .Z(n6937) );
  NAND U6938 ( .A(n6939), .B(n6938), .Z(n6934) );
  ANDN U6939 ( .B(B[29]), .A(n57), .Z(n6718) );
  XNOR U6940 ( .A(n6726), .B(n6940), .Z(n6719) );
  XNOR U6941 ( .A(n6725), .B(n6723), .Z(n6940) );
  AND U6942 ( .A(n6941), .B(n6942), .Z(n6723) );
  NANDN U6943 ( .A(n6943), .B(n6944), .Z(n6942) );
  NANDN U6944 ( .A(n6945), .B(n6946), .Z(n6944) );
  NANDN U6945 ( .A(n6946), .B(n6945), .Z(n6941) );
  ANDN U6946 ( .B(B[30]), .A(n58), .Z(n6725) );
  XNOR U6947 ( .A(n6733), .B(n6947), .Z(n6726) );
  XNOR U6948 ( .A(n6732), .B(n6730), .Z(n6947) );
  AND U6949 ( .A(n6948), .B(n6949), .Z(n6730) );
  NANDN U6950 ( .A(n6950), .B(n6951), .Z(n6949) );
  OR U6951 ( .A(n6952), .B(n6953), .Z(n6951) );
  NAND U6952 ( .A(n6953), .B(n6952), .Z(n6948) );
  ANDN U6953 ( .B(B[31]), .A(n59), .Z(n6732) );
  XNOR U6954 ( .A(n6740), .B(n6954), .Z(n6733) );
  XNOR U6955 ( .A(n6739), .B(n6737), .Z(n6954) );
  AND U6956 ( .A(n6955), .B(n6956), .Z(n6737) );
  NANDN U6957 ( .A(n6957), .B(n6958), .Z(n6956) );
  NANDN U6958 ( .A(n6959), .B(n6960), .Z(n6958) );
  NANDN U6959 ( .A(n6960), .B(n6959), .Z(n6955) );
  ANDN U6960 ( .B(B[32]), .A(n60), .Z(n6739) );
  XNOR U6961 ( .A(n6747), .B(n6961), .Z(n6740) );
  XNOR U6962 ( .A(n6746), .B(n6744), .Z(n6961) );
  AND U6963 ( .A(n6962), .B(n6963), .Z(n6744) );
  NANDN U6964 ( .A(n6964), .B(n6965), .Z(n6963) );
  OR U6965 ( .A(n6966), .B(n6967), .Z(n6965) );
  NAND U6966 ( .A(n6967), .B(n6966), .Z(n6962) );
  ANDN U6967 ( .B(B[33]), .A(n61), .Z(n6746) );
  XNOR U6968 ( .A(n6754), .B(n6968), .Z(n6747) );
  XNOR U6969 ( .A(n6753), .B(n6751), .Z(n6968) );
  AND U6970 ( .A(n6969), .B(n6970), .Z(n6751) );
  NANDN U6971 ( .A(n6971), .B(n6972), .Z(n6970) );
  NANDN U6972 ( .A(n6973), .B(n6974), .Z(n6972) );
  NANDN U6973 ( .A(n6974), .B(n6973), .Z(n6969) );
  ANDN U6974 ( .B(B[34]), .A(n62), .Z(n6753) );
  XNOR U6975 ( .A(n6761), .B(n6975), .Z(n6754) );
  XNOR U6976 ( .A(n6760), .B(n6758), .Z(n6975) );
  AND U6977 ( .A(n6976), .B(n6977), .Z(n6758) );
  NANDN U6978 ( .A(n6978), .B(n6979), .Z(n6977) );
  OR U6979 ( .A(n6980), .B(n6981), .Z(n6979) );
  NAND U6980 ( .A(n6981), .B(n6980), .Z(n6976) );
  ANDN U6981 ( .B(B[35]), .A(n63), .Z(n6760) );
  XNOR U6982 ( .A(n6768), .B(n6982), .Z(n6761) );
  XNOR U6983 ( .A(n6767), .B(n6765), .Z(n6982) );
  AND U6984 ( .A(n6983), .B(n6984), .Z(n6765) );
  NANDN U6985 ( .A(n6985), .B(n6986), .Z(n6984) );
  NANDN U6986 ( .A(n6987), .B(n6988), .Z(n6986) );
  NANDN U6987 ( .A(n6988), .B(n6987), .Z(n6983) );
  ANDN U6988 ( .B(B[36]), .A(n64), .Z(n6767) );
  XNOR U6989 ( .A(n6775), .B(n6989), .Z(n6768) );
  XNOR U6990 ( .A(n6774), .B(n6772), .Z(n6989) );
  AND U6991 ( .A(n6990), .B(n6991), .Z(n6772) );
  NANDN U6992 ( .A(n6992), .B(n6993), .Z(n6991) );
  OR U6993 ( .A(n6994), .B(n6995), .Z(n6993) );
  NAND U6994 ( .A(n6995), .B(n6994), .Z(n6990) );
  ANDN U6995 ( .B(B[37]), .A(n65), .Z(n6774) );
  XNOR U6996 ( .A(n6782), .B(n6996), .Z(n6775) );
  XNOR U6997 ( .A(n6781), .B(n6779), .Z(n6996) );
  AND U6998 ( .A(n6997), .B(n6998), .Z(n6779) );
  NANDN U6999 ( .A(n6999), .B(n7000), .Z(n6998) );
  NANDN U7000 ( .A(n7001), .B(n7002), .Z(n7000) );
  NANDN U7001 ( .A(n7002), .B(n7001), .Z(n6997) );
  ANDN U7002 ( .B(B[38]), .A(n66), .Z(n6781) );
  XNOR U7003 ( .A(n6789), .B(n7003), .Z(n6782) );
  XNOR U7004 ( .A(n6788), .B(n6786), .Z(n7003) );
  AND U7005 ( .A(n7004), .B(n7005), .Z(n6786) );
  NANDN U7006 ( .A(n7006), .B(n7007), .Z(n7005) );
  OR U7007 ( .A(n7008), .B(n7009), .Z(n7007) );
  NAND U7008 ( .A(n7009), .B(n7008), .Z(n7004) );
  ANDN U7009 ( .B(B[39]), .A(n67), .Z(n6788) );
  XNOR U7010 ( .A(n6796), .B(n7010), .Z(n6789) );
  XNOR U7011 ( .A(n6795), .B(n6793), .Z(n7010) );
  AND U7012 ( .A(n7011), .B(n7012), .Z(n6793) );
  NANDN U7013 ( .A(n7013), .B(n7014), .Z(n7012) );
  NANDN U7014 ( .A(n7015), .B(n7016), .Z(n7014) );
  NANDN U7015 ( .A(n7016), .B(n7015), .Z(n7011) );
  ANDN U7016 ( .B(B[40]), .A(n68), .Z(n6795) );
  XNOR U7017 ( .A(n6803), .B(n7017), .Z(n6796) );
  XNOR U7018 ( .A(n6802), .B(n6800), .Z(n7017) );
  AND U7019 ( .A(n7018), .B(n7019), .Z(n6800) );
  NANDN U7020 ( .A(n7020), .B(n7021), .Z(n7019) );
  OR U7021 ( .A(n7022), .B(n7023), .Z(n7021) );
  NAND U7022 ( .A(n7023), .B(n7022), .Z(n7018) );
  ANDN U7023 ( .B(B[41]), .A(n69), .Z(n6802) );
  XNOR U7024 ( .A(n6810), .B(n7024), .Z(n6803) );
  XNOR U7025 ( .A(n6809), .B(n6807), .Z(n7024) );
  AND U7026 ( .A(n7025), .B(n7026), .Z(n6807) );
  NANDN U7027 ( .A(n7027), .B(n7028), .Z(n7026) );
  NANDN U7028 ( .A(n7029), .B(n7030), .Z(n7028) );
  NANDN U7029 ( .A(n7030), .B(n7029), .Z(n7025) );
  ANDN U7030 ( .B(B[42]), .A(n70), .Z(n6809) );
  XNOR U7031 ( .A(n6817), .B(n7031), .Z(n6810) );
  XNOR U7032 ( .A(n6816), .B(n6814), .Z(n7031) );
  AND U7033 ( .A(n7032), .B(n7033), .Z(n6814) );
  NANDN U7034 ( .A(n7034), .B(n7035), .Z(n7033) );
  OR U7035 ( .A(n7036), .B(n7037), .Z(n7035) );
  NAND U7036 ( .A(n7037), .B(n7036), .Z(n7032) );
  ANDN U7037 ( .B(B[43]), .A(n71), .Z(n6816) );
  XNOR U7038 ( .A(n6824), .B(n7038), .Z(n6817) );
  XNOR U7039 ( .A(n6823), .B(n6821), .Z(n7038) );
  AND U7040 ( .A(n7039), .B(n7040), .Z(n6821) );
  NANDN U7041 ( .A(n7041), .B(n7042), .Z(n7040) );
  NANDN U7042 ( .A(n7043), .B(n7044), .Z(n7042) );
  NANDN U7043 ( .A(n7044), .B(n7043), .Z(n7039) );
  ANDN U7044 ( .B(B[44]), .A(n72), .Z(n6823) );
  XNOR U7045 ( .A(n6831), .B(n7045), .Z(n6824) );
  XNOR U7046 ( .A(n6830), .B(n6828), .Z(n7045) );
  AND U7047 ( .A(n7046), .B(n7047), .Z(n6828) );
  NANDN U7048 ( .A(n7048), .B(n7049), .Z(n7047) );
  OR U7049 ( .A(n7050), .B(n7051), .Z(n7049) );
  NAND U7050 ( .A(n7051), .B(n7050), .Z(n7046) );
  ANDN U7051 ( .B(B[45]), .A(n73), .Z(n6830) );
  XNOR U7052 ( .A(n6838), .B(n7052), .Z(n6831) );
  XNOR U7053 ( .A(n6837), .B(n6835), .Z(n7052) );
  AND U7054 ( .A(n7053), .B(n7054), .Z(n6835) );
  NANDN U7055 ( .A(n7055), .B(n7056), .Z(n7054) );
  NANDN U7056 ( .A(n7057), .B(n7058), .Z(n7056) );
  NANDN U7057 ( .A(n7058), .B(n7057), .Z(n7053) );
  ANDN U7058 ( .B(B[46]), .A(n74), .Z(n6837) );
  XNOR U7059 ( .A(n6845), .B(n7059), .Z(n6838) );
  XNOR U7060 ( .A(n6844), .B(n6842), .Z(n7059) );
  AND U7061 ( .A(n7060), .B(n7061), .Z(n6842) );
  NANDN U7062 ( .A(n7062), .B(n7063), .Z(n7061) );
  OR U7063 ( .A(n7064), .B(n7065), .Z(n7063) );
  NAND U7064 ( .A(n7065), .B(n7064), .Z(n7060) );
  ANDN U7065 ( .B(B[47]), .A(n75), .Z(n6844) );
  XNOR U7066 ( .A(n6852), .B(n7066), .Z(n6845) );
  XNOR U7067 ( .A(n6851), .B(n6849), .Z(n7066) );
  AND U7068 ( .A(n7067), .B(n7068), .Z(n6849) );
  NANDN U7069 ( .A(n7069), .B(n7070), .Z(n7068) );
  NANDN U7070 ( .A(n7071), .B(n7072), .Z(n7070) );
  NANDN U7071 ( .A(n7072), .B(n7071), .Z(n7067) );
  ANDN U7072 ( .B(B[48]), .A(n76), .Z(n6851) );
  XNOR U7073 ( .A(n6859), .B(n7073), .Z(n6852) );
  XNOR U7074 ( .A(n6858), .B(n6856), .Z(n7073) );
  AND U7075 ( .A(n7074), .B(n7075), .Z(n6856) );
  NANDN U7076 ( .A(n7076), .B(n7077), .Z(n7075) );
  OR U7077 ( .A(n7078), .B(n7079), .Z(n7077) );
  NAND U7078 ( .A(n7079), .B(n7078), .Z(n7074) );
  ANDN U7079 ( .B(B[49]), .A(n77), .Z(n6858) );
  XNOR U7080 ( .A(n6866), .B(n7080), .Z(n6859) );
  XNOR U7081 ( .A(n6865), .B(n6863), .Z(n7080) );
  AND U7082 ( .A(n7081), .B(n7082), .Z(n6863) );
  NANDN U7083 ( .A(n7083), .B(n7084), .Z(n7082) );
  NANDN U7084 ( .A(n7085), .B(n7086), .Z(n7084) );
  NANDN U7085 ( .A(n7086), .B(n7085), .Z(n7081) );
  ANDN U7086 ( .B(B[50]), .A(n78), .Z(n6865) );
  XNOR U7087 ( .A(n6873), .B(n7087), .Z(n6866) );
  XNOR U7088 ( .A(n6872), .B(n6870), .Z(n7087) );
  AND U7089 ( .A(n7088), .B(n7089), .Z(n6870) );
  NANDN U7090 ( .A(n7090), .B(n7091), .Z(n7089) );
  OR U7091 ( .A(n7092), .B(n7093), .Z(n7091) );
  NAND U7092 ( .A(n7093), .B(n7092), .Z(n7088) );
  ANDN U7093 ( .B(B[51]), .A(n79), .Z(n6872) );
  XNOR U7094 ( .A(n6880), .B(n7094), .Z(n6873) );
  XNOR U7095 ( .A(n6879), .B(n6877), .Z(n7094) );
  AND U7096 ( .A(n7095), .B(n7096), .Z(n6877) );
  NANDN U7097 ( .A(n7097), .B(n7098), .Z(n7096) );
  NANDN U7098 ( .A(n7099), .B(n7100), .Z(n7098) );
  NANDN U7099 ( .A(n7100), .B(n7099), .Z(n7095) );
  ANDN U7100 ( .B(B[52]), .A(n80), .Z(n6879) );
  XNOR U7101 ( .A(n6887), .B(n7101), .Z(n6880) );
  XNOR U7102 ( .A(n6886), .B(n6884), .Z(n7101) );
  AND U7103 ( .A(n7102), .B(n7103), .Z(n6884) );
  NANDN U7104 ( .A(n7104), .B(n7105), .Z(n7103) );
  OR U7105 ( .A(n7106), .B(n7107), .Z(n7105) );
  NAND U7106 ( .A(n7107), .B(n7106), .Z(n7102) );
  ANDN U7107 ( .B(B[53]), .A(n81), .Z(n6886) );
  XNOR U7108 ( .A(n6894), .B(n7108), .Z(n6887) );
  XNOR U7109 ( .A(n6893), .B(n6891), .Z(n7108) );
  AND U7110 ( .A(n7109), .B(n7110), .Z(n6891) );
  NANDN U7111 ( .A(n7111), .B(n7112), .Z(n7110) );
  NAND U7112 ( .A(n7113), .B(n7114), .Z(n7112) );
  ANDN U7113 ( .B(B[54]), .A(n82), .Z(n6893) );
  XOR U7114 ( .A(n6900), .B(n7115), .Z(n6894) );
  XNOR U7115 ( .A(n6898), .B(n6901), .Z(n7115) );
  NAND U7116 ( .A(A[2]), .B(B[55]), .Z(n6901) );
  NANDN U7117 ( .A(n7116), .B(n7117), .Z(n6898) );
  AND U7118 ( .A(A[0]), .B(B[56]), .Z(n7117) );
  XNOR U7119 ( .A(n6903), .B(n7118), .Z(n6900) );
  NAND U7120 ( .A(A[0]), .B(B[57]), .Z(n7118) );
  NAND U7121 ( .A(B[56]), .B(A[1]), .Z(n6903) );
  NAND U7122 ( .A(n7119), .B(n7120), .Z(n173) );
  NANDN U7123 ( .A(n7121), .B(n7122), .Z(n7120) );
  OR U7124 ( .A(n7123), .B(n7124), .Z(n7122) );
  NAND U7125 ( .A(n7124), .B(n7123), .Z(n7119) );
  XOR U7126 ( .A(n175), .B(n174), .Z(\A1[54] ) );
  XOR U7127 ( .A(n7124), .B(n7125), .Z(n174) );
  XNOR U7128 ( .A(n7123), .B(n7121), .Z(n7125) );
  AND U7129 ( .A(n7126), .B(n7127), .Z(n7121) );
  NANDN U7130 ( .A(n7128), .B(n7129), .Z(n7127) );
  NANDN U7131 ( .A(n7130), .B(n7131), .Z(n7129) );
  NANDN U7132 ( .A(n7131), .B(n7130), .Z(n7126) );
  ANDN U7133 ( .B(B[25]), .A(n54), .Z(n7123) );
  XNOR U7134 ( .A(n6918), .B(n7132), .Z(n7124) );
  XNOR U7135 ( .A(n6917), .B(n6915), .Z(n7132) );
  AND U7136 ( .A(n7133), .B(n7134), .Z(n6915) );
  NANDN U7137 ( .A(n7135), .B(n7136), .Z(n7134) );
  OR U7138 ( .A(n7137), .B(n7138), .Z(n7136) );
  NAND U7139 ( .A(n7138), .B(n7137), .Z(n7133) );
  ANDN U7140 ( .B(B[26]), .A(n55), .Z(n6917) );
  XNOR U7141 ( .A(n6925), .B(n7139), .Z(n6918) );
  XNOR U7142 ( .A(n6924), .B(n6922), .Z(n7139) );
  AND U7143 ( .A(n7140), .B(n7141), .Z(n6922) );
  NANDN U7144 ( .A(n7142), .B(n7143), .Z(n7141) );
  NANDN U7145 ( .A(n7144), .B(n7145), .Z(n7143) );
  NANDN U7146 ( .A(n7145), .B(n7144), .Z(n7140) );
  ANDN U7147 ( .B(B[27]), .A(n56), .Z(n6924) );
  XNOR U7148 ( .A(n6932), .B(n7146), .Z(n6925) );
  XNOR U7149 ( .A(n6931), .B(n6929), .Z(n7146) );
  AND U7150 ( .A(n7147), .B(n7148), .Z(n6929) );
  NANDN U7151 ( .A(n7149), .B(n7150), .Z(n7148) );
  OR U7152 ( .A(n7151), .B(n7152), .Z(n7150) );
  NAND U7153 ( .A(n7152), .B(n7151), .Z(n7147) );
  ANDN U7154 ( .B(B[28]), .A(n57), .Z(n6931) );
  XNOR U7155 ( .A(n6939), .B(n7153), .Z(n6932) );
  XNOR U7156 ( .A(n6938), .B(n6936), .Z(n7153) );
  AND U7157 ( .A(n7154), .B(n7155), .Z(n6936) );
  NANDN U7158 ( .A(n7156), .B(n7157), .Z(n7155) );
  NANDN U7159 ( .A(n7158), .B(n7159), .Z(n7157) );
  NANDN U7160 ( .A(n7159), .B(n7158), .Z(n7154) );
  ANDN U7161 ( .B(B[29]), .A(n58), .Z(n6938) );
  XNOR U7162 ( .A(n6946), .B(n7160), .Z(n6939) );
  XNOR U7163 ( .A(n6945), .B(n6943), .Z(n7160) );
  AND U7164 ( .A(n7161), .B(n7162), .Z(n6943) );
  NANDN U7165 ( .A(n7163), .B(n7164), .Z(n7162) );
  OR U7166 ( .A(n7165), .B(n7166), .Z(n7164) );
  NAND U7167 ( .A(n7166), .B(n7165), .Z(n7161) );
  ANDN U7168 ( .B(B[30]), .A(n59), .Z(n6945) );
  XNOR U7169 ( .A(n6953), .B(n7167), .Z(n6946) );
  XNOR U7170 ( .A(n6952), .B(n6950), .Z(n7167) );
  AND U7171 ( .A(n7168), .B(n7169), .Z(n6950) );
  NANDN U7172 ( .A(n7170), .B(n7171), .Z(n7169) );
  NANDN U7173 ( .A(n7172), .B(n7173), .Z(n7171) );
  NANDN U7174 ( .A(n7173), .B(n7172), .Z(n7168) );
  ANDN U7175 ( .B(B[31]), .A(n60), .Z(n6952) );
  XNOR U7176 ( .A(n6960), .B(n7174), .Z(n6953) );
  XNOR U7177 ( .A(n6959), .B(n6957), .Z(n7174) );
  AND U7178 ( .A(n7175), .B(n7176), .Z(n6957) );
  NANDN U7179 ( .A(n7177), .B(n7178), .Z(n7176) );
  OR U7180 ( .A(n7179), .B(n7180), .Z(n7178) );
  NAND U7181 ( .A(n7180), .B(n7179), .Z(n7175) );
  ANDN U7182 ( .B(B[32]), .A(n61), .Z(n6959) );
  XNOR U7183 ( .A(n6967), .B(n7181), .Z(n6960) );
  XNOR U7184 ( .A(n6966), .B(n6964), .Z(n7181) );
  AND U7185 ( .A(n7182), .B(n7183), .Z(n6964) );
  NANDN U7186 ( .A(n7184), .B(n7185), .Z(n7183) );
  NANDN U7187 ( .A(n7186), .B(n7187), .Z(n7185) );
  NANDN U7188 ( .A(n7187), .B(n7186), .Z(n7182) );
  ANDN U7189 ( .B(B[33]), .A(n62), .Z(n6966) );
  XNOR U7190 ( .A(n6974), .B(n7188), .Z(n6967) );
  XNOR U7191 ( .A(n6973), .B(n6971), .Z(n7188) );
  AND U7192 ( .A(n7189), .B(n7190), .Z(n6971) );
  NANDN U7193 ( .A(n7191), .B(n7192), .Z(n7190) );
  OR U7194 ( .A(n7193), .B(n7194), .Z(n7192) );
  NAND U7195 ( .A(n7194), .B(n7193), .Z(n7189) );
  ANDN U7196 ( .B(B[34]), .A(n63), .Z(n6973) );
  XNOR U7197 ( .A(n6981), .B(n7195), .Z(n6974) );
  XNOR U7198 ( .A(n6980), .B(n6978), .Z(n7195) );
  AND U7199 ( .A(n7196), .B(n7197), .Z(n6978) );
  NANDN U7200 ( .A(n7198), .B(n7199), .Z(n7197) );
  NANDN U7201 ( .A(n7200), .B(n7201), .Z(n7199) );
  NANDN U7202 ( .A(n7201), .B(n7200), .Z(n7196) );
  ANDN U7203 ( .B(B[35]), .A(n64), .Z(n6980) );
  XNOR U7204 ( .A(n6988), .B(n7202), .Z(n6981) );
  XNOR U7205 ( .A(n6987), .B(n6985), .Z(n7202) );
  AND U7206 ( .A(n7203), .B(n7204), .Z(n6985) );
  NANDN U7207 ( .A(n7205), .B(n7206), .Z(n7204) );
  OR U7208 ( .A(n7207), .B(n7208), .Z(n7206) );
  NAND U7209 ( .A(n7208), .B(n7207), .Z(n7203) );
  ANDN U7210 ( .B(B[36]), .A(n65), .Z(n6987) );
  XNOR U7211 ( .A(n6995), .B(n7209), .Z(n6988) );
  XNOR U7212 ( .A(n6994), .B(n6992), .Z(n7209) );
  AND U7213 ( .A(n7210), .B(n7211), .Z(n6992) );
  NANDN U7214 ( .A(n7212), .B(n7213), .Z(n7211) );
  NANDN U7215 ( .A(n7214), .B(n7215), .Z(n7213) );
  NANDN U7216 ( .A(n7215), .B(n7214), .Z(n7210) );
  ANDN U7217 ( .B(B[37]), .A(n66), .Z(n6994) );
  XNOR U7218 ( .A(n7002), .B(n7216), .Z(n6995) );
  XNOR U7219 ( .A(n7001), .B(n6999), .Z(n7216) );
  AND U7220 ( .A(n7217), .B(n7218), .Z(n6999) );
  NANDN U7221 ( .A(n7219), .B(n7220), .Z(n7218) );
  OR U7222 ( .A(n7221), .B(n7222), .Z(n7220) );
  NAND U7223 ( .A(n7222), .B(n7221), .Z(n7217) );
  ANDN U7224 ( .B(B[38]), .A(n67), .Z(n7001) );
  XNOR U7225 ( .A(n7009), .B(n7223), .Z(n7002) );
  XNOR U7226 ( .A(n7008), .B(n7006), .Z(n7223) );
  AND U7227 ( .A(n7224), .B(n7225), .Z(n7006) );
  NANDN U7228 ( .A(n7226), .B(n7227), .Z(n7225) );
  NANDN U7229 ( .A(n7228), .B(n7229), .Z(n7227) );
  NANDN U7230 ( .A(n7229), .B(n7228), .Z(n7224) );
  ANDN U7231 ( .B(B[39]), .A(n68), .Z(n7008) );
  XNOR U7232 ( .A(n7016), .B(n7230), .Z(n7009) );
  XNOR U7233 ( .A(n7015), .B(n7013), .Z(n7230) );
  AND U7234 ( .A(n7231), .B(n7232), .Z(n7013) );
  NANDN U7235 ( .A(n7233), .B(n7234), .Z(n7232) );
  OR U7236 ( .A(n7235), .B(n7236), .Z(n7234) );
  NAND U7237 ( .A(n7236), .B(n7235), .Z(n7231) );
  ANDN U7238 ( .B(B[40]), .A(n69), .Z(n7015) );
  XNOR U7239 ( .A(n7023), .B(n7237), .Z(n7016) );
  XNOR U7240 ( .A(n7022), .B(n7020), .Z(n7237) );
  AND U7241 ( .A(n7238), .B(n7239), .Z(n7020) );
  NANDN U7242 ( .A(n7240), .B(n7241), .Z(n7239) );
  NANDN U7243 ( .A(n7242), .B(n7243), .Z(n7241) );
  NANDN U7244 ( .A(n7243), .B(n7242), .Z(n7238) );
  ANDN U7245 ( .B(B[41]), .A(n70), .Z(n7022) );
  XNOR U7246 ( .A(n7030), .B(n7244), .Z(n7023) );
  XNOR U7247 ( .A(n7029), .B(n7027), .Z(n7244) );
  AND U7248 ( .A(n7245), .B(n7246), .Z(n7027) );
  NANDN U7249 ( .A(n7247), .B(n7248), .Z(n7246) );
  OR U7250 ( .A(n7249), .B(n7250), .Z(n7248) );
  NAND U7251 ( .A(n7250), .B(n7249), .Z(n7245) );
  ANDN U7252 ( .B(B[42]), .A(n71), .Z(n7029) );
  XNOR U7253 ( .A(n7037), .B(n7251), .Z(n7030) );
  XNOR U7254 ( .A(n7036), .B(n7034), .Z(n7251) );
  AND U7255 ( .A(n7252), .B(n7253), .Z(n7034) );
  NANDN U7256 ( .A(n7254), .B(n7255), .Z(n7253) );
  NANDN U7257 ( .A(n7256), .B(n7257), .Z(n7255) );
  NANDN U7258 ( .A(n7257), .B(n7256), .Z(n7252) );
  ANDN U7259 ( .B(B[43]), .A(n72), .Z(n7036) );
  XNOR U7260 ( .A(n7044), .B(n7258), .Z(n7037) );
  XNOR U7261 ( .A(n7043), .B(n7041), .Z(n7258) );
  AND U7262 ( .A(n7259), .B(n7260), .Z(n7041) );
  NANDN U7263 ( .A(n7261), .B(n7262), .Z(n7260) );
  OR U7264 ( .A(n7263), .B(n7264), .Z(n7262) );
  NAND U7265 ( .A(n7264), .B(n7263), .Z(n7259) );
  ANDN U7266 ( .B(B[44]), .A(n73), .Z(n7043) );
  XNOR U7267 ( .A(n7051), .B(n7265), .Z(n7044) );
  XNOR U7268 ( .A(n7050), .B(n7048), .Z(n7265) );
  AND U7269 ( .A(n7266), .B(n7267), .Z(n7048) );
  NANDN U7270 ( .A(n7268), .B(n7269), .Z(n7267) );
  NANDN U7271 ( .A(n7270), .B(n7271), .Z(n7269) );
  NANDN U7272 ( .A(n7271), .B(n7270), .Z(n7266) );
  ANDN U7273 ( .B(B[45]), .A(n74), .Z(n7050) );
  XNOR U7274 ( .A(n7058), .B(n7272), .Z(n7051) );
  XNOR U7275 ( .A(n7057), .B(n7055), .Z(n7272) );
  AND U7276 ( .A(n7273), .B(n7274), .Z(n7055) );
  NANDN U7277 ( .A(n7275), .B(n7276), .Z(n7274) );
  OR U7278 ( .A(n7277), .B(n7278), .Z(n7276) );
  NAND U7279 ( .A(n7278), .B(n7277), .Z(n7273) );
  ANDN U7280 ( .B(B[46]), .A(n75), .Z(n7057) );
  XNOR U7281 ( .A(n7065), .B(n7279), .Z(n7058) );
  XNOR U7282 ( .A(n7064), .B(n7062), .Z(n7279) );
  AND U7283 ( .A(n7280), .B(n7281), .Z(n7062) );
  NANDN U7284 ( .A(n7282), .B(n7283), .Z(n7281) );
  NANDN U7285 ( .A(n7284), .B(n7285), .Z(n7283) );
  NANDN U7286 ( .A(n7285), .B(n7284), .Z(n7280) );
  ANDN U7287 ( .B(B[47]), .A(n76), .Z(n7064) );
  XNOR U7288 ( .A(n7072), .B(n7286), .Z(n7065) );
  XNOR U7289 ( .A(n7071), .B(n7069), .Z(n7286) );
  AND U7290 ( .A(n7287), .B(n7288), .Z(n7069) );
  NANDN U7291 ( .A(n7289), .B(n7290), .Z(n7288) );
  OR U7292 ( .A(n7291), .B(n7292), .Z(n7290) );
  NAND U7293 ( .A(n7292), .B(n7291), .Z(n7287) );
  ANDN U7294 ( .B(B[48]), .A(n77), .Z(n7071) );
  XNOR U7295 ( .A(n7079), .B(n7293), .Z(n7072) );
  XNOR U7296 ( .A(n7078), .B(n7076), .Z(n7293) );
  AND U7297 ( .A(n7294), .B(n7295), .Z(n7076) );
  NANDN U7298 ( .A(n7296), .B(n7297), .Z(n7295) );
  NANDN U7299 ( .A(n7298), .B(n7299), .Z(n7297) );
  NANDN U7300 ( .A(n7299), .B(n7298), .Z(n7294) );
  ANDN U7301 ( .B(B[49]), .A(n78), .Z(n7078) );
  XNOR U7302 ( .A(n7086), .B(n7300), .Z(n7079) );
  XNOR U7303 ( .A(n7085), .B(n7083), .Z(n7300) );
  AND U7304 ( .A(n7301), .B(n7302), .Z(n7083) );
  NANDN U7305 ( .A(n7303), .B(n7304), .Z(n7302) );
  OR U7306 ( .A(n7305), .B(n7306), .Z(n7304) );
  NAND U7307 ( .A(n7306), .B(n7305), .Z(n7301) );
  ANDN U7308 ( .B(B[50]), .A(n79), .Z(n7085) );
  XNOR U7309 ( .A(n7093), .B(n7307), .Z(n7086) );
  XNOR U7310 ( .A(n7092), .B(n7090), .Z(n7307) );
  AND U7311 ( .A(n7308), .B(n7309), .Z(n7090) );
  NANDN U7312 ( .A(n7310), .B(n7311), .Z(n7309) );
  NANDN U7313 ( .A(n7312), .B(n7313), .Z(n7311) );
  NANDN U7314 ( .A(n7313), .B(n7312), .Z(n7308) );
  ANDN U7315 ( .B(B[51]), .A(n80), .Z(n7092) );
  XNOR U7316 ( .A(n7100), .B(n7314), .Z(n7093) );
  XNOR U7317 ( .A(n7099), .B(n7097), .Z(n7314) );
  AND U7318 ( .A(n7315), .B(n7316), .Z(n7097) );
  NANDN U7319 ( .A(n7317), .B(n7318), .Z(n7316) );
  OR U7320 ( .A(n7319), .B(n7320), .Z(n7318) );
  NAND U7321 ( .A(n7320), .B(n7319), .Z(n7315) );
  ANDN U7322 ( .B(B[52]), .A(n81), .Z(n7099) );
  XNOR U7323 ( .A(n7107), .B(n7321), .Z(n7100) );
  XNOR U7324 ( .A(n7106), .B(n7104), .Z(n7321) );
  AND U7325 ( .A(n7322), .B(n7323), .Z(n7104) );
  NANDN U7326 ( .A(n7324), .B(n7325), .Z(n7323) );
  NAND U7327 ( .A(n7326), .B(n7327), .Z(n7325) );
  ANDN U7328 ( .B(B[53]), .A(n82), .Z(n7106) );
  XOR U7329 ( .A(n7113), .B(n7328), .Z(n7107) );
  XNOR U7330 ( .A(n7111), .B(n7114), .Z(n7328) );
  NAND U7331 ( .A(A[2]), .B(B[54]), .Z(n7114) );
  NANDN U7332 ( .A(n7329), .B(n7330), .Z(n7111) );
  AND U7333 ( .A(A[0]), .B(B[55]), .Z(n7330) );
  XNOR U7334 ( .A(n7116), .B(n7331), .Z(n7113) );
  NAND U7335 ( .A(A[0]), .B(B[56]), .Z(n7331) );
  NAND U7336 ( .A(B[55]), .B(A[1]), .Z(n7116) );
  NAND U7337 ( .A(n7332), .B(n7333), .Z(n175) );
  NANDN U7338 ( .A(n7334), .B(n7335), .Z(n7333) );
  OR U7339 ( .A(n7336), .B(n7337), .Z(n7335) );
  NAND U7340 ( .A(n7337), .B(n7336), .Z(n7332) );
  XOR U7341 ( .A(n177), .B(n176), .Z(\A1[53] ) );
  XOR U7342 ( .A(n7337), .B(n7338), .Z(n176) );
  XNOR U7343 ( .A(n7336), .B(n7334), .Z(n7338) );
  AND U7344 ( .A(n7339), .B(n7340), .Z(n7334) );
  NANDN U7345 ( .A(n7341), .B(n7342), .Z(n7340) );
  NANDN U7346 ( .A(n7343), .B(n7344), .Z(n7342) );
  NANDN U7347 ( .A(n7344), .B(n7343), .Z(n7339) );
  ANDN U7348 ( .B(B[24]), .A(n54), .Z(n7336) );
  XNOR U7349 ( .A(n7131), .B(n7345), .Z(n7337) );
  XNOR U7350 ( .A(n7130), .B(n7128), .Z(n7345) );
  AND U7351 ( .A(n7346), .B(n7347), .Z(n7128) );
  NANDN U7352 ( .A(n7348), .B(n7349), .Z(n7347) );
  OR U7353 ( .A(n7350), .B(n7351), .Z(n7349) );
  NAND U7354 ( .A(n7351), .B(n7350), .Z(n7346) );
  ANDN U7355 ( .B(B[25]), .A(n55), .Z(n7130) );
  XNOR U7356 ( .A(n7138), .B(n7352), .Z(n7131) );
  XNOR U7357 ( .A(n7137), .B(n7135), .Z(n7352) );
  AND U7358 ( .A(n7353), .B(n7354), .Z(n7135) );
  NANDN U7359 ( .A(n7355), .B(n7356), .Z(n7354) );
  NANDN U7360 ( .A(n7357), .B(n7358), .Z(n7356) );
  NANDN U7361 ( .A(n7358), .B(n7357), .Z(n7353) );
  ANDN U7362 ( .B(B[26]), .A(n56), .Z(n7137) );
  XNOR U7363 ( .A(n7145), .B(n7359), .Z(n7138) );
  XNOR U7364 ( .A(n7144), .B(n7142), .Z(n7359) );
  AND U7365 ( .A(n7360), .B(n7361), .Z(n7142) );
  NANDN U7366 ( .A(n7362), .B(n7363), .Z(n7361) );
  OR U7367 ( .A(n7364), .B(n7365), .Z(n7363) );
  NAND U7368 ( .A(n7365), .B(n7364), .Z(n7360) );
  ANDN U7369 ( .B(B[27]), .A(n57), .Z(n7144) );
  XNOR U7370 ( .A(n7152), .B(n7366), .Z(n7145) );
  XNOR U7371 ( .A(n7151), .B(n7149), .Z(n7366) );
  AND U7372 ( .A(n7367), .B(n7368), .Z(n7149) );
  NANDN U7373 ( .A(n7369), .B(n7370), .Z(n7368) );
  NANDN U7374 ( .A(n7371), .B(n7372), .Z(n7370) );
  NANDN U7375 ( .A(n7372), .B(n7371), .Z(n7367) );
  ANDN U7376 ( .B(B[28]), .A(n58), .Z(n7151) );
  XNOR U7377 ( .A(n7159), .B(n7373), .Z(n7152) );
  XNOR U7378 ( .A(n7158), .B(n7156), .Z(n7373) );
  AND U7379 ( .A(n7374), .B(n7375), .Z(n7156) );
  NANDN U7380 ( .A(n7376), .B(n7377), .Z(n7375) );
  OR U7381 ( .A(n7378), .B(n7379), .Z(n7377) );
  NAND U7382 ( .A(n7379), .B(n7378), .Z(n7374) );
  ANDN U7383 ( .B(B[29]), .A(n59), .Z(n7158) );
  XNOR U7384 ( .A(n7166), .B(n7380), .Z(n7159) );
  XNOR U7385 ( .A(n7165), .B(n7163), .Z(n7380) );
  AND U7386 ( .A(n7381), .B(n7382), .Z(n7163) );
  NANDN U7387 ( .A(n7383), .B(n7384), .Z(n7382) );
  NANDN U7388 ( .A(n7385), .B(n7386), .Z(n7384) );
  NANDN U7389 ( .A(n7386), .B(n7385), .Z(n7381) );
  ANDN U7390 ( .B(B[30]), .A(n60), .Z(n7165) );
  XNOR U7391 ( .A(n7173), .B(n7387), .Z(n7166) );
  XNOR U7392 ( .A(n7172), .B(n7170), .Z(n7387) );
  AND U7393 ( .A(n7388), .B(n7389), .Z(n7170) );
  NANDN U7394 ( .A(n7390), .B(n7391), .Z(n7389) );
  OR U7395 ( .A(n7392), .B(n7393), .Z(n7391) );
  NAND U7396 ( .A(n7393), .B(n7392), .Z(n7388) );
  ANDN U7397 ( .B(B[31]), .A(n61), .Z(n7172) );
  XNOR U7398 ( .A(n7180), .B(n7394), .Z(n7173) );
  XNOR U7399 ( .A(n7179), .B(n7177), .Z(n7394) );
  AND U7400 ( .A(n7395), .B(n7396), .Z(n7177) );
  NANDN U7401 ( .A(n7397), .B(n7398), .Z(n7396) );
  NANDN U7402 ( .A(n7399), .B(n7400), .Z(n7398) );
  NANDN U7403 ( .A(n7400), .B(n7399), .Z(n7395) );
  ANDN U7404 ( .B(B[32]), .A(n62), .Z(n7179) );
  XNOR U7405 ( .A(n7187), .B(n7401), .Z(n7180) );
  XNOR U7406 ( .A(n7186), .B(n7184), .Z(n7401) );
  AND U7407 ( .A(n7402), .B(n7403), .Z(n7184) );
  NANDN U7408 ( .A(n7404), .B(n7405), .Z(n7403) );
  OR U7409 ( .A(n7406), .B(n7407), .Z(n7405) );
  NAND U7410 ( .A(n7407), .B(n7406), .Z(n7402) );
  ANDN U7411 ( .B(B[33]), .A(n63), .Z(n7186) );
  XNOR U7412 ( .A(n7194), .B(n7408), .Z(n7187) );
  XNOR U7413 ( .A(n7193), .B(n7191), .Z(n7408) );
  AND U7414 ( .A(n7409), .B(n7410), .Z(n7191) );
  NANDN U7415 ( .A(n7411), .B(n7412), .Z(n7410) );
  NANDN U7416 ( .A(n7413), .B(n7414), .Z(n7412) );
  NANDN U7417 ( .A(n7414), .B(n7413), .Z(n7409) );
  ANDN U7418 ( .B(B[34]), .A(n64), .Z(n7193) );
  XNOR U7419 ( .A(n7201), .B(n7415), .Z(n7194) );
  XNOR U7420 ( .A(n7200), .B(n7198), .Z(n7415) );
  AND U7421 ( .A(n7416), .B(n7417), .Z(n7198) );
  NANDN U7422 ( .A(n7418), .B(n7419), .Z(n7417) );
  OR U7423 ( .A(n7420), .B(n7421), .Z(n7419) );
  NAND U7424 ( .A(n7421), .B(n7420), .Z(n7416) );
  ANDN U7425 ( .B(B[35]), .A(n65), .Z(n7200) );
  XNOR U7426 ( .A(n7208), .B(n7422), .Z(n7201) );
  XNOR U7427 ( .A(n7207), .B(n7205), .Z(n7422) );
  AND U7428 ( .A(n7423), .B(n7424), .Z(n7205) );
  NANDN U7429 ( .A(n7425), .B(n7426), .Z(n7424) );
  NANDN U7430 ( .A(n7427), .B(n7428), .Z(n7426) );
  NANDN U7431 ( .A(n7428), .B(n7427), .Z(n7423) );
  ANDN U7432 ( .B(B[36]), .A(n66), .Z(n7207) );
  XNOR U7433 ( .A(n7215), .B(n7429), .Z(n7208) );
  XNOR U7434 ( .A(n7214), .B(n7212), .Z(n7429) );
  AND U7435 ( .A(n7430), .B(n7431), .Z(n7212) );
  NANDN U7436 ( .A(n7432), .B(n7433), .Z(n7431) );
  OR U7437 ( .A(n7434), .B(n7435), .Z(n7433) );
  NAND U7438 ( .A(n7435), .B(n7434), .Z(n7430) );
  ANDN U7439 ( .B(B[37]), .A(n67), .Z(n7214) );
  XNOR U7440 ( .A(n7222), .B(n7436), .Z(n7215) );
  XNOR U7441 ( .A(n7221), .B(n7219), .Z(n7436) );
  AND U7442 ( .A(n7437), .B(n7438), .Z(n7219) );
  NANDN U7443 ( .A(n7439), .B(n7440), .Z(n7438) );
  NANDN U7444 ( .A(n7441), .B(n7442), .Z(n7440) );
  NANDN U7445 ( .A(n7442), .B(n7441), .Z(n7437) );
  ANDN U7446 ( .B(B[38]), .A(n68), .Z(n7221) );
  XNOR U7447 ( .A(n7229), .B(n7443), .Z(n7222) );
  XNOR U7448 ( .A(n7228), .B(n7226), .Z(n7443) );
  AND U7449 ( .A(n7444), .B(n7445), .Z(n7226) );
  NANDN U7450 ( .A(n7446), .B(n7447), .Z(n7445) );
  OR U7451 ( .A(n7448), .B(n7449), .Z(n7447) );
  NAND U7452 ( .A(n7449), .B(n7448), .Z(n7444) );
  ANDN U7453 ( .B(B[39]), .A(n69), .Z(n7228) );
  XNOR U7454 ( .A(n7236), .B(n7450), .Z(n7229) );
  XNOR U7455 ( .A(n7235), .B(n7233), .Z(n7450) );
  AND U7456 ( .A(n7451), .B(n7452), .Z(n7233) );
  NANDN U7457 ( .A(n7453), .B(n7454), .Z(n7452) );
  NANDN U7458 ( .A(n7455), .B(n7456), .Z(n7454) );
  NANDN U7459 ( .A(n7456), .B(n7455), .Z(n7451) );
  ANDN U7460 ( .B(B[40]), .A(n70), .Z(n7235) );
  XNOR U7461 ( .A(n7243), .B(n7457), .Z(n7236) );
  XNOR U7462 ( .A(n7242), .B(n7240), .Z(n7457) );
  AND U7463 ( .A(n7458), .B(n7459), .Z(n7240) );
  NANDN U7464 ( .A(n7460), .B(n7461), .Z(n7459) );
  OR U7465 ( .A(n7462), .B(n7463), .Z(n7461) );
  NAND U7466 ( .A(n7463), .B(n7462), .Z(n7458) );
  ANDN U7467 ( .B(B[41]), .A(n71), .Z(n7242) );
  XNOR U7468 ( .A(n7250), .B(n7464), .Z(n7243) );
  XNOR U7469 ( .A(n7249), .B(n7247), .Z(n7464) );
  AND U7470 ( .A(n7465), .B(n7466), .Z(n7247) );
  NANDN U7471 ( .A(n7467), .B(n7468), .Z(n7466) );
  NANDN U7472 ( .A(n7469), .B(n7470), .Z(n7468) );
  NANDN U7473 ( .A(n7470), .B(n7469), .Z(n7465) );
  ANDN U7474 ( .B(B[42]), .A(n72), .Z(n7249) );
  XNOR U7475 ( .A(n7257), .B(n7471), .Z(n7250) );
  XNOR U7476 ( .A(n7256), .B(n7254), .Z(n7471) );
  AND U7477 ( .A(n7472), .B(n7473), .Z(n7254) );
  NANDN U7478 ( .A(n7474), .B(n7475), .Z(n7473) );
  OR U7479 ( .A(n7476), .B(n7477), .Z(n7475) );
  NAND U7480 ( .A(n7477), .B(n7476), .Z(n7472) );
  ANDN U7481 ( .B(B[43]), .A(n73), .Z(n7256) );
  XNOR U7482 ( .A(n7264), .B(n7478), .Z(n7257) );
  XNOR U7483 ( .A(n7263), .B(n7261), .Z(n7478) );
  AND U7484 ( .A(n7479), .B(n7480), .Z(n7261) );
  NANDN U7485 ( .A(n7481), .B(n7482), .Z(n7480) );
  NANDN U7486 ( .A(n7483), .B(n7484), .Z(n7482) );
  NANDN U7487 ( .A(n7484), .B(n7483), .Z(n7479) );
  ANDN U7488 ( .B(B[44]), .A(n74), .Z(n7263) );
  XNOR U7489 ( .A(n7271), .B(n7485), .Z(n7264) );
  XNOR U7490 ( .A(n7270), .B(n7268), .Z(n7485) );
  AND U7491 ( .A(n7486), .B(n7487), .Z(n7268) );
  NANDN U7492 ( .A(n7488), .B(n7489), .Z(n7487) );
  OR U7493 ( .A(n7490), .B(n7491), .Z(n7489) );
  NAND U7494 ( .A(n7491), .B(n7490), .Z(n7486) );
  ANDN U7495 ( .B(B[45]), .A(n75), .Z(n7270) );
  XNOR U7496 ( .A(n7278), .B(n7492), .Z(n7271) );
  XNOR U7497 ( .A(n7277), .B(n7275), .Z(n7492) );
  AND U7498 ( .A(n7493), .B(n7494), .Z(n7275) );
  NANDN U7499 ( .A(n7495), .B(n7496), .Z(n7494) );
  NANDN U7500 ( .A(n7497), .B(n7498), .Z(n7496) );
  NANDN U7501 ( .A(n7498), .B(n7497), .Z(n7493) );
  ANDN U7502 ( .B(B[46]), .A(n76), .Z(n7277) );
  XNOR U7503 ( .A(n7285), .B(n7499), .Z(n7278) );
  XNOR U7504 ( .A(n7284), .B(n7282), .Z(n7499) );
  AND U7505 ( .A(n7500), .B(n7501), .Z(n7282) );
  NANDN U7506 ( .A(n7502), .B(n7503), .Z(n7501) );
  OR U7507 ( .A(n7504), .B(n7505), .Z(n7503) );
  NAND U7508 ( .A(n7505), .B(n7504), .Z(n7500) );
  ANDN U7509 ( .B(B[47]), .A(n77), .Z(n7284) );
  XNOR U7510 ( .A(n7292), .B(n7506), .Z(n7285) );
  XNOR U7511 ( .A(n7291), .B(n7289), .Z(n7506) );
  AND U7512 ( .A(n7507), .B(n7508), .Z(n7289) );
  NANDN U7513 ( .A(n7509), .B(n7510), .Z(n7508) );
  NANDN U7514 ( .A(n7511), .B(n7512), .Z(n7510) );
  NANDN U7515 ( .A(n7512), .B(n7511), .Z(n7507) );
  ANDN U7516 ( .B(B[48]), .A(n78), .Z(n7291) );
  XNOR U7517 ( .A(n7299), .B(n7513), .Z(n7292) );
  XNOR U7518 ( .A(n7298), .B(n7296), .Z(n7513) );
  AND U7519 ( .A(n7514), .B(n7515), .Z(n7296) );
  NANDN U7520 ( .A(n7516), .B(n7517), .Z(n7515) );
  OR U7521 ( .A(n7518), .B(n7519), .Z(n7517) );
  NAND U7522 ( .A(n7519), .B(n7518), .Z(n7514) );
  ANDN U7523 ( .B(B[49]), .A(n79), .Z(n7298) );
  XNOR U7524 ( .A(n7306), .B(n7520), .Z(n7299) );
  XNOR U7525 ( .A(n7305), .B(n7303), .Z(n7520) );
  AND U7526 ( .A(n7521), .B(n7522), .Z(n7303) );
  NANDN U7527 ( .A(n7523), .B(n7524), .Z(n7522) );
  NANDN U7528 ( .A(n7525), .B(n7526), .Z(n7524) );
  NANDN U7529 ( .A(n7526), .B(n7525), .Z(n7521) );
  ANDN U7530 ( .B(B[50]), .A(n80), .Z(n7305) );
  XNOR U7531 ( .A(n7313), .B(n7527), .Z(n7306) );
  XNOR U7532 ( .A(n7312), .B(n7310), .Z(n7527) );
  AND U7533 ( .A(n7528), .B(n7529), .Z(n7310) );
  NANDN U7534 ( .A(n7530), .B(n7531), .Z(n7529) );
  OR U7535 ( .A(n7532), .B(n7533), .Z(n7531) );
  NAND U7536 ( .A(n7533), .B(n7532), .Z(n7528) );
  ANDN U7537 ( .B(B[51]), .A(n81), .Z(n7312) );
  XNOR U7538 ( .A(n7320), .B(n7534), .Z(n7313) );
  XNOR U7539 ( .A(n7319), .B(n7317), .Z(n7534) );
  AND U7540 ( .A(n7535), .B(n7536), .Z(n7317) );
  NANDN U7541 ( .A(n7537), .B(n7538), .Z(n7536) );
  NAND U7542 ( .A(n7539), .B(n7540), .Z(n7538) );
  ANDN U7543 ( .B(B[52]), .A(n82), .Z(n7319) );
  XOR U7544 ( .A(n7326), .B(n7541), .Z(n7320) );
  XNOR U7545 ( .A(n7324), .B(n7327), .Z(n7541) );
  NAND U7546 ( .A(A[2]), .B(B[53]), .Z(n7327) );
  NANDN U7547 ( .A(n7542), .B(n7543), .Z(n7324) );
  AND U7548 ( .A(A[0]), .B(B[54]), .Z(n7543) );
  XNOR U7549 ( .A(n7329), .B(n7544), .Z(n7326) );
  NAND U7550 ( .A(A[0]), .B(B[55]), .Z(n7544) );
  NAND U7551 ( .A(B[54]), .B(A[1]), .Z(n7329) );
  NAND U7552 ( .A(n7545), .B(n7546), .Z(n177) );
  NANDN U7553 ( .A(n7547), .B(n7548), .Z(n7546) );
  OR U7554 ( .A(n7549), .B(n7550), .Z(n7548) );
  NAND U7555 ( .A(n7550), .B(n7549), .Z(n7545) );
  XOR U7556 ( .A(n179), .B(n178), .Z(\A1[52] ) );
  XOR U7557 ( .A(n7550), .B(n7551), .Z(n178) );
  XNOR U7558 ( .A(n7549), .B(n7547), .Z(n7551) );
  AND U7559 ( .A(n7552), .B(n7553), .Z(n7547) );
  NANDN U7560 ( .A(n7554), .B(n7555), .Z(n7553) );
  NANDN U7561 ( .A(n7556), .B(n7557), .Z(n7555) );
  NANDN U7562 ( .A(n7557), .B(n7556), .Z(n7552) );
  ANDN U7563 ( .B(B[23]), .A(n54), .Z(n7549) );
  XNOR U7564 ( .A(n7344), .B(n7558), .Z(n7550) );
  XNOR U7565 ( .A(n7343), .B(n7341), .Z(n7558) );
  AND U7566 ( .A(n7559), .B(n7560), .Z(n7341) );
  NANDN U7567 ( .A(n7561), .B(n7562), .Z(n7560) );
  OR U7568 ( .A(n7563), .B(n7564), .Z(n7562) );
  NAND U7569 ( .A(n7564), .B(n7563), .Z(n7559) );
  ANDN U7570 ( .B(B[24]), .A(n55), .Z(n7343) );
  XNOR U7571 ( .A(n7351), .B(n7565), .Z(n7344) );
  XNOR U7572 ( .A(n7350), .B(n7348), .Z(n7565) );
  AND U7573 ( .A(n7566), .B(n7567), .Z(n7348) );
  NANDN U7574 ( .A(n7568), .B(n7569), .Z(n7567) );
  NANDN U7575 ( .A(n7570), .B(n7571), .Z(n7569) );
  NANDN U7576 ( .A(n7571), .B(n7570), .Z(n7566) );
  ANDN U7577 ( .B(B[25]), .A(n56), .Z(n7350) );
  XNOR U7578 ( .A(n7358), .B(n7572), .Z(n7351) );
  XNOR U7579 ( .A(n7357), .B(n7355), .Z(n7572) );
  AND U7580 ( .A(n7573), .B(n7574), .Z(n7355) );
  NANDN U7581 ( .A(n7575), .B(n7576), .Z(n7574) );
  OR U7582 ( .A(n7577), .B(n7578), .Z(n7576) );
  NAND U7583 ( .A(n7578), .B(n7577), .Z(n7573) );
  ANDN U7584 ( .B(B[26]), .A(n57), .Z(n7357) );
  XNOR U7585 ( .A(n7365), .B(n7579), .Z(n7358) );
  XNOR U7586 ( .A(n7364), .B(n7362), .Z(n7579) );
  AND U7587 ( .A(n7580), .B(n7581), .Z(n7362) );
  NANDN U7588 ( .A(n7582), .B(n7583), .Z(n7581) );
  NANDN U7589 ( .A(n7584), .B(n7585), .Z(n7583) );
  NANDN U7590 ( .A(n7585), .B(n7584), .Z(n7580) );
  ANDN U7591 ( .B(B[27]), .A(n58), .Z(n7364) );
  XNOR U7592 ( .A(n7372), .B(n7586), .Z(n7365) );
  XNOR U7593 ( .A(n7371), .B(n7369), .Z(n7586) );
  AND U7594 ( .A(n7587), .B(n7588), .Z(n7369) );
  NANDN U7595 ( .A(n7589), .B(n7590), .Z(n7588) );
  OR U7596 ( .A(n7591), .B(n7592), .Z(n7590) );
  NAND U7597 ( .A(n7592), .B(n7591), .Z(n7587) );
  ANDN U7598 ( .B(B[28]), .A(n59), .Z(n7371) );
  XNOR U7599 ( .A(n7379), .B(n7593), .Z(n7372) );
  XNOR U7600 ( .A(n7378), .B(n7376), .Z(n7593) );
  AND U7601 ( .A(n7594), .B(n7595), .Z(n7376) );
  NANDN U7602 ( .A(n7596), .B(n7597), .Z(n7595) );
  NANDN U7603 ( .A(n7598), .B(n7599), .Z(n7597) );
  NANDN U7604 ( .A(n7599), .B(n7598), .Z(n7594) );
  ANDN U7605 ( .B(B[29]), .A(n60), .Z(n7378) );
  XNOR U7606 ( .A(n7386), .B(n7600), .Z(n7379) );
  XNOR U7607 ( .A(n7385), .B(n7383), .Z(n7600) );
  AND U7608 ( .A(n7601), .B(n7602), .Z(n7383) );
  NANDN U7609 ( .A(n7603), .B(n7604), .Z(n7602) );
  OR U7610 ( .A(n7605), .B(n7606), .Z(n7604) );
  NAND U7611 ( .A(n7606), .B(n7605), .Z(n7601) );
  ANDN U7612 ( .B(B[30]), .A(n61), .Z(n7385) );
  XNOR U7613 ( .A(n7393), .B(n7607), .Z(n7386) );
  XNOR U7614 ( .A(n7392), .B(n7390), .Z(n7607) );
  AND U7615 ( .A(n7608), .B(n7609), .Z(n7390) );
  NANDN U7616 ( .A(n7610), .B(n7611), .Z(n7609) );
  NANDN U7617 ( .A(n7612), .B(n7613), .Z(n7611) );
  NANDN U7618 ( .A(n7613), .B(n7612), .Z(n7608) );
  ANDN U7619 ( .B(B[31]), .A(n62), .Z(n7392) );
  XNOR U7620 ( .A(n7400), .B(n7614), .Z(n7393) );
  XNOR U7621 ( .A(n7399), .B(n7397), .Z(n7614) );
  AND U7622 ( .A(n7615), .B(n7616), .Z(n7397) );
  NANDN U7623 ( .A(n7617), .B(n7618), .Z(n7616) );
  OR U7624 ( .A(n7619), .B(n7620), .Z(n7618) );
  NAND U7625 ( .A(n7620), .B(n7619), .Z(n7615) );
  ANDN U7626 ( .B(B[32]), .A(n63), .Z(n7399) );
  XNOR U7627 ( .A(n7407), .B(n7621), .Z(n7400) );
  XNOR U7628 ( .A(n7406), .B(n7404), .Z(n7621) );
  AND U7629 ( .A(n7622), .B(n7623), .Z(n7404) );
  NANDN U7630 ( .A(n7624), .B(n7625), .Z(n7623) );
  NANDN U7631 ( .A(n7626), .B(n7627), .Z(n7625) );
  NANDN U7632 ( .A(n7627), .B(n7626), .Z(n7622) );
  ANDN U7633 ( .B(B[33]), .A(n64), .Z(n7406) );
  XNOR U7634 ( .A(n7414), .B(n7628), .Z(n7407) );
  XNOR U7635 ( .A(n7413), .B(n7411), .Z(n7628) );
  AND U7636 ( .A(n7629), .B(n7630), .Z(n7411) );
  NANDN U7637 ( .A(n7631), .B(n7632), .Z(n7630) );
  OR U7638 ( .A(n7633), .B(n7634), .Z(n7632) );
  NAND U7639 ( .A(n7634), .B(n7633), .Z(n7629) );
  ANDN U7640 ( .B(B[34]), .A(n65), .Z(n7413) );
  XNOR U7641 ( .A(n7421), .B(n7635), .Z(n7414) );
  XNOR U7642 ( .A(n7420), .B(n7418), .Z(n7635) );
  AND U7643 ( .A(n7636), .B(n7637), .Z(n7418) );
  NANDN U7644 ( .A(n7638), .B(n7639), .Z(n7637) );
  NANDN U7645 ( .A(n7640), .B(n7641), .Z(n7639) );
  NANDN U7646 ( .A(n7641), .B(n7640), .Z(n7636) );
  ANDN U7647 ( .B(B[35]), .A(n66), .Z(n7420) );
  XNOR U7648 ( .A(n7428), .B(n7642), .Z(n7421) );
  XNOR U7649 ( .A(n7427), .B(n7425), .Z(n7642) );
  AND U7650 ( .A(n7643), .B(n7644), .Z(n7425) );
  NANDN U7651 ( .A(n7645), .B(n7646), .Z(n7644) );
  OR U7652 ( .A(n7647), .B(n7648), .Z(n7646) );
  NAND U7653 ( .A(n7648), .B(n7647), .Z(n7643) );
  ANDN U7654 ( .B(B[36]), .A(n67), .Z(n7427) );
  XNOR U7655 ( .A(n7435), .B(n7649), .Z(n7428) );
  XNOR U7656 ( .A(n7434), .B(n7432), .Z(n7649) );
  AND U7657 ( .A(n7650), .B(n7651), .Z(n7432) );
  NANDN U7658 ( .A(n7652), .B(n7653), .Z(n7651) );
  NANDN U7659 ( .A(n7654), .B(n7655), .Z(n7653) );
  NANDN U7660 ( .A(n7655), .B(n7654), .Z(n7650) );
  ANDN U7661 ( .B(B[37]), .A(n68), .Z(n7434) );
  XNOR U7662 ( .A(n7442), .B(n7656), .Z(n7435) );
  XNOR U7663 ( .A(n7441), .B(n7439), .Z(n7656) );
  AND U7664 ( .A(n7657), .B(n7658), .Z(n7439) );
  NANDN U7665 ( .A(n7659), .B(n7660), .Z(n7658) );
  OR U7666 ( .A(n7661), .B(n7662), .Z(n7660) );
  NAND U7667 ( .A(n7662), .B(n7661), .Z(n7657) );
  ANDN U7668 ( .B(B[38]), .A(n69), .Z(n7441) );
  XNOR U7669 ( .A(n7449), .B(n7663), .Z(n7442) );
  XNOR U7670 ( .A(n7448), .B(n7446), .Z(n7663) );
  AND U7671 ( .A(n7664), .B(n7665), .Z(n7446) );
  NANDN U7672 ( .A(n7666), .B(n7667), .Z(n7665) );
  NANDN U7673 ( .A(n7668), .B(n7669), .Z(n7667) );
  NANDN U7674 ( .A(n7669), .B(n7668), .Z(n7664) );
  ANDN U7675 ( .B(B[39]), .A(n70), .Z(n7448) );
  XNOR U7676 ( .A(n7456), .B(n7670), .Z(n7449) );
  XNOR U7677 ( .A(n7455), .B(n7453), .Z(n7670) );
  AND U7678 ( .A(n7671), .B(n7672), .Z(n7453) );
  NANDN U7679 ( .A(n7673), .B(n7674), .Z(n7672) );
  OR U7680 ( .A(n7675), .B(n7676), .Z(n7674) );
  NAND U7681 ( .A(n7676), .B(n7675), .Z(n7671) );
  ANDN U7682 ( .B(B[40]), .A(n71), .Z(n7455) );
  XNOR U7683 ( .A(n7463), .B(n7677), .Z(n7456) );
  XNOR U7684 ( .A(n7462), .B(n7460), .Z(n7677) );
  AND U7685 ( .A(n7678), .B(n7679), .Z(n7460) );
  NANDN U7686 ( .A(n7680), .B(n7681), .Z(n7679) );
  NANDN U7687 ( .A(n7682), .B(n7683), .Z(n7681) );
  NANDN U7688 ( .A(n7683), .B(n7682), .Z(n7678) );
  ANDN U7689 ( .B(B[41]), .A(n72), .Z(n7462) );
  XNOR U7690 ( .A(n7470), .B(n7684), .Z(n7463) );
  XNOR U7691 ( .A(n7469), .B(n7467), .Z(n7684) );
  AND U7692 ( .A(n7685), .B(n7686), .Z(n7467) );
  NANDN U7693 ( .A(n7687), .B(n7688), .Z(n7686) );
  OR U7694 ( .A(n7689), .B(n7690), .Z(n7688) );
  NAND U7695 ( .A(n7690), .B(n7689), .Z(n7685) );
  ANDN U7696 ( .B(B[42]), .A(n73), .Z(n7469) );
  XNOR U7697 ( .A(n7477), .B(n7691), .Z(n7470) );
  XNOR U7698 ( .A(n7476), .B(n7474), .Z(n7691) );
  AND U7699 ( .A(n7692), .B(n7693), .Z(n7474) );
  NANDN U7700 ( .A(n7694), .B(n7695), .Z(n7693) );
  NANDN U7701 ( .A(n7696), .B(n7697), .Z(n7695) );
  NANDN U7702 ( .A(n7697), .B(n7696), .Z(n7692) );
  ANDN U7703 ( .B(B[43]), .A(n74), .Z(n7476) );
  XNOR U7704 ( .A(n7484), .B(n7698), .Z(n7477) );
  XNOR U7705 ( .A(n7483), .B(n7481), .Z(n7698) );
  AND U7706 ( .A(n7699), .B(n7700), .Z(n7481) );
  NANDN U7707 ( .A(n7701), .B(n7702), .Z(n7700) );
  OR U7708 ( .A(n7703), .B(n7704), .Z(n7702) );
  NAND U7709 ( .A(n7704), .B(n7703), .Z(n7699) );
  ANDN U7710 ( .B(B[44]), .A(n75), .Z(n7483) );
  XNOR U7711 ( .A(n7491), .B(n7705), .Z(n7484) );
  XNOR U7712 ( .A(n7490), .B(n7488), .Z(n7705) );
  AND U7713 ( .A(n7706), .B(n7707), .Z(n7488) );
  NANDN U7714 ( .A(n7708), .B(n7709), .Z(n7707) );
  NANDN U7715 ( .A(n7710), .B(n7711), .Z(n7709) );
  NANDN U7716 ( .A(n7711), .B(n7710), .Z(n7706) );
  ANDN U7717 ( .B(B[45]), .A(n76), .Z(n7490) );
  XNOR U7718 ( .A(n7498), .B(n7712), .Z(n7491) );
  XNOR U7719 ( .A(n7497), .B(n7495), .Z(n7712) );
  AND U7720 ( .A(n7713), .B(n7714), .Z(n7495) );
  NANDN U7721 ( .A(n7715), .B(n7716), .Z(n7714) );
  OR U7722 ( .A(n7717), .B(n7718), .Z(n7716) );
  NAND U7723 ( .A(n7718), .B(n7717), .Z(n7713) );
  ANDN U7724 ( .B(B[46]), .A(n77), .Z(n7497) );
  XNOR U7725 ( .A(n7505), .B(n7719), .Z(n7498) );
  XNOR U7726 ( .A(n7504), .B(n7502), .Z(n7719) );
  AND U7727 ( .A(n7720), .B(n7721), .Z(n7502) );
  NANDN U7728 ( .A(n7722), .B(n7723), .Z(n7721) );
  NANDN U7729 ( .A(n7724), .B(n7725), .Z(n7723) );
  NANDN U7730 ( .A(n7725), .B(n7724), .Z(n7720) );
  ANDN U7731 ( .B(B[47]), .A(n78), .Z(n7504) );
  XNOR U7732 ( .A(n7512), .B(n7726), .Z(n7505) );
  XNOR U7733 ( .A(n7511), .B(n7509), .Z(n7726) );
  AND U7734 ( .A(n7727), .B(n7728), .Z(n7509) );
  NANDN U7735 ( .A(n7729), .B(n7730), .Z(n7728) );
  OR U7736 ( .A(n7731), .B(n7732), .Z(n7730) );
  NAND U7737 ( .A(n7732), .B(n7731), .Z(n7727) );
  ANDN U7738 ( .B(B[48]), .A(n79), .Z(n7511) );
  XNOR U7739 ( .A(n7519), .B(n7733), .Z(n7512) );
  XNOR U7740 ( .A(n7518), .B(n7516), .Z(n7733) );
  AND U7741 ( .A(n7734), .B(n7735), .Z(n7516) );
  NANDN U7742 ( .A(n7736), .B(n7737), .Z(n7735) );
  NANDN U7743 ( .A(n7738), .B(n7739), .Z(n7737) );
  NANDN U7744 ( .A(n7739), .B(n7738), .Z(n7734) );
  ANDN U7745 ( .B(B[49]), .A(n80), .Z(n7518) );
  XNOR U7746 ( .A(n7526), .B(n7740), .Z(n7519) );
  XNOR U7747 ( .A(n7525), .B(n7523), .Z(n7740) );
  AND U7748 ( .A(n7741), .B(n7742), .Z(n7523) );
  NANDN U7749 ( .A(n7743), .B(n7744), .Z(n7742) );
  OR U7750 ( .A(n7745), .B(n7746), .Z(n7744) );
  NAND U7751 ( .A(n7746), .B(n7745), .Z(n7741) );
  ANDN U7752 ( .B(B[50]), .A(n81), .Z(n7525) );
  XNOR U7753 ( .A(n7533), .B(n7747), .Z(n7526) );
  XNOR U7754 ( .A(n7532), .B(n7530), .Z(n7747) );
  AND U7755 ( .A(n7748), .B(n7749), .Z(n7530) );
  NANDN U7756 ( .A(n7750), .B(n7751), .Z(n7749) );
  NAND U7757 ( .A(n7752), .B(n7753), .Z(n7751) );
  ANDN U7758 ( .B(B[51]), .A(n82), .Z(n7532) );
  XOR U7759 ( .A(n7539), .B(n7754), .Z(n7533) );
  XNOR U7760 ( .A(n7537), .B(n7540), .Z(n7754) );
  NAND U7761 ( .A(A[2]), .B(B[52]), .Z(n7540) );
  NANDN U7762 ( .A(n7755), .B(n7756), .Z(n7537) );
  AND U7763 ( .A(A[0]), .B(B[53]), .Z(n7756) );
  XNOR U7764 ( .A(n7542), .B(n7757), .Z(n7539) );
  NAND U7765 ( .A(A[0]), .B(B[54]), .Z(n7757) );
  NAND U7766 ( .A(B[53]), .B(A[1]), .Z(n7542) );
  NAND U7767 ( .A(n7758), .B(n7759), .Z(n179) );
  NANDN U7768 ( .A(n7760), .B(n7761), .Z(n7759) );
  OR U7769 ( .A(n7762), .B(n7763), .Z(n7761) );
  NAND U7770 ( .A(n7763), .B(n7762), .Z(n7758) );
  XOR U7771 ( .A(n181), .B(n180), .Z(\A1[51] ) );
  XOR U7772 ( .A(n7763), .B(n7764), .Z(n180) );
  XNOR U7773 ( .A(n7762), .B(n7760), .Z(n7764) );
  AND U7774 ( .A(n7765), .B(n7766), .Z(n7760) );
  NANDN U7775 ( .A(n7767), .B(n7768), .Z(n7766) );
  NANDN U7776 ( .A(n7769), .B(n7770), .Z(n7768) );
  NANDN U7777 ( .A(n7770), .B(n7769), .Z(n7765) );
  ANDN U7778 ( .B(B[22]), .A(n54), .Z(n7762) );
  XNOR U7779 ( .A(n7557), .B(n7771), .Z(n7763) );
  XNOR U7780 ( .A(n7556), .B(n7554), .Z(n7771) );
  AND U7781 ( .A(n7772), .B(n7773), .Z(n7554) );
  NANDN U7782 ( .A(n7774), .B(n7775), .Z(n7773) );
  OR U7783 ( .A(n7776), .B(n7777), .Z(n7775) );
  NAND U7784 ( .A(n7777), .B(n7776), .Z(n7772) );
  ANDN U7785 ( .B(B[23]), .A(n55), .Z(n7556) );
  XNOR U7786 ( .A(n7564), .B(n7778), .Z(n7557) );
  XNOR U7787 ( .A(n7563), .B(n7561), .Z(n7778) );
  AND U7788 ( .A(n7779), .B(n7780), .Z(n7561) );
  NANDN U7789 ( .A(n7781), .B(n7782), .Z(n7780) );
  NANDN U7790 ( .A(n7783), .B(n7784), .Z(n7782) );
  NANDN U7791 ( .A(n7784), .B(n7783), .Z(n7779) );
  ANDN U7792 ( .B(B[24]), .A(n56), .Z(n7563) );
  XNOR U7793 ( .A(n7571), .B(n7785), .Z(n7564) );
  XNOR U7794 ( .A(n7570), .B(n7568), .Z(n7785) );
  AND U7795 ( .A(n7786), .B(n7787), .Z(n7568) );
  NANDN U7796 ( .A(n7788), .B(n7789), .Z(n7787) );
  OR U7797 ( .A(n7790), .B(n7791), .Z(n7789) );
  NAND U7798 ( .A(n7791), .B(n7790), .Z(n7786) );
  ANDN U7799 ( .B(B[25]), .A(n57), .Z(n7570) );
  XNOR U7800 ( .A(n7578), .B(n7792), .Z(n7571) );
  XNOR U7801 ( .A(n7577), .B(n7575), .Z(n7792) );
  AND U7802 ( .A(n7793), .B(n7794), .Z(n7575) );
  NANDN U7803 ( .A(n7795), .B(n7796), .Z(n7794) );
  NANDN U7804 ( .A(n7797), .B(n7798), .Z(n7796) );
  NANDN U7805 ( .A(n7798), .B(n7797), .Z(n7793) );
  ANDN U7806 ( .B(B[26]), .A(n58), .Z(n7577) );
  XNOR U7807 ( .A(n7585), .B(n7799), .Z(n7578) );
  XNOR U7808 ( .A(n7584), .B(n7582), .Z(n7799) );
  AND U7809 ( .A(n7800), .B(n7801), .Z(n7582) );
  NANDN U7810 ( .A(n7802), .B(n7803), .Z(n7801) );
  OR U7811 ( .A(n7804), .B(n7805), .Z(n7803) );
  NAND U7812 ( .A(n7805), .B(n7804), .Z(n7800) );
  ANDN U7813 ( .B(B[27]), .A(n59), .Z(n7584) );
  XNOR U7814 ( .A(n7592), .B(n7806), .Z(n7585) );
  XNOR U7815 ( .A(n7591), .B(n7589), .Z(n7806) );
  AND U7816 ( .A(n7807), .B(n7808), .Z(n7589) );
  NANDN U7817 ( .A(n7809), .B(n7810), .Z(n7808) );
  NANDN U7818 ( .A(n7811), .B(n7812), .Z(n7810) );
  NANDN U7819 ( .A(n7812), .B(n7811), .Z(n7807) );
  ANDN U7820 ( .B(B[28]), .A(n60), .Z(n7591) );
  XNOR U7821 ( .A(n7599), .B(n7813), .Z(n7592) );
  XNOR U7822 ( .A(n7598), .B(n7596), .Z(n7813) );
  AND U7823 ( .A(n7814), .B(n7815), .Z(n7596) );
  NANDN U7824 ( .A(n7816), .B(n7817), .Z(n7815) );
  OR U7825 ( .A(n7818), .B(n7819), .Z(n7817) );
  NAND U7826 ( .A(n7819), .B(n7818), .Z(n7814) );
  ANDN U7827 ( .B(B[29]), .A(n61), .Z(n7598) );
  XNOR U7828 ( .A(n7606), .B(n7820), .Z(n7599) );
  XNOR U7829 ( .A(n7605), .B(n7603), .Z(n7820) );
  AND U7830 ( .A(n7821), .B(n7822), .Z(n7603) );
  NANDN U7831 ( .A(n7823), .B(n7824), .Z(n7822) );
  NANDN U7832 ( .A(n7825), .B(n7826), .Z(n7824) );
  NANDN U7833 ( .A(n7826), .B(n7825), .Z(n7821) );
  ANDN U7834 ( .B(B[30]), .A(n62), .Z(n7605) );
  XNOR U7835 ( .A(n7613), .B(n7827), .Z(n7606) );
  XNOR U7836 ( .A(n7612), .B(n7610), .Z(n7827) );
  AND U7837 ( .A(n7828), .B(n7829), .Z(n7610) );
  NANDN U7838 ( .A(n7830), .B(n7831), .Z(n7829) );
  OR U7839 ( .A(n7832), .B(n7833), .Z(n7831) );
  NAND U7840 ( .A(n7833), .B(n7832), .Z(n7828) );
  ANDN U7841 ( .B(B[31]), .A(n63), .Z(n7612) );
  XNOR U7842 ( .A(n7620), .B(n7834), .Z(n7613) );
  XNOR U7843 ( .A(n7619), .B(n7617), .Z(n7834) );
  AND U7844 ( .A(n7835), .B(n7836), .Z(n7617) );
  NANDN U7845 ( .A(n7837), .B(n7838), .Z(n7836) );
  NANDN U7846 ( .A(n7839), .B(n7840), .Z(n7838) );
  NANDN U7847 ( .A(n7840), .B(n7839), .Z(n7835) );
  ANDN U7848 ( .B(B[32]), .A(n64), .Z(n7619) );
  XNOR U7849 ( .A(n7627), .B(n7841), .Z(n7620) );
  XNOR U7850 ( .A(n7626), .B(n7624), .Z(n7841) );
  AND U7851 ( .A(n7842), .B(n7843), .Z(n7624) );
  NANDN U7852 ( .A(n7844), .B(n7845), .Z(n7843) );
  OR U7853 ( .A(n7846), .B(n7847), .Z(n7845) );
  NAND U7854 ( .A(n7847), .B(n7846), .Z(n7842) );
  ANDN U7855 ( .B(B[33]), .A(n65), .Z(n7626) );
  XNOR U7856 ( .A(n7634), .B(n7848), .Z(n7627) );
  XNOR U7857 ( .A(n7633), .B(n7631), .Z(n7848) );
  AND U7858 ( .A(n7849), .B(n7850), .Z(n7631) );
  NANDN U7859 ( .A(n7851), .B(n7852), .Z(n7850) );
  NANDN U7860 ( .A(n7853), .B(n7854), .Z(n7852) );
  NANDN U7861 ( .A(n7854), .B(n7853), .Z(n7849) );
  ANDN U7862 ( .B(B[34]), .A(n66), .Z(n7633) );
  XNOR U7863 ( .A(n7641), .B(n7855), .Z(n7634) );
  XNOR U7864 ( .A(n7640), .B(n7638), .Z(n7855) );
  AND U7865 ( .A(n7856), .B(n7857), .Z(n7638) );
  NANDN U7866 ( .A(n7858), .B(n7859), .Z(n7857) );
  OR U7867 ( .A(n7860), .B(n7861), .Z(n7859) );
  NAND U7868 ( .A(n7861), .B(n7860), .Z(n7856) );
  ANDN U7869 ( .B(B[35]), .A(n67), .Z(n7640) );
  XNOR U7870 ( .A(n7648), .B(n7862), .Z(n7641) );
  XNOR U7871 ( .A(n7647), .B(n7645), .Z(n7862) );
  AND U7872 ( .A(n7863), .B(n7864), .Z(n7645) );
  NANDN U7873 ( .A(n7865), .B(n7866), .Z(n7864) );
  NANDN U7874 ( .A(n7867), .B(n7868), .Z(n7866) );
  NANDN U7875 ( .A(n7868), .B(n7867), .Z(n7863) );
  ANDN U7876 ( .B(B[36]), .A(n68), .Z(n7647) );
  XNOR U7877 ( .A(n7655), .B(n7869), .Z(n7648) );
  XNOR U7878 ( .A(n7654), .B(n7652), .Z(n7869) );
  AND U7879 ( .A(n7870), .B(n7871), .Z(n7652) );
  NANDN U7880 ( .A(n7872), .B(n7873), .Z(n7871) );
  OR U7881 ( .A(n7874), .B(n7875), .Z(n7873) );
  NAND U7882 ( .A(n7875), .B(n7874), .Z(n7870) );
  ANDN U7883 ( .B(B[37]), .A(n69), .Z(n7654) );
  XNOR U7884 ( .A(n7662), .B(n7876), .Z(n7655) );
  XNOR U7885 ( .A(n7661), .B(n7659), .Z(n7876) );
  AND U7886 ( .A(n7877), .B(n7878), .Z(n7659) );
  NANDN U7887 ( .A(n7879), .B(n7880), .Z(n7878) );
  NANDN U7888 ( .A(n7881), .B(n7882), .Z(n7880) );
  NANDN U7889 ( .A(n7882), .B(n7881), .Z(n7877) );
  ANDN U7890 ( .B(B[38]), .A(n70), .Z(n7661) );
  XNOR U7891 ( .A(n7669), .B(n7883), .Z(n7662) );
  XNOR U7892 ( .A(n7668), .B(n7666), .Z(n7883) );
  AND U7893 ( .A(n7884), .B(n7885), .Z(n7666) );
  NANDN U7894 ( .A(n7886), .B(n7887), .Z(n7885) );
  OR U7895 ( .A(n7888), .B(n7889), .Z(n7887) );
  NAND U7896 ( .A(n7889), .B(n7888), .Z(n7884) );
  ANDN U7897 ( .B(B[39]), .A(n71), .Z(n7668) );
  XNOR U7898 ( .A(n7676), .B(n7890), .Z(n7669) );
  XNOR U7899 ( .A(n7675), .B(n7673), .Z(n7890) );
  AND U7900 ( .A(n7891), .B(n7892), .Z(n7673) );
  NANDN U7901 ( .A(n7893), .B(n7894), .Z(n7892) );
  NANDN U7902 ( .A(n7895), .B(n7896), .Z(n7894) );
  NANDN U7903 ( .A(n7896), .B(n7895), .Z(n7891) );
  ANDN U7904 ( .B(B[40]), .A(n72), .Z(n7675) );
  XNOR U7905 ( .A(n7683), .B(n7897), .Z(n7676) );
  XNOR U7906 ( .A(n7682), .B(n7680), .Z(n7897) );
  AND U7907 ( .A(n7898), .B(n7899), .Z(n7680) );
  NANDN U7908 ( .A(n7900), .B(n7901), .Z(n7899) );
  OR U7909 ( .A(n7902), .B(n7903), .Z(n7901) );
  NAND U7910 ( .A(n7903), .B(n7902), .Z(n7898) );
  ANDN U7911 ( .B(B[41]), .A(n73), .Z(n7682) );
  XNOR U7912 ( .A(n7690), .B(n7904), .Z(n7683) );
  XNOR U7913 ( .A(n7689), .B(n7687), .Z(n7904) );
  AND U7914 ( .A(n7905), .B(n7906), .Z(n7687) );
  NANDN U7915 ( .A(n7907), .B(n7908), .Z(n7906) );
  NANDN U7916 ( .A(n7909), .B(n7910), .Z(n7908) );
  NANDN U7917 ( .A(n7910), .B(n7909), .Z(n7905) );
  ANDN U7918 ( .B(B[42]), .A(n74), .Z(n7689) );
  XNOR U7919 ( .A(n7697), .B(n7911), .Z(n7690) );
  XNOR U7920 ( .A(n7696), .B(n7694), .Z(n7911) );
  AND U7921 ( .A(n7912), .B(n7913), .Z(n7694) );
  NANDN U7922 ( .A(n7914), .B(n7915), .Z(n7913) );
  OR U7923 ( .A(n7916), .B(n7917), .Z(n7915) );
  NAND U7924 ( .A(n7917), .B(n7916), .Z(n7912) );
  ANDN U7925 ( .B(B[43]), .A(n75), .Z(n7696) );
  XNOR U7926 ( .A(n7704), .B(n7918), .Z(n7697) );
  XNOR U7927 ( .A(n7703), .B(n7701), .Z(n7918) );
  AND U7928 ( .A(n7919), .B(n7920), .Z(n7701) );
  NANDN U7929 ( .A(n7921), .B(n7922), .Z(n7920) );
  NANDN U7930 ( .A(n7923), .B(n7924), .Z(n7922) );
  NANDN U7931 ( .A(n7924), .B(n7923), .Z(n7919) );
  ANDN U7932 ( .B(B[44]), .A(n76), .Z(n7703) );
  XNOR U7933 ( .A(n7711), .B(n7925), .Z(n7704) );
  XNOR U7934 ( .A(n7710), .B(n7708), .Z(n7925) );
  AND U7935 ( .A(n7926), .B(n7927), .Z(n7708) );
  NANDN U7936 ( .A(n7928), .B(n7929), .Z(n7927) );
  OR U7937 ( .A(n7930), .B(n7931), .Z(n7929) );
  NAND U7938 ( .A(n7931), .B(n7930), .Z(n7926) );
  ANDN U7939 ( .B(B[45]), .A(n77), .Z(n7710) );
  XNOR U7940 ( .A(n7718), .B(n7932), .Z(n7711) );
  XNOR U7941 ( .A(n7717), .B(n7715), .Z(n7932) );
  AND U7942 ( .A(n7933), .B(n7934), .Z(n7715) );
  NANDN U7943 ( .A(n7935), .B(n7936), .Z(n7934) );
  NANDN U7944 ( .A(n7937), .B(n7938), .Z(n7936) );
  NANDN U7945 ( .A(n7938), .B(n7937), .Z(n7933) );
  ANDN U7946 ( .B(B[46]), .A(n78), .Z(n7717) );
  XNOR U7947 ( .A(n7725), .B(n7939), .Z(n7718) );
  XNOR U7948 ( .A(n7724), .B(n7722), .Z(n7939) );
  AND U7949 ( .A(n7940), .B(n7941), .Z(n7722) );
  NANDN U7950 ( .A(n7942), .B(n7943), .Z(n7941) );
  OR U7951 ( .A(n7944), .B(n7945), .Z(n7943) );
  NAND U7952 ( .A(n7945), .B(n7944), .Z(n7940) );
  ANDN U7953 ( .B(B[47]), .A(n79), .Z(n7724) );
  XNOR U7954 ( .A(n7732), .B(n7946), .Z(n7725) );
  XNOR U7955 ( .A(n7731), .B(n7729), .Z(n7946) );
  AND U7956 ( .A(n7947), .B(n7948), .Z(n7729) );
  NANDN U7957 ( .A(n7949), .B(n7950), .Z(n7948) );
  NANDN U7958 ( .A(n7951), .B(n7952), .Z(n7950) );
  NANDN U7959 ( .A(n7952), .B(n7951), .Z(n7947) );
  ANDN U7960 ( .B(B[48]), .A(n80), .Z(n7731) );
  XNOR U7961 ( .A(n7739), .B(n7953), .Z(n7732) );
  XNOR U7962 ( .A(n7738), .B(n7736), .Z(n7953) );
  AND U7963 ( .A(n7954), .B(n7955), .Z(n7736) );
  NANDN U7964 ( .A(n7956), .B(n7957), .Z(n7955) );
  OR U7965 ( .A(n7958), .B(n7959), .Z(n7957) );
  NAND U7966 ( .A(n7959), .B(n7958), .Z(n7954) );
  ANDN U7967 ( .B(B[49]), .A(n81), .Z(n7738) );
  XNOR U7968 ( .A(n7746), .B(n7960), .Z(n7739) );
  XNOR U7969 ( .A(n7745), .B(n7743), .Z(n7960) );
  AND U7970 ( .A(n7961), .B(n7962), .Z(n7743) );
  NANDN U7971 ( .A(n7963), .B(n7964), .Z(n7962) );
  NAND U7972 ( .A(n7965), .B(n7966), .Z(n7964) );
  ANDN U7973 ( .B(B[50]), .A(n82), .Z(n7745) );
  XOR U7974 ( .A(n7752), .B(n7967), .Z(n7746) );
  XNOR U7975 ( .A(n7750), .B(n7753), .Z(n7967) );
  NAND U7976 ( .A(A[2]), .B(B[51]), .Z(n7753) );
  NANDN U7977 ( .A(n7968), .B(n7969), .Z(n7750) );
  AND U7978 ( .A(A[0]), .B(B[52]), .Z(n7969) );
  XNOR U7979 ( .A(n7755), .B(n7970), .Z(n7752) );
  NAND U7980 ( .A(A[0]), .B(B[53]), .Z(n7970) );
  NAND U7981 ( .A(B[52]), .B(A[1]), .Z(n7755) );
  NAND U7982 ( .A(n7971), .B(n7972), .Z(n181) );
  NANDN U7983 ( .A(n7973), .B(n7974), .Z(n7972) );
  OR U7984 ( .A(n7975), .B(n7976), .Z(n7974) );
  NAND U7985 ( .A(n7976), .B(n7975), .Z(n7971) );
  XOR U7986 ( .A(n183), .B(n182), .Z(\A1[50] ) );
  XOR U7987 ( .A(n7976), .B(n7977), .Z(n182) );
  XNOR U7988 ( .A(n7975), .B(n7973), .Z(n7977) );
  AND U7989 ( .A(n7978), .B(n7979), .Z(n7973) );
  NANDN U7990 ( .A(n7980), .B(n7981), .Z(n7979) );
  NANDN U7991 ( .A(n7982), .B(n7983), .Z(n7981) );
  NANDN U7992 ( .A(n7983), .B(n7982), .Z(n7978) );
  ANDN U7993 ( .B(B[21]), .A(n54), .Z(n7975) );
  XNOR U7994 ( .A(n7770), .B(n7984), .Z(n7976) );
  XNOR U7995 ( .A(n7769), .B(n7767), .Z(n7984) );
  AND U7996 ( .A(n7985), .B(n7986), .Z(n7767) );
  NANDN U7997 ( .A(n7987), .B(n7988), .Z(n7986) );
  OR U7998 ( .A(n7989), .B(n7990), .Z(n7988) );
  NAND U7999 ( .A(n7990), .B(n7989), .Z(n7985) );
  ANDN U8000 ( .B(B[22]), .A(n55), .Z(n7769) );
  XNOR U8001 ( .A(n7777), .B(n7991), .Z(n7770) );
  XNOR U8002 ( .A(n7776), .B(n7774), .Z(n7991) );
  AND U8003 ( .A(n7992), .B(n7993), .Z(n7774) );
  NANDN U8004 ( .A(n7994), .B(n7995), .Z(n7993) );
  NANDN U8005 ( .A(n7996), .B(n7997), .Z(n7995) );
  NANDN U8006 ( .A(n7997), .B(n7996), .Z(n7992) );
  ANDN U8007 ( .B(B[23]), .A(n56), .Z(n7776) );
  XNOR U8008 ( .A(n7784), .B(n7998), .Z(n7777) );
  XNOR U8009 ( .A(n7783), .B(n7781), .Z(n7998) );
  AND U8010 ( .A(n7999), .B(n8000), .Z(n7781) );
  NANDN U8011 ( .A(n8001), .B(n8002), .Z(n8000) );
  OR U8012 ( .A(n8003), .B(n8004), .Z(n8002) );
  NAND U8013 ( .A(n8004), .B(n8003), .Z(n7999) );
  ANDN U8014 ( .B(B[24]), .A(n57), .Z(n7783) );
  XNOR U8015 ( .A(n7791), .B(n8005), .Z(n7784) );
  XNOR U8016 ( .A(n7790), .B(n7788), .Z(n8005) );
  AND U8017 ( .A(n8006), .B(n8007), .Z(n7788) );
  NANDN U8018 ( .A(n8008), .B(n8009), .Z(n8007) );
  NANDN U8019 ( .A(n8010), .B(n8011), .Z(n8009) );
  NANDN U8020 ( .A(n8011), .B(n8010), .Z(n8006) );
  ANDN U8021 ( .B(B[25]), .A(n58), .Z(n7790) );
  XNOR U8022 ( .A(n7798), .B(n8012), .Z(n7791) );
  XNOR U8023 ( .A(n7797), .B(n7795), .Z(n8012) );
  AND U8024 ( .A(n8013), .B(n8014), .Z(n7795) );
  NANDN U8025 ( .A(n8015), .B(n8016), .Z(n8014) );
  OR U8026 ( .A(n8017), .B(n8018), .Z(n8016) );
  NAND U8027 ( .A(n8018), .B(n8017), .Z(n8013) );
  ANDN U8028 ( .B(B[26]), .A(n59), .Z(n7797) );
  XNOR U8029 ( .A(n7805), .B(n8019), .Z(n7798) );
  XNOR U8030 ( .A(n7804), .B(n7802), .Z(n8019) );
  AND U8031 ( .A(n8020), .B(n8021), .Z(n7802) );
  NANDN U8032 ( .A(n8022), .B(n8023), .Z(n8021) );
  NANDN U8033 ( .A(n8024), .B(n8025), .Z(n8023) );
  NANDN U8034 ( .A(n8025), .B(n8024), .Z(n8020) );
  ANDN U8035 ( .B(B[27]), .A(n60), .Z(n7804) );
  XNOR U8036 ( .A(n7812), .B(n8026), .Z(n7805) );
  XNOR U8037 ( .A(n7811), .B(n7809), .Z(n8026) );
  AND U8038 ( .A(n8027), .B(n8028), .Z(n7809) );
  NANDN U8039 ( .A(n8029), .B(n8030), .Z(n8028) );
  OR U8040 ( .A(n8031), .B(n8032), .Z(n8030) );
  NAND U8041 ( .A(n8032), .B(n8031), .Z(n8027) );
  ANDN U8042 ( .B(B[28]), .A(n61), .Z(n7811) );
  XNOR U8043 ( .A(n7819), .B(n8033), .Z(n7812) );
  XNOR U8044 ( .A(n7818), .B(n7816), .Z(n8033) );
  AND U8045 ( .A(n8034), .B(n8035), .Z(n7816) );
  NANDN U8046 ( .A(n8036), .B(n8037), .Z(n8035) );
  NANDN U8047 ( .A(n8038), .B(n8039), .Z(n8037) );
  NANDN U8048 ( .A(n8039), .B(n8038), .Z(n8034) );
  ANDN U8049 ( .B(B[29]), .A(n62), .Z(n7818) );
  XNOR U8050 ( .A(n7826), .B(n8040), .Z(n7819) );
  XNOR U8051 ( .A(n7825), .B(n7823), .Z(n8040) );
  AND U8052 ( .A(n8041), .B(n8042), .Z(n7823) );
  NANDN U8053 ( .A(n8043), .B(n8044), .Z(n8042) );
  OR U8054 ( .A(n8045), .B(n8046), .Z(n8044) );
  NAND U8055 ( .A(n8046), .B(n8045), .Z(n8041) );
  ANDN U8056 ( .B(B[30]), .A(n63), .Z(n7825) );
  XNOR U8057 ( .A(n7833), .B(n8047), .Z(n7826) );
  XNOR U8058 ( .A(n7832), .B(n7830), .Z(n8047) );
  AND U8059 ( .A(n8048), .B(n8049), .Z(n7830) );
  NANDN U8060 ( .A(n8050), .B(n8051), .Z(n8049) );
  NANDN U8061 ( .A(n8052), .B(n8053), .Z(n8051) );
  NANDN U8062 ( .A(n8053), .B(n8052), .Z(n8048) );
  ANDN U8063 ( .B(B[31]), .A(n64), .Z(n7832) );
  XNOR U8064 ( .A(n7840), .B(n8054), .Z(n7833) );
  XNOR U8065 ( .A(n7839), .B(n7837), .Z(n8054) );
  AND U8066 ( .A(n8055), .B(n8056), .Z(n7837) );
  NANDN U8067 ( .A(n8057), .B(n8058), .Z(n8056) );
  OR U8068 ( .A(n8059), .B(n8060), .Z(n8058) );
  NAND U8069 ( .A(n8060), .B(n8059), .Z(n8055) );
  ANDN U8070 ( .B(B[32]), .A(n65), .Z(n7839) );
  XNOR U8071 ( .A(n7847), .B(n8061), .Z(n7840) );
  XNOR U8072 ( .A(n7846), .B(n7844), .Z(n8061) );
  AND U8073 ( .A(n8062), .B(n8063), .Z(n7844) );
  NANDN U8074 ( .A(n8064), .B(n8065), .Z(n8063) );
  NANDN U8075 ( .A(n8066), .B(n8067), .Z(n8065) );
  NANDN U8076 ( .A(n8067), .B(n8066), .Z(n8062) );
  ANDN U8077 ( .B(B[33]), .A(n66), .Z(n7846) );
  XNOR U8078 ( .A(n7854), .B(n8068), .Z(n7847) );
  XNOR U8079 ( .A(n7853), .B(n7851), .Z(n8068) );
  AND U8080 ( .A(n8069), .B(n8070), .Z(n7851) );
  NANDN U8081 ( .A(n8071), .B(n8072), .Z(n8070) );
  OR U8082 ( .A(n8073), .B(n8074), .Z(n8072) );
  NAND U8083 ( .A(n8074), .B(n8073), .Z(n8069) );
  ANDN U8084 ( .B(B[34]), .A(n67), .Z(n7853) );
  XNOR U8085 ( .A(n7861), .B(n8075), .Z(n7854) );
  XNOR U8086 ( .A(n7860), .B(n7858), .Z(n8075) );
  AND U8087 ( .A(n8076), .B(n8077), .Z(n7858) );
  NANDN U8088 ( .A(n8078), .B(n8079), .Z(n8077) );
  NANDN U8089 ( .A(n8080), .B(n8081), .Z(n8079) );
  NANDN U8090 ( .A(n8081), .B(n8080), .Z(n8076) );
  ANDN U8091 ( .B(B[35]), .A(n68), .Z(n7860) );
  XNOR U8092 ( .A(n7868), .B(n8082), .Z(n7861) );
  XNOR U8093 ( .A(n7867), .B(n7865), .Z(n8082) );
  AND U8094 ( .A(n8083), .B(n8084), .Z(n7865) );
  NANDN U8095 ( .A(n8085), .B(n8086), .Z(n8084) );
  OR U8096 ( .A(n8087), .B(n8088), .Z(n8086) );
  NAND U8097 ( .A(n8088), .B(n8087), .Z(n8083) );
  ANDN U8098 ( .B(B[36]), .A(n69), .Z(n7867) );
  XNOR U8099 ( .A(n7875), .B(n8089), .Z(n7868) );
  XNOR U8100 ( .A(n7874), .B(n7872), .Z(n8089) );
  AND U8101 ( .A(n8090), .B(n8091), .Z(n7872) );
  NANDN U8102 ( .A(n8092), .B(n8093), .Z(n8091) );
  NANDN U8103 ( .A(n8094), .B(n8095), .Z(n8093) );
  NANDN U8104 ( .A(n8095), .B(n8094), .Z(n8090) );
  ANDN U8105 ( .B(B[37]), .A(n70), .Z(n7874) );
  XNOR U8106 ( .A(n7882), .B(n8096), .Z(n7875) );
  XNOR U8107 ( .A(n7881), .B(n7879), .Z(n8096) );
  AND U8108 ( .A(n8097), .B(n8098), .Z(n7879) );
  NANDN U8109 ( .A(n8099), .B(n8100), .Z(n8098) );
  OR U8110 ( .A(n8101), .B(n8102), .Z(n8100) );
  NAND U8111 ( .A(n8102), .B(n8101), .Z(n8097) );
  ANDN U8112 ( .B(B[38]), .A(n71), .Z(n7881) );
  XNOR U8113 ( .A(n7889), .B(n8103), .Z(n7882) );
  XNOR U8114 ( .A(n7888), .B(n7886), .Z(n8103) );
  AND U8115 ( .A(n8104), .B(n8105), .Z(n7886) );
  NANDN U8116 ( .A(n8106), .B(n8107), .Z(n8105) );
  NANDN U8117 ( .A(n8108), .B(n8109), .Z(n8107) );
  NANDN U8118 ( .A(n8109), .B(n8108), .Z(n8104) );
  ANDN U8119 ( .B(B[39]), .A(n72), .Z(n7888) );
  XNOR U8120 ( .A(n7896), .B(n8110), .Z(n7889) );
  XNOR U8121 ( .A(n7895), .B(n7893), .Z(n8110) );
  AND U8122 ( .A(n8111), .B(n8112), .Z(n7893) );
  NANDN U8123 ( .A(n8113), .B(n8114), .Z(n8112) );
  OR U8124 ( .A(n8115), .B(n8116), .Z(n8114) );
  NAND U8125 ( .A(n8116), .B(n8115), .Z(n8111) );
  ANDN U8126 ( .B(B[40]), .A(n73), .Z(n7895) );
  XNOR U8127 ( .A(n7903), .B(n8117), .Z(n7896) );
  XNOR U8128 ( .A(n7902), .B(n7900), .Z(n8117) );
  AND U8129 ( .A(n8118), .B(n8119), .Z(n7900) );
  NANDN U8130 ( .A(n8120), .B(n8121), .Z(n8119) );
  NANDN U8131 ( .A(n8122), .B(n8123), .Z(n8121) );
  NANDN U8132 ( .A(n8123), .B(n8122), .Z(n8118) );
  ANDN U8133 ( .B(B[41]), .A(n74), .Z(n7902) );
  XNOR U8134 ( .A(n7910), .B(n8124), .Z(n7903) );
  XNOR U8135 ( .A(n7909), .B(n7907), .Z(n8124) );
  AND U8136 ( .A(n8125), .B(n8126), .Z(n7907) );
  NANDN U8137 ( .A(n8127), .B(n8128), .Z(n8126) );
  OR U8138 ( .A(n8129), .B(n8130), .Z(n8128) );
  NAND U8139 ( .A(n8130), .B(n8129), .Z(n8125) );
  ANDN U8140 ( .B(B[42]), .A(n75), .Z(n7909) );
  XNOR U8141 ( .A(n7917), .B(n8131), .Z(n7910) );
  XNOR U8142 ( .A(n7916), .B(n7914), .Z(n8131) );
  AND U8143 ( .A(n8132), .B(n8133), .Z(n7914) );
  NANDN U8144 ( .A(n8134), .B(n8135), .Z(n8133) );
  NANDN U8145 ( .A(n8136), .B(n8137), .Z(n8135) );
  NANDN U8146 ( .A(n8137), .B(n8136), .Z(n8132) );
  ANDN U8147 ( .B(B[43]), .A(n76), .Z(n7916) );
  XNOR U8148 ( .A(n7924), .B(n8138), .Z(n7917) );
  XNOR U8149 ( .A(n7923), .B(n7921), .Z(n8138) );
  AND U8150 ( .A(n8139), .B(n8140), .Z(n7921) );
  NANDN U8151 ( .A(n8141), .B(n8142), .Z(n8140) );
  OR U8152 ( .A(n8143), .B(n8144), .Z(n8142) );
  NAND U8153 ( .A(n8144), .B(n8143), .Z(n8139) );
  ANDN U8154 ( .B(B[44]), .A(n77), .Z(n7923) );
  XNOR U8155 ( .A(n7931), .B(n8145), .Z(n7924) );
  XNOR U8156 ( .A(n7930), .B(n7928), .Z(n8145) );
  AND U8157 ( .A(n8146), .B(n8147), .Z(n7928) );
  NANDN U8158 ( .A(n8148), .B(n8149), .Z(n8147) );
  NANDN U8159 ( .A(n8150), .B(n8151), .Z(n8149) );
  NANDN U8160 ( .A(n8151), .B(n8150), .Z(n8146) );
  ANDN U8161 ( .B(B[45]), .A(n78), .Z(n7930) );
  XNOR U8162 ( .A(n7938), .B(n8152), .Z(n7931) );
  XNOR U8163 ( .A(n7937), .B(n7935), .Z(n8152) );
  AND U8164 ( .A(n8153), .B(n8154), .Z(n7935) );
  NANDN U8165 ( .A(n8155), .B(n8156), .Z(n8154) );
  OR U8166 ( .A(n8157), .B(n8158), .Z(n8156) );
  NAND U8167 ( .A(n8158), .B(n8157), .Z(n8153) );
  ANDN U8168 ( .B(B[46]), .A(n79), .Z(n7937) );
  XNOR U8169 ( .A(n7945), .B(n8159), .Z(n7938) );
  XNOR U8170 ( .A(n7944), .B(n7942), .Z(n8159) );
  AND U8171 ( .A(n8160), .B(n8161), .Z(n7942) );
  NANDN U8172 ( .A(n8162), .B(n8163), .Z(n8161) );
  NANDN U8173 ( .A(n8164), .B(n8165), .Z(n8163) );
  NANDN U8174 ( .A(n8165), .B(n8164), .Z(n8160) );
  ANDN U8175 ( .B(B[47]), .A(n80), .Z(n7944) );
  XNOR U8176 ( .A(n7952), .B(n8166), .Z(n7945) );
  XNOR U8177 ( .A(n7951), .B(n7949), .Z(n8166) );
  AND U8178 ( .A(n8167), .B(n8168), .Z(n7949) );
  NANDN U8179 ( .A(n8169), .B(n8170), .Z(n8168) );
  OR U8180 ( .A(n8171), .B(n8172), .Z(n8170) );
  NAND U8181 ( .A(n8172), .B(n8171), .Z(n8167) );
  ANDN U8182 ( .B(B[48]), .A(n81), .Z(n7951) );
  XNOR U8183 ( .A(n7959), .B(n8173), .Z(n7952) );
  XNOR U8184 ( .A(n7958), .B(n7956), .Z(n8173) );
  AND U8185 ( .A(n8174), .B(n8175), .Z(n7956) );
  NANDN U8186 ( .A(n8176), .B(n8177), .Z(n8175) );
  NAND U8187 ( .A(n8178), .B(n8179), .Z(n8177) );
  ANDN U8188 ( .B(B[49]), .A(n82), .Z(n7958) );
  XOR U8189 ( .A(n7965), .B(n8180), .Z(n7959) );
  XNOR U8190 ( .A(n7963), .B(n7966), .Z(n8180) );
  NAND U8191 ( .A(A[2]), .B(B[50]), .Z(n7966) );
  NANDN U8192 ( .A(n8181), .B(n8182), .Z(n7963) );
  AND U8193 ( .A(A[0]), .B(B[51]), .Z(n8182) );
  XNOR U8194 ( .A(n7968), .B(n8183), .Z(n7965) );
  NAND U8195 ( .A(A[0]), .B(B[52]), .Z(n8183) );
  NAND U8196 ( .A(B[51]), .B(A[1]), .Z(n7968) );
  NAND U8197 ( .A(n8184), .B(n8185), .Z(n183) );
  NANDN U8198 ( .A(n8186), .B(n8187), .Z(n8185) );
  OR U8199 ( .A(n8188), .B(n8189), .Z(n8187) );
  NAND U8200 ( .A(n8189), .B(n8188), .Z(n8184) );
  XNOR U8201 ( .A(n8190), .B(n8191), .Z(\A1[4] ) );
  XNOR U8202 ( .A(n8192), .B(n8193), .Z(n8191) );
  XOR U8203 ( .A(n185), .B(n184), .Z(\A1[49] ) );
  XOR U8204 ( .A(n8189), .B(n8194), .Z(n184) );
  XNOR U8205 ( .A(n8188), .B(n8186), .Z(n8194) );
  AND U8206 ( .A(n8195), .B(n8196), .Z(n8186) );
  NANDN U8207 ( .A(n8197), .B(n8198), .Z(n8196) );
  NANDN U8208 ( .A(n8199), .B(n8200), .Z(n8198) );
  NANDN U8209 ( .A(n8200), .B(n8199), .Z(n8195) );
  ANDN U8210 ( .B(B[20]), .A(n54), .Z(n8188) );
  XNOR U8211 ( .A(n7983), .B(n8201), .Z(n8189) );
  XNOR U8212 ( .A(n7982), .B(n7980), .Z(n8201) );
  AND U8213 ( .A(n8202), .B(n8203), .Z(n7980) );
  NANDN U8214 ( .A(n8204), .B(n8205), .Z(n8203) );
  OR U8215 ( .A(n8206), .B(n8207), .Z(n8205) );
  NAND U8216 ( .A(n8207), .B(n8206), .Z(n8202) );
  ANDN U8217 ( .B(B[21]), .A(n55), .Z(n7982) );
  XNOR U8218 ( .A(n7990), .B(n8208), .Z(n7983) );
  XNOR U8219 ( .A(n7989), .B(n7987), .Z(n8208) );
  AND U8220 ( .A(n8209), .B(n8210), .Z(n7987) );
  NANDN U8221 ( .A(n8211), .B(n8212), .Z(n8210) );
  NANDN U8222 ( .A(n8213), .B(n8214), .Z(n8212) );
  NANDN U8223 ( .A(n8214), .B(n8213), .Z(n8209) );
  ANDN U8224 ( .B(B[22]), .A(n56), .Z(n7989) );
  XNOR U8225 ( .A(n7997), .B(n8215), .Z(n7990) );
  XNOR U8226 ( .A(n7996), .B(n7994), .Z(n8215) );
  AND U8227 ( .A(n8216), .B(n8217), .Z(n7994) );
  NANDN U8228 ( .A(n8218), .B(n8219), .Z(n8217) );
  OR U8229 ( .A(n8220), .B(n8221), .Z(n8219) );
  NAND U8230 ( .A(n8221), .B(n8220), .Z(n8216) );
  ANDN U8231 ( .B(B[23]), .A(n57), .Z(n7996) );
  XNOR U8232 ( .A(n8004), .B(n8222), .Z(n7997) );
  XNOR U8233 ( .A(n8003), .B(n8001), .Z(n8222) );
  AND U8234 ( .A(n8223), .B(n8224), .Z(n8001) );
  NANDN U8235 ( .A(n8225), .B(n8226), .Z(n8224) );
  NANDN U8236 ( .A(n8227), .B(n8228), .Z(n8226) );
  NANDN U8237 ( .A(n8228), .B(n8227), .Z(n8223) );
  ANDN U8238 ( .B(B[24]), .A(n58), .Z(n8003) );
  XNOR U8239 ( .A(n8011), .B(n8229), .Z(n8004) );
  XNOR U8240 ( .A(n8010), .B(n8008), .Z(n8229) );
  AND U8241 ( .A(n8230), .B(n8231), .Z(n8008) );
  NANDN U8242 ( .A(n8232), .B(n8233), .Z(n8231) );
  OR U8243 ( .A(n8234), .B(n8235), .Z(n8233) );
  NAND U8244 ( .A(n8235), .B(n8234), .Z(n8230) );
  ANDN U8245 ( .B(B[25]), .A(n59), .Z(n8010) );
  XNOR U8246 ( .A(n8018), .B(n8236), .Z(n8011) );
  XNOR U8247 ( .A(n8017), .B(n8015), .Z(n8236) );
  AND U8248 ( .A(n8237), .B(n8238), .Z(n8015) );
  NANDN U8249 ( .A(n8239), .B(n8240), .Z(n8238) );
  NANDN U8250 ( .A(n8241), .B(n8242), .Z(n8240) );
  NANDN U8251 ( .A(n8242), .B(n8241), .Z(n8237) );
  ANDN U8252 ( .B(B[26]), .A(n60), .Z(n8017) );
  XNOR U8253 ( .A(n8025), .B(n8243), .Z(n8018) );
  XNOR U8254 ( .A(n8024), .B(n8022), .Z(n8243) );
  AND U8255 ( .A(n8244), .B(n8245), .Z(n8022) );
  NANDN U8256 ( .A(n8246), .B(n8247), .Z(n8245) );
  OR U8257 ( .A(n8248), .B(n8249), .Z(n8247) );
  NAND U8258 ( .A(n8249), .B(n8248), .Z(n8244) );
  ANDN U8259 ( .B(B[27]), .A(n61), .Z(n8024) );
  XNOR U8260 ( .A(n8032), .B(n8250), .Z(n8025) );
  XNOR U8261 ( .A(n8031), .B(n8029), .Z(n8250) );
  AND U8262 ( .A(n8251), .B(n8252), .Z(n8029) );
  NANDN U8263 ( .A(n8253), .B(n8254), .Z(n8252) );
  NANDN U8264 ( .A(n8255), .B(n8256), .Z(n8254) );
  NANDN U8265 ( .A(n8256), .B(n8255), .Z(n8251) );
  ANDN U8266 ( .B(B[28]), .A(n62), .Z(n8031) );
  XNOR U8267 ( .A(n8039), .B(n8257), .Z(n8032) );
  XNOR U8268 ( .A(n8038), .B(n8036), .Z(n8257) );
  AND U8269 ( .A(n8258), .B(n8259), .Z(n8036) );
  NANDN U8270 ( .A(n8260), .B(n8261), .Z(n8259) );
  OR U8271 ( .A(n8262), .B(n8263), .Z(n8261) );
  NAND U8272 ( .A(n8263), .B(n8262), .Z(n8258) );
  ANDN U8273 ( .B(B[29]), .A(n63), .Z(n8038) );
  XNOR U8274 ( .A(n8046), .B(n8264), .Z(n8039) );
  XNOR U8275 ( .A(n8045), .B(n8043), .Z(n8264) );
  AND U8276 ( .A(n8265), .B(n8266), .Z(n8043) );
  NANDN U8277 ( .A(n8267), .B(n8268), .Z(n8266) );
  NANDN U8278 ( .A(n8269), .B(n8270), .Z(n8268) );
  NANDN U8279 ( .A(n8270), .B(n8269), .Z(n8265) );
  ANDN U8280 ( .B(B[30]), .A(n64), .Z(n8045) );
  XNOR U8281 ( .A(n8053), .B(n8271), .Z(n8046) );
  XNOR U8282 ( .A(n8052), .B(n8050), .Z(n8271) );
  AND U8283 ( .A(n8272), .B(n8273), .Z(n8050) );
  NANDN U8284 ( .A(n8274), .B(n8275), .Z(n8273) );
  OR U8285 ( .A(n8276), .B(n8277), .Z(n8275) );
  NAND U8286 ( .A(n8277), .B(n8276), .Z(n8272) );
  ANDN U8287 ( .B(B[31]), .A(n65), .Z(n8052) );
  XNOR U8288 ( .A(n8060), .B(n8278), .Z(n8053) );
  XNOR U8289 ( .A(n8059), .B(n8057), .Z(n8278) );
  AND U8290 ( .A(n8279), .B(n8280), .Z(n8057) );
  NANDN U8291 ( .A(n8281), .B(n8282), .Z(n8280) );
  NANDN U8292 ( .A(n8283), .B(n8284), .Z(n8282) );
  NANDN U8293 ( .A(n8284), .B(n8283), .Z(n8279) );
  ANDN U8294 ( .B(B[32]), .A(n66), .Z(n8059) );
  XNOR U8295 ( .A(n8067), .B(n8285), .Z(n8060) );
  XNOR U8296 ( .A(n8066), .B(n8064), .Z(n8285) );
  AND U8297 ( .A(n8286), .B(n8287), .Z(n8064) );
  NANDN U8298 ( .A(n8288), .B(n8289), .Z(n8287) );
  OR U8299 ( .A(n8290), .B(n8291), .Z(n8289) );
  NAND U8300 ( .A(n8291), .B(n8290), .Z(n8286) );
  ANDN U8301 ( .B(B[33]), .A(n67), .Z(n8066) );
  XNOR U8302 ( .A(n8074), .B(n8292), .Z(n8067) );
  XNOR U8303 ( .A(n8073), .B(n8071), .Z(n8292) );
  AND U8304 ( .A(n8293), .B(n8294), .Z(n8071) );
  NANDN U8305 ( .A(n8295), .B(n8296), .Z(n8294) );
  NANDN U8306 ( .A(n8297), .B(n8298), .Z(n8296) );
  NANDN U8307 ( .A(n8298), .B(n8297), .Z(n8293) );
  ANDN U8308 ( .B(B[34]), .A(n68), .Z(n8073) );
  XNOR U8309 ( .A(n8081), .B(n8299), .Z(n8074) );
  XNOR U8310 ( .A(n8080), .B(n8078), .Z(n8299) );
  AND U8311 ( .A(n8300), .B(n8301), .Z(n8078) );
  NANDN U8312 ( .A(n8302), .B(n8303), .Z(n8301) );
  OR U8313 ( .A(n8304), .B(n8305), .Z(n8303) );
  NAND U8314 ( .A(n8305), .B(n8304), .Z(n8300) );
  ANDN U8315 ( .B(B[35]), .A(n69), .Z(n8080) );
  XNOR U8316 ( .A(n8088), .B(n8306), .Z(n8081) );
  XNOR U8317 ( .A(n8087), .B(n8085), .Z(n8306) );
  AND U8318 ( .A(n8307), .B(n8308), .Z(n8085) );
  NANDN U8319 ( .A(n8309), .B(n8310), .Z(n8308) );
  NANDN U8320 ( .A(n8311), .B(n8312), .Z(n8310) );
  NANDN U8321 ( .A(n8312), .B(n8311), .Z(n8307) );
  ANDN U8322 ( .B(B[36]), .A(n70), .Z(n8087) );
  XNOR U8323 ( .A(n8095), .B(n8313), .Z(n8088) );
  XNOR U8324 ( .A(n8094), .B(n8092), .Z(n8313) );
  AND U8325 ( .A(n8314), .B(n8315), .Z(n8092) );
  NANDN U8326 ( .A(n8316), .B(n8317), .Z(n8315) );
  OR U8327 ( .A(n8318), .B(n8319), .Z(n8317) );
  NAND U8328 ( .A(n8319), .B(n8318), .Z(n8314) );
  ANDN U8329 ( .B(B[37]), .A(n71), .Z(n8094) );
  XNOR U8330 ( .A(n8102), .B(n8320), .Z(n8095) );
  XNOR U8331 ( .A(n8101), .B(n8099), .Z(n8320) );
  AND U8332 ( .A(n8321), .B(n8322), .Z(n8099) );
  NANDN U8333 ( .A(n8323), .B(n8324), .Z(n8322) );
  NANDN U8334 ( .A(n8325), .B(n8326), .Z(n8324) );
  NANDN U8335 ( .A(n8326), .B(n8325), .Z(n8321) );
  ANDN U8336 ( .B(B[38]), .A(n72), .Z(n8101) );
  XNOR U8337 ( .A(n8109), .B(n8327), .Z(n8102) );
  XNOR U8338 ( .A(n8108), .B(n8106), .Z(n8327) );
  AND U8339 ( .A(n8328), .B(n8329), .Z(n8106) );
  NANDN U8340 ( .A(n8330), .B(n8331), .Z(n8329) );
  OR U8341 ( .A(n8332), .B(n8333), .Z(n8331) );
  NAND U8342 ( .A(n8333), .B(n8332), .Z(n8328) );
  ANDN U8343 ( .B(B[39]), .A(n73), .Z(n8108) );
  XNOR U8344 ( .A(n8116), .B(n8334), .Z(n8109) );
  XNOR U8345 ( .A(n8115), .B(n8113), .Z(n8334) );
  AND U8346 ( .A(n8335), .B(n8336), .Z(n8113) );
  NANDN U8347 ( .A(n8337), .B(n8338), .Z(n8336) );
  NANDN U8348 ( .A(n8339), .B(n8340), .Z(n8338) );
  NANDN U8349 ( .A(n8340), .B(n8339), .Z(n8335) );
  ANDN U8350 ( .B(B[40]), .A(n74), .Z(n8115) );
  XNOR U8351 ( .A(n8123), .B(n8341), .Z(n8116) );
  XNOR U8352 ( .A(n8122), .B(n8120), .Z(n8341) );
  AND U8353 ( .A(n8342), .B(n8343), .Z(n8120) );
  NANDN U8354 ( .A(n8344), .B(n8345), .Z(n8343) );
  OR U8355 ( .A(n8346), .B(n8347), .Z(n8345) );
  NAND U8356 ( .A(n8347), .B(n8346), .Z(n8342) );
  ANDN U8357 ( .B(B[41]), .A(n75), .Z(n8122) );
  XNOR U8358 ( .A(n8130), .B(n8348), .Z(n8123) );
  XNOR U8359 ( .A(n8129), .B(n8127), .Z(n8348) );
  AND U8360 ( .A(n8349), .B(n8350), .Z(n8127) );
  NANDN U8361 ( .A(n8351), .B(n8352), .Z(n8350) );
  NANDN U8362 ( .A(n8353), .B(n8354), .Z(n8352) );
  NANDN U8363 ( .A(n8354), .B(n8353), .Z(n8349) );
  ANDN U8364 ( .B(B[42]), .A(n76), .Z(n8129) );
  XNOR U8365 ( .A(n8137), .B(n8355), .Z(n8130) );
  XNOR U8366 ( .A(n8136), .B(n8134), .Z(n8355) );
  AND U8367 ( .A(n8356), .B(n8357), .Z(n8134) );
  NANDN U8368 ( .A(n8358), .B(n8359), .Z(n8357) );
  OR U8369 ( .A(n8360), .B(n8361), .Z(n8359) );
  NAND U8370 ( .A(n8361), .B(n8360), .Z(n8356) );
  ANDN U8371 ( .B(B[43]), .A(n77), .Z(n8136) );
  XNOR U8372 ( .A(n8144), .B(n8362), .Z(n8137) );
  XNOR U8373 ( .A(n8143), .B(n8141), .Z(n8362) );
  AND U8374 ( .A(n8363), .B(n8364), .Z(n8141) );
  NANDN U8375 ( .A(n8365), .B(n8366), .Z(n8364) );
  NANDN U8376 ( .A(n8367), .B(n8368), .Z(n8366) );
  NANDN U8377 ( .A(n8368), .B(n8367), .Z(n8363) );
  ANDN U8378 ( .B(B[44]), .A(n78), .Z(n8143) );
  XNOR U8379 ( .A(n8151), .B(n8369), .Z(n8144) );
  XNOR U8380 ( .A(n8150), .B(n8148), .Z(n8369) );
  AND U8381 ( .A(n8370), .B(n8371), .Z(n8148) );
  NANDN U8382 ( .A(n8372), .B(n8373), .Z(n8371) );
  OR U8383 ( .A(n8374), .B(n8375), .Z(n8373) );
  NAND U8384 ( .A(n8375), .B(n8374), .Z(n8370) );
  ANDN U8385 ( .B(B[45]), .A(n79), .Z(n8150) );
  XNOR U8386 ( .A(n8158), .B(n8376), .Z(n8151) );
  XNOR U8387 ( .A(n8157), .B(n8155), .Z(n8376) );
  AND U8388 ( .A(n8377), .B(n8378), .Z(n8155) );
  NANDN U8389 ( .A(n8379), .B(n8380), .Z(n8378) );
  NANDN U8390 ( .A(n8381), .B(n8382), .Z(n8380) );
  NANDN U8391 ( .A(n8382), .B(n8381), .Z(n8377) );
  ANDN U8392 ( .B(B[46]), .A(n80), .Z(n8157) );
  XNOR U8393 ( .A(n8165), .B(n8383), .Z(n8158) );
  XNOR U8394 ( .A(n8164), .B(n8162), .Z(n8383) );
  AND U8395 ( .A(n8384), .B(n8385), .Z(n8162) );
  NANDN U8396 ( .A(n8386), .B(n8387), .Z(n8385) );
  OR U8397 ( .A(n8388), .B(n8389), .Z(n8387) );
  NAND U8398 ( .A(n8389), .B(n8388), .Z(n8384) );
  ANDN U8399 ( .B(B[47]), .A(n81), .Z(n8164) );
  XNOR U8400 ( .A(n8172), .B(n8390), .Z(n8165) );
  XNOR U8401 ( .A(n8171), .B(n8169), .Z(n8390) );
  AND U8402 ( .A(n8391), .B(n8392), .Z(n8169) );
  NANDN U8403 ( .A(n8393), .B(n8394), .Z(n8392) );
  NAND U8404 ( .A(n8395), .B(n8396), .Z(n8394) );
  ANDN U8405 ( .B(B[48]), .A(n82), .Z(n8171) );
  XOR U8406 ( .A(n8178), .B(n8397), .Z(n8172) );
  XNOR U8407 ( .A(n8176), .B(n8179), .Z(n8397) );
  NAND U8408 ( .A(A[2]), .B(B[49]), .Z(n8179) );
  NANDN U8409 ( .A(n8398), .B(n8399), .Z(n8176) );
  AND U8410 ( .A(A[0]), .B(B[50]), .Z(n8399) );
  XNOR U8411 ( .A(n8181), .B(n8400), .Z(n8178) );
  NAND U8412 ( .A(A[0]), .B(B[51]), .Z(n8400) );
  NAND U8413 ( .A(B[50]), .B(A[1]), .Z(n8181) );
  NAND U8414 ( .A(n8401), .B(n8402), .Z(n185) );
  NANDN U8415 ( .A(n8403), .B(n8404), .Z(n8402) );
  OR U8416 ( .A(n8405), .B(n8406), .Z(n8404) );
  NAND U8417 ( .A(n8406), .B(n8405), .Z(n8401) );
  XOR U8418 ( .A(n187), .B(n186), .Z(\A1[48] ) );
  XOR U8419 ( .A(n8406), .B(n8407), .Z(n186) );
  XNOR U8420 ( .A(n8405), .B(n8403), .Z(n8407) );
  AND U8421 ( .A(n8408), .B(n8409), .Z(n8403) );
  NANDN U8422 ( .A(n8410), .B(n8411), .Z(n8409) );
  NANDN U8423 ( .A(n8412), .B(n8413), .Z(n8411) );
  NANDN U8424 ( .A(n8413), .B(n8412), .Z(n8408) );
  ANDN U8425 ( .B(B[19]), .A(n54), .Z(n8405) );
  XNOR U8426 ( .A(n8200), .B(n8414), .Z(n8406) );
  XNOR U8427 ( .A(n8199), .B(n8197), .Z(n8414) );
  AND U8428 ( .A(n8415), .B(n8416), .Z(n8197) );
  NANDN U8429 ( .A(n8417), .B(n8418), .Z(n8416) );
  OR U8430 ( .A(n8419), .B(n8420), .Z(n8418) );
  NAND U8431 ( .A(n8420), .B(n8419), .Z(n8415) );
  ANDN U8432 ( .B(B[20]), .A(n55), .Z(n8199) );
  XNOR U8433 ( .A(n8207), .B(n8421), .Z(n8200) );
  XNOR U8434 ( .A(n8206), .B(n8204), .Z(n8421) );
  AND U8435 ( .A(n8422), .B(n8423), .Z(n8204) );
  NANDN U8436 ( .A(n8424), .B(n8425), .Z(n8423) );
  NANDN U8437 ( .A(n8426), .B(n8427), .Z(n8425) );
  NANDN U8438 ( .A(n8427), .B(n8426), .Z(n8422) );
  ANDN U8439 ( .B(B[21]), .A(n56), .Z(n8206) );
  XNOR U8440 ( .A(n8214), .B(n8428), .Z(n8207) );
  XNOR U8441 ( .A(n8213), .B(n8211), .Z(n8428) );
  AND U8442 ( .A(n8429), .B(n8430), .Z(n8211) );
  NANDN U8443 ( .A(n8431), .B(n8432), .Z(n8430) );
  OR U8444 ( .A(n8433), .B(n8434), .Z(n8432) );
  NAND U8445 ( .A(n8434), .B(n8433), .Z(n8429) );
  ANDN U8446 ( .B(B[22]), .A(n57), .Z(n8213) );
  XNOR U8447 ( .A(n8221), .B(n8435), .Z(n8214) );
  XNOR U8448 ( .A(n8220), .B(n8218), .Z(n8435) );
  AND U8449 ( .A(n8436), .B(n8437), .Z(n8218) );
  NANDN U8450 ( .A(n8438), .B(n8439), .Z(n8437) );
  NANDN U8451 ( .A(n8440), .B(n8441), .Z(n8439) );
  NANDN U8452 ( .A(n8441), .B(n8440), .Z(n8436) );
  ANDN U8453 ( .B(B[23]), .A(n58), .Z(n8220) );
  XNOR U8454 ( .A(n8228), .B(n8442), .Z(n8221) );
  XNOR U8455 ( .A(n8227), .B(n8225), .Z(n8442) );
  AND U8456 ( .A(n8443), .B(n8444), .Z(n8225) );
  NANDN U8457 ( .A(n8445), .B(n8446), .Z(n8444) );
  OR U8458 ( .A(n8447), .B(n8448), .Z(n8446) );
  NAND U8459 ( .A(n8448), .B(n8447), .Z(n8443) );
  ANDN U8460 ( .B(B[24]), .A(n59), .Z(n8227) );
  XNOR U8461 ( .A(n8235), .B(n8449), .Z(n8228) );
  XNOR U8462 ( .A(n8234), .B(n8232), .Z(n8449) );
  AND U8463 ( .A(n8450), .B(n8451), .Z(n8232) );
  NANDN U8464 ( .A(n8452), .B(n8453), .Z(n8451) );
  NANDN U8465 ( .A(n8454), .B(n8455), .Z(n8453) );
  NANDN U8466 ( .A(n8455), .B(n8454), .Z(n8450) );
  ANDN U8467 ( .B(B[25]), .A(n60), .Z(n8234) );
  XNOR U8468 ( .A(n8242), .B(n8456), .Z(n8235) );
  XNOR U8469 ( .A(n8241), .B(n8239), .Z(n8456) );
  AND U8470 ( .A(n8457), .B(n8458), .Z(n8239) );
  NANDN U8471 ( .A(n8459), .B(n8460), .Z(n8458) );
  OR U8472 ( .A(n8461), .B(n8462), .Z(n8460) );
  NAND U8473 ( .A(n8462), .B(n8461), .Z(n8457) );
  ANDN U8474 ( .B(B[26]), .A(n61), .Z(n8241) );
  XNOR U8475 ( .A(n8249), .B(n8463), .Z(n8242) );
  XNOR U8476 ( .A(n8248), .B(n8246), .Z(n8463) );
  AND U8477 ( .A(n8464), .B(n8465), .Z(n8246) );
  NANDN U8478 ( .A(n8466), .B(n8467), .Z(n8465) );
  NANDN U8479 ( .A(n8468), .B(n8469), .Z(n8467) );
  NANDN U8480 ( .A(n8469), .B(n8468), .Z(n8464) );
  ANDN U8481 ( .B(B[27]), .A(n62), .Z(n8248) );
  XNOR U8482 ( .A(n8256), .B(n8470), .Z(n8249) );
  XNOR U8483 ( .A(n8255), .B(n8253), .Z(n8470) );
  AND U8484 ( .A(n8471), .B(n8472), .Z(n8253) );
  NANDN U8485 ( .A(n8473), .B(n8474), .Z(n8472) );
  OR U8486 ( .A(n8475), .B(n8476), .Z(n8474) );
  NAND U8487 ( .A(n8476), .B(n8475), .Z(n8471) );
  ANDN U8488 ( .B(B[28]), .A(n63), .Z(n8255) );
  XNOR U8489 ( .A(n8263), .B(n8477), .Z(n8256) );
  XNOR U8490 ( .A(n8262), .B(n8260), .Z(n8477) );
  AND U8491 ( .A(n8478), .B(n8479), .Z(n8260) );
  NANDN U8492 ( .A(n8480), .B(n8481), .Z(n8479) );
  NANDN U8493 ( .A(n8482), .B(n8483), .Z(n8481) );
  NANDN U8494 ( .A(n8483), .B(n8482), .Z(n8478) );
  ANDN U8495 ( .B(B[29]), .A(n64), .Z(n8262) );
  XNOR U8496 ( .A(n8270), .B(n8484), .Z(n8263) );
  XNOR U8497 ( .A(n8269), .B(n8267), .Z(n8484) );
  AND U8498 ( .A(n8485), .B(n8486), .Z(n8267) );
  NANDN U8499 ( .A(n8487), .B(n8488), .Z(n8486) );
  OR U8500 ( .A(n8489), .B(n8490), .Z(n8488) );
  NAND U8501 ( .A(n8490), .B(n8489), .Z(n8485) );
  ANDN U8502 ( .B(B[30]), .A(n65), .Z(n8269) );
  XNOR U8503 ( .A(n8277), .B(n8491), .Z(n8270) );
  XNOR U8504 ( .A(n8276), .B(n8274), .Z(n8491) );
  AND U8505 ( .A(n8492), .B(n8493), .Z(n8274) );
  NANDN U8506 ( .A(n8494), .B(n8495), .Z(n8493) );
  NANDN U8507 ( .A(n8496), .B(n8497), .Z(n8495) );
  NANDN U8508 ( .A(n8497), .B(n8496), .Z(n8492) );
  ANDN U8509 ( .B(B[31]), .A(n66), .Z(n8276) );
  XNOR U8510 ( .A(n8284), .B(n8498), .Z(n8277) );
  XNOR U8511 ( .A(n8283), .B(n8281), .Z(n8498) );
  AND U8512 ( .A(n8499), .B(n8500), .Z(n8281) );
  NANDN U8513 ( .A(n8501), .B(n8502), .Z(n8500) );
  OR U8514 ( .A(n8503), .B(n8504), .Z(n8502) );
  NAND U8515 ( .A(n8504), .B(n8503), .Z(n8499) );
  ANDN U8516 ( .B(B[32]), .A(n67), .Z(n8283) );
  XNOR U8517 ( .A(n8291), .B(n8505), .Z(n8284) );
  XNOR U8518 ( .A(n8290), .B(n8288), .Z(n8505) );
  AND U8519 ( .A(n8506), .B(n8507), .Z(n8288) );
  NANDN U8520 ( .A(n8508), .B(n8509), .Z(n8507) );
  NANDN U8521 ( .A(n8510), .B(n8511), .Z(n8509) );
  NANDN U8522 ( .A(n8511), .B(n8510), .Z(n8506) );
  ANDN U8523 ( .B(B[33]), .A(n68), .Z(n8290) );
  XNOR U8524 ( .A(n8298), .B(n8512), .Z(n8291) );
  XNOR U8525 ( .A(n8297), .B(n8295), .Z(n8512) );
  AND U8526 ( .A(n8513), .B(n8514), .Z(n8295) );
  NANDN U8527 ( .A(n8515), .B(n8516), .Z(n8514) );
  OR U8528 ( .A(n8517), .B(n8518), .Z(n8516) );
  NAND U8529 ( .A(n8518), .B(n8517), .Z(n8513) );
  ANDN U8530 ( .B(B[34]), .A(n69), .Z(n8297) );
  XNOR U8531 ( .A(n8305), .B(n8519), .Z(n8298) );
  XNOR U8532 ( .A(n8304), .B(n8302), .Z(n8519) );
  AND U8533 ( .A(n8520), .B(n8521), .Z(n8302) );
  NANDN U8534 ( .A(n8522), .B(n8523), .Z(n8521) );
  NANDN U8535 ( .A(n8524), .B(n8525), .Z(n8523) );
  NANDN U8536 ( .A(n8525), .B(n8524), .Z(n8520) );
  ANDN U8537 ( .B(B[35]), .A(n70), .Z(n8304) );
  XNOR U8538 ( .A(n8312), .B(n8526), .Z(n8305) );
  XNOR U8539 ( .A(n8311), .B(n8309), .Z(n8526) );
  AND U8540 ( .A(n8527), .B(n8528), .Z(n8309) );
  NANDN U8541 ( .A(n8529), .B(n8530), .Z(n8528) );
  OR U8542 ( .A(n8531), .B(n8532), .Z(n8530) );
  NAND U8543 ( .A(n8532), .B(n8531), .Z(n8527) );
  ANDN U8544 ( .B(B[36]), .A(n71), .Z(n8311) );
  XNOR U8545 ( .A(n8319), .B(n8533), .Z(n8312) );
  XNOR U8546 ( .A(n8318), .B(n8316), .Z(n8533) );
  AND U8547 ( .A(n8534), .B(n8535), .Z(n8316) );
  NANDN U8548 ( .A(n8536), .B(n8537), .Z(n8535) );
  NANDN U8549 ( .A(n8538), .B(n8539), .Z(n8537) );
  NANDN U8550 ( .A(n8539), .B(n8538), .Z(n8534) );
  ANDN U8551 ( .B(B[37]), .A(n72), .Z(n8318) );
  XNOR U8552 ( .A(n8326), .B(n8540), .Z(n8319) );
  XNOR U8553 ( .A(n8325), .B(n8323), .Z(n8540) );
  AND U8554 ( .A(n8541), .B(n8542), .Z(n8323) );
  NANDN U8555 ( .A(n8543), .B(n8544), .Z(n8542) );
  OR U8556 ( .A(n8545), .B(n8546), .Z(n8544) );
  NAND U8557 ( .A(n8546), .B(n8545), .Z(n8541) );
  ANDN U8558 ( .B(B[38]), .A(n73), .Z(n8325) );
  XNOR U8559 ( .A(n8333), .B(n8547), .Z(n8326) );
  XNOR U8560 ( .A(n8332), .B(n8330), .Z(n8547) );
  AND U8561 ( .A(n8548), .B(n8549), .Z(n8330) );
  NANDN U8562 ( .A(n8550), .B(n8551), .Z(n8549) );
  NANDN U8563 ( .A(n8552), .B(n8553), .Z(n8551) );
  NANDN U8564 ( .A(n8553), .B(n8552), .Z(n8548) );
  ANDN U8565 ( .B(B[39]), .A(n74), .Z(n8332) );
  XNOR U8566 ( .A(n8340), .B(n8554), .Z(n8333) );
  XNOR U8567 ( .A(n8339), .B(n8337), .Z(n8554) );
  AND U8568 ( .A(n8555), .B(n8556), .Z(n8337) );
  NANDN U8569 ( .A(n8557), .B(n8558), .Z(n8556) );
  OR U8570 ( .A(n8559), .B(n8560), .Z(n8558) );
  NAND U8571 ( .A(n8560), .B(n8559), .Z(n8555) );
  ANDN U8572 ( .B(B[40]), .A(n75), .Z(n8339) );
  XNOR U8573 ( .A(n8347), .B(n8561), .Z(n8340) );
  XNOR U8574 ( .A(n8346), .B(n8344), .Z(n8561) );
  AND U8575 ( .A(n8562), .B(n8563), .Z(n8344) );
  NANDN U8576 ( .A(n8564), .B(n8565), .Z(n8563) );
  NANDN U8577 ( .A(n8566), .B(n8567), .Z(n8565) );
  NANDN U8578 ( .A(n8567), .B(n8566), .Z(n8562) );
  ANDN U8579 ( .B(B[41]), .A(n76), .Z(n8346) );
  XNOR U8580 ( .A(n8354), .B(n8568), .Z(n8347) );
  XNOR U8581 ( .A(n8353), .B(n8351), .Z(n8568) );
  AND U8582 ( .A(n8569), .B(n8570), .Z(n8351) );
  NANDN U8583 ( .A(n8571), .B(n8572), .Z(n8570) );
  OR U8584 ( .A(n8573), .B(n8574), .Z(n8572) );
  NAND U8585 ( .A(n8574), .B(n8573), .Z(n8569) );
  ANDN U8586 ( .B(B[42]), .A(n77), .Z(n8353) );
  XNOR U8587 ( .A(n8361), .B(n8575), .Z(n8354) );
  XNOR U8588 ( .A(n8360), .B(n8358), .Z(n8575) );
  AND U8589 ( .A(n8576), .B(n8577), .Z(n8358) );
  NANDN U8590 ( .A(n8578), .B(n8579), .Z(n8577) );
  NANDN U8591 ( .A(n8580), .B(n8581), .Z(n8579) );
  NANDN U8592 ( .A(n8581), .B(n8580), .Z(n8576) );
  ANDN U8593 ( .B(B[43]), .A(n78), .Z(n8360) );
  XNOR U8594 ( .A(n8368), .B(n8582), .Z(n8361) );
  XNOR U8595 ( .A(n8367), .B(n8365), .Z(n8582) );
  AND U8596 ( .A(n8583), .B(n8584), .Z(n8365) );
  NANDN U8597 ( .A(n8585), .B(n8586), .Z(n8584) );
  OR U8598 ( .A(n8587), .B(n8588), .Z(n8586) );
  NAND U8599 ( .A(n8588), .B(n8587), .Z(n8583) );
  ANDN U8600 ( .B(B[44]), .A(n79), .Z(n8367) );
  XNOR U8601 ( .A(n8375), .B(n8589), .Z(n8368) );
  XNOR U8602 ( .A(n8374), .B(n8372), .Z(n8589) );
  AND U8603 ( .A(n8590), .B(n8591), .Z(n8372) );
  NANDN U8604 ( .A(n8592), .B(n8593), .Z(n8591) );
  NANDN U8605 ( .A(n8594), .B(n8595), .Z(n8593) );
  NANDN U8606 ( .A(n8595), .B(n8594), .Z(n8590) );
  ANDN U8607 ( .B(B[45]), .A(n80), .Z(n8374) );
  XNOR U8608 ( .A(n8382), .B(n8596), .Z(n8375) );
  XNOR U8609 ( .A(n8381), .B(n8379), .Z(n8596) );
  AND U8610 ( .A(n8597), .B(n8598), .Z(n8379) );
  NANDN U8611 ( .A(n8599), .B(n8600), .Z(n8598) );
  OR U8612 ( .A(n8601), .B(n8602), .Z(n8600) );
  NAND U8613 ( .A(n8602), .B(n8601), .Z(n8597) );
  ANDN U8614 ( .B(B[46]), .A(n81), .Z(n8381) );
  XNOR U8615 ( .A(n8389), .B(n8603), .Z(n8382) );
  XNOR U8616 ( .A(n8388), .B(n8386), .Z(n8603) );
  AND U8617 ( .A(n8604), .B(n8605), .Z(n8386) );
  NANDN U8618 ( .A(n8606), .B(n8607), .Z(n8605) );
  NAND U8619 ( .A(n8608), .B(n8609), .Z(n8607) );
  ANDN U8620 ( .B(B[47]), .A(n82), .Z(n8388) );
  XOR U8621 ( .A(n8395), .B(n8610), .Z(n8389) );
  XNOR U8622 ( .A(n8393), .B(n8396), .Z(n8610) );
  NAND U8623 ( .A(A[2]), .B(B[48]), .Z(n8396) );
  NANDN U8624 ( .A(n8611), .B(n8612), .Z(n8393) );
  AND U8625 ( .A(A[0]), .B(B[49]), .Z(n8612) );
  XNOR U8626 ( .A(n8398), .B(n8613), .Z(n8395) );
  NAND U8627 ( .A(A[0]), .B(B[50]), .Z(n8613) );
  NAND U8628 ( .A(B[49]), .B(A[1]), .Z(n8398) );
  NAND U8629 ( .A(n8614), .B(n8615), .Z(n187) );
  NANDN U8630 ( .A(n8616), .B(n8617), .Z(n8615) );
  OR U8631 ( .A(n8618), .B(n8619), .Z(n8617) );
  NAND U8632 ( .A(n8619), .B(n8618), .Z(n8614) );
  XOR U8633 ( .A(n189), .B(n188), .Z(\A1[47] ) );
  XOR U8634 ( .A(n8619), .B(n8620), .Z(n188) );
  XNOR U8635 ( .A(n8618), .B(n8616), .Z(n8620) );
  AND U8636 ( .A(n8621), .B(n8622), .Z(n8616) );
  NANDN U8637 ( .A(n8623), .B(n8624), .Z(n8622) );
  NANDN U8638 ( .A(n8625), .B(n8626), .Z(n8624) );
  NANDN U8639 ( .A(n8626), .B(n8625), .Z(n8621) );
  ANDN U8640 ( .B(B[18]), .A(n54), .Z(n8618) );
  XNOR U8641 ( .A(n8413), .B(n8627), .Z(n8619) );
  XNOR U8642 ( .A(n8412), .B(n8410), .Z(n8627) );
  AND U8643 ( .A(n8628), .B(n8629), .Z(n8410) );
  NANDN U8644 ( .A(n8630), .B(n8631), .Z(n8629) );
  OR U8645 ( .A(n8632), .B(n8633), .Z(n8631) );
  NAND U8646 ( .A(n8633), .B(n8632), .Z(n8628) );
  ANDN U8647 ( .B(B[19]), .A(n55), .Z(n8412) );
  XNOR U8648 ( .A(n8420), .B(n8634), .Z(n8413) );
  XNOR U8649 ( .A(n8419), .B(n8417), .Z(n8634) );
  AND U8650 ( .A(n8635), .B(n8636), .Z(n8417) );
  NANDN U8651 ( .A(n8637), .B(n8638), .Z(n8636) );
  NANDN U8652 ( .A(n8639), .B(n8640), .Z(n8638) );
  NANDN U8653 ( .A(n8640), .B(n8639), .Z(n8635) );
  ANDN U8654 ( .B(B[20]), .A(n56), .Z(n8419) );
  XNOR U8655 ( .A(n8427), .B(n8641), .Z(n8420) );
  XNOR U8656 ( .A(n8426), .B(n8424), .Z(n8641) );
  AND U8657 ( .A(n8642), .B(n8643), .Z(n8424) );
  NANDN U8658 ( .A(n8644), .B(n8645), .Z(n8643) );
  OR U8659 ( .A(n8646), .B(n8647), .Z(n8645) );
  NAND U8660 ( .A(n8647), .B(n8646), .Z(n8642) );
  ANDN U8661 ( .B(B[21]), .A(n57), .Z(n8426) );
  XNOR U8662 ( .A(n8434), .B(n8648), .Z(n8427) );
  XNOR U8663 ( .A(n8433), .B(n8431), .Z(n8648) );
  AND U8664 ( .A(n8649), .B(n8650), .Z(n8431) );
  NANDN U8665 ( .A(n8651), .B(n8652), .Z(n8650) );
  NANDN U8666 ( .A(n8653), .B(n8654), .Z(n8652) );
  NANDN U8667 ( .A(n8654), .B(n8653), .Z(n8649) );
  ANDN U8668 ( .B(B[22]), .A(n58), .Z(n8433) );
  XNOR U8669 ( .A(n8441), .B(n8655), .Z(n8434) );
  XNOR U8670 ( .A(n8440), .B(n8438), .Z(n8655) );
  AND U8671 ( .A(n8656), .B(n8657), .Z(n8438) );
  NANDN U8672 ( .A(n8658), .B(n8659), .Z(n8657) );
  OR U8673 ( .A(n8660), .B(n8661), .Z(n8659) );
  NAND U8674 ( .A(n8661), .B(n8660), .Z(n8656) );
  ANDN U8675 ( .B(B[23]), .A(n59), .Z(n8440) );
  XNOR U8676 ( .A(n8448), .B(n8662), .Z(n8441) );
  XNOR U8677 ( .A(n8447), .B(n8445), .Z(n8662) );
  AND U8678 ( .A(n8663), .B(n8664), .Z(n8445) );
  NANDN U8679 ( .A(n8665), .B(n8666), .Z(n8664) );
  NANDN U8680 ( .A(n8667), .B(n8668), .Z(n8666) );
  NANDN U8681 ( .A(n8668), .B(n8667), .Z(n8663) );
  ANDN U8682 ( .B(B[24]), .A(n60), .Z(n8447) );
  XNOR U8683 ( .A(n8455), .B(n8669), .Z(n8448) );
  XNOR U8684 ( .A(n8454), .B(n8452), .Z(n8669) );
  AND U8685 ( .A(n8670), .B(n8671), .Z(n8452) );
  NANDN U8686 ( .A(n8672), .B(n8673), .Z(n8671) );
  OR U8687 ( .A(n8674), .B(n8675), .Z(n8673) );
  NAND U8688 ( .A(n8675), .B(n8674), .Z(n8670) );
  ANDN U8689 ( .B(B[25]), .A(n61), .Z(n8454) );
  XNOR U8690 ( .A(n8462), .B(n8676), .Z(n8455) );
  XNOR U8691 ( .A(n8461), .B(n8459), .Z(n8676) );
  AND U8692 ( .A(n8677), .B(n8678), .Z(n8459) );
  NANDN U8693 ( .A(n8679), .B(n8680), .Z(n8678) );
  NANDN U8694 ( .A(n8681), .B(n8682), .Z(n8680) );
  NANDN U8695 ( .A(n8682), .B(n8681), .Z(n8677) );
  ANDN U8696 ( .B(B[26]), .A(n62), .Z(n8461) );
  XNOR U8697 ( .A(n8469), .B(n8683), .Z(n8462) );
  XNOR U8698 ( .A(n8468), .B(n8466), .Z(n8683) );
  AND U8699 ( .A(n8684), .B(n8685), .Z(n8466) );
  NANDN U8700 ( .A(n8686), .B(n8687), .Z(n8685) );
  OR U8701 ( .A(n8688), .B(n8689), .Z(n8687) );
  NAND U8702 ( .A(n8689), .B(n8688), .Z(n8684) );
  ANDN U8703 ( .B(B[27]), .A(n63), .Z(n8468) );
  XNOR U8704 ( .A(n8476), .B(n8690), .Z(n8469) );
  XNOR U8705 ( .A(n8475), .B(n8473), .Z(n8690) );
  AND U8706 ( .A(n8691), .B(n8692), .Z(n8473) );
  NANDN U8707 ( .A(n8693), .B(n8694), .Z(n8692) );
  NANDN U8708 ( .A(n8695), .B(n8696), .Z(n8694) );
  NANDN U8709 ( .A(n8696), .B(n8695), .Z(n8691) );
  ANDN U8710 ( .B(B[28]), .A(n64), .Z(n8475) );
  XNOR U8711 ( .A(n8483), .B(n8697), .Z(n8476) );
  XNOR U8712 ( .A(n8482), .B(n8480), .Z(n8697) );
  AND U8713 ( .A(n8698), .B(n8699), .Z(n8480) );
  NANDN U8714 ( .A(n8700), .B(n8701), .Z(n8699) );
  OR U8715 ( .A(n8702), .B(n8703), .Z(n8701) );
  NAND U8716 ( .A(n8703), .B(n8702), .Z(n8698) );
  ANDN U8717 ( .B(B[29]), .A(n65), .Z(n8482) );
  XNOR U8718 ( .A(n8490), .B(n8704), .Z(n8483) );
  XNOR U8719 ( .A(n8489), .B(n8487), .Z(n8704) );
  AND U8720 ( .A(n8705), .B(n8706), .Z(n8487) );
  NANDN U8721 ( .A(n8707), .B(n8708), .Z(n8706) );
  NANDN U8722 ( .A(n8709), .B(n8710), .Z(n8708) );
  NANDN U8723 ( .A(n8710), .B(n8709), .Z(n8705) );
  ANDN U8724 ( .B(B[30]), .A(n66), .Z(n8489) );
  XNOR U8725 ( .A(n8497), .B(n8711), .Z(n8490) );
  XNOR U8726 ( .A(n8496), .B(n8494), .Z(n8711) );
  AND U8727 ( .A(n8712), .B(n8713), .Z(n8494) );
  NANDN U8728 ( .A(n8714), .B(n8715), .Z(n8713) );
  OR U8729 ( .A(n8716), .B(n8717), .Z(n8715) );
  NAND U8730 ( .A(n8717), .B(n8716), .Z(n8712) );
  ANDN U8731 ( .B(B[31]), .A(n67), .Z(n8496) );
  XNOR U8732 ( .A(n8504), .B(n8718), .Z(n8497) );
  XNOR U8733 ( .A(n8503), .B(n8501), .Z(n8718) );
  AND U8734 ( .A(n8719), .B(n8720), .Z(n8501) );
  NANDN U8735 ( .A(n8721), .B(n8722), .Z(n8720) );
  NANDN U8736 ( .A(n8723), .B(n8724), .Z(n8722) );
  NANDN U8737 ( .A(n8724), .B(n8723), .Z(n8719) );
  ANDN U8738 ( .B(B[32]), .A(n68), .Z(n8503) );
  XNOR U8739 ( .A(n8511), .B(n8725), .Z(n8504) );
  XNOR U8740 ( .A(n8510), .B(n8508), .Z(n8725) );
  AND U8741 ( .A(n8726), .B(n8727), .Z(n8508) );
  NANDN U8742 ( .A(n8728), .B(n8729), .Z(n8727) );
  OR U8743 ( .A(n8730), .B(n8731), .Z(n8729) );
  NAND U8744 ( .A(n8731), .B(n8730), .Z(n8726) );
  ANDN U8745 ( .B(B[33]), .A(n69), .Z(n8510) );
  XNOR U8746 ( .A(n8518), .B(n8732), .Z(n8511) );
  XNOR U8747 ( .A(n8517), .B(n8515), .Z(n8732) );
  AND U8748 ( .A(n8733), .B(n8734), .Z(n8515) );
  NANDN U8749 ( .A(n8735), .B(n8736), .Z(n8734) );
  NANDN U8750 ( .A(n8737), .B(n8738), .Z(n8736) );
  NANDN U8751 ( .A(n8738), .B(n8737), .Z(n8733) );
  ANDN U8752 ( .B(B[34]), .A(n70), .Z(n8517) );
  XNOR U8753 ( .A(n8525), .B(n8739), .Z(n8518) );
  XNOR U8754 ( .A(n8524), .B(n8522), .Z(n8739) );
  AND U8755 ( .A(n8740), .B(n8741), .Z(n8522) );
  NANDN U8756 ( .A(n8742), .B(n8743), .Z(n8741) );
  OR U8757 ( .A(n8744), .B(n8745), .Z(n8743) );
  NAND U8758 ( .A(n8745), .B(n8744), .Z(n8740) );
  ANDN U8759 ( .B(B[35]), .A(n71), .Z(n8524) );
  XNOR U8760 ( .A(n8532), .B(n8746), .Z(n8525) );
  XNOR U8761 ( .A(n8531), .B(n8529), .Z(n8746) );
  AND U8762 ( .A(n8747), .B(n8748), .Z(n8529) );
  NANDN U8763 ( .A(n8749), .B(n8750), .Z(n8748) );
  NANDN U8764 ( .A(n8751), .B(n8752), .Z(n8750) );
  NANDN U8765 ( .A(n8752), .B(n8751), .Z(n8747) );
  ANDN U8766 ( .B(B[36]), .A(n72), .Z(n8531) );
  XNOR U8767 ( .A(n8539), .B(n8753), .Z(n8532) );
  XNOR U8768 ( .A(n8538), .B(n8536), .Z(n8753) );
  AND U8769 ( .A(n8754), .B(n8755), .Z(n8536) );
  NANDN U8770 ( .A(n8756), .B(n8757), .Z(n8755) );
  OR U8771 ( .A(n8758), .B(n8759), .Z(n8757) );
  NAND U8772 ( .A(n8759), .B(n8758), .Z(n8754) );
  ANDN U8773 ( .B(B[37]), .A(n73), .Z(n8538) );
  XNOR U8774 ( .A(n8546), .B(n8760), .Z(n8539) );
  XNOR U8775 ( .A(n8545), .B(n8543), .Z(n8760) );
  AND U8776 ( .A(n8761), .B(n8762), .Z(n8543) );
  NANDN U8777 ( .A(n8763), .B(n8764), .Z(n8762) );
  NANDN U8778 ( .A(n8765), .B(n8766), .Z(n8764) );
  NANDN U8779 ( .A(n8766), .B(n8765), .Z(n8761) );
  ANDN U8780 ( .B(B[38]), .A(n74), .Z(n8545) );
  XNOR U8781 ( .A(n8553), .B(n8767), .Z(n8546) );
  XNOR U8782 ( .A(n8552), .B(n8550), .Z(n8767) );
  AND U8783 ( .A(n8768), .B(n8769), .Z(n8550) );
  NANDN U8784 ( .A(n8770), .B(n8771), .Z(n8769) );
  OR U8785 ( .A(n8772), .B(n8773), .Z(n8771) );
  NAND U8786 ( .A(n8773), .B(n8772), .Z(n8768) );
  ANDN U8787 ( .B(B[39]), .A(n75), .Z(n8552) );
  XNOR U8788 ( .A(n8560), .B(n8774), .Z(n8553) );
  XNOR U8789 ( .A(n8559), .B(n8557), .Z(n8774) );
  AND U8790 ( .A(n8775), .B(n8776), .Z(n8557) );
  NANDN U8791 ( .A(n8777), .B(n8778), .Z(n8776) );
  NANDN U8792 ( .A(n8779), .B(n8780), .Z(n8778) );
  NANDN U8793 ( .A(n8780), .B(n8779), .Z(n8775) );
  ANDN U8794 ( .B(B[40]), .A(n76), .Z(n8559) );
  XNOR U8795 ( .A(n8567), .B(n8781), .Z(n8560) );
  XNOR U8796 ( .A(n8566), .B(n8564), .Z(n8781) );
  AND U8797 ( .A(n8782), .B(n8783), .Z(n8564) );
  NANDN U8798 ( .A(n8784), .B(n8785), .Z(n8783) );
  OR U8799 ( .A(n8786), .B(n8787), .Z(n8785) );
  NAND U8800 ( .A(n8787), .B(n8786), .Z(n8782) );
  ANDN U8801 ( .B(B[41]), .A(n77), .Z(n8566) );
  XNOR U8802 ( .A(n8574), .B(n8788), .Z(n8567) );
  XNOR U8803 ( .A(n8573), .B(n8571), .Z(n8788) );
  AND U8804 ( .A(n8789), .B(n8790), .Z(n8571) );
  NANDN U8805 ( .A(n8791), .B(n8792), .Z(n8790) );
  NANDN U8806 ( .A(n8793), .B(n8794), .Z(n8792) );
  NANDN U8807 ( .A(n8794), .B(n8793), .Z(n8789) );
  ANDN U8808 ( .B(B[42]), .A(n78), .Z(n8573) );
  XNOR U8809 ( .A(n8581), .B(n8795), .Z(n8574) );
  XNOR U8810 ( .A(n8580), .B(n8578), .Z(n8795) );
  AND U8811 ( .A(n8796), .B(n8797), .Z(n8578) );
  NANDN U8812 ( .A(n8798), .B(n8799), .Z(n8797) );
  OR U8813 ( .A(n8800), .B(n8801), .Z(n8799) );
  NAND U8814 ( .A(n8801), .B(n8800), .Z(n8796) );
  ANDN U8815 ( .B(B[43]), .A(n79), .Z(n8580) );
  XNOR U8816 ( .A(n8588), .B(n8802), .Z(n8581) );
  XNOR U8817 ( .A(n8587), .B(n8585), .Z(n8802) );
  AND U8818 ( .A(n8803), .B(n8804), .Z(n8585) );
  NANDN U8819 ( .A(n8805), .B(n8806), .Z(n8804) );
  NANDN U8820 ( .A(n8807), .B(n8808), .Z(n8806) );
  NANDN U8821 ( .A(n8808), .B(n8807), .Z(n8803) );
  ANDN U8822 ( .B(B[44]), .A(n80), .Z(n8587) );
  XNOR U8823 ( .A(n8595), .B(n8809), .Z(n8588) );
  XNOR U8824 ( .A(n8594), .B(n8592), .Z(n8809) );
  AND U8825 ( .A(n8810), .B(n8811), .Z(n8592) );
  NANDN U8826 ( .A(n8812), .B(n8813), .Z(n8811) );
  OR U8827 ( .A(n8814), .B(n8815), .Z(n8813) );
  NAND U8828 ( .A(n8815), .B(n8814), .Z(n8810) );
  ANDN U8829 ( .B(B[45]), .A(n81), .Z(n8594) );
  XNOR U8830 ( .A(n8602), .B(n8816), .Z(n8595) );
  XNOR U8831 ( .A(n8601), .B(n8599), .Z(n8816) );
  AND U8832 ( .A(n8817), .B(n8818), .Z(n8599) );
  NANDN U8833 ( .A(n8819), .B(n8820), .Z(n8818) );
  NAND U8834 ( .A(n8821), .B(n8822), .Z(n8820) );
  ANDN U8835 ( .B(B[46]), .A(n82), .Z(n8601) );
  XOR U8836 ( .A(n8608), .B(n8823), .Z(n8602) );
  XNOR U8837 ( .A(n8606), .B(n8609), .Z(n8823) );
  NAND U8838 ( .A(A[2]), .B(B[47]), .Z(n8609) );
  NANDN U8839 ( .A(n8824), .B(n8825), .Z(n8606) );
  AND U8840 ( .A(A[0]), .B(B[48]), .Z(n8825) );
  XNOR U8841 ( .A(n8611), .B(n8826), .Z(n8608) );
  NAND U8842 ( .A(A[0]), .B(B[49]), .Z(n8826) );
  NAND U8843 ( .A(B[48]), .B(A[1]), .Z(n8611) );
  NAND U8844 ( .A(n8827), .B(n8828), .Z(n189) );
  NANDN U8845 ( .A(n8829), .B(n8830), .Z(n8828) );
  OR U8846 ( .A(n8831), .B(n8832), .Z(n8830) );
  NAND U8847 ( .A(n8832), .B(n8831), .Z(n8827) );
  XOR U8848 ( .A(n191), .B(n190), .Z(\A1[46] ) );
  XOR U8849 ( .A(n8832), .B(n8833), .Z(n190) );
  XNOR U8850 ( .A(n8831), .B(n8829), .Z(n8833) );
  AND U8851 ( .A(n8834), .B(n8835), .Z(n8829) );
  NANDN U8852 ( .A(n8836), .B(n8837), .Z(n8835) );
  NANDN U8853 ( .A(n8838), .B(n8839), .Z(n8837) );
  NANDN U8854 ( .A(n8839), .B(n8838), .Z(n8834) );
  ANDN U8855 ( .B(B[17]), .A(n54), .Z(n8831) );
  XNOR U8856 ( .A(n8626), .B(n8840), .Z(n8832) );
  XNOR U8857 ( .A(n8625), .B(n8623), .Z(n8840) );
  AND U8858 ( .A(n8841), .B(n8842), .Z(n8623) );
  NANDN U8859 ( .A(n8843), .B(n8844), .Z(n8842) );
  OR U8860 ( .A(n8845), .B(n8846), .Z(n8844) );
  NAND U8861 ( .A(n8846), .B(n8845), .Z(n8841) );
  ANDN U8862 ( .B(B[18]), .A(n55), .Z(n8625) );
  XNOR U8863 ( .A(n8633), .B(n8847), .Z(n8626) );
  XNOR U8864 ( .A(n8632), .B(n8630), .Z(n8847) );
  AND U8865 ( .A(n8848), .B(n8849), .Z(n8630) );
  NANDN U8866 ( .A(n8850), .B(n8851), .Z(n8849) );
  NANDN U8867 ( .A(n8852), .B(n8853), .Z(n8851) );
  NANDN U8868 ( .A(n8853), .B(n8852), .Z(n8848) );
  ANDN U8869 ( .B(B[19]), .A(n56), .Z(n8632) );
  XNOR U8870 ( .A(n8640), .B(n8854), .Z(n8633) );
  XNOR U8871 ( .A(n8639), .B(n8637), .Z(n8854) );
  AND U8872 ( .A(n8855), .B(n8856), .Z(n8637) );
  NANDN U8873 ( .A(n8857), .B(n8858), .Z(n8856) );
  OR U8874 ( .A(n8859), .B(n8860), .Z(n8858) );
  NAND U8875 ( .A(n8860), .B(n8859), .Z(n8855) );
  ANDN U8876 ( .B(B[20]), .A(n57), .Z(n8639) );
  XNOR U8877 ( .A(n8647), .B(n8861), .Z(n8640) );
  XNOR U8878 ( .A(n8646), .B(n8644), .Z(n8861) );
  AND U8879 ( .A(n8862), .B(n8863), .Z(n8644) );
  NANDN U8880 ( .A(n8864), .B(n8865), .Z(n8863) );
  NANDN U8881 ( .A(n8866), .B(n8867), .Z(n8865) );
  NANDN U8882 ( .A(n8867), .B(n8866), .Z(n8862) );
  ANDN U8883 ( .B(B[21]), .A(n58), .Z(n8646) );
  XNOR U8884 ( .A(n8654), .B(n8868), .Z(n8647) );
  XNOR U8885 ( .A(n8653), .B(n8651), .Z(n8868) );
  AND U8886 ( .A(n8869), .B(n8870), .Z(n8651) );
  NANDN U8887 ( .A(n8871), .B(n8872), .Z(n8870) );
  OR U8888 ( .A(n8873), .B(n8874), .Z(n8872) );
  NAND U8889 ( .A(n8874), .B(n8873), .Z(n8869) );
  ANDN U8890 ( .B(B[22]), .A(n59), .Z(n8653) );
  XNOR U8891 ( .A(n8661), .B(n8875), .Z(n8654) );
  XNOR U8892 ( .A(n8660), .B(n8658), .Z(n8875) );
  AND U8893 ( .A(n8876), .B(n8877), .Z(n8658) );
  NANDN U8894 ( .A(n8878), .B(n8879), .Z(n8877) );
  NANDN U8895 ( .A(n8880), .B(n8881), .Z(n8879) );
  NANDN U8896 ( .A(n8881), .B(n8880), .Z(n8876) );
  ANDN U8897 ( .B(B[23]), .A(n60), .Z(n8660) );
  XNOR U8898 ( .A(n8668), .B(n8882), .Z(n8661) );
  XNOR U8899 ( .A(n8667), .B(n8665), .Z(n8882) );
  AND U8900 ( .A(n8883), .B(n8884), .Z(n8665) );
  NANDN U8901 ( .A(n8885), .B(n8886), .Z(n8884) );
  OR U8902 ( .A(n8887), .B(n8888), .Z(n8886) );
  NAND U8903 ( .A(n8888), .B(n8887), .Z(n8883) );
  ANDN U8904 ( .B(B[24]), .A(n61), .Z(n8667) );
  XNOR U8905 ( .A(n8675), .B(n8889), .Z(n8668) );
  XNOR U8906 ( .A(n8674), .B(n8672), .Z(n8889) );
  AND U8907 ( .A(n8890), .B(n8891), .Z(n8672) );
  NANDN U8908 ( .A(n8892), .B(n8893), .Z(n8891) );
  NANDN U8909 ( .A(n8894), .B(n8895), .Z(n8893) );
  NANDN U8910 ( .A(n8895), .B(n8894), .Z(n8890) );
  ANDN U8911 ( .B(B[25]), .A(n62), .Z(n8674) );
  XNOR U8912 ( .A(n8682), .B(n8896), .Z(n8675) );
  XNOR U8913 ( .A(n8681), .B(n8679), .Z(n8896) );
  AND U8914 ( .A(n8897), .B(n8898), .Z(n8679) );
  NANDN U8915 ( .A(n8899), .B(n8900), .Z(n8898) );
  OR U8916 ( .A(n8901), .B(n8902), .Z(n8900) );
  NAND U8917 ( .A(n8902), .B(n8901), .Z(n8897) );
  ANDN U8918 ( .B(B[26]), .A(n63), .Z(n8681) );
  XNOR U8919 ( .A(n8689), .B(n8903), .Z(n8682) );
  XNOR U8920 ( .A(n8688), .B(n8686), .Z(n8903) );
  AND U8921 ( .A(n8904), .B(n8905), .Z(n8686) );
  NANDN U8922 ( .A(n8906), .B(n8907), .Z(n8905) );
  NANDN U8923 ( .A(n8908), .B(n8909), .Z(n8907) );
  NANDN U8924 ( .A(n8909), .B(n8908), .Z(n8904) );
  ANDN U8925 ( .B(B[27]), .A(n64), .Z(n8688) );
  XNOR U8926 ( .A(n8696), .B(n8910), .Z(n8689) );
  XNOR U8927 ( .A(n8695), .B(n8693), .Z(n8910) );
  AND U8928 ( .A(n8911), .B(n8912), .Z(n8693) );
  NANDN U8929 ( .A(n8913), .B(n8914), .Z(n8912) );
  OR U8930 ( .A(n8915), .B(n8916), .Z(n8914) );
  NAND U8931 ( .A(n8916), .B(n8915), .Z(n8911) );
  ANDN U8932 ( .B(B[28]), .A(n65), .Z(n8695) );
  XNOR U8933 ( .A(n8703), .B(n8917), .Z(n8696) );
  XNOR U8934 ( .A(n8702), .B(n8700), .Z(n8917) );
  AND U8935 ( .A(n8918), .B(n8919), .Z(n8700) );
  NANDN U8936 ( .A(n8920), .B(n8921), .Z(n8919) );
  NANDN U8937 ( .A(n8922), .B(n8923), .Z(n8921) );
  NANDN U8938 ( .A(n8923), .B(n8922), .Z(n8918) );
  ANDN U8939 ( .B(B[29]), .A(n66), .Z(n8702) );
  XNOR U8940 ( .A(n8710), .B(n8924), .Z(n8703) );
  XNOR U8941 ( .A(n8709), .B(n8707), .Z(n8924) );
  AND U8942 ( .A(n8925), .B(n8926), .Z(n8707) );
  NANDN U8943 ( .A(n8927), .B(n8928), .Z(n8926) );
  OR U8944 ( .A(n8929), .B(n8930), .Z(n8928) );
  NAND U8945 ( .A(n8930), .B(n8929), .Z(n8925) );
  ANDN U8946 ( .B(B[30]), .A(n67), .Z(n8709) );
  XNOR U8947 ( .A(n8717), .B(n8931), .Z(n8710) );
  XNOR U8948 ( .A(n8716), .B(n8714), .Z(n8931) );
  AND U8949 ( .A(n8932), .B(n8933), .Z(n8714) );
  NANDN U8950 ( .A(n8934), .B(n8935), .Z(n8933) );
  NANDN U8951 ( .A(n8936), .B(n8937), .Z(n8935) );
  NANDN U8952 ( .A(n8937), .B(n8936), .Z(n8932) );
  ANDN U8953 ( .B(B[31]), .A(n68), .Z(n8716) );
  XNOR U8954 ( .A(n8724), .B(n8938), .Z(n8717) );
  XNOR U8955 ( .A(n8723), .B(n8721), .Z(n8938) );
  AND U8956 ( .A(n8939), .B(n8940), .Z(n8721) );
  NANDN U8957 ( .A(n8941), .B(n8942), .Z(n8940) );
  OR U8958 ( .A(n8943), .B(n8944), .Z(n8942) );
  NAND U8959 ( .A(n8944), .B(n8943), .Z(n8939) );
  ANDN U8960 ( .B(B[32]), .A(n69), .Z(n8723) );
  XNOR U8961 ( .A(n8731), .B(n8945), .Z(n8724) );
  XNOR U8962 ( .A(n8730), .B(n8728), .Z(n8945) );
  AND U8963 ( .A(n8946), .B(n8947), .Z(n8728) );
  NANDN U8964 ( .A(n8948), .B(n8949), .Z(n8947) );
  NANDN U8965 ( .A(n8950), .B(n8951), .Z(n8949) );
  NANDN U8966 ( .A(n8951), .B(n8950), .Z(n8946) );
  ANDN U8967 ( .B(B[33]), .A(n70), .Z(n8730) );
  XNOR U8968 ( .A(n8738), .B(n8952), .Z(n8731) );
  XNOR U8969 ( .A(n8737), .B(n8735), .Z(n8952) );
  AND U8970 ( .A(n8953), .B(n8954), .Z(n8735) );
  NANDN U8971 ( .A(n8955), .B(n8956), .Z(n8954) );
  OR U8972 ( .A(n8957), .B(n8958), .Z(n8956) );
  NAND U8973 ( .A(n8958), .B(n8957), .Z(n8953) );
  ANDN U8974 ( .B(B[34]), .A(n71), .Z(n8737) );
  XNOR U8975 ( .A(n8745), .B(n8959), .Z(n8738) );
  XNOR U8976 ( .A(n8744), .B(n8742), .Z(n8959) );
  AND U8977 ( .A(n8960), .B(n8961), .Z(n8742) );
  NANDN U8978 ( .A(n8962), .B(n8963), .Z(n8961) );
  NANDN U8979 ( .A(n8964), .B(n8965), .Z(n8963) );
  NANDN U8980 ( .A(n8965), .B(n8964), .Z(n8960) );
  ANDN U8981 ( .B(B[35]), .A(n72), .Z(n8744) );
  XNOR U8982 ( .A(n8752), .B(n8966), .Z(n8745) );
  XNOR U8983 ( .A(n8751), .B(n8749), .Z(n8966) );
  AND U8984 ( .A(n8967), .B(n8968), .Z(n8749) );
  NANDN U8985 ( .A(n8969), .B(n8970), .Z(n8968) );
  OR U8986 ( .A(n8971), .B(n8972), .Z(n8970) );
  NAND U8987 ( .A(n8972), .B(n8971), .Z(n8967) );
  ANDN U8988 ( .B(B[36]), .A(n73), .Z(n8751) );
  XNOR U8989 ( .A(n8759), .B(n8973), .Z(n8752) );
  XNOR U8990 ( .A(n8758), .B(n8756), .Z(n8973) );
  AND U8991 ( .A(n8974), .B(n8975), .Z(n8756) );
  NANDN U8992 ( .A(n8976), .B(n8977), .Z(n8975) );
  NANDN U8993 ( .A(n8978), .B(n8979), .Z(n8977) );
  NANDN U8994 ( .A(n8979), .B(n8978), .Z(n8974) );
  ANDN U8995 ( .B(B[37]), .A(n74), .Z(n8758) );
  XNOR U8996 ( .A(n8766), .B(n8980), .Z(n8759) );
  XNOR U8997 ( .A(n8765), .B(n8763), .Z(n8980) );
  AND U8998 ( .A(n8981), .B(n8982), .Z(n8763) );
  NANDN U8999 ( .A(n8983), .B(n8984), .Z(n8982) );
  OR U9000 ( .A(n8985), .B(n8986), .Z(n8984) );
  NAND U9001 ( .A(n8986), .B(n8985), .Z(n8981) );
  ANDN U9002 ( .B(B[38]), .A(n75), .Z(n8765) );
  XNOR U9003 ( .A(n8773), .B(n8987), .Z(n8766) );
  XNOR U9004 ( .A(n8772), .B(n8770), .Z(n8987) );
  AND U9005 ( .A(n8988), .B(n8989), .Z(n8770) );
  NANDN U9006 ( .A(n8990), .B(n8991), .Z(n8989) );
  NANDN U9007 ( .A(n8992), .B(n8993), .Z(n8991) );
  NANDN U9008 ( .A(n8993), .B(n8992), .Z(n8988) );
  ANDN U9009 ( .B(B[39]), .A(n76), .Z(n8772) );
  XNOR U9010 ( .A(n8780), .B(n8994), .Z(n8773) );
  XNOR U9011 ( .A(n8779), .B(n8777), .Z(n8994) );
  AND U9012 ( .A(n8995), .B(n8996), .Z(n8777) );
  NANDN U9013 ( .A(n8997), .B(n8998), .Z(n8996) );
  OR U9014 ( .A(n8999), .B(n9000), .Z(n8998) );
  NAND U9015 ( .A(n9000), .B(n8999), .Z(n8995) );
  ANDN U9016 ( .B(B[40]), .A(n77), .Z(n8779) );
  XNOR U9017 ( .A(n8787), .B(n9001), .Z(n8780) );
  XNOR U9018 ( .A(n8786), .B(n8784), .Z(n9001) );
  AND U9019 ( .A(n9002), .B(n9003), .Z(n8784) );
  NANDN U9020 ( .A(n9004), .B(n9005), .Z(n9003) );
  NANDN U9021 ( .A(n9006), .B(n9007), .Z(n9005) );
  NANDN U9022 ( .A(n9007), .B(n9006), .Z(n9002) );
  ANDN U9023 ( .B(B[41]), .A(n78), .Z(n8786) );
  XNOR U9024 ( .A(n8794), .B(n9008), .Z(n8787) );
  XNOR U9025 ( .A(n8793), .B(n8791), .Z(n9008) );
  AND U9026 ( .A(n9009), .B(n9010), .Z(n8791) );
  NANDN U9027 ( .A(n9011), .B(n9012), .Z(n9010) );
  OR U9028 ( .A(n9013), .B(n9014), .Z(n9012) );
  NAND U9029 ( .A(n9014), .B(n9013), .Z(n9009) );
  ANDN U9030 ( .B(B[42]), .A(n79), .Z(n8793) );
  XNOR U9031 ( .A(n8801), .B(n9015), .Z(n8794) );
  XNOR U9032 ( .A(n8800), .B(n8798), .Z(n9015) );
  AND U9033 ( .A(n9016), .B(n9017), .Z(n8798) );
  NANDN U9034 ( .A(n9018), .B(n9019), .Z(n9017) );
  NANDN U9035 ( .A(n9020), .B(n9021), .Z(n9019) );
  NANDN U9036 ( .A(n9021), .B(n9020), .Z(n9016) );
  ANDN U9037 ( .B(B[43]), .A(n80), .Z(n8800) );
  XNOR U9038 ( .A(n8808), .B(n9022), .Z(n8801) );
  XNOR U9039 ( .A(n8807), .B(n8805), .Z(n9022) );
  AND U9040 ( .A(n9023), .B(n9024), .Z(n8805) );
  NANDN U9041 ( .A(n9025), .B(n9026), .Z(n9024) );
  OR U9042 ( .A(n9027), .B(n9028), .Z(n9026) );
  NAND U9043 ( .A(n9028), .B(n9027), .Z(n9023) );
  ANDN U9044 ( .B(B[44]), .A(n81), .Z(n8807) );
  XNOR U9045 ( .A(n8815), .B(n9029), .Z(n8808) );
  XNOR U9046 ( .A(n8814), .B(n8812), .Z(n9029) );
  AND U9047 ( .A(n9030), .B(n9031), .Z(n8812) );
  NANDN U9048 ( .A(n9032), .B(n9033), .Z(n9031) );
  NAND U9049 ( .A(n9034), .B(n9035), .Z(n9033) );
  ANDN U9050 ( .B(B[45]), .A(n82), .Z(n8814) );
  XOR U9051 ( .A(n8821), .B(n9036), .Z(n8815) );
  XNOR U9052 ( .A(n8819), .B(n8822), .Z(n9036) );
  NAND U9053 ( .A(A[2]), .B(B[46]), .Z(n8822) );
  NANDN U9054 ( .A(n9037), .B(n9038), .Z(n8819) );
  AND U9055 ( .A(A[0]), .B(B[47]), .Z(n9038) );
  XNOR U9056 ( .A(n8824), .B(n9039), .Z(n8821) );
  NAND U9057 ( .A(A[0]), .B(B[48]), .Z(n9039) );
  NAND U9058 ( .A(B[47]), .B(A[1]), .Z(n8824) );
  NAND U9059 ( .A(n9040), .B(n9041), .Z(n191) );
  NANDN U9060 ( .A(n9042), .B(n9043), .Z(n9041) );
  OR U9061 ( .A(n9044), .B(n9045), .Z(n9043) );
  NAND U9062 ( .A(n9045), .B(n9044), .Z(n9040) );
  XOR U9063 ( .A(n193), .B(n192), .Z(\A1[45] ) );
  XOR U9064 ( .A(n9045), .B(n9046), .Z(n192) );
  XNOR U9065 ( .A(n9044), .B(n9042), .Z(n9046) );
  AND U9066 ( .A(n9047), .B(n9048), .Z(n9042) );
  NANDN U9067 ( .A(n9049), .B(n9050), .Z(n9048) );
  NANDN U9068 ( .A(n9051), .B(n9052), .Z(n9050) );
  NANDN U9069 ( .A(n9052), .B(n9051), .Z(n9047) );
  ANDN U9070 ( .B(B[16]), .A(n54), .Z(n9044) );
  XNOR U9071 ( .A(n8839), .B(n9053), .Z(n9045) );
  XNOR U9072 ( .A(n8838), .B(n8836), .Z(n9053) );
  AND U9073 ( .A(n9054), .B(n9055), .Z(n8836) );
  NANDN U9074 ( .A(n9056), .B(n9057), .Z(n9055) );
  OR U9075 ( .A(n9058), .B(n9059), .Z(n9057) );
  NAND U9076 ( .A(n9059), .B(n9058), .Z(n9054) );
  ANDN U9077 ( .B(B[17]), .A(n55), .Z(n8838) );
  XNOR U9078 ( .A(n8846), .B(n9060), .Z(n8839) );
  XNOR U9079 ( .A(n8845), .B(n8843), .Z(n9060) );
  AND U9080 ( .A(n9061), .B(n9062), .Z(n8843) );
  NANDN U9081 ( .A(n9063), .B(n9064), .Z(n9062) );
  NANDN U9082 ( .A(n9065), .B(n9066), .Z(n9064) );
  NANDN U9083 ( .A(n9066), .B(n9065), .Z(n9061) );
  ANDN U9084 ( .B(B[18]), .A(n56), .Z(n8845) );
  XNOR U9085 ( .A(n8853), .B(n9067), .Z(n8846) );
  XNOR U9086 ( .A(n8852), .B(n8850), .Z(n9067) );
  AND U9087 ( .A(n9068), .B(n9069), .Z(n8850) );
  NANDN U9088 ( .A(n9070), .B(n9071), .Z(n9069) );
  OR U9089 ( .A(n9072), .B(n9073), .Z(n9071) );
  NAND U9090 ( .A(n9073), .B(n9072), .Z(n9068) );
  ANDN U9091 ( .B(B[19]), .A(n57), .Z(n8852) );
  XNOR U9092 ( .A(n8860), .B(n9074), .Z(n8853) );
  XNOR U9093 ( .A(n8859), .B(n8857), .Z(n9074) );
  AND U9094 ( .A(n9075), .B(n9076), .Z(n8857) );
  NANDN U9095 ( .A(n9077), .B(n9078), .Z(n9076) );
  NANDN U9096 ( .A(n9079), .B(n9080), .Z(n9078) );
  NANDN U9097 ( .A(n9080), .B(n9079), .Z(n9075) );
  ANDN U9098 ( .B(B[20]), .A(n58), .Z(n8859) );
  XNOR U9099 ( .A(n8867), .B(n9081), .Z(n8860) );
  XNOR U9100 ( .A(n8866), .B(n8864), .Z(n9081) );
  AND U9101 ( .A(n9082), .B(n9083), .Z(n8864) );
  NANDN U9102 ( .A(n9084), .B(n9085), .Z(n9083) );
  OR U9103 ( .A(n9086), .B(n9087), .Z(n9085) );
  NAND U9104 ( .A(n9087), .B(n9086), .Z(n9082) );
  ANDN U9105 ( .B(B[21]), .A(n59), .Z(n8866) );
  XNOR U9106 ( .A(n8874), .B(n9088), .Z(n8867) );
  XNOR U9107 ( .A(n8873), .B(n8871), .Z(n9088) );
  AND U9108 ( .A(n9089), .B(n9090), .Z(n8871) );
  NANDN U9109 ( .A(n9091), .B(n9092), .Z(n9090) );
  NANDN U9110 ( .A(n9093), .B(n9094), .Z(n9092) );
  NANDN U9111 ( .A(n9094), .B(n9093), .Z(n9089) );
  ANDN U9112 ( .B(B[22]), .A(n60), .Z(n8873) );
  XNOR U9113 ( .A(n8881), .B(n9095), .Z(n8874) );
  XNOR U9114 ( .A(n8880), .B(n8878), .Z(n9095) );
  AND U9115 ( .A(n9096), .B(n9097), .Z(n8878) );
  NANDN U9116 ( .A(n9098), .B(n9099), .Z(n9097) );
  OR U9117 ( .A(n9100), .B(n9101), .Z(n9099) );
  NAND U9118 ( .A(n9101), .B(n9100), .Z(n9096) );
  ANDN U9119 ( .B(B[23]), .A(n61), .Z(n8880) );
  XNOR U9120 ( .A(n8888), .B(n9102), .Z(n8881) );
  XNOR U9121 ( .A(n8887), .B(n8885), .Z(n9102) );
  AND U9122 ( .A(n9103), .B(n9104), .Z(n8885) );
  NANDN U9123 ( .A(n9105), .B(n9106), .Z(n9104) );
  NANDN U9124 ( .A(n9107), .B(n9108), .Z(n9106) );
  NANDN U9125 ( .A(n9108), .B(n9107), .Z(n9103) );
  ANDN U9126 ( .B(B[24]), .A(n62), .Z(n8887) );
  XNOR U9127 ( .A(n8895), .B(n9109), .Z(n8888) );
  XNOR U9128 ( .A(n8894), .B(n8892), .Z(n9109) );
  AND U9129 ( .A(n9110), .B(n9111), .Z(n8892) );
  NANDN U9130 ( .A(n9112), .B(n9113), .Z(n9111) );
  OR U9131 ( .A(n9114), .B(n9115), .Z(n9113) );
  NAND U9132 ( .A(n9115), .B(n9114), .Z(n9110) );
  ANDN U9133 ( .B(B[25]), .A(n63), .Z(n8894) );
  XNOR U9134 ( .A(n8902), .B(n9116), .Z(n8895) );
  XNOR U9135 ( .A(n8901), .B(n8899), .Z(n9116) );
  AND U9136 ( .A(n9117), .B(n9118), .Z(n8899) );
  NANDN U9137 ( .A(n9119), .B(n9120), .Z(n9118) );
  NANDN U9138 ( .A(n9121), .B(n9122), .Z(n9120) );
  NANDN U9139 ( .A(n9122), .B(n9121), .Z(n9117) );
  ANDN U9140 ( .B(B[26]), .A(n64), .Z(n8901) );
  XNOR U9141 ( .A(n8909), .B(n9123), .Z(n8902) );
  XNOR U9142 ( .A(n8908), .B(n8906), .Z(n9123) );
  AND U9143 ( .A(n9124), .B(n9125), .Z(n8906) );
  NANDN U9144 ( .A(n9126), .B(n9127), .Z(n9125) );
  OR U9145 ( .A(n9128), .B(n9129), .Z(n9127) );
  NAND U9146 ( .A(n9129), .B(n9128), .Z(n9124) );
  ANDN U9147 ( .B(B[27]), .A(n65), .Z(n8908) );
  XNOR U9148 ( .A(n8916), .B(n9130), .Z(n8909) );
  XNOR U9149 ( .A(n8915), .B(n8913), .Z(n9130) );
  AND U9150 ( .A(n9131), .B(n9132), .Z(n8913) );
  NANDN U9151 ( .A(n9133), .B(n9134), .Z(n9132) );
  NANDN U9152 ( .A(n9135), .B(n9136), .Z(n9134) );
  NANDN U9153 ( .A(n9136), .B(n9135), .Z(n9131) );
  ANDN U9154 ( .B(B[28]), .A(n66), .Z(n8915) );
  XNOR U9155 ( .A(n8923), .B(n9137), .Z(n8916) );
  XNOR U9156 ( .A(n8922), .B(n8920), .Z(n9137) );
  AND U9157 ( .A(n9138), .B(n9139), .Z(n8920) );
  NANDN U9158 ( .A(n9140), .B(n9141), .Z(n9139) );
  OR U9159 ( .A(n9142), .B(n9143), .Z(n9141) );
  NAND U9160 ( .A(n9143), .B(n9142), .Z(n9138) );
  ANDN U9161 ( .B(B[29]), .A(n67), .Z(n8922) );
  XNOR U9162 ( .A(n8930), .B(n9144), .Z(n8923) );
  XNOR U9163 ( .A(n8929), .B(n8927), .Z(n9144) );
  AND U9164 ( .A(n9145), .B(n9146), .Z(n8927) );
  NANDN U9165 ( .A(n9147), .B(n9148), .Z(n9146) );
  NANDN U9166 ( .A(n9149), .B(n9150), .Z(n9148) );
  NANDN U9167 ( .A(n9150), .B(n9149), .Z(n9145) );
  ANDN U9168 ( .B(B[30]), .A(n68), .Z(n8929) );
  XNOR U9169 ( .A(n8937), .B(n9151), .Z(n8930) );
  XNOR U9170 ( .A(n8936), .B(n8934), .Z(n9151) );
  AND U9171 ( .A(n9152), .B(n9153), .Z(n8934) );
  NANDN U9172 ( .A(n9154), .B(n9155), .Z(n9153) );
  OR U9173 ( .A(n9156), .B(n9157), .Z(n9155) );
  NAND U9174 ( .A(n9157), .B(n9156), .Z(n9152) );
  ANDN U9175 ( .B(B[31]), .A(n69), .Z(n8936) );
  XNOR U9176 ( .A(n8944), .B(n9158), .Z(n8937) );
  XNOR U9177 ( .A(n8943), .B(n8941), .Z(n9158) );
  AND U9178 ( .A(n9159), .B(n9160), .Z(n8941) );
  NANDN U9179 ( .A(n9161), .B(n9162), .Z(n9160) );
  NANDN U9180 ( .A(n9163), .B(n9164), .Z(n9162) );
  NANDN U9181 ( .A(n9164), .B(n9163), .Z(n9159) );
  ANDN U9182 ( .B(B[32]), .A(n70), .Z(n8943) );
  XNOR U9183 ( .A(n8951), .B(n9165), .Z(n8944) );
  XNOR U9184 ( .A(n8950), .B(n8948), .Z(n9165) );
  AND U9185 ( .A(n9166), .B(n9167), .Z(n8948) );
  NANDN U9186 ( .A(n9168), .B(n9169), .Z(n9167) );
  OR U9187 ( .A(n9170), .B(n9171), .Z(n9169) );
  NAND U9188 ( .A(n9171), .B(n9170), .Z(n9166) );
  ANDN U9189 ( .B(B[33]), .A(n71), .Z(n8950) );
  XNOR U9190 ( .A(n8958), .B(n9172), .Z(n8951) );
  XNOR U9191 ( .A(n8957), .B(n8955), .Z(n9172) );
  AND U9192 ( .A(n9173), .B(n9174), .Z(n8955) );
  NANDN U9193 ( .A(n9175), .B(n9176), .Z(n9174) );
  NANDN U9194 ( .A(n9177), .B(n9178), .Z(n9176) );
  NANDN U9195 ( .A(n9178), .B(n9177), .Z(n9173) );
  ANDN U9196 ( .B(B[34]), .A(n72), .Z(n8957) );
  XNOR U9197 ( .A(n8965), .B(n9179), .Z(n8958) );
  XNOR U9198 ( .A(n8964), .B(n8962), .Z(n9179) );
  AND U9199 ( .A(n9180), .B(n9181), .Z(n8962) );
  NANDN U9200 ( .A(n9182), .B(n9183), .Z(n9181) );
  OR U9201 ( .A(n9184), .B(n9185), .Z(n9183) );
  NAND U9202 ( .A(n9185), .B(n9184), .Z(n9180) );
  ANDN U9203 ( .B(B[35]), .A(n73), .Z(n8964) );
  XNOR U9204 ( .A(n8972), .B(n9186), .Z(n8965) );
  XNOR U9205 ( .A(n8971), .B(n8969), .Z(n9186) );
  AND U9206 ( .A(n9187), .B(n9188), .Z(n8969) );
  NANDN U9207 ( .A(n9189), .B(n9190), .Z(n9188) );
  NANDN U9208 ( .A(n9191), .B(n9192), .Z(n9190) );
  NANDN U9209 ( .A(n9192), .B(n9191), .Z(n9187) );
  ANDN U9210 ( .B(B[36]), .A(n74), .Z(n8971) );
  XNOR U9211 ( .A(n8979), .B(n9193), .Z(n8972) );
  XNOR U9212 ( .A(n8978), .B(n8976), .Z(n9193) );
  AND U9213 ( .A(n9194), .B(n9195), .Z(n8976) );
  NANDN U9214 ( .A(n9196), .B(n9197), .Z(n9195) );
  OR U9215 ( .A(n9198), .B(n9199), .Z(n9197) );
  NAND U9216 ( .A(n9199), .B(n9198), .Z(n9194) );
  ANDN U9217 ( .B(B[37]), .A(n75), .Z(n8978) );
  XNOR U9218 ( .A(n8986), .B(n9200), .Z(n8979) );
  XNOR U9219 ( .A(n8985), .B(n8983), .Z(n9200) );
  AND U9220 ( .A(n9201), .B(n9202), .Z(n8983) );
  NANDN U9221 ( .A(n9203), .B(n9204), .Z(n9202) );
  NANDN U9222 ( .A(n9205), .B(n9206), .Z(n9204) );
  NANDN U9223 ( .A(n9206), .B(n9205), .Z(n9201) );
  ANDN U9224 ( .B(B[38]), .A(n76), .Z(n8985) );
  XNOR U9225 ( .A(n8993), .B(n9207), .Z(n8986) );
  XNOR U9226 ( .A(n8992), .B(n8990), .Z(n9207) );
  AND U9227 ( .A(n9208), .B(n9209), .Z(n8990) );
  NANDN U9228 ( .A(n9210), .B(n9211), .Z(n9209) );
  OR U9229 ( .A(n9212), .B(n9213), .Z(n9211) );
  NAND U9230 ( .A(n9213), .B(n9212), .Z(n9208) );
  ANDN U9231 ( .B(B[39]), .A(n77), .Z(n8992) );
  XNOR U9232 ( .A(n9000), .B(n9214), .Z(n8993) );
  XNOR U9233 ( .A(n8999), .B(n8997), .Z(n9214) );
  AND U9234 ( .A(n9215), .B(n9216), .Z(n8997) );
  NANDN U9235 ( .A(n9217), .B(n9218), .Z(n9216) );
  NANDN U9236 ( .A(n9219), .B(n9220), .Z(n9218) );
  NANDN U9237 ( .A(n9220), .B(n9219), .Z(n9215) );
  ANDN U9238 ( .B(B[40]), .A(n78), .Z(n8999) );
  XNOR U9239 ( .A(n9007), .B(n9221), .Z(n9000) );
  XNOR U9240 ( .A(n9006), .B(n9004), .Z(n9221) );
  AND U9241 ( .A(n9222), .B(n9223), .Z(n9004) );
  NANDN U9242 ( .A(n9224), .B(n9225), .Z(n9223) );
  OR U9243 ( .A(n9226), .B(n9227), .Z(n9225) );
  NAND U9244 ( .A(n9227), .B(n9226), .Z(n9222) );
  ANDN U9245 ( .B(B[41]), .A(n79), .Z(n9006) );
  XNOR U9246 ( .A(n9014), .B(n9228), .Z(n9007) );
  XNOR U9247 ( .A(n9013), .B(n9011), .Z(n9228) );
  AND U9248 ( .A(n9229), .B(n9230), .Z(n9011) );
  NANDN U9249 ( .A(n9231), .B(n9232), .Z(n9230) );
  NANDN U9250 ( .A(n9233), .B(n9234), .Z(n9232) );
  NANDN U9251 ( .A(n9234), .B(n9233), .Z(n9229) );
  ANDN U9252 ( .B(B[42]), .A(n80), .Z(n9013) );
  XNOR U9253 ( .A(n9021), .B(n9235), .Z(n9014) );
  XNOR U9254 ( .A(n9020), .B(n9018), .Z(n9235) );
  AND U9255 ( .A(n9236), .B(n9237), .Z(n9018) );
  NANDN U9256 ( .A(n9238), .B(n9239), .Z(n9237) );
  OR U9257 ( .A(n9240), .B(n9241), .Z(n9239) );
  NAND U9258 ( .A(n9241), .B(n9240), .Z(n9236) );
  ANDN U9259 ( .B(B[43]), .A(n81), .Z(n9020) );
  XNOR U9260 ( .A(n9028), .B(n9242), .Z(n9021) );
  XNOR U9261 ( .A(n9027), .B(n9025), .Z(n9242) );
  AND U9262 ( .A(n9243), .B(n9244), .Z(n9025) );
  NANDN U9263 ( .A(n9245), .B(n9246), .Z(n9244) );
  NAND U9264 ( .A(n9247), .B(n9248), .Z(n9246) );
  ANDN U9265 ( .B(B[44]), .A(n82), .Z(n9027) );
  XOR U9266 ( .A(n9034), .B(n9249), .Z(n9028) );
  XNOR U9267 ( .A(n9032), .B(n9035), .Z(n9249) );
  NAND U9268 ( .A(A[2]), .B(B[45]), .Z(n9035) );
  NANDN U9269 ( .A(n9250), .B(n9251), .Z(n9032) );
  AND U9270 ( .A(A[0]), .B(B[46]), .Z(n9251) );
  XNOR U9271 ( .A(n9037), .B(n9252), .Z(n9034) );
  NAND U9272 ( .A(A[0]), .B(B[47]), .Z(n9252) );
  NAND U9273 ( .A(B[46]), .B(A[1]), .Z(n9037) );
  NAND U9274 ( .A(n9253), .B(n9254), .Z(n193) );
  NANDN U9275 ( .A(n9255), .B(n9256), .Z(n9254) );
  OR U9276 ( .A(n9257), .B(n9258), .Z(n9256) );
  NAND U9277 ( .A(n9258), .B(n9257), .Z(n9253) );
  XOR U9278 ( .A(n195), .B(n194), .Z(\A1[44] ) );
  XOR U9279 ( .A(n9258), .B(n9259), .Z(n194) );
  XNOR U9280 ( .A(n9257), .B(n9255), .Z(n9259) );
  AND U9281 ( .A(n9260), .B(n9261), .Z(n9255) );
  NANDN U9282 ( .A(n9262), .B(n9263), .Z(n9261) );
  NANDN U9283 ( .A(n9264), .B(n9265), .Z(n9263) );
  NANDN U9284 ( .A(n9265), .B(n9264), .Z(n9260) );
  ANDN U9285 ( .B(B[15]), .A(n54), .Z(n9257) );
  XNOR U9286 ( .A(n9052), .B(n9266), .Z(n9258) );
  XNOR U9287 ( .A(n9051), .B(n9049), .Z(n9266) );
  AND U9288 ( .A(n9267), .B(n9268), .Z(n9049) );
  NANDN U9289 ( .A(n9269), .B(n9270), .Z(n9268) );
  OR U9290 ( .A(n9271), .B(n9272), .Z(n9270) );
  NAND U9291 ( .A(n9272), .B(n9271), .Z(n9267) );
  ANDN U9292 ( .B(B[16]), .A(n55), .Z(n9051) );
  XNOR U9293 ( .A(n9059), .B(n9273), .Z(n9052) );
  XNOR U9294 ( .A(n9058), .B(n9056), .Z(n9273) );
  AND U9295 ( .A(n9274), .B(n9275), .Z(n9056) );
  NANDN U9296 ( .A(n9276), .B(n9277), .Z(n9275) );
  NANDN U9297 ( .A(n9278), .B(n9279), .Z(n9277) );
  NANDN U9298 ( .A(n9279), .B(n9278), .Z(n9274) );
  ANDN U9299 ( .B(B[17]), .A(n56), .Z(n9058) );
  XNOR U9300 ( .A(n9066), .B(n9280), .Z(n9059) );
  XNOR U9301 ( .A(n9065), .B(n9063), .Z(n9280) );
  AND U9302 ( .A(n9281), .B(n9282), .Z(n9063) );
  NANDN U9303 ( .A(n9283), .B(n9284), .Z(n9282) );
  OR U9304 ( .A(n9285), .B(n9286), .Z(n9284) );
  NAND U9305 ( .A(n9286), .B(n9285), .Z(n9281) );
  ANDN U9306 ( .B(B[18]), .A(n57), .Z(n9065) );
  XNOR U9307 ( .A(n9073), .B(n9287), .Z(n9066) );
  XNOR U9308 ( .A(n9072), .B(n9070), .Z(n9287) );
  AND U9309 ( .A(n9288), .B(n9289), .Z(n9070) );
  NANDN U9310 ( .A(n9290), .B(n9291), .Z(n9289) );
  NANDN U9311 ( .A(n9292), .B(n9293), .Z(n9291) );
  NANDN U9312 ( .A(n9293), .B(n9292), .Z(n9288) );
  ANDN U9313 ( .B(B[19]), .A(n58), .Z(n9072) );
  XNOR U9314 ( .A(n9080), .B(n9294), .Z(n9073) );
  XNOR U9315 ( .A(n9079), .B(n9077), .Z(n9294) );
  AND U9316 ( .A(n9295), .B(n9296), .Z(n9077) );
  NANDN U9317 ( .A(n9297), .B(n9298), .Z(n9296) );
  OR U9318 ( .A(n9299), .B(n9300), .Z(n9298) );
  NAND U9319 ( .A(n9300), .B(n9299), .Z(n9295) );
  ANDN U9320 ( .B(B[20]), .A(n59), .Z(n9079) );
  XNOR U9321 ( .A(n9087), .B(n9301), .Z(n9080) );
  XNOR U9322 ( .A(n9086), .B(n9084), .Z(n9301) );
  AND U9323 ( .A(n9302), .B(n9303), .Z(n9084) );
  NANDN U9324 ( .A(n9304), .B(n9305), .Z(n9303) );
  NANDN U9325 ( .A(n9306), .B(n9307), .Z(n9305) );
  NANDN U9326 ( .A(n9307), .B(n9306), .Z(n9302) );
  ANDN U9327 ( .B(B[21]), .A(n60), .Z(n9086) );
  XNOR U9328 ( .A(n9094), .B(n9308), .Z(n9087) );
  XNOR U9329 ( .A(n9093), .B(n9091), .Z(n9308) );
  AND U9330 ( .A(n9309), .B(n9310), .Z(n9091) );
  NANDN U9331 ( .A(n9311), .B(n9312), .Z(n9310) );
  OR U9332 ( .A(n9313), .B(n9314), .Z(n9312) );
  NAND U9333 ( .A(n9314), .B(n9313), .Z(n9309) );
  ANDN U9334 ( .B(B[22]), .A(n61), .Z(n9093) );
  XNOR U9335 ( .A(n9101), .B(n9315), .Z(n9094) );
  XNOR U9336 ( .A(n9100), .B(n9098), .Z(n9315) );
  AND U9337 ( .A(n9316), .B(n9317), .Z(n9098) );
  NANDN U9338 ( .A(n9318), .B(n9319), .Z(n9317) );
  NANDN U9339 ( .A(n9320), .B(n9321), .Z(n9319) );
  NANDN U9340 ( .A(n9321), .B(n9320), .Z(n9316) );
  ANDN U9341 ( .B(B[23]), .A(n62), .Z(n9100) );
  XNOR U9342 ( .A(n9108), .B(n9322), .Z(n9101) );
  XNOR U9343 ( .A(n9107), .B(n9105), .Z(n9322) );
  AND U9344 ( .A(n9323), .B(n9324), .Z(n9105) );
  NANDN U9345 ( .A(n9325), .B(n9326), .Z(n9324) );
  OR U9346 ( .A(n9327), .B(n9328), .Z(n9326) );
  NAND U9347 ( .A(n9328), .B(n9327), .Z(n9323) );
  ANDN U9348 ( .B(B[24]), .A(n63), .Z(n9107) );
  XNOR U9349 ( .A(n9115), .B(n9329), .Z(n9108) );
  XNOR U9350 ( .A(n9114), .B(n9112), .Z(n9329) );
  AND U9351 ( .A(n9330), .B(n9331), .Z(n9112) );
  NANDN U9352 ( .A(n9332), .B(n9333), .Z(n9331) );
  NANDN U9353 ( .A(n9334), .B(n9335), .Z(n9333) );
  NANDN U9354 ( .A(n9335), .B(n9334), .Z(n9330) );
  ANDN U9355 ( .B(B[25]), .A(n64), .Z(n9114) );
  XNOR U9356 ( .A(n9122), .B(n9336), .Z(n9115) );
  XNOR U9357 ( .A(n9121), .B(n9119), .Z(n9336) );
  AND U9358 ( .A(n9337), .B(n9338), .Z(n9119) );
  NANDN U9359 ( .A(n9339), .B(n9340), .Z(n9338) );
  OR U9360 ( .A(n9341), .B(n9342), .Z(n9340) );
  NAND U9361 ( .A(n9342), .B(n9341), .Z(n9337) );
  ANDN U9362 ( .B(B[26]), .A(n65), .Z(n9121) );
  XNOR U9363 ( .A(n9129), .B(n9343), .Z(n9122) );
  XNOR U9364 ( .A(n9128), .B(n9126), .Z(n9343) );
  AND U9365 ( .A(n9344), .B(n9345), .Z(n9126) );
  NANDN U9366 ( .A(n9346), .B(n9347), .Z(n9345) );
  NANDN U9367 ( .A(n9348), .B(n9349), .Z(n9347) );
  NANDN U9368 ( .A(n9349), .B(n9348), .Z(n9344) );
  ANDN U9369 ( .B(B[27]), .A(n66), .Z(n9128) );
  XNOR U9370 ( .A(n9136), .B(n9350), .Z(n9129) );
  XNOR U9371 ( .A(n9135), .B(n9133), .Z(n9350) );
  AND U9372 ( .A(n9351), .B(n9352), .Z(n9133) );
  NANDN U9373 ( .A(n9353), .B(n9354), .Z(n9352) );
  OR U9374 ( .A(n9355), .B(n9356), .Z(n9354) );
  NAND U9375 ( .A(n9356), .B(n9355), .Z(n9351) );
  ANDN U9376 ( .B(B[28]), .A(n67), .Z(n9135) );
  XNOR U9377 ( .A(n9143), .B(n9357), .Z(n9136) );
  XNOR U9378 ( .A(n9142), .B(n9140), .Z(n9357) );
  AND U9379 ( .A(n9358), .B(n9359), .Z(n9140) );
  NANDN U9380 ( .A(n9360), .B(n9361), .Z(n9359) );
  NANDN U9381 ( .A(n9362), .B(n9363), .Z(n9361) );
  NANDN U9382 ( .A(n9363), .B(n9362), .Z(n9358) );
  ANDN U9383 ( .B(B[29]), .A(n68), .Z(n9142) );
  XNOR U9384 ( .A(n9150), .B(n9364), .Z(n9143) );
  XNOR U9385 ( .A(n9149), .B(n9147), .Z(n9364) );
  AND U9386 ( .A(n9365), .B(n9366), .Z(n9147) );
  NANDN U9387 ( .A(n9367), .B(n9368), .Z(n9366) );
  OR U9388 ( .A(n9369), .B(n9370), .Z(n9368) );
  NAND U9389 ( .A(n9370), .B(n9369), .Z(n9365) );
  ANDN U9390 ( .B(B[30]), .A(n69), .Z(n9149) );
  XNOR U9391 ( .A(n9157), .B(n9371), .Z(n9150) );
  XNOR U9392 ( .A(n9156), .B(n9154), .Z(n9371) );
  AND U9393 ( .A(n9372), .B(n9373), .Z(n9154) );
  NANDN U9394 ( .A(n9374), .B(n9375), .Z(n9373) );
  NANDN U9395 ( .A(n9376), .B(n9377), .Z(n9375) );
  NANDN U9396 ( .A(n9377), .B(n9376), .Z(n9372) );
  ANDN U9397 ( .B(B[31]), .A(n70), .Z(n9156) );
  XNOR U9398 ( .A(n9164), .B(n9378), .Z(n9157) );
  XNOR U9399 ( .A(n9163), .B(n9161), .Z(n9378) );
  AND U9400 ( .A(n9379), .B(n9380), .Z(n9161) );
  NANDN U9401 ( .A(n9381), .B(n9382), .Z(n9380) );
  OR U9402 ( .A(n9383), .B(n9384), .Z(n9382) );
  NAND U9403 ( .A(n9384), .B(n9383), .Z(n9379) );
  ANDN U9404 ( .B(B[32]), .A(n71), .Z(n9163) );
  XNOR U9405 ( .A(n9171), .B(n9385), .Z(n9164) );
  XNOR U9406 ( .A(n9170), .B(n9168), .Z(n9385) );
  AND U9407 ( .A(n9386), .B(n9387), .Z(n9168) );
  NANDN U9408 ( .A(n9388), .B(n9389), .Z(n9387) );
  NANDN U9409 ( .A(n9390), .B(n9391), .Z(n9389) );
  NANDN U9410 ( .A(n9391), .B(n9390), .Z(n9386) );
  ANDN U9411 ( .B(B[33]), .A(n72), .Z(n9170) );
  XNOR U9412 ( .A(n9178), .B(n9392), .Z(n9171) );
  XNOR U9413 ( .A(n9177), .B(n9175), .Z(n9392) );
  AND U9414 ( .A(n9393), .B(n9394), .Z(n9175) );
  NANDN U9415 ( .A(n9395), .B(n9396), .Z(n9394) );
  OR U9416 ( .A(n9397), .B(n9398), .Z(n9396) );
  NAND U9417 ( .A(n9398), .B(n9397), .Z(n9393) );
  ANDN U9418 ( .B(B[34]), .A(n73), .Z(n9177) );
  XNOR U9419 ( .A(n9185), .B(n9399), .Z(n9178) );
  XNOR U9420 ( .A(n9184), .B(n9182), .Z(n9399) );
  AND U9421 ( .A(n9400), .B(n9401), .Z(n9182) );
  NANDN U9422 ( .A(n9402), .B(n9403), .Z(n9401) );
  NANDN U9423 ( .A(n9404), .B(n9405), .Z(n9403) );
  NANDN U9424 ( .A(n9405), .B(n9404), .Z(n9400) );
  ANDN U9425 ( .B(B[35]), .A(n74), .Z(n9184) );
  XNOR U9426 ( .A(n9192), .B(n9406), .Z(n9185) );
  XNOR U9427 ( .A(n9191), .B(n9189), .Z(n9406) );
  AND U9428 ( .A(n9407), .B(n9408), .Z(n9189) );
  NANDN U9429 ( .A(n9409), .B(n9410), .Z(n9408) );
  OR U9430 ( .A(n9411), .B(n9412), .Z(n9410) );
  NAND U9431 ( .A(n9412), .B(n9411), .Z(n9407) );
  ANDN U9432 ( .B(B[36]), .A(n75), .Z(n9191) );
  XNOR U9433 ( .A(n9199), .B(n9413), .Z(n9192) );
  XNOR U9434 ( .A(n9198), .B(n9196), .Z(n9413) );
  AND U9435 ( .A(n9414), .B(n9415), .Z(n9196) );
  NANDN U9436 ( .A(n9416), .B(n9417), .Z(n9415) );
  NANDN U9437 ( .A(n9418), .B(n9419), .Z(n9417) );
  NANDN U9438 ( .A(n9419), .B(n9418), .Z(n9414) );
  ANDN U9439 ( .B(B[37]), .A(n76), .Z(n9198) );
  XNOR U9440 ( .A(n9206), .B(n9420), .Z(n9199) );
  XNOR U9441 ( .A(n9205), .B(n9203), .Z(n9420) );
  AND U9442 ( .A(n9421), .B(n9422), .Z(n9203) );
  NANDN U9443 ( .A(n9423), .B(n9424), .Z(n9422) );
  OR U9444 ( .A(n9425), .B(n9426), .Z(n9424) );
  NAND U9445 ( .A(n9426), .B(n9425), .Z(n9421) );
  ANDN U9446 ( .B(B[38]), .A(n77), .Z(n9205) );
  XNOR U9447 ( .A(n9213), .B(n9427), .Z(n9206) );
  XNOR U9448 ( .A(n9212), .B(n9210), .Z(n9427) );
  AND U9449 ( .A(n9428), .B(n9429), .Z(n9210) );
  NANDN U9450 ( .A(n9430), .B(n9431), .Z(n9429) );
  NANDN U9451 ( .A(n9432), .B(n9433), .Z(n9431) );
  NANDN U9452 ( .A(n9433), .B(n9432), .Z(n9428) );
  ANDN U9453 ( .B(B[39]), .A(n78), .Z(n9212) );
  XNOR U9454 ( .A(n9220), .B(n9434), .Z(n9213) );
  XNOR U9455 ( .A(n9219), .B(n9217), .Z(n9434) );
  AND U9456 ( .A(n9435), .B(n9436), .Z(n9217) );
  NANDN U9457 ( .A(n9437), .B(n9438), .Z(n9436) );
  OR U9458 ( .A(n9439), .B(n9440), .Z(n9438) );
  NAND U9459 ( .A(n9440), .B(n9439), .Z(n9435) );
  ANDN U9460 ( .B(B[40]), .A(n79), .Z(n9219) );
  XNOR U9461 ( .A(n9227), .B(n9441), .Z(n9220) );
  XNOR U9462 ( .A(n9226), .B(n9224), .Z(n9441) );
  AND U9463 ( .A(n9442), .B(n9443), .Z(n9224) );
  NANDN U9464 ( .A(n9444), .B(n9445), .Z(n9443) );
  NANDN U9465 ( .A(n9446), .B(n9447), .Z(n9445) );
  NANDN U9466 ( .A(n9447), .B(n9446), .Z(n9442) );
  ANDN U9467 ( .B(B[41]), .A(n80), .Z(n9226) );
  XNOR U9468 ( .A(n9234), .B(n9448), .Z(n9227) );
  XNOR U9469 ( .A(n9233), .B(n9231), .Z(n9448) );
  AND U9470 ( .A(n9449), .B(n9450), .Z(n9231) );
  NANDN U9471 ( .A(n9451), .B(n9452), .Z(n9450) );
  OR U9472 ( .A(n9453), .B(n9454), .Z(n9452) );
  NAND U9473 ( .A(n9454), .B(n9453), .Z(n9449) );
  ANDN U9474 ( .B(B[42]), .A(n81), .Z(n9233) );
  XNOR U9475 ( .A(n9241), .B(n9455), .Z(n9234) );
  XNOR U9476 ( .A(n9240), .B(n9238), .Z(n9455) );
  AND U9477 ( .A(n9456), .B(n9457), .Z(n9238) );
  NANDN U9478 ( .A(n9458), .B(n9459), .Z(n9457) );
  NAND U9479 ( .A(n9460), .B(n9461), .Z(n9459) );
  ANDN U9480 ( .B(B[43]), .A(n82), .Z(n9240) );
  XOR U9481 ( .A(n9247), .B(n9462), .Z(n9241) );
  XNOR U9482 ( .A(n9245), .B(n9248), .Z(n9462) );
  NAND U9483 ( .A(A[2]), .B(B[44]), .Z(n9248) );
  NANDN U9484 ( .A(n9463), .B(n9464), .Z(n9245) );
  AND U9485 ( .A(A[0]), .B(B[45]), .Z(n9464) );
  XNOR U9486 ( .A(n9250), .B(n9465), .Z(n9247) );
  NAND U9487 ( .A(A[0]), .B(B[46]), .Z(n9465) );
  NAND U9488 ( .A(B[45]), .B(A[1]), .Z(n9250) );
  NAND U9489 ( .A(n9466), .B(n9467), .Z(n195) );
  NANDN U9490 ( .A(n9468), .B(n9469), .Z(n9467) );
  OR U9491 ( .A(n9470), .B(n9471), .Z(n9469) );
  NAND U9492 ( .A(n9471), .B(n9470), .Z(n9466) );
  XOR U9493 ( .A(n197), .B(n196), .Z(\A1[43] ) );
  XOR U9494 ( .A(n9471), .B(n9472), .Z(n196) );
  XNOR U9495 ( .A(n9470), .B(n9468), .Z(n9472) );
  AND U9496 ( .A(n9473), .B(n9474), .Z(n9468) );
  NANDN U9497 ( .A(n9475), .B(n9476), .Z(n9474) );
  NANDN U9498 ( .A(n9477), .B(n9478), .Z(n9476) );
  NANDN U9499 ( .A(n9478), .B(n9477), .Z(n9473) );
  ANDN U9500 ( .B(B[14]), .A(n54), .Z(n9470) );
  XNOR U9501 ( .A(n9265), .B(n9479), .Z(n9471) );
  XNOR U9502 ( .A(n9264), .B(n9262), .Z(n9479) );
  AND U9503 ( .A(n9480), .B(n9481), .Z(n9262) );
  NANDN U9504 ( .A(n9482), .B(n9483), .Z(n9481) );
  OR U9505 ( .A(n9484), .B(n9485), .Z(n9483) );
  NAND U9506 ( .A(n9485), .B(n9484), .Z(n9480) );
  ANDN U9507 ( .B(B[15]), .A(n55), .Z(n9264) );
  XNOR U9508 ( .A(n9272), .B(n9486), .Z(n9265) );
  XNOR U9509 ( .A(n9271), .B(n9269), .Z(n9486) );
  AND U9510 ( .A(n9487), .B(n9488), .Z(n9269) );
  NANDN U9511 ( .A(n9489), .B(n9490), .Z(n9488) );
  NANDN U9512 ( .A(n9491), .B(n9492), .Z(n9490) );
  NANDN U9513 ( .A(n9492), .B(n9491), .Z(n9487) );
  ANDN U9514 ( .B(B[16]), .A(n56), .Z(n9271) );
  XNOR U9515 ( .A(n9279), .B(n9493), .Z(n9272) );
  XNOR U9516 ( .A(n9278), .B(n9276), .Z(n9493) );
  AND U9517 ( .A(n9494), .B(n9495), .Z(n9276) );
  NANDN U9518 ( .A(n9496), .B(n9497), .Z(n9495) );
  OR U9519 ( .A(n9498), .B(n9499), .Z(n9497) );
  NAND U9520 ( .A(n9499), .B(n9498), .Z(n9494) );
  ANDN U9521 ( .B(B[17]), .A(n57), .Z(n9278) );
  XNOR U9522 ( .A(n9286), .B(n9500), .Z(n9279) );
  XNOR U9523 ( .A(n9285), .B(n9283), .Z(n9500) );
  AND U9524 ( .A(n9501), .B(n9502), .Z(n9283) );
  NANDN U9525 ( .A(n9503), .B(n9504), .Z(n9502) );
  NANDN U9526 ( .A(n9505), .B(n9506), .Z(n9504) );
  NANDN U9527 ( .A(n9506), .B(n9505), .Z(n9501) );
  ANDN U9528 ( .B(B[18]), .A(n58), .Z(n9285) );
  XNOR U9529 ( .A(n9293), .B(n9507), .Z(n9286) );
  XNOR U9530 ( .A(n9292), .B(n9290), .Z(n9507) );
  AND U9531 ( .A(n9508), .B(n9509), .Z(n9290) );
  NANDN U9532 ( .A(n9510), .B(n9511), .Z(n9509) );
  OR U9533 ( .A(n9512), .B(n9513), .Z(n9511) );
  NAND U9534 ( .A(n9513), .B(n9512), .Z(n9508) );
  ANDN U9535 ( .B(B[19]), .A(n59), .Z(n9292) );
  XNOR U9536 ( .A(n9300), .B(n9514), .Z(n9293) );
  XNOR U9537 ( .A(n9299), .B(n9297), .Z(n9514) );
  AND U9538 ( .A(n9515), .B(n9516), .Z(n9297) );
  NANDN U9539 ( .A(n9517), .B(n9518), .Z(n9516) );
  NANDN U9540 ( .A(n9519), .B(n9520), .Z(n9518) );
  NANDN U9541 ( .A(n9520), .B(n9519), .Z(n9515) );
  ANDN U9542 ( .B(B[20]), .A(n60), .Z(n9299) );
  XNOR U9543 ( .A(n9307), .B(n9521), .Z(n9300) );
  XNOR U9544 ( .A(n9306), .B(n9304), .Z(n9521) );
  AND U9545 ( .A(n9522), .B(n9523), .Z(n9304) );
  NANDN U9546 ( .A(n9524), .B(n9525), .Z(n9523) );
  OR U9547 ( .A(n9526), .B(n9527), .Z(n9525) );
  NAND U9548 ( .A(n9527), .B(n9526), .Z(n9522) );
  ANDN U9549 ( .B(B[21]), .A(n61), .Z(n9306) );
  XNOR U9550 ( .A(n9314), .B(n9528), .Z(n9307) );
  XNOR U9551 ( .A(n9313), .B(n9311), .Z(n9528) );
  AND U9552 ( .A(n9529), .B(n9530), .Z(n9311) );
  NANDN U9553 ( .A(n9531), .B(n9532), .Z(n9530) );
  NANDN U9554 ( .A(n9533), .B(n9534), .Z(n9532) );
  NANDN U9555 ( .A(n9534), .B(n9533), .Z(n9529) );
  ANDN U9556 ( .B(B[22]), .A(n62), .Z(n9313) );
  XNOR U9557 ( .A(n9321), .B(n9535), .Z(n9314) );
  XNOR U9558 ( .A(n9320), .B(n9318), .Z(n9535) );
  AND U9559 ( .A(n9536), .B(n9537), .Z(n9318) );
  NANDN U9560 ( .A(n9538), .B(n9539), .Z(n9537) );
  OR U9561 ( .A(n9540), .B(n9541), .Z(n9539) );
  NAND U9562 ( .A(n9541), .B(n9540), .Z(n9536) );
  ANDN U9563 ( .B(B[23]), .A(n63), .Z(n9320) );
  XNOR U9564 ( .A(n9328), .B(n9542), .Z(n9321) );
  XNOR U9565 ( .A(n9327), .B(n9325), .Z(n9542) );
  AND U9566 ( .A(n9543), .B(n9544), .Z(n9325) );
  NANDN U9567 ( .A(n9545), .B(n9546), .Z(n9544) );
  NANDN U9568 ( .A(n9547), .B(n9548), .Z(n9546) );
  NANDN U9569 ( .A(n9548), .B(n9547), .Z(n9543) );
  ANDN U9570 ( .B(B[24]), .A(n64), .Z(n9327) );
  XNOR U9571 ( .A(n9335), .B(n9549), .Z(n9328) );
  XNOR U9572 ( .A(n9334), .B(n9332), .Z(n9549) );
  AND U9573 ( .A(n9550), .B(n9551), .Z(n9332) );
  NANDN U9574 ( .A(n9552), .B(n9553), .Z(n9551) );
  OR U9575 ( .A(n9554), .B(n9555), .Z(n9553) );
  NAND U9576 ( .A(n9555), .B(n9554), .Z(n9550) );
  ANDN U9577 ( .B(B[25]), .A(n65), .Z(n9334) );
  XNOR U9578 ( .A(n9342), .B(n9556), .Z(n9335) );
  XNOR U9579 ( .A(n9341), .B(n9339), .Z(n9556) );
  AND U9580 ( .A(n9557), .B(n9558), .Z(n9339) );
  NANDN U9581 ( .A(n9559), .B(n9560), .Z(n9558) );
  NANDN U9582 ( .A(n9561), .B(n9562), .Z(n9560) );
  NANDN U9583 ( .A(n9562), .B(n9561), .Z(n9557) );
  ANDN U9584 ( .B(B[26]), .A(n66), .Z(n9341) );
  XNOR U9585 ( .A(n9349), .B(n9563), .Z(n9342) );
  XNOR U9586 ( .A(n9348), .B(n9346), .Z(n9563) );
  AND U9587 ( .A(n9564), .B(n9565), .Z(n9346) );
  NANDN U9588 ( .A(n9566), .B(n9567), .Z(n9565) );
  OR U9589 ( .A(n9568), .B(n9569), .Z(n9567) );
  NAND U9590 ( .A(n9569), .B(n9568), .Z(n9564) );
  ANDN U9591 ( .B(B[27]), .A(n67), .Z(n9348) );
  XNOR U9592 ( .A(n9356), .B(n9570), .Z(n9349) );
  XNOR U9593 ( .A(n9355), .B(n9353), .Z(n9570) );
  AND U9594 ( .A(n9571), .B(n9572), .Z(n9353) );
  NANDN U9595 ( .A(n9573), .B(n9574), .Z(n9572) );
  NANDN U9596 ( .A(n9575), .B(n9576), .Z(n9574) );
  NANDN U9597 ( .A(n9576), .B(n9575), .Z(n9571) );
  ANDN U9598 ( .B(B[28]), .A(n68), .Z(n9355) );
  XNOR U9599 ( .A(n9363), .B(n9577), .Z(n9356) );
  XNOR U9600 ( .A(n9362), .B(n9360), .Z(n9577) );
  AND U9601 ( .A(n9578), .B(n9579), .Z(n9360) );
  NANDN U9602 ( .A(n9580), .B(n9581), .Z(n9579) );
  OR U9603 ( .A(n9582), .B(n9583), .Z(n9581) );
  NAND U9604 ( .A(n9583), .B(n9582), .Z(n9578) );
  ANDN U9605 ( .B(B[29]), .A(n69), .Z(n9362) );
  XNOR U9606 ( .A(n9370), .B(n9584), .Z(n9363) );
  XNOR U9607 ( .A(n9369), .B(n9367), .Z(n9584) );
  AND U9608 ( .A(n9585), .B(n9586), .Z(n9367) );
  NANDN U9609 ( .A(n9587), .B(n9588), .Z(n9586) );
  NANDN U9610 ( .A(n9589), .B(n9590), .Z(n9588) );
  NANDN U9611 ( .A(n9590), .B(n9589), .Z(n9585) );
  ANDN U9612 ( .B(B[30]), .A(n70), .Z(n9369) );
  XNOR U9613 ( .A(n9377), .B(n9591), .Z(n9370) );
  XNOR U9614 ( .A(n9376), .B(n9374), .Z(n9591) );
  AND U9615 ( .A(n9592), .B(n9593), .Z(n9374) );
  NANDN U9616 ( .A(n9594), .B(n9595), .Z(n9593) );
  OR U9617 ( .A(n9596), .B(n9597), .Z(n9595) );
  NAND U9618 ( .A(n9597), .B(n9596), .Z(n9592) );
  ANDN U9619 ( .B(B[31]), .A(n71), .Z(n9376) );
  XNOR U9620 ( .A(n9384), .B(n9598), .Z(n9377) );
  XNOR U9621 ( .A(n9383), .B(n9381), .Z(n9598) );
  AND U9622 ( .A(n9599), .B(n9600), .Z(n9381) );
  NANDN U9623 ( .A(n9601), .B(n9602), .Z(n9600) );
  NANDN U9624 ( .A(n9603), .B(n9604), .Z(n9602) );
  NANDN U9625 ( .A(n9604), .B(n9603), .Z(n9599) );
  ANDN U9626 ( .B(B[32]), .A(n72), .Z(n9383) );
  XNOR U9627 ( .A(n9391), .B(n9605), .Z(n9384) );
  XNOR U9628 ( .A(n9390), .B(n9388), .Z(n9605) );
  AND U9629 ( .A(n9606), .B(n9607), .Z(n9388) );
  NANDN U9630 ( .A(n9608), .B(n9609), .Z(n9607) );
  OR U9631 ( .A(n9610), .B(n9611), .Z(n9609) );
  NAND U9632 ( .A(n9611), .B(n9610), .Z(n9606) );
  ANDN U9633 ( .B(B[33]), .A(n73), .Z(n9390) );
  XNOR U9634 ( .A(n9398), .B(n9612), .Z(n9391) );
  XNOR U9635 ( .A(n9397), .B(n9395), .Z(n9612) );
  AND U9636 ( .A(n9613), .B(n9614), .Z(n9395) );
  NANDN U9637 ( .A(n9615), .B(n9616), .Z(n9614) );
  NANDN U9638 ( .A(n9617), .B(n9618), .Z(n9616) );
  NANDN U9639 ( .A(n9618), .B(n9617), .Z(n9613) );
  ANDN U9640 ( .B(B[34]), .A(n74), .Z(n9397) );
  XNOR U9641 ( .A(n9405), .B(n9619), .Z(n9398) );
  XNOR U9642 ( .A(n9404), .B(n9402), .Z(n9619) );
  AND U9643 ( .A(n9620), .B(n9621), .Z(n9402) );
  NANDN U9644 ( .A(n9622), .B(n9623), .Z(n9621) );
  OR U9645 ( .A(n9624), .B(n9625), .Z(n9623) );
  NAND U9646 ( .A(n9625), .B(n9624), .Z(n9620) );
  ANDN U9647 ( .B(B[35]), .A(n75), .Z(n9404) );
  XNOR U9648 ( .A(n9412), .B(n9626), .Z(n9405) );
  XNOR U9649 ( .A(n9411), .B(n9409), .Z(n9626) );
  AND U9650 ( .A(n9627), .B(n9628), .Z(n9409) );
  NANDN U9651 ( .A(n9629), .B(n9630), .Z(n9628) );
  NANDN U9652 ( .A(n9631), .B(n9632), .Z(n9630) );
  NANDN U9653 ( .A(n9632), .B(n9631), .Z(n9627) );
  ANDN U9654 ( .B(B[36]), .A(n76), .Z(n9411) );
  XNOR U9655 ( .A(n9419), .B(n9633), .Z(n9412) );
  XNOR U9656 ( .A(n9418), .B(n9416), .Z(n9633) );
  AND U9657 ( .A(n9634), .B(n9635), .Z(n9416) );
  NANDN U9658 ( .A(n9636), .B(n9637), .Z(n9635) );
  OR U9659 ( .A(n9638), .B(n9639), .Z(n9637) );
  NAND U9660 ( .A(n9639), .B(n9638), .Z(n9634) );
  ANDN U9661 ( .B(B[37]), .A(n77), .Z(n9418) );
  XNOR U9662 ( .A(n9426), .B(n9640), .Z(n9419) );
  XNOR U9663 ( .A(n9425), .B(n9423), .Z(n9640) );
  AND U9664 ( .A(n9641), .B(n9642), .Z(n9423) );
  NANDN U9665 ( .A(n9643), .B(n9644), .Z(n9642) );
  NANDN U9666 ( .A(n9645), .B(n9646), .Z(n9644) );
  NANDN U9667 ( .A(n9646), .B(n9645), .Z(n9641) );
  ANDN U9668 ( .B(B[38]), .A(n78), .Z(n9425) );
  XNOR U9669 ( .A(n9433), .B(n9647), .Z(n9426) );
  XNOR U9670 ( .A(n9432), .B(n9430), .Z(n9647) );
  AND U9671 ( .A(n9648), .B(n9649), .Z(n9430) );
  NANDN U9672 ( .A(n9650), .B(n9651), .Z(n9649) );
  OR U9673 ( .A(n9652), .B(n9653), .Z(n9651) );
  NAND U9674 ( .A(n9653), .B(n9652), .Z(n9648) );
  ANDN U9675 ( .B(B[39]), .A(n79), .Z(n9432) );
  XNOR U9676 ( .A(n9440), .B(n9654), .Z(n9433) );
  XNOR U9677 ( .A(n9439), .B(n9437), .Z(n9654) );
  AND U9678 ( .A(n9655), .B(n9656), .Z(n9437) );
  NANDN U9679 ( .A(n9657), .B(n9658), .Z(n9656) );
  NANDN U9680 ( .A(n9659), .B(n9660), .Z(n9658) );
  NANDN U9681 ( .A(n9660), .B(n9659), .Z(n9655) );
  ANDN U9682 ( .B(B[40]), .A(n80), .Z(n9439) );
  XNOR U9683 ( .A(n9447), .B(n9661), .Z(n9440) );
  XNOR U9684 ( .A(n9446), .B(n9444), .Z(n9661) );
  AND U9685 ( .A(n9662), .B(n9663), .Z(n9444) );
  NANDN U9686 ( .A(n9664), .B(n9665), .Z(n9663) );
  OR U9687 ( .A(n9666), .B(n9667), .Z(n9665) );
  NAND U9688 ( .A(n9667), .B(n9666), .Z(n9662) );
  ANDN U9689 ( .B(B[41]), .A(n81), .Z(n9446) );
  XNOR U9690 ( .A(n9454), .B(n9668), .Z(n9447) );
  XNOR U9691 ( .A(n9453), .B(n9451), .Z(n9668) );
  AND U9692 ( .A(n9669), .B(n9670), .Z(n9451) );
  NANDN U9693 ( .A(n9671), .B(n9672), .Z(n9670) );
  NAND U9694 ( .A(n9673), .B(n9674), .Z(n9672) );
  ANDN U9695 ( .B(B[42]), .A(n82), .Z(n9453) );
  XOR U9696 ( .A(n9460), .B(n9675), .Z(n9454) );
  XNOR U9697 ( .A(n9458), .B(n9461), .Z(n9675) );
  NAND U9698 ( .A(A[2]), .B(B[43]), .Z(n9461) );
  NANDN U9699 ( .A(n9676), .B(n9677), .Z(n9458) );
  AND U9700 ( .A(A[0]), .B(B[44]), .Z(n9677) );
  XNOR U9701 ( .A(n9463), .B(n9678), .Z(n9460) );
  NAND U9702 ( .A(A[0]), .B(B[45]), .Z(n9678) );
  NAND U9703 ( .A(B[44]), .B(A[1]), .Z(n9463) );
  NAND U9704 ( .A(n9679), .B(n9680), .Z(n197) );
  NANDN U9705 ( .A(n9681), .B(n9682), .Z(n9680) );
  OR U9706 ( .A(n9683), .B(n9684), .Z(n9682) );
  NAND U9707 ( .A(n9684), .B(n9683), .Z(n9679) );
  XOR U9708 ( .A(n199), .B(n198), .Z(\A1[42] ) );
  XOR U9709 ( .A(n9684), .B(n9685), .Z(n198) );
  XNOR U9710 ( .A(n9683), .B(n9681), .Z(n9685) );
  AND U9711 ( .A(n9686), .B(n9687), .Z(n9681) );
  NANDN U9712 ( .A(n9688), .B(n9689), .Z(n9687) );
  NANDN U9713 ( .A(n9690), .B(n9691), .Z(n9689) );
  NANDN U9714 ( .A(n9691), .B(n9690), .Z(n9686) );
  ANDN U9715 ( .B(B[13]), .A(n54), .Z(n9683) );
  XNOR U9716 ( .A(n9478), .B(n9692), .Z(n9684) );
  XNOR U9717 ( .A(n9477), .B(n9475), .Z(n9692) );
  AND U9718 ( .A(n9693), .B(n9694), .Z(n9475) );
  NANDN U9719 ( .A(n9695), .B(n9696), .Z(n9694) );
  OR U9720 ( .A(n9697), .B(n9698), .Z(n9696) );
  NAND U9721 ( .A(n9698), .B(n9697), .Z(n9693) );
  ANDN U9722 ( .B(B[14]), .A(n55), .Z(n9477) );
  XNOR U9723 ( .A(n9485), .B(n9699), .Z(n9478) );
  XNOR U9724 ( .A(n9484), .B(n9482), .Z(n9699) );
  AND U9725 ( .A(n9700), .B(n9701), .Z(n9482) );
  NANDN U9726 ( .A(n9702), .B(n9703), .Z(n9701) );
  NANDN U9727 ( .A(n9704), .B(n9705), .Z(n9703) );
  NANDN U9728 ( .A(n9705), .B(n9704), .Z(n9700) );
  ANDN U9729 ( .B(B[15]), .A(n56), .Z(n9484) );
  XNOR U9730 ( .A(n9492), .B(n9706), .Z(n9485) );
  XNOR U9731 ( .A(n9491), .B(n9489), .Z(n9706) );
  AND U9732 ( .A(n9707), .B(n9708), .Z(n9489) );
  NANDN U9733 ( .A(n9709), .B(n9710), .Z(n9708) );
  OR U9734 ( .A(n9711), .B(n9712), .Z(n9710) );
  NAND U9735 ( .A(n9712), .B(n9711), .Z(n9707) );
  ANDN U9736 ( .B(B[16]), .A(n57), .Z(n9491) );
  XNOR U9737 ( .A(n9499), .B(n9713), .Z(n9492) );
  XNOR U9738 ( .A(n9498), .B(n9496), .Z(n9713) );
  AND U9739 ( .A(n9714), .B(n9715), .Z(n9496) );
  NANDN U9740 ( .A(n9716), .B(n9717), .Z(n9715) );
  NANDN U9741 ( .A(n9718), .B(n9719), .Z(n9717) );
  NANDN U9742 ( .A(n9719), .B(n9718), .Z(n9714) );
  ANDN U9743 ( .B(B[17]), .A(n58), .Z(n9498) );
  XNOR U9744 ( .A(n9506), .B(n9720), .Z(n9499) );
  XNOR U9745 ( .A(n9505), .B(n9503), .Z(n9720) );
  AND U9746 ( .A(n9721), .B(n9722), .Z(n9503) );
  NANDN U9747 ( .A(n9723), .B(n9724), .Z(n9722) );
  OR U9748 ( .A(n9725), .B(n9726), .Z(n9724) );
  NAND U9749 ( .A(n9726), .B(n9725), .Z(n9721) );
  ANDN U9750 ( .B(B[18]), .A(n59), .Z(n9505) );
  XNOR U9751 ( .A(n9513), .B(n9727), .Z(n9506) );
  XNOR U9752 ( .A(n9512), .B(n9510), .Z(n9727) );
  AND U9753 ( .A(n9728), .B(n9729), .Z(n9510) );
  NANDN U9754 ( .A(n9730), .B(n9731), .Z(n9729) );
  NANDN U9755 ( .A(n9732), .B(n9733), .Z(n9731) );
  NANDN U9756 ( .A(n9733), .B(n9732), .Z(n9728) );
  ANDN U9757 ( .B(B[19]), .A(n60), .Z(n9512) );
  XNOR U9758 ( .A(n9520), .B(n9734), .Z(n9513) );
  XNOR U9759 ( .A(n9519), .B(n9517), .Z(n9734) );
  AND U9760 ( .A(n9735), .B(n9736), .Z(n9517) );
  NANDN U9761 ( .A(n9737), .B(n9738), .Z(n9736) );
  OR U9762 ( .A(n9739), .B(n9740), .Z(n9738) );
  NAND U9763 ( .A(n9740), .B(n9739), .Z(n9735) );
  ANDN U9764 ( .B(B[20]), .A(n61), .Z(n9519) );
  XNOR U9765 ( .A(n9527), .B(n9741), .Z(n9520) );
  XNOR U9766 ( .A(n9526), .B(n9524), .Z(n9741) );
  AND U9767 ( .A(n9742), .B(n9743), .Z(n9524) );
  NANDN U9768 ( .A(n9744), .B(n9745), .Z(n9743) );
  NANDN U9769 ( .A(n9746), .B(n9747), .Z(n9745) );
  NANDN U9770 ( .A(n9747), .B(n9746), .Z(n9742) );
  ANDN U9771 ( .B(B[21]), .A(n62), .Z(n9526) );
  XNOR U9772 ( .A(n9534), .B(n9748), .Z(n9527) );
  XNOR U9773 ( .A(n9533), .B(n9531), .Z(n9748) );
  AND U9774 ( .A(n9749), .B(n9750), .Z(n9531) );
  NANDN U9775 ( .A(n9751), .B(n9752), .Z(n9750) );
  OR U9776 ( .A(n9753), .B(n9754), .Z(n9752) );
  NAND U9777 ( .A(n9754), .B(n9753), .Z(n9749) );
  ANDN U9778 ( .B(B[22]), .A(n63), .Z(n9533) );
  XNOR U9779 ( .A(n9541), .B(n9755), .Z(n9534) );
  XNOR U9780 ( .A(n9540), .B(n9538), .Z(n9755) );
  AND U9781 ( .A(n9756), .B(n9757), .Z(n9538) );
  NANDN U9782 ( .A(n9758), .B(n9759), .Z(n9757) );
  NANDN U9783 ( .A(n9760), .B(n9761), .Z(n9759) );
  NANDN U9784 ( .A(n9761), .B(n9760), .Z(n9756) );
  ANDN U9785 ( .B(B[23]), .A(n64), .Z(n9540) );
  XNOR U9786 ( .A(n9548), .B(n9762), .Z(n9541) );
  XNOR U9787 ( .A(n9547), .B(n9545), .Z(n9762) );
  AND U9788 ( .A(n9763), .B(n9764), .Z(n9545) );
  NANDN U9789 ( .A(n9765), .B(n9766), .Z(n9764) );
  OR U9790 ( .A(n9767), .B(n9768), .Z(n9766) );
  NAND U9791 ( .A(n9768), .B(n9767), .Z(n9763) );
  ANDN U9792 ( .B(B[24]), .A(n65), .Z(n9547) );
  XNOR U9793 ( .A(n9555), .B(n9769), .Z(n9548) );
  XNOR U9794 ( .A(n9554), .B(n9552), .Z(n9769) );
  AND U9795 ( .A(n9770), .B(n9771), .Z(n9552) );
  NANDN U9796 ( .A(n9772), .B(n9773), .Z(n9771) );
  NANDN U9797 ( .A(n9774), .B(n9775), .Z(n9773) );
  NANDN U9798 ( .A(n9775), .B(n9774), .Z(n9770) );
  ANDN U9799 ( .B(B[25]), .A(n66), .Z(n9554) );
  XNOR U9800 ( .A(n9562), .B(n9776), .Z(n9555) );
  XNOR U9801 ( .A(n9561), .B(n9559), .Z(n9776) );
  AND U9802 ( .A(n9777), .B(n9778), .Z(n9559) );
  NANDN U9803 ( .A(n9779), .B(n9780), .Z(n9778) );
  OR U9804 ( .A(n9781), .B(n9782), .Z(n9780) );
  NAND U9805 ( .A(n9782), .B(n9781), .Z(n9777) );
  ANDN U9806 ( .B(B[26]), .A(n67), .Z(n9561) );
  XNOR U9807 ( .A(n9569), .B(n9783), .Z(n9562) );
  XNOR U9808 ( .A(n9568), .B(n9566), .Z(n9783) );
  AND U9809 ( .A(n9784), .B(n9785), .Z(n9566) );
  NANDN U9810 ( .A(n9786), .B(n9787), .Z(n9785) );
  NANDN U9811 ( .A(n9788), .B(n9789), .Z(n9787) );
  NANDN U9812 ( .A(n9789), .B(n9788), .Z(n9784) );
  ANDN U9813 ( .B(B[27]), .A(n68), .Z(n9568) );
  XNOR U9814 ( .A(n9576), .B(n9790), .Z(n9569) );
  XNOR U9815 ( .A(n9575), .B(n9573), .Z(n9790) );
  AND U9816 ( .A(n9791), .B(n9792), .Z(n9573) );
  NANDN U9817 ( .A(n9793), .B(n9794), .Z(n9792) );
  OR U9818 ( .A(n9795), .B(n9796), .Z(n9794) );
  NAND U9819 ( .A(n9796), .B(n9795), .Z(n9791) );
  ANDN U9820 ( .B(B[28]), .A(n69), .Z(n9575) );
  XNOR U9821 ( .A(n9583), .B(n9797), .Z(n9576) );
  XNOR U9822 ( .A(n9582), .B(n9580), .Z(n9797) );
  AND U9823 ( .A(n9798), .B(n9799), .Z(n9580) );
  NANDN U9824 ( .A(n9800), .B(n9801), .Z(n9799) );
  NANDN U9825 ( .A(n9802), .B(n9803), .Z(n9801) );
  NANDN U9826 ( .A(n9803), .B(n9802), .Z(n9798) );
  ANDN U9827 ( .B(B[29]), .A(n70), .Z(n9582) );
  XNOR U9828 ( .A(n9590), .B(n9804), .Z(n9583) );
  XNOR U9829 ( .A(n9589), .B(n9587), .Z(n9804) );
  AND U9830 ( .A(n9805), .B(n9806), .Z(n9587) );
  NANDN U9831 ( .A(n9807), .B(n9808), .Z(n9806) );
  OR U9832 ( .A(n9809), .B(n9810), .Z(n9808) );
  NAND U9833 ( .A(n9810), .B(n9809), .Z(n9805) );
  ANDN U9834 ( .B(B[30]), .A(n71), .Z(n9589) );
  XNOR U9835 ( .A(n9597), .B(n9811), .Z(n9590) );
  XNOR U9836 ( .A(n9596), .B(n9594), .Z(n9811) );
  AND U9837 ( .A(n9812), .B(n9813), .Z(n9594) );
  NANDN U9838 ( .A(n9814), .B(n9815), .Z(n9813) );
  NANDN U9839 ( .A(n9816), .B(n9817), .Z(n9815) );
  NANDN U9840 ( .A(n9817), .B(n9816), .Z(n9812) );
  ANDN U9841 ( .B(B[31]), .A(n72), .Z(n9596) );
  XNOR U9842 ( .A(n9604), .B(n9818), .Z(n9597) );
  XNOR U9843 ( .A(n9603), .B(n9601), .Z(n9818) );
  AND U9844 ( .A(n9819), .B(n9820), .Z(n9601) );
  NANDN U9845 ( .A(n9821), .B(n9822), .Z(n9820) );
  OR U9846 ( .A(n9823), .B(n9824), .Z(n9822) );
  NAND U9847 ( .A(n9824), .B(n9823), .Z(n9819) );
  ANDN U9848 ( .B(B[32]), .A(n73), .Z(n9603) );
  XNOR U9849 ( .A(n9611), .B(n9825), .Z(n9604) );
  XNOR U9850 ( .A(n9610), .B(n9608), .Z(n9825) );
  AND U9851 ( .A(n9826), .B(n9827), .Z(n9608) );
  NANDN U9852 ( .A(n9828), .B(n9829), .Z(n9827) );
  NANDN U9853 ( .A(n9830), .B(n9831), .Z(n9829) );
  NANDN U9854 ( .A(n9831), .B(n9830), .Z(n9826) );
  ANDN U9855 ( .B(B[33]), .A(n74), .Z(n9610) );
  XNOR U9856 ( .A(n9618), .B(n9832), .Z(n9611) );
  XNOR U9857 ( .A(n9617), .B(n9615), .Z(n9832) );
  AND U9858 ( .A(n9833), .B(n9834), .Z(n9615) );
  NANDN U9859 ( .A(n9835), .B(n9836), .Z(n9834) );
  OR U9860 ( .A(n9837), .B(n9838), .Z(n9836) );
  NAND U9861 ( .A(n9838), .B(n9837), .Z(n9833) );
  ANDN U9862 ( .B(B[34]), .A(n75), .Z(n9617) );
  XNOR U9863 ( .A(n9625), .B(n9839), .Z(n9618) );
  XNOR U9864 ( .A(n9624), .B(n9622), .Z(n9839) );
  AND U9865 ( .A(n9840), .B(n9841), .Z(n9622) );
  NANDN U9866 ( .A(n9842), .B(n9843), .Z(n9841) );
  NANDN U9867 ( .A(n9844), .B(n9845), .Z(n9843) );
  NANDN U9868 ( .A(n9845), .B(n9844), .Z(n9840) );
  ANDN U9869 ( .B(B[35]), .A(n76), .Z(n9624) );
  XNOR U9870 ( .A(n9632), .B(n9846), .Z(n9625) );
  XNOR U9871 ( .A(n9631), .B(n9629), .Z(n9846) );
  AND U9872 ( .A(n9847), .B(n9848), .Z(n9629) );
  NANDN U9873 ( .A(n9849), .B(n9850), .Z(n9848) );
  OR U9874 ( .A(n9851), .B(n9852), .Z(n9850) );
  NAND U9875 ( .A(n9852), .B(n9851), .Z(n9847) );
  ANDN U9876 ( .B(B[36]), .A(n77), .Z(n9631) );
  XNOR U9877 ( .A(n9639), .B(n9853), .Z(n9632) );
  XNOR U9878 ( .A(n9638), .B(n9636), .Z(n9853) );
  AND U9879 ( .A(n9854), .B(n9855), .Z(n9636) );
  NANDN U9880 ( .A(n9856), .B(n9857), .Z(n9855) );
  NANDN U9881 ( .A(n9858), .B(n9859), .Z(n9857) );
  NANDN U9882 ( .A(n9859), .B(n9858), .Z(n9854) );
  ANDN U9883 ( .B(B[37]), .A(n78), .Z(n9638) );
  XNOR U9884 ( .A(n9646), .B(n9860), .Z(n9639) );
  XNOR U9885 ( .A(n9645), .B(n9643), .Z(n9860) );
  AND U9886 ( .A(n9861), .B(n9862), .Z(n9643) );
  NANDN U9887 ( .A(n9863), .B(n9864), .Z(n9862) );
  OR U9888 ( .A(n9865), .B(n9866), .Z(n9864) );
  NAND U9889 ( .A(n9866), .B(n9865), .Z(n9861) );
  ANDN U9890 ( .B(B[38]), .A(n79), .Z(n9645) );
  XNOR U9891 ( .A(n9653), .B(n9867), .Z(n9646) );
  XNOR U9892 ( .A(n9652), .B(n9650), .Z(n9867) );
  AND U9893 ( .A(n9868), .B(n9869), .Z(n9650) );
  NANDN U9894 ( .A(n9870), .B(n9871), .Z(n9869) );
  NANDN U9895 ( .A(n9872), .B(n9873), .Z(n9871) );
  NANDN U9896 ( .A(n9873), .B(n9872), .Z(n9868) );
  ANDN U9897 ( .B(B[39]), .A(n80), .Z(n9652) );
  XNOR U9898 ( .A(n9660), .B(n9874), .Z(n9653) );
  XNOR U9899 ( .A(n9659), .B(n9657), .Z(n9874) );
  AND U9900 ( .A(n9875), .B(n9876), .Z(n9657) );
  NANDN U9901 ( .A(n9877), .B(n9878), .Z(n9876) );
  OR U9902 ( .A(n9879), .B(n9880), .Z(n9878) );
  NAND U9903 ( .A(n9880), .B(n9879), .Z(n9875) );
  ANDN U9904 ( .B(B[40]), .A(n81), .Z(n9659) );
  XNOR U9905 ( .A(n9667), .B(n9881), .Z(n9660) );
  XNOR U9906 ( .A(n9666), .B(n9664), .Z(n9881) );
  AND U9907 ( .A(n9882), .B(n9883), .Z(n9664) );
  NANDN U9908 ( .A(n9884), .B(n9885), .Z(n9883) );
  NAND U9909 ( .A(n9886), .B(n9887), .Z(n9885) );
  ANDN U9910 ( .B(B[41]), .A(n82), .Z(n9666) );
  XOR U9911 ( .A(n9673), .B(n9888), .Z(n9667) );
  XNOR U9912 ( .A(n9671), .B(n9674), .Z(n9888) );
  NAND U9913 ( .A(A[2]), .B(B[42]), .Z(n9674) );
  NANDN U9914 ( .A(n9889), .B(n9890), .Z(n9671) );
  AND U9915 ( .A(A[0]), .B(B[43]), .Z(n9890) );
  XNOR U9916 ( .A(n9676), .B(n9891), .Z(n9673) );
  NAND U9917 ( .A(A[0]), .B(B[44]), .Z(n9891) );
  NAND U9918 ( .A(B[43]), .B(A[1]), .Z(n9676) );
  NAND U9919 ( .A(n9892), .B(n9893), .Z(n199) );
  NANDN U9920 ( .A(n9894), .B(n9895), .Z(n9893) );
  OR U9921 ( .A(n9896), .B(n9897), .Z(n9895) );
  NAND U9922 ( .A(n9897), .B(n9896), .Z(n9892) );
  XOR U9923 ( .A(n201), .B(n200), .Z(\A1[41] ) );
  XOR U9924 ( .A(n9897), .B(n9898), .Z(n200) );
  XNOR U9925 ( .A(n9896), .B(n9894), .Z(n9898) );
  AND U9926 ( .A(n9899), .B(n9900), .Z(n9894) );
  NANDN U9927 ( .A(n9901), .B(n9902), .Z(n9900) );
  NANDN U9928 ( .A(n9903), .B(n9904), .Z(n9902) );
  NANDN U9929 ( .A(n9904), .B(n9903), .Z(n9899) );
  ANDN U9930 ( .B(B[12]), .A(n54), .Z(n9896) );
  XNOR U9931 ( .A(n9691), .B(n9905), .Z(n9897) );
  XNOR U9932 ( .A(n9690), .B(n9688), .Z(n9905) );
  AND U9933 ( .A(n9906), .B(n9907), .Z(n9688) );
  NANDN U9934 ( .A(n9908), .B(n9909), .Z(n9907) );
  OR U9935 ( .A(n9910), .B(n9911), .Z(n9909) );
  NAND U9936 ( .A(n9911), .B(n9910), .Z(n9906) );
  ANDN U9937 ( .B(B[13]), .A(n55), .Z(n9690) );
  XNOR U9938 ( .A(n9698), .B(n9912), .Z(n9691) );
  XNOR U9939 ( .A(n9697), .B(n9695), .Z(n9912) );
  AND U9940 ( .A(n9913), .B(n9914), .Z(n9695) );
  NANDN U9941 ( .A(n9915), .B(n9916), .Z(n9914) );
  NANDN U9942 ( .A(n9917), .B(n9918), .Z(n9916) );
  NANDN U9943 ( .A(n9918), .B(n9917), .Z(n9913) );
  ANDN U9944 ( .B(B[14]), .A(n56), .Z(n9697) );
  XNOR U9945 ( .A(n9705), .B(n9919), .Z(n9698) );
  XNOR U9946 ( .A(n9704), .B(n9702), .Z(n9919) );
  AND U9947 ( .A(n9920), .B(n9921), .Z(n9702) );
  NANDN U9948 ( .A(n9922), .B(n9923), .Z(n9921) );
  OR U9949 ( .A(n9924), .B(n9925), .Z(n9923) );
  NAND U9950 ( .A(n9925), .B(n9924), .Z(n9920) );
  ANDN U9951 ( .B(B[15]), .A(n57), .Z(n9704) );
  XNOR U9952 ( .A(n9712), .B(n9926), .Z(n9705) );
  XNOR U9953 ( .A(n9711), .B(n9709), .Z(n9926) );
  AND U9954 ( .A(n9927), .B(n9928), .Z(n9709) );
  NANDN U9955 ( .A(n9929), .B(n9930), .Z(n9928) );
  NANDN U9956 ( .A(n9931), .B(n9932), .Z(n9930) );
  NANDN U9957 ( .A(n9932), .B(n9931), .Z(n9927) );
  ANDN U9958 ( .B(B[16]), .A(n58), .Z(n9711) );
  XNOR U9959 ( .A(n9719), .B(n9933), .Z(n9712) );
  XNOR U9960 ( .A(n9718), .B(n9716), .Z(n9933) );
  AND U9961 ( .A(n9934), .B(n9935), .Z(n9716) );
  NANDN U9962 ( .A(n9936), .B(n9937), .Z(n9935) );
  OR U9963 ( .A(n9938), .B(n9939), .Z(n9937) );
  NAND U9964 ( .A(n9939), .B(n9938), .Z(n9934) );
  ANDN U9965 ( .B(B[17]), .A(n59), .Z(n9718) );
  XNOR U9966 ( .A(n9726), .B(n9940), .Z(n9719) );
  XNOR U9967 ( .A(n9725), .B(n9723), .Z(n9940) );
  AND U9968 ( .A(n9941), .B(n9942), .Z(n9723) );
  NANDN U9969 ( .A(n9943), .B(n9944), .Z(n9942) );
  NANDN U9970 ( .A(n9945), .B(n9946), .Z(n9944) );
  NANDN U9971 ( .A(n9946), .B(n9945), .Z(n9941) );
  ANDN U9972 ( .B(B[18]), .A(n60), .Z(n9725) );
  XNOR U9973 ( .A(n9733), .B(n9947), .Z(n9726) );
  XNOR U9974 ( .A(n9732), .B(n9730), .Z(n9947) );
  AND U9975 ( .A(n9948), .B(n9949), .Z(n9730) );
  NANDN U9976 ( .A(n9950), .B(n9951), .Z(n9949) );
  OR U9977 ( .A(n9952), .B(n9953), .Z(n9951) );
  NAND U9978 ( .A(n9953), .B(n9952), .Z(n9948) );
  ANDN U9979 ( .B(B[19]), .A(n61), .Z(n9732) );
  XNOR U9980 ( .A(n9740), .B(n9954), .Z(n9733) );
  XNOR U9981 ( .A(n9739), .B(n9737), .Z(n9954) );
  AND U9982 ( .A(n9955), .B(n9956), .Z(n9737) );
  NANDN U9983 ( .A(n9957), .B(n9958), .Z(n9956) );
  NANDN U9984 ( .A(n9959), .B(n9960), .Z(n9958) );
  NANDN U9985 ( .A(n9960), .B(n9959), .Z(n9955) );
  ANDN U9986 ( .B(B[20]), .A(n62), .Z(n9739) );
  XNOR U9987 ( .A(n9747), .B(n9961), .Z(n9740) );
  XNOR U9988 ( .A(n9746), .B(n9744), .Z(n9961) );
  AND U9989 ( .A(n9962), .B(n9963), .Z(n9744) );
  NANDN U9990 ( .A(n9964), .B(n9965), .Z(n9963) );
  OR U9991 ( .A(n9966), .B(n9967), .Z(n9965) );
  NAND U9992 ( .A(n9967), .B(n9966), .Z(n9962) );
  ANDN U9993 ( .B(B[21]), .A(n63), .Z(n9746) );
  XNOR U9994 ( .A(n9754), .B(n9968), .Z(n9747) );
  XNOR U9995 ( .A(n9753), .B(n9751), .Z(n9968) );
  AND U9996 ( .A(n9969), .B(n9970), .Z(n9751) );
  NANDN U9997 ( .A(n9971), .B(n9972), .Z(n9970) );
  NANDN U9998 ( .A(n9973), .B(n9974), .Z(n9972) );
  NANDN U9999 ( .A(n9974), .B(n9973), .Z(n9969) );
  ANDN U10000 ( .B(B[22]), .A(n64), .Z(n9753) );
  XNOR U10001 ( .A(n9761), .B(n9975), .Z(n9754) );
  XNOR U10002 ( .A(n9760), .B(n9758), .Z(n9975) );
  AND U10003 ( .A(n9976), .B(n9977), .Z(n9758) );
  NANDN U10004 ( .A(n9978), .B(n9979), .Z(n9977) );
  OR U10005 ( .A(n9980), .B(n9981), .Z(n9979) );
  NAND U10006 ( .A(n9981), .B(n9980), .Z(n9976) );
  ANDN U10007 ( .B(B[23]), .A(n65), .Z(n9760) );
  XNOR U10008 ( .A(n9768), .B(n9982), .Z(n9761) );
  XNOR U10009 ( .A(n9767), .B(n9765), .Z(n9982) );
  AND U10010 ( .A(n9983), .B(n9984), .Z(n9765) );
  NANDN U10011 ( .A(n9985), .B(n9986), .Z(n9984) );
  NANDN U10012 ( .A(n9987), .B(n9988), .Z(n9986) );
  NANDN U10013 ( .A(n9988), .B(n9987), .Z(n9983) );
  ANDN U10014 ( .B(B[24]), .A(n66), .Z(n9767) );
  XNOR U10015 ( .A(n9775), .B(n9989), .Z(n9768) );
  XNOR U10016 ( .A(n9774), .B(n9772), .Z(n9989) );
  AND U10017 ( .A(n9990), .B(n9991), .Z(n9772) );
  NANDN U10018 ( .A(n9992), .B(n9993), .Z(n9991) );
  OR U10019 ( .A(n9994), .B(n9995), .Z(n9993) );
  NAND U10020 ( .A(n9995), .B(n9994), .Z(n9990) );
  ANDN U10021 ( .B(B[25]), .A(n67), .Z(n9774) );
  XNOR U10022 ( .A(n9782), .B(n9996), .Z(n9775) );
  XNOR U10023 ( .A(n9781), .B(n9779), .Z(n9996) );
  AND U10024 ( .A(n9997), .B(n9998), .Z(n9779) );
  NANDN U10025 ( .A(n9999), .B(n10000), .Z(n9998) );
  NANDN U10026 ( .A(n10001), .B(n10002), .Z(n10000) );
  NANDN U10027 ( .A(n10002), .B(n10001), .Z(n9997) );
  ANDN U10028 ( .B(B[26]), .A(n68), .Z(n9781) );
  XNOR U10029 ( .A(n9789), .B(n10003), .Z(n9782) );
  XNOR U10030 ( .A(n9788), .B(n9786), .Z(n10003) );
  AND U10031 ( .A(n10004), .B(n10005), .Z(n9786) );
  NANDN U10032 ( .A(n10006), .B(n10007), .Z(n10005) );
  OR U10033 ( .A(n10008), .B(n10009), .Z(n10007) );
  NAND U10034 ( .A(n10009), .B(n10008), .Z(n10004) );
  ANDN U10035 ( .B(B[27]), .A(n69), .Z(n9788) );
  XNOR U10036 ( .A(n9796), .B(n10010), .Z(n9789) );
  XNOR U10037 ( .A(n9795), .B(n9793), .Z(n10010) );
  AND U10038 ( .A(n10011), .B(n10012), .Z(n9793) );
  NANDN U10039 ( .A(n10013), .B(n10014), .Z(n10012) );
  NANDN U10040 ( .A(n10015), .B(n10016), .Z(n10014) );
  NANDN U10041 ( .A(n10016), .B(n10015), .Z(n10011) );
  ANDN U10042 ( .B(B[28]), .A(n70), .Z(n9795) );
  XNOR U10043 ( .A(n9803), .B(n10017), .Z(n9796) );
  XNOR U10044 ( .A(n9802), .B(n9800), .Z(n10017) );
  AND U10045 ( .A(n10018), .B(n10019), .Z(n9800) );
  NANDN U10046 ( .A(n10020), .B(n10021), .Z(n10019) );
  OR U10047 ( .A(n10022), .B(n10023), .Z(n10021) );
  NAND U10048 ( .A(n10023), .B(n10022), .Z(n10018) );
  ANDN U10049 ( .B(B[29]), .A(n71), .Z(n9802) );
  XNOR U10050 ( .A(n9810), .B(n10024), .Z(n9803) );
  XNOR U10051 ( .A(n9809), .B(n9807), .Z(n10024) );
  AND U10052 ( .A(n10025), .B(n10026), .Z(n9807) );
  NANDN U10053 ( .A(n10027), .B(n10028), .Z(n10026) );
  NANDN U10054 ( .A(n10029), .B(n10030), .Z(n10028) );
  NANDN U10055 ( .A(n10030), .B(n10029), .Z(n10025) );
  ANDN U10056 ( .B(B[30]), .A(n72), .Z(n9809) );
  XNOR U10057 ( .A(n9817), .B(n10031), .Z(n9810) );
  XNOR U10058 ( .A(n9816), .B(n9814), .Z(n10031) );
  AND U10059 ( .A(n10032), .B(n10033), .Z(n9814) );
  NANDN U10060 ( .A(n10034), .B(n10035), .Z(n10033) );
  OR U10061 ( .A(n10036), .B(n10037), .Z(n10035) );
  NAND U10062 ( .A(n10037), .B(n10036), .Z(n10032) );
  ANDN U10063 ( .B(B[31]), .A(n73), .Z(n9816) );
  XNOR U10064 ( .A(n9824), .B(n10038), .Z(n9817) );
  XNOR U10065 ( .A(n9823), .B(n9821), .Z(n10038) );
  AND U10066 ( .A(n10039), .B(n10040), .Z(n9821) );
  NANDN U10067 ( .A(n10041), .B(n10042), .Z(n10040) );
  NANDN U10068 ( .A(n10043), .B(n10044), .Z(n10042) );
  NANDN U10069 ( .A(n10044), .B(n10043), .Z(n10039) );
  ANDN U10070 ( .B(B[32]), .A(n74), .Z(n9823) );
  XNOR U10071 ( .A(n9831), .B(n10045), .Z(n9824) );
  XNOR U10072 ( .A(n9830), .B(n9828), .Z(n10045) );
  AND U10073 ( .A(n10046), .B(n10047), .Z(n9828) );
  NANDN U10074 ( .A(n10048), .B(n10049), .Z(n10047) );
  OR U10075 ( .A(n10050), .B(n10051), .Z(n10049) );
  NAND U10076 ( .A(n10051), .B(n10050), .Z(n10046) );
  ANDN U10077 ( .B(B[33]), .A(n75), .Z(n9830) );
  XNOR U10078 ( .A(n9838), .B(n10052), .Z(n9831) );
  XNOR U10079 ( .A(n9837), .B(n9835), .Z(n10052) );
  AND U10080 ( .A(n10053), .B(n10054), .Z(n9835) );
  NANDN U10081 ( .A(n10055), .B(n10056), .Z(n10054) );
  NANDN U10082 ( .A(n10057), .B(n10058), .Z(n10056) );
  NANDN U10083 ( .A(n10058), .B(n10057), .Z(n10053) );
  ANDN U10084 ( .B(B[34]), .A(n76), .Z(n9837) );
  XNOR U10085 ( .A(n9845), .B(n10059), .Z(n9838) );
  XNOR U10086 ( .A(n9844), .B(n9842), .Z(n10059) );
  AND U10087 ( .A(n10060), .B(n10061), .Z(n9842) );
  NANDN U10088 ( .A(n10062), .B(n10063), .Z(n10061) );
  OR U10089 ( .A(n10064), .B(n10065), .Z(n10063) );
  NAND U10090 ( .A(n10065), .B(n10064), .Z(n10060) );
  ANDN U10091 ( .B(B[35]), .A(n77), .Z(n9844) );
  XNOR U10092 ( .A(n9852), .B(n10066), .Z(n9845) );
  XNOR U10093 ( .A(n9851), .B(n9849), .Z(n10066) );
  AND U10094 ( .A(n10067), .B(n10068), .Z(n9849) );
  NANDN U10095 ( .A(n10069), .B(n10070), .Z(n10068) );
  NANDN U10096 ( .A(n10071), .B(n10072), .Z(n10070) );
  NANDN U10097 ( .A(n10072), .B(n10071), .Z(n10067) );
  ANDN U10098 ( .B(B[36]), .A(n78), .Z(n9851) );
  XNOR U10099 ( .A(n9859), .B(n10073), .Z(n9852) );
  XNOR U10100 ( .A(n9858), .B(n9856), .Z(n10073) );
  AND U10101 ( .A(n10074), .B(n10075), .Z(n9856) );
  NANDN U10102 ( .A(n10076), .B(n10077), .Z(n10075) );
  OR U10103 ( .A(n10078), .B(n10079), .Z(n10077) );
  NAND U10104 ( .A(n10079), .B(n10078), .Z(n10074) );
  ANDN U10105 ( .B(B[37]), .A(n79), .Z(n9858) );
  XNOR U10106 ( .A(n9866), .B(n10080), .Z(n9859) );
  XNOR U10107 ( .A(n9865), .B(n9863), .Z(n10080) );
  AND U10108 ( .A(n10081), .B(n10082), .Z(n9863) );
  NANDN U10109 ( .A(n10083), .B(n10084), .Z(n10082) );
  NANDN U10110 ( .A(n10085), .B(n10086), .Z(n10084) );
  NANDN U10111 ( .A(n10086), .B(n10085), .Z(n10081) );
  ANDN U10112 ( .B(B[38]), .A(n80), .Z(n9865) );
  XNOR U10113 ( .A(n9873), .B(n10087), .Z(n9866) );
  XNOR U10114 ( .A(n9872), .B(n9870), .Z(n10087) );
  AND U10115 ( .A(n10088), .B(n10089), .Z(n9870) );
  NANDN U10116 ( .A(n10090), .B(n10091), .Z(n10089) );
  OR U10117 ( .A(n10092), .B(n10093), .Z(n10091) );
  NAND U10118 ( .A(n10093), .B(n10092), .Z(n10088) );
  ANDN U10119 ( .B(B[39]), .A(n81), .Z(n9872) );
  XNOR U10120 ( .A(n9880), .B(n10094), .Z(n9873) );
  XNOR U10121 ( .A(n9879), .B(n9877), .Z(n10094) );
  AND U10122 ( .A(n10095), .B(n10096), .Z(n9877) );
  NANDN U10123 ( .A(n10097), .B(n10098), .Z(n10096) );
  NAND U10124 ( .A(n10099), .B(n10100), .Z(n10098) );
  ANDN U10125 ( .B(B[40]), .A(n82), .Z(n9879) );
  XOR U10126 ( .A(n9886), .B(n10101), .Z(n9880) );
  XNOR U10127 ( .A(n9884), .B(n9887), .Z(n10101) );
  NAND U10128 ( .A(A[2]), .B(B[41]), .Z(n9887) );
  NANDN U10129 ( .A(n10102), .B(n10103), .Z(n9884) );
  AND U10130 ( .A(A[0]), .B(B[42]), .Z(n10103) );
  XNOR U10131 ( .A(n9889), .B(n10104), .Z(n9886) );
  NAND U10132 ( .A(A[0]), .B(B[43]), .Z(n10104) );
  NAND U10133 ( .A(B[42]), .B(A[1]), .Z(n9889) );
  NAND U10134 ( .A(n10105), .B(n10106), .Z(n201) );
  NANDN U10135 ( .A(n10107), .B(n10108), .Z(n10106) );
  OR U10136 ( .A(n10109), .B(n10110), .Z(n10108) );
  NAND U10137 ( .A(n10110), .B(n10109), .Z(n10105) );
  XOR U10138 ( .A(n203), .B(n202), .Z(\A1[40] ) );
  XOR U10139 ( .A(n10110), .B(n10111), .Z(n202) );
  XNOR U10140 ( .A(n10109), .B(n10107), .Z(n10111) );
  AND U10141 ( .A(n10112), .B(n10113), .Z(n10107) );
  NANDN U10142 ( .A(n10114), .B(n10115), .Z(n10113) );
  NANDN U10143 ( .A(n10116), .B(n10117), .Z(n10115) );
  NANDN U10144 ( .A(n10117), .B(n10116), .Z(n10112) );
  ANDN U10145 ( .B(B[11]), .A(n54), .Z(n10109) );
  XNOR U10146 ( .A(n9904), .B(n10118), .Z(n10110) );
  XNOR U10147 ( .A(n9903), .B(n9901), .Z(n10118) );
  AND U10148 ( .A(n10119), .B(n10120), .Z(n9901) );
  NANDN U10149 ( .A(n10121), .B(n10122), .Z(n10120) );
  OR U10150 ( .A(n10123), .B(n10124), .Z(n10122) );
  NAND U10151 ( .A(n10124), .B(n10123), .Z(n10119) );
  ANDN U10152 ( .B(B[12]), .A(n55), .Z(n9903) );
  XNOR U10153 ( .A(n9911), .B(n10125), .Z(n9904) );
  XNOR U10154 ( .A(n9910), .B(n9908), .Z(n10125) );
  AND U10155 ( .A(n10126), .B(n10127), .Z(n9908) );
  NANDN U10156 ( .A(n10128), .B(n10129), .Z(n10127) );
  NANDN U10157 ( .A(n10130), .B(n10131), .Z(n10129) );
  NANDN U10158 ( .A(n10131), .B(n10130), .Z(n10126) );
  ANDN U10159 ( .B(B[13]), .A(n56), .Z(n9910) );
  XNOR U10160 ( .A(n9918), .B(n10132), .Z(n9911) );
  XNOR U10161 ( .A(n9917), .B(n9915), .Z(n10132) );
  AND U10162 ( .A(n10133), .B(n10134), .Z(n9915) );
  NANDN U10163 ( .A(n10135), .B(n10136), .Z(n10134) );
  OR U10164 ( .A(n10137), .B(n10138), .Z(n10136) );
  NAND U10165 ( .A(n10138), .B(n10137), .Z(n10133) );
  ANDN U10166 ( .B(B[14]), .A(n57), .Z(n9917) );
  XNOR U10167 ( .A(n9925), .B(n10139), .Z(n9918) );
  XNOR U10168 ( .A(n9924), .B(n9922), .Z(n10139) );
  AND U10169 ( .A(n10140), .B(n10141), .Z(n9922) );
  NANDN U10170 ( .A(n10142), .B(n10143), .Z(n10141) );
  NANDN U10171 ( .A(n10144), .B(n10145), .Z(n10143) );
  NANDN U10172 ( .A(n10145), .B(n10144), .Z(n10140) );
  ANDN U10173 ( .B(B[15]), .A(n58), .Z(n9924) );
  XNOR U10174 ( .A(n9932), .B(n10146), .Z(n9925) );
  XNOR U10175 ( .A(n9931), .B(n9929), .Z(n10146) );
  AND U10176 ( .A(n10147), .B(n10148), .Z(n9929) );
  NANDN U10177 ( .A(n10149), .B(n10150), .Z(n10148) );
  OR U10178 ( .A(n10151), .B(n10152), .Z(n10150) );
  NAND U10179 ( .A(n10152), .B(n10151), .Z(n10147) );
  ANDN U10180 ( .B(B[16]), .A(n59), .Z(n9931) );
  XNOR U10181 ( .A(n9939), .B(n10153), .Z(n9932) );
  XNOR U10182 ( .A(n9938), .B(n9936), .Z(n10153) );
  AND U10183 ( .A(n10154), .B(n10155), .Z(n9936) );
  NANDN U10184 ( .A(n10156), .B(n10157), .Z(n10155) );
  NANDN U10185 ( .A(n10158), .B(n10159), .Z(n10157) );
  NANDN U10186 ( .A(n10159), .B(n10158), .Z(n10154) );
  ANDN U10187 ( .B(B[17]), .A(n60), .Z(n9938) );
  XNOR U10188 ( .A(n9946), .B(n10160), .Z(n9939) );
  XNOR U10189 ( .A(n9945), .B(n9943), .Z(n10160) );
  AND U10190 ( .A(n10161), .B(n10162), .Z(n9943) );
  NANDN U10191 ( .A(n10163), .B(n10164), .Z(n10162) );
  OR U10192 ( .A(n10165), .B(n10166), .Z(n10164) );
  NAND U10193 ( .A(n10166), .B(n10165), .Z(n10161) );
  ANDN U10194 ( .B(B[18]), .A(n61), .Z(n9945) );
  XNOR U10195 ( .A(n9953), .B(n10167), .Z(n9946) );
  XNOR U10196 ( .A(n9952), .B(n9950), .Z(n10167) );
  AND U10197 ( .A(n10168), .B(n10169), .Z(n9950) );
  NANDN U10198 ( .A(n10170), .B(n10171), .Z(n10169) );
  NANDN U10199 ( .A(n10172), .B(n10173), .Z(n10171) );
  NANDN U10200 ( .A(n10173), .B(n10172), .Z(n10168) );
  ANDN U10201 ( .B(B[19]), .A(n62), .Z(n9952) );
  XNOR U10202 ( .A(n9960), .B(n10174), .Z(n9953) );
  XNOR U10203 ( .A(n9959), .B(n9957), .Z(n10174) );
  AND U10204 ( .A(n10175), .B(n10176), .Z(n9957) );
  NANDN U10205 ( .A(n10177), .B(n10178), .Z(n10176) );
  OR U10206 ( .A(n10179), .B(n10180), .Z(n10178) );
  NAND U10207 ( .A(n10180), .B(n10179), .Z(n10175) );
  ANDN U10208 ( .B(B[20]), .A(n63), .Z(n9959) );
  XNOR U10209 ( .A(n9967), .B(n10181), .Z(n9960) );
  XNOR U10210 ( .A(n9966), .B(n9964), .Z(n10181) );
  AND U10211 ( .A(n10182), .B(n10183), .Z(n9964) );
  NANDN U10212 ( .A(n10184), .B(n10185), .Z(n10183) );
  NANDN U10213 ( .A(n10186), .B(n10187), .Z(n10185) );
  NANDN U10214 ( .A(n10187), .B(n10186), .Z(n10182) );
  ANDN U10215 ( .B(B[21]), .A(n64), .Z(n9966) );
  XNOR U10216 ( .A(n9974), .B(n10188), .Z(n9967) );
  XNOR U10217 ( .A(n9973), .B(n9971), .Z(n10188) );
  AND U10218 ( .A(n10189), .B(n10190), .Z(n9971) );
  NANDN U10219 ( .A(n10191), .B(n10192), .Z(n10190) );
  OR U10220 ( .A(n10193), .B(n10194), .Z(n10192) );
  NAND U10221 ( .A(n10194), .B(n10193), .Z(n10189) );
  ANDN U10222 ( .B(B[22]), .A(n65), .Z(n9973) );
  XNOR U10223 ( .A(n9981), .B(n10195), .Z(n9974) );
  XNOR U10224 ( .A(n9980), .B(n9978), .Z(n10195) );
  AND U10225 ( .A(n10196), .B(n10197), .Z(n9978) );
  NANDN U10226 ( .A(n10198), .B(n10199), .Z(n10197) );
  NANDN U10227 ( .A(n10200), .B(n10201), .Z(n10199) );
  NANDN U10228 ( .A(n10201), .B(n10200), .Z(n10196) );
  ANDN U10229 ( .B(B[23]), .A(n66), .Z(n9980) );
  XNOR U10230 ( .A(n9988), .B(n10202), .Z(n9981) );
  XNOR U10231 ( .A(n9987), .B(n9985), .Z(n10202) );
  AND U10232 ( .A(n10203), .B(n10204), .Z(n9985) );
  NANDN U10233 ( .A(n10205), .B(n10206), .Z(n10204) );
  OR U10234 ( .A(n10207), .B(n10208), .Z(n10206) );
  NAND U10235 ( .A(n10208), .B(n10207), .Z(n10203) );
  ANDN U10236 ( .B(B[24]), .A(n67), .Z(n9987) );
  XNOR U10237 ( .A(n9995), .B(n10209), .Z(n9988) );
  XNOR U10238 ( .A(n9994), .B(n9992), .Z(n10209) );
  AND U10239 ( .A(n10210), .B(n10211), .Z(n9992) );
  NANDN U10240 ( .A(n10212), .B(n10213), .Z(n10211) );
  NANDN U10241 ( .A(n10214), .B(n10215), .Z(n10213) );
  NANDN U10242 ( .A(n10215), .B(n10214), .Z(n10210) );
  ANDN U10243 ( .B(B[25]), .A(n68), .Z(n9994) );
  XNOR U10244 ( .A(n10002), .B(n10216), .Z(n9995) );
  XNOR U10245 ( .A(n10001), .B(n9999), .Z(n10216) );
  AND U10246 ( .A(n10217), .B(n10218), .Z(n9999) );
  NANDN U10247 ( .A(n10219), .B(n10220), .Z(n10218) );
  OR U10248 ( .A(n10221), .B(n10222), .Z(n10220) );
  NAND U10249 ( .A(n10222), .B(n10221), .Z(n10217) );
  ANDN U10250 ( .B(B[26]), .A(n69), .Z(n10001) );
  XNOR U10251 ( .A(n10009), .B(n10223), .Z(n10002) );
  XNOR U10252 ( .A(n10008), .B(n10006), .Z(n10223) );
  AND U10253 ( .A(n10224), .B(n10225), .Z(n10006) );
  NANDN U10254 ( .A(n10226), .B(n10227), .Z(n10225) );
  NANDN U10255 ( .A(n10228), .B(n10229), .Z(n10227) );
  NANDN U10256 ( .A(n10229), .B(n10228), .Z(n10224) );
  ANDN U10257 ( .B(B[27]), .A(n70), .Z(n10008) );
  XNOR U10258 ( .A(n10016), .B(n10230), .Z(n10009) );
  XNOR U10259 ( .A(n10015), .B(n10013), .Z(n10230) );
  AND U10260 ( .A(n10231), .B(n10232), .Z(n10013) );
  NANDN U10261 ( .A(n10233), .B(n10234), .Z(n10232) );
  OR U10262 ( .A(n10235), .B(n10236), .Z(n10234) );
  NAND U10263 ( .A(n10236), .B(n10235), .Z(n10231) );
  ANDN U10264 ( .B(B[28]), .A(n71), .Z(n10015) );
  XNOR U10265 ( .A(n10023), .B(n10237), .Z(n10016) );
  XNOR U10266 ( .A(n10022), .B(n10020), .Z(n10237) );
  AND U10267 ( .A(n10238), .B(n10239), .Z(n10020) );
  NANDN U10268 ( .A(n10240), .B(n10241), .Z(n10239) );
  NANDN U10269 ( .A(n10242), .B(n10243), .Z(n10241) );
  NANDN U10270 ( .A(n10243), .B(n10242), .Z(n10238) );
  ANDN U10271 ( .B(B[29]), .A(n72), .Z(n10022) );
  XNOR U10272 ( .A(n10030), .B(n10244), .Z(n10023) );
  XNOR U10273 ( .A(n10029), .B(n10027), .Z(n10244) );
  AND U10274 ( .A(n10245), .B(n10246), .Z(n10027) );
  NANDN U10275 ( .A(n10247), .B(n10248), .Z(n10246) );
  OR U10276 ( .A(n10249), .B(n10250), .Z(n10248) );
  NAND U10277 ( .A(n10250), .B(n10249), .Z(n10245) );
  ANDN U10278 ( .B(B[30]), .A(n73), .Z(n10029) );
  XNOR U10279 ( .A(n10037), .B(n10251), .Z(n10030) );
  XNOR U10280 ( .A(n10036), .B(n10034), .Z(n10251) );
  AND U10281 ( .A(n10252), .B(n10253), .Z(n10034) );
  NANDN U10282 ( .A(n10254), .B(n10255), .Z(n10253) );
  NANDN U10283 ( .A(n10256), .B(n10257), .Z(n10255) );
  NANDN U10284 ( .A(n10257), .B(n10256), .Z(n10252) );
  ANDN U10285 ( .B(B[31]), .A(n74), .Z(n10036) );
  XNOR U10286 ( .A(n10044), .B(n10258), .Z(n10037) );
  XNOR U10287 ( .A(n10043), .B(n10041), .Z(n10258) );
  AND U10288 ( .A(n10259), .B(n10260), .Z(n10041) );
  NANDN U10289 ( .A(n10261), .B(n10262), .Z(n10260) );
  OR U10290 ( .A(n10263), .B(n10264), .Z(n10262) );
  NAND U10291 ( .A(n10264), .B(n10263), .Z(n10259) );
  ANDN U10292 ( .B(B[32]), .A(n75), .Z(n10043) );
  XNOR U10293 ( .A(n10051), .B(n10265), .Z(n10044) );
  XNOR U10294 ( .A(n10050), .B(n10048), .Z(n10265) );
  AND U10295 ( .A(n10266), .B(n10267), .Z(n10048) );
  NANDN U10296 ( .A(n10268), .B(n10269), .Z(n10267) );
  NANDN U10297 ( .A(n10270), .B(n10271), .Z(n10269) );
  NANDN U10298 ( .A(n10271), .B(n10270), .Z(n10266) );
  ANDN U10299 ( .B(B[33]), .A(n76), .Z(n10050) );
  XNOR U10300 ( .A(n10058), .B(n10272), .Z(n10051) );
  XNOR U10301 ( .A(n10057), .B(n10055), .Z(n10272) );
  AND U10302 ( .A(n10273), .B(n10274), .Z(n10055) );
  NANDN U10303 ( .A(n10275), .B(n10276), .Z(n10274) );
  OR U10304 ( .A(n10277), .B(n10278), .Z(n10276) );
  NAND U10305 ( .A(n10278), .B(n10277), .Z(n10273) );
  ANDN U10306 ( .B(B[34]), .A(n77), .Z(n10057) );
  XNOR U10307 ( .A(n10065), .B(n10279), .Z(n10058) );
  XNOR U10308 ( .A(n10064), .B(n10062), .Z(n10279) );
  AND U10309 ( .A(n10280), .B(n10281), .Z(n10062) );
  NANDN U10310 ( .A(n10282), .B(n10283), .Z(n10281) );
  NANDN U10311 ( .A(n10284), .B(n10285), .Z(n10283) );
  NANDN U10312 ( .A(n10285), .B(n10284), .Z(n10280) );
  ANDN U10313 ( .B(B[35]), .A(n78), .Z(n10064) );
  XNOR U10314 ( .A(n10072), .B(n10286), .Z(n10065) );
  XNOR U10315 ( .A(n10071), .B(n10069), .Z(n10286) );
  AND U10316 ( .A(n10287), .B(n10288), .Z(n10069) );
  NANDN U10317 ( .A(n10289), .B(n10290), .Z(n10288) );
  OR U10318 ( .A(n10291), .B(n10292), .Z(n10290) );
  NAND U10319 ( .A(n10292), .B(n10291), .Z(n10287) );
  ANDN U10320 ( .B(B[36]), .A(n79), .Z(n10071) );
  XNOR U10321 ( .A(n10079), .B(n10293), .Z(n10072) );
  XNOR U10322 ( .A(n10078), .B(n10076), .Z(n10293) );
  AND U10323 ( .A(n10294), .B(n10295), .Z(n10076) );
  NANDN U10324 ( .A(n10296), .B(n10297), .Z(n10295) );
  NANDN U10325 ( .A(n10298), .B(n10299), .Z(n10297) );
  NANDN U10326 ( .A(n10299), .B(n10298), .Z(n10294) );
  ANDN U10327 ( .B(B[37]), .A(n80), .Z(n10078) );
  XNOR U10328 ( .A(n10086), .B(n10300), .Z(n10079) );
  XNOR U10329 ( .A(n10085), .B(n10083), .Z(n10300) );
  AND U10330 ( .A(n10301), .B(n10302), .Z(n10083) );
  NANDN U10331 ( .A(n10303), .B(n10304), .Z(n10302) );
  OR U10332 ( .A(n10305), .B(n10306), .Z(n10304) );
  NAND U10333 ( .A(n10306), .B(n10305), .Z(n10301) );
  ANDN U10334 ( .B(B[38]), .A(n81), .Z(n10085) );
  XNOR U10335 ( .A(n10093), .B(n10307), .Z(n10086) );
  XNOR U10336 ( .A(n10092), .B(n10090), .Z(n10307) );
  AND U10337 ( .A(n10308), .B(n10309), .Z(n10090) );
  NANDN U10338 ( .A(n10310), .B(n10311), .Z(n10309) );
  NAND U10339 ( .A(n10312), .B(n10313), .Z(n10311) );
  ANDN U10340 ( .B(B[39]), .A(n82), .Z(n10092) );
  XOR U10341 ( .A(n10099), .B(n10314), .Z(n10093) );
  XNOR U10342 ( .A(n10097), .B(n10100), .Z(n10314) );
  NAND U10343 ( .A(A[2]), .B(B[40]), .Z(n10100) );
  NANDN U10344 ( .A(n10315), .B(n10316), .Z(n10097) );
  AND U10345 ( .A(A[0]), .B(B[41]), .Z(n10316) );
  XNOR U10346 ( .A(n10102), .B(n10317), .Z(n10099) );
  NAND U10347 ( .A(A[0]), .B(B[42]), .Z(n10317) );
  NAND U10348 ( .A(B[41]), .B(A[1]), .Z(n10102) );
  NAND U10349 ( .A(n10318), .B(n10319), .Z(n203) );
  NANDN U10350 ( .A(n10320), .B(n10321), .Z(n10319) );
  OR U10351 ( .A(n10322), .B(n10323), .Z(n10321) );
  NAND U10352 ( .A(n10323), .B(n10322), .Z(n10318) );
  XOR U10353 ( .A(n10324), .B(n10325), .Z(\A1[3] ) );
  XNOR U10354 ( .A(n10326), .B(n52), .Z(n10325) );
  XOR U10355 ( .A(n205), .B(n204), .Z(\A1[39] ) );
  XOR U10356 ( .A(n10323), .B(n10327), .Z(n204) );
  XNOR U10357 ( .A(n10322), .B(n10320), .Z(n10327) );
  AND U10358 ( .A(n10328), .B(n10329), .Z(n10320) );
  NANDN U10359 ( .A(n10330), .B(n10331), .Z(n10329) );
  NANDN U10360 ( .A(n10332), .B(n10333), .Z(n10331) );
  NANDN U10361 ( .A(n10333), .B(n10332), .Z(n10328) );
  ANDN U10362 ( .B(B[10]), .A(n54), .Z(n10322) );
  XNOR U10363 ( .A(n10117), .B(n10334), .Z(n10323) );
  XNOR U10364 ( .A(n10116), .B(n10114), .Z(n10334) );
  AND U10365 ( .A(n10335), .B(n10336), .Z(n10114) );
  NANDN U10366 ( .A(n10337), .B(n10338), .Z(n10336) );
  OR U10367 ( .A(n10339), .B(n10340), .Z(n10338) );
  NAND U10368 ( .A(n10340), .B(n10339), .Z(n10335) );
  ANDN U10369 ( .B(B[11]), .A(n55), .Z(n10116) );
  XNOR U10370 ( .A(n10124), .B(n10341), .Z(n10117) );
  XNOR U10371 ( .A(n10123), .B(n10121), .Z(n10341) );
  AND U10372 ( .A(n10342), .B(n10343), .Z(n10121) );
  NANDN U10373 ( .A(n10344), .B(n10345), .Z(n10343) );
  NANDN U10374 ( .A(n10346), .B(n10347), .Z(n10345) );
  NANDN U10375 ( .A(n10347), .B(n10346), .Z(n10342) );
  ANDN U10376 ( .B(B[12]), .A(n56), .Z(n10123) );
  XNOR U10377 ( .A(n10131), .B(n10348), .Z(n10124) );
  XNOR U10378 ( .A(n10130), .B(n10128), .Z(n10348) );
  AND U10379 ( .A(n10349), .B(n10350), .Z(n10128) );
  NANDN U10380 ( .A(n10351), .B(n10352), .Z(n10350) );
  OR U10381 ( .A(n10353), .B(n10354), .Z(n10352) );
  NAND U10382 ( .A(n10354), .B(n10353), .Z(n10349) );
  ANDN U10383 ( .B(B[13]), .A(n57), .Z(n10130) );
  XNOR U10384 ( .A(n10138), .B(n10355), .Z(n10131) );
  XNOR U10385 ( .A(n10137), .B(n10135), .Z(n10355) );
  AND U10386 ( .A(n10356), .B(n10357), .Z(n10135) );
  NANDN U10387 ( .A(n10358), .B(n10359), .Z(n10357) );
  NANDN U10388 ( .A(n10360), .B(n10361), .Z(n10359) );
  NANDN U10389 ( .A(n10361), .B(n10360), .Z(n10356) );
  ANDN U10390 ( .B(B[14]), .A(n58), .Z(n10137) );
  XNOR U10391 ( .A(n10145), .B(n10362), .Z(n10138) );
  XNOR U10392 ( .A(n10144), .B(n10142), .Z(n10362) );
  AND U10393 ( .A(n10363), .B(n10364), .Z(n10142) );
  NANDN U10394 ( .A(n10365), .B(n10366), .Z(n10364) );
  OR U10395 ( .A(n10367), .B(n10368), .Z(n10366) );
  NAND U10396 ( .A(n10368), .B(n10367), .Z(n10363) );
  ANDN U10397 ( .B(B[15]), .A(n59), .Z(n10144) );
  XNOR U10398 ( .A(n10152), .B(n10369), .Z(n10145) );
  XNOR U10399 ( .A(n10151), .B(n10149), .Z(n10369) );
  AND U10400 ( .A(n10370), .B(n10371), .Z(n10149) );
  NANDN U10401 ( .A(n10372), .B(n10373), .Z(n10371) );
  NANDN U10402 ( .A(n10374), .B(n10375), .Z(n10373) );
  NANDN U10403 ( .A(n10375), .B(n10374), .Z(n10370) );
  ANDN U10404 ( .B(B[16]), .A(n60), .Z(n10151) );
  XNOR U10405 ( .A(n10159), .B(n10376), .Z(n10152) );
  XNOR U10406 ( .A(n10158), .B(n10156), .Z(n10376) );
  AND U10407 ( .A(n10377), .B(n10378), .Z(n10156) );
  NANDN U10408 ( .A(n10379), .B(n10380), .Z(n10378) );
  OR U10409 ( .A(n10381), .B(n10382), .Z(n10380) );
  NAND U10410 ( .A(n10382), .B(n10381), .Z(n10377) );
  ANDN U10411 ( .B(B[17]), .A(n61), .Z(n10158) );
  XNOR U10412 ( .A(n10166), .B(n10383), .Z(n10159) );
  XNOR U10413 ( .A(n10165), .B(n10163), .Z(n10383) );
  AND U10414 ( .A(n10384), .B(n10385), .Z(n10163) );
  NANDN U10415 ( .A(n10386), .B(n10387), .Z(n10385) );
  NANDN U10416 ( .A(n10388), .B(n10389), .Z(n10387) );
  NANDN U10417 ( .A(n10389), .B(n10388), .Z(n10384) );
  ANDN U10418 ( .B(B[18]), .A(n62), .Z(n10165) );
  XNOR U10419 ( .A(n10173), .B(n10390), .Z(n10166) );
  XNOR U10420 ( .A(n10172), .B(n10170), .Z(n10390) );
  AND U10421 ( .A(n10391), .B(n10392), .Z(n10170) );
  NANDN U10422 ( .A(n10393), .B(n10394), .Z(n10392) );
  OR U10423 ( .A(n10395), .B(n10396), .Z(n10394) );
  NAND U10424 ( .A(n10396), .B(n10395), .Z(n10391) );
  ANDN U10425 ( .B(B[19]), .A(n63), .Z(n10172) );
  XNOR U10426 ( .A(n10180), .B(n10397), .Z(n10173) );
  XNOR U10427 ( .A(n10179), .B(n10177), .Z(n10397) );
  AND U10428 ( .A(n10398), .B(n10399), .Z(n10177) );
  NANDN U10429 ( .A(n10400), .B(n10401), .Z(n10399) );
  NANDN U10430 ( .A(n10402), .B(n10403), .Z(n10401) );
  NANDN U10431 ( .A(n10403), .B(n10402), .Z(n10398) );
  ANDN U10432 ( .B(B[20]), .A(n64), .Z(n10179) );
  XNOR U10433 ( .A(n10187), .B(n10404), .Z(n10180) );
  XNOR U10434 ( .A(n10186), .B(n10184), .Z(n10404) );
  AND U10435 ( .A(n10405), .B(n10406), .Z(n10184) );
  NANDN U10436 ( .A(n10407), .B(n10408), .Z(n10406) );
  OR U10437 ( .A(n10409), .B(n10410), .Z(n10408) );
  NAND U10438 ( .A(n10410), .B(n10409), .Z(n10405) );
  ANDN U10439 ( .B(B[21]), .A(n65), .Z(n10186) );
  XNOR U10440 ( .A(n10194), .B(n10411), .Z(n10187) );
  XNOR U10441 ( .A(n10193), .B(n10191), .Z(n10411) );
  AND U10442 ( .A(n10412), .B(n10413), .Z(n10191) );
  NANDN U10443 ( .A(n10414), .B(n10415), .Z(n10413) );
  NANDN U10444 ( .A(n10416), .B(n10417), .Z(n10415) );
  NANDN U10445 ( .A(n10417), .B(n10416), .Z(n10412) );
  ANDN U10446 ( .B(B[22]), .A(n66), .Z(n10193) );
  XNOR U10447 ( .A(n10201), .B(n10418), .Z(n10194) );
  XNOR U10448 ( .A(n10200), .B(n10198), .Z(n10418) );
  AND U10449 ( .A(n10419), .B(n10420), .Z(n10198) );
  NANDN U10450 ( .A(n10421), .B(n10422), .Z(n10420) );
  OR U10451 ( .A(n10423), .B(n10424), .Z(n10422) );
  NAND U10452 ( .A(n10424), .B(n10423), .Z(n10419) );
  ANDN U10453 ( .B(B[23]), .A(n67), .Z(n10200) );
  XNOR U10454 ( .A(n10208), .B(n10425), .Z(n10201) );
  XNOR U10455 ( .A(n10207), .B(n10205), .Z(n10425) );
  AND U10456 ( .A(n10426), .B(n10427), .Z(n10205) );
  NANDN U10457 ( .A(n10428), .B(n10429), .Z(n10427) );
  NANDN U10458 ( .A(n10430), .B(n10431), .Z(n10429) );
  NANDN U10459 ( .A(n10431), .B(n10430), .Z(n10426) );
  ANDN U10460 ( .B(B[24]), .A(n68), .Z(n10207) );
  XNOR U10461 ( .A(n10215), .B(n10432), .Z(n10208) );
  XNOR U10462 ( .A(n10214), .B(n10212), .Z(n10432) );
  AND U10463 ( .A(n10433), .B(n10434), .Z(n10212) );
  NANDN U10464 ( .A(n10435), .B(n10436), .Z(n10434) );
  OR U10465 ( .A(n10437), .B(n10438), .Z(n10436) );
  NAND U10466 ( .A(n10438), .B(n10437), .Z(n10433) );
  ANDN U10467 ( .B(B[25]), .A(n69), .Z(n10214) );
  XNOR U10468 ( .A(n10222), .B(n10439), .Z(n10215) );
  XNOR U10469 ( .A(n10221), .B(n10219), .Z(n10439) );
  AND U10470 ( .A(n10440), .B(n10441), .Z(n10219) );
  NANDN U10471 ( .A(n10442), .B(n10443), .Z(n10441) );
  NANDN U10472 ( .A(n10444), .B(n10445), .Z(n10443) );
  NANDN U10473 ( .A(n10445), .B(n10444), .Z(n10440) );
  ANDN U10474 ( .B(B[26]), .A(n70), .Z(n10221) );
  XNOR U10475 ( .A(n10229), .B(n10446), .Z(n10222) );
  XNOR U10476 ( .A(n10228), .B(n10226), .Z(n10446) );
  AND U10477 ( .A(n10447), .B(n10448), .Z(n10226) );
  NANDN U10478 ( .A(n10449), .B(n10450), .Z(n10448) );
  OR U10479 ( .A(n10451), .B(n10452), .Z(n10450) );
  NAND U10480 ( .A(n10452), .B(n10451), .Z(n10447) );
  ANDN U10481 ( .B(B[27]), .A(n71), .Z(n10228) );
  XNOR U10482 ( .A(n10236), .B(n10453), .Z(n10229) );
  XNOR U10483 ( .A(n10235), .B(n10233), .Z(n10453) );
  AND U10484 ( .A(n10454), .B(n10455), .Z(n10233) );
  NANDN U10485 ( .A(n10456), .B(n10457), .Z(n10455) );
  NANDN U10486 ( .A(n10458), .B(n10459), .Z(n10457) );
  NANDN U10487 ( .A(n10459), .B(n10458), .Z(n10454) );
  ANDN U10488 ( .B(B[28]), .A(n72), .Z(n10235) );
  XNOR U10489 ( .A(n10243), .B(n10460), .Z(n10236) );
  XNOR U10490 ( .A(n10242), .B(n10240), .Z(n10460) );
  AND U10491 ( .A(n10461), .B(n10462), .Z(n10240) );
  NANDN U10492 ( .A(n10463), .B(n10464), .Z(n10462) );
  OR U10493 ( .A(n10465), .B(n10466), .Z(n10464) );
  NAND U10494 ( .A(n10466), .B(n10465), .Z(n10461) );
  ANDN U10495 ( .B(B[29]), .A(n73), .Z(n10242) );
  XNOR U10496 ( .A(n10250), .B(n10467), .Z(n10243) );
  XNOR U10497 ( .A(n10249), .B(n10247), .Z(n10467) );
  AND U10498 ( .A(n10468), .B(n10469), .Z(n10247) );
  NANDN U10499 ( .A(n10470), .B(n10471), .Z(n10469) );
  NANDN U10500 ( .A(n10472), .B(n10473), .Z(n10471) );
  NANDN U10501 ( .A(n10473), .B(n10472), .Z(n10468) );
  ANDN U10502 ( .B(B[30]), .A(n74), .Z(n10249) );
  XNOR U10503 ( .A(n10257), .B(n10474), .Z(n10250) );
  XNOR U10504 ( .A(n10256), .B(n10254), .Z(n10474) );
  AND U10505 ( .A(n10475), .B(n10476), .Z(n10254) );
  NANDN U10506 ( .A(n10477), .B(n10478), .Z(n10476) );
  OR U10507 ( .A(n10479), .B(n10480), .Z(n10478) );
  NAND U10508 ( .A(n10480), .B(n10479), .Z(n10475) );
  ANDN U10509 ( .B(B[31]), .A(n75), .Z(n10256) );
  XNOR U10510 ( .A(n10264), .B(n10481), .Z(n10257) );
  XNOR U10511 ( .A(n10263), .B(n10261), .Z(n10481) );
  AND U10512 ( .A(n10482), .B(n10483), .Z(n10261) );
  NANDN U10513 ( .A(n10484), .B(n10485), .Z(n10483) );
  NANDN U10514 ( .A(n10486), .B(n10487), .Z(n10485) );
  NANDN U10515 ( .A(n10487), .B(n10486), .Z(n10482) );
  ANDN U10516 ( .B(B[32]), .A(n76), .Z(n10263) );
  XNOR U10517 ( .A(n10271), .B(n10488), .Z(n10264) );
  XNOR U10518 ( .A(n10270), .B(n10268), .Z(n10488) );
  AND U10519 ( .A(n10489), .B(n10490), .Z(n10268) );
  NANDN U10520 ( .A(n10491), .B(n10492), .Z(n10490) );
  OR U10521 ( .A(n10493), .B(n10494), .Z(n10492) );
  NAND U10522 ( .A(n10494), .B(n10493), .Z(n10489) );
  ANDN U10523 ( .B(B[33]), .A(n77), .Z(n10270) );
  XNOR U10524 ( .A(n10278), .B(n10495), .Z(n10271) );
  XNOR U10525 ( .A(n10277), .B(n10275), .Z(n10495) );
  AND U10526 ( .A(n10496), .B(n10497), .Z(n10275) );
  NANDN U10527 ( .A(n10498), .B(n10499), .Z(n10497) );
  NANDN U10528 ( .A(n10500), .B(n10501), .Z(n10499) );
  NANDN U10529 ( .A(n10501), .B(n10500), .Z(n10496) );
  ANDN U10530 ( .B(B[34]), .A(n78), .Z(n10277) );
  XNOR U10531 ( .A(n10285), .B(n10502), .Z(n10278) );
  XNOR U10532 ( .A(n10284), .B(n10282), .Z(n10502) );
  AND U10533 ( .A(n10503), .B(n10504), .Z(n10282) );
  NANDN U10534 ( .A(n10505), .B(n10506), .Z(n10504) );
  OR U10535 ( .A(n10507), .B(n10508), .Z(n10506) );
  NAND U10536 ( .A(n10508), .B(n10507), .Z(n10503) );
  ANDN U10537 ( .B(B[35]), .A(n79), .Z(n10284) );
  XNOR U10538 ( .A(n10292), .B(n10509), .Z(n10285) );
  XNOR U10539 ( .A(n10291), .B(n10289), .Z(n10509) );
  AND U10540 ( .A(n10510), .B(n10511), .Z(n10289) );
  NANDN U10541 ( .A(n10512), .B(n10513), .Z(n10511) );
  NANDN U10542 ( .A(n10514), .B(n10515), .Z(n10513) );
  NANDN U10543 ( .A(n10515), .B(n10514), .Z(n10510) );
  ANDN U10544 ( .B(B[36]), .A(n80), .Z(n10291) );
  XNOR U10545 ( .A(n10299), .B(n10516), .Z(n10292) );
  XNOR U10546 ( .A(n10298), .B(n10296), .Z(n10516) );
  AND U10547 ( .A(n10517), .B(n10518), .Z(n10296) );
  NANDN U10548 ( .A(n10519), .B(n10520), .Z(n10518) );
  OR U10549 ( .A(n10521), .B(n10522), .Z(n10520) );
  NAND U10550 ( .A(n10522), .B(n10521), .Z(n10517) );
  ANDN U10551 ( .B(B[37]), .A(n81), .Z(n10298) );
  XNOR U10552 ( .A(n10306), .B(n10523), .Z(n10299) );
  XNOR U10553 ( .A(n10305), .B(n10303), .Z(n10523) );
  AND U10554 ( .A(n10524), .B(n10525), .Z(n10303) );
  NANDN U10555 ( .A(n10526), .B(n10527), .Z(n10525) );
  NAND U10556 ( .A(n10528), .B(n10529), .Z(n10527) );
  ANDN U10557 ( .B(B[38]), .A(n82), .Z(n10305) );
  XOR U10558 ( .A(n10312), .B(n10530), .Z(n10306) );
  XNOR U10559 ( .A(n10310), .B(n10313), .Z(n10530) );
  NAND U10560 ( .A(A[2]), .B(B[39]), .Z(n10313) );
  NANDN U10561 ( .A(n10531), .B(n10532), .Z(n10310) );
  AND U10562 ( .A(A[0]), .B(B[40]), .Z(n10532) );
  XNOR U10563 ( .A(n10315), .B(n10533), .Z(n10312) );
  NAND U10564 ( .A(A[0]), .B(B[41]), .Z(n10533) );
  NAND U10565 ( .A(B[40]), .B(A[1]), .Z(n10315) );
  NAND U10566 ( .A(n10534), .B(n10535), .Z(n205) );
  NANDN U10567 ( .A(n10536), .B(n10537), .Z(n10535) );
  OR U10568 ( .A(n10538), .B(n10539), .Z(n10537) );
  NAND U10569 ( .A(n10539), .B(n10538), .Z(n10534) );
  XOR U10570 ( .A(n207), .B(n206), .Z(\A1[38] ) );
  XOR U10571 ( .A(n10539), .B(n10540), .Z(n206) );
  XNOR U10572 ( .A(n10538), .B(n10536), .Z(n10540) );
  AND U10573 ( .A(n10541), .B(n10542), .Z(n10536) );
  NANDN U10574 ( .A(n10543), .B(n10544), .Z(n10542) );
  NANDN U10575 ( .A(n10545), .B(n10546), .Z(n10544) );
  NANDN U10576 ( .A(n10546), .B(n10545), .Z(n10541) );
  ANDN U10577 ( .B(B[9]), .A(n54), .Z(n10538) );
  XNOR U10578 ( .A(n10333), .B(n10547), .Z(n10539) );
  XNOR U10579 ( .A(n10332), .B(n10330), .Z(n10547) );
  AND U10580 ( .A(n10548), .B(n10549), .Z(n10330) );
  NANDN U10581 ( .A(n10550), .B(n10551), .Z(n10549) );
  OR U10582 ( .A(n10552), .B(n10553), .Z(n10551) );
  NAND U10583 ( .A(n10553), .B(n10552), .Z(n10548) );
  ANDN U10584 ( .B(B[10]), .A(n55), .Z(n10332) );
  XNOR U10585 ( .A(n10340), .B(n10554), .Z(n10333) );
  XNOR U10586 ( .A(n10339), .B(n10337), .Z(n10554) );
  AND U10587 ( .A(n10555), .B(n10556), .Z(n10337) );
  NANDN U10588 ( .A(n10557), .B(n10558), .Z(n10556) );
  NANDN U10589 ( .A(n10559), .B(n10560), .Z(n10558) );
  NANDN U10590 ( .A(n10560), .B(n10559), .Z(n10555) );
  ANDN U10591 ( .B(B[11]), .A(n56), .Z(n10339) );
  XNOR U10592 ( .A(n10347), .B(n10561), .Z(n10340) );
  XNOR U10593 ( .A(n10346), .B(n10344), .Z(n10561) );
  AND U10594 ( .A(n10562), .B(n10563), .Z(n10344) );
  NANDN U10595 ( .A(n10564), .B(n10565), .Z(n10563) );
  OR U10596 ( .A(n10566), .B(n10567), .Z(n10565) );
  NAND U10597 ( .A(n10567), .B(n10566), .Z(n10562) );
  ANDN U10598 ( .B(B[12]), .A(n57), .Z(n10346) );
  XNOR U10599 ( .A(n10354), .B(n10568), .Z(n10347) );
  XNOR U10600 ( .A(n10353), .B(n10351), .Z(n10568) );
  AND U10601 ( .A(n10569), .B(n10570), .Z(n10351) );
  NANDN U10602 ( .A(n10571), .B(n10572), .Z(n10570) );
  NANDN U10603 ( .A(n10573), .B(n10574), .Z(n10572) );
  NANDN U10604 ( .A(n10574), .B(n10573), .Z(n10569) );
  ANDN U10605 ( .B(B[13]), .A(n58), .Z(n10353) );
  XNOR U10606 ( .A(n10361), .B(n10575), .Z(n10354) );
  XNOR U10607 ( .A(n10360), .B(n10358), .Z(n10575) );
  AND U10608 ( .A(n10576), .B(n10577), .Z(n10358) );
  NANDN U10609 ( .A(n10578), .B(n10579), .Z(n10577) );
  OR U10610 ( .A(n10580), .B(n10581), .Z(n10579) );
  NAND U10611 ( .A(n10581), .B(n10580), .Z(n10576) );
  ANDN U10612 ( .B(B[14]), .A(n59), .Z(n10360) );
  XNOR U10613 ( .A(n10368), .B(n10582), .Z(n10361) );
  XNOR U10614 ( .A(n10367), .B(n10365), .Z(n10582) );
  AND U10615 ( .A(n10583), .B(n10584), .Z(n10365) );
  NANDN U10616 ( .A(n10585), .B(n10586), .Z(n10584) );
  NANDN U10617 ( .A(n10587), .B(n10588), .Z(n10586) );
  NANDN U10618 ( .A(n10588), .B(n10587), .Z(n10583) );
  ANDN U10619 ( .B(B[15]), .A(n60), .Z(n10367) );
  XNOR U10620 ( .A(n10375), .B(n10589), .Z(n10368) );
  XNOR U10621 ( .A(n10374), .B(n10372), .Z(n10589) );
  AND U10622 ( .A(n10590), .B(n10591), .Z(n10372) );
  NANDN U10623 ( .A(n10592), .B(n10593), .Z(n10591) );
  OR U10624 ( .A(n10594), .B(n10595), .Z(n10593) );
  NAND U10625 ( .A(n10595), .B(n10594), .Z(n10590) );
  ANDN U10626 ( .B(B[16]), .A(n61), .Z(n10374) );
  XNOR U10627 ( .A(n10382), .B(n10596), .Z(n10375) );
  XNOR U10628 ( .A(n10381), .B(n10379), .Z(n10596) );
  AND U10629 ( .A(n10597), .B(n10598), .Z(n10379) );
  NANDN U10630 ( .A(n10599), .B(n10600), .Z(n10598) );
  NANDN U10631 ( .A(n10601), .B(n10602), .Z(n10600) );
  NANDN U10632 ( .A(n10602), .B(n10601), .Z(n10597) );
  ANDN U10633 ( .B(B[17]), .A(n62), .Z(n10381) );
  XNOR U10634 ( .A(n10389), .B(n10603), .Z(n10382) );
  XNOR U10635 ( .A(n10388), .B(n10386), .Z(n10603) );
  AND U10636 ( .A(n10604), .B(n10605), .Z(n10386) );
  NANDN U10637 ( .A(n10606), .B(n10607), .Z(n10605) );
  OR U10638 ( .A(n10608), .B(n10609), .Z(n10607) );
  NAND U10639 ( .A(n10609), .B(n10608), .Z(n10604) );
  ANDN U10640 ( .B(B[18]), .A(n63), .Z(n10388) );
  XNOR U10641 ( .A(n10396), .B(n10610), .Z(n10389) );
  XNOR U10642 ( .A(n10395), .B(n10393), .Z(n10610) );
  AND U10643 ( .A(n10611), .B(n10612), .Z(n10393) );
  NANDN U10644 ( .A(n10613), .B(n10614), .Z(n10612) );
  NANDN U10645 ( .A(n10615), .B(n10616), .Z(n10614) );
  NANDN U10646 ( .A(n10616), .B(n10615), .Z(n10611) );
  ANDN U10647 ( .B(B[19]), .A(n64), .Z(n10395) );
  XNOR U10648 ( .A(n10403), .B(n10617), .Z(n10396) );
  XNOR U10649 ( .A(n10402), .B(n10400), .Z(n10617) );
  AND U10650 ( .A(n10618), .B(n10619), .Z(n10400) );
  NANDN U10651 ( .A(n10620), .B(n10621), .Z(n10619) );
  OR U10652 ( .A(n10622), .B(n10623), .Z(n10621) );
  NAND U10653 ( .A(n10623), .B(n10622), .Z(n10618) );
  ANDN U10654 ( .B(B[20]), .A(n65), .Z(n10402) );
  XNOR U10655 ( .A(n10410), .B(n10624), .Z(n10403) );
  XNOR U10656 ( .A(n10409), .B(n10407), .Z(n10624) );
  AND U10657 ( .A(n10625), .B(n10626), .Z(n10407) );
  NANDN U10658 ( .A(n10627), .B(n10628), .Z(n10626) );
  NANDN U10659 ( .A(n10629), .B(n10630), .Z(n10628) );
  NANDN U10660 ( .A(n10630), .B(n10629), .Z(n10625) );
  ANDN U10661 ( .B(B[21]), .A(n66), .Z(n10409) );
  XNOR U10662 ( .A(n10417), .B(n10631), .Z(n10410) );
  XNOR U10663 ( .A(n10416), .B(n10414), .Z(n10631) );
  AND U10664 ( .A(n10632), .B(n10633), .Z(n10414) );
  NANDN U10665 ( .A(n10634), .B(n10635), .Z(n10633) );
  OR U10666 ( .A(n10636), .B(n10637), .Z(n10635) );
  NAND U10667 ( .A(n10637), .B(n10636), .Z(n10632) );
  ANDN U10668 ( .B(B[22]), .A(n67), .Z(n10416) );
  XNOR U10669 ( .A(n10424), .B(n10638), .Z(n10417) );
  XNOR U10670 ( .A(n10423), .B(n10421), .Z(n10638) );
  AND U10671 ( .A(n10639), .B(n10640), .Z(n10421) );
  NANDN U10672 ( .A(n10641), .B(n10642), .Z(n10640) );
  NANDN U10673 ( .A(n10643), .B(n10644), .Z(n10642) );
  NANDN U10674 ( .A(n10644), .B(n10643), .Z(n10639) );
  ANDN U10675 ( .B(B[23]), .A(n68), .Z(n10423) );
  XNOR U10676 ( .A(n10431), .B(n10645), .Z(n10424) );
  XNOR U10677 ( .A(n10430), .B(n10428), .Z(n10645) );
  AND U10678 ( .A(n10646), .B(n10647), .Z(n10428) );
  NANDN U10679 ( .A(n10648), .B(n10649), .Z(n10647) );
  OR U10680 ( .A(n10650), .B(n10651), .Z(n10649) );
  NAND U10681 ( .A(n10651), .B(n10650), .Z(n10646) );
  ANDN U10682 ( .B(B[24]), .A(n69), .Z(n10430) );
  XNOR U10683 ( .A(n10438), .B(n10652), .Z(n10431) );
  XNOR U10684 ( .A(n10437), .B(n10435), .Z(n10652) );
  AND U10685 ( .A(n10653), .B(n10654), .Z(n10435) );
  NANDN U10686 ( .A(n10655), .B(n10656), .Z(n10654) );
  NANDN U10687 ( .A(n10657), .B(n10658), .Z(n10656) );
  NANDN U10688 ( .A(n10658), .B(n10657), .Z(n10653) );
  ANDN U10689 ( .B(B[25]), .A(n70), .Z(n10437) );
  XNOR U10690 ( .A(n10445), .B(n10659), .Z(n10438) );
  XNOR U10691 ( .A(n10444), .B(n10442), .Z(n10659) );
  AND U10692 ( .A(n10660), .B(n10661), .Z(n10442) );
  NANDN U10693 ( .A(n10662), .B(n10663), .Z(n10661) );
  OR U10694 ( .A(n10664), .B(n10665), .Z(n10663) );
  NAND U10695 ( .A(n10665), .B(n10664), .Z(n10660) );
  ANDN U10696 ( .B(B[26]), .A(n71), .Z(n10444) );
  XNOR U10697 ( .A(n10452), .B(n10666), .Z(n10445) );
  XNOR U10698 ( .A(n10451), .B(n10449), .Z(n10666) );
  AND U10699 ( .A(n10667), .B(n10668), .Z(n10449) );
  NANDN U10700 ( .A(n10669), .B(n10670), .Z(n10668) );
  NANDN U10701 ( .A(n10671), .B(n10672), .Z(n10670) );
  NANDN U10702 ( .A(n10672), .B(n10671), .Z(n10667) );
  ANDN U10703 ( .B(B[27]), .A(n72), .Z(n10451) );
  XNOR U10704 ( .A(n10459), .B(n10673), .Z(n10452) );
  XNOR U10705 ( .A(n10458), .B(n10456), .Z(n10673) );
  AND U10706 ( .A(n10674), .B(n10675), .Z(n10456) );
  NANDN U10707 ( .A(n10676), .B(n10677), .Z(n10675) );
  OR U10708 ( .A(n10678), .B(n10679), .Z(n10677) );
  NAND U10709 ( .A(n10679), .B(n10678), .Z(n10674) );
  ANDN U10710 ( .B(B[28]), .A(n73), .Z(n10458) );
  XNOR U10711 ( .A(n10466), .B(n10680), .Z(n10459) );
  XNOR U10712 ( .A(n10465), .B(n10463), .Z(n10680) );
  AND U10713 ( .A(n10681), .B(n10682), .Z(n10463) );
  NANDN U10714 ( .A(n10683), .B(n10684), .Z(n10682) );
  NANDN U10715 ( .A(n10685), .B(n10686), .Z(n10684) );
  NANDN U10716 ( .A(n10686), .B(n10685), .Z(n10681) );
  ANDN U10717 ( .B(B[29]), .A(n74), .Z(n10465) );
  XNOR U10718 ( .A(n10473), .B(n10687), .Z(n10466) );
  XNOR U10719 ( .A(n10472), .B(n10470), .Z(n10687) );
  AND U10720 ( .A(n10688), .B(n10689), .Z(n10470) );
  NANDN U10721 ( .A(n10690), .B(n10691), .Z(n10689) );
  OR U10722 ( .A(n10692), .B(n10693), .Z(n10691) );
  NAND U10723 ( .A(n10693), .B(n10692), .Z(n10688) );
  ANDN U10724 ( .B(B[30]), .A(n75), .Z(n10472) );
  XNOR U10725 ( .A(n10480), .B(n10694), .Z(n10473) );
  XNOR U10726 ( .A(n10479), .B(n10477), .Z(n10694) );
  AND U10727 ( .A(n10695), .B(n10696), .Z(n10477) );
  NANDN U10728 ( .A(n10697), .B(n10698), .Z(n10696) );
  NANDN U10729 ( .A(n10699), .B(n10700), .Z(n10698) );
  NANDN U10730 ( .A(n10700), .B(n10699), .Z(n10695) );
  ANDN U10731 ( .B(B[31]), .A(n76), .Z(n10479) );
  XNOR U10732 ( .A(n10487), .B(n10701), .Z(n10480) );
  XNOR U10733 ( .A(n10486), .B(n10484), .Z(n10701) );
  AND U10734 ( .A(n10702), .B(n10703), .Z(n10484) );
  NANDN U10735 ( .A(n10704), .B(n10705), .Z(n10703) );
  OR U10736 ( .A(n10706), .B(n10707), .Z(n10705) );
  NAND U10737 ( .A(n10707), .B(n10706), .Z(n10702) );
  ANDN U10738 ( .B(B[32]), .A(n77), .Z(n10486) );
  XNOR U10739 ( .A(n10494), .B(n10708), .Z(n10487) );
  XNOR U10740 ( .A(n10493), .B(n10491), .Z(n10708) );
  AND U10741 ( .A(n10709), .B(n10710), .Z(n10491) );
  NANDN U10742 ( .A(n10711), .B(n10712), .Z(n10710) );
  NANDN U10743 ( .A(n10713), .B(n10714), .Z(n10712) );
  NANDN U10744 ( .A(n10714), .B(n10713), .Z(n10709) );
  ANDN U10745 ( .B(B[33]), .A(n78), .Z(n10493) );
  XNOR U10746 ( .A(n10501), .B(n10715), .Z(n10494) );
  XNOR U10747 ( .A(n10500), .B(n10498), .Z(n10715) );
  AND U10748 ( .A(n10716), .B(n10717), .Z(n10498) );
  NANDN U10749 ( .A(n10718), .B(n10719), .Z(n10717) );
  OR U10750 ( .A(n10720), .B(n10721), .Z(n10719) );
  NAND U10751 ( .A(n10721), .B(n10720), .Z(n10716) );
  ANDN U10752 ( .B(B[34]), .A(n79), .Z(n10500) );
  XNOR U10753 ( .A(n10508), .B(n10722), .Z(n10501) );
  XNOR U10754 ( .A(n10507), .B(n10505), .Z(n10722) );
  AND U10755 ( .A(n10723), .B(n10724), .Z(n10505) );
  NANDN U10756 ( .A(n10725), .B(n10726), .Z(n10724) );
  NANDN U10757 ( .A(n10727), .B(n10728), .Z(n10726) );
  NANDN U10758 ( .A(n10728), .B(n10727), .Z(n10723) );
  ANDN U10759 ( .B(B[35]), .A(n80), .Z(n10507) );
  XNOR U10760 ( .A(n10515), .B(n10729), .Z(n10508) );
  XNOR U10761 ( .A(n10514), .B(n10512), .Z(n10729) );
  AND U10762 ( .A(n10730), .B(n10731), .Z(n10512) );
  NANDN U10763 ( .A(n10732), .B(n10733), .Z(n10731) );
  OR U10764 ( .A(n10734), .B(n10735), .Z(n10733) );
  NAND U10765 ( .A(n10735), .B(n10734), .Z(n10730) );
  ANDN U10766 ( .B(B[36]), .A(n81), .Z(n10514) );
  XNOR U10767 ( .A(n10522), .B(n10736), .Z(n10515) );
  XNOR U10768 ( .A(n10521), .B(n10519), .Z(n10736) );
  AND U10769 ( .A(n10737), .B(n10738), .Z(n10519) );
  NANDN U10770 ( .A(n10739), .B(n10740), .Z(n10738) );
  NAND U10771 ( .A(n10741), .B(n10742), .Z(n10740) );
  ANDN U10772 ( .B(B[37]), .A(n82), .Z(n10521) );
  XOR U10773 ( .A(n10528), .B(n10743), .Z(n10522) );
  XNOR U10774 ( .A(n10526), .B(n10529), .Z(n10743) );
  NAND U10775 ( .A(A[2]), .B(B[38]), .Z(n10529) );
  NANDN U10776 ( .A(n10744), .B(n10745), .Z(n10526) );
  AND U10777 ( .A(A[0]), .B(B[39]), .Z(n10745) );
  XNOR U10778 ( .A(n10531), .B(n10746), .Z(n10528) );
  NAND U10779 ( .A(A[0]), .B(B[40]), .Z(n10746) );
  NAND U10780 ( .A(B[39]), .B(A[1]), .Z(n10531) );
  NAND U10781 ( .A(n10747), .B(n10748), .Z(n207) );
  NANDN U10782 ( .A(n10749), .B(n10750), .Z(n10748) );
  OR U10783 ( .A(n10751), .B(n10752), .Z(n10750) );
  NAND U10784 ( .A(n10752), .B(n10751), .Z(n10747) );
  XOR U10785 ( .A(n209), .B(n208), .Z(\A1[37] ) );
  XOR U10786 ( .A(n10752), .B(n10753), .Z(n208) );
  XNOR U10787 ( .A(n10751), .B(n10749), .Z(n10753) );
  AND U10788 ( .A(n10754), .B(n10755), .Z(n10749) );
  NANDN U10789 ( .A(n10756), .B(n10757), .Z(n10755) );
  NANDN U10790 ( .A(n10758), .B(n10759), .Z(n10757) );
  NANDN U10791 ( .A(n10759), .B(n10758), .Z(n10754) );
  ANDN U10792 ( .B(B[8]), .A(n54), .Z(n10751) );
  XNOR U10793 ( .A(n10546), .B(n10760), .Z(n10752) );
  XNOR U10794 ( .A(n10545), .B(n10543), .Z(n10760) );
  AND U10795 ( .A(n10761), .B(n10762), .Z(n10543) );
  NANDN U10796 ( .A(n10763), .B(n10764), .Z(n10762) );
  OR U10797 ( .A(n10765), .B(n10766), .Z(n10764) );
  NAND U10798 ( .A(n10766), .B(n10765), .Z(n10761) );
  ANDN U10799 ( .B(B[9]), .A(n55), .Z(n10545) );
  XNOR U10800 ( .A(n10553), .B(n10767), .Z(n10546) );
  XNOR U10801 ( .A(n10552), .B(n10550), .Z(n10767) );
  AND U10802 ( .A(n10768), .B(n10769), .Z(n10550) );
  NANDN U10803 ( .A(n10770), .B(n10771), .Z(n10769) );
  NANDN U10804 ( .A(n10772), .B(n10773), .Z(n10771) );
  NANDN U10805 ( .A(n10773), .B(n10772), .Z(n10768) );
  ANDN U10806 ( .B(B[10]), .A(n56), .Z(n10552) );
  XNOR U10807 ( .A(n10560), .B(n10774), .Z(n10553) );
  XNOR U10808 ( .A(n10559), .B(n10557), .Z(n10774) );
  AND U10809 ( .A(n10775), .B(n10776), .Z(n10557) );
  NANDN U10810 ( .A(n10777), .B(n10778), .Z(n10776) );
  OR U10811 ( .A(n10779), .B(n10780), .Z(n10778) );
  NAND U10812 ( .A(n10780), .B(n10779), .Z(n10775) );
  ANDN U10813 ( .B(B[11]), .A(n57), .Z(n10559) );
  XNOR U10814 ( .A(n10567), .B(n10781), .Z(n10560) );
  XNOR U10815 ( .A(n10566), .B(n10564), .Z(n10781) );
  AND U10816 ( .A(n10782), .B(n10783), .Z(n10564) );
  NANDN U10817 ( .A(n10784), .B(n10785), .Z(n10783) );
  NANDN U10818 ( .A(n10786), .B(n10787), .Z(n10785) );
  NANDN U10819 ( .A(n10787), .B(n10786), .Z(n10782) );
  ANDN U10820 ( .B(B[12]), .A(n58), .Z(n10566) );
  XNOR U10821 ( .A(n10574), .B(n10788), .Z(n10567) );
  XNOR U10822 ( .A(n10573), .B(n10571), .Z(n10788) );
  AND U10823 ( .A(n10789), .B(n10790), .Z(n10571) );
  NANDN U10824 ( .A(n10791), .B(n10792), .Z(n10790) );
  OR U10825 ( .A(n10793), .B(n10794), .Z(n10792) );
  NAND U10826 ( .A(n10794), .B(n10793), .Z(n10789) );
  ANDN U10827 ( .B(B[13]), .A(n59), .Z(n10573) );
  XNOR U10828 ( .A(n10581), .B(n10795), .Z(n10574) );
  XNOR U10829 ( .A(n10580), .B(n10578), .Z(n10795) );
  AND U10830 ( .A(n10796), .B(n10797), .Z(n10578) );
  NANDN U10831 ( .A(n10798), .B(n10799), .Z(n10797) );
  NANDN U10832 ( .A(n10800), .B(n10801), .Z(n10799) );
  NANDN U10833 ( .A(n10801), .B(n10800), .Z(n10796) );
  ANDN U10834 ( .B(B[14]), .A(n60), .Z(n10580) );
  XNOR U10835 ( .A(n10588), .B(n10802), .Z(n10581) );
  XNOR U10836 ( .A(n10587), .B(n10585), .Z(n10802) );
  AND U10837 ( .A(n10803), .B(n10804), .Z(n10585) );
  NANDN U10838 ( .A(n10805), .B(n10806), .Z(n10804) );
  OR U10839 ( .A(n10807), .B(n10808), .Z(n10806) );
  NAND U10840 ( .A(n10808), .B(n10807), .Z(n10803) );
  ANDN U10841 ( .B(B[15]), .A(n61), .Z(n10587) );
  XNOR U10842 ( .A(n10595), .B(n10809), .Z(n10588) );
  XNOR U10843 ( .A(n10594), .B(n10592), .Z(n10809) );
  AND U10844 ( .A(n10810), .B(n10811), .Z(n10592) );
  NANDN U10845 ( .A(n10812), .B(n10813), .Z(n10811) );
  NANDN U10846 ( .A(n10814), .B(n10815), .Z(n10813) );
  NANDN U10847 ( .A(n10815), .B(n10814), .Z(n10810) );
  ANDN U10848 ( .B(B[16]), .A(n62), .Z(n10594) );
  XNOR U10849 ( .A(n10602), .B(n10816), .Z(n10595) );
  XNOR U10850 ( .A(n10601), .B(n10599), .Z(n10816) );
  AND U10851 ( .A(n10817), .B(n10818), .Z(n10599) );
  NANDN U10852 ( .A(n10819), .B(n10820), .Z(n10818) );
  OR U10853 ( .A(n10821), .B(n10822), .Z(n10820) );
  NAND U10854 ( .A(n10822), .B(n10821), .Z(n10817) );
  ANDN U10855 ( .B(B[17]), .A(n63), .Z(n10601) );
  XNOR U10856 ( .A(n10609), .B(n10823), .Z(n10602) );
  XNOR U10857 ( .A(n10608), .B(n10606), .Z(n10823) );
  AND U10858 ( .A(n10824), .B(n10825), .Z(n10606) );
  NANDN U10859 ( .A(n10826), .B(n10827), .Z(n10825) );
  NANDN U10860 ( .A(n10828), .B(n10829), .Z(n10827) );
  NANDN U10861 ( .A(n10829), .B(n10828), .Z(n10824) );
  ANDN U10862 ( .B(B[18]), .A(n64), .Z(n10608) );
  XNOR U10863 ( .A(n10616), .B(n10830), .Z(n10609) );
  XNOR U10864 ( .A(n10615), .B(n10613), .Z(n10830) );
  AND U10865 ( .A(n10831), .B(n10832), .Z(n10613) );
  NANDN U10866 ( .A(n10833), .B(n10834), .Z(n10832) );
  OR U10867 ( .A(n10835), .B(n10836), .Z(n10834) );
  NAND U10868 ( .A(n10836), .B(n10835), .Z(n10831) );
  ANDN U10869 ( .B(B[19]), .A(n65), .Z(n10615) );
  XNOR U10870 ( .A(n10623), .B(n10837), .Z(n10616) );
  XNOR U10871 ( .A(n10622), .B(n10620), .Z(n10837) );
  AND U10872 ( .A(n10838), .B(n10839), .Z(n10620) );
  NANDN U10873 ( .A(n10840), .B(n10841), .Z(n10839) );
  NANDN U10874 ( .A(n10842), .B(n10843), .Z(n10841) );
  NANDN U10875 ( .A(n10843), .B(n10842), .Z(n10838) );
  ANDN U10876 ( .B(B[20]), .A(n66), .Z(n10622) );
  XNOR U10877 ( .A(n10630), .B(n10844), .Z(n10623) );
  XNOR U10878 ( .A(n10629), .B(n10627), .Z(n10844) );
  AND U10879 ( .A(n10845), .B(n10846), .Z(n10627) );
  NANDN U10880 ( .A(n10847), .B(n10848), .Z(n10846) );
  OR U10881 ( .A(n10849), .B(n10850), .Z(n10848) );
  NAND U10882 ( .A(n10850), .B(n10849), .Z(n10845) );
  ANDN U10883 ( .B(B[21]), .A(n67), .Z(n10629) );
  XNOR U10884 ( .A(n10637), .B(n10851), .Z(n10630) );
  XNOR U10885 ( .A(n10636), .B(n10634), .Z(n10851) );
  AND U10886 ( .A(n10852), .B(n10853), .Z(n10634) );
  NANDN U10887 ( .A(n10854), .B(n10855), .Z(n10853) );
  NANDN U10888 ( .A(n10856), .B(n10857), .Z(n10855) );
  NANDN U10889 ( .A(n10857), .B(n10856), .Z(n10852) );
  ANDN U10890 ( .B(B[22]), .A(n68), .Z(n10636) );
  XNOR U10891 ( .A(n10644), .B(n10858), .Z(n10637) );
  XNOR U10892 ( .A(n10643), .B(n10641), .Z(n10858) );
  AND U10893 ( .A(n10859), .B(n10860), .Z(n10641) );
  NANDN U10894 ( .A(n10861), .B(n10862), .Z(n10860) );
  OR U10895 ( .A(n10863), .B(n10864), .Z(n10862) );
  NAND U10896 ( .A(n10864), .B(n10863), .Z(n10859) );
  ANDN U10897 ( .B(B[23]), .A(n69), .Z(n10643) );
  XNOR U10898 ( .A(n10651), .B(n10865), .Z(n10644) );
  XNOR U10899 ( .A(n10650), .B(n10648), .Z(n10865) );
  AND U10900 ( .A(n10866), .B(n10867), .Z(n10648) );
  NANDN U10901 ( .A(n10868), .B(n10869), .Z(n10867) );
  NANDN U10902 ( .A(n10870), .B(n10871), .Z(n10869) );
  NANDN U10903 ( .A(n10871), .B(n10870), .Z(n10866) );
  ANDN U10904 ( .B(B[24]), .A(n70), .Z(n10650) );
  XNOR U10905 ( .A(n10658), .B(n10872), .Z(n10651) );
  XNOR U10906 ( .A(n10657), .B(n10655), .Z(n10872) );
  AND U10907 ( .A(n10873), .B(n10874), .Z(n10655) );
  NANDN U10908 ( .A(n10875), .B(n10876), .Z(n10874) );
  OR U10909 ( .A(n10877), .B(n10878), .Z(n10876) );
  NAND U10910 ( .A(n10878), .B(n10877), .Z(n10873) );
  ANDN U10911 ( .B(B[25]), .A(n71), .Z(n10657) );
  XNOR U10912 ( .A(n10665), .B(n10879), .Z(n10658) );
  XNOR U10913 ( .A(n10664), .B(n10662), .Z(n10879) );
  AND U10914 ( .A(n10880), .B(n10881), .Z(n10662) );
  NANDN U10915 ( .A(n10882), .B(n10883), .Z(n10881) );
  NANDN U10916 ( .A(n10884), .B(n10885), .Z(n10883) );
  NANDN U10917 ( .A(n10885), .B(n10884), .Z(n10880) );
  ANDN U10918 ( .B(B[26]), .A(n72), .Z(n10664) );
  XNOR U10919 ( .A(n10672), .B(n10886), .Z(n10665) );
  XNOR U10920 ( .A(n10671), .B(n10669), .Z(n10886) );
  AND U10921 ( .A(n10887), .B(n10888), .Z(n10669) );
  NANDN U10922 ( .A(n10889), .B(n10890), .Z(n10888) );
  OR U10923 ( .A(n10891), .B(n10892), .Z(n10890) );
  NAND U10924 ( .A(n10892), .B(n10891), .Z(n10887) );
  ANDN U10925 ( .B(B[27]), .A(n73), .Z(n10671) );
  XNOR U10926 ( .A(n10679), .B(n10893), .Z(n10672) );
  XNOR U10927 ( .A(n10678), .B(n10676), .Z(n10893) );
  AND U10928 ( .A(n10894), .B(n10895), .Z(n10676) );
  NANDN U10929 ( .A(n10896), .B(n10897), .Z(n10895) );
  NANDN U10930 ( .A(n10898), .B(n10899), .Z(n10897) );
  NANDN U10931 ( .A(n10899), .B(n10898), .Z(n10894) );
  ANDN U10932 ( .B(B[28]), .A(n74), .Z(n10678) );
  XNOR U10933 ( .A(n10686), .B(n10900), .Z(n10679) );
  XNOR U10934 ( .A(n10685), .B(n10683), .Z(n10900) );
  AND U10935 ( .A(n10901), .B(n10902), .Z(n10683) );
  NANDN U10936 ( .A(n10903), .B(n10904), .Z(n10902) );
  OR U10937 ( .A(n10905), .B(n10906), .Z(n10904) );
  NAND U10938 ( .A(n10906), .B(n10905), .Z(n10901) );
  ANDN U10939 ( .B(B[29]), .A(n75), .Z(n10685) );
  XNOR U10940 ( .A(n10693), .B(n10907), .Z(n10686) );
  XNOR U10941 ( .A(n10692), .B(n10690), .Z(n10907) );
  AND U10942 ( .A(n10908), .B(n10909), .Z(n10690) );
  NANDN U10943 ( .A(n10910), .B(n10911), .Z(n10909) );
  NANDN U10944 ( .A(n10912), .B(n10913), .Z(n10911) );
  NANDN U10945 ( .A(n10913), .B(n10912), .Z(n10908) );
  ANDN U10946 ( .B(B[30]), .A(n76), .Z(n10692) );
  XNOR U10947 ( .A(n10700), .B(n10914), .Z(n10693) );
  XNOR U10948 ( .A(n10699), .B(n10697), .Z(n10914) );
  AND U10949 ( .A(n10915), .B(n10916), .Z(n10697) );
  NANDN U10950 ( .A(n10917), .B(n10918), .Z(n10916) );
  OR U10951 ( .A(n10919), .B(n10920), .Z(n10918) );
  NAND U10952 ( .A(n10920), .B(n10919), .Z(n10915) );
  ANDN U10953 ( .B(B[31]), .A(n77), .Z(n10699) );
  XNOR U10954 ( .A(n10707), .B(n10921), .Z(n10700) );
  XNOR U10955 ( .A(n10706), .B(n10704), .Z(n10921) );
  AND U10956 ( .A(n10922), .B(n10923), .Z(n10704) );
  NANDN U10957 ( .A(n10924), .B(n10925), .Z(n10923) );
  NANDN U10958 ( .A(n10926), .B(n10927), .Z(n10925) );
  NANDN U10959 ( .A(n10927), .B(n10926), .Z(n10922) );
  ANDN U10960 ( .B(B[32]), .A(n78), .Z(n10706) );
  XNOR U10961 ( .A(n10714), .B(n10928), .Z(n10707) );
  XNOR U10962 ( .A(n10713), .B(n10711), .Z(n10928) );
  AND U10963 ( .A(n10929), .B(n10930), .Z(n10711) );
  NANDN U10964 ( .A(n10931), .B(n10932), .Z(n10930) );
  OR U10965 ( .A(n10933), .B(n10934), .Z(n10932) );
  NAND U10966 ( .A(n10934), .B(n10933), .Z(n10929) );
  ANDN U10967 ( .B(B[33]), .A(n79), .Z(n10713) );
  XNOR U10968 ( .A(n10721), .B(n10935), .Z(n10714) );
  XNOR U10969 ( .A(n10720), .B(n10718), .Z(n10935) );
  AND U10970 ( .A(n10936), .B(n10937), .Z(n10718) );
  NANDN U10971 ( .A(n10938), .B(n10939), .Z(n10937) );
  NANDN U10972 ( .A(n10940), .B(n10941), .Z(n10939) );
  NANDN U10973 ( .A(n10941), .B(n10940), .Z(n10936) );
  ANDN U10974 ( .B(B[34]), .A(n80), .Z(n10720) );
  XNOR U10975 ( .A(n10728), .B(n10942), .Z(n10721) );
  XNOR U10976 ( .A(n10727), .B(n10725), .Z(n10942) );
  AND U10977 ( .A(n10943), .B(n10944), .Z(n10725) );
  NANDN U10978 ( .A(n10945), .B(n10946), .Z(n10944) );
  OR U10979 ( .A(n10947), .B(n10948), .Z(n10946) );
  NAND U10980 ( .A(n10948), .B(n10947), .Z(n10943) );
  ANDN U10981 ( .B(B[35]), .A(n81), .Z(n10727) );
  XNOR U10982 ( .A(n10735), .B(n10949), .Z(n10728) );
  XNOR U10983 ( .A(n10734), .B(n10732), .Z(n10949) );
  AND U10984 ( .A(n10950), .B(n10951), .Z(n10732) );
  NANDN U10985 ( .A(n10952), .B(n10953), .Z(n10951) );
  NAND U10986 ( .A(n10954), .B(n10955), .Z(n10953) );
  ANDN U10987 ( .B(B[36]), .A(n82), .Z(n10734) );
  XOR U10988 ( .A(n10741), .B(n10956), .Z(n10735) );
  XNOR U10989 ( .A(n10739), .B(n10742), .Z(n10956) );
  NAND U10990 ( .A(A[2]), .B(B[37]), .Z(n10742) );
  NANDN U10991 ( .A(n10957), .B(n10958), .Z(n10739) );
  AND U10992 ( .A(A[0]), .B(B[38]), .Z(n10958) );
  XNOR U10993 ( .A(n10744), .B(n10959), .Z(n10741) );
  NAND U10994 ( .A(A[0]), .B(B[39]), .Z(n10959) );
  NAND U10995 ( .A(B[38]), .B(A[1]), .Z(n10744) );
  NAND U10996 ( .A(n10960), .B(n10961), .Z(n209) );
  NANDN U10997 ( .A(n10962), .B(n10963), .Z(n10961) );
  OR U10998 ( .A(n10964), .B(n10965), .Z(n10963) );
  NAND U10999 ( .A(n10965), .B(n10964), .Z(n10960) );
  XOR U11000 ( .A(n211), .B(n210), .Z(\A1[36] ) );
  XOR U11001 ( .A(n10965), .B(n10966), .Z(n210) );
  XNOR U11002 ( .A(n10964), .B(n10962), .Z(n10966) );
  AND U11003 ( .A(n10967), .B(n10968), .Z(n10962) );
  NANDN U11004 ( .A(n10969), .B(n10970), .Z(n10968) );
  NANDN U11005 ( .A(n10971), .B(n10972), .Z(n10970) );
  NANDN U11006 ( .A(n10972), .B(n10971), .Z(n10967) );
  ANDN U11007 ( .B(B[7]), .A(n54), .Z(n10964) );
  XNOR U11008 ( .A(n10759), .B(n10973), .Z(n10965) );
  XNOR U11009 ( .A(n10758), .B(n10756), .Z(n10973) );
  AND U11010 ( .A(n10974), .B(n10975), .Z(n10756) );
  NANDN U11011 ( .A(n10976), .B(n10977), .Z(n10975) );
  OR U11012 ( .A(n10978), .B(n10979), .Z(n10977) );
  NAND U11013 ( .A(n10979), .B(n10978), .Z(n10974) );
  ANDN U11014 ( .B(B[8]), .A(n55), .Z(n10758) );
  XNOR U11015 ( .A(n10766), .B(n10980), .Z(n10759) );
  XNOR U11016 ( .A(n10765), .B(n10763), .Z(n10980) );
  AND U11017 ( .A(n10981), .B(n10982), .Z(n10763) );
  NANDN U11018 ( .A(n10983), .B(n10984), .Z(n10982) );
  NANDN U11019 ( .A(n10985), .B(n10986), .Z(n10984) );
  NANDN U11020 ( .A(n10986), .B(n10985), .Z(n10981) );
  ANDN U11021 ( .B(B[9]), .A(n56), .Z(n10765) );
  XNOR U11022 ( .A(n10773), .B(n10987), .Z(n10766) );
  XNOR U11023 ( .A(n10772), .B(n10770), .Z(n10987) );
  AND U11024 ( .A(n10988), .B(n10989), .Z(n10770) );
  NANDN U11025 ( .A(n10990), .B(n10991), .Z(n10989) );
  OR U11026 ( .A(n10992), .B(n10993), .Z(n10991) );
  NAND U11027 ( .A(n10993), .B(n10992), .Z(n10988) );
  ANDN U11028 ( .B(B[10]), .A(n57), .Z(n10772) );
  XNOR U11029 ( .A(n10780), .B(n10994), .Z(n10773) );
  XNOR U11030 ( .A(n10779), .B(n10777), .Z(n10994) );
  AND U11031 ( .A(n10995), .B(n10996), .Z(n10777) );
  NANDN U11032 ( .A(n10997), .B(n10998), .Z(n10996) );
  NANDN U11033 ( .A(n10999), .B(n11000), .Z(n10998) );
  NANDN U11034 ( .A(n11000), .B(n10999), .Z(n10995) );
  ANDN U11035 ( .B(B[11]), .A(n58), .Z(n10779) );
  XNOR U11036 ( .A(n10787), .B(n11001), .Z(n10780) );
  XNOR U11037 ( .A(n10786), .B(n10784), .Z(n11001) );
  AND U11038 ( .A(n11002), .B(n11003), .Z(n10784) );
  NANDN U11039 ( .A(n11004), .B(n11005), .Z(n11003) );
  OR U11040 ( .A(n11006), .B(n11007), .Z(n11005) );
  NAND U11041 ( .A(n11007), .B(n11006), .Z(n11002) );
  ANDN U11042 ( .B(B[12]), .A(n59), .Z(n10786) );
  XNOR U11043 ( .A(n10794), .B(n11008), .Z(n10787) );
  XNOR U11044 ( .A(n10793), .B(n10791), .Z(n11008) );
  AND U11045 ( .A(n11009), .B(n11010), .Z(n10791) );
  NANDN U11046 ( .A(n11011), .B(n11012), .Z(n11010) );
  NANDN U11047 ( .A(n11013), .B(n11014), .Z(n11012) );
  NANDN U11048 ( .A(n11014), .B(n11013), .Z(n11009) );
  ANDN U11049 ( .B(B[13]), .A(n60), .Z(n10793) );
  XNOR U11050 ( .A(n10801), .B(n11015), .Z(n10794) );
  XNOR U11051 ( .A(n10800), .B(n10798), .Z(n11015) );
  AND U11052 ( .A(n11016), .B(n11017), .Z(n10798) );
  NANDN U11053 ( .A(n11018), .B(n11019), .Z(n11017) );
  OR U11054 ( .A(n11020), .B(n11021), .Z(n11019) );
  NAND U11055 ( .A(n11021), .B(n11020), .Z(n11016) );
  ANDN U11056 ( .B(B[14]), .A(n61), .Z(n10800) );
  XNOR U11057 ( .A(n10808), .B(n11022), .Z(n10801) );
  XNOR U11058 ( .A(n10807), .B(n10805), .Z(n11022) );
  AND U11059 ( .A(n11023), .B(n11024), .Z(n10805) );
  NANDN U11060 ( .A(n11025), .B(n11026), .Z(n11024) );
  NANDN U11061 ( .A(n11027), .B(n11028), .Z(n11026) );
  NANDN U11062 ( .A(n11028), .B(n11027), .Z(n11023) );
  ANDN U11063 ( .B(B[15]), .A(n62), .Z(n10807) );
  XNOR U11064 ( .A(n10815), .B(n11029), .Z(n10808) );
  XNOR U11065 ( .A(n10814), .B(n10812), .Z(n11029) );
  AND U11066 ( .A(n11030), .B(n11031), .Z(n10812) );
  NANDN U11067 ( .A(n11032), .B(n11033), .Z(n11031) );
  OR U11068 ( .A(n11034), .B(n11035), .Z(n11033) );
  NAND U11069 ( .A(n11035), .B(n11034), .Z(n11030) );
  ANDN U11070 ( .B(B[16]), .A(n63), .Z(n10814) );
  XNOR U11071 ( .A(n10822), .B(n11036), .Z(n10815) );
  XNOR U11072 ( .A(n10821), .B(n10819), .Z(n11036) );
  AND U11073 ( .A(n11037), .B(n11038), .Z(n10819) );
  NANDN U11074 ( .A(n11039), .B(n11040), .Z(n11038) );
  NANDN U11075 ( .A(n11041), .B(n11042), .Z(n11040) );
  NANDN U11076 ( .A(n11042), .B(n11041), .Z(n11037) );
  ANDN U11077 ( .B(B[17]), .A(n64), .Z(n10821) );
  XNOR U11078 ( .A(n10829), .B(n11043), .Z(n10822) );
  XNOR U11079 ( .A(n10828), .B(n10826), .Z(n11043) );
  AND U11080 ( .A(n11044), .B(n11045), .Z(n10826) );
  NANDN U11081 ( .A(n11046), .B(n11047), .Z(n11045) );
  OR U11082 ( .A(n11048), .B(n11049), .Z(n11047) );
  NAND U11083 ( .A(n11049), .B(n11048), .Z(n11044) );
  ANDN U11084 ( .B(B[18]), .A(n65), .Z(n10828) );
  XNOR U11085 ( .A(n10836), .B(n11050), .Z(n10829) );
  XNOR U11086 ( .A(n10835), .B(n10833), .Z(n11050) );
  AND U11087 ( .A(n11051), .B(n11052), .Z(n10833) );
  NANDN U11088 ( .A(n11053), .B(n11054), .Z(n11052) );
  NANDN U11089 ( .A(n11055), .B(n11056), .Z(n11054) );
  NANDN U11090 ( .A(n11056), .B(n11055), .Z(n11051) );
  ANDN U11091 ( .B(B[19]), .A(n66), .Z(n10835) );
  XNOR U11092 ( .A(n10843), .B(n11057), .Z(n10836) );
  XNOR U11093 ( .A(n10842), .B(n10840), .Z(n11057) );
  AND U11094 ( .A(n11058), .B(n11059), .Z(n10840) );
  NANDN U11095 ( .A(n11060), .B(n11061), .Z(n11059) );
  OR U11096 ( .A(n11062), .B(n11063), .Z(n11061) );
  NAND U11097 ( .A(n11063), .B(n11062), .Z(n11058) );
  ANDN U11098 ( .B(B[20]), .A(n67), .Z(n10842) );
  XNOR U11099 ( .A(n10850), .B(n11064), .Z(n10843) );
  XNOR U11100 ( .A(n10849), .B(n10847), .Z(n11064) );
  AND U11101 ( .A(n11065), .B(n11066), .Z(n10847) );
  NANDN U11102 ( .A(n11067), .B(n11068), .Z(n11066) );
  NANDN U11103 ( .A(n11069), .B(n11070), .Z(n11068) );
  NANDN U11104 ( .A(n11070), .B(n11069), .Z(n11065) );
  ANDN U11105 ( .B(B[21]), .A(n68), .Z(n10849) );
  XNOR U11106 ( .A(n10857), .B(n11071), .Z(n10850) );
  XNOR U11107 ( .A(n10856), .B(n10854), .Z(n11071) );
  AND U11108 ( .A(n11072), .B(n11073), .Z(n10854) );
  NANDN U11109 ( .A(n11074), .B(n11075), .Z(n11073) );
  OR U11110 ( .A(n11076), .B(n11077), .Z(n11075) );
  NAND U11111 ( .A(n11077), .B(n11076), .Z(n11072) );
  ANDN U11112 ( .B(B[22]), .A(n69), .Z(n10856) );
  XNOR U11113 ( .A(n10864), .B(n11078), .Z(n10857) );
  XNOR U11114 ( .A(n10863), .B(n10861), .Z(n11078) );
  AND U11115 ( .A(n11079), .B(n11080), .Z(n10861) );
  NANDN U11116 ( .A(n11081), .B(n11082), .Z(n11080) );
  NANDN U11117 ( .A(n11083), .B(n11084), .Z(n11082) );
  NANDN U11118 ( .A(n11084), .B(n11083), .Z(n11079) );
  ANDN U11119 ( .B(B[23]), .A(n70), .Z(n10863) );
  XNOR U11120 ( .A(n10871), .B(n11085), .Z(n10864) );
  XNOR U11121 ( .A(n10870), .B(n10868), .Z(n11085) );
  AND U11122 ( .A(n11086), .B(n11087), .Z(n10868) );
  NANDN U11123 ( .A(n11088), .B(n11089), .Z(n11087) );
  OR U11124 ( .A(n11090), .B(n11091), .Z(n11089) );
  NAND U11125 ( .A(n11091), .B(n11090), .Z(n11086) );
  ANDN U11126 ( .B(B[24]), .A(n71), .Z(n10870) );
  XNOR U11127 ( .A(n10878), .B(n11092), .Z(n10871) );
  XNOR U11128 ( .A(n10877), .B(n10875), .Z(n11092) );
  AND U11129 ( .A(n11093), .B(n11094), .Z(n10875) );
  NANDN U11130 ( .A(n11095), .B(n11096), .Z(n11094) );
  NANDN U11131 ( .A(n11097), .B(n11098), .Z(n11096) );
  NANDN U11132 ( .A(n11098), .B(n11097), .Z(n11093) );
  ANDN U11133 ( .B(B[25]), .A(n72), .Z(n10877) );
  XNOR U11134 ( .A(n10885), .B(n11099), .Z(n10878) );
  XNOR U11135 ( .A(n10884), .B(n10882), .Z(n11099) );
  AND U11136 ( .A(n11100), .B(n11101), .Z(n10882) );
  NANDN U11137 ( .A(n11102), .B(n11103), .Z(n11101) );
  OR U11138 ( .A(n11104), .B(n11105), .Z(n11103) );
  NAND U11139 ( .A(n11105), .B(n11104), .Z(n11100) );
  ANDN U11140 ( .B(B[26]), .A(n73), .Z(n10884) );
  XNOR U11141 ( .A(n10892), .B(n11106), .Z(n10885) );
  XNOR U11142 ( .A(n10891), .B(n10889), .Z(n11106) );
  AND U11143 ( .A(n11107), .B(n11108), .Z(n10889) );
  NANDN U11144 ( .A(n11109), .B(n11110), .Z(n11108) );
  NANDN U11145 ( .A(n11111), .B(n11112), .Z(n11110) );
  NANDN U11146 ( .A(n11112), .B(n11111), .Z(n11107) );
  ANDN U11147 ( .B(B[27]), .A(n74), .Z(n10891) );
  XNOR U11148 ( .A(n10899), .B(n11113), .Z(n10892) );
  XNOR U11149 ( .A(n10898), .B(n10896), .Z(n11113) );
  AND U11150 ( .A(n11114), .B(n11115), .Z(n10896) );
  NANDN U11151 ( .A(n11116), .B(n11117), .Z(n11115) );
  OR U11152 ( .A(n11118), .B(n11119), .Z(n11117) );
  NAND U11153 ( .A(n11119), .B(n11118), .Z(n11114) );
  ANDN U11154 ( .B(B[28]), .A(n75), .Z(n10898) );
  XNOR U11155 ( .A(n10906), .B(n11120), .Z(n10899) );
  XNOR U11156 ( .A(n10905), .B(n10903), .Z(n11120) );
  AND U11157 ( .A(n11121), .B(n11122), .Z(n10903) );
  NANDN U11158 ( .A(n11123), .B(n11124), .Z(n11122) );
  NANDN U11159 ( .A(n11125), .B(n11126), .Z(n11124) );
  NANDN U11160 ( .A(n11126), .B(n11125), .Z(n11121) );
  ANDN U11161 ( .B(B[29]), .A(n76), .Z(n10905) );
  XNOR U11162 ( .A(n10913), .B(n11127), .Z(n10906) );
  XNOR U11163 ( .A(n10912), .B(n10910), .Z(n11127) );
  AND U11164 ( .A(n11128), .B(n11129), .Z(n10910) );
  NANDN U11165 ( .A(n11130), .B(n11131), .Z(n11129) );
  OR U11166 ( .A(n11132), .B(n11133), .Z(n11131) );
  NAND U11167 ( .A(n11133), .B(n11132), .Z(n11128) );
  ANDN U11168 ( .B(B[30]), .A(n77), .Z(n10912) );
  XNOR U11169 ( .A(n10920), .B(n11134), .Z(n10913) );
  XNOR U11170 ( .A(n10919), .B(n10917), .Z(n11134) );
  AND U11171 ( .A(n11135), .B(n11136), .Z(n10917) );
  NANDN U11172 ( .A(n11137), .B(n11138), .Z(n11136) );
  NANDN U11173 ( .A(n11139), .B(n11140), .Z(n11138) );
  NANDN U11174 ( .A(n11140), .B(n11139), .Z(n11135) );
  ANDN U11175 ( .B(B[31]), .A(n78), .Z(n10919) );
  XNOR U11176 ( .A(n10927), .B(n11141), .Z(n10920) );
  XNOR U11177 ( .A(n10926), .B(n10924), .Z(n11141) );
  AND U11178 ( .A(n11142), .B(n11143), .Z(n10924) );
  NANDN U11179 ( .A(n11144), .B(n11145), .Z(n11143) );
  OR U11180 ( .A(n11146), .B(n11147), .Z(n11145) );
  NAND U11181 ( .A(n11147), .B(n11146), .Z(n11142) );
  ANDN U11182 ( .B(B[32]), .A(n79), .Z(n10926) );
  XNOR U11183 ( .A(n10934), .B(n11148), .Z(n10927) );
  XNOR U11184 ( .A(n10933), .B(n10931), .Z(n11148) );
  AND U11185 ( .A(n11149), .B(n11150), .Z(n10931) );
  NANDN U11186 ( .A(n11151), .B(n11152), .Z(n11150) );
  NANDN U11187 ( .A(n11153), .B(n11154), .Z(n11152) );
  NANDN U11188 ( .A(n11154), .B(n11153), .Z(n11149) );
  ANDN U11189 ( .B(B[33]), .A(n80), .Z(n10933) );
  XNOR U11190 ( .A(n10941), .B(n11155), .Z(n10934) );
  XNOR U11191 ( .A(n10940), .B(n10938), .Z(n11155) );
  AND U11192 ( .A(n11156), .B(n11157), .Z(n10938) );
  NANDN U11193 ( .A(n11158), .B(n11159), .Z(n11157) );
  OR U11194 ( .A(n11160), .B(n11161), .Z(n11159) );
  NAND U11195 ( .A(n11161), .B(n11160), .Z(n11156) );
  ANDN U11196 ( .B(B[34]), .A(n81), .Z(n10940) );
  XNOR U11197 ( .A(n10948), .B(n11162), .Z(n10941) );
  XNOR U11198 ( .A(n10947), .B(n10945), .Z(n11162) );
  AND U11199 ( .A(n11163), .B(n11164), .Z(n10945) );
  NANDN U11200 ( .A(n11165), .B(n11166), .Z(n11164) );
  NAND U11201 ( .A(n11167), .B(n11168), .Z(n11166) );
  ANDN U11202 ( .B(B[35]), .A(n82), .Z(n10947) );
  XOR U11203 ( .A(n10954), .B(n11169), .Z(n10948) );
  XNOR U11204 ( .A(n10952), .B(n10955), .Z(n11169) );
  NAND U11205 ( .A(A[2]), .B(B[36]), .Z(n10955) );
  NANDN U11206 ( .A(n11170), .B(n11171), .Z(n10952) );
  AND U11207 ( .A(A[0]), .B(B[37]), .Z(n11171) );
  XNOR U11208 ( .A(n10957), .B(n11172), .Z(n10954) );
  NAND U11209 ( .A(A[0]), .B(B[38]), .Z(n11172) );
  NAND U11210 ( .A(B[37]), .B(A[1]), .Z(n10957) );
  NAND U11211 ( .A(n11173), .B(n11174), .Z(n211) );
  NANDN U11212 ( .A(n11175), .B(n11176), .Z(n11174) );
  OR U11213 ( .A(n11177), .B(n11178), .Z(n11176) );
  NAND U11214 ( .A(n11178), .B(n11177), .Z(n11173) );
  XOR U11215 ( .A(n213), .B(n212), .Z(\A1[35] ) );
  XOR U11216 ( .A(n11178), .B(n11179), .Z(n212) );
  XNOR U11217 ( .A(n11177), .B(n11175), .Z(n11179) );
  AND U11218 ( .A(n11180), .B(n11181), .Z(n11175) );
  NANDN U11219 ( .A(n11182), .B(n11183), .Z(n11181) );
  NANDN U11220 ( .A(n11184), .B(n11185), .Z(n11183) );
  NANDN U11221 ( .A(n11185), .B(n11184), .Z(n11180) );
  ANDN U11222 ( .B(B[6]), .A(n54), .Z(n11177) );
  XNOR U11223 ( .A(n10972), .B(n11186), .Z(n11178) );
  XNOR U11224 ( .A(n10971), .B(n10969), .Z(n11186) );
  AND U11225 ( .A(n11187), .B(n11188), .Z(n10969) );
  NANDN U11226 ( .A(n11189), .B(n11190), .Z(n11188) );
  OR U11227 ( .A(n11191), .B(n11192), .Z(n11190) );
  NAND U11228 ( .A(n11192), .B(n11191), .Z(n11187) );
  ANDN U11229 ( .B(B[7]), .A(n55), .Z(n10971) );
  XNOR U11230 ( .A(n10979), .B(n11193), .Z(n10972) );
  XNOR U11231 ( .A(n10978), .B(n10976), .Z(n11193) );
  AND U11232 ( .A(n11194), .B(n11195), .Z(n10976) );
  NANDN U11233 ( .A(n11196), .B(n11197), .Z(n11195) );
  NANDN U11234 ( .A(n11198), .B(n11199), .Z(n11197) );
  NANDN U11235 ( .A(n11199), .B(n11198), .Z(n11194) );
  ANDN U11236 ( .B(B[8]), .A(n56), .Z(n10978) );
  XNOR U11237 ( .A(n10986), .B(n11200), .Z(n10979) );
  XNOR U11238 ( .A(n10985), .B(n10983), .Z(n11200) );
  AND U11239 ( .A(n11201), .B(n11202), .Z(n10983) );
  NANDN U11240 ( .A(n11203), .B(n11204), .Z(n11202) );
  OR U11241 ( .A(n11205), .B(n11206), .Z(n11204) );
  NAND U11242 ( .A(n11206), .B(n11205), .Z(n11201) );
  ANDN U11243 ( .B(B[9]), .A(n57), .Z(n10985) );
  XNOR U11244 ( .A(n10993), .B(n11207), .Z(n10986) );
  XNOR U11245 ( .A(n10992), .B(n10990), .Z(n11207) );
  AND U11246 ( .A(n11208), .B(n11209), .Z(n10990) );
  NANDN U11247 ( .A(n11210), .B(n11211), .Z(n11209) );
  NANDN U11248 ( .A(n11212), .B(n11213), .Z(n11211) );
  NANDN U11249 ( .A(n11213), .B(n11212), .Z(n11208) );
  ANDN U11250 ( .B(B[10]), .A(n58), .Z(n10992) );
  XNOR U11251 ( .A(n11000), .B(n11214), .Z(n10993) );
  XNOR U11252 ( .A(n10999), .B(n10997), .Z(n11214) );
  AND U11253 ( .A(n11215), .B(n11216), .Z(n10997) );
  NANDN U11254 ( .A(n11217), .B(n11218), .Z(n11216) );
  OR U11255 ( .A(n11219), .B(n11220), .Z(n11218) );
  NAND U11256 ( .A(n11220), .B(n11219), .Z(n11215) );
  ANDN U11257 ( .B(B[11]), .A(n59), .Z(n10999) );
  XNOR U11258 ( .A(n11007), .B(n11221), .Z(n11000) );
  XNOR U11259 ( .A(n11006), .B(n11004), .Z(n11221) );
  AND U11260 ( .A(n11222), .B(n11223), .Z(n11004) );
  NANDN U11261 ( .A(n11224), .B(n11225), .Z(n11223) );
  NANDN U11262 ( .A(n11226), .B(n11227), .Z(n11225) );
  NANDN U11263 ( .A(n11227), .B(n11226), .Z(n11222) );
  ANDN U11264 ( .B(B[12]), .A(n60), .Z(n11006) );
  XNOR U11265 ( .A(n11014), .B(n11228), .Z(n11007) );
  XNOR U11266 ( .A(n11013), .B(n11011), .Z(n11228) );
  AND U11267 ( .A(n11229), .B(n11230), .Z(n11011) );
  NANDN U11268 ( .A(n11231), .B(n11232), .Z(n11230) );
  OR U11269 ( .A(n11233), .B(n11234), .Z(n11232) );
  NAND U11270 ( .A(n11234), .B(n11233), .Z(n11229) );
  ANDN U11271 ( .B(B[13]), .A(n61), .Z(n11013) );
  XNOR U11272 ( .A(n11021), .B(n11235), .Z(n11014) );
  XNOR U11273 ( .A(n11020), .B(n11018), .Z(n11235) );
  AND U11274 ( .A(n11236), .B(n11237), .Z(n11018) );
  NANDN U11275 ( .A(n11238), .B(n11239), .Z(n11237) );
  NANDN U11276 ( .A(n11240), .B(n11241), .Z(n11239) );
  NANDN U11277 ( .A(n11241), .B(n11240), .Z(n11236) );
  ANDN U11278 ( .B(B[14]), .A(n62), .Z(n11020) );
  XNOR U11279 ( .A(n11028), .B(n11242), .Z(n11021) );
  XNOR U11280 ( .A(n11027), .B(n11025), .Z(n11242) );
  AND U11281 ( .A(n11243), .B(n11244), .Z(n11025) );
  NANDN U11282 ( .A(n11245), .B(n11246), .Z(n11244) );
  OR U11283 ( .A(n11247), .B(n11248), .Z(n11246) );
  NAND U11284 ( .A(n11248), .B(n11247), .Z(n11243) );
  ANDN U11285 ( .B(B[15]), .A(n63), .Z(n11027) );
  XNOR U11286 ( .A(n11035), .B(n11249), .Z(n11028) );
  XNOR U11287 ( .A(n11034), .B(n11032), .Z(n11249) );
  AND U11288 ( .A(n11250), .B(n11251), .Z(n11032) );
  NANDN U11289 ( .A(n11252), .B(n11253), .Z(n11251) );
  NANDN U11290 ( .A(n11254), .B(n11255), .Z(n11253) );
  NANDN U11291 ( .A(n11255), .B(n11254), .Z(n11250) );
  ANDN U11292 ( .B(B[16]), .A(n64), .Z(n11034) );
  XNOR U11293 ( .A(n11042), .B(n11256), .Z(n11035) );
  XNOR U11294 ( .A(n11041), .B(n11039), .Z(n11256) );
  AND U11295 ( .A(n11257), .B(n11258), .Z(n11039) );
  NANDN U11296 ( .A(n11259), .B(n11260), .Z(n11258) );
  OR U11297 ( .A(n11261), .B(n11262), .Z(n11260) );
  NAND U11298 ( .A(n11262), .B(n11261), .Z(n11257) );
  ANDN U11299 ( .B(B[17]), .A(n65), .Z(n11041) );
  XNOR U11300 ( .A(n11049), .B(n11263), .Z(n11042) );
  XNOR U11301 ( .A(n11048), .B(n11046), .Z(n11263) );
  AND U11302 ( .A(n11264), .B(n11265), .Z(n11046) );
  NANDN U11303 ( .A(n11266), .B(n11267), .Z(n11265) );
  NANDN U11304 ( .A(n11268), .B(n11269), .Z(n11267) );
  NANDN U11305 ( .A(n11269), .B(n11268), .Z(n11264) );
  ANDN U11306 ( .B(B[18]), .A(n66), .Z(n11048) );
  XNOR U11307 ( .A(n11056), .B(n11270), .Z(n11049) );
  XNOR U11308 ( .A(n11055), .B(n11053), .Z(n11270) );
  AND U11309 ( .A(n11271), .B(n11272), .Z(n11053) );
  NANDN U11310 ( .A(n11273), .B(n11274), .Z(n11272) );
  OR U11311 ( .A(n11275), .B(n11276), .Z(n11274) );
  NAND U11312 ( .A(n11276), .B(n11275), .Z(n11271) );
  ANDN U11313 ( .B(B[19]), .A(n67), .Z(n11055) );
  XNOR U11314 ( .A(n11063), .B(n11277), .Z(n11056) );
  XNOR U11315 ( .A(n11062), .B(n11060), .Z(n11277) );
  AND U11316 ( .A(n11278), .B(n11279), .Z(n11060) );
  NANDN U11317 ( .A(n11280), .B(n11281), .Z(n11279) );
  NANDN U11318 ( .A(n11282), .B(n11283), .Z(n11281) );
  NANDN U11319 ( .A(n11283), .B(n11282), .Z(n11278) );
  ANDN U11320 ( .B(B[20]), .A(n68), .Z(n11062) );
  XNOR U11321 ( .A(n11070), .B(n11284), .Z(n11063) );
  XNOR U11322 ( .A(n11069), .B(n11067), .Z(n11284) );
  AND U11323 ( .A(n11285), .B(n11286), .Z(n11067) );
  NANDN U11324 ( .A(n11287), .B(n11288), .Z(n11286) );
  OR U11325 ( .A(n11289), .B(n11290), .Z(n11288) );
  NAND U11326 ( .A(n11290), .B(n11289), .Z(n11285) );
  ANDN U11327 ( .B(B[21]), .A(n69), .Z(n11069) );
  XNOR U11328 ( .A(n11077), .B(n11291), .Z(n11070) );
  XNOR U11329 ( .A(n11076), .B(n11074), .Z(n11291) );
  AND U11330 ( .A(n11292), .B(n11293), .Z(n11074) );
  NANDN U11331 ( .A(n11294), .B(n11295), .Z(n11293) );
  NANDN U11332 ( .A(n11296), .B(n11297), .Z(n11295) );
  NANDN U11333 ( .A(n11297), .B(n11296), .Z(n11292) );
  ANDN U11334 ( .B(B[22]), .A(n70), .Z(n11076) );
  XNOR U11335 ( .A(n11084), .B(n11298), .Z(n11077) );
  XNOR U11336 ( .A(n11083), .B(n11081), .Z(n11298) );
  AND U11337 ( .A(n11299), .B(n11300), .Z(n11081) );
  NANDN U11338 ( .A(n11301), .B(n11302), .Z(n11300) );
  OR U11339 ( .A(n11303), .B(n11304), .Z(n11302) );
  NAND U11340 ( .A(n11304), .B(n11303), .Z(n11299) );
  ANDN U11341 ( .B(B[23]), .A(n71), .Z(n11083) );
  XNOR U11342 ( .A(n11091), .B(n11305), .Z(n11084) );
  XNOR U11343 ( .A(n11090), .B(n11088), .Z(n11305) );
  AND U11344 ( .A(n11306), .B(n11307), .Z(n11088) );
  NANDN U11345 ( .A(n11308), .B(n11309), .Z(n11307) );
  NANDN U11346 ( .A(n11310), .B(n11311), .Z(n11309) );
  NANDN U11347 ( .A(n11311), .B(n11310), .Z(n11306) );
  ANDN U11348 ( .B(B[24]), .A(n72), .Z(n11090) );
  XNOR U11349 ( .A(n11098), .B(n11312), .Z(n11091) );
  XNOR U11350 ( .A(n11097), .B(n11095), .Z(n11312) );
  AND U11351 ( .A(n11313), .B(n11314), .Z(n11095) );
  NANDN U11352 ( .A(n11315), .B(n11316), .Z(n11314) );
  OR U11353 ( .A(n11317), .B(n11318), .Z(n11316) );
  NAND U11354 ( .A(n11318), .B(n11317), .Z(n11313) );
  ANDN U11355 ( .B(B[25]), .A(n73), .Z(n11097) );
  XNOR U11356 ( .A(n11105), .B(n11319), .Z(n11098) );
  XNOR U11357 ( .A(n11104), .B(n11102), .Z(n11319) );
  AND U11358 ( .A(n11320), .B(n11321), .Z(n11102) );
  NANDN U11359 ( .A(n11322), .B(n11323), .Z(n11321) );
  NANDN U11360 ( .A(n11324), .B(n11325), .Z(n11323) );
  NANDN U11361 ( .A(n11325), .B(n11324), .Z(n11320) );
  ANDN U11362 ( .B(B[26]), .A(n74), .Z(n11104) );
  XNOR U11363 ( .A(n11112), .B(n11326), .Z(n11105) );
  XNOR U11364 ( .A(n11111), .B(n11109), .Z(n11326) );
  AND U11365 ( .A(n11327), .B(n11328), .Z(n11109) );
  NANDN U11366 ( .A(n11329), .B(n11330), .Z(n11328) );
  OR U11367 ( .A(n11331), .B(n11332), .Z(n11330) );
  NAND U11368 ( .A(n11332), .B(n11331), .Z(n11327) );
  ANDN U11369 ( .B(B[27]), .A(n75), .Z(n11111) );
  XNOR U11370 ( .A(n11119), .B(n11333), .Z(n11112) );
  XNOR U11371 ( .A(n11118), .B(n11116), .Z(n11333) );
  AND U11372 ( .A(n11334), .B(n11335), .Z(n11116) );
  NANDN U11373 ( .A(n11336), .B(n11337), .Z(n11335) );
  NANDN U11374 ( .A(n11338), .B(n11339), .Z(n11337) );
  NANDN U11375 ( .A(n11339), .B(n11338), .Z(n11334) );
  ANDN U11376 ( .B(B[28]), .A(n76), .Z(n11118) );
  XNOR U11377 ( .A(n11126), .B(n11340), .Z(n11119) );
  XNOR U11378 ( .A(n11125), .B(n11123), .Z(n11340) );
  AND U11379 ( .A(n11341), .B(n11342), .Z(n11123) );
  NANDN U11380 ( .A(n11343), .B(n11344), .Z(n11342) );
  OR U11381 ( .A(n11345), .B(n11346), .Z(n11344) );
  NAND U11382 ( .A(n11346), .B(n11345), .Z(n11341) );
  ANDN U11383 ( .B(B[29]), .A(n77), .Z(n11125) );
  XNOR U11384 ( .A(n11133), .B(n11347), .Z(n11126) );
  XNOR U11385 ( .A(n11132), .B(n11130), .Z(n11347) );
  AND U11386 ( .A(n11348), .B(n11349), .Z(n11130) );
  NANDN U11387 ( .A(n11350), .B(n11351), .Z(n11349) );
  NANDN U11388 ( .A(n11352), .B(n11353), .Z(n11351) );
  NANDN U11389 ( .A(n11353), .B(n11352), .Z(n11348) );
  ANDN U11390 ( .B(B[30]), .A(n78), .Z(n11132) );
  XNOR U11391 ( .A(n11140), .B(n11354), .Z(n11133) );
  XNOR U11392 ( .A(n11139), .B(n11137), .Z(n11354) );
  AND U11393 ( .A(n11355), .B(n11356), .Z(n11137) );
  NANDN U11394 ( .A(n11357), .B(n11358), .Z(n11356) );
  OR U11395 ( .A(n11359), .B(n11360), .Z(n11358) );
  NAND U11396 ( .A(n11360), .B(n11359), .Z(n11355) );
  ANDN U11397 ( .B(B[31]), .A(n79), .Z(n11139) );
  XNOR U11398 ( .A(n11147), .B(n11361), .Z(n11140) );
  XNOR U11399 ( .A(n11146), .B(n11144), .Z(n11361) );
  AND U11400 ( .A(n11362), .B(n11363), .Z(n11144) );
  NANDN U11401 ( .A(n11364), .B(n11365), .Z(n11363) );
  NANDN U11402 ( .A(n11366), .B(n11367), .Z(n11365) );
  NANDN U11403 ( .A(n11367), .B(n11366), .Z(n11362) );
  ANDN U11404 ( .B(B[32]), .A(n80), .Z(n11146) );
  XNOR U11405 ( .A(n11154), .B(n11368), .Z(n11147) );
  XNOR U11406 ( .A(n11153), .B(n11151), .Z(n11368) );
  AND U11407 ( .A(n11369), .B(n11370), .Z(n11151) );
  NANDN U11408 ( .A(n11371), .B(n11372), .Z(n11370) );
  OR U11409 ( .A(n11373), .B(n11374), .Z(n11372) );
  NAND U11410 ( .A(n11374), .B(n11373), .Z(n11369) );
  ANDN U11411 ( .B(B[33]), .A(n81), .Z(n11153) );
  XNOR U11412 ( .A(n11161), .B(n11375), .Z(n11154) );
  XNOR U11413 ( .A(n11160), .B(n11158), .Z(n11375) );
  AND U11414 ( .A(n11376), .B(n11377), .Z(n11158) );
  NANDN U11415 ( .A(n11378), .B(n11379), .Z(n11377) );
  NAND U11416 ( .A(n11380), .B(n11381), .Z(n11379) );
  ANDN U11417 ( .B(B[34]), .A(n82), .Z(n11160) );
  XOR U11418 ( .A(n11167), .B(n11382), .Z(n11161) );
  XNOR U11419 ( .A(n11165), .B(n11168), .Z(n11382) );
  NAND U11420 ( .A(A[2]), .B(B[35]), .Z(n11168) );
  NANDN U11421 ( .A(n11383), .B(n11384), .Z(n11165) );
  AND U11422 ( .A(A[0]), .B(B[36]), .Z(n11384) );
  XNOR U11423 ( .A(n11170), .B(n11385), .Z(n11167) );
  NAND U11424 ( .A(A[0]), .B(B[37]), .Z(n11385) );
  NAND U11425 ( .A(B[36]), .B(A[1]), .Z(n11170) );
  NAND U11426 ( .A(n11386), .B(n11387), .Z(n213) );
  NANDN U11427 ( .A(n11388), .B(n11389), .Z(n11387) );
  OR U11428 ( .A(n11390), .B(n11391), .Z(n11389) );
  NAND U11429 ( .A(n11391), .B(n11390), .Z(n11386) );
  XOR U11430 ( .A(n215), .B(n214), .Z(\A1[34] ) );
  XOR U11431 ( .A(n11391), .B(n11392), .Z(n214) );
  XNOR U11432 ( .A(n11390), .B(n11388), .Z(n11392) );
  AND U11433 ( .A(n11393), .B(n11394), .Z(n11388) );
  NANDN U11434 ( .A(n11395), .B(n11396), .Z(n11394) );
  NANDN U11435 ( .A(n11397), .B(n11398), .Z(n11396) );
  NANDN U11436 ( .A(n11398), .B(n11397), .Z(n11393) );
  ANDN U11437 ( .B(B[5]), .A(n54), .Z(n11390) );
  XNOR U11438 ( .A(n11185), .B(n11399), .Z(n11391) );
  XNOR U11439 ( .A(n11184), .B(n11182), .Z(n11399) );
  AND U11440 ( .A(n11400), .B(n11401), .Z(n11182) );
  NANDN U11441 ( .A(n11402), .B(n11403), .Z(n11401) );
  OR U11442 ( .A(n11404), .B(n11405), .Z(n11403) );
  NAND U11443 ( .A(n11405), .B(n11404), .Z(n11400) );
  ANDN U11444 ( .B(B[6]), .A(n55), .Z(n11184) );
  XNOR U11445 ( .A(n11192), .B(n11406), .Z(n11185) );
  XNOR U11446 ( .A(n11191), .B(n11189), .Z(n11406) );
  AND U11447 ( .A(n11407), .B(n11408), .Z(n11189) );
  NANDN U11448 ( .A(n11409), .B(n11410), .Z(n11408) );
  NANDN U11449 ( .A(n11411), .B(n11412), .Z(n11410) );
  NANDN U11450 ( .A(n11412), .B(n11411), .Z(n11407) );
  ANDN U11451 ( .B(B[7]), .A(n56), .Z(n11191) );
  XNOR U11452 ( .A(n11199), .B(n11413), .Z(n11192) );
  XNOR U11453 ( .A(n11198), .B(n11196), .Z(n11413) );
  AND U11454 ( .A(n11414), .B(n11415), .Z(n11196) );
  NANDN U11455 ( .A(n11416), .B(n11417), .Z(n11415) );
  OR U11456 ( .A(n11418), .B(n11419), .Z(n11417) );
  NAND U11457 ( .A(n11419), .B(n11418), .Z(n11414) );
  ANDN U11458 ( .B(B[8]), .A(n57), .Z(n11198) );
  XNOR U11459 ( .A(n11206), .B(n11420), .Z(n11199) );
  XNOR U11460 ( .A(n11205), .B(n11203), .Z(n11420) );
  AND U11461 ( .A(n11421), .B(n11422), .Z(n11203) );
  NANDN U11462 ( .A(n11423), .B(n11424), .Z(n11422) );
  NANDN U11463 ( .A(n11425), .B(n11426), .Z(n11424) );
  NANDN U11464 ( .A(n11426), .B(n11425), .Z(n11421) );
  ANDN U11465 ( .B(B[9]), .A(n58), .Z(n11205) );
  XNOR U11466 ( .A(n11213), .B(n11427), .Z(n11206) );
  XNOR U11467 ( .A(n11212), .B(n11210), .Z(n11427) );
  AND U11468 ( .A(n11428), .B(n11429), .Z(n11210) );
  NANDN U11469 ( .A(n11430), .B(n11431), .Z(n11429) );
  OR U11470 ( .A(n11432), .B(n11433), .Z(n11431) );
  NAND U11471 ( .A(n11433), .B(n11432), .Z(n11428) );
  ANDN U11472 ( .B(B[10]), .A(n59), .Z(n11212) );
  XNOR U11473 ( .A(n11220), .B(n11434), .Z(n11213) );
  XNOR U11474 ( .A(n11219), .B(n11217), .Z(n11434) );
  AND U11475 ( .A(n11435), .B(n11436), .Z(n11217) );
  NANDN U11476 ( .A(n11437), .B(n11438), .Z(n11436) );
  NANDN U11477 ( .A(n11439), .B(n11440), .Z(n11438) );
  NANDN U11478 ( .A(n11440), .B(n11439), .Z(n11435) );
  ANDN U11479 ( .B(B[11]), .A(n60), .Z(n11219) );
  XNOR U11480 ( .A(n11227), .B(n11441), .Z(n11220) );
  XNOR U11481 ( .A(n11226), .B(n11224), .Z(n11441) );
  AND U11482 ( .A(n11442), .B(n11443), .Z(n11224) );
  NANDN U11483 ( .A(n11444), .B(n11445), .Z(n11443) );
  OR U11484 ( .A(n11446), .B(n11447), .Z(n11445) );
  NAND U11485 ( .A(n11447), .B(n11446), .Z(n11442) );
  ANDN U11486 ( .B(B[12]), .A(n61), .Z(n11226) );
  XNOR U11487 ( .A(n11234), .B(n11448), .Z(n11227) );
  XNOR U11488 ( .A(n11233), .B(n11231), .Z(n11448) );
  AND U11489 ( .A(n11449), .B(n11450), .Z(n11231) );
  NANDN U11490 ( .A(n11451), .B(n11452), .Z(n11450) );
  NANDN U11491 ( .A(n11453), .B(n11454), .Z(n11452) );
  NANDN U11492 ( .A(n11454), .B(n11453), .Z(n11449) );
  ANDN U11493 ( .B(B[13]), .A(n62), .Z(n11233) );
  XNOR U11494 ( .A(n11241), .B(n11455), .Z(n11234) );
  XNOR U11495 ( .A(n11240), .B(n11238), .Z(n11455) );
  AND U11496 ( .A(n11456), .B(n11457), .Z(n11238) );
  NANDN U11497 ( .A(n11458), .B(n11459), .Z(n11457) );
  OR U11498 ( .A(n11460), .B(n11461), .Z(n11459) );
  NAND U11499 ( .A(n11461), .B(n11460), .Z(n11456) );
  ANDN U11500 ( .B(B[14]), .A(n63), .Z(n11240) );
  XNOR U11501 ( .A(n11248), .B(n11462), .Z(n11241) );
  XNOR U11502 ( .A(n11247), .B(n11245), .Z(n11462) );
  AND U11503 ( .A(n11463), .B(n11464), .Z(n11245) );
  NANDN U11504 ( .A(n11465), .B(n11466), .Z(n11464) );
  NANDN U11505 ( .A(n11467), .B(n11468), .Z(n11466) );
  NANDN U11506 ( .A(n11468), .B(n11467), .Z(n11463) );
  ANDN U11507 ( .B(B[15]), .A(n64), .Z(n11247) );
  XNOR U11508 ( .A(n11255), .B(n11469), .Z(n11248) );
  XNOR U11509 ( .A(n11254), .B(n11252), .Z(n11469) );
  AND U11510 ( .A(n11470), .B(n11471), .Z(n11252) );
  NANDN U11511 ( .A(n11472), .B(n11473), .Z(n11471) );
  OR U11512 ( .A(n11474), .B(n11475), .Z(n11473) );
  NAND U11513 ( .A(n11475), .B(n11474), .Z(n11470) );
  ANDN U11514 ( .B(B[16]), .A(n65), .Z(n11254) );
  XNOR U11515 ( .A(n11262), .B(n11476), .Z(n11255) );
  XNOR U11516 ( .A(n11261), .B(n11259), .Z(n11476) );
  AND U11517 ( .A(n11477), .B(n11478), .Z(n11259) );
  NANDN U11518 ( .A(n11479), .B(n11480), .Z(n11478) );
  NANDN U11519 ( .A(n11481), .B(n11482), .Z(n11480) );
  NANDN U11520 ( .A(n11482), .B(n11481), .Z(n11477) );
  ANDN U11521 ( .B(B[17]), .A(n66), .Z(n11261) );
  XNOR U11522 ( .A(n11269), .B(n11483), .Z(n11262) );
  XNOR U11523 ( .A(n11268), .B(n11266), .Z(n11483) );
  AND U11524 ( .A(n11484), .B(n11485), .Z(n11266) );
  NANDN U11525 ( .A(n11486), .B(n11487), .Z(n11485) );
  OR U11526 ( .A(n11488), .B(n11489), .Z(n11487) );
  NAND U11527 ( .A(n11489), .B(n11488), .Z(n11484) );
  ANDN U11528 ( .B(B[18]), .A(n67), .Z(n11268) );
  XNOR U11529 ( .A(n11276), .B(n11490), .Z(n11269) );
  XNOR U11530 ( .A(n11275), .B(n11273), .Z(n11490) );
  AND U11531 ( .A(n11491), .B(n11492), .Z(n11273) );
  NANDN U11532 ( .A(n11493), .B(n11494), .Z(n11492) );
  NANDN U11533 ( .A(n11495), .B(n11496), .Z(n11494) );
  NANDN U11534 ( .A(n11496), .B(n11495), .Z(n11491) );
  ANDN U11535 ( .B(B[19]), .A(n68), .Z(n11275) );
  XNOR U11536 ( .A(n11283), .B(n11497), .Z(n11276) );
  XNOR U11537 ( .A(n11282), .B(n11280), .Z(n11497) );
  AND U11538 ( .A(n11498), .B(n11499), .Z(n11280) );
  NANDN U11539 ( .A(n11500), .B(n11501), .Z(n11499) );
  OR U11540 ( .A(n11502), .B(n11503), .Z(n11501) );
  NAND U11541 ( .A(n11503), .B(n11502), .Z(n11498) );
  ANDN U11542 ( .B(B[20]), .A(n69), .Z(n11282) );
  XNOR U11543 ( .A(n11290), .B(n11504), .Z(n11283) );
  XNOR U11544 ( .A(n11289), .B(n11287), .Z(n11504) );
  AND U11545 ( .A(n11505), .B(n11506), .Z(n11287) );
  NANDN U11546 ( .A(n11507), .B(n11508), .Z(n11506) );
  NANDN U11547 ( .A(n11509), .B(n11510), .Z(n11508) );
  NANDN U11548 ( .A(n11510), .B(n11509), .Z(n11505) );
  ANDN U11549 ( .B(B[21]), .A(n70), .Z(n11289) );
  XNOR U11550 ( .A(n11297), .B(n11511), .Z(n11290) );
  XNOR U11551 ( .A(n11296), .B(n11294), .Z(n11511) );
  AND U11552 ( .A(n11512), .B(n11513), .Z(n11294) );
  NANDN U11553 ( .A(n11514), .B(n11515), .Z(n11513) );
  OR U11554 ( .A(n11516), .B(n11517), .Z(n11515) );
  NAND U11555 ( .A(n11517), .B(n11516), .Z(n11512) );
  ANDN U11556 ( .B(B[22]), .A(n71), .Z(n11296) );
  XNOR U11557 ( .A(n11304), .B(n11518), .Z(n11297) );
  XNOR U11558 ( .A(n11303), .B(n11301), .Z(n11518) );
  AND U11559 ( .A(n11519), .B(n11520), .Z(n11301) );
  NANDN U11560 ( .A(n11521), .B(n11522), .Z(n11520) );
  NANDN U11561 ( .A(n11523), .B(n11524), .Z(n11522) );
  NANDN U11562 ( .A(n11524), .B(n11523), .Z(n11519) );
  ANDN U11563 ( .B(B[23]), .A(n72), .Z(n11303) );
  XNOR U11564 ( .A(n11311), .B(n11525), .Z(n11304) );
  XNOR U11565 ( .A(n11310), .B(n11308), .Z(n11525) );
  AND U11566 ( .A(n11526), .B(n11527), .Z(n11308) );
  NANDN U11567 ( .A(n11528), .B(n11529), .Z(n11527) );
  OR U11568 ( .A(n11530), .B(n11531), .Z(n11529) );
  NAND U11569 ( .A(n11531), .B(n11530), .Z(n11526) );
  ANDN U11570 ( .B(B[24]), .A(n73), .Z(n11310) );
  XNOR U11571 ( .A(n11318), .B(n11532), .Z(n11311) );
  XNOR U11572 ( .A(n11317), .B(n11315), .Z(n11532) );
  AND U11573 ( .A(n11533), .B(n11534), .Z(n11315) );
  NANDN U11574 ( .A(n11535), .B(n11536), .Z(n11534) );
  NANDN U11575 ( .A(n11537), .B(n11538), .Z(n11536) );
  NANDN U11576 ( .A(n11538), .B(n11537), .Z(n11533) );
  ANDN U11577 ( .B(B[25]), .A(n74), .Z(n11317) );
  XNOR U11578 ( .A(n11325), .B(n11539), .Z(n11318) );
  XNOR U11579 ( .A(n11324), .B(n11322), .Z(n11539) );
  AND U11580 ( .A(n11540), .B(n11541), .Z(n11322) );
  NANDN U11581 ( .A(n11542), .B(n11543), .Z(n11541) );
  OR U11582 ( .A(n11544), .B(n11545), .Z(n11543) );
  NAND U11583 ( .A(n11545), .B(n11544), .Z(n11540) );
  ANDN U11584 ( .B(B[26]), .A(n75), .Z(n11324) );
  XNOR U11585 ( .A(n11332), .B(n11546), .Z(n11325) );
  XNOR U11586 ( .A(n11331), .B(n11329), .Z(n11546) );
  AND U11587 ( .A(n11547), .B(n11548), .Z(n11329) );
  NANDN U11588 ( .A(n11549), .B(n11550), .Z(n11548) );
  NANDN U11589 ( .A(n11551), .B(n11552), .Z(n11550) );
  NANDN U11590 ( .A(n11552), .B(n11551), .Z(n11547) );
  ANDN U11591 ( .B(B[27]), .A(n76), .Z(n11331) );
  XNOR U11592 ( .A(n11339), .B(n11553), .Z(n11332) );
  XNOR U11593 ( .A(n11338), .B(n11336), .Z(n11553) );
  AND U11594 ( .A(n11554), .B(n11555), .Z(n11336) );
  NANDN U11595 ( .A(n11556), .B(n11557), .Z(n11555) );
  OR U11596 ( .A(n11558), .B(n11559), .Z(n11557) );
  NAND U11597 ( .A(n11559), .B(n11558), .Z(n11554) );
  ANDN U11598 ( .B(B[28]), .A(n77), .Z(n11338) );
  XNOR U11599 ( .A(n11346), .B(n11560), .Z(n11339) );
  XNOR U11600 ( .A(n11345), .B(n11343), .Z(n11560) );
  AND U11601 ( .A(n11561), .B(n11562), .Z(n11343) );
  NANDN U11602 ( .A(n11563), .B(n11564), .Z(n11562) );
  NANDN U11603 ( .A(n11565), .B(n11566), .Z(n11564) );
  NANDN U11604 ( .A(n11566), .B(n11565), .Z(n11561) );
  ANDN U11605 ( .B(B[29]), .A(n78), .Z(n11345) );
  XNOR U11606 ( .A(n11353), .B(n11567), .Z(n11346) );
  XNOR U11607 ( .A(n11352), .B(n11350), .Z(n11567) );
  AND U11608 ( .A(n11568), .B(n11569), .Z(n11350) );
  NANDN U11609 ( .A(n11570), .B(n11571), .Z(n11569) );
  OR U11610 ( .A(n11572), .B(n11573), .Z(n11571) );
  NAND U11611 ( .A(n11573), .B(n11572), .Z(n11568) );
  ANDN U11612 ( .B(B[30]), .A(n79), .Z(n11352) );
  XNOR U11613 ( .A(n11360), .B(n11574), .Z(n11353) );
  XNOR U11614 ( .A(n11359), .B(n11357), .Z(n11574) );
  AND U11615 ( .A(n11575), .B(n11576), .Z(n11357) );
  NANDN U11616 ( .A(n11577), .B(n11578), .Z(n11576) );
  NANDN U11617 ( .A(n11579), .B(n11580), .Z(n11578) );
  NANDN U11618 ( .A(n11580), .B(n11579), .Z(n11575) );
  ANDN U11619 ( .B(B[31]), .A(n80), .Z(n11359) );
  XNOR U11620 ( .A(n11367), .B(n11581), .Z(n11360) );
  XNOR U11621 ( .A(n11366), .B(n11364), .Z(n11581) );
  AND U11622 ( .A(n11582), .B(n11583), .Z(n11364) );
  NANDN U11623 ( .A(n11584), .B(n11585), .Z(n11583) );
  OR U11624 ( .A(n11586), .B(n11587), .Z(n11585) );
  NAND U11625 ( .A(n11587), .B(n11586), .Z(n11582) );
  ANDN U11626 ( .B(B[32]), .A(n81), .Z(n11366) );
  XNOR U11627 ( .A(n11374), .B(n11588), .Z(n11367) );
  XNOR U11628 ( .A(n11373), .B(n11371), .Z(n11588) );
  AND U11629 ( .A(n11589), .B(n11590), .Z(n11371) );
  NANDN U11630 ( .A(n11591), .B(n11592), .Z(n11590) );
  NAND U11631 ( .A(n11593), .B(n11594), .Z(n11592) );
  ANDN U11632 ( .B(B[33]), .A(n82), .Z(n11373) );
  XOR U11633 ( .A(n11380), .B(n11595), .Z(n11374) );
  XNOR U11634 ( .A(n11378), .B(n11381), .Z(n11595) );
  NAND U11635 ( .A(A[2]), .B(B[34]), .Z(n11381) );
  NANDN U11636 ( .A(n11596), .B(n11597), .Z(n11378) );
  AND U11637 ( .A(A[0]), .B(B[35]), .Z(n11597) );
  XNOR U11638 ( .A(n11383), .B(n11598), .Z(n11380) );
  NAND U11639 ( .A(A[0]), .B(B[36]), .Z(n11598) );
  NAND U11640 ( .A(B[35]), .B(A[1]), .Z(n11383) );
  NAND U11641 ( .A(n11599), .B(n11600), .Z(n215) );
  NANDN U11642 ( .A(n11601), .B(n11602), .Z(n11600) );
  OR U11643 ( .A(n11603), .B(n11604), .Z(n11602) );
  NAND U11644 ( .A(n11604), .B(n11603), .Z(n11599) );
  XOR U11645 ( .A(n217), .B(n216), .Z(\A1[33] ) );
  XOR U11646 ( .A(n11604), .B(n11605), .Z(n216) );
  XNOR U11647 ( .A(n11603), .B(n11601), .Z(n11605) );
  AND U11648 ( .A(n11606), .B(n11607), .Z(n11601) );
  NANDN U11649 ( .A(n11608), .B(n11609), .Z(n11607) );
  NANDN U11650 ( .A(n11610), .B(n11611), .Z(n11609) );
  NANDN U11651 ( .A(n11611), .B(n11610), .Z(n11606) );
  ANDN U11652 ( .B(B[4]), .A(n54), .Z(n11603) );
  XNOR U11653 ( .A(n11398), .B(n11612), .Z(n11604) );
  XNOR U11654 ( .A(n11397), .B(n11395), .Z(n11612) );
  AND U11655 ( .A(n11613), .B(n11614), .Z(n11395) );
  NANDN U11656 ( .A(n11615), .B(n11616), .Z(n11614) );
  OR U11657 ( .A(n11617), .B(n11618), .Z(n11616) );
  NAND U11658 ( .A(n11618), .B(n11617), .Z(n11613) );
  ANDN U11659 ( .B(B[5]), .A(n55), .Z(n11397) );
  XNOR U11660 ( .A(n11405), .B(n11619), .Z(n11398) );
  XNOR U11661 ( .A(n11404), .B(n11402), .Z(n11619) );
  AND U11662 ( .A(n11620), .B(n11621), .Z(n11402) );
  NANDN U11663 ( .A(n11622), .B(n11623), .Z(n11621) );
  NANDN U11664 ( .A(n11624), .B(n11625), .Z(n11623) );
  NANDN U11665 ( .A(n11625), .B(n11624), .Z(n11620) );
  ANDN U11666 ( .B(B[6]), .A(n56), .Z(n11404) );
  XNOR U11667 ( .A(n11412), .B(n11626), .Z(n11405) );
  XNOR U11668 ( .A(n11411), .B(n11409), .Z(n11626) );
  AND U11669 ( .A(n11627), .B(n11628), .Z(n11409) );
  NANDN U11670 ( .A(n11629), .B(n11630), .Z(n11628) );
  OR U11671 ( .A(n11631), .B(n11632), .Z(n11630) );
  NAND U11672 ( .A(n11632), .B(n11631), .Z(n11627) );
  ANDN U11673 ( .B(B[7]), .A(n57), .Z(n11411) );
  XNOR U11674 ( .A(n11419), .B(n11633), .Z(n11412) );
  XNOR U11675 ( .A(n11418), .B(n11416), .Z(n11633) );
  AND U11676 ( .A(n11634), .B(n11635), .Z(n11416) );
  NANDN U11677 ( .A(n11636), .B(n11637), .Z(n11635) );
  NANDN U11678 ( .A(n11638), .B(n11639), .Z(n11637) );
  NANDN U11679 ( .A(n11639), .B(n11638), .Z(n11634) );
  ANDN U11680 ( .B(B[8]), .A(n58), .Z(n11418) );
  XNOR U11681 ( .A(n11426), .B(n11640), .Z(n11419) );
  XNOR U11682 ( .A(n11425), .B(n11423), .Z(n11640) );
  AND U11683 ( .A(n11641), .B(n11642), .Z(n11423) );
  NANDN U11684 ( .A(n11643), .B(n11644), .Z(n11642) );
  OR U11685 ( .A(n11645), .B(n11646), .Z(n11644) );
  NAND U11686 ( .A(n11646), .B(n11645), .Z(n11641) );
  ANDN U11687 ( .B(B[9]), .A(n59), .Z(n11425) );
  XNOR U11688 ( .A(n11433), .B(n11647), .Z(n11426) );
  XNOR U11689 ( .A(n11432), .B(n11430), .Z(n11647) );
  AND U11690 ( .A(n11648), .B(n11649), .Z(n11430) );
  NANDN U11691 ( .A(n11650), .B(n11651), .Z(n11649) );
  NANDN U11692 ( .A(n11652), .B(n11653), .Z(n11651) );
  NANDN U11693 ( .A(n11653), .B(n11652), .Z(n11648) );
  ANDN U11694 ( .B(B[10]), .A(n60), .Z(n11432) );
  XNOR U11695 ( .A(n11440), .B(n11654), .Z(n11433) );
  XNOR U11696 ( .A(n11439), .B(n11437), .Z(n11654) );
  AND U11697 ( .A(n11655), .B(n11656), .Z(n11437) );
  NANDN U11698 ( .A(n11657), .B(n11658), .Z(n11656) );
  OR U11699 ( .A(n11659), .B(n11660), .Z(n11658) );
  NAND U11700 ( .A(n11660), .B(n11659), .Z(n11655) );
  ANDN U11701 ( .B(B[11]), .A(n61), .Z(n11439) );
  XNOR U11702 ( .A(n11447), .B(n11661), .Z(n11440) );
  XNOR U11703 ( .A(n11446), .B(n11444), .Z(n11661) );
  AND U11704 ( .A(n11662), .B(n11663), .Z(n11444) );
  NANDN U11705 ( .A(n11664), .B(n11665), .Z(n11663) );
  NANDN U11706 ( .A(n11666), .B(n11667), .Z(n11665) );
  NANDN U11707 ( .A(n11667), .B(n11666), .Z(n11662) );
  ANDN U11708 ( .B(B[12]), .A(n62), .Z(n11446) );
  XNOR U11709 ( .A(n11454), .B(n11668), .Z(n11447) );
  XNOR U11710 ( .A(n11453), .B(n11451), .Z(n11668) );
  AND U11711 ( .A(n11669), .B(n11670), .Z(n11451) );
  NANDN U11712 ( .A(n11671), .B(n11672), .Z(n11670) );
  OR U11713 ( .A(n11673), .B(n11674), .Z(n11672) );
  NAND U11714 ( .A(n11674), .B(n11673), .Z(n11669) );
  ANDN U11715 ( .B(B[13]), .A(n63), .Z(n11453) );
  XNOR U11716 ( .A(n11461), .B(n11675), .Z(n11454) );
  XNOR U11717 ( .A(n11460), .B(n11458), .Z(n11675) );
  AND U11718 ( .A(n11676), .B(n11677), .Z(n11458) );
  NANDN U11719 ( .A(n11678), .B(n11679), .Z(n11677) );
  NANDN U11720 ( .A(n11680), .B(n11681), .Z(n11679) );
  NANDN U11721 ( .A(n11681), .B(n11680), .Z(n11676) );
  ANDN U11722 ( .B(B[14]), .A(n64), .Z(n11460) );
  XNOR U11723 ( .A(n11468), .B(n11682), .Z(n11461) );
  XNOR U11724 ( .A(n11467), .B(n11465), .Z(n11682) );
  AND U11725 ( .A(n11683), .B(n11684), .Z(n11465) );
  NANDN U11726 ( .A(n11685), .B(n11686), .Z(n11684) );
  OR U11727 ( .A(n11687), .B(n11688), .Z(n11686) );
  NAND U11728 ( .A(n11688), .B(n11687), .Z(n11683) );
  ANDN U11729 ( .B(B[15]), .A(n65), .Z(n11467) );
  XNOR U11730 ( .A(n11475), .B(n11689), .Z(n11468) );
  XNOR U11731 ( .A(n11474), .B(n11472), .Z(n11689) );
  AND U11732 ( .A(n11690), .B(n11691), .Z(n11472) );
  NANDN U11733 ( .A(n11692), .B(n11693), .Z(n11691) );
  NANDN U11734 ( .A(n11694), .B(n11695), .Z(n11693) );
  NANDN U11735 ( .A(n11695), .B(n11694), .Z(n11690) );
  ANDN U11736 ( .B(B[16]), .A(n66), .Z(n11474) );
  XNOR U11737 ( .A(n11482), .B(n11696), .Z(n11475) );
  XNOR U11738 ( .A(n11481), .B(n11479), .Z(n11696) );
  AND U11739 ( .A(n11697), .B(n11698), .Z(n11479) );
  NANDN U11740 ( .A(n11699), .B(n11700), .Z(n11698) );
  OR U11741 ( .A(n11701), .B(n11702), .Z(n11700) );
  NAND U11742 ( .A(n11702), .B(n11701), .Z(n11697) );
  ANDN U11743 ( .B(B[17]), .A(n67), .Z(n11481) );
  XNOR U11744 ( .A(n11489), .B(n11703), .Z(n11482) );
  XNOR U11745 ( .A(n11488), .B(n11486), .Z(n11703) );
  AND U11746 ( .A(n11704), .B(n11705), .Z(n11486) );
  NANDN U11747 ( .A(n11706), .B(n11707), .Z(n11705) );
  NANDN U11748 ( .A(n11708), .B(n11709), .Z(n11707) );
  NANDN U11749 ( .A(n11709), .B(n11708), .Z(n11704) );
  ANDN U11750 ( .B(B[18]), .A(n68), .Z(n11488) );
  XNOR U11751 ( .A(n11496), .B(n11710), .Z(n11489) );
  XNOR U11752 ( .A(n11495), .B(n11493), .Z(n11710) );
  AND U11753 ( .A(n11711), .B(n11712), .Z(n11493) );
  NANDN U11754 ( .A(n11713), .B(n11714), .Z(n11712) );
  OR U11755 ( .A(n11715), .B(n11716), .Z(n11714) );
  NAND U11756 ( .A(n11716), .B(n11715), .Z(n11711) );
  ANDN U11757 ( .B(B[19]), .A(n69), .Z(n11495) );
  XNOR U11758 ( .A(n11503), .B(n11717), .Z(n11496) );
  XNOR U11759 ( .A(n11502), .B(n11500), .Z(n11717) );
  AND U11760 ( .A(n11718), .B(n11719), .Z(n11500) );
  NANDN U11761 ( .A(n11720), .B(n11721), .Z(n11719) );
  NANDN U11762 ( .A(n11722), .B(n11723), .Z(n11721) );
  NANDN U11763 ( .A(n11723), .B(n11722), .Z(n11718) );
  ANDN U11764 ( .B(B[20]), .A(n70), .Z(n11502) );
  XNOR U11765 ( .A(n11510), .B(n11724), .Z(n11503) );
  XNOR U11766 ( .A(n11509), .B(n11507), .Z(n11724) );
  AND U11767 ( .A(n11725), .B(n11726), .Z(n11507) );
  NANDN U11768 ( .A(n11727), .B(n11728), .Z(n11726) );
  OR U11769 ( .A(n11729), .B(n11730), .Z(n11728) );
  NAND U11770 ( .A(n11730), .B(n11729), .Z(n11725) );
  ANDN U11771 ( .B(B[21]), .A(n71), .Z(n11509) );
  XNOR U11772 ( .A(n11517), .B(n11731), .Z(n11510) );
  XNOR U11773 ( .A(n11516), .B(n11514), .Z(n11731) );
  AND U11774 ( .A(n11732), .B(n11733), .Z(n11514) );
  NANDN U11775 ( .A(n11734), .B(n11735), .Z(n11733) );
  NANDN U11776 ( .A(n11736), .B(n11737), .Z(n11735) );
  NANDN U11777 ( .A(n11737), .B(n11736), .Z(n11732) );
  ANDN U11778 ( .B(B[22]), .A(n72), .Z(n11516) );
  XNOR U11779 ( .A(n11524), .B(n11738), .Z(n11517) );
  XNOR U11780 ( .A(n11523), .B(n11521), .Z(n11738) );
  AND U11781 ( .A(n11739), .B(n11740), .Z(n11521) );
  NANDN U11782 ( .A(n11741), .B(n11742), .Z(n11740) );
  OR U11783 ( .A(n11743), .B(n11744), .Z(n11742) );
  NAND U11784 ( .A(n11744), .B(n11743), .Z(n11739) );
  ANDN U11785 ( .B(B[23]), .A(n73), .Z(n11523) );
  XNOR U11786 ( .A(n11531), .B(n11745), .Z(n11524) );
  XNOR U11787 ( .A(n11530), .B(n11528), .Z(n11745) );
  AND U11788 ( .A(n11746), .B(n11747), .Z(n11528) );
  NANDN U11789 ( .A(n11748), .B(n11749), .Z(n11747) );
  NANDN U11790 ( .A(n11750), .B(n11751), .Z(n11749) );
  NANDN U11791 ( .A(n11751), .B(n11750), .Z(n11746) );
  ANDN U11792 ( .B(B[24]), .A(n74), .Z(n11530) );
  XNOR U11793 ( .A(n11538), .B(n11752), .Z(n11531) );
  XNOR U11794 ( .A(n11537), .B(n11535), .Z(n11752) );
  AND U11795 ( .A(n11753), .B(n11754), .Z(n11535) );
  NANDN U11796 ( .A(n11755), .B(n11756), .Z(n11754) );
  OR U11797 ( .A(n11757), .B(n11758), .Z(n11756) );
  NAND U11798 ( .A(n11758), .B(n11757), .Z(n11753) );
  ANDN U11799 ( .B(B[25]), .A(n75), .Z(n11537) );
  XNOR U11800 ( .A(n11545), .B(n11759), .Z(n11538) );
  XNOR U11801 ( .A(n11544), .B(n11542), .Z(n11759) );
  AND U11802 ( .A(n11760), .B(n11761), .Z(n11542) );
  NANDN U11803 ( .A(n11762), .B(n11763), .Z(n11761) );
  NANDN U11804 ( .A(n11764), .B(n11765), .Z(n11763) );
  NANDN U11805 ( .A(n11765), .B(n11764), .Z(n11760) );
  ANDN U11806 ( .B(B[26]), .A(n76), .Z(n11544) );
  XNOR U11807 ( .A(n11552), .B(n11766), .Z(n11545) );
  XNOR U11808 ( .A(n11551), .B(n11549), .Z(n11766) );
  AND U11809 ( .A(n11767), .B(n11768), .Z(n11549) );
  NANDN U11810 ( .A(n11769), .B(n11770), .Z(n11768) );
  OR U11811 ( .A(n11771), .B(n11772), .Z(n11770) );
  NAND U11812 ( .A(n11772), .B(n11771), .Z(n11767) );
  ANDN U11813 ( .B(B[27]), .A(n77), .Z(n11551) );
  XNOR U11814 ( .A(n11559), .B(n11773), .Z(n11552) );
  XNOR U11815 ( .A(n11558), .B(n11556), .Z(n11773) );
  AND U11816 ( .A(n11774), .B(n11775), .Z(n11556) );
  NANDN U11817 ( .A(n11776), .B(n11777), .Z(n11775) );
  NANDN U11818 ( .A(n11778), .B(n11779), .Z(n11777) );
  NANDN U11819 ( .A(n11779), .B(n11778), .Z(n11774) );
  ANDN U11820 ( .B(B[28]), .A(n78), .Z(n11558) );
  XNOR U11821 ( .A(n11566), .B(n11780), .Z(n11559) );
  XNOR U11822 ( .A(n11565), .B(n11563), .Z(n11780) );
  AND U11823 ( .A(n11781), .B(n11782), .Z(n11563) );
  NANDN U11824 ( .A(n11783), .B(n11784), .Z(n11782) );
  OR U11825 ( .A(n11785), .B(n11786), .Z(n11784) );
  NAND U11826 ( .A(n11786), .B(n11785), .Z(n11781) );
  ANDN U11827 ( .B(B[29]), .A(n79), .Z(n11565) );
  XNOR U11828 ( .A(n11573), .B(n11787), .Z(n11566) );
  XNOR U11829 ( .A(n11572), .B(n11570), .Z(n11787) );
  AND U11830 ( .A(n11788), .B(n11789), .Z(n11570) );
  NANDN U11831 ( .A(n11790), .B(n11791), .Z(n11789) );
  NANDN U11832 ( .A(n11792), .B(n11793), .Z(n11791) );
  NANDN U11833 ( .A(n11793), .B(n11792), .Z(n11788) );
  ANDN U11834 ( .B(B[30]), .A(n80), .Z(n11572) );
  XNOR U11835 ( .A(n11580), .B(n11794), .Z(n11573) );
  XNOR U11836 ( .A(n11579), .B(n11577), .Z(n11794) );
  AND U11837 ( .A(n11795), .B(n11796), .Z(n11577) );
  NANDN U11838 ( .A(n11797), .B(n11798), .Z(n11796) );
  OR U11839 ( .A(n11799), .B(n11800), .Z(n11798) );
  NAND U11840 ( .A(n11800), .B(n11799), .Z(n11795) );
  ANDN U11841 ( .B(B[31]), .A(n81), .Z(n11579) );
  XNOR U11842 ( .A(n11587), .B(n11801), .Z(n11580) );
  XNOR U11843 ( .A(n11586), .B(n11584), .Z(n11801) );
  AND U11844 ( .A(n11802), .B(n11803), .Z(n11584) );
  NANDN U11845 ( .A(n11804), .B(n11805), .Z(n11803) );
  NAND U11846 ( .A(n11806), .B(n11807), .Z(n11805) );
  ANDN U11847 ( .B(B[32]), .A(n82), .Z(n11586) );
  XOR U11848 ( .A(n11593), .B(n11808), .Z(n11587) );
  XNOR U11849 ( .A(n11591), .B(n11594), .Z(n11808) );
  NAND U11850 ( .A(A[2]), .B(B[33]), .Z(n11594) );
  NANDN U11851 ( .A(n11809), .B(n11810), .Z(n11591) );
  AND U11852 ( .A(A[0]), .B(B[34]), .Z(n11810) );
  XNOR U11853 ( .A(n11596), .B(n11811), .Z(n11593) );
  NAND U11854 ( .A(A[0]), .B(B[35]), .Z(n11811) );
  NAND U11855 ( .A(B[34]), .B(A[1]), .Z(n11596) );
  NAND U11856 ( .A(n11812), .B(n11813), .Z(n217) );
  NANDN U11857 ( .A(n11814), .B(n11815), .Z(n11813) );
  OR U11858 ( .A(n11816), .B(n11817), .Z(n11815) );
  NAND U11859 ( .A(n11817), .B(n11816), .Z(n11812) );
  XOR U11860 ( .A(n219), .B(n218), .Z(\A1[32] ) );
  XOR U11861 ( .A(n11817), .B(n11818), .Z(n218) );
  XNOR U11862 ( .A(n11816), .B(n11814), .Z(n11818) );
  AND U11863 ( .A(n11819), .B(n11820), .Z(n11814) );
  NANDN U11864 ( .A(n11821), .B(n11822), .Z(n11820) );
  NANDN U11865 ( .A(n11823), .B(n11824), .Z(n11822) );
  NANDN U11866 ( .A(n11824), .B(n11823), .Z(n11819) );
  ANDN U11867 ( .B(B[3]), .A(n54), .Z(n11816) );
  XNOR U11868 ( .A(n11611), .B(n11825), .Z(n11817) );
  XNOR U11869 ( .A(n11610), .B(n11608), .Z(n11825) );
  AND U11870 ( .A(n11826), .B(n11827), .Z(n11608) );
  NANDN U11871 ( .A(n11828), .B(n11829), .Z(n11827) );
  OR U11872 ( .A(n11830), .B(n11831), .Z(n11829) );
  NAND U11873 ( .A(n11831), .B(n11830), .Z(n11826) );
  ANDN U11874 ( .B(B[4]), .A(n55), .Z(n11610) );
  XNOR U11875 ( .A(n11618), .B(n11832), .Z(n11611) );
  XNOR U11876 ( .A(n11617), .B(n11615), .Z(n11832) );
  AND U11877 ( .A(n11833), .B(n11834), .Z(n11615) );
  NANDN U11878 ( .A(n11835), .B(n11836), .Z(n11834) );
  NANDN U11879 ( .A(n11837), .B(n11838), .Z(n11836) );
  NANDN U11880 ( .A(n11838), .B(n11837), .Z(n11833) );
  ANDN U11881 ( .B(B[5]), .A(n56), .Z(n11617) );
  XNOR U11882 ( .A(n11625), .B(n11839), .Z(n11618) );
  XNOR U11883 ( .A(n11624), .B(n11622), .Z(n11839) );
  AND U11884 ( .A(n11840), .B(n11841), .Z(n11622) );
  NANDN U11885 ( .A(n11842), .B(n11843), .Z(n11841) );
  OR U11886 ( .A(n11844), .B(n11845), .Z(n11843) );
  NAND U11887 ( .A(n11845), .B(n11844), .Z(n11840) );
  ANDN U11888 ( .B(B[6]), .A(n57), .Z(n11624) );
  XNOR U11889 ( .A(n11632), .B(n11846), .Z(n11625) );
  XNOR U11890 ( .A(n11631), .B(n11629), .Z(n11846) );
  AND U11891 ( .A(n11847), .B(n11848), .Z(n11629) );
  NANDN U11892 ( .A(n11849), .B(n11850), .Z(n11848) );
  NANDN U11893 ( .A(n11851), .B(n11852), .Z(n11850) );
  NANDN U11894 ( .A(n11852), .B(n11851), .Z(n11847) );
  ANDN U11895 ( .B(B[7]), .A(n58), .Z(n11631) );
  XNOR U11896 ( .A(n11639), .B(n11853), .Z(n11632) );
  XNOR U11897 ( .A(n11638), .B(n11636), .Z(n11853) );
  AND U11898 ( .A(n11854), .B(n11855), .Z(n11636) );
  NANDN U11899 ( .A(n11856), .B(n11857), .Z(n11855) );
  OR U11900 ( .A(n11858), .B(n11859), .Z(n11857) );
  NAND U11901 ( .A(n11859), .B(n11858), .Z(n11854) );
  ANDN U11902 ( .B(B[8]), .A(n59), .Z(n11638) );
  XNOR U11903 ( .A(n11646), .B(n11860), .Z(n11639) );
  XNOR U11904 ( .A(n11645), .B(n11643), .Z(n11860) );
  AND U11905 ( .A(n11861), .B(n11862), .Z(n11643) );
  NANDN U11906 ( .A(n11863), .B(n11864), .Z(n11862) );
  NANDN U11907 ( .A(n11865), .B(n11866), .Z(n11864) );
  NANDN U11908 ( .A(n11866), .B(n11865), .Z(n11861) );
  ANDN U11909 ( .B(B[9]), .A(n60), .Z(n11645) );
  XNOR U11910 ( .A(n11653), .B(n11867), .Z(n11646) );
  XNOR U11911 ( .A(n11652), .B(n11650), .Z(n11867) );
  AND U11912 ( .A(n11868), .B(n11869), .Z(n11650) );
  NANDN U11913 ( .A(n11870), .B(n11871), .Z(n11869) );
  OR U11914 ( .A(n11872), .B(n11873), .Z(n11871) );
  NAND U11915 ( .A(n11873), .B(n11872), .Z(n11868) );
  ANDN U11916 ( .B(B[10]), .A(n61), .Z(n11652) );
  XNOR U11917 ( .A(n11660), .B(n11874), .Z(n11653) );
  XNOR U11918 ( .A(n11659), .B(n11657), .Z(n11874) );
  AND U11919 ( .A(n11875), .B(n11876), .Z(n11657) );
  NANDN U11920 ( .A(n11877), .B(n11878), .Z(n11876) );
  NANDN U11921 ( .A(n11879), .B(n11880), .Z(n11878) );
  NANDN U11922 ( .A(n11880), .B(n11879), .Z(n11875) );
  ANDN U11923 ( .B(B[11]), .A(n62), .Z(n11659) );
  XNOR U11924 ( .A(n11667), .B(n11881), .Z(n11660) );
  XNOR U11925 ( .A(n11666), .B(n11664), .Z(n11881) );
  AND U11926 ( .A(n11882), .B(n11883), .Z(n11664) );
  NANDN U11927 ( .A(n11884), .B(n11885), .Z(n11883) );
  OR U11928 ( .A(n11886), .B(n11887), .Z(n11885) );
  NAND U11929 ( .A(n11887), .B(n11886), .Z(n11882) );
  ANDN U11930 ( .B(B[12]), .A(n63), .Z(n11666) );
  XNOR U11931 ( .A(n11674), .B(n11888), .Z(n11667) );
  XNOR U11932 ( .A(n11673), .B(n11671), .Z(n11888) );
  AND U11933 ( .A(n11889), .B(n11890), .Z(n11671) );
  NANDN U11934 ( .A(n11891), .B(n11892), .Z(n11890) );
  NANDN U11935 ( .A(n11893), .B(n11894), .Z(n11892) );
  NANDN U11936 ( .A(n11894), .B(n11893), .Z(n11889) );
  ANDN U11937 ( .B(B[13]), .A(n64), .Z(n11673) );
  XNOR U11938 ( .A(n11681), .B(n11895), .Z(n11674) );
  XNOR U11939 ( .A(n11680), .B(n11678), .Z(n11895) );
  AND U11940 ( .A(n11896), .B(n11897), .Z(n11678) );
  NANDN U11941 ( .A(n11898), .B(n11899), .Z(n11897) );
  OR U11942 ( .A(n11900), .B(n11901), .Z(n11899) );
  NAND U11943 ( .A(n11901), .B(n11900), .Z(n11896) );
  ANDN U11944 ( .B(B[14]), .A(n65), .Z(n11680) );
  XNOR U11945 ( .A(n11688), .B(n11902), .Z(n11681) );
  XNOR U11946 ( .A(n11687), .B(n11685), .Z(n11902) );
  AND U11947 ( .A(n11903), .B(n11904), .Z(n11685) );
  NANDN U11948 ( .A(n11905), .B(n11906), .Z(n11904) );
  NANDN U11949 ( .A(n11907), .B(n11908), .Z(n11906) );
  NANDN U11950 ( .A(n11908), .B(n11907), .Z(n11903) );
  ANDN U11951 ( .B(B[15]), .A(n66), .Z(n11687) );
  XNOR U11952 ( .A(n11695), .B(n11909), .Z(n11688) );
  XNOR U11953 ( .A(n11694), .B(n11692), .Z(n11909) );
  AND U11954 ( .A(n11910), .B(n11911), .Z(n11692) );
  NANDN U11955 ( .A(n11912), .B(n11913), .Z(n11911) );
  OR U11956 ( .A(n11914), .B(n11915), .Z(n11913) );
  NAND U11957 ( .A(n11915), .B(n11914), .Z(n11910) );
  ANDN U11958 ( .B(B[16]), .A(n67), .Z(n11694) );
  XNOR U11959 ( .A(n11702), .B(n11916), .Z(n11695) );
  XNOR U11960 ( .A(n11701), .B(n11699), .Z(n11916) );
  AND U11961 ( .A(n11917), .B(n11918), .Z(n11699) );
  NANDN U11962 ( .A(n11919), .B(n11920), .Z(n11918) );
  NANDN U11963 ( .A(n11921), .B(n11922), .Z(n11920) );
  NANDN U11964 ( .A(n11922), .B(n11921), .Z(n11917) );
  ANDN U11965 ( .B(B[17]), .A(n68), .Z(n11701) );
  XNOR U11966 ( .A(n11709), .B(n11923), .Z(n11702) );
  XNOR U11967 ( .A(n11708), .B(n11706), .Z(n11923) );
  AND U11968 ( .A(n11924), .B(n11925), .Z(n11706) );
  NANDN U11969 ( .A(n11926), .B(n11927), .Z(n11925) );
  OR U11970 ( .A(n11928), .B(n11929), .Z(n11927) );
  NAND U11971 ( .A(n11929), .B(n11928), .Z(n11924) );
  ANDN U11972 ( .B(B[18]), .A(n69), .Z(n11708) );
  XNOR U11973 ( .A(n11716), .B(n11930), .Z(n11709) );
  XNOR U11974 ( .A(n11715), .B(n11713), .Z(n11930) );
  AND U11975 ( .A(n11931), .B(n11932), .Z(n11713) );
  NANDN U11976 ( .A(n11933), .B(n11934), .Z(n11932) );
  NANDN U11977 ( .A(n11935), .B(n11936), .Z(n11934) );
  NANDN U11978 ( .A(n11936), .B(n11935), .Z(n11931) );
  ANDN U11979 ( .B(B[19]), .A(n70), .Z(n11715) );
  XNOR U11980 ( .A(n11723), .B(n11937), .Z(n11716) );
  XNOR U11981 ( .A(n11722), .B(n11720), .Z(n11937) );
  AND U11982 ( .A(n11938), .B(n11939), .Z(n11720) );
  NANDN U11983 ( .A(n11940), .B(n11941), .Z(n11939) );
  OR U11984 ( .A(n11942), .B(n11943), .Z(n11941) );
  NAND U11985 ( .A(n11943), .B(n11942), .Z(n11938) );
  ANDN U11986 ( .B(B[20]), .A(n71), .Z(n11722) );
  XNOR U11987 ( .A(n11730), .B(n11944), .Z(n11723) );
  XNOR U11988 ( .A(n11729), .B(n11727), .Z(n11944) );
  AND U11989 ( .A(n11945), .B(n11946), .Z(n11727) );
  NANDN U11990 ( .A(n11947), .B(n11948), .Z(n11946) );
  NANDN U11991 ( .A(n11949), .B(n11950), .Z(n11948) );
  NANDN U11992 ( .A(n11950), .B(n11949), .Z(n11945) );
  ANDN U11993 ( .B(B[21]), .A(n72), .Z(n11729) );
  XNOR U11994 ( .A(n11737), .B(n11951), .Z(n11730) );
  XNOR U11995 ( .A(n11736), .B(n11734), .Z(n11951) );
  AND U11996 ( .A(n11952), .B(n11953), .Z(n11734) );
  NANDN U11997 ( .A(n11954), .B(n11955), .Z(n11953) );
  OR U11998 ( .A(n11956), .B(n11957), .Z(n11955) );
  NAND U11999 ( .A(n11957), .B(n11956), .Z(n11952) );
  ANDN U12000 ( .B(B[22]), .A(n73), .Z(n11736) );
  XNOR U12001 ( .A(n11744), .B(n11958), .Z(n11737) );
  XNOR U12002 ( .A(n11743), .B(n11741), .Z(n11958) );
  AND U12003 ( .A(n11959), .B(n11960), .Z(n11741) );
  NANDN U12004 ( .A(n11961), .B(n11962), .Z(n11960) );
  NANDN U12005 ( .A(n11963), .B(n11964), .Z(n11962) );
  NANDN U12006 ( .A(n11964), .B(n11963), .Z(n11959) );
  ANDN U12007 ( .B(B[23]), .A(n74), .Z(n11743) );
  XNOR U12008 ( .A(n11751), .B(n11965), .Z(n11744) );
  XNOR U12009 ( .A(n11750), .B(n11748), .Z(n11965) );
  AND U12010 ( .A(n11966), .B(n11967), .Z(n11748) );
  NANDN U12011 ( .A(n11968), .B(n11969), .Z(n11967) );
  OR U12012 ( .A(n11970), .B(n11971), .Z(n11969) );
  NAND U12013 ( .A(n11971), .B(n11970), .Z(n11966) );
  ANDN U12014 ( .B(B[24]), .A(n75), .Z(n11750) );
  XNOR U12015 ( .A(n11758), .B(n11972), .Z(n11751) );
  XNOR U12016 ( .A(n11757), .B(n11755), .Z(n11972) );
  AND U12017 ( .A(n11973), .B(n11974), .Z(n11755) );
  NANDN U12018 ( .A(n11975), .B(n11976), .Z(n11974) );
  NANDN U12019 ( .A(n11977), .B(n11978), .Z(n11976) );
  NANDN U12020 ( .A(n11978), .B(n11977), .Z(n11973) );
  ANDN U12021 ( .B(B[25]), .A(n76), .Z(n11757) );
  XNOR U12022 ( .A(n11765), .B(n11979), .Z(n11758) );
  XNOR U12023 ( .A(n11764), .B(n11762), .Z(n11979) );
  AND U12024 ( .A(n11980), .B(n11981), .Z(n11762) );
  NANDN U12025 ( .A(n11982), .B(n11983), .Z(n11981) );
  OR U12026 ( .A(n11984), .B(n11985), .Z(n11983) );
  NAND U12027 ( .A(n11985), .B(n11984), .Z(n11980) );
  ANDN U12028 ( .B(B[26]), .A(n77), .Z(n11764) );
  XNOR U12029 ( .A(n11772), .B(n11986), .Z(n11765) );
  XNOR U12030 ( .A(n11771), .B(n11769), .Z(n11986) );
  AND U12031 ( .A(n11987), .B(n11988), .Z(n11769) );
  NANDN U12032 ( .A(n11989), .B(n11990), .Z(n11988) );
  NANDN U12033 ( .A(n11991), .B(n11992), .Z(n11990) );
  NANDN U12034 ( .A(n11992), .B(n11991), .Z(n11987) );
  ANDN U12035 ( .B(B[27]), .A(n78), .Z(n11771) );
  XNOR U12036 ( .A(n11779), .B(n11993), .Z(n11772) );
  XNOR U12037 ( .A(n11778), .B(n11776), .Z(n11993) );
  AND U12038 ( .A(n11994), .B(n11995), .Z(n11776) );
  NANDN U12039 ( .A(n11996), .B(n11997), .Z(n11995) );
  OR U12040 ( .A(n11998), .B(n11999), .Z(n11997) );
  NAND U12041 ( .A(n11999), .B(n11998), .Z(n11994) );
  ANDN U12042 ( .B(B[28]), .A(n79), .Z(n11778) );
  XNOR U12043 ( .A(n11786), .B(n12000), .Z(n11779) );
  XNOR U12044 ( .A(n11785), .B(n11783), .Z(n12000) );
  AND U12045 ( .A(n12001), .B(n12002), .Z(n11783) );
  NANDN U12046 ( .A(n12003), .B(n12004), .Z(n12002) );
  NANDN U12047 ( .A(n12005), .B(n12006), .Z(n12004) );
  NANDN U12048 ( .A(n12006), .B(n12005), .Z(n12001) );
  ANDN U12049 ( .B(B[29]), .A(n80), .Z(n11785) );
  XNOR U12050 ( .A(n11793), .B(n12007), .Z(n11786) );
  XNOR U12051 ( .A(n11792), .B(n11790), .Z(n12007) );
  AND U12052 ( .A(n12008), .B(n12009), .Z(n11790) );
  NANDN U12053 ( .A(n12010), .B(n12011), .Z(n12009) );
  OR U12054 ( .A(n12012), .B(n12013), .Z(n12011) );
  NAND U12055 ( .A(n12013), .B(n12012), .Z(n12008) );
  ANDN U12056 ( .B(B[30]), .A(n81), .Z(n11792) );
  XNOR U12057 ( .A(n11800), .B(n12014), .Z(n11793) );
  XNOR U12058 ( .A(n11799), .B(n11797), .Z(n12014) );
  AND U12059 ( .A(n12015), .B(n12016), .Z(n11797) );
  NANDN U12060 ( .A(n12017), .B(n12018), .Z(n12016) );
  NAND U12061 ( .A(n12019), .B(n12020), .Z(n12018) );
  ANDN U12062 ( .B(B[31]), .A(n82), .Z(n11799) );
  XOR U12063 ( .A(n11806), .B(n12021), .Z(n11800) );
  XNOR U12064 ( .A(n11804), .B(n11807), .Z(n12021) );
  NAND U12065 ( .A(A[2]), .B(B[32]), .Z(n11807) );
  NANDN U12066 ( .A(n12022), .B(n12023), .Z(n11804) );
  AND U12067 ( .A(A[0]), .B(B[33]), .Z(n12023) );
  XNOR U12068 ( .A(n11809), .B(n12024), .Z(n11806) );
  NAND U12069 ( .A(A[0]), .B(B[34]), .Z(n12024) );
  NAND U12070 ( .A(B[33]), .B(A[1]), .Z(n11809) );
  NAND U12071 ( .A(n12025), .B(n12026), .Z(n219) );
  NANDN U12072 ( .A(n12027), .B(n12028), .Z(n12026) );
  OR U12073 ( .A(n12029), .B(n12030), .Z(n12028) );
  NAND U12074 ( .A(n12030), .B(n12029), .Z(n12025) );
  XOR U12075 ( .A(n221), .B(n220), .Z(\A1[31] ) );
  XOR U12076 ( .A(n12030), .B(n12031), .Z(n220) );
  XNOR U12077 ( .A(n12029), .B(n12027), .Z(n12031) );
  AND U12078 ( .A(n12032), .B(n12033), .Z(n12027) );
  NANDN U12079 ( .A(n12034), .B(n12035), .Z(n12033) );
  NANDN U12080 ( .A(n12036), .B(n12037), .Z(n12035) );
  NANDN U12081 ( .A(n12037), .B(n12036), .Z(n12032) );
  ANDN U12082 ( .B(B[2]), .A(n54), .Z(n12029) );
  XNOR U12083 ( .A(n11824), .B(n12038), .Z(n12030) );
  XNOR U12084 ( .A(n11823), .B(n11821), .Z(n12038) );
  AND U12085 ( .A(n12039), .B(n12040), .Z(n11821) );
  NANDN U12086 ( .A(n12041), .B(n12042), .Z(n12040) );
  OR U12087 ( .A(n12043), .B(n12044), .Z(n12042) );
  NAND U12088 ( .A(n12044), .B(n12043), .Z(n12039) );
  ANDN U12089 ( .B(B[3]), .A(n55), .Z(n11823) );
  XNOR U12090 ( .A(n11831), .B(n12045), .Z(n11824) );
  XNOR U12091 ( .A(n11830), .B(n11828), .Z(n12045) );
  AND U12092 ( .A(n12046), .B(n12047), .Z(n11828) );
  NANDN U12093 ( .A(n12048), .B(n12049), .Z(n12047) );
  NANDN U12094 ( .A(n12050), .B(n12051), .Z(n12049) );
  NANDN U12095 ( .A(n12051), .B(n12050), .Z(n12046) );
  ANDN U12096 ( .B(B[4]), .A(n56), .Z(n11830) );
  XNOR U12097 ( .A(n11838), .B(n12052), .Z(n11831) );
  XNOR U12098 ( .A(n11837), .B(n11835), .Z(n12052) );
  AND U12099 ( .A(n12053), .B(n12054), .Z(n11835) );
  NANDN U12100 ( .A(n12055), .B(n12056), .Z(n12054) );
  OR U12101 ( .A(n12057), .B(n12058), .Z(n12056) );
  NAND U12102 ( .A(n12058), .B(n12057), .Z(n12053) );
  ANDN U12103 ( .B(B[5]), .A(n57), .Z(n11837) );
  XNOR U12104 ( .A(n11845), .B(n12059), .Z(n11838) );
  XNOR U12105 ( .A(n11844), .B(n11842), .Z(n12059) );
  AND U12106 ( .A(n12060), .B(n12061), .Z(n11842) );
  NANDN U12107 ( .A(n12062), .B(n12063), .Z(n12061) );
  NANDN U12108 ( .A(n12064), .B(n12065), .Z(n12063) );
  NANDN U12109 ( .A(n12065), .B(n12064), .Z(n12060) );
  ANDN U12110 ( .B(B[6]), .A(n58), .Z(n11844) );
  XNOR U12111 ( .A(n11852), .B(n12066), .Z(n11845) );
  XNOR U12112 ( .A(n11851), .B(n11849), .Z(n12066) );
  AND U12113 ( .A(n12067), .B(n12068), .Z(n11849) );
  NANDN U12114 ( .A(n12069), .B(n12070), .Z(n12068) );
  OR U12115 ( .A(n12071), .B(n12072), .Z(n12070) );
  NAND U12116 ( .A(n12072), .B(n12071), .Z(n12067) );
  ANDN U12117 ( .B(B[7]), .A(n59), .Z(n11851) );
  XNOR U12118 ( .A(n11859), .B(n12073), .Z(n11852) );
  XNOR U12119 ( .A(n11858), .B(n11856), .Z(n12073) );
  AND U12120 ( .A(n12074), .B(n12075), .Z(n11856) );
  NANDN U12121 ( .A(n12076), .B(n12077), .Z(n12075) );
  NANDN U12122 ( .A(n12078), .B(n12079), .Z(n12077) );
  NANDN U12123 ( .A(n12079), .B(n12078), .Z(n12074) );
  ANDN U12124 ( .B(B[8]), .A(n60), .Z(n11858) );
  XNOR U12125 ( .A(n11866), .B(n12080), .Z(n11859) );
  XNOR U12126 ( .A(n11865), .B(n11863), .Z(n12080) );
  AND U12127 ( .A(n12081), .B(n12082), .Z(n11863) );
  NANDN U12128 ( .A(n12083), .B(n12084), .Z(n12082) );
  OR U12129 ( .A(n12085), .B(n12086), .Z(n12084) );
  NAND U12130 ( .A(n12086), .B(n12085), .Z(n12081) );
  ANDN U12131 ( .B(B[9]), .A(n61), .Z(n11865) );
  XNOR U12132 ( .A(n11873), .B(n12087), .Z(n11866) );
  XNOR U12133 ( .A(n11872), .B(n11870), .Z(n12087) );
  AND U12134 ( .A(n12088), .B(n12089), .Z(n11870) );
  NANDN U12135 ( .A(n12090), .B(n12091), .Z(n12089) );
  NANDN U12136 ( .A(n12092), .B(n12093), .Z(n12091) );
  NANDN U12137 ( .A(n12093), .B(n12092), .Z(n12088) );
  ANDN U12138 ( .B(B[10]), .A(n62), .Z(n11872) );
  XNOR U12139 ( .A(n11880), .B(n12094), .Z(n11873) );
  XNOR U12140 ( .A(n11879), .B(n11877), .Z(n12094) );
  AND U12141 ( .A(n12095), .B(n12096), .Z(n11877) );
  NANDN U12142 ( .A(n12097), .B(n12098), .Z(n12096) );
  OR U12143 ( .A(n12099), .B(n12100), .Z(n12098) );
  NAND U12144 ( .A(n12100), .B(n12099), .Z(n12095) );
  ANDN U12145 ( .B(B[11]), .A(n63), .Z(n11879) );
  XNOR U12146 ( .A(n11887), .B(n12101), .Z(n11880) );
  XNOR U12147 ( .A(n11886), .B(n11884), .Z(n12101) );
  AND U12148 ( .A(n12102), .B(n12103), .Z(n11884) );
  NANDN U12149 ( .A(n12104), .B(n12105), .Z(n12103) );
  NANDN U12150 ( .A(n12106), .B(n12107), .Z(n12105) );
  NANDN U12151 ( .A(n12107), .B(n12106), .Z(n12102) );
  ANDN U12152 ( .B(B[12]), .A(n64), .Z(n11886) );
  XNOR U12153 ( .A(n11894), .B(n12108), .Z(n11887) );
  XNOR U12154 ( .A(n11893), .B(n11891), .Z(n12108) );
  AND U12155 ( .A(n12109), .B(n12110), .Z(n11891) );
  NANDN U12156 ( .A(n12111), .B(n12112), .Z(n12110) );
  OR U12157 ( .A(n12113), .B(n12114), .Z(n12112) );
  NAND U12158 ( .A(n12114), .B(n12113), .Z(n12109) );
  ANDN U12159 ( .B(B[13]), .A(n65), .Z(n11893) );
  XNOR U12160 ( .A(n11901), .B(n12115), .Z(n11894) );
  XNOR U12161 ( .A(n11900), .B(n11898), .Z(n12115) );
  AND U12162 ( .A(n12116), .B(n12117), .Z(n11898) );
  NANDN U12163 ( .A(n12118), .B(n12119), .Z(n12117) );
  NANDN U12164 ( .A(n12120), .B(n12121), .Z(n12119) );
  NANDN U12165 ( .A(n12121), .B(n12120), .Z(n12116) );
  ANDN U12166 ( .B(B[14]), .A(n66), .Z(n11900) );
  XNOR U12167 ( .A(n11908), .B(n12122), .Z(n11901) );
  XNOR U12168 ( .A(n11907), .B(n11905), .Z(n12122) );
  AND U12169 ( .A(n12123), .B(n12124), .Z(n11905) );
  NANDN U12170 ( .A(n12125), .B(n12126), .Z(n12124) );
  OR U12171 ( .A(n12127), .B(n12128), .Z(n12126) );
  NAND U12172 ( .A(n12128), .B(n12127), .Z(n12123) );
  ANDN U12173 ( .B(B[15]), .A(n67), .Z(n11907) );
  XNOR U12174 ( .A(n11915), .B(n12129), .Z(n11908) );
  XNOR U12175 ( .A(n11914), .B(n11912), .Z(n12129) );
  AND U12176 ( .A(n12130), .B(n12131), .Z(n11912) );
  NANDN U12177 ( .A(n12132), .B(n12133), .Z(n12131) );
  NANDN U12178 ( .A(n12134), .B(n12135), .Z(n12133) );
  NANDN U12179 ( .A(n12135), .B(n12134), .Z(n12130) );
  ANDN U12180 ( .B(B[16]), .A(n68), .Z(n11914) );
  XNOR U12181 ( .A(n11922), .B(n12136), .Z(n11915) );
  XNOR U12182 ( .A(n11921), .B(n11919), .Z(n12136) );
  AND U12183 ( .A(n12137), .B(n12138), .Z(n11919) );
  NANDN U12184 ( .A(n12139), .B(n12140), .Z(n12138) );
  OR U12185 ( .A(n12141), .B(n12142), .Z(n12140) );
  NAND U12186 ( .A(n12142), .B(n12141), .Z(n12137) );
  ANDN U12187 ( .B(B[17]), .A(n69), .Z(n11921) );
  XNOR U12188 ( .A(n11929), .B(n12143), .Z(n11922) );
  XNOR U12189 ( .A(n11928), .B(n11926), .Z(n12143) );
  AND U12190 ( .A(n12144), .B(n12145), .Z(n11926) );
  NANDN U12191 ( .A(n12146), .B(n12147), .Z(n12145) );
  NANDN U12192 ( .A(n12148), .B(n12149), .Z(n12147) );
  NANDN U12193 ( .A(n12149), .B(n12148), .Z(n12144) );
  ANDN U12194 ( .B(B[18]), .A(n70), .Z(n11928) );
  XNOR U12195 ( .A(n11936), .B(n12150), .Z(n11929) );
  XNOR U12196 ( .A(n11935), .B(n11933), .Z(n12150) );
  AND U12197 ( .A(n12151), .B(n12152), .Z(n11933) );
  NANDN U12198 ( .A(n12153), .B(n12154), .Z(n12152) );
  OR U12199 ( .A(n12155), .B(n12156), .Z(n12154) );
  NAND U12200 ( .A(n12156), .B(n12155), .Z(n12151) );
  ANDN U12201 ( .B(B[19]), .A(n71), .Z(n11935) );
  XNOR U12202 ( .A(n11943), .B(n12157), .Z(n11936) );
  XNOR U12203 ( .A(n11942), .B(n11940), .Z(n12157) );
  AND U12204 ( .A(n12158), .B(n12159), .Z(n11940) );
  NANDN U12205 ( .A(n12160), .B(n12161), .Z(n12159) );
  NANDN U12206 ( .A(n12162), .B(n12163), .Z(n12161) );
  NANDN U12207 ( .A(n12163), .B(n12162), .Z(n12158) );
  ANDN U12208 ( .B(B[20]), .A(n72), .Z(n11942) );
  XNOR U12209 ( .A(n11950), .B(n12164), .Z(n11943) );
  XNOR U12210 ( .A(n11949), .B(n11947), .Z(n12164) );
  AND U12211 ( .A(n12165), .B(n12166), .Z(n11947) );
  NANDN U12212 ( .A(n12167), .B(n12168), .Z(n12166) );
  OR U12213 ( .A(n12169), .B(n12170), .Z(n12168) );
  NAND U12214 ( .A(n12170), .B(n12169), .Z(n12165) );
  ANDN U12215 ( .B(B[21]), .A(n73), .Z(n11949) );
  XNOR U12216 ( .A(n11957), .B(n12171), .Z(n11950) );
  XNOR U12217 ( .A(n11956), .B(n11954), .Z(n12171) );
  AND U12218 ( .A(n12172), .B(n12173), .Z(n11954) );
  NANDN U12219 ( .A(n12174), .B(n12175), .Z(n12173) );
  NANDN U12220 ( .A(n12176), .B(n12177), .Z(n12175) );
  NANDN U12221 ( .A(n12177), .B(n12176), .Z(n12172) );
  ANDN U12222 ( .B(B[22]), .A(n74), .Z(n11956) );
  XNOR U12223 ( .A(n11964), .B(n12178), .Z(n11957) );
  XNOR U12224 ( .A(n11963), .B(n11961), .Z(n12178) );
  AND U12225 ( .A(n12179), .B(n12180), .Z(n11961) );
  NANDN U12226 ( .A(n12181), .B(n12182), .Z(n12180) );
  OR U12227 ( .A(n12183), .B(n12184), .Z(n12182) );
  NAND U12228 ( .A(n12184), .B(n12183), .Z(n12179) );
  ANDN U12229 ( .B(B[23]), .A(n75), .Z(n11963) );
  XNOR U12230 ( .A(n11971), .B(n12185), .Z(n11964) );
  XNOR U12231 ( .A(n11970), .B(n11968), .Z(n12185) );
  AND U12232 ( .A(n12186), .B(n12187), .Z(n11968) );
  NANDN U12233 ( .A(n12188), .B(n12189), .Z(n12187) );
  NANDN U12234 ( .A(n12190), .B(n12191), .Z(n12189) );
  NANDN U12235 ( .A(n12191), .B(n12190), .Z(n12186) );
  ANDN U12236 ( .B(B[24]), .A(n76), .Z(n11970) );
  XNOR U12237 ( .A(n11978), .B(n12192), .Z(n11971) );
  XNOR U12238 ( .A(n11977), .B(n11975), .Z(n12192) );
  AND U12239 ( .A(n12193), .B(n12194), .Z(n11975) );
  NANDN U12240 ( .A(n12195), .B(n12196), .Z(n12194) );
  OR U12241 ( .A(n12197), .B(n12198), .Z(n12196) );
  NAND U12242 ( .A(n12198), .B(n12197), .Z(n12193) );
  ANDN U12243 ( .B(B[25]), .A(n77), .Z(n11977) );
  XNOR U12244 ( .A(n11985), .B(n12199), .Z(n11978) );
  XNOR U12245 ( .A(n11984), .B(n11982), .Z(n12199) );
  AND U12246 ( .A(n12200), .B(n12201), .Z(n11982) );
  NANDN U12247 ( .A(n12202), .B(n12203), .Z(n12201) );
  NANDN U12248 ( .A(n12204), .B(n12205), .Z(n12203) );
  NANDN U12249 ( .A(n12205), .B(n12204), .Z(n12200) );
  ANDN U12250 ( .B(B[26]), .A(n78), .Z(n11984) );
  XNOR U12251 ( .A(n11992), .B(n12206), .Z(n11985) );
  XNOR U12252 ( .A(n11991), .B(n11989), .Z(n12206) );
  AND U12253 ( .A(n12207), .B(n12208), .Z(n11989) );
  NANDN U12254 ( .A(n12209), .B(n12210), .Z(n12208) );
  OR U12255 ( .A(n12211), .B(n12212), .Z(n12210) );
  NAND U12256 ( .A(n12212), .B(n12211), .Z(n12207) );
  ANDN U12257 ( .B(B[27]), .A(n79), .Z(n11991) );
  XNOR U12258 ( .A(n11999), .B(n12213), .Z(n11992) );
  XNOR U12259 ( .A(n11998), .B(n11996), .Z(n12213) );
  AND U12260 ( .A(n12214), .B(n12215), .Z(n11996) );
  NANDN U12261 ( .A(n12216), .B(n12217), .Z(n12215) );
  NANDN U12262 ( .A(n12218), .B(n12219), .Z(n12217) );
  NANDN U12263 ( .A(n12219), .B(n12218), .Z(n12214) );
  ANDN U12264 ( .B(B[28]), .A(n80), .Z(n11998) );
  XNOR U12265 ( .A(n12006), .B(n12220), .Z(n11999) );
  XNOR U12266 ( .A(n12005), .B(n12003), .Z(n12220) );
  AND U12267 ( .A(n12221), .B(n12222), .Z(n12003) );
  NANDN U12268 ( .A(n12223), .B(n12224), .Z(n12222) );
  OR U12269 ( .A(n12225), .B(n12226), .Z(n12224) );
  NAND U12270 ( .A(n12226), .B(n12225), .Z(n12221) );
  ANDN U12271 ( .B(B[29]), .A(n81), .Z(n12005) );
  XNOR U12272 ( .A(n12013), .B(n12227), .Z(n12006) );
  XNOR U12273 ( .A(n12012), .B(n12010), .Z(n12227) );
  AND U12274 ( .A(n12228), .B(n12229), .Z(n12010) );
  NANDN U12275 ( .A(n12230), .B(n12231), .Z(n12229) );
  NAND U12276 ( .A(n12232), .B(n12233), .Z(n12231) );
  ANDN U12277 ( .B(B[30]), .A(n82), .Z(n12012) );
  XOR U12278 ( .A(n12019), .B(n12234), .Z(n12013) );
  XNOR U12279 ( .A(n12017), .B(n12020), .Z(n12234) );
  NAND U12280 ( .A(A[2]), .B(B[31]), .Z(n12020) );
  NANDN U12281 ( .A(n12235), .B(n12236), .Z(n12017) );
  AND U12282 ( .A(A[0]), .B(B[32]), .Z(n12236) );
  XNOR U12283 ( .A(n12022), .B(n12237), .Z(n12019) );
  NAND U12284 ( .A(A[0]), .B(B[33]), .Z(n12237) );
  NAND U12285 ( .A(B[32]), .B(A[1]), .Z(n12022) );
  NAND U12286 ( .A(n12238), .B(n12239), .Z(n221) );
  NANDN U12287 ( .A(n12240), .B(n12241), .Z(n12239) );
  OR U12288 ( .A(n12242), .B(n12243), .Z(n12241) );
  NAND U12289 ( .A(n12243), .B(n12242), .Z(n12238) );
  XOR U12290 ( .A(n223), .B(n222), .Z(\A1[30] ) );
  XOR U12291 ( .A(n12243), .B(n12244), .Z(n222) );
  XNOR U12292 ( .A(n12242), .B(n12240), .Z(n12244) );
  AND U12293 ( .A(n12245), .B(n12246), .Z(n12240) );
  NANDN U12294 ( .A(n12247), .B(n12248), .Z(n12246) );
  NANDN U12295 ( .A(n12249), .B(n12250), .Z(n12248) );
  NANDN U12296 ( .A(n12250), .B(n12249), .Z(n12245) );
  ANDN U12297 ( .B(B[1]), .A(n54), .Z(n12242) );
  XNOR U12298 ( .A(n12037), .B(n12251), .Z(n12243) );
  XNOR U12299 ( .A(n12036), .B(n12034), .Z(n12251) );
  AND U12300 ( .A(n12252), .B(n12253), .Z(n12034) );
  NANDN U12301 ( .A(n12254), .B(n12255), .Z(n12253) );
  OR U12302 ( .A(n12256), .B(n12257), .Z(n12255) );
  NAND U12303 ( .A(n12257), .B(n12256), .Z(n12252) );
  ANDN U12304 ( .B(B[2]), .A(n55), .Z(n12036) );
  XNOR U12305 ( .A(n12044), .B(n12258), .Z(n12037) );
  XNOR U12306 ( .A(n12043), .B(n12041), .Z(n12258) );
  AND U12307 ( .A(n12259), .B(n12260), .Z(n12041) );
  NANDN U12308 ( .A(n12261), .B(n12262), .Z(n12260) );
  NANDN U12309 ( .A(n12263), .B(n12264), .Z(n12262) );
  NANDN U12310 ( .A(n12264), .B(n12263), .Z(n12259) );
  ANDN U12311 ( .B(B[3]), .A(n56), .Z(n12043) );
  XNOR U12312 ( .A(n12051), .B(n12265), .Z(n12044) );
  XNOR U12313 ( .A(n12050), .B(n12048), .Z(n12265) );
  AND U12314 ( .A(n12266), .B(n12267), .Z(n12048) );
  NANDN U12315 ( .A(n12268), .B(n12269), .Z(n12267) );
  OR U12316 ( .A(n12270), .B(n12271), .Z(n12269) );
  NAND U12317 ( .A(n12271), .B(n12270), .Z(n12266) );
  ANDN U12318 ( .B(B[4]), .A(n57), .Z(n12050) );
  XNOR U12319 ( .A(n12058), .B(n12272), .Z(n12051) );
  XNOR U12320 ( .A(n12057), .B(n12055), .Z(n12272) );
  AND U12321 ( .A(n12273), .B(n12274), .Z(n12055) );
  NANDN U12322 ( .A(n12275), .B(n12276), .Z(n12274) );
  NANDN U12323 ( .A(n12277), .B(n12278), .Z(n12276) );
  NANDN U12324 ( .A(n12278), .B(n12277), .Z(n12273) );
  ANDN U12325 ( .B(B[5]), .A(n58), .Z(n12057) );
  XNOR U12326 ( .A(n12065), .B(n12279), .Z(n12058) );
  XNOR U12327 ( .A(n12064), .B(n12062), .Z(n12279) );
  AND U12328 ( .A(n12280), .B(n12281), .Z(n12062) );
  NANDN U12329 ( .A(n12282), .B(n12283), .Z(n12281) );
  OR U12330 ( .A(n12284), .B(n12285), .Z(n12283) );
  NAND U12331 ( .A(n12285), .B(n12284), .Z(n12280) );
  ANDN U12332 ( .B(B[6]), .A(n59), .Z(n12064) );
  XNOR U12333 ( .A(n12072), .B(n12286), .Z(n12065) );
  XNOR U12334 ( .A(n12071), .B(n12069), .Z(n12286) );
  AND U12335 ( .A(n12287), .B(n12288), .Z(n12069) );
  NANDN U12336 ( .A(n12289), .B(n12290), .Z(n12288) );
  NANDN U12337 ( .A(n12291), .B(n12292), .Z(n12290) );
  NANDN U12338 ( .A(n12292), .B(n12291), .Z(n12287) );
  ANDN U12339 ( .B(B[7]), .A(n60), .Z(n12071) );
  XNOR U12340 ( .A(n12079), .B(n12293), .Z(n12072) );
  XNOR U12341 ( .A(n12078), .B(n12076), .Z(n12293) );
  AND U12342 ( .A(n12294), .B(n12295), .Z(n12076) );
  NANDN U12343 ( .A(n12296), .B(n12297), .Z(n12295) );
  OR U12344 ( .A(n12298), .B(n12299), .Z(n12297) );
  NAND U12345 ( .A(n12299), .B(n12298), .Z(n12294) );
  ANDN U12346 ( .B(B[8]), .A(n61), .Z(n12078) );
  XNOR U12347 ( .A(n12086), .B(n12300), .Z(n12079) );
  XNOR U12348 ( .A(n12085), .B(n12083), .Z(n12300) );
  AND U12349 ( .A(n12301), .B(n12302), .Z(n12083) );
  NANDN U12350 ( .A(n12303), .B(n12304), .Z(n12302) );
  NANDN U12351 ( .A(n12305), .B(n12306), .Z(n12304) );
  NANDN U12352 ( .A(n12306), .B(n12305), .Z(n12301) );
  ANDN U12353 ( .B(B[9]), .A(n62), .Z(n12085) );
  XNOR U12354 ( .A(n12093), .B(n12307), .Z(n12086) );
  XNOR U12355 ( .A(n12092), .B(n12090), .Z(n12307) );
  AND U12356 ( .A(n12308), .B(n12309), .Z(n12090) );
  NANDN U12357 ( .A(n12310), .B(n12311), .Z(n12309) );
  OR U12358 ( .A(n12312), .B(n12313), .Z(n12311) );
  NAND U12359 ( .A(n12313), .B(n12312), .Z(n12308) );
  ANDN U12360 ( .B(B[10]), .A(n63), .Z(n12092) );
  XNOR U12361 ( .A(n12100), .B(n12314), .Z(n12093) );
  XNOR U12362 ( .A(n12099), .B(n12097), .Z(n12314) );
  AND U12363 ( .A(n12315), .B(n12316), .Z(n12097) );
  NANDN U12364 ( .A(n12317), .B(n12318), .Z(n12316) );
  NANDN U12365 ( .A(n12319), .B(n12320), .Z(n12318) );
  NANDN U12366 ( .A(n12320), .B(n12319), .Z(n12315) );
  ANDN U12367 ( .B(B[11]), .A(n64), .Z(n12099) );
  XNOR U12368 ( .A(n12107), .B(n12321), .Z(n12100) );
  XNOR U12369 ( .A(n12106), .B(n12104), .Z(n12321) );
  AND U12370 ( .A(n12322), .B(n12323), .Z(n12104) );
  NANDN U12371 ( .A(n12324), .B(n12325), .Z(n12323) );
  OR U12372 ( .A(n12326), .B(n12327), .Z(n12325) );
  NAND U12373 ( .A(n12327), .B(n12326), .Z(n12322) );
  ANDN U12374 ( .B(B[12]), .A(n65), .Z(n12106) );
  XNOR U12375 ( .A(n12114), .B(n12328), .Z(n12107) );
  XNOR U12376 ( .A(n12113), .B(n12111), .Z(n12328) );
  AND U12377 ( .A(n12329), .B(n12330), .Z(n12111) );
  NANDN U12378 ( .A(n12331), .B(n12332), .Z(n12330) );
  NANDN U12379 ( .A(n12333), .B(n12334), .Z(n12332) );
  NANDN U12380 ( .A(n12334), .B(n12333), .Z(n12329) );
  ANDN U12381 ( .B(B[13]), .A(n66), .Z(n12113) );
  XNOR U12382 ( .A(n12121), .B(n12335), .Z(n12114) );
  XNOR U12383 ( .A(n12120), .B(n12118), .Z(n12335) );
  AND U12384 ( .A(n12336), .B(n12337), .Z(n12118) );
  NANDN U12385 ( .A(n12338), .B(n12339), .Z(n12337) );
  OR U12386 ( .A(n12340), .B(n12341), .Z(n12339) );
  NAND U12387 ( .A(n12341), .B(n12340), .Z(n12336) );
  ANDN U12388 ( .B(B[14]), .A(n67), .Z(n12120) );
  XNOR U12389 ( .A(n12128), .B(n12342), .Z(n12121) );
  XNOR U12390 ( .A(n12127), .B(n12125), .Z(n12342) );
  AND U12391 ( .A(n12343), .B(n12344), .Z(n12125) );
  NANDN U12392 ( .A(n12345), .B(n12346), .Z(n12344) );
  NANDN U12393 ( .A(n12347), .B(n12348), .Z(n12346) );
  NANDN U12394 ( .A(n12348), .B(n12347), .Z(n12343) );
  ANDN U12395 ( .B(B[15]), .A(n68), .Z(n12127) );
  XNOR U12396 ( .A(n12135), .B(n12349), .Z(n12128) );
  XNOR U12397 ( .A(n12134), .B(n12132), .Z(n12349) );
  AND U12398 ( .A(n12350), .B(n12351), .Z(n12132) );
  NANDN U12399 ( .A(n12352), .B(n12353), .Z(n12351) );
  OR U12400 ( .A(n12354), .B(n12355), .Z(n12353) );
  NAND U12401 ( .A(n12355), .B(n12354), .Z(n12350) );
  ANDN U12402 ( .B(B[16]), .A(n69), .Z(n12134) );
  XNOR U12403 ( .A(n12142), .B(n12356), .Z(n12135) );
  XNOR U12404 ( .A(n12141), .B(n12139), .Z(n12356) );
  AND U12405 ( .A(n12357), .B(n12358), .Z(n12139) );
  NANDN U12406 ( .A(n12359), .B(n12360), .Z(n12358) );
  NANDN U12407 ( .A(n12361), .B(n12362), .Z(n12360) );
  NANDN U12408 ( .A(n12362), .B(n12361), .Z(n12357) );
  ANDN U12409 ( .B(B[17]), .A(n70), .Z(n12141) );
  XNOR U12410 ( .A(n12149), .B(n12363), .Z(n12142) );
  XNOR U12411 ( .A(n12148), .B(n12146), .Z(n12363) );
  AND U12412 ( .A(n12364), .B(n12365), .Z(n12146) );
  NANDN U12413 ( .A(n12366), .B(n12367), .Z(n12365) );
  OR U12414 ( .A(n12368), .B(n12369), .Z(n12367) );
  NAND U12415 ( .A(n12369), .B(n12368), .Z(n12364) );
  ANDN U12416 ( .B(B[18]), .A(n71), .Z(n12148) );
  XNOR U12417 ( .A(n12156), .B(n12370), .Z(n12149) );
  XNOR U12418 ( .A(n12155), .B(n12153), .Z(n12370) );
  AND U12419 ( .A(n12371), .B(n12372), .Z(n12153) );
  NANDN U12420 ( .A(n12373), .B(n12374), .Z(n12372) );
  NANDN U12421 ( .A(n12375), .B(n12376), .Z(n12374) );
  NANDN U12422 ( .A(n12376), .B(n12375), .Z(n12371) );
  ANDN U12423 ( .B(B[19]), .A(n72), .Z(n12155) );
  XNOR U12424 ( .A(n12163), .B(n12377), .Z(n12156) );
  XNOR U12425 ( .A(n12162), .B(n12160), .Z(n12377) );
  AND U12426 ( .A(n12378), .B(n12379), .Z(n12160) );
  NANDN U12427 ( .A(n12380), .B(n12381), .Z(n12379) );
  OR U12428 ( .A(n12382), .B(n12383), .Z(n12381) );
  NAND U12429 ( .A(n12383), .B(n12382), .Z(n12378) );
  ANDN U12430 ( .B(B[20]), .A(n73), .Z(n12162) );
  XNOR U12431 ( .A(n12170), .B(n12384), .Z(n12163) );
  XNOR U12432 ( .A(n12169), .B(n12167), .Z(n12384) );
  AND U12433 ( .A(n12385), .B(n12386), .Z(n12167) );
  NANDN U12434 ( .A(n12387), .B(n12388), .Z(n12386) );
  NANDN U12435 ( .A(n12389), .B(n12390), .Z(n12388) );
  NANDN U12436 ( .A(n12390), .B(n12389), .Z(n12385) );
  ANDN U12437 ( .B(B[21]), .A(n74), .Z(n12169) );
  XNOR U12438 ( .A(n12177), .B(n12391), .Z(n12170) );
  XNOR U12439 ( .A(n12176), .B(n12174), .Z(n12391) );
  AND U12440 ( .A(n12392), .B(n12393), .Z(n12174) );
  NANDN U12441 ( .A(n12394), .B(n12395), .Z(n12393) );
  OR U12442 ( .A(n12396), .B(n12397), .Z(n12395) );
  NAND U12443 ( .A(n12397), .B(n12396), .Z(n12392) );
  ANDN U12444 ( .B(B[22]), .A(n75), .Z(n12176) );
  XNOR U12445 ( .A(n12184), .B(n12398), .Z(n12177) );
  XNOR U12446 ( .A(n12183), .B(n12181), .Z(n12398) );
  AND U12447 ( .A(n12399), .B(n12400), .Z(n12181) );
  NANDN U12448 ( .A(n12401), .B(n12402), .Z(n12400) );
  NANDN U12449 ( .A(n12403), .B(n12404), .Z(n12402) );
  NANDN U12450 ( .A(n12404), .B(n12403), .Z(n12399) );
  ANDN U12451 ( .B(B[23]), .A(n76), .Z(n12183) );
  XNOR U12452 ( .A(n12191), .B(n12405), .Z(n12184) );
  XNOR U12453 ( .A(n12190), .B(n12188), .Z(n12405) );
  AND U12454 ( .A(n12406), .B(n12407), .Z(n12188) );
  NANDN U12455 ( .A(n12408), .B(n12409), .Z(n12407) );
  OR U12456 ( .A(n12410), .B(n12411), .Z(n12409) );
  NAND U12457 ( .A(n12411), .B(n12410), .Z(n12406) );
  ANDN U12458 ( .B(B[24]), .A(n77), .Z(n12190) );
  XNOR U12459 ( .A(n12198), .B(n12412), .Z(n12191) );
  XNOR U12460 ( .A(n12197), .B(n12195), .Z(n12412) );
  AND U12461 ( .A(n12413), .B(n12414), .Z(n12195) );
  NANDN U12462 ( .A(n12415), .B(n12416), .Z(n12414) );
  NANDN U12463 ( .A(n12417), .B(n12418), .Z(n12416) );
  NANDN U12464 ( .A(n12418), .B(n12417), .Z(n12413) );
  ANDN U12465 ( .B(B[25]), .A(n78), .Z(n12197) );
  XNOR U12466 ( .A(n12205), .B(n12419), .Z(n12198) );
  XNOR U12467 ( .A(n12204), .B(n12202), .Z(n12419) );
  AND U12468 ( .A(n12420), .B(n12421), .Z(n12202) );
  NANDN U12469 ( .A(n12422), .B(n12423), .Z(n12421) );
  OR U12470 ( .A(n12424), .B(n12425), .Z(n12423) );
  NAND U12471 ( .A(n12425), .B(n12424), .Z(n12420) );
  ANDN U12472 ( .B(B[26]), .A(n79), .Z(n12204) );
  XNOR U12473 ( .A(n12212), .B(n12426), .Z(n12205) );
  XNOR U12474 ( .A(n12211), .B(n12209), .Z(n12426) );
  AND U12475 ( .A(n12427), .B(n12428), .Z(n12209) );
  NANDN U12476 ( .A(n12429), .B(n12430), .Z(n12428) );
  NANDN U12477 ( .A(n12431), .B(n12432), .Z(n12430) );
  NANDN U12478 ( .A(n12432), .B(n12431), .Z(n12427) );
  ANDN U12479 ( .B(B[27]), .A(n80), .Z(n12211) );
  XNOR U12480 ( .A(n12219), .B(n12433), .Z(n12212) );
  XNOR U12481 ( .A(n12218), .B(n12216), .Z(n12433) );
  AND U12482 ( .A(n12434), .B(n12435), .Z(n12216) );
  NANDN U12483 ( .A(n12436), .B(n12437), .Z(n12435) );
  OR U12484 ( .A(n12438), .B(n12439), .Z(n12437) );
  NAND U12485 ( .A(n12439), .B(n12438), .Z(n12434) );
  ANDN U12486 ( .B(B[28]), .A(n81), .Z(n12218) );
  XNOR U12487 ( .A(n12226), .B(n12440), .Z(n12219) );
  XNOR U12488 ( .A(n12225), .B(n12223), .Z(n12440) );
  AND U12489 ( .A(n12441), .B(n12442), .Z(n12223) );
  NANDN U12490 ( .A(n12443), .B(n12444), .Z(n12442) );
  NAND U12491 ( .A(n12445), .B(n12446), .Z(n12444) );
  ANDN U12492 ( .B(B[29]), .A(n82), .Z(n12225) );
  XOR U12493 ( .A(n12232), .B(n12447), .Z(n12226) );
  XNOR U12494 ( .A(n12230), .B(n12233), .Z(n12447) );
  NAND U12495 ( .A(A[2]), .B(B[30]), .Z(n12233) );
  NANDN U12496 ( .A(n12448), .B(n12449), .Z(n12230) );
  AND U12497 ( .A(A[0]), .B(B[31]), .Z(n12449) );
  XNOR U12498 ( .A(n12235), .B(n12450), .Z(n12232) );
  NAND U12499 ( .A(A[0]), .B(B[32]), .Z(n12450) );
  NAND U12500 ( .A(B[31]), .B(A[1]), .Z(n12235) );
  NAND U12501 ( .A(n12451), .B(n12452), .Z(n223) );
  NANDN U12502 ( .A(n12453), .B(n12454), .Z(n12452) );
  OR U12503 ( .A(n12455), .B(n12456), .Z(n12454) );
  NAND U12504 ( .A(n12456), .B(n12455), .Z(n12451) );
  XNOR U12505 ( .A(n12457), .B(n12458), .Z(\A1[2] ) );
  XNOR U12506 ( .A(n12459), .B(n12460), .Z(n12458) );
  XOR U12507 ( .A(n12456), .B(n12461), .Z(\A1[29] ) );
  XNOR U12508 ( .A(n12455), .B(n12453), .Z(n12461) );
  AND U12509 ( .A(n12462), .B(n12463), .Z(n12453) );
  NAND U12510 ( .A(n12464), .B(n12465), .Z(n12463) );
  NANDN U12511 ( .A(n12466), .B(n12467), .Z(n12464) );
  NANDN U12512 ( .A(n12467), .B(n12466), .Z(n12462) );
  ANDN U12513 ( .B(B[0]), .A(n54), .Z(n12455) );
  XNOR U12514 ( .A(n12250), .B(n12468), .Z(n12456) );
  XNOR U12515 ( .A(n12249), .B(n12247), .Z(n12468) );
  AND U12516 ( .A(n12469), .B(n12470), .Z(n12247) );
  NANDN U12517 ( .A(n12471), .B(n12472), .Z(n12470) );
  OR U12518 ( .A(n12473), .B(n12474), .Z(n12472) );
  NAND U12519 ( .A(n12474), .B(n12473), .Z(n12469) );
  ANDN U12520 ( .B(B[1]), .A(n55), .Z(n12249) );
  XNOR U12521 ( .A(n12257), .B(n12475), .Z(n12250) );
  XNOR U12522 ( .A(n12256), .B(n12254), .Z(n12475) );
  AND U12523 ( .A(n12476), .B(n12477), .Z(n12254) );
  NANDN U12524 ( .A(n12478), .B(n12479), .Z(n12477) );
  NANDN U12525 ( .A(n12480), .B(n12481), .Z(n12479) );
  NANDN U12526 ( .A(n12481), .B(n12480), .Z(n12476) );
  ANDN U12527 ( .B(B[2]), .A(n56), .Z(n12256) );
  XNOR U12528 ( .A(n12264), .B(n12482), .Z(n12257) );
  XNOR U12529 ( .A(n12263), .B(n12261), .Z(n12482) );
  AND U12530 ( .A(n12483), .B(n12484), .Z(n12261) );
  NANDN U12531 ( .A(n12485), .B(n12486), .Z(n12484) );
  OR U12532 ( .A(n12487), .B(n12488), .Z(n12486) );
  NAND U12533 ( .A(n12488), .B(n12487), .Z(n12483) );
  ANDN U12534 ( .B(B[3]), .A(n57), .Z(n12263) );
  XNOR U12535 ( .A(n12271), .B(n12489), .Z(n12264) );
  XNOR U12536 ( .A(n12270), .B(n12268), .Z(n12489) );
  AND U12537 ( .A(n12490), .B(n12491), .Z(n12268) );
  NANDN U12538 ( .A(n12492), .B(n12493), .Z(n12491) );
  NANDN U12539 ( .A(n12494), .B(n12495), .Z(n12493) );
  NANDN U12540 ( .A(n12495), .B(n12494), .Z(n12490) );
  ANDN U12541 ( .B(B[4]), .A(n58), .Z(n12270) );
  XNOR U12542 ( .A(n12278), .B(n12496), .Z(n12271) );
  XNOR U12543 ( .A(n12277), .B(n12275), .Z(n12496) );
  AND U12544 ( .A(n12497), .B(n12498), .Z(n12275) );
  NANDN U12545 ( .A(n12499), .B(n12500), .Z(n12498) );
  OR U12546 ( .A(n12501), .B(n12502), .Z(n12500) );
  NAND U12547 ( .A(n12502), .B(n12501), .Z(n12497) );
  ANDN U12548 ( .B(B[5]), .A(n59), .Z(n12277) );
  XNOR U12549 ( .A(n12285), .B(n12503), .Z(n12278) );
  XNOR U12550 ( .A(n12284), .B(n12282), .Z(n12503) );
  AND U12551 ( .A(n12504), .B(n12505), .Z(n12282) );
  NANDN U12552 ( .A(n12506), .B(n12507), .Z(n12505) );
  NANDN U12553 ( .A(n12508), .B(n12509), .Z(n12507) );
  NANDN U12554 ( .A(n12509), .B(n12508), .Z(n12504) );
  ANDN U12555 ( .B(B[6]), .A(n60), .Z(n12284) );
  XNOR U12556 ( .A(n12292), .B(n12510), .Z(n12285) );
  XNOR U12557 ( .A(n12291), .B(n12289), .Z(n12510) );
  AND U12558 ( .A(n12511), .B(n12512), .Z(n12289) );
  NANDN U12559 ( .A(n12513), .B(n12514), .Z(n12512) );
  OR U12560 ( .A(n12515), .B(n12516), .Z(n12514) );
  NAND U12561 ( .A(n12516), .B(n12515), .Z(n12511) );
  ANDN U12562 ( .B(B[7]), .A(n61), .Z(n12291) );
  XNOR U12563 ( .A(n12299), .B(n12517), .Z(n12292) );
  XNOR U12564 ( .A(n12298), .B(n12296), .Z(n12517) );
  AND U12565 ( .A(n12518), .B(n12519), .Z(n12296) );
  NANDN U12566 ( .A(n12520), .B(n12521), .Z(n12519) );
  NANDN U12567 ( .A(n12522), .B(n12523), .Z(n12521) );
  NANDN U12568 ( .A(n12523), .B(n12522), .Z(n12518) );
  ANDN U12569 ( .B(B[8]), .A(n62), .Z(n12298) );
  XNOR U12570 ( .A(n12306), .B(n12524), .Z(n12299) );
  XNOR U12571 ( .A(n12305), .B(n12303), .Z(n12524) );
  AND U12572 ( .A(n12525), .B(n12526), .Z(n12303) );
  NANDN U12573 ( .A(n12527), .B(n12528), .Z(n12526) );
  OR U12574 ( .A(n12529), .B(n12530), .Z(n12528) );
  NAND U12575 ( .A(n12530), .B(n12529), .Z(n12525) );
  ANDN U12576 ( .B(B[9]), .A(n63), .Z(n12305) );
  XNOR U12577 ( .A(n12313), .B(n12531), .Z(n12306) );
  XNOR U12578 ( .A(n12312), .B(n12310), .Z(n12531) );
  AND U12579 ( .A(n12532), .B(n12533), .Z(n12310) );
  NANDN U12580 ( .A(n12534), .B(n12535), .Z(n12533) );
  NANDN U12581 ( .A(n12536), .B(n12537), .Z(n12535) );
  NANDN U12582 ( .A(n12537), .B(n12536), .Z(n12532) );
  ANDN U12583 ( .B(B[10]), .A(n64), .Z(n12312) );
  XNOR U12584 ( .A(n12320), .B(n12538), .Z(n12313) );
  XNOR U12585 ( .A(n12319), .B(n12317), .Z(n12538) );
  AND U12586 ( .A(n12539), .B(n12540), .Z(n12317) );
  NANDN U12587 ( .A(n12541), .B(n12542), .Z(n12540) );
  OR U12588 ( .A(n12543), .B(n12544), .Z(n12542) );
  NAND U12589 ( .A(n12544), .B(n12543), .Z(n12539) );
  ANDN U12590 ( .B(B[11]), .A(n65), .Z(n12319) );
  XNOR U12591 ( .A(n12327), .B(n12545), .Z(n12320) );
  XNOR U12592 ( .A(n12326), .B(n12324), .Z(n12545) );
  AND U12593 ( .A(n12546), .B(n12547), .Z(n12324) );
  NANDN U12594 ( .A(n12548), .B(n12549), .Z(n12547) );
  NANDN U12595 ( .A(n12550), .B(n12551), .Z(n12549) );
  NANDN U12596 ( .A(n12551), .B(n12550), .Z(n12546) );
  ANDN U12597 ( .B(B[12]), .A(n66), .Z(n12326) );
  XNOR U12598 ( .A(n12334), .B(n12552), .Z(n12327) );
  XNOR U12599 ( .A(n12333), .B(n12331), .Z(n12552) );
  AND U12600 ( .A(n12553), .B(n12554), .Z(n12331) );
  NANDN U12601 ( .A(n12555), .B(n12556), .Z(n12554) );
  OR U12602 ( .A(n12557), .B(n12558), .Z(n12556) );
  NAND U12603 ( .A(n12558), .B(n12557), .Z(n12553) );
  ANDN U12604 ( .B(B[13]), .A(n67), .Z(n12333) );
  XNOR U12605 ( .A(n12341), .B(n12559), .Z(n12334) );
  XNOR U12606 ( .A(n12340), .B(n12338), .Z(n12559) );
  AND U12607 ( .A(n12560), .B(n12561), .Z(n12338) );
  NANDN U12608 ( .A(n12562), .B(n12563), .Z(n12561) );
  NANDN U12609 ( .A(n12564), .B(n12565), .Z(n12563) );
  NANDN U12610 ( .A(n12565), .B(n12564), .Z(n12560) );
  ANDN U12611 ( .B(B[14]), .A(n68), .Z(n12340) );
  XNOR U12612 ( .A(n12348), .B(n12566), .Z(n12341) );
  XNOR U12613 ( .A(n12347), .B(n12345), .Z(n12566) );
  AND U12614 ( .A(n12567), .B(n12568), .Z(n12345) );
  NANDN U12615 ( .A(n12569), .B(n12570), .Z(n12568) );
  OR U12616 ( .A(n12571), .B(n12572), .Z(n12570) );
  NAND U12617 ( .A(n12572), .B(n12571), .Z(n12567) );
  ANDN U12618 ( .B(B[15]), .A(n69), .Z(n12347) );
  XNOR U12619 ( .A(n12355), .B(n12573), .Z(n12348) );
  XNOR U12620 ( .A(n12354), .B(n12352), .Z(n12573) );
  AND U12621 ( .A(n12574), .B(n12575), .Z(n12352) );
  NANDN U12622 ( .A(n12576), .B(n12577), .Z(n12575) );
  NANDN U12623 ( .A(n12578), .B(n12579), .Z(n12577) );
  NANDN U12624 ( .A(n12579), .B(n12578), .Z(n12574) );
  ANDN U12625 ( .B(B[16]), .A(n70), .Z(n12354) );
  XNOR U12626 ( .A(n12362), .B(n12580), .Z(n12355) );
  XNOR U12627 ( .A(n12361), .B(n12359), .Z(n12580) );
  AND U12628 ( .A(n12581), .B(n12582), .Z(n12359) );
  NANDN U12629 ( .A(n12583), .B(n12584), .Z(n12582) );
  OR U12630 ( .A(n12585), .B(n12586), .Z(n12584) );
  NAND U12631 ( .A(n12586), .B(n12585), .Z(n12581) );
  ANDN U12632 ( .B(B[17]), .A(n71), .Z(n12361) );
  XNOR U12633 ( .A(n12369), .B(n12587), .Z(n12362) );
  XNOR U12634 ( .A(n12368), .B(n12366), .Z(n12587) );
  AND U12635 ( .A(n12588), .B(n12589), .Z(n12366) );
  NANDN U12636 ( .A(n12590), .B(n12591), .Z(n12589) );
  NANDN U12637 ( .A(n12592), .B(n12593), .Z(n12591) );
  NANDN U12638 ( .A(n12593), .B(n12592), .Z(n12588) );
  ANDN U12639 ( .B(B[18]), .A(n72), .Z(n12368) );
  XNOR U12640 ( .A(n12376), .B(n12594), .Z(n12369) );
  XNOR U12641 ( .A(n12375), .B(n12373), .Z(n12594) );
  AND U12642 ( .A(n12595), .B(n12596), .Z(n12373) );
  NANDN U12643 ( .A(n12597), .B(n12598), .Z(n12596) );
  OR U12644 ( .A(n12599), .B(n12600), .Z(n12598) );
  NAND U12645 ( .A(n12600), .B(n12599), .Z(n12595) );
  ANDN U12646 ( .B(B[19]), .A(n73), .Z(n12375) );
  XNOR U12647 ( .A(n12383), .B(n12601), .Z(n12376) );
  XNOR U12648 ( .A(n12382), .B(n12380), .Z(n12601) );
  AND U12649 ( .A(n12602), .B(n12603), .Z(n12380) );
  NANDN U12650 ( .A(n12604), .B(n12605), .Z(n12603) );
  NANDN U12651 ( .A(n12606), .B(n12607), .Z(n12605) );
  NANDN U12652 ( .A(n12607), .B(n12606), .Z(n12602) );
  ANDN U12653 ( .B(B[20]), .A(n74), .Z(n12382) );
  XNOR U12654 ( .A(n12390), .B(n12608), .Z(n12383) );
  XNOR U12655 ( .A(n12389), .B(n12387), .Z(n12608) );
  AND U12656 ( .A(n12609), .B(n12610), .Z(n12387) );
  NANDN U12657 ( .A(n12611), .B(n12612), .Z(n12610) );
  OR U12658 ( .A(n12613), .B(n12614), .Z(n12612) );
  NAND U12659 ( .A(n12614), .B(n12613), .Z(n12609) );
  ANDN U12660 ( .B(B[21]), .A(n75), .Z(n12389) );
  XNOR U12661 ( .A(n12397), .B(n12615), .Z(n12390) );
  XNOR U12662 ( .A(n12396), .B(n12394), .Z(n12615) );
  AND U12663 ( .A(n12616), .B(n12617), .Z(n12394) );
  NANDN U12664 ( .A(n12618), .B(n12619), .Z(n12617) );
  NANDN U12665 ( .A(n12620), .B(n12621), .Z(n12619) );
  NANDN U12666 ( .A(n12621), .B(n12620), .Z(n12616) );
  ANDN U12667 ( .B(B[22]), .A(n76), .Z(n12396) );
  XNOR U12668 ( .A(n12404), .B(n12622), .Z(n12397) );
  XNOR U12669 ( .A(n12403), .B(n12401), .Z(n12622) );
  AND U12670 ( .A(n12623), .B(n12624), .Z(n12401) );
  NANDN U12671 ( .A(n12625), .B(n12626), .Z(n12624) );
  OR U12672 ( .A(n12627), .B(n12628), .Z(n12626) );
  NAND U12673 ( .A(n12628), .B(n12627), .Z(n12623) );
  ANDN U12674 ( .B(B[23]), .A(n77), .Z(n12403) );
  XNOR U12675 ( .A(n12411), .B(n12629), .Z(n12404) );
  XNOR U12676 ( .A(n12410), .B(n12408), .Z(n12629) );
  AND U12677 ( .A(n12630), .B(n12631), .Z(n12408) );
  NANDN U12678 ( .A(n12632), .B(n12633), .Z(n12631) );
  NANDN U12679 ( .A(n12634), .B(n12635), .Z(n12633) );
  NANDN U12680 ( .A(n12635), .B(n12634), .Z(n12630) );
  ANDN U12681 ( .B(B[24]), .A(n78), .Z(n12410) );
  XNOR U12682 ( .A(n12418), .B(n12636), .Z(n12411) );
  XNOR U12683 ( .A(n12417), .B(n12415), .Z(n12636) );
  AND U12684 ( .A(n12637), .B(n12638), .Z(n12415) );
  NANDN U12685 ( .A(n12639), .B(n12640), .Z(n12638) );
  OR U12686 ( .A(n12641), .B(n12642), .Z(n12640) );
  NAND U12687 ( .A(n12642), .B(n12641), .Z(n12637) );
  ANDN U12688 ( .B(B[25]), .A(n79), .Z(n12417) );
  XNOR U12689 ( .A(n12425), .B(n12643), .Z(n12418) );
  XNOR U12690 ( .A(n12424), .B(n12422), .Z(n12643) );
  AND U12691 ( .A(n12644), .B(n12645), .Z(n12422) );
  NANDN U12692 ( .A(n12646), .B(n12647), .Z(n12645) );
  NANDN U12693 ( .A(n12648), .B(n12649), .Z(n12647) );
  NANDN U12694 ( .A(n12649), .B(n12648), .Z(n12644) );
  ANDN U12695 ( .B(B[26]), .A(n80), .Z(n12424) );
  XNOR U12696 ( .A(n12432), .B(n12650), .Z(n12425) );
  XNOR U12697 ( .A(n12431), .B(n12429), .Z(n12650) );
  AND U12698 ( .A(n12651), .B(n12652), .Z(n12429) );
  NANDN U12699 ( .A(n12653), .B(n12654), .Z(n12652) );
  OR U12700 ( .A(n12655), .B(n12656), .Z(n12654) );
  NAND U12701 ( .A(n12656), .B(n12655), .Z(n12651) );
  ANDN U12702 ( .B(B[27]), .A(n81), .Z(n12431) );
  XNOR U12703 ( .A(n12439), .B(n12657), .Z(n12432) );
  XNOR U12704 ( .A(n12438), .B(n12436), .Z(n12657) );
  AND U12705 ( .A(n12658), .B(n12659), .Z(n12436) );
  NANDN U12706 ( .A(n12660), .B(n12661), .Z(n12659) );
  NAND U12707 ( .A(n12662), .B(n12663), .Z(n12661) );
  ANDN U12708 ( .B(B[28]), .A(n82), .Z(n12438) );
  XOR U12709 ( .A(n12445), .B(n12664), .Z(n12439) );
  XNOR U12710 ( .A(n12443), .B(n12446), .Z(n12664) );
  NAND U12711 ( .A(A[2]), .B(B[29]), .Z(n12446) );
  NANDN U12712 ( .A(n12665), .B(n12666), .Z(n12443) );
  AND U12713 ( .A(A[0]), .B(B[30]), .Z(n12666) );
  XNOR U12714 ( .A(n12448), .B(n12667), .Z(n12445) );
  NAND U12715 ( .A(A[0]), .B(B[31]), .Z(n12667) );
  NAND U12716 ( .A(B[30]), .B(A[1]), .Z(n12448) );
  XOR U12717 ( .A(n12467), .B(n12668), .Z(\A1[28] ) );
  XNOR U12718 ( .A(n12466), .B(n12465), .Z(n12668) );
  NAND U12719 ( .A(n12669), .B(n12670), .Z(n12465) );
  NANDN U12720 ( .A(n12671), .B(n12672), .Z(n12670) );
  OR U12721 ( .A(n12673), .B(n12674), .Z(n12672) );
  NAND U12722 ( .A(n12674), .B(n12673), .Z(n12669) );
  ANDN U12723 ( .B(B[0]), .A(n55), .Z(n12466) );
  XNOR U12724 ( .A(n12474), .B(n12675), .Z(n12467) );
  XNOR U12725 ( .A(n12473), .B(n12471), .Z(n12675) );
  AND U12726 ( .A(n12676), .B(n12677), .Z(n12471) );
  NANDN U12727 ( .A(n12678), .B(n12679), .Z(n12677) );
  NANDN U12728 ( .A(n12680), .B(n12681), .Z(n12679) );
  NANDN U12729 ( .A(n12681), .B(n12680), .Z(n12676) );
  ANDN U12730 ( .B(B[1]), .A(n56), .Z(n12473) );
  XNOR U12731 ( .A(n12481), .B(n12682), .Z(n12474) );
  XNOR U12732 ( .A(n12480), .B(n12478), .Z(n12682) );
  AND U12733 ( .A(n12683), .B(n12684), .Z(n12478) );
  NANDN U12734 ( .A(n12685), .B(n12686), .Z(n12684) );
  OR U12735 ( .A(n12687), .B(n12688), .Z(n12686) );
  NAND U12736 ( .A(n12688), .B(n12687), .Z(n12683) );
  ANDN U12737 ( .B(B[2]), .A(n57), .Z(n12480) );
  XNOR U12738 ( .A(n12488), .B(n12689), .Z(n12481) );
  XNOR U12739 ( .A(n12487), .B(n12485), .Z(n12689) );
  AND U12740 ( .A(n12690), .B(n12691), .Z(n12485) );
  NANDN U12741 ( .A(n12692), .B(n12693), .Z(n12691) );
  NANDN U12742 ( .A(n12694), .B(n12695), .Z(n12693) );
  NANDN U12743 ( .A(n12695), .B(n12694), .Z(n12690) );
  ANDN U12744 ( .B(B[3]), .A(n58), .Z(n12487) );
  XNOR U12745 ( .A(n12495), .B(n12696), .Z(n12488) );
  XNOR U12746 ( .A(n12494), .B(n12492), .Z(n12696) );
  AND U12747 ( .A(n12697), .B(n12698), .Z(n12492) );
  NANDN U12748 ( .A(n12699), .B(n12700), .Z(n12698) );
  OR U12749 ( .A(n12701), .B(n12702), .Z(n12700) );
  NAND U12750 ( .A(n12702), .B(n12701), .Z(n12697) );
  ANDN U12751 ( .B(B[4]), .A(n59), .Z(n12494) );
  XNOR U12752 ( .A(n12502), .B(n12703), .Z(n12495) );
  XNOR U12753 ( .A(n12501), .B(n12499), .Z(n12703) );
  AND U12754 ( .A(n12704), .B(n12705), .Z(n12499) );
  NANDN U12755 ( .A(n12706), .B(n12707), .Z(n12705) );
  NANDN U12756 ( .A(n12708), .B(n12709), .Z(n12707) );
  NANDN U12757 ( .A(n12709), .B(n12708), .Z(n12704) );
  ANDN U12758 ( .B(B[5]), .A(n60), .Z(n12501) );
  XNOR U12759 ( .A(n12509), .B(n12710), .Z(n12502) );
  XNOR U12760 ( .A(n12508), .B(n12506), .Z(n12710) );
  AND U12761 ( .A(n12711), .B(n12712), .Z(n12506) );
  NANDN U12762 ( .A(n12713), .B(n12714), .Z(n12712) );
  OR U12763 ( .A(n12715), .B(n12716), .Z(n12714) );
  NAND U12764 ( .A(n12716), .B(n12715), .Z(n12711) );
  ANDN U12765 ( .B(B[6]), .A(n61), .Z(n12508) );
  XNOR U12766 ( .A(n12516), .B(n12717), .Z(n12509) );
  XNOR U12767 ( .A(n12515), .B(n12513), .Z(n12717) );
  AND U12768 ( .A(n12718), .B(n12719), .Z(n12513) );
  NANDN U12769 ( .A(n12720), .B(n12721), .Z(n12719) );
  NANDN U12770 ( .A(n12722), .B(n12723), .Z(n12721) );
  NANDN U12771 ( .A(n12723), .B(n12722), .Z(n12718) );
  ANDN U12772 ( .B(B[7]), .A(n62), .Z(n12515) );
  XNOR U12773 ( .A(n12523), .B(n12724), .Z(n12516) );
  XNOR U12774 ( .A(n12522), .B(n12520), .Z(n12724) );
  AND U12775 ( .A(n12725), .B(n12726), .Z(n12520) );
  NANDN U12776 ( .A(n12727), .B(n12728), .Z(n12726) );
  OR U12777 ( .A(n12729), .B(n12730), .Z(n12728) );
  NAND U12778 ( .A(n12730), .B(n12729), .Z(n12725) );
  ANDN U12779 ( .B(B[8]), .A(n63), .Z(n12522) );
  XNOR U12780 ( .A(n12530), .B(n12731), .Z(n12523) );
  XNOR U12781 ( .A(n12529), .B(n12527), .Z(n12731) );
  AND U12782 ( .A(n12732), .B(n12733), .Z(n12527) );
  NANDN U12783 ( .A(n12734), .B(n12735), .Z(n12733) );
  NANDN U12784 ( .A(n12736), .B(n12737), .Z(n12735) );
  NANDN U12785 ( .A(n12737), .B(n12736), .Z(n12732) );
  ANDN U12786 ( .B(B[9]), .A(n64), .Z(n12529) );
  XNOR U12787 ( .A(n12537), .B(n12738), .Z(n12530) );
  XNOR U12788 ( .A(n12536), .B(n12534), .Z(n12738) );
  AND U12789 ( .A(n12739), .B(n12740), .Z(n12534) );
  NANDN U12790 ( .A(n12741), .B(n12742), .Z(n12740) );
  OR U12791 ( .A(n12743), .B(n12744), .Z(n12742) );
  NAND U12792 ( .A(n12744), .B(n12743), .Z(n12739) );
  ANDN U12793 ( .B(B[10]), .A(n65), .Z(n12536) );
  XNOR U12794 ( .A(n12544), .B(n12745), .Z(n12537) );
  XNOR U12795 ( .A(n12543), .B(n12541), .Z(n12745) );
  AND U12796 ( .A(n12746), .B(n12747), .Z(n12541) );
  NANDN U12797 ( .A(n12748), .B(n12749), .Z(n12747) );
  NANDN U12798 ( .A(n12750), .B(n12751), .Z(n12749) );
  NANDN U12799 ( .A(n12751), .B(n12750), .Z(n12746) );
  ANDN U12800 ( .B(B[11]), .A(n66), .Z(n12543) );
  XNOR U12801 ( .A(n12551), .B(n12752), .Z(n12544) );
  XNOR U12802 ( .A(n12550), .B(n12548), .Z(n12752) );
  AND U12803 ( .A(n12753), .B(n12754), .Z(n12548) );
  NANDN U12804 ( .A(n12755), .B(n12756), .Z(n12754) );
  OR U12805 ( .A(n12757), .B(n12758), .Z(n12756) );
  NAND U12806 ( .A(n12758), .B(n12757), .Z(n12753) );
  ANDN U12807 ( .B(B[12]), .A(n67), .Z(n12550) );
  XNOR U12808 ( .A(n12558), .B(n12759), .Z(n12551) );
  XNOR U12809 ( .A(n12557), .B(n12555), .Z(n12759) );
  AND U12810 ( .A(n12760), .B(n12761), .Z(n12555) );
  NANDN U12811 ( .A(n12762), .B(n12763), .Z(n12761) );
  NANDN U12812 ( .A(n12764), .B(n12765), .Z(n12763) );
  NANDN U12813 ( .A(n12765), .B(n12764), .Z(n12760) );
  ANDN U12814 ( .B(B[13]), .A(n68), .Z(n12557) );
  XNOR U12815 ( .A(n12565), .B(n12766), .Z(n12558) );
  XNOR U12816 ( .A(n12564), .B(n12562), .Z(n12766) );
  AND U12817 ( .A(n12767), .B(n12768), .Z(n12562) );
  NANDN U12818 ( .A(n12769), .B(n12770), .Z(n12768) );
  OR U12819 ( .A(n12771), .B(n12772), .Z(n12770) );
  NAND U12820 ( .A(n12772), .B(n12771), .Z(n12767) );
  ANDN U12821 ( .B(B[14]), .A(n69), .Z(n12564) );
  XNOR U12822 ( .A(n12572), .B(n12773), .Z(n12565) );
  XNOR U12823 ( .A(n12571), .B(n12569), .Z(n12773) );
  AND U12824 ( .A(n12774), .B(n12775), .Z(n12569) );
  NANDN U12825 ( .A(n12776), .B(n12777), .Z(n12775) );
  NANDN U12826 ( .A(n12778), .B(n12779), .Z(n12777) );
  NANDN U12827 ( .A(n12779), .B(n12778), .Z(n12774) );
  ANDN U12828 ( .B(B[15]), .A(n70), .Z(n12571) );
  XNOR U12829 ( .A(n12579), .B(n12780), .Z(n12572) );
  XNOR U12830 ( .A(n12578), .B(n12576), .Z(n12780) );
  AND U12831 ( .A(n12781), .B(n12782), .Z(n12576) );
  NANDN U12832 ( .A(n12783), .B(n12784), .Z(n12782) );
  OR U12833 ( .A(n12785), .B(n12786), .Z(n12784) );
  NAND U12834 ( .A(n12786), .B(n12785), .Z(n12781) );
  ANDN U12835 ( .B(B[16]), .A(n71), .Z(n12578) );
  XNOR U12836 ( .A(n12586), .B(n12787), .Z(n12579) );
  XNOR U12837 ( .A(n12585), .B(n12583), .Z(n12787) );
  AND U12838 ( .A(n12788), .B(n12789), .Z(n12583) );
  NANDN U12839 ( .A(n12790), .B(n12791), .Z(n12789) );
  NANDN U12840 ( .A(n12792), .B(n12793), .Z(n12791) );
  NANDN U12841 ( .A(n12793), .B(n12792), .Z(n12788) );
  ANDN U12842 ( .B(B[17]), .A(n72), .Z(n12585) );
  XNOR U12843 ( .A(n12593), .B(n12794), .Z(n12586) );
  XNOR U12844 ( .A(n12592), .B(n12590), .Z(n12794) );
  AND U12845 ( .A(n12795), .B(n12796), .Z(n12590) );
  NANDN U12846 ( .A(n12797), .B(n12798), .Z(n12796) );
  OR U12847 ( .A(n12799), .B(n12800), .Z(n12798) );
  NAND U12848 ( .A(n12800), .B(n12799), .Z(n12795) );
  ANDN U12849 ( .B(B[18]), .A(n73), .Z(n12592) );
  XNOR U12850 ( .A(n12600), .B(n12801), .Z(n12593) );
  XNOR U12851 ( .A(n12599), .B(n12597), .Z(n12801) );
  AND U12852 ( .A(n12802), .B(n12803), .Z(n12597) );
  NANDN U12853 ( .A(n12804), .B(n12805), .Z(n12803) );
  NANDN U12854 ( .A(n12806), .B(n12807), .Z(n12805) );
  NANDN U12855 ( .A(n12807), .B(n12806), .Z(n12802) );
  ANDN U12856 ( .B(B[19]), .A(n74), .Z(n12599) );
  XNOR U12857 ( .A(n12607), .B(n12808), .Z(n12600) );
  XNOR U12858 ( .A(n12606), .B(n12604), .Z(n12808) );
  AND U12859 ( .A(n12809), .B(n12810), .Z(n12604) );
  NANDN U12860 ( .A(n12811), .B(n12812), .Z(n12810) );
  OR U12861 ( .A(n12813), .B(n12814), .Z(n12812) );
  NAND U12862 ( .A(n12814), .B(n12813), .Z(n12809) );
  ANDN U12863 ( .B(B[20]), .A(n75), .Z(n12606) );
  XNOR U12864 ( .A(n12614), .B(n12815), .Z(n12607) );
  XNOR U12865 ( .A(n12613), .B(n12611), .Z(n12815) );
  AND U12866 ( .A(n12816), .B(n12817), .Z(n12611) );
  NANDN U12867 ( .A(n12818), .B(n12819), .Z(n12817) );
  NANDN U12868 ( .A(n12820), .B(n12821), .Z(n12819) );
  NANDN U12869 ( .A(n12821), .B(n12820), .Z(n12816) );
  ANDN U12870 ( .B(B[21]), .A(n76), .Z(n12613) );
  XNOR U12871 ( .A(n12621), .B(n12822), .Z(n12614) );
  XNOR U12872 ( .A(n12620), .B(n12618), .Z(n12822) );
  AND U12873 ( .A(n12823), .B(n12824), .Z(n12618) );
  NANDN U12874 ( .A(n12825), .B(n12826), .Z(n12824) );
  OR U12875 ( .A(n12827), .B(n12828), .Z(n12826) );
  NAND U12876 ( .A(n12828), .B(n12827), .Z(n12823) );
  ANDN U12877 ( .B(B[22]), .A(n77), .Z(n12620) );
  XNOR U12878 ( .A(n12628), .B(n12829), .Z(n12621) );
  XNOR U12879 ( .A(n12627), .B(n12625), .Z(n12829) );
  AND U12880 ( .A(n12830), .B(n12831), .Z(n12625) );
  NANDN U12881 ( .A(n12832), .B(n12833), .Z(n12831) );
  NANDN U12882 ( .A(n12834), .B(n12835), .Z(n12833) );
  NANDN U12883 ( .A(n12835), .B(n12834), .Z(n12830) );
  ANDN U12884 ( .B(B[23]), .A(n78), .Z(n12627) );
  XNOR U12885 ( .A(n12635), .B(n12836), .Z(n12628) );
  XNOR U12886 ( .A(n12634), .B(n12632), .Z(n12836) );
  AND U12887 ( .A(n12837), .B(n12838), .Z(n12632) );
  NANDN U12888 ( .A(n12839), .B(n12840), .Z(n12838) );
  OR U12889 ( .A(n12841), .B(n12842), .Z(n12840) );
  NAND U12890 ( .A(n12842), .B(n12841), .Z(n12837) );
  ANDN U12891 ( .B(B[24]), .A(n79), .Z(n12634) );
  XNOR U12892 ( .A(n12642), .B(n12843), .Z(n12635) );
  XNOR U12893 ( .A(n12641), .B(n12639), .Z(n12843) );
  AND U12894 ( .A(n12844), .B(n12845), .Z(n12639) );
  NANDN U12895 ( .A(n12846), .B(n12847), .Z(n12845) );
  NANDN U12896 ( .A(n12848), .B(n12849), .Z(n12847) );
  NANDN U12897 ( .A(n12849), .B(n12848), .Z(n12844) );
  ANDN U12898 ( .B(B[25]), .A(n80), .Z(n12641) );
  XNOR U12899 ( .A(n12649), .B(n12850), .Z(n12642) );
  XNOR U12900 ( .A(n12648), .B(n12646), .Z(n12850) );
  AND U12901 ( .A(n12851), .B(n12852), .Z(n12646) );
  NANDN U12902 ( .A(n12853), .B(n12854), .Z(n12852) );
  OR U12903 ( .A(n12855), .B(n12856), .Z(n12854) );
  NAND U12904 ( .A(n12856), .B(n12855), .Z(n12851) );
  ANDN U12905 ( .B(B[26]), .A(n81), .Z(n12648) );
  XNOR U12906 ( .A(n12656), .B(n12857), .Z(n12649) );
  XNOR U12907 ( .A(n12655), .B(n12653), .Z(n12857) );
  AND U12908 ( .A(n12858), .B(n12859), .Z(n12653) );
  NANDN U12909 ( .A(n12860), .B(n12861), .Z(n12859) );
  NAND U12910 ( .A(n12862), .B(n12863), .Z(n12861) );
  ANDN U12911 ( .B(B[27]), .A(n82), .Z(n12655) );
  XOR U12912 ( .A(n12662), .B(n12864), .Z(n12656) );
  XNOR U12913 ( .A(n12660), .B(n12663), .Z(n12864) );
  NAND U12914 ( .A(A[2]), .B(B[28]), .Z(n12663) );
  NANDN U12915 ( .A(n12865), .B(n12866), .Z(n12660) );
  AND U12916 ( .A(A[0]), .B(B[29]), .Z(n12866) );
  XNOR U12917 ( .A(n12665), .B(n12867), .Z(n12662) );
  NAND U12918 ( .A(A[0]), .B(B[30]), .Z(n12867) );
  NAND U12919 ( .A(B[29]), .B(A[1]), .Z(n12665) );
  XNOR U12921 ( .A(n224), .B(n12868), .Z(\A1[284] ) );
  NAND U12922 ( .A(A[31]), .B(B[255]), .Z(n12868) );
  NAND U12923 ( .A(n12869), .B(n12870), .Z(n224) );
  NAND U12924 ( .A(n12871), .B(n12872), .Z(n12870) );
  NANDN U12925 ( .A(n12873), .B(n12874), .Z(n12871) );
  NANDN U12926 ( .A(n12874), .B(n12873), .Z(n12869) );
  XOR U12927 ( .A(n226), .B(n225), .Z(\A1[283] ) );
  XNOR U12928 ( .A(n12872), .B(n12875), .Z(n225) );
  XOR U12929 ( .A(n12873), .B(n12874), .Z(n12875) );
  NAND U12930 ( .A(A[30]), .B(B[255]), .Z(n12874) );
  AND U12931 ( .A(B[254]), .B(A[31]), .Z(n12873) );
  NAND U12932 ( .A(n12876), .B(n12877), .Z(n12872) );
  NAND U12933 ( .A(n12878), .B(n12879), .Z(n12877) );
  NANDN U12934 ( .A(n12880), .B(n12881), .Z(n12878) );
  NANDN U12935 ( .A(n12881), .B(n12880), .Z(n12876) );
  NAND U12936 ( .A(n12882), .B(n12883), .Z(n226) );
  NANDN U12937 ( .A(n12884), .B(n12885), .Z(n12883) );
  NAND U12938 ( .A(n12887), .B(n12886), .Z(n12882) );
  XOR U12939 ( .A(n228), .B(n227), .Z(\A1[282] ) );
  XOR U12940 ( .A(n12887), .B(n12888), .Z(n227) );
  XNOR U12941 ( .A(n12886), .B(n12884), .Z(n12888) );
  AND U12942 ( .A(n12889), .B(n12890), .Z(n12884) );
  NANDN U12943 ( .A(n12891), .B(n12892), .Z(n12890) );
  NANDN U12944 ( .A(n12893), .B(n12894), .Z(n12892) );
  NANDN U12945 ( .A(n12894), .B(n12893), .Z(n12889) );
  ANDN U12946 ( .B(B[253]), .A(n54), .Z(n12886) );
  XNOR U12947 ( .A(n12879), .B(n12895), .Z(n12887) );
  XOR U12948 ( .A(n12880), .B(n12881), .Z(n12895) );
  NAND U12949 ( .A(A[29]), .B(B[255]), .Z(n12881) );
  AND U12950 ( .A(B[254]), .B(A[30]), .Z(n12880) );
  NAND U12951 ( .A(n12896), .B(n12897), .Z(n12879) );
  NAND U12952 ( .A(n12898), .B(n12899), .Z(n12897) );
  NANDN U12953 ( .A(n12900), .B(n12901), .Z(n12898) );
  NANDN U12954 ( .A(n12901), .B(n12900), .Z(n12896) );
  NAND U12955 ( .A(n12902), .B(n12903), .Z(n228) );
  NANDN U12956 ( .A(n12904), .B(n12905), .Z(n12903) );
  OR U12957 ( .A(n12906), .B(n12907), .Z(n12905) );
  NAND U12958 ( .A(n12907), .B(n12906), .Z(n12902) );
  XOR U12959 ( .A(n230), .B(n229), .Z(\A1[281] ) );
  XOR U12960 ( .A(n12907), .B(n12908), .Z(n229) );
  XNOR U12961 ( .A(n12906), .B(n12904), .Z(n12908) );
  AND U12962 ( .A(n12909), .B(n12910), .Z(n12904) );
  NANDN U12963 ( .A(n12911), .B(n12912), .Z(n12910) );
  OR U12964 ( .A(n12913), .B(n12914), .Z(n12912) );
  NAND U12965 ( .A(n12914), .B(n12913), .Z(n12909) );
  ANDN U12966 ( .B(B[252]), .A(n54), .Z(n12906) );
  XNOR U12967 ( .A(n12894), .B(n12915), .Z(n12907) );
  XNOR U12968 ( .A(n12893), .B(n12891), .Z(n12915) );
  AND U12969 ( .A(n12916), .B(n12917), .Z(n12891) );
  NANDN U12970 ( .A(n12918), .B(n12919), .Z(n12917) );
  NANDN U12971 ( .A(n12920), .B(n12921), .Z(n12919) );
  NANDN U12972 ( .A(n12921), .B(n12920), .Z(n12916) );
  ANDN U12973 ( .B(B[253]), .A(n55), .Z(n12893) );
  XOR U12974 ( .A(n12899), .B(n12922), .Z(n12894) );
  XOR U12975 ( .A(n12900), .B(n12901), .Z(n12922) );
  NAND U12976 ( .A(A[28]), .B(B[255]), .Z(n12901) );
  AND U12977 ( .A(B[254]), .B(A[29]), .Z(n12900) );
  NAND U12978 ( .A(n12923), .B(n12924), .Z(n12899) );
  NAND U12979 ( .A(n12925), .B(n12926), .Z(n12924) );
  NANDN U12980 ( .A(n12927), .B(n12928), .Z(n12925) );
  NANDN U12981 ( .A(n12928), .B(n12927), .Z(n12923) );
  NAND U12982 ( .A(n12929), .B(n12930), .Z(n230) );
  NANDN U12983 ( .A(n12931), .B(n12932), .Z(n12930) );
  NAND U12984 ( .A(n12934), .B(n12933), .Z(n12929) );
  XOR U12985 ( .A(n232), .B(n231), .Z(\A1[280] ) );
  XOR U12986 ( .A(n12934), .B(n12935), .Z(n231) );
  XNOR U12987 ( .A(n12933), .B(n12931), .Z(n12935) );
  AND U12988 ( .A(n12936), .B(n12937), .Z(n12931) );
  NANDN U12989 ( .A(n12938), .B(n12939), .Z(n12937) );
  NANDN U12990 ( .A(n12940), .B(n12941), .Z(n12939) );
  NANDN U12991 ( .A(n12941), .B(n12940), .Z(n12936) );
  ANDN U12992 ( .B(B[251]), .A(n54), .Z(n12933) );
  XOR U12993 ( .A(n12914), .B(n12942), .Z(n12934) );
  XNOR U12994 ( .A(n12913), .B(n12911), .Z(n12942) );
  AND U12995 ( .A(n12943), .B(n12944), .Z(n12911) );
  NANDN U12996 ( .A(n12945), .B(n12946), .Z(n12944) );
  OR U12997 ( .A(n12947), .B(n12948), .Z(n12946) );
  NAND U12998 ( .A(n12948), .B(n12947), .Z(n12943) );
  ANDN U12999 ( .B(B[252]), .A(n55), .Z(n12913) );
  XNOR U13000 ( .A(n12921), .B(n12949), .Z(n12914) );
  XNOR U13001 ( .A(n12920), .B(n12918), .Z(n12949) );
  AND U13002 ( .A(n12950), .B(n12951), .Z(n12918) );
  NANDN U13003 ( .A(n12952), .B(n12953), .Z(n12951) );
  NANDN U13004 ( .A(n12954), .B(n12955), .Z(n12953) );
  NANDN U13005 ( .A(n12955), .B(n12954), .Z(n12950) );
  ANDN U13006 ( .B(B[253]), .A(n56), .Z(n12920) );
  XOR U13007 ( .A(n12926), .B(n12956), .Z(n12921) );
  XOR U13008 ( .A(n12927), .B(n12928), .Z(n12956) );
  NAND U13009 ( .A(A[27]), .B(B[255]), .Z(n12928) );
  AND U13010 ( .A(B[254]), .B(A[28]), .Z(n12927) );
  NAND U13011 ( .A(n12957), .B(n12958), .Z(n12926) );
  NAND U13012 ( .A(n12959), .B(n12960), .Z(n12958) );
  NANDN U13013 ( .A(n12961), .B(n12962), .Z(n12959) );
  NANDN U13014 ( .A(n12962), .B(n12961), .Z(n12957) );
  NAND U13015 ( .A(n12963), .B(n12964), .Z(n232) );
  NANDN U13016 ( .A(n12965), .B(n12966), .Z(n12964) );
  OR U13017 ( .A(n12967), .B(n12968), .Z(n12966) );
  NAND U13018 ( .A(n12968), .B(n12967), .Z(n12963) );
  XOR U13019 ( .A(n12674), .B(n12969), .Z(\A1[27] ) );
  XNOR U13020 ( .A(n12673), .B(n12671), .Z(n12969) );
  AND U13021 ( .A(n12970), .B(n12971), .Z(n12671) );
  NAND U13022 ( .A(n12972), .B(n12973), .Z(n12971) );
  NANDN U13023 ( .A(n12974), .B(n12975), .Z(n12972) );
  NANDN U13024 ( .A(n12975), .B(n12974), .Z(n12970) );
  ANDN U13025 ( .B(B[0]), .A(n56), .Z(n12673) );
  XNOR U13026 ( .A(n12681), .B(n12976), .Z(n12674) );
  XNOR U13027 ( .A(n12680), .B(n12678), .Z(n12976) );
  AND U13028 ( .A(n12977), .B(n12978), .Z(n12678) );
  NANDN U13029 ( .A(n12979), .B(n12980), .Z(n12978) );
  OR U13030 ( .A(n12981), .B(n12982), .Z(n12980) );
  NAND U13031 ( .A(n12982), .B(n12981), .Z(n12977) );
  ANDN U13032 ( .B(B[1]), .A(n57), .Z(n12680) );
  XNOR U13033 ( .A(n12688), .B(n12983), .Z(n12681) );
  XNOR U13034 ( .A(n12687), .B(n12685), .Z(n12983) );
  AND U13035 ( .A(n12984), .B(n12985), .Z(n12685) );
  NANDN U13036 ( .A(n12986), .B(n12987), .Z(n12985) );
  NANDN U13037 ( .A(n12988), .B(n12989), .Z(n12987) );
  NANDN U13038 ( .A(n12989), .B(n12988), .Z(n12984) );
  ANDN U13039 ( .B(B[2]), .A(n58), .Z(n12687) );
  XNOR U13040 ( .A(n12695), .B(n12990), .Z(n12688) );
  XNOR U13041 ( .A(n12694), .B(n12692), .Z(n12990) );
  AND U13042 ( .A(n12991), .B(n12992), .Z(n12692) );
  NANDN U13043 ( .A(n12993), .B(n12994), .Z(n12992) );
  OR U13044 ( .A(n12995), .B(n12996), .Z(n12994) );
  NAND U13045 ( .A(n12996), .B(n12995), .Z(n12991) );
  ANDN U13046 ( .B(B[3]), .A(n59), .Z(n12694) );
  XNOR U13047 ( .A(n12702), .B(n12997), .Z(n12695) );
  XNOR U13048 ( .A(n12701), .B(n12699), .Z(n12997) );
  AND U13049 ( .A(n12998), .B(n12999), .Z(n12699) );
  NANDN U13050 ( .A(n13000), .B(n13001), .Z(n12999) );
  NANDN U13051 ( .A(n13002), .B(n13003), .Z(n13001) );
  NANDN U13052 ( .A(n13003), .B(n13002), .Z(n12998) );
  ANDN U13053 ( .B(B[4]), .A(n60), .Z(n12701) );
  XNOR U13054 ( .A(n12709), .B(n13004), .Z(n12702) );
  XNOR U13055 ( .A(n12708), .B(n12706), .Z(n13004) );
  AND U13056 ( .A(n13005), .B(n13006), .Z(n12706) );
  NANDN U13057 ( .A(n13007), .B(n13008), .Z(n13006) );
  OR U13058 ( .A(n13009), .B(n13010), .Z(n13008) );
  NAND U13059 ( .A(n13010), .B(n13009), .Z(n13005) );
  ANDN U13060 ( .B(B[5]), .A(n61), .Z(n12708) );
  XNOR U13061 ( .A(n12716), .B(n13011), .Z(n12709) );
  XNOR U13062 ( .A(n12715), .B(n12713), .Z(n13011) );
  AND U13063 ( .A(n13012), .B(n13013), .Z(n12713) );
  NANDN U13064 ( .A(n13014), .B(n13015), .Z(n13013) );
  NANDN U13065 ( .A(n13016), .B(n13017), .Z(n13015) );
  NANDN U13066 ( .A(n13017), .B(n13016), .Z(n13012) );
  ANDN U13067 ( .B(B[6]), .A(n62), .Z(n12715) );
  XNOR U13068 ( .A(n12723), .B(n13018), .Z(n12716) );
  XNOR U13069 ( .A(n12722), .B(n12720), .Z(n13018) );
  AND U13070 ( .A(n13019), .B(n13020), .Z(n12720) );
  NANDN U13071 ( .A(n13021), .B(n13022), .Z(n13020) );
  OR U13072 ( .A(n13023), .B(n13024), .Z(n13022) );
  NAND U13073 ( .A(n13024), .B(n13023), .Z(n13019) );
  ANDN U13074 ( .B(B[7]), .A(n63), .Z(n12722) );
  XNOR U13075 ( .A(n12730), .B(n13025), .Z(n12723) );
  XNOR U13076 ( .A(n12729), .B(n12727), .Z(n13025) );
  AND U13077 ( .A(n13026), .B(n13027), .Z(n12727) );
  NANDN U13078 ( .A(n13028), .B(n13029), .Z(n13027) );
  NANDN U13079 ( .A(n13030), .B(n13031), .Z(n13029) );
  NANDN U13080 ( .A(n13031), .B(n13030), .Z(n13026) );
  ANDN U13081 ( .B(B[8]), .A(n64), .Z(n12729) );
  XNOR U13082 ( .A(n12737), .B(n13032), .Z(n12730) );
  XNOR U13083 ( .A(n12736), .B(n12734), .Z(n13032) );
  AND U13084 ( .A(n13033), .B(n13034), .Z(n12734) );
  NANDN U13085 ( .A(n13035), .B(n13036), .Z(n13034) );
  OR U13086 ( .A(n13037), .B(n13038), .Z(n13036) );
  NAND U13087 ( .A(n13038), .B(n13037), .Z(n13033) );
  ANDN U13088 ( .B(B[9]), .A(n65), .Z(n12736) );
  XNOR U13089 ( .A(n12744), .B(n13039), .Z(n12737) );
  XNOR U13090 ( .A(n12743), .B(n12741), .Z(n13039) );
  AND U13091 ( .A(n13040), .B(n13041), .Z(n12741) );
  NANDN U13092 ( .A(n13042), .B(n13043), .Z(n13041) );
  NANDN U13093 ( .A(n13044), .B(n13045), .Z(n13043) );
  NANDN U13094 ( .A(n13045), .B(n13044), .Z(n13040) );
  ANDN U13095 ( .B(B[10]), .A(n66), .Z(n12743) );
  XNOR U13096 ( .A(n12751), .B(n13046), .Z(n12744) );
  XNOR U13097 ( .A(n12750), .B(n12748), .Z(n13046) );
  AND U13098 ( .A(n13047), .B(n13048), .Z(n12748) );
  NANDN U13099 ( .A(n13049), .B(n13050), .Z(n13048) );
  OR U13100 ( .A(n13051), .B(n13052), .Z(n13050) );
  NAND U13101 ( .A(n13052), .B(n13051), .Z(n13047) );
  ANDN U13102 ( .B(B[11]), .A(n67), .Z(n12750) );
  XNOR U13103 ( .A(n12758), .B(n13053), .Z(n12751) );
  XNOR U13104 ( .A(n12757), .B(n12755), .Z(n13053) );
  AND U13105 ( .A(n13054), .B(n13055), .Z(n12755) );
  NANDN U13106 ( .A(n13056), .B(n13057), .Z(n13055) );
  NANDN U13107 ( .A(n13058), .B(n13059), .Z(n13057) );
  NANDN U13108 ( .A(n13059), .B(n13058), .Z(n13054) );
  ANDN U13109 ( .B(B[12]), .A(n68), .Z(n12757) );
  XNOR U13110 ( .A(n12765), .B(n13060), .Z(n12758) );
  XNOR U13111 ( .A(n12764), .B(n12762), .Z(n13060) );
  AND U13112 ( .A(n13061), .B(n13062), .Z(n12762) );
  NANDN U13113 ( .A(n13063), .B(n13064), .Z(n13062) );
  OR U13114 ( .A(n13065), .B(n13066), .Z(n13064) );
  NAND U13115 ( .A(n13066), .B(n13065), .Z(n13061) );
  ANDN U13116 ( .B(B[13]), .A(n69), .Z(n12764) );
  XNOR U13117 ( .A(n12772), .B(n13067), .Z(n12765) );
  XNOR U13118 ( .A(n12771), .B(n12769), .Z(n13067) );
  AND U13119 ( .A(n13068), .B(n13069), .Z(n12769) );
  NANDN U13120 ( .A(n13070), .B(n13071), .Z(n13069) );
  NANDN U13121 ( .A(n13072), .B(n13073), .Z(n13071) );
  NANDN U13122 ( .A(n13073), .B(n13072), .Z(n13068) );
  ANDN U13123 ( .B(B[14]), .A(n70), .Z(n12771) );
  XNOR U13124 ( .A(n12779), .B(n13074), .Z(n12772) );
  XNOR U13125 ( .A(n12778), .B(n12776), .Z(n13074) );
  AND U13126 ( .A(n13075), .B(n13076), .Z(n12776) );
  NANDN U13127 ( .A(n13077), .B(n13078), .Z(n13076) );
  OR U13128 ( .A(n13079), .B(n13080), .Z(n13078) );
  NAND U13129 ( .A(n13080), .B(n13079), .Z(n13075) );
  ANDN U13130 ( .B(B[15]), .A(n71), .Z(n12778) );
  XNOR U13131 ( .A(n12786), .B(n13081), .Z(n12779) );
  XNOR U13132 ( .A(n12785), .B(n12783), .Z(n13081) );
  AND U13133 ( .A(n13082), .B(n13083), .Z(n12783) );
  NANDN U13134 ( .A(n13084), .B(n13085), .Z(n13083) );
  NANDN U13135 ( .A(n13086), .B(n13087), .Z(n13085) );
  NANDN U13136 ( .A(n13087), .B(n13086), .Z(n13082) );
  ANDN U13137 ( .B(B[16]), .A(n72), .Z(n12785) );
  XNOR U13138 ( .A(n12793), .B(n13088), .Z(n12786) );
  XNOR U13139 ( .A(n12792), .B(n12790), .Z(n13088) );
  AND U13140 ( .A(n13089), .B(n13090), .Z(n12790) );
  NANDN U13141 ( .A(n13091), .B(n13092), .Z(n13090) );
  OR U13142 ( .A(n13093), .B(n13094), .Z(n13092) );
  NAND U13143 ( .A(n13094), .B(n13093), .Z(n13089) );
  ANDN U13144 ( .B(B[17]), .A(n73), .Z(n12792) );
  XNOR U13145 ( .A(n12800), .B(n13095), .Z(n12793) );
  XNOR U13146 ( .A(n12799), .B(n12797), .Z(n13095) );
  AND U13147 ( .A(n13096), .B(n13097), .Z(n12797) );
  NANDN U13148 ( .A(n13098), .B(n13099), .Z(n13097) );
  NANDN U13149 ( .A(n13100), .B(n13101), .Z(n13099) );
  NANDN U13150 ( .A(n13101), .B(n13100), .Z(n13096) );
  ANDN U13151 ( .B(B[18]), .A(n74), .Z(n12799) );
  XNOR U13152 ( .A(n12807), .B(n13102), .Z(n12800) );
  XNOR U13153 ( .A(n12806), .B(n12804), .Z(n13102) );
  AND U13154 ( .A(n13103), .B(n13104), .Z(n12804) );
  NANDN U13155 ( .A(n13105), .B(n13106), .Z(n13104) );
  OR U13156 ( .A(n13107), .B(n13108), .Z(n13106) );
  NAND U13157 ( .A(n13108), .B(n13107), .Z(n13103) );
  ANDN U13158 ( .B(B[19]), .A(n75), .Z(n12806) );
  XNOR U13159 ( .A(n12814), .B(n13109), .Z(n12807) );
  XNOR U13160 ( .A(n12813), .B(n12811), .Z(n13109) );
  AND U13161 ( .A(n13110), .B(n13111), .Z(n12811) );
  NANDN U13162 ( .A(n13112), .B(n13113), .Z(n13111) );
  NANDN U13163 ( .A(n13114), .B(n13115), .Z(n13113) );
  NANDN U13164 ( .A(n13115), .B(n13114), .Z(n13110) );
  ANDN U13165 ( .B(B[20]), .A(n76), .Z(n12813) );
  XNOR U13166 ( .A(n12821), .B(n13116), .Z(n12814) );
  XNOR U13167 ( .A(n12820), .B(n12818), .Z(n13116) );
  AND U13168 ( .A(n13117), .B(n13118), .Z(n12818) );
  NANDN U13169 ( .A(n13119), .B(n13120), .Z(n13118) );
  OR U13170 ( .A(n13121), .B(n13122), .Z(n13120) );
  NAND U13171 ( .A(n13122), .B(n13121), .Z(n13117) );
  ANDN U13172 ( .B(B[21]), .A(n77), .Z(n12820) );
  XNOR U13173 ( .A(n12828), .B(n13123), .Z(n12821) );
  XNOR U13174 ( .A(n12827), .B(n12825), .Z(n13123) );
  AND U13175 ( .A(n13124), .B(n13125), .Z(n12825) );
  NANDN U13176 ( .A(n13126), .B(n13127), .Z(n13125) );
  NANDN U13177 ( .A(n13128), .B(n13129), .Z(n13127) );
  NANDN U13178 ( .A(n13129), .B(n13128), .Z(n13124) );
  ANDN U13179 ( .B(B[22]), .A(n78), .Z(n12827) );
  XNOR U13180 ( .A(n12835), .B(n13130), .Z(n12828) );
  XNOR U13181 ( .A(n12834), .B(n12832), .Z(n13130) );
  AND U13182 ( .A(n13131), .B(n13132), .Z(n12832) );
  NANDN U13183 ( .A(n13133), .B(n13134), .Z(n13132) );
  OR U13184 ( .A(n13135), .B(n13136), .Z(n13134) );
  NAND U13185 ( .A(n13136), .B(n13135), .Z(n13131) );
  ANDN U13186 ( .B(B[23]), .A(n79), .Z(n12834) );
  XNOR U13187 ( .A(n12842), .B(n13137), .Z(n12835) );
  XNOR U13188 ( .A(n12841), .B(n12839), .Z(n13137) );
  AND U13189 ( .A(n13138), .B(n13139), .Z(n12839) );
  NANDN U13190 ( .A(n13140), .B(n13141), .Z(n13139) );
  NANDN U13191 ( .A(n13142), .B(n13143), .Z(n13141) );
  NANDN U13192 ( .A(n13143), .B(n13142), .Z(n13138) );
  ANDN U13193 ( .B(B[24]), .A(n80), .Z(n12841) );
  XNOR U13194 ( .A(n12849), .B(n13144), .Z(n12842) );
  XNOR U13195 ( .A(n12848), .B(n12846), .Z(n13144) );
  AND U13196 ( .A(n13145), .B(n13146), .Z(n12846) );
  NANDN U13197 ( .A(n13147), .B(n13148), .Z(n13146) );
  OR U13198 ( .A(n13149), .B(n13150), .Z(n13148) );
  NAND U13199 ( .A(n13150), .B(n13149), .Z(n13145) );
  ANDN U13200 ( .B(B[25]), .A(n81), .Z(n12848) );
  XNOR U13201 ( .A(n12856), .B(n13151), .Z(n12849) );
  XNOR U13202 ( .A(n12855), .B(n12853), .Z(n13151) );
  AND U13203 ( .A(n13152), .B(n13153), .Z(n12853) );
  NANDN U13204 ( .A(n13154), .B(n13155), .Z(n13153) );
  NAND U13205 ( .A(n13156), .B(n13157), .Z(n13155) );
  ANDN U13206 ( .B(B[26]), .A(n82), .Z(n12855) );
  XOR U13207 ( .A(n12862), .B(n13158), .Z(n12856) );
  XNOR U13208 ( .A(n12860), .B(n12863), .Z(n13158) );
  NAND U13209 ( .A(A[2]), .B(B[27]), .Z(n12863) );
  NANDN U13210 ( .A(n13159), .B(n13160), .Z(n12860) );
  AND U13211 ( .A(A[0]), .B(B[28]), .Z(n13160) );
  XNOR U13212 ( .A(n12865), .B(n13161), .Z(n12862) );
  NAND U13213 ( .A(A[0]), .B(B[29]), .Z(n13161) );
  NAND U13214 ( .A(B[28]), .B(A[1]), .Z(n12865) );
  XOR U13215 ( .A(n234), .B(n233), .Z(\A1[279] ) );
  XOR U13216 ( .A(n12968), .B(n13162), .Z(n233) );
  XNOR U13217 ( .A(n12967), .B(n12965), .Z(n13162) );
  AND U13218 ( .A(n13163), .B(n13164), .Z(n12965) );
  NANDN U13219 ( .A(n13165), .B(n13166), .Z(n13164) );
  OR U13220 ( .A(n13167), .B(n13168), .Z(n13166) );
  NAND U13221 ( .A(n13168), .B(n13167), .Z(n13163) );
  ANDN U13222 ( .B(B[250]), .A(n54), .Z(n12967) );
  XNOR U13223 ( .A(n12941), .B(n13169), .Z(n12968) );
  XNOR U13224 ( .A(n12940), .B(n12938), .Z(n13169) );
  AND U13225 ( .A(n13170), .B(n13171), .Z(n12938) );
  NANDN U13226 ( .A(n13172), .B(n13173), .Z(n13171) );
  NANDN U13227 ( .A(n13174), .B(n13175), .Z(n13173) );
  NANDN U13228 ( .A(n13175), .B(n13174), .Z(n13170) );
  ANDN U13229 ( .B(B[251]), .A(n55), .Z(n12940) );
  XNOR U13230 ( .A(n12948), .B(n13176), .Z(n12941) );
  XNOR U13231 ( .A(n12947), .B(n12945), .Z(n13176) );
  AND U13232 ( .A(n13177), .B(n13178), .Z(n12945) );
  NANDN U13233 ( .A(n13179), .B(n13180), .Z(n13178) );
  OR U13234 ( .A(n13181), .B(n13182), .Z(n13180) );
  NAND U13235 ( .A(n13182), .B(n13181), .Z(n13177) );
  ANDN U13236 ( .B(B[252]), .A(n56), .Z(n12947) );
  XNOR U13237 ( .A(n12955), .B(n13183), .Z(n12948) );
  XNOR U13238 ( .A(n12954), .B(n12952), .Z(n13183) );
  AND U13239 ( .A(n13184), .B(n13185), .Z(n12952) );
  NANDN U13240 ( .A(n13186), .B(n13187), .Z(n13185) );
  NANDN U13241 ( .A(n13188), .B(n13189), .Z(n13187) );
  NANDN U13242 ( .A(n13189), .B(n13188), .Z(n13184) );
  ANDN U13243 ( .B(B[253]), .A(n57), .Z(n12954) );
  XOR U13244 ( .A(n12960), .B(n13190), .Z(n12955) );
  XOR U13245 ( .A(n12961), .B(n12962), .Z(n13190) );
  NAND U13246 ( .A(A[26]), .B(B[255]), .Z(n12962) );
  AND U13247 ( .A(B[254]), .B(A[27]), .Z(n12961) );
  NAND U13248 ( .A(n13191), .B(n13192), .Z(n12960) );
  NAND U13249 ( .A(n13193), .B(n13194), .Z(n13192) );
  NANDN U13250 ( .A(n13195), .B(n13196), .Z(n13193) );
  NANDN U13251 ( .A(n13196), .B(n13195), .Z(n13191) );
  NAND U13252 ( .A(n13197), .B(n13198), .Z(n234) );
  NANDN U13253 ( .A(n13199), .B(n13200), .Z(n13198) );
  NAND U13254 ( .A(n13202), .B(n13201), .Z(n13197) );
  XOR U13255 ( .A(n236), .B(n235), .Z(\A1[278] ) );
  XOR U13256 ( .A(n13202), .B(n13203), .Z(n235) );
  XNOR U13257 ( .A(n13201), .B(n13199), .Z(n13203) );
  AND U13258 ( .A(n13204), .B(n13205), .Z(n13199) );
  NANDN U13259 ( .A(n13206), .B(n13207), .Z(n13205) );
  NANDN U13260 ( .A(n13208), .B(n13209), .Z(n13207) );
  NANDN U13261 ( .A(n13209), .B(n13208), .Z(n13204) );
  ANDN U13262 ( .B(B[249]), .A(n54), .Z(n13201) );
  XOR U13263 ( .A(n13168), .B(n13210), .Z(n13202) );
  XNOR U13264 ( .A(n13167), .B(n13165), .Z(n13210) );
  AND U13265 ( .A(n13211), .B(n13212), .Z(n13165) );
  NANDN U13266 ( .A(n13213), .B(n13214), .Z(n13212) );
  OR U13267 ( .A(n13215), .B(n13216), .Z(n13214) );
  NAND U13268 ( .A(n13216), .B(n13215), .Z(n13211) );
  ANDN U13269 ( .B(B[250]), .A(n55), .Z(n13167) );
  XNOR U13270 ( .A(n13175), .B(n13217), .Z(n13168) );
  XNOR U13271 ( .A(n13174), .B(n13172), .Z(n13217) );
  AND U13272 ( .A(n13218), .B(n13219), .Z(n13172) );
  NANDN U13273 ( .A(n13220), .B(n13221), .Z(n13219) );
  NANDN U13274 ( .A(n13222), .B(n13223), .Z(n13221) );
  NANDN U13275 ( .A(n13223), .B(n13222), .Z(n13218) );
  ANDN U13276 ( .B(B[251]), .A(n56), .Z(n13174) );
  XNOR U13277 ( .A(n13182), .B(n13224), .Z(n13175) );
  XNOR U13278 ( .A(n13181), .B(n13179), .Z(n13224) );
  AND U13279 ( .A(n13225), .B(n13226), .Z(n13179) );
  NANDN U13280 ( .A(n13227), .B(n13228), .Z(n13226) );
  OR U13281 ( .A(n13229), .B(n13230), .Z(n13228) );
  NAND U13282 ( .A(n13230), .B(n13229), .Z(n13225) );
  ANDN U13283 ( .B(B[252]), .A(n57), .Z(n13181) );
  XNOR U13284 ( .A(n13189), .B(n13231), .Z(n13182) );
  XNOR U13285 ( .A(n13188), .B(n13186), .Z(n13231) );
  AND U13286 ( .A(n13232), .B(n13233), .Z(n13186) );
  NANDN U13287 ( .A(n13234), .B(n13235), .Z(n13233) );
  NANDN U13288 ( .A(n13236), .B(n13237), .Z(n13235) );
  NANDN U13289 ( .A(n13237), .B(n13236), .Z(n13232) );
  ANDN U13290 ( .B(B[253]), .A(n58), .Z(n13188) );
  XOR U13291 ( .A(n13194), .B(n13238), .Z(n13189) );
  XOR U13292 ( .A(n13195), .B(n13196), .Z(n13238) );
  NAND U13293 ( .A(A[25]), .B(B[255]), .Z(n13196) );
  AND U13294 ( .A(B[254]), .B(A[26]), .Z(n13195) );
  NAND U13295 ( .A(n13239), .B(n13240), .Z(n13194) );
  NAND U13296 ( .A(n13241), .B(n13242), .Z(n13240) );
  NANDN U13297 ( .A(n13243), .B(n13244), .Z(n13241) );
  NANDN U13298 ( .A(n13244), .B(n13243), .Z(n13239) );
  NAND U13299 ( .A(n13245), .B(n13246), .Z(n236) );
  NANDN U13300 ( .A(n13247), .B(n13248), .Z(n13246) );
  OR U13301 ( .A(n13249), .B(n13250), .Z(n13248) );
  NAND U13302 ( .A(n13250), .B(n13249), .Z(n13245) );
  XOR U13303 ( .A(n238), .B(n237), .Z(\A1[277] ) );
  XOR U13304 ( .A(n13250), .B(n13251), .Z(n237) );
  XNOR U13305 ( .A(n13249), .B(n13247), .Z(n13251) );
  AND U13306 ( .A(n13252), .B(n13253), .Z(n13247) );
  NANDN U13307 ( .A(n13254), .B(n13255), .Z(n13253) );
  OR U13308 ( .A(n13256), .B(n13257), .Z(n13255) );
  NAND U13309 ( .A(n13257), .B(n13256), .Z(n13252) );
  ANDN U13310 ( .B(B[248]), .A(n54), .Z(n13249) );
  XNOR U13311 ( .A(n13209), .B(n13258), .Z(n13250) );
  XNOR U13312 ( .A(n13208), .B(n13206), .Z(n13258) );
  AND U13313 ( .A(n13259), .B(n13260), .Z(n13206) );
  NANDN U13314 ( .A(n13261), .B(n13262), .Z(n13260) );
  NANDN U13315 ( .A(n13263), .B(n13264), .Z(n13262) );
  NANDN U13316 ( .A(n13264), .B(n13263), .Z(n13259) );
  ANDN U13317 ( .B(B[249]), .A(n55), .Z(n13208) );
  XNOR U13318 ( .A(n13216), .B(n13265), .Z(n13209) );
  XNOR U13319 ( .A(n13215), .B(n13213), .Z(n13265) );
  AND U13320 ( .A(n13266), .B(n13267), .Z(n13213) );
  NANDN U13321 ( .A(n13268), .B(n13269), .Z(n13267) );
  OR U13322 ( .A(n13270), .B(n13271), .Z(n13269) );
  NAND U13323 ( .A(n13271), .B(n13270), .Z(n13266) );
  ANDN U13324 ( .B(B[250]), .A(n56), .Z(n13215) );
  XNOR U13325 ( .A(n13223), .B(n13272), .Z(n13216) );
  XNOR U13326 ( .A(n13222), .B(n13220), .Z(n13272) );
  AND U13327 ( .A(n13273), .B(n13274), .Z(n13220) );
  NANDN U13328 ( .A(n13275), .B(n13276), .Z(n13274) );
  NANDN U13329 ( .A(n13277), .B(n13278), .Z(n13276) );
  NANDN U13330 ( .A(n13278), .B(n13277), .Z(n13273) );
  ANDN U13331 ( .B(B[251]), .A(n57), .Z(n13222) );
  XNOR U13332 ( .A(n13230), .B(n13279), .Z(n13223) );
  XNOR U13333 ( .A(n13229), .B(n13227), .Z(n13279) );
  AND U13334 ( .A(n13280), .B(n13281), .Z(n13227) );
  NANDN U13335 ( .A(n13282), .B(n13283), .Z(n13281) );
  OR U13336 ( .A(n13284), .B(n13285), .Z(n13283) );
  NAND U13337 ( .A(n13285), .B(n13284), .Z(n13280) );
  ANDN U13338 ( .B(B[252]), .A(n58), .Z(n13229) );
  XNOR U13339 ( .A(n13237), .B(n13286), .Z(n13230) );
  XNOR U13340 ( .A(n13236), .B(n13234), .Z(n13286) );
  AND U13341 ( .A(n13287), .B(n13288), .Z(n13234) );
  NANDN U13342 ( .A(n13289), .B(n13290), .Z(n13288) );
  NANDN U13343 ( .A(n13291), .B(n13292), .Z(n13290) );
  NANDN U13344 ( .A(n13292), .B(n13291), .Z(n13287) );
  ANDN U13345 ( .B(B[253]), .A(n59), .Z(n13236) );
  XOR U13346 ( .A(n13242), .B(n13293), .Z(n13237) );
  XOR U13347 ( .A(n13243), .B(n13244), .Z(n13293) );
  NAND U13348 ( .A(A[24]), .B(B[255]), .Z(n13244) );
  AND U13349 ( .A(B[254]), .B(A[25]), .Z(n13243) );
  NAND U13350 ( .A(n13294), .B(n13295), .Z(n13242) );
  NAND U13351 ( .A(n13296), .B(n13297), .Z(n13295) );
  NANDN U13352 ( .A(n13298), .B(n13299), .Z(n13296) );
  NANDN U13353 ( .A(n13299), .B(n13298), .Z(n13294) );
  NAND U13354 ( .A(n13300), .B(n13301), .Z(n238) );
  NANDN U13355 ( .A(n13302), .B(n13303), .Z(n13301) );
  NAND U13356 ( .A(n13305), .B(n13304), .Z(n13300) );
  XOR U13357 ( .A(n240), .B(n239), .Z(\A1[276] ) );
  XOR U13358 ( .A(n13305), .B(n13306), .Z(n239) );
  XNOR U13359 ( .A(n13304), .B(n13302), .Z(n13306) );
  AND U13360 ( .A(n13307), .B(n13308), .Z(n13302) );
  NANDN U13361 ( .A(n13309), .B(n13310), .Z(n13308) );
  NANDN U13362 ( .A(n13311), .B(n13312), .Z(n13310) );
  NANDN U13363 ( .A(n13312), .B(n13311), .Z(n13307) );
  ANDN U13364 ( .B(B[247]), .A(n54), .Z(n13304) );
  XOR U13365 ( .A(n13257), .B(n13313), .Z(n13305) );
  XNOR U13366 ( .A(n13256), .B(n13254), .Z(n13313) );
  AND U13367 ( .A(n13314), .B(n13315), .Z(n13254) );
  NANDN U13368 ( .A(n13316), .B(n13317), .Z(n13315) );
  OR U13369 ( .A(n13318), .B(n13319), .Z(n13317) );
  NAND U13370 ( .A(n13319), .B(n13318), .Z(n13314) );
  ANDN U13371 ( .B(B[248]), .A(n55), .Z(n13256) );
  XNOR U13372 ( .A(n13264), .B(n13320), .Z(n13257) );
  XNOR U13373 ( .A(n13263), .B(n13261), .Z(n13320) );
  AND U13374 ( .A(n13321), .B(n13322), .Z(n13261) );
  NANDN U13375 ( .A(n13323), .B(n13324), .Z(n13322) );
  NANDN U13376 ( .A(n13325), .B(n13326), .Z(n13324) );
  NANDN U13377 ( .A(n13326), .B(n13325), .Z(n13321) );
  ANDN U13378 ( .B(B[249]), .A(n56), .Z(n13263) );
  XNOR U13379 ( .A(n13271), .B(n13327), .Z(n13264) );
  XNOR U13380 ( .A(n13270), .B(n13268), .Z(n13327) );
  AND U13381 ( .A(n13328), .B(n13329), .Z(n13268) );
  NANDN U13382 ( .A(n13330), .B(n13331), .Z(n13329) );
  OR U13383 ( .A(n13332), .B(n13333), .Z(n13331) );
  NAND U13384 ( .A(n13333), .B(n13332), .Z(n13328) );
  ANDN U13385 ( .B(B[250]), .A(n57), .Z(n13270) );
  XNOR U13386 ( .A(n13278), .B(n13334), .Z(n13271) );
  XNOR U13387 ( .A(n13277), .B(n13275), .Z(n13334) );
  AND U13388 ( .A(n13335), .B(n13336), .Z(n13275) );
  NANDN U13389 ( .A(n13337), .B(n13338), .Z(n13336) );
  NANDN U13390 ( .A(n13339), .B(n13340), .Z(n13338) );
  NANDN U13391 ( .A(n13340), .B(n13339), .Z(n13335) );
  ANDN U13392 ( .B(B[251]), .A(n58), .Z(n13277) );
  XNOR U13393 ( .A(n13285), .B(n13341), .Z(n13278) );
  XNOR U13394 ( .A(n13284), .B(n13282), .Z(n13341) );
  AND U13395 ( .A(n13342), .B(n13343), .Z(n13282) );
  NANDN U13396 ( .A(n13344), .B(n13345), .Z(n13343) );
  OR U13397 ( .A(n13346), .B(n13347), .Z(n13345) );
  NAND U13398 ( .A(n13347), .B(n13346), .Z(n13342) );
  ANDN U13399 ( .B(B[252]), .A(n59), .Z(n13284) );
  XNOR U13400 ( .A(n13292), .B(n13348), .Z(n13285) );
  XNOR U13401 ( .A(n13291), .B(n13289), .Z(n13348) );
  AND U13402 ( .A(n13349), .B(n13350), .Z(n13289) );
  NANDN U13403 ( .A(n13351), .B(n13352), .Z(n13350) );
  NANDN U13404 ( .A(n13353), .B(n13354), .Z(n13352) );
  NANDN U13405 ( .A(n13354), .B(n13353), .Z(n13349) );
  ANDN U13406 ( .B(B[253]), .A(n60), .Z(n13291) );
  XOR U13407 ( .A(n13297), .B(n13355), .Z(n13292) );
  XOR U13408 ( .A(n13298), .B(n13299), .Z(n13355) );
  NAND U13409 ( .A(A[23]), .B(B[255]), .Z(n13299) );
  AND U13410 ( .A(B[254]), .B(A[24]), .Z(n13298) );
  NAND U13411 ( .A(n13356), .B(n13357), .Z(n13297) );
  NAND U13412 ( .A(n13358), .B(n13359), .Z(n13357) );
  NANDN U13413 ( .A(n13360), .B(n13361), .Z(n13358) );
  NANDN U13414 ( .A(n13361), .B(n13360), .Z(n13356) );
  NAND U13415 ( .A(n13362), .B(n13363), .Z(n240) );
  NANDN U13416 ( .A(n13364), .B(n13365), .Z(n13363) );
  OR U13417 ( .A(n13366), .B(n13367), .Z(n13365) );
  NAND U13418 ( .A(n13367), .B(n13366), .Z(n13362) );
  XOR U13419 ( .A(n242), .B(n241), .Z(\A1[275] ) );
  XOR U13420 ( .A(n13367), .B(n13368), .Z(n241) );
  XNOR U13421 ( .A(n13366), .B(n13364), .Z(n13368) );
  AND U13422 ( .A(n13369), .B(n13370), .Z(n13364) );
  NANDN U13423 ( .A(n13371), .B(n13372), .Z(n13370) );
  OR U13424 ( .A(n13373), .B(n13374), .Z(n13372) );
  NAND U13425 ( .A(n13374), .B(n13373), .Z(n13369) );
  ANDN U13426 ( .B(B[246]), .A(n54), .Z(n13366) );
  XNOR U13427 ( .A(n13312), .B(n13375), .Z(n13367) );
  XNOR U13428 ( .A(n13311), .B(n13309), .Z(n13375) );
  AND U13429 ( .A(n13376), .B(n13377), .Z(n13309) );
  NANDN U13430 ( .A(n13378), .B(n13379), .Z(n13377) );
  NANDN U13431 ( .A(n13380), .B(n13381), .Z(n13379) );
  NANDN U13432 ( .A(n13381), .B(n13380), .Z(n13376) );
  ANDN U13433 ( .B(B[247]), .A(n55), .Z(n13311) );
  XNOR U13434 ( .A(n13319), .B(n13382), .Z(n13312) );
  XNOR U13435 ( .A(n13318), .B(n13316), .Z(n13382) );
  AND U13436 ( .A(n13383), .B(n13384), .Z(n13316) );
  NANDN U13437 ( .A(n13385), .B(n13386), .Z(n13384) );
  OR U13438 ( .A(n13387), .B(n13388), .Z(n13386) );
  NAND U13439 ( .A(n13388), .B(n13387), .Z(n13383) );
  ANDN U13440 ( .B(B[248]), .A(n56), .Z(n13318) );
  XNOR U13441 ( .A(n13326), .B(n13389), .Z(n13319) );
  XNOR U13442 ( .A(n13325), .B(n13323), .Z(n13389) );
  AND U13443 ( .A(n13390), .B(n13391), .Z(n13323) );
  NANDN U13444 ( .A(n13392), .B(n13393), .Z(n13391) );
  NANDN U13445 ( .A(n13394), .B(n13395), .Z(n13393) );
  NANDN U13446 ( .A(n13395), .B(n13394), .Z(n13390) );
  ANDN U13447 ( .B(B[249]), .A(n57), .Z(n13325) );
  XNOR U13448 ( .A(n13333), .B(n13396), .Z(n13326) );
  XNOR U13449 ( .A(n13332), .B(n13330), .Z(n13396) );
  AND U13450 ( .A(n13397), .B(n13398), .Z(n13330) );
  NANDN U13451 ( .A(n13399), .B(n13400), .Z(n13398) );
  OR U13452 ( .A(n13401), .B(n13402), .Z(n13400) );
  NAND U13453 ( .A(n13402), .B(n13401), .Z(n13397) );
  ANDN U13454 ( .B(B[250]), .A(n58), .Z(n13332) );
  XNOR U13455 ( .A(n13340), .B(n13403), .Z(n13333) );
  XNOR U13456 ( .A(n13339), .B(n13337), .Z(n13403) );
  AND U13457 ( .A(n13404), .B(n13405), .Z(n13337) );
  NANDN U13458 ( .A(n13406), .B(n13407), .Z(n13405) );
  NANDN U13459 ( .A(n13408), .B(n13409), .Z(n13407) );
  NANDN U13460 ( .A(n13409), .B(n13408), .Z(n13404) );
  ANDN U13461 ( .B(B[251]), .A(n59), .Z(n13339) );
  XNOR U13462 ( .A(n13347), .B(n13410), .Z(n13340) );
  XNOR U13463 ( .A(n13346), .B(n13344), .Z(n13410) );
  AND U13464 ( .A(n13411), .B(n13412), .Z(n13344) );
  NANDN U13465 ( .A(n13413), .B(n13414), .Z(n13412) );
  OR U13466 ( .A(n13415), .B(n13416), .Z(n13414) );
  NAND U13467 ( .A(n13416), .B(n13415), .Z(n13411) );
  ANDN U13468 ( .B(B[252]), .A(n60), .Z(n13346) );
  XNOR U13469 ( .A(n13354), .B(n13417), .Z(n13347) );
  XNOR U13470 ( .A(n13353), .B(n13351), .Z(n13417) );
  AND U13471 ( .A(n13418), .B(n13419), .Z(n13351) );
  NANDN U13472 ( .A(n13420), .B(n13421), .Z(n13419) );
  NANDN U13473 ( .A(n13422), .B(n13423), .Z(n13421) );
  NANDN U13474 ( .A(n13423), .B(n13422), .Z(n13418) );
  ANDN U13475 ( .B(B[253]), .A(n61), .Z(n13353) );
  XOR U13476 ( .A(n13359), .B(n13424), .Z(n13354) );
  XOR U13477 ( .A(n13360), .B(n13361), .Z(n13424) );
  NAND U13478 ( .A(A[22]), .B(B[255]), .Z(n13361) );
  AND U13479 ( .A(B[254]), .B(A[23]), .Z(n13360) );
  NAND U13480 ( .A(n13425), .B(n13426), .Z(n13359) );
  NAND U13481 ( .A(n13427), .B(n13428), .Z(n13426) );
  NANDN U13482 ( .A(n13429), .B(n13430), .Z(n13427) );
  NANDN U13483 ( .A(n13430), .B(n13429), .Z(n13425) );
  NAND U13484 ( .A(n13431), .B(n13432), .Z(n242) );
  NANDN U13485 ( .A(n13433), .B(n13434), .Z(n13432) );
  NAND U13486 ( .A(n13436), .B(n13435), .Z(n13431) );
  XOR U13487 ( .A(n244), .B(n243), .Z(\A1[274] ) );
  XOR U13488 ( .A(n13436), .B(n13437), .Z(n243) );
  XNOR U13489 ( .A(n13435), .B(n13433), .Z(n13437) );
  AND U13490 ( .A(n13438), .B(n13439), .Z(n13433) );
  NANDN U13491 ( .A(n13440), .B(n13441), .Z(n13439) );
  NANDN U13492 ( .A(n13442), .B(n13443), .Z(n13441) );
  NANDN U13493 ( .A(n13443), .B(n13442), .Z(n13438) );
  ANDN U13494 ( .B(B[245]), .A(n54), .Z(n13435) );
  XOR U13495 ( .A(n13374), .B(n13444), .Z(n13436) );
  XNOR U13496 ( .A(n13373), .B(n13371), .Z(n13444) );
  AND U13497 ( .A(n13445), .B(n13446), .Z(n13371) );
  NANDN U13498 ( .A(n13447), .B(n13448), .Z(n13446) );
  OR U13499 ( .A(n13449), .B(n13450), .Z(n13448) );
  NAND U13500 ( .A(n13450), .B(n13449), .Z(n13445) );
  ANDN U13501 ( .B(B[246]), .A(n55), .Z(n13373) );
  XNOR U13502 ( .A(n13381), .B(n13451), .Z(n13374) );
  XNOR U13503 ( .A(n13380), .B(n13378), .Z(n13451) );
  AND U13504 ( .A(n13452), .B(n13453), .Z(n13378) );
  NANDN U13505 ( .A(n13454), .B(n13455), .Z(n13453) );
  NANDN U13506 ( .A(n13456), .B(n13457), .Z(n13455) );
  NANDN U13507 ( .A(n13457), .B(n13456), .Z(n13452) );
  ANDN U13508 ( .B(B[247]), .A(n56), .Z(n13380) );
  XNOR U13509 ( .A(n13388), .B(n13458), .Z(n13381) );
  XNOR U13510 ( .A(n13387), .B(n13385), .Z(n13458) );
  AND U13511 ( .A(n13459), .B(n13460), .Z(n13385) );
  NANDN U13512 ( .A(n13461), .B(n13462), .Z(n13460) );
  OR U13513 ( .A(n13463), .B(n13464), .Z(n13462) );
  NAND U13514 ( .A(n13464), .B(n13463), .Z(n13459) );
  ANDN U13515 ( .B(B[248]), .A(n57), .Z(n13387) );
  XNOR U13516 ( .A(n13395), .B(n13465), .Z(n13388) );
  XNOR U13517 ( .A(n13394), .B(n13392), .Z(n13465) );
  AND U13518 ( .A(n13466), .B(n13467), .Z(n13392) );
  NANDN U13519 ( .A(n13468), .B(n13469), .Z(n13467) );
  NANDN U13520 ( .A(n13470), .B(n13471), .Z(n13469) );
  NANDN U13521 ( .A(n13471), .B(n13470), .Z(n13466) );
  ANDN U13522 ( .B(B[249]), .A(n58), .Z(n13394) );
  XNOR U13523 ( .A(n13402), .B(n13472), .Z(n13395) );
  XNOR U13524 ( .A(n13401), .B(n13399), .Z(n13472) );
  AND U13525 ( .A(n13473), .B(n13474), .Z(n13399) );
  NANDN U13526 ( .A(n13475), .B(n13476), .Z(n13474) );
  OR U13527 ( .A(n13477), .B(n13478), .Z(n13476) );
  NAND U13528 ( .A(n13478), .B(n13477), .Z(n13473) );
  ANDN U13529 ( .B(B[250]), .A(n59), .Z(n13401) );
  XNOR U13530 ( .A(n13409), .B(n13479), .Z(n13402) );
  XNOR U13531 ( .A(n13408), .B(n13406), .Z(n13479) );
  AND U13532 ( .A(n13480), .B(n13481), .Z(n13406) );
  NANDN U13533 ( .A(n13482), .B(n13483), .Z(n13481) );
  NANDN U13534 ( .A(n13484), .B(n13485), .Z(n13483) );
  NANDN U13535 ( .A(n13485), .B(n13484), .Z(n13480) );
  ANDN U13536 ( .B(B[251]), .A(n60), .Z(n13408) );
  XNOR U13537 ( .A(n13416), .B(n13486), .Z(n13409) );
  XNOR U13538 ( .A(n13415), .B(n13413), .Z(n13486) );
  AND U13539 ( .A(n13487), .B(n13488), .Z(n13413) );
  NANDN U13540 ( .A(n13489), .B(n13490), .Z(n13488) );
  OR U13541 ( .A(n13491), .B(n13492), .Z(n13490) );
  NAND U13542 ( .A(n13492), .B(n13491), .Z(n13487) );
  ANDN U13543 ( .B(B[252]), .A(n61), .Z(n13415) );
  XNOR U13544 ( .A(n13423), .B(n13493), .Z(n13416) );
  XNOR U13545 ( .A(n13422), .B(n13420), .Z(n13493) );
  AND U13546 ( .A(n13494), .B(n13495), .Z(n13420) );
  NANDN U13547 ( .A(n13496), .B(n13497), .Z(n13495) );
  NANDN U13548 ( .A(n13498), .B(n13499), .Z(n13497) );
  NANDN U13549 ( .A(n13499), .B(n13498), .Z(n13494) );
  ANDN U13550 ( .B(B[253]), .A(n62), .Z(n13422) );
  XOR U13551 ( .A(n13428), .B(n13500), .Z(n13423) );
  XOR U13552 ( .A(n13429), .B(n13430), .Z(n13500) );
  NAND U13553 ( .A(A[21]), .B(B[255]), .Z(n13430) );
  AND U13554 ( .A(B[254]), .B(A[22]), .Z(n13429) );
  NAND U13555 ( .A(n13501), .B(n13502), .Z(n13428) );
  NAND U13556 ( .A(n13503), .B(n13504), .Z(n13502) );
  NANDN U13557 ( .A(n13505), .B(n13506), .Z(n13503) );
  NANDN U13558 ( .A(n13506), .B(n13505), .Z(n13501) );
  NAND U13559 ( .A(n13507), .B(n13508), .Z(n244) );
  NANDN U13560 ( .A(n13509), .B(n13510), .Z(n13508) );
  OR U13561 ( .A(n13511), .B(n13512), .Z(n13510) );
  NAND U13562 ( .A(n13512), .B(n13511), .Z(n13507) );
  XOR U13563 ( .A(n246), .B(n245), .Z(\A1[273] ) );
  XOR U13564 ( .A(n13512), .B(n13513), .Z(n245) );
  XNOR U13565 ( .A(n13511), .B(n13509), .Z(n13513) );
  AND U13566 ( .A(n13514), .B(n13515), .Z(n13509) );
  NANDN U13567 ( .A(n13516), .B(n13517), .Z(n13515) );
  OR U13568 ( .A(n13518), .B(n13519), .Z(n13517) );
  NAND U13569 ( .A(n13519), .B(n13518), .Z(n13514) );
  ANDN U13570 ( .B(B[244]), .A(n54), .Z(n13511) );
  XNOR U13571 ( .A(n13443), .B(n13520), .Z(n13512) );
  XNOR U13572 ( .A(n13442), .B(n13440), .Z(n13520) );
  AND U13573 ( .A(n13521), .B(n13522), .Z(n13440) );
  NANDN U13574 ( .A(n13523), .B(n13524), .Z(n13522) );
  NANDN U13575 ( .A(n13525), .B(n13526), .Z(n13524) );
  NANDN U13576 ( .A(n13526), .B(n13525), .Z(n13521) );
  ANDN U13577 ( .B(B[245]), .A(n55), .Z(n13442) );
  XNOR U13578 ( .A(n13450), .B(n13527), .Z(n13443) );
  XNOR U13579 ( .A(n13449), .B(n13447), .Z(n13527) );
  AND U13580 ( .A(n13528), .B(n13529), .Z(n13447) );
  NANDN U13581 ( .A(n13530), .B(n13531), .Z(n13529) );
  OR U13582 ( .A(n13532), .B(n13533), .Z(n13531) );
  NAND U13583 ( .A(n13533), .B(n13532), .Z(n13528) );
  ANDN U13584 ( .B(B[246]), .A(n56), .Z(n13449) );
  XNOR U13585 ( .A(n13457), .B(n13534), .Z(n13450) );
  XNOR U13586 ( .A(n13456), .B(n13454), .Z(n13534) );
  AND U13587 ( .A(n13535), .B(n13536), .Z(n13454) );
  NANDN U13588 ( .A(n13537), .B(n13538), .Z(n13536) );
  NANDN U13589 ( .A(n13539), .B(n13540), .Z(n13538) );
  NANDN U13590 ( .A(n13540), .B(n13539), .Z(n13535) );
  ANDN U13591 ( .B(B[247]), .A(n57), .Z(n13456) );
  XNOR U13592 ( .A(n13464), .B(n13541), .Z(n13457) );
  XNOR U13593 ( .A(n13463), .B(n13461), .Z(n13541) );
  AND U13594 ( .A(n13542), .B(n13543), .Z(n13461) );
  NANDN U13595 ( .A(n13544), .B(n13545), .Z(n13543) );
  OR U13596 ( .A(n13546), .B(n13547), .Z(n13545) );
  NAND U13597 ( .A(n13547), .B(n13546), .Z(n13542) );
  ANDN U13598 ( .B(B[248]), .A(n58), .Z(n13463) );
  XNOR U13599 ( .A(n13471), .B(n13548), .Z(n13464) );
  XNOR U13600 ( .A(n13470), .B(n13468), .Z(n13548) );
  AND U13601 ( .A(n13549), .B(n13550), .Z(n13468) );
  NANDN U13602 ( .A(n13551), .B(n13552), .Z(n13550) );
  NANDN U13603 ( .A(n13553), .B(n13554), .Z(n13552) );
  NANDN U13604 ( .A(n13554), .B(n13553), .Z(n13549) );
  ANDN U13605 ( .B(B[249]), .A(n59), .Z(n13470) );
  XNOR U13606 ( .A(n13478), .B(n13555), .Z(n13471) );
  XNOR U13607 ( .A(n13477), .B(n13475), .Z(n13555) );
  AND U13608 ( .A(n13556), .B(n13557), .Z(n13475) );
  NANDN U13609 ( .A(n13558), .B(n13559), .Z(n13557) );
  OR U13610 ( .A(n13560), .B(n13561), .Z(n13559) );
  NAND U13611 ( .A(n13561), .B(n13560), .Z(n13556) );
  ANDN U13612 ( .B(B[250]), .A(n60), .Z(n13477) );
  XNOR U13613 ( .A(n13485), .B(n13562), .Z(n13478) );
  XNOR U13614 ( .A(n13484), .B(n13482), .Z(n13562) );
  AND U13615 ( .A(n13563), .B(n13564), .Z(n13482) );
  NANDN U13616 ( .A(n13565), .B(n13566), .Z(n13564) );
  NANDN U13617 ( .A(n13567), .B(n13568), .Z(n13566) );
  NANDN U13618 ( .A(n13568), .B(n13567), .Z(n13563) );
  ANDN U13619 ( .B(B[251]), .A(n61), .Z(n13484) );
  XNOR U13620 ( .A(n13492), .B(n13569), .Z(n13485) );
  XNOR U13621 ( .A(n13491), .B(n13489), .Z(n13569) );
  AND U13622 ( .A(n13570), .B(n13571), .Z(n13489) );
  NANDN U13623 ( .A(n13572), .B(n13573), .Z(n13571) );
  OR U13624 ( .A(n13574), .B(n13575), .Z(n13573) );
  NAND U13625 ( .A(n13575), .B(n13574), .Z(n13570) );
  ANDN U13626 ( .B(B[252]), .A(n62), .Z(n13491) );
  XNOR U13627 ( .A(n13499), .B(n13576), .Z(n13492) );
  XNOR U13628 ( .A(n13498), .B(n13496), .Z(n13576) );
  AND U13629 ( .A(n13577), .B(n13578), .Z(n13496) );
  NANDN U13630 ( .A(n13579), .B(n13580), .Z(n13578) );
  NANDN U13631 ( .A(n13581), .B(n13582), .Z(n13580) );
  NANDN U13632 ( .A(n13582), .B(n13581), .Z(n13577) );
  ANDN U13633 ( .B(B[253]), .A(n63), .Z(n13498) );
  XOR U13634 ( .A(n13504), .B(n13583), .Z(n13499) );
  XOR U13635 ( .A(n13505), .B(n13506), .Z(n13583) );
  NAND U13636 ( .A(A[20]), .B(B[255]), .Z(n13506) );
  AND U13637 ( .A(B[254]), .B(A[21]), .Z(n13505) );
  NAND U13638 ( .A(n13584), .B(n13585), .Z(n13504) );
  NAND U13639 ( .A(n13586), .B(n13587), .Z(n13585) );
  NANDN U13640 ( .A(n13588), .B(n13589), .Z(n13586) );
  NANDN U13641 ( .A(n13589), .B(n13588), .Z(n13584) );
  NAND U13642 ( .A(n13590), .B(n13591), .Z(n246) );
  NANDN U13643 ( .A(n13592), .B(n13593), .Z(n13591) );
  NAND U13644 ( .A(n13595), .B(n13594), .Z(n13590) );
  XOR U13645 ( .A(n248), .B(n247), .Z(\A1[272] ) );
  XOR U13646 ( .A(n13595), .B(n13596), .Z(n247) );
  XNOR U13647 ( .A(n13594), .B(n13592), .Z(n13596) );
  AND U13648 ( .A(n13597), .B(n13598), .Z(n13592) );
  NANDN U13649 ( .A(n13599), .B(n13600), .Z(n13598) );
  NANDN U13650 ( .A(n13601), .B(n13602), .Z(n13600) );
  NANDN U13651 ( .A(n13602), .B(n13601), .Z(n13597) );
  ANDN U13652 ( .B(B[243]), .A(n54), .Z(n13594) );
  XOR U13653 ( .A(n13519), .B(n13603), .Z(n13595) );
  XNOR U13654 ( .A(n13518), .B(n13516), .Z(n13603) );
  AND U13655 ( .A(n13604), .B(n13605), .Z(n13516) );
  NANDN U13656 ( .A(n13606), .B(n13607), .Z(n13605) );
  OR U13657 ( .A(n13608), .B(n13609), .Z(n13607) );
  NAND U13658 ( .A(n13609), .B(n13608), .Z(n13604) );
  ANDN U13659 ( .B(B[244]), .A(n55), .Z(n13518) );
  XNOR U13660 ( .A(n13526), .B(n13610), .Z(n13519) );
  XNOR U13661 ( .A(n13525), .B(n13523), .Z(n13610) );
  AND U13662 ( .A(n13611), .B(n13612), .Z(n13523) );
  NANDN U13663 ( .A(n13613), .B(n13614), .Z(n13612) );
  NANDN U13664 ( .A(n13615), .B(n13616), .Z(n13614) );
  NANDN U13665 ( .A(n13616), .B(n13615), .Z(n13611) );
  ANDN U13666 ( .B(B[245]), .A(n56), .Z(n13525) );
  XNOR U13667 ( .A(n13533), .B(n13617), .Z(n13526) );
  XNOR U13668 ( .A(n13532), .B(n13530), .Z(n13617) );
  AND U13669 ( .A(n13618), .B(n13619), .Z(n13530) );
  NANDN U13670 ( .A(n13620), .B(n13621), .Z(n13619) );
  OR U13671 ( .A(n13622), .B(n13623), .Z(n13621) );
  NAND U13672 ( .A(n13623), .B(n13622), .Z(n13618) );
  ANDN U13673 ( .B(B[246]), .A(n57), .Z(n13532) );
  XNOR U13674 ( .A(n13540), .B(n13624), .Z(n13533) );
  XNOR U13675 ( .A(n13539), .B(n13537), .Z(n13624) );
  AND U13676 ( .A(n13625), .B(n13626), .Z(n13537) );
  NANDN U13677 ( .A(n13627), .B(n13628), .Z(n13626) );
  NANDN U13678 ( .A(n13629), .B(n13630), .Z(n13628) );
  NANDN U13679 ( .A(n13630), .B(n13629), .Z(n13625) );
  ANDN U13680 ( .B(B[247]), .A(n58), .Z(n13539) );
  XNOR U13681 ( .A(n13547), .B(n13631), .Z(n13540) );
  XNOR U13682 ( .A(n13546), .B(n13544), .Z(n13631) );
  AND U13683 ( .A(n13632), .B(n13633), .Z(n13544) );
  NANDN U13684 ( .A(n13634), .B(n13635), .Z(n13633) );
  OR U13685 ( .A(n13636), .B(n13637), .Z(n13635) );
  NAND U13686 ( .A(n13637), .B(n13636), .Z(n13632) );
  ANDN U13687 ( .B(B[248]), .A(n59), .Z(n13546) );
  XNOR U13688 ( .A(n13554), .B(n13638), .Z(n13547) );
  XNOR U13689 ( .A(n13553), .B(n13551), .Z(n13638) );
  AND U13690 ( .A(n13639), .B(n13640), .Z(n13551) );
  NANDN U13691 ( .A(n13641), .B(n13642), .Z(n13640) );
  NANDN U13692 ( .A(n13643), .B(n13644), .Z(n13642) );
  NANDN U13693 ( .A(n13644), .B(n13643), .Z(n13639) );
  ANDN U13694 ( .B(B[249]), .A(n60), .Z(n13553) );
  XNOR U13695 ( .A(n13561), .B(n13645), .Z(n13554) );
  XNOR U13696 ( .A(n13560), .B(n13558), .Z(n13645) );
  AND U13697 ( .A(n13646), .B(n13647), .Z(n13558) );
  NANDN U13698 ( .A(n13648), .B(n13649), .Z(n13647) );
  OR U13699 ( .A(n13650), .B(n13651), .Z(n13649) );
  NAND U13700 ( .A(n13651), .B(n13650), .Z(n13646) );
  ANDN U13701 ( .B(B[250]), .A(n61), .Z(n13560) );
  XNOR U13702 ( .A(n13568), .B(n13652), .Z(n13561) );
  XNOR U13703 ( .A(n13567), .B(n13565), .Z(n13652) );
  AND U13704 ( .A(n13653), .B(n13654), .Z(n13565) );
  NANDN U13705 ( .A(n13655), .B(n13656), .Z(n13654) );
  NANDN U13706 ( .A(n13657), .B(n13658), .Z(n13656) );
  NANDN U13707 ( .A(n13658), .B(n13657), .Z(n13653) );
  ANDN U13708 ( .B(B[251]), .A(n62), .Z(n13567) );
  XNOR U13709 ( .A(n13575), .B(n13659), .Z(n13568) );
  XNOR U13710 ( .A(n13574), .B(n13572), .Z(n13659) );
  AND U13711 ( .A(n13660), .B(n13661), .Z(n13572) );
  NANDN U13712 ( .A(n13662), .B(n13663), .Z(n13661) );
  OR U13713 ( .A(n13664), .B(n13665), .Z(n13663) );
  NAND U13714 ( .A(n13665), .B(n13664), .Z(n13660) );
  ANDN U13715 ( .B(B[252]), .A(n63), .Z(n13574) );
  XNOR U13716 ( .A(n13582), .B(n13666), .Z(n13575) );
  XNOR U13717 ( .A(n13581), .B(n13579), .Z(n13666) );
  AND U13718 ( .A(n13667), .B(n13668), .Z(n13579) );
  NANDN U13719 ( .A(n13669), .B(n13670), .Z(n13668) );
  NANDN U13720 ( .A(n13671), .B(n13672), .Z(n13670) );
  NANDN U13721 ( .A(n13672), .B(n13671), .Z(n13667) );
  ANDN U13722 ( .B(B[253]), .A(n64), .Z(n13581) );
  XOR U13723 ( .A(n13587), .B(n13673), .Z(n13582) );
  XOR U13724 ( .A(n13588), .B(n13589), .Z(n13673) );
  NAND U13725 ( .A(A[19]), .B(B[255]), .Z(n13589) );
  AND U13726 ( .A(B[254]), .B(A[20]), .Z(n13588) );
  NAND U13727 ( .A(n13674), .B(n13675), .Z(n13587) );
  NAND U13728 ( .A(n13676), .B(n13677), .Z(n13675) );
  NANDN U13729 ( .A(n13678), .B(n13679), .Z(n13676) );
  NANDN U13730 ( .A(n13679), .B(n13678), .Z(n13674) );
  NAND U13731 ( .A(n13680), .B(n13681), .Z(n248) );
  NANDN U13732 ( .A(n13682), .B(n13683), .Z(n13681) );
  OR U13733 ( .A(n13684), .B(n13685), .Z(n13683) );
  NAND U13734 ( .A(n13685), .B(n13684), .Z(n13680) );
  XOR U13735 ( .A(n250), .B(n249), .Z(\A1[271] ) );
  XOR U13736 ( .A(n13685), .B(n13686), .Z(n249) );
  XNOR U13737 ( .A(n13684), .B(n13682), .Z(n13686) );
  AND U13738 ( .A(n13687), .B(n13688), .Z(n13682) );
  NANDN U13739 ( .A(n13689), .B(n13690), .Z(n13688) );
  OR U13740 ( .A(n13691), .B(n13692), .Z(n13690) );
  NAND U13741 ( .A(n13692), .B(n13691), .Z(n13687) );
  ANDN U13742 ( .B(B[242]), .A(n54), .Z(n13684) );
  XNOR U13743 ( .A(n13602), .B(n13693), .Z(n13685) );
  XNOR U13744 ( .A(n13601), .B(n13599), .Z(n13693) );
  AND U13745 ( .A(n13694), .B(n13695), .Z(n13599) );
  NANDN U13746 ( .A(n13696), .B(n13697), .Z(n13695) );
  NANDN U13747 ( .A(n13698), .B(n13699), .Z(n13697) );
  NANDN U13748 ( .A(n13699), .B(n13698), .Z(n13694) );
  ANDN U13749 ( .B(B[243]), .A(n55), .Z(n13601) );
  XNOR U13750 ( .A(n13609), .B(n13700), .Z(n13602) );
  XNOR U13751 ( .A(n13608), .B(n13606), .Z(n13700) );
  AND U13752 ( .A(n13701), .B(n13702), .Z(n13606) );
  NANDN U13753 ( .A(n13703), .B(n13704), .Z(n13702) );
  OR U13754 ( .A(n13705), .B(n13706), .Z(n13704) );
  NAND U13755 ( .A(n13706), .B(n13705), .Z(n13701) );
  ANDN U13756 ( .B(B[244]), .A(n56), .Z(n13608) );
  XNOR U13757 ( .A(n13616), .B(n13707), .Z(n13609) );
  XNOR U13758 ( .A(n13615), .B(n13613), .Z(n13707) );
  AND U13759 ( .A(n13708), .B(n13709), .Z(n13613) );
  NANDN U13760 ( .A(n13710), .B(n13711), .Z(n13709) );
  NANDN U13761 ( .A(n13712), .B(n13713), .Z(n13711) );
  NANDN U13762 ( .A(n13713), .B(n13712), .Z(n13708) );
  ANDN U13763 ( .B(B[245]), .A(n57), .Z(n13615) );
  XNOR U13764 ( .A(n13623), .B(n13714), .Z(n13616) );
  XNOR U13765 ( .A(n13622), .B(n13620), .Z(n13714) );
  AND U13766 ( .A(n13715), .B(n13716), .Z(n13620) );
  NANDN U13767 ( .A(n13717), .B(n13718), .Z(n13716) );
  OR U13768 ( .A(n13719), .B(n13720), .Z(n13718) );
  NAND U13769 ( .A(n13720), .B(n13719), .Z(n13715) );
  ANDN U13770 ( .B(B[246]), .A(n58), .Z(n13622) );
  XNOR U13771 ( .A(n13630), .B(n13721), .Z(n13623) );
  XNOR U13772 ( .A(n13629), .B(n13627), .Z(n13721) );
  AND U13773 ( .A(n13722), .B(n13723), .Z(n13627) );
  NANDN U13774 ( .A(n13724), .B(n13725), .Z(n13723) );
  NANDN U13775 ( .A(n13726), .B(n13727), .Z(n13725) );
  NANDN U13776 ( .A(n13727), .B(n13726), .Z(n13722) );
  ANDN U13777 ( .B(B[247]), .A(n59), .Z(n13629) );
  XNOR U13778 ( .A(n13637), .B(n13728), .Z(n13630) );
  XNOR U13779 ( .A(n13636), .B(n13634), .Z(n13728) );
  AND U13780 ( .A(n13729), .B(n13730), .Z(n13634) );
  NANDN U13781 ( .A(n13731), .B(n13732), .Z(n13730) );
  OR U13782 ( .A(n13733), .B(n13734), .Z(n13732) );
  NAND U13783 ( .A(n13734), .B(n13733), .Z(n13729) );
  ANDN U13784 ( .B(B[248]), .A(n60), .Z(n13636) );
  XNOR U13785 ( .A(n13644), .B(n13735), .Z(n13637) );
  XNOR U13786 ( .A(n13643), .B(n13641), .Z(n13735) );
  AND U13787 ( .A(n13736), .B(n13737), .Z(n13641) );
  NANDN U13788 ( .A(n13738), .B(n13739), .Z(n13737) );
  NANDN U13789 ( .A(n13740), .B(n13741), .Z(n13739) );
  NANDN U13790 ( .A(n13741), .B(n13740), .Z(n13736) );
  ANDN U13791 ( .B(B[249]), .A(n61), .Z(n13643) );
  XNOR U13792 ( .A(n13651), .B(n13742), .Z(n13644) );
  XNOR U13793 ( .A(n13650), .B(n13648), .Z(n13742) );
  AND U13794 ( .A(n13743), .B(n13744), .Z(n13648) );
  NANDN U13795 ( .A(n13745), .B(n13746), .Z(n13744) );
  OR U13796 ( .A(n13747), .B(n13748), .Z(n13746) );
  NAND U13797 ( .A(n13748), .B(n13747), .Z(n13743) );
  ANDN U13798 ( .B(B[250]), .A(n62), .Z(n13650) );
  XNOR U13799 ( .A(n13658), .B(n13749), .Z(n13651) );
  XNOR U13800 ( .A(n13657), .B(n13655), .Z(n13749) );
  AND U13801 ( .A(n13750), .B(n13751), .Z(n13655) );
  NANDN U13802 ( .A(n13752), .B(n13753), .Z(n13751) );
  NANDN U13803 ( .A(n13754), .B(n13755), .Z(n13753) );
  NANDN U13804 ( .A(n13755), .B(n13754), .Z(n13750) );
  ANDN U13805 ( .B(B[251]), .A(n63), .Z(n13657) );
  XNOR U13806 ( .A(n13665), .B(n13756), .Z(n13658) );
  XNOR U13807 ( .A(n13664), .B(n13662), .Z(n13756) );
  AND U13808 ( .A(n13757), .B(n13758), .Z(n13662) );
  NANDN U13809 ( .A(n13759), .B(n13760), .Z(n13758) );
  OR U13810 ( .A(n13761), .B(n13762), .Z(n13760) );
  NAND U13811 ( .A(n13762), .B(n13761), .Z(n13757) );
  ANDN U13812 ( .B(B[252]), .A(n64), .Z(n13664) );
  XNOR U13813 ( .A(n13672), .B(n13763), .Z(n13665) );
  XNOR U13814 ( .A(n13671), .B(n13669), .Z(n13763) );
  AND U13815 ( .A(n13764), .B(n13765), .Z(n13669) );
  NANDN U13816 ( .A(n13766), .B(n13767), .Z(n13765) );
  NANDN U13817 ( .A(n13768), .B(n13769), .Z(n13767) );
  NANDN U13818 ( .A(n13769), .B(n13768), .Z(n13764) );
  ANDN U13819 ( .B(B[253]), .A(n65), .Z(n13671) );
  XOR U13820 ( .A(n13677), .B(n13770), .Z(n13672) );
  XOR U13821 ( .A(n13678), .B(n13679), .Z(n13770) );
  NAND U13822 ( .A(A[18]), .B(B[255]), .Z(n13679) );
  AND U13823 ( .A(B[254]), .B(A[19]), .Z(n13678) );
  NAND U13824 ( .A(n13771), .B(n13772), .Z(n13677) );
  NAND U13825 ( .A(n13773), .B(n13774), .Z(n13772) );
  NANDN U13826 ( .A(n13775), .B(n13776), .Z(n13773) );
  NANDN U13827 ( .A(n13776), .B(n13775), .Z(n13771) );
  NAND U13828 ( .A(n13777), .B(n13778), .Z(n250) );
  NANDN U13829 ( .A(n13779), .B(n13780), .Z(n13778) );
  NAND U13830 ( .A(n13782), .B(n13781), .Z(n13777) );
  XOR U13831 ( .A(n252), .B(n251), .Z(\A1[270] ) );
  XOR U13832 ( .A(n13782), .B(n13783), .Z(n251) );
  XNOR U13833 ( .A(n13781), .B(n13779), .Z(n13783) );
  AND U13834 ( .A(n13784), .B(n13785), .Z(n13779) );
  NANDN U13835 ( .A(n13786), .B(n13787), .Z(n13785) );
  NANDN U13836 ( .A(n13788), .B(n13789), .Z(n13787) );
  NANDN U13837 ( .A(n13789), .B(n13788), .Z(n13784) );
  ANDN U13838 ( .B(B[241]), .A(n54), .Z(n13781) );
  XOR U13839 ( .A(n13692), .B(n13790), .Z(n13782) );
  XNOR U13840 ( .A(n13691), .B(n13689), .Z(n13790) );
  AND U13841 ( .A(n13791), .B(n13792), .Z(n13689) );
  NANDN U13842 ( .A(n13793), .B(n13794), .Z(n13792) );
  OR U13843 ( .A(n13795), .B(n13796), .Z(n13794) );
  NAND U13844 ( .A(n13796), .B(n13795), .Z(n13791) );
  ANDN U13845 ( .B(B[242]), .A(n55), .Z(n13691) );
  XNOR U13846 ( .A(n13699), .B(n13797), .Z(n13692) );
  XNOR U13847 ( .A(n13698), .B(n13696), .Z(n13797) );
  AND U13848 ( .A(n13798), .B(n13799), .Z(n13696) );
  NANDN U13849 ( .A(n13800), .B(n13801), .Z(n13799) );
  NANDN U13850 ( .A(n13802), .B(n13803), .Z(n13801) );
  NANDN U13851 ( .A(n13803), .B(n13802), .Z(n13798) );
  ANDN U13852 ( .B(B[243]), .A(n56), .Z(n13698) );
  XNOR U13853 ( .A(n13706), .B(n13804), .Z(n13699) );
  XNOR U13854 ( .A(n13705), .B(n13703), .Z(n13804) );
  AND U13855 ( .A(n13805), .B(n13806), .Z(n13703) );
  NANDN U13856 ( .A(n13807), .B(n13808), .Z(n13806) );
  OR U13857 ( .A(n13809), .B(n13810), .Z(n13808) );
  NAND U13858 ( .A(n13810), .B(n13809), .Z(n13805) );
  ANDN U13859 ( .B(B[244]), .A(n57), .Z(n13705) );
  XNOR U13860 ( .A(n13713), .B(n13811), .Z(n13706) );
  XNOR U13861 ( .A(n13712), .B(n13710), .Z(n13811) );
  AND U13862 ( .A(n13812), .B(n13813), .Z(n13710) );
  NANDN U13863 ( .A(n13814), .B(n13815), .Z(n13813) );
  NANDN U13864 ( .A(n13816), .B(n13817), .Z(n13815) );
  NANDN U13865 ( .A(n13817), .B(n13816), .Z(n13812) );
  ANDN U13866 ( .B(B[245]), .A(n58), .Z(n13712) );
  XNOR U13867 ( .A(n13720), .B(n13818), .Z(n13713) );
  XNOR U13868 ( .A(n13719), .B(n13717), .Z(n13818) );
  AND U13869 ( .A(n13819), .B(n13820), .Z(n13717) );
  NANDN U13870 ( .A(n13821), .B(n13822), .Z(n13820) );
  OR U13871 ( .A(n13823), .B(n13824), .Z(n13822) );
  NAND U13872 ( .A(n13824), .B(n13823), .Z(n13819) );
  ANDN U13873 ( .B(B[246]), .A(n59), .Z(n13719) );
  XNOR U13874 ( .A(n13727), .B(n13825), .Z(n13720) );
  XNOR U13875 ( .A(n13726), .B(n13724), .Z(n13825) );
  AND U13876 ( .A(n13826), .B(n13827), .Z(n13724) );
  NANDN U13877 ( .A(n13828), .B(n13829), .Z(n13827) );
  NANDN U13878 ( .A(n13830), .B(n13831), .Z(n13829) );
  NANDN U13879 ( .A(n13831), .B(n13830), .Z(n13826) );
  ANDN U13880 ( .B(B[247]), .A(n60), .Z(n13726) );
  XNOR U13881 ( .A(n13734), .B(n13832), .Z(n13727) );
  XNOR U13882 ( .A(n13733), .B(n13731), .Z(n13832) );
  AND U13883 ( .A(n13833), .B(n13834), .Z(n13731) );
  NANDN U13884 ( .A(n13835), .B(n13836), .Z(n13834) );
  OR U13885 ( .A(n13837), .B(n13838), .Z(n13836) );
  NAND U13886 ( .A(n13838), .B(n13837), .Z(n13833) );
  ANDN U13887 ( .B(B[248]), .A(n61), .Z(n13733) );
  XNOR U13888 ( .A(n13741), .B(n13839), .Z(n13734) );
  XNOR U13889 ( .A(n13740), .B(n13738), .Z(n13839) );
  AND U13890 ( .A(n13840), .B(n13841), .Z(n13738) );
  NANDN U13891 ( .A(n13842), .B(n13843), .Z(n13841) );
  NANDN U13892 ( .A(n13844), .B(n13845), .Z(n13843) );
  NANDN U13893 ( .A(n13845), .B(n13844), .Z(n13840) );
  ANDN U13894 ( .B(B[249]), .A(n62), .Z(n13740) );
  XNOR U13895 ( .A(n13748), .B(n13846), .Z(n13741) );
  XNOR U13896 ( .A(n13747), .B(n13745), .Z(n13846) );
  AND U13897 ( .A(n13847), .B(n13848), .Z(n13745) );
  NANDN U13898 ( .A(n13849), .B(n13850), .Z(n13848) );
  OR U13899 ( .A(n13851), .B(n13852), .Z(n13850) );
  NAND U13900 ( .A(n13852), .B(n13851), .Z(n13847) );
  ANDN U13901 ( .B(B[250]), .A(n63), .Z(n13747) );
  XNOR U13902 ( .A(n13755), .B(n13853), .Z(n13748) );
  XNOR U13903 ( .A(n13754), .B(n13752), .Z(n13853) );
  AND U13904 ( .A(n13854), .B(n13855), .Z(n13752) );
  NANDN U13905 ( .A(n13856), .B(n13857), .Z(n13855) );
  NANDN U13906 ( .A(n13858), .B(n13859), .Z(n13857) );
  NANDN U13907 ( .A(n13859), .B(n13858), .Z(n13854) );
  ANDN U13908 ( .B(B[251]), .A(n64), .Z(n13754) );
  XNOR U13909 ( .A(n13762), .B(n13860), .Z(n13755) );
  XNOR U13910 ( .A(n13761), .B(n13759), .Z(n13860) );
  AND U13911 ( .A(n13861), .B(n13862), .Z(n13759) );
  NANDN U13912 ( .A(n13863), .B(n13864), .Z(n13862) );
  OR U13913 ( .A(n13865), .B(n13866), .Z(n13864) );
  NAND U13914 ( .A(n13866), .B(n13865), .Z(n13861) );
  ANDN U13915 ( .B(B[252]), .A(n65), .Z(n13761) );
  XNOR U13916 ( .A(n13769), .B(n13867), .Z(n13762) );
  XNOR U13917 ( .A(n13768), .B(n13766), .Z(n13867) );
  AND U13918 ( .A(n13868), .B(n13869), .Z(n13766) );
  NANDN U13919 ( .A(n13870), .B(n13871), .Z(n13869) );
  NANDN U13920 ( .A(n13872), .B(n13873), .Z(n13871) );
  NANDN U13921 ( .A(n13873), .B(n13872), .Z(n13868) );
  ANDN U13922 ( .B(B[253]), .A(n66), .Z(n13768) );
  XOR U13923 ( .A(n13774), .B(n13874), .Z(n13769) );
  XOR U13924 ( .A(n13775), .B(n13776), .Z(n13874) );
  NAND U13925 ( .A(A[17]), .B(B[255]), .Z(n13776) );
  AND U13926 ( .A(B[254]), .B(A[18]), .Z(n13775) );
  NAND U13927 ( .A(n13875), .B(n13876), .Z(n13774) );
  NAND U13928 ( .A(n13877), .B(n13878), .Z(n13876) );
  NANDN U13929 ( .A(n13879), .B(n13880), .Z(n13877) );
  NANDN U13930 ( .A(n13880), .B(n13879), .Z(n13875) );
  NAND U13931 ( .A(n13881), .B(n13882), .Z(n252) );
  NANDN U13932 ( .A(n13883), .B(n13884), .Z(n13882) );
  OR U13933 ( .A(n13885), .B(n13886), .Z(n13884) );
  NAND U13934 ( .A(n13886), .B(n13885), .Z(n13881) );
  XOR U13935 ( .A(n12975), .B(n13887), .Z(\A1[26] ) );
  XNOR U13936 ( .A(n12974), .B(n12973), .Z(n13887) );
  NAND U13937 ( .A(n13888), .B(n13889), .Z(n12973) );
  NANDN U13938 ( .A(n13890), .B(n13891), .Z(n13889) );
  OR U13939 ( .A(n13892), .B(n13893), .Z(n13891) );
  NAND U13940 ( .A(n13893), .B(n13892), .Z(n13888) );
  ANDN U13941 ( .B(B[0]), .A(n57), .Z(n12974) );
  XNOR U13942 ( .A(n12982), .B(n13894), .Z(n12975) );
  XNOR U13943 ( .A(n12981), .B(n12979), .Z(n13894) );
  AND U13944 ( .A(n13895), .B(n13896), .Z(n12979) );
  NANDN U13945 ( .A(n13897), .B(n13898), .Z(n13896) );
  NANDN U13946 ( .A(n13899), .B(n13900), .Z(n13898) );
  NANDN U13947 ( .A(n13900), .B(n13899), .Z(n13895) );
  ANDN U13948 ( .B(B[1]), .A(n58), .Z(n12981) );
  XNOR U13949 ( .A(n12989), .B(n13901), .Z(n12982) );
  XNOR U13950 ( .A(n12988), .B(n12986), .Z(n13901) );
  AND U13951 ( .A(n13902), .B(n13903), .Z(n12986) );
  NANDN U13952 ( .A(n13904), .B(n13905), .Z(n13903) );
  OR U13953 ( .A(n13906), .B(n13907), .Z(n13905) );
  NAND U13954 ( .A(n13907), .B(n13906), .Z(n13902) );
  ANDN U13955 ( .B(B[2]), .A(n59), .Z(n12988) );
  XNOR U13956 ( .A(n12996), .B(n13908), .Z(n12989) );
  XNOR U13957 ( .A(n12995), .B(n12993), .Z(n13908) );
  AND U13958 ( .A(n13909), .B(n13910), .Z(n12993) );
  NANDN U13959 ( .A(n13911), .B(n13912), .Z(n13910) );
  NANDN U13960 ( .A(n13913), .B(n13914), .Z(n13912) );
  NANDN U13961 ( .A(n13914), .B(n13913), .Z(n13909) );
  ANDN U13962 ( .B(B[3]), .A(n60), .Z(n12995) );
  XNOR U13963 ( .A(n13003), .B(n13915), .Z(n12996) );
  XNOR U13964 ( .A(n13002), .B(n13000), .Z(n13915) );
  AND U13965 ( .A(n13916), .B(n13917), .Z(n13000) );
  NANDN U13966 ( .A(n13918), .B(n13919), .Z(n13917) );
  OR U13967 ( .A(n13920), .B(n13921), .Z(n13919) );
  NAND U13968 ( .A(n13921), .B(n13920), .Z(n13916) );
  ANDN U13969 ( .B(B[4]), .A(n61), .Z(n13002) );
  XNOR U13970 ( .A(n13010), .B(n13922), .Z(n13003) );
  XNOR U13971 ( .A(n13009), .B(n13007), .Z(n13922) );
  AND U13972 ( .A(n13923), .B(n13924), .Z(n13007) );
  NANDN U13973 ( .A(n13925), .B(n13926), .Z(n13924) );
  NANDN U13974 ( .A(n13927), .B(n13928), .Z(n13926) );
  NANDN U13975 ( .A(n13928), .B(n13927), .Z(n13923) );
  ANDN U13976 ( .B(B[5]), .A(n62), .Z(n13009) );
  XNOR U13977 ( .A(n13017), .B(n13929), .Z(n13010) );
  XNOR U13978 ( .A(n13016), .B(n13014), .Z(n13929) );
  AND U13979 ( .A(n13930), .B(n13931), .Z(n13014) );
  NANDN U13980 ( .A(n13932), .B(n13933), .Z(n13931) );
  OR U13981 ( .A(n13934), .B(n13935), .Z(n13933) );
  NAND U13982 ( .A(n13935), .B(n13934), .Z(n13930) );
  ANDN U13983 ( .B(B[6]), .A(n63), .Z(n13016) );
  XNOR U13984 ( .A(n13024), .B(n13936), .Z(n13017) );
  XNOR U13985 ( .A(n13023), .B(n13021), .Z(n13936) );
  AND U13986 ( .A(n13937), .B(n13938), .Z(n13021) );
  NANDN U13987 ( .A(n13939), .B(n13940), .Z(n13938) );
  NANDN U13988 ( .A(n13941), .B(n13942), .Z(n13940) );
  NANDN U13989 ( .A(n13942), .B(n13941), .Z(n13937) );
  ANDN U13990 ( .B(B[7]), .A(n64), .Z(n13023) );
  XNOR U13991 ( .A(n13031), .B(n13943), .Z(n13024) );
  XNOR U13992 ( .A(n13030), .B(n13028), .Z(n13943) );
  AND U13993 ( .A(n13944), .B(n13945), .Z(n13028) );
  NANDN U13994 ( .A(n13946), .B(n13947), .Z(n13945) );
  OR U13995 ( .A(n13948), .B(n13949), .Z(n13947) );
  NAND U13996 ( .A(n13949), .B(n13948), .Z(n13944) );
  ANDN U13997 ( .B(B[8]), .A(n65), .Z(n13030) );
  XNOR U13998 ( .A(n13038), .B(n13950), .Z(n13031) );
  XNOR U13999 ( .A(n13037), .B(n13035), .Z(n13950) );
  AND U14000 ( .A(n13951), .B(n13952), .Z(n13035) );
  NANDN U14001 ( .A(n13953), .B(n13954), .Z(n13952) );
  NANDN U14002 ( .A(n13955), .B(n13956), .Z(n13954) );
  NANDN U14003 ( .A(n13956), .B(n13955), .Z(n13951) );
  ANDN U14004 ( .B(B[9]), .A(n66), .Z(n13037) );
  XNOR U14005 ( .A(n13045), .B(n13957), .Z(n13038) );
  XNOR U14006 ( .A(n13044), .B(n13042), .Z(n13957) );
  AND U14007 ( .A(n13958), .B(n13959), .Z(n13042) );
  NANDN U14008 ( .A(n13960), .B(n13961), .Z(n13959) );
  OR U14009 ( .A(n13962), .B(n13963), .Z(n13961) );
  NAND U14010 ( .A(n13963), .B(n13962), .Z(n13958) );
  ANDN U14011 ( .B(B[10]), .A(n67), .Z(n13044) );
  XNOR U14012 ( .A(n13052), .B(n13964), .Z(n13045) );
  XNOR U14013 ( .A(n13051), .B(n13049), .Z(n13964) );
  AND U14014 ( .A(n13965), .B(n13966), .Z(n13049) );
  NANDN U14015 ( .A(n13967), .B(n13968), .Z(n13966) );
  NANDN U14016 ( .A(n13969), .B(n13970), .Z(n13968) );
  NANDN U14017 ( .A(n13970), .B(n13969), .Z(n13965) );
  ANDN U14018 ( .B(B[11]), .A(n68), .Z(n13051) );
  XNOR U14019 ( .A(n13059), .B(n13971), .Z(n13052) );
  XNOR U14020 ( .A(n13058), .B(n13056), .Z(n13971) );
  AND U14021 ( .A(n13972), .B(n13973), .Z(n13056) );
  NANDN U14022 ( .A(n13974), .B(n13975), .Z(n13973) );
  OR U14023 ( .A(n13976), .B(n13977), .Z(n13975) );
  NAND U14024 ( .A(n13977), .B(n13976), .Z(n13972) );
  ANDN U14025 ( .B(B[12]), .A(n69), .Z(n13058) );
  XNOR U14026 ( .A(n13066), .B(n13978), .Z(n13059) );
  XNOR U14027 ( .A(n13065), .B(n13063), .Z(n13978) );
  AND U14028 ( .A(n13979), .B(n13980), .Z(n13063) );
  NANDN U14029 ( .A(n13981), .B(n13982), .Z(n13980) );
  NANDN U14030 ( .A(n13983), .B(n13984), .Z(n13982) );
  NANDN U14031 ( .A(n13984), .B(n13983), .Z(n13979) );
  ANDN U14032 ( .B(B[13]), .A(n70), .Z(n13065) );
  XNOR U14033 ( .A(n13073), .B(n13985), .Z(n13066) );
  XNOR U14034 ( .A(n13072), .B(n13070), .Z(n13985) );
  AND U14035 ( .A(n13986), .B(n13987), .Z(n13070) );
  NANDN U14036 ( .A(n13988), .B(n13989), .Z(n13987) );
  OR U14037 ( .A(n13990), .B(n13991), .Z(n13989) );
  NAND U14038 ( .A(n13991), .B(n13990), .Z(n13986) );
  ANDN U14039 ( .B(B[14]), .A(n71), .Z(n13072) );
  XNOR U14040 ( .A(n13080), .B(n13992), .Z(n13073) );
  XNOR U14041 ( .A(n13079), .B(n13077), .Z(n13992) );
  AND U14042 ( .A(n13993), .B(n13994), .Z(n13077) );
  NANDN U14043 ( .A(n13995), .B(n13996), .Z(n13994) );
  NANDN U14044 ( .A(n13997), .B(n13998), .Z(n13996) );
  NANDN U14045 ( .A(n13998), .B(n13997), .Z(n13993) );
  ANDN U14046 ( .B(B[15]), .A(n72), .Z(n13079) );
  XNOR U14047 ( .A(n13087), .B(n13999), .Z(n13080) );
  XNOR U14048 ( .A(n13086), .B(n13084), .Z(n13999) );
  AND U14049 ( .A(n14000), .B(n14001), .Z(n13084) );
  NANDN U14050 ( .A(n14002), .B(n14003), .Z(n14001) );
  OR U14051 ( .A(n14004), .B(n14005), .Z(n14003) );
  NAND U14052 ( .A(n14005), .B(n14004), .Z(n14000) );
  ANDN U14053 ( .B(B[16]), .A(n73), .Z(n13086) );
  XNOR U14054 ( .A(n13094), .B(n14006), .Z(n13087) );
  XNOR U14055 ( .A(n13093), .B(n13091), .Z(n14006) );
  AND U14056 ( .A(n14007), .B(n14008), .Z(n13091) );
  NANDN U14057 ( .A(n14009), .B(n14010), .Z(n14008) );
  NANDN U14058 ( .A(n14011), .B(n14012), .Z(n14010) );
  NANDN U14059 ( .A(n14012), .B(n14011), .Z(n14007) );
  ANDN U14060 ( .B(B[17]), .A(n74), .Z(n13093) );
  XNOR U14061 ( .A(n13101), .B(n14013), .Z(n13094) );
  XNOR U14062 ( .A(n13100), .B(n13098), .Z(n14013) );
  AND U14063 ( .A(n14014), .B(n14015), .Z(n13098) );
  NANDN U14064 ( .A(n14016), .B(n14017), .Z(n14015) );
  OR U14065 ( .A(n14018), .B(n14019), .Z(n14017) );
  NAND U14066 ( .A(n14019), .B(n14018), .Z(n14014) );
  ANDN U14067 ( .B(B[18]), .A(n75), .Z(n13100) );
  XNOR U14068 ( .A(n13108), .B(n14020), .Z(n13101) );
  XNOR U14069 ( .A(n13107), .B(n13105), .Z(n14020) );
  AND U14070 ( .A(n14021), .B(n14022), .Z(n13105) );
  NANDN U14071 ( .A(n14023), .B(n14024), .Z(n14022) );
  NANDN U14072 ( .A(n14025), .B(n14026), .Z(n14024) );
  NANDN U14073 ( .A(n14026), .B(n14025), .Z(n14021) );
  ANDN U14074 ( .B(B[19]), .A(n76), .Z(n13107) );
  XNOR U14075 ( .A(n13115), .B(n14027), .Z(n13108) );
  XNOR U14076 ( .A(n13114), .B(n13112), .Z(n14027) );
  AND U14077 ( .A(n14028), .B(n14029), .Z(n13112) );
  NANDN U14078 ( .A(n14030), .B(n14031), .Z(n14029) );
  OR U14079 ( .A(n14032), .B(n14033), .Z(n14031) );
  NAND U14080 ( .A(n14033), .B(n14032), .Z(n14028) );
  ANDN U14081 ( .B(B[20]), .A(n77), .Z(n13114) );
  XNOR U14082 ( .A(n13122), .B(n14034), .Z(n13115) );
  XNOR U14083 ( .A(n13121), .B(n13119), .Z(n14034) );
  AND U14084 ( .A(n14035), .B(n14036), .Z(n13119) );
  NANDN U14085 ( .A(n14037), .B(n14038), .Z(n14036) );
  NANDN U14086 ( .A(n14039), .B(n14040), .Z(n14038) );
  NANDN U14087 ( .A(n14040), .B(n14039), .Z(n14035) );
  ANDN U14088 ( .B(B[21]), .A(n78), .Z(n13121) );
  XNOR U14089 ( .A(n13129), .B(n14041), .Z(n13122) );
  XNOR U14090 ( .A(n13128), .B(n13126), .Z(n14041) );
  AND U14091 ( .A(n14042), .B(n14043), .Z(n13126) );
  NANDN U14092 ( .A(n14044), .B(n14045), .Z(n14043) );
  OR U14093 ( .A(n14046), .B(n14047), .Z(n14045) );
  NAND U14094 ( .A(n14047), .B(n14046), .Z(n14042) );
  ANDN U14095 ( .B(B[22]), .A(n79), .Z(n13128) );
  XNOR U14096 ( .A(n13136), .B(n14048), .Z(n13129) );
  XNOR U14097 ( .A(n13135), .B(n13133), .Z(n14048) );
  AND U14098 ( .A(n14049), .B(n14050), .Z(n13133) );
  NANDN U14099 ( .A(n14051), .B(n14052), .Z(n14050) );
  NANDN U14100 ( .A(n14053), .B(n14054), .Z(n14052) );
  NANDN U14101 ( .A(n14054), .B(n14053), .Z(n14049) );
  ANDN U14102 ( .B(B[23]), .A(n80), .Z(n13135) );
  XNOR U14103 ( .A(n13143), .B(n14055), .Z(n13136) );
  XNOR U14104 ( .A(n13142), .B(n13140), .Z(n14055) );
  AND U14105 ( .A(n14056), .B(n14057), .Z(n13140) );
  NANDN U14106 ( .A(n14058), .B(n14059), .Z(n14057) );
  OR U14107 ( .A(n14060), .B(n14061), .Z(n14059) );
  NAND U14108 ( .A(n14061), .B(n14060), .Z(n14056) );
  ANDN U14109 ( .B(B[24]), .A(n81), .Z(n13142) );
  XNOR U14110 ( .A(n13150), .B(n14062), .Z(n13143) );
  XNOR U14111 ( .A(n13149), .B(n13147), .Z(n14062) );
  AND U14112 ( .A(n14063), .B(n14064), .Z(n13147) );
  NANDN U14113 ( .A(n14065), .B(n14066), .Z(n14064) );
  NAND U14114 ( .A(n14067), .B(n14068), .Z(n14066) );
  ANDN U14115 ( .B(B[25]), .A(n82), .Z(n13149) );
  XOR U14116 ( .A(n13156), .B(n14069), .Z(n13150) );
  XNOR U14117 ( .A(n13154), .B(n13157), .Z(n14069) );
  NAND U14118 ( .A(A[2]), .B(B[26]), .Z(n13157) );
  NANDN U14119 ( .A(n14070), .B(n14071), .Z(n13154) );
  AND U14120 ( .A(A[0]), .B(B[27]), .Z(n14071) );
  XNOR U14121 ( .A(n13159), .B(n14072), .Z(n13156) );
  NAND U14122 ( .A(A[0]), .B(B[28]), .Z(n14072) );
  NAND U14123 ( .A(B[27]), .B(A[1]), .Z(n13159) );
  XOR U14124 ( .A(n254), .B(n253), .Z(\A1[269] ) );
  XOR U14125 ( .A(n13886), .B(n14073), .Z(n253) );
  XNOR U14126 ( .A(n13885), .B(n13883), .Z(n14073) );
  AND U14127 ( .A(n14074), .B(n14075), .Z(n13883) );
  NANDN U14128 ( .A(n14076), .B(n14077), .Z(n14075) );
  OR U14129 ( .A(n14078), .B(n14079), .Z(n14077) );
  NAND U14130 ( .A(n14079), .B(n14078), .Z(n14074) );
  ANDN U14131 ( .B(B[240]), .A(n54), .Z(n13885) );
  XNOR U14132 ( .A(n13789), .B(n14080), .Z(n13886) );
  XNOR U14133 ( .A(n13788), .B(n13786), .Z(n14080) );
  AND U14134 ( .A(n14081), .B(n14082), .Z(n13786) );
  NANDN U14135 ( .A(n14083), .B(n14084), .Z(n14082) );
  NANDN U14136 ( .A(n14085), .B(n14086), .Z(n14084) );
  NANDN U14137 ( .A(n14086), .B(n14085), .Z(n14081) );
  ANDN U14138 ( .B(B[241]), .A(n55), .Z(n13788) );
  XNOR U14139 ( .A(n13796), .B(n14087), .Z(n13789) );
  XNOR U14140 ( .A(n13795), .B(n13793), .Z(n14087) );
  AND U14141 ( .A(n14088), .B(n14089), .Z(n13793) );
  NANDN U14142 ( .A(n14090), .B(n14091), .Z(n14089) );
  OR U14143 ( .A(n14092), .B(n14093), .Z(n14091) );
  NAND U14144 ( .A(n14093), .B(n14092), .Z(n14088) );
  ANDN U14145 ( .B(B[242]), .A(n56), .Z(n13795) );
  XNOR U14146 ( .A(n13803), .B(n14094), .Z(n13796) );
  XNOR U14147 ( .A(n13802), .B(n13800), .Z(n14094) );
  AND U14148 ( .A(n14095), .B(n14096), .Z(n13800) );
  NANDN U14149 ( .A(n14097), .B(n14098), .Z(n14096) );
  NANDN U14150 ( .A(n14099), .B(n14100), .Z(n14098) );
  NANDN U14151 ( .A(n14100), .B(n14099), .Z(n14095) );
  ANDN U14152 ( .B(B[243]), .A(n57), .Z(n13802) );
  XNOR U14153 ( .A(n13810), .B(n14101), .Z(n13803) );
  XNOR U14154 ( .A(n13809), .B(n13807), .Z(n14101) );
  AND U14155 ( .A(n14102), .B(n14103), .Z(n13807) );
  NANDN U14156 ( .A(n14104), .B(n14105), .Z(n14103) );
  OR U14157 ( .A(n14106), .B(n14107), .Z(n14105) );
  NAND U14158 ( .A(n14107), .B(n14106), .Z(n14102) );
  ANDN U14159 ( .B(B[244]), .A(n58), .Z(n13809) );
  XNOR U14160 ( .A(n13817), .B(n14108), .Z(n13810) );
  XNOR U14161 ( .A(n13816), .B(n13814), .Z(n14108) );
  AND U14162 ( .A(n14109), .B(n14110), .Z(n13814) );
  NANDN U14163 ( .A(n14111), .B(n14112), .Z(n14110) );
  NANDN U14164 ( .A(n14113), .B(n14114), .Z(n14112) );
  NANDN U14165 ( .A(n14114), .B(n14113), .Z(n14109) );
  ANDN U14166 ( .B(B[245]), .A(n59), .Z(n13816) );
  XNOR U14167 ( .A(n13824), .B(n14115), .Z(n13817) );
  XNOR U14168 ( .A(n13823), .B(n13821), .Z(n14115) );
  AND U14169 ( .A(n14116), .B(n14117), .Z(n13821) );
  NANDN U14170 ( .A(n14118), .B(n14119), .Z(n14117) );
  OR U14171 ( .A(n14120), .B(n14121), .Z(n14119) );
  NAND U14172 ( .A(n14121), .B(n14120), .Z(n14116) );
  ANDN U14173 ( .B(B[246]), .A(n60), .Z(n13823) );
  XNOR U14174 ( .A(n13831), .B(n14122), .Z(n13824) );
  XNOR U14175 ( .A(n13830), .B(n13828), .Z(n14122) );
  AND U14176 ( .A(n14123), .B(n14124), .Z(n13828) );
  NANDN U14177 ( .A(n14125), .B(n14126), .Z(n14124) );
  NANDN U14178 ( .A(n14127), .B(n14128), .Z(n14126) );
  NANDN U14179 ( .A(n14128), .B(n14127), .Z(n14123) );
  ANDN U14180 ( .B(B[247]), .A(n61), .Z(n13830) );
  XNOR U14181 ( .A(n13838), .B(n14129), .Z(n13831) );
  XNOR U14182 ( .A(n13837), .B(n13835), .Z(n14129) );
  AND U14183 ( .A(n14130), .B(n14131), .Z(n13835) );
  NANDN U14184 ( .A(n14132), .B(n14133), .Z(n14131) );
  OR U14185 ( .A(n14134), .B(n14135), .Z(n14133) );
  NAND U14186 ( .A(n14135), .B(n14134), .Z(n14130) );
  ANDN U14187 ( .B(B[248]), .A(n62), .Z(n13837) );
  XNOR U14188 ( .A(n13845), .B(n14136), .Z(n13838) );
  XNOR U14189 ( .A(n13844), .B(n13842), .Z(n14136) );
  AND U14190 ( .A(n14137), .B(n14138), .Z(n13842) );
  NANDN U14191 ( .A(n14139), .B(n14140), .Z(n14138) );
  NANDN U14192 ( .A(n14141), .B(n14142), .Z(n14140) );
  NANDN U14193 ( .A(n14142), .B(n14141), .Z(n14137) );
  ANDN U14194 ( .B(B[249]), .A(n63), .Z(n13844) );
  XNOR U14195 ( .A(n13852), .B(n14143), .Z(n13845) );
  XNOR U14196 ( .A(n13851), .B(n13849), .Z(n14143) );
  AND U14197 ( .A(n14144), .B(n14145), .Z(n13849) );
  NANDN U14198 ( .A(n14146), .B(n14147), .Z(n14145) );
  OR U14199 ( .A(n14148), .B(n14149), .Z(n14147) );
  NAND U14200 ( .A(n14149), .B(n14148), .Z(n14144) );
  ANDN U14201 ( .B(B[250]), .A(n64), .Z(n13851) );
  XNOR U14202 ( .A(n13859), .B(n14150), .Z(n13852) );
  XNOR U14203 ( .A(n13858), .B(n13856), .Z(n14150) );
  AND U14204 ( .A(n14151), .B(n14152), .Z(n13856) );
  NANDN U14205 ( .A(n14153), .B(n14154), .Z(n14152) );
  NANDN U14206 ( .A(n14155), .B(n14156), .Z(n14154) );
  NANDN U14207 ( .A(n14156), .B(n14155), .Z(n14151) );
  ANDN U14208 ( .B(B[251]), .A(n65), .Z(n13858) );
  XNOR U14209 ( .A(n13866), .B(n14157), .Z(n13859) );
  XNOR U14210 ( .A(n13865), .B(n13863), .Z(n14157) );
  AND U14211 ( .A(n14158), .B(n14159), .Z(n13863) );
  NANDN U14212 ( .A(n14160), .B(n14161), .Z(n14159) );
  OR U14213 ( .A(n14162), .B(n14163), .Z(n14161) );
  NAND U14214 ( .A(n14163), .B(n14162), .Z(n14158) );
  ANDN U14215 ( .B(B[252]), .A(n66), .Z(n13865) );
  XNOR U14216 ( .A(n13873), .B(n14164), .Z(n13866) );
  XNOR U14217 ( .A(n13872), .B(n13870), .Z(n14164) );
  AND U14218 ( .A(n14165), .B(n14166), .Z(n13870) );
  NANDN U14219 ( .A(n14167), .B(n14168), .Z(n14166) );
  NANDN U14220 ( .A(n14169), .B(n14170), .Z(n14168) );
  NANDN U14221 ( .A(n14170), .B(n14169), .Z(n14165) );
  ANDN U14222 ( .B(B[253]), .A(n67), .Z(n13872) );
  XOR U14223 ( .A(n13878), .B(n14171), .Z(n13873) );
  XOR U14224 ( .A(n13879), .B(n13880), .Z(n14171) );
  NAND U14225 ( .A(A[16]), .B(B[255]), .Z(n13880) );
  AND U14226 ( .A(B[254]), .B(A[17]), .Z(n13879) );
  NAND U14227 ( .A(n14172), .B(n14173), .Z(n13878) );
  NAND U14228 ( .A(n14174), .B(n14175), .Z(n14173) );
  NANDN U14229 ( .A(n14176), .B(n14177), .Z(n14174) );
  NANDN U14230 ( .A(n14177), .B(n14176), .Z(n14172) );
  NAND U14231 ( .A(n14178), .B(n14179), .Z(n254) );
  NANDN U14232 ( .A(n14180), .B(n14181), .Z(n14179) );
  NAND U14233 ( .A(n14183), .B(n14182), .Z(n14178) );
  XOR U14234 ( .A(n256), .B(n255), .Z(\A1[268] ) );
  XOR U14235 ( .A(n14183), .B(n14184), .Z(n255) );
  XNOR U14236 ( .A(n14182), .B(n14180), .Z(n14184) );
  AND U14237 ( .A(n14185), .B(n14186), .Z(n14180) );
  NANDN U14238 ( .A(n14187), .B(n14188), .Z(n14186) );
  NANDN U14239 ( .A(n14189), .B(n14190), .Z(n14188) );
  NANDN U14240 ( .A(n14190), .B(n14189), .Z(n14185) );
  ANDN U14241 ( .B(B[239]), .A(n54), .Z(n14182) );
  XOR U14242 ( .A(n14079), .B(n14191), .Z(n14183) );
  XNOR U14243 ( .A(n14078), .B(n14076), .Z(n14191) );
  AND U14244 ( .A(n14192), .B(n14193), .Z(n14076) );
  NANDN U14245 ( .A(n14194), .B(n14195), .Z(n14193) );
  OR U14246 ( .A(n14196), .B(n14197), .Z(n14195) );
  NAND U14247 ( .A(n14197), .B(n14196), .Z(n14192) );
  ANDN U14248 ( .B(B[240]), .A(n55), .Z(n14078) );
  XNOR U14249 ( .A(n14086), .B(n14198), .Z(n14079) );
  XNOR U14250 ( .A(n14085), .B(n14083), .Z(n14198) );
  AND U14251 ( .A(n14199), .B(n14200), .Z(n14083) );
  NANDN U14252 ( .A(n14201), .B(n14202), .Z(n14200) );
  NANDN U14253 ( .A(n14203), .B(n14204), .Z(n14202) );
  NANDN U14254 ( .A(n14204), .B(n14203), .Z(n14199) );
  ANDN U14255 ( .B(B[241]), .A(n56), .Z(n14085) );
  XNOR U14256 ( .A(n14093), .B(n14205), .Z(n14086) );
  XNOR U14257 ( .A(n14092), .B(n14090), .Z(n14205) );
  AND U14258 ( .A(n14206), .B(n14207), .Z(n14090) );
  NANDN U14259 ( .A(n14208), .B(n14209), .Z(n14207) );
  OR U14260 ( .A(n14210), .B(n14211), .Z(n14209) );
  NAND U14261 ( .A(n14211), .B(n14210), .Z(n14206) );
  ANDN U14262 ( .B(B[242]), .A(n57), .Z(n14092) );
  XNOR U14263 ( .A(n14100), .B(n14212), .Z(n14093) );
  XNOR U14264 ( .A(n14099), .B(n14097), .Z(n14212) );
  AND U14265 ( .A(n14213), .B(n14214), .Z(n14097) );
  NANDN U14266 ( .A(n14215), .B(n14216), .Z(n14214) );
  NANDN U14267 ( .A(n14217), .B(n14218), .Z(n14216) );
  NANDN U14268 ( .A(n14218), .B(n14217), .Z(n14213) );
  ANDN U14269 ( .B(B[243]), .A(n58), .Z(n14099) );
  XNOR U14270 ( .A(n14107), .B(n14219), .Z(n14100) );
  XNOR U14271 ( .A(n14106), .B(n14104), .Z(n14219) );
  AND U14272 ( .A(n14220), .B(n14221), .Z(n14104) );
  NANDN U14273 ( .A(n14222), .B(n14223), .Z(n14221) );
  OR U14274 ( .A(n14224), .B(n14225), .Z(n14223) );
  NAND U14275 ( .A(n14225), .B(n14224), .Z(n14220) );
  ANDN U14276 ( .B(B[244]), .A(n59), .Z(n14106) );
  XNOR U14277 ( .A(n14114), .B(n14226), .Z(n14107) );
  XNOR U14278 ( .A(n14113), .B(n14111), .Z(n14226) );
  AND U14279 ( .A(n14227), .B(n14228), .Z(n14111) );
  NANDN U14280 ( .A(n14229), .B(n14230), .Z(n14228) );
  NANDN U14281 ( .A(n14231), .B(n14232), .Z(n14230) );
  NANDN U14282 ( .A(n14232), .B(n14231), .Z(n14227) );
  ANDN U14283 ( .B(B[245]), .A(n60), .Z(n14113) );
  XNOR U14284 ( .A(n14121), .B(n14233), .Z(n14114) );
  XNOR U14285 ( .A(n14120), .B(n14118), .Z(n14233) );
  AND U14286 ( .A(n14234), .B(n14235), .Z(n14118) );
  NANDN U14287 ( .A(n14236), .B(n14237), .Z(n14235) );
  OR U14288 ( .A(n14238), .B(n14239), .Z(n14237) );
  NAND U14289 ( .A(n14239), .B(n14238), .Z(n14234) );
  ANDN U14290 ( .B(B[246]), .A(n61), .Z(n14120) );
  XNOR U14291 ( .A(n14128), .B(n14240), .Z(n14121) );
  XNOR U14292 ( .A(n14127), .B(n14125), .Z(n14240) );
  AND U14293 ( .A(n14241), .B(n14242), .Z(n14125) );
  NANDN U14294 ( .A(n14243), .B(n14244), .Z(n14242) );
  NANDN U14295 ( .A(n14245), .B(n14246), .Z(n14244) );
  NANDN U14296 ( .A(n14246), .B(n14245), .Z(n14241) );
  ANDN U14297 ( .B(B[247]), .A(n62), .Z(n14127) );
  XNOR U14298 ( .A(n14135), .B(n14247), .Z(n14128) );
  XNOR U14299 ( .A(n14134), .B(n14132), .Z(n14247) );
  AND U14300 ( .A(n14248), .B(n14249), .Z(n14132) );
  NANDN U14301 ( .A(n14250), .B(n14251), .Z(n14249) );
  OR U14302 ( .A(n14252), .B(n14253), .Z(n14251) );
  NAND U14303 ( .A(n14253), .B(n14252), .Z(n14248) );
  ANDN U14304 ( .B(B[248]), .A(n63), .Z(n14134) );
  XNOR U14305 ( .A(n14142), .B(n14254), .Z(n14135) );
  XNOR U14306 ( .A(n14141), .B(n14139), .Z(n14254) );
  AND U14307 ( .A(n14255), .B(n14256), .Z(n14139) );
  NANDN U14308 ( .A(n14257), .B(n14258), .Z(n14256) );
  NANDN U14309 ( .A(n14259), .B(n14260), .Z(n14258) );
  NANDN U14310 ( .A(n14260), .B(n14259), .Z(n14255) );
  ANDN U14311 ( .B(B[249]), .A(n64), .Z(n14141) );
  XNOR U14312 ( .A(n14149), .B(n14261), .Z(n14142) );
  XNOR U14313 ( .A(n14148), .B(n14146), .Z(n14261) );
  AND U14314 ( .A(n14262), .B(n14263), .Z(n14146) );
  NANDN U14315 ( .A(n14264), .B(n14265), .Z(n14263) );
  OR U14316 ( .A(n14266), .B(n14267), .Z(n14265) );
  NAND U14317 ( .A(n14267), .B(n14266), .Z(n14262) );
  ANDN U14318 ( .B(B[250]), .A(n65), .Z(n14148) );
  XNOR U14319 ( .A(n14156), .B(n14268), .Z(n14149) );
  XNOR U14320 ( .A(n14155), .B(n14153), .Z(n14268) );
  AND U14321 ( .A(n14269), .B(n14270), .Z(n14153) );
  NANDN U14322 ( .A(n14271), .B(n14272), .Z(n14270) );
  NANDN U14323 ( .A(n14273), .B(n14274), .Z(n14272) );
  NANDN U14324 ( .A(n14274), .B(n14273), .Z(n14269) );
  ANDN U14325 ( .B(B[251]), .A(n66), .Z(n14155) );
  XNOR U14326 ( .A(n14163), .B(n14275), .Z(n14156) );
  XNOR U14327 ( .A(n14162), .B(n14160), .Z(n14275) );
  AND U14328 ( .A(n14276), .B(n14277), .Z(n14160) );
  NANDN U14329 ( .A(n14278), .B(n14279), .Z(n14277) );
  OR U14330 ( .A(n14280), .B(n14281), .Z(n14279) );
  NAND U14331 ( .A(n14281), .B(n14280), .Z(n14276) );
  ANDN U14332 ( .B(B[252]), .A(n67), .Z(n14162) );
  XNOR U14333 ( .A(n14170), .B(n14282), .Z(n14163) );
  XNOR U14334 ( .A(n14169), .B(n14167), .Z(n14282) );
  AND U14335 ( .A(n14283), .B(n14284), .Z(n14167) );
  NANDN U14336 ( .A(n14285), .B(n14286), .Z(n14284) );
  NANDN U14337 ( .A(n14287), .B(n14288), .Z(n14286) );
  NANDN U14338 ( .A(n14288), .B(n14287), .Z(n14283) );
  ANDN U14339 ( .B(B[253]), .A(n68), .Z(n14169) );
  XOR U14340 ( .A(n14175), .B(n14289), .Z(n14170) );
  XOR U14341 ( .A(n14176), .B(n14177), .Z(n14289) );
  NAND U14342 ( .A(A[15]), .B(B[255]), .Z(n14177) );
  AND U14343 ( .A(B[254]), .B(A[16]), .Z(n14176) );
  NAND U14344 ( .A(n14290), .B(n14291), .Z(n14175) );
  NAND U14345 ( .A(n14292), .B(n14293), .Z(n14291) );
  NANDN U14346 ( .A(n14294), .B(n14295), .Z(n14292) );
  NANDN U14347 ( .A(n14295), .B(n14294), .Z(n14290) );
  NAND U14348 ( .A(n14296), .B(n14297), .Z(n256) );
  NANDN U14349 ( .A(n14298), .B(n14299), .Z(n14297) );
  OR U14350 ( .A(n14300), .B(n14301), .Z(n14299) );
  NAND U14351 ( .A(n14301), .B(n14300), .Z(n14296) );
  XOR U14352 ( .A(n258), .B(n257), .Z(\A1[267] ) );
  XOR U14353 ( .A(n14301), .B(n14302), .Z(n257) );
  XNOR U14354 ( .A(n14300), .B(n14298), .Z(n14302) );
  AND U14355 ( .A(n14303), .B(n14304), .Z(n14298) );
  NANDN U14356 ( .A(n14305), .B(n14306), .Z(n14304) );
  OR U14357 ( .A(n14307), .B(n14308), .Z(n14306) );
  NAND U14358 ( .A(n14308), .B(n14307), .Z(n14303) );
  ANDN U14359 ( .B(B[238]), .A(n54), .Z(n14300) );
  XNOR U14360 ( .A(n14190), .B(n14309), .Z(n14301) );
  XNOR U14361 ( .A(n14189), .B(n14187), .Z(n14309) );
  AND U14362 ( .A(n14310), .B(n14311), .Z(n14187) );
  NANDN U14363 ( .A(n14312), .B(n14313), .Z(n14311) );
  NANDN U14364 ( .A(n14314), .B(n14315), .Z(n14313) );
  NANDN U14365 ( .A(n14315), .B(n14314), .Z(n14310) );
  ANDN U14366 ( .B(B[239]), .A(n55), .Z(n14189) );
  XNOR U14367 ( .A(n14197), .B(n14316), .Z(n14190) );
  XNOR U14368 ( .A(n14196), .B(n14194), .Z(n14316) );
  AND U14369 ( .A(n14317), .B(n14318), .Z(n14194) );
  NANDN U14370 ( .A(n14319), .B(n14320), .Z(n14318) );
  OR U14371 ( .A(n14321), .B(n14322), .Z(n14320) );
  NAND U14372 ( .A(n14322), .B(n14321), .Z(n14317) );
  ANDN U14373 ( .B(B[240]), .A(n56), .Z(n14196) );
  XNOR U14374 ( .A(n14204), .B(n14323), .Z(n14197) );
  XNOR U14375 ( .A(n14203), .B(n14201), .Z(n14323) );
  AND U14376 ( .A(n14324), .B(n14325), .Z(n14201) );
  NANDN U14377 ( .A(n14326), .B(n14327), .Z(n14325) );
  NANDN U14378 ( .A(n14328), .B(n14329), .Z(n14327) );
  NANDN U14379 ( .A(n14329), .B(n14328), .Z(n14324) );
  ANDN U14380 ( .B(B[241]), .A(n57), .Z(n14203) );
  XNOR U14381 ( .A(n14211), .B(n14330), .Z(n14204) );
  XNOR U14382 ( .A(n14210), .B(n14208), .Z(n14330) );
  AND U14383 ( .A(n14331), .B(n14332), .Z(n14208) );
  NANDN U14384 ( .A(n14333), .B(n14334), .Z(n14332) );
  OR U14385 ( .A(n14335), .B(n14336), .Z(n14334) );
  NAND U14386 ( .A(n14336), .B(n14335), .Z(n14331) );
  ANDN U14387 ( .B(B[242]), .A(n58), .Z(n14210) );
  XNOR U14388 ( .A(n14218), .B(n14337), .Z(n14211) );
  XNOR U14389 ( .A(n14217), .B(n14215), .Z(n14337) );
  AND U14390 ( .A(n14338), .B(n14339), .Z(n14215) );
  NANDN U14391 ( .A(n14340), .B(n14341), .Z(n14339) );
  NANDN U14392 ( .A(n14342), .B(n14343), .Z(n14341) );
  NANDN U14393 ( .A(n14343), .B(n14342), .Z(n14338) );
  ANDN U14394 ( .B(B[243]), .A(n59), .Z(n14217) );
  XNOR U14395 ( .A(n14225), .B(n14344), .Z(n14218) );
  XNOR U14396 ( .A(n14224), .B(n14222), .Z(n14344) );
  AND U14397 ( .A(n14345), .B(n14346), .Z(n14222) );
  NANDN U14398 ( .A(n14347), .B(n14348), .Z(n14346) );
  OR U14399 ( .A(n14349), .B(n14350), .Z(n14348) );
  NAND U14400 ( .A(n14350), .B(n14349), .Z(n14345) );
  ANDN U14401 ( .B(B[244]), .A(n60), .Z(n14224) );
  XNOR U14402 ( .A(n14232), .B(n14351), .Z(n14225) );
  XNOR U14403 ( .A(n14231), .B(n14229), .Z(n14351) );
  AND U14404 ( .A(n14352), .B(n14353), .Z(n14229) );
  NANDN U14405 ( .A(n14354), .B(n14355), .Z(n14353) );
  NANDN U14406 ( .A(n14356), .B(n14357), .Z(n14355) );
  NANDN U14407 ( .A(n14357), .B(n14356), .Z(n14352) );
  ANDN U14408 ( .B(B[245]), .A(n61), .Z(n14231) );
  XNOR U14409 ( .A(n14239), .B(n14358), .Z(n14232) );
  XNOR U14410 ( .A(n14238), .B(n14236), .Z(n14358) );
  AND U14411 ( .A(n14359), .B(n14360), .Z(n14236) );
  NANDN U14412 ( .A(n14361), .B(n14362), .Z(n14360) );
  OR U14413 ( .A(n14363), .B(n14364), .Z(n14362) );
  NAND U14414 ( .A(n14364), .B(n14363), .Z(n14359) );
  ANDN U14415 ( .B(B[246]), .A(n62), .Z(n14238) );
  XNOR U14416 ( .A(n14246), .B(n14365), .Z(n14239) );
  XNOR U14417 ( .A(n14245), .B(n14243), .Z(n14365) );
  AND U14418 ( .A(n14366), .B(n14367), .Z(n14243) );
  NANDN U14419 ( .A(n14368), .B(n14369), .Z(n14367) );
  NANDN U14420 ( .A(n14370), .B(n14371), .Z(n14369) );
  NANDN U14421 ( .A(n14371), .B(n14370), .Z(n14366) );
  ANDN U14422 ( .B(B[247]), .A(n63), .Z(n14245) );
  XNOR U14423 ( .A(n14253), .B(n14372), .Z(n14246) );
  XNOR U14424 ( .A(n14252), .B(n14250), .Z(n14372) );
  AND U14425 ( .A(n14373), .B(n14374), .Z(n14250) );
  NANDN U14426 ( .A(n14375), .B(n14376), .Z(n14374) );
  OR U14427 ( .A(n14377), .B(n14378), .Z(n14376) );
  NAND U14428 ( .A(n14378), .B(n14377), .Z(n14373) );
  ANDN U14429 ( .B(B[248]), .A(n64), .Z(n14252) );
  XNOR U14430 ( .A(n14260), .B(n14379), .Z(n14253) );
  XNOR U14431 ( .A(n14259), .B(n14257), .Z(n14379) );
  AND U14432 ( .A(n14380), .B(n14381), .Z(n14257) );
  NANDN U14433 ( .A(n14382), .B(n14383), .Z(n14381) );
  NANDN U14434 ( .A(n14384), .B(n14385), .Z(n14383) );
  NANDN U14435 ( .A(n14385), .B(n14384), .Z(n14380) );
  ANDN U14436 ( .B(B[249]), .A(n65), .Z(n14259) );
  XNOR U14437 ( .A(n14267), .B(n14386), .Z(n14260) );
  XNOR U14438 ( .A(n14266), .B(n14264), .Z(n14386) );
  AND U14439 ( .A(n14387), .B(n14388), .Z(n14264) );
  NANDN U14440 ( .A(n14389), .B(n14390), .Z(n14388) );
  OR U14441 ( .A(n14391), .B(n14392), .Z(n14390) );
  NAND U14442 ( .A(n14392), .B(n14391), .Z(n14387) );
  ANDN U14443 ( .B(B[250]), .A(n66), .Z(n14266) );
  XNOR U14444 ( .A(n14274), .B(n14393), .Z(n14267) );
  XNOR U14445 ( .A(n14273), .B(n14271), .Z(n14393) );
  AND U14446 ( .A(n14394), .B(n14395), .Z(n14271) );
  NANDN U14447 ( .A(n14396), .B(n14397), .Z(n14395) );
  NANDN U14448 ( .A(n14398), .B(n14399), .Z(n14397) );
  NANDN U14449 ( .A(n14399), .B(n14398), .Z(n14394) );
  ANDN U14450 ( .B(B[251]), .A(n67), .Z(n14273) );
  XNOR U14451 ( .A(n14281), .B(n14400), .Z(n14274) );
  XNOR U14452 ( .A(n14280), .B(n14278), .Z(n14400) );
  AND U14453 ( .A(n14401), .B(n14402), .Z(n14278) );
  NANDN U14454 ( .A(n14403), .B(n14404), .Z(n14402) );
  OR U14455 ( .A(n14405), .B(n14406), .Z(n14404) );
  NAND U14456 ( .A(n14406), .B(n14405), .Z(n14401) );
  ANDN U14457 ( .B(B[252]), .A(n68), .Z(n14280) );
  XNOR U14458 ( .A(n14288), .B(n14407), .Z(n14281) );
  XNOR U14459 ( .A(n14287), .B(n14285), .Z(n14407) );
  AND U14460 ( .A(n14408), .B(n14409), .Z(n14285) );
  NANDN U14461 ( .A(n14410), .B(n14411), .Z(n14409) );
  NANDN U14462 ( .A(n14412), .B(n14413), .Z(n14411) );
  NANDN U14463 ( .A(n14413), .B(n14412), .Z(n14408) );
  ANDN U14464 ( .B(B[253]), .A(n69), .Z(n14287) );
  XOR U14465 ( .A(n14293), .B(n14414), .Z(n14288) );
  XOR U14466 ( .A(n14294), .B(n14295), .Z(n14414) );
  NAND U14467 ( .A(A[14]), .B(B[255]), .Z(n14295) );
  AND U14468 ( .A(B[254]), .B(A[15]), .Z(n14294) );
  NAND U14469 ( .A(n14415), .B(n14416), .Z(n14293) );
  NAND U14470 ( .A(n14417), .B(n14418), .Z(n14416) );
  NANDN U14471 ( .A(n14419), .B(n14420), .Z(n14417) );
  NANDN U14472 ( .A(n14420), .B(n14419), .Z(n14415) );
  NAND U14473 ( .A(n14421), .B(n14422), .Z(n258) );
  NANDN U14474 ( .A(n14423), .B(n14424), .Z(n14422) );
  NAND U14475 ( .A(n14426), .B(n14425), .Z(n14421) );
  XOR U14476 ( .A(n260), .B(n259), .Z(\A1[266] ) );
  XOR U14477 ( .A(n14426), .B(n14427), .Z(n259) );
  XNOR U14478 ( .A(n14425), .B(n14423), .Z(n14427) );
  AND U14479 ( .A(n14428), .B(n14429), .Z(n14423) );
  NANDN U14480 ( .A(n14430), .B(n14431), .Z(n14429) );
  NANDN U14481 ( .A(n14432), .B(n14433), .Z(n14431) );
  NANDN U14482 ( .A(n14433), .B(n14432), .Z(n14428) );
  ANDN U14483 ( .B(B[237]), .A(n54), .Z(n14425) );
  XOR U14484 ( .A(n14308), .B(n14434), .Z(n14426) );
  XNOR U14485 ( .A(n14307), .B(n14305), .Z(n14434) );
  AND U14486 ( .A(n14435), .B(n14436), .Z(n14305) );
  NANDN U14487 ( .A(n14437), .B(n14438), .Z(n14436) );
  OR U14488 ( .A(n14439), .B(n14440), .Z(n14438) );
  NAND U14489 ( .A(n14440), .B(n14439), .Z(n14435) );
  ANDN U14490 ( .B(B[238]), .A(n55), .Z(n14307) );
  XNOR U14491 ( .A(n14315), .B(n14441), .Z(n14308) );
  XNOR U14492 ( .A(n14314), .B(n14312), .Z(n14441) );
  AND U14493 ( .A(n14442), .B(n14443), .Z(n14312) );
  NANDN U14494 ( .A(n14444), .B(n14445), .Z(n14443) );
  NANDN U14495 ( .A(n14446), .B(n14447), .Z(n14445) );
  NANDN U14496 ( .A(n14447), .B(n14446), .Z(n14442) );
  ANDN U14497 ( .B(B[239]), .A(n56), .Z(n14314) );
  XNOR U14498 ( .A(n14322), .B(n14448), .Z(n14315) );
  XNOR U14499 ( .A(n14321), .B(n14319), .Z(n14448) );
  AND U14500 ( .A(n14449), .B(n14450), .Z(n14319) );
  NANDN U14501 ( .A(n14451), .B(n14452), .Z(n14450) );
  OR U14502 ( .A(n14453), .B(n14454), .Z(n14452) );
  NAND U14503 ( .A(n14454), .B(n14453), .Z(n14449) );
  ANDN U14504 ( .B(B[240]), .A(n57), .Z(n14321) );
  XNOR U14505 ( .A(n14329), .B(n14455), .Z(n14322) );
  XNOR U14506 ( .A(n14328), .B(n14326), .Z(n14455) );
  AND U14507 ( .A(n14456), .B(n14457), .Z(n14326) );
  NANDN U14508 ( .A(n14458), .B(n14459), .Z(n14457) );
  NANDN U14509 ( .A(n14460), .B(n14461), .Z(n14459) );
  NANDN U14510 ( .A(n14461), .B(n14460), .Z(n14456) );
  ANDN U14511 ( .B(B[241]), .A(n58), .Z(n14328) );
  XNOR U14512 ( .A(n14336), .B(n14462), .Z(n14329) );
  XNOR U14513 ( .A(n14335), .B(n14333), .Z(n14462) );
  AND U14514 ( .A(n14463), .B(n14464), .Z(n14333) );
  NANDN U14515 ( .A(n14465), .B(n14466), .Z(n14464) );
  OR U14516 ( .A(n14467), .B(n14468), .Z(n14466) );
  NAND U14517 ( .A(n14468), .B(n14467), .Z(n14463) );
  ANDN U14518 ( .B(B[242]), .A(n59), .Z(n14335) );
  XNOR U14519 ( .A(n14343), .B(n14469), .Z(n14336) );
  XNOR U14520 ( .A(n14342), .B(n14340), .Z(n14469) );
  AND U14521 ( .A(n14470), .B(n14471), .Z(n14340) );
  NANDN U14522 ( .A(n14472), .B(n14473), .Z(n14471) );
  NANDN U14523 ( .A(n14474), .B(n14475), .Z(n14473) );
  NANDN U14524 ( .A(n14475), .B(n14474), .Z(n14470) );
  ANDN U14525 ( .B(B[243]), .A(n60), .Z(n14342) );
  XNOR U14526 ( .A(n14350), .B(n14476), .Z(n14343) );
  XNOR U14527 ( .A(n14349), .B(n14347), .Z(n14476) );
  AND U14528 ( .A(n14477), .B(n14478), .Z(n14347) );
  NANDN U14529 ( .A(n14479), .B(n14480), .Z(n14478) );
  OR U14530 ( .A(n14481), .B(n14482), .Z(n14480) );
  NAND U14531 ( .A(n14482), .B(n14481), .Z(n14477) );
  ANDN U14532 ( .B(B[244]), .A(n61), .Z(n14349) );
  XNOR U14533 ( .A(n14357), .B(n14483), .Z(n14350) );
  XNOR U14534 ( .A(n14356), .B(n14354), .Z(n14483) );
  AND U14535 ( .A(n14484), .B(n14485), .Z(n14354) );
  NANDN U14536 ( .A(n14486), .B(n14487), .Z(n14485) );
  NANDN U14537 ( .A(n14488), .B(n14489), .Z(n14487) );
  NANDN U14538 ( .A(n14489), .B(n14488), .Z(n14484) );
  ANDN U14539 ( .B(B[245]), .A(n62), .Z(n14356) );
  XNOR U14540 ( .A(n14364), .B(n14490), .Z(n14357) );
  XNOR U14541 ( .A(n14363), .B(n14361), .Z(n14490) );
  AND U14542 ( .A(n14491), .B(n14492), .Z(n14361) );
  NANDN U14543 ( .A(n14493), .B(n14494), .Z(n14492) );
  OR U14544 ( .A(n14495), .B(n14496), .Z(n14494) );
  NAND U14545 ( .A(n14496), .B(n14495), .Z(n14491) );
  ANDN U14546 ( .B(B[246]), .A(n63), .Z(n14363) );
  XNOR U14547 ( .A(n14371), .B(n14497), .Z(n14364) );
  XNOR U14548 ( .A(n14370), .B(n14368), .Z(n14497) );
  AND U14549 ( .A(n14498), .B(n14499), .Z(n14368) );
  NANDN U14550 ( .A(n14500), .B(n14501), .Z(n14499) );
  NANDN U14551 ( .A(n14502), .B(n14503), .Z(n14501) );
  NANDN U14552 ( .A(n14503), .B(n14502), .Z(n14498) );
  ANDN U14553 ( .B(B[247]), .A(n64), .Z(n14370) );
  XNOR U14554 ( .A(n14378), .B(n14504), .Z(n14371) );
  XNOR U14555 ( .A(n14377), .B(n14375), .Z(n14504) );
  AND U14556 ( .A(n14505), .B(n14506), .Z(n14375) );
  NANDN U14557 ( .A(n14507), .B(n14508), .Z(n14506) );
  OR U14558 ( .A(n14509), .B(n14510), .Z(n14508) );
  NAND U14559 ( .A(n14510), .B(n14509), .Z(n14505) );
  ANDN U14560 ( .B(B[248]), .A(n65), .Z(n14377) );
  XNOR U14561 ( .A(n14385), .B(n14511), .Z(n14378) );
  XNOR U14562 ( .A(n14384), .B(n14382), .Z(n14511) );
  AND U14563 ( .A(n14512), .B(n14513), .Z(n14382) );
  NANDN U14564 ( .A(n14514), .B(n14515), .Z(n14513) );
  NANDN U14565 ( .A(n14516), .B(n14517), .Z(n14515) );
  NANDN U14566 ( .A(n14517), .B(n14516), .Z(n14512) );
  ANDN U14567 ( .B(B[249]), .A(n66), .Z(n14384) );
  XNOR U14568 ( .A(n14392), .B(n14518), .Z(n14385) );
  XNOR U14569 ( .A(n14391), .B(n14389), .Z(n14518) );
  AND U14570 ( .A(n14519), .B(n14520), .Z(n14389) );
  NANDN U14571 ( .A(n14521), .B(n14522), .Z(n14520) );
  OR U14572 ( .A(n14523), .B(n14524), .Z(n14522) );
  NAND U14573 ( .A(n14524), .B(n14523), .Z(n14519) );
  ANDN U14574 ( .B(B[250]), .A(n67), .Z(n14391) );
  XNOR U14575 ( .A(n14399), .B(n14525), .Z(n14392) );
  XNOR U14576 ( .A(n14398), .B(n14396), .Z(n14525) );
  AND U14577 ( .A(n14526), .B(n14527), .Z(n14396) );
  NANDN U14578 ( .A(n14528), .B(n14529), .Z(n14527) );
  NANDN U14579 ( .A(n14530), .B(n14531), .Z(n14529) );
  NANDN U14580 ( .A(n14531), .B(n14530), .Z(n14526) );
  ANDN U14581 ( .B(B[251]), .A(n68), .Z(n14398) );
  XNOR U14582 ( .A(n14406), .B(n14532), .Z(n14399) );
  XNOR U14583 ( .A(n14405), .B(n14403), .Z(n14532) );
  AND U14584 ( .A(n14533), .B(n14534), .Z(n14403) );
  NANDN U14585 ( .A(n14535), .B(n14536), .Z(n14534) );
  OR U14586 ( .A(n14537), .B(n14538), .Z(n14536) );
  NAND U14587 ( .A(n14538), .B(n14537), .Z(n14533) );
  ANDN U14588 ( .B(B[252]), .A(n69), .Z(n14405) );
  XNOR U14589 ( .A(n14413), .B(n14539), .Z(n14406) );
  XNOR U14590 ( .A(n14412), .B(n14410), .Z(n14539) );
  AND U14591 ( .A(n14540), .B(n14541), .Z(n14410) );
  NANDN U14592 ( .A(n14542), .B(n14543), .Z(n14541) );
  NANDN U14593 ( .A(n14544), .B(n14545), .Z(n14543) );
  NANDN U14594 ( .A(n14545), .B(n14544), .Z(n14540) );
  ANDN U14595 ( .B(B[253]), .A(n70), .Z(n14412) );
  XOR U14596 ( .A(n14418), .B(n14546), .Z(n14413) );
  XOR U14597 ( .A(n14419), .B(n14420), .Z(n14546) );
  NAND U14598 ( .A(A[13]), .B(B[255]), .Z(n14420) );
  AND U14599 ( .A(B[254]), .B(A[14]), .Z(n14419) );
  NAND U14600 ( .A(n14547), .B(n14548), .Z(n14418) );
  NAND U14601 ( .A(n14549), .B(n14550), .Z(n14548) );
  NANDN U14602 ( .A(n14551), .B(n14552), .Z(n14549) );
  NANDN U14603 ( .A(n14552), .B(n14551), .Z(n14547) );
  NAND U14604 ( .A(n14553), .B(n14554), .Z(n260) );
  NANDN U14605 ( .A(n14555), .B(n14556), .Z(n14554) );
  OR U14606 ( .A(n14557), .B(n14558), .Z(n14556) );
  NAND U14607 ( .A(n14558), .B(n14557), .Z(n14553) );
  XOR U14608 ( .A(n262), .B(n261), .Z(\A1[265] ) );
  XOR U14609 ( .A(n14558), .B(n14559), .Z(n261) );
  XNOR U14610 ( .A(n14557), .B(n14555), .Z(n14559) );
  AND U14611 ( .A(n14560), .B(n14561), .Z(n14555) );
  NANDN U14612 ( .A(n14562), .B(n14563), .Z(n14561) );
  OR U14613 ( .A(n14564), .B(n14565), .Z(n14563) );
  NAND U14614 ( .A(n14565), .B(n14564), .Z(n14560) );
  ANDN U14615 ( .B(B[236]), .A(n54), .Z(n14557) );
  XNOR U14616 ( .A(n14433), .B(n14566), .Z(n14558) );
  XNOR U14617 ( .A(n14432), .B(n14430), .Z(n14566) );
  AND U14618 ( .A(n14567), .B(n14568), .Z(n14430) );
  NANDN U14619 ( .A(n14569), .B(n14570), .Z(n14568) );
  NANDN U14620 ( .A(n14571), .B(n14572), .Z(n14570) );
  NANDN U14621 ( .A(n14572), .B(n14571), .Z(n14567) );
  ANDN U14622 ( .B(B[237]), .A(n55), .Z(n14432) );
  XNOR U14623 ( .A(n14440), .B(n14573), .Z(n14433) );
  XNOR U14624 ( .A(n14439), .B(n14437), .Z(n14573) );
  AND U14625 ( .A(n14574), .B(n14575), .Z(n14437) );
  NANDN U14626 ( .A(n14576), .B(n14577), .Z(n14575) );
  OR U14627 ( .A(n14578), .B(n14579), .Z(n14577) );
  NAND U14628 ( .A(n14579), .B(n14578), .Z(n14574) );
  ANDN U14629 ( .B(B[238]), .A(n56), .Z(n14439) );
  XNOR U14630 ( .A(n14447), .B(n14580), .Z(n14440) );
  XNOR U14631 ( .A(n14446), .B(n14444), .Z(n14580) );
  AND U14632 ( .A(n14581), .B(n14582), .Z(n14444) );
  NANDN U14633 ( .A(n14583), .B(n14584), .Z(n14582) );
  NANDN U14634 ( .A(n14585), .B(n14586), .Z(n14584) );
  NANDN U14635 ( .A(n14586), .B(n14585), .Z(n14581) );
  ANDN U14636 ( .B(B[239]), .A(n57), .Z(n14446) );
  XNOR U14637 ( .A(n14454), .B(n14587), .Z(n14447) );
  XNOR U14638 ( .A(n14453), .B(n14451), .Z(n14587) );
  AND U14639 ( .A(n14588), .B(n14589), .Z(n14451) );
  NANDN U14640 ( .A(n14590), .B(n14591), .Z(n14589) );
  OR U14641 ( .A(n14592), .B(n14593), .Z(n14591) );
  NAND U14642 ( .A(n14593), .B(n14592), .Z(n14588) );
  ANDN U14643 ( .B(B[240]), .A(n58), .Z(n14453) );
  XNOR U14644 ( .A(n14461), .B(n14594), .Z(n14454) );
  XNOR U14645 ( .A(n14460), .B(n14458), .Z(n14594) );
  AND U14646 ( .A(n14595), .B(n14596), .Z(n14458) );
  NANDN U14647 ( .A(n14597), .B(n14598), .Z(n14596) );
  NANDN U14648 ( .A(n14599), .B(n14600), .Z(n14598) );
  NANDN U14649 ( .A(n14600), .B(n14599), .Z(n14595) );
  ANDN U14650 ( .B(B[241]), .A(n59), .Z(n14460) );
  XNOR U14651 ( .A(n14468), .B(n14601), .Z(n14461) );
  XNOR U14652 ( .A(n14467), .B(n14465), .Z(n14601) );
  AND U14653 ( .A(n14602), .B(n14603), .Z(n14465) );
  NANDN U14654 ( .A(n14604), .B(n14605), .Z(n14603) );
  OR U14655 ( .A(n14606), .B(n14607), .Z(n14605) );
  NAND U14656 ( .A(n14607), .B(n14606), .Z(n14602) );
  ANDN U14657 ( .B(B[242]), .A(n60), .Z(n14467) );
  XNOR U14658 ( .A(n14475), .B(n14608), .Z(n14468) );
  XNOR U14659 ( .A(n14474), .B(n14472), .Z(n14608) );
  AND U14660 ( .A(n14609), .B(n14610), .Z(n14472) );
  NANDN U14661 ( .A(n14611), .B(n14612), .Z(n14610) );
  NANDN U14662 ( .A(n14613), .B(n14614), .Z(n14612) );
  NANDN U14663 ( .A(n14614), .B(n14613), .Z(n14609) );
  ANDN U14664 ( .B(B[243]), .A(n61), .Z(n14474) );
  XNOR U14665 ( .A(n14482), .B(n14615), .Z(n14475) );
  XNOR U14666 ( .A(n14481), .B(n14479), .Z(n14615) );
  AND U14667 ( .A(n14616), .B(n14617), .Z(n14479) );
  NANDN U14668 ( .A(n14618), .B(n14619), .Z(n14617) );
  OR U14669 ( .A(n14620), .B(n14621), .Z(n14619) );
  NAND U14670 ( .A(n14621), .B(n14620), .Z(n14616) );
  ANDN U14671 ( .B(B[244]), .A(n62), .Z(n14481) );
  XNOR U14672 ( .A(n14489), .B(n14622), .Z(n14482) );
  XNOR U14673 ( .A(n14488), .B(n14486), .Z(n14622) );
  AND U14674 ( .A(n14623), .B(n14624), .Z(n14486) );
  NANDN U14675 ( .A(n14625), .B(n14626), .Z(n14624) );
  NANDN U14676 ( .A(n14627), .B(n14628), .Z(n14626) );
  NANDN U14677 ( .A(n14628), .B(n14627), .Z(n14623) );
  ANDN U14678 ( .B(B[245]), .A(n63), .Z(n14488) );
  XNOR U14679 ( .A(n14496), .B(n14629), .Z(n14489) );
  XNOR U14680 ( .A(n14495), .B(n14493), .Z(n14629) );
  AND U14681 ( .A(n14630), .B(n14631), .Z(n14493) );
  NANDN U14682 ( .A(n14632), .B(n14633), .Z(n14631) );
  OR U14683 ( .A(n14634), .B(n14635), .Z(n14633) );
  NAND U14684 ( .A(n14635), .B(n14634), .Z(n14630) );
  ANDN U14685 ( .B(B[246]), .A(n64), .Z(n14495) );
  XNOR U14686 ( .A(n14503), .B(n14636), .Z(n14496) );
  XNOR U14687 ( .A(n14502), .B(n14500), .Z(n14636) );
  AND U14688 ( .A(n14637), .B(n14638), .Z(n14500) );
  NANDN U14689 ( .A(n14639), .B(n14640), .Z(n14638) );
  NANDN U14690 ( .A(n14641), .B(n14642), .Z(n14640) );
  NANDN U14691 ( .A(n14642), .B(n14641), .Z(n14637) );
  ANDN U14692 ( .B(B[247]), .A(n65), .Z(n14502) );
  XNOR U14693 ( .A(n14510), .B(n14643), .Z(n14503) );
  XNOR U14694 ( .A(n14509), .B(n14507), .Z(n14643) );
  AND U14695 ( .A(n14644), .B(n14645), .Z(n14507) );
  NANDN U14696 ( .A(n14646), .B(n14647), .Z(n14645) );
  OR U14697 ( .A(n14648), .B(n14649), .Z(n14647) );
  NAND U14698 ( .A(n14649), .B(n14648), .Z(n14644) );
  ANDN U14699 ( .B(B[248]), .A(n66), .Z(n14509) );
  XNOR U14700 ( .A(n14517), .B(n14650), .Z(n14510) );
  XNOR U14701 ( .A(n14516), .B(n14514), .Z(n14650) );
  AND U14702 ( .A(n14651), .B(n14652), .Z(n14514) );
  NANDN U14703 ( .A(n14653), .B(n14654), .Z(n14652) );
  NANDN U14704 ( .A(n14655), .B(n14656), .Z(n14654) );
  NANDN U14705 ( .A(n14656), .B(n14655), .Z(n14651) );
  ANDN U14706 ( .B(B[249]), .A(n67), .Z(n14516) );
  XNOR U14707 ( .A(n14524), .B(n14657), .Z(n14517) );
  XNOR U14708 ( .A(n14523), .B(n14521), .Z(n14657) );
  AND U14709 ( .A(n14658), .B(n14659), .Z(n14521) );
  NANDN U14710 ( .A(n14660), .B(n14661), .Z(n14659) );
  OR U14711 ( .A(n14662), .B(n14663), .Z(n14661) );
  NAND U14712 ( .A(n14663), .B(n14662), .Z(n14658) );
  ANDN U14713 ( .B(B[250]), .A(n68), .Z(n14523) );
  XNOR U14714 ( .A(n14531), .B(n14664), .Z(n14524) );
  XNOR U14715 ( .A(n14530), .B(n14528), .Z(n14664) );
  AND U14716 ( .A(n14665), .B(n14666), .Z(n14528) );
  NANDN U14717 ( .A(n14667), .B(n14668), .Z(n14666) );
  NANDN U14718 ( .A(n14669), .B(n14670), .Z(n14668) );
  NANDN U14719 ( .A(n14670), .B(n14669), .Z(n14665) );
  ANDN U14720 ( .B(B[251]), .A(n69), .Z(n14530) );
  XNOR U14721 ( .A(n14538), .B(n14671), .Z(n14531) );
  XNOR U14722 ( .A(n14537), .B(n14535), .Z(n14671) );
  AND U14723 ( .A(n14672), .B(n14673), .Z(n14535) );
  NANDN U14724 ( .A(n14674), .B(n14675), .Z(n14673) );
  OR U14725 ( .A(n14676), .B(n14677), .Z(n14675) );
  NAND U14726 ( .A(n14677), .B(n14676), .Z(n14672) );
  ANDN U14727 ( .B(B[252]), .A(n70), .Z(n14537) );
  XNOR U14728 ( .A(n14545), .B(n14678), .Z(n14538) );
  XNOR U14729 ( .A(n14544), .B(n14542), .Z(n14678) );
  AND U14730 ( .A(n14679), .B(n14680), .Z(n14542) );
  NANDN U14731 ( .A(n14681), .B(n14682), .Z(n14680) );
  NANDN U14732 ( .A(n14683), .B(n14684), .Z(n14682) );
  NANDN U14733 ( .A(n14684), .B(n14683), .Z(n14679) );
  ANDN U14734 ( .B(B[253]), .A(n71), .Z(n14544) );
  XOR U14735 ( .A(n14550), .B(n14685), .Z(n14545) );
  XOR U14736 ( .A(n14551), .B(n14552), .Z(n14685) );
  NAND U14737 ( .A(A[12]), .B(B[255]), .Z(n14552) );
  AND U14738 ( .A(B[254]), .B(A[13]), .Z(n14551) );
  NAND U14739 ( .A(n14686), .B(n14687), .Z(n14550) );
  NAND U14740 ( .A(n14688), .B(n14689), .Z(n14687) );
  NANDN U14741 ( .A(n14690), .B(n14691), .Z(n14688) );
  NANDN U14742 ( .A(n14691), .B(n14690), .Z(n14686) );
  NAND U14743 ( .A(n14692), .B(n14693), .Z(n262) );
  NANDN U14744 ( .A(n14694), .B(n14695), .Z(n14693) );
  NAND U14745 ( .A(n14697), .B(n14696), .Z(n14692) );
  XOR U14746 ( .A(n264), .B(n263), .Z(\A1[264] ) );
  XOR U14747 ( .A(n14697), .B(n14698), .Z(n263) );
  XNOR U14748 ( .A(n14696), .B(n14694), .Z(n14698) );
  AND U14749 ( .A(n14699), .B(n14700), .Z(n14694) );
  NANDN U14750 ( .A(n14701), .B(n14702), .Z(n14700) );
  NANDN U14751 ( .A(n14703), .B(n14704), .Z(n14702) );
  NANDN U14752 ( .A(n14704), .B(n14703), .Z(n14699) );
  ANDN U14753 ( .B(B[235]), .A(n54), .Z(n14696) );
  XOR U14754 ( .A(n14565), .B(n14705), .Z(n14697) );
  XNOR U14755 ( .A(n14564), .B(n14562), .Z(n14705) );
  AND U14756 ( .A(n14706), .B(n14707), .Z(n14562) );
  NANDN U14757 ( .A(n14708), .B(n14709), .Z(n14707) );
  OR U14758 ( .A(n14710), .B(n14711), .Z(n14709) );
  NAND U14759 ( .A(n14711), .B(n14710), .Z(n14706) );
  ANDN U14760 ( .B(B[236]), .A(n55), .Z(n14564) );
  XNOR U14761 ( .A(n14572), .B(n14712), .Z(n14565) );
  XNOR U14762 ( .A(n14571), .B(n14569), .Z(n14712) );
  AND U14763 ( .A(n14713), .B(n14714), .Z(n14569) );
  NANDN U14764 ( .A(n14715), .B(n14716), .Z(n14714) );
  NANDN U14765 ( .A(n14717), .B(n14718), .Z(n14716) );
  NANDN U14766 ( .A(n14718), .B(n14717), .Z(n14713) );
  ANDN U14767 ( .B(B[237]), .A(n56), .Z(n14571) );
  XNOR U14768 ( .A(n14579), .B(n14719), .Z(n14572) );
  XNOR U14769 ( .A(n14578), .B(n14576), .Z(n14719) );
  AND U14770 ( .A(n14720), .B(n14721), .Z(n14576) );
  NANDN U14771 ( .A(n14722), .B(n14723), .Z(n14721) );
  OR U14772 ( .A(n14724), .B(n14725), .Z(n14723) );
  NAND U14773 ( .A(n14725), .B(n14724), .Z(n14720) );
  ANDN U14774 ( .B(B[238]), .A(n57), .Z(n14578) );
  XNOR U14775 ( .A(n14586), .B(n14726), .Z(n14579) );
  XNOR U14776 ( .A(n14585), .B(n14583), .Z(n14726) );
  AND U14777 ( .A(n14727), .B(n14728), .Z(n14583) );
  NANDN U14778 ( .A(n14729), .B(n14730), .Z(n14728) );
  NANDN U14779 ( .A(n14731), .B(n14732), .Z(n14730) );
  NANDN U14780 ( .A(n14732), .B(n14731), .Z(n14727) );
  ANDN U14781 ( .B(B[239]), .A(n58), .Z(n14585) );
  XNOR U14782 ( .A(n14593), .B(n14733), .Z(n14586) );
  XNOR U14783 ( .A(n14592), .B(n14590), .Z(n14733) );
  AND U14784 ( .A(n14734), .B(n14735), .Z(n14590) );
  NANDN U14785 ( .A(n14736), .B(n14737), .Z(n14735) );
  OR U14786 ( .A(n14738), .B(n14739), .Z(n14737) );
  NAND U14787 ( .A(n14739), .B(n14738), .Z(n14734) );
  ANDN U14788 ( .B(B[240]), .A(n59), .Z(n14592) );
  XNOR U14789 ( .A(n14600), .B(n14740), .Z(n14593) );
  XNOR U14790 ( .A(n14599), .B(n14597), .Z(n14740) );
  AND U14791 ( .A(n14741), .B(n14742), .Z(n14597) );
  NANDN U14792 ( .A(n14743), .B(n14744), .Z(n14742) );
  NANDN U14793 ( .A(n14745), .B(n14746), .Z(n14744) );
  NANDN U14794 ( .A(n14746), .B(n14745), .Z(n14741) );
  ANDN U14795 ( .B(B[241]), .A(n60), .Z(n14599) );
  XNOR U14796 ( .A(n14607), .B(n14747), .Z(n14600) );
  XNOR U14797 ( .A(n14606), .B(n14604), .Z(n14747) );
  AND U14798 ( .A(n14748), .B(n14749), .Z(n14604) );
  NANDN U14799 ( .A(n14750), .B(n14751), .Z(n14749) );
  OR U14800 ( .A(n14752), .B(n14753), .Z(n14751) );
  NAND U14801 ( .A(n14753), .B(n14752), .Z(n14748) );
  ANDN U14802 ( .B(B[242]), .A(n61), .Z(n14606) );
  XNOR U14803 ( .A(n14614), .B(n14754), .Z(n14607) );
  XNOR U14804 ( .A(n14613), .B(n14611), .Z(n14754) );
  AND U14805 ( .A(n14755), .B(n14756), .Z(n14611) );
  NANDN U14806 ( .A(n14757), .B(n14758), .Z(n14756) );
  NANDN U14807 ( .A(n14759), .B(n14760), .Z(n14758) );
  NANDN U14808 ( .A(n14760), .B(n14759), .Z(n14755) );
  ANDN U14809 ( .B(B[243]), .A(n62), .Z(n14613) );
  XNOR U14810 ( .A(n14621), .B(n14761), .Z(n14614) );
  XNOR U14811 ( .A(n14620), .B(n14618), .Z(n14761) );
  AND U14812 ( .A(n14762), .B(n14763), .Z(n14618) );
  NANDN U14813 ( .A(n14764), .B(n14765), .Z(n14763) );
  OR U14814 ( .A(n14766), .B(n14767), .Z(n14765) );
  NAND U14815 ( .A(n14767), .B(n14766), .Z(n14762) );
  ANDN U14816 ( .B(B[244]), .A(n63), .Z(n14620) );
  XNOR U14817 ( .A(n14628), .B(n14768), .Z(n14621) );
  XNOR U14818 ( .A(n14627), .B(n14625), .Z(n14768) );
  AND U14819 ( .A(n14769), .B(n14770), .Z(n14625) );
  NANDN U14820 ( .A(n14771), .B(n14772), .Z(n14770) );
  NANDN U14821 ( .A(n14773), .B(n14774), .Z(n14772) );
  NANDN U14822 ( .A(n14774), .B(n14773), .Z(n14769) );
  ANDN U14823 ( .B(B[245]), .A(n64), .Z(n14627) );
  XNOR U14824 ( .A(n14635), .B(n14775), .Z(n14628) );
  XNOR U14825 ( .A(n14634), .B(n14632), .Z(n14775) );
  AND U14826 ( .A(n14776), .B(n14777), .Z(n14632) );
  NANDN U14827 ( .A(n14778), .B(n14779), .Z(n14777) );
  OR U14828 ( .A(n14780), .B(n14781), .Z(n14779) );
  NAND U14829 ( .A(n14781), .B(n14780), .Z(n14776) );
  ANDN U14830 ( .B(B[246]), .A(n65), .Z(n14634) );
  XNOR U14831 ( .A(n14642), .B(n14782), .Z(n14635) );
  XNOR U14832 ( .A(n14641), .B(n14639), .Z(n14782) );
  AND U14833 ( .A(n14783), .B(n14784), .Z(n14639) );
  NANDN U14834 ( .A(n14785), .B(n14786), .Z(n14784) );
  NANDN U14835 ( .A(n14787), .B(n14788), .Z(n14786) );
  NANDN U14836 ( .A(n14788), .B(n14787), .Z(n14783) );
  ANDN U14837 ( .B(B[247]), .A(n66), .Z(n14641) );
  XNOR U14838 ( .A(n14649), .B(n14789), .Z(n14642) );
  XNOR U14839 ( .A(n14648), .B(n14646), .Z(n14789) );
  AND U14840 ( .A(n14790), .B(n14791), .Z(n14646) );
  NANDN U14841 ( .A(n14792), .B(n14793), .Z(n14791) );
  OR U14842 ( .A(n14794), .B(n14795), .Z(n14793) );
  NAND U14843 ( .A(n14795), .B(n14794), .Z(n14790) );
  ANDN U14844 ( .B(B[248]), .A(n67), .Z(n14648) );
  XNOR U14845 ( .A(n14656), .B(n14796), .Z(n14649) );
  XNOR U14846 ( .A(n14655), .B(n14653), .Z(n14796) );
  AND U14847 ( .A(n14797), .B(n14798), .Z(n14653) );
  NANDN U14848 ( .A(n14799), .B(n14800), .Z(n14798) );
  NANDN U14849 ( .A(n14801), .B(n14802), .Z(n14800) );
  NANDN U14850 ( .A(n14802), .B(n14801), .Z(n14797) );
  ANDN U14851 ( .B(B[249]), .A(n68), .Z(n14655) );
  XNOR U14852 ( .A(n14663), .B(n14803), .Z(n14656) );
  XNOR U14853 ( .A(n14662), .B(n14660), .Z(n14803) );
  AND U14854 ( .A(n14804), .B(n14805), .Z(n14660) );
  NANDN U14855 ( .A(n14806), .B(n14807), .Z(n14805) );
  OR U14856 ( .A(n14808), .B(n14809), .Z(n14807) );
  NAND U14857 ( .A(n14809), .B(n14808), .Z(n14804) );
  ANDN U14858 ( .B(B[250]), .A(n69), .Z(n14662) );
  XNOR U14859 ( .A(n14670), .B(n14810), .Z(n14663) );
  XNOR U14860 ( .A(n14669), .B(n14667), .Z(n14810) );
  AND U14861 ( .A(n14811), .B(n14812), .Z(n14667) );
  NANDN U14862 ( .A(n14813), .B(n14814), .Z(n14812) );
  NANDN U14863 ( .A(n14815), .B(n14816), .Z(n14814) );
  NANDN U14864 ( .A(n14816), .B(n14815), .Z(n14811) );
  ANDN U14865 ( .B(B[251]), .A(n70), .Z(n14669) );
  XNOR U14866 ( .A(n14677), .B(n14817), .Z(n14670) );
  XNOR U14867 ( .A(n14676), .B(n14674), .Z(n14817) );
  AND U14868 ( .A(n14818), .B(n14819), .Z(n14674) );
  NANDN U14869 ( .A(n14820), .B(n14821), .Z(n14819) );
  OR U14870 ( .A(n14822), .B(n14823), .Z(n14821) );
  NAND U14871 ( .A(n14823), .B(n14822), .Z(n14818) );
  ANDN U14872 ( .B(B[252]), .A(n71), .Z(n14676) );
  XNOR U14873 ( .A(n14684), .B(n14824), .Z(n14677) );
  XNOR U14874 ( .A(n14683), .B(n14681), .Z(n14824) );
  AND U14875 ( .A(n14825), .B(n14826), .Z(n14681) );
  NANDN U14876 ( .A(n14827), .B(n14828), .Z(n14826) );
  NANDN U14877 ( .A(n14829), .B(n14830), .Z(n14828) );
  NANDN U14878 ( .A(n14830), .B(n14829), .Z(n14825) );
  ANDN U14879 ( .B(B[253]), .A(n72), .Z(n14683) );
  XOR U14880 ( .A(n14689), .B(n14831), .Z(n14684) );
  XOR U14881 ( .A(n14690), .B(n14691), .Z(n14831) );
  NAND U14882 ( .A(A[11]), .B(B[255]), .Z(n14691) );
  AND U14883 ( .A(B[254]), .B(A[12]), .Z(n14690) );
  NAND U14884 ( .A(n14832), .B(n14833), .Z(n14689) );
  NAND U14885 ( .A(n14834), .B(n14835), .Z(n14833) );
  NANDN U14886 ( .A(n14836), .B(n14837), .Z(n14834) );
  NANDN U14887 ( .A(n14837), .B(n14836), .Z(n14832) );
  NAND U14888 ( .A(n14838), .B(n14839), .Z(n264) );
  NANDN U14889 ( .A(n14840), .B(n14841), .Z(n14839) );
  OR U14890 ( .A(n14842), .B(n14843), .Z(n14841) );
  NAND U14891 ( .A(n14843), .B(n14842), .Z(n14838) );
  XOR U14892 ( .A(n266), .B(n265), .Z(\A1[263] ) );
  XOR U14893 ( .A(n14843), .B(n14844), .Z(n265) );
  XNOR U14894 ( .A(n14842), .B(n14840), .Z(n14844) );
  AND U14895 ( .A(n14845), .B(n14846), .Z(n14840) );
  NANDN U14896 ( .A(n14847), .B(n14848), .Z(n14846) );
  OR U14897 ( .A(n14849), .B(n14850), .Z(n14848) );
  NAND U14898 ( .A(n14850), .B(n14849), .Z(n14845) );
  ANDN U14899 ( .B(B[234]), .A(n54), .Z(n14842) );
  XNOR U14900 ( .A(n14704), .B(n14851), .Z(n14843) );
  XNOR U14901 ( .A(n14703), .B(n14701), .Z(n14851) );
  AND U14902 ( .A(n14852), .B(n14853), .Z(n14701) );
  NANDN U14903 ( .A(n14854), .B(n14855), .Z(n14853) );
  NANDN U14904 ( .A(n14856), .B(n14857), .Z(n14855) );
  NANDN U14905 ( .A(n14857), .B(n14856), .Z(n14852) );
  ANDN U14906 ( .B(B[235]), .A(n55), .Z(n14703) );
  XNOR U14907 ( .A(n14711), .B(n14858), .Z(n14704) );
  XNOR U14908 ( .A(n14710), .B(n14708), .Z(n14858) );
  AND U14909 ( .A(n14859), .B(n14860), .Z(n14708) );
  NANDN U14910 ( .A(n14861), .B(n14862), .Z(n14860) );
  OR U14911 ( .A(n14863), .B(n14864), .Z(n14862) );
  NAND U14912 ( .A(n14864), .B(n14863), .Z(n14859) );
  ANDN U14913 ( .B(B[236]), .A(n56), .Z(n14710) );
  XNOR U14914 ( .A(n14718), .B(n14865), .Z(n14711) );
  XNOR U14915 ( .A(n14717), .B(n14715), .Z(n14865) );
  AND U14916 ( .A(n14866), .B(n14867), .Z(n14715) );
  NANDN U14917 ( .A(n14868), .B(n14869), .Z(n14867) );
  NANDN U14918 ( .A(n14870), .B(n14871), .Z(n14869) );
  NANDN U14919 ( .A(n14871), .B(n14870), .Z(n14866) );
  ANDN U14920 ( .B(B[237]), .A(n57), .Z(n14717) );
  XNOR U14921 ( .A(n14725), .B(n14872), .Z(n14718) );
  XNOR U14922 ( .A(n14724), .B(n14722), .Z(n14872) );
  AND U14923 ( .A(n14873), .B(n14874), .Z(n14722) );
  NANDN U14924 ( .A(n14875), .B(n14876), .Z(n14874) );
  OR U14925 ( .A(n14877), .B(n14878), .Z(n14876) );
  NAND U14926 ( .A(n14878), .B(n14877), .Z(n14873) );
  ANDN U14927 ( .B(B[238]), .A(n58), .Z(n14724) );
  XNOR U14928 ( .A(n14732), .B(n14879), .Z(n14725) );
  XNOR U14929 ( .A(n14731), .B(n14729), .Z(n14879) );
  AND U14930 ( .A(n14880), .B(n14881), .Z(n14729) );
  NANDN U14931 ( .A(n14882), .B(n14883), .Z(n14881) );
  NANDN U14932 ( .A(n14884), .B(n14885), .Z(n14883) );
  NANDN U14933 ( .A(n14885), .B(n14884), .Z(n14880) );
  ANDN U14934 ( .B(B[239]), .A(n59), .Z(n14731) );
  XNOR U14935 ( .A(n14739), .B(n14886), .Z(n14732) );
  XNOR U14936 ( .A(n14738), .B(n14736), .Z(n14886) );
  AND U14937 ( .A(n14887), .B(n14888), .Z(n14736) );
  NANDN U14938 ( .A(n14889), .B(n14890), .Z(n14888) );
  OR U14939 ( .A(n14891), .B(n14892), .Z(n14890) );
  NAND U14940 ( .A(n14892), .B(n14891), .Z(n14887) );
  ANDN U14941 ( .B(B[240]), .A(n60), .Z(n14738) );
  XNOR U14942 ( .A(n14746), .B(n14893), .Z(n14739) );
  XNOR U14943 ( .A(n14745), .B(n14743), .Z(n14893) );
  AND U14944 ( .A(n14894), .B(n14895), .Z(n14743) );
  NANDN U14945 ( .A(n14896), .B(n14897), .Z(n14895) );
  NANDN U14946 ( .A(n14898), .B(n14899), .Z(n14897) );
  NANDN U14947 ( .A(n14899), .B(n14898), .Z(n14894) );
  ANDN U14948 ( .B(B[241]), .A(n61), .Z(n14745) );
  XNOR U14949 ( .A(n14753), .B(n14900), .Z(n14746) );
  XNOR U14950 ( .A(n14752), .B(n14750), .Z(n14900) );
  AND U14951 ( .A(n14901), .B(n14902), .Z(n14750) );
  NANDN U14952 ( .A(n14903), .B(n14904), .Z(n14902) );
  OR U14953 ( .A(n14905), .B(n14906), .Z(n14904) );
  NAND U14954 ( .A(n14906), .B(n14905), .Z(n14901) );
  ANDN U14955 ( .B(B[242]), .A(n62), .Z(n14752) );
  XNOR U14956 ( .A(n14760), .B(n14907), .Z(n14753) );
  XNOR U14957 ( .A(n14759), .B(n14757), .Z(n14907) );
  AND U14958 ( .A(n14908), .B(n14909), .Z(n14757) );
  NANDN U14959 ( .A(n14910), .B(n14911), .Z(n14909) );
  NANDN U14960 ( .A(n14912), .B(n14913), .Z(n14911) );
  NANDN U14961 ( .A(n14913), .B(n14912), .Z(n14908) );
  ANDN U14962 ( .B(B[243]), .A(n63), .Z(n14759) );
  XNOR U14963 ( .A(n14767), .B(n14914), .Z(n14760) );
  XNOR U14964 ( .A(n14766), .B(n14764), .Z(n14914) );
  AND U14965 ( .A(n14915), .B(n14916), .Z(n14764) );
  NANDN U14966 ( .A(n14917), .B(n14918), .Z(n14916) );
  OR U14967 ( .A(n14919), .B(n14920), .Z(n14918) );
  NAND U14968 ( .A(n14920), .B(n14919), .Z(n14915) );
  ANDN U14969 ( .B(B[244]), .A(n64), .Z(n14766) );
  XNOR U14970 ( .A(n14774), .B(n14921), .Z(n14767) );
  XNOR U14971 ( .A(n14773), .B(n14771), .Z(n14921) );
  AND U14972 ( .A(n14922), .B(n14923), .Z(n14771) );
  NANDN U14973 ( .A(n14924), .B(n14925), .Z(n14923) );
  NANDN U14974 ( .A(n14926), .B(n14927), .Z(n14925) );
  NANDN U14975 ( .A(n14927), .B(n14926), .Z(n14922) );
  ANDN U14976 ( .B(B[245]), .A(n65), .Z(n14773) );
  XNOR U14977 ( .A(n14781), .B(n14928), .Z(n14774) );
  XNOR U14978 ( .A(n14780), .B(n14778), .Z(n14928) );
  AND U14979 ( .A(n14929), .B(n14930), .Z(n14778) );
  NANDN U14980 ( .A(n14931), .B(n14932), .Z(n14930) );
  OR U14981 ( .A(n14933), .B(n14934), .Z(n14932) );
  NAND U14982 ( .A(n14934), .B(n14933), .Z(n14929) );
  ANDN U14983 ( .B(B[246]), .A(n66), .Z(n14780) );
  XNOR U14984 ( .A(n14788), .B(n14935), .Z(n14781) );
  XNOR U14985 ( .A(n14787), .B(n14785), .Z(n14935) );
  AND U14986 ( .A(n14936), .B(n14937), .Z(n14785) );
  NANDN U14987 ( .A(n14938), .B(n14939), .Z(n14937) );
  NANDN U14988 ( .A(n14940), .B(n14941), .Z(n14939) );
  NANDN U14989 ( .A(n14941), .B(n14940), .Z(n14936) );
  ANDN U14990 ( .B(B[247]), .A(n67), .Z(n14787) );
  XNOR U14991 ( .A(n14795), .B(n14942), .Z(n14788) );
  XNOR U14992 ( .A(n14794), .B(n14792), .Z(n14942) );
  AND U14993 ( .A(n14943), .B(n14944), .Z(n14792) );
  NANDN U14994 ( .A(n14945), .B(n14946), .Z(n14944) );
  OR U14995 ( .A(n14947), .B(n14948), .Z(n14946) );
  NAND U14996 ( .A(n14948), .B(n14947), .Z(n14943) );
  ANDN U14997 ( .B(B[248]), .A(n68), .Z(n14794) );
  XNOR U14998 ( .A(n14802), .B(n14949), .Z(n14795) );
  XNOR U14999 ( .A(n14801), .B(n14799), .Z(n14949) );
  AND U15000 ( .A(n14950), .B(n14951), .Z(n14799) );
  NANDN U15001 ( .A(n14952), .B(n14953), .Z(n14951) );
  NANDN U15002 ( .A(n14954), .B(n14955), .Z(n14953) );
  NANDN U15003 ( .A(n14955), .B(n14954), .Z(n14950) );
  ANDN U15004 ( .B(B[249]), .A(n69), .Z(n14801) );
  XNOR U15005 ( .A(n14809), .B(n14956), .Z(n14802) );
  XNOR U15006 ( .A(n14808), .B(n14806), .Z(n14956) );
  AND U15007 ( .A(n14957), .B(n14958), .Z(n14806) );
  NANDN U15008 ( .A(n14959), .B(n14960), .Z(n14958) );
  OR U15009 ( .A(n14961), .B(n14962), .Z(n14960) );
  NAND U15010 ( .A(n14962), .B(n14961), .Z(n14957) );
  ANDN U15011 ( .B(B[250]), .A(n70), .Z(n14808) );
  XNOR U15012 ( .A(n14816), .B(n14963), .Z(n14809) );
  XNOR U15013 ( .A(n14815), .B(n14813), .Z(n14963) );
  AND U15014 ( .A(n14964), .B(n14965), .Z(n14813) );
  NANDN U15015 ( .A(n14966), .B(n14967), .Z(n14965) );
  NANDN U15016 ( .A(n14968), .B(n14969), .Z(n14967) );
  NANDN U15017 ( .A(n14969), .B(n14968), .Z(n14964) );
  ANDN U15018 ( .B(B[251]), .A(n71), .Z(n14815) );
  XNOR U15019 ( .A(n14823), .B(n14970), .Z(n14816) );
  XNOR U15020 ( .A(n14822), .B(n14820), .Z(n14970) );
  AND U15021 ( .A(n14971), .B(n14972), .Z(n14820) );
  NANDN U15022 ( .A(n14973), .B(n14974), .Z(n14972) );
  OR U15023 ( .A(n14975), .B(n14976), .Z(n14974) );
  NAND U15024 ( .A(n14976), .B(n14975), .Z(n14971) );
  ANDN U15025 ( .B(B[252]), .A(n72), .Z(n14822) );
  XNOR U15026 ( .A(n14830), .B(n14977), .Z(n14823) );
  XNOR U15027 ( .A(n14829), .B(n14827), .Z(n14977) );
  AND U15028 ( .A(n14978), .B(n14979), .Z(n14827) );
  NANDN U15029 ( .A(n14980), .B(n14981), .Z(n14979) );
  NANDN U15030 ( .A(n14982), .B(n14983), .Z(n14981) );
  NANDN U15031 ( .A(n14983), .B(n14982), .Z(n14978) );
  ANDN U15032 ( .B(B[253]), .A(n73), .Z(n14829) );
  XOR U15033 ( .A(n14835), .B(n14984), .Z(n14830) );
  XOR U15034 ( .A(n14836), .B(n14837), .Z(n14984) );
  NAND U15035 ( .A(A[10]), .B(B[255]), .Z(n14837) );
  AND U15036 ( .A(B[254]), .B(A[11]), .Z(n14836) );
  NAND U15037 ( .A(n14985), .B(n14986), .Z(n14835) );
  NAND U15038 ( .A(n14987), .B(n14988), .Z(n14986) );
  NANDN U15039 ( .A(n14989), .B(n14990), .Z(n14987) );
  NANDN U15040 ( .A(n14990), .B(n14989), .Z(n14985) );
  NAND U15041 ( .A(n14991), .B(n14992), .Z(n266) );
  NANDN U15042 ( .A(n14993), .B(n14994), .Z(n14992) );
  NAND U15043 ( .A(n14996), .B(n14995), .Z(n14991) );
  XOR U15044 ( .A(n268), .B(n267), .Z(\A1[262] ) );
  XOR U15045 ( .A(n14996), .B(n14997), .Z(n267) );
  XNOR U15046 ( .A(n14995), .B(n14993), .Z(n14997) );
  AND U15047 ( .A(n14998), .B(n14999), .Z(n14993) );
  NANDN U15048 ( .A(n15000), .B(n15001), .Z(n14999) );
  NANDN U15049 ( .A(n15002), .B(n15003), .Z(n15001) );
  NANDN U15050 ( .A(n15003), .B(n15002), .Z(n14998) );
  ANDN U15051 ( .B(B[233]), .A(n54), .Z(n14995) );
  XOR U15052 ( .A(n14850), .B(n15004), .Z(n14996) );
  XNOR U15053 ( .A(n14849), .B(n14847), .Z(n15004) );
  AND U15054 ( .A(n15005), .B(n15006), .Z(n14847) );
  NANDN U15055 ( .A(n15007), .B(n15008), .Z(n15006) );
  OR U15056 ( .A(n15009), .B(n15010), .Z(n15008) );
  NAND U15057 ( .A(n15010), .B(n15009), .Z(n15005) );
  ANDN U15058 ( .B(B[234]), .A(n55), .Z(n14849) );
  XNOR U15059 ( .A(n14857), .B(n15011), .Z(n14850) );
  XNOR U15060 ( .A(n14856), .B(n14854), .Z(n15011) );
  AND U15061 ( .A(n15012), .B(n15013), .Z(n14854) );
  NANDN U15062 ( .A(n15014), .B(n15015), .Z(n15013) );
  NANDN U15063 ( .A(n15016), .B(n15017), .Z(n15015) );
  NANDN U15064 ( .A(n15017), .B(n15016), .Z(n15012) );
  ANDN U15065 ( .B(B[235]), .A(n56), .Z(n14856) );
  XNOR U15066 ( .A(n14864), .B(n15018), .Z(n14857) );
  XNOR U15067 ( .A(n14863), .B(n14861), .Z(n15018) );
  AND U15068 ( .A(n15019), .B(n15020), .Z(n14861) );
  NANDN U15069 ( .A(n15021), .B(n15022), .Z(n15020) );
  OR U15070 ( .A(n15023), .B(n15024), .Z(n15022) );
  NAND U15071 ( .A(n15024), .B(n15023), .Z(n15019) );
  ANDN U15072 ( .B(B[236]), .A(n57), .Z(n14863) );
  XNOR U15073 ( .A(n14871), .B(n15025), .Z(n14864) );
  XNOR U15074 ( .A(n14870), .B(n14868), .Z(n15025) );
  AND U15075 ( .A(n15026), .B(n15027), .Z(n14868) );
  NANDN U15076 ( .A(n15028), .B(n15029), .Z(n15027) );
  NANDN U15077 ( .A(n15030), .B(n15031), .Z(n15029) );
  NANDN U15078 ( .A(n15031), .B(n15030), .Z(n15026) );
  ANDN U15079 ( .B(B[237]), .A(n58), .Z(n14870) );
  XNOR U15080 ( .A(n14878), .B(n15032), .Z(n14871) );
  XNOR U15081 ( .A(n14877), .B(n14875), .Z(n15032) );
  AND U15082 ( .A(n15033), .B(n15034), .Z(n14875) );
  NANDN U15083 ( .A(n15035), .B(n15036), .Z(n15034) );
  OR U15084 ( .A(n15037), .B(n15038), .Z(n15036) );
  NAND U15085 ( .A(n15038), .B(n15037), .Z(n15033) );
  ANDN U15086 ( .B(B[238]), .A(n59), .Z(n14877) );
  XNOR U15087 ( .A(n14885), .B(n15039), .Z(n14878) );
  XNOR U15088 ( .A(n14884), .B(n14882), .Z(n15039) );
  AND U15089 ( .A(n15040), .B(n15041), .Z(n14882) );
  NANDN U15090 ( .A(n15042), .B(n15043), .Z(n15041) );
  NANDN U15091 ( .A(n15044), .B(n15045), .Z(n15043) );
  NANDN U15092 ( .A(n15045), .B(n15044), .Z(n15040) );
  ANDN U15093 ( .B(B[239]), .A(n60), .Z(n14884) );
  XNOR U15094 ( .A(n14892), .B(n15046), .Z(n14885) );
  XNOR U15095 ( .A(n14891), .B(n14889), .Z(n15046) );
  AND U15096 ( .A(n15047), .B(n15048), .Z(n14889) );
  NANDN U15097 ( .A(n15049), .B(n15050), .Z(n15048) );
  OR U15098 ( .A(n15051), .B(n15052), .Z(n15050) );
  NAND U15099 ( .A(n15052), .B(n15051), .Z(n15047) );
  ANDN U15100 ( .B(B[240]), .A(n61), .Z(n14891) );
  XNOR U15101 ( .A(n14899), .B(n15053), .Z(n14892) );
  XNOR U15102 ( .A(n14898), .B(n14896), .Z(n15053) );
  AND U15103 ( .A(n15054), .B(n15055), .Z(n14896) );
  NANDN U15104 ( .A(n15056), .B(n15057), .Z(n15055) );
  NANDN U15105 ( .A(n15058), .B(n15059), .Z(n15057) );
  NANDN U15106 ( .A(n15059), .B(n15058), .Z(n15054) );
  ANDN U15107 ( .B(B[241]), .A(n62), .Z(n14898) );
  XNOR U15108 ( .A(n14906), .B(n15060), .Z(n14899) );
  XNOR U15109 ( .A(n14905), .B(n14903), .Z(n15060) );
  AND U15110 ( .A(n15061), .B(n15062), .Z(n14903) );
  NANDN U15111 ( .A(n15063), .B(n15064), .Z(n15062) );
  OR U15112 ( .A(n15065), .B(n15066), .Z(n15064) );
  NAND U15113 ( .A(n15066), .B(n15065), .Z(n15061) );
  ANDN U15114 ( .B(B[242]), .A(n63), .Z(n14905) );
  XNOR U15115 ( .A(n14913), .B(n15067), .Z(n14906) );
  XNOR U15116 ( .A(n14912), .B(n14910), .Z(n15067) );
  AND U15117 ( .A(n15068), .B(n15069), .Z(n14910) );
  NANDN U15118 ( .A(n15070), .B(n15071), .Z(n15069) );
  NANDN U15119 ( .A(n15072), .B(n15073), .Z(n15071) );
  NANDN U15120 ( .A(n15073), .B(n15072), .Z(n15068) );
  ANDN U15121 ( .B(B[243]), .A(n64), .Z(n14912) );
  XNOR U15122 ( .A(n14920), .B(n15074), .Z(n14913) );
  XNOR U15123 ( .A(n14919), .B(n14917), .Z(n15074) );
  AND U15124 ( .A(n15075), .B(n15076), .Z(n14917) );
  NANDN U15125 ( .A(n15077), .B(n15078), .Z(n15076) );
  OR U15126 ( .A(n15079), .B(n15080), .Z(n15078) );
  NAND U15127 ( .A(n15080), .B(n15079), .Z(n15075) );
  ANDN U15128 ( .B(B[244]), .A(n65), .Z(n14919) );
  XNOR U15129 ( .A(n14927), .B(n15081), .Z(n14920) );
  XNOR U15130 ( .A(n14926), .B(n14924), .Z(n15081) );
  AND U15131 ( .A(n15082), .B(n15083), .Z(n14924) );
  NANDN U15132 ( .A(n15084), .B(n15085), .Z(n15083) );
  NANDN U15133 ( .A(n15086), .B(n15087), .Z(n15085) );
  NANDN U15134 ( .A(n15087), .B(n15086), .Z(n15082) );
  ANDN U15135 ( .B(B[245]), .A(n66), .Z(n14926) );
  XNOR U15136 ( .A(n14934), .B(n15088), .Z(n14927) );
  XNOR U15137 ( .A(n14933), .B(n14931), .Z(n15088) );
  AND U15138 ( .A(n15089), .B(n15090), .Z(n14931) );
  NANDN U15139 ( .A(n15091), .B(n15092), .Z(n15090) );
  OR U15140 ( .A(n15093), .B(n15094), .Z(n15092) );
  NAND U15141 ( .A(n15094), .B(n15093), .Z(n15089) );
  ANDN U15142 ( .B(B[246]), .A(n67), .Z(n14933) );
  XNOR U15143 ( .A(n14941), .B(n15095), .Z(n14934) );
  XNOR U15144 ( .A(n14940), .B(n14938), .Z(n15095) );
  AND U15145 ( .A(n15096), .B(n15097), .Z(n14938) );
  NANDN U15146 ( .A(n15098), .B(n15099), .Z(n15097) );
  NANDN U15147 ( .A(n15100), .B(n15101), .Z(n15099) );
  NANDN U15148 ( .A(n15101), .B(n15100), .Z(n15096) );
  ANDN U15149 ( .B(B[247]), .A(n68), .Z(n14940) );
  XNOR U15150 ( .A(n14948), .B(n15102), .Z(n14941) );
  XNOR U15151 ( .A(n14947), .B(n14945), .Z(n15102) );
  AND U15152 ( .A(n15103), .B(n15104), .Z(n14945) );
  NANDN U15153 ( .A(n15105), .B(n15106), .Z(n15104) );
  OR U15154 ( .A(n15107), .B(n15108), .Z(n15106) );
  NAND U15155 ( .A(n15108), .B(n15107), .Z(n15103) );
  ANDN U15156 ( .B(B[248]), .A(n69), .Z(n14947) );
  XNOR U15157 ( .A(n14955), .B(n15109), .Z(n14948) );
  XNOR U15158 ( .A(n14954), .B(n14952), .Z(n15109) );
  AND U15159 ( .A(n15110), .B(n15111), .Z(n14952) );
  NANDN U15160 ( .A(n15112), .B(n15113), .Z(n15111) );
  NANDN U15161 ( .A(n15114), .B(n15115), .Z(n15113) );
  NANDN U15162 ( .A(n15115), .B(n15114), .Z(n15110) );
  ANDN U15163 ( .B(B[249]), .A(n70), .Z(n14954) );
  XNOR U15164 ( .A(n14962), .B(n15116), .Z(n14955) );
  XNOR U15165 ( .A(n14961), .B(n14959), .Z(n15116) );
  AND U15166 ( .A(n15117), .B(n15118), .Z(n14959) );
  NANDN U15167 ( .A(n15119), .B(n15120), .Z(n15118) );
  OR U15168 ( .A(n15121), .B(n15122), .Z(n15120) );
  NAND U15169 ( .A(n15122), .B(n15121), .Z(n15117) );
  ANDN U15170 ( .B(B[250]), .A(n71), .Z(n14961) );
  XNOR U15171 ( .A(n14969), .B(n15123), .Z(n14962) );
  XNOR U15172 ( .A(n14968), .B(n14966), .Z(n15123) );
  AND U15173 ( .A(n15124), .B(n15125), .Z(n14966) );
  NANDN U15174 ( .A(n15126), .B(n15127), .Z(n15125) );
  NANDN U15175 ( .A(n15128), .B(n15129), .Z(n15127) );
  NANDN U15176 ( .A(n15129), .B(n15128), .Z(n15124) );
  ANDN U15177 ( .B(B[251]), .A(n72), .Z(n14968) );
  XNOR U15178 ( .A(n14976), .B(n15130), .Z(n14969) );
  XNOR U15179 ( .A(n14975), .B(n14973), .Z(n15130) );
  AND U15180 ( .A(n15131), .B(n15132), .Z(n14973) );
  NANDN U15181 ( .A(n15133), .B(n15134), .Z(n15132) );
  OR U15182 ( .A(n15135), .B(n15136), .Z(n15134) );
  NAND U15183 ( .A(n15136), .B(n15135), .Z(n15131) );
  ANDN U15184 ( .B(B[252]), .A(n73), .Z(n14975) );
  XNOR U15185 ( .A(n14983), .B(n15137), .Z(n14976) );
  XNOR U15186 ( .A(n14982), .B(n14980), .Z(n15137) );
  AND U15187 ( .A(n15138), .B(n15139), .Z(n14980) );
  NANDN U15188 ( .A(n15140), .B(n15141), .Z(n15139) );
  NANDN U15189 ( .A(n15142), .B(n15143), .Z(n15141) );
  NANDN U15190 ( .A(n15143), .B(n15142), .Z(n15138) );
  ANDN U15191 ( .B(B[253]), .A(n74), .Z(n14982) );
  XOR U15192 ( .A(n14988), .B(n15144), .Z(n14983) );
  XOR U15193 ( .A(n14989), .B(n14990), .Z(n15144) );
  NAND U15194 ( .A(A[9]), .B(B[255]), .Z(n14990) );
  AND U15195 ( .A(B[254]), .B(A[10]), .Z(n14989) );
  NAND U15196 ( .A(n15145), .B(n15146), .Z(n14988) );
  NAND U15197 ( .A(n15147), .B(n15148), .Z(n15146) );
  NANDN U15198 ( .A(n15149), .B(n15150), .Z(n15147) );
  NANDN U15199 ( .A(n15150), .B(n15149), .Z(n15145) );
  NAND U15200 ( .A(n15151), .B(n15152), .Z(n268) );
  NANDN U15201 ( .A(n15153), .B(n15154), .Z(n15152) );
  OR U15202 ( .A(n15155), .B(n15156), .Z(n15154) );
  NAND U15203 ( .A(n15156), .B(n15155), .Z(n15151) );
  XOR U15204 ( .A(n270), .B(n269), .Z(\A1[261] ) );
  XOR U15205 ( .A(n15156), .B(n15157), .Z(n269) );
  XNOR U15206 ( .A(n15155), .B(n15153), .Z(n15157) );
  AND U15207 ( .A(n15158), .B(n15159), .Z(n15153) );
  NANDN U15208 ( .A(n15160), .B(n15161), .Z(n15159) );
  OR U15209 ( .A(n15162), .B(n15163), .Z(n15161) );
  NAND U15210 ( .A(n15163), .B(n15162), .Z(n15158) );
  ANDN U15211 ( .B(B[232]), .A(n54), .Z(n15155) );
  XNOR U15212 ( .A(n15003), .B(n15164), .Z(n15156) );
  XNOR U15213 ( .A(n15002), .B(n15000), .Z(n15164) );
  AND U15214 ( .A(n15165), .B(n15166), .Z(n15000) );
  NANDN U15215 ( .A(n15167), .B(n15168), .Z(n15166) );
  NANDN U15216 ( .A(n15169), .B(n15170), .Z(n15168) );
  NANDN U15217 ( .A(n15170), .B(n15169), .Z(n15165) );
  ANDN U15218 ( .B(B[233]), .A(n55), .Z(n15002) );
  XNOR U15219 ( .A(n15010), .B(n15171), .Z(n15003) );
  XNOR U15220 ( .A(n15009), .B(n15007), .Z(n15171) );
  AND U15221 ( .A(n15172), .B(n15173), .Z(n15007) );
  NANDN U15222 ( .A(n15174), .B(n15175), .Z(n15173) );
  OR U15223 ( .A(n15176), .B(n15177), .Z(n15175) );
  NAND U15224 ( .A(n15177), .B(n15176), .Z(n15172) );
  ANDN U15225 ( .B(B[234]), .A(n56), .Z(n15009) );
  XNOR U15226 ( .A(n15017), .B(n15178), .Z(n15010) );
  XNOR U15227 ( .A(n15016), .B(n15014), .Z(n15178) );
  AND U15228 ( .A(n15179), .B(n15180), .Z(n15014) );
  NANDN U15229 ( .A(n15181), .B(n15182), .Z(n15180) );
  NANDN U15230 ( .A(n15183), .B(n15184), .Z(n15182) );
  NANDN U15231 ( .A(n15184), .B(n15183), .Z(n15179) );
  ANDN U15232 ( .B(B[235]), .A(n57), .Z(n15016) );
  XNOR U15233 ( .A(n15024), .B(n15185), .Z(n15017) );
  XNOR U15234 ( .A(n15023), .B(n15021), .Z(n15185) );
  AND U15235 ( .A(n15186), .B(n15187), .Z(n15021) );
  NANDN U15236 ( .A(n15188), .B(n15189), .Z(n15187) );
  OR U15237 ( .A(n15190), .B(n15191), .Z(n15189) );
  NAND U15238 ( .A(n15191), .B(n15190), .Z(n15186) );
  ANDN U15239 ( .B(B[236]), .A(n58), .Z(n15023) );
  XNOR U15240 ( .A(n15031), .B(n15192), .Z(n15024) );
  XNOR U15241 ( .A(n15030), .B(n15028), .Z(n15192) );
  AND U15242 ( .A(n15193), .B(n15194), .Z(n15028) );
  NANDN U15243 ( .A(n15195), .B(n15196), .Z(n15194) );
  NANDN U15244 ( .A(n15197), .B(n15198), .Z(n15196) );
  NANDN U15245 ( .A(n15198), .B(n15197), .Z(n15193) );
  ANDN U15246 ( .B(B[237]), .A(n59), .Z(n15030) );
  XNOR U15247 ( .A(n15038), .B(n15199), .Z(n15031) );
  XNOR U15248 ( .A(n15037), .B(n15035), .Z(n15199) );
  AND U15249 ( .A(n15200), .B(n15201), .Z(n15035) );
  NANDN U15250 ( .A(n15202), .B(n15203), .Z(n15201) );
  OR U15251 ( .A(n15204), .B(n15205), .Z(n15203) );
  NAND U15252 ( .A(n15205), .B(n15204), .Z(n15200) );
  ANDN U15253 ( .B(B[238]), .A(n60), .Z(n15037) );
  XNOR U15254 ( .A(n15045), .B(n15206), .Z(n15038) );
  XNOR U15255 ( .A(n15044), .B(n15042), .Z(n15206) );
  AND U15256 ( .A(n15207), .B(n15208), .Z(n15042) );
  NANDN U15257 ( .A(n15209), .B(n15210), .Z(n15208) );
  NANDN U15258 ( .A(n15211), .B(n15212), .Z(n15210) );
  NANDN U15259 ( .A(n15212), .B(n15211), .Z(n15207) );
  ANDN U15260 ( .B(B[239]), .A(n61), .Z(n15044) );
  XNOR U15261 ( .A(n15052), .B(n15213), .Z(n15045) );
  XNOR U15262 ( .A(n15051), .B(n15049), .Z(n15213) );
  AND U15263 ( .A(n15214), .B(n15215), .Z(n15049) );
  NANDN U15264 ( .A(n15216), .B(n15217), .Z(n15215) );
  OR U15265 ( .A(n15218), .B(n15219), .Z(n15217) );
  NAND U15266 ( .A(n15219), .B(n15218), .Z(n15214) );
  ANDN U15267 ( .B(B[240]), .A(n62), .Z(n15051) );
  XNOR U15268 ( .A(n15059), .B(n15220), .Z(n15052) );
  XNOR U15269 ( .A(n15058), .B(n15056), .Z(n15220) );
  AND U15270 ( .A(n15221), .B(n15222), .Z(n15056) );
  NANDN U15271 ( .A(n15223), .B(n15224), .Z(n15222) );
  NANDN U15272 ( .A(n15225), .B(n15226), .Z(n15224) );
  NANDN U15273 ( .A(n15226), .B(n15225), .Z(n15221) );
  ANDN U15274 ( .B(B[241]), .A(n63), .Z(n15058) );
  XNOR U15275 ( .A(n15066), .B(n15227), .Z(n15059) );
  XNOR U15276 ( .A(n15065), .B(n15063), .Z(n15227) );
  AND U15277 ( .A(n15228), .B(n15229), .Z(n15063) );
  NANDN U15278 ( .A(n15230), .B(n15231), .Z(n15229) );
  OR U15279 ( .A(n15232), .B(n15233), .Z(n15231) );
  NAND U15280 ( .A(n15233), .B(n15232), .Z(n15228) );
  ANDN U15281 ( .B(B[242]), .A(n64), .Z(n15065) );
  XNOR U15282 ( .A(n15073), .B(n15234), .Z(n15066) );
  XNOR U15283 ( .A(n15072), .B(n15070), .Z(n15234) );
  AND U15284 ( .A(n15235), .B(n15236), .Z(n15070) );
  NANDN U15285 ( .A(n15237), .B(n15238), .Z(n15236) );
  NANDN U15286 ( .A(n15239), .B(n15240), .Z(n15238) );
  NANDN U15287 ( .A(n15240), .B(n15239), .Z(n15235) );
  ANDN U15288 ( .B(B[243]), .A(n65), .Z(n15072) );
  XNOR U15289 ( .A(n15080), .B(n15241), .Z(n15073) );
  XNOR U15290 ( .A(n15079), .B(n15077), .Z(n15241) );
  AND U15291 ( .A(n15242), .B(n15243), .Z(n15077) );
  NANDN U15292 ( .A(n15244), .B(n15245), .Z(n15243) );
  OR U15293 ( .A(n15246), .B(n15247), .Z(n15245) );
  NAND U15294 ( .A(n15247), .B(n15246), .Z(n15242) );
  ANDN U15295 ( .B(B[244]), .A(n66), .Z(n15079) );
  XNOR U15296 ( .A(n15087), .B(n15248), .Z(n15080) );
  XNOR U15297 ( .A(n15086), .B(n15084), .Z(n15248) );
  AND U15298 ( .A(n15249), .B(n15250), .Z(n15084) );
  NANDN U15299 ( .A(n15251), .B(n15252), .Z(n15250) );
  NANDN U15300 ( .A(n15253), .B(n15254), .Z(n15252) );
  NANDN U15301 ( .A(n15254), .B(n15253), .Z(n15249) );
  ANDN U15302 ( .B(B[245]), .A(n67), .Z(n15086) );
  XNOR U15303 ( .A(n15094), .B(n15255), .Z(n15087) );
  XNOR U15304 ( .A(n15093), .B(n15091), .Z(n15255) );
  AND U15305 ( .A(n15256), .B(n15257), .Z(n15091) );
  NANDN U15306 ( .A(n15258), .B(n15259), .Z(n15257) );
  OR U15307 ( .A(n15260), .B(n15261), .Z(n15259) );
  NAND U15308 ( .A(n15261), .B(n15260), .Z(n15256) );
  ANDN U15309 ( .B(B[246]), .A(n68), .Z(n15093) );
  XNOR U15310 ( .A(n15101), .B(n15262), .Z(n15094) );
  XNOR U15311 ( .A(n15100), .B(n15098), .Z(n15262) );
  AND U15312 ( .A(n15263), .B(n15264), .Z(n15098) );
  NANDN U15313 ( .A(n15265), .B(n15266), .Z(n15264) );
  NANDN U15314 ( .A(n15267), .B(n15268), .Z(n15266) );
  NANDN U15315 ( .A(n15268), .B(n15267), .Z(n15263) );
  ANDN U15316 ( .B(B[247]), .A(n69), .Z(n15100) );
  XNOR U15317 ( .A(n15108), .B(n15269), .Z(n15101) );
  XNOR U15318 ( .A(n15107), .B(n15105), .Z(n15269) );
  AND U15319 ( .A(n15270), .B(n15271), .Z(n15105) );
  NANDN U15320 ( .A(n15272), .B(n15273), .Z(n15271) );
  OR U15321 ( .A(n15274), .B(n15275), .Z(n15273) );
  NAND U15322 ( .A(n15275), .B(n15274), .Z(n15270) );
  ANDN U15323 ( .B(B[248]), .A(n70), .Z(n15107) );
  XNOR U15324 ( .A(n15115), .B(n15276), .Z(n15108) );
  XNOR U15325 ( .A(n15114), .B(n15112), .Z(n15276) );
  AND U15326 ( .A(n15277), .B(n15278), .Z(n15112) );
  NANDN U15327 ( .A(n15279), .B(n15280), .Z(n15278) );
  NANDN U15328 ( .A(n15281), .B(n15282), .Z(n15280) );
  NANDN U15329 ( .A(n15282), .B(n15281), .Z(n15277) );
  ANDN U15330 ( .B(B[249]), .A(n71), .Z(n15114) );
  XNOR U15331 ( .A(n15122), .B(n15283), .Z(n15115) );
  XNOR U15332 ( .A(n15121), .B(n15119), .Z(n15283) );
  AND U15333 ( .A(n15284), .B(n15285), .Z(n15119) );
  NANDN U15334 ( .A(n15286), .B(n15287), .Z(n15285) );
  OR U15335 ( .A(n15288), .B(n15289), .Z(n15287) );
  NAND U15336 ( .A(n15289), .B(n15288), .Z(n15284) );
  ANDN U15337 ( .B(B[250]), .A(n72), .Z(n15121) );
  XNOR U15338 ( .A(n15129), .B(n15290), .Z(n15122) );
  XNOR U15339 ( .A(n15128), .B(n15126), .Z(n15290) );
  AND U15340 ( .A(n15291), .B(n15292), .Z(n15126) );
  NANDN U15341 ( .A(n15293), .B(n15294), .Z(n15292) );
  NANDN U15342 ( .A(n15295), .B(n15296), .Z(n15294) );
  NANDN U15343 ( .A(n15296), .B(n15295), .Z(n15291) );
  ANDN U15344 ( .B(B[251]), .A(n73), .Z(n15128) );
  XNOR U15345 ( .A(n15136), .B(n15297), .Z(n15129) );
  XNOR U15346 ( .A(n15135), .B(n15133), .Z(n15297) );
  AND U15347 ( .A(n15298), .B(n15299), .Z(n15133) );
  NANDN U15348 ( .A(n15300), .B(n15301), .Z(n15299) );
  OR U15349 ( .A(n15302), .B(n15303), .Z(n15301) );
  NAND U15350 ( .A(n15303), .B(n15302), .Z(n15298) );
  ANDN U15351 ( .B(B[252]), .A(n74), .Z(n15135) );
  XNOR U15352 ( .A(n15143), .B(n15304), .Z(n15136) );
  XNOR U15353 ( .A(n15142), .B(n15140), .Z(n15304) );
  AND U15354 ( .A(n15305), .B(n15306), .Z(n15140) );
  NANDN U15355 ( .A(n15307), .B(n15308), .Z(n15306) );
  NANDN U15356 ( .A(n15309), .B(n15310), .Z(n15308) );
  NANDN U15357 ( .A(n15310), .B(n15309), .Z(n15305) );
  ANDN U15358 ( .B(B[253]), .A(n75), .Z(n15142) );
  XOR U15359 ( .A(n15148), .B(n15311), .Z(n15143) );
  XOR U15360 ( .A(n15149), .B(n15150), .Z(n15311) );
  NAND U15361 ( .A(A[8]), .B(B[255]), .Z(n15150) );
  AND U15362 ( .A(B[254]), .B(A[9]), .Z(n15149) );
  NAND U15363 ( .A(n15312), .B(n15313), .Z(n15148) );
  NAND U15364 ( .A(n15314), .B(n15315), .Z(n15313) );
  NANDN U15365 ( .A(n15316), .B(n15317), .Z(n15314) );
  NANDN U15366 ( .A(n15317), .B(n15316), .Z(n15312) );
  NAND U15367 ( .A(n15318), .B(n15319), .Z(n270) );
  NANDN U15368 ( .A(n15320), .B(n15321), .Z(n15319) );
  NAND U15369 ( .A(n15323), .B(n15322), .Z(n15318) );
  XOR U15370 ( .A(n272), .B(n271), .Z(\A1[260] ) );
  XOR U15371 ( .A(n15323), .B(n15324), .Z(n271) );
  XNOR U15372 ( .A(n15322), .B(n15320), .Z(n15324) );
  AND U15373 ( .A(n15325), .B(n15326), .Z(n15320) );
  NANDN U15374 ( .A(n15327), .B(n15328), .Z(n15326) );
  NANDN U15375 ( .A(n15329), .B(n15330), .Z(n15328) );
  NANDN U15376 ( .A(n15330), .B(n15329), .Z(n15325) );
  ANDN U15377 ( .B(B[231]), .A(n54), .Z(n15322) );
  XOR U15378 ( .A(n15163), .B(n15331), .Z(n15323) );
  XNOR U15379 ( .A(n15162), .B(n15160), .Z(n15331) );
  AND U15380 ( .A(n15332), .B(n15333), .Z(n15160) );
  NANDN U15381 ( .A(n15334), .B(n15335), .Z(n15333) );
  OR U15382 ( .A(n15336), .B(n15337), .Z(n15335) );
  NAND U15383 ( .A(n15337), .B(n15336), .Z(n15332) );
  ANDN U15384 ( .B(B[232]), .A(n55), .Z(n15162) );
  XNOR U15385 ( .A(n15170), .B(n15338), .Z(n15163) );
  XNOR U15386 ( .A(n15169), .B(n15167), .Z(n15338) );
  AND U15387 ( .A(n15339), .B(n15340), .Z(n15167) );
  NANDN U15388 ( .A(n15341), .B(n15342), .Z(n15340) );
  NANDN U15389 ( .A(n15343), .B(n15344), .Z(n15342) );
  NANDN U15390 ( .A(n15344), .B(n15343), .Z(n15339) );
  ANDN U15391 ( .B(B[233]), .A(n56), .Z(n15169) );
  XNOR U15392 ( .A(n15177), .B(n15345), .Z(n15170) );
  XNOR U15393 ( .A(n15176), .B(n15174), .Z(n15345) );
  AND U15394 ( .A(n15346), .B(n15347), .Z(n15174) );
  NANDN U15395 ( .A(n15348), .B(n15349), .Z(n15347) );
  OR U15396 ( .A(n15350), .B(n15351), .Z(n15349) );
  NAND U15397 ( .A(n15351), .B(n15350), .Z(n15346) );
  ANDN U15398 ( .B(B[234]), .A(n57), .Z(n15176) );
  XNOR U15399 ( .A(n15184), .B(n15352), .Z(n15177) );
  XNOR U15400 ( .A(n15183), .B(n15181), .Z(n15352) );
  AND U15401 ( .A(n15353), .B(n15354), .Z(n15181) );
  NANDN U15402 ( .A(n15355), .B(n15356), .Z(n15354) );
  NANDN U15403 ( .A(n15357), .B(n15358), .Z(n15356) );
  NANDN U15404 ( .A(n15358), .B(n15357), .Z(n15353) );
  ANDN U15405 ( .B(B[235]), .A(n58), .Z(n15183) );
  XNOR U15406 ( .A(n15191), .B(n15359), .Z(n15184) );
  XNOR U15407 ( .A(n15190), .B(n15188), .Z(n15359) );
  AND U15408 ( .A(n15360), .B(n15361), .Z(n15188) );
  NANDN U15409 ( .A(n15362), .B(n15363), .Z(n15361) );
  OR U15410 ( .A(n15364), .B(n15365), .Z(n15363) );
  NAND U15411 ( .A(n15365), .B(n15364), .Z(n15360) );
  ANDN U15412 ( .B(B[236]), .A(n59), .Z(n15190) );
  XNOR U15413 ( .A(n15198), .B(n15366), .Z(n15191) );
  XNOR U15414 ( .A(n15197), .B(n15195), .Z(n15366) );
  AND U15415 ( .A(n15367), .B(n15368), .Z(n15195) );
  NANDN U15416 ( .A(n15369), .B(n15370), .Z(n15368) );
  NANDN U15417 ( .A(n15371), .B(n15372), .Z(n15370) );
  NANDN U15418 ( .A(n15372), .B(n15371), .Z(n15367) );
  ANDN U15419 ( .B(B[237]), .A(n60), .Z(n15197) );
  XNOR U15420 ( .A(n15205), .B(n15373), .Z(n15198) );
  XNOR U15421 ( .A(n15204), .B(n15202), .Z(n15373) );
  AND U15422 ( .A(n15374), .B(n15375), .Z(n15202) );
  NANDN U15423 ( .A(n15376), .B(n15377), .Z(n15375) );
  OR U15424 ( .A(n15378), .B(n15379), .Z(n15377) );
  NAND U15425 ( .A(n15379), .B(n15378), .Z(n15374) );
  ANDN U15426 ( .B(B[238]), .A(n61), .Z(n15204) );
  XNOR U15427 ( .A(n15212), .B(n15380), .Z(n15205) );
  XNOR U15428 ( .A(n15211), .B(n15209), .Z(n15380) );
  AND U15429 ( .A(n15381), .B(n15382), .Z(n15209) );
  NANDN U15430 ( .A(n15383), .B(n15384), .Z(n15382) );
  NANDN U15431 ( .A(n15385), .B(n15386), .Z(n15384) );
  NANDN U15432 ( .A(n15386), .B(n15385), .Z(n15381) );
  ANDN U15433 ( .B(B[239]), .A(n62), .Z(n15211) );
  XNOR U15434 ( .A(n15219), .B(n15387), .Z(n15212) );
  XNOR U15435 ( .A(n15218), .B(n15216), .Z(n15387) );
  AND U15436 ( .A(n15388), .B(n15389), .Z(n15216) );
  NANDN U15437 ( .A(n15390), .B(n15391), .Z(n15389) );
  OR U15438 ( .A(n15392), .B(n15393), .Z(n15391) );
  NAND U15439 ( .A(n15393), .B(n15392), .Z(n15388) );
  ANDN U15440 ( .B(B[240]), .A(n63), .Z(n15218) );
  XNOR U15441 ( .A(n15226), .B(n15394), .Z(n15219) );
  XNOR U15442 ( .A(n15225), .B(n15223), .Z(n15394) );
  AND U15443 ( .A(n15395), .B(n15396), .Z(n15223) );
  NANDN U15444 ( .A(n15397), .B(n15398), .Z(n15396) );
  NANDN U15445 ( .A(n15399), .B(n15400), .Z(n15398) );
  NANDN U15446 ( .A(n15400), .B(n15399), .Z(n15395) );
  ANDN U15447 ( .B(B[241]), .A(n64), .Z(n15225) );
  XNOR U15448 ( .A(n15233), .B(n15401), .Z(n15226) );
  XNOR U15449 ( .A(n15232), .B(n15230), .Z(n15401) );
  AND U15450 ( .A(n15402), .B(n15403), .Z(n15230) );
  NANDN U15451 ( .A(n15404), .B(n15405), .Z(n15403) );
  OR U15452 ( .A(n15406), .B(n15407), .Z(n15405) );
  NAND U15453 ( .A(n15407), .B(n15406), .Z(n15402) );
  ANDN U15454 ( .B(B[242]), .A(n65), .Z(n15232) );
  XNOR U15455 ( .A(n15240), .B(n15408), .Z(n15233) );
  XNOR U15456 ( .A(n15239), .B(n15237), .Z(n15408) );
  AND U15457 ( .A(n15409), .B(n15410), .Z(n15237) );
  NANDN U15458 ( .A(n15411), .B(n15412), .Z(n15410) );
  NANDN U15459 ( .A(n15413), .B(n15414), .Z(n15412) );
  NANDN U15460 ( .A(n15414), .B(n15413), .Z(n15409) );
  ANDN U15461 ( .B(B[243]), .A(n66), .Z(n15239) );
  XNOR U15462 ( .A(n15247), .B(n15415), .Z(n15240) );
  XNOR U15463 ( .A(n15246), .B(n15244), .Z(n15415) );
  AND U15464 ( .A(n15416), .B(n15417), .Z(n15244) );
  NANDN U15465 ( .A(n15418), .B(n15419), .Z(n15417) );
  OR U15466 ( .A(n15420), .B(n15421), .Z(n15419) );
  NAND U15467 ( .A(n15421), .B(n15420), .Z(n15416) );
  ANDN U15468 ( .B(B[244]), .A(n67), .Z(n15246) );
  XNOR U15469 ( .A(n15254), .B(n15422), .Z(n15247) );
  XNOR U15470 ( .A(n15253), .B(n15251), .Z(n15422) );
  AND U15471 ( .A(n15423), .B(n15424), .Z(n15251) );
  NANDN U15472 ( .A(n15425), .B(n15426), .Z(n15424) );
  NANDN U15473 ( .A(n15427), .B(n15428), .Z(n15426) );
  NANDN U15474 ( .A(n15428), .B(n15427), .Z(n15423) );
  ANDN U15475 ( .B(B[245]), .A(n68), .Z(n15253) );
  XNOR U15476 ( .A(n15261), .B(n15429), .Z(n15254) );
  XNOR U15477 ( .A(n15260), .B(n15258), .Z(n15429) );
  AND U15478 ( .A(n15430), .B(n15431), .Z(n15258) );
  NANDN U15479 ( .A(n15432), .B(n15433), .Z(n15431) );
  OR U15480 ( .A(n15434), .B(n15435), .Z(n15433) );
  NAND U15481 ( .A(n15435), .B(n15434), .Z(n15430) );
  ANDN U15482 ( .B(B[246]), .A(n69), .Z(n15260) );
  XNOR U15483 ( .A(n15268), .B(n15436), .Z(n15261) );
  XNOR U15484 ( .A(n15267), .B(n15265), .Z(n15436) );
  AND U15485 ( .A(n15437), .B(n15438), .Z(n15265) );
  NANDN U15486 ( .A(n15439), .B(n15440), .Z(n15438) );
  NANDN U15487 ( .A(n15441), .B(n15442), .Z(n15440) );
  NANDN U15488 ( .A(n15442), .B(n15441), .Z(n15437) );
  ANDN U15489 ( .B(B[247]), .A(n70), .Z(n15267) );
  XNOR U15490 ( .A(n15275), .B(n15443), .Z(n15268) );
  XNOR U15491 ( .A(n15274), .B(n15272), .Z(n15443) );
  AND U15492 ( .A(n15444), .B(n15445), .Z(n15272) );
  NANDN U15493 ( .A(n15446), .B(n15447), .Z(n15445) );
  OR U15494 ( .A(n15448), .B(n15449), .Z(n15447) );
  NAND U15495 ( .A(n15449), .B(n15448), .Z(n15444) );
  ANDN U15496 ( .B(B[248]), .A(n71), .Z(n15274) );
  XNOR U15497 ( .A(n15282), .B(n15450), .Z(n15275) );
  XNOR U15498 ( .A(n15281), .B(n15279), .Z(n15450) );
  AND U15499 ( .A(n15451), .B(n15452), .Z(n15279) );
  NANDN U15500 ( .A(n15453), .B(n15454), .Z(n15452) );
  NANDN U15501 ( .A(n15455), .B(n15456), .Z(n15454) );
  NANDN U15502 ( .A(n15456), .B(n15455), .Z(n15451) );
  ANDN U15503 ( .B(B[249]), .A(n72), .Z(n15281) );
  XNOR U15504 ( .A(n15289), .B(n15457), .Z(n15282) );
  XNOR U15505 ( .A(n15288), .B(n15286), .Z(n15457) );
  AND U15506 ( .A(n15458), .B(n15459), .Z(n15286) );
  NANDN U15507 ( .A(n15460), .B(n15461), .Z(n15459) );
  OR U15508 ( .A(n15462), .B(n15463), .Z(n15461) );
  NAND U15509 ( .A(n15463), .B(n15462), .Z(n15458) );
  ANDN U15510 ( .B(B[250]), .A(n73), .Z(n15288) );
  XNOR U15511 ( .A(n15296), .B(n15464), .Z(n15289) );
  XNOR U15512 ( .A(n15295), .B(n15293), .Z(n15464) );
  AND U15513 ( .A(n15465), .B(n15466), .Z(n15293) );
  NANDN U15514 ( .A(n15467), .B(n15468), .Z(n15466) );
  NANDN U15515 ( .A(n15469), .B(n15470), .Z(n15468) );
  NANDN U15516 ( .A(n15470), .B(n15469), .Z(n15465) );
  ANDN U15517 ( .B(B[251]), .A(n74), .Z(n15295) );
  XNOR U15518 ( .A(n15303), .B(n15471), .Z(n15296) );
  XNOR U15519 ( .A(n15302), .B(n15300), .Z(n15471) );
  AND U15520 ( .A(n15472), .B(n15473), .Z(n15300) );
  NANDN U15521 ( .A(n15474), .B(n15475), .Z(n15473) );
  OR U15522 ( .A(n15476), .B(n15477), .Z(n15475) );
  NAND U15523 ( .A(n15477), .B(n15476), .Z(n15472) );
  ANDN U15524 ( .B(B[252]), .A(n75), .Z(n15302) );
  XNOR U15525 ( .A(n15310), .B(n15478), .Z(n15303) );
  XNOR U15526 ( .A(n15309), .B(n15307), .Z(n15478) );
  AND U15527 ( .A(n15479), .B(n15480), .Z(n15307) );
  NANDN U15528 ( .A(n15481), .B(n15482), .Z(n15480) );
  NANDN U15529 ( .A(n15483), .B(n15484), .Z(n15482) );
  NANDN U15530 ( .A(n15484), .B(n15483), .Z(n15479) );
  ANDN U15531 ( .B(B[253]), .A(n76), .Z(n15309) );
  XOR U15532 ( .A(n15315), .B(n15485), .Z(n15310) );
  XOR U15533 ( .A(n15316), .B(n15317), .Z(n15485) );
  NAND U15534 ( .A(A[7]), .B(B[255]), .Z(n15317) );
  AND U15535 ( .A(B[254]), .B(A[8]), .Z(n15316) );
  NAND U15536 ( .A(n15486), .B(n15487), .Z(n15315) );
  NAND U15537 ( .A(n15488), .B(n15489), .Z(n15487) );
  NANDN U15538 ( .A(n15490), .B(n15491), .Z(n15488) );
  NANDN U15539 ( .A(n15491), .B(n15490), .Z(n15486) );
  NAND U15540 ( .A(n15492), .B(n15493), .Z(n272) );
  NANDN U15541 ( .A(n15494), .B(n15495), .Z(n15493) );
  OR U15542 ( .A(n15496), .B(n15497), .Z(n15495) );
  NAND U15543 ( .A(n15497), .B(n15496), .Z(n15492) );
  XOR U15544 ( .A(n13893), .B(n15498), .Z(\A1[25] ) );
  XNOR U15545 ( .A(n13892), .B(n13890), .Z(n15498) );
  AND U15546 ( .A(n15499), .B(n15500), .Z(n13890) );
  NAND U15547 ( .A(n15501), .B(n15502), .Z(n15500) );
  NANDN U15548 ( .A(n15503), .B(n15504), .Z(n15501) );
  NANDN U15549 ( .A(n15504), .B(n15503), .Z(n15499) );
  ANDN U15550 ( .B(B[0]), .A(n58), .Z(n13892) );
  XNOR U15551 ( .A(n13900), .B(n15505), .Z(n13893) );
  XNOR U15552 ( .A(n13899), .B(n13897), .Z(n15505) );
  AND U15553 ( .A(n15506), .B(n15507), .Z(n13897) );
  NANDN U15554 ( .A(n15508), .B(n15509), .Z(n15507) );
  OR U15555 ( .A(n15510), .B(n15511), .Z(n15509) );
  NAND U15556 ( .A(n15511), .B(n15510), .Z(n15506) );
  ANDN U15557 ( .B(B[1]), .A(n59), .Z(n13899) );
  XNOR U15558 ( .A(n13907), .B(n15512), .Z(n13900) );
  XNOR U15559 ( .A(n13906), .B(n13904), .Z(n15512) );
  AND U15560 ( .A(n15513), .B(n15514), .Z(n13904) );
  NANDN U15561 ( .A(n15515), .B(n15516), .Z(n15514) );
  NANDN U15562 ( .A(n15517), .B(n15518), .Z(n15516) );
  NANDN U15563 ( .A(n15518), .B(n15517), .Z(n15513) );
  ANDN U15564 ( .B(B[2]), .A(n60), .Z(n13906) );
  XNOR U15565 ( .A(n13914), .B(n15519), .Z(n13907) );
  XNOR U15566 ( .A(n13913), .B(n13911), .Z(n15519) );
  AND U15567 ( .A(n15520), .B(n15521), .Z(n13911) );
  NANDN U15568 ( .A(n15522), .B(n15523), .Z(n15521) );
  OR U15569 ( .A(n15524), .B(n15525), .Z(n15523) );
  NAND U15570 ( .A(n15525), .B(n15524), .Z(n15520) );
  ANDN U15571 ( .B(B[3]), .A(n61), .Z(n13913) );
  XNOR U15572 ( .A(n13921), .B(n15526), .Z(n13914) );
  XNOR U15573 ( .A(n13920), .B(n13918), .Z(n15526) );
  AND U15574 ( .A(n15527), .B(n15528), .Z(n13918) );
  NANDN U15575 ( .A(n15529), .B(n15530), .Z(n15528) );
  NANDN U15576 ( .A(n15531), .B(n15532), .Z(n15530) );
  NANDN U15577 ( .A(n15532), .B(n15531), .Z(n15527) );
  ANDN U15578 ( .B(B[4]), .A(n62), .Z(n13920) );
  XNOR U15579 ( .A(n13928), .B(n15533), .Z(n13921) );
  XNOR U15580 ( .A(n13927), .B(n13925), .Z(n15533) );
  AND U15581 ( .A(n15534), .B(n15535), .Z(n13925) );
  NANDN U15582 ( .A(n15536), .B(n15537), .Z(n15535) );
  OR U15583 ( .A(n15538), .B(n15539), .Z(n15537) );
  NAND U15584 ( .A(n15539), .B(n15538), .Z(n15534) );
  ANDN U15585 ( .B(B[5]), .A(n63), .Z(n13927) );
  XNOR U15586 ( .A(n13935), .B(n15540), .Z(n13928) );
  XNOR U15587 ( .A(n13934), .B(n13932), .Z(n15540) );
  AND U15588 ( .A(n15541), .B(n15542), .Z(n13932) );
  NANDN U15589 ( .A(n15543), .B(n15544), .Z(n15542) );
  NANDN U15590 ( .A(n15545), .B(n15546), .Z(n15544) );
  NANDN U15591 ( .A(n15546), .B(n15545), .Z(n15541) );
  ANDN U15592 ( .B(B[6]), .A(n64), .Z(n13934) );
  XNOR U15593 ( .A(n13942), .B(n15547), .Z(n13935) );
  XNOR U15594 ( .A(n13941), .B(n13939), .Z(n15547) );
  AND U15595 ( .A(n15548), .B(n15549), .Z(n13939) );
  NANDN U15596 ( .A(n15550), .B(n15551), .Z(n15549) );
  OR U15597 ( .A(n15552), .B(n15553), .Z(n15551) );
  NAND U15598 ( .A(n15553), .B(n15552), .Z(n15548) );
  ANDN U15599 ( .B(B[7]), .A(n65), .Z(n13941) );
  XNOR U15600 ( .A(n13949), .B(n15554), .Z(n13942) );
  XNOR U15601 ( .A(n13948), .B(n13946), .Z(n15554) );
  AND U15602 ( .A(n15555), .B(n15556), .Z(n13946) );
  NANDN U15603 ( .A(n15557), .B(n15558), .Z(n15556) );
  NANDN U15604 ( .A(n15559), .B(n15560), .Z(n15558) );
  NANDN U15605 ( .A(n15560), .B(n15559), .Z(n15555) );
  ANDN U15606 ( .B(B[8]), .A(n66), .Z(n13948) );
  XNOR U15607 ( .A(n13956), .B(n15561), .Z(n13949) );
  XNOR U15608 ( .A(n13955), .B(n13953), .Z(n15561) );
  AND U15609 ( .A(n15562), .B(n15563), .Z(n13953) );
  NANDN U15610 ( .A(n15564), .B(n15565), .Z(n15563) );
  OR U15611 ( .A(n15566), .B(n15567), .Z(n15565) );
  NAND U15612 ( .A(n15567), .B(n15566), .Z(n15562) );
  ANDN U15613 ( .B(B[9]), .A(n67), .Z(n13955) );
  XNOR U15614 ( .A(n13963), .B(n15568), .Z(n13956) );
  XNOR U15615 ( .A(n13962), .B(n13960), .Z(n15568) );
  AND U15616 ( .A(n15569), .B(n15570), .Z(n13960) );
  NANDN U15617 ( .A(n15571), .B(n15572), .Z(n15570) );
  NANDN U15618 ( .A(n15573), .B(n15574), .Z(n15572) );
  NANDN U15619 ( .A(n15574), .B(n15573), .Z(n15569) );
  ANDN U15620 ( .B(B[10]), .A(n68), .Z(n13962) );
  XNOR U15621 ( .A(n13970), .B(n15575), .Z(n13963) );
  XNOR U15622 ( .A(n13969), .B(n13967), .Z(n15575) );
  AND U15623 ( .A(n15576), .B(n15577), .Z(n13967) );
  NANDN U15624 ( .A(n15578), .B(n15579), .Z(n15577) );
  OR U15625 ( .A(n15580), .B(n15581), .Z(n15579) );
  NAND U15626 ( .A(n15581), .B(n15580), .Z(n15576) );
  ANDN U15627 ( .B(B[11]), .A(n69), .Z(n13969) );
  XNOR U15628 ( .A(n13977), .B(n15582), .Z(n13970) );
  XNOR U15629 ( .A(n13976), .B(n13974), .Z(n15582) );
  AND U15630 ( .A(n15583), .B(n15584), .Z(n13974) );
  NANDN U15631 ( .A(n15585), .B(n15586), .Z(n15584) );
  NANDN U15632 ( .A(n15587), .B(n15588), .Z(n15586) );
  NANDN U15633 ( .A(n15588), .B(n15587), .Z(n15583) );
  ANDN U15634 ( .B(B[12]), .A(n70), .Z(n13976) );
  XNOR U15635 ( .A(n13984), .B(n15589), .Z(n13977) );
  XNOR U15636 ( .A(n13983), .B(n13981), .Z(n15589) );
  AND U15637 ( .A(n15590), .B(n15591), .Z(n13981) );
  NANDN U15638 ( .A(n15592), .B(n15593), .Z(n15591) );
  OR U15639 ( .A(n15594), .B(n15595), .Z(n15593) );
  NAND U15640 ( .A(n15595), .B(n15594), .Z(n15590) );
  ANDN U15641 ( .B(B[13]), .A(n71), .Z(n13983) );
  XNOR U15642 ( .A(n13991), .B(n15596), .Z(n13984) );
  XNOR U15643 ( .A(n13990), .B(n13988), .Z(n15596) );
  AND U15644 ( .A(n15597), .B(n15598), .Z(n13988) );
  NANDN U15645 ( .A(n15599), .B(n15600), .Z(n15598) );
  NANDN U15646 ( .A(n15601), .B(n15602), .Z(n15600) );
  NANDN U15647 ( .A(n15602), .B(n15601), .Z(n15597) );
  ANDN U15648 ( .B(B[14]), .A(n72), .Z(n13990) );
  XNOR U15649 ( .A(n13998), .B(n15603), .Z(n13991) );
  XNOR U15650 ( .A(n13997), .B(n13995), .Z(n15603) );
  AND U15651 ( .A(n15604), .B(n15605), .Z(n13995) );
  NANDN U15652 ( .A(n15606), .B(n15607), .Z(n15605) );
  OR U15653 ( .A(n15608), .B(n15609), .Z(n15607) );
  NAND U15654 ( .A(n15609), .B(n15608), .Z(n15604) );
  ANDN U15655 ( .B(B[15]), .A(n73), .Z(n13997) );
  XNOR U15656 ( .A(n14005), .B(n15610), .Z(n13998) );
  XNOR U15657 ( .A(n14004), .B(n14002), .Z(n15610) );
  AND U15658 ( .A(n15611), .B(n15612), .Z(n14002) );
  NANDN U15659 ( .A(n15613), .B(n15614), .Z(n15612) );
  NANDN U15660 ( .A(n15615), .B(n15616), .Z(n15614) );
  NANDN U15661 ( .A(n15616), .B(n15615), .Z(n15611) );
  ANDN U15662 ( .B(B[16]), .A(n74), .Z(n14004) );
  XNOR U15663 ( .A(n14012), .B(n15617), .Z(n14005) );
  XNOR U15664 ( .A(n14011), .B(n14009), .Z(n15617) );
  AND U15665 ( .A(n15618), .B(n15619), .Z(n14009) );
  NANDN U15666 ( .A(n15620), .B(n15621), .Z(n15619) );
  OR U15667 ( .A(n15622), .B(n15623), .Z(n15621) );
  NAND U15668 ( .A(n15623), .B(n15622), .Z(n15618) );
  ANDN U15669 ( .B(B[17]), .A(n75), .Z(n14011) );
  XNOR U15670 ( .A(n14019), .B(n15624), .Z(n14012) );
  XNOR U15671 ( .A(n14018), .B(n14016), .Z(n15624) );
  AND U15672 ( .A(n15625), .B(n15626), .Z(n14016) );
  NANDN U15673 ( .A(n15627), .B(n15628), .Z(n15626) );
  NANDN U15674 ( .A(n15629), .B(n15630), .Z(n15628) );
  NANDN U15675 ( .A(n15630), .B(n15629), .Z(n15625) );
  ANDN U15676 ( .B(B[18]), .A(n76), .Z(n14018) );
  XNOR U15677 ( .A(n14026), .B(n15631), .Z(n14019) );
  XNOR U15678 ( .A(n14025), .B(n14023), .Z(n15631) );
  AND U15679 ( .A(n15632), .B(n15633), .Z(n14023) );
  NANDN U15680 ( .A(n15634), .B(n15635), .Z(n15633) );
  OR U15681 ( .A(n15636), .B(n15637), .Z(n15635) );
  NAND U15682 ( .A(n15637), .B(n15636), .Z(n15632) );
  ANDN U15683 ( .B(B[19]), .A(n77), .Z(n14025) );
  XNOR U15684 ( .A(n14033), .B(n15638), .Z(n14026) );
  XNOR U15685 ( .A(n14032), .B(n14030), .Z(n15638) );
  AND U15686 ( .A(n15639), .B(n15640), .Z(n14030) );
  NANDN U15687 ( .A(n15641), .B(n15642), .Z(n15640) );
  NANDN U15688 ( .A(n15643), .B(n15644), .Z(n15642) );
  NANDN U15689 ( .A(n15644), .B(n15643), .Z(n15639) );
  ANDN U15690 ( .B(B[20]), .A(n78), .Z(n14032) );
  XNOR U15691 ( .A(n14040), .B(n15645), .Z(n14033) );
  XNOR U15692 ( .A(n14039), .B(n14037), .Z(n15645) );
  AND U15693 ( .A(n15646), .B(n15647), .Z(n14037) );
  NANDN U15694 ( .A(n15648), .B(n15649), .Z(n15647) );
  OR U15695 ( .A(n15650), .B(n15651), .Z(n15649) );
  NAND U15696 ( .A(n15651), .B(n15650), .Z(n15646) );
  ANDN U15697 ( .B(B[21]), .A(n79), .Z(n14039) );
  XNOR U15698 ( .A(n14047), .B(n15652), .Z(n14040) );
  XNOR U15699 ( .A(n14046), .B(n14044), .Z(n15652) );
  AND U15700 ( .A(n15653), .B(n15654), .Z(n14044) );
  NANDN U15701 ( .A(n15655), .B(n15656), .Z(n15654) );
  NANDN U15702 ( .A(n15657), .B(n15658), .Z(n15656) );
  NANDN U15703 ( .A(n15658), .B(n15657), .Z(n15653) );
  ANDN U15704 ( .B(B[22]), .A(n80), .Z(n14046) );
  XNOR U15705 ( .A(n14054), .B(n15659), .Z(n14047) );
  XNOR U15706 ( .A(n14053), .B(n14051), .Z(n15659) );
  AND U15707 ( .A(n15660), .B(n15661), .Z(n14051) );
  NANDN U15708 ( .A(n15662), .B(n15663), .Z(n15661) );
  OR U15709 ( .A(n15664), .B(n15665), .Z(n15663) );
  NAND U15710 ( .A(n15665), .B(n15664), .Z(n15660) );
  ANDN U15711 ( .B(B[23]), .A(n81), .Z(n14053) );
  XNOR U15712 ( .A(n14061), .B(n15666), .Z(n14054) );
  XNOR U15713 ( .A(n14060), .B(n14058), .Z(n15666) );
  AND U15714 ( .A(n15667), .B(n15668), .Z(n14058) );
  NANDN U15715 ( .A(n15669), .B(n15670), .Z(n15668) );
  NAND U15716 ( .A(n15671), .B(n15672), .Z(n15670) );
  ANDN U15717 ( .B(B[24]), .A(n82), .Z(n14060) );
  XOR U15718 ( .A(n14067), .B(n15673), .Z(n14061) );
  XNOR U15719 ( .A(n14065), .B(n14068), .Z(n15673) );
  NAND U15720 ( .A(A[2]), .B(B[25]), .Z(n14068) );
  NANDN U15721 ( .A(n15674), .B(n15675), .Z(n14065) );
  AND U15722 ( .A(A[0]), .B(B[26]), .Z(n15675) );
  XNOR U15723 ( .A(n14070), .B(n15676), .Z(n14067) );
  NAND U15724 ( .A(A[0]), .B(B[27]), .Z(n15676) );
  NAND U15725 ( .A(B[26]), .B(A[1]), .Z(n14070) );
  XOR U15726 ( .A(n274), .B(n273), .Z(\A1[259] ) );
  XOR U15727 ( .A(n15497), .B(n15677), .Z(n273) );
  XNOR U15728 ( .A(n15496), .B(n15494), .Z(n15677) );
  AND U15729 ( .A(n15678), .B(n15679), .Z(n15494) );
  NANDN U15730 ( .A(n15680), .B(n15681), .Z(n15679) );
  OR U15731 ( .A(n15682), .B(n15683), .Z(n15681) );
  NAND U15732 ( .A(n15683), .B(n15682), .Z(n15678) );
  ANDN U15733 ( .B(B[230]), .A(n54), .Z(n15496) );
  XNOR U15734 ( .A(n15330), .B(n15684), .Z(n15497) );
  XNOR U15735 ( .A(n15329), .B(n15327), .Z(n15684) );
  AND U15736 ( .A(n15685), .B(n15686), .Z(n15327) );
  NANDN U15737 ( .A(n15687), .B(n15688), .Z(n15686) );
  NANDN U15738 ( .A(n15689), .B(n15690), .Z(n15688) );
  NANDN U15739 ( .A(n15690), .B(n15689), .Z(n15685) );
  ANDN U15740 ( .B(B[231]), .A(n55), .Z(n15329) );
  XNOR U15741 ( .A(n15337), .B(n15691), .Z(n15330) );
  XNOR U15742 ( .A(n15336), .B(n15334), .Z(n15691) );
  AND U15743 ( .A(n15692), .B(n15693), .Z(n15334) );
  NANDN U15744 ( .A(n15694), .B(n15695), .Z(n15693) );
  OR U15745 ( .A(n15696), .B(n15697), .Z(n15695) );
  NAND U15746 ( .A(n15697), .B(n15696), .Z(n15692) );
  ANDN U15747 ( .B(B[232]), .A(n56), .Z(n15336) );
  XNOR U15748 ( .A(n15344), .B(n15698), .Z(n15337) );
  XNOR U15749 ( .A(n15343), .B(n15341), .Z(n15698) );
  AND U15750 ( .A(n15699), .B(n15700), .Z(n15341) );
  NANDN U15751 ( .A(n15701), .B(n15702), .Z(n15700) );
  NANDN U15752 ( .A(n15703), .B(n15704), .Z(n15702) );
  NANDN U15753 ( .A(n15704), .B(n15703), .Z(n15699) );
  ANDN U15754 ( .B(B[233]), .A(n57), .Z(n15343) );
  XNOR U15755 ( .A(n15351), .B(n15705), .Z(n15344) );
  XNOR U15756 ( .A(n15350), .B(n15348), .Z(n15705) );
  AND U15757 ( .A(n15706), .B(n15707), .Z(n15348) );
  NANDN U15758 ( .A(n15708), .B(n15709), .Z(n15707) );
  OR U15759 ( .A(n15710), .B(n15711), .Z(n15709) );
  NAND U15760 ( .A(n15711), .B(n15710), .Z(n15706) );
  ANDN U15761 ( .B(B[234]), .A(n58), .Z(n15350) );
  XNOR U15762 ( .A(n15358), .B(n15712), .Z(n15351) );
  XNOR U15763 ( .A(n15357), .B(n15355), .Z(n15712) );
  AND U15764 ( .A(n15713), .B(n15714), .Z(n15355) );
  NANDN U15765 ( .A(n15715), .B(n15716), .Z(n15714) );
  NANDN U15766 ( .A(n15717), .B(n15718), .Z(n15716) );
  NANDN U15767 ( .A(n15718), .B(n15717), .Z(n15713) );
  ANDN U15768 ( .B(B[235]), .A(n59), .Z(n15357) );
  XNOR U15769 ( .A(n15365), .B(n15719), .Z(n15358) );
  XNOR U15770 ( .A(n15364), .B(n15362), .Z(n15719) );
  AND U15771 ( .A(n15720), .B(n15721), .Z(n15362) );
  NANDN U15772 ( .A(n15722), .B(n15723), .Z(n15721) );
  OR U15773 ( .A(n15724), .B(n15725), .Z(n15723) );
  NAND U15774 ( .A(n15725), .B(n15724), .Z(n15720) );
  ANDN U15775 ( .B(B[236]), .A(n60), .Z(n15364) );
  XNOR U15776 ( .A(n15372), .B(n15726), .Z(n15365) );
  XNOR U15777 ( .A(n15371), .B(n15369), .Z(n15726) );
  AND U15778 ( .A(n15727), .B(n15728), .Z(n15369) );
  NANDN U15779 ( .A(n15729), .B(n15730), .Z(n15728) );
  NANDN U15780 ( .A(n15731), .B(n15732), .Z(n15730) );
  NANDN U15781 ( .A(n15732), .B(n15731), .Z(n15727) );
  ANDN U15782 ( .B(B[237]), .A(n61), .Z(n15371) );
  XNOR U15783 ( .A(n15379), .B(n15733), .Z(n15372) );
  XNOR U15784 ( .A(n15378), .B(n15376), .Z(n15733) );
  AND U15785 ( .A(n15734), .B(n15735), .Z(n15376) );
  NANDN U15786 ( .A(n15736), .B(n15737), .Z(n15735) );
  OR U15787 ( .A(n15738), .B(n15739), .Z(n15737) );
  NAND U15788 ( .A(n15739), .B(n15738), .Z(n15734) );
  ANDN U15789 ( .B(B[238]), .A(n62), .Z(n15378) );
  XNOR U15790 ( .A(n15386), .B(n15740), .Z(n15379) );
  XNOR U15791 ( .A(n15385), .B(n15383), .Z(n15740) );
  AND U15792 ( .A(n15741), .B(n15742), .Z(n15383) );
  NANDN U15793 ( .A(n15743), .B(n15744), .Z(n15742) );
  NANDN U15794 ( .A(n15745), .B(n15746), .Z(n15744) );
  NANDN U15795 ( .A(n15746), .B(n15745), .Z(n15741) );
  ANDN U15796 ( .B(B[239]), .A(n63), .Z(n15385) );
  XNOR U15797 ( .A(n15393), .B(n15747), .Z(n15386) );
  XNOR U15798 ( .A(n15392), .B(n15390), .Z(n15747) );
  AND U15799 ( .A(n15748), .B(n15749), .Z(n15390) );
  NANDN U15800 ( .A(n15750), .B(n15751), .Z(n15749) );
  OR U15801 ( .A(n15752), .B(n15753), .Z(n15751) );
  NAND U15802 ( .A(n15753), .B(n15752), .Z(n15748) );
  ANDN U15803 ( .B(B[240]), .A(n64), .Z(n15392) );
  XNOR U15804 ( .A(n15400), .B(n15754), .Z(n15393) );
  XNOR U15805 ( .A(n15399), .B(n15397), .Z(n15754) );
  AND U15806 ( .A(n15755), .B(n15756), .Z(n15397) );
  NANDN U15807 ( .A(n15757), .B(n15758), .Z(n15756) );
  NANDN U15808 ( .A(n15759), .B(n15760), .Z(n15758) );
  NANDN U15809 ( .A(n15760), .B(n15759), .Z(n15755) );
  ANDN U15810 ( .B(B[241]), .A(n65), .Z(n15399) );
  XNOR U15811 ( .A(n15407), .B(n15761), .Z(n15400) );
  XNOR U15812 ( .A(n15406), .B(n15404), .Z(n15761) );
  AND U15813 ( .A(n15762), .B(n15763), .Z(n15404) );
  NANDN U15814 ( .A(n15764), .B(n15765), .Z(n15763) );
  OR U15815 ( .A(n15766), .B(n15767), .Z(n15765) );
  NAND U15816 ( .A(n15767), .B(n15766), .Z(n15762) );
  ANDN U15817 ( .B(B[242]), .A(n66), .Z(n15406) );
  XNOR U15818 ( .A(n15414), .B(n15768), .Z(n15407) );
  XNOR U15819 ( .A(n15413), .B(n15411), .Z(n15768) );
  AND U15820 ( .A(n15769), .B(n15770), .Z(n15411) );
  NANDN U15821 ( .A(n15771), .B(n15772), .Z(n15770) );
  NANDN U15822 ( .A(n15773), .B(n15774), .Z(n15772) );
  NANDN U15823 ( .A(n15774), .B(n15773), .Z(n15769) );
  ANDN U15824 ( .B(B[243]), .A(n67), .Z(n15413) );
  XNOR U15825 ( .A(n15421), .B(n15775), .Z(n15414) );
  XNOR U15826 ( .A(n15420), .B(n15418), .Z(n15775) );
  AND U15827 ( .A(n15776), .B(n15777), .Z(n15418) );
  NANDN U15828 ( .A(n15778), .B(n15779), .Z(n15777) );
  OR U15829 ( .A(n15780), .B(n15781), .Z(n15779) );
  NAND U15830 ( .A(n15781), .B(n15780), .Z(n15776) );
  ANDN U15831 ( .B(B[244]), .A(n68), .Z(n15420) );
  XNOR U15832 ( .A(n15428), .B(n15782), .Z(n15421) );
  XNOR U15833 ( .A(n15427), .B(n15425), .Z(n15782) );
  AND U15834 ( .A(n15783), .B(n15784), .Z(n15425) );
  NANDN U15835 ( .A(n15785), .B(n15786), .Z(n15784) );
  NANDN U15836 ( .A(n15787), .B(n15788), .Z(n15786) );
  NANDN U15837 ( .A(n15788), .B(n15787), .Z(n15783) );
  ANDN U15838 ( .B(B[245]), .A(n69), .Z(n15427) );
  XNOR U15839 ( .A(n15435), .B(n15789), .Z(n15428) );
  XNOR U15840 ( .A(n15434), .B(n15432), .Z(n15789) );
  AND U15841 ( .A(n15790), .B(n15791), .Z(n15432) );
  NANDN U15842 ( .A(n15792), .B(n15793), .Z(n15791) );
  OR U15843 ( .A(n15794), .B(n15795), .Z(n15793) );
  NAND U15844 ( .A(n15795), .B(n15794), .Z(n15790) );
  ANDN U15845 ( .B(B[246]), .A(n70), .Z(n15434) );
  XNOR U15846 ( .A(n15442), .B(n15796), .Z(n15435) );
  XNOR U15847 ( .A(n15441), .B(n15439), .Z(n15796) );
  AND U15848 ( .A(n15797), .B(n15798), .Z(n15439) );
  NANDN U15849 ( .A(n15799), .B(n15800), .Z(n15798) );
  NANDN U15850 ( .A(n15801), .B(n15802), .Z(n15800) );
  NANDN U15851 ( .A(n15802), .B(n15801), .Z(n15797) );
  ANDN U15852 ( .B(B[247]), .A(n71), .Z(n15441) );
  XNOR U15853 ( .A(n15449), .B(n15803), .Z(n15442) );
  XNOR U15854 ( .A(n15448), .B(n15446), .Z(n15803) );
  AND U15855 ( .A(n15804), .B(n15805), .Z(n15446) );
  NANDN U15856 ( .A(n15806), .B(n15807), .Z(n15805) );
  OR U15857 ( .A(n15808), .B(n15809), .Z(n15807) );
  NAND U15858 ( .A(n15809), .B(n15808), .Z(n15804) );
  ANDN U15859 ( .B(B[248]), .A(n72), .Z(n15448) );
  XNOR U15860 ( .A(n15456), .B(n15810), .Z(n15449) );
  XNOR U15861 ( .A(n15455), .B(n15453), .Z(n15810) );
  AND U15862 ( .A(n15811), .B(n15812), .Z(n15453) );
  NANDN U15863 ( .A(n15813), .B(n15814), .Z(n15812) );
  NANDN U15864 ( .A(n15815), .B(n15816), .Z(n15814) );
  NANDN U15865 ( .A(n15816), .B(n15815), .Z(n15811) );
  ANDN U15866 ( .B(B[249]), .A(n73), .Z(n15455) );
  XNOR U15867 ( .A(n15463), .B(n15817), .Z(n15456) );
  XNOR U15868 ( .A(n15462), .B(n15460), .Z(n15817) );
  AND U15869 ( .A(n15818), .B(n15819), .Z(n15460) );
  NANDN U15870 ( .A(n15820), .B(n15821), .Z(n15819) );
  OR U15871 ( .A(n15822), .B(n15823), .Z(n15821) );
  NAND U15872 ( .A(n15823), .B(n15822), .Z(n15818) );
  ANDN U15873 ( .B(B[250]), .A(n74), .Z(n15462) );
  XNOR U15874 ( .A(n15470), .B(n15824), .Z(n15463) );
  XNOR U15875 ( .A(n15469), .B(n15467), .Z(n15824) );
  AND U15876 ( .A(n15825), .B(n15826), .Z(n15467) );
  NANDN U15877 ( .A(n15827), .B(n15828), .Z(n15826) );
  NANDN U15878 ( .A(n15829), .B(n15830), .Z(n15828) );
  NANDN U15879 ( .A(n15830), .B(n15829), .Z(n15825) );
  ANDN U15880 ( .B(B[251]), .A(n75), .Z(n15469) );
  XNOR U15881 ( .A(n15477), .B(n15831), .Z(n15470) );
  XNOR U15882 ( .A(n15476), .B(n15474), .Z(n15831) );
  AND U15883 ( .A(n15832), .B(n15833), .Z(n15474) );
  NANDN U15884 ( .A(n15834), .B(n15835), .Z(n15833) );
  OR U15885 ( .A(n15836), .B(n15837), .Z(n15835) );
  NAND U15886 ( .A(n15837), .B(n15836), .Z(n15832) );
  ANDN U15887 ( .B(B[252]), .A(n76), .Z(n15476) );
  XNOR U15888 ( .A(n15484), .B(n15838), .Z(n15477) );
  XNOR U15889 ( .A(n15483), .B(n15481), .Z(n15838) );
  AND U15890 ( .A(n15839), .B(n15840), .Z(n15481) );
  NANDN U15891 ( .A(n15841), .B(n15842), .Z(n15840) );
  NANDN U15892 ( .A(n15843), .B(n15844), .Z(n15842) );
  NANDN U15893 ( .A(n15844), .B(n15843), .Z(n15839) );
  ANDN U15894 ( .B(B[253]), .A(n77), .Z(n15483) );
  XOR U15895 ( .A(n15489), .B(n15845), .Z(n15484) );
  XOR U15896 ( .A(n15490), .B(n15491), .Z(n15845) );
  NAND U15897 ( .A(A[6]), .B(B[255]), .Z(n15491) );
  AND U15898 ( .A(B[254]), .B(A[7]), .Z(n15490) );
  NAND U15899 ( .A(n15846), .B(n15847), .Z(n15489) );
  NAND U15900 ( .A(n15848), .B(n15849), .Z(n15847) );
  NANDN U15901 ( .A(n15850), .B(n15851), .Z(n15848) );
  NANDN U15902 ( .A(n15851), .B(n15850), .Z(n15846) );
  NAND U15903 ( .A(n15852), .B(n15853), .Z(n274) );
  NANDN U15904 ( .A(n15854), .B(n15855), .Z(n15853) );
  NAND U15905 ( .A(n15857), .B(n15856), .Z(n15852) );
  XOR U15906 ( .A(n276), .B(n275), .Z(\A1[258] ) );
  XOR U15907 ( .A(n15857), .B(n15858), .Z(n275) );
  XNOR U15908 ( .A(n15856), .B(n15854), .Z(n15858) );
  AND U15909 ( .A(n15859), .B(n15860), .Z(n15854) );
  NANDN U15910 ( .A(n15861), .B(n15862), .Z(n15860) );
  NANDN U15911 ( .A(n15863), .B(n15864), .Z(n15862) );
  NANDN U15912 ( .A(n15864), .B(n15863), .Z(n15859) );
  ANDN U15913 ( .B(B[229]), .A(n54), .Z(n15856) );
  XOR U15914 ( .A(n15683), .B(n15865), .Z(n15857) );
  XNOR U15915 ( .A(n15682), .B(n15680), .Z(n15865) );
  AND U15916 ( .A(n15866), .B(n15867), .Z(n15680) );
  NANDN U15917 ( .A(n15868), .B(n15869), .Z(n15867) );
  OR U15918 ( .A(n15870), .B(n15871), .Z(n15869) );
  NAND U15919 ( .A(n15871), .B(n15870), .Z(n15866) );
  ANDN U15920 ( .B(B[230]), .A(n55), .Z(n15682) );
  XNOR U15921 ( .A(n15690), .B(n15872), .Z(n15683) );
  XNOR U15922 ( .A(n15689), .B(n15687), .Z(n15872) );
  AND U15923 ( .A(n15873), .B(n15874), .Z(n15687) );
  NANDN U15924 ( .A(n15875), .B(n15876), .Z(n15874) );
  NANDN U15925 ( .A(n15877), .B(n15878), .Z(n15876) );
  NANDN U15926 ( .A(n15878), .B(n15877), .Z(n15873) );
  ANDN U15927 ( .B(B[231]), .A(n56), .Z(n15689) );
  XNOR U15928 ( .A(n15697), .B(n15879), .Z(n15690) );
  XNOR U15929 ( .A(n15696), .B(n15694), .Z(n15879) );
  AND U15930 ( .A(n15880), .B(n15881), .Z(n15694) );
  NANDN U15931 ( .A(n15882), .B(n15883), .Z(n15881) );
  OR U15932 ( .A(n15884), .B(n15885), .Z(n15883) );
  NAND U15933 ( .A(n15885), .B(n15884), .Z(n15880) );
  ANDN U15934 ( .B(B[232]), .A(n57), .Z(n15696) );
  XNOR U15935 ( .A(n15704), .B(n15886), .Z(n15697) );
  XNOR U15936 ( .A(n15703), .B(n15701), .Z(n15886) );
  AND U15937 ( .A(n15887), .B(n15888), .Z(n15701) );
  NANDN U15938 ( .A(n15889), .B(n15890), .Z(n15888) );
  NANDN U15939 ( .A(n15891), .B(n15892), .Z(n15890) );
  NANDN U15940 ( .A(n15892), .B(n15891), .Z(n15887) );
  ANDN U15941 ( .B(B[233]), .A(n58), .Z(n15703) );
  XNOR U15942 ( .A(n15711), .B(n15893), .Z(n15704) );
  XNOR U15943 ( .A(n15710), .B(n15708), .Z(n15893) );
  AND U15944 ( .A(n15894), .B(n15895), .Z(n15708) );
  NANDN U15945 ( .A(n15896), .B(n15897), .Z(n15895) );
  OR U15946 ( .A(n15898), .B(n15899), .Z(n15897) );
  NAND U15947 ( .A(n15899), .B(n15898), .Z(n15894) );
  ANDN U15948 ( .B(B[234]), .A(n59), .Z(n15710) );
  XNOR U15949 ( .A(n15718), .B(n15900), .Z(n15711) );
  XNOR U15950 ( .A(n15717), .B(n15715), .Z(n15900) );
  AND U15951 ( .A(n15901), .B(n15902), .Z(n15715) );
  NANDN U15952 ( .A(n15903), .B(n15904), .Z(n15902) );
  NANDN U15953 ( .A(n15905), .B(n15906), .Z(n15904) );
  NANDN U15954 ( .A(n15906), .B(n15905), .Z(n15901) );
  ANDN U15955 ( .B(B[235]), .A(n60), .Z(n15717) );
  XNOR U15956 ( .A(n15725), .B(n15907), .Z(n15718) );
  XNOR U15957 ( .A(n15724), .B(n15722), .Z(n15907) );
  AND U15958 ( .A(n15908), .B(n15909), .Z(n15722) );
  NANDN U15959 ( .A(n15910), .B(n15911), .Z(n15909) );
  OR U15960 ( .A(n15912), .B(n15913), .Z(n15911) );
  NAND U15961 ( .A(n15913), .B(n15912), .Z(n15908) );
  ANDN U15962 ( .B(B[236]), .A(n61), .Z(n15724) );
  XNOR U15963 ( .A(n15732), .B(n15914), .Z(n15725) );
  XNOR U15964 ( .A(n15731), .B(n15729), .Z(n15914) );
  AND U15965 ( .A(n15915), .B(n15916), .Z(n15729) );
  NANDN U15966 ( .A(n15917), .B(n15918), .Z(n15916) );
  NANDN U15967 ( .A(n15919), .B(n15920), .Z(n15918) );
  NANDN U15968 ( .A(n15920), .B(n15919), .Z(n15915) );
  ANDN U15969 ( .B(B[237]), .A(n62), .Z(n15731) );
  XNOR U15970 ( .A(n15739), .B(n15921), .Z(n15732) );
  XNOR U15971 ( .A(n15738), .B(n15736), .Z(n15921) );
  AND U15972 ( .A(n15922), .B(n15923), .Z(n15736) );
  NANDN U15973 ( .A(n15924), .B(n15925), .Z(n15923) );
  OR U15974 ( .A(n15926), .B(n15927), .Z(n15925) );
  NAND U15975 ( .A(n15927), .B(n15926), .Z(n15922) );
  ANDN U15976 ( .B(B[238]), .A(n63), .Z(n15738) );
  XNOR U15977 ( .A(n15746), .B(n15928), .Z(n15739) );
  XNOR U15978 ( .A(n15745), .B(n15743), .Z(n15928) );
  AND U15979 ( .A(n15929), .B(n15930), .Z(n15743) );
  NANDN U15980 ( .A(n15931), .B(n15932), .Z(n15930) );
  NANDN U15981 ( .A(n15933), .B(n15934), .Z(n15932) );
  NANDN U15982 ( .A(n15934), .B(n15933), .Z(n15929) );
  ANDN U15983 ( .B(B[239]), .A(n64), .Z(n15745) );
  XNOR U15984 ( .A(n15753), .B(n15935), .Z(n15746) );
  XNOR U15985 ( .A(n15752), .B(n15750), .Z(n15935) );
  AND U15986 ( .A(n15936), .B(n15937), .Z(n15750) );
  NANDN U15987 ( .A(n15938), .B(n15939), .Z(n15937) );
  OR U15988 ( .A(n15940), .B(n15941), .Z(n15939) );
  NAND U15989 ( .A(n15941), .B(n15940), .Z(n15936) );
  ANDN U15990 ( .B(B[240]), .A(n65), .Z(n15752) );
  XNOR U15991 ( .A(n15760), .B(n15942), .Z(n15753) );
  XNOR U15992 ( .A(n15759), .B(n15757), .Z(n15942) );
  AND U15993 ( .A(n15943), .B(n15944), .Z(n15757) );
  NANDN U15994 ( .A(n15945), .B(n15946), .Z(n15944) );
  NANDN U15995 ( .A(n15947), .B(n15948), .Z(n15946) );
  NANDN U15996 ( .A(n15948), .B(n15947), .Z(n15943) );
  ANDN U15997 ( .B(B[241]), .A(n66), .Z(n15759) );
  XNOR U15998 ( .A(n15767), .B(n15949), .Z(n15760) );
  XNOR U15999 ( .A(n15766), .B(n15764), .Z(n15949) );
  AND U16000 ( .A(n15950), .B(n15951), .Z(n15764) );
  NANDN U16001 ( .A(n15952), .B(n15953), .Z(n15951) );
  OR U16002 ( .A(n15954), .B(n15955), .Z(n15953) );
  NAND U16003 ( .A(n15955), .B(n15954), .Z(n15950) );
  ANDN U16004 ( .B(B[242]), .A(n67), .Z(n15766) );
  XNOR U16005 ( .A(n15774), .B(n15956), .Z(n15767) );
  XNOR U16006 ( .A(n15773), .B(n15771), .Z(n15956) );
  AND U16007 ( .A(n15957), .B(n15958), .Z(n15771) );
  NANDN U16008 ( .A(n15959), .B(n15960), .Z(n15958) );
  NANDN U16009 ( .A(n15961), .B(n15962), .Z(n15960) );
  NANDN U16010 ( .A(n15962), .B(n15961), .Z(n15957) );
  ANDN U16011 ( .B(B[243]), .A(n68), .Z(n15773) );
  XNOR U16012 ( .A(n15781), .B(n15963), .Z(n15774) );
  XNOR U16013 ( .A(n15780), .B(n15778), .Z(n15963) );
  AND U16014 ( .A(n15964), .B(n15965), .Z(n15778) );
  NANDN U16015 ( .A(n15966), .B(n15967), .Z(n15965) );
  OR U16016 ( .A(n15968), .B(n15969), .Z(n15967) );
  NAND U16017 ( .A(n15969), .B(n15968), .Z(n15964) );
  ANDN U16018 ( .B(B[244]), .A(n69), .Z(n15780) );
  XNOR U16019 ( .A(n15788), .B(n15970), .Z(n15781) );
  XNOR U16020 ( .A(n15787), .B(n15785), .Z(n15970) );
  AND U16021 ( .A(n15971), .B(n15972), .Z(n15785) );
  NANDN U16022 ( .A(n15973), .B(n15974), .Z(n15972) );
  NANDN U16023 ( .A(n15975), .B(n15976), .Z(n15974) );
  NANDN U16024 ( .A(n15976), .B(n15975), .Z(n15971) );
  ANDN U16025 ( .B(B[245]), .A(n70), .Z(n15787) );
  XNOR U16026 ( .A(n15795), .B(n15977), .Z(n15788) );
  XNOR U16027 ( .A(n15794), .B(n15792), .Z(n15977) );
  AND U16028 ( .A(n15978), .B(n15979), .Z(n15792) );
  NANDN U16029 ( .A(n15980), .B(n15981), .Z(n15979) );
  OR U16030 ( .A(n15982), .B(n15983), .Z(n15981) );
  NAND U16031 ( .A(n15983), .B(n15982), .Z(n15978) );
  ANDN U16032 ( .B(B[246]), .A(n71), .Z(n15794) );
  XNOR U16033 ( .A(n15802), .B(n15984), .Z(n15795) );
  XNOR U16034 ( .A(n15801), .B(n15799), .Z(n15984) );
  AND U16035 ( .A(n15985), .B(n15986), .Z(n15799) );
  NANDN U16036 ( .A(n15987), .B(n15988), .Z(n15986) );
  NANDN U16037 ( .A(n15989), .B(n15990), .Z(n15988) );
  NANDN U16038 ( .A(n15990), .B(n15989), .Z(n15985) );
  ANDN U16039 ( .B(B[247]), .A(n72), .Z(n15801) );
  XNOR U16040 ( .A(n15809), .B(n15991), .Z(n15802) );
  XNOR U16041 ( .A(n15808), .B(n15806), .Z(n15991) );
  AND U16042 ( .A(n15992), .B(n15993), .Z(n15806) );
  NANDN U16043 ( .A(n15994), .B(n15995), .Z(n15993) );
  OR U16044 ( .A(n15996), .B(n15997), .Z(n15995) );
  NAND U16045 ( .A(n15997), .B(n15996), .Z(n15992) );
  ANDN U16046 ( .B(B[248]), .A(n73), .Z(n15808) );
  XNOR U16047 ( .A(n15816), .B(n15998), .Z(n15809) );
  XNOR U16048 ( .A(n15815), .B(n15813), .Z(n15998) );
  AND U16049 ( .A(n15999), .B(n16000), .Z(n15813) );
  NANDN U16050 ( .A(n16001), .B(n16002), .Z(n16000) );
  NANDN U16051 ( .A(n16003), .B(n16004), .Z(n16002) );
  NANDN U16052 ( .A(n16004), .B(n16003), .Z(n15999) );
  ANDN U16053 ( .B(B[249]), .A(n74), .Z(n15815) );
  XNOR U16054 ( .A(n15823), .B(n16005), .Z(n15816) );
  XNOR U16055 ( .A(n15822), .B(n15820), .Z(n16005) );
  AND U16056 ( .A(n16006), .B(n16007), .Z(n15820) );
  NANDN U16057 ( .A(n16008), .B(n16009), .Z(n16007) );
  OR U16058 ( .A(n16010), .B(n16011), .Z(n16009) );
  NAND U16059 ( .A(n16011), .B(n16010), .Z(n16006) );
  ANDN U16060 ( .B(B[250]), .A(n75), .Z(n15822) );
  XNOR U16061 ( .A(n15830), .B(n16012), .Z(n15823) );
  XNOR U16062 ( .A(n15829), .B(n15827), .Z(n16012) );
  AND U16063 ( .A(n16013), .B(n16014), .Z(n15827) );
  NANDN U16064 ( .A(n16015), .B(n16016), .Z(n16014) );
  NANDN U16065 ( .A(n16017), .B(n16018), .Z(n16016) );
  NANDN U16066 ( .A(n16018), .B(n16017), .Z(n16013) );
  ANDN U16067 ( .B(B[251]), .A(n76), .Z(n15829) );
  XNOR U16068 ( .A(n15837), .B(n16019), .Z(n15830) );
  XNOR U16069 ( .A(n15836), .B(n15834), .Z(n16019) );
  AND U16070 ( .A(n16020), .B(n16021), .Z(n15834) );
  NANDN U16071 ( .A(n16022), .B(n16023), .Z(n16021) );
  OR U16072 ( .A(n16024), .B(n16025), .Z(n16023) );
  NAND U16073 ( .A(n16025), .B(n16024), .Z(n16020) );
  ANDN U16074 ( .B(B[252]), .A(n77), .Z(n15836) );
  XNOR U16075 ( .A(n15844), .B(n16026), .Z(n15837) );
  XNOR U16076 ( .A(n15843), .B(n15841), .Z(n16026) );
  AND U16077 ( .A(n16027), .B(n16028), .Z(n15841) );
  NANDN U16078 ( .A(n16029), .B(n16030), .Z(n16028) );
  NANDN U16079 ( .A(n16031), .B(n16032), .Z(n16030) );
  NANDN U16080 ( .A(n16032), .B(n16031), .Z(n16027) );
  ANDN U16081 ( .B(B[253]), .A(n78), .Z(n15843) );
  XOR U16082 ( .A(n15849), .B(n16033), .Z(n15844) );
  XOR U16083 ( .A(n15850), .B(n15851), .Z(n16033) );
  NAND U16084 ( .A(A[5]), .B(B[255]), .Z(n15851) );
  AND U16085 ( .A(B[254]), .B(A[6]), .Z(n15850) );
  NAND U16086 ( .A(n16034), .B(n16035), .Z(n15849) );
  NAND U16087 ( .A(n16036), .B(n16037), .Z(n16035) );
  NANDN U16088 ( .A(n16038), .B(n16039), .Z(n16036) );
  NANDN U16089 ( .A(n16039), .B(n16038), .Z(n16034) );
  NAND U16090 ( .A(n16040), .B(n16041), .Z(n276) );
  NANDN U16091 ( .A(n16042), .B(n16043), .Z(n16041) );
  OR U16092 ( .A(n16044), .B(n16045), .Z(n16043) );
  NAND U16093 ( .A(n16045), .B(n16044), .Z(n16040) );
  XOR U16094 ( .A(n278), .B(n277), .Z(\A1[257] ) );
  XOR U16095 ( .A(n16045), .B(n16046), .Z(n277) );
  XNOR U16096 ( .A(n16044), .B(n16042), .Z(n16046) );
  AND U16097 ( .A(n16047), .B(n16048), .Z(n16042) );
  NANDN U16098 ( .A(n16049), .B(n16050), .Z(n16048) );
  OR U16099 ( .A(n16051), .B(n16052), .Z(n16050) );
  NAND U16100 ( .A(n16052), .B(n16051), .Z(n16047) );
  ANDN U16101 ( .B(B[228]), .A(n54), .Z(n16044) );
  XNOR U16102 ( .A(n15864), .B(n16053), .Z(n16045) );
  XNOR U16103 ( .A(n15863), .B(n15861), .Z(n16053) );
  AND U16104 ( .A(n16054), .B(n16055), .Z(n15861) );
  NANDN U16105 ( .A(n16056), .B(n16057), .Z(n16055) );
  NANDN U16106 ( .A(n16058), .B(n16059), .Z(n16057) );
  NANDN U16107 ( .A(n16059), .B(n16058), .Z(n16054) );
  ANDN U16108 ( .B(B[229]), .A(n55), .Z(n15863) );
  XNOR U16109 ( .A(n15871), .B(n16060), .Z(n15864) );
  XNOR U16110 ( .A(n15870), .B(n15868), .Z(n16060) );
  AND U16111 ( .A(n16061), .B(n16062), .Z(n15868) );
  NANDN U16112 ( .A(n16063), .B(n16064), .Z(n16062) );
  OR U16113 ( .A(n16065), .B(n16066), .Z(n16064) );
  NAND U16114 ( .A(n16066), .B(n16065), .Z(n16061) );
  ANDN U16115 ( .B(B[230]), .A(n56), .Z(n15870) );
  XNOR U16116 ( .A(n15878), .B(n16067), .Z(n15871) );
  XNOR U16117 ( .A(n15877), .B(n15875), .Z(n16067) );
  AND U16118 ( .A(n16068), .B(n16069), .Z(n15875) );
  NANDN U16119 ( .A(n16070), .B(n16071), .Z(n16069) );
  NANDN U16120 ( .A(n16072), .B(n16073), .Z(n16071) );
  NANDN U16121 ( .A(n16073), .B(n16072), .Z(n16068) );
  ANDN U16122 ( .B(B[231]), .A(n57), .Z(n15877) );
  XNOR U16123 ( .A(n15885), .B(n16074), .Z(n15878) );
  XNOR U16124 ( .A(n15884), .B(n15882), .Z(n16074) );
  AND U16125 ( .A(n16075), .B(n16076), .Z(n15882) );
  NANDN U16126 ( .A(n16077), .B(n16078), .Z(n16076) );
  OR U16127 ( .A(n16079), .B(n16080), .Z(n16078) );
  NAND U16128 ( .A(n16080), .B(n16079), .Z(n16075) );
  ANDN U16129 ( .B(B[232]), .A(n58), .Z(n15884) );
  XNOR U16130 ( .A(n15892), .B(n16081), .Z(n15885) );
  XNOR U16131 ( .A(n15891), .B(n15889), .Z(n16081) );
  AND U16132 ( .A(n16082), .B(n16083), .Z(n15889) );
  NANDN U16133 ( .A(n16084), .B(n16085), .Z(n16083) );
  NANDN U16134 ( .A(n16086), .B(n16087), .Z(n16085) );
  NANDN U16135 ( .A(n16087), .B(n16086), .Z(n16082) );
  ANDN U16136 ( .B(B[233]), .A(n59), .Z(n15891) );
  XNOR U16137 ( .A(n15899), .B(n16088), .Z(n15892) );
  XNOR U16138 ( .A(n15898), .B(n15896), .Z(n16088) );
  AND U16139 ( .A(n16089), .B(n16090), .Z(n15896) );
  NANDN U16140 ( .A(n16091), .B(n16092), .Z(n16090) );
  OR U16141 ( .A(n16093), .B(n16094), .Z(n16092) );
  NAND U16142 ( .A(n16094), .B(n16093), .Z(n16089) );
  ANDN U16143 ( .B(B[234]), .A(n60), .Z(n15898) );
  XNOR U16144 ( .A(n15906), .B(n16095), .Z(n15899) );
  XNOR U16145 ( .A(n15905), .B(n15903), .Z(n16095) );
  AND U16146 ( .A(n16096), .B(n16097), .Z(n15903) );
  NANDN U16147 ( .A(n16098), .B(n16099), .Z(n16097) );
  NANDN U16148 ( .A(n16100), .B(n16101), .Z(n16099) );
  NANDN U16149 ( .A(n16101), .B(n16100), .Z(n16096) );
  ANDN U16150 ( .B(B[235]), .A(n61), .Z(n15905) );
  XNOR U16151 ( .A(n15913), .B(n16102), .Z(n15906) );
  XNOR U16152 ( .A(n15912), .B(n15910), .Z(n16102) );
  AND U16153 ( .A(n16103), .B(n16104), .Z(n15910) );
  NANDN U16154 ( .A(n16105), .B(n16106), .Z(n16104) );
  OR U16155 ( .A(n16107), .B(n16108), .Z(n16106) );
  NAND U16156 ( .A(n16108), .B(n16107), .Z(n16103) );
  ANDN U16157 ( .B(B[236]), .A(n62), .Z(n15912) );
  XNOR U16158 ( .A(n15920), .B(n16109), .Z(n15913) );
  XNOR U16159 ( .A(n15919), .B(n15917), .Z(n16109) );
  AND U16160 ( .A(n16110), .B(n16111), .Z(n15917) );
  NANDN U16161 ( .A(n16112), .B(n16113), .Z(n16111) );
  NANDN U16162 ( .A(n16114), .B(n16115), .Z(n16113) );
  NANDN U16163 ( .A(n16115), .B(n16114), .Z(n16110) );
  ANDN U16164 ( .B(B[237]), .A(n63), .Z(n15919) );
  XNOR U16165 ( .A(n15927), .B(n16116), .Z(n15920) );
  XNOR U16166 ( .A(n15926), .B(n15924), .Z(n16116) );
  AND U16167 ( .A(n16117), .B(n16118), .Z(n15924) );
  NANDN U16168 ( .A(n16119), .B(n16120), .Z(n16118) );
  OR U16169 ( .A(n16121), .B(n16122), .Z(n16120) );
  NAND U16170 ( .A(n16122), .B(n16121), .Z(n16117) );
  ANDN U16171 ( .B(B[238]), .A(n64), .Z(n15926) );
  XNOR U16172 ( .A(n15934), .B(n16123), .Z(n15927) );
  XNOR U16173 ( .A(n15933), .B(n15931), .Z(n16123) );
  AND U16174 ( .A(n16124), .B(n16125), .Z(n15931) );
  NANDN U16175 ( .A(n16126), .B(n16127), .Z(n16125) );
  NANDN U16176 ( .A(n16128), .B(n16129), .Z(n16127) );
  NANDN U16177 ( .A(n16129), .B(n16128), .Z(n16124) );
  ANDN U16178 ( .B(B[239]), .A(n65), .Z(n15933) );
  XNOR U16179 ( .A(n15941), .B(n16130), .Z(n15934) );
  XNOR U16180 ( .A(n15940), .B(n15938), .Z(n16130) );
  AND U16181 ( .A(n16131), .B(n16132), .Z(n15938) );
  NANDN U16182 ( .A(n16133), .B(n16134), .Z(n16132) );
  OR U16183 ( .A(n16135), .B(n16136), .Z(n16134) );
  NAND U16184 ( .A(n16136), .B(n16135), .Z(n16131) );
  ANDN U16185 ( .B(B[240]), .A(n66), .Z(n15940) );
  XNOR U16186 ( .A(n15948), .B(n16137), .Z(n15941) );
  XNOR U16187 ( .A(n15947), .B(n15945), .Z(n16137) );
  AND U16188 ( .A(n16138), .B(n16139), .Z(n15945) );
  NANDN U16189 ( .A(n16140), .B(n16141), .Z(n16139) );
  NANDN U16190 ( .A(n16142), .B(n16143), .Z(n16141) );
  NANDN U16191 ( .A(n16143), .B(n16142), .Z(n16138) );
  ANDN U16192 ( .B(B[241]), .A(n67), .Z(n15947) );
  XNOR U16193 ( .A(n15955), .B(n16144), .Z(n15948) );
  XNOR U16194 ( .A(n15954), .B(n15952), .Z(n16144) );
  AND U16195 ( .A(n16145), .B(n16146), .Z(n15952) );
  NANDN U16196 ( .A(n16147), .B(n16148), .Z(n16146) );
  OR U16197 ( .A(n16149), .B(n16150), .Z(n16148) );
  NAND U16198 ( .A(n16150), .B(n16149), .Z(n16145) );
  ANDN U16199 ( .B(B[242]), .A(n68), .Z(n15954) );
  XNOR U16200 ( .A(n15962), .B(n16151), .Z(n15955) );
  XNOR U16201 ( .A(n15961), .B(n15959), .Z(n16151) );
  AND U16202 ( .A(n16152), .B(n16153), .Z(n15959) );
  NANDN U16203 ( .A(n16154), .B(n16155), .Z(n16153) );
  NANDN U16204 ( .A(n16156), .B(n16157), .Z(n16155) );
  NANDN U16205 ( .A(n16157), .B(n16156), .Z(n16152) );
  ANDN U16206 ( .B(B[243]), .A(n69), .Z(n15961) );
  XNOR U16207 ( .A(n15969), .B(n16158), .Z(n15962) );
  XNOR U16208 ( .A(n15968), .B(n15966), .Z(n16158) );
  AND U16209 ( .A(n16159), .B(n16160), .Z(n15966) );
  NANDN U16210 ( .A(n16161), .B(n16162), .Z(n16160) );
  OR U16211 ( .A(n16163), .B(n16164), .Z(n16162) );
  NAND U16212 ( .A(n16164), .B(n16163), .Z(n16159) );
  ANDN U16213 ( .B(B[244]), .A(n70), .Z(n15968) );
  XNOR U16214 ( .A(n15976), .B(n16165), .Z(n15969) );
  XNOR U16215 ( .A(n15975), .B(n15973), .Z(n16165) );
  AND U16216 ( .A(n16166), .B(n16167), .Z(n15973) );
  NANDN U16217 ( .A(n16168), .B(n16169), .Z(n16167) );
  NANDN U16218 ( .A(n16170), .B(n16171), .Z(n16169) );
  NANDN U16219 ( .A(n16171), .B(n16170), .Z(n16166) );
  ANDN U16220 ( .B(B[245]), .A(n71), .Z(n15975) );
  XNOR U16221 ( .A(n15983), .B(n16172), .Z(n15976) );
  XNOR U16222 ( .A(n15982), .B(n15980), .Z(n16172) );
  AND U16223 ( .A(n16173), .B(n16174), .Z(n15980) );
  NANDN U16224 ( .A(n16175), .B(n16176), .Z(n16174) );
  OR U16225 ( .A(n16177), .B(n16178), .Z(n16176) );
  NAND U16226 ( .A(n16178), .B(n16177), .Z(n16173) );
  ANDN U16227 ( .B(B[246]), .A(n72), .Z(n15982) );
  XNOR U16228 ( .A(n15990), .B(n16179), .Z(n15983) );
  XNOR U16229 ( .A(n15989), .B(n15987), .Z(n16179) );
  AND U16230 ( .A(n16180), .B(n16181), .Z(n15987) );
  NANDN U16231 ( .A(n16182), .B(n16183), .Z(n16181) );
  NANDN U16232 ( .A(n16184), .B(n16185), .Z(n16183) );
  NANDN U16233 ( .A(n16185), .B(n16184), .Z(n16180) );
  ANDN U16234 ( .B(B[247]), .A(n73), .Z(n15989) );
  XNOR U16235 ( .A(n15997), .B(n16186), .Z(n15990) );
  XNOR U16236 ( .A(n15996), .B(n15994), .Z(n16186) );
  AND U16237 ( .A(n16187), .B(n16188), .Z(n15994) );
  NANDN U16238 ( .A(n16189), .B(n16190), .Z(n16188) );
  OR U16239 ( .A(n16191), .B(n16192), .Z(n16190) );
  NAND U16240 ( .A(n16192), .B(n16191), .Z(n16187) );
  ANDN U16241 ( .B(B[248]), .A(n74), .Z(n15996) );
  XNOR U16242 ( .A(n16004), .B(n16193), .Z(n15997) );
  XNOR U16243 ( .A(n16003), .B(n16001), .Z(n16193) );
  AND U16244 ( .A(n16194), .B(n16195), .Z(n16001) );
  NANDN U16245 ( .A(n16196), .B(n16197), .Z(n16195) );
  NANDN U16246 ( .A(n16198), .B(n16199), .Z(n16197) );
  NANDN U16247 ( .A(n16199), .B(n16198), .Z(n16194) );
  ANDN U16248 ( .B(B[249]), .A(n75), .Z(n16003) );
  XNOR U16249 ( .A(n16011), .B(n16200), .Z(n16004) );
  XNOR U16250 ( .A(n16010), .B(n16008), .Z(n16200) );
  AND U16251 ( .A(n16201), .B(n16202), .Z(n16008) );
  NANDN U16252 ( .A(n16203), .B(n16204), .Z(n16202) );
  OR U16253 ( .A(n16205), .B(n16206), .Z(n16204) );
  NAND U16254 ( .A(n16206), .B(n16205), .Z(n16201) );
  ANDN U16255 ( .B(B[250]), .A(n76), .Z(n16010) );
  XNOR U16256 ( .A(n16018), .B(n16207), .Z(n16011) );
  XNOR U16257 ( .A(n16017), .B(n16015), .Z(n16207) );
  AND U16258 ( .A(n16208), .B(n16209), .Z(n16015) );
  NANDN U16259 ( .A(n16210), .B(n16211), .Z(n16209) );
  NANDN U16260 ( .A(n16212), .B(n16213), .Z(n16211) );
  NANDN U16261 ( .A(n16213), .B(n16212), .Z(n16208) );
  ANDN U16262 ( .B(B[251]), .A(n77), .Z(n16017) );
  XNOR U16263 ( .A(n16025), .B(n16214), .Z(n16018) );
  XNOR U16264 ( .A(n16024), .B(n16022), .Z(n16214) );
  AND U16265 ( .A(n16215), .B(n16216), .Z(n16022) );
  NANDN U16266 ( .A(n16217), .B(n16218), .Z(n16216) );
  OR U16267 ( .A(n16219), .B(n16220), .Z(n16218) );
  NAND U16268 ( .A(n16220), .B(n16219), .Z(n16215) );
  ANDN U16269 ( .B(B[252]), .A(n78), .Z(n16024) );
  XNOR U16270 ( .A(n16032), .B(n16221), .Z(n16025) );
  XNOR U16271 ( .A(n16031), .B(n16029), .Z(n16221) );
  AND U16272 ( .A(n16222), .B(n16223), .Z(n16029) );
  NANDN U16273 ( .A(n16224), .B(n16225), .Z(n16223) );
  NANDN U16274 ( .A(n16226), .B(n16227), .Z(n16225) );
  NANDN U16275 ( .A(n16227), .B(n16226), .Z(n16222) );
  ANDN U16276 ( .B(B[253]), .A(n79), .Z(n16031) );
  XOR U16277 ( .A(n16037), .B(n16228), .Z(n16032) );
  XOR U16278 ( .A(n16038), .B(n16039), .Z(n16228) );
  NAND U16279 ( .A(A[4]), .B(B[255]), .Z(n16039) );
  AND U16280 ( .A(B[254]), .B(A[5]), .Z(n16038) );
  NAND U16281 ( .A(n16229), .B(n16230), .Z(n16037) );
  NAND U16282 ( .A(n16231), .B(n16232), .Z(n16230) );
  NANDN U16283 ( .A(n16233), .B(n16234), .Z(n16231) );
  NANDN U16284 ( .A(n16234), .B(n16233), .Z(n16229) );
  NAND U16285 ( .A(n16235), .B(n16236), .Z(n278) );
  NANDN U16286 ( .A(n16237), .B(n16238), .Z(n16236) );
  NAND U16287 ( .A(n16240), .B(n16239), .Z(n16235) );
  XOR U16288 ( .A(n280), .B(n279), .Z(\A1[256] ) );
  XOR U16289 ( .A(n16240), .B(n16241), .Z(n279) );
  XNOR U16290 ( .A(n16239), .B(n16237), .Z(n16241) );
  AND U16291 ( .A(n16242), .B(n16243), .Z(n16237) );
  NANDN U16292 ( .A(n16244), .B(n16245), .Z(n16243) );
  NANDN U16293 ( .A(n16246), .B(n16247), .Z(n16245) );
  NANDN U16294 ( .A(n16247), .B(n16246), .Z(n16242) );
  ANDN U16295 ( .B(B[227]), .A(n54), .Z(n16239) );
  XOR U16296 ( .A(n16052), .B(n16248), .Z(n16240) );
  XNOR U16297 ( .A(n16051), .B(n16049), .Z(n16248) );
  AND U16298 ( .A(n16249), .B(n16250), .Z(n16049) );
  NANDN U16299 ( .A(n16251), .B(n16252), .Z(n16250) );
  OR U16300 ( .A(n16253), .B(n16254), .Z(n16252) );
  NAND U16301 ( .A(n16254), .B(n16253), .Z(n16249) );
  ANDN U16302 ( .B(B[228]), .A(n55), .Z(n16051) );
  XNOR U16303 ( .A(n16059), .B(n16255), .Z(n16052) );
  XNOR U16304 ( .A(n16058), .B(n16056), .Z(n16255) );
  AND U16305 ( .A(n16256), .B(n16257), .Z(n16056) );
  NANDN U16306 ( .A(n16258), .B(n16259), .Z(n16257) );
  NANDN U16307 ( .A(n16260), .B(n16261), .Z(n16259) );
  NANDN U16308 ( .A(n16261), .B(n16260), .Z(n16256) );
  ANDN U16309 ( .B(B[229]), .A(n56), .Z(n16058) );
  XNOR U16310 ( .A(n16066), .B(n16262), .Z(n16059) );
  XNOR U16311 ( .A(n16065), .B(n16063), .Z(n16262) );
  AND U16312 ( .A(n16263), .B(n16264), .Z(n16063) );
  NANDN U16313 ( .A(n16265), .B(n16266), .Z(n16264) );
  OR U16314 ( .A(n16267), .B(n16268), .Z(n16266) );
  NAND U16315 ( .A(n16268), .B(n16267), .Z(n16263) );
  ANDN U16316 ( .B(B[230]), .A(n57), .Z(n16065) );
  XNOR U16317 ( .A(n16073), .B(n16269), .Z(n16066) );
  XNOR U16318 ( .A(n16072), .B(n16070), .Z(n16269) );
  AND U16319 ( .A(n16270), .B(n16271), .Z(n16070) );
  NANDN U16320 ( .A(n16272), .B(n16273), .Z(n16271) );
  NANDN U16321 ( .A(n16274), .B(n16275), .Z(n16273) );
  NANDN U16322 ( .A(n16275), .B(n16274), .Z(n16270) );
  ANDN U16323 ( .B(B[231]), .A(n58), .Z(n16072) );
  XNOR U16324 ( .A(n16080), .B(n16276), .Z(n16073) );
  XNOR U16325 ( .A(n16079), .B(n16077), .Z(n16276) );
  AND U16326 ( .A(n16277), .B(n16278), .Z(n16077) );
  NANDN U16327 ( .A(n16279), .B(n16280), .Z(n16278) );
  OR U16328 ( .A(n16281), .B(n16282), .Z(n16280) );
  NAND U16329 ( .A(n16282), .B(n16281), .Z(n16277) );
  ANDN U16330 ( .B(B[232]), .A(n59), .Z(n16079) );
  XNOR U16331 ( .A(n16087), .B(n16283), .Z(n16080) );
  XNOR U16332 ( .A(n16086), .B(n16084), .Z(n16283) );
  AND U16333 ( .A(n16284), .B(n16285), .Z(n16084) );
  NANDN U16334 ( .A(n16286), .B(n16287), .Z(n16285) );
  NANDN U16335 ( .A(n16288), .B(n16289), .Z(n16287) );
  NANDN U16336 ( .A(n16289), .B(n16288), .Z(n16284) );
  ANDN U16337 ( .B(B[233]), .A(n60), .Z(n16086) );
  XNOR U16338 ( .A(n16094), .B(n16290), .Z(n16087) );
  XNOR U16339 ( .A(n16093), .B(n16091), .Z(n16290) );
  AND U16340 ( .A(n16291), .B(n16292), .Z(n16091) );
  NANDN U16341 ( .A(n16293), .B(n16294), .Z(n16292) );
  OR U16342 ( .A(n16295), .B(n16296), .Z(n16294) );
  NAND U16343 ( .A(n16296), .B(n16295), .Z(n16291) );
  ANDN U16344 ( .B(B[234]), .A(n61), .Z(n16093) );
  XNOR U16345 ( .A(n16101), .B(n16297), .Z(n16094) );
  XNOR U16346 ( .A(n16100), .B(n16098), .Z(n16297) );
  AND U16347 ( .A(n16298), .B(n16299), .Z(n16098) );
  NANDN U16348 ( .A(n16300), .B(n16301), .Z(n16299) );
  NANDN U16349 ( .A(n16302), .B(n16303), .Z(n16301) );
  NANDN U16350 ( .A(n16303), .B(n16302), .Z(n16298) );
  ANDN U16351 ( .B(B[235]), .A(n62), .Z(n16100) );
  XNOR U16352 ( .A(n16108), .B(n16304), .Z(n16101) );
  XNOR U16353 ( .A(n16107), .B(n16105), .Z(n16304) );
  AND U16354 ( .A(n16305), .B(n16306), .Z(n16105) );
  NANDN U16355 ( .A(n16307), .B(n16308), .Z(n16306) );
  OR U16356 ( .A(n16309), .B(n16310), .Z(n16308) );
  NAND U16357 ( .A(n16310), .B(n16309), .Z(n16305) );
  ANDN U16358 ( .B(B[236]), .A(n63), .Z(n16107) );
  XNOR U16359 ( .A(n16115), .B(n16311), .Z(n16108) );
  XNOR U16360 ( .A(n16114), .B(n16112), .Z(n16311) );
  AND U16361 ( .A(n16312), .B(n16313), .Z(n16112) );
  NANDN U16362 ( .A(n16314), .B(n16315), .Z(n16313) );
  NANDN U16363 ( .A(n16316), .B(n16317), .Z(n16315) );
  NANDN U16364 ( .A(n16317), .B(n16316), .Z(n16312) );
  ANDN U16365 ( .B(B[237]), .A(n64), .Z(n16114) );
  XNOR U16366 ( .A(n16122), .B(n16318), .Z(n16115) );
  XNOR U16367 ( .A(n16121), .B(n16119), .Z(n16318) );
  AND U16368 ( .A(n16319), .B(n16320), .Z(n16119) );
  NANDN U16369 ( .A(n16321), .B(n16322), .Z(n16320) );
  OR U16370 ( .A(n16323), .B(n16324), .Z(n16322) );
  NAND U16371 ( .A(n16324), .B(n16323), .Z(n16319) );
  ANDN U16372 ( .B(B[238]), .A(n65), .Z(n16121) );
  XNOR U16373 ( .A(n16129), .B(n16325), .Z(n16122) );
  XNOR U16374 ( .A(n16128), .B(n16126), .Z(n16325) );
  AND U16375 ( .A(n16326), .B(n16327), .Z(n16126) );
  NANDN U16376 ( .A(n16328), .B(n16329), .Z(n16327) );
  NANDN U16377 ( .A(n16330), .B(n16331), .Z(n16329) );
  NANDN U16378 ( .A(n16331), .B(n16330), .Z(n16326) );
  ANDN U16379 ( .B(B[239]), .A(n66), .Z(n16128) );
  XNOR U16380 ( .A(n16136), .B(n16332), .Z(n16129) );
  XNOR U16381 ( .A(n16135), .B(n16133), .Z(n16332) );
  AND U16382 ( .A(n16333), .B(n16334), .Z(n16133) );
  NANDN U16383 ( .A(n16335), .B(n16336), .Z(n16334) );
  OR U16384 ( .A(n16337), .B(n16338), .Z(n16336) );
  NAND U16385 ( .A(n16338), .B(n16337), .Z(n16333) );
  ANDN U16386 ( .B(B[240]), .A(n67), .Z(n16135) );
  XNOR U16387 ( .A(n16143), .B(n16339), .Z(n16136) );
  XNOR U16388 ( .A(n16142), .B(n16140), .Z(n16339) );
  AND U16389 ( .A(n16340), .B(n16341), .Z(n16140) );
  NANDN U16390 ( .A(n16342), .B(n16343), .Z(n16341) );
  NANDN U16391 ( .A(n16344), .B(n16345), .Z(n16343) );
  NANDN U16392 ( .A(n16345), .B(n16344), .Z(n16340) );
  ANDN U16393 ( .B(B[241]), .A(n68), .Z(n16142) );
  XNOR U16394 ( .A(n16150), .B(n16346), .Z(n16143) );
  XNOR U16395 ( .A(n16149), .B(n16147), .Z(n16346) );
  AND U16396 ( .A(n16347), .B(n16348), .Z(n16147) );
  NANDN U16397 ( .A(n16349), .B(n16350), .Z(n16348) );
  OR U16398 ( .A(n16351), .B(n16352), .Z(n16350) );
  NAND U16399 ( .A(n16352), .B(n16351), .Z(n16347) );
  ANDN U16400 ( .B(B[242]), .A(n69), .Z(n16149) );
  XNOR U16401 ( .A(n16157), .B(n16353), .Z(n16150) );
  XNOR U16402 ( .A(n16156), .B(n16154), .Z(n16353) );
  AND U16403 ( .A(n16354), .B(n16355), .Z(n16154) );
  NANDN U16404 ( .A(n16356), .B(n16357), .Z(n16355) );
  NANDN U16405 ( .A(n16358), .B(n16359), .Z(n16357) );
  NANDN U16406 ( .A(n16359), .B(n16358), .Z(n16354) );
  ANDN U16407 ( .B(B[243]), .A(n70), .Z(n16156) );
  XNOR U16408 ( .A(n16164), .B(n16360), .Z(n16157) );
  XNOR U16409 ( .A(n16163), .B(n16161), .Z(n16360) );
  AND U16410 ( .A(n16361), .B(n16362), .Z(n16161) );
  NANDN U16411 ( .A(n16363), .B(n16364), .Z(n16362) );
  OR U16412 ( .A(n16365), .B(n16366), .Z(n16364) );
  NAND U16413 ( .A(n16366), .B(n16365), .Z(n16361) );
  ANDN U16414 ( .B(B[244]), .A(n71), .Z(n16163) );
  XNOR U16415 ( .A(n16171), .B(n16367), .Z(n16164) );
  XNOR U16416 ( .A(n16170), .B(n16168), .Z(n16367) );
  AND U16417 ( .A(n16368), .B(n16369), .Z(n16168) );
  NANDN U16418 ( .A(n16370), .B(n16371), .Z(n16369) );
  NANDN U16419 ( .A(n16372), .B(n16373), .Z(n16371) );
  NANDN U16420 ( .A(n16373), .B(n16372), .Z(n16368) );
  ANDN U16421 ( .B(B[245]), .A(n72), .Z(n16170) );
  XNOR U16422 ( .A(n16178), .B(n16374), .Z(n16171) );
  XNOR U16423 ( .A(n16177), .B(n16175), .Z(n16374) );
  AND U16424 ( .A(n16375), .B(n16376), .Z(n16175) );
  NANDN U16425 ( .A(n16377), .B(n16378), .Z(n16376) );
  OR U16426 ( .A(n16379), .B(n16380), .Z(n16378) );
  NAND U16427 ( .A(n16380), .B(n16379), .Z(n16375) );
  ANDN U16428 ( .B(B[246]), .A(n73), .Z(n16177) );
  XNOR U16429 ( .A(n16185), .B(n16381), .Z(n16178) );
  XNOR U16430 ( .A(n16184), .B(n16182), .Z(n16381) );
  AND U16431 ( .A(n16382), .B(n16383), .Z(n16182) );
  NANDN U16432 ( .A(n16384), .B(n16385), .Z(n16383) );
  NANDN U16433 ( .A(n16386), .B(n16387), .Z(n16385) );
  NANDN U16434 ( .A(n16387), .B(n16386), .Z(n16382) );
  ANDN U16435 ( .B(B[247]), .A(n74), .Z(n16184) );
  XNOR U16436 ( .A(n16192), .B(n16388), .Z(n16185) );
  XNOR U16437 ( .A(n16191), .B(n16189), .Z(n16388) );
  AND U16438 ( .A(n16389), .B(n16390), .Z(n16189) );
  NANDN U16439 ( .A(n16391), .B(n16392), .Z(n16390) );
  OR U16440 ( .A(n16393), .B(n16394), .Z(n16392) );
  NAND U16441 ( .A(n16394), .B(n16393), .Z(n16389) );
  ANDN U16442 ( .B(B[248]), .A(n75), .Z(n16191) );
  XNOR U16443 ( .A(n16199), .B(n16395), .Z(n16192) );
  XNOR U16444 ( .A(n16198), .B(n16196), .Z(n16395) );
  AND U16445 ( .A(n16396), .B(n16397), .Z(n16196) );
  NANDN U16446 ( .A(n16398), .B(n16399), .Z(n16397) );
  NANDN U16447 ( .A(n16400), .B(n16401), .Z(n16399) );
  NANDN U16448 ( .A(n16401), .B(n16400), .Z(n16396) );
  ANDN U16449 ( .B(B[249]), .A(n76), .Z(n16198) );
  XNOR U16450 ( .A(n16206), .B(n16402), .Z(n16199) );
  XNOR U16451 ( .A(n16205), .B(n16203), .Z(n16402) );
  AND U16452 ( .A(n16403), .B(n16404), .Z(n16203) );
  NANDN U16453 ( .A(n16405), .B(n16406), .Z(n16404) );
  OR U16454 ( .A(n16407), .B(n16408), .Z(n16406) );
  NAND U16455 ( .A(n16408), .B(n16407), .Z(n16403) );
  ANDN U16456 ( .B(B[250]), .A(n77), .Z(n16205) );
  XNOR U16457 ( .A(n16213), .B(n16409), .Z(n16206) );
  XNOR U16458 ( .A(n16212), .B(n16210), .Z(n16409) );
  AND U16459 ( .A(n16410), .B(n16411), .Z(n16210) );
  NANDN U16460 ( .A(n16412), .B(n16413), .Z(n16411) );
  NANDN U16461 ( .A(n16414), .B(n16415), .Z(n16413) );
  NANDN U16462 ( .A(n16415), .B(n16414), .Z(n16410) );
  ANDN U16463 ( .B(B[251]), .A(n78), .Z(n16212) );
  XNOR U16464 ( .A(n16220), .B(n16416), .Z(n16213) );
  XNOR U16465 ( .A(n16219), .B(n16217), .Z(n16416) );
  AND U16466 ( .A(n16417), .B(n16418), .Z(n16217) );
  NANDN U16467 ( .A(n16419), .B(n16420), .Z(n16418) );
  OR U16468 ( .A(n16421), .B(n16422), .Z(n16420) );
  NAND U16469 ( .A(n16422), .B(n16421), .Z(n16417) );
  ANDN U16470 ( .B(B[252]), .A(n79), .Z(n16219) );
  XNOR U16471 ( .A(n16227), .B(n16423), .Z(n16220) );
  XNOR U16472 ( .A(n16226), .B(n16224), .Z(n16423) );
  AND U16473 ( .A(n16424), .B(n16425), .Z(n16224) );
  NANDN U16474 ( .A(n16426), .B(n16427), .Z(n16425) );
  NANDN U16475 ( .A(n16428), .B(n16429), .Z(n16427) );
  NANDN U16476 ( .A(n16429), .B(n16428), .Z(n16424) );
  ANDN U16477 ( .B(B[253]), .A(n80), .Z(n16226) );
  XOR U16478 ( .A(n16232), .B(n16430), .Z(n16227) );
  XOR U16479 ( .A(n16233), .B(n16234), .Z(n16430) );
  NAND U16480 ( .A(A[3]), .B(B[255]), .Z(n16234) );
  AND U16481 ( .A(B[254]), .B(A[4]), .Z(n16233) );
  NAND U16482 ( .A(n16431), .B(n16432), .Z(n16232) );
  NANDN U16483 ( .A(n16434), .B(n16435), .Z(n16433) );
  NANDN U16484 ( .A(n16435), .B(n16434), .Z(n16431) );
  NAND U16485 ( .A(n16437), .B(n16438), .Z(n280) );
  NANDN U16486 ( .A(n16439), .B(n16440), .Z(n16438) );
  OR U16487 ( .A(n16441), .B(n16442), .Z(n16440) );
  NAND U16488 ( .A(n16442), .B(n16441), .Z(n16437) );
  XOR U16489 ( .A(n282), .B(n281), .Z(\A1[255] ) );
  XOR U16490 ( .A(n16442), .B(n16443), .Z(n281) );
  XNOR U16491 ( .A(n16441), .B(n16439), .Z(n16443) );
  AND U16492 ( .A(n16444), .B(n16445), .Z(n16439) );
  NANDN U16493 ( .A(n16446), .B(n16447), .Z(n16445) );
  NANDN U16494 ( .A(n16448), .B(n16449), .Z(n16447) );
  NANDN U16495 ( .A(n16449), .B(n16448), .Z(n16444) );
  ANDN U16496 ( .B(B[226]), .A(n54), .Z(n16441) );
  XNOR U16497 ( .A(n16247), .B(n16450), .Z(n16442) );
  XNOR U16498 ( .A(n16246), .B(n16244), .Z(n16450) );
  AND U16499 ( .A(n16451), .B(n16452), .Z(n16244) );
  NANDN U16500 ( .A(n16453), .B(n16454), .Z(n16452) );
  OR U16501 ( .A(n16455), .B(n16456), .Z(n16454) );
  NAND U16502 ( .A(n16456), .B(n16455), .Z(n16451) );
  ANDN U16503 ( .B(B[227]), .A(n55), .Z(n16246) );
  XNOR U16504 ( .A(n16254), .B(n16457), .Z(n16247) );
  XNOR U16505 ( .A(n16253), .B(n16251), .Z(n16457) );
  AND U16506 ( .A(n16458), .B(n16459), .Z(n16251) );
  NANDN U16507 ( .A(n16460), .B(n16461), .Z(n16459) );
  NANDN U16508 ( .A(n16462), .B(n16463), .Z(n16461) );
  NANDN U16509 ( .A(n16463), .B(n16462), .Z(n16458) );
  ANDN U16510 ( .B(B[228]), .A(n56), .Z(n16253) );
  XNOR U16511 ( .A(n16261), .B(n16464), .Z(n16254) );
  XNOR U16512 ( .A(n16260), .B(n16258), .Z(n16464) );
  AND U16513 ( .A(n16465), .B(n16466), .Z(n16258) );
  NANDN U16514 ( .A(n16467), .B(n16468), .Z(n16466) );
  OR U16515 ( .A(n16469), .B(n16470), .Z(n16468) );
  NAND U16516 ( .A(n16470), .B(n16469), .Z(n16465) );
  ANDN U16517 ( .B(B[229]), .A(n57), .Z(n16260) );
  XNOR U16518 ( .A(n16268), .B(n16471), .Z(n16261) );
  XNOR U16519 ( .A(n16267), .B(n16265), .Z(n16471) );
  AND U16520 ( .A(n16472), .B(n16473), .Z(n16265) );
  NANDN U16521 ( .A(n16474), .B(n16475), .Z(n16473) );
  NANDN U16522 ( .A(n16476), .B(n16477), .Z(n16475) );
  NANDN U16523 ( .A(n16477), .B(n16476), .Z(n16472) );
  ANDN U16524 ( .B(B[230]), .A(n58), .Z(n16267) );
  XNOR U16525 ( .A(n16275), .B(n16478), .Z(n16268) );
  XNOR U16526 ( .A(n16274), .B(n16272), .Z(n16478) );
  AND U16527 ( .A(n16479), .B(n16480), .Z(n16272) );
  NANDN U16528 ( .A(n16481), .B(n16482), .Z(n16480) );
  OR U16529 ( .A(n16483), .B(n16484), .Z(n16482) );
  NAND U16530 ( .A(n16484), .B(n16483), .Z(n16479) );
  ANDN U16531 ( .B(B[231]), .A(n59), .Z(n16274) );
  XNOR U16532 ( .A(n16282), .B(n16485), .Z(n16275) );
  XNOR U16533 ( .A(n16281), .B(n16279), .Z(n16485) );
  AND U16534 ( .A(n16486), .B(n16487), .Z(n16279) );
  NANDN U16535 ( .A(n16488), .B(n16489), .Z(n16487) );
  NANDN U16536 ( .A(n16490), .B(n16491), .Z(n16489) );
  NANDN U16537 ( .A(n16491), .B(n16490), .Z(n16486) );
  ANDN U16538 ( .B(B[232]), .A(n60), .Z(n16281) );
  XNOR U16539 ( .A(n16289), .B(n16492), .Z(n16282) );
  XNOR U16540 ( .A(n16288), .B(n16286), .Z(n16492) );
  AND U16541 ( .A(n16493), .B(n16494), .Z(n16286) );
  NANDN U16542 ( .A(n16495), .B(n16496), .Z(n16494) );
  OR U16543 ( .A(n16497), .B(n16498), .Z(n16496) );
  NAND U16544 ( .A(n16498), .B(n16497), .Z(n16493) );
  ANDN U16545 ( .B(B[233]), .A(n61), .Z(n16288) );
  XNOR U16546 ( .A(n16296), .B(n16499), .Z(n16289) );
  XNOR U16547 ( .A(n16295), .B(n16293), .Z(n16499) );
  AND U16548 ( .A(n16500), .B(n16501), .Z(n16293) );
  NANDN U16549 ( .A(n16502), .B(n16503), .Z(n16501) );
  NANDN U16550 ( .A(n16504), .B(n16505), .Z(n16503) );
  NANDN U16551 ( .A(n16505), .B(n16504), .Z(n16500) );
  ANDN U16552 ( .B(B[234]), .A(n62), .Z(n16295) );
  XNOR U16553 ( .A(n16303), .B(n16506), .Z(n16296) );
  XNOR U16554 ( .A(n16302), .B(n16300), .Z(n16506) );
  AND U16555 ( .A(n16507), .B(n16508), .Z(n16300) );
  NANDN U16556 ( .A(n16509), .B(n16510), .Z(n16508) );
  OR U16557 ( .A(n16511), .B(n16512), .Z(n16510) );
  NAND U16558 ( .A(n16512), .B(n16511), .Z(n16507) );
  ANDN U16559 ( .B(B[235]), .A(n63), .Z(n16302) );
  XNOR U16560 ( .A(n16310), .B(n16513), .Z(n16303) );
  XNOR U16561 ( .A(n16309), .B(n16307), .Z(n16513) );
  AND U16562 ( .A(n16514), .B(n16515), .Z(n16307) );
  NANDN U16563 ( .A(n16516), .B(n16517), .Z(n16515) );
  NANDN U16564 ( .A(n16518), .B(n16519), .Z(n16517) );
  NANDN U16565 ( .A(n16519), .B(n16518), .Z(n16514) );
  ANDN U16566 ( .B(B[236]), .A(n64), .Z(n16309) );
  XNOR U16567 ( .A(n16317), .B(n16520), .Z(n16310) );
  XNOR U16568 ( .A(n16316), .B(n16314), .Z(n16520) );
  AND U16569 ( .A(n16521), .B(n16522), .Z(n16314) );
  NANDN U16570 ( .A(n16523), .B(n16524), .Z(n16522) );
  OR U16571 ( .A(n16525), .B(n16526), .Z(n16524) );
  NAND U16572 ( .A(n16526), .B(n16525), .Z(n16521) );
  ANDN U16573 ( .B(B[237]), .A(n65), .Z(n16316) );
  XNOR U16574 ( .A(n16324), .B(n16527), .Z(n16317) );
  XNOR U16575 ( .A(n16323), .B(n16321), .Z(n16527) );
  AND U16576 ( .A(n16528), .B(n16529), .Z(n16321) );
  NANDN U16577 ( .A(n16530), .B(n16531), .Z(n16529) );
  NANDN U16578 ( .A(n16532), .B(n16533), .Z(n16531) );
  NANDN U16579 ( .A(n16533), .B(n16532), .Z(n16528) );
  ANDN U16580 ( .B(B[238]), .A(n66), .Z(n16323) );
  XNOR U16581 ( .A(n16331), .B(n16534), .Z(n16324) );
  XNOR U16582 ( .A(n16330), .B(n16328), .Z(n16534) );
  AND U16583 ( .A(n16535), .B(n16536), .Z(n16328) );
  NANDN U16584 ( .A(n16537), .B(n16538), .Z(n16536) );
  OR U16585 ( .A(n16539), .B(n16540), .Z(n16538) );
  NAND U16586 ( .A(n16540), .B(n16539), .Z(n16535) );
  ANDN U16587 ( .B(B[239]), .A(n67), .Z(n16330) );
  XNOR U16588 ( .A(n16338), .B(n16541), .Z(n16331) );
  XNOR U16589 ( .A(n16337), .B(n16335), .Z(n16541) );
  AND U16590 ( .A(n16542), .B(n16543), .Z(n16335) );
  NANDN U16591 ( .A(n16544), .B(n16545), .Z(n16543) );
  NANDN U16592 ( .A(n16546), .B(n16547), .Z(n16545) );
  NANDN U16593 ( .A(n16547), .B(n16546), .Z(n16542) );
  ANDN U16594 ( .B(B[240]), .A(n68), .Z(n16337) );
  XNOR U16595 ( .A(n16345), .B(n16548), .Z(n16338) );
  XNOR U16596 ( .A(n16344), .B(n16342), .Z(n16548) );
  AND U16597 ( .A(n16549), .B(n16550), .Z(n16342) );
  NANDN U16598 ( .A(n16551), .B(n16552), .Z(n16550) );
  OR U16599 ( .A(n16553), .B(n16554), .Z(n16552) );
  NAND U16600 ( .A(n16554), .B(n16553), .Z(n16549) );
  ANDN U16601 ( .B(B[241]), .A(n69), .Z(n16344) );
  XNOR U16602 ( .A(n16352), .B(n16555), .Z(n16345) );
  XNOR U16603 ( .A(n16351), .B(n16349), .Z(n16555) );
  AND U16604 ( .A(n16556), .B(n16557), .Z(n16349) );
  NANDN U16605 ( .A(n16558), .B(n16559), .Z(n16557) );
  NANDN U16606 ( .A(n16560), .B(n16561), .Z(n16559) );
  NANDN U16607 ( .A(n16561), .B(n16560), .Z(n16556) );
  ANDN U16608 ( .B(B[242]), .A(n70), .Z(n16351) );
  XNOR U16609 ( .A(n16359), .B(n16562), .Z(n16352) );
  XNOR U16610 ( .A(n16358), .B(n16356), .Z(n16562) );
  AND U16611 ( .A(n16563), .B(n16564), .Z(n16356) );
  NANDN U16612 ( .A(n16565), .B(n16566), .Z(n16564) );
  OR U16613 ( .A(n16567), .B(n16568), .Z(n16566) );
  NAND U16614 ( .A(n16568), .B(n16567), .Z(n16563) );
  ANDN U16615 ( .B(B[243]), .A(n71), .Z(n16358) );
  XNOR U16616 ( .A(n16366), .B(n16569), .Z(n16359) );
  XNOR U16617 ( .A(n16365), .B(n16363), .Z(n16569) );
  AND U16618 ( .A(n16570), .B(n16571), .Z(n16363) );
  NANDN U16619 ( .A(n16572), .B(n16573), .Z(n16571) );
  NANDN U16620 ( .A(n16574), .B(n16575), .Z(n16573) );
  NANDN U16621 ( .A(n16575), .B(n16574), .Z(n16570) );
  ANDN U16622 ( .B(B[244]), .A(n72), .Z(n16365) );
  XNOR U16623 ( .A(n16373), .B(n16576), .Z(n16366) );
  XNOR U16624 ( .A(n16372), .B(n16370), .Z(n16576) );
  AND U16625 ( .A(n16577), .B(n16578), .Z(n16370) );
  NANDN U16626 ( .A(n16579), .B(n16580), .Z(n16578) );
  OR U16627 ( .A(n16581), .B(n16582), .Z(n16580) );
  NAND U16628 ( .A(n16582), .B(n16581), .Z(n16577) );
  ANDN U16629 ( .B(B[245]), .A(n73), .Z(n16372) );
  XNOR U16630 ( .A(n16380), .B(n16583), .Z(n16373) );
  XNOR U16631 ( .A(n16379), .B(n16377), .Z(n16583) );
  AND U16632 ( .A(n16584), .B(n16585), .Z(n16377) );
  NANDN U16633 ( .A(n16586), .B(n16587), .Z(n16585) );
  NANDN U16634 ( .A(n16588), .B(n16589), .Z(n16587) );
  NANDN U16635 ( .A(n16589), .B(n16588), .Z(n16584) );
  ANDN U16636 ( .B(B[246]), .A(n74), .Z(n16379) );
  XNOR U16637 ( .A(n16387), .B(n16590), .Z(n16380) );
  XNOR U16638 ( .A(n16386), .B(n16384), .Z(n16590) );
  AND U16639 ( .A(n16591), .B(n16592), .Z(n16384) );
  NANDN U16640 ( .A(n16593), .B(n16594), .Z(n16592) );
  OR U16641 ( .A(n16595), .B(n16596), .Z(n16594) );
  NAND U16642 ( .A(n16596), .B(n16595), .Z(n16591) );
  ANDN U16643 ( .B(B[247]), .A(n75), .Z(n16386) );
  XNOR U16644 ( .A(n16394), .B(n16597), .Z(n16387) );
  XNOR U16645 ( .A(n16393), .B(n16391), .Z(n16597) );
  AND U16646 ( .A(n16598), .B(n16599), .Z(n16391) );
  NANDN U16647 ( .A(n16600), .B(n16601), .Z(n16599) );
  NANDN U16648 ( .A(n16602), .B(n16603), .Z(n16601) );
  NANDN U16649 ( .A(n16603), .B(n16602), .Z(n16598) );
  ANDN U16650 ( .B(B[248]), .A(n76), .Z(n16393) );
  XNOR U16651 ( .A(n16401), .B(n16604), .Z(n16394) );
  XNOR U16652 ( .A(n16400), .B(n16398), .Z(n16604) );
  AND U16653 ( .A(n16605), .B(n16606), .Z(n16398) );
  NANDN U16654 ( .A(n16607), .B(n16608), .Z(n16606) );
  OR U16655 ( .A(n16609), .B(n16610), .Z(n16608) );
  NAND U16656 ( .A(n16610), .B(n16609), .Z(n16605) );
  ANDN U16657 ( .B(B[249]), .A(n77), .Z(n16400) );
  XNOR U16658 ( .A(n16408), .B(n16611), .Z(n16401) );
  XNOR U16659 ( .A(n16407), .B(n16405), .Z(n16611) );
  AND U16660 ( .A(n16612), .B(n16613), .Z(n16405) );
  NANDN U16661 ( .A(n16614), .B(n16615), .Z(n16613) );
  NANDN U16662 ( .A(n16616), .B(n16617), .Z(n16615) );
  NANDN U16663 ( .A(n16617), .B(n16616), .Z(n16612) );
  ANDN U16664 ( .B(B[250]), .A(n78), .Z(n16407) );
  XNOR U16665 ( .A(n16415), .B(n16618), .Z(n16408) );
  XNOR U16666 ( .A(n16414), .B(n16412), .Z(n16618) );
  AND U16667 ( .A(n16619), .B(n16620), .Z(n16412) );
  NANDN U16668 ( .A(n16621), .B(n16622), .Z(n16620) );
  OR U16669 ( .A(n16623), .B(n16624), .Z(n16622) );
  NAND U16670 ( .A(n16624), .B(n16623), .Z(n16619) );
  ANDN U16671 ( .B(B[251]), .A(n79), .Z(n16414) );
  XNOR U16672 ( .A(n16422), .B(n16625), .Z(n16415) );
  XNOR U16673 ( .A(n16421), .B(n16419), .Z(n16625) );
  AND U16674 ( .A(n16626), .B(n16627), .Z(n16419) );
  NANDN U16675 ( .A(n16628), .B(n16629), .Z(n16627) );
  NANDN U16676 ( .A(n16630), .B(n16631), .Z(n16629) );
  NANDN U16677 ( .A(n16631), .B(n16630), .Z(n16626) );
  ANDN U16678 ( .B(B[252]), .A(n80), .Z(n16421) );
  XNOR U16679 ( .A(n16429), .B(n16632), .Z(n16422) );
  XNOR U16680 ( .A(n16428), .B(n16426), .Z(n16632) );
  AND U16681 ( .A(n16633), .B(n16634), .Z(n16426) );
  NANDN U16682 ( .A(n16635), .B(n16636), .Z(n16634) );
  NANDN U16683 ( .A(n16637), .B(n16638), .Z(n16636) );
  NAND U16684 ( .A(n3), .B(n16637), .Z(n16633) );
  ANDN U16685 ( .B(B[253]), .A(n81), .Z(n16428) );
  XNOR U16686 ( .A(n16436), .B(n16639), .Z(n16429) );
  XOR U16687 ( .A(n16434), .B(n16435), .Z(n16639) );
  NAND U16688 ( .A(B[255]), .B(A[2]), .Z(n16435) );
  AND U16689 ( .A(B[254]), .B(A[3]), .Z(n16434) );
  AND U16690 ( .A(n16640), .B(n16641), .Z(n16436) );
  OR U16691 ( .A(n16642), .B(n16643), .Z(n16640) );
  NAND U16692 ( .A(n16644), .B(n16645), .Z(n282) );
  NANDN U16693 ( .A(n16646), .B(n16647), .Z(n16645) );
  OR U16694 ( .A(n16648), .B(n16649), .Z(n16647) );
  NAND U16695 ( .A(n16649), .B(n16648), .Z(n16644) );
  XOR U16696 ( .A(n284), .B(n283), .Z(\A1[254] ) );
  XOR U16697 ( .A(n16649), .B(n16650), .Z(n283) );
  XNOR U16698 ( .A(n16648), .B(n16646), .Z(n16650) );
  AND U16699 ( .A(n16651), .B(n16652), .Z(n16646) );
  NANDN U16700 ( .A(n16653), .B(n16654), .Z(n16652) );
  NANDN U16701 ( .A(n16655), .B(n16656), .Z(n16654) );
  NANDN U16702 ( .A(n16656), .B(n16655), .Z(n16651) );
  ANDN U16703 ( .B(B[225]), .A(n54), .Z(n16648) );
  XNOR U16704 ( .A(n16449), .B(n16657), .Z(n16649) );
  XNOR U16705 ( .A(n16448), .B(n16446), .Z(n16657) );
  AND U16706 ( .A(n16658), .B(n16659), .Z(n16446) );
  NANDN U16707 ( .A(n16660), .B(n16661), .Z(n16659) );
  OR U16708 ( .A(n16662), .B(n16663), .Z(n16661) );
  NAND U16709 ( .A(n16663), .B(n16662), .Z(n16658) );
  ANDN U16710 ( .B(B[226]), .A(n55), .Z(n16448) );
  XNOR U16711 ( .A(n16456), .B(n16664), .Z(n16449) );
  XNOR U16712 ( .A(n16455), .B(n16453), .Z(n16664) );
  AND U16713 ( .A(n16665), .B(n16666), .Z(n16453) );
  NANDN U16714 ( .A(n16667), .B(n16668), .Z(n16666) );
  NANDN U16715 ( .A(n16669), .B(n16670), .Z(n16668) );
  NANDN U16716 ( .A(n16670), .B(n16669), .Z(n16665) );
  ANDN U16717 ( .B(B[227]), .A(n56), .Z(n16455) );
  XNOR U16718 ( .A(n16463), .B(n16671), .Z(n16456) );
  XNOR U16719 ( .A(n16462), .B(n16460), .Z(n16671) );
  AND U16720 ( .A(n16672), .B(n16673), .Z(n16460) );
  NANDN U16721 ( .A(n16674), .B(n16675), .Z(n16673) );
  OR U16722 ( .A(n16676), .B(n16677), .Z(n16675) );
  NAND U16723 ( .A(n16677), .B(n16676), .Z(n16672) );
  ANDN U16724 ( .B(B[228]), .A(n57), .Z(n16462) );
  XNOR U16725 ( .A(n16470), .B(n16678), .Z(n16463) );
  XNOR U16726 ( .A(n16469), .B(n16467), .Z(n16678) );
  AND U16727 ( .A(n16679), .B(n16680), .Z(n16467) );
  NANDN U16728 ( .A(n16681), .B(n16682), .Z(n16680) );
  NANDN U16729 ( .A(n16683), .B(n16684), .Z(n16682) );
  NANDN U16730 ( .A(n16684), .B(n16683), .Z(n16679) );
  ANDN U16731 ( .B(B[229]), .A(n58), .Z(n16469) );
  XNOR U16732 ( .A(n16477), .B(n16685), .Z(n16470) );
  XNOR U16733 ( .A(n16476), .B(n16474), .Z(n16685) );
  AND U16734 ( .A(n16686), .B(n16687), .Z(n16474) );
  NANDN U16735 ( .A(n16688), .B(n16689), .Z(n16687) );
  OR U16736 ( .A(n16690), .B(n16691), .Z(n16689) );
  NAND U16737 ( .A(n16691), .B(n16690), .Z(n16686) );
  ANDN U16738 ( .B(B[230]), .A(n59), .Z(n16476) );
  XNOR U16739 ( .A(n16484), .B(n16692), .Z(n16477) );
  XNOR U16740 ( .A(n16483), .B(n16481), .Z(n16692) );
  AND U16741 ( .A(n16693), .B(n16694), .Z(n16481) );
  NANDN U16742 ( .A(n16695), .B(n16696), .Z(n16694) );
  NANDN U16743 ( .A(n16697), .B(n16698), .Z(n16696) );
  NANDN U16744 ( .A(n16698), .B(n16697), .Z(n16693) );
  ANDN U16745 ( .B(B[231]), .A(n60), .Z(n16483) );
  XNOR U16746 ( .A(n16491), .B(n16699), .Z(n16484) );
  XNOR U16747 ( .A(n16490), .B(n16488), .Z(n16699) );
  AND U16748 ( .A(n16700), .B(n16701), .Z(n16488) );
  NANDN U16749 ( .A(n16702), .B(n16703), .Z(n16701) );
  OR U16750 ( .A(n16704), .B(n16705), .Z(n16703) );
  NAND U16751 ( .A(n16705), .B(n16704), .Z(n16700) );
  ANDN U16752 ( .B(B[232]), .A(n61), .Z(n16490) );
  XNOR U16753 ( .A(n16498), .B(n16706), .Z(n16491) );
  XNOR U16754 ( .A(n16497), .B(n16495), .Z(n16706) );
  AND U16755 ( .A(n16707), .B(n16708), .Z(n16495) );
  NANDN U16756 ( .A(n16709), .B(n16710), .Z(n16708) );
  NANDN U16757 ( .A(n16711), .B(n16712), .Z(n16710) );
  NANDN U16758 ( .A(n16712), .B(n16711), .Z(n16707) );
  ANDN U16759 ( .B(B[233]), .A(n62), .Z(n16497) );
  XNOR U16760 ( .A(n16505), .B(n16713), .Z(n16498) );
  XNOR U16761 ( .A(n16504), .B(n16502), .Z(n16713) );
  AND U16762 ( .A(n16714), .B(n16715), .Z(n16502) );
  NANDN U16763 ( .A(n16716), .B(n16717), .Z(n16715) );
  OR U16764 ( .A(n16718), .B(n16719), .Z(n16717) );
  NAND U16765 ( .A(n16719), .B(n16718), .Z(n16714) );
  ANDN U16766 ( .B(B[234]), .A(n63), .Z(n16504) );
  XNOR U16767 ( .A(n16512), .B(n16720), .Z(n16505) );
  XNOR U16768 ( .A(n16511), .B(n16509), .Z(n16720) );
  AND U16769 ( .A(n16721), .B(n16722), .Z(n16509) );
  NANDN U16770 ( .A(n16723), .B(n16724), .Z(n16722) );
  NANDN U16771 ( .A(n16725), .B(n16726), .Z(n16724) );
  NANDN U16772 ( .A(n16726), .B(n16725), .Z(n16721) );
  ANDN U16773 ( .B(B[235]), .A(n64), .Z(n16511) );
  XNOR U16774 ( .A(n16519), .B(n16727), .Z(n16512) );
  XNOR U16775 ( .A(n16518), .B(n16516), .Z(n16727) );
  AND U16776 ( .A(n16728), .B(n16729), .Z(n16516) );
  NANDN U16777 ( .A(n16730), .B(n16731), .Z(n16729) );
  OR U16778 ( .A(n16732), .B(n16733), .Z(n16731) );
  NAND U16779 ( .A(n16733), .B(n16732), .Z(n16728) );
  ANDN U16780 ( .B(B[236]), .A(n65), .Z(n16518) );
  XNOR U16781 ( .A(n16526), .B(n16734), .Z(n16519) );
  XNOR U16782 ( .A(n16525), .B(n16523), .Z(n16734) );
  AND U16783 ( .A(n16735), .B(n16736), .Z(n16523) );
  NANDN U16784 ( .A(n16737), .B(n16738), .Z(n16736) );
  NANDN U16785 ( .A(n16739), .B(n16740), .Z(n16738) );
  NANDN U16786 ( .A(n16740), .B(n16739), .Z(n16735) );
  ANDN U16787 ( .B(B[237]), .A(n66), .Z(n16525) );
  XNOR U16788 ( .A(n16533), .B(n16741), .Z(n16526) );
  XNOR U16789 ( .A(n16532), .B(n16530), .Z(n16741) );
  AND U16790 ( .A(n16742), .B(n16743), .Z(n16530) );
  NANDN U16791 ( .A(n16744), .B(n16745), .Z(n16743) );
  OR U16792 ( .A(n16746), .B(n16747), .Z(n16745) );
  NAND U16793 ( .A(n16747), .B(n16746), .Z(n16742) );
  ANDN U16794 ( .B(B[238]), .A(n67), .Z(n16532) );
  XNOR U16795 ( .A(n16540), .B(n16748), .Z(n16533) );
  XNOR U16796 ( .A(n16539), .B(n16537), .Z(n16748) );
  AND U16797 ( .A(n16749), .B(n16750), .Z(n16537) );
  NANDN U16798 ( .A(n16751), .B(n16752), .Z(n16750) );
  NANDN U16799 ( .A(n16753), .B(n16754), .Z(n16752) );
  NANDN U16800 ( .A(n16754), .B(n16753), .Z(n16749) );
  ANDN U16801 ( .B(B[239]), .A(n68), .Z(n16539) );
  XNOR U16802 ( .A(n16547), .B(n16755), .Z(n16540) );
  XNOR U16803 ( .A(n16546), .B(n16544), .Z(n16755) );
  AND U16804 ( .A(n16756), .B(n16757), .Z(n16544) );
  NANDN U16805 ( .A(n16758), .B(n16759), .Z(n16757) );
  OR U16806 ( .A(n16760), .B(n16761), .Z(n16759) );
  NAND U16807 ( .A(n16761), .B(n16760), .Z(n16756) );
  ANDN U16808 ( .B(B[240]), .A(n69), .Z(n16546) );
  XNOR U16809 ( .A(n16554), .B(n16762), .Z(n16547) );
  XNOR U16810 ( .A(n16553), .B(n16551), .Z(n16762) );
  AND U16811 ( .A(n16763), .B(n16764), .Z(n16551) );
  NANDN U16812 ( .A(n16765), .B(n16766), .Z(n16764) );
  NANDN U16813 ( .A(n16767), .B(n16768), .Z(n16766) );
  NANDN U16814 ( .A(n16768), .B(n16767), .Z(n16763) );
  ANDN U16815 ( .B(B[241]), .A(n70), .Z(n16553) );
  XNOR U16816 ( .A(n16561), .B(n16769), .Z(n16554) );
  XNOR U16817 ( .A(n16560), .B(n16558), .Z(n16769) );
  AND U16818 ( .A(n16770), .B(n16771), .Z(n16558) );
  NANDN U16819 ( .A(n16772), .B(n16773), .Z(n16771) );
  OR U16820 ( .A(n16774), .B(n16775), .Z(n16773) );
  NAND U16821 ( .A(n16775), .B(n16774), .Z(n16770) );
  ANDN U16822 ( .B(B[242]), .A(n71), .Z(n16560) );
  XNOR U16823 ( .A(n16568), .B(n16776), .Z(n16561) );
  XNOR U16824 ( .A(n16567), .B(n16565), .Z(n16776) );
  AND U16825 ( .A(n16777), .B(n16778), .Z(n16565) );
  NANDN U16826 ( .A(n16779), .B(n16780), .Z(n16778) );
  NANDN U16827 ( .A(n16781), .B(n16782), .Z(n16780) );
  NANDN U16828 ( .A(n16782), .B(n16781), .Z(n16777) );
  ANDN U16829 ( .B(B[243]), .A(n72), .Z(n16567) );
  XNOR U16830 ( .A(n16575), .B(n16783), .Z(n16568) );
  XNOR U16831 ( .A(n16574), .B(n16572), .Z(n16783) );
  AND U16832 ( .A(n16784), .B(n16785), .Z(n16572) );
  NANDN U16833 ( .A(n16786), .B(n16787), .Z(n16785) );
  OR U16834 ( .A(n16788), .B(n16789), .Z(n16787) );
  NAND U16835 ( .A(n16789), .B(n16788), .Z(n16784) );
  ANDN U16836 ( .B(B[244]), .A(n73), .Z(n16574) );
  XNOR U16837 ( .A(n16582), .B(n16790), .Z(n16575) );
  XNOR U16838 ( .A(n16581), .B(n16579), .Z(n16790) );
  AND U16839 ( .A(n16791), .B(n16792), .Z(n16579) );
  NANDN U16840 ( .A(n16793), .B(n16794), .Z(n16792) );
  NANDN U16841 ( .A(n16795), .B(n16796), .Z(n16794) );
  NANDN U16842 ( .A(n16796), .B(n16795), .Z(n16791) );
  ANDN U16843 ( .B(B[245]), .A(n74), .Z(n16581) );
  XNOR U16844 ( .A(n16589), .B(n16797), .Z(n16582) );
  XNOR U16845 ( .A(n16588), .B(n16586), .Z(n16797) );
  AND U16846 ( .A(n16798), .B(n16799), .Z(n16586) );
  NANDN U16847 ( .A(n16800), .B(n16801), .Z(n16799) );
  OR U16848 ( .A(n16802), .B(n16803), .Z(n16801) );
  NAND U16849 ( .A(n16803), .B(n16802), .Z(n16798) );
  ANDN U16850 ( .B(B[246]), .A(n75), .Z(n16588) );
  XNOR U16851 ( .A(n16596), .B(n16804), .Z(n16589) );
  XNOR U16852 ( .A(n16595), .B(n16593), .Z(n16804) );
  AND U16853 ( .A(n16805), .B(n16806), .Z(n16593) );
  NANDN U16854 ( .A(n16807), .B(n16808), .Z(n16806) );
  NANDN U16855 ( .A(n16809), .B(n16810), .Z(n16808) );
  NANDN U16856 ( .A(n16810), .B(n16809), .Z(n16805) );
  ANDN U16857 ( .B(B[247]), .A(n76), .Z(n16595) );
  XNOR U16858 ( .A(n16603), .B(n16811), .Z(n16596) );
  XNOR U16859 ( .A(n16602), .B(n16600), .Z(n16811) );
  AND U16860 ( .A(n16812), .B(n16813), .Z(n16600) );
  NANDN U16861 ( .A(n16814), .B(n16815), .Z(n16813) );
  OR U16862 ( .A(n16816), .B(n16817), .Z(n16815) );
  NAND U16863 ( .A(n16817), .B(n16816), .Z(n16812) );
  ANDN U16864 ( .B(B[248]), .A(n77), .Z(n16602) );
  XNOR U16865 ( .A(n16610), .B(n16818), .Z(n16603) );
  XNOR U16866 ( .A(n16609), .B(n16607), .Z(n16818) );
  AND U16867 ( .A(n16819), .B(n16820), .Z(n16607) );
  NANDN U16868 ( .A(n16821), .B(n16822), .Z(n16820) );
  NANDN U16869 ( .A(n16823), .B(n16824), .Z(n16822) );
  NANDN U16870 ( .A(n16824), .B(n16823), .Z(n16819) );
  ANDN U16871 ( .B(B[249]), .A(n78), .Z(n16609) );
  XNOR U16872 ( .A(n16617), .B(n16825), .Z(n16610) );
  XNOR U16873 ( .A(n16616), .B(n16614), .Z(n16825) );
  AND U16874 ( .A(n16826), .B(n16827), .Z(n16614) );
  NANDN U16875 ( .A(n16828), .B(n16829), .Z(n16827) );
  OR U16876 ( .A(n16830), .B(n16831), .Z(n16829) );
  NAND U16877 ( .A(n16831), .B(n16830), .Z(n16826) );
  ANDN U16878 ( .B(B[250]), .A(n79), .Z(n16616) );
  XNOR U16879 ( .A(n16624), .B(n16832), .Z(n16617) );
  XNOR U16880 ( .A(n16623), .B(n16621), .Z(n16832) );
  AND U16881 ( .A(n16833), .B(n16834), .Z(n16621) );
  NANDN U16882 ( .A(n16835), .B(n16836), .Z(n16834) );
  NANDN U16883 ( .A(n16837), .B(n16838), .Z(n16836) );
  NANDN U16884 ( .A(n16838), .B(n16837), .Z(n16833) );
  ANDN U16885 ( .B(B[251]), .A(n80), .Z(n16623) );
  XNOR U16886 ( .A(n16631), .B(n16839), .Z(n16624) );
  XNOR U16887 ( .A(n16630), .B(n16628), .Z(n16839) );
  AND U16888 ( .A(n16840), .B(n16841), .Z(n16628) );
  NANDN U16889 ( .A(n16842), .B(n16843), .Z(n16841) );
  OR U16890 ( .A(n16844), .B(n16845), .Z(n16843) );
  NAND U16891 ( .A(n16845), .B(n16844), .Z(n16840) );
  ANDN U16892 ( .B(B[252]), .A(n81), .Z(n16630) );
  XNOR U16893 ( .A(n3), .B(n16846), .Z(n16631) );
  XNOR U16894 ( .A(n16637), .B(n16635), .Z(n16846) );
  AND U16895 ( .A(n16847), .B(n16848), .Z(n16635) );
  NANDN U16896 ( .A(n16849), .B(n16850), .Z(n16848) );
  NAND U16897 ( .A(n16851), .B(n16852), .Z(n16850) );
  ANDN U16898 ( .B(B[253]), .A(n82), .Z(n16637) );
  XNOR U16899 ( .A(n16643), .B(n16853), .Z(n16638) );
  XNOR U16900 ( .A(n16641), .B(n16642), .Z(n16853) );
  NAND U16901 ( .A(A[2]), .B(B[254]), .Z(n16642) );
  ANDN U16902 ( .B(A[0]), .A(n16855), .Z(n16854) );
  NAND U16903 ( .A(B[255]), .B(A[1]), .Z(n16643) );
  NAND U16904 ( .A(n16856), .B(n16857), .Z(n284) );
  NANDN U16905 ( .A(n16858), .B(n16859), .Z(n16857) );
  OR U16906 ( .A(n16860), .B(n16861), .Z(n16859) );
  NAND U16907 ( .A(n16861), .B(n16860), .Z(n16856) );
  XOR U16908 ( .A(n286), .B(n285), .Z(\A1[253] ) );
  XOR U16909 ( .A(n16861), .B(n16862), .Z(n285) );
  XNOR U16910 ( .A(n16860), .B(n16858), .Z(n16862) );
  AND U16911 ( .A(n16863), .B(n16864), .Z(n16858) );
  NANDN U16912 ( .A(n16865), .B(n16866), .Z(n16864) );
  NANDN U16913 ( .A(n16867), .B(n16868), .Z(n16866) );
  NANDN U16914 ( .A(n16868), .B(n16867), .Z(n16863) );
  ANDN U16915 ( .B(B[224]), .A(n54), .Z(n16860) );
  XNOR U16916 ( .A(n16656), .B(n16869), .Z(n16861) );
  XNOR U16917 ( .A(n16655), .B(n16653), .Z(n16869) );
  AND U16918 ( .A(n16870), .B(n16871), .Z(n16653) );
  NANDN U16919 ( .A(n16872), .B(n16873), .Z(n16871) );
  OR U16920 ( .A(n16874), .B(n16875), .Z(n16873) );
  NAND U16921 ( .A(n16875), .B(n16874), .Z(n16870) );
  ANDN U16922 ( .B(B[225]), .A(n55), .Z(n16655) );
  XNOR U16923 ( .A(n16663), .B(n16876), .Z(n16656) );
  XNOR U16924 ( .A(n16662), .B(n16660), .Z(n16876) );
  AND U16925 ( .A(n16877), .B(n16878), .Z(n16660) );
  NANDN U16926 ( .A(n16879), .B(n16880), .Z(n16878) );
  NANDN U16927 ( .A(n16881), .B(n16882), .Z(n16880) );
  NANDN U16928 ( .A(n16882), .B(n16881), .Z(n16877) );
  ANDN U16929 ( .B(B[226]), .A(n56), .Z(n16662) );
  XNOR U16930 ( .A(n16670), .B(n16883), .Z(n16663) );
  XNOR U16931 ( .A(n16669), .B(n16667), .Z(n16883) );
  AND U16932 ( .A(n16884), .B(n16885), .Z(n16667) );
  NANDN U16933 ( .A(n16886), .B(n16887), .Z(n16885) );
  OR U16934 ( .A(n16888), .B(n16889), .Z(n16887) );
  NAND U16935 ( .A(n16889), .B(n16888), .Z(n16884) );
  ANDN U16936 ( .B(B[227]), .A(n57), .Z(n16669) );
  XNOR U16937 ( .A(n16677), .B(n16890), .Z(n16670) );
  XNOR U16938 ( .A(n16676), .B(n16674), .Z(n16890) );
  AND U16939 ( .A(n16891), .B(n16892), .Z(n16674) );
  NANDN U16940 ( .A(n16893), .B(n16894), .Z(n16892) );
  NANDN U16941 ( .A(n16895), .B(n16896), .Z(n16894) );
  NANDN U16942 ( .A(n16896), .B(n16895), .Z(n16891) );
  ANDN U16943 ( .B(B[228]), .A(n58), .Z(n16676) );
  XNOR U16944 ( .A(n16684), .B(n16897), .Z(n16677) );
  XNOR U16945 ( .A(n16683), .B(n16681), .Z(n16897) );
  AND U16946 ( .A(n16898), .B(n16899), .Z(n16681) );
  NANDN U16947 ( .A(n16900), .B(n16901), .Z(n16899) );
  OR U16948 ( .A(n16902), .B(n16903), .Z(n16901) );
  NAND U16949 ( .A(n16903), .B(n16902), .Z(n16898) );
  ANDN U16950 ( .B(B[229]), .A(n59), .Z(n16683) );
  XNOR U16951 ( .A(n16691), .B(n16904), .Z(n16684) );
  XNOR U16952 ( .A(n16690), .B(n16688), .Z(n16904) );
  AND U16953 ( .A(n16905), .B(n16906), .Z(n16688) );
  NANDN U16954 ( .A(n16907), .B(n16908), .Z(n16906) );
  NANDN U16955 ( .A(n16909), .B(n16910), .Z(n16908) );
  NANDN U16956 ( .A(n16910), .B(n16909), .Z(n16905) );
  ANDN U16957 ( .B(B[230]), .A(n60), .Z(n16690) );
  XNOR U16958 ( .A(n16698), .B(n16911), .Z(n16691) );
  XNOR U16959 ( .A(n16697), .B(n16695), .Z(n16911) );
  AND U16960 ( .A(n16912), .B(n16913), .Z(n16695) );
  NANDN U16961 ( .A(n16914), .B(n16915), .Z(n16913) );
  OR U16962 ( .A(n16916), .B(n16917), .Z(n16915) );
  NAND U16963 ( .A(n16917), .B(n16916), .Z(n16912) );
  ANDN U16964 ( .B(B[231]), .A(n61), .Z(n16697) );
  XNOR U16965 ( .A(n16705), .B(n16918), .Z(n16698) );
  XNOR U16966 ( .A(n16704), .B(n16702), .Z(n16918) );
  AND U16967 ( .A(n16919), .B(n16920), .Z(n16702) );
  NANDN U16968 ( .A(n16921), .B(n16922), .Z(n16920) );
  NANDN U16969 ( .A(n16923), .B(n16924), .Z(n16922) );
  NANDN U16970 ( .A(n16924), .B(n16923), .Z(n16919) );
  ANDN U16971 ( .B(B[232]), .A(n62), .Z(n16704) );
  XNOR U16972 ( .A(n16712), .B(n16925), .Z(n16705) );
  XNOR U16973 ( .A(n16711), .B(n16709), .Z(n16925) );
  AND U16974 ( .A(n16926), .B(n16927), .Z(n16709) );
  NANDN U16975 ( .A(n16928), .B(n16929), .Z(n16927) );
  OR U16976 ( .A(n16930), .B(n16931), .Z(n16929) );
  NAND U16977 ( .A(n16931), .B(n16930), .Z(n16926) );
  ANDN U16978 ( .B(B[233]), .A(n63), .Z(n16711) );
  XNOR U16979 ( .A(n16719), .B(n16932), .Z(n16712) );
  XNOR U16980 ( .A(n16718), .B(n16716), .Z(n16932) );
  AND U16981 ( .A(n16933), .B(n16934), .Z(n16716) );
  NANDN U16982 ( .A(n16935), .B(n16936), .Z(n16934) );
  NANDN U16983 ( .A(n16937), .B(n16938), .Z(n16936) );
  NANDN U16984 ( .A(n16938), .B(n16937), .Z(n16933) );
  ANDN U16985 ( .B(B[234]), .A(n64), .Z(n16718) );
  XNOR U16986 ( .A(n16726), .B(n16939), .Z(n16719) );
  XNOR U16987 ( .A(n16725), .B(n16723), .Z(n16939) );
  AND U16988 ( .A(n16940), .B(n16941), .Z(n16723) );
  NANDN U16989 ( .A(n16942), .B(n16943), .Z(n16941) );
  OR U16990 ( .A(n16944), .B(n16945), .Z(n16943) );
  NAND U16991 ( .A(n16945), .B(n16944), .Z(n16940) );
  ANDN U16992 ( .B(B[235]), .A(n65), .Z(n16725) );
  XNOR U16993 ( .A(n16733), .B(n16946), .Z(n16726) );
  XNOR U16994 ( .A(n16732), .B(n16730), .Z(n16946) );
  AND U16995 ( .A(n16947), .B(n16948), .Z(n16730) );
  NANDN U16996 ( .A(n16949), .B(n16950), .Z(n16948) );
  NANDN U16997 ( .A(n16951), .B(n16952), .Z(n16950) );
  NANDN U16998 ( .A(n16952), .B(n16951), .Z(n16947) );
  ANDN U16999 ( .B(B[236]), .A(n66), .Z(n16732) );
  XNOR U17000 ( .A(n16740), .B(n16953), .Z(n16733) );
  XNOR U17001 ( .A(n16739), .B(n16737), .Z(n16953) );
  AND U17002 ( .A(n16954), .B(n16955), .Z(n16737) );
  NANDN U17003 ( .A(n16956), .B(n16957), .Z(n16955) );
  OR U17004 ( .A(n16958), .B(n16959), .Z(n16957) );
  NAND U17005 ( .A(n16959), .B(n16958), .Z(n16954) );
  ANDN U17006 ( .B(B[237]), .A(n67), .Z(n16739) );
  XNOR U17007 ( .A(n16747), .B(n16960), .Z(n16740) );
  XNOR U17008 ( .A(n16746), .B(n16744), .Z(n16960) );
  AND U17009 ( .A(n16961), .B(n16962), .Z(n16744) );
  NANDN U17010 ( .A(n16963), .B(n16964), .Z(n16962) );
  NANDN U17011 ( .A(n16965), .B(n16966), .Z(n16964) );
  NANDN U17012 ( .A(n16966), .B(n16965), .Z(n16961) );
  ANDN U17013 ( .B(B[238]), .A(n68), .Z(n16746) );
  XNOR U17014 ( .A(n16754), .B(n16967), .Z(n16747) );
  XNOR U17015 ( .A(n16753), .B(n16751), .Z(n16967) );
  AND U17016 ( .A(n16968), .B(n16969), .Z(n16751) );
  NANDN U17017 ( .A(n16970), .B(n16971), .Z(n16969) );
  OR U17018 ( .A(n16972), .B(n16973), .Z(n16971) );
  NAND U17019 ( .A(n16973), .B(n16972), .Z(n16968) );
  ANDN U17020 ( .B(B[239]), .A(n69), .Z(n16753) );
  XNOR U17021 ( .A(n16761), .B(n16974), .Z(n16754) );
  XNOR U17022 ( .A(n16760), .B(n16758), .Z(n16974) );
  AND U17023 ( .A(n16975), .B(n16976), .Z(n16758) );
  NANDN U17024 ( .A(n16977), .B(n16978), .Z(n16976) );
  NANDN U17025 ( .A(n16979), .B(n16980), .Z(n16978) );
  NANDN U17026 ( .A(n16980), .B(n16979), .Z(n16975) );
  ANDN U17027 ( .B(B[240]), .A(n70), .Z(n16760) );
  XNOR U17028 ( .A(n16768), .B(n16981), .Z(n16761) );
  XNOR U17029 ( .A(n16767), .B(n16765), .Z(n16981) );
  AND U17030 ( .A(n16982), .B(n16983), .Z(n16765) );
  NANDN U17031 ( .A(n16984), .B(n16985), .Z(n16983) );
  OR U17032 ( .A(n16986), .B(n16987), .Z(n16985) );
  NAND U17033 ( .A(n16987), .B(n16986), .Z(n16982) );
  ANDN U17034 ( .B(B[241]), .A(n71), .Z(n16767) );
  XNOR U17035 ( .A(n16775), .B(n16988), .Z(n16768) );
  XNOR U17036 ( .A(n16774), .B(n16772), .Z(n16988) );
  AND U17037 ( .A(n16989), .B(n16990), .Z(n16772) );
  NANDN U17038 ( .A(n16991), .B(n16992), .Z(n16990) );
  NANDN U17039 ( .A(n16993), .B(n16994), .Z(n16992) );
  NANDN U17040 ( .A(n16994), .B(n16993), .Z(n16989) );
  ANDN U17041 ( .B(B[242]), .A(n72), .Z(n16774) );
  XNOR U17042 ( .A(n16782), .B(n16995), .Z(n16775) );
  XNOR U17043 ( .A(n16781), .B(n16779), .Z(n16995) );
  AND U17044 ( .A(n16996), .B(n16997), .Z(n16779) );
  NANDN U17045 ( .A(n16998), .B(n16999), .Z(n16997) );
  OR U17046 ( .A(n17000), .B(n17001), .Z(n16999) );
  NAND U17047 ( .A(n17001), .B(n17000), .Z(n16996) );
  ANDN U17048 ( .B(B[243]), .A(n73), .Z(n16781) );
  XNOR U17049 ( .A(n16789), .B(n17002), .Z(n16782) );
  XNOR U17050 ( .A(n16788), .B(n16786), .Z(n17002) );
  AND U17051 ( .A(n17003), .B(n17004), .Z(n16786) );
  NANDN U17052 ( .A(n17005), .B(n17006), .Z(n17004) );
  NANDN U17053 ( .A(n17007), .B(n17008), .Z(n17006) );
  NANDN U17054 ( .A(n17008), .B(n17007), .Z(n17003) );
  ANDN U17055 ( .B(B[244]), .A(n74), .Z(n16788) );
  XNOR U17056 ( .A(n16796), .B(n17009), .Z(n16789) );
  XNOR U17057 ( .A(n16795), .B(n16793), .Z(n17009) );
  AND U17058 ( .A(n17010), .B(n17011), .Z(n16793) );
  NANDN U17059 ( .A(n17012), .B(n17013), .Z(n17011) );
  OR U17060 ( .A(n17014), .B(n17015), .Z(n17013) );
  NAND U17061 ( .A(n17015), .B(n17014), .Z(n17010) );
  ANDN U17062 ( .B(B[245]), .A(n75), .Z(n16795) );
  XNOR U17063 ( .A(n16803), .B(n17016), .Z(n16796) );
  XNOR U17064 ( .A(n16802), .B(n16800), .Z(n17016) );
  AND U17065 ( .A(n17017), .B(n17018), .Z(n16800) );
  NANDN U17066 ( .A(n17019), .B(n17020), .Z(n17018) );
  NANDN U17067 ( .A(n17021), .B(n17022), .Z(n17020) );
  NANDN U17068 ( .A(n17022), .B(n17021), .Z(n17017) );
  ANDN U17069 ( .B(B[246]), .A(n76), .Z(n16802) );
  XNOR U17070 ( .A(n16810), .B(n17023), .Z(n16803) );
  XNOR U17071 ( .A(n16809), .B(n16807), .Z(n17023) );
  AND U17072 ( .A(n17024), .B(n17025), .Z(n16807) );
  NANDN U17073 ( .A(n17026), .B(n17027), .Z(n17025) );
  OR U17074 ( .A(n17028), .B(n17029), .Z(n17027) );
  NAND U17075 ( .A(n17029), .B(n17028), .Z(n17024) );
  ANDN U17076 ( .B(B[247]), .A(n77), .Z(n16809) );
  XNOR U17077 ( .A(n16817), .B(n17030), .Z(n16810) );
  XNOR U17078 ( .A(n16816), .B(n16814), .Z(n17030) );
  AND U17079 ( .A(n17031), .B(n17032), .Z(n16814) );
  NANDN U17080 ( .A(n17033), .B(n17034), .Z(n17032) );
  NANDN U17081 ( .A(n17035), .B(n17036), .Z(n17034) );
  NANDN U17082 ( .A(n17036), .B(n17035), .Z(n17031) );
  ANDN U17083 ( .B(B[248]), .A(n78), .Z(n16816) );
  XNOR U17084 ( .A(n16824), .B(n17037), .Z(n16817) );
  XNOR U17085 ( .A(n16823), .B(n16821), .Z(n17037) );
  AND U17086 ( .A(n17038), .B(n17039), .Z(n16821) );
  NANDN U17087 ( .A(n17040), .B(n17041), .Z(n17039) );
  OR U17088 ( .A(n17042), .B(n17043), .Z(n17041) );
  NAND U17089 ( .A(n17043), .B(n17042), .Z(n17038) );
  ANDN U17090 ( .B(B[249]), .A(n79), .Z(n16823) );
  XNOR U17091 ( .A(n16831), .B(n17044), .Z(n16824) );
  XNOR U17092 ( .A(n16830), .B(n16828), .Z(n17044) );
  AND U17093 ( .A(n17045), .B(n17046), .Z(n16828) );
  NANDN U17094 ( .A(n17047), .B(n17048), .Z(n17046) );
  NANDN U17095 ( .A(n17049), .B(n17050), .Z(n17048) );
  NANDN U17096 ( .A(n17050), .B(n17049), .Z(n17045) );
  ANDN U17097 ( .B(B[250]), .A(n80), .Z(n16830) );
  XNOR U17098 ( .A(n16838), .B(n17051), .Z(n16831) );
  XNOR U17099 ( .A(n16837), .B(n16835), .Z(n17051) );
  AND U17100 ( .A(n17052), .B(n17053), .Z(n16835) );
  NANDN U17101 ( .A(n17054), .B(n17055), .Z(n17053) );
  OR U17102 ( .A(n17056), .B(n17057), .Z(n17055) );
  NAND U17103 ( .A(n17057), .B(n17056), .Z(n17052) );
  ANDN U17104 ( .B(B[251]), .A(n81), .Z(n16837) );
  XNOR U17105 ( .A(n16845), .B(n17058), .Z(n16838) );
  XNOR U17106 ( .A(n16844), .B(n16842), .Z(n17058) );
  AND U17107 ( .A(n17059), .B(n17060), .Z(n16842) );
  NANDN U17108 ( .A(n17061), .B(n17062), .Z(n17060) );
  NAND U17109 ( .A(n17063), .B(n17064), .Z(n17062) );
  ANDN U17110 ( .B(B[252]), .A(n82), .Z(n16844) );
  XOR U17111 ( .A(n16851), .B(n17065), .Z(n16845) );
  XNOR U17112 ( .A(n16849), .B(n16852), .Z(n17065) );
  NAND U17113 ( .A(A[2]), .B(B[253]), .Z(n16852) );
  NANDN U17114 ( .A(n17066), .B(n17067), .Z(n16849) );
  AND U17115 ( .A(A[0]), .B(B[254]), .Z(n17067) );
  XNOR U17116 ( .A(n16855), .B(n17068), .Z(n16851) );
  NAND U17117 ( .A(B[255]), .B(A[0]), .Z(n17068) );
  NAND U17118 ( .A(B[254]), .B(A[1]), .Z(n16855) );
  NAND U17119 ( .A(n17069), .B(n17070), .Z(n286) );
  NANDN U17120 ( .A(n17071), .B(n17072), .Z(n17070) );
  OR U17121 ( .A(n17073), .B(n17074), .Z(n17072) );
  NAND U17122 ( .A(n17074), .B(n17073), .Z(n17069) );
  XOR U17123 ( .A(n288), .B(n287), .Z(\A1[252] ) );
  XOR U17124 ( .A(n17074), .B(n17075), .Z(n287) );
  XNOR U17125 ( .A(n17073), .B(n17071), .Z(n17075) );
  AND U17126 ( .A(n17076), .B(n17077), .Z(n17071) );
  NANDN U17127 ( .A(n17078), .B(n17079), .Z(n17077) );
  NANDN U17128 ( .A(n17080), .B(n17081), .Z(n17079) );
  NANDN U17129 ( .A(n17081), .B(n17080), .Z(n17076) );
  ANDN U17130 ( .B(B[223]), .A(n54), .Z(n17073) );
  XNOR U17131 ( .A(n16868), .B(n17082), .Z(n17074) );
  XNOR U17132 ( .A(n16867), .B(n16865), .Z(n17082) );
  AND U17133 ( .A(n17083), .B(n17084), .Z(n16865) );
  NANDN U17134 ( .A(n17085), .B(n17086), .Z(n17084) );
  OR U17135 ( .A(n17087), .B(n17088), .Z(n17086) );
  NAND U17136 ( .A(n17088), .B(n17087), .Z(n17083) );
  ANDN U17137 ( .B(B[224]), .A(n55), .Z(n16867) );
  XNOR U17138 ( .A(n16875), .B(n17089), .Z(n16868) );
  XNOR U17139 ( .A(n16874), .B(n16872), .Z(n17089) );
  AND U17140 ( .A(n17090), .B(n17091), .Z(n16872) );
  NANDN U17141 ( .A(n17092), .B(n17093), .Z(n17091) );
  NANDN U17142 ( .A(n17094), .B(n17095), .Z(n17093) );
  NANDN U17143 ( .A(n17095), .B(n17094), .Z(n17090) );
  ANDN U17144 ( .B(B[225]), .A(n56), .Z(n16874) );
  XNOR U17145 ( .A(n16882), .B(n17096), .Z(n16875) );
  XNOR U17146 ( .A(n16881), .B(n16879), .Z(n17096) );
  AND U17147 ( .A(n17097), .B(n17098), .Z(n16879) );
  NANDN U17148 ( .A(n17099), .B(n17100), .Z(n17098) );
  OR U17149 ( .A(n17101), .B(n17102), .Z(n17100) );
  NAND U17150 ( .A(n17102), .B(n17101), .Z(n17097) );
  ANDN U17151 ( .B(B[226]), .A(n57), .Z(n16881) );
  XNOR U17152 ( .A(n16889), .B(n17103), .Z(n16882) );
  XNOR U17153 ( .A(n16888), .B(n16886), .Z(n17103) );
  AND U17154 ( .A(n17104), .B(n17105), .Z(n16886) );
  NANDN U17155 ( .A(n17106), .B(n17107), .Z(n17105) );
  NANDN U17156 ( .A(n17108), .B(n17109), .Z(n17107) );
  NANDN U17157 ( .A(n17109), .B(n17108), .Z(n17104) );
  ANDN U17158 ( .B(B[227]), .A(n58), .Z(n16888) );
  XNOR U17159 ( .A(n16896), .B(n17110), .Z(n16889) );
  XNOR U17160 ( .A(n16895), .B(n16893), .Z(n17110) );
  AND U17161 ( .A(n17111), .B(n17112), .Z(n16893) );
  NANDN U17162 ( .A(n17113), .B(n17114), .Z(n17112) );
  OR U17163 ( .A(n17115), .B(n17116), .Z(n17114) );
  NAND U17164 ( .A(n17116), .B(n17115), .Z(n17111) );
  ANDN U17165 ( .B(B[228]), .A(n59), .Z(n16895) );
  XNOR U17166 ( .A(n16903), .B(n17117), .Z(n16896) );
  XNOR U17167 ( .A(n16902), .B(n16900), .Z(n17117) );
  AND U17168 ( .A(n17118), .B(n17119), .Z(n16900) );
  NANDN U17169 ( .A(n17120), .B(n17121), .Z(n17119) );
  NANDN U17170 ( .A(n17122), .B(n17123), .Z(n17121) );
  NANDN U17171 ( .A(n17123), .B(n17122), .Z(n17118) );
  ANDN U17172 ( .B(B[229]), .A(n60), .Z(n16902) );
  XNOR U17173 ( .A(n16910), .B(n17124), .Z(n16903) );
  XNOR U17174 ( .A(n16909), .B(n16907), .Z(n17124) );
  AND U17175 ( .A(n17125), .B(n17126), .Z(n16907) );
  NANDN U17176 ( .A(n17127), .B(n17128), .Z(n17126) );
  OR U17177 ( .A(n17129), .B(n17130), .Z(n17128) );
  NAND U17178 ( .A(n17130), .B(n17129), .Z(n17125) );
  ANDN U17179 ( .B(B[230]), .A(n61), .Z(n16909) );
  XNOR U17180 ( .A(n16917), .B(n17131), .Z(n16910) );
  XNOR U17181 ( .A(n16916), .B(n16914), .Z(n17131) );
  AND U17182 ( .A(n17132), .B(n17133), .Z(n16914) );
  NANDN U17183 ( .A(n17134), .B(n17135), .Z(n17133) );
  NANDN U17184 ( .A(n17136), .B(n17137), .Z(n17135) );
  NANDN U17185 ( .A(n17137), .B(n17136), .Z(n17132) );
  ANDN U17186 ( .B(B[231]), .A(n62), .Z(n16916) );
  XNOR U17187 ( .A(n16924), .B(n17138), .Z(n16917) );
  XNOR U17188 ( .A(n16923), .B(n16921), .Z(n17138) );
  AND U17189 ( .A(n17139), .B(n17140), .Z(n16921) );
  NANDN U17190 ( .A(n17141), .B(n17142), .Z(n17140) );
  OR U17191 ( .A(n17143), .B(n17144), .Z(n17142) );
  NAND U17192 ( .A(n17144), .B(n17143), .Z(n17139) );
  ANDN U17193 ( .B(B[232]), .A(n63), .Z(n16923) );
  XNOR U17194 ( .A(n16931), .B(n17145), .Z(n16924) );
  XNOR U17195 ( .A(n16930), .B(n16928), .Z(n17145) );
  AND U17196 ( .A(n17146), .B(n17147), .Z(n16928) );
  NANDN U17197 ( .A(n17148), .B(n17149), .Z(n17147) );
  NANDN U17198 ( .A(n17150), .B(n17151), .Z(n17149) );
  NANDN U17199 ( .A(n17151), .B(n17150), .Z(n17146) );
  ANDN U17200 ( .B(B[233]), .A(n64), .Z(n16930) );
  XNOR U17201 ( .A(n16938), .B(n17152), .Z(n16931) );
  XNOR U17202 ( .A(n16937), .B(n16935), .Z(n17152) );
  AND U17203 ( .A(n17153), .B(n17154), .Z(n16935) );
  NANDN U17204 ( .A(n17155), .B(n17156), .Z(n17154) );
  OR U17205 ( .A(n17157), .B(n17158), .Z(n17156) );
  NAND U17206 ( .A(n17158), .B(n17157), .Z(n17153) );
  ANDN U17207 ( .B(B[234]), .A(n65), .Z(n16937) );
  XNOR U17208 ( .A(n16945), .B(n17159), .Z(n16938) );
  XNOR U17209 ( .A(n16944), .B(n16942), .Z(n17159) );
  AND U17210 ( .A(n17160), .B(n17161), .Z(n16942) );
  NANDN U17211 ( .A(n17162), .B(n17163), .Z(n17161) );
  NANDN U17212 ( .A(n17164), .B(n17165), .Z(n17163) );
  NANDN U17213 ( .A(n17165), .B(n17164), .Z(n17160) );
  ANDN U17214 ( .B(B[235]), .A(n66), .Z(n16944) );
  XNOR U17215 ( .A(n16952), .B(n17166), .Z(n16945) );
  XNOR U17216 ( .A(n16951), .B(n16949), .Z(n17166) );
  AND U17217 ( .A(n17167), .B(n17168), .Z(n16949) );
  NANDN U17218 ( .A(n17169), .B(n17170), .Z(n17168) );
  OR U17219 ( .A(n17171), .B(n17172), .Z(n17170) );
  NAND U17220 ( .A(n17172), .B(n17171), .Z(n17167) );
  ANDN U17221 ( .B(B[236]), .A(n67), .Z(n16951) );
  XNOR U17222 ( .A(n16959), .B(n17173), .Z(n16952) );
  XNOR U17223 ( .A(n16958), .B(n16956), .Z(n17173) );
  AND U17224 ( .A(n17174), .B(n17175), .Z(n16956) );
  NANDN U17225 ( .A(n17176), .B(n17177), .Z(n17175) );
  NANDN U17226 ( .A(n17178), .B(n17179), .Z(n17177) );
  NANDN U17227 ( .A(n17179), .B(n17178), .Z(n17174) );
  ANDN U17228 ( .B(B[237]), .A(n68), .Z(n16958) );
  XNOR U17229 ( .A(n16966), .B(n17180), .Z(n16959) );
  XNOR U17230 ( .A(n16965), .B(n16963), .Z(n17180) );
  AND U17231 ( .A(n17181), .B(n17182), .Z(n16963) );
  NANDN U17232 ( .A(n17183), .B(n17184), .Z(n17182) );
  OR U17233 ( .A(n17185), .B(n17186), .Z(n17184) );
  NAND U17234 ( .A(n17186), .B(n17185), .Z(n17181) );
  ANDN U17235 ( .B(B[238]), .A(n69), .Z(n16965) );
  XNOR U17236 ( .A(n16973), .B(n17187), .Z(n16966) );
  XNOR U17237 ( .A(n16972), .B(n16970), .Z(n17187) );
  AND U17238 ( .A(n17188), .B(n17189), .Z(n16970) );
  NANDN U17239 ( .A(n17190), .B(n17191), .Z(n17189) );
  NANDN U17240 ( .A(n17192), .B(n17193), .Z(n17191) );
  NANDN U17241 ( .A(n17193), .B(n17192), .Z(n17188) );
  ANDN U17242 ( .B(B[239]), .A(n70), .Z(n16972) );
  XNOR U17243 ( .A(n16980), .B(n17194), .Z(n16973) );
  XNOR U17244 ( .A(n16979), .B(n16977), .Z(n17194) );
  AND U17245 ( .A(n17195), .B(n17196), .Z(n16977) );
  NANDN U17246 ( .A(n17197), .B(n17198), .Z(n17196) );
  OR U17247 ( .A(n17199), .B(n17200), .Z(n17198) );
  NAND U17248 ( .A(n17200), .B(n17199), .Z(n17195) );
  ANDN U17249 ( .B(B[240]), .A(n71), .Z(n16979) );
  XNOR U17250 ( .A(n16987), .B(n17201), .Z(n16980) );
  XNOR U17251 ( .A(n16986), .B(n16984), .Z(n17201) );
  AND U17252 ( .A(n17202), .B(n17203), .Z(n16984) );
  NANDN U17253 ( .A(n17204), .B(n17205), .Z(n17203) );
  NANDN U17254 ( .A(n17206), .B(n17207), .Z(n17205) );
  NANDN U17255 ( .A(n17207), .B(n17206), .Z(n17202) );
  ANDN U17256 ( .B(B[241]), .A(n72), .Z(n16986) );
  XNOR U17257 ( .A(n16994), .B(n17208), .Z(n16987) );
  XNOR U17258 ( .A(n16993), .B(n16991), .Z(n17208) );
  AND U17259 ( .A(n17209), .B(n17210), .Z(n16991) );
  NANDN U17260 ( .A(n17211), .B(n17212), .Z(n17210) );
  OR U17261 ( .A(n17213), .B(n17214), .Z(n17212) );
  NAND U17262 ( .A(n17214), .B(n17213), .Z(n17209) );
  ANDN U17263 ( .B(B[242]), .A(n73), .Z(n16993) );
  XNOR U17264 ( .A(n17001), .B(n17215), .Z(n16994) );
  XNOR U17265 ( .A(n17000), .B(n16998), .Z(n17215) );
  AND U17266 ( .A(n17216), .B(n17217), .Z(n16998) );
  NANDN U17267 ( .A(n17218), .B(n17219), .Z(n17217) );
  NANDN U17268 ( .A(n17220), .B(n17221), .Z(n17219) );
  NANDN U17269 ( .A(n17221), .B(n17220), .Z(n17216) );
  ANDN U17270 ( .B(B[243]), .A(n74), .Z(n17000) );
  XNOR U17271 ( .A(n17008), .B(n17222), .Z(n17001) );
  XNOR U17272 ( .A(n17007), .B(n17005), .Z(n17222) );
  AND U17273 ( .A(n17223), .B(n17224), .Z(n17005) );
  NANDN U17274 ( .A(n17225), .B(n17226), .Z(n17224) );
  OR U17275 ( .A(n17227), .B(n17228), .Z(n17226) );
  NAND U17276 ( .A(n17228), .B(n17227), .Z(n17223) );
  ANDN U17277 ( .B(B[244]), .A(n75), .Z(n17007) );
  XNOR U17278 ( .A(n17015), .B(n17229), .Z(n17008) );
  XNOR U17279 ( .A(n17014), .B(n17012), .Z(n17229) );
  AND U17280 ( .A(n17230), .B(n17231), .Z(n17012) );
  NANDN U17281 ( .A(n17232), .B(n17233), .Z(n17231) );
  NANDN U17282 ( .A(n17234), .B(n17235), .Z(n17233) );
  NANDN U17283 ( .A(n17235), .B(n17234), .Z(n17230) );
  ANDN U17284 ( .B(B[245]), .A(n76), .Z(n17014) );
  XNOR U17285 ( .A(n17022), .B(n17236), .Z(n17015) );
  XNOR U17286 ( .A(n17021), .B(n17019), .Z(n17236) );
  AND U17287 ( .A(n17237), .B(n17238), .Z(n17019) );
  NANDN U17288 ( .A(n17239), .B(n17240), .Z(n17238) );
  OR U17289 ( .A(n17241), .B(n17242), .Z(n17240) );
  NAND U17290 ( .A(n17242), .B(n17241), .Z(n17237) );
  ANDN U17291 ( .B(B[246]), .A(n77), .Z(n17021) );
  XNOR U17292 ( .A(n17029), .B(n17243), .Z(n17022) );
  XNOR U17293 ( .A(n17028), .B(n17026), .Z(n17243) );
  AND U17294 ( .A(n17244), .B(n17245), .Z(n17026) );
  NANDN U17295 ( .A(n17246), .B(n17247), .Z(n17245) );
  NANDN U17296 ( .A(n17248), .B(n17249), .Z(n17247) );
  NANDN U17297 ( .A(n17249), .B(n17248), .Z(n17244) );
  ANDN U17298 ( .B(B[247]), .A(n78), .Z(n17028) );
  XNOR U17299 ( .A(n17036), .B(n17250), .Z(n17029) );
  XNOR U17300 ( .A(n17035), .B(n17033), .Z(n17250) );
  AND U17301 ( .A(n17251), .B(n17252), .Z(n17033) );
  NANDN U17302 ( .A(n17253), .B(n17254), .Z(n17252) );
  OR U17303 ( .A(n17255), .B(n17256), .Z(n17254) );
  NAND U17304 ( .A(n17256), .B(n17255), .Z(n17251) );
  ANDN U17305 ( .B(B[248]), .A(n79), .Z(n17035) );
  XNOR U17306 ( .A(n17043), .B(n17257), .Z(n17036) );
  XNOR U17307 ( .A(n17042), .B(n17040), .Z(n17257) );
  AND U17308 ( .A(n17258), .B(n17259), .Z(n17040) );
  NANDN U17309 ( .A(n17260), .B(n17261), .Z(n17259) );
  NANDN U17310 ( .A(n17262), .B(n17263), .Z(n17261) );
  NANDN U17311 ( .A(n17263), .B(n17262), .Z(n17258) );
  ANDN U17312 ( .B(B[249]), .A(n80), .Z(n17042) );
  XNOR U17313 ( .A(n17050), .B(n17264), .Z(n17043) );
  XNOR U17314 ( .A(n17049), .B(n17047), .Z(n17264) );
  AND U17315 ( .A(n17265), .B(n17266), .Z(n17047) );
  NANDN U17316 ( .A(n17267), .B(n17268), .Z(n17266) );
  OR U17317 ( .A(n17269), .B(n17270), .Z(n17268) );
  NAND U17318 ( .A(n17270), .B(n17269), .Z(n17265) );
  ANDN U17319 ( .B(B[250]), .A(n81), .Z(n17049) );
  XNOR U17320 ( .A(n17057), .B(n17271), .Z(n17050) );
  XNOR U17321 ( .A(n17056), .B(n17054), .Z(n17271) );
  AND U17322 ( .A(n17272), .B(n17273), .Z(n17054) );
  NANDN U17323 ( .A(n17274), .B(n17275), .Z(n17273) );
  NAND U17324 ( .A(n17276), .B(n17277), .Z(n17275) );
  ANDN U17325 ( .B(B[251]), .A(n82), .Z(n17056) );
  XOR U17326 ( .A(n17063), .B(n17278), .Z(n17057) );
  XNOR U17327 ( .A(n17061), .B(n17064), .Z(n17278) );
  NAND U17328 ( .A(A[2]), .B(B[252]), .Z(n17064) );
  NANDN U17329 ( .A(n17279), .B(n17280), .Z(n17061) );
  AND U17330 ( .A(A[0]), .B(B[253]), .Z(n17280) );
  XNOR U17331 ( .A(n17066), .B(n17281), .Z(n17063) );
  NAND U17332 ( .A(A[0]), .B(B[254]), .Z(n17281) );
  NAND U17333 ( .A(B[253]), .B(A[1]), .Z(n17066) );
  NAND U17334 ( .A(n17282), .B(n17283), .Z(n288) );
  NANDN U17335 ( .A(n17284), .B(n17285), .Z(n17283) );
  OR U17336 ( .A(n17286), .B(n17287), .Z(n17285) );
  NAND U17337 ( .A(n17287), .B(n17286), .Z(n17282) );
  XOR U17338 ( .A(n290), .B(n289), .Z(\A1[251] ) );
  XOR U17339 ( .A(n17287), .B(n17288), .Z(n289) );
  XNOR U17340 ( .A(n17286), .B(n17284), .Z(n17288) );
  AND U17341 ( .A(n17289), .B(n17290), .Z(n17284) );
  NANDN U17342 ( .A(n17291), .B(n17292), .Z(n17290) );
  NANDN U17343 ( .A(n17293), .B(n17294), .Z(n17292) );
  NANDN U17344 ( .A(n17294), .B(n17293), .Z(n17289) );
  ANDN U17345 ( .B(B[222]), .A(n54), .Z(n17286) );
  XNOR U17346 ( .A(n17081), .B(n17295), .Z(n17287) );
  XNOR U17347 ( .A(n17080), .B(n17078), .Z(n17295) );
  AND U17348 ( .A(n17296), .B(n17297), .Z(n17078) );
  NANDN U17349 ( .A(n17298), .B(n17299), .Z(n17297) );
  OR U17350 ( .A(n17300), .B(n17301), .Z(n17299) );
  NAND U17351 ( .A(n17301), .B(n17300), .Z(n17296) );
  ANDN U17352 ( .B(B[223]), .A(n55), .Z(n17080) );
  XNOR U17353 ( .A(n17088), .B(n17302), .Z(n17081) );
  XNOR U17354 ( .A(n17087), .B(n17085), .Z(n17302) );
  AND U17355 ( .A(n17303), .B(n17304), .Z(n17085) );
  NANDN U17356 ( .A(n17305), .B(n17306), .Z(n17304) );
  NANDN U17357 ( .A(n17307), .B(n17308), .Z(n17306) );
  NANDN U17358 ( .A(n17308), .B(n17307), .Z(n17303) );
  ANDN U17359 ( .B(B[224]), .A(n56), .Z(n17087) );
  XNOR U17360 ( .A(n17095), .B(n17309), .Z(n17088) );
  XNOR U17361 ( .A(n17094), .B(n17092), .Z(n17309) );
  AND U17362 ( .A(n17310), .B(n17311), .Z(n17092) );
  NANDN U17363 ( .A(n17312), .B(n17313), .Z(n17311) );
  OR U17364 ( .A(n17314), .B(n17315), .Z(n17313) );
  NAND U17365 ( .A(n17315), .B(n17314), .Z(n17310) );
  ANDN U17366 ( .B(B[225]), .A(n57), .Z(n17094) );
  XNOR U17367 ( .A(n17102), .B(n17316), .Z(n17095) );
  XNOR U17368 ( .A(n17101), .B(n17099), .Z(n17316) );
  AND U17369 ( .A(n17317), .B(n17318), .Z(n17099) );
  NANDN U17370 ( .A(n17319), .B(n17320), .Z(n17318) );
  NANDN U17371 ( .A(n17321), .B(n17322), .Z(n17320) );
  NANDN U17372 ( .A(n17322), .B(n17321), .Z(n17317) );
  ANDN U17373 ( .B(B[226]), .A(n58), .Z(n17101) );
  XNOR U17374 ( .A(n17109), .B(n17323), .Z(n17102) );
  XNOR U17375 ( .A(n17108), .B(n17106), .Z(n17323) );
  AND U17376 ( .A(n17324), .B(n17325), .Z(n17106) );
  NANDN U17377 ( .A(n17326), .B(n17327), .Z(n17325) );
  OR U17378 ( .A(n17328), .B(n17329), .Z(n17327) );
  NAND U17379 ( .A(n17329), .B(n17328), .Z(n17324) );
  ANDN U17380 ( .B(B[227]), .A(n59), .Z(n17108) );
  XNOR U17381 ( .A(n17116), .B(n17330), .Z(n17109) );
  XNOR U17382 ( .A(n17115), .B(n17113), .Z(n17330) );
  AND U17383 ( .A(n17331), .B(n17332), .Z(n17113) );
  NANDN U17384 ( .A(n17333), .B(n17334), .Z(n17332) );
  NANDN U17385 ( .A(n17335), .B(n17336), .Z(n17334) );
  NANDN U17386 ( .A(n17336), .B(n17335), .Z(n17331) );
  ANDN U17387 ( .B(B[228]), .A(n60), .Z(n17115) );
  XNOR U17388 ( .A(n17123), .B(n17337), .Z(n17116) );
  XNOR U17389 ( .A(n17122), .B(n17120), .Z(n17337) );
  AND U17390 ( .A(n17338), .B(n17339), .Z(n17120) );
  NANDN U17391 ( .A(n17340), .B(n17341), .Z(n17339) );
  OR U17392 ( .A(n17342), .B(n17343), .Z(n17341) );
  NAND U17393 ( .A(n17343), .B(n17342), .Z(n17338) );
  ANDN U17394 ( .B(B[229]), .A(n61), .Z(n17122) );
  XNOR U17395 ( .A(n17130), .B(n17344), .Z(n17123) );
  XNOR U17396 ( .A(n17129), .B(n17127), .Z(n17344) );
  AND U17397 ( .A(n17345), .B(n17346), .Z(n17127) );
  NANDN U17398 ( .A(n17347), .B(n17348), .Z(n17346) );
  NANDN U17399 ( .A(n17349), .B(n17350), .Z(n17348) );
  NANDN U17400 ( .A(n17350), .B(n17349), .Z(n17345) );
  ANDN U17401 ( .B(B[230]), .A(n62), .Z(n17129) );
  XNOR U17402 ( .A(n17137), .B(n17351), .Z(n17130) );
  XNOR U17403 ( .A(n17136), .B(n17134), .Z(n17351) );
  AND U17404 ( .A(n17352), .B(n17353), .Z(n17134) );
  NANDN U17405 ( .A(n17354), .B(n17355), .Z(n17353) );
  OR U17406 ( .A(n17356), .B(n17357), .Z(n17355) );
  NAND U17407 ( .A(n17357), .B(n17356), .Z(n17352) );
  ANDN U17408 ( .B(B[231]), .A(n63), .Z(n17136) );
  XNOR U17409 ( .A(n17144), .B(n17358), .Z(n17137) );
  XNOR U17410 ( .A(n17143), .B(n17141), .Z(n17358) );
  AND U17411 ( .A(n17359), .B(n17360), .Z(n17141) );
  NANDN U17412 ( .A(n17361), .B(n17362), .Z(n17360) );
  NANDN U17413 ( .A(n17363), .B(n17364), .Z(n17362) );
  NANDN U17414 ( .A(n17364), .B(n17363), .Z(n17359) );
  ANDN U17415 ( .B(B[232]), .A(n64), .Z(n17143) );
  XNOR U17416 ( .A(n17151), .B(n17365), .Z(n17144) );
  XNOR U17417 ( .A(n17150), .B(n17148), .Z(n17365) );
  AND U17418 ( .A(n17366), .B(n17367), .Z(n17148) );
  NANDN U17419 ( .A(n17368), .B(n17369), .Z(n17367) );
  OR U17420 ( .A(n17370), .B(n17371), .Z(n17369) );
  NAND U17421 ( .A(n17371), .B(n17370), .Z(n17366) );
  ANDN U17422 ( .B(B[233]), .A(n65), .Z(n17150) );
  XNOR U17423 ( .A(n17158), .B(n17372), .Z(n17151) );
  XNOR U17424 ( .A(n17157), .B(n17155), .Z(n17372) );
  AND U17425 ( .A(n17373), .B(n17374), .Z(n17155) );
  NANDN U17426 ( .A(n17375), .B(n17376), .Z(n17374) );
  NANDN U17427 ( .A(n17377), .B(n17378), .Z(n17376) );
  NANDN U17428 ( .A(n17378), .B(n17377), .Z(n17373) );
  ANDN U17429 ( .B(B[234]), .A(n66), .Z(n17157) );
  XNOR U17430 ( .A(n17165), .B(n17379), .Z(n17158) );
  XNOR U17431 ( .A(n17164), .B(n17162), .Z(n17379) );
  AND U17432 ( .A(n17380), .B(n17381), .Z(n17162) );
  NANDN U17433 ( .A(n17382), .B(n17383), .Z(n17381) );
  OR U17434 ( .A(n17384), .B(n17385), .Z(n17383) );
  NAND U17435 ( .A(n17385), .B(n17384), .Z(n17380) );
  ANDN U17436 ( .B(B[235]), .A(n67), .Z(n17164) );
  XNOR U17437 ( .A(n17172), .B(n17386), .Z(n17165) );
  XNOR U17438 ( .A(n17171), .B(n17169), .Z(n17386) );
  AND U17439 ( .A(n17387), .B(n17388), .Z(n17169) );
  NANDN U17440 ( .A(n17389), .B(n17390), .Z(n17388) );
  NANDN U17441 ( .A(n17391), .B(n17392), .Z(n17390) );
  NANDN U17442 ( .A(n17392), .B(n17391), .Z(n17387) );
  ANDN U17443 ( .B(B[236]), .A(n68), .Z(n17171) );
  XNOR U17444 ( .A(n17179), .B(n17393), .Z(n17172) );
  XNOR U17445 ( .A(n17178), .B(n17176), .Z(n17393) );
  AND U17446 ( .A(n17394), .B(n17395), .Z(n17176) );
  NANDN U17447 ( .A(n17396), .B(n17397), .Z(n17395) );
  OR U17448 ( .A(n17398), .B(n17399), .Z(n17397) );
  NAND U17449 ( .A(n17399), .B(n17398), .Z(n17394) );
  ANDN U17450 ( .B(B[237]), .A(n69), .Z(n17178) );
  XNOR U17451 ( .A(n17186), .B(n17400), .Z(n17179) );
  XNOR U17452 ( .A(n17185), .B(n17183), .Z(n17400) );
  AND U17453 ( .A(n17401), .B(n17402), .Z(n17183) );
  NANDN U17454 ( .A(n17403), .B(n17404), .Z(n17402) );
  NANDN U17455 ( .A(n17405), .B(n17406), .Z(n17404) );
  NANDN U17456 ( .A(n17406), .B(n17405), .Z(n17401) );
  ANDN U17457 ( .B(B[238]), .A(n70), .Z(n17185) );
  XNOR U17458 ( .A(n17193), .B(n17407), .Z(n17186) );
  XNOR U17459 ( .A(n17192), .B(n17190), .Z(n17407) );
  AND U17460 ( .A(n17408), .B(n17409), .Z(n17190) );
  NANDN U17461 ( .A(n17410), .B(n17411), .Z(n17409) );
  OR U17462 ( .A(n17412), .B(n17413), .Z(n17411) );
  NAND U17463 ( .A(n17413), .B(n17412), .Z(n17408) );
  ANDN U17464 ( .B(B[239]), .A(n71), .Z(n17192) );
  XNOR U17465 ( .A(n17200), .B(n17414), .Z(n17193) );
  XNOR U17466 ( .A(n17199), .B(n17197), .Z(n17414) );
  AND U17467 ( .A(n17415), .B(n17416), .Z(n17197) );
  NANDN U17468 ( .A(n17417), .B(n17418), .Z(n17416) );
  NANDN U17469 ( .A(n17419), .B(n17420), .Z(n17418) );
  NANDN U17470 ( .A(n17420), .B(n17419), .Z(n17415) );
  ANDN U17471 ( .B(B[240]), .A(n72), .Z(n17199) );
  XNOR U17472 ( .A(n17207), .B(n17421), .Z(n17200) );
  XNOR U17473 ( .A(n17206), .B(n17204), .Z(n17421) );
  AND U17474 ( .A(n17422), .B(n17423), .Z(n17204) );
  NANDN U17475 ( .A(n17424), .B(n17425), .Z(n17423) );
  OR U17476 ( .A(n17426), .B(n17427), .Z(n17425) );
  NAND U17477 ( .A(n17427), .B(n17426), .Z(n17422) );
  ANDN U17478 ( .B(B[241]), .A(n73), .Z(n17206) );
  XNOR U17479 ( .A(n17214), .B(n17428), .Z(n17207) );
  XNOR U17480 ( .A(n17213), .B(n17211), .Z(n17428) );
  AND U17481 ( .A(n17429), .B(n17430), .Z(n17211) );
  NANDN U17482 ( .A(n17431), .B(n17432), .Z(n17430) );
  NANDN U17483 ( .A(n17433), .B(n17434), .Z(n17432) );
  NANDN U17484 ( .A(n17434), .B(n17433), .Z(n17429) );
  ANDN U17485 ( .B(B[242]), .A(n74), .Z(n17213) );
  XNOR U17486 ( .A(n17221), .B(n17435), .Z(n17214) );
  XNOR U17487 ( .A(n17220), .B(n17218), .Z(n17435) );
  AND U17488 ( .A(n17436), .B(n17437), .Z(n17218) );
  NANDN U17489 ( .A(n17438), .B(n17439), .Z(n17437) );
  OR U17490 ( .A(n17440), .B(n17441), .Z(n17439) );
  NAND U17491 ( .A(n17441), .B(n17440), .Z(n17436) );
  ANDN U17492 ( .B(B[243]), .A(n75), .Z(n17220) );
  XNOR U17493 ( .A(n17228), .B(n17442), .Z(n17221) );
  XNOR U17494 ( .A(n17227), .B(n17225), .Z(n17442) );
  AND U17495 ( .A(n17443), .B(n17444), .Z(n17225) );
  NANDN U17496 ( .A(n17445), .B(n17446), .Z(n17444) );
  NANDN U17497 ( .A(n17447), .B(n17448), .Z(n17446) );
  NANDN U17498 ( .A(n17448), .B(n17447), .Z(n17443) );
  ANDN U17499 ( .B(B[244]), .A(n76), .Z(n17227) );
  XNOR U17500 ( .A(n17235), .B(n17449), .Z(n17228) );
  XNOR U17501 ( .A(n17234), .B(n17232), .Z(n17449) );
  AND U17502 ( .A(n17450), .B(n17451), .Z(n17232) );
  NANDN U17503 ( .A(n17452), .B(n17453), .Z(n17451) );
  OR U17504 ( .A(n17454), .B(n17455), .Z(n17453) );
  NAND U17505 ( .A(n17455), .B(n17454), .Z(n17450) );
  ANDN U17506 ( .B(B[245]), .A(n77), .Z(n17234) );
  XNOR U17507 ( .A(n17242), .B(n17456), .Z(n17235) );
  XNOR U17508 ( .A(n17241), .B(n17239), .Z(n17456) );
  AND U17509 ( .A(n17457), .B(n17458), .Z(n17239) );
  NANDN U17510 ( .A(n17459), .B(n17460), .Z(n17458) );
  NANDN U17511 ( .A(n17461), .B(n17462), .Z(n17460) );
  NANDN U17512 ( .A(n17462), .B(n17461), .Z(n17457) );
  ANDN U17513 ( .B(B[246]), .A(n78), .Z(n17241) );
  XNOR U17514 ( .A(n17249), .B(n17463), .Z(n17242) );
  XNOR U17515 ( .A(n17248), .B(n17246), .Z(n17463) );
  AND U17516 ( .A(n17464), .B(n17465), .Z(n17246) );
  NANDN U17517 ( .A(n17466), .B(n17467), .Z(n17465) );
  OR U17518 ( .A(n17468), .B(n17469), .Z(n17467) );
  NAND U17519 ( .A(n17469), .B(n17468), .Z(n17464) );
  ANDN U17520 ( .B(B[247]), .A(n79), .Z(n17248) );
  XNOR U17521 ( .A(n17256), .B(n17470), .Z(n17249) );
  XNOR U17522 ( .A(n17255), .B(n17253), .Z(n17470) );
  AND U17523 ( .A(n17471), .B(n17472), .Z(n17253) );
  NANDN U17524 ( .A(n17473), .B(n17474), .Z(n17472) );
  NANDN U17525 ( .A(n17475), .B(n17476), .Z(n17474) );
  NANDN U17526 ( .A(n17476), .B(n17475), .Z(n17471) );
  ANDN U17527 ( .B(B[248]), .A(n80), .Z(n17255) );
  XNOR U17528 ( .A(n17263), .B(n17477), .Z(n17256) );
  XNOR U17529 ( .A(n17262), .B(n17260), .Z(n17477) );
  AND U17530 ( .A(n17478), .B(n17479), .Z(n17260) );
  NANDN U17531 ( .A(n17480), .B(n17481), .Z(n17479) );
  OR U17532 ( .A(n17482), .B(n17483), .Z(n17481) );
  NAND U17533 ( .A(n17483), .B(n17482), .Z(n17478) );
  ANDN U17534 ( .B(B[249]), .A(n81), .Z(n17262) );
  XNOR U17535 ( .A(n17270), .B(n17484), .Z(n17263) );
  XNOR U17536 ( .A(n17269), .B(n17267), .Z(n17484) );
  AND U17537 ( .A(n17485), .B(n17486), .Z(n17267) );
  NANDN U17538 ( .A(n17487), .B(n17488), .Z(n17486) );
  NAND U17539 ( .A(n17489), .B(n17490), .Z(n17488) );
  ANDN U17540 ( .B(B[250]), .A(n82), .Z(n17269) );
  XOR U17541 ( .A(n17276), .B(n17491), .Z(n17270) );
  XNOR U17542 ( .A(n17274), .B(n17277), .Z(n17491) );
  NAND U17543 ( .A(A[2]), .B(B[251]), .Z(n17277) );
  NANDN U17544 ( .A(n17492), .B(n17493), .Z(n17274) );
  AND U17545 ( .A(A[0]), .B(B[252]), .Z(n17493) );
  XNOR U17546 ( .A(n17279), .B(n17494), .Z(n17276) );
  NAND U17547 ( .A(A[0]), .B(B[253]), .Z(n17494) );
  NAND U17548 ( .A(B[252]), .B(A[1]), .Z(n17279) );
  NAND U17549 ( .A(n17495), .B(n17496), .Z(n290) );
  NANDN U17550 ( .A(n17497), .B(n17498), .Z(n17496) );
  OR U17551 ( .A(n17499), .B(n17500), .Z(n17498) );
  NAND U17552 ( .A(n17500), .B(n17499), .Z(n17495) );
  XOR U17553 ( .A(n292), .B(n291), .Z(\A1[250] ) );
  XOR U17554 ( .A(n17500), .B(n17501), .Z(n291) );
  XNOR U17555 ( .A(n17499), .B(n17497), .Z(n17501) );
  AND U17556 ( .A(n17502), .B(n17503), .Z(n17497) );
  NANDN U17557 ( .A(n17504), .B(n17505), .Z(n17503) );
  NANDN U17558 ( .A(n17506), .B(n17507), .Z(n17505) );
  NANDN U17559 ( .A(n17507), .B(n17506), .Z(n17502) );
  ANDN U17560 ( .B(B[221]), .A(n54), .Z(n17499) );
  XNOR U17561 ( .A(n17294), .B(n17508), .Z(n17500) );
  XNOR U17562 ( .A(n17293), .B(n17291), .Z(n17508) );
  AND U17563 ( .A(n17509), .B(n17510), .Z(n17291) );
  NANDN U17564 ( .A(n17511), .B(n17512), .Z(n17510) );
  OR U17565 ( .A(n17513), .B(n17514), .Z(n17512) );
  NAND U17566 ( .A(n17514), .B(n17513), .Z(n17509) );
  ANDN U17567 ( .B(B[222]), .A(n55), .Z(n17293) );
  XNOR U17568 ( .A(n17301), .B(n17515), .Z(n17294) );
  XNOR U17569 ( .A(n17300), .B(n17298), .Z(n17515) );
  AND U17570 ( .A(n17516), .B(n17517), .Z(n17298) );
  NANDN U17571 ( .A(n17518), .B(n17519), .Z(n17517) );
  NANDN U17572 ( .A(n17520), .B(n17521), .Z(n17519) );
  NANDN U17573 ( .A(n17521), .B(n17520), .Z(n17516) );
  ANDN U17574 ( .B(B[223]), .A(n56), .Z(n17300) );
  XNOR U17575 ( .A(n17308), .B(n17522), .Z(n17301) );
  XNOR U17576 ( .A(n17307), .B(n17305), .Z(n17522) );
  AND U17577 ( .A(n17523), .B(n17524), .Z(n17305) );
  NANDN U17578 ( .A(n17525), .B(n17526), .Z(n17524) );
  OR U17579 ( .A(n17527), .B(n17528), .Z(n17526) );
  NAND U17580 ( .A(n17528), .B(n17527), .Z(n17523) );
  ANDN U17581 ( .B(B[224]), .A(n57), .Z(n17307) );
  XNOR U17582 ( .A(n17315), .B(n17529), .Z(n17308) );
  XNOR U17583 ( .A(n17314), .B(n17312), .Z(n17529) );
  AND U17584 ( .A(n17530), .B(n17531), .Z(n17312) );
  NANDN U17585 ( .A(n17532), .B(n17533), .Z(n17531) );
  NANDN U17586 ( .A(n17534), .B(n17535), .Z(n17533) );
  NANDN U17587 ( .A(n17535), .B(n17534), .Z(n17530) );
  ANDN U17588 ( .B(B[225]), .A(n58), .Z(n17314) );
  XNOR U17589 ( .A(n17322), .B(n17536), .Z(n17315) );
  XNOR U17590 ( .A(n17321), .B(n17319), .Z(n17536) );
  AND U17591 ( .A(n17537), .B(n17538), .Z(n17319) );
  NANDN U17592 ( .A(n17539), .B(n17540), .Z(n17538) );
  OR U17593 ( .A(n17541), .B(n17542), .Z(n17540) );
  NAND U17594 ( .A(n17542), .B(n17541), .Z(n17537) );
  ANDN U17595 ( .B(B[226]), .A(n59), .Z(n17321) );
  XNOR U17596 ( .A(n17329), .B(n17543), .Z(n17322) );
  XNOR U17597 ( .A(n17328), .B(n17326), .Z(n17543) );
  AND U17598 ( .A(n17544), .B(n17545), .Z(n17326) );
  NANDN U17599 ( .A(n17546), .B(n17547), .Z(n17545) );
  NANDN U17600 ( .A(n17548), .B(n17549), .Z(n17547) );
  NANDN U17601 ( .A(n17549), .B(n17548), .Z(n17544) );
  ANDN U17602 ( .B(B[227]), .A(n60), .Z(n17328) );
  XNOR U17603 ( .A(n17336), .B(n17550), .Z(n17329) );
  XNOR U17604 ( .A(n17335), .B(n17333), .Z(n17550) );
  AND U17605 ( .A(n17551), .B(n17552), .Z(n17333) );
  NANDN U17606 ( .A(n17553), .B(n17554), .Z(n17552) );
  OR U17607 ( .A(n17555), .B(n17556), .Z(n17554) );
  NAND U17608 ( .A(n17556), .B(n17555), .Z(n17551) );
  ANDN U17609 ( .B(B[228]), .A(n61), .Z(n17335) );
  XNOR U17610 ( .A(n17343), .B(n17557), .Z(n17336) );
  XNOR U17611 ( .A(n17342), .B(n17340), .Z(n17557) );
  AND U17612 ( .A(n17558), .B(n17559), .Z(n17340) );
  NANDN U17613 ( .A(n17560), .B(n17561), .Z(n17559) );
  NANDN U17614 ( .A(n17562), .B(n17563), .Z(n17561) );
  NANDN U17615 ( .A(n17563), .B(n17562), .Z(n17558) );
  ANDN U17616 ( .B(B[229]), .A(n62), .Z(n17342) );
  XNOR U17617 ( .A(n17350), .B(n17564), .Z(n17343) );
  XNOR U17618 ( .A(n17349), .B(n17347), .Z(n17564) );
  AND U17619 ( .A(n17565), .B(n17566), .Z(n17347) );
  NANDN U17620 ( .A(n17567), .B(n17568), .Z(n17566) );
  OR U17621 ( .A(n17569), .B(n17570), .Z(n17568) );
  NAND U17622 ( .A(n17570), .B(n17569), .Z(n17565) );
  ANDN U17623 ( .B(B[230]), .A(n63), .Z(n17349) );
  XNOR U17624 ( .A(n17357), .B(n17571), .Z(n17350) );
  XNOR U17625 ( .A(n17356), .B(n17354), .Z(n17571) );
  AND U17626 ( .A(n17572), .B(n17573), .Z(n17354) );
  NANDN U17627 ( .A(n17574), .B(n17575), .Z(n17573) );
  NANDN U17628 ( .A(n17576), .B(n17577), .Z(n17575) );
  NANDN U17629 ( .A(n17577), .B(n17576), .Z(n17572) );
  ANDN U17630 ( .B(B[231]), .A(n64), .Z(n17356) );
  XNOR U17631 ( .A(n17364), .B(n17578), .Z(n17357) );
  XNOR U17632 ( .A(n17363), .B(n17361), .Z(n17578) );
  AND U17633 ( .A(n17579), .B(n17580), .Z(n17361) );
  NANDN U17634 ( .A(n17581), .B(n17582), .Z(n17580) );
  OR U17635 ( .A(n17583), .B(n17584), .Z(n17582) );
  NAND U17636 ( .A(n17584), .B(n17583), .Z(n17579) );
  ANDN U17637 ( .B(B[232]), .A(n65), .Z(n17363) );
  XNOR U17638 ( .A(n17371), .B(n17585), .Z(n17364) );
  XNOR U17639 ( .A(n17370), .B(n17368), .Z(n17585) );
  AND U17640 ( .A(n17586), .B(n17587), .Z(n17368) );
  NANDN U17641 ( .A(n17588), .B(n17589), .Z(n17587) );
  NANDN U17642 ( .A(n17590), .B(n17591), .Z(n17589) );
  NANDN U17643 ( .A(n17591), .B(n17590), .Z(n17586) );
  ANDN U17644 ( .B(B[233]), .A(n66), .Z(n17370) );
  XNOR U17645 ( .A(n17378), .B(n17592), .Z(n17371) );
  XNOR U17646 ( .A(n17377), .B(n17375), .Z(n17592) );
  AND U17647 ( .A(n17593), .B(n17594), .Z(n17375) );
  NANDN U17648 ( .A(n17595), .B(n17596), .Z(n17594) );
  OR U17649 ( .A(n17597), .B(n17598), .Z(n17596) );
  NAND U17650 ( .A(n17598), .B(n17597), .Z(n17593) );
  ANDN U17651 ( .B(B[234]), .A(n67), .Z(n17377) );
  XNOR U17652 ( .A(n17385), .B(n17599), .Z(n17378) );
  XNOR U17653 ( .A(n17384), .B(n17382), .Z(n17599) );
  AND U17654 ( .A(n17600), .B(n17601), .Z(n17382) );
  NANDN U17655 ( .A(n17602), .B(n17603), .Z(n17601) );
  NANDN U17656 ( .A(n17604), .B(n17605), .Z(n17603) );
  NANDN U17657 ( .A(n17605), .B(n17604), .Z(n17600) );
  ANDN U17658 ( .B(B[235]), .A(n68), .Z(n17384) );
  XNOR U17659 ( .A(n17392), .B(n17606), .Z(n17385) );
  XNOR U17660 ( .A(n17391), .B(n17389), .Z(n17606) );
  AND U17661 ( .A(n17607), .B(n17608), .Z(n17389) );
  NANDN U17662 ( .A(n17609), .B(n17610), .Z(n17608) );
  OR U17663 ( .A(n17611), .B(n17612), .Z(n17610) );
  NAND U17664 ( .A(n17612), .B(n17611), .Z(n17607) );
  ANDN U17665 ( .B(B[236]), .A(n69), .Z(n17391) );
  XNOR U17666 ( .A(n17399), .B(n17613), .Z(n17392) );
  XNOR U17667 ( .A(n17398), .B(n17396), .Z(n17613) );
  AND U17668 ( .A(n17614), .B(n17615), .Z(n17396) );
  NANDN U17669 ( .A(n17616), .B(n17617), .Z(n17615) );
  NANDN U17670 ( .A(n17618), .B(n17619), .Z(n17617) );
  NANDN U17671 ( .A(n17619), .B(n17618), .Z(n17614) );
  ANDN U17672 ( .B(B[237]), .A(n70), .Z(n17398) );
  XNOR U17673 ( .A(n17406), .B(n17620), .Z(n17399) );
  XNOR U17674 ( .A(n17405), .B(n17403), .Z(n17620) );
  AND U17675 ( .A(n17621), .B(n17622), .Z(n17403) );
  NANDN U17676 ( .A(n17623), .B(n17624), .Z(n17622) );
  OR U17677 ( .A(n17625), .B(n17626), .Z(n17624) );
  NAND U17678 ( .A(n17626), .B(n17625), .Z(n17621) );
  ANDN U17679 ( .B(B[238]), .A(n71), .Z(n17405) );
  XNOR U17680 ( .A(n17413), .B(n17627), .Z(n17406) );
  XNOR U17681 ( .A(n17412), .B(n17410), .Z(n17627) );
  AND U17682 ( .A(n17628), .B(n17629), .Z(n17410) );
  NANDN U17683 ( .A(n17630), .B(n17631), .Z(n17629) );
  NANDN U17684 ( .A(n17632), .B(n17633), .Z(n17631) );
  NANDN U17685 ( .A(n17633), .B(n17632), .Z(n17628) );
  ANDN U17686 ( .B(B[239]), .A(n72), .Z(n17412) );
  XNOR U17687 ( .A(n17420), .B(n17634), .Z(n17413) );
  XNOR U17688 ( .A(n17419), .B(n17417), .Z(n17634) );
  AND U17689 ( .A(n17635), .B(n17636), .Z(n17417) );
  NANDN U17690 ( .A(n17637), .B(n17638), .Z(n17636) );
  OR U17691 ( .A(n17639), .B(n17640), .Z(n17638) );
  NAND U17692 ( .A(n17640), .B(n17639), .Z(n17635) );
  ANDN U17693 ( .B(B[240]), .A(n73), .Z(n17419) );
  XNOR U17694 ( .A(n17427), .B(n17641), .Z(n17420) );
  XNOR U17695 ( .A(n17426), .B(n17424), .Z(n17641) );
  AND U17696 ( .A(n17642), .B(n17643), .Z(n17424) );
  NANDN U17697 ( .A(n17644), .B(n17645), .Z(n17643) );
  NANDN U17698 ( .A(n17646), .B(n17647), .Z(n17645) );
  NANDN U17699 ( .A(n17647), .B(n17646), .Z(n17642) );
  ANDN U17700 ( .B(B[241]), .A(n74), .Z(n17426) );
  XNOR U17701 ( .A(n17434), .B(n17648), .Z(n17427) );
  XNOR U17702 ( .A(n17433), .B(n17431), .Z(n17648) );
  AND U17703 ( .A(n17649), .B(n17650), .Z(n17431) );
  NANDN U17704 ( .A(n17651), .B(n17652), .Z(n17650) );
  OR U17705 ( .A(n17653), .B(n17654), .Z(n17652) );
  NAND U17706 ( .A(n17654), .B(n17653), .Z(n17649) );
  ANDN U17707 ( .B(B[242]), .A(n75), .Z(n17433) );
  XNOR U17708 ( .A(n17441), .B(n17655), .Z(n17434) );
  XNOR U17709 ( .A(n17440), .B(n17438), .Z(n17655) );
  AND U17710 ( .A(n17656), .B(n17657), .Z(n17438) );
  NANDN U17711 ( .A(n17658), .B(n17659), .Z(n17657) );
  NANDN U17712 ( .A(n17660), .B(n17661), .Z(n17659) );
  NANDN U17713 ( .A(n17661), .B(n17660), .Z(n17656) );
  ANDN U17714 ( .B(B[243]), .A(n76), .Z(n17440) );
  XNOR U17715 ( .A(n17448), .B(n17662), .Z(n17441) );
  XNOR U17716 ( .A(n17447), .B(n17445), .Z(n17662) );
  AND U17717 ( .A(n17663), .B(n17664), .Z(n17445) );
  NANDN U17718 ( .A(n17665), .B(n17666), .Z(n17664) );
  OR U17719 ( .A(n17667), .B(n17668), .Z(n17666) );
  NAND U17720 ( .A(n17668), .B(n17667), .Z(n17663) );
  ANDN U17721 ( .B(B[244]), .A(n77), .Z(n17447) );
  XNOR U17722 ( .A(n17455), .B(n17669), .Z(n17448) );
  XNOR U17723 ( .A(n17454), .B(n17452), .Z(n17669) );
  AND U17724 ( .A(n17670), .B(n17671), .Z(n17452) );
  NANDN U17725 ( .A(n17672), .B(n17673), .Z(n17671) );
  NANDN U17726 ( .A(n17674), .B(n17675), .Z(n17673) );
  NANDN U17727 ( .A(n17675), .B(n17674), .Z(n17670) );
  ANDN U17728 ( .B(B[245]), .A(n78), .Z(n17454) );
  XNOR U17729 ( .A(n17462), .B(n17676), .Z(n17455) );
  XNOR U17730 ( .A(n17461), .B(n17459), .Z(n17676) );
  AND U17731 ( .A(n17677), .B(n17678), .Z(n17459) );
  NANDN U17732 ( .A(n17679), .B(n17680), .Z(n17678) );
  OR U17733 ( .A(n17681), .B(n17682), .Z(n17680) );
  NAND U17734 ( .A(n17682), .B(n17681), .Z(n17677) );
  ANDN U17735 ( .B(B[246]), .A(n79), .Z(n17461) );
  XNOR U17736 ( .A(n17469), .B(n17683), .Z(n17462) );
  XNOR U17737 ( .A(n17468), .B(n17466), .Z(n17683) );
  AND U17738 ( .A(n17684), .B(n17685), .Z(n17466) );
  NANDN U17739 ( .A(n17686), .B(n17687), .Z(n17685) );
  NANDN U17740 ( .A(n17688), .B(n17689), .Z(n17687) );
  NANDN U17741 ( .A(n17689), .B(n17688), .Z(n17684) );
  ANDN U17742 ( .B(B[247]), .A(n80), .Z(n17468) );
  XNOR U17743 ( .A(n17476), .B(n17690), .Z(n17469) );
  XNOR U17744 ( .A(n17475), .B(n17473), .Z(n17690) );
  AND U17745 ( .A(n17691), .B(n17692), .Z(n17473) );
  NANDN U17746 ( .A(n17693), .B(n17694), .Z(n17692) );
  OR U17747 ( .A(n17695), .B(n17696), .Z(n17694) );
  NAND U17748 ( .A(n17696), .B(n17695), .Z(n17691) );
  ANDN U17749 ( .B(B[248]), .A(n81), .Z(n17475) );
  XNOR U17750 ( .A(n17483), .B(n17697), .Z(n17476) );
  XNOR U17751 ( .A(n17482), .B(n17480), .Z(n17697) );
  AND U17752 ( .A(n17698), .B(n17699), .Z(n17480) );
  NANDN U17753 ( .A(n17700), .B(n17701), .Z(n17699) );
  NAND U17754 ( .A(n17702), .B(n17703), .Z(n17701) );
  ANDN U17755 ( .B(B[249]), .A(n82), .Z(n17482) );
  XOR U17756 ( .A(n17489), .B(n17704), .Z(n17483) );
  XNOR U17757 ( .A(n17487), .B(n17490), .Z(n17704) );
  NAND U17758 ( .A(A[2]), .B(B[250]), .Z(n17490) );
  NANDN U17759 ( .A(n17705), .B(n17706), .Z(n17487) );
  AND U17760 ( .A(A[0]), .B(B[251]), .Z(n17706) );
  XNOR U17761 ( .A(n17492), .B(n17707), .Z(n17489) );
  NAND U17762 ( .A(A[0]), .B(B[252]), .Z(n17707) );
  NAND U17763 ( .A(B[251]), .B(A[1]), .Z(n17492) );
  NAND U17764 ( .A(n17708), .B(n17709), .Z(n292) );
  NANDN U17765 ( .A(n17710), .B(n17711), .Z(n17709) );
  OR U17766 ( .A(n17712), .B(n17713), .Z(n17711) );
  NAND U17767 ( .A(n17713), .B(n17712), .Z(n17708) );
  XOR U17768 ( .A(n15504), .B(n17714), .Z(\A1[24] ) );
  XNOR U17769 ( .A(n15503), .B(n15502), .Z(n17714) );
  NAND U17770 ( .A(n17715), .B(n17716), .Z(n15502) );
  NANDN U17771 ( .A(n17717), .B(n17718), .Z(n17716) );
  OR U17772 ( .A(n17719), .B(n17720), .Z(n17718) );
  NAND U17773 ( .A(n17720), .B(n17719), .Z(n17715) );
  ANDN U17774 ( .B(B[0]), .A(n59), .Z(n15503) );
  XNOR U17775 ( .A(n15511), .B(n17721), .Z(n15504) );
  XNOR U17776 ( .A(n15510), .B(n15508), .Z(n17721) );
  AND U17777 ( .A(n17722), .B(n17723), .Z(n15508) );
  NANDN U17778 ( .A(n17724), .B(n17725), .Z(n17723) );
  NANDN U17779 ( .A(n17726), .B(n17727), .Z(n17725) );
  NANDN U17780 ( .A(n17727), .B(n17726), .Z(n17722) );
  ANDN U17781 ( .B(B[1]), .A(n60), .Z(n15510) );
  XNOR U17782 ( .A(n15518), .B(n17728), .Z(n15511) );
  XNOR U17783 ( .A(n15517), .B(n15515), .Z(n17728) );
  AND U17784 ( .A(n17729), .B(n17730), .Z(n15515) );
  NANDN U17785 ( .A(n17731), .B(n17732), .Z(n17730) );
  OR U17786 ( .A(n17733), .B(n17734), .Z(n17732) );
  NAND U17787 ( .A(n17734), .B(n17733), .Z(n17729) );
  ANDN U17788 ( .B(B[2]), .A(n61), .Z(n15517) );
  XNOR U17789 ( .A(n15525), .B(n17735), .Z(n15518) );
  XNOR U17790 ( .A(n15524), .B(n15522), .Z(n17735) );
  AND U17791 ( .A(n17736), .B(n17737), .Z(n15522) );
  NANDN U17792 ( .A(n17738), .B(n17739), .Z(n17737) );
  NANDN U17793 ( .A(n17740), .B(n17741), .Z(n17739) );
  NANDN U17794 ( .A(n17741), .B(n17740), .Z(n17736) );
  ANDN U17795 ( .B(B[3]), .A(n62), .Z(n15524) );
  XNOR U17796 ( .A(n15532), .B(n17742), .Z(n15525) );
  XNOR U17797 ( .A(n15531), .B(n15529), .Z(n17742) );
  AND U17798 ( .A(n17743), .B(n17744), .Z(n15529) );
  NANDN U17799 ( .A(n17745), .B(n17746), .Z(n17744) );
  OR U17800 ( .A(n17747), .B(n17748), .Z(n17746) );
  NAND U17801 ( .A(n17748), .B(n17747), .Z(n17743) );
  ANDN U17802 ( .B(B[4]), .A(n63), .Z(n15531) );
  XNOR U17803 ( .A(n15539), .B(n17749), .Z(n15532) );
  XNOR U17804 ( .A(n15538), .B(n15536), .Z(n17749) );
  AND U17805 ( .A(n17750), .B(n17751), .Z(n15536) );
  NANDN U17806 ( .A(n17752), .B(n17753), .Z(n17751) );
  NANDN U17807 ( .A(n17754), .B(n17755), .Z(n17753) );
  NANDN U17808 ( .A(n17755), .B(n17754), .Z(n17750) );
  ANDN U17809 ( .B(B[5]), .A(n64), .Z(n15538) );
  XNOR U17810 ( .A(n15546), .B(n17756), .Z(n15539) );
  XNOR U17811 ( .A(n15545), .B(n15543), .Z(n17756) );
  AND U17812 ( .A(n17757), .B(n17758), .Z(n15543) );
  NANDN U17813 ( .A(n17759), .B(n17760), .Z(n17758) );
  OR U17814 ( .A(n17761), .B(n17762), .Z(n17760) );
  NAND U17815 ( .A(n17762), .B(n17761), .Z(n17757) );
  ANDN U17816 ( .B(B[6]), .A(n65), .Z(n15545) );
  XNOR U17817 ( .A(n15553), .B(n17763), .Z(n15546) );
  XNOR U17818 ( .A(n15552), .B(n15550), .Z(n17763) );
  AND U17819 ( .A(n17764), .B(n17765), .Z(n15550) );
  NANDN U17820 ( .A(n17766), .B(n17767), .Z(n17765) );
  NANDN U17821 ( .A(n17768), .B(n17769), .Z(n17767) );
  NANDN U17822 ( .A(n17769), .B(n17768), .Z(n17764) );
  ANDN U17823 ( .B(B[7]), .A(n66), .Z(n15552) );
  XNOR U17824 ( .A(n15560), .B(n17770), .Z(n15553) );
  XNOR U17825 ( .A(n15559), .B(n15557), .Z(n17770) );
  AND U17826 ( .A(n17771), .B(n17772), .Z(n15557) );
  NANDN U17827 ( .A(n17773), .B(n17774), .Z(n17772) );
  OR U17828 ( .A(n17775), .B(n17776), .Z(n17774) );
  NAND U17829 ( .A(n17776), .B(n17775), .Z(n17771) );
  ANDN U17830 ( .B(B[8]), .A(n67), .Z(n15559) );
  XNOR U17831 ( .A(n15567), .B(n17777), .Z(n15560) );
  XNOR U17832 ( .A(n15566), .B(n15564), .Z(n17777) );
  AND U17833 ( .A(n17778), .B(n17779), .Z(n15564) );
  NANDN U17834 ( .A(n17780), .B(n17781), .Z(n17779) );
  NANDN U17835 ( .A(n17782), .B(n17783), .Z(n17781) );
  NANDN U17836 ( .A(n17783), .B(n17782), .Z(n17778) );
  ANDN U17837 ( .B(B[9]), .A(n68), .Z(n15566) );
  XNOR U17838 ( .A(n15574), .B(n17784), .Z(n15567) );
  XNOR U17839 ( .A(n15573), .B(n15571), .Z(n17784) );
  AND U17840 ( .A(n17785), .B(n17786), .Z(n15571) );
  NANDN U17841 ( .A(n17787), .B(n17788), .Z(n17786) );
  OR U17842 ( .A(n17789), .B(n17790), .Z(n17788) );
  NAND U17843 ( .A(n17790), .B(n17789), .Z(n17785) );
  ANDN U17844 ( .B(B[10]), .A(n69), .Z(n15573) );
  XNOR U17845 ( .A(n15581), .B(n17791), .Z(n15574) );
  XNOR U17846 ( .A(n15580), .B(n15578), .Z(n17791) );
  AND U17847 ( .A(n17792), .B(n17793), .Z(n15578) );
  NANDN U17848 ( .A(n17794), .B(n17795), .Z(n17793) );
  NANDN U17849 ( .A(n17796), .B(n17797), .Z(n17795) );
  NANDN U17850 ( .A(n17797), .B(n17796), .Z(n17792) );
  ANDN U17851 ( .B(B[11]), .A(n70), .Z(n15580) );
  XNOR U17852 ( .A(n15588), .B(n17798), .Z(n15581) );
  XNOR U17853 ( .A(n15587), .B(n15585), .Z(n17798) );
  AND U17854 ( .A(n17799), .B(n17800), .Z(n15585) );
  NANDN U17855 ( .A(n17801), .B(n17802), .Z(n17800) );
  OR U17856 ( .A(n17803), .B(n17804), .Z(n17802) );
  NAND U17857 ( .A(n17804), .B(n17803), .Z(n17799) );
  ANDN U17858 ( .B(B[12]), .A(n71), .Z(n15587) );
  XNOR U17859 ( .A(n15595), .B(n17805), .Z(n15588) );
  XNOR U17860 ( .A(n15594), .B(n15592), .Z(n17805) );
  AND U17861 ( .A(n17806), .B(n17807), .Z(n15592) );
  NANDN U17862 ( .A(n17808), .B(n17809), .Z(n17807) );
  NANDN U17863 ( .A(n17810), .B(n17811), .Z(n17809) );
  NANDN U17864 ( .A(n17811), .B(n17810), .Z(n17806) );
  ANDN U17865 ( .B(B[13]), .A(n72), .Z(n15594) );
  XNOR U17866 ( .A(n15602), .B(n17812), .Z(n15595) );
  XNOR U17867 ( .A(n15601), .B(n15599), .Z(n17812) );
  AND U17868 ( .A(n17813), .B(n17814), .Z(n15599) );
  NANDN U17869 ( .A(n17815), .B(n17816), .Z(n17814) );
  OR U17870 ( .A(n17817), .B(n17818), .Z(n17816) );
  NAND U17871 ( .A(n17818), .B(n17817), .Z(n17813) );
  ANDN U17872 ( .B(B[14]), .A(n73), .Z(n15601) );
  XNOR U17873 ( .A(n15609), .B(n17819), .Z(n15602) );
  XNOR U17874 ( .A(n15608), .B(n15606), .Z(n17819) );
  AND U17875 ( .A(n17820), .B(n17821), .Z(n15606) );
  NANDN U17876 ( .A(n17822), .B(n17823), .Z(n17821) );
  NANDN U17877 ( .A(n17824), .B(n17825), .Z(n17823) );
  NANDN U17878 ( .A(n17825), .B(n17824), .Z(n17820) );
  ANDN U17879 ( .B(B[15]), .A(n74), .Z(n15608) );
  XNOR U17880 ( .A(n15616), .B(n17826), .Z(n15609) );
  XNOR U17881 ( .A(n15615), .B(n15613), .Z(n17826) );
  AND U17882 ( .A(n17827), .B(n17828), .Z(n15613) );
  NANDN U17883 ( .A(n17829), .B(n17830), .Z(n17828) );
  OR U17884 ( .A(n17831), .B(n17832), .Z(n17830) );
  NAND U17885 ( .A(n17832), .B(n17831), .Z(n17827) );
  ANDN U17886 ( .B(B[16]), .A(n75), .Z(n15615) );
  XNOR U17887 ( .A(n15623), .B(n17833), .Z(n15616) );
  XNOR U17888 ( .A(n15622), .B(n15620), .Z(n17833) );
  AND U17889 ( .A(n17834), .B(n17835), .Z(n15620) );
  NANDN U17890 ( .A(n17836), .B(n17837), .Z(n17835) );
  NANDN U17891 ( .A(n17838), .B(n17839), .Z(n17837) );
  NANDN U17892 ( .A(n17839), .B(n17838), .Z(n17834) );
  ANDN U17893 ( .B(B[17]), .A(n76), .Z(n15622) );
  XNOR U17894 ( .A(n15630), .B(n17840), .Z(n15623) );
  XNOR U17895 ( .A(n15629), .B(n15627), .Z(n17840) );
  AND U17896 ( .A(n17841), .B(n17842), .Z(n15627) );
  NANDN U17897 ( .A(n17843), .B(n17844), .Z(n17842) );
  OR U17898 ( .A(n17845), .B(n17846), .Z(n17844) );
  NAND U17899 ( .A(n17846), .B(n17845), .Z(n17841) );
  ANDN U17900 ( .B(B[18]), .A(n77), .Z(n15629) );
  XNOR U17901 ( .A(n15637), .B(n17847), .Z(n15630) );
  XNOR U17902 ( .A(n15636), .B(n15634), .Z(n17847) );
  AND U17903 ( .A(n17848), .B(n17849), .Z(n15634) );
  NANDN U17904 ( .A(n17850), .B(n17851), .Z(n17849) );
  NANDN U17905 ( .A(n17852), .B(n17853), .Z(n17851) );
  NANDN U17906 ( .A(n17853), .B(n17852), .Z(n17848) );
  ANDN U17907 ( .B(B[19]), .A(n78), .Z(n15636) );
  XNOR U17908 ( .A(n15644), .B(n17854), .Z(n15637) );
  XNOR U17909 ( .A(n15643), .B(n15641), .Z(n17854) );
  AND U17910 ( .A(n17855), .B(n17856), .Z(n15641) );
  NANDN U17911 ( .A(n17857), .B(n17858), .Z(n17856) );
  OR U17912 ( .A(n17859), .B(n17860), .Z(n17858) );
  NAND U17913 ( .A(n17860), .B(n17859), .Z(n17855) );
  ANDN U17914 ( .B(B[20]), .A(n79), .Z(n15643) );
  XNOR U17915 ( .A(n15651), .B(n17861), .Z(n15644) );
  XNOR U17916 ( .A(n15650), .B(n15648), .Z(n17861) );
  AND U17917 ( .A(n17862), .B(n17863), .Z(n15648) );
  NANDN U17918 ( .A(n17864), .B(n17865), .Z(n17863) );
  NANDN U17919 ( .A(n17866), .B(n17867), .Z(n17865) );
  NANDN U17920 ( .A(n17867), .B(n17866), .Z(n17862) );
  ANDN U17921 ( .B(B[21]), .A(n80), .Z(n15650) );
  XNOR U17922 ( .A(n15658), .B(n17868), .Z(n15651) );
  XNOR U17923 ( .A(n15657), .B(n15655), .Z(n17868) );
  AND U17924 ( .A(n17869), .B(n17870), .Z(n15655) );
  NANDN U17925 ( .A(n17871), .B(n17872), .Z(n17870) );
  OR U17926 ( .A(n17873), .B(n17874), .Z(n17872) );
  NAND U17927 ( .A(n17874), .B(n17873), .Z(n17869) );
  ANDN U17928 ( .B(B[22]), .A(n81), .Z(n15657) );
  XNOR U17929 ( .A(n15665), .B(n17875), .Z(n15658) );
  XNOR U17930 ( .A(n15664), .B(n15662), .Z(n17875) );
  AND U17931 ( .A(n17876), .B(n17877), .Z(n15662) );
  NANDN U17932 ( .A(n17878), .B(n17879), .Z(n17877) );
  NAND U17933 ( .A(n17880), .B(n17881), .Z(n17879) );
  ANDN U17934 ( .B(B[23]), .A(n82), .Z(n15664) );
  XOR U17935 ( .A(n15671), .B(n17882), .Z(n15665) );
  XNOR U17936 ( .A(n15669), .B(n15672), .Z(n17882) );
  NAND U17937 ( .A(A[2]), .B(B[24]), .Z(n15672) );
  NANDN U17938 ( .A(n17883), .B(n17884), .Z(n15669) );
  AND U17939 ( .A(A[0]), .B(B[25]), .Z(n17884) );
  XNOR U17940 ( .A(n15674), .B(n17885), .Z(n15671) );
  NAND U17941 ( .A(A[0]), .B(B[26]), .Z(n17885) );
  NAND U17942 ( .A(B[25]), .B(A[1]), .Z(n15674) );
  XOR U17943 ( .A(n294), .B(n293), .Z(\A1[249] ) );
  XOR U17944 ( .A(n17713), .B(n17886), .Z(n293) );
  XNOR U17945 ( .A(n17712), .B(n17710), .Z(n17886) );
  AND U17946 ( .A(n17887), .B(n17888), .Z(n17710) );
  NANDN U17947 ( .A(n17889), .B(n17890), .Z(n17888) );
  NANDN U17948 ( .A(n17891), .B(n17892), .Z(n17890) );
  NANDN U17949 ( .A(n17892), .B(n17891), .Z(n17887) );
  ANDN U17950 ( .B(B[220]), .A(n54), .Z(n17712) );
  XNOR U17951 ( .A(n17507), .B(n17893), .Z(n17713) );
  XNOR U17952 ( .A(n17506), .B(n17504), .Z(n17893) );
  AND U17953 ( .A(n17894), .B(n17895), .Z(n17504) );
  NANDN U17954 ( .A(n17896), .B(n17897), .Z(n17895) );
  OR U17955 ( .A(n17898), .B(n17899), .Z(n17897) );
  NAND U17956 ( .A(n17899), .B(n17898), .Z(n17894) );
  ANDN U17957 ( .B(B[221]), .A(n55), .Z(n17506) );
  XNOR U17958 ( .A(n17514), .B(n17900), .Z(n17507) );
  XNOR U17959 ( .A(n17513), .B(n17511), .Z(n17900) );
  AND U17960 ( .A(n17901), .B(n17902), .Z(n17511) );
  NANDN U17961 ( .A(n17903), .B(n17904), .Z(n17902) );
  NANDN U17962 ( .A(n17905), .B(n17906), .Z(n17904) );
  NANDN U17963 ( .A(n17906), .B(n17905), .Z(n17901) );
  ANDN U17964 ( .B(B[222]), .A(n56), .Z(n17513) );
  XNOR U17965 ( .A(n17521), .B(n17907), .Z(n17514) );
  XNOR U17966 ( .A(n17520), .B(n17518), .Z(n17907) );
  AND U17967 ( .A(n17908), .B(n17909), .Z(n17518) );
  NANDN U17968 ( .A(n17910), .B(n17911), .Z(n17909) );
  OR U17969 ( .A(n17912), .B(n17913), .Z(n17911) );
  NAND U17970 ( .A(n17913), .B(n17912), .Z(n17908) );
  ANDN U17971 ( .B(B[223]), .A(n57), .Z(n17520) );
  XNOR U17972 ( .A(n17528), .B(n17914), .Z(n17521) );
  XNOR U17973 ( .A(n17527), .B(n17525), .Z(n17914) );
  AND U17974 ( .A(n17915), .B(n17916), .Z(n17525) );
  NANDN U17975 ( .A(n17917), .B(n17918), .Z(n17916) );
  NANDN U17976 ( .A(n17919), .B(n17920), .Z(n17918) );
  NANDN U17977 ( .A(n17920), .B(n17919), .Z(n17915) );
  ANDN U17978 ( .B(B[224]), .A(n58), .Z(n17527) );
  XNOR U17979 ( .A(n17535), .B(n17921), .Z(n17528) );
  XNOR U17980 ( .A(n17534), .B(n17532), .Z(n17921) );
  AND U17981 ( .A(n17922), .B(n17923), .Z(n17532) );
  NANDN U17982 ( .A(n17924), .B(n17925), .Z(n17923) );
  OR U17983 ( .A(n17926), .B(n17927), .Z(n17925) );
  NAND U17984 ( .A(n17927), .B(n17926), .Z(n17922) );
  ANDN U17985 ( .B(B[225]), .A(n59), .Z(n17534) );
  XNOR U17986 ( .A(n17542), .B(n17928), .Z(n17535) );
  XNOR U17987 ( .A(n17541), .B(n17539), .Z(n17928) );
  AND U17988 ( .A(n17929), .B(n17930), .Z(n17539) );
  NANDN U17989 ( .A(n17931), .B(n17932), .Z(n17930) );
  NANDN U17990 ( .A(n17933), .B(n17934), .Z(n17932) );
  NANDN U17991 ( .A(n17934), .B(n17933), .Z(n17929) );
  ANDN U17992 ( .B(B[226]), .A(n60), .Z(n17541) );
  XNOR U17993 ( .A(n17549), .B(n17935), .Z(n17542) );
  XNOR U17994 ( .A(n17548), .B(n17546), .Z(n17935) );
  AND U17995 ( .A(n17936), .B(n17937), .Z(n17546) );
  NANDN U17996 ( .A(n17938), .B(n17939), .Z(n17937) );
  OR U17997 ( .A(n17940), .B(n17941), .Z(n17939) );
  NAND U17998 ( .A(n17941), .B(n17940), .Z(n17936) );
  ANDN U17999 ( .B(B[227]), .A(n61), .Z(n17548) );
  XNOR U18000 ( .A(n17556), .B(n17942), .Z(n17549) );
  XNOR U18001 ( .A(n17555), .B(n17553), .Z(n17942) );
  AND U18002 ( .A(n17943), .B(n17944), .Z(n17553) );
  NANDN U18003 ( .A(n17945), .B(n17946), .Z(n17944) );
  NANDN U18004 ( .A(n17947), .B(n17948), .Z(n17946) );
  NANDN U18005 ( .A(n17948), .B(n17947), .Z(n17943) );
  ANDN U18006 ( .B(B[228]), .A(n62), .Z(n17555) );
  XNOR U18007 ( .A(n17563), .B(n17949), .Z(n17556) );
  XNOR U18008 ( .A(n17562), .B(n17560), .Z(n17949) );
  AND U18009 ( .A(n17950), .B(n17951), .Z(n17560) );
  NANDN U18010 ( .A(n17952), .B(n17953), .Z(n17951) );
  OR U18011 ( .A(n17954), .B(n17955), .Z(n17953) );
  NAND U18012 ( .A(n17955), .B(n17954), .Z(n17950) );
  ANDN U18013 ( .B(B[229]), .A(n63), .Z(n17562) );
  XNOR U18014 ( .A(n17570), .B(n17956), .Z(n17563) );
  XNOR U18015 ( .A(n17569), .B(n17567), .Z(n17956) );
  AND U18016 ( .A(n17957), .B(n17958), .Z(n17567) );
  NANDN U18017 ( .A(n17959), .B(n17960), .Z(n17958) );
  NANDN U18018 ( .A(n17961), .B(n17962), .Z(n17960) );
  NANDN U18019 ( .A(n17962), .B(n17961), .Z(n17957) );
  ANDN U18020 ( .B(B[230]), .A(n64), .Z(n17569) );
  XNOR U18021 ( .A(n17577), .B(n17963), .Z(n17570) );
  XNOR U18022 ( .A(n17576), .B(n17574), .Z(n17963) );
  AND U18023 ( .A(n17964), .B(n17965), .Z(n17574) );
  NANDN U18024 ( .A(n17966), .B(n17967), .Z(n17965) );
  OR U18025 ( .A(n17968), .B(n17969), .Z(n17967) );
  NAND U18026 ( .A(n17969), .B(n17968), .Z(n17964) );
  ANDN U18027 ( .B(B[231]), .A(n65), .Z(n17576) );
  XNOR U18028 ( .A(n17584), .B(n17970), .Z(n17577) );
  XNOR U18029 ( .A(n17583), .B(n17581), .Z(n17970) );
  AND U18030 ( .A(n17971), .B(n17972), .Z(n17581) );
  NANDN U18031 ( .A(n17973), .B(n17974), .Z(n17972) );
  NANDN U18032 ( .A(n17975), .B(n17976), .Z(n17974) );
  NANDN U18033 ( .A(n17976), .B(n17975), .Z(n17971) );
  ANDN U18034 ( .B(B[232]), .A(n66), .Z(n17583) );
  XNOR U18035 ( .A(n17591), .B(n17977), .Z(n17584) );
  XNOR U18036 ( .A(n17590), .B(n17588), .Z(n17977) );
  AND U18037 ( .A(n17978), .B(n17979), .Z(n17588) );
  NANDN U18038 ( .A(n17980), .B(n17981), .Z(n17979) );
  OR U18039 ( .A(n17982), .B(n17983), .Z(n17981) );
  NAND U18040 ( .A(n17983), .B(n17982), .Z(n17978) );
  ANDN U18041 ( .B(B[233]), .A(n67), .Z(n17590) );
  XNOR U18042 ( .A(n17598), .B(n17984), .Z(n17591) );
  XNOR U18043 ( .A(n17597), .B(n17595), .Z(n17984) );
  AND U18044 ( .A(n17985), .B(n17986), .Z(n17595) );
  NANDN U18045 ( .A(n17987), .B(n17988), .Z(n17986) );
  NANDN U18046 ( .A(n17989), .B(n17990), .Z(n17988) );
  NANDN U18047 ( .A(n17990), .B(n17989), .Z(n17985) );
  ANDN U18048 ( .B(B[234]), .A(n68), .Z(n17597) );
  XNOR U18049 ( .A(n17605), .B(n17991), .Z(n17598) );
  XNOR U18050 ( .A(n17604), .B(n17602), .Z(n17991) );
  AND U18051 ( .A(n17992), .B(n17993), .Z(n17602) );
  NANDN U18052 ( .A(n17994), .B(n17995), .Z(n17993) );
  OR U18053 ( .A(n17996), .B(n17997), .Z(n17995) );
  NAND U18054 ( .A(n17997), .B(n17996), .Z(n17992) );
  ANDN U18055 ( .B(B[235]), .A(n69), .Z(n17604) );
  XNOR U18056 ( .A(n17612), .B(n17998), .Z(n17605) );
  XNOR U18057 ( .A(n17611), .B(n17609), .Z(n17998) );
  AND U18058 ( .A(n17999), .B(n18000), .Z(n17609) );
  NANDN U18059 ( .A(n18001), .B(n18002), .Z(n18000) );
  NANDN U18060 ( .A(n18003), .B(n18004), .Z(n18002) );
  NANDN U18061 ( .A(n18004), .B(n18003), .Z(n17999) );
  ANDN U18062 ( .B(B[236]), .A(n70), .Z(n17611) );
  XNOR U18063 ( .A(n17619), .B(n18005), .Z(n17612) );
  XNOR U18064 ( .A(n17618), .B(n17616), .Z(n18005) );
  AND U18065 ( .A(n18006), .B(n18007), .Z(n17616) );
  NANDN U18066 ( .A(n18008), .B(n18009), .Z(n18007) );
  OR U18067 ( .A(n18010), .B(n18011), .Z(n18009) );
  NAND U18068 ( .A(n18011), .B(n18010), .Z(n18006) );
  ANDN U18069 ( .B(B[237]), .A(n71), .Z(n17618) );
  XNOR U18070 ( .A(n17626), .B(n18012), .Z(n17619) );
  XNOR U18071 ( .A(n17625), .B(n17623), .Z(n18012) );
  AND U18072 ( .A(n18013), .B(n18014), .Z(n17623) );
  NANDN U18073 ( .A(n18015), .B(n18016), .Z(n18014) );
  NANDN U18074 ( .A(n18017), .B(n18018), .Z(n18016) );
  NANDN U18075 ( .A(n18018), .B(n18017), .Z(n18013) );
  ANDN U18076 ( .B(B[238]), .A(n72), .Z(n17625) );
  XNOR U18077 ( .A(n17633), .B(n18019), .Z(n17626) );
  XNOR U18078 ( .A(n17632), .B(n17630), .Z(n18019) );
  AND U18079 ( .A(n18020), .B(n18021), .Z(n17630) );
  NANDN U18080 ( .A(n18022), .B(n18023), .Z(n18021) );
  OR U18081 ( .A(n18024), .B(n18025), .Z(n18023) );
  NAND U18082 ( .A(n18025), .B(n18024), .Z(n18020) );
  ANDN U18083 ( .B(B[239]), .A(n73), .Z(n17632) );
  XNOR U18084 ( .A(n17640), .B(n18026), .Z(n17633) );
  XNOR U18085 ( .A(n17639), .B(n17637), .Z(n18026) );
  AND U18086 ( .A(n18027), .B(n18028), .Z(n17637) );
  NANDN U18087 ( .A(n18029), .B(n18030), .Z(n18028) );
  NANDN U18088 ( .A(n18031), .B(n18032), .Z(n18030) );
  NANDN U18089 ( .A(n18032), .B(n18031), .Z(n18027) );
  ANDN U18090 ( .B(B[240]), .A(n74), .Z(n17639) );
  XNOR U18091 ( .A(n17647), .B(n18033), .Z(n17640) );
  XNOR U18092 ( .A(n17646), .B(n17644), .Z(n18033) );
  AND U18093 ( .A(n18034), .B(n18035), .Z(n17644) );
  NANDN U18094 ( .A(n18036), .B(n18037), .Z(n18035) );
  OR U18095 ( .A(n18038), .B(n18039), .Z(n18037) );
  NAND U18096 ( .A(n18039), .B(n18038), .Z(n18034) );
  ANDN U18097 ( .B(B[241]), .A(n75), .Z(n17646) );
  XNOR U18098 ( .A(n17654), .B(n18040), .Z(n17647) );
  XNOR U18099 ( .A(n17653), .B(n17651), .Z(n18040) );
  AND U18100 ( .A(n18041), .B(n18042), .Z(n17651) );
  NANDN U18101 ( .A(n18043), .B(n18044), .Z(n18042) );
  NANDN U18102 ( .A(n18045), .B(n18046), .Z(n18044) );
  NANDN U18103 ( .A(n18046), .B(n18045), .Z(n18041) );
  ANDN U18104 ( .B(B[242]), .A(n76), .Z(n17653) );
  XNOR U18105 ( .A(n17661), .B(n18047), .Z(n17654) );
  XNOR U18106 ( .A(n17660), .B(n17658), .Z(n18047) );
  AND U18107 ( .A(n18048), .B(n18049), .Z(n17658) );
  NANDN U18108 ( .A(n18050), .B(n18051), .Z(n18049) );
  OR U18109 ( .A(n18052), .B(n18053), .Z(n18051) );
  NAND U18110 ( .A(n18053), .B(n18052), .Z(n18048) );
  ANDN U18111 ( .B(B[243]), .A(n77), .Z(n17660) );
  XNOR U18112 ( .A(n17668), .B(n18054), .Z(n17661) );
  XNOR U18113 ( .A(n17667), .B(n17665), .Z(n18054) );
  AND U18114 ( .A(n18055), .B(n18056), .Z(n17665) );
  NANDN U18115 ( .A(n18057), .B(n18058), .Z(n18056) );
  NANDN U18116 ( .A(n18059), .B(n18060), .Z(n18058) );
  NANDN U18117 ( .A(n18060), .B(n18059), .Z(n18055) );
  ANDN U18118 ( .B(B[244]), .A(n78), .Z(n17667) );
  XNOR U18119 ( .A(n17675), .B(n18061), .Z(n17668) );
  XNOR U18120 ( .A(n17674), .B(n17672), .Z(n18061) );
  AND U18121 ( .A(n18062), .B(n18063), .Z(n17672) );
  NANDN U18122 ( .A(n18064), .B(n18065), .Z(n18063) );
  OR U18123 ( .A(n18066), .B(n18067), .Z(n18065) );
  NAND U18124 ( .A(n18067), .B(n18066), .Z(n18062) );
  ANDN U18125 ( .B(B[245]), .A(n79), .Z(n17674) );
  XNOR U18126 ( .A(n17682), .B(n18068), .Z(n17675) );
  XNOR U18127 ( .A(n17681), .B(n17679), .Z(n18068) );
  AND U18128 ( .A(n18069), .B(n18070), .Z(n17679) );
  NANDN U18129 ( .A(n18071), .B(n18072), .Z(n18070) );
  NANDN U18130 ( .A(n18073), .B(n18074), .Z(n18072) );
  NANDN U18131 ( .A(n18074), .B(n18073), .Z(n18069) );
  ANDN U18132 ( .B(B[246]), .A(n80), .Z(n17681) );
  XNOR U18133 ( .A(n17689), .B(n18075), .Z(n17682) );
  XNOR U18134 ( .A(n17688), .B(n17686), .Z(n18075) );
  AND U18135 ( .A(n18076), .B(n18077), .Z(n17686) );
  NANDN U18136 ( .A(n18078), .B(n18079), .Z(n18077) );
  OR U18137 ( .A(n18080), .B(n18081), .Z(n18079) );
  NAND U18138 ( .A(n18081), .B(n18080), .Z(n18076) );
  ANDN U18139 ( .B(B[247]), .A(n81), .Z(n17688) );
  XNOR U18140 ( .A(n17696), .B(n18082), .Z(n17689) );
  XNOR U18141 ( .A(n17695), .B(n17693), .Z(n18082) );
  AND U18142 ( .A(n18083), .B(n18084), .Z(n17693) );
  NANDN U18143 ( .A(n18085), .B(n18086), .Z(n18084) );
  NAND U18144 ( .A(n18087), .B(n18088), .Z(n18086) );
  ANDN U18145 ( .B(B[248]), .A(n82), .Z(n17695) );
  XOR U18146 ( .A(n17702), .B(n18089), .Z(n17696) );
  XNOR U18147 ( .A(n17700), .B(n17703), .Z(n18089) );
  NAND U18148 ( .A(A[2]), .B(B[249]), .Z(n17703) );
  NANDN U18149 ( .A(n18090), .B(n18091), .Z(n17700) );
  AND U18150 ( .A(A[0]), .B(B[250]), .Z(n18091) );
  XNOR U18151 ( .A(n17705), .B(n18092), .Z(n17702) );
  NAND U18152 ( .A(A[0]), .B(B[251]), .Z(n18092) );
  NAND U18153 ( .A(B[250]), .B(A[1]), .Z(n17705) );
  NAND U18154 ( .A(n18093), .B(n18094), .Z(n294) );
  NANDN U18155 ( .A(n18095), .B(n18096), .Z(n18094) );
  OR U18156 ( .A(n18097), .B(n18098), .Z(n18096) );
  NAND U18157 ( .A(n18098), .B(n18097), .Z(n18093) );
  XOR U18158 ( .A(n296), .B(n295), .Z(\A1[248] ) );
  XOR U18159 ( .A(n18098), .B(n18099), .Z(n295) );
  XNOR U18160 ( .A(n18097), .B(n18095), .Z(n18099) );
  AND U18161 ( .A(n18100), .B(n18101), .Z(n18095) );
  NANDN U18162 ( .A(n18102), .B(n18103), .Z(n18101) );
  NANDN U18163 ( .A(n18104), .B(n18105), .Z(n18103) );
  NANDN U18164 ( .A(n18105), .B(n18104), .Z(n18100) );
  ANDN U18165 ( .B(B[219]), .A(n54), .Z(n18097) );
  XNOR U18166 ( .A(n17892), .B(n18106), .Z(n18098) );
  XNOR U18167 ( .A(n17891), .B(n17889), .Z(n18106) );
  AND U18168 ( .A(n18107), .B(n18108), .Z(n17889) );
  NANDN U18169 ( .A(n18109), .B(n18110), .Z(n18108) );
  OR U18170 ( .A(n18111), .B(n18112), .Z(n18110) );
  NAND U18171 ( .A(n18112), .B(n18111), .Z(n18107) );
  ANDN U18172 ( .B(B[220]), .A(n55), .Z(n17891) );
  XNOR U18173 ( .A(n17899), .B(n18113), .Z(n17892) );
  XNOR U18174 ( .A(n17898), .B(n17896), .Z(n18113) );
  AND U18175 ( .A(n18114), .B(n18115), .Z(n17896) );
  NANDN U18176 ( .A(n18116), .B(n18117), .Z(n18115) );
  NANDN U18177 ( .A(n18118), .B(n18119), .Z(n18117) );
  NANDN U18178 ( .A(n18119), .B(n18118), .Z(n18114) );
  ANDN U18179 ( .B(B[221]), .A(n56), .Z(n17898) );
  XNOR U18180 ( .A(n17906), .B(n18120), .Z(n17899) );
  XNOR U18181 ( .A(n17905), .B(n17903), .Z(n18120) );
  AND U18182 ( .A(n18121), .B(n18122), .Z(n17903) );
  NANDN U18183 ( .A(n18123), .B(n18124), .Z(n18122) );
  OR U18184 ( .A(n18125), .B(n18126), .Z(n18124) );
  NAND U18185 ( .A(n18126), .B(n18125), .Z(n18121) );
  ANDN U18186 ( .B(B[222]), .A(n57), .Z(n17905) );
  XNOR U18187 ( .A(n17913), .B(n18127), .Z(n17906) );
  XNOR U18188 ( .A(n17912), .B(n17910), .Z(n18127) );
  AND U18189 ( .A(n18128), .B(n18129), .Z(n17910) );
  NANDN U18190 ( .A(n18130), .B(n18131), .Z(n18129) );
  NANDN U18191 ( .A(n18132), .B(n18133), .Z(n18131) );
  NANDN U18192 ( .A(n18133), .B(n18132), .Z(n18128) );
  ANDN U18193 ( .B(B[223]), .A(n58), .Z(n17912) );
  XNOR U18194 ( .A(n17920), .B(n18134), .Z(n17913) );
  XNOR U18195 ( .A(n17919), .B(n17917), .Z(n18134) );
  AND U18196 ( .A(n18135), .B(n18136), .Z(n17917) );
  NANDN U18197 ( .A(n18137), .B(n18138), .Z(n18136) );
  OR U18198 ( .A(n18139), .B(n18140), .Z(n18138) );
  NAND U18199 ( .A(n18140), .B(n18139), .Z(n18135) );
  ANDN U18200 ( .B(B[224]), .A(n59), .Z(n17919) );
  XNOR U18201 ( .A(n17927), .B(n18141), .Z(n17920) );
  XNOR U18202 ( .A(n17926), .B(n17924), .Z(n18141) );
  AND U18203 ( .A(n18142), .B(n18143), .Z(n17924) );
  NANDN U18204 ( .A(n18144), .B(n18145), .Z(n18143) );
  NANDN U18205 ( .A(n18146), .B(n18147), .Z(n18145) );
  NANDN U18206 ( .A(n18147), .B(n18146), .Z(n18142) );
  ANDN U18207 ( .B(B[225]), .A(n60), .Z(n17926) );
  XNOR U18208 ( .A(n17934), .B(n18148), .Z(n17927) );
  XNOR U18209 ( .A(n17933), .B(n17931), .Z(n18148) );
  AND U18210 ( .A(n18149), .B(n18150), .Z(n17931) );
  NANDN U18211 ( .A(n18151), .B(n18152), .Z(n18150) );
  OR U18212 ( .A(n18153), .B(n18154), .Z(n18152) );
  NAND U18213 ( .A(n18154), .B(n18153), .Z(n18149) );
  ANDN U18214 ( .B(B[226]), .A(n61), .Z(n17933) );
  XNOR U18215 ( .A(n17941), .B(n18155), .Z(n17934) );
  XNOR U18216 ( .A(n17940), .B(n17938), .Z(n18155) );
  AND U18217 ( .A(n18156), .B(n18157), .Z(n17938) );
  NANDN U18218 ( .A(n18158), .B(n18159), .Z(n18157) );
  NANDN U18219 ( .A(n18160), .B(n18161), .Z(n18159) );
  NANDN U18220 ( .A(n18161), .B(n18160), .Z(n18156) );
  ANDN U18221 ( .B(B[227]), .A(n62), .Z(n17940) );
  XNOR U18222 ( .A(n17948), .B(n18162), .Z(n17941) );
  XNOR U18223 ( .A(n17947), .B(n17945), .Z(n18162) );
  AND U18224 ( .A(n18163), .B(n18164), .Z(n17945) );
  NANDN U18225 ( .A(n18165), .B(n18166), .Z(n18164) );
  OR U18226 ( .A(n18167), .B(n18168), .Z(n18166) );
  NAND U18227 ( .A(n18168), .B(n18167), .Z(n18163) );
  ANDN U18228 ( .B(B[228]), .A(n63), .Z(n17947) );
  XNOR U18229 ( .A(n17955), .B(n18169), .Z(n17948) );
  XNOR U18230 ( .A(n17954), .B(n17952), .Z(n18169) );
  AND U18231 ( .A(n18170), .B(n18171), .Z(n17952) );
  NANDN U18232 ( .A(n18172), .B(n18173), .Z(n18171) );
  NANDN U18233 ( .A(n18174), .B(n18175), .Z(n18173) );
  NANDN U18234 ( .A(n18175), .B(n18174), .Z(n18170) );
  ANDN U18235 ( .B(B[229]), .A(n64), .Z(n17954) );
  XNOR U18236 ( .A(n17962), .B(n18176), .Z(n17955) );
  XNOR U18237 ( .A(n17961), .B(n17959), .Z(n18176) );
  AND U18238 ( .A(n18177), .B(n18178), .Z(n17959) );
  NANDN U18239 ( .A(n18179), .B(n18180), .Z(n18178) );
  OR U18240 ( .A(n18181), .B(n18182), .Z(n18180) );
  NAND U18241 ( .A(n18182), .B(n18181), .Z(n18177) );
  ANDN U18242 ( .B(B[230]), .A(n65), .Z(n17961) );
  XNOR U18243 ( .A(n17969), .B(n18183), .Z(n17962) );
  XNOR U18244 ( .A(n17968), .B(n17966), .Z(n18183) );
  AND U18245 ( .A(n18184), .B(n18185), .Z(n17966) );
  NANDN U18246 ( .A(n18186), .B(n18187), .Z(n18185) );
  NANDN U18247 ( .A(n18188), .B(n18189), .Z(n18187) );
  NANDN U18248 ( .A(n18189), .B(n18188), .Z(n18184) );
  ANDN U18249 ( .B(B[231]), .A(n66), .Z(n17968) );
  XNOR U18250 ( .A(n17976), .B(n18190), .Z(n17969) );
  XNOR U18251 ( .A(n17975), .B(n17973), .Z(n18190) );
  AND U18252 ( .A(n18191), .B(n18192), .Z(n17973) );
  NANDN U18253 ( .A(n18193), .B(n18194), .Z(n18192) );
  OR U18254 ( .A(n18195), .B(n18196), .Z(n18194) );
  NAND U18255 ( .A(n18196), .B(n18195), .Z(n18191) );
  ANDN U18256 ( .B(B[232]), .A(n67), .Z(n17975) );
  XNOR U18257 ( .A(n17983), .B(n18197), .Z(n17976) );
  XNOR U18258 ( .A(n17982), .B(n17980), .Z(n18197) );
  AND U18259 ( .A(n18198), .B(n18199), .Z(n17980) );
  NANDN U18260 ( .A(n18200), .B(n18201), .Z(n18199) );
  NANDN U18261 ( .A(n18202), .B(n18203), .Z(n18201) );
  NANDN U18262 ( .A(n18203), .B(n18202), .Z(n18198) );
  ANDN U18263 ( .B(B[233]), .A(n68), .Z(n17982) );
  XNOR U18264 ( .A(n17990), .B(n18204), .Z(n17983) );
  XNOR U18265 ( .A(n17989), .B(n17987), .Z(n18204) );
  AND U18266 ( .A(n18205), .B(n18206), .Z(n17987) );
  NANDN U18267 ( .A(n18207), .B(n18208), .Z(n18206) );
  OR U18268 ( .A(n18209), .B(n18210), .Z(n18208) );
  NAND U18269 ( .A(n18210), .B(n18209), .Z(n18205) );
  ANDN U18270 ( .B(B[234]), .A(n69), .Z(n17989) );
  XNOR U18271 ( .A(n17997), .B(n18211), .Z(n17990) );
  XNOR U18272 ( .A(n17996), .B(n17994), .Z(n18211) );
  AND U18273 ( .A(n18212), .B(n18213), .Z(n17994) );
  NANDN U18274 ( .A(n18214), .B(n18215), .Z(n18213) );
  NANDN U18275 ( .A(n18216), .B(n18217), .Z(n18215) );
  NANDN U18276 ( .A(n18217), .B(n18216), .Z(n18212) );
  ANDN U18277 ( .B(B[235]), .A(n70), .Z(n17996) );
  XNOR U18278 ( .A(n18004), .B(n18218), .Z(n17997) );
  XNOR U18279 ( .A(n18003), .B(n18001), .Z(n18218) );
  AND U18280 ( .A(n18219), .B(n18220), .Z(n18001) );
  NANDN U18281 ( .A(n18221), .B(n18222), .Z(n18220) );
  OR U18282 ( .A(n18223), .B(n18224), .Z(n18222) );
  NAND U18283 ( .A(n18224), .B(n18223), .Z(n18219) );
  ANDN U18284 ( .B(B[236]), .A(n71), .Z(n18003) );
  XNOR U18285 ( .A(n18011), .B(n18225), .Z(n18004) );
  XNOR U18286 ( .A(n18010), .B(n18008), .Z(n18225) );
  AND U18287 ( .A(n18226), .B(n18227), .Z(n18008) );
  NANDN U18288 ( .A(n18228), .B(n18229), .Z(n18227) );
  NANDN U18289 ( .A(n18230), .B(n18231), .Z(n18229) );
  NANDN U18290 ( .A(n18231), .B(n18230), .Z(n18226) );
  ANDN U18291 ( .B(B[237]), .A(n72), .Z(n18010) );
  XNOR U18292 ( .A(n18018), .B(n18232), .Z(n18011) );
  XNOR U18293 ( .A(n18017), .B(n18015), .Z(n18232) );
  AND U18294 ( .A(n18233), .B(n18234), .Z(n18015) );
  NANDN U18295 ( .A(n18235), .B(n18236), .Z(n18234) );
  OR U18296 ( .A(n18237), .B(n18238), .Z(n18236) );
  NAND U18297 ( .A(n18238), .B(n18237), .Z(n18233) );
  ANDN U18298 ( .B(B[238]), .A(n73), .Z(n18017) );
  XNOR U18299 ( .A(n18025), .B(n18239), .Z(n18018) );
  XNOR U18300 ( .A(n18024), .B(n18022), .Z(n18239) );
  AND U18301 ( .A(n18240), .B(n18241), .Z(n18022) );
  NANDN U18302 ( .A(n18242), .B(n18243), .Z(n18241) );
  NANDN U18303 ( .A(n18244), .B(n18245), .Z(n18243) );
  NANDN U18304 ( .A(n18245), .B(n18244), .Z(n18240) );
  ANDN U18305 ( .B(B[239]), .A(n74), .Z(n18024) );
  XNOR U18306 ( .A(n18032), .B(n18246), .Z(n18025) );
  XNOR U18307 ( .A(n18031), .B(n18029), .Z(n18246) );
  AND U18308 ( .A(n18247), .B(n18248), .Z(n18029) );
  NANDN U18309 ( .A(n18249), .B(n18250), .Z(n18248) );
  OR U18310 ( .A(n18251), .B(n18252), .Z(n18250) );
  NAND U18311 ( .A(n18252), .B(n18251), .Z(n18247) );
  ANDN U18312 ( .B(B[240]), .A(n75), .Z(n18031) );
  XNOR U18313 ( .A(n18039), .B(n18253), .Z(n18032) );
  XNOR U18314 ( .A(n18038), .B(n18036), .Z(n18253) );
  AND U18315 ( .A(n18254), .B(n18255), .Z(n18036) );
  NANDN U18316 ( .A(n18256), .B(n18257), .Z(n18255) );
  NANDN U18317 ( .A(n18258), .B(n18259), .Z(n18257) );
  NANDN U18318 ( .A(n18259), .B(n18258), .Z(n18254) );
  ANDN U18319 ( .B(B[241]), .A(n76), .Z(n18038) );
  XNOR U18320 ( .A(n18046), .B(n18260), .Z(n18039) );
  XNOR U18321 ( .A(n18045), .B(n18043), .Z(n18260) );
  AND U18322 ( .A(n18261), .B(n18262), .Z(n18043) );
  NANDN U18323 ( .A(n18263), .B(n18264), .Z(n18262) );
  OR U18324 ( .A(n18265), .B(n18266), .Z(n18264) );
  NAND U18325 ( .A(n18266), .B(n18265), .Z(n18261) );
  ANDN U18326 ( .B(B[242]), .A(n77), .Z(n18045) );
  XNOR U18327 ( .A(n18053), .B(n18267), .Z(n18046) );
  XNOR U18328 ( .A(n18052), .B(n18050), .Z(n18267) );
  AND U18329 ( .A(n18268), .B(n18269), .Z(n18050) );
  NANDN U18330 ( .A(n18270), .B(n18271), .Z(n18269) );
  NANDN U18331 ( .A(n18272), .B(n18273), .Z(n18271) );
  NANDN U18332 ( .A(n18273), .B(n18272), .Z(n18268) );
  ANDN U18333 ( .B(B[243]), .A(n78), .Z(n18052) );
  XNOR U18334 ( .A(n18060), .B(n18274), .Z(n18053) );
  XNOR U18335 ( .A(n18059), .B(n18057), .Z(n18274) );
  AND U18336 ( .A(n18275), .B(n18276), .Z(n18057) );
  NANDN U18337 ( .A(n18277), .B(n18278), .Z(n18276) );
  OR U18338 ( .A(n18279), .B(n18280), .Z(n18278) );
  NAND U18339 ( .A(n18280), .B(n18279), .Z(n18275) );
  ANDN U18340 ( .B(B[244]), .A(n79), .Z(n18059) );
  XNOR U18341 ( .A(n18067), .B(n18281), .Z(n18060) );
  XNOR U18342 ( .A(n18066), .B(n18064), .Z(n18281) );
  AND U18343 ( .A(n18282), .B(n18283), .Z(n18064) );
  NANDN U18344 ( .A(n18284), .B(n18285), .Z(n18283) );
  NANDN U18345 ( .A(n18286), .B(n18287), .Z(n18285) );
  NANDN U18346 ( .A(n18287), .B(n18286), .Z(n18282) );
  ANDN U18347 ( .B(B[245]), .A(n80), .Z(n18066) );
  XNOR U18348 ( .A(n18074), .B(n18288), .Z(n18067) );
  XNOR U18349 ( .A(n18073), .B(n18071), .Z(n18288) );
  AND U18350 ( .A(n18289), .B(n18290), .Z(n18071) );
  NANDN U18351 ( .A(n18291), .B(n18292), .Z(n18290) );
  OR U18352 ( .A(n18293), .B(n18294), .Z(n18292) );
  NAND U18353 ( .A(n18294), .B(n18293), .Z(n18289) );
  ANDN U18354 ( .B(B[246]), .A(n81), .Z(n18073) );
  XNOR U18355 ( .A(n18081), .B(n18295), .Z(n18074) );
  XNOR U18356 ( .A(n18080), .B(n18078), .Z(n18295) );
  AND U18357 ( .A(n18296), .B(n18297), .Z(n18078) );
  NANDN U18358 ( .A(n18298), .B(n18299), .Z(n18297) );
  NAND U18359 ( .A(n18300), .B(n18301), .Z(n18299) );
  ANDN U18360 ( .B(B[247]), .A(n82), .Z(n18080) );
  XOR U18361 ( .A(n18087), .B(n18302), .Z(n18081) );
  XNOR U18362 ( .A(n18085), .B(n18088), .Z(n18302) );
  NAND U18363 ( .A(A[2]), .B(B[248]), .Z(n18088) );
  NANDN U18364 ( .A(n18303), .B(n18304), .Z(n18085) );
  AND U18365 ( .A(A[0]), .B(B[249]), .Z(n18304) );
  XNOR U18366 ( .A(n18090), .B(n18305), .Z(n18087) );
  NAND U18367 ( .A(A[0]), .B(B[250]), .Z(n18305) );
  NAND U18368 ( .A(B[249]), .B(A[1]), .Z(n18090) );
  NAND U18369 ( .A(n18306), .B(n18307), .Z(n296) );
  NANDN U18370 ( .A(n18308), .B(n18309), .Z(n18307) );
  OR U18371 ( .A(n18310), .B(n18311), .Z(n18309) );
  NAND U18372 ( .A(n18311), .B(n18310), .Z(n18306) );
  XOR U18373 ( .A(n298), .B(n297), .Z(\A1[247] ) );
  XOR U18374 ( .A(n18311), .B(n18312), .Z(n297) );
  XNOR U18375 ( .A(n18310), .B(n18308), .Z(n18312) );
  AND U18376 ( .A(n18313), .B(n18314), .Z(n18308) );
  NANDN U18377 ( .A(n18315), .B(n18316), .Z(n18314) );
  NANDN U18378 ( .A(n18317), .B(n18318), .Z(n18316) );
  NANDN U18379 ( .A(n18318), .B(n18317), .Z(n18313) );
  ANDN U18380 ( .B(B[218]), .A(n54), .Z(n18310) );
  XNOR U18381 ( .A(n18105), .B(n18319), .Z(n18311) );
  XNOR U18382 ( .A(n18104), .B(n18102), .Z(n18319) );
  AND U18383 ( .A(n18320), .B(n18321), .Z(n18102) );
  NANDN U18384 ( .A(n18322), .B(n18323), .Z(n18321) );
  OR U18385 ( .A(n18324), .B(n18325), .Z(n18323) );
  NAND U18386 ( .A(n18325), .B(n18324), .Z(n18320) );
  ANDN U18387 ( .B(B[219]), .A(n55), .Z(n18104) );
  XNOR U18388 ( .A(n18112), .B(n18326), .Z(n18105) );
  XNOR U18389 ( .A(n18111), .B(n18109), .Z(n18326) );
  AND U18390 ( .A(n18327), .B(n18328), .Z(n18109) );
  NANDN U18391 ( .A(n18329), .B(n18330), .Z(n18328) );
  NANDN U18392 ( .A(n18331), .B(n18332), .Z(n18330) );
  NANDN U18393 ( .A(n18332), .B(n18331), .Z(n18327) );
  ANDN U18394 ( .B(B[220]), .A(n56), .Z(n18111) );
  XNOR U18395 ( .A(n18119), .B(n18333), .Z(n18112) );
  XNOR U18396 ( .A(n18118), .B(n18116), .Z(n18333) );
  AND U18397 ( .A(n18334), .B(n18335), .Z(n18116) );
  NANDN U18398 ( .A(n18336), .B(n18337), .Z(n18335) );
  OR U18399 ( .A(n18338), .B(n18339), .Z(n18337) );
  NAND U18400 ( .A(n18339), .B(n18338), .Z(n18334) );
  ANDN U18401 ( .B(B[221]), .A(n57), .Z(n18118) );
  XNOR U18402 ( .A(n18126), .B(n18340), .Z(n18119) );
  XNOR U18403 ( .A(n18125), .B(n18123), .Z(n18340) );
  AND U18404 ( .A(n18341), .B(n18342), .Z(n18123) );
  NANDN U18405 ( .A(n18343), .B(n18344), .Z(n18342) );
  NANDN U18406 ( .A(n18345), .B(n18346), .Z(n18344) );
  NANDN U18407 ( .A(n18346), .B(n18345), .Z(n18341) );
  ANDN U18408 ( .B(B[222]), .A(n58), .Z(n18125) );
  XNOR U18409 ( .A(n18133), .B(n18347), .Z(n18126) );
  XNOR U18410 ( .A(n18132), .B(n18130), .Z(n18347) );
  AND U18411 ( .A(n18348), .B(n18349), .Z(n18130) );
  NANDN U18412 ( .A(n18350), .B(n18351), .Z(n18349) );
  OR U18413 ( .A(n18352), .B(n18353), .Z(n18351) );
  NAND U18414 ( .A(n18353), .B(n18352), .Z(n18348) );
  ANDN U18415 ( .B(B[223]), .A(n59), .Z(n18132) );
  XNOR U18416 ( .A(n18140), .B(n18354), .Z(n18133) );
  XNOR U18417 ( .A(n18139), .B(n18137), .Z(n18354) );
  AND U18418 ( .A(n18355), .B(n18356), .Z(n18137) );
  NANDN U18419 ( .A(n18357), .B(n18358), .Z(n18356) );
  NANDN U18420 ( .A(n18359), .B(n18360), .Z(n18358) );
  NANDN U18421 ( .A(n18360), .B(n18359), .Z(n18355) );
  ANDN U18422 ( .B(B[224]), .A(n60), .Z(n18139) );
  XNOR U18423 ( .A(n18147), .B(n18361), .Z(n18140) );
  XNOR U18424 ( .A(n18146), .B(n18144), .Z(n18361) );
  AND U18425 ( .A(n18362), .B(n18363), .Z(n18144) );
  NANDN U18426 ( .A(n18364), .B(n18365), .Z(n18363) );
  OR U18427 ( .A(n18366), .B(n18367), .Z(n18365) );
  NAND U18428 ( .A(n18367), .B(n18366), .Z(n18362) );
  ANDN U18429 ( .B(B[225]), .A(n61), .Z(n18146) );
  XNOR U18430 ( .A(n18154), .B(n18368), .Z(n18147) );
  XNOR U18431 ( .A(n18153), .B(n18151), .Z(n18368) );
  AND U18432 ( .A(n18369), .B(n18370), .Z(n18151) );
  NANDN U18433 ( .A(n18371), .B(n18372), .Z(n18370) );
  NANDN U18434 ( .A(n18373), .B(n18374), .Z(n18372) );
  NANDN U18435 ( .A(n18374), .B(n18373), .Z(n18369) );
  ANDN U18436 ( .B(B[226]), .A(n62), .Z(n18153) );
  XNOR U18437 ( .A(n18161), .B(n18375), .Z(n18154) );
  XNOR U18438 ( .A(n18160), .B(n18158), .Z(n18375) );
  AND U18439 ( .A(n18376), .B(n18377), .Z(n18158) );
  NANDN U18440 ( .A(n18378), .B(n18379), .Z(n18377) );
  OR U18441 ( .A(n18380), .B(n18381), .Z(n18379) );
  NAND U18442 ( .A(n18381), .B(n18380), .Z(n18376) );
  ANDN U18443 ( .B(B[227]), .A(n63), .Z(n18160) );
  XNOR U18444 ( .A(n18168), .B(n18382), .Z(n18161) );
  XNOR U18445 ( .A(n18167), .B(n18165), .Z(n18382) );
  AND U18446 ( .A(n18383), .B(n18384), .Z(n18165) );
  NANDN U18447 ( .A(n18385), .B(n18386), .Z(n18384) );
  NANDN U18448 ( .A(n18387), .B(n18388), .Z(n18386) );
  NANDN U18449 ( .A(n18388), .B(n18387), .Z(n18383) );
  ANDN U18450 ( .B(B[228]), .A(n64), .Z(n18167) );
  XNOR U18451 ( .A(n18175), .B(n18389), .Z(n18168) );
  XNOR U18452 ( .A(n18174), .B(n18172), .Z(n18389) );
  AND U18453 ( .A(n18390), .B(n18391), .Z(n18172) );
  NANDN U18454 ( .A(n18392), .B(n18393), .Z(n18391) );
  OR U18455 ( .A(n18394), .B(n18395), .Z(n18393) );
  NAND U18456 ( .A(n18395), .B(n18394), .Z(n18390) );
  ANDN U18457 ( .B(B[229]), .A(n65), .Z(n18174) );
  XNOR U18458 ( .A(n18182), .B(n18396), .Z(n18175) );
  XNOR U18459 ( .A(n18181), .B(n18179), .Z(n18396) );
  AND U18460 ( .A(n18397), .B(n18398), .Z(n18179) );
  NANDN U18461 ( .A(n18399), .B(n18400), .Z(n18398) );
  NANDN U18462 ( .A(n18401), .B(n18402), .Z(n18400) );
  NANDN U18463 ( .A(n18402), .B(n18401), .Z(n18397) );
  ANDN U18464 ( .B(B[230]), .A(n66), .Z(n18181) );
  XNOR U18465 ( .A(n18189), .B(n18403), .Z(n18182) );
  XNOR U18466 ( .A(n18188), .B(n18186), .Z(n18403) );
  AND U18467 ( .A(n18404), .B(n18405), .Z(n18186) );
  NANDN U18468 ( .A(n18406), .B(n18407), .Z(n18405) );
  OR U18469 ( .A(n18408), .B(n18409), .Z(n18407) );
  NAND U18470 ( .A(n18409), .B(n18408), .Z(n18404) );
  ANDN U18471 ( .B(B[231]), .A(n67), .Z(n18188) );
  XNOR U18472 ( .A(n18196), .B(n18410), .Z(n18189) );
  XNOR U18473 ( .A(n18195), .B(n18193), .Z(n18410) );
  AND U18474 ( .A(n18411), .B(n18412), .Z(n18193) );
  NANDN U18475 ( .A(n18413), .B(n18414), .Z(n18412) );
  NANDN U18476 ( .A(n18415), .B(n18416), .Z(n18414) );
  NANDN U18477 ( .A(n18416), .B(n18415), .Z(n18411) );
  ANDN U18478 ( .B(B[232]), .A(n68), .Z(n18195) );
  XNOR U18479 ( .A(n18203), .B(n18417), .Z(n18196) );
  XNOR U18480 ( .A(n18202), .B(n18200), .Z(n18417) );
  AND U18481 ( .A(n18418), .B(n18419), .Z(n18200) );
  NANDN U18482 ( .A(n18420), .B(n18421), .Z(n18419) );
  OR U18483 ( .A(n18422), .B(n18423), .Z(n18421) );
  NAND U18484 ( .A(n18423), .B(n18422), .Z(n18418) );
  ANDN U18485 ( .B(B[233]), .A(n69), .Z(n18202) );
  XNOR U18486 ( .A(n18210), .B(n18424), .Z(n18203) );
  XNOR U18487 ( .A(n18209), .B(n18207), .Z(n18424) );
  AND U18488 ( .A(n18425), .B(n18426), .Z(n18207) );
  NANDN U18489 ( .A(n18427), .B(n18428), .Z(n18426) );
  NANDN U18490 ( .A(n18429), .B(n18430), .Z(n18428) );
  NANDN U18491 ( .A(n18430), .B(n18429), .Z(n18425) );
  ANDN U18492 ( .B(B[234]), .A(n70), .Z(n18209) );
  XNOR U18493 ( .A(n18217), .B(n18431), .Z(n18210) );
  XNOR U18494 ( .A(n18216), .B(n18214), .Z(n18431) );
  AND U18495 ( .A(n18432), .B(n18433), .Z(n18214) );
  NANDN U18496 ( .A(n18434), .B(n18435), .Z(n18433) );
  OR U18497 ( .A(n18436), .B(n18437), .Z(n18435) );
  NAND U18498 ( .A(n18437), .B(n18436), .Z(n18432) );
  ANDN U18499 ( .B(B[235]), .A(n71), .Z(n18216) );
  XNOR U18500 ( .A(n18224), .B(n18438), .Z(n18217) );
  XNOR U18501 ( .A(n18223), .B(n18221), .Z(n18438) );
  AND U18502 ( .A(n18439), .B(n18440), .Z(n18221) );
  NANDN U18503 ( .A(n18441), .B(n18442), .Z(n18440) );
  NANDN U18504 ( .A(n18443), .B(n18444), .Z(n18442) );
  NANDN U18505 ( .A(n18444), .B(n18443), .Z(n18439) );
  ANDN U18506 ( .B(B[236]), .A(n72), .Z(n18223) );
  XNOR U18507 ( .A(n18231), .B(n18445), .Z(n18224) );
  XNOR U18508 ( .A(n18230), .B(n18228), .Z(n18445) );
  AND U18509 ( .A(n18446), .B(n18447), .Z(n18228) );
  NANDN U18510 ( .A(n18448), .B(n18449), .Z(n18447) );
  OR U18511 ( .A(n18450), .B(n18451), .Z(n18449) );
  NAND U18512 ( .A(n18451), .B(n18450), .Z(n18446) );
  ANDN U18513 ( .B(B[237]), .A(n73), .Z(n18230) );
  XNOR U18514 ( .A(n18238), .B(n18452), .Z(n18231) );
  XNOR U18515 ( .A(n18237), .B(n18235), .Z(n18452) );
  AND U18516 ( .A(n18453), .B(n18454), .Z(n18235) );
  NANDN U18517 ( .A(n18455), .B(n18456), .Z(n18454) );
  NANDN U18518 ( .A(n18457), .B(n18458), .Z(n18456) );
  NANDN U18519 ( .A(n18458), .B(n18457), .Z(n18453) );
  ANDN U18520 ( .B(B[238]), .A(n74), .Z(n18237) );
  XNOR U18521 ( .A(n18245), .B(n18459), .Z(n18238) );
  XNOR U18522 ( .A(n18244), .B(n18242), .Z(n18459) );
  AND U18523 ( .A(n18460), .B(n18461), .Z(n18242) );
  NANDN U18524 ( .A(n18462), .B(n18463), .Z(n18461) );
  OR U18525 ( .A(n18464), .B(n18465), .Z(n18463) );
  NAND U18526 ( .A(n18465), .B(n18464), .Z(n18460) );
  ANDN U18527 ( .B(B[239]), .A(n75), .Z(n18244) );
  XNOR U18528 ( .A(n18252), .B(n18466), .Z(n18245) );
  XNOR U18529 ( .A(n18251), .B(n18249), .Z(n18466) );
  AND U18530 ( .A(n18467), .B(n18468), .Z(n18249) );
  NANDN U18531 ( .A(n18469), .B(n18470), .Z(n18468) );
  NANDN U18532 ( .A(n18471), .B(n18472), .Z(n18470) );
  NANDN U18533 ( .A(n18472), .B(n18471), .Z(n18467) );
  ANDN U18534 ( .B(B[240]), .A(n76), .Z(n18251) );
  XNOR U18535 ( .A(n18259), .B(n18473), .Z(n18252) );
  XNOR U18536 ( .A(n18258), .B(n18256), .Z(n18473) );
  AND U18537 ( .A(n18474), .B(n18475), .Z(n18256) );
  NANDN U18538 ( .A(n18476), .B(n18477), .Z(n18475) );
  OR U18539 ( .A(n18478), .B(n18479), .Z(n18477) );
  NAND U18540 ( .A(n18479), .B(n18478), .Z(n18474) );
  ANDN U18541 ( .B(B[241]), .A(n77), .Z(n18258) );
  XNOR U18542 ( .A(n18266), .B(n18480), .Z(n18259) );
  XNOR U18543 ( .A(n18265), .B(n18263), .Z(n18480) );
  AND U18544 ( .A(n18481), .B(n18482), .Z(n18263) );
  NANDN U18545 ( .A(n18483), .B(n18484), .Z(n18482) );
  NANDN U18546 ( .A(n18485), .B(n18486), .Z(n18484) );
  NANDN U18547 ( .A(n18486), .B(n18485), .Z(n18481) );
  ANDN U18548 ( .B(B[242]), .A(n78), .Z(n18265) );
  XNOR U18549 ( .A(n18273), .B(n18487), .Z(n18266) );
  XNOR U18550 ( .A(n18272), .B(n18270), .Z(n18487) );
  AND U18551 ( .A(n18488), .B(n18489), .Z(n18270) );
  NANDN U18552 ( .A(n18490), .B(n18491), .Z(n18489) );
  OR U18553 ( .A(n18492), .B(n18493), .Z(n18491) );
  NAND U18554 ( .A(n18493), .B(n18492), .Z(n18488) );
  ANDN U18555 ( .B(B[243]), .A(n79), .Z(n18272) );
  XNOR U18556 ( .A(n18280), .B(n18494), .Z(n18273) );
  XNOR U18557 ( .A(n18279), .B(n18277), .Z(n18494) );
  AND U18558 ( .A(n18495), .B(n18496), .Z(n18277) );
  NANDN U18559 ( .A(n18497), .B(n18498), .Z(n18496) );
  NANDN U18560 ( .A(n18499), .B(n18500), .Z(n18498) );
  NANDN U18561 ( .A(n18500), .B(n18499), .Z(n18495) );
  ANDN U18562 ( .B(B[244]), .A(n80), .Z(n18279) );
  XNOR U18563 ( .A(n18287), .B(n18501), .Z(n18280) );
  XNOR U18564 ( .A(n18286), .B(n18284), .Z(n18501) );
  AND U18565 ( .A(n18502), .B(n18503), .Z(n18284) );
  NANDN U18566 ( .A(n18504), .B(n18505), .Z(n18503) );
  OR U18567 ( .A(n18506), .B(n18507), .Z(n18505) );
  NAND U18568 ( .A(n18507), .B(n18506), .Z(n18502) );
  ANDN U18569 ( .B(B[245]), .A(n81), .Z(n18286) );
  XNOR U18570 ( .A(n18294), .B(n18508), .Z(n18287) );
  XNOR U18571 ( .A(n18293), .B(n18291), .Z(n18508) );
  AND U18572 ( .A(n18509), .B(n18510), .Z(n18291) );
  NANDN U18573 ( .A(n18511), .B(n18512), .Z(n18510) );
  NAND U18574 ( .A(n18513), .B(n18514), .Z(n18512) );
  ANDN U18575 ( .B(B[246]), .A(n82), .Z(n18293) );
  XOR U18576 ( .A(n18300), .B(n18515), .Z(n18294) );
  XNOR U18577 ( .A(n18298), .B(n18301), .Z(n18515) );
  NAND U18578 ( .A(A[2]), .B(B[247]), .Z(n18301) );
  NANDN U18579 ( .A(n18516), .B(n18517), .Z(n18298) );
  AND U18580 ( .A(A[0]), .B(B[248]), .Z(n18517) );
  XNOR U18581 ( .A(n18303), .B(n18518), .Z(n18300) );
  NAND U18582 ( .A(A[0]), .B(B[249]), .Z(n18518) );
  NAND U18583 ( .A(B[248]), .B(A[1]), .Z(n18303) );
  NAND U18584 ( .A(n18519), .B(n18520), .Z(n298) );
  NANDN U18585 ( .A(n18521), .B(n18522), .Z(n18520) );
  OR U18586 ( .A(n18523), .B(n18524), .Z(n18522) );
  NAND U18587 ( .A(n18524), .B(n18523), .Z(n18519) );
  XOR U18588 ( .A(n300), .B(n299), .Z(\A1[246] ) );
  XOR U18589 ( .A(n18524), .B(n18525), .Z(n299) );
  XNOR U18590 ( .A(n18523), .B(n18521), .Z(n18525) );
  AND U18591 ( .A(n18526), .B(n18527), .Z(n18521) );
  NANDN U18592 ( .A(n18528), .B(n18529), .Z(n18527) );
  NANDN U18593 ( .A(n18530), .B(n18531), .Z(n18529) );
  NANDN U18594 ( .A(n18531), .B(n18530), .Z(n18526) );
  ANDN U18595 ( .B(B[217]), .A(n54), .Z(n18523) );
  XNOR U18596 ( .A(n18318), .B(n18532), .Z(n18524) );
  XNOR U18597 ( .A(n18317), .B(n18315), .Z(n18532) );
  AND U18598 ( .A(n18533), .B(n18534), .Z(n18315) );
  NANDN U18599 ( .A(n18535), .B(n18536), .Z(n18534) );
  OR U18600 ( .A(n18537), .B(n18538), .Z(n18536) );
  NAND U18601 ( .A(n18538), .B(n18537), .Z(n18533) );
  ANDN U18602 ( .B(B[218]), .A(n55), .Z(n18317) );
  XNOR U18603 ( .A(n18325), .B(n18539), .Z(n18318) );
  XNOR U18604 ( .A(n18324), .B(n18322), .Z(n18539) );
  AND U18605 ( .A(n18540), .B(n18541), .Z(n18322) );
  NANDN U18606 ( .A(n18542), .B(n18543), .Z(n18541) );
  NANDN U18607 ( .A(n18544), .B(n18545), .Z(n18543) );
  NANDN U18608 ( .A(n18545), .B(n18544), .Z(n18540) );
  ANDN U18609 ( .B(B[219]), .A(n56), .Z(n18324) );
  XNOR U18610 ( .A(n18332), .B(n18546), .Z(n18325) );
  XNOR U18611 ( .A(n18331), .B(n18329), .Z(n18546) );
  AND U18612 ( .A(n18547), .B(n18548), .Z(n18329) );
  NANDN U18613 ( .A(n18549), .B(n18550), .Z(n18548) );
  OR U18614 ( .A(n18551), .B(n18552), .Z(n18550) );
  NAND U18615 ( .A(n18552), .B(n18551), .Z(n18547) );
  ANDN U18616 ( .B(B[220]), .A(n57), .Z(n18331) );
  XNOR U18617 ( .A(n18339), .B(n18553), .Z(n18332) );
  XNOR U18618 ( .A(n18338), .B(n18336), .Z(n18553) );
  AND U18619 ( .A(n18554), .B(n18555), .Z(n18336) );
  NANDN U18620 ( .A(n18556), .B(n18557), .Z(n18555) );
  NANDN U18621 ( .A(n18558), .B(n18559), .Z(n18557) );
  NANDN U18622 ( .A(n18559), .B(n18558), .Z(n18554) );
  ANDN U18623 ( .B(B[221]), .A(n58), .Z(n18338) );
  XNOR U18624 ( .A(n18346), .B(n18560), .Z(n18339) );
  XNOR U18625 ( .A(n18345), .B(n18343), .Z(n18560) );
  AND U18626 ( .A(n18561), .B(n18562), .Z(n18343) );
  NANDN U18627 ( .A(n18563), .B(n18564), .Z(n18562) );
  OR U18628 ( .A(n18565), .B(n18566), .Z(n18564) );
  NAND U18629 ( .A(n18566), .B(n18565), .Z(n18561) );
  ANDN U18630 ( .B(B[222]), .A(n59), .Z(n18345) );
  XNOR U18631 ( .A(n18353), .B(n18567), .Z(n18346) );
  XNOR U18632 ( .A(n18352), .B(n18350), .Z(n18567) );
  AND U18633 ( .A(n18568), .B(n18569), .Z(n18350) );
  NANDN U18634 ( .A(n18570), .B(n18571), .Z(n18569) );
  NANDN U18635 ( .A(n18572), .B(n18573), .Z(n18571) );
  NANDN U18636 ( .A(n18573), .B(n18572), .Z(n18568) );
  ANDN U18637 ( .B(B[223]), .A(n60), .Z(n18352) );
  XNOR U18638 ( .A(n18360), .B(n18574), .Z(n18353) );
  XNOR U18639 ( .A(n18359), .B(n18357), .Z(n18574) );
  AND U18640 ( .A(n18575), .B(n18576), .Z(n18357) );
  NANDN U18641 ( .A(n18577), .B(n18578), .Z(n18576) );
  OR U18642 ( .A(n18579), .B(n18580), .Z(n18578) );
  NAND U18643 ( .A(n18580), .B(n18579), .Z(n18575) );
  ANDN U18644 ( .B(B[224]), .A(n61), .Z(n18359) );
  XNOR U18645 ( .A(n18367), .B(n18581), .Z(n18360) );
  XNOR U18646 ( .A(n18366), .B(n18364), .Z(n18581) );
  AND U18647 ( .A(n18582), .B(n18583), .Z(n18364) );
  NANDN U18648 ( .A(n18584), .B(n18585), .Z(n18583) );
  NANDN U18649 ( .A(n18586), .B(n18587), .Z(n18585) );
  NANDN U18650 ( .A(n18587), .B(n18586), .Z(n18582) );
  ANDN U18651 ( .B(B[225]), .A(n62), .Z(n18366) );
  XNOR U18652 ( .A(n18374), .B(n18588), .Z(n18367) );
  XNOR U18653 ( .A(n18373), .B(n18371), .Z(n18588) );
  AND U18654 ( .A(n18589), .B(n18590), .Z(n18371) );
  NANDN U18655 ( .A(n18591), .B(n18592), .Z(n18590) );
  OR U18656 ( .A(n18593), .B(n18594), .Z(n18592) );
  NAND U18657 ( .A(n18594), .B(n18593), .Z(n18589) );
  ANDN U18658 ( .B(B[226]), .A(n63), .Z(n18373) );
  XNOR U18659 ( .A(n18381), .B(n18595), .Z(n18374) );
  XNOR U18660 ( .A(n18380), .B(n18378), .Z(n18595) );
  AND U18661 ( .A(n18596), .B(n18597), .Z(n18378) );
  NANDN U18662 ( .A(n18598), .B(n18599), .Z(n18597) );
  NANDN U18663 ( .A(n18600), .B(n18601), .Z(n18599) );
  NANDN U18664 ( .A(n18601), .B(n18600), .Z(n18596) );
  ANDN U18665 ( .B(B[227]), .A(n64), .Z(n18380) );
  XNOR U18666 ( .A(n18388), .B(n18602), .Z(n18381) );
  XNOR U18667 ( .A(n18387), .B(n18385), .Z(n18602) );
  AND U18668 ( .A(n18603), .B(n18604), .Z(n18385) );
  NANDN U18669 ( .A(n18605), .B(n18606), .Z(n18604) );
  OR U18670 ( .A(n18607), .B(n18608), .Z(n18606) );
  NAND U18671 ( .A(n18608), .B(n18607), .Z(n18603) );
  ANDN U18672 ( .B(B[228]), .A(n65), .Z(n18387) );
  XNOR U18673 ( .A(n18395), .B(n18609), .Z(n18388) );
  XNOR U18674 ( .A(n18394), .B(n18392), .Z(n18609) );
  AND U18675 ( .A(n18610), .B(n18611), .Z(n18392) );
  NANDN U18676 ( .A(n18612), .B(n18613), .Z(n18611) );
  NANDN U18677 ( .A(n18614), .B(n18615), .Z(n18613) );
  NANDN U18678 ( .A(n18615), .B(n18614), .Z(n18610) );
  ANDN U18679 ( .B(B[229]), .A(n66), .Z(n18394) );
  XNOR U18680 ( .A(n18402), .B(n18616), .Z(n18395) );
  XNOR U18681 ( .A(n18401), .B(n18399), .Z(n18616) );
  AND U18682 ( .A(n18617), .B(n18618), .Z(n18399) );
  NANDN U18683 ( .A(n18619), .B(n18620), .Z(n18618) );
  OR U18684 ( .A(n18621), .B(n18622), .Z(n18620) );
  NAND U18685 ( .A(n18622), .B(n18621), .Z(n18617) );
  ANDN U18686 ( .B(B[230]), .A(n67), .Z(n18401) );
  XNOR U18687 ( .A(n18409), .B(n18623), .Z(n18402) );
  XNOR U18688 ( .A(n18408), .B(n18406), .Z(n18623) );
  AND U18689 ( .A(n18624), .B(n18625), .Z(n18406) );
  NANDN U18690 ( .A(n18626), .B(n18627), .Z(n18625) );
  NANDN U18691 ( .A(n18628), .B(n18629), .Z(n18627) );
  NANDN U18692 ( .A(n18629), .B(n18628), .Z(n18624) );
  ANDN U18693 ( .B(B[231]), .A(n68), .Z(n18408) );
  XNOR U18694 ( .A(n18416), .B(n18630), .Z(n18409) );
  XNOR U18695 ( .A(n18415), .B(n18413), .Z(n18630) );
  AND U18696 ( .A(n18631), .B(n18632), .Z(n18413) );
  NANDN U18697 ( .A(n18633), .B(n18634), .Z(n18632) );
  OR U18698 ( .A(n18635), .B(n18636), .Z(n18634) );
  NAND U18699 ( .A(n18636), .B(n18635), .Z(n18631) );
  ANDN U18700 ( .B(B[232]), .A(n69), .Z(n18415) );
  XNOR U18701 ( .A(n18423), .B(n18637), .Z(n18416) );
  XNOR U18702 ( .A(n18422), .B(n18420), .Z(n18637) );
  AND U18703 ( .A(n18638), .B(n18639), .Z(n18420) );
  NANDN U18704 ( .A(n18640), .B(n18641), .Z(n18639) );
  NANDN U18705 ( .A(n18642), .B(n18643), .Z(n18641) );
  NANDN U18706 ( .A(n18643), .B(n18642), .Z(n18638) );
  ANDN U18707 ( .B(B[233]), .A(n70), .Z(n18422) );
  XNOR U18708 ( .A(n18430), .B(n18644), .Z(n18423) );
  XNOR U18709 ( .A(n18429), .B(n18427), .Z(n18644) );
  AND U18710 ( .A(n18645), .B(n18646), .Z(n18427) );
  NANDN U18711 ( .A(n18647), .B(n18648), .Z(n18646) );
  OR U18712 ( .A(n18649), .B(n18650), .Z(n18648) );
  NAND U18713 ( .A(n18650), .B(n18649), .Z(n18645) );
  ANDN U18714 ( .B(B[234]), .A(n71), .Z(n18429) );
  XNOR U18715 ( .A(n18437), .B(n18651), .Z(n18430) );
  XNOR U18716 ( .A(n18436), .B(n18434), .Z(n18651) );
  AND U18717 ( .A(n18652), .B(n18653), .Z(n18434) );
  NANDN U18718 ( .A(n18654), .B(n18655), .Z(n18653) );
  NANDN U18719 ( .A(n18656), .B(n18657), .Z(n18655) );
  NANDN U18720 ( .A(n18657), .B(n18656), .Z(n18652) );
  ANDN U18721 ( .B(B[235]), .A(n72), .Z(n18436) );
  XNOR U18722 ( .A(n18444), .B(n18658), .Z(n18437) );
  XNOR U18723 ( .A(n18443), .B(n18441), .Z(n18658) );
  AND U18724 ( .A(n18659), .B(n18660), .Z(n18441) );
  NANDN U18725 ( .A(n18661), .B(n18662), .Z(n18660) );
  OR U18726 ( .A(n18663), .B(n18664), .Z(n18662) );
  NAND U18727 ( .A(n18664), .B(n18663), .Z(n18659) );
  ANDN U18728 ( .B(B[236]), .A(n73), .Z(n18443) );
  XNOR U18729 ( .A(n18451), .B(n18665), .Z(n18444) );
  XNOR U18730 ( .A(n18450), .B(n18448), .Z(n18665) );
  AND U18731 ( .A(n18666), .B(n18667), .Z(n18448) );
  NANDN U18732 ( .A(n18668), .B(n18669), .Z(n18667) );
  NANDN U18733 ( .A(n18670), .B(n18671), .Z(n18669) );
  NANDN U18734 ( .A(n18671), .B(n18670), .Z(n18666) );
  ANDN U18735 ( .B(B[237]), .A(n74), .Z(n18450) );
  XNOR U18736 ( .A(n18458), .B(n18672), .Z(n18451) );
  XNOR U18737 ( .A(n18457), .B(n18455), .Z(n18672) );
  AND U18738 ( .A(n18673), .B(n18674), .Z(n18455) );
  NANDN U18739 ( .A(n18675), .B(n18676), .Z(n18674) );
  OR U18740 ( .A(n18677), .B(n18678), .Z(n18676) );
  NAND U18741 ( .A(n18678), .B(n18677), .Z(n18673) );
  ANDN U18742 ( .B(B[238]), .A(n75), .Z(n18457) );
  XNOR U18743 ( .A(n18465), .B(n18679), .Z(n18458) );
  XNOR U18744 ( .A(n18464), .B(n18462), .Z(n18679) );
  AND U18745 ( .A(n18680), .B(n18681), .Z(n18462) );
  NANDN U18746 ( .A(n18682), .B(n18683), .Z(n18681) );
  NANDN U18747 ( .A(n18684), .B(n18685), .Z(n18683) );
  NANDN U18748 ( .A(n18685), .B(n18684), .Z(n18680) );
  ANDN U18749 ( .B(B[239]), .A(n76), .Z(n18464) );
  XNOR U18750 ( .A(n18472), .B(n18686), .Z(n18465) );
  XNOR U18751 ( .A(n18471), .B(n18469), .Z(n18686) );
  AND U18752 ( .A(n18687), .B(n18688), .Z(n18469) );
  NANDN U18753 ( .A(n18689), .B(n18690), .Z(n18688) );
  OR U18754 ( .A(n18691), .B(n18692), .Z(n18690) );
  NAND U18755 ( .A(n18692), .B(n18691), .Z(n18687) );
  ANDN U18756 ( .B(B[240]), .A(n77), .Z(n18471) );
  XNOR U18757 ( .A(n18479), .B(n18693), .Z(n18472) );
  XNOR U18758 ( .A(n18478), .B(n18476), .Z(n18693) );
  AND U18759 ( .A(n18694), .B(n18695), .Z(n18476) );
  NANDN U18760 ( .A(n18696), .B(n18697), .Z(n18695) );
  NANDN U18761 ( .A(n18698), .B(n18699), .Z(n18697) );
  NANDN U18762 ( .A(n18699), .B(n18698), .Z(n18694) );
  ANDN U18763 ( .B(B[241]), .A(n78), .Z(n18478) );
  XNOR U18764 ( .A(n18486), .B(n18700), .Z(n18479) );
  XNOR U18765 ( .A(n18485), .B(n18483), .Z(n18700) );
  AND U18766 ( .A(n18701), .B(n18702), .Z(n18483) );
  NANDN U18767 ( .A(n18703), .B(n18704), .Z(n18702) );
  OR U18768 ( .A(n18705), .B(n18706), .Z(n18704) );
  NAND U18769 ( .A(n18706), .B(n18705), .Z(n18701) );
  ANDN U18770 ( .B(B[242]), .A(n79), .Z(n18485) );
  XNOR U18771 ( .A(n18493), .B(n18707), .Z(n18486) );
  XNOR U18772 ( .A(n18492), .B(n18490), .Z(n18707) );
  AND U18773 ( .A(n18708), .B(n18709), .Z(n18490) );
  NANDN U18774 ( .A(n18710), .B(n18711), .Z(n18709) );
  NANDN U18775 ( .A(n18712), .B(n18713), .Z(n18711) );
  NANDN U18776 ( .A(n18713), .B(n18712), .Z(n18708) );
  ANDN U18777 ( .B(B[243]), .A(n80), .Z(n18492) );
  XNOR U18778 ( .A(n18500), .B(n18714), .Z(n18493) );
  XNOR U18779 ( .A(n18499), .B(n18497), .Z(n18714) );
  AND U18780 ( .A(n18715), .B(n18716), .Z(n18497) );
  NANDN U18781 ( .A(n18717), .B(n18718), .Z(n18716) );
  OR U18782 ( .A(n18719), .B(n18720), .Z(n18718) );
  NAND U18783 ( .A(n18720), .B(n18719), .Z(n18715) );
  ANDN U18784 ( .B(B[244]), .A(n81), .Z(n18499) );
  XNOR U18785 ( .A(n18507), .B(n18721), .Z(n18500) );
  XNOR U18786 ( .A(n18506), .B(n18504), .Z(n18721) );
  AND U18787 ( .A(n18722), .B(n18723), .Z(n18504) );
  NANDN U18788 ( .A(n18724), .B(n18725), .Z(n18723) );
  NAND U18789 ( .A(n18726), .B(n18727), .Z(n18725) );
  ANDN U18790 ( .B(B[245]), .A(n82), .Z(n18506) );
  XOR U18791 ( .A(n18513), .B(n18728), .Z(n18507) );
  XNOR U18792 ( .A(n18511), .B(n18514), .Z(n18728) );
  NAND U18793 ( .A(A[2]), .B(B[246]), .Z(n18514) );
  NANDN U18794 ( .A(n18729), .B(n18730), .Z(n18511) );
  AND U18795 ( .A(A[0]), .B(B[247]), .Z(n18730) );
  XNOR U18796 ( .A(n18516), .B(n18731), .Z(n18513) );
  NAND U18797 ( .A(A[0]), .B(B[248]), .Z(n18731) );
  NAND U18798 ( .A(B[247]), .B(A[1]), .Z(n18516) );
  NAND U18799 ( .A(n18732), .B(n18733), .Z(n300) );
  NANDN U18800 ( .A(n18734), .B(n18735), .Z(n18733) );
  OR U18801 ( .A(n18736), .B(n18737), .Z(n18735) );
  NAND U18802 ( .A(n18737), .B(n18736), .Z(n18732) );
  XOR U18803 ( .A(n302), .B(n301), .Z(\A1[245] ) );
  XOR U18804 ( .A(n18737), .B(n18738), .Z(n301) );
  XNOR U18805 ( .A(n18736), .B(n18734), .Z(n18738) );
  AND U18806 ( .A(n18739), .B(n18740), .Z(n18734) );
  NANDN U18807 ( .A(n18741), .B(n18742), .Z(n18740) );
  NANDN U18808 ( .A(n18743), .B(n18744), .Z(n18742) );
  NANDN U18809 ( .A(n18744), .B(n18743), .Z(n18739) );
  ANDN U18810 ( .B(B[216]), .A(n54), .Z(n18736) );
  XNOR U18811 ( .A(n18531), .B(n18745), .Z(n18737) );
  XNOR U18812 ( .A(n18530), .B(n18528), .Z(n18745) );
  AND U18813 ( .A(n18746), .B(n18747), .Z(n18528) );
  NANDN U18814 ( .A(n18748), .B(n18749), .Z(n18747) );
  OR U18815 ( .A(n18750), .B(n18751), .Z(n18749) );
  NAND U18816 ( .A(n18751), .B(n18750), .Z(n18746) );
  ANDN U18817 ( .B(B[217]), .A(n55), .Z(n18530) );
  XNOR U18818 ( .A(n18538), .B(n18752), .Z(n18531) );
  XNOR U18819 ( .A(n18537), .B(n18535), .Z(n18752) );
  AND U18820 ( .A(n18753), .B(n18754), .Z(n18535) );
  NANDN U18821 ( .A(n18755), .B(n18756), .Z(n18754) );
  NANDN U18822 ( .A(n18757), .B(n18758), .Z(n18756) );
  NANDN U18823 ( .A(n18758), .B(n18757), .Z(n18753) );
  ANDN U18824 ( .B(B[218]), .A(n56), .Z(n18537) );
  XNOR U18825 ( .A(n18545), .B(n18759), .Z(n18538) );
  XNOR U18826 ( .A(n18544), .B(n18542), .Z(n18759) );
  AND U18827 ( .A(n18760), .B(n18761), .Z(n18542) );
  NANDN U18828 ( .A(n18762), .B(n18763), .Z(n18761) );
  OR U18829 ( .A(n18764), .B(n18765), .Z(n18763) );
  NAND U18830 ( .A(n18765), .B(n18764), .Z(n18760) );
  ANDN U18831 ( .B(B[219]), .A(n57), .Z(n18544) );
  XNOR U18832 ( .A(n18552), .B(n18766), .Z(n18545) );
  XNOR U18833 ( .A(n18551), .B(n18549), .Z(n18766) );
  AND U18834 ( .A(n18767), .B(n18768), .Z(n18549) );
  NANDN U18835 ( .A(n18769), .B(n18770), .Z(n18768) );
  NANDN U18836 ( .A(n18771), .B(n18772), .Z(n18770) );
  NANDN U18837 ( .A(n18772), .B(n18771), .Z(n18767) );
  ANDN U18838 ( .B(B[220]), .A(n58), .Z(n18551) );
  XNOR U18839 ( .A(n18559), .B(n18773), .Z(n18552) );
  XNOR U18840 ( .A(n18558), .B(n18556), .Z(n18773) );
  AND U18841 ( .A(n18774), .B(n18775), .Z(n18556) );
  NANDN U18842 ( .A(n18776), .B(n18777), .Z(n18775) );
  OR U18843 ( .A(n18778), .B(n18779), .Z(n18777) );
  NAND U18844 ( .A(n18779), .B(n18778), .Z(n18774) );
  ANDN U18845 ( .B(B[221]), .A(n59), .Z(n18558) );
  XNOR U18846 ( .A(n18566), .B(n18780), .Z(n18559) );
  XNOR U18847 ( .A(n18565), .B(n18563), .Z(n18780) );
  AND U18848 ( .A(n18781), .B(n18782), .Z(n18563) );
  NANDN U18849 ( .A(n18783), .B(n18784), .Z(n18782) );
  NANDN U18850 ( .A(n18785), .B(n18786), .Z(n18784) );
  NANDN U18851 ( .A(n18786), .B(n18785), .Z(n18781) );
  ANDN U18852 ( .B(B[222]), .A(n60), .Z(n18565) );
  XNOR U18853 ( .A(n18573), .B(n18787), .Z(n18566) );
  XNOR U18854 ( .A(n18572), .B(n18570), .Z(n18787) );
  AND U18855 ( .A(n18788), .B(n18789), .Z(n18570) );
  NANDN U18856 ( .A(n18790), .B(n18791), .Z(n18789) );
  OR U18857 ( .A(n18792), .B(n18793), .Z(n18791) );
  NAND U18858 ( .A(n18793), .B(n18792), .Z(n18788) );
  ANDN U18859 ( .B(B[223]), .A(n61), .Z(n18572) );
  XNOR U18860 ( .A(n18580), .B(n18794), .Z(n18573) );
  XNOR U18861 ( .A(n18579), .B(n18577), .Z(n18794) );
  AND U18862 ( .A(n18795), .B(n18796), .Z(n18577) );
  NANDN U18863 ( .A(n18797), .B(n18798), .Z(n18796) );
  NANDN U18864 ( .A(n18799), .B(n18800), .Z(n18798) );
  NANDN U18865 ( .A(n18800), .B(n18799), .Z(n18795) );
  ANDN U18866 ( .B(B[224]), .A(n62), .Z(n18579) );
  XNOR U18867 ( .A(n18587), .B(n18801), .Z(n18580) );
  XNOR U18868 ( .A(n18586), .B(n18584), .Z(n18801) );
  AND U18869 ( .A(n18802), .B(n18803), .Z(n18584) );
  NANDN U18870 ( .A(n18804), .B(n18805), .Z(n18803) );
  OR U18871 ( .A(n18806), .B(n18807), .Z(n18805) );
  NAND U18872 ( .A(n18807), .B(n18806), .Z(n18802) );
  ANDN U18873 ( .B(B[225]), .A(n63), .Z(n18586) );
  XNOR U18874 ( .A(n18594), .B(n18808), .Z(n18587) );
  XNOR U18875 ( .A(n18593), .B(n18591), .Z(n18808) );
  AND U18876 ( .A(n18809), .B(n18810), .Z(n18591) );
  NANDN U18877 ( .A(n18811), .B(n18812), .Z(n18810) );
  NANDN U18878 ( .A(n18813), .B(n18814), .Z(n18812) );
  NANDN U18879 ( .A(n18814), .B(n18813), .Z(n18809) );
  ANDN U18880 ( .B(B[226]), .A(n64), .Z(n18593) );
  XNOR U18881 ( .A(n18601), .B(n18815), .Z(n18594) );
  XNOR U18882 ( .A(n18600), .B(n18598), .Z(n18815) );
  AND U18883 ( .A(n18816), .B(n18817), .Z(n18598) );
  NANDN U18884 ( .A(n18818), .B(n18819), .Z(n18817) );
  OR U18885 ( .A(n18820), .B(n18821), .Z(n18819) );
  NAND U18886 ( .A(n18821), .B(n18820), .Z(n18816) );
  ANDN U18887 ( .B(B[227]), .A(n65), .Z(n18600) );
  XNOR U18888 ( .A(n18608), .B(n18822), .Z(n18601) );
  XNOR U18889 ( .A(n18607), .B(n18605), .Z(n18822) );
  AND U18890 ( .A(n18823), .B(n18824), .Z(n18605) );
  NANDN U18891 ( .A(n18825), .B(n18826), .Z(n18824) );
  NANDN U18892 ( .A(n18827), .B(n18828), .Z(n18826) );
  NANDN U18893 ( .A(n18828), .B(n18827), .Z(n18823) );
  ANDN U18894 ( .B(B[228]), .A(n66), .Z(n18607) );
  XNOR U18895 ( .A(n18615), .B(n18829), .Z(n18608) );
  XNOR U18896 ( .A(n18614), .B(n18612), .Z(n18829) );
  AND U18897 ( .A(n18830), .B(n18831), .Z(n18612) );
  NANDN U18898 ( .A(n18832), .B(n18833), .Z(n18831) );
  OR U18899 ( .A(n18834), .B(n18835), .Z(n18833) );
  NAND U18900 ( .A(n18835), .B(n18834), .Z(n18830) );
  ANDN U18901 ( .B(B[229]), .A(n67), .Z(n18614) );
  XNOR U18902 ( .A(n18622), .B(n18836), .Z(n18615) );
  XNOR U18903 ( .A(n18621), .B(n18619), .Z(n18836) );
  AND U18904 ( .A(n18837), .B(n18838), .Z(n18619) );
  NANDN U18905 ( .A(n18839), .B(n18840), .Z(n18838) );
  NANDN U18906 ( .A(n18841), .B(n18842), .Z(n18840) );
  NANDN U18907 ( .A(n18842), .B(n18841), .Z(n18837) );
  ANDN U18908 ( .B(B[230]), .A(n68), .Z(n18621) );
  XNOR U18909 ( .A(n18629), .B(n18843), .Z(n18622) );
  XNOR U18910 ( .A(n18628), .B(n18626), .Z(n18843) );
  AND U18911 ( .A(n18844), .B(n18845), .Z(n18626) );
  NANDN U18912 ( .A(n18846), .B(n18847), .Z(n18845) );
  OR U18913 ( .A(n18848), .B(n18849), .Z(n18847) );
  NAND U18914 ( .A(n18849), .B(n18848), .Z(n18844) );
  ANDN U18915 ( .B(B[231]), .A(n69), .Z(n18628) );
  XNOR U18916 ( .A(n18636), .B(n18850), .Z(n18629) );
  XNOR U18917 ( .A(n18635), .B(n18633), .Z(n18850) );
  AND U18918 ( .A(n18851), .B(n18852), .Z(n18633) );
  NANDN U18919 ( .A(n18853), .B(n18854), .Z(n18852) );
  NANDN U18920 ( .A(n18855), .B(n18856), .Z(n18854) );
  NANDN U18921 ( .A(n18856), .B(n18855), .Z(n18851) );
  ANDN U18922 ( .B(B[232]), .A(n70), .Z(n18635) );
  XNOR U18923 ( .A(n18643), .B(n18857), .Z(n18636) );
  XNOR U18924 ( .A(n18642), .B(n18640), .Z(n18857) );
  AND U18925 ( .A(n18858), .B(n18859), .Z(n18640) );
  NANDN U18926 ( .A(n18860), .B(n18861), .Z(n18859) );
  OR U18927 ( .A(n18862), .B(n18863), .Z(n18861) );
  NAND U18928 ( .A(n18863), .B(n18862), .Z(n18858) );
  ANDN U18929 ( .B(B[233]), .A(n71), .Z(n18642) );
  XNOR U18930 ( .A(n18650), .B(n18864), .Z(n18643) );
  XNOR U18931 ( .A(n18649), .B(n18647), .Z(n18864) );
  AND U18932 ( .A(n18865), .B(n18866), .Z(n18647) );
  NANDN U18933 ( .A(n18867), .B(n18868), .Z(n18866) );
  NANDN U18934 ( .A(n18869), .B(n18870), .Z(n18868) );
  NANDN U18935 ( .A(n18870), .B(n18869), .Z(n18865) );
  ANDN U18936 ( .B(B[234]), .A(n72), .Z(n18649) );
  XNOR U18937 ( .A(n18657), .B(n18871), .Z(n18650) );
  XNOR U18938 ( .A(n18656), .B(n18654), .Z(n18871) );
  AND U18939 ( .A(n18872), .B(n18873), .Z(n18654) );
  NANDN U18940 ( .A(n18874), .B(n18875), .Z(n18873) );
  OR U18941 ( .A(n18876), .B(n18877), .Z(n18875) );
  NAND U18942 ( .A(n18877), .B(n18876), .Z(n18872) );
  ANDN U18943 ( .B(B[235]), .A(n73), .Z(n18656) );
  XNOR U18944 ( .A(n18664), .B(n18878), .Z(n18657) );
  XNOR U18945 ( .A(n18663), .B(n18661), .Z(n18878) );
  AND U18946 ( .A(n18879), .B(n18880), .Z(n18661) );
  NANDN U18947 ( .A(n18881), .B(n18882), .Z(n18880) );
  NANDN U18948 ( .A(n18883), .B(n18884), .Z(n18882) );
  NANDN U18949 ( .A(n18884), .B(n18883), .Z(n18879) );
  ANDN U18950 ( .B(B[236]), .A(n74), .Z(n18663) );
  XNOR U18951 ( .A(n18671), .B(n18885), .Z(n18664) );
  XNOR U18952 ( .A(n18670), .B(n18668), .Z(n18885) );
  AND U18953 ( .A(n18886), .B(n18887), .Z(n18668) );
  NANDN U18954 ( .A(n18888), .B(n18889), .Z(n18887) );
  OR U18955 ( .A(n18890), .B(n18891), .Z(n18889) );
  NAND U18956 ( .A(n18891), .B(n18890), .Z(n18886) );
  ANDN U18957 ( .B(B[237]), .A(n75), .Z(n18670) );
  XNOR U18958 ( .A(n18678), .B(n18892), .Z(n18671) );
  XNOR U18959 ( .A(n18677), .B(n18675), .Z(n18892) );
  AND U18960 ( .A(n18893), .B(n18894), .Z(n18675) );
  NANDN U18961 ( .A(n18895), .B(n18896), .Z(n18894) );
  NANDN U18962 ( .A(n18897), .B(n18898), .Z(n18896) );
  NANDN U18963 ( .A(n18898), .B(n18897), .Z(n18893) );
  ANDN U18964 ( .B(B[238]), .A(n76), .Z(n18677) );
  XNOR U18965 ( .A(n18685), .B(n18899), .Z(n18678) );
  XNOR U18966 ( .A(n18684), .B(n18682), .Z(n18899) );
  AND U18967 ( .A(n18900), .B(n18901), .Z(n18682) );
  NANDN U18968 ( .A(n18902), .B(n18903), .Z(n18901) );
  OR U18969 ( .A(n18904), .B(n18905), .Z(n18903) );
  NAND U18970 ( .A(n18905), .B(n18904), .Z(n18900) );
  ANDN U18971 ( .B(B[239]), .A(n77), .Z(n18684) );
  XNOR U18972 ( .A(n18692), .B(n18906), .Z(n18685) );
  XNOR U18973 ( .A(n18691), .B(n18689), .Z(n18906) );
  AND U18974 ( .A(n18907), .B(n18908), .Z(n18689) );
  NANDN U18975 ( .A(n18909), .B(n18910), .Z(n18908) );
  NANDN U18976 ( .A(n18911), .B(n18912), .Z(n18910) );
  NANDN U18977 ( .A(n18912), .B(n18911), .Z(n18907) );
  ANDN U18978 ( .B(B[240]), .A(n78), .Z(n18691) );
  XNOR U18979 ( .A(n18699), .B(n18913), .Z(n18692) );
  XNOR U18980 ( .A(n18698), .B(n18696), .Z(n18913) );
  AND U18981 ( .A(n18914), .B(n18915), .Z(n18696) );
  NANDN U18982 ( .A(n18916), .B(n18917), .Z(n18915) );
  OR U18983 ( .A(n18918), .B(n18919), .Z(n18917) );
  NAND U18984 ( .A(n18919), .B(n18918), .Z(n18914) );
  ANDN U18985 ( .B(B[241]), .A(n79), .Z(n18698) );
  XNOR U18986 ( .A(n18706), .B(n18920), .Z(n18699) );
  XNOR U18987 ( .A(n18705), .B(n18703), .Z(n18920) );
  AND U18988 ( .A(n18921), .B(n18922), .Z(n18703) );
  NANDN U18989 ( .A(n18923), .B(n18924), .Z(n18922) );
  NANDN U18990 ( .A(n18925), .B(n18926), .Z(n18924) );
  NANDN U18991 ( .A(n18926), .B(n18925), .Z(n18921) );
  ANDN U18992 ( .B(B[242]), .A(n80), .Z(n18705) );
  XNOR U18993 ( .A(n18713), .B(n18927), .Z(n18706) );
  XNOR U18994 ( .A(n18712), .B(n18710), .Z(n18927) );
  AND U18995 ( .A(n18928), .B(n18929), .Z(n18710) );
  NANDN U18996 ( .A(n18930), .B(n18931), .Z(n18929) );
  OR U18997 ( .A(n18932), .B(n18933), .Z(n18931) );
  NAND U18998 ( .A(n18933), .B(n18932), .Z(n18928) );
  ANDN U18999 ( .B(B[243]), .A(n81), .Z(n18712) );
  XNOR U19000 ( .A(n18720), .B(n18934), .Z(n18713) );
  XNOR U19001 ( .A(n18719), .B(n18717), .Z(n18934) );
  AND U19002 ( .A(n18935), .B(n18936), .Z(n18717) );
  NANDN U19003 ( .A(n18937), .B(n18938), .Z(n18936) );
  NAND U19004 ( .A(n18939), .B(n18940), .Z(n18938) );
  ANDN U19005 ( .B(B[244]), .A(n82), .Z(n18719) );
  XOR U19006 ( .A(n18726), .B(n18941), .Z(n18720) );
  XNOR U19007 ( .A(n18724), .B(n18727), .Z(n18941) );
  NAND U19008 ( .A(A[2]), .B(B[245]), .Z(n18727) );
  NANDN U19009 ( .A(n18942), .B(n18943), .Z(n18724) );
  AND U19010 ( .A(A[0]), .B(B[246]), .Z(n18943) );
  XNOR U19011 ( .A(n18729), .B(n18944), .Z(n18726) );
  NAND U19012 ( .A(A[0]), .B(B[247]), .Z(n18944) );
  NAND U19013 ( .A(B[246]), .B(A[1]), .Z(n18729) );
  NAND U19014 ( .A(n18945), .B(n18946), .Z(n302) );
  NANDN U19015 ( .A(n18947), .B(n18948), .Z(n18946) );
  OR U19016 ( .A(n18949), .B(n18950), .Z(n18948) );
  NAND U19017 ( .A(n18950), .B(n18949), .Z(n18945) );
  XOR U19018 ( .A(n304), .B(n303), .Z(\A1[244] ) );
  XOR U19019 ( .A(n18950), .B(n18951), .Z(n303) );
  XNOR U19020 ( .A(n18949), .B(n18947), .Z(n18951) );
  AND U19021 ( .A(n18952), .B(n18953), .Z(n18947) );
  NANDN U19022 ( .A(n18954), .B(n18955), .Z(n18953) );
  NANDN U19023 ( .A(n18956), .B(n18957), .Z(n18955) );
  NANDN U19024 ( .A(n18957), .B(n18956), .Z(n18952) );
  ANDN U19025 ( .B(B[215]), .A(n54), .Z(n18949) );
  XNOR U19026 ( .A(n18744), .B(n18958), .Z(n18950) );
  XNOR U19027 ( .A(n18743), .B(n18741), .Z(n18958) );
  AND U19028 ( .A(n18959), .B(n18960), .Z(n18741) );
  NANDN U19029 ( .A(n18961), .B(n18962), .Z(n18960) );
  OR U19030 ( .A(n18963), .B(n18964), .Z(n18962) );
  NAND U19031 ( .A(n18964), .B(n18963), .Z(n18959) );
  ANDN U19032 ( .B(B[216]), .A(n55), .Z(n18743) );
  XNOR U19033 ( .A(n18751), .B(n18965), .Z(n18744) );
  XNOR U19034 ( .A(n18750), .B(n18748), .Z(n18965) );
  AND U19035 ( .A(n18966), .B(n18967), .Z(n18748) );
  NANDN U19036 ( .A(n18968), .B(n18969), .Z(n18967) );
  NANDN U19037 ( .A(n18970), .B(n18971), .Z(n18969) );
  NANDN U19038 ( .A(n18971), .B(n18970), .Z(n18966) );
  ANDN U19039 ( .B(B[217]), .A(n56), .Z(n18750) );
  XNOR U19040 ( .A(n18758), .B(n18972), .Z(n18751) );
  XNOR U19041 ( .A(n18757), .B(n18755), .Z(n18972) );
  AND U19042 ( .A(n18973), .B(n18974), .Z(n18755) );
  NANDN U19043 ( .A(n18975), .B(n18976), .Z(n18974) );
  OR U19044 ( .A(n18977), .B(n18978), .Z(n18976) );
  NAND U19045 ( .A(n18978), .B(n18977), .Z(n18973) );
  ANDN U19046 ( .B(B[218]), .A(n57), .Z(n18757) );
  XNOR U19047 ( .A(n18765), .B(n18979), .Z(n18758) );
  XNOR U19048 ( .A(n18764), .B(n18762), .Z(n18979) );
  AND U19049 ( .A(n18980), .B(n18981), .Z(n18762) );
  NANDN U19050 ( .A(n18982), .B(n18983), .Z(n18981) );
  NANDN U19051 ( .A(n18984), .B(n18985), .Z(n18983) );
  NANDN U19052 ( .A(n18985), .B(n18984), .Z(n18980) );
  ANDN U19053 ( .B(B[219]), .A(n58), .Z(n18764) );
  XNOR U19054 ( .A(n18772), .B(n18986), .Z(n18765) );
  XNOR U19055 ( .A(n18771), .B(n18769), .Z(n18986) );
  AND U19056 ( .A(n18987), .B(n18988), .Z(n18769) );
  NANDN U19057 ( .A(n18989), .B(n18990), .Z(n18988) );
  OR U19058 ( .A(n18991), .B(n18992), .Z(n18990) );
  NAND U19059 ( .A(n18992), .B(n18991), .Z(n18987) );
  ANDN U19060 ( .B(B[220]), .A(n59), .Z(n18771) );
  XNOR U19061 ( .A(n18779), .B(n18993), .Z(n18772) );
  XNOR U19062 ( .A(n18778), .B(n18776), .Z(n18993) );
  AND U19063 ( .A(n18994), .B(n18995), .Z(n18776) );
  NANDN U19064 ( .A(n18996), .B(n18997), .Z(n18995) );
  NANDN U19065 ( .A(n18998), .B(n18999), .Z(n18997) );
  NANDN U19066 ( .A(n18999), .B(n18998), .Z(n18994) );
  ANDN U19067 ( .B(B[221]), .A(n60), .Z(n18778) );
  XNOR U19068 ( .A(n18786), .B(n19000), .Z(n18779) );
  XNOR U19069 ( .A(n18785), .B(n18783), .Z(n19000) );
  AND U19070 ( .A(n19001), .B(n19002), .Z(n18783) );
  NANDN U19071 ( .A(n19003), .B(n19004), .Z(n19002) );
  OR U19072 ( .A(n19005), .B(n19006), .Z(n19004) );
  NAND U19073 ( .A(n19006), .B(n19005), .Z(n19001) );
  ANDN U19074 ( .B(B[222]), .A(n61), .Z(n18785) );
  XNOR U19075 ( .A(n18793), .B(n19007), .Z(n18786) );
  XNOR U19076 ( .A(n18792), .B(n18790), .Z(n19007) );
  AND U19077 ( .A(n19008), .B(n19009), .Z(n18790) );
  NANDN U19078 ( .A(n19010), .B(n19011), .Z(n19009) );
  NANDN U19079 ( .A(n19012), .B(n19013), .Z(n19011) );
  NANDN U19080 ( .A(n19013), .B(n19012), .Z(n19008) );
  ANDN U19081 ( .B(B[223]), .A(n62), .Z(n18792) );
  XNOR U19082 ( .A(n18800), .B(n19014), .Z(n18793) );
  XNOR U19083 ( .A(n18799), .B(n18797), .Z(n19014) );
  AND U19084 ( .A(n19015), .B(n19016), .Z(n18797) );
  NANDN U19085 ( .A(n19017), .B(n19018), .Z(n19016) );
  OR U19086 ( .A(n19019), .B(n19020), .Z(n19018) );
  NAND U19087 ( .A(n19020), .B(n19019), .Z(n19015) );
  ANDN U19088 ( .B(B[224]), .A(n63), .Z(n18799) );
  XNOR U19089 ( .A(n18807), .B(n19021), .Z(n18800) );
  XNOR U19090 ( .A(n18806), .B(n18804), .Z(n19021) );
  AND U19091 ( .A(n19022), .B(n19023), .Z(n18804) );
  NANDN U19092 ( .A(n19024), .B(n19025), .Z(n19023) );
  NANDN U19093 ( .A(n19026), .B(n19027), .Z(n19025) );
  NANDN U19094 ( .A(n19027), .B(n19026), .Z(n19022) );
  ANDN U19095 ( .B(B[225]), .A(n64), .Z(n18806) );
  XNOR U19096 ( .A(n18814), .B(n19028), .Z(n18807) );
  XNOR U19097 ( .A(n18813), .B(n18811), .Z(n19028) );
  AND U19098 ( .A(n19029), .B(n19030), .Z(n18811) );
  NANDN U19099 ( .A(n19031), .B(n19032), .Z(n19030) );
  OR U19100 ( .A(n19033), .B(n19034), .Z(n19032) );
  NAND U19101 ( .A(n19034), .B(n19033), .Z(n19029) );
  ANDN U19102 ( .B(B[226]), .A(n65), .Z(n18813) );
  XNOR U19103 ( .A(n18821), .B(n19035), .Z(n18814) );
  XNOR U19104 ( .A(n18820), .B(n18818), .Z(n19035) );
  AND U19105 ( .A(n19036), .B(n19037), .Z(n18818) );
  NANDN U19106 ( .A(n19038), .B(n19039), .Z(n19037) );
  NANDN U19107 ( .A(n19040), .B(n19041), .Z(n19039) );
  NANDN U19108 ( .A(n19041), .B(n19040), .Z(n19036) );
  ANDN U19109 ( .B(B[227]), .A(n66), .Z(n18820) );
  XNOR U19110 ( .A(n18828), .B(n19042), .Z(n18821) );
  XNOR U19111 ( .A(n18827), .B(n18825), .Z(n19042) );
  AND U19112 ( .A(n19043), .B(n19044), .Z(n18825) );
  NANDN U19113 ( .A(n19045), .B(n19046), .Z(n19044) );
  OR U19114 ( .A(n19047), .B(n19048), .Z(n19046) );
  NAND U19115 ( .A(n19048), .B(n19047), .Z(n19043) );
  ANDN U19116 ( .B(B[228]), .A(n67), .Z(n18827) );
  XNOR U19117 ( .A(n18835), .B(n19049), .Z(n18828) );
  XNOR U19118 ( .A(n18834), .B(n18832), .Z(n19049) );
  AND U19119 ( .A(n19050), .B(n19051), .Z(n18832) );
  NANDN U19120 ( .A(n19052), .B(n19053), .Z(n19051) );
  NANDN U19121 ( .A(n19054), .B(n19055), .Z(n19053) );
  NANDN U19122 ( .A(n19055), .B(n19054), .Z(n19050) );
  ANDN U19123 ( .B(B[229]), .A(n68), .Z(n18834) );
  XNOR U19124 ( .A(n18842), .B(n19056), .Z(n18835) );
  XNOR U19125 ( .A(n18841), .B(n18839), .Z(n19056) );
  AND U19126 ( .A(n19057), .B(n19058), .Z(n18839) );
  NANDN U19127 ( .A(n19059), .B(n19060), .Z(n19058) );
  OR U19128 ( .A(n19061), .B(n19062), .Z(n19060) );
  NAND U19129 ( .A(n19062), .B(n19061), .Z(n19057) );
  ANDN U19130 ( .B(B[230]), .A(n69), .Z(n18841) );
  XNOR U19131 ( .A(n18849), .B(n19063), .Z(n18842) );
  XNOR U19132 ( .A(n18848), .B(n18846), .Z(n19063) );
  AND U19133 ( .A(n19064), .B(n19065), .Z(n18846) );
  NANDN U19134 ( .A(n19066), .B(n19067), .Z(n19065) );
  NANDN U19135 ( .A(n19068), .B(n19069), .Z(n19067) );
  NANDN U19136 ( .A(n19069), .B(n19068), .Z(n19064) );
  ANDN U19137 ( .B(B[231]), .A(n70), .Z(n18848) );
  XNOR U19138 ( .A(n18856), .B(n19070), .Z(n18849) );
  XNOR U19139 ( .A(n18855), .B(n18853), .Z(n19070) );
  AND U19140 ( .A(n19071), .B(n19072), .Z(n18853) );
  NANDN U19141 ( .A(n19073), .B(n19074), .Z(n19072) );
  OR U19142 ( .A(n19075), .B(n19076), .Z(n19074) );
  NAND U19143 ( .A(n19076), .B(n19075), .Z(n19071) );
  ANDN U19144 ( .B(B[232]), .A(n71), .Z(n18855) );
  XNOR U19145 ( .A(n18863), .B(n19077), .Z(n18856) );
  XNOR U19146 ( .A(n18862), .B(n18860), .Z(n19077) );
  AND U19147 ( .A(n19078), .B(n19079), .Z(n18860) );
  NANDN U19148 ( .A(n19080), .B(n19081), .Z(n19079) );
  NANDN U19149 ( .A(n19082), .B(n19083), .Z(n19081) );
  NANDN U19150 ( .A(n19083), .B(n19082), .Z(n19078) );
  ANDN U19151 ( .B(B[233]), .A(n72), .Z(n18862) );
  XNOR U19152 ( .A(n18870), .B(n19084), .Z(n18863) );
  XNOR U19153 ( .A(n18869), .B(n18867), .Z(n19084) );
  AND U19154 ( .A(n19085), .B(n19086), .Z(n18867) );
  NANDN U19155 ( .A(n19087), .B(n19088), .Z(n19086) );
  OR U19156 ( .A(n19089), .B(n19090), .Z(n19088) );
  NAND U19157 ( .A(n19090), .B(n19089), .Z(n19085) );
  ANDN U19158 ( .B(B[234]), .A(n73), .Z(n18869) );
  XNOR U19159 ( .A(n18877), .B(n19091), .Z(n18870) );
  XNOR U19160 ( .A(n18876), .B(n18874), .Z(n19091) );
  AND U19161 ( .A(n19092), .B(n19093), .Z(n18874) );
  NANDN U19162 ( .A(n19094), .B(n19095), .Z(n19093) );
  NANDN U19163 ( .A(n19096), .B(n19097), .Z(n19095) );
  NANDN U19164 ( .A(n19097), .B(n19096), .Z(n19092) );
  ANDN U19165 ( .B(B[235]), .A(n74), .Z(n18876) );
  XNOR U19166 ( .A(n18884), .B(n19098), .Z(n18877) );
  XNOR U19167 ( .A(n18883), .B(n18881), .Z(n19098) );
  AND U19168 ( .A(n19099), .B(n19100), .Z(n18881) );
  NANDN U19169 ( .A(n19101), .B(n19102), .Z(n19100) );
  OR U19170 ( .A(n19103), .B(n19104), .Z(n19102) );
  NAND U19171 ( .A(n19104), .B(n19103), .Z(n19099) );
  ANDN U19172 ( .B(B[236]), .A(n75), .Z(n18883) );
  XNOR U19173 ( .A(n18891), .B(n19105), .Z(n18884) );
  XNOR U19174 ( .A(n18890), .B(n18888), .Z(n19105) );
  AND U19175 ( .A(n19106), .B(n19107), .Z(n18888) );
  NANDN U19176 ( .A(n19108), .B(n19109), .Z(n19107) );
  NANDN U19177 ( .A(n19110), .B(n19111), .Z(n19109) );
  NANDN U19178 ( .A(n19111), .B(n19110), .Z(n19106) );
  ANDN U19179 ( .B(B[237]), .A(n76), .Z(n18890) );
  XNOR U19180 ( .A(n18898), .B(n19112), .Z(n18891) );
  XNOR U19181 ( .A(n18897), .B(n18895), .Z(n19112) );
  AND U19182 ( .A(n19113), .B(n19114), .Z(n18895) );
  NANDN U19183 ( .A(n19115), .B(n19116), .Z(n19114) );
  OR U19184 ( .A(n19117), .B(n19118), .Z(n19116) );
  NAND U19185 ( .A(n19118), .B(n19117), .Z(n19113) );
  ANDN U19186 ( .B(B[238]), .A(n77), .Z(n18897) );
  XNOR U19187 ( .A(n18905), .B(n19119), .Z(n18898) );
  XNOR U19188 ( .A(n18904), .B(n18902), .Z(n19119) );
  AND U19189 ( .A(n19120), .B(n19121), .Z(n18902) );
  NANDN U19190 ( .A(n19122), .B(n19123), .Z(n19121) );
  NANDN U19191 ( .A(n19124), .B(n19125), .Z(n19123) );
  NANDN U19192 ( .A(n19125), .B(n19124), .Z(n19120) );
  ANDN U19193 ( .B(B[239]), .A(n78), .Z(n18904) );
  XNOR U19194 ( .A(n18912), .B(n19126), .Z(n18905) );
  XNOR U19195 ( .A(n18911), .B(n18909), .Z(n19126) );
  AND U19196 ( .A(n19127), .B(n19128), .Z(n18909) );
  NANDN U19197 ( .A(n19129), .B(n19130), .Z(n19128) );
  OR U19198 ( .A(n19131), .B(n19132), .Z(n19130) );
  NAND U19199 ( .A(n19132), .B(n19131), .Z(n19127) );
  ANDN U19200 ( .B(B[240]), .A(n79), .Z(n18911) );
  XNOR U19201 ( .A(n18919), .B(n19133), .Z(n18912) );
  XNOR U19202 ( .A(n18918), .B(n18916), .Z(n19133) );
  AND U19203 ( .A(n19134), .B(n19135), .Z(n18916) );
  NANDN U19204 ( .A(n19136), .B(n19137), .Z(n19135) );
  NANDN U19205 ( .A(n19138), .B(n19139), .Z(n19137) );
  NANDN U19206 ( .A(n19139), .B(n19138), .Z(n19134) );
  ANDN U19207 ( .B(B[241]), .A(n80), .Z(n18918) );
  XNOR U19208 ( .A(n18926), .B(n19140), .Z(n18919) );
  XNOR U19209 ( .A(n18925), .B(n18923), .Z(n19140) );
  AND U19210 ( .A(n19141), .B(n19142), .Z(n18923) );
  NANDN U19211 ( .A(n19143), .B(n19144), .Z(n19142) );
  OR U19212 ( .A(n19145), .B(n19146), .Z(n19144) );
  NAND U19213 ( .A(n19146), .B(n19145), .Z(n19141) );
  ANDN U19214 ( .B(B[242]), .A(n81), .Z(n18925) );
  XNOR U19215 ( .A(n18933), .B(n19147), .Z(n18926) );
  XNOR U19216 ( .A(n18932), .B(n18930), .Z(n19147) );
  AND U19217 ( .A(n19148), .B(n19149), .Z(n18930) );
  NANDN U19218 ( .A(n19150), .B(n19151), .Z(n19149) );
  NAND U19219 ( .A(n19152), .B(n19153), .Z(n19151) );
  ANDN U19220 ( .B(B[243]), .A(n82), .Z(n18932) );
  XOR U19221 ( .A(n18939), .B(n19154), .Z(n18933) );
  XNOR U19222 ( .A(n18937), .B(n18940), .Z(n19154) );
  NAND U19223 ( .A(A[2]), .B(B[244]), .Z(n18940) );
  NANDN U19224 ( .A(n19155), .B(n19156), .Z(n18937) );
  AND U19225 ( .A(A[0]), .B(B[245]), .Z(n19156) );
  XNOR U19226 ( .A(n18942), .B(n19157), .Z(n18939) );
  NAND U19227 ( .A(A[0]), .B(B[246]), .Z(n19157) );
  NAND U19228 ( .A(B[245]), .B(A[1]), .Z(n18942) );
  NAND U19229 ( .A(n19158), .B(n19159), .Z(n304) );
  NANDN U19230 ( .A(n19160), .B(n19161), .Z(n19159) );
  OR U19231 ( .A(n19162), .B(n19163), .Z(n19161) );
  NAND U19232 ( .A(n19163), .B(n19162), .Z(n19158) );
  XOR U19233 ( .A(n306), .B(n305), .Z(\A1[243] ) );
  XOR U19234 ( .A(n19163), .B(n19164), .Z(n305) );
  XNOR U19235 ( .A(n19162), .B(n19160), .Z(n19164) );
  AND U19236 ( .A(n19165), .B(n19166), .Z(n19160) );
  NANDN U19237 ( .A(n19167), .B(n19168), .Z(n19166) );
  NANDN U19238 ( .A(n19169), .B(n19170), .Z(n19168) );
  NANDN U19239 ( .A(n19170), .B(n19169), .Z(n19165) );
  ANDN U19240 ( .B(B[214]), .A(n54), .Z(n19162) );
  XNOR U19241 ( .A(n18957), .B(n19171), .Z(n19163) );
  XNOR U19242 ( .A(n18956), .B(n18954), .Z(n19171) );
  AND U19243 ( .A(n19172), .B(n19173), .Z(n18954) );
  NANDN U19244 ( .A(n19174), .B(n19175), .Z(n19173) );
  OR U19245 ( .A(n19176), .B(n19177), .Z(n19175) );
  NAND U19246 ( .A(n19177), .B(n19176), .Z(n19172) );
  ANDN U19247 ( .B(B[215]), .A(n55), .Z(n18956) );
  XNOR U19248 ( .A(n18964), .B(n19178), .Z(n18957) );
  XNOR U19249 ( .A(n18963), .B(n18961), .Z(n19178) );
  AND U19250 ( .A(n19179), .B(n19180), .Z(n18961) );
  NANDN U19251 ( .A(n19181), .B(n19182), .Z(n19180) );
  NANDN U19252 ( .A(n19183), .B(n19184), .Z(n19182) );
  NANDN U19253 ( .A(n19184), .B(n19183), .Z(n19179) );
  ANDN U19254 ( .B(B[216]), .A(n56), .Z(n18963) );
  XNOR U19255 ( .A(n18971), .B(n19185), .Z(n18964) );
  XNOR U19256 ( .A(n18970), .B(n18968), .Z(n19185) );
  AND U19257 ( .A(n19186), .B(n19187), .Z(n18968) );
  NANDN U19258 ( .A(n19188), .B(n19189), .Z(n19187) );
  OR U19259 ( .A(n19190), .B(n19191), .Z(n19189) );
  NAND U19260 ( .A(n19191), .B(n19190), .Z(n19186) );
  ANDN U19261 ( .B(B[217]), .A(n57), .Z(n18970) );
  XNOR U19262 ( .A(n18978), .B(n19192), .Z(n18971) );
  XNOR U19263 ( .A(n18977), .B(n18975), .Z(n19192) );
  AND U19264 ( .A(n19193), .B(n19194), .Z(n18975) );
  NANDN U19265 ( .A(n19195), .B(n19196), .Z(n19194) );
  NANDN U19266 ( .A(n19197), .B(n19198), .Z(n19196) );
  NANDN U19267 ( .A(n19198), .B(n19197), .Z(n19193) );
  ANDN U19268 ( .B(B[218]), .A(n58), .Z(n18977) );
  XNOR U19269 ( .A(n18985), .B(n19199), .Z(n18978) );
  XNOR U19270 ( .A(n18984), .B(n18982), .Z(n19199) );
  AND U19271 ( .A(n19200), .B(n19201), .Z(n18982) );
  NANDN U19272 ( .A(n19202), .B(n19203), .Z(n19201) );
  OR U19273 ( .A(n19204), .B(n19205), .Z(n19203) );
  NAND U19274 ( .A(n19205), .B(n19204), .Z(n19200) );
  ANDN U19275 ( .B(B[219]), .A(n59), .Z(n18984) );
  XNOR U19276 ( .A(n18992), .B(n19206), .Z(n18985) );
  XNOR U19277 ( .A(n18991), .B(n18989), .Z(n19206) );
  AND U19278 ( .A(n19207), .B(n19208), .Z(n18989) );
  NANDN U19279 ( .A(n19209), .B(n19210), .Z(n19208) );
  NANDN U19280 ( .A(n19211), .B(n19212), .Z(n19210) );
  NANDN U19281 ( .A(n19212), .B(n19211), .Z(n19207) );
  ANDN U19282 ( .B(B[220]), .A(n60), .Z(n18991) );
  XNOR U19283 ( .A(n18999), .B(n19213), .Z(n18992) );
  XNOR U19284 ( .A(n18998), .B(n18996), .Z(n19213) );
  AND U19285 ( .A(n19214), .B(n19215), .Z(n18996) );
  NANDN U19286 ( .A(n19216), .B(n19217), .Z(n19215) );
  OR U19287 ( .A(n19218), .B(n19219), .Z(n19217) );
  NAND U19288 ( .A(n19219), .B(n19218), .Z(n19214) );
  ANDN U19289 ( .B(B[221]), .A(n61), .Z(n18998) );
  XNOR U19290 ( .A(n19006), .B(n19220), .Z(n18999) );
  XNOR U19291 ( .A(n19005), .B(n19003), .Z(n19220) );
  AND U19292 ( .A(n19221), .B(n19222), .Z(n19003) );
  NANDN U19293 ( .A(n19223), .B(n19224), .Z(n19222) );
  NANDN U19294 ( .A(n19225), .B(n19226), .Z(n19224) );
  NANDN U19295 ( .A(n19226), .B(n19225), .Z(n19221) );
  ANDN U19296 ( .B(B[222]), .A(n62), .Z(n19005) );
  XNOR U19297 ( .A(n19013), .B(n19227), .Z(n19006) );
  XNOR U19298 ( .A(n19012), .B(n19010), .Z(n19227) );
  AND U19299 ( .A(n19228), .B(n19229), .Z(n19010) );
  NANDN U19300 ( .A(n19230), .B(n19231), .Z(n19229) );
  OR U19301 ( .A(n19232), .B(n19233), .Z(n19231) );
  NAND U19302 ( .A(n19233), .B(n19232), .Z(n19228) );
  ANDN U19303 ( .B(B[223]), .A(n63), .Z(n19012) );
  XNOR U19304 ( .A(n19020), .B(n19234), .Z(n19013) );
  XNOR U19305 ( .A(n19019), .B(n19017), .Z(n19234) );
  AND U19306 ( .A(n19235), .B(n19236), .Z(n19017) );
  NANDN U19307 ( .A(n19237), .B(n19238), .Z(n19236) );
  NANDN U19308 ( .A(n19239), .B(n19240), .Z(n19238) );
  NANDN U19309 ( .A(n19240), .B(n19239), .Z(n19235) );
  ANDN U19310 ( .B(B[224]), .A(n64), .Z(n19019) );
  XNOR U19311 ( .A(n19027), .B(n19241), .Z(n19020) );
  XNOR U19312 ( .A(n19026), .B(n19024), .Z(n19241) );
  AND U19313 ( .A(n19242), .B(n19243), .Z(n19024) );
  NANDN U19314 ( .A(n19244), .B(n19245), .Z(n19243) );
  OR U19315 ( .A(n19246), .B(n19247), .Z(n19245) );
  NAND U19316 ( .A(n19247), .B(n19246), .Z(n19242) );
  ANDN U19317 ( .B(B[225]), .A(n65), .Z(n19026) );
  XNOR U19318 ( .A(n19034), .B(n19248), .Z(n19027) );
  XNOR U19319 ( .A(n19033), .B(n19031), .Z(n19248) );
  AND U19320 ( .A(n19249), .B(n19250), .Z(n19031) );
  NANDN U19321 ( .A(n19251), .B(n19252), .Z(n19250) );
  NANDN U19322 ( .A(n19253), .B(n19254), .Z(n19252) );
  NANDN U19323 ( .A(n19254), .B(n19253), .Z(n19249) );
  ANDN U19324 ( .B(B[226]), .A(n66), .Z(n19033) );
  XNOR U19325 ( .A(n19041), .B(n19255), .Z(n19034) );
  XNOR U19326 ( .A(n19040), .B(n19038), .Z(n19255) );
  AND U19327 ( .A(n19256), .B(n19257), .Z(n19038) );
  NANDN U19328 ( .A(n19258), .B(n19259), .Z(n19257) );
  OR U19329 ( .A(n19260), .B(n19261), .Z(n19259) );
  NAND U19330 ( .A(n19261), .B(n19260), .Z(n19256) );
  ANDN U19331 ( .B(B[227]), .A(n67), .Z(n19040) );
  XNOR U19332 ( .A(n19048), .B(n19262), .Z(n19041) );
  XNOR U19333 ( .A(n19047), .B(n19045), .Z(n19262) );
  AND U19334 ( .A(n19263), .B(n19264), .Z(n19045) );
  NANDN U19335 ( .A(n19265), .B(n19266), .Z(n19264) );
  NANDN U19336 ( .A(n19267), .B(n19268), .Z(n19266) );
  NANDN U19337 ( .A(n19268), .B(n19267), .Z(n19263) );
  ANDN U19338 ( .B(B[228]), .A(n68), .Z(n19047) );
  XNOR U19339 ( .A(n19055), .B(n19269), .Z(n19048) );
  XNOR U19340 ( .A(n19054), .B(n19052), .Z(n19269) );
  AND U19341 ( .A(n19270), .B(n19271), .Z(n19052) );
  NANDN U19342 ( .A(n19272), .B(n19273), .Z(n19271) );
  OR U19343 ( .A(n19274), .B(n19275), .Z(n19273) );
  NAND U19344 ( .A(n19275), .B(n19274), .Z(n19270) );
  ANDN U19345 ( .B(B[229]), .A(n69), .Z(n19054) );
  XNOR U19346 ( .A(n19062), .B(n19276), .Z(n19055) );
  XNOR U19347 ( .A(n19061), .B(n19059), .Z(n19276) );
  AND U19348 ( .A(n19277), .B(n19278), .Z(n19059) );
  NANDN U19349 ( .A(n19279), .B(n19280), .Z(n19278) );
  NANDN U19350 ( .A(n19281), .B(n19282), .Z(n19280) );
  NANDN U19351 ( .A(n19282), .B(n19281), .Z(n19277) );
  ANDN U19352 ( .B(B[230]), .A(n70), .Z(n19061) );
  XNOR U19353 ( .A(n19069), .B(n19283), .Z(n19062) );
  XNOR U19354 ( .A(n19068), .B(n19066), .Z(n19283) );
  AND U19355 ( .A(n19284), .B(n19285), .Z(n19066) );
  NANDN U19356 ( .A(n19286), .B(n19287), .Z(n19285) );
  OR U19357 ( .A(n19288), .B(n19289), .Z(n19287) );
  NAND U19358 ( .A(n19289), .B(n19288), .Z(n19284) );
  ANDN U19359 ( .B(B[231]), .A(n71), .Z(n19068) );
  XNOR U19360 ( .A(n19076), .B(n19290), .Z(n19069) );
  XNOR U19361 ( .A(n19075), .B(n19073), .Z(n19290) );
  AND U19362 ( .A(n19291), .B(n19292), .Z(n19073) );
  NANDN U19363 ( .A(n19293), .B(n19294), .Z(n19292) );
  NANDN U19364 ( .A(n19295), .B(n19296), .Z(n19294) );
  NANDN U19365 ( .A(n19296), .B(n19295), .Z(n19291) );
  ANDN U19366 ( .B(B[232]), .A(n72), .Z(n19075) );
  XNOR U19367 ( .A(n19083), .B(n19297), .Z(n19076) );
  XNOR U19368 ( .A(n19082), .B(n19080), .Z(n19297) );
  AND U19369 ( .A(n19298), .B(n19299), .Z(n19080) );
  NANDN U19370 ( .A(n19300), .B(n19301), .Z(n19299) );
  OR U19371 ( .A(n19302), .B(n19303), .Z(n19301) );
  NAND U19372 ( .A(n19303), .B(n19302), .Z(n19298) );
  ANDN U19373 ( .B(B[233]), .A(n73), .Z(n19082) );
  XNOR U19374 ( .A(n19090), .B(n19304), .Z(n19083) );
  XNOR U19375 ( .A(n19089), .B(n19087), .Z(n19304) );
  AND U19376 ( .A(n19305), .B(n19306), .Z(n19087) );
  NANDN U19377 ( .A(n19307), .B(n19308), .Z(n19306) );
  NANDN U19378 ( .A(n19309), .B(n19310), .Z(n19308) );
  NANDN U19379 ( .A(n19310), .B(n19309), .Z(n19305) );
  ANDN U19380 ( .B(B[234]), .A(n74), .Z(n19089) );
  XNOR U19381 ( .A(n19097), .B(n19311), .Z(n19090) );
  XNOR U19382 ( .A(n19096), .B(n19094), .Z(n19311) );
  AND U19383 ( .A(n19312), .B(n19313), .Z(n19094) );
  NANDN U19384 ( .A(n19314), .B(n19315), .Z(n19313) );
  OR U19385 ( .A(n19316), .B(n19317), .Z(n19315) );
  NAND U19386 ( .A(n19317), .B(n19316), .Z(n19312) );
  ANDN U19387 ( .B(B[235]), .A(n75), .Z(n19096) );
  XNOR U19388 ( .A(n19104), .B(n19318), .Z(n19097) );
  XNOR U19389 ( .A(n19103), .B(n19101), .Z(n19318) );
  AND U19390 ( .A(n19319), .B(n19320), .Z(n19101) );
  NANDN U19391 ( .A(n19321), .B(n19322), .Z(n19320) );
  NANDN U19392 ( .A(n19323), .B(n19324), .Z(n19322) );
  NANDN U19393 ( .A(n19324), .B(n19323), .Z(n19319) );
  ANDN U19394 ( .B(B[236]), .A(n76), .Z(n19103) );
  XNOR U19395 ( .A(n19111), .B(n19325), .Z(n19104) );
  XNOR U19396 ( .A(n19110), .B(n19108), .Z(n19325) );
  AND U19397 ( .A(n19326), .B(n19327), .Z(n19108) );
  NANDN U19398 ( .A(n19328), .B(n19329), .Z(n19327) );
  OR U19399 ( .A(n19330), .B(n19331), .Z(n19329) );
  NAND U19400 ( .A(n19331), .B(n19330), .Z(n19326) );
  ANDN U19401 ( .B(B[237]), .A(n77), .Z(n19110) );
  XNOR U19402 ( .A(n19118), .B(n19332), .Z(n19111) );
  XNOR U19403 ( .A(n19117), .B(n19115), .Z(n19332) );
  AND U19404 ( .A(n19333), .B(n19334), .Z(n19115) );
  NANDN U19405 ( .A(n19335), .B(n19336), .Z(n19334) );
  NANDN U19406 ( .A(n19337), .B(n19338), .Z(n19336) );
  NANDN U19407 ( .A(n19338), .B(n19337), .Z(n19333) );
  ANDN U19408 ( .B(B[238]), .A(n78), .Z(n19117) );
  XNOR U19409 ( .A(n19125), .B(n19339), .Z(n19118) );
  XNOR U19410 ( .A(n19124), .B(n19122), .Z(n19339) );
  AND U19411 ( .A(n19340), .B(n19341), .Z(n19122) );
  NANDN U19412 ( .A(n19342), .B(n19343), .Z(n19341) );
  OR U19413 ( .A(n19344), .B(n19345), .Z(n19343) );
  NAND U19414 ( .A(n19345), .B(n19344), .Z(n19340) );
  ANDN U19415 ( .B(B[239]), .A(n79), .Z(n19124) );
  XNOR U19416 ( .A(n19132), .B(n19346), .Z(n19125) );
  XNOR U19417 ( .A(n19131), .B(n19129), .Z(n19346) );
  AND U19418 ( .A(n19347), .B(n19348), .Z(n19129) );
  NANDN U19419 ( .A(n19349), .B(n19350), .Z(n19348) );
  NANDN U19420 ( .A(n19351), .B(n19352), .Z(n19350) );
  NANDN U19421 ( .A(n19352), .B(n19351), .Z(n19347) );
  ANDN U19422 ( .B(B[240]), .A(n80), .Z(n19131) );
  XNOR U19423 ( .A(n19139), .B(n19353), .Z(n19132) );
  XNOR U19424 ( .A(n19138), .B(n19136), .Z(n19353) );
  AND U19425 ( .A(n19354), .B(n19355), .Z(n19136) );
  NANDN U19426 ( .A(n19356), .B(n19357), .Z(n19355) );
  OR U19427 ( .A(n19358), .B(n19359), .Z(n19357) );
  NAND U19428 ( .A(n19359), .B(n19358), .Z(n19354) );
  ANDN U19429 ( .B(B[241]), .A(n81), .Z(n19138) );
  XNOR U19430 ( .A(n19146), .B(n19360), .Z(n19139) );
  XNOR U19431 ( .A(n19145), .B(n19143), .Z(n19360) );
  AND U19432 ( .A(n19361), .B(n19362), .Z(n19143) );
  NANDN U19433 ( .A(n19363), .B(n19364), .Z(n19362) );
  NAND U19434 ( .A(n19365), .B(n19366), .Z(n19364) );
  ANDN U19435 ( .B(B[242]), .A(n82), .Z(n19145) );
  XOR U19436 ( .A(n19152), .B(n19367), .Z(n19146) );
  XNOR U19437 ( .A(n19150), .B(n19153), .Z(n19367) );
  NAND U19438 ( .A(A[2]), .B(B[243]), .Z(n19153) );
  NANDN U19439 ( .A(n19368), .B(n19369), .Z(n19150) );
  AND U19440 ( .A(A[0]), .B(B[244]), .Z(n19369) );
  XNOR U19441 ( .A(n19155), .B(n19370), .Z(n19152) );
  NAND U19442 ( .A(A[0]), .B(B[245]), .Z(n19370) );
  NAND U19443 ( .A(B[244]), .B(A[1]), .Z(n19155) );
  NAND U19444 ( .A(n19371), .B(n19372), .Z(n306) );
  NANDN U19445 ( .A(n19373), .B(n19374), .Z(n19372) );
  OR U19446 ( .A(n19375), .B(n19376), .Z(n19374) );
  NAND U19447 ( .A(n19376), .B(n19375), .Z(n19371) );
  XOR U19448 ( .A(n308), .B(n307), .Z(\A1[242] ) );
  XOR U19449 ( .A(n19376), .B(n19377), .Z(n307) );
  XNOR U19450 ( .A(n19375), .B(n19373), .Z(n19377) );
  AND U19451 ( .A(n19378), .B(n19379), .Z(n19373) );
  NANDN U19452 ( .A(n19380), .B(n19381), .Z(n19379) );
  NANDN U19453 ( .A(n19382), .B(n19383), .Z(n19381) );
  NANDN U19454 ( .A(n19383), .B(n19382), .Z(n19378) );
  ANDN U19455 ( .B(B[213]), .A(n54), .Z(n19375) );
  XNOR U19456 ( .A(n19170), .B(n19384), .Z(n19376) );
  XNOR U19457 ( .A(n19169), .B(n19167), .Z(n19384) );
  AND U19458 ( .A(n19385), .B(n19386), .Z(n19167) );
  NANDN U19459 ( .A(n19387), .B(n19388), .Z(n19386) );
  OR U19460 ( .A(n19389), .B(n19390), .Z(n19388) );
  NAND U19461 ( .A(n19390), .B(n19389), .Z(n19385) );
  ANDN U19462 ( .B(B[214]), .A(n55), .Z(n19169) );
  XNOR U19463 ( .A(n19177), .B(n19391), .Z(n19170) );
  XNOR U19464 ( .A(n19176), .B(n19174), .Z(n19391) );
  AND U19465 ( .A(n19392), .B(n19393), .Z(n19174) );
  NANDN U19466 ( .A(n19394), .B(n19395), .Z(n19393) );
  NANDN U19467 ( .A(n19396), .B(n19397), .Z(n19395) );
  NANDN U19468 ( .A(n19397), .B(n19396), .Z(n19392) );
  ANDN U19469 ( .B(B[215]), .A(n56), .Z(n19176) );
  XNOR U19470 ( .A(n19184), .B(n19398), .Z(n19177) );
  XNOR U19471 ( .A(n19183), .B(n19181), .Z(n19398) );
  AND U19472 ( .A(n19399), .B(n19400), .Z(n19181) );
  NANDN U19473 ( .A(n19401), .B(n19402), .Z(n19400) );
  OR U19474 ( .A(n19403), .B(n19404), .Z(n19402) );
  NAND U19475 ( .A(n19404), .B(n19403), .Z(n19399) );
  ANDN U19476 ( .B(B[216]), .A(n57), .Z(n19183) );
  XNOR U19477 ( .A(n19191), .B(n19405), .Z(n19184) );
  XNOR U19478 ( .A(n19190), .B(n19188), .Z(n19405) );
  AND U19479 ( .A(n19406), .B(n19407), .Z(n19188) );
  NANDN U19480 ( .A(n19408), .B(n19409), .Z(n19407) );
  NANDN U19481 ( .A(n19410), .B(n19411), .Z(n19409) );
  NANDN U19482 ( .A(n19411), .B(n19410), .Z(n19406) );
  ANDN U19483 ( .B(B[217]), .A(n58), .Z(n19190) );
  XNOR U19484 ( .A(n19198), .B(n19412), .Z(n19191) );
  XNOR U19485 ( .A(n19197), .B(n19195), .Z(n19412) );
  AND U19486 ( .A(n19413), .B(n19414), .Z(n19195) );
  NANDN U19487 ( .A(n19415), .B(n19416), .Z(n19414) );
  OR U19488 ( .A(n19417), .B(n19418), .Z(n19416) );
  NAND U19489 ( .A(n19418), .B(n19417), .Z(n19413) );
  ANDN U19490 ( .B(B[218]), .A(n59), .Z(n19197) );
  XNOR U19491 ( .A(n19205), .B(n19419), .Z(n19198) );
  XNOR U19492 ( .A(n19204), .B(n19202), .Z(n19419) );
  AND U19493 ( .A(n19420), .B(n19421), .Z(n19202) );
  NANDN U19494 ( .A(n19422), .B(n19423), .Z(n19421) );
  NANDN U19495 ( .A(n19424), .B(n19425), .Z(n19423) );
  NANDN U19496 ( .A(n19425), .B(n19424), .Z(n19420) );
  ANDN U19497 ( .B(B[219]), .A(n60), .Z(n19204) );
  XNOR U19498 ( .A(n19212), .B(n19426), .Z(n19205) );
  XNOR U19499 ( .A(n19211), .B(n19209), .Z(n19426) );
  AND U19500 ( .A(n19427), .B(n19428), .Z(n19209) );
  NANDN U19501 ( .A(n19429), .B(n19430), .Z(n19428) );
  OR U19502 ( .A(n19431), .B(n19432), .Z(n19430) );
  NAND U19503 ( .A(n19432), .B(n19431), .Z(n19427) );
  ANDN U19504 ( .B(B[220]), .A(n61), .Z(n19211) );
  XNOR U19505 ( .A(n19219), .B(n19433), .Z(n19212) );
  XNOR U19506 ( .A(n19218), .B(n19216), .Z(n19433) );
  AND U19507 ( .A(n19434), .B(n19435), .Z(n19216) );
  NANDN U19508 ( .A(n19436), .B(n19437), .Z(n19435) );
  NANDN U19509 ( .A(n19438), .B(n19439), .Z(n19437) );
  NANDN U19510 ( .A(n19439), .B(n19438), .Z(n19434) );
  ANDN U19511 ( .B(B[221]), .A(n62), .Z(n19218) );
  XNOR U19512 ( .A(n19226), .B(n19440), .Z(n19219) );
  XNOR U19513 ( .A(n19225), .B(n19223), .Z(n19440) );
  AND U19514 ( .A(n19441), .B(n19442), .Z(n19223) );
  NANDN U19515 ( .A(n19443), .B(n19444), .Z(n19442) );
  OR U19516 ( .A(n19445), .B(n19446), .Z(n19444) );
  NAND U19517 ( .A(n19446), .B(n19445), .Z(n19441) );
  ANDN U19518 ( .B(B[222]), .A(n63), .Z(n19225) );
  XNOR U19519 ( .A(n19233), .B(n19447), .Z(n19226) );
  XNOR U19520 ( .A(n19232), .B(n19230), .Z(n19447) );
  AND U19521 ( .A(n19448), .B(n19449), .Z(n19230) );
  NANDN U19522 ( .A(n19450), .B(n19451), .Z(n19449) );
  NANDN U19523 ( .A(n19452), .B(n19453), .Z(n19451) );
  NANDN U19524 ( .A(n19453), .B(n19452), .Z(n19448) );
  ANDN U19525 ( .B(B[223]), .A(n64), .Z(n19232) );
  XNOR U19526 ( .A(n19240), .B(n19454), .Z(n19233) );
  XNOR U19527 ( .A(n19239), .B(n19237), .Z(n19454) );
  AND U19528 ( .A(n19455), .B(n19456), .Z(n19237) );
  NANDN U19529 ( .A(n19457), .B(n19458), .Z(n19456) );
  OR U19530 ( .A(n19459), .B(n19460), .Z(n19458) );
  NAND U19531 ( .A(n19460), .B(n19459), .Z(n19455) );
  ANDN U19532 ( .B(B[224]), .A(n65), .Z(n19239) );
  XNOR U19533 ( .A(n19247), .B(n19461), .Z(n19240) );
  XNOR U19534 ( .A(n19246), .B(n19244), .Z(n19461) );
  AND U19535 ( .A(n19462), .B(n19463), .Z(n19244) );
  NANDN U19536 ( .A(n19464), .B(n19465), .Z(n19463) );
  NANDN U19537 ( .A(n19466), .B(n19467), .Z(n19465) );
  NANDN U19538 ( .A(n19467), .B(n19466), .Z(n19462) );
  ANDN U19539 ( .B(B[225]), .A(n66), .Z(n19246) );
  XNOR U19540 ( .A(n19254), .B(n19468), .Z(n19247) );
  XNOR U19541 ( .A(n19253), .B(n19251), .Z(n19468) );
  AND U19542 ( .A(n19469), .B(n19470), .Z(n19251) );
  NANDN U19543 ( .A(n19471), .B(n19472), .Z(n19470) );
  OR U19544 ( .A(n19473), .B(n19474), .Z(n19472) );
  NAND U19545 ( .A(n19474), .B(n19473), .Z(n19469) );
  ANDN U19546 ( .B(B[226]), .A(n67), .Z(n19253) );
  XNOR U19547 ( .A(n19261), .B(n19475), .Z(n19254) );
  XNOR U19548 ( .A(n19260), .B(n19258), .Z(n19475) );
  AND U19549 ( .A(n19476), .B(n19477), .Z(n19258) );
  NANDN U19550 ( .A(n19478), .B(n19479), .Z(n19477) );
  NANDN U19551 ( .A(n19480), .B(n19481), .Z(n19479) );
  NANDN U19552 ( .A(n19481), .B(n19480), .Z(n19476) );
  ANDN U19553 ( .B(B[227]), .A(n68), .Z(n19260) );
  XNOR U19554 ( .A(n19268), .B(n19482), .Z(n19261) );
  XNOR U19555 ( .A(n19267), .B(n19265), .Z(n19482) );
  AND U19556 ( .A(n19483), .B(n19484), .Z(n19265) );
  NANDN U19557 ( .A(n19485), .B(n19486), .Z(n19484) );
  OR U19558 ( .A(n19487), .B(n19488), .Z(n19486) );
  NAND U19559 ( .A(n19488), .B(n19487), .Z(n19483) );
  ANDN U19560 ( .B(B[228]), .A(n69), .Z(n19267) );
  XNOR U19561 ( .A(n19275), .B(n19489), .Z(n19268) );
  XNOR U19562 ( .A(n19274), .B(n19272), .Z(n19489) );
  AND U19563 ( .A(n19490), .B(n19491), .Z(n19272) );
  NANDN U19564 ( .A(n19492), .B(n19493), .Z(n19491) );
  NANDN U19565 ( .A(n19494), .B(n19495), .Z(n19493) );
  NANDN U19566 ( .A(n19495), .B(n19494), .Z(n19490) );
  ANDN U19567 ( .B(B[229]), .A(n70), .Z(n19274) );
  XNOR U19568 ( .A(n19282), .B(n19496), .Z(n19275) );
  XNOR U19569 ( .A(n19281), .B(n19279), .Z(n19496) );
  AND U19570 ( .A(n19497), .B(n19498), .Z(n19279) );
  NANDN U19571 ( .A(n19499), .B(n19500), .Z(n19498) );
  OR U19572 ( .A(n19501), .B(n19502), .Z(n19500) );
  NAND U19573 ( .A(n19502), .B(n19501), .Z(n19497) );
  ANDN U19574 ( .B(B[230]), .A(n71), .Z(n19281) );
  XNOR U19575 ( .A(n19289), .B(n19503), .Z(n19282) );
  XNOR U19576 ( .A(n19288), .B(n19286), .Z(n19503) );
  AND U19577 ( .A(n19504), .B(n19505), .Z(n19286) );
  NANDN U19578 ( .A(n19506), .B(n19507), .Z(n19505) );
  NANDN U19579 ( .A(n19508), .B(n19509), .Z(n19507) );
  NANDN U19580 ( .A(n19509), .B(n19508), .Z(n19504) );
  ANDN U19581 ( .B(B[231]), .A(n72), .Z(n19288) );
  XNOR U19582 ( .A(n19296), .B(n19510), .Z(n19289) );
  XNOR U19583 ( .A(n19295), .B(n19293), .Z(n19510) );
  AND U19584 ( .A(n19511), .B(n19512), .Z(n19293) );
  NANDN U19585 ( .A(n19513), .B(n19514), .Z(n19512) );
  OR U19586 ( .A(n19515), .B(n19516), .Z(n19514) );
  NAND U19587 ( .A(n19516), .B(n19515), .Z(n19511) );
  ANDN U19588 ( .B(B[232]), .A(n73), .Z(n19295) );
  XNOR U19589 ( .A(n19303), .B(n19517), .Z(n19296) );
  XNOR U19590 ( .A(n19302), .B(n19300), .Z(n19517) );
  AND U19591 ( .A(n19518), .B(n19519), .Z(n19300) );
  NANDN U19592 ( .A(n19520), .B(n19521), .Z(n19519) );
  NANDN U19593 ( .A(n19522), .B(n19523), .Z(n19521) );
  NANDN U19594 ( .A(n19523), .B(n19522), .Z(n19518) );
  ANDN U19595 ( .B(B[233]), .A(n74), .Z(n19302) );
  XNOR U19596 ( .A(n19310), .B(n19524), .Z(n19303) );
  XNOR U19597 ( .A(n19309), .B(n19307), .Z(n19524) );
  AND U19598 ( .A(n19525), .B(n19526), .Z(n19307) );
  NANDN U19599 ( .A(n19527), .B(n19528), .Z(n19526) );
  OR U19600 ( .A(n19529), .B(n19530), .Z(n19528) );
  NAND U19601 ( .A(n19530), .B(n19529), .Z(n19525) );
  ANDN U19602 ( .B(B[234]), .A(n75), .Z(n19309) );
  XNOR U19603 ( .A(n19317), .B(n19531), .Z(n19310) );
  XNOR U19604 ( .A(n19316), .B(n19314), .Z(n19531) );
  AND U19605 ( .A(n19532), .B(n19533), .Z(n19314) );
  NANDN U19606 ( .A(n19534), .B(n19535), .Z(n19533) );
  NANDN U19607 ( .A(n19536), .B(n19537), .Z(n19535) );
  NANDN U19608 ( .A(n19537), .B(n19536), .Z(n19532) );
  ANDN U19609 ( .B(B[235]), .A(n76), .Z(n19316) );
  XNOR U19610 ( .A(n19324), .B(n19538), .Z(n19317) );
  XNOR U19611 ( .A(n19323), .B(n19321), .Z(n19538) );
  AND U19612 ( .A(n19539), .B(n19540), .Z(n19321) );
  NANDN U19613 ( .A(n19541), .B(n19542), .Z(n19540) );
  OR U19614 ( .A(n19543), .B(n19544), .Z(n19542) );
  NAND U19615 ( .A(n19544), .B(n19543), .Z(n19539) );
  ANDN U19616 ( .B(B[236]), .A(n77), .Z(n19323) );
  XNOR U19617 ( .A(n19331), .B(n19545), .Z(n19324) );
  XNOR U19618 ( .A(n19330), .B(n19328), .Z(n19545) );
  AND U19619 ( .A(n19546), .B(n19547), .Z(n19328) );
  NANDN U19620 ( .A(n19548), .B(n19549), .Z(n19547) );
  NANDN U19621 ( .A(n19550), .B(n19551), .Z(n19549) );
  NANDN U19622 ( .A(n19551), .B(n19550), .Z(n19546) );
  ANDN U19623 ( .B(B[237]), .A(n78), .Z(n19330) );
  XNOR U19624 ( .A(n19338), .B(n19552), .Z(n19331) );
  XNOR U19625 ( .A(n19337), .B(n19335), .Z(n19552) );
  AND U19626 ( .A(n19553), .B(n19554), .Z(n19335) );
  NANDN U19627 ( .A(n19555), .B(n19556), .Z(n19554) );
  OR U19628 ( .A(n19557), .B(n19558), .Z(n19556) );
  NAND U19629 ( .A(n19558), .B(n19557), .Z(n19553) );
  ANDN U19630 ( .B(B[238]), .A(n79), .Z(n19337) );
  XNOR U19631 ( .A(n19345), .B(n19559), .Z(n19338) );
  XNOR U19632 ( .A(n19344), .B(n19342), .Z(n19559) );
  AND U19633 ( .A(n19560), .B(n19561), .Z(n19342) );
  NANDN U19634 ( .A(n19562), .B(n19563), .Z(n19561) );
  NANDN U19635 ( .A(n19564), .B(n19565), .Z(n19563) );
  NANDN U19636 ( .A(n19565), .B(n19564), .Z(n19560) );
  ANDN U19637 ( .B(B[239]), .A(n80), .Z(n19344) );
  XNOR U19638 ( .A(n19352), .B(n19566), .Z(n19345) );
  XNOR U19639 ( .A(n19351), .B(n19349), .Z(n19566) );
  AND U19640 ( .A(n19567), .B(n19568), .Z(n19349) );
  NANDN U19641 ( .A(n19569), .B(n19570), .Z(n19568) );
  OR U19642 ( .A(n19571), .B(n19572), .Z(n19570) );
  NAND U19643 ( .A(n19572), .B(n19571), .Z(n19567) );
  ANDN U19644 ( .B(B[240]), .A(n81), .Z(n19351) );
  XNOR U19645 ( .A(n19359), .B(n19573), .Z(n19352) );
  XNOR U19646 ( .A(n19358), .B(n19356), .Z(n19573) );
  AND U19647 ( .A(n19574), .B(n19575), .Z(n19356) );
  NANDN U19648 ( .A(n19576), .B(n19577), .Z(n19575) );
  NAND U19649 ( .A(n19578), .B(n19579), .Z(n19577) );
  ANDN U19650 ( .B(B[241]), .A(n82), .Z(n19358) );
  XOR U19651 ( .A(n19365), .B(n19580), .Z(n19359) );
  XNOR U19652 ( .A(n19363), .B(n19366), .Z(n19580) );
  NAND U19653 ( .A(A[2]), .B(B[242]), .Z(n19366) );
  NANDN U19654 ( .A(n19581), .B(n19582), .Z(n19363) );
  AND U19655 ( .A(A[0]), .B(B[243]), .Z(n19582) );
  XNOR U19656 ( .A(n19368), .B(n19583), .Z(n19365) );
  NAND U19657 ( .A(A[0]), .B(B[244]), .Z(n19583) );
  NAND U19658 ( .A(B[243]), .B(A[1]), .Z(n19368) );
  NAND U19659 ( .A(n19584), .B(n19585), .Z(n308) );
  NANDN U19660 ( .A(n19586), .B(n19587), .Z(n19585) );
  OR U19661 ( .A(n19588), .B(n19589), .Z(n19587) );
  NAND U19662 ( .A(n19589), .B(n19588), .Z(n19584) );
  XOR U19663 ( .A(n310), .B(n309), .Z(\A1[241] ) );
  XOR U19664 ( .A(n19589), .B(n19590), .Z(n309) );
  XNOR U19665 ( .A(n19588), .B(n19586), .Z(n19590) );
  AND U19666 ( .A(n19591), .B(n19592), .Z(n19586) );
  NANDN U19667 ( .A(n19593), .B(n19594), .Z(n19592) );
  NANDN U19668 ( .A(n19595), .B(n19596), .Z(n19594) );
  NANDN U19669 ( .A(n19596), .B(n19595), .Z(n19591) );
  ANDN U19670 ( .B(B[212]), .A(n54), .Z(n19588) );
  XNOR U19671 ( .A(n19383), .B(n19597), .Z(n19589) );
  XNOR U19672 ( .A(n19382), .B(n19380), .Z(n19597) );
  AND U19673 ( .A(n19598), .B(n19599), .Z(n19380) );
  NANDN U19674 ( .A(n19600), .B(n19601), .Z(n19599) );
  OR U19675 ( .A(n19602), .B(n19603), .Z(n19601) );
  NAND U19676 ( .A(n19603), .B(n19602), .Z(n19598) );
  ANDN U19677 ( .B(B[213]), .A(n55), .Z(n19382) );
  XNOR U19678 ( .A(n19390), .B(n19604), .Z(n19383) );
  XNOR U19679 ( .A(n19389), .B(n19387), .Z(n19604) );
  AND U19680 ( .A(n19605), .B(n19606), .Z(n19387) );
  NANDN U19681 ( .A(n19607), .B(n19608), .Z(n19606) );
  NANDN U19682 ( .A(n19609), .B(n19610), .Z(n19608) );
  NANDN U19683 ( .A(n19610), .B(n19609), .Z(n19605) );
  ANDN U19684 ( .B(B[214]), .A(n56), .Z(n19389) );
  XNOR U19685 ( .A(n19397), .B(n19611), .Z(n19390) );
  XNOR U19686 ( .A(n19396), .B(n19394), .Z(n19611) );
  AND U19687 ( .A(n19612), .B(n19613), .Z(n19394) );
  NANDN U19688 ( .A(n19614), .B(n19615), .Z(n19613) );
  OR U19689 ( .A(n19616), .B(n19617), .Z(n19615) );
  NAND U19690 ( .A(n19617), .B(n19616), .Z(n19612) );
  ANDN U19691 ( .B(B[215]), .A(n57), .Z(n19396) );
  XNOR U19692 ( .A(n19404), .B(n19618), .Z(n19397) );
  XNOR U19693 ( .A(n19403), .B(n19401), .Z(n19618) );
  AND U19694 ( .A(n19619), .B(n19620), .Z(n19401) );
  NANDN U19695 ( .A(n19621), .B(n19622), .Z(n19620) );
  NANDN U19696 ( .A(n19623), .B(n19624), .Z(n19622) );
  NANDN U19697 ( .A(n19624), .B(n19623), .Z(n19619) );
  ANDN U19698 ( .B(B[216]), .A(n58), .Z(n19403) );
  XNOR U19699 ( .A(n19411), .B(n19625), .Z(n19404) );
  XNOR U19700 ( .A(n19410), .B(n19408), .Z(n19625) );
  AND U19701 ( .A(n19626), .B(n19627), .Z(n19408) );
  NANDN U19702 ( .A(n19628), .B(n19629), .Z(n19627) );
  OR U19703 ( .A(n19630), .B(n19631), .Z(n19629) );
  NAND U19704 ( .A(n19631), .B(n19630), .Z(n19626) );
  ANDN U19705 ( .B(B[217]), .A(n59), .Z(n19410) );
  XNOR U19706 ( .A(n19418), .B(n19632), .Z(n19411) );
  XNOR U19707 ( .A(n19417), .B(n19415), .Z(n19632) );
  AND U19708 ( .A(n19633), .B(n19634), .Z(n19415) );
  NANDN U19709 ( .A(n19635), .B(n19636), .Z(n19634) );
  NANDN U19710 ( .A(n19637), .B(n19638), .Z(n19636) );
  NANDN U19711 ( .A(n19638), .B(n19637), .Z(n19633) );
  ANDN U19712 ( .B(B[218]), .A(n60), .Z(n19417) );
  XNOR U19713 ( .A(n19425), .B(n19639), .Z(n19418) );
  XNOR U19714 ( .A(n19424), .B(n19422), .Z(n19639) );
  AND U19715 ( .A(n19640), .B(n19641), .Z(n19422) );
  NANDN U19716 ( .A(n19642), .B(n19643), .Z(n19641) );
  OR U19717 ( .A(n19644), .B(n19645), .Z(n19643) );
  NAND U19718 ( .A(n19645), .B(n19644), .Z(n19640) );
  ANDN U19719 ( .B(B[219]), .A(n61), .Z(n19424) );
  XNOR U19720 ( .A(n19432), .B(n19646), .Z(n19425) );
  XNOR U19721 ( .A(n19431), .B(n19429), .Z(n19646) );
  AND U19722 ( .A(n19647), .B(n19648), .Z(n19429) );
  NANDN U19723 ( .A(n19649), .B(n19650), .Z(n19648) );
  NANDN U19724 ( .A(n19651), .B(n19652), .Z(n19650) );
  NANDN U19725 ( .A(n19652), .B(n19651), .Z(n19647) );
  ANDN U19726 ( .B(B[220]), .A(n62), .Z(n19431) );
  XNOR U19727 ( .A(n19439), .B(n19653), .Z(n19432) );
  XNOR U19728 ( .A(n19438), .B(n19436), .Z(n19653) );
  AND U19729 ( .A(n19654), .B(n19655), .Z(n19436) );
  NANDN U19730 ( .A(n19656), .B(n19657), .Z(n19655) );
  OR U19731 ( .A(n19658), .B(n19659), .Z(n19657) );
  NAND U19732 ( .A(n19659), .B(n19658), .Z(n19654) );
  ANDN U19733 ( .B(B[221]), .A(n63), .Z(n19438) );
  XNOR U19734 ( .A(n19446), .B(n19660), .Z(n19439) );
  XNOR U19735 ( .A(n19445), .B(n19443), .Z(n19660) );
  AND U19736 ( .A(n19661), .B(n19662), .Z(n19443) );
  NANDN U19737 ( .A(n19663), .B(n19664), .Z(n19662) );
  NANDN U19738 ( .A(n19665), .B(n19666), .Z(n19664) );
  NANDN U19739 ( .A(n19666), .B(n19665), .Z(n19661) );
  ANDN U19740 ( .B(B[222]), .A(n64), .Z(n19445) );
  XNOR U19741 ( .A(n19453), .B(n19667), .Z(n19446) );
  XNOR U19742 ( .A(n19452), .B(n19450), .Z(n19667) );
  AND U19743 ( .A(n19668), .B(n19669), .Z(n19450) );
  NANDN U19744 ( .A(n19670), .B(n19671), .Z(n19669) );
  OR U19745 ( .A(n19672), .B(n19673), .Z(n19671) );
  NAND U19746 ( .A(n19673), .B(n19672), .Z(n19668) );
  ANDN U19747 ( .B(B[223]), .A(n65), .Z(n19452) );
  XNOR U19748 ( .A(n19460), .B(n19674), .Z(n19453) );
  XNOR U19749 ( .A(n19459), .B(n19457), .Z(n19674) );
  AND U19750 ( .A(n19675), .B(n19676), .Z(n19457) );
  NANDN U19751 ( .A(n19677), .B(n19678), .Z(n19676) );
  NANDN U19752 ( .A(n19679), .B(n19680), .Z(n19678) );
  NANDN U19753 ( .A(n19680), .B(n19679), .Z(n19675) );
  ANDN U19754 ( .B(B[224]), .A(n66), .Z(n19459) );
  XNOR U19755 ( .A(n19467), .B(n19681), .Z(n19460) );
  XNOR U19756 ( .A(n19466), .B(n19464), .Z(n19681) );
  AND U19757 ( .A(n19682), .B(n19683), .Z(n19464) );
  NANDN U19758 ( .A(n19684), .B(n19685), .Z(n19683) );
  OR U19759 ( .A(n19686), .B(n19687), .Z(n19685) );
  NAND U19760 ( .A(n19687), .B(n19686), .Z(n19682) );
  ANDN U19761 ( .B(B[225]), .A(n67), .Z(n19466) );
  XNOR U19762 ( .A(n19474), .B(n19688), .Z(n19467) );
  XNOR U19763 ( .A(n19473), .B(n19471), .Z(n19688) );
  AND U19764 ( .A(n19689), .B(n19690), .Z(n19471) );
  NANDN U19765 ( .A(n19691), .B(n19692), .Z(n19690) );
  NANDN U19766 ( .A(n19693), .B(n19694), .Z(n19692) );
  NANDN U19767 ( .A(n19694), .B(n19693), .Z(n19689) );
  ANDN U19768 ( .B(B[226]), .A(n68), .Z(n19473) );
  XNOR U19769 ( .A(n19481), .B(n19695), .Z(n19474) );
  XNOR U19770 ( .A(n19480), .B(n19478), .Z(n19695) );
  AND U19771 ( .A(n19696), .B(n19697), .Z(n19478) );
  NANDN U19772 ( .A(n19698), .B(n19699), .Z(n19697) );
  OR U19773 ( .A(n19700), .B(n19701), .Z(n19699) );
  NAND U19774 ( .A(n19701), .B(n19700), .Z(n19696) );
  ANDN U19775 ( .B(B[227]), .A(n69), .Z(n19480) );
  XNOR U19776 ( .A(n19488), .B(n19702), .Z(n19481) );
  XNOR U19777 ( .A(n19487), .B(n19485), .Z(n19702) );
  AND U19778 ( .A(n19703), .B(n19704), .Z(n19485) );
  NANDN U19779 ( .A(n19705), .B(n19706), .Z(n19704) );
  NANDN U19780 ( .A(n19707), .B(n19708), .Z(n19706) );
  NANDN U19781 ( .A(n19708), .B(n19707), .Z(n19703) );
  ANDN U19782 ( .B(B[228]), .A(n70), .Z(n19487) );
  XNOR U19783 ( .A(n19495), .B(n19709), .Z(n19488) );
  XNOR U19784 ( .A(n19494), .B(n19492), .Z(n19709) );
  AND U19785 ( .A(n19710), .B(n19711), .Z(n19492) );
  NANDN U19786 ( .A(n19712), .B(n19713), .Z(n19711) );
  OR U19787 ( .A(n19714), .B(n19715), .Z(n19713) );
  NAND U19788 ( .A(n19715), .B(n19714), .Z(n19710) );
  ANDN U19789 ( .B(B[229]), .A(n71), .Z(n19494) );
  XNOR U19790 ( .A(n19502), .B(n19716), .Z(n19495) );
  XNOR U19791 ( .A(n19501), .B(n19499), .Z(n19716) );
  AND U19792 ( .A(n19717), .B(n19718), .Z(n19499) );
  NANDN U19793 ( .A(n19719), .B(n19720), .Z(n19718) );
  NANDN U19794 ( .A(n19721), .B(n19722), .Z(n19720) );
  NANDN U19795 ( .A(n19722), .B(n19721), .Z(n19717) );
  ANDN U19796 ( .B(B[230]), .A(n72), .Z(n19501) );
  XNOR U19797 ( .A(n19509), .B(n19723), .Z(n19502) );
  XNOR U19798 ( .A(n19508), .B(n19506), .Z(n19723) );
  AND U19799 ( .A(n19724), .B(n19725), .Z(n19506) );
  NANDN U19800 ( .A(n19726), .B(n19727), .Z(n19725) );
  OR U19801 ( .A(n19728), .B(n19729), .Z(n19727) );
  NAND U19802 ( .A(n19729), .B(n19728), .Z(n19724) );
  ANDN U19803 ( .B(B[231]), .A(n73), .Z(n19508) );
  XNOR U19804 ( .A(n19516), .B(n19730), .Z(n19509) );
  XNOR U19805 ( .A(n19515), .B(n19513), .Z(n19730) );
  AND U19806 ( .A(n19731), .B(n19732), .Z(n19513) );
  NANDN U19807 ( .A(n19733), .B(n19734), .Z(n19732) );
  NANDN U19808 ( .A(n19735), .B(n19736), .Z(n19734) );
  NANDN U19809 ( .A(n19736), .B(n19735), .Z(n19731) );
  ANDN U19810 ( .B(B[232]), .A(n74), .Z(n19515) );
  XNOR U19811 ( .A(n19523), .B(n19737), .Z(n19516) );
  XNOR U19812 ( .A(n19522), .B(n19520), .Z(n19737) );
  AND U19813 ( .A(n19738), .B(n19739), .Z(n19520) );
  NANDN U19814 ( .A(n19740), .B(n19741), .Z(n19739) );
  OR U19815 ( .A(n19742), .B(n19743), .Z(n19741) );
  NAND U19816 ( .A(n19743), .B(n19742), .Z(n19738) );
  ANDN U19817 ( .B(B[233]), .A(n75), .Z(n19522) );
  XNOR U19818 ( .A(n19530), .B(n19744), .Z(n19523) );
  XNOR U19819 ( .A(n19529), .B(n19527), .Z(n19744) );
  AND U19820 ( .A(n19745), .B(n19746), .Z(n19527) );
  NANDN U19821 ( .A(n19747), .B(n19748), .Z(n19746) );
  NANDN U19822 ( .A(n19749), .B(n19750), .Z(n19748) );
  NANDN U19823 ( .A(n19750), .B(n19749), .Z(n19745) );
  ANDN U19824 ( .B(B[234]), .A(n76), .Z(n19529) );
  XNOR U19825 ( .A(n19537), .B(n19751), .Z(n19530) );
  XNOR U19826 ( .A(n19536), .B(n19534), .Z(n19751) );
  AND U19827 ( .A(n19752), .B(n19753), .Z(n19534) );
  NANDN U19828 ( .A(n19754), .B(n19755), .Z(n19753) );
  OR U19829 ( .A(n19756), .B(n19757), .Z(n19755) );
  NAND U19830 ( .A(n19757), .B(n19756), .Z(n19752) );
  ANDN U19831 ( .B(B[235]), .A(n77), .Z(n19536) );
  XNOR U19832 ( .A(n19544), .B(n19758), .Z(n19537) );
  XNOR U19833 ( .A(n19543), .B(n19541), .Z(n19758) );
  AND U19834 ( .A(n19759), .B(n19760), .Z(n19541) );
  NANDN U19835 ( .A(n19761), .B(n19762), .Z(n19760) );
  NANDN U19836 ( .A(n19763), .B(n19764), .Z(n19762) );
  NANDN U19837 ( .A(n19764), .B(n19763), .Z(n19759) );
  ANDN U19838 ( .B(B[236]), .A(n78), .Z(n19543) );
  XNOR U19839 ( .A(n19551), .B(n19765), .Z(n19544) );
  XNOR U19840 ( .A(n19550), .B(n19548), .Z(n19765) );
  AND U19841 ( .A(n19766), .B(n19767), .Z(n19548) );
  NANDN U19842 ( .A(n19768), .B(n19769), .Z(n19767) );
  OR U19843 ( .A(n19770), .B(n19771), .Z(n19769) );
  NAND U19844 ( .A(n19771), .B(n19770), .Z(n19766) );
  ANDN U19845 ( .B(B[237]), .A(n79), .Z(n19550) );
  XNOR U19846 ( .A(n19558), .B(n19772), .Z(n19551) );
  XNOR U19847 ( .A(n19557), .B(n19555), .Z(n19772) );
  AND U19848 ( .A(n19773), .B(n19774), .Z(n19555) );
  NANDN U19849 ( .A(n19775), .B(n19776), .Z(n19774) );
  NANDN U19850 ( .A(n19777), .B(n19778), .Z(n19776) );
  NANDN U19851 ( .A(n19778), .B(n19777), .Z(n19773) );
  ANDN U19852 ( .B(B[238]), .A(n80), .Z(n19557) );
  XNOR U19853 ( .A(n19565), .B(n19779), .Z(n19558) );
  XNOR U19854 ( .A(n19564), .B(n19562), .Z(n19779) );
  AND U19855 ( .A(n19780), .B(n19781), .Z(n19562) );
  NANDN U19856 ( .A(n19782), .B(n19783), .Z(n19781) );
  OR U19857 ( .A(n19784), .B(n19785), .Z(n19783) );
  NAND U19858 ( .A(n19785), .B(n19784), .Z(n19780) );
  ANDN U19859 ( .B(B[239]), .A(n81), .Z(n19564) );
  XNOR U19860 ( .A(n19572), .B(n19786), .Z(n19565) );
  XNOR U19861 ( .A(n19571), .B(n19569), .Z(n19786) );
  AND U19862 ( .A(n19787), .B(n19788), .Z(n19569) );
  NANDN U19863 ( .A(n19789), .B(n19790), .Z(n19788) );
  NAND U19864 ( .A(n19791), .B(n19792), .Z(n19790) );
  ANDN U19865 ( .B(B[240]), .A(n82), .Z(n19571) );
  XOR U19866 ( .A(n19578), .B(n19793), .Z(n19572) );
  XNOR U19867 ( .A(n19576), .B(n19579), .Z(n19793) );
  NAND U19868 ( .A(A[2]), .B(B[241]), .Z(n19579) );
  NANDN U19869 ( .A(n19794), .B(n19795), .Z(n19576) );
  AND U19870 ( .A(A[0]), .B(B[242]), .Z(n19795) );
  XNOR U19871 ( .A(n19581), .B(n19796), .Z(n19578) );
  NAND U19872 ( .A(A[0]), .B(B[243]), .Z(n19796) );
  NAND U19873 ( .A(B[242]), .B(A[1]), .Z(n19581) );
  NAND U19874 ( .A(n19797), .B(n19798), .Z(n310) );
  NANDN U19875 ( .A(n19799), .B(n19800), .Z(n19798) );
  OR U19876 ( .A(n19801), .B(n19802), .Z(n19800) );
  NAND U19877 ( .A(n19802), .B(n19801), .Z(n19797) );
  XOR U19878 ( .A(n312), .B(n311), .Z(\A1[240] ) );
  XOR U19879 ( .A(n19802), .B(n19803), .Z(n311) );
  XNOR U19880 ( .A(n19801), .B(n19799), .Z(n19803) );
  AND U19881 ( .A(n19804), .B(n19805), .Z(n19799) );
  NANDN U19882 ( .A(n19806), .B(n19807), .Z(n19805) );
  NANDN U19883 ( .A(n19808), .B(n19809), .Z(n19807) );
  NANDN U19884 ( .A(n19809), .B(n19808), .Z(n19804) );
  ANDN U19885 ( .B(B[211]), .A(n54), .Z(n19801) );
  XNOR U19886 ( .A(n19596), .B(n19810), .Z(n19802) );
  XNOR U19887 ( .A(n19595), .B(n19593), .Z(n19810) );
  AND U19888 ( .A(n19811), .B(n19812), .Z(n19593) );
  NANDN U19889 ( .A(n19813), .B(n19814), .Z(n19812) );
  OR U19890 ( .A(n19815), .B(n19816), .Z(n19814) );
  NAND U19891 ( .A(n19816), .B(n19815), .Z(n19811) );
  ANDN U19892 ( .B(B[212]), .A(n55), .Z(n19595) );
  XNOR U19893 ( .A(n19603), .B(n19817), .Z(n19596) );
  XNOR U19894 ( .A(n19602), .B(n19600), .Z(n19817) );
  AND U19895 ( .A(n19818), .B(n19819), .Z(n19600) );
  NANDN U19896 ( .A(n19820), .B(n19821), .Z(n19819) );
  NANDN U19897 ( .A(n19822), .B(n19823), .Z(n19821) );
  NANDN U19898 ( .A(n19823), .B(n19822), .Z(n19818) );
  ANDN U19899 ( .B(B[213]), .A(n56), .Z(n19602) );
  XNOR U19900 ( .A(n19610), .B(n19824), .Z(n19603) );
  XNOR U19901 ( .A(n19609), .B(n19607), .Z(n19824) );
  AND U19902 ( .A(n19825), .B(n19826), .Z(n19607) );
  NANDN U19903 ( .A(n19827), .B(n19828), .Z(n19826) );
  OR U19904 ( .A(n19829), .B(n19830), .Z(n19828) );
  NAND U19905 ( .A(n19830), .B(n19829), .Z(n19825) );
  ANDN U19906 ( .B(B[214]), .A(n57), .Z(n19609) );
  XNOR U19907 ( .A(n19617), .B(n19831), .Z(n19610) );
  XNOR U19908 ( .A(n19616), .B(n19614), .Z(n19831) );
  AND U19909 ( .A(n19832), .B(n19833), .Z(n19614) );
  NANDN U19910 ( .A(n19834), .B(n19835), .Z(n19833) );
  NANDN U19911 ( .A(n19836), .B(n19837), .Z(n19835) );
  NANDN U19912 ( .A(n19837), .B(n19836), .Z(n19832) );
  ANDN U19913 ( .B(B[215]), .A(n58), .Z(n19616) );
  XNOR U19914 ( .A(n19624), .B(n19838), .Z(n19617) );
  XNOR U19915 ( .A(n19623), .B(n19621), .Z(n19838) );
  AND U19916 ( .A(n19839), .B(n19840), .Z(n19621) );
  NANDN U19917 ( .A(n19841), .B(n19842), .Z(n19840) );
  OR U19918 ( .A(n19843), .B(n19844), .Z(n19842) );
  NAND U19919 ( .A(n19844), .B(n19843), .Z(n19839) );
  ANDN U19920 ( .B(B[216]), .A(n59), .Z(n19623) );
  XNOR U19921 ( .A(n19631), .B(n19845), .Z(n19624) );
  XNOR U19922 ( .A(n19630), .B(n19628), .Z(n19845) );
  AND U19923 ( .A(n19846), .B(n19847), .Z(n19628) );
  NANDN U19924 ( .A(n19848), .B(n19849), .Z(n19847) );
  NANDN U19925 ( .A(n19850), .B(n19851), .Z(n19849) );
  NANDN U19926 ( .A(n19851), .B(n19850), .Z(n19846) );
  ANDN U19927 ( .B(B[217]), .A(n60), .Z(n19630) );
  XNOR U19928 ( .A(n19638), .B(n19852), .Z(n19631) );
  XNOR U19929 ( .A(n19637), .B(n19635), .Z(n19852) );
  AND U19930 ( .A(n19853), .B(n19854), .Z(n19635) );
  NANDN U19931 ( .A(n19855), .B(n19856), .Z(n19854) );
  OR U19932 ( .A(n19857), .B(n19858), .Z(n19856) );
  NAND U19933 ( .A(n19858), .B(n19857), .Z(n19853) );
  ANDN U19934 ( .B(B[218]), .A(n61), .Z(n19637) );
  XNOR U19935 ( .A(n19645), .B(n19859), .Z(n19638) );
  XNOR U19936 ( .A(n19644), .B(n19642), .Z(n19859) );
  AND U19937 ( .A(n19860), .B(n19861), .Z(n19642) );
  NANDN U19938 ( .A(n19862), .B(n19863), .Z(n19861) );
  NANDN U19939 ( .A(n19864), .B(n19865), .Z(n19863) );
  NANDN U19940 ( .A(n19865), .B(n19864), .Z(n19860) );
  ANDN U19941 ( .B(B[219]), .A(n62), .Z(n19644) );
  XNOR U19942 ( .A(n19652), .B(n19866), .Z(n19645) );
  XNOR U19943 ( .A(n19651), .B(n19649), .Z(n19866) );
  AND U19944 ( .A(n19867), .B(n19868), .Z(n19649) );
  NANDN U19945 ( .A(n19869), .B(n19870), .Z(n19868) );
  OR U19946 ( .A(n19871), .B(n19872), .Z(n19870) );
  NAND U19947 ( .A(n19872), .B(n19871), .Z(n19867) );
  ANDN U19948 ( .B(B[220]), .A(n63), .Z(n19651) );
  XNOR U19949 ( .A(n19659), .B(n19873), .Z(n19652) );
  XNOR U19950 ( .A(n19658), .B(n19656), .Z(n19873) );
  AND U19951 ( .A(n19874), .B(n19875), .Z(n19656) );
  NANDN U19952 ( .A(n19876), .B(n19877), .Z(n19875) );
  NANDN U19953 ( .A(n19878), .B(n19879), .Z(n19877) );
  NANDN U19954 ( .A(n19879), .B(n19878), .Z(n19874) );
  ANDN U19955 ( .B(B[221]), .A(n64), .Z(n19658) );
  XNOR U19956 ( .A(n19666), .B(n19880), .Z(n19659) );
  XNOR U19957 ( .A(n19665), .B(n19663), .Z(n19880) );
  AND U19958 ( .A(n19881), .B(n19882), .Z(n19663) );
  NANDN U19959 ( .A(n19883), .B(n19884), .Z(n19882) );
  OR U19960 ( .A(n19885), .B(n19886), .Z(n19884) );
  NAND U19961 ( .A(n19886), .B(n19885), .Z(n19881) );
  ANDN U19962 ( .B(B[222]), .A(n65), .Z(n19665) );
  XNOR U19963 ( .A(n19673), .B(n19887), .Z(n19666) );
  XNOR U19964 ( .A(n19672), .B(n19670), .Z(n19887) );
  AND U19965 ( .A(n19888), .B(n19889), .Z(n19670) );
  NANDN U19966 ( .A(n19890), .B(n19891), .Z(n19889) );
  NANDN U19967 ( .A(n19892), .B(n19893), .Z(n19891) );
  NANDN U19968 ( .A(n19893), .B(n19892), .Z(n19888) );
  ANDN U19969 ( .B(B[223]), .A(n66), .Z(n19672) );
  XNOR U19970 ( .A(n19680), .B(n19894), .Z(n19673) );
  XNOR U19971 ( .A(n19679), .B(n19677), .Z(n19894) );
  AND U19972 ( .A(n19895), .B(n19896), .Z(n19677) );
  NANDN U19973 ( .A(n19897), .B(n19898), .Z(n19896) );
  OR U19974 ( .A(n19899), .B(n19900), .Z(n19898) );
  NAND U19975 ( .A(n19900), .B(n19899), .Z(n19895) );
  ANDN U19976 ( .B(B[224]), .A(n67), .Z(n19679) );
  XNOR U19977 ( .A(n19687), .B(n19901), .Z(n19680) );
  XNOR U19978 ( .A(n19686), .B(n19684), .Z(n19901) );
  AND U19979 ( .A(n19902), .B(n19903), .Z(n19684) );
  NANDN U19980 ( .A(n19904), .B(n19905), .Z(n19903) );
  NANDN U19981 ( .A(n19906), .B(n19907), .Z(n19905) );
  NANDN U19982 ( .A(n19907), .B(n19906), .Z(n19902) );
  ANDN U19983 ( .B(B[225]), .A(n68), .Z(n19686) );
  XNOR U19984 ( .A(n19694), .B(n19908), .Z(n19687) );
  XNOR U19985 ( .A(n19693), .B(n19691), .Z(n19908) );
  AND U19986 ( .A(n19909), .B(n19910), .Z(n19691) );
  NANDN U19987 ( .A(n19911), .B(n19912), .Z(n19910) );
  OR U19988 ( .A(n19913), .B(n19914), .Z(n19912) );
  NAND U19989 ( .A(n19914), .B(n19913), .Z(n19909) );
  ANDN U19990 ( .B(B[226]), .A(n69), .Z(n19693) );
  XNOR U19991 ( .A(n19701), .B(n19915), .Z(n19694) );
  XNOR U19992 ( .A(n19700), .B(n19698), .Z(n19915) );
  AND U19993 ( .A(n19916), .B(n19917), .Z(n19698) );
  NANDN U19994 ( .A(n19918), .B(n19919), .Z(n19917) );
  NANDN U19995 ( .A(n19920), .B(n19921), .Z(n19919) );
  NANDN U19996 ( .A(n19921), .B(n19920), .Z(n19916) );
  ANDN U19997 ( .B(B[227]), .A(n70), .Z(n19700) );
  XNOR U19998 ( .A(n19708), .B(n19922), .Z(n19701) );
  XNOR U19999 ( .A(n19707), .B(n19705), .Z(n19922) );
  AND U20000 ( .A(n19923), .B(n19924), .Z(n19705) );
  NANDN U20001 ( .A(n19925), .B(n19926), .Z(n19924) );
  OR U20002 ( .A(n19927), .B(n19928), .Z(n19926) );
  NAND U20003 ( .A(n19928), .B(n19927), .Z(n19923) );
  ANDN U20004 ( .B(B[228]), .A(n71), .Z(n19707) );
  XNOR U20005 ( .A(n19715), .B(n19929), .Z(n19708) );
  XNOR U20006 ( .A(n19714), .B(n19712), .Z(n19929) );
  AND U20007 ( .A(n19930), .B(n19931), .Z(n19712) );
  NANDN U20008 ( .A(n19932), .B(n19933), .Z(n19931) );
  NANDN U20009 ( .A(n19934), .B(n19935), .Z(n19933) );
  NANDN U20010 ( .A(n19935), .B(n19934), .Z(n19930) );
  ANDN U20011 ( .B(B[229]), .A(n72), .Z(n19714) );
  XNOR U20012 ( .A(n19722), .B(n19936), .Z(n19715) );
  XNOR U20013 ( .A(n19721), .B(n19719), .Z(n19936) );
  AND U20014 ( .A(n19937), .B(n19938), .Z(n19719) );
  NANDN U20015 ( .A(n19939), .B(n19940), .Z(n19938) );
  OR U20016 ( .A(n19941), .B(n19942), .Z(n19940) );
  NAND U20017 ( .A(n19942), .B(n19941), .Z(n19937) );
  ANDN U20018 ( .B(B[230]), .A(n73), .Z(n19721) );
  XNOR U20019 ( .A(n19729), .B(n19943), .Z(n19722) );
  XNOR U20020 ( .A(n19728), .B(n19726), .Z(n19943) );
  AND U20021 ( .A(n19944), .B(n19945), .Z(n19726) );
  NANDN U20022 ( .A(n19946), .B(n19947), .Z(n19945) );
  NANDN U20023 ( .A(n19948), .B(n19949), .Z(n19947) );
  NANDN U20024 ( .A(n19949), .B(n19948), .Z(n19944) );
  ANDN U20025 ( .B(B[231]), .A(n74), .Z(n19728) );
  XNOR U20026 ( .A(n19736), .B(n19950), .Z(n19729) );
  XNOR U20027 ( .A(n19735), .B(n19733), .Z(n19950) );
  AND U20028 ( .A(n19951), .B(n19952), .Z(n19733) );
  NANDN U20029 ( .A(n19953), .B(n19954), .Z(n19952) );
  OR U20030 ( .A(n19955), .B(n19956), .Z(n19954) );
  NAND U20031 ( .A(n19956), .B(n19955), .Z(n19951) );
  ANDN U20032 ( .B(B[232]), .A(n75), .Z(n19735) );
  XNOR U20033 ( .A(n19743), .B(n19957), .Z(n19736) );
  XNOR U20034 ( .A(n19742), .B(n19740), .Z(n19957) );
  AND U20035 ( .A(n19958), .B(n19959), .Z(n19740) );
  NANDN U20036 ( .A(n19960), .B(n19961), .Z(n19959) );
  NANDN U20037 ( .A(n19962), .B(n19963), .Z(n19961) );
  NANDN U20038 ( .A(n19963), .B(n19962), .Z(n19958) );
  ANDN U20039 ( .B(B[233]), .A(n76), .Z(n19742) );
  XNOR U20040 ( .A(n19750), .B(n19964), .Z(n19743) );
  XNOR U20041 ( .A(n19749), .B(n19747), .Z(n19964) );
  AND U20042 ( .A(n19965), .B(n19966), .Z(n19747) );
  NANDN U20043 ( .A(n19967), .B(n19968), .Z(n19966) );
  OR U20044 ( .A(n19969), .B(n19970), .Z(n19968) );
  NAND U20045 ( .A(n19970), .B(n19969), .Z(n19965) );
  ANDN U20046 ( .B(B[234]), .A(n77), .Z(n19749) );
  XNOR U20047 ( .A(n19757), .B(n19971), .Z(n19750) );
  XNOR U20048 ( .A(n19756), .B(n19754), .Z(n19971) );
  AND U20049 ( .A(n19972), .B(n19973), .Z(n19754) );
  NANDN U20050 ( .A(n19974), .B(n19975), .Z(n19973) );
  NANDN U20051 ( .A(n19976), .B(n19977), .Z(n19975) );
  NANDN U20052 ( .A(n19977), .B(n19976), .Z(n19972) );
  ANDN U20053 ( .B(B[235]), .A(n78), .Z(n19756) );
  XNOR U20054 ( .A(n19764), .B(n19978), .Z(n19757) );
  XNOR U20055 ( .A(n19763), .B(n19761), .Z(n19978) );
  AND U20056 ( .A(n19979), .B(n19980), .Z(n19761) );
  NANDN U20057 ( .A(n19981), .B(n19982), .Z(n19980) );
  OR U20058 ( .A(n19983), .B(n19984), .Z(n19982) );
  NAND U20059 ( .A(n19984), .B(n19983), .Z(n19979) );
  ANDN U20060 ( .B(B[236]), .A(n79), .Z(n19763) );
  XNOR U20061 ( .A(n19771), .B(n19985), .Z(n19764) );
  XNOR U20062 ( .A(n19770), .B(n19768), .Z(n19985) );
  AND U20063 ( .A(n19986), .B(n19987), .Z(n19768) );
  NANDN U20064 ( .A(n19988), .B(n19989), .Z(n19987) );
  NANDN U20065 ( .A(n19990), .B(n19991), .Z(n19989) );
  NANDN U20066 ( .A(n19991), .B(n19990), .Z(n19986) );
  ANDN U20067 ( .B(B[237]), .A(n80), .Z(n19770) );
  XNOR U20068 ( .A(n19778), .B(n19992), .Z(n19771) );
  XNOR U20069 ( .A(n19777), .B(n19775), .Z(n19992) );
  AND U20070 ( .A(n19993), .B(n19994), .Z(n19775) );
  NANDN U20071 ( .A(n19995), .B(n19996), .Z(n19994) );
  OR U20072 ( .A(n19997), .B(n19998), .Z(n19996) );
  NAND U20073 ( .A(n19998), .B(n19997), .Z(n19993) );
  ANDN U20074 ( .B(B[238]), .A(n81), .Z(n19777) );
  XNOR U20075 ( .A(n19785), .B(n19999), .Z(n19778) );
  XNOR U20076 ( .A(n19784), .B(n19782), .Z(n19999) );
  AND U20077 ( .A(n20000), .B(n20001), .Z(n19782) );
  NANDN U20078 ( .A(n20002), .B(n20003), .Z(n20001) );
  NAND U20079 ( .A(n20004), .B(n20005), .Z(n20003) );
  ANDN U20080 ( .B(B[239]), .A(n82), .Z(n19784) );
  XOR U20081 ( .A(n19791), .B(n20006), .Z(n19785) );
  XNOR U20082 ( .A(n19789), .B(n19792), .Z(n20006) );
  NAND U20083 ( .A(A[2]), .B(B[240]), .Z(n19792) );
  NANDN U20084 ( .A(n20007), .B(n20008), .Z(n19789) );
  AND U20085 ( .A(A[0]), .B(B[241]), .Z(n20008) );
  XNOR U20086 ( .A(n19794), .B(n20009), .Z(n19791) );
  NAND U20087 ( .A(A[0]), .B(B[242]), .Z(n20009) );
  NAND U20088 ( .A(B[241]), .B(A[1]), .Z(n19794) );
  NAND U20089 ( .A(n20010), .B(n20011), .Z(n312) );
  NANDN U20090 ( .A(n20012), .B(n20013), .Z(n20011) );
  OR U20091 ( .A(n20014), .B(n20015), .Z(n20013) );
  NAND U20092 ( .A(n20015), .B(n20014), .Z(n20010) );
  XOR U20093 ( .A(n17720), .B(n20016), .Z(\A1[23] ) );
  XNOR U20094 ( .A(n17719), .B(n17717), .Z(n20016) );
  AND U20095 ( .A(n20017), .B(n20018), .Z(n17717) );
  NAND U20096 ( .A(n20019), .B(n20020), .Z(n20018) );
  NANDN U20097 ( .A(n20021), .B(n20022), .Z(n20019) );
  NANDN U20098 ( .A(n20022), .B(n20021), .Z(n20017) );
  ANDN U20099 ( .B(B[0]), .A(n60), .Z(n17719) );
  XNOR U20100 ( .A(n17727), .B(n20023), .Z(n17720) );
  XNOR U20101 ( .A(n17726), .B(n17724), .Z(n20023) );
  AND U20102 ( .A(n20024), .B(n20025), .Z(n17724) );
  NANDN U20103 ( .A(n20026), .B(n20027), .Z(n20025) );
  OR U20104 ( .A(n20028), .B(n20029), .Z(n20027) );
  NAND U20105 ( .A(n20029), .B(n20028), .Z(n20024) );
  ANDN U20106 ( .B(B[1]), .A(n61), .Z(n17726) );
  XNOR U20107 ( .A(n17734), .B(n20030), .Z(n17727) );
  XNOR U20108 ( .A(n17733), .B(n17731), .Z(n20030) );
  AND U20109 ( .A(n20031), .B(n20032), .Z(n17731) );
  NANDN U20110 ( .A(n20033), .B(n20034), .Z(n20032) );
  NANDN U20111 ( .A(n20035), .B(n20036), .Z(n20034) );
  NANDN U20112 ( .A(n20036), .B(n20035), .Z(n20031) );
  ANDN U20113 ( .B(B[2]), .A(n62), .Z(n17733) );
  XNOR U20114 ( .A(n17741), .B(n20037), .Z(n17734) );
  XNOR U20115 ( .A(n17740), .B(n17738), .Z(n20037) );
  AND U20116 ( .A(n20038), .B(n20039), .Z(n17738) );
  NANDN U20117 ( .A(n20040), .B(n20041), .Z(n20039) );
  OR U20118 ( .A(n20042), .B(n20043), .Z(n20041) );
  NAND U20119 ( .A(n20043), .B(n20042), .Z(n20038) );
  ANDN U20120 ( .B(B[3]), .A(n63), .Z(n17740) );
  XNOR U20121 ( .A(n17748), .B(n20044), .Z(n17741) );
  XNOR U20122 ( .A(n17747), .B(n17745), .Z(n20044) );
  AND U20123 ( .A(n20045), .B(n20046), .Z(n17745) );
  NANDN U20124 ( .A(n20047), .B(n20048), .Z(n20046) );
  NANDN U20125 ( .A(n20049), .B(n20050), .Z(n20048) );
  NANDN U20126 ( .A(n20050), .B(n20049), .Z(n20045) );
  ANDN U20127 ( .B(B[4]), .A(n64), .Z(n17747) );
  XNOR U20128 ( .A(n17755), .B(n20051), .Z(n17748) );
  XNOR U20129 ( .A(n17754), .B(n17752), .Z(n20051) );
  AND U20130 ( .A(n20052), .B(n20053), .Z(n17752) );
  NANDN U20131 ( .A(n20054), .B(n20055), .Z(n20053) );
  OR U20132 ( .A(n20056), .B(n20057), .Z(n20055) );
  NAND U20133 ( .A(n20057), .B(n20056), .Z(n20052) );
  ANDN U20134 ( .B(B[5]), .A(n65), .Z(n17754) );
  XNOR U20135 ( .A(n17762), .B(n20058), .Z(n17755) );
  XNOR U20136 ( .A(n17761), .B(n17759), .Z(n20058) );
  AND U20137 ( .A(n20059), .B(n20060), .Z(n17759) );
  NANDN U20138 ( .A(n20061), .B(n20062), .Z(n20060) );
  NANDN U20139 ( .A(n20063), .B(n20064), .Z(n20062) );
  NANDN U20140 ( .A(n20064), .B(n20063), .Z(n20059) );
  ANDN U20141 ( .B(B[6]), .A(n66), .Z(n17761) );
  XNOR U20142 ( .A(n17769), .B(n20065), .Z(n17762) );
  XNOR U20143 ( .A(n17768), .B(n17766), .Z(n20065) );
  AND U20144 ( .A(n20066), .B(n20067), .Z(n17766) );
  NANDN U20145 ( .A(n20068), .B(n20069), .Z(n20067) );
  OR U20146 ( .A(n20070), .B(n20071), .Z(n20069) );
  NAND U20147 ( .A(n20071), .B(n20070), .Z(n20066) );
  ANDN U20148 ( .B(B[7]), .A(n67), .Z(n17768) );
  XNOR U20149 ( .A(n17776), .B(n20072), .Z(n17769) );
  XNOR U20150 ( .A(n17775), .B(n17773), .Z(n20072) );
  AND U20151 ( .A(n20073), .B(n20074), .Z(n17773) );
  NANDN U20152 ( .A(n20075), .B(n20076), .Z(n20074) );
  NANDN U20153 ( .A(n20077), .B(n20078), .Z(n20076) );
  NANDN U20154 ( .A(n20078), .B(n20077), .Z(n20073) );
  ANDN U20155 ( .B(B[8]), .A(n68), .Z(n17775) );
  XNOR U20156 ( .A(n17783), .B(n20079), .Z(n17776) );
  XNOR U20157 ( .A(n17782), .B(n17780), .Z(n20079) );
  AND U20158 ( .A(n20080), .B(n20081), .Z(n17780) );
  NANDN U20159 ( .A(n20082), .B(n20083), .Z(n20081) );
  OR U20160 ( .A(n20084), .B(n20085), .Z(n20083) );
  NAND U20161 ( .A(n20085), .B(n20084), .Z(n20080) );
  ANDN U20162 ( .B(B[9]), .A(n69), .Z(n17782) );
  XNOR U20163 ( .A(n17790), .B(n20086), .Z(n17783) );
  XNOR U20164 ( .A(n17789), .B(n17787), .Z(n20086) );
  AND U20165 ( .A(n20087), .B(n20088), .Z(n17787) );
  NANDN U20166 ( .A(n20089), .B(n20090), .Z(n20088) );
  NANDN U20167 ( .A(n20091), .B(n20092), .Z(n20090) );
  NANDN U20168 ( .A(n20092), .B(n20091), .Z(n20087) );
  ANDN U20169 ( .B(B[10]), .A(n70), .Z(n17789) );
  XNOR U20170 ( .A(n17797), .B(n20093), .Z(n17790) );
  XNOR U20171 ( .A(n17796), .B(n17794), .Z(n20093) );
  AND U20172 ( .A(n20094), .B(n20095), .Z(n17794) );
  NANDN U20173 ( .A(n20096), .B(n20097), .Z(n20095) );
  OR U20174 ( .A(n20098), .B(n20099), .Z(n20097) );
  NAND U20175 ( .A(n20099), .B(n20098), .Z(n20094) );
  ANDN U20176 ( .B(B[11]), .A(n71), .Z(n17796) );
  XNOR U20177 ( .A(n17804), .B(n20100), .Z(n17797) );
  XNOR U20178 ( .A(n17803), .B(n17801), .Z(n20100) );
  AND U20179 ( .A(n20101), .B(n20102), .Z(n17801) );
  NANDN U20180 ( .A(n20103), .B(n20104), .Z(n20102) );
  NANDN U20181 ( .A(n20105), .B(n20106), .Z(n20104) );
  NANDN U20182 ( .A(n20106), .B(n20105), .Z(n20101) );
  ANDN U20183 ( .B(B[12]), .A(n72), .Z(n17803) );
  XNOR U20184 ( .A(n17811), .B(n20107), .Z(n17804) );
  XNOR U20185 ( .A(n17810), .B(n17808), .Z(n20107) );
  AND U20186 ( .A(n20108), .B(n20109), .Z(n17808) );
  NANDN U20187 ( .A(n20110), .B(n20111), .Z(n20109) );
  OR U20188 ( .A(n20112), .B(n20113), .Z(n20111) );
  NAND U20189 ( .A(n20113), .B(n20112), .Z(n20108) );
  ANDN U20190 ( .B(B[13]), .A(n73), .Z(n17810) );
  XNOR U20191 ( .A(n17818), .B(n20114), .Z(n17811) );
  XNOR U20192 ( .A(n17817), .B(n17815), .Z(n20114) );
  AND U20193 ( .A(n20115), .B(n20116), .Z(n17815) );
  NANDN U20194 ( .A(n20117), .B(n20118), .Z(n20116) );
  NANDN U20195 ( .A(n20119), .B(n20120), .Z(n20118) );
  NANDN U20196 ( .A(n20120), .B(n20119), .Z(n20115) );
  ANDN U20197 ( .B(B[14]), .A(n74), .Z(n17817) );
  XNOR U20198 ( .A(n17825), .B(n20121), .Z(n17818) );
  XNOR U20199 ( .A(n17824), .B(n17822), .Z(n20121) );
  AND U20200 ( .A(n20122), .B(n20123), .Z(n17822) );
  NANDN U20201 ( .A(n20124), .B(n20125), .Z(n20123) );
  OR U20202 ( .A(n20126), .B(n20127), .Z(n20125) );
  NAND U20203 ( .A(n20127), .B(n20126), .Z(n20122) );
  ANDN U20204 ( .B(B[15]), .A(n75), .Z(n17824) );
  XNOR U20205 ( .A(n17832), .B(n20128), .Z(n17825) );
  XNOR U20206 ( .A(n17831), .B(n17829), .Z(n20128) );
  AND U20207 ( .A(n20129), .B(n20130), .Z(n17829) );
  NANDN U20208 ( .A(n20131), .B(n20132), .Z(n20130) );
  NANDN U20209 ( .A(n20133), .B(n20134), .Z(n20132) );
  NANDN U20210 ( .A(n20134), .B(n20133), .Z(n20129) );
  ANDN U20211 ( .B(B[16]), .A(n76), .Z(n17831) );
  XNOR U20212 ( .A(n17839), .B(n20135), .Z(n17832) );
  XNOR U20213 ( .A(n17838), .B(n17836), .Z(n20135) );
  AND U20214 ( .A(n20136), .B(n20137), .Z(n17836) );
  NANDN U20215 ( .A(n20138), .B(n20139), .Z(n20137) );
  OR U20216 ( .A(n20140), .B(n20141), .Z(n20139) );
  NAND U20217 ( .A(n20141), .B(n20140), .Z(n20136) );
  ANDN U20218 ( .B(B[17]), .A(n77), .Z(n17838) );
  XNOR U20219 ( .A(n17846), .B(n20142), .Z(n17839) );
  XNOR U20220 ( .A(n17845), .B(n17843), .Z(n20142) );
  AND U20221 ( .A(n20143), .B(n20144), .Z(n17843) );
  NANDN U20222 ( .A(n20145), .B(n20146), .Z(n20144) );
  NANDN U20223 ( .A(n20147), .B(n20148), .Z(n20146) );
  NANDN U20224 ( .A(n20148), .B(n20147), .Z(n20143) );
  ANDN U20225 ( .B(B[18]), .A(n78), .Z(n17845) );
  XNOR U20226 ( .A(n17853), .B(n20149), .Z(n17846) );
  XNOR U20227 ( .A(n17852), .B(n17850), .Z(n20149) );
  AND U20228 ( .A(n20150), .B(n20151), .Z(n17850) );
  NANDN U20229 ( .A(n20152), .B(n20153), .Z(n20151) );
  OR U20230 ( .A(n20154), .B(n20155), .Z(n20153) );
  NAND U20231 ( .A(n20155), .B(n20154), .Z(n20150) );
  ANDN U20232 ( .B(B[19]), .A(n79), .Z(n17852) );
  XNOR U20233 ( .A(n17860), .B(n20156), .Z(n17853) );
  XNOR U20234 ( .A(n17859), .B(n17857), .Z(n20156) );
  AND U20235 ( .A(n20157), .B(n20158), .Z(n17857) );
  NANDN U20236 ( .A(n20159), .B(n20160), .Z(n20158) );
  NANDN U20237 ( .A(n20161), .B(n20162), .Z(n20160) );
  NANDN U20238 ( .A(n20162), .B(n20161), .Z(n20157) );
  ANDN U20239 ( .B(B[20]), .A(n80), .Z(n17859) );
  XNOR U20240 ( .A(n17867), .B(n20163), .Z(n17860) );
  XNOR U20241 ( .A(n17866), .B(n17864), .Z(n20163) );
  AND U20242 ( .A(n20164), .B(n20165), .Z(n17864) );
  NANDN U20243 ( .A(n20166), .B(n20167), .Z(n20165) );
  OR U20244 ( .A(n20168), .B(n20169), .Z(n20167) );
  NAND U20245 ( .A(n20169), .B(n20168), .Z(n20164) );
  ANDN U20246 ( .B(B[21]), .A(n81), .Z(n17866) );
  XNOR U20247 ( .A(n17874), .B(n20170), .Z(n17867) );
  XNOR U20248 ( .A(n17873), .B(n17871), .Z(n20170) );
  AND U20249 ( .A(n20171), .B(n20172), .Z(n17871) );
  NANDN U20250 ( .A(n20173), .B(n20174), .Z(n20172) );
  NAND U20251 ( .A(n20175), .B(n20176), .Z(n20174) );
  ANDN U20252 ( .B(B[22]), .A(n82), .Z(n17873) );
  XOR U20253 ( .A(n17880), .B(n20177), .Z(n17874) );
  XNOR U20254 ( .A(n17878), .B(n17881), .Z(n20177) );
  NAND U20255 ( .A(A[2]), .B(B[23]), .Z(n17881) );
  NANDN U20256 ( .A(n20178), .B(n20179), .Z(n17878) );
  AND U20257 ( .A(A[0]), .B(B[24]), .Z(n20179) );
  XNOR U20258 ( .A(n17883), .B(n20180), .Z(n17880) );
  NAND U20259 ( .A(A[0]), .B(B[25]), .Z(n20180) );
  NAND U20260 ( .A(B[24]), .B(A[1]), .Z(n17883) );
  XOR U20261 ( .A(n314), .B(n313), .Z(\A1[239] ) );
  XOR U20262 ( .A(n20015), .B(n20181), .Z(n313) );
  XNOR U20263 ( .A(n20014), .B(n20012), .Z(n20181) );
  AND U20264 ( .A(n20182), .B(n20183), .Z(n20012) );
  NANDN U20265 ( .A(n20184), .B(n20185), .Z(n20183) );
  NANDN U20266 ( .A(n20186), .B(n20187), .Z(n20185) );
  NANDN U20267 ( .A(n20187), .B(n20186), .Z(n20182) );
  ANDN U20268 ( .B(B[210]), .A(n54), .Z(n20014) );
  XNOR U20269 ( .A(n19809), .B(n20188), .Z(n20015) );
  XNOR U20270 ( .A(n19808), .B(n19806), .Z(n20188) );
  AND U20271 ( .A(n20189), .B(n20190), .Z(n19806) );
  NANDN U20272 ( .A(n20191), .B(n20192), .Z(n20190) );
  OR U20273 ( .A(n20193), .B(n20194), .Z(n20192) );
  NAND U20274 ( .A(n20194), .B(n20193), .Z(n20189) );
  ANDN U20275 ( .B(B[211]), .A(n55), .Z(n19808) );
  XNOR U20276 ( .A(n19816), .B(n20195), .Z(n19809) );
  XNOR U20277 ( .A(n19815), .B(n19813), .Z(n20195) );
  AND U20278 ( .A(n20196), .B(n20197), .Z(n19813) );
  NANDN U20279 ( .A(n20198), .B(n20199), .Z(n20197) );
  NANDN U20280 ( .A(n20200), .B(n20201), .Z(n20199) );
  NANDN U20281 ( .A(n20201), .B(n20200), .Z(n20196) );
  ANDN U20282 ( .B(B[212]), .A(n56), .Z(n19815) );
  XNOR U20283 ( .A(n19823), .B(n20202), .Z(n19816) );
  XNOR U20284 ( .A(n19822), .B(n19820), .Z(n20202) );
  AND U20285 ( .A(n20203), .B(n20204), .Z(n19820) );
  NANDN U20286 ( .A(n20205), .B(n20206), .Z(n20204) );
  OR U20287 ( .A(n20207), .B(n20208), .Z(n20206) );
  NAND U20288 ( .A(n20208), .B(n20207), .Z(n20203) );
  ANDN U20289 ( .B(B[213]), .A(n57), .Z(n19822) );
  XNOR U20290 ( .A(n19830), .B(n20209), .Z(n19823) );
  XNOR U20291 ( .A(n19829), .B(n19827), .Z(n20209) );
  AND U20292 ( .A(n20210), .B(n20211), .Z(n19827) );
  NANDN U20293 ( .A(n20212), .B(n20213), .Z(n20211) );
  NANDN U20294 ( .A(n20214), .B(n20215), .Z(n20213) );
  NANDN U20295 ( .A(n20215), .B(n20214), .Z(n20210) );
  ANDN U20296 ( .B(B[214]), .A(n58), .Z(n19829) );
  XNOR U20297 ( .A(n19837), .B(n20216), .Z(n19830) );
  XNOR U20298 ( .A(n19836), .B(n19834), .Z(n20216) );
  AND U20299 ( .A(n20217), .B(n20218), .Z(n19834) );
  NANDN U20300 ( .A(n20219), .B(n20220), .Z(n20218) );
  OR U20301 ( .A(n20221), .B(n20222), .Z(n20220) );
  NAND U20302 ( .A(n20222), .B(n20221), .Z(n20217) );
  ANDN U20303 ( .B(B[215]), .A(n59), .Z(n19836) );
  XNOR U20304 ( .A(n19844), .B(n20223), .Z(n19837) );
  XNOR U20305 ( .A(n19843), .B(n19841), .Z(n20223) );
  AND U20306 ( .A(n20224), .B(n20225), .Z(n19841) );
  NANDN U20307 ( .A(n20226), .B(n20227), .Z(n20225) );
  NANDN U20308 ( .A(n20228), .B(n20229), .Z(n20227) );
  NANDN U20309 ( .A(n20229), .B(n20228), .Z(n20224) );
  ANDN U20310 ( .B(B[216]), .A(n60), .Z(n19843) );
  XNOR U20311 ( .A(n19851), .B(n20230), .Z(n19844) );
  XNOR U20312 ( .A(n19850), .B(n19848), .Z(n20230) );
  AND U20313 ( .A(n20231), .B(n20232), .Z(n19848) );
  NANDN U20314 ( .A(n20233), .B(n20234), .Z(n20232) );
  OR U20315 ( .A(n20235), .B(n20236), .Z(n20234) );
  NAND U20316 ( .A(n20236), .B(n20235), .Z(n20231) );
  ANDN U20317 ( .B(B[217]), .A(n61), .Z(n19850) );
  XNOR U20318 ( .A(n19858), .B(n20237), .Z(n19851) );
  XNOR U20319 ( .A(n19857), .B(n19855), .Z(n20237) );
  AND U20320 ( .A(n20238), .B(n20239), .Z(n19855) );
  NANDN U20321 ( .A(n20240), .B(n20241), .Z(n20239) );
  NANDN U20322 ( .A(n20242), .B(n20243), .Z(n20241) );
  NANDN U20323 ( .A(n20243), .B(n20242), .Z(n20238) );
  ANDN U20324 ( .B(B[218]), .A(n62), .Z(n19857) );
  XNOR U20325 ( .A(n19865), .B(n20244), .Z(n19858) );
  XNOR U20326 ( .A(n19864), .B(n19862), .Z(n20244) );
  AND U20327 ( .A(n20245), .B(n20246), .Z(n19862) );
  NANDN U20328 ( .A(n20247), .B(n20248), .Z(n20246) );
  OR U20329 ( .A(n20249), .B(n20250), .Z(n20248) );
  NAND U20330 ( .A(n20250), .B(n20249), .Z(n20245) );
  ANDN U20331 ( .B(B[219]), .A(n63), .Z(n19864) );
  XNOR U20332 ( .A(n19872), .B(n20251), .Z(n19865) );
  XNOR U20333 ( .A(n19871), .B(n19869), .Z(n20251) );
  AND U20334 ( .A(n20252), .B(n20253), .Z(n19869) );
  NANDN U20335 ( .A(n20254), .B(n20255), .Z(n20253) );
  NANDN U20336 ( .A(n20256), .B(n20257), .Z(n20255) );
  NANDN U20337 ( .A(n20257), .B(n20256), .Z(n20252) );
  ANDN U20338 ( .B(B[220]), .A(n64), .Z(n19871) );
  XNOR U20339 ( .A(n19879), .B(n20258), .Z(n19872) );
  XNOR U20340 ( .A(n19878), .B(n19876), .Z(n20258) );
  AND U20341 ( .A(n20259), .B(n20260), .Z(n19876) );
  NANDN U20342 ( .A(n20261), .B(n20262), .Z(n20260) );
  OR U20343 ( .A(n20263), .B(n20264), .Z(n20262) );
  NAND U20344 ( .A(n20264), .B(n20263), .Z(n20259) );
  ANDN U20345 ( .B(B[221]), .A(n65), .Z(n19878) );
  XNOR U20346 ( .A(n19886), .B(n20265), .Z(n19879) );
  XNOR U20347 ( .A(n19885), .B(n19883), .Z(n20265) );
  AND U20348 ( .A(n20266), .B(n20267), .Z(n19883) );
  NANDN U20349 ( .A(n20268), .B(n20269), .Z(n20267) );
  NANDN U20350 ( .A(n20270), .B(n20271), .Z(n20269) );
  NANDN U20351 ( .A(n20271), .B(n20270), .Z(n20266) );
  ANDN U20352 ( .B(B[222]), .A(n66), .Z(n19885) );
  XNOR U20353 ( .A(n19893), .B(n20272), .Z(n19886) );
  XNOR U20354 ( .A(n19892), .B(n19890), .Z(n20272) );
  AND U20355 ( .A(n20273), .B(n20274), .Z(n19890) );
  NANDN U20356 ( .A(n20275), .B(n20276), .Z(n20274) );
  OR U20357 ( .A(n20277), .B(n20278), .Z(n20276) );
  NAND U20358 ( .A(n20278), .B(n20277), .Z(n20273) );
  ANDN U20359 ( .B(B[223]), .A(n67), .Z(n19892) );
  XNOR U20360 ( .A(n19900), .B(n20279), .Z(n19893) );
  XNOR U20361 ( .A(n19899), .B(n19897), .Z(n20279) );
  AND U20362 ( .A(n20280), .B(n20281), .Z(n19897) );
  NANDN U20363 ( .A(n20282), .B(n20283), .Z(n20281) );
  NANDN U20364 ( .A(n20284), .B(n20285), .Z(n20283) );
  NANDN U20365 ( .A(n20285), .B(n20284), .Z(n20280) );
  ANDN U20366 ( .B(B[224]), .A(n68), .Z(n19899) );
  XNOR U20367 ( .A(n19907), .B(n20286), .Z(n19900) );
  XNOR U20368 ( .A(n19906), .B(n19904), .Z(n20286) );
  AND U20369 ( .A(n20287), .B(n20288), .Z(n19904) );
  NANDN U20370 ( .A(n20289), .B(n20290), .Z(n20288) );
  OR U20371 ( .A(n20291), .B(n20292), .Z(n20290) );
  NAND U20372 ( .A(n20292), .B(n20291), .Z(n20287) );
  ANDN U20373 ( .B(B[225]), .A(n69), .Z(n19906) );
  XNOR U20374 ( .A(n19914), .B(n20293), .Z(n19907) );
  XNOR U20375 ( .A(n19913), .B(n19911), .Z(n20293) );
  AND U20376 ( .A(n20294), .B(n20295), .Z(n19911) );
  NANDN U20377 ( .A(n20296), .B(n20297), .Z(n20295) );
  NANDN U20378 ( .A(n20298), .B(n20299), .Z(n20297) );
  NANDN U20379 ( .A(n20299), .B(n20298), .Z(n20294) );
  ANDN U20380 ( .B(B[226]), .A(n70), .Z(n19913) );
  XNOR U20381 ( .A(n19921), .B(n20300), .Z(n19914) );
  XNOR U20382 ( .A(n19920), .B(n19918), .Z(n20300) );
  AND U20383 ( .A(n20301), .B(n20302), .Z(n19918) );
  NANDN U20384 ( .A(n20303), .B(n20304), .Z(n20302) );
  OR U20385 ( .A(n20305), .B(n20306), .Z(n20304) );
  NAND U20386 ( .A(n20306), .B(n20305), .Z(n20301) );
  ANDN U20387 ( .B(B[227]), .A(n71), .Z(n19920) );
  XNOR U20388 ( .A(n19928), .B(n20307), .Z(n19921) );
  XNOR U20389 ( .A(n19927), .B(n19925), .Z(n20307) );
  AND U20390 ( .A(n20308), .B(n20309), .Z(n19925) );
  NANDN U20391 ( .A(n20310), .B(n20311), .Z(n20309) );
  NANDN U20392 ( .A(n20312), .B(n20313), .Z(n20311) );
  NANDN U20393 ( .A(n20313), .B(n20312), .Z(n20308) );
  ANDN U20394 ( .B(B[228]), .A(n72), .Z(n19927) );
  XNOR U20395 ( .A(n19935), .B(n20314), .Z(n19928) );
  XNOR U20396 ( .A(n19934), .B(n19932), .Z(n20314) );
  AND U20397 ( .A(n20315), .B(n20316), .Z(n19932) );
  NANDN U20398 ( .A(n20317), .B(n20318), .Z(n20316) );
  OR U20399 ( .A(n20319), .B(n20320), .Z(n20318) );
  NAND U20400 ( .A(n20320), .B(n20319), .Z(n20315) );
  ANDN U20401 ( .B(B[229]), .A(n73), .Z(n19934) );
  XNOR U20402 ( .A(n19942), .B(n20321), .Z(n19935) );
  XNOR U20403 ( .A(n19941), .B(n19939), .Z(n20321) );
  AND U20404 ( .A(n20322), .B(n20323), .Z(n19939) );
  NANDN U20405 ( .A(n20324), .B(n20325), .Z(n20323) );
  NANDN U20406 ( .A(n20326), .B(n20327), .Z(n20325) );
  NANDN U20407 ( .A(n20327), .B(n20326), .Z(n20322) );
  ANDN U20408 ( .B(B[230]), .A(n74), .Z(n19941) );
  XNOR U20409 ( .A(n19949), .B(n20328), .Z(n19942) );
  XNOR U20410 ( .A(n19948), .B(n19946), .Z(n20328) );
  AND U20411 ( .A(n20329), .B(n20330), .Z(n19946) );
  NANDN U20412 ( .A(n20331), .B(n20332), .Z(n20330) );
  OR U20413 ( .A(n20333), .B(n20334), .Z(n20332) );
  NAND U20414 ( .A(n20334), .B(n20333), .Z(n20329) );
  ANDN U20415 ( .B(B[231]), .A(n75), .Z(n19948) );
  XNOR U20416 ( .A(n19956), .B(n20335), .Z(n19949) );
  XNOR U20417 ( .A(n19955), .B(n19953), .Z(n20335) );
  AND U20418 ( .A(n20336), .B(n20337), .Z(n19953) );
  NANDN U20419 ( .A(n20338), .B(n20339), .Z(n20337) );
  NANDN U20420 ( .A(n20340), .B(n20341), .Z(n20339) );
  NANDN U20421 ( .A(n20341), .B(n20340), .Z(n20336) );
  ANDN U20422 ( .B(B[232]), .A(n76), .Z(n19955) );
  XNOR U20423 ( .A(n19963), .B(n20342), .Z(n19956) );
  XNOR U20424 ( .A(n19962), .B(n19960), .Z(n20342) );
  AND U20425 ( .A(n20343), .B(n20344), .Z(n19960) );
  NANDN U20426 ( .A(n20345), .B(n20346), .Z(n20344) );
  OR U20427 ( .A(n20347), .B(n20348), .Z(n20346) );
  NAND U20428 ( .A(n20348), .B(n20347), .Z(n20343) );
  ANDN U20429 ( .B(B[233]), .A(n77), .Z(n19962) );
  XNOR U20430 ( .A(n19970), .B(n20349), .Z(n19963) );
  XNOR U20431 ( .A(n19969), .B(n19967), .Z(n20349) );
  AND U20432 ( .A(n20350), .B(n20351), .Z(n19967) );
  NANDN U20433 ( .A(n20352), .B(n20353), .Z(n20351) );
  NANDN U20434 ( .A(n20354), .B(n20355), .Z(n20353) );
  NANDN U20435 ( .A(n20355), .B(n20354), .Z(n20350) );
  ANDN U20436 ( .B(B[234]), .A(n78), .Z(n19969) );
  XNOR U20437 ( .A(n19977), .B(n20356), .Z(n19970) );
  XNOR U20438 ( .A(n19976), .B(n19974), .Z(n20356) );
  AND U20439 ( .A(n20357), .B(n20358), .Z(n19974) );
  NANDN U20440 ( .A(n20359), .B(n20360), .Z(n20358) );
  OR U20441 ( .A(n20361), .B(n20362), .Z(n20360) );
  NAND U20442 ( .A(n20362), .B(n20361), .Z(n20357) );
  ANDN U20443 ( .B(B[235]), .A(n79), .Z(n19976) );
  XNOR U20444 ( .A(n19984), .B(n20363), .Z(n19977) );
  XNOR U20445 ( .A(n19983), .B(n19981), .Z(n20363) );
  AND U20446 ( .A(n20364), .B(n20365), .Z(n19981) );
  NANDN U20447 ( .A(n20366), .B(n20367), .Z(n20365) );
  NANDN U20448 ( .A(n20368), .B(n20369), .Z(n20367) );
  NANDN U20449 ( .A(n20369), .B(n20368), .Z(n20364) );
  ANDN U20450 ( .B(B[236]), .A(n80), .Z(n19983) );
  XNOR U20451 ( .A(n19991), .B(n20370), .Z(n19984) );
  XNOR U20452 ( .A(n19990), .B(n19988), .Z(n20370) );
  AND U20453 ( .A(n20371), .B(n20372), .Z(n19988) );
  NANDN U20454 ( .A(n20373), .B(n20374), .Z(n20372) );
  OR U20455 ( .A(n20375), .B(n20376), .Z(n20374) );
  NAND U20456 ( .A(n20376), .B(n20375), .Z(n20371) );
  ANDN U20457 ( .B(B[237]), .A(n81), .Z(n19990) );
  XNOR U20458 ( .A(n19998), .B(n20377), .Z(n19991) );
  XNOR U20459 ( .A(n19997), .B(n19995), .Z(n20377) );
  AND U20460 ( .A(n20378), .B(n20379), .Z(n19995) );
  NANDN U20461 ( .A(n20380), .B(n20381), .Z(n20379) );
  NAND U20462 ( .A(n20382), .B(n20383), .Z(n20381) );
  ANDN U20463 ( .B(B[238]), .A(n82), .Z(n19997) );
  XOR U20464 ( .A(n20004), .B(n20384), .Z(n19998) );
  XNOR U20465 ( .A(n20002), .B(n20005), .Z(n20384) );
  NAND U20466 ( .A(A[2]), .B(B[239]), .Z(n20005) );
  NANDN U20467 ( .A(n20385), .B(n20386), .Z(n20002) );
  AND U20468 ( .A(A[0]), .B(B[240]), .Z(n20386) );
  XNOR U20469 ( .A(n20007), .B(n20387), .Z(n20004) );
  NAND U20470 ( .A(A[0]), .B(B[241]), .Z(n20387) );
  NAND U20471 ( .A(B[240]), .B(A[1]), .Z(n20007) );
  NAND U20472 ( .A(n20388), .B(n20389), .Z(n314) );
  NANDN U20473 ( .A(n20390), .B(n20391), .Z(n20389) );
  OR U20474 ( .A(n20392), .B(n20393), .Z(n20391) );
  NAND U20475 ( .A(n20393), .B(n20392), .Z(n20388) );
  XOR U20476 ( .A(n316), .B(n315), .Z(\A1[238] ) );
  XOR U20477 ( .A(n20393), .B(n20394), .Z(n315) );
  XNOR U20478 ( .A(n20392), .B(n20390), .Z(n20394) );
  AND U20479 ( .A(n20395), .B(n20396), .Z(n20390) );
  NANDN U20480 ( .A(n20397), .B(n20398), .Z(n20396) );
  NANDN U20481 ( .A(n20399), .B(n20400), .Z(n20398) );
  NANDN U20482 ( .A(n20400), .B(n20399), .Z(n20395) );
  ANDN U20483 ( .B(B[209]), .A(n54), .Z(n20392) );
  XNOR U20484 ( .A(n20187), .B(n20401), .Z(n20393) );
  XNOR U20485 ( .A(n20186), .B(n20184), .Z(n20401) );
  AND U20486 ( .A(n20402), .B(n20403), .Z(n20184) );
  NANDN U20487 ( .A(n20404), .B(n20405), .Z(n20403) );
  OR U20488 ( .A(n20406), .B(n20407), .Z(n20405) );
  NAND U20489 ( .A(n20407), .B(n20406), .Z(n20402) );
  ANDN U20490 ( .B(B[210]), .A(n55), .Z(n20186) );
  XNOR U20491 ( .A(n20194), .B(n20408), .Z(n20187) );
  XNOR U20492 ( .A(n20193), .B(n20191), .Z(n20408) );
  AND U20493 ( .A(n20409), .B(n20410), .Z(n20191) );
  NANDN U20494 ( .A(n20411), .B(n20412), .Z(n20410) );
  NANDN U20495 ( .A(n20413), .B(n20414), .Z(n20412) );
  NANDN U20496 ( .A(n20414), .B(n20413), .Z(n20409) );
  ANDN U20497 ( .B(B[211]), .A(n56), .Z(n20193) );
  XNOR U20498 ( .A(n20201), .B(n20415), .Z(n20194) );
  XNOR U20499 ( .A(n20200), .B(n20198), .Z(n20415) );
  AND U20500 ( .A(n20416), .B(n20417), .Z(n20198) );
  NANDN U20501 ( .A(n20418), .B(n20419), .Z(n20417) );
  OR U20502 ( .A(n20420), .B(n20421), .Z(n20419) );
  NAND U20503 ( .A(n20421), .B(n20420), .Z(n20416) );
  ANDN U20504 ( .B(B[212]), .A(n57), .Z(n20200) );
  XNOR U20505 ( .A(n20208), .B(n20422), .Z(n20201) );
  XNOR U20506 ( .A(n20207), .B(n20205), .Z(n20422) );
  AND U20507 ( .A(n20423), .B(n20424), .Z(n20205) );
  NANDN U20508 ( .A(n20425), .B(n20426), .Z(n20424) );
  NANDN U20509 ( .A(n20427), .B(n20428), .Z(n20426) );
  NANDN U20510 ( .A(n20428), .B(n20427), .Z(n20423) );
  ANDN U20511 ( .B(B[213]), .A(n58), .Z(n20207) );
  XNOR U20512 ( .A(n20215), .B(n20429), .Z(n20208) );
  XNOR U20513 ( .A(n20214), .B(n20212), .Z(n20429) );
  AND U20514 ( .A(n20430), .B(n20431), .Z(n20212) );
  NANDN U20515 ( .A(n20432), .B(n20433), .Z(n20431) );
  OR U20516 ( .A(n20434), .B(n20435), .Z(n20433) );
  NAND U20517 ( .A(n20435), .B(n20434), .Z(n20430) );
  ANDN U20518 ( .B(B[214]), .A(n59), .Z(n20214) );
  XNOR U20519 ( .A(n20222), .B(n20436), .Z(n20215) );
  XNOR U20520 ( .A(n20221), .B(n20219), .Z(n20436) );
  AND U20521 ( .A(n20437), .B(n20438), .Z(n20219) );
  NANDN U20522 ( .A(n20439), .B(n20440), .Z(n20438) );
  NANDN U20523 ( .A(n20441), .B(n20442), .Z(n20440) );
  NANDN U20524 ( .A(n20442), .B(n20441), .Z(n20437) );
  ANDN U20525 ( .B(B[215]), .A(n60), .Z(n20221) );
  XNOR U20526 ( .A(n20229), .B(n20443), .Z(n20222) );
  XNOR U20527 ( .A(n20228), .B(n20226), .Z(n20443) );
  AND U20528 ( .A(n20444), .B(n20445), .Z(n20226) );
  NANDN U20529 ( .A(n20446), .B(n20447), .Z(n20445) );
  OR U20530 ( .A(n20448), .B(n20449), .Z(n20447) );
  NAND U20531 ( .A(n20449), .B(n20448), .Z(n20444) );
  ANDN U20532 ( .B(B[216]), .A(n61), .Z(n20228) );
  XNOR U20533 ( .A(n20236), .B(n20450), .Z(n20229) );
  XNOR U20534 ( .A(n20235), .B(n20233), .Z(n20450) );
  AND U20535 ( .A(n20451), .B(n20452), .Z(n20233) );
  NANDN U20536 ( .A(n20453), .B(n20454), .Z(n20452) );
  NANDN U20537 ( .A(n20455), .B(n20456), .Z(n20454) );
  NANDN U20538 ( .A(n20456), .B(n20455), .Z(n20451) );
  ANDN U20539 ( .B(B[217]), .A(n62), .Z(n20235) );
  XNOR U20540 ( .A(n20243), .B(n20457), .Z(n20236) );
  XNOR U20541 ( .A(n20242), .B(n20240), .Z(n20457) );
  AND U20542 ( .A(n20458), .B(n20459), .Z(n20240) );
  NANDN U20543 ( .A(n20460), .B(n20461), .Z(n20459) );
  OR U20544 ( .A(n20462), .B(n20463), .Z(n20461) );
  NAND U20545 ( .A(n20463), .B(n20462), .Z(n20458) );
  ANDN U20546 ( .B(B[218]), .A(n63), .Z(n20242) );
  XNOR U20547 ( .A(n20250), .B(n20464), .Z(n20243) );
  XNOR U20548 ( .A(n20249), .B(n20247), .Z(n20464) );
  AND U20549 ( .A(n20465), .B(n20466), .Z(n20247) );
  NANDN U20550 ( .A(n20467), .B(n20468), .Z(n20466) );
  NANDN U20551 ( .A(n20469), .B(n20470), .Z(n20468) );
  NANDN U20552 ( .A(n20470), .B(n20469), .Z(n20465) );
  ANDN U20553 ( .B(B[219]), .A(n64), .Z(n20249) );
  XNOR U20554 ( .A(n20257), .B(n20471), .Z(n20250) );
  XNOR U20555 ( .A(n20256), .B(n20254), .Z(n20471) );
  AND U20556 ( .A(n20472), .B(n20473), .Z(n20254) );
  NANDN U20557 ( .A(n20474), .B(n20475), .Z(n20473) );
  OR U20558 ( .A(n20476), .B(n20477), .Z(n20475) );
  NAND U20559 ( .A(n20477), .B(n20476), .Z(n20472) );
  ANDN U20560 ( .B(B[220]), .A(n65), .Z(n20256) );
  XNOR U20561 ( .A(n20264), .B(n20478), .Z(n20257) );
  XNOR U20562 ( .A(n20263), .B(n20261), .Z(n20478) );
  AND U20563 ( .A(n20479), .B(n20480), .Z(n20261) );
  NANDN U20564 ( .A(n20481), .B(n20482), .Z(n20480) );
  NANDN U20565 ( .A(n20483), .B(n20484), .Z(n20482) );
  NANDN U20566 ( .A(n20484), .B(n20483), .Z(n20479) );
  ANDN U20567 ( .B(B[221]), .A(n66), .Z(n20263) );
  XNOR U20568 ( .A(n20271), .B(n20485), .Z(n20264) );
  XNOR U20569 ( .A(n20270), .B(n20268), .Z(n20485) );
  AND U20570 ( .A(n20486), .B(n20487), .Z(n20268) );
  NANDN U20571 ( .A(n20488), .B(n20489), .Z(n20487) );
  OR U20572 ( .A(n20490), .B(n20491), .Z(n20489) );
  NAND U20573 ( .A(n20491), .B(n20490), .Z(n20486) );
  ANDN U20574 ( .B(B[222]), .A(n67), .Z(n20270) );
  XNOR U20575 ( .A(n20278), .B(n20492), .Z(n20271) );
  XNOR U20576 ( .A(n20277), .B(n20275), .Z(n20492) );
  AND U20577 ( .A(n20493), .B(n20494), .Z(n20275) );
  NANDN U20578 ( .A(n20495), .B(n20496), .Z(n20494) );
  NANDN U20579 ( .A(n20497), .B(n20498), .Z(n20496) );
  NANDN U20580 ( .A(n20498), .B(n20497), .Z(n20493) );
  ANDN U20581 ( .B(B[223]), .A(n68), .Z(n20277) );
  XNOR U20582 ( .A(n20285), .B(n20499), .Z(n20278) );
  XNOR U20583 ( .A(n20284), .B(n20282), .Z(n20499) );
  AND U20584 ( .A(n20500), .B(n20501), .Z(n20282) );
  NANDN U20585 ( .A(n20502), .B(n20503), .Z(n20501) );
  OR U20586 ( .A(n20504), .B(n20505), .Z(n20503) );
  NAND U20587 ( .A(n20505), .B(n20504), .Z(n20500) );
  ANDN U20588 ( .B(B[224]), .A(n69), .Z(n20284) );
  XNOR U20589 ( .A(n20292), .B(n20506), .Z(n20285) );
  XNOR U20590 ( .A(n20291), .B(n20289), .Z(n20506) );
  AND U20591 ( .A(n20507), .B(n20508), .Z(n20289) );
  NANDN U20592 ( .A(n20509), .B(n20510), .Z(n20508) );
  NANDN U20593 ( .A(n20511), .B(n20512), .Z(n20510) );
  NANDN U20594 ( .A(n20512), .B(n20511), .Z(n20507) );
  ANDN U20595 ( .B(B[225]), .A(n70), .Z(n20291) );
  XNOR U20596 ( .A(n20299), .B(n20513), .Z(n20292) );
  XNOR U20597 ( .A(n20298), .B(n20296), .Z(n20513) );
  AND U20598 ( .A(n20514), .B(n20515), .Z(n20296) );
  NANDN U20599 ( .A(n20516), .B(n20517), .Z(n20515) );
  OR U20600 ( .A(n20518), .B(n20519), .Z(n20517) );
  NAND U20601 ( .A(n20519), .B(n20518), .Z(n20514) );
  ANDN U20602 ( .B(B[226]), .A(n71), .Z(n20298) );
  XNOR U20603 ( .A(n20306), .B(n20520), .Z(n20299) );
  XNOR U20604 ( .A(n20305), .B(n20303), .Z(n20520) );
  AND U20605 ( .A(n20521), .B(n20522), .Z(n20303) );
  NANDN U20606 ( .A(n20523), .B(n20524), .Z(n20522) );
  NANDN U20607 ( .A(n20525), .B(n20526), .Z(n20524) );
  NANDN U20608 ( .A(n20526), .B(n20525), .Z(n20521) );
  ANDN U20609 ( .B(B[227]), .A(n72), .Z(n20305) );
  XNOR U20610 ( .A(n20313), .B(n20527), .Z(n20306) );
  XNOR U20611 ( .A(n20312), .B(n20310), .Z(n20527) );
  AND U20612 ( .A(n20528), .B(n20529), .Z(n20310) );
  NANDN U20613 ( .A(n20530), .B(n20531), .Z(n20529) );
  OR U20614 ( .A(n20532), .B(n20533), .Z(n20531) );
  NAND U20615 ( .A(n20533), .B(n20532), .Z(n20528) );
  ANDN U20616 ( .B(B[228]), .A(n73), .Z(n20312) );
  XNOR U20617 ( .A(n20320), .B(n20534), .Z(n20313) );
  XNOR U20618 ( .A(n20319), .B(n20317), .Z(n20534) );
  AND U20619 ( .A(n20535), .B(n20536), .Z(n20317) );
  NANDN U20620 ( .A(n20537), .B(n20538), .Z(n20536) );
  NANDN U20621 ( .A(n20539), .B(n20540), .Z(n20538) );
  NANDN U20622 ( .A(n20540), .B(n20539), .Z(n20535) );
  ANDN U20623 ( .B(B[229]), .A(n74), .Z(n20319) );
  XNOR U20624 ( .A(n20327), .B(n20541), .Z(n20320) );
  XNOR U20625 ( .A(n20326), .B(n20324), .Z(n20541) );
  AND U20626 ( .A(n20542), .B(n20543), .Z(n20324) );
  NANDN U20627 ( .A(n20544), .B(n20545), .Z(n20543) );
  OR U20628 ( .A(n20546), .B(n20547), .Z(n20545) );
  NAND U20629 ( .A(n20547), .B(n20546), .Z(n20542) );
  ANDN U20630 ( .B(B[230]), .A(n75), .Z(n20326) );
  XNOR U20631 ( .A(n20334), .B(n20548), .Z(n20327) );
  XNOR U20632 ( .A(n20333), .B(n20331), .Z(n20548) );
  AND U20633 ( .A(n20549), .B(n20550), .Z(n20331) );
  NANDN U20634 ( .A(n20551), .B(n20552), .Z(n20550) );
  NANDN U20635 ( .A(n20553), .B(n20554), .Z(n20552) );
  NANDN U20636 ( .A(n20554), .B(n20553), .Z(n20549) );
  ANDN U20637 ( .B(B[231]), .A(n76), .Z(n20333) );
  XNOR U20638 ( .A(n20341), .B(n20555), .Z(n20334) );
  XNOR U20639 ( .A(n20340), .B(n20338), .Z(n20555) );
  AND U20640 ( .A(n20556), .B(n20557), .Z(n20338) );
  NANDN U20641 ( .A(n20558), .B(n20559), .Z(n20557) );
  OR U20642 ( .A(n20560), .B(n20561), .Z(n20559) );
  NAND U20643 ( .A(n20561), .B(n20560), .Z(n20556) );
  ANDN U20644 ( .B(B[232]), .A(n77), .Z(n20340) );
  XNOR U20645 ( .A(n20348), .B(n20562), .Z(n20341) );
  XNOR U20646 ( .A(n20347), .B(n20345), .Z(n20562) );
  AND U20647 ( .A(n20563), .B(n20564), .Z(n20345) );
  NANDN U20648 ( .A(n20565), .B(n20566), .Z(n20564) );
  NANDN U20649 ( .A(n20567), .B(n20568), .Z(n20566) );
  NANDN U20650 ( .A(n20568), .B(n20567), .Z(n20563) );
  ANDN U20651 ( .B(B[233]), .A(n78), .Z(n20347) );
  XNOR U20652 ( .A(n20355), .B(n20569), .Z(n20348) );
  XNOR U20653 ( .A(n20354), .B(n20352), .Z(n20569) );
  AND U20654 ( .A(n20570), .B(n20571), .Z(n20352) );
  NANDN U20655 ( .A(n20572), .B(n20573), .Z(n20571) );
  OR U20656 ( .A(n20574), .B(n20575), .Z(n20573) );
  NAND U20657 ( .A(n20575), .B(n20574), .Z(n20570) );
  ANDN U20658 ( .B(B[234]), .A(n79), .Z(n20354) );
  XNOR U20659 ( .A(n20362), .B(n20576), .Z(n20355) );
  XNOR U20660 ( .A(n20361), .B(n20359), .Z(n20576) );
  AND U20661 ( .A(n20577), .B(n20578), .Z(n20359) );
  NANDN U20662 ( .A(n20579), .B(n20580), .Z(n20578) );
  NANDN U20663 ( .A(n20581), .B(n20582), .Z(n20580) );
  NANDN U20664 ( .A(n20582), .B(n20581), .Z(n20577) );
  ANDN U20665 ( .B(B[235]), .A(n80), .Z(n20361) );
  XNOR U20666 ( .A(n20369), .B(n20583), .Z(n20362) );
  XNOR U20667 ( .A(n20368), .B(n20366), .Z(n20583) );
  AND U20668 ( .A(n20584), .B(n20585), .Z(n20366) );
  NANDN U20669 ( .A(n20586), .B(n20587), .Z(n20585) );
  OR U20670 ( .A(n20588), .B(n20589), .Z(n20587) );
  NAND U20671 ( .A(n20589), .B(n20588), .Z(n20584) );
  ANDN U20672 ( .B(B[236]), .A(n81), .Z(n20368) );
  XNOR U20673 ( .A(n20376), .B(n20590), .Z(n20369) );
  XNOR U20674 ( .A(n20375), .B(n20373), .Z(n20590) );
  AND U20675 ( .A(n20591), .B(n20592), .Z(n20373) );
  NANDN U20676 ( .A(n20593), .B(n20594), .Z(n20592) );
  NAND U20677 ( .A(n20595), .B(n20596), .Z(n20594) );
  ANDN U20678 ( .B(B[237]), .A(n82), .Z(n20375) );
  XOR U20679 ( .A(n20382), .B(n20597), .Z(n20376) );
  XNOR U20680 ( .A(n20380), .B(n20383), .Z(n20597) );
  NAND U20681 ( .A(A[2]), .B(B[238]), .Z(n20383) );
  NANDN U20682 ( .A(n20598), .B(n20599), .Z(n20380) );
  AND U20683 ( .A(A[0]), .B(B[239]), .Z(n20599) );
  XNOR U20684 ( .A(n20385), .B(n20600), .Z(n20382) );
  NAND U20685 ( .A(A[0]), .B(B[240]), .Z(n20600) );
  NAND U20686 ( .A(B[239]), .B(A[1]), .Z(n20385) );
  NAND U20687 ( .A(n20601), .B(n20602), .Z(n316) );
  NANDN U20688 ( .A(n20603), .B(n20604), .Z(n20602) );
  OR U20689 ( .A(n20605), .B(n20606), .Z(n20604) );
  NAND U20690 ( .A(n20606), .B(n20605), .Z(n20601) );
  XOR U20691 ( .A(n318), .B(n317), .Z(\A1[237] ) );
  XOR U20692 ( .A(n20606), .B(n20607), .Z(n317) );
  XNOR U20693 ( .A(n20605), .B(n20603), .Z(n20607) );
  AND U20694 ( .A(n20608), .B(n20609), .Z(n20603) );
  NANDN U20695 ( .A(n20610), .B(n20611), .Z(n20609) );
  NANDN U20696 ( .A(n20612), .B(n20613), .Z(n20611) );
  NANDN U20697 ( .A(n20613), .B(n20612), .Z(n20608) );
  ANDN U20698 ( .B(B[208]), .A(n54), .Z(n20605) );
  XNOR U20699 ( .A(n20400), .B(n20614), .Z(n20606) );
  XNOR U20700 ( .A(n20399), .B(n20397), .Z(n20614) );
  AND U20701 ( .A(n20615), .B(n20616), .Z(n20397) );
  NANDN U20702 ( .A(n20617), .B(n20618), .Z(n20616) );
  OR U20703 ( .A(n20619), .B(n20620), .Z(n20618) );
  NAND U20704 ( .A(n20620), .B(n20619), .Z(n20615) );
  ANDN U20705 ( .B(B[209]), .A(n55), .Z(n20399) );
  XNOR U20706 ( .A(n20407), .B(n20621), .Z(n20400) );
  XNOR U20707 ( .A(n20406), .B(n20404), .Z(n20621) );
  AND U20708 ( .A(n20622), .B(n20623), .Z(n20404) );
  NANDN U20709 ( .A(n20624), .B(n20625), .Z(n20623) );
  NANDN U20710 ( .A(n20626), .B(n20627), .Z(n20625) );
  NANDN U20711 ( .A(n20627), .B(n20626), .Z(n20622) );
  ANDN U20712 ( .B(B[210]), .A(n56), .Z(n20406) );
  XNOR U20713 ( .A(n20414), .B(n20628), .Z(n20407) );
  XNOR U20714 ( .A(n20413), .B(n20411), .Z(n20628) );
  AND U20715 ( .A(n20629), .B(n20630), .Z(n20411) );
  NANDN U20716 ( .A(n20631), .B(n20632), .Z(n20630) );
  OR U20717 ( .A(n20633), .B(n20634), .Z(n20632) );
  NAND U20718 ( .A(n20634), .B(n20633), .Z(n20629) );
  ANDN U20719 ( .B(B[211]), .A(n57), .Z(n20413) );
  XNOR U20720 ( .A(n20421), .B(n20635), .Z(n20414) );
  XNOR U20721 ( .A(n20420), .B(n20418), .Z(n20635) );
  AND U20722 ( .A(n20636), .B(n20637), .Z(n20418) );
  NANDN U20723 ( .A(n20638), .B(n20639), .Z(n20637) );
  NANDN U20724 ( .A(n20640), .B(n20641), .Z(n20639) );
  NANDN U20725 ( .A(n20641), .B(n20640), .Z(n20636) );
  ANDN U20726 ( .B(B[212]), .A(n58), .Z(n20420) );
  XNOR U20727 ( .A(n20428), .B(n20642), .Z(n20421) );
  XNOR U20728 ( .A(n20427), .B(n20425), .Z(n20642) );
  AND U20729 ( .A(n20643), .B(n20644), .Z(n20425) );
  NANDN U20730 ( .A(n20645), .B(n20646), .Z(n20644) );
  OR U20731 ( .A(n20647), .B(n20648), .Z(n20646) );
  NAND U20732 ( .A(n20648), .B(n20647), .Z(n20643) );
  ANDN U20733 ( .B(B[213]), .A(n59), .Z(n20427) );
  XNOR U20734 ( .A(n20435), .B(n20649), .Z(n20428) );
  XNOR U20735 ( .A(n20434), .B(n20432), .Z(n20649) );
  AND U20736 ( .A(n20650), .B(n20651), .Z(n20432) );
  NANDN U20737 ( .A(n20652), .B(n20653), .Z(n20651) );
  NANDN U20738 ( .A(n20654), .B(n20655), .Z(n20653) );
  NANDN U20739 ( .A(n20655), .B(n20654), .Z(n20650) );
  ANDN U20740 ( .B(B[214]), .A(n60), .Z(n20434) );
  XNOR U20741 ( .A(n20442), .B(n20656), .Z(n20435) );
  XNOR U20742 ( .A(n20441), .B(n20439), .Z(n20656) );
  AND U20743 ( .A(n20657), .B(n20658), .Z(n20439) );
  NANDN U20744 ( .A(n20659), .B(n20660), .Z(n20658) );
  OR U20745 ( .A(n20661), .B(n20662), .Z(n20660) );
  NAND U20746 ( .A(n20662), .B(n20661), .Z(n20657) );
  ANDN U20747 ( .B(B[215]), .A(n61), .Z(n20441) );
  XNOR U20748 ( .A(n20449), .B(n20663), .Z(n20442) );
  XNOR U20749 ( .A(n20448), .B(n20446), .Z(n20663) );
  AND U20750 ( .A(n20664), .B(n20665), .Z(n20446) );
  NANDN U20751 ( .A(n20666), .B(n20667), .Z(n20665) );
  NANDN U20752 ( .A(n20668), .B(n20669), .Z(n20667) );
  NANDN U20753 ( .A(n20669), .B(n20668), .Z(n20664) );
  ANDN U20754 ( .B(B[216]), .A(n62), .Z(n20448) );
  XNOR U20755 ( .A(n20456), .B(n20670), .Z(n20449) );
  XNOR U20756 ( .A(n20455), .B(n20453), .Z(n20670) );
  AND U20757 ( .A(n20671), .B(n20672), .Z(n20453) );
  NANDN U20758 ( .A(n20673), .B(n20674), .Z(n20672) );
  OR U20759 ( .A(n20675), .B(n20676), .Z(n20674) );
  NAND U20760 ( .A(n20676), .B(n20675), .Z(n20671) );
  ANDN U20761 ( .B(B[217]), .A(n63), .Z(n20455) );
  XNOR U20762 ( .A(n20463), .B(n20677), .Z(n20456) );
  XNOR U20763 ( .A(n20462), .B(n20460), .Z(n20677) );
  AND U20764 ( .A(n20678), .B(n20679), .Z(n20460) );
  NANDN U20765 ( .A(n20680), .B(n20681), .Z(n20679) );
  NANDN U20766 ( .A(n20682), .B(n20683), .Z(n20681) );
  NANDN U20767 ( .A(n20683), .B(n20682), .Z(n20678) );
  ANDN U20768 ( .B(B[218]), .A(n64), .Z(n20462) );
  XNOR U20769 ( .A(n20470), .B(n20684), .Z(n20463) );
  XNOR U20770 ( .A(n20469), .B(n20467), .Z(n20684) );
  AND U20771 ( .A(n20685), .B(n20686), .Z(n20467) );
  NANDN U20772 ( .A(n20687), .B(n20688), .Z(n20686) );
  OR U20773 ( .A(n20689), .B(n20690), .Z(n20688) );
  NAND U20774 ( .A(n20690), .B(n20689), .Z(n20685) );
  ANDN U20775 ( .B(B[219]), .A(n65), .Z(n20469) );
  XNOR U20776 ( .A(n20477), .B(n20691), .Z(n20470) );
  XNOR U20777 ( .A(n20476), .B(n20474), .Z(n20691) );
  AND U20778 ( .A(n20692), .B(n20693), .Z(n20474) );
  NANDN U20779 ( .A(n20694), .B(n20695), .Z(n20693) );
  NANDN U20780 ( .A(n20696), .B(n20697), .Z(n20695) );
  NANDN U20781 ( .A(n20697), .B(n20696), .Z(n20692) );
  ANDN U20782 ( .B(B[220]), .A(n66), .Z(n20476) );
  XNOR U20783 ( .A(n20484), .B(n20698), .Z(n20477) );
  XNOR U20784 ( .A(n20483), .B(n20481), .Z(n20698) );
  AND U20785 ( .A(n20699), .B(n20700), .Z(n20481) );
  NANDN U20786 ( .A(n20701), .B(n20702), .Z(n20700) );
  OR U20787 ( .A(n20703), .B(n20704), .Z(n20702) );
  NAND U20788 ( .A(n20704), .B(n20703), .Z(n20699) );
  ANDN U20789 ( .B(B[221]), .A(n67), .Z(n20483) );
  XNOR U20790 ( .A(n20491), .B(n20705), .Z(n20484) );
  XNOR U20791 ( .A(n20490), .B(n20488), .Z(n20705) );
  AND U20792 ( .A(n20706), .B(n20707), .Z(n20488) );
  NANDN U20793 ( .A(n20708), .B(n20709), .Z(n20707) );
  NANDN U20794 ( .A(n20710), .B(n20711), .Z(n20709) );
  NANDN U20795 ( .A(n20711), .B(n20710), .Z(n20706) );
  ANDN U20796 ( .B(B[222]), .A(n68), .Z(n20490) );
  XNOR U20797 ( .A(n20498), .B(n20712), .Z(n20491) );
  XNOR U20798 ( .A(n20497), .B(n20495), .Z(n20712) );
  AND U20799 ( .A(n20713), .B(n20714), .Z(n20495) );
  NANDN U20800 ( .A(n20715), .B(n20716), .Z(n20714) );
  OR U20801 ( .A(n20717), .B(n20718), .Z(n20716) );
  NAND U20802 ( .A(n20718), .B(n20717), .Z(n20713) );
  ANDN U20803 ( .B(B[223]), .A(n69), .Z(n20497) );
  XNOR U20804 ( .A(n20505), .B(n20719), .Z(n20498) );
  XNOR U20805 ( .A(n20504), .B(n20502), .Z(n20719) );
  AND U20806 ( .A(n20720), .B(n20721), .Z(n20502) );
  NANDN U20807 ( .A(n20722), .B(n20723), .Z(n20721) );
  NANDN U20808 ( .A(n20724), .B(n20725), .Z(n20723) );
  NANDN U20809 ( .A(n20725), .B(n20724), .Z(n20720) );
  ANDN U20810 ( .B(B[224]), .A(n70), .Z(n20504) );
  XNOR U20811 ( .A(n20512), .B(n20726), .Z(n20505) );
  XNOR U20812 ( .A(n20511), .B(n20509), .Z(n20726) );
  AND U20813 ( .A(n20727), .B(n20728), .Z(n20509) );
  NANDN U20814 ( .A(n20729), .B(n20730), .Z(n20728) );
  OR U20815 ( .A(n20731), .B(n20732), .Z(n20730) );
  NAND U20816 ( .A(n20732), .B(n20731), .Z(n20727) );
  ANDN U20817 ( .B(B[225]), .A(n71), .Z(n20511) );
  XNOR U20818 ( .A(n20519), .B(n20733), .Z(n20512) );
  XNOR U20819 ( .A(n20518), .B(n20516), .Z(n20733) );
  AND U20820 ( .A(n20734), .B(n20735), .Z(n20516) );
  NANDN U20821 ( .A(n20736), .B(n20737), .Z(n20735) );
  NANDN U20822 ( .A(n20738), .B(n20739), .Z(n20737) );
  NANDN U20823 ( .A(n20739), .B(n20738), .Z(n20734) );
  ANDN U20824 ( .B(B[226]), .A(n72), .Z(n20518) );
  XNOR U20825 ( .A(n20526), .B(n20740), .Z(n20519) );
  XNOR U20826 ( .A(n20525), .B(n20523), .Z(n20740) );
  AND U20827 ( .A(n20741), .B(n20742), .Z(n20523) );
  NANDN U20828 ( .A(n20743), .B(n20744), .Z(n20742) );
  OR U20829 ( .A(n20745), .B(n20746), .Z(n20744) );
  NAND U20830 ( .A(n20746), .B(n20745), .Z(n20741) );
  ANDN U20831 ( .B(B[227]), .A(n73), .Z(n20525) );
  XNOR U20832 ( .A(n20533), .B(n20747), .Z(n20526) );
  XNOR U20833 ( .A(n20532), .B(n20530), .Z(n20747) );
  AND U20834 ( .A(n20748), .B(n20749), .Z(n20530) );
  NANDN U20835 ( .A(n20750), .B(n20751), .Z(n20749) );
  NANDN U20836 ( .A(n20752), .B(n20753), .Z(n20751) );
  NANDN U20837 ( .A(n20753), .B(n20752), .Z(n20748) );
  ANDN U20838 ( .B(B[228]), .A(n74), .Z(n20532) );
  XNOR U20839 ( .A(n20540), .B(n20754), .Z(n20533) );
  XNOR U20840 ( .A(n20539), .B(n20537), .Z(n20754) );
  AND U20841 ( .A(n20755), .B(n20756), .Z(n20537) );
  NANDN U20842 ( .A(n20757), .B(n20758), .Z(n20756) );
  OR U20843 ( .A(n20759), .B(n20760), .Z(n20758) );
  NAND U20844 ( .A(n20760), .B(n20759), .Z(n20755) );
  ANDN U20845 ( .B(B[229]), .A(n75), .Z(n20539) );
  XNOR U20846 ( .A(n20547), .B(n20761), .Z(n20540) );
  XNOR U20847 ( .A(n20546), .B(n20544), .Z(n20761) );
  AND U20848 ( .A(n20762), .B(n20763), .Z(n20544) );
  NANDN U20849 ( .A(n20764), .B(n20765), .Z(n20763) );
  NANDN U20850 ( .A(n20766), .B(n20767), .Z(n20765) );
  NANDN U20851 ( .A(n20767), .B(n20766), .Z(n20762) );
  ANDN U20852 ( .B(B[230]), .A(n76), .Z(n20546) );
  XNOR U20853 ( .A(n20554), .B(n20768), .Z(n20547) );
  XNOR U20854 ( .A(n20553), .B(n20551), .Z(n20768) );
  AND U20855 ( .A(n20769), .B(n20770), .Z(n20551) );
  NANDN U20856 ( .A(n20771), .B(n20772), .Z(n20770) );
  OR U20857 ( .A(n20773), .B(n20774), .Z(n20772) );
  NAND U20858 ( .A(n20774), .B(n20773), .Z(n20769) );
  ANDN U20859 ( .B(B[231]), .A(n77), .Z(n20553) );
  XNOR U20860 ( .A(n20561), .B(n20775), .Z(n20554) );
  XNOR U20861 ( .A(n20560), .B(n20558), .Z(n20775) );
  AND U20862 ( .A(n20776), .B(n20777), .Z(n20558) );
  NANDN U20863 ( .A(n20778), .B(n20779), .Z(n20777) );
  NANDN U20864 ( .A(n20780), .B(n20781), .Z(n20779) );
  NANDN U20865 ( .A(n20781), .B(n20780), .Z(n20776) );
  ANDN U20866 ( .B(B[232]), .A(n78), .Z(n20560) );
  XNOR U20867 ( .A(n20568), .B(n20782), .Z(n20561) );
  XNOR U20868 ( .A(n20567), .B(n20565), .Z(n20782) );
  AND U20869 ( .A(n20783), .B(n20784), .Z(n20565) );
  NANDN U20870 ( .A(n20785), .B(n20786), .Z(n20784) );
  OR U20871 ( .A(n20787), .B(n20788), .Z(n20786) );
  NAND U20872 ( .A(n20788), .B(n20787), .Z(n20783) );
  ANDN U20873 ( .B(B[233]), .A(n79), .Z(n20567) );
  XNOR U20874 ( .A(n20575), .B(n20789), .Z(n20568) );
  XNOR U20875 ( .A(n20574), .B(n20572), .Z(n20789) );
  AND U20876 ( .A(n20790), .B(n20791), .Z(n20572) );
  NANDN U20877 ( .A(n20792), .B(n20793), .Z(n20791) );
  NANDN U20878 ( .A(n20794), .B(n20795), .Z(n20793) );
  NANDN U20879 ( .A(n20795), .B(n20794), .Z(n20790) );
  ANDN U20880 ( .B(B[234]), .A(n80), .Z(n20574) );
  XNOR U20881 ( .A(n20582), .B(n20796), .Z(n20575) );
  XNOR U20882 ( .A(n20581), .B(n20579), .Z(n20796) );
  AND U20883 ( .A(n20797), .B(n20798), .Z(n20579) );
  NANDN U20884 ( .A(n20799), .B(n20800), .Z(n20798) );
  OR U20885 ( .A(n20801), .B(n20802), .Z(n20800) );
  NAND U20886 ( .A(n20802), .B(n20801), .Z(n20797) );
  ANDN U20887 ( .B(B[235]), .A(n81), .Z(n20581) );
  XNOR U20888 ( .A(n20589), .B(n20803), .Z(n20582) );
  XNOR U20889 ( .A(n20588), .B(n20586), .Z(n20803) );
  AND U20890 ( .A(n20804), .B(n20805), .Z(n20586) );
  NANDN U20891 ( .A(n20806), .B(n20807), .Z(n20805) );
  NAND U20892 ( .A(n20808), .B(n20809), .Z(n20807) );
  ANDN U20893 ( .B(B[236]), .A(n82), .Z(n20588) );
  XOR U20894 ( .A(n20595), .B(n20810), .Z(n20589) );
  XNOR U20895 ( .A(n20593), .B(n20596), .Z(n20810) );
  NAND U20896 ( .A(A[2]), .B(B[237]), .Z(n20596) );
  NANDN U20897 ( .A(n20811), .B(n20812), .Z(n20593) );
  AND U20898 ( .A(A[0]), .B(B[238]), .Z(n20812) );
  XNOR U20899 ( .A(n20598), .B(n20813), .Z(n20595) );
  NAND U20900 ( .A(A[0]), .B(B[239]), .Z(n20813) );
  NAND U20901 ( .A(B[238]), .B(A[1]), .Z(n20598) );
  NAND U20902 ( .A(n20814), .B(n20815), .Z(n318) );
  NANDN U20903 ( .A(n20816), .B(n20817), .Z(n20815) );
  OR U20904 ( .A(n20818), .B(n20819), .Z(n20817) );
  NAND U20905 ( .A(n20819), .B(n20818), .Z(n20814) );
  XOR U20906 ( .A(n320), .B(n319), .Z(\A1[236] ) );
  XOR U20907 ( .A(n20819), .B(n20820), .Z(n319) );
  XNOR U20908 ( .A(n20818), .B(n20816), .Z(n20820) );
  AND U20909 ( .A(n20821), .B(n20822), .Z(n20816) );
  NANDN U20910 ( .A(n20823), .B(n20824), .Z(n20822) );
  NANDN U20911 ( .A(n20825), .B(n20826), .Z(n20824) );
  NANDN U20912 ( .A(n20826), .B(n20825), .Z(n20821) );
  ANDN U20913 ( .B(B[207]), .A(n54), .Z(n20818) );
  XNOR U20914 ( .A(n20613), .B(n20827), .Z(n20819) );
  XNOR U20915 ( .A(n20612), .B(n20610), .Z(n20827) );
  AND U20916 ( .A(n20828), .B(n20829), .Z(n20610) );
  NANDN U20917 ( .A(n20830), .B(n20831), .Z(n20829) );
  OR U20918 ( .A(n20832), .B(n20833), .Z(n20831) );
  NAND U20919 ( .A(n20833), .B(n20832), .Z(n20828) );
  ANDN U20920 ( .B(B[208]), .A(n55), .Z(n20612) );
  XNOR U20921 ( .A(n20620), .B(n20834), .Z(n20613) );
  XNOR U20922 ( .A(n20619), .B(n20617), .Z(n20834) );
  AND U20923 ( .A(n20835), .B(n20836), .Z(n20617) );
  NANDN U20924 ( .A(n20837), .B(n20838), .Z(n20836) );
  NANDN U20925 ( .A(n20839), .B(n20840), .Z(n20838) );
  NANDN U20926 ( .A(n20840), .B(n20839), .Z(n20835) );
  ANDN U20927 ( .B(B[209]), .A(n56), .Z(n20619) );
  XNOR U20928 ( .A(n20627), .B(n20841), .Z(n20620) );
  XNOR U20929 ( .A(n20626), .B(n20624), .Z(n20841) );
  AND U20930 ( .A(n20842), .B(n20843), .Z(n20624) );
  NANDN U20931 ( .A(n20844), .B(n20845), .Z(n20843) );
  OR U20932 ( .A(n20846), .B(n20847), .Z(n20845) );
  NAND U20933 ( .A(n20847), .B(n20846), .Z(n20842) );
  ANDN U20934 ( .B(B[210]), .A(n57), .Z(n20626) );
  XNOR U20935 ( .A(n20634), .B(n20848), .Z(n20627) );
  XNOR U20936 ( .A(n20633), .B(n20631), .Z(n20848) );
  AND U20937 ( .A(n20849), .B(n20850), .Z(n20631) );
  NANDN U20938 ( .A(n20851), .B(n20852), .Z(n20850) );
  NANDN U20939 ( .A(n20853), .B(n20854), .Z(n20852) );
  NANDN U20940 ( .A(n20854), .B(n20853), .Z(n20849) );
  ANDN U20941 ( .B(B[211]), .A(n58), .Z(n20633) );
  XNOR U20942 ( .A(n20641), .B(n20855), .Z(n20634) );
  XNOR U20943 ( .A(n20640), .B(n20638), .Z(n20855) );
  AND U20944 ( .A(n20856), .B(n20857), .Z(n20638) );
  NANDN U20945 ( .A(n20858), .B(n20859), .Z(n20857) );
  OR U20946 ( .A(n20860), .B(n20861), .Z(n20859) );
  NAND U20947 ( .A(n20861), .B(n20860), .Z(n20856) );
  ANDN U20948 ( .B(B[212]), .A(n59), .Z(n20640) );
  XNOR U20949 ( .A(n20648), .B(n20862), .Z(n20641) );
  XNOR U20950 ( .A(n20647), .B(n20645), .Z(n20862) );
  AND U20951 ( .A(n20863), .B(n20864), .Z(n20645) );
  NANDN U20952 ( .A(n20865), .B(n20866), .Z(n20864) );
  NANDN U20953 ( .A(n20867), .B(n20868), .Z(n20866) );
  NANDN U20954 ( .A(n20868), .B(n20867), .Z(n20863) );
  ANDN U20955 ( .B(B[213]), .A(n60), .Z(n20647) );
  XNOR U20956 ( .A(n20655), .B(n20869), .Z(n20648) );
  XNOR U20957 ( .A(n20654), .B(n20652), .Z(n20869) );
  AND U20958 ( .A(n20870), .B(n20871), .Z(n20652) );
  NANDN U20959 ( .A(n20872), .B(n20873), .Z(n20871) );
  OR U20960 ( .A(n20874), .B(n20875), .Z(n20873) );
  NAND U20961 ( .A(n20875), .B(n20874), .Z(n20870) );
  ANDN U20962 ( .B(B[214]), .A(n61), .Z(n20654) );
  XNOR U20963 ( .A(n20662), .B(n20876), .Z(n20655) );
  XNOR U20964 ( .A(n20661), .B(n20659), .Z(n20876) );
  AND U20965 ( .A(n20877), .B(n20878), .Z(n20659) );
  NANDN U20966 ( .A(n20879), .B(n20880), .Z(n20878) );
  NANDN U20967 ( .A(n20881), .B(n20882), .Z(n20880) );
  NANDN U20968 ( .A(n20882), .B(n20881), .Z(n20877) );
  ANDN U20969 ( .B(B[215]), .A(n62), .Z(n20661) );
  XNOR U20970 ( .A(n20669), .B(n20883), .Z(n20662) );
  XNOR U20971 ( .A(n20668), .B(n20666), .Z(n20883) );
  AND U20972 ( .A(n20884), .B(n20885), .Z(n20666) );
  NANDN U20973 ( .A(n20886), .B(n20887), .Z(n20885) );
  OR U20974 ( .A(n20888), .B(n20889), .Z(n20887) );
  NAND U20975 ( .A(n20889), .B(n20888), .Z(n20884) );
  ANDN U20976 ( .B(B[216]), .A(n63), .Z(n20668) );
  XNOR U20977 ( .A(n20676), .B(n20890), .Z(n20669) );
  XNOR U20978 ( .A(n20675), .B(n20673), .Z(n20890) );
  AND U20979 ( .A(n20891), .B(n20892), .Z(n20673) );
  NANDN U20980 ( .A(n20893), .B(n20894), .Z(n20892) );
  NANDN U20981 ( .A(n20895), .B(n20896), .Z(n20894) );
  NANDN U20982 ( .A(n20896), .B(n20895), .Z(n20891) );
  ANDN U20983 ( .B(B[217]), .A(n64), .Z(n20675) );
  XNOR U20984 ( .A(n20683), .B(n20897), .Z(n20676) );
  XNOR U20985 ( .A(n20682), .B(n20680), .Z(n20897) );
  AND U20986 ( .A(n20898), .B(n20899), .Z(n20680) );
  NANDN U20987 ( .A(n20900), .B(n20901), .Z(n20899) );
  OR U20988 ( .A(n20902), .B(n20903), .Z(n20901) );
  NAND U20989 ( .A(n20903), .B(n20902), .Z(n20898) );
  ANDN U20990 ( .B(B[218]), .A(n65), .Z(n20682) );
  XNOR U20991 ( .A(n20690), .B(n20904), .Z(n20683) );
  XNOR U20992 ( .A(n20689), .B(n20687), .Z(n20904) );
  AND U20993 ( .A(n20905), .B(n20906), .Z(n20687) );
  NANDN U20994 ( .A(n20907), .B(n20908), .Z(n20906) );
  NANDN U20995 ( .A(n20909), .B(n20910), .Z(n20908) );
  NANDN U20996 ( .A(n20910), .B(n20909), .Z(n20905) );
  ANDN U20997 ( .B(B[219]), .A(n66), .Z(n20689) );
  XNOR U20998 ( .A(n20697), .B(n20911), .Z(n20690) );
  XNOR U20999 ( .A(n20696), .B(n20694), .Z(n20911) );
  AND U21000 ( .A(n20912), .B(n20913), .Z(n20694) );
  NANDN U21001 ( .A(n20914), .B(n20915), .Z(n20913) );
  OR U21002 ( .A(n20916), .B(n20917), .Z(n20915) );
  NAND U21003 ( .A(n20917), .B(n20916), .Z(n20912) );
  ANDN U21004 ( .B(B[220]), .A(n67), .Z(n20696) );
  XNOR U21005 ( .A(n20704), .B(n20918), .Z(n20697) );
  XNOR U21006 ( .A(n20703), .B(n20701), .Z(n20918) );
  AND U21007 ( .A(n20919), .B(n20920), .Z(n20701) );
  NANDN U21008 ( .A(n20921), .B(n20922), .Z(n20920) );
  NANDN U21009 ( .A(n20923), .B(n20924), .Z(n20922) );
  NANDN U21010 ( .A(n20924), .B(n20923), .Z(n20919) );
  ANDN U21011 ( .B(B[221]), .A(n68), .Z(n20703) );
  XNOR U21012 ( .A(n20711), .B(n20925), .Z(n20704) );
  XNOR U21013 ( .A(n20710), .B(n20708), .Z(n20925) );
  AND U21014 ( .A(n20926), .B(n20927), .Z(n20708) );
  NANDN U21015 ( .A(n20928), .B(n20929), .Z(n20927) );
  OR U21016 ( .A(n20930), .B(n20931), .Z(n20929) );
  NAND U21017 ( .A(n20931), .B(n20930), .Z(n20926) );
  ANDN U21018 ( .B(B[222]), .A(n69), .Z(n20710) );
  XNOR U21019 ( .A(n20718), .B(n20932), .Z(n20711) );
  XNOR U21020 ( .A(n20717), .B(n20715), .Z(n20932) );
  AND U21021 ( .A(n20933), .B(n20934), .Z(n20715) );
  NANDN U21022 ( .A(n20935), .B(n20936), .Z(n20934) );
  NANDN U21023 ( .A(n20937), .B(n20938), .Z(n20936) );
  NANDN U21024 ( .A(n20938), .B(n20937), .Z(n20933) );
  ANDN U21025 ( .B(B[223]), .A(n70), .Z(n20717) );
  XNOR U21026 ( .A(n20725), .B(n20939), .Z(n20718) );
  XNOR U21027 ( .A(n20724), .B(n20722), .Z(n20939) );
  AND U21028 ( .A(n20940), .B(n20941), .Z(n20722) );
  NANDN U21029 ( .A(n20942), .B(n20943), .Z(n20941) );
  OR U21030 ( .A(n20944), .B(n20945), .Z(n20943) );
  NAND U21031 ( .A(n20945), .B(n20944), .Z(n20940) );
  ANDN U21032 ( .B(B[224]), .A(n71), .Z(n20724) );
  XNOR U21033 ( .A(n20732), .B(n20946), .Z(n20725) );
  XNOR U21034 ( .A(n20731), .B(n20729), .Z(n20946) );
  AND U21035 ( .A(n20947), .B(n20948), .Z(n20729) );
  NANDN U21036 ( .A(n20949), .B(n20950), .Z(n20948) );
  NANDN U21037 ( .A(n20951), .B(n20952), .Z(n20950) );
  NANDN U21038 ( .A(n20952), .B(n20951), .Z(n20947) );
  ANDN U21039 ( .B(B[225]), .A(n72), .Z(n20731) );
  XNOR U21040 ( .A(n20739), .B(n20953), .Z(n20732) );
  XNOR U21041 ( .A(n20738), .B(n20736), .Z(n20953) );
  AND U21042 ( .A(n20954), .B(n20955), .Z(n20736) );
  NANDN U21043 ( .A(n20956), .B(n20957), .Z(n20955) );
  OR U21044 ( .A(n20958), .B(n20959), .Z(n20957) );
  NAND U21045 ( .A(n20959), .B(n20958), .Z(n20954) );
  ANDN U21046 ( .B(B[226]), .A(n73), .Z(n20738) );
  XNOR U21047 ( .A(n20746), .B(n20960), .Z(n20739) );
  XNOR U21048 ( .A(n20745), .B(n20743), .Z(n20960) );
  AND U21049 ( .A(n20961), .B(n20962), .Z(n20743) );
  NANDN U21050 ( .A(n20963), .B(n20964), .Z(n20962) );
  NANDN U21051 ( .A(n20965), .B(n20966), .Z(n20964) );
  NANDN U21052 ( .A(n20966), .B(n20965), .Z(n20961) );
  ANDN U21053 ( .B(B[227]), .A(n74), .Z(n20745) );
  XNOR U21054 ( .A(n20753), .B(n20967), .Z(n20746) );
  XNOR U21055 ( .A(n20752), .B(n20750), .Z(n20967) );
  AND U21056 ( .A(n20968), .B(n20969), .Z(n20750) );
  NANDN U21057 ( .A(n20970), .B(n20971), .Z(n20969) );
  OR U21058 ( .A(n20972), .B(n20973), .Z(n20971) );
  NAND U21059 ( .A(n20973), .B(n20972), .Z(n20968) );
  ANDN U21060 ( .B(B[228]), .A(n75), .Z(n20752) );
  XNOR U21061 ( .A(n20760), .B(n20974), .Z(n20753) );
  XNOR U21062 ( .A(n20759), .B(n20757), .Z(n20974) );
  AND U21063 ( .A(n20975), .B(n20976), .Z(n20757) );
  NANDN U21064 ( .A(n20977), .B(n20978), .Z(n20976) );
  NANDN U21065 ( .A(n20979), .B(n20980), .Z(n20978) );
  NANDN U21066 ( .A(n20980), .B(n20979), .Z(n20975) );
  ANDN U21067 ( .B(B[229]), .A(n76), .Z(n20759) );
  XNOR U21068 ( .A(n20767), .B(n20981), .Z(n20760) );
  XNOR U21069 ( .A(n20766), .B(n20764), .Z(n20981) );
  AND U21070 ( .A(n20982), .B(n20983), .Z(n20764) );
  NANDN U21071 ( .A(n20984), .B(n20985), .Z(n20983) );
  OR U21072 ( .A(n20986), .B(n20987), .Z(n20985) );
  NAND U21073 ( .A(n20987), .B(n20986), .Z(n20982) );
  ANDN U21074 ( .B(B[230]), .A(n77), .Z(n20766) );
  XNOR U21075 ( .A(n20774), .B(n20988), .Z(n20767) );
  XNOR U21076 ( .A(n20773), .B(n20771), .Z(n20988) );
  AND U21077 ( .A(n20989), .B(n20990), .Z(n20771) );
  NANDN U21078 ( .A(n20991), .B(n20992), .Z(n20990) );
  NANDN U21079 ( .A(n20993), .B(n20994), .Z(n20992) );
  NANDN U21080 ( .A(n20994), .B(n20993), .Z(n20989) );
  ANDN U21081 ( .B(B[231]), .A(n78), .Z(n20773) );
  XNOR U21082 ( .A(n20781), .B(n20995), .Z(n20774) );
  XNOR U21083 ( .A(n20780), .B(n20778), .Z(n20995) );
  AND U21084 ( .A(n20996), .B(n20997), .Z(n20778) );
  NANDN U21085 ( .A(n20998), .B(n20999), .Z(n20997) );
  OR U21086 ( .A(n21000), .B(n21001), .Z(n20999) );
  NAND U21087 ( .A(n21001), .B(n21000), .Z(n20996) );
  ANDN U21088 ( .B(B[232]), .A(n79), .Z(n20780) );
  XNOR U21089 ( .A(n20788), .B(n21002), .Z(n20781) );
  XNOR U21090 ( .A(n20787), .B(n20785), .Z(n21002) );
  AND U21091 ( .A(n21003), .B(n21004), .Z(n20785) );
  NANDN U21092 ( .A(n21005), .B(n21006), .Z(n21004) );
  NANDN U21093 ( .A(n21007), .B(n21008), .Z(n21006) );
  NANDN U21094 ( .A(n21008), .B(n21007), .Z(n21003) );
  ANDN U21095 ( .B(B[233]), .A(n80), .Z(n20787) );
  XNOR U21096 ( .A(n20795), .B(n21009), .Z(n20788) );
  XNOR U21097 ( .A(n20794), .B(n20792), .Z(n21009) );
  AND U21098 ( .A(n21010), .B(n21011), .Z(n20792) );
  NANDN U21099 ( .A(n21012), .B(n21013), .Z(n21011) );
  OR U21100 ( .A(n21014), .B(n21015), .Z(n21013) );
  NAND U21101 ( .A(n21015), .B(n21014), .Z(n21010) );
  ANDN U21102 ( .B(B[234]), .A(n81), .Z(n20794) );
  XNOR U21103 ( .A(n20802), .B(n21016), .Z(n20795) );
  XNOR U21104 ( .A(n20801), .B(n20799), .Z(n21016) );
  AND U21105 ( .A(n21017), .B(n21018), .Z(n20799) );
  NANDN U21106 ( .A(n21019), .B(n21020), .Z(n21018) );
  NAND U21107 ( .A(n21021), .B(n21022), .Z(n21020) );
  ANDN U21108 ( .B(B[235]), .A(n82), .Z(n20801) );
  XOR U21109 ( .A(n20808), .B(n21023), .Z(n20802) );
  XNOR U21110 ( .A(n20806), .B(n20809), .Z(n21023) );
  NAND U21111 ( .A(A[2]), .B(B[236]), .Z(n20809) );
  NANDN U21112 ( .A(n21024), .B(n21025), .Z(n20806) );
  AND U21113 ( .A(A[0]), .B(B[237]), .Z(n21025) );
  XNOR U21114 ( .A(n20811), .B(n21026), .Z(n20808) );
  NAND U21115 ( .A(A[0]), .B(B[238]), .Z(n21026) );
  NAND U21116 ( .A(B[237]), .B(A[1]), .Z(n20811) );
  NAND U21117 ( .A(n21027), .B(n21028), .Z(n320) );
  NANDN U21118 ( .A(n21029), .B(n21030), .Z(n21028) );
  OR U21119 ( .A(n21031), .B(n21032), .Z(n21030) );
  NAND U21120 ( .A(n21032), .B(n21031), .Z(n21027) );
  XOR U21121 ( .A(n322), .B(n321), .Z(\A1[235] ) );
  XOR U21122 ( .A(n21032), .B(n21033), .Z(n321) );
  XNOR U21123 ( .A(n21031), .B(n21029), .Z(n21033) );
  AND U21124 ( .A(n21034), .B(n21035), .Z(n21029) );
  NANDN U21125 ( .A(n21036), .B(n21037), .Z(n21035) );
  NANDN U21126 ( .A(n21038), .B(n21039), .Z(n21037) );
  NANDN U21127 ( .A(n21039), .B(n21038), .Z(n21034) );
  ANDN U21128 ( .B(B[206]), .A(n54), .Z(n21031) );
  XNOR U21129 ( .A(n20826), .B(n21040), .Z(n21032) );
  XNOR U21130 ( .A(n20825), .B(n20823), .Z(n21040) );
  AND U21131 ( .A(n21041), .B(n21042), .Z(n20823) );
  NANDN U21132 ( .A(n21043), .B(n21044), .Z(n21042) );
  OR U21133 ( .A(n21045), .B(n21046), .Z(n21044) );
  NAND U21134 ( .A(n21046), .B(n21045), .Z(n21041) );
  ANDN U21135 ( .B(B[207]), .A(n55), .Z(n20825) );
  XNOR U21136 ( .A(n20833), .B(n21047), .Z(n20826) );
  XNOR U21137 ( .A(n20832), .B(n20830), .Z(n21047) );
  AND U21138 ( .A(n21048), .B(n21049), .Z(n20830) );
  NANDN U21139 ( .A(n21050), .B(n21051), .Z(n21049) );
  NANDN U21140 ( .A(n21052), .B(n21053), .Z(n21051) );
  NANDN U21141 ( .A(n21053), .B(n21052), .Z(n21048) );
  ANDN U21142 ( .B(B[208]), .A(n56), .Z(n20832) );
  XNOR U21143 ( .A(n20840), .B(n21054), .Z(n20833) );
  XNOR U21144 ( .A(n20839), .B(n20837), .Z(n21054) );
  AND U21145 ( .A(n21055), .B(n21056), .Z(n20837) );
  NANDN U21146 ( .A(n21057), .B(n21058), .Z(n21056) );
  OR U21147 ( .A(n21059), .B(n21060), .Z(n21058) );
  NAND U21148 ( .A(n21060), .B(n21059), .Z(n21055) );
  ANDN U21149 ( .B(B[209]), .A(n57), .Z(n20839) );
  XNOR U21150 ( .A(n20847), .B(n21061), .Z(n20840) );
  XNOR U21151 ( .A(n20846), .B(n20844), .Z(n21061) );
  AND U21152 ( .A(n21062), .B(n21063), .Z(n20844) );
  NANDN U21153 ( .A(n21064), .B(n21065), .Z(n21063) );
  NANDN U21154 ( .A(n21066), .B(n21067), .Z(n21065) );
  NANDN U21155 ( .A(n21067), .B(n21066), .Z(n21062) );
  ANDN U21156 ( .B(B[210]), .A(n58), .Z(n20846) );
  XNOR U21157 ( .A(n20854), .B(n21068), .Z(n20847) );
  XNOR U21158 ( .A(n20853), .B(n20851), .Z(n21068) );
  AND U21159 ( .A(n21069), .B(n21070), .Z(n20851) );
  NANDN U21160 ( .A(n21071), .B(n21072), .Z(n21070) );
  OR U21161 ( .A(n21073), .B(n21074), .Z(n21072) );
  NAND U21162 ( .A(n21074), .B(n21073), .Z(n21069) );
  ANDN U21163 ( .B(B[211]), .A(n59), .Z(n20853) );
  XNOR U21164 ( .A(n20861), .B(n21075), .Z(n20854) );
  XNOR U21165 ( .A(n20860), .B(n20858), .Z(n21075) );
  AND U21166 ( .A(n21076), .B(n21077), .Z(n20858) );
  NANDN U21167 ( .A(n21078), .B(n21079), .Z(n21077) );
  NANDN U21168 ( .A(n21080), .B(n21081), .Z(n21079) );
  NANDN U21169 ( .A(n21081), .B(n21080), .Z(n21076) );
  ANDN U21170 ( .B(B[212]), .A(n60), .Z(n20860) );
  XNOR U21171 ( .A(n20868), .B(n21082), .Z(n20861) );
  XNOR U21172 ( .A(n20867), .B(n20865), .Z(n21082) );
  AND U21173 ( .A(n21083), .B(n21084), .Z(n20865) );
  NANDN U21174 ( .A(n21085), .B(n21086), .Z(n21084) );
  OR U21175 ( .A(n21087), .B(n21088), .Z(n21086) );
  NAND U21176 ( .A(n21088), .B(n21087), .Z(n21083) );
  ANDN U21177 ( .B(B[213]), .A(n61), .Z(n20867) );
  XNOR U21178 ( .A(n20875), .B(n21089), .Z(n20868) );
  XNOR U21179 ( .A(n20874), .B(n20872), .Z(n21089) );
  AND U21180 ( .A(n21090), .B(n21091), .Z(n20872) );
  NANDN U21181 ( .A(n21092), .B(n21093), .Z(n21091) );
  NANDN U21182 ( .A(n21094), .B(n21095), .Z(n21093) );
  NANDN U21183 ( .A(n21095), .B(n21094), .Z(n21090) );
  ANDN U21184 ( .B(B[214]), .A(n62), .Z(n20874) );
  XNOR U21185 ( .A(n20882), .B(n21096), .Z(n20875) );
  XNOR U21186 ( .A(n20881), .B(n20879), .Z(n21096) );
  AND U21187 ( .A(n21097), .B(n21098), .Z(n20879) );
  NANDN U21188 ( .A(n21099), .B(n21100), .Z(n21098) );
  OR U21189 ( .A(n21101), .B(n21102), .Z(n21100) );
  NAND U21190 ( .A(n21102), .B(n21101), .Z(n21097) );
  ANDN U21191 ( .B(B[215]), .A(n63), .Z(n20881) );
  XNOR U21192 ( .A(n20889), .B(n21103), .Z(n20882) );
  XNOR U21193 ( .A(n20888), .B(n20886), .Z(n21103) );
  AND U21194 ( .A(n21104), .B(n21105), .Z(n20886) );
  NANDN U21195 ( .A(n21106), .B(n21107), .Z(n21105) );
  NANDN U21196 ( .A(n21108), .B(n21109), .Z(n21107) );
  NANDN U21197 ( .A(n21109), .B(n21108), .Z(n21104) );
  ANDN U21198 ( .B(B[216]), .A(n64), .Z(n20888) );
  XNOR U21199 ( .A(n20896), .B(n21110), .Z(n20889) );
  XNOR U21200 ( .A(n20895), .B(n20893), .Z(n21110) );
  AND U21201 ( .A(n21111), .B(n21112), .Z(n20893) );
  NANDN U21202 ( .A(n21113), .B(n21114), .Z(n21112) );
  OR U21203 ( .A(n21115), .B(n21116), .Z(n21114) );
  NAND U21204 ( .A(n21116), .B(n21115), .Z(n21111) );
  ANDN U21205 ( .B(B[217]), .A(n65), .Z(n20895) );
  XNOR U21206 ( .A(n20903), .B(n21117), .Z(n20896) );
  XNOR U21207 ( .A(n20902), .B(n20900), .Z(n21117) );
  AND U21208 ( .A(n21118), .B(n21119), .Z(n20900) );
  NANDN U21209 ( .A(n21120), .B(n21121), .Z(n21119) );
  NANDN U21210 ( .A(n21122), .B(n21123), .Z(n21121) );
  NANDN U21211 ( .A(n21123), .B(n21122), .Z(n21118) );
  ANDN U21212 ( .B(B[218]), .A(n66), .Z(n20902) );
  XNOR U21213 ( .A(n20910), .B(n21124), .Z(n20903) );
  XNOR U21214 ( .A(n20909), .B(n20907), .Z(n21124) );
  AND U21215 ( .A(n21125), .B(n21126), .Z(n20907) );
  NANDN U21216 ( .A(n21127), .B(n21128), .Z(n21126) );
  OR U21217 ( .A(n21129), .B(n21130), .Z(n21128) );
  NAND U21218 ( .A(n21130), .B(n21129), .Z(n21125) );
  ANDN U21219 ( .B(B[219]), .A(n67), .Z(n20909) );
  XNOR U21220 ( .A(n20917), .B(n21131), .Z(n20910) );
  XNOR U21221 ( .A(n20916), .B(n20914), .Z(n21131) );
  AND U21222 ( .A(n21132), .B(n21133), .Z(n20914) );
  NANDN U21223 ( .A(n21134), .B(n21135), .Z(n21133) );
  NANDN U21224 ( .A(n21136), .B(n21137), .Z(n21135) );
  NANDN U21225 ( .A(n21137), .B(n21136), .Z(n21132) );
  ANDN U21226 ( .B(B[220]), .A(n68), .Z(n20916) );
  XNOR U21227 ( .A(n20924), .B(n21138), .Z(n20917) );
  XNOR U21228 ( .A(n20923), .B(n20921), .Z(n21138) );
  AND U21229 ( .A(n21139), .B(n21140), .Z(n20921) );
  NANDN U21230 ( .A(n21141), .B(n21142), .Z(n21140) );
  OR U21231 ( .A(n21143), .B(n21144), .Z(n21142) );
  NAND U21232 ( .A(n21144), .B(n21143), .Z(n21139) );
  ANDN U21233 ( .B(B[221]), .A(n69), .Z(n20923) );
  XNOR U21234 ( .A(n20931), .B(n21145), .Z(n20924) );
  XNOR U21235 ( .A(n20930), .B(n20928), .Z(n21145) );
  AND U21236 ( .A(n21146), .B(n21147), .Z(n20928) );
  NANDN U21237 ( .A(n21148), .B(n21149), .Z(n21147) );
  NANDN U21238 ( .A(n21150), .B(n21151), .Z(n21149) );
  NANDN U21239 ( .A(n21151), .B(n21150), .Z(n21146) );
  ANDN U21240 ( .B(B[222]), .A(n70), .Z(n20930) );
  XNOR U21241 ( .A(n20938), .B(n21152), .Z(n20931) );
  XNOR U21242 ( .A(n20937), .B(n20935), .Z(n21152) );
  AND U21243 ( .A(n21153), .B(n21154), .Z(n20935) );
  NANDN U21244 ( .A(n21155), .B(n21156), .Z(n21154) );
  OR U21245 ( .A(n21157), .B(n21158), .Z(n21156) );
  NAND U21246 ( .A(n21158), .B(n21157), .Z(n21153) );
  ANDN U21247 ( .B(B[223]), .A(n71), .Z(n20937) );
  XNOR U21248 ( .A(n20945), .B(n21159), .Z(n20938) );
  XNOR U21249 ( .A(n20944), .B(n20942), .Z(n21159) );
  AND U21250 ( .A(n21160), .B(n21161), .Z(n20942) );
  NANDN U21251 ( .A(n21162), .B(n21163), .Z(n21161) );
  NANDN U21252 ( .A(n21164), .B(n21165), .Z(n21163) );
  NANDN U21253 ( .A(n21165), .B(n21164), .Z(n21160) );
  ANDN U21254 ( .B(B[224]), .A(n72), .Z(n20944) );
  XNOR U21255 ( .A(n20952), .B(n21166), .Z(n20945) );
  XNOR U21256 ( .A(n20951), .B(n20949), .Z(n21166) );
  AND U21257 ( .A(n21167), .B(n21168), .Z(n20949) );
  NANDN U21258 ( .A(n21169), .B(n21170), .Z(n21168) );
  OR U21259 ( .A(n21171), .B(n21172), .Z(n21170) );
  NAND U21260 ( .A(n21172), .B(n21171), .Z(n21167) );
  ANDN U21261 ( .B(B[225]), .A(n73), .Z(n20951) );
  XNOR U21262 ( .A(n20959), .B(n21173), .Z(n20952) );
  XNOR U21263 ( .A(n20958), .B(n20956), .Z(n21173) );
  AND U21264 ( .A(n21174), .B(n21175), .Z(n20956) );
  NANDN U21265 ( .A(n21176), .B(n21177), .Z(n21175) );
  NANDN U21266 ( .A(n21178), .B(n21179), .Z(n21177) );
  NANDN U21267 ( .A(n21179), .B(n21178), .Z(n21174) );
  ANDN U21268 ( .B(B[226]), .A(n74), .Z(n20958) );
  XNOR U21269 ( .A(n20966), .B(n21180), .Z(n20959) );
  XNOR U21270 ( .A(n20965), .B(n20963), .Z(n21180) );
  AND U21271 ( .A(n21181), .B(n21182), .Z(n20963) );
  NANDN U21272 ( .A(n21183), .B(n21184), .Z(n21182) );
  OR U21273 ( .A(n21185), .B(n21186), .Z(n21184) );
  NAND U21274 ( .A(n21186), .B(n21185), .Z(n21181) );
  ANDN U21275 ( .B(B[227]), .A(n75), .Z(n20965) );
  XNOR U21276 ( .A(n20973), .B(n21187), .Z(n20966) );
  XNOR U21277 ( .A(n20972), .B(n20970), .Z(n21187) );
  AND U21278 ( .A(n21188), .B(n21189), .Z(n20970) );
  NANDN U21279 ( .A(n21190), .B(n21191), .Z(n21189) );
  NANDN U21280 ( .A(n21192), .B(n21193), .Z(n21191) );
  NANDN U21281 ( .A(n21193), .B(n21192), .Z(n21188) );
  ANDN U21282 ( .B(B[228]), .A(n76), .Z(n20972) );
  XNOR U21283 ( .A(n20980), .B(n21194), .Z(n20973) );
  XNOR U21284 ( .A(n20979), .B(n20977), .Z(n21194) );
  AND U21285 ( .A(n21195), .B(n21196), .Z(n20977) );
  NANDN U21286 ( .A(n21197), .B(n21198), .Z(n21196) );
  OR U21287 ( .A(n21199), .B(n21200), .Z(n21198) );
  NAND U21288 ( .A(n21200), .B(n21199), .Z(n21195) );
  ANDN U21289 ( .B(B[229]), .A(n77), .Z(n20979) );
  XNOR U21290 ( .A(n20987), .B(n21201), .Z(n20980) );
  XNOR U21291 ( .A(n20986), .B(n20984), .Z(n21201) );
  AND U21292 ( .A(n21202), .B(n21203), .Z(n20984) );
  NANDN U21293 ( .A(n21204), .B(n21205), .Z(n21203) );
  NANDN U21294 ( .A(n21206), .B(n21207), .Z(n21205) );
  NANDN U21295 ( .A(n21207), .B(n21206), .Z(n21202) );
  ANDN U21296 ( .B(B[230]), .A(n78), .Z(n20986) );
  XNOR U21297 ( .A(n20994), .B(n21208), .Z(n20987) );
  XNOR U21298 ( .A(n20993), .B(n20991), .Z(n21208) );
  AND U21299 ( .A(n21209), .B(n21210), .Z(n20991) );
  NANDN U21300 ( .A(n21211), .B(n21212), .Z(n21210) );
  OR U21301 ( .A(n21213), .B(n21214), .Z(n21212) );
  NAND U21302 ( .A(n21214), .B(n21213), .Z(n21209) );
  ANDN U21303 ( .B(B[231]), .A(n79), .Z(n20993) );
  XNOR U21304 ( .A(n21001), .B(n21215), .Z(n20994) );
  XNOR U21305 ( .A(n21000), .B(n20998), .Z(n21215) );
  AND U21306 ( .A(n21216), .B(n21217), .Z(n20998) );
  NANDN U21307 ( .A(n21218), .B(n21219), .Z(n21217) );
  NANDN U21308 ( .A(n21220), .B(n21221), .Z(n21219) );
  NANDN U21309 ( .A(n21221), .B(n21220), .Z(n21216) );
  ANDN U21310 ( .B(B[232]), .A(n80), .Z(n21000) );
  XNOR U21311 ( .A(n21008), .B(n21222), .Z(n21001) );
  XNOR U21312 ( .A(n21007), .B(n21005), .Z(n21222) );
  AND U21313 ( .A(n21223), .B(n21224), .Z(n21005) );
  NANDN U21314 ( .A(n21225), .B(n21226), .Z(n21224) );
  OR U21315 ( .A(n21227), .B(n21228), .Z(n21226) );
  NAND U21316 ( .A(n21228), .B(n21227), .Z(n21223) );
  ANDN U21317 ( .B(B[233]), .A(n81), .Z(n21007) );
  XNOR U21318 ( .A(n21015), .B(n21229), .Z(n21008) );
  XNOR U21319 ( .A(n21014), .B(n21012), .Z(n21229) );
  AND U21320 ( .A(n21230), .B(n21231), .Z(n21012) );
  NANDN U21321 ( .A(n21232), .B(n21233), .Z(n21231) );
  NAND U21322 ( .A(n21234), .B(n21235), .Z(n21233) );
  ANDN U21323 ( .B(B[234]), .A(n82), .Z(n21014) );
  XOR U21324 ( .A(n21021), .B(n21236), .Z(n21015) );
  XNOR U21325 ( .A(n21019), .B(n21022), .Z(n21236) );
  NAND U21326 ( .A(A[2]), .B(B[235]), .Z(n21022) );
  NANDN U21327 ( .A(n21237), .B(n21238), .Z(n21019) );
  AND U21328 ( .A(A[0]), .B(B[236]), .Z(n21238) );
  XNOR U21329 ( .A(n21024), .B(n21239), .Z(n21021) );
  NAND U21330 ( .A(A[0]), .B(B[237]), .Z(n21239) );
  NAND U21331 ( .A(B[236]), .B(A[1]), .Z(n21024) );
  NAND U21332 ( .A(n21240), .B(n21241), .Z(n322) );
  NANDN U21333 ( .A(n21242), .B(n21243), .Z(n21241) );
  OR U21334 ( .A(n21244), .B(n21245), .Z(n21243) );
  NAND U21335 ( .A(n21245), .B(n21244), .Z(n21240) );
  XOR U21336 ( .A(n324), .B(n323), .Z(\A1[234] ) );
  XOR U21337 ( .A(n21245), .B(n21246), .Z(n323) );
  XNOR U21338 ( .A(n21244), .B(n21242), .Z(n21246) );
  AND U21339 ( .A(n21247), .B(n21248), .Z(n21242) );
  NANDN U21340 ( .A(n21249), .B(n21250), .Z(n21248) );
  NANDN U21341 ( .A(n21251), .B(n21252), .Z(n21250) );
  NANDN U21342 ( .A(n21252), .B(n21251), .Z(n21247) );
  ANDN U21343 ( .B(B[205]), .A(n54), .Z(n21244) );
  XNOR U21344 ( .A(n21039), .B(n21253), .Z(n21245) );
  XNOR U21345 ( .A(n21038), .B(n21036), .Z(n21253) );
  AND U21346 ( .A(n21254), .B(n21255), .Z(n21036) );
  NANDN U21347 ( .A(n21256), .B(n21257), .Z(n21255) );
  OR U21348 ( .A(n21258), .B(n21259), .Z(n21257) );
  NAND U21349 ( .A(n21259), .B(n21258), .Z(n21254) );
  ANDN U21350 ( .B(B[206]), .A(n55), .Z(n21038) );
  XNOR U21351 ( .A(n21046), .B(n21260), .Z(n21039) );
  XNOR U21352 ( .A(n21045), .B(n21043), .Z(n21260) );
  AND U21353 ( .A(n21261), .B(n21262), .Z(n21043) );
  NANDN U21354 ( .A(n21263), .B(n21264), .Z(n21262) );
  NANDN U21355 ( .A(n21265), .B(n21266), .Z(n21264) );
  NANDN U21356 ( .A(n21266), .B(n21265), .Z(n21261) );
  ANDN U21357 ( .B(B[207]), .A(n56), .Z(n21045) );
  XNOR U21358 ( .A(n21053), .B(n21267), .Z(n21046) );
  XNOR U21359 ( .A(n21052), .B(n21050), .Z(n21267) );
  AND U21360 ( .A(n21268), .B(n21269), .Z(n21050) );
  NANDN U21361 ( .A(n21270), .B(n21271), .Z(n21269) );
  OR U21362 ( .A(n21272), .B(n21273), .Z(n21271) );
  NAND U21363 ( .A(n21273), .B(n21272), .Z(n21268) );
  ANDN U21364 ( .B(B[208]), .A(n57), .Z(n21052) );
  XNOR U21365 ( .A(n21060), .B(n21274), .Z(n21053) );
  XNOR U21366 ( .A(n21059), .B(n21057), .Z(n21274) );
  AND U21367 ( .A(n21275), .B(n21276), .Z(n21057) );
  NANDN U21368 ( .A(n21277), .B(n21278), .Z(n21276) );
  NANDN U21369 ( .A(n21279), .B(n21280), .Z(n21278) );
  NANDN U21370 ( .A(n21280), .B(n21279), .Z(n21275) );
  ANDN U21371 ( .B(B[209]), .A(n58), .Z(n21059) );
  XNOR U21372 ( .A(n21067), .B(n21281), .Z(n21060) );
  XNOR U21373 ( .A(n21066), .B(n21064), .Z(n21281) );
  AND U21374 ( .A(n21282), .B(n21283), .Z(n21064) );
  NANDN U21375 ( .A(n21284), .B(n21285), .Z(n21283) );
  OR U21376 ( .A(n21286), .B(n21287), .Z(n21285) );
  NAND U21377 ( .A(n21287), .B(n21286), .Z(n21282) );
  ANDN U21378 ( .B(B[210]), .A(n59), .Z(n21066) );
  XNOR U21379 ( .A(n21074), .B(n21288), .Z(n21067) );
  XNOR U21380 ( .A(n21073), .B(n21071), .Z(n21288) );
  AND U21381 ( .A(n21289), .B(n21290), .Z(n21071) );
  NANDN U21382 ( .A(n21291), .B(n21292), .Z(n21290) );
  NANDN U21383 ( .A(n21293), .B(n21294), .Z(n21292) );
  NANDN U21384 ( .A(n21294), .B(n21293), .Z(n21289) );
  ANDN U21385 ( .B(B[211]), .A(n60), .Z(n21073) );
  XNOR U21386 ( .A(n21081), .B(n21295), .Z(n21074) );
  XNOR U21387 ( .A(n21080), .B(n21078), .Z(n21295) );
  AND U21388 ( .A(n21296), .B(n21297), .Z(n21078) );
  NANDN U21389 ( .A(n21298), .B(n21299), .Z(n21297) );
  OR U21390 ( .A(n21300), .B(n21301), .Z(n21299) );
  NAND U21391 ( .A(n21301), .B(n21300), .Z(n21296) );
  ANDN U21392 ( .B(B[212]), .A(n61), .Z(n21080) );
  XNOR U21393 ( .A(n21088), .B(n21302), .Z(n21081) );
  XNOR U21394 ( .A(n21087), .B(n21085), .Z(n21302) );
  AND U21395 ( .A(n21303), .B(n21304), .Z(n21085) );
  NANDN U21396 ( .A(n21305), .B(n21306), .Z(n21304) );
  NANDN U21397 ( .A(n21307), .B(n21308), .Z(n21306) );
  NANDN U21398 ( .A(n21308), .B(n21307), .Z(n21303) );
  ANDN U21399 ( .B(B[213]), .A(n62), .Z(n21087) );
  XNOR U21400 ( .A(n21095), .B(n21309), .Z(n21088) );
  XNOR U21401 ( .A(n21094), .B(n21092), .Z(n21309) );
  AND U21402 ( .A(n21310), .B(n21311), .Z(n21092) );
  NANDN U21403 ( .A(n21312), .B(n21313), .Z(n21311) );
  OR U21404 ( .A(n21314), .B(n21315), .Z(n21313) );
  NAND U21405 ( .A(n21315), .B(n21314), .Z(n21310) );
  ANDN U21406 ( .B(B[214]), .A(n63), .Z(n21094) );
  XNOR U21407 ( .A(n21102), .B(n21316), .Z(n21095) );
  XNOR U21408 ( .A(n21101), .B(n21099), .Z(n21316) );
  AND U21409 ( .A(n21317), .B(n21318), .Z(n21099) );
  NANDN U21410 ( .A(n21319), .B(n21320), .Z(n21318) );
  NANDN U21411 ( .A(n21321), .B(n21322), .Z(n21320) );
  NANDN U21412 ( .A(n21322), .B(n21321), .Z(n21317) );
  ANDN U21413 ( .B(B[215]), .A(n64), .Z(n21101) );
  XNOR U21414 ( .A(n21109), .B(n21323), .Z(n21102) );
  XNOR U21415 ( .A(n21108), .B(n21106), .Z(n21323) );
  AND U21416 ( .A(n21324), .B(n21325), .Z(n21106) );
  NANDN U21417 ( .A(n21326), .B(n21327), .Z(n21325) );
  OR U21418 ( .A(n21328), .B(n21329), .Z(n21327) );
  NAND U21419 ( .A(n21329), .B(n21328), .Z(n21324) );
  ANDN U21420 ( .B(B[216]), .A(n65), .Z(n21108) );
  XNOR U21421 ( .A(n21116), .B(n21330), .Z(n21109) );
  XNOR U21422 ( .A(n21115), .B(n21113), .Z(n21330) );
  AND U21423 ( .A(n21331), .B(n21332), .Z(n21113) );
  NANDN U21424 ( .A(n21333), .B(n21334), .Z(n21332) );
  NANDN U21425 ( .A(n21335), .B(n21336), .Z(n21334) );
  NANDN U21426 ( .A(n21336), .B(n21335), .Z(n21331) );
  ANDN U21427 ( .B(B[217]), .A(n66), .Z(n21115) );
  XNOR U21428 ( .A(n21123), .B(n21337), .Z(n21116) );
  XNOR U21429 ( .A(n21122), .B(n21120), .Z(n21337) );
  AND U21430 ( .A(n21338), .B(n21339), .Z(n21120) );
  NANDN U21431 ( .A(n21340), .B(n21341), .Z(n21339) );
  OR U21432 ( .A(n21342), .B(n21343), .Z(n21341) );
  NAND U21433 ( .A(n21343), .B(n21342), .Z(n21338) );
  ANDN U21434 ( .B(B[218]), .A(n67), .Z(n21122) );
  XNOR U21435 ( .A(n21130), .B(n21344), .Z(n21123) );
  XNOR U21436 ( .A(n21129), .B(n21127), .Z(n21344) );
  AND U21437 ( .A(n21345), .B(n21346), .Z(n21127) );
  NANDN U21438 ( .A(n21347), .B(n21348), .Z(n21346) );
  NANDN U21439 ( .A(n21349), .B(n21350), .Z(n21348) );
  NANDN U21440 ( .A(n21350), .B(n21349), .Z(n21345) );
  ANDN U21441 ( .B(B[219]), .A(n68), .Z(n21129) );
  XNOR U21442 ( .A(n21137), .B(n21351), .Z(n21130) );
  XNOR U21443 ( .A(n21136), .B(n21134), .Z(n21351) );
  AND U21444 ( .A(n21352), .B(n21353), .Z(n21134) );
  NANDN U21445 ( .A(n21354), .B(n21355), .Z(n21353) );
  OR U21446 ( .A(n21356), .B(n21357), .Z(n21355) );
  NAND U21447 ( .A(n21357), .B(n21356), .Z(n21352) );
  ANDN U21448 ( .B(B[220]), .A(n69), .Z(n21136) );
  XNOR U21449 ( .A(n21144), .B(n21358), .Z(n21137) );
  XNOR U21450 ( .A(n21143), .B(n21141), .Z(n21358) );
  AND U21451 ( .A(n21359), .B(n21360), .Z(n21141) );
  NANDN U21452 ( .A(n21361), .B(n21362), .Z(n21360) );
  NANDN U21453 ( .A(n21363), .B(n21364), .Z(n21362) );
  NANDN U21454 ( .A(n21364), .B(n21363), .Z(n21359) );
  ANDN U21455 ( .B(B[221]), .A(n70), .Z(n21143) );
  XNOR U21456 ( .A(n21151), .B(n21365), .Z(n21144) );
  XNOR U21457 ( .A(n21150), .B(n21148), .Z(n21365) );
  AND U21458 ( .A(n21366), .B(n21367), .Z(n21148) );
  NANDN U21459 ( .A(n21368), .B(n21369), .Z(n21367) );
  OR U21460 ( .A(n21370), .B(n21371), .Z(n21369) );
  NAND U21461 ( .A(n21371), .B(n21370), .Z(n21366) );
  ANDN U21462 ( .B(B[222]), .A(n71), .Z(n21150) );
  XNOR U21463 ( .A(n21158), .B(n21372), .Z(n21151) );
  XNOR U21464 ( .A(n21157), .B(n21155), .Z(n21372) );
  AND U21465 ( .A(n21373), .B(n21374), .Z(n21155) );
  NANDN U21466 ( .A(n21375), .B(n21376), .Z(n21374) );
  NANDN U21467 ( .A(n21377), .B(n21378), .Z(n21376) );
  NANDN U21468 ( .A(n21378), .B(n21377), .Z(n21373) );
  ANDN U21469 ( .B(B[223]), .A(n72), .Z(n21157) );
  XNOR U21470 ( .A(n21165), .B(n21379), .Z(n21158) );
  XNOR U21471 ( .A(n21164), .B(n21162), .Z(n21379) );
  AND U21472 ( .A(n21380), .B(n21381), .Z(n21162) );
  NANDN U21473 ( .A(n21382), .B(n21383), .Z(n21381) );
  OR U21474 ( .A(n21384), .B(n21385), .Z(n21383) );
  NAND U21475 ( .A(n21385), .B(n21384), .Z(n21380) );
  ANDN U21476 ( .B(B[224]), .A(n73), .Z(n21164) );
  XNOR U21477 ( .A(n21172), .B(n21386), .Z(n21165) );
  XNOR U21478 ( .A(n21171), .B(n21169), .Z(n21386) );
  AND U21479 ( .A(n21387), .B(n21388), .Z(n21169) );
  NANDN U21480 ( .A(n21389), .B(n21390), .Z(n21388) );
  NANDN U21481 ( .A(n21391), .B(n21392), .Z(n21390) );
  NANDN U21482 ( .A(n21392), .B(n21391), .Z(n21387) );
  ANDN U21483 ( .B(B[225]), .A(n74), .Z(n21171) );
  XNOR U21484 ( .A(n21179), .B(n21393), .Z(n21172) );
  XNOR U21485 ( .A(n21178), .B(n21176), .Z(n21393) );
  AND U21486 ( .A(n21394), .B(n21395), .Z(n21176) );
  NANDN U21487 ( .A(n21396), .B(n21397), .Z(n21395) );
  OR U21488 ( .A(n21398), .B(n21399), .Z(n21397) );
  NAND U21489 ( .A(n21399), .B(n21398), .Z(n21394) );
  ANDN U21490 ( .B(B[226]), .A(n75), .Z(n21178) );
  XNOR U21491 ( .A(n21186), .B(n21400), .Z(n21179) );
  XNOR U21492 ( .A(n21185), .B(n21183), .Z(n21400) );
  AND U21493 ( .A(n21401), .B(n21402), .Z(n21183) );
  NANDN U21494 ( .A(n21403), .B(n21404), .Z(n21402) );
  NANDN U21495 ( .A(n21405), .B(n21406), .Z(n21404) );
  NANDN U21496 ( .A(n21406), .B(n21405), .Z(n21401) );
  ANDN U21497 ( .B(B[227]), .A(n76), .Z(n21185) );
  XNOR U21498 ( .A(n21193), .B(n21407), .Z(n21186) );
  XNOR U21499 ( .A(n21192), .B(n21190), .Z(n21407) );
  AND U21500 ( .A(n21408), .B(n21409), .Z(n21190) );
  NANDN U21501 ( .A(n21410), .B(n21411), .Z(n21409) );
  OR U21502 ( .A(n21412), .B(n21413), .Z(n21411) );
  NAND U21503 ( .A(n21413), .B(n21412), .Z(n21408) );
  ANDN U21504 ( .B(B[228]), .A(n77), .Z(n21192) );
  XNOR U21505 ( .A(n21200), .B(n21414), .Z(n21193) );
  XNOR U21506 ( .A(n21199), .B(n21197), .Z(n21414) );
  AND U21507 ( .A(n21415), .B(n21416), .Z(n21197) );
  NANDN U21508 ( .A(n21417), .B(n21418), .Z(n21416) );
  NANDN U21509 ( .A(n21419), .B(n21420), .Z(n21418) );
  NANDN U21510 ( .A(n21420), .B(n21419), .Z(n21415) );
  ANDN U21511 ( .B(B[229]), .A(n78), .Z(n21199) );
  XNOR U21512 ( .A(n21207), .B(n21421), .Z(n21200) );
  XNOR U21513 ( .A(n21206), .B(n21204), .Z(n21421) );
  AND U21514 ( .A(n21422), .B(n21423), .Z(n21204) );
  NANDN U21515 ( .A(n21424), .B(n21425), .Z(n21423) );
  OR U21516 ( .A(n21426), .B(n21427), .Z(n21425) );
  NAND U21517 ( .A(n21427), .B(n21426), .Z(n21422) );
  ANDN U21518 ( .B(B[230]), .A(n79), .Z(n21206) );
  XNOR U21519 ( .A(n21214), .B(n21428), .Z(n21207) );
  XNOR U21520 ( .A(n21213), .B(n21211), .Z(n21428) );
  AND U21521 ( .A(n21429), .B(n21430), .Z(n21211) );
  NANDN U21522 ( .A(n21431), .B(n21432), .Z(n21430) );
  NANDN U21523 ( .A(n21433), .B(n21434), .Z(n21432) );
  NANDN U21524 ( .A(n21434), .B(n21433), .Z(n21429) );
  ANDN U21525 ( .B(B[231]), .A(n80), .Z(n21213) );
  XNOR U21526 ( .A(n21221), .B(n21435), .Z(n21214) );
  XNOR U21527 ( .A(n21220), .B(n21218), .Z(n21435) );
  AND U21528 ( .A(n21436), .B(n21437), .Z(n21218) );
  NANDN U21529 ( .A(n21438), .B(n21439), .Z(n21437) );
  OR U21530 ( .A(n21440), .B(n21441), .Z(n21439) );
  NAND U21531 ( .A(n21441), .B(n21440), .Z(n21436) );
  ANDN U21532 ( .B(B[232]), .A(n81), .Z(n21220) );
  XNOR U21533 ( .A(n21228), .B(n21442), .Z(n21221) );
  XNOR U21534 ( .A(n21227), .B(n21225), .Z(n21442) );
  AND U21535 ( .A(n21443), .B(n21444), .Z(n21225) );
  NANDN U21536 ( .A(n21445), .B(n21446), .Z(n21444) );
  NAND U21537 ( .A(n21447), .B(n21448), .Z(n21446) );
  ANDN U21538 ( .B(B[233]), .A(n82), .Z(n21227) );
  XOR U21539 ( .A(n21234), .B(n21449), .Z(n21228) );
  XNOR U21540 ( .A(n21232), .B(n21235), .Z(n21449) );
  NAND U21541 ( .A(A[2]), .B(B[234]), .Z(n21235) );
  NANDN U21542 ( .A(n21450), .B(n21451), .Z(n21232) );
  AND U21543 ( .A(A[0]), .B(B[235]), .Z(n21451) );
  XNOR U21544 ( .A(n21237), .B(n21452), .Z(n21234) );
  NAND U21545 ( .A(A[0]), .B(B[236]), .Z(n21452) );
  NAND U21546 ( .A(B[235]), .B(A[1]), .Z(n21237) );
  NAND U21547 ( .A(n21453), .B(n21454), .Z(n324) );
  NANDN U21548 ( .A(n21455), .B(n21456), .Z(n21454) );
  OR U21549 ( .A(n21457), .B(n21458), .Z(n21456) );
  NAND U21550 ( .A(n21458), .B(n21457), .Z(n21453) );
  XOR U21551 ( .A(n326), .B(n325), .Z(\A1[233] ) );
  XOR U21552 ( .A(n21458), .B(n21459), .Z(n325) );
  XNOR U21553 ( .A(n21457), .B(n21455), .Z(n21459) );
  AND U21554 ( .A(n21460), .B(n21461), .Z(n21455) );
  NANDN U21555 ( .A(n21462), .B(n21463), .Z(n21461) );
  NANDN U21556 ( .A(n21464), .B(n21465), .Z(n21463) );
  NANDN U21557 ( .A(n21465), .B(n21464), .Z(n21460) );
  ANDN U21558 ( .B(B[204]), .A(n54), .Z(n21457) );
  XNOR U21559 ( .A(n21252), .B(n21466), .Z(n21458) );
  XNOR U21560 ( .A(n21251), .B(n21249), .Z(n21466) );
  AND U21561 ( .A(n21467), .B(n21468), .Z(n21249) );
  NANDN U21562 ( .A(n21469), .B(n21470), .Z(n21468) );
  OR U21563 ( .A(n21471), .B(n21472), .Z(n21470) );
  NAND U21564 ( .A(n21472), .B(n21471), .Z(n21467) );
  ANDN U21565 ( .B(B[205]), .A(n55), .Z(n21251) );
  XNOR U21566 ( .A(n21259), .B(n21473), .Z(n21252) );
  XNOR U21567 ( .A(n21258), .B(n21256), .Z(n21473) );
  AND U21568 ( .A(n21474), .B(n21475), .Z(n21256) );
  NANDN U21569 ( .A(n21476), .B(n21477), .Z(n21475) );
  NANDN U21570 ( .A(n21478), .B(n21479), .Z(n21477) );
  NANDN U21571 ( .A(n21479), .B(n21478), .Z(n21474) );
  ANDN U21572 ( .B(B[206]), .A(n56), .Z(n21258) );
  XNOR U21573 ( .A(n21266), .B(n21480), .Z(n21259) );
  XNOR U21574 ( .A(n21265), .B(n21263), .Z(n21480) );
  AND U21575 ( .A(n21481), .B(n21482), .Z(n21263) );
  NANDN U21576 ( .A(n21483), .B(n21484), .Z(n21482) );
  OR U21577 ( .A(n21485), .B(n21486), .Z(n21484) );
  NAND U21578 ( .A(n21486), .B(n21485), .Z(n21481) );
  ANDN U21579 ( .B(B[207]), .A(n57), .Z(n21265) );
  XNOR U21580 ( .A(n21273), .B(n21487), .Z(n21266) );
  XNOR U21581 ( .A(n21272), .B(n21270), .Z(n21487) );
  AND U21582 ( .A(n21488), .B(n21489), .Z(n21270) );
  NANDN U21583 ( .A(n21490), .B(n21491), .Z(n21489) );
  NANDN U21584 ( .A(n21492), .B(n21493), .Z(n21491) );
  NANDN U21585 ( .A(n21493), .B(n21492), .Z(n21488) );
  ANDN U21586 ( .B(B[208]), .A(n58), .Z(n21272) );
  XNOR U21587 ( .A(n21280), .B(n21494), .Z(n21273) );
  XNOR U21588 ( .A(n21279), .B(n21277), .Z(n21494) );
  AND U21589 ( .A(n21495), .B(n21496), .Z(n21277) );
  NANDN U21590 ( .A(n21497), .B(n21498), .Z(n21496) );
  OR U21591 ( .A(n21499), .B(n21500), .Z(n21498) );
  NAND U21592 ( .A(n21500), .B(n21499), .Z(n21495) );
  ANDN U21593 ( .B(B[209]), .A(n59), .Z(n21279) );
  XNOR U21594 ( .A(n21287), .B(n21501), .Z(n21280) );
  XNOR U21595 ( .A(n21286), .B(n21284), .Z(n21501) );
  AND U21596 ( .A(n21502), .B(n21503), .Z(n21284) );
  NANDN U21597 ( .A(n21504), .B(n21505), .Z(n21503) );
  NANDN U21598 ( .A(n21506), .B(n21507), .Z(n21505) );
  NANDN U21599 ( .A(n21507), .B(n21506), .Z(n21502) );
  ANDN U21600 ( .B(B[210]), .A(n60), .Z(n21286) );
  XNOR U21601 ( .A(n21294), .B(n21508), .Z(n21287) );
  XNOR U21602 ( .A(n21293), .B(n21291), .Z(n21508) );
  AND U21603 ( .A(n21509), .B(n21510), .Z(n21291) );
  NANDN U21604 ( .A(n21511), .B(n21512), .Z(n21510) );
  OR U21605 ( .A(n21513), .B(n21514), .Z(n21512) );
  NAND U21606 ( .A(n21514), .B(n21513), .Z(n21509) );
  ANDN U21607 ( .B(B[211]), .A(n61), .Z(n21293) );
  XNOR U21608 ( .A(n21301), .B(n21515), .Z(n21294) );
  XNOR U21609 ( .A(n21300), .B(n21298), .Z(n21515) );
  AND U21610 ( .A(n21516), .B(n21517), .Z(n21298) );
  NANDN U21611 ( .A(n21518), .B(n21519), .Z(n21517) );
  NANDN U21612 ( .A(n21520), .B(n21521), .Z(n21519) );
  NANDN U21613 ( .A(n21521), .B(n21520), .Z(n21516) );
  ANDN U21614 ( .B(B[212]), .A(n62), .Z(n21300) );
  XNOR U21615 ( .A(n21308), .B(n21522), .Z(n21301) );
  XNOR U21616 ( .A(n21307), .B(n21305), .Z(n21522) );
  AND U21617 ( .A(n21523), .B(n21524), .Z(n21305) );
  NANDN U21618 ( .A(n21525), .B(n21526), .Z(n21524) );
  OR U21619 ( .A(n21527), .B(n21528), .Z(n21526) );
  NAND U21620 ( .A(n21528), .B(n21527), .Z(n21523) );
  ANDN U21621 ( .B(B[213]), .A(n63), .Z(n21307) );
  XNOR U21622 ( .A(n21315), .B(n21529), .Z(n21308) );
  XNOR U21623 ( .A(n21314), .B(n21312), .Z(n21529) );
  AND U21624 ( .A(n21530), .B(n21531), .Z(n21312) );
  NANDN U21625 ( .A(n21532), .B(n21533), .Z(n21531) );
  NANDN U21626 ( .A(n21534), .B(n21535), .Z(n21533) );
  NANDN U21627 ( .A(n21535), .B(n21534), .Z(n21530) );
  ANDN U21628 ( .B(B[214]), .A(n64), .Z(n21314) );
  XNOR U21629 ( .A(n21322), .B(n21536), .Z(n21315) );
  XNOR U21630 ( .A(n21321), .B(n21319), .Z(n21536) );
  AND U21631 ( .A(n21537), .B(n21538), .Z(n21319) );
  NANDN U21632 ( .A(n21539), .B(n21540), .Z(n21538) );
  OR U21633 ( .A(n21541), .B(n21542), .Z(n21540) );
  NAND U21634 ( .A(n21542), .B(n21541), .Z(n21537) );
  ANDN U21635 ( .B(B[215]), .A(n65), .Z(n21321) );
  XNOR U21636 ( .A(n21329), .B(n21543), .Z(n21322) );
  XNOR U21637 ( .A(n21328), .B(n21326), .Z(n21543) );
  AND U21638 ( .A(n21544), .B(n21545), .Z(n21326) );
  NANDN U21639 ( .A(n21546), .B(n21547), .Z(n21545) );
  NANDN U21640 ( .A(n21548), .B(n21549), .Z(n21547) );
  NANDN U21641 ( .A(n21549), .B(n21548), .Z(n21544) );
  ANDN U21642 ( .B(B[216]), .A(n66), .Z(n21328) );
  XNOR U21643 ( .A(n21336), .B(n21550), .Z(n21329) );
  XNOR U21644 ( .A(n21335), .B(n21333), .Z(n21550) );
  AND U21645 ( .A(n21551), .B(n21552), .Z(n21333) );
  NANDN U21646 ( .A(n21553), .B(n21554), .Z(n21552) );
  OR U21647 ( .A(n21555), .B(n21556), .Z(n21554) );
  NAND U21648 ( .A(n21556), .B(n21555), .Z(n21551) );
  ANDN U21649 ( .B(B[217]), .A(n67), .Z(n21335) );
  XNOR U21650 ( .A(n21343), .B(n21557), .Z(n21336) );
  XNOR U21651 ( .A(n21342), .B(n21340), .Z(n21557) );
  AND U21652 ( .A(n21558), .B(n21559), .Z(n21340) );
  NANDN U21653 ( .A(n21560), .B(n21561), .Z(n21559) );
  NANDN U21654 ( .A(n21562), .B(n21563), .Z(n21561) );
  NANDN U21655 ( .A(n21563), .B(n21562), .Z(n21558) );
  ANDN U21656 ( .B(B[218]), .A(n68), .Z(n21342) );
  XNOR U21657 ( .A(n21350), .B(n21564), .Z(n21343) );
  XNOR U21658 ( .A(n21349), .B(n21347), .Z(n21564) );
  AND U21659 ( .A(n21565), .B(n21566), .Z(n21347) );
  NANDN U21660 ( .A(n21567), .B(n21568), .Z(n21566) );
  OR U21661 ( .A(n21569), .B(n21570), .Z(n21568) );
  NAND U21662 ( .A(n21570), .B(n21569), .Z(n21565) );
  ANDN U21663 ( .B(B[219]), .A(n69), .Z(n21349) );
  XNOR U21664 ( .A(n21357), .B(n21571), .Z(n21350) );
  XNOR U21665 ( .A(n21356), .B(n21354), .Z(n21571) );
  AND U21666 ( .A(n21572), .B(n21573), .Z(n21354) );
  NANDN U21667 ( .A(n21574), .B(n21575), .Z(n21573) );
  NANDN U21668 ( .A(n21576), .B(n21577), .Z(n21575) );
  NANDN U21669 ( .A(n21577), .B(n21576), .Z(n21572) );
  ANDN U21670 ( .B(B[220]), .A(n70), .Z(n21356) );
  XNOR U21671 ( .A(n21364), .B(n21578), .Z(n21357) );
  XNOR U21672 ( .A(n21363), .B(n21361), .Z(n21578) );
  AND U21673 ( .A(n21579), .B(n21580), .Z(n21361) );
  NANDN U21674 ( .A(n21581), .B(n21582), .Z(n21580) );
  OR U21675 ( .A(n21583), .B(n21584), .Z(n21582) );
  NAND U21676 ( .A(n21584), .B(n21583), .Z(n21579) );
  ANDN U21677 ( .B(B[221]), .A(n71), .Z(n21363) );
  XNOR U21678 ( .A(n21371), .B(n21585), .Z(n21364) );
  XNOR U21679 ( .A(n21370), .B(n21368), .Z(n21585) );
  AND U21680 ( .A(n21586), .B(n21587), .Z(n21368) );
  NANDN U21681 ( .A(n21588), .B(n21589), .Z(n21587) );
  NANDN U21682 ( .A(n21590), .B(n21591), .Z(n21589) );
  NANDN U21683 ( .A(n21591), .B(n21590), .Z(n21586) );
  ANDN U21684 ( .B(B[222]), .A(n72), .Z(n21370) );
  XNOR U21685 ( .A(n21378), .B(n21592), .Z(n21371) );
  XNOR U21686 ( .A(n21377), .B(n21375), .Z(n21592) );
  AND U21687 ( .A(n21593), .B(n21594), .Z(n21375) );
  NANDN U21688 ( .A(n21595), .B(n21596), .Z(n21594) );
  OR U21689 ( .A(n21597), .B(n21598), .Z(n21596) );
  NAND U21690 ( .A(n21598), .B(n21597), .Z(n21593) );
  ANDN U21691 ( .B(B[223]), .A(n73), .Z(n21377) );
  XNOR U21692 ( .A(n21385), .B(n21599), .Z(n21378) );
  XNOR U21693 ( .A(n21384), .B(n21382), .Z(n21599) );
  AND U21694 ( .A(n21600), .B(n21601), .Z(n21382) );
  NANDN U21695 ( .A(n21602), .B(n21603), .Z(n21601) );
  NANDN U21696 ( .A(n21604), .B(n21605), .Z(n21603) );
  NANDN U21697 ( .A(n21605), .B(n21604), .Z(n21600) );
  ANDN U21698 ( .B(B[224]), .A(n74), .Z(n21384) );
  XNOR U21699 ( .A(n21392), .B(n21606), .Z(n21385) );
  XNOR U21700 ( .A(n21391), .B(n21389), .Z(n21606) );
  AND U21701 ( .A(n21607), .B(n21608), .Z(n21389) );
  NANDN U21702 ( .A(n21609), .B(n21610), .Z(n21608) );
  OR U21703 ( .A(n21611), .B(n21612), .Z(n21610) );
  NAND U21704 ( .A(n21612), .B(n21611), .Z(n21607) );
  ANDN U21705 ( .B(B[225]), .A(n75), .Z(n21391) );
  XNOR U21706 ( .A(n21399), .B(n21613), .Z(n21392) );
  XNOR U21707 ( .A(n21398), .B(n21396), .Z(n21613) );
  AND U21708 ( .A(n21614), .B(n21615), .Z(n21396) );
  NANDN U21709 ( .A(n21616), .B(n21617), .Z(n21615) );
  NANDN U21710 ( .A(n21618), .B(n21619), .Z(n21617) );
  NANDN U21711 ( .A(n21619), .B(n21618), .Z(n21614) );
  ANDN U21712 ( .B(B[226]), .A(n76), .Z(n21398) );
  XNOR U21713 ( .A(n21406), .B(n21620), .Z(n21399) );
  XNOR U21714 ( .A(n21405), .B(n21403), .Z(n21620) );
  AND U21715 ( .A(n21621), .B(n21622), .Z(n21403) );
  NANDN U21716 ( .A(n21623), .B(n21624), .Z(n21622) );
  OR U21717 ( .A(n21625), .B(n21626), .Z(n21624) );
  NAND U21718 ( .A(n21626), .B(n21625), .Z(n21621) );
  ANDN U21719 ( .B(B[227]), .A(n77), .Z(n21405) );
  XNOR U21720 ( .A(n21413), .B(n21627), .Z(n21406) );
  XNOR U21721 ( .A(n21412), .B(n21410), .Z(n21627) );
  AND U21722 ( .A(n21628), .B(n21629), .Z(n21410) );
  NANDN U21723 ( .A(n21630), .B(n21631), .Z(n21629) );
  NANDN U21724 ( .A(n21632), .B(n21633), .Z(n21631) );
  NANDN U21725 ( .A(n21633), .B(n21632), .Z(n21628) );
  ANDN U21726 ( .B(B[228]), .A(n78), .Z(n21412) );
  XNOR U21727 ( .A(n21420), .B(n21634), .Z(n21413) );
  XNOR U21728 ( .A(n21419), .B(n21417), .Z(n21634) );
  AND U21729 ( .A(n21635), .B(n21636), .Z(n21417) );
  NANDN U21730 ( .A(n21637), .B(n21638), .Z(n21636) );
  OR U21731 ( .A(n21639), .B(n21640), .Z(n21638) );
  NAND U21732 ( .A(n21640), .B(n21639), .Z(n21635) );
  ANDN U21733 ( .B(B[229]), .A(n79), .Z(n21419) );
  XNOR U21734 ( .A(n21427), .B(n21641), .Z(n21420) );
  XNOR U21735 ( .A(n21426), .B(n21424), .Z(n21641) );
  AND U21736 ( .A(n21642), .B(n21643), .Z(n21424) );
  NANDN U21737 ( .A(n21644), .B(n21645), .Z(n21643) );
  NANDN U21738 ( .A(n21646), .B(n21647), .Z(n21645) );
  NANDN U21739 ( .A(n21647), .B(n21646), .Z(n21642) );
  ANDN U21740 ( .B(B[230]), .A(n80), .Z(n21426) );
  XNOR U21741 ( .A(n21434), .B(n21648), .Z(n21427) );
  XNOR U21742 ( .A(n21433), .B(n21431), .Z(n21648) );
  AND U21743 ( .A(n21649), .B(n21650), .Z(n21431) );
  NANDN U21744 ( .A(n21651), .B(n21652), .Z(n21650) );
  OR U21745 ( .A(n21653), .B(n21654), .Z(n21652) );
  NAND U21746 ( .A(n21654), .B(n21653), .Z(n21649) );
  ANDN U21747 ( .B(B[231]), .A(n81), .Z(n21433) );
  XNOR U21748 ( .A(n21441), .B(n21655), .Z(n21434) );
  XNOR U21749 ( .A(n21440), .B(n21438), .Z(n21655) );
  AND U21750 ( .A(n21656), .B(n21657), .Z(n21438) );
  NANDN U21751 ( .A(n21658), .B(n21659), .Z(n21657) );
  NAND U21752 ( .A(n21660), .B(n21661), .Z(n21659) );
  ANDN U21753 ( .B(B[232]), .A(n82), .Z(n21440) );
  XOR U21754 ( .A(n21447), .B(n21662), .Z(n21441) );
  XNOR U21755 ( .A(n21445), .B(n21448), .Z(n21662) );
  NAND U21756 ( .A(A[2]), .B(B[233]), .Z(n21448) );
  NANDN U21757 ( .A(n21663), .B(n21664), .Z(n21445) );
  AND U21758 ( .A(A[0]), .B(B[234]), .Z(n21664) );
  XNOR U21759 ( .A(n21450), .B(n21665), .Z(n21447) );
  NAND U21760 ( .A(A[0]), .B(B[235]), .Z(n21665) );
  NAND U21761 ( .A(B[234]), .B(A[1]), .Z(n21450) );
  NAND U21762 ( .A(n21666), .B(n21667), .Z(n326) );
  NANDN U21763 ( .A(n21668), .B(n21669), .Z(n21667) );
  OR U21764 ( .A(n21670), .B(n21671), .Z(n21669) );
  NAND U21765 ( .A(n21671), .B(n21670), .Z(n21666) );
  XOR U21766 ( .A(n328), .B(n327), .Z(\A1[232] ) );
  XOR U21767 ( .A(n21671), .B(n21672), .Z(n327) );
  XNOR U21768 ( .A(n21670), .B(n21668), .Z(n21672) );
  AND U21769 ( .A(n21673), .B(n21674), .Z(n21668) );
  NANDN U21770 ( .A(n21675), .B(n21676), .Z(n21674) );
  NANDN U21771 ( .A(n21677), .B(n21678), .Z(n21676) );
  NANDN U21772 ( .A(n21678), .B(n21677), .Z(n21673) );
  ANDN U21773 ( .B(B[203]), .A(n54), .Z(n21670) );
  XNOR U21774 ( .A(n21465), .B(n21679), .Z(n21671) );
  XNOR U21775 ( .A(n21464), .B(n21462), .Z(n21679) );
  AND U21776 ( .A(n21680), .B(n21681), .Z(n21462) );
  NANDN U21777 ( .A(n21682), .B(n21683), .Z(n21681) );
  OR U21778 ( .A(n21684), .B(n21685), .Z(n21683) );
  NAND U21779 ( .A(n21685), .B(n21684), .Z(n21680) );
  ANDN U21780 ( .B(B[204]), .A(n55), .Z(n21464) );
  XNOR U21781 ( .A(n21472), .B(n21686), .Z(n21465) );
  XNOR U21782 ( .A(n21471), .B(n21469), .Z(n21686) );
  AND U21783 ( .A(n21687), .B(n21688), .Z(n21469) );
  NANDN U21784 ( .A(n21689), .B(n21690), .Z(n21688) );
  NANDN U21785 ( .A(n21691), .B(n21692), .Z(n21690) );
  NANDN U21786 ( .A(n21692), .B(n21691), .Z(n21687) );
  ANDN U21787 ( .B(B[205]), .A(n56), .Z(n21471) );
  XNOR U21788 ( .A(n21479), .B(n21693), .Z(n21472) );
  XNOR U21789 ( .A(n21478), .B(n21476), .Z(n21693) );
  AND U21790 ( .A(n21694), .B(n21695), .Z(n21476) );
  NANDN U21791 ( .A(n21696), .B(n21697), .Z(n21695) );
  OR U21792 ( .A(n21698), .B(n21699), .Z(n21697) );
  NAND U21793 ( .A(n21699), .B(n21698), .Z(n21694) );
  ANDN U21794 ( .B(B[206]), .A(n57), .Z(n21478) );
  XNOR U21795 ( .A(n21486), .B(n21700), .Z(n21479) );
  XNOR U21796 ( .A(n21485), .B(n21483), .Z(n21700) );
  AND U21797 ( .A(n21701), .B(n21702), .Z(n21483) );
  NANDN U21798 ( .A(n21703), .B(n21704), .Z(n21702) );
  NANDN U21799 ( .A(n21705), .B(n21706), .Z(n21704) );
  NANDN U21800 ( .A(n21706), .B(n21705), .Z(n21701) );
  ANDN U21801 ( .B(B[207]), .A(n58), .Z(n21485) );
  XNOR U21802 ( .A(n21493), .B(n21707), .Z(n21486) );
  XNOR U21803 ( .A(n21492), .B(n21490), .Z(n21707) );
  AND U21804 ( .A(n21708), .B(n21709), .Z(n21490) );
  NANDN U21805 ( .A(n21710), .B(n21711), .Z(n21709) );
  OR U21806 ( .A(n21712), .B(n21713), .Z(n21711) );
  NAND U21807 ( .A(n21713), .B(n21712), .Z(n21708) );
  ANDN U21808 ( .B(B[208]), .A(n59), .Z(n21492) );
  XNOR U21809 ( .A(n21500), .B(n21714), .Z(n21493) );
  XNOR U21810 ( .A(n21499), .B(n21497), .Z(n21714) );
  AND U21811 ( .A(n21715), .B(n21716), .Z(n21497) );
  NANDN U21812 ( .A(n21717), .B(n21718), .Z(n21716) );
  NANDN U21813 ( .A(n21719), .B(n21720), .Z(n21718) );
  NANDN U21814 ( .A(n21720), .B(n21719), .Z(n21715) );
  ANDN U21815 ( .B(B[209]), .A(n60), .Z(n21499) );
  XNOR U21816 ( .A(n21507), .B(n21721), .Z(n21500) );
  XNOR U21817 ( .A(n21506), .B(n21504), .Z(n21721) );
  AND U21818 ( .A(n21722), .B(n21723), .Z(n21504) );
  NANDN U21819 ( .A(n21724), .B(n21725), .Z(n21723) );
  OR U21820 ( .A(n21726), .B(n21727), .Z(n21725) );
  NAND U21821 ( .A(n21727), .B(n21726), .Z(n21722) );
  ANDN U21822 ( .B(B[210]), .A(n61), .Z(n21506) );
  XNOR U21823 ( .A(n21514), .B(n21728), .Z(n21507) );
  XNOR U21824 ( .A(n21513), .B(n21511), .Z(n21728) );
  AND U21825 ( .A(n21729), .B(n21730), .Z(n21511) );
  NANDN U21826 ( .A(n21731), .B(n21732), .Z(n21730) );
  NANDN U21827 ( .A(n21733), .B(n21734), .Z(n21732) );
  NANDN U21828 ( .A(n21734), .B(n21733), .Z(n21729) );
  ANDN U21829 ( .B(B[211]), .A(n62), .Z(n21513) );
  XNOR U21830 ( .A(n21521), .B(n21735), .Z(n21514) );
  XNOR U21831 ( .A(n21520), .B(n21518), .Z(n21735) );
  AND U21832 ( .A(n21736), .B(n21737), .Z(n21518) );
  NANDN U21833 ( .A(n21738), .B(n21739), .Z(n21737) );
  OR U21834 ( .A(n21740), .B(n21741), .Z(n21739) );
  NAND U21835 ( .A(n21741), .B(n21740), .Z(n21736) );
  ANDN U21836 ( .B(B[212]), .A(n63), .Z(n21520) );
  XNOR U21837 ( .A(n21528), .B(n21742), .Z(n21521) );
  XNOR U21838 ( .A(n21527), .B(n21525), .Z(n21742) );
  AND U21839 ( .A(n21743), .B(n21744), .Z(n21525) );
  NANDN U21840 ( .A(n21745), .B(n21746), .Z(n21744) );
  NANDN U21841 ( .A(n21747), .B(n21748), .Z(n21746) );
  NANDN U21842 ( .A(n21748), .B(n21747), .Z(n21743) );
  ANDN U21843 ( .B(B[213]), .A(n64), .Z(n21527) );
  XNOR U21844 ( .A(n21535), .B(n21749), .Z(n21528) );
  XNOR U21845 ( .A(n21534), .B(n21532), .Z(n21749) );
  AND U21846 ( .A(n21750), .B(n21751), .Z(n21532) );
  NANDN U21847 ( .A(n21752), .B(n21753), .Z(n21751) );
  OR U21848 ( .A(n21754), .B(n21755), .Z(n21753) );
  NAND U21849 ( .A(n21755), .B(n21754), .Z(n21750) );
  ANDN U21850 ( .B(B[214]), .A(n65), .Z(n21534) );
  XNOR U21851 ( .A(n21542), .B(n21756), .Z(n21535) );
  XNOR U21852 ( .A(n21541), .B(n21539), .Z(n21756) );
  AND U21853 ( .A(n21757), .B(n21758), .Z(n21539) );
  NANDN U21854 ( .A(n21759), .B(n21760), .Z(n21758) );
  NANDN U21855 ( .A(n21761), .B(n21762), .Z(n21760) );
  NANDN U21856 ( .A(n21762), .B(n21761), .Z(n21757) );
  ANDN U21857 ( .B(B[215]), .A(n66), .Z(n21541) );
  XNOR U21858 ( .A(n21549), .B(n21763), .Z(n21542) );
  XNOR U21859 ( .A(n21548), .B(n21546), .Z(n21763) );
  AND U21860 ( .A(n21764), .B(n21765), .Z(n21546) );
  NANDN U21861 ( .A(n21766), .B(n21767), .Z(n21765) );
  OR U21862 ( .A(n21768), .B(n21769), .Z(n21767) );
  NAND U21863 ( .A(n21769), .B(n21768), .Z(n21764) );
  ANDN U21864 ( .B(B[216]), .A(n67), .Z(n21548) );
  XNOR U21865 ( .A(n21556), .B(n21770), .Z(n21549) );
  XNOR U21866 ( .A(n21555), .B(n21553), .Z(n21770) );
  AND U21867 ( .A(n21771), .B(n21772), .Z(n21553) );
  NANDN U21868 ( .A(n21773), .B(n21774), .Z(n21772) );
  NANDN U21869 ( .A(n21775), .B(n21776), .Z(n21774) );
  NANDN U21870 ( .A(n21776), .B(n21775), .Z(n21771) );
  ANDN U21871 ( .B(B[217]), .A(n68), .Z(n21555) );
  XNOR U21872 ( .A(n21563), .B(n21777), .Z(n21556) );
  XNOR U21873 ( .A(n21562), .B(n21560), .Z(n21777) );
  AND U21874 ( .A(n21778), .B(n21779), .Z(n21560) );
  NANDN U21875 ( .A(n21780), .B(n21781), .Z(n21779) );
  OR U21876 ( .A(n21782), .B(n21783), .Z(n21781) );
  NAND U21877 ( .A(n21783), .B(n21782), .Z(n21778) );
  ANDN U21878 ( .B(B[218]), .A(n69), .Z(n21562) );
  XNOR U21879 ( .A(n21570), .B(n21784), .Z(n21563) );
  XNOR U21880 ( .A(n21569), .B(n21567), .Z(n21784) );
  AND U21881 ( .A(n21785), .B(n21786), .Z(n21567) );
  NANDN U21882 ( .A(n21787), .B(n21788), .Z(n21786) );
  NANDN U21883 ( .A(n21789), .B(n21790), .Z(n21788) );
  NANDN U21884 ( .A(n21790), .B(n21789), .Z(n21785) );
  ANDN U21885 ( .B(B[219]), .A(n70), .Z(n21569) );
  XNOR U21886 ( .A(n21577), .B(n21791), .Z(n21570) );
  XNOR U21887 ( .A(n21576), .B(n21574), .Z(n21791) );
  AND U21888 ( .A(n21792), .B(n21793), .Z(n21574) );
  NANDN U21889 ( .A(n21794), .B(n21795), .Z(n21793) );
  OR U21890 ( .A(n21796), .B(n21797), .Z(n21795) );
  NAND U21891 ( .A(n21797), .B(n21796), .Z(n21792) );
  ANDN U21892 ( .B(B[220]), .A(n71), .Z(n21576) );
  XNOR U21893 ( .A(n21584), .B(n21798), .Z(n21577) );
  XNOR U21894 ( .A(n21583), .B(n21581), .Z(n21798) );
  AND U21895 ( .A(n21799), .B(n21800), .Z(n21581) );
  NANDN U21896 ( .A(n21801), .B(n21802), .Z(n21800) );
  NANDN U21897 ( .A(n21803), .B(n21804), .Z(n21802) );
  NANDN U21898 ( .A(n21804), .B(n21803), .Z(n21799) );
  ANDN U21899 ( .B(B[221]), .A(n72), .Z(n21583) );
  XNOR U21900 ( .A(n21591), .B(n21805), .Z(n21584) );
  XNOR U21901 ( .A(n21590), .B(n21588), .Z(n21805) );
  AND U21902 ( .A(n21806), .B(n21807), .Z(n21588) );
  NANDN U21903 ( .A(n21808), .B(n21809), .Z(n21807) );
  OR U21904 ( .A(n21810), .B(n21811), .Z(n21809) );
  NAND U21905 ( .A(n21811), .B(n21810), .Z(n21806) );
  ANDN U21906 ( .B(B[222]), .A(n73), .Z(n21590) );
  XNOR U21907 ( .A(n21598), .B(n21812), .Z(n21591) );
  XNOR U21908 ( .A(n21597), .B(n21595), .Z(n21812) );
  AND U21909 ( .A(n21813), .B(n21814), .Z(n21595) );
  NANDN U21910 ( .A(n21815), .B(n21816), .Z(n21814) );
  NANDN U21911 ( .A(n21817), .B(n21818), .Z(n21816) );
  NANDN U21912 ( .A(n21818), .B(n21817), .Z(n21813) );
  ANDN U21913 ( .B(B[223]), .A(n74), .Z(n21597) );
  XNOR U21914 ( .A(n21605), .B(n21819), .Z(n21598) );
  XNOR U21915 ( .A(n21604), .B(n21602), .Z(n21819) );
  AND U21916 ( .A(n21820), .B(n21821), .Z(n21602) );
  NANDN U21917 ( .A(n21822), .B(n21823), .Z(n21821) );
  OR U21918 ( .A(n21824), .B(n21825), .Z(n21823) );
  NAND U21919 ( .A(n21825), .B(n21824), .Z(n21820) );
  ANDN U21920 ( .B(B[224]), .A(n75), .Z(n21604) );
  XNOR U21921 ( .A(n21612), .B(n21826), .Z(n21605) );
  XNOR U21922 ( .A(n21611), .B(n21609), .Z(n21826) );
  AND U21923 ( .A(n21827), .B(n21828), .Z(n21609) );
  NANDN U21924 ( .A(n21829), .B(n21830), .Z(n21828) );
  NANDN U21925 ( .A(n21831), .B(n21832), .Z(n21830) );
  NANDN U21926 ( .A(n21832), .B(n21831), .Z(n21827) );
  ANDN U21927 ( .B(B[225]), .A(n76), .Z(n21611) );
  XNOR U21928 ( .A(n21619), .B(n21833), .Z(n21612) );
  XNOR U21929 ( .A(n21618), .B(n21616), .Z(n21833) );
  AND U21930 ( .A(n21834), .B(n21835), .Z(n21616) );
  NANDN U21931 ( .A(n21836), .B(n21837), .Z(n21835) );
  OR U21932 ( .A(n21838), .B(n21839), .Z(n21837) );
  NAND U21933 ( .A(n21839), .B(n21838), .Z(n21834) );
  ANDN U21934 ( .B(B[226]), .A(n77), .Z(n21618) );
  XNOR U21935 ( .A(n21626), .B(n21840), .Z(n21619) );
  XNOR U21936 ( .A(n21625), .B(n21623), .Z(n21840) );
  AND U21937 ( .A(n21841), .B(n21842), .Z(n21623) );
  NANDN U21938 ( .A(n21843), .B(n21844), .Z(n21842) );
  NANDN U21939 ( .A(n21845), .B(n21846), .Z(n21844) );
  NANDN U21940 ( .A(n21846), .B(n21845), .Z(n21841) );
  ANDN U21941 ( .B(B[227]), .A(n78), .Z(n21625) );
  XNOR U21942 ( .A(n21633), .B(n21847), .Z(n21626) );
  XNOR U21943 ( .A(n21632), .B(n21630), .Z(n21847) );
  AND U21944 ( .A(n21848), .B(n21849), .Z(n21630) );
  NANDN U21945 ( .A(n21850), .B(n21851), .Z(n21849) );
  OR U21946 ( .A(n21852), .B(n21853), .Z(n21851) );
  NAND U21947 ( .A(n21853), .B(n21852), .Z(n21848) );
  ANDN U21948 ( .B(B[228]), .A(n79), .Z(n21632) );
  XNOR U21949 ( .A(n21640), .B(n21854), .Z(n21633) );
  XNOR U21950 ( .A(n21639), .B(n21637), .Z(n21854) );
  AND U21951 ( .A(n21855), .B(n21856), .Z(n21637) );
  NANDN U21952 ( .A(n21857), .B(n21858), .Z(n21856) );
  NANDN U21953 ( .A(n21859), .B(n21860), .Z(n21858) );
  NANDN U21954 ( .A(n21860), .B(n21859), .Z(n21855) );
  ANDN U21955 ( .B(B[229]), .A(n80), .Z(n21639) );
  XNOR U21956 ( .A(n21647), .B(n21861), .Z(n21640) );
  XNOR U21957 ( .A(n21646), .B(n21644), .Z(n21861) );
  AND U21958 ( .A(n21862), .B(n21863), .Z(n21644) );
  NANDN U21959 ( .A(n21864), .B(n21865), .Z(n21863) );
  OR U21960 ( .A(n21866), .B(n21867), .Z(n21865) );
  NAND U21961 ( .A(n21867), .B(n21866), .Z(n21862) );
  ANDN U21962 ( .B(B[230]), .A(n81), .Z(n21646) );
  XNOR U21963 ( .A(n21654), .B(n21868), .Z(n21647) );
  XNOR U21964 ( .A(n21653), .B(n21651), .Z(n21868) );
  AND U21965 ( .A(n21869), .B(n21870), .Z(n21651) );
  NANDN U21966 ( .A(n21871), .B(n21872), .Z(n21870) );
  NAND U21967 ( .A(n21873), .B(n21874), .Z(n21872) );
  ANDN U21968 ( .B(B[231]), .A(n82), .Z(n21653) );
  XOR U21969 ( .A(n21660), .B(n21875), .Z(n21654) );
  XNOR U21970 ( .A(n21658), .B(n21661), .Z(n21875) );
  NAND U21971 ( .A(A[2]), .B(B[232]), .Z(n21661) );
  NANDN U21972 ( .A(n21876), .B(n21877), .Z(n21658) );
  AND U21973 ( .A(A[0]), .B(B[233]), .Z(n21877) );
  XNOR U21974 ( .A(n21663), .B(n21878), .Z(n21660) );
  NAND U21975 ( .A(A[0]), .B(B[234]), .Z(n21878) );
  NAND U21976 ( .A(B[233]), .B(A[1]), .Z(n21663) );
  NAND U21977 ( .A(n21879), .B(n21880), .Z(n328) );
  NANDN U21978 ( .A(n21881), .B(n21882), .Z(n21880) );
  OR U21979 ( .A(n21883), .B(n21884), .Z(n21882) );
  NAND U21980 ( .A(n21884), .B(n21883), .Z(n21879) );
  XOR U21981 ( .A(n330), .B(n329), .Z(\A1[231] ) );
  XOR U21982 ( .A(n21884), .B(n21885), .Z(n329) );
  XNOR U21983 ( .A(n21883), .B(n21881), .Z(n21885) );
  AND U21984 ( .A(n21886), .B(n21887), .Z(n21881) );
  NANDN U21985 ( .A(n21888), .B(n21889), .Z(n21887) );
  NANDN U21986 ( .A(n21890), .B(n21891), .Z(n21889) );
  NANDN U21987 ( .A(n21891), .B(n21890), .Z(n21886) );
  ANDN U21988 ( .B(B[202]), .A(n54), .Z(n21883) );
  XNOR U21989 ( .A(n21678), .B(n21892), .Z(n21884) );
  XNOR U21990 ( .A(n21677), .B(n21675), .Z(n21892) );
  AND U21991 ( .A(n21893), .B(n21894), .Z(n21675) );
  NANDN U21992 ( .A(n21895), .B(n21896), .Z(n21894) );
  OR U21993 ( .A(n21897), .B(n21898), .Z(n21896) );
  NAND U21994 ( .A(n21898), .B(n21897), .Z(n21893) );
  ANDN U21995 ( .B(B[203]), .A(n55), .Z(n21677) );
  XNOR U21996 ( .A(n21685), .B(n21899), .Z(n21678) );
  XNOR U21997 ( .A(n21684), .B(n21682), .Z(n21899) );
  AND U21998 ( .A(n21900), .B(n21901), .Z(n21682) );
  NANDN U21999 ( .A(n21902), .B(n21903), .Z(n21901) );
  NANDN U22000 ( .A(n21904), .B(n21905), .Z(n21903) );
  NANDN U22001 ( .A(n21905), .B(n21904), .Z(n21900) );
  ANDN U22002 ( .B(B[204]), .A(n56), .Z(n21684) );
  XNOR U22003 ( .A(n21692), .B(n21906), .Z(n21685) );
  XNOR U22004 ( .A(n21691), .B(n21689), .Z(n21906) );
  AND U22005 ( .A(n21907), .B(n21908), .Z(n21689) );
  NANDN U22006 ( .A(n21909), .B(n21910), .Z(n21908) );
  OR U22007 ( .A(n21911), .B(n21912), .Z(n21910) );
  NAND U22008 ( .A(n21912), .B(n21911), .Z(n21907) );
  ANDN U22009 ( .B(B[205]), .A(n57), .Z(n21691) );
  XNOR U22010 ( .A(n21699), .B(n21913), .Z(n21692) );
  XNOR U22011 ( .A(n21698), .B(n21696), .Z(n21913) );
  AND U22012 ( .A(n21914), .B(n21915), .Z(n21696) );
  NANDN U22013 ( .A(n21916), .B(n21917), .Z(n21915) );
  NANDN U22014 ( .A(n21918), .B(n21919), .Z(n21917) );
  NANDN U22015 ( .A(n21919), .B(n21918), .Z(n21914) );
  ANDN U22016 ( .B(B[206]), .A(n58), .Z(n21698) );
  XNOR U22017 ( .A(n21706), .B(n21920), .Z(n21699) );
  XNOR U22018 ( .A(n21705), .B(n21703), .Z(n21920) );
  AND U22019 ( .A(n21921), .B(n21922), .Z(n21703) );
  NANDN U22020 ( .A(n21923), .B(n21924), .Z(n21922) );
  OR U22021 ( .A(n21925), .B(n21926), .Z(n21924) );
  NAND U22022 ( .A(n21926), .B(n21925), .Z(n21921) );
  ANDN U22023 ( .B(B[207]), .A(n59), .Z(n21705) );
  XNOR U22024 ( .A(n21713), .B(n21927), .Z(n21706) );
  XNOR U22025 ( .A(n21712), .B(n21710), .Z(n21927) );
  AND U22026 ( .A(n21928), .B(n21929), .Z(n21710) );
  NANDN U22027 ( .A(n21930), .B(n21931), .Z(n21929) );
  NANDN U22028 ( .A(n21932), .B(n21933), .Z(n21931) );
  NANDN U22029 ( .A(n21933), .B(n21932), .Z(n21928) );
  ANDN U22030 ( .B(B[208]), .A(n60), .Z(n21712) );
  XNOR U22031 ( .A(n21720), .B(n21934), .Z(n21713) );
  XNOR U22032 ( .A(n21719), .B(n21717), .Z(n21934) );
  AND U22033 ( .A(n21935), .B(n21936), .Z(n21717) );
  NANDN U22034 ( .A(n21937), .B(n21938), .Z(n21936) );
  OR U22035 ( .A(n21939), .B(n21940), .Z(n21938) );
  NAND U22036 ( .A(n21940), .B(n21939), .Z(n21935) );
  ANDN U22037 ( .B(B[209]), .A(n61), .Z(n21719) );
  XNOR U22038 ( .A(n21727), .B(n21941), .Z(n21720) );
  XNOR U22039 ( .A(n21726), .B(n21724), .Z(n21941) );
  AND U22040 ( .A(n21942), .B(n21943), .Z(n21724) );
  NANDN U22041 ( .A(n21944), .B(n21945), .Z(n21943) );
  NANDN U22042 ( .A(n21946), .B(n21947), .Z(n21945) );
  NANDN U22043 ( .A(n21947), .B(n21946), .Z(n21942) );
  ANDN U22044 ( .B(B[210]), .A(n62), .Z(n21726) );
  XNOR U22045 ( .A(n21734), .B(n21948), .Z(n21727) );
  XNOR U22046 ( .A(n21733), .B(n21731), .Z(n21948) );
  AND U22047 ( .A(n21949), .B(n21950), .Z(n21731) );
  NANDN U22048 ( .A(n21951), .B(n21952), .Z(n21950) );
  OR U22049 ( .A(n21953), .B(n21954), .Z(n21952) );
  NAND U22050 ( .A(n21954), .B(n21953), .Z(n21949) );
  ANDN U22051 ( .B(B[211]), .A(n63), .Z(n21733) );
  XNOR U22052 ( .A(n21741), .B(n21955), .Z(n21734) );
  XNOR U22053 ( .A(n21740), .B(n21738), .Z(n21955) );
  AND U22054 ( .A(n21956), .B(n21957), .Z(n21738) );
  NANDN U22055 ( .A(n21958), .B(n21959), .Z(n21957) );
  NANDN U22056 ( .A(n21960), .B(n21961), .Z(n21959) );
  NANDN U22057 ( .A(n21961), .B(n21960), .Z(n21956) );
  ANDN U22058 ( .B(B[212]), .A(n64), .Z(n21740) );
  XNOR U22059 ( .A(n21748), .B(n21962), .Z(n21741) );
  XNOR U22060 ( .A(n21747), .B(n21745), .Z(n21962) );
  AND U22061 ( .A(n21963), .B(n21964), .Z(n21745) );
  NANDN U22062 ( .A(n21965), .B(n21966), .Z(n21964) );
  OR U22063 ( .A(n21967), .B(n21968), .Z(n21966) );
  NAND U22064 ( .A(n21968), .B(n21967), .Z(n21963) );
  ANDN U22065 ( .B(B[213]), .A(n65), .Z(n21747) );
  XNOR U22066 ( .A(n21755), .B(n21969), .Z(n21748) );
  XNOR U22067 ( .A(n21754), .B(n21752), .Z(n21969) );
  AND U22068 ( .A(n21970), .B(n21971), .Z(n21752) );
  NANDN U22069 ( .A(n21972), .B(n21973), .Z(n21971) );
  NANDN U22070 ( .A(n21974), .B(n21975), .Z(n21973) );
  NANDN U22071 ( .A(n21975), .B(n21974), .Z(n21970) );
  ANDN U22072 ( .B(B[214]), .A(n66), .Z(n21754) );
  XNOR U22073 ( .A(n21762), .B(n21976), .Z(n21755) );
  XNOR U22074 ( .A(n21761), .B(n21759), .Z(n21976) );
  AND U22075 ( .A(n21977), .B(n21978), .Z(n21759) );
  NANDN U22076 ( .A(n21979), .B(n21980), .Z(n21978) );
  OR U22077 ( .A(n21981), .B(n21982), .Z(n21980) );
  NAND U22078 ( .A(n21982), .B(n21981), .Z(n21977) );
  ANDN U22079 ( .B(B[215]), .A(n67), .Z(n21761) );
  XNOR U22080 ( .A(n21769), .B(n21983), .Z(n21762) );
  XNOR U22081 ( .A(n21768), .B(n21766), .Z(n21983) );
  AND U22082 ( .A(n21984), .B(n21985), .Z(n21766) );
  NANDN U22083 ( .A(n21986), .B(n21987), .Z(n21985) );
  NANDN U22084 ( .A(n21988), .B(n21989), .Z(n21987) );
  NANDN U22085 ( .A(n21989), .B(n21988), .Z(n21984) );
  ANDN U22086 ( .B(B[216]), .A(n68), .Z(n21768) );
  XNOR U22087 ( .A(n21776), .B(n21990), .Z(n21769) );
  XNOR U22088 ( .A(n21775), .B(n21773), .Z(n21990) );
  AND U22089 ( .A(n21991), .B(n21992), .Z(n21773) );
  NANDN U22090 ( .A(n21993), .B(n21994), .Z(n21992) );
  OR U22091 ( .A(n21995), .B(n21996), .Z(n21994) );
  NAND U22092 ( .A(n21996), .B(n21995), .Z(n21991) );
  ANDN U22093 ( .B(B[217]), .A(n69), .Z(n21775) );
  XNOR U22094 ( .A(n21783), .B(n21997), .Z(n21776) );
  XNOR U22095 ( .A(n21782), .B(n21780), .Z(n21997) );
  AND U22096 ( .A(n21998), .B(n21999), .Z(n21780) );
  NANDN U22097 ( .A(n22000), .B(n22001), .Z(n21999) );
  NANDN U22098 ( .A(n22002), .B(n22003), .Z(n22001) );
  NANDN U22099 ( .A(n22003), .B(n22002), .Z(n21998) );
  ANDN U22100 ( .B(B[218]), .A(n70), .Z(n21782) );
  XNOR U22101 ( .A(n21790), .B(n22004), .Z(n21783) );
  XNOR U22102 ( .A(n21789), .B(n21787), .Z(n22004) );
  AND U22103 ( .A(n22005), .B(n22006), .Z(n21787) );
  NANDN U22104 ( .A(n22007), .B(n22008), .Z(n22006) );
  OR U22105 ( .A(n22009), .B(n22010), .Z(n22008) );
  NAND U22106 ( .A(n22010), .B(n22009), .Z(n22005) );
  ANDN U22107 ( .B(B[219]), .A(n71), .Z(n21789) );
  XNOR U22108 ( .A(n21797), .B(n22011), .Z(n21790) );
  XNOR U22109 ( .A(n21796), .B(n21794), .Z(n22011) );
  AND U22110 ( .A(n22012), .B(n22013), .Z(n21794) );
  NANDN U22111 ( .A(n22014), .B(n22015), .Z(n22013) );
  NANDN U22112 ( .A(n22016), .B(n22017), .Z(n22015) );
  NANDN U22113 ( .A(n22017), .B(n22016), .Z(n22012) );
  ANDN U22114 ( .B(B[220]), .A(n72), .Z(n21796) );
  XNOR U22115 ( .A(n21804), .B(n22018), .Z(n21797) );
  XNOR U22116 ( .A(n21803), .B(n21801), .Z(n22018) );
  AND U22117 ( .A(n22019), .B(n22020), .Z(n21801) );
  NANDN U22118 ( .A(n22021), .B(n22022), .Z(n22020) );
  OR U22119 ( .A(n22023), .B(n22024), .Z(n22022) );
  NAND U22120 ( .A(n22024), .B(n22023), .Z(n22019) );
  ANDN U22121 ( .B(B[221]), .A(n73), .Z(n21803) );
  XNOR U22122 ( .A(n21811), .B(n22025), .Z(n21804) );
  XNOR U22123 ( .A(n21810), .B(n21808), .Z(n22025) );
  AND U22124 ( .A(n22026), .B(n22027), .Z(n21808) );
  NANDN U22125 ( .A(n22028), .B(n22029), .Z(n22027) );
  NANDN U22126 ( .A(n22030), .B(n22031), .Z(n22029) );
  NANDN U22127 ( .A(n22031), .B(n22030), .Z(n22026) );
  ANDN U22128 ( .B(B[222]), .A(n74), .Z(n21810) );
  XNOR U22129 ( .A(n21818), .B(n22032), .Z(n21811) );
  XNOR U22130 ( .A(n21817), .B(n21815), .Z(n22032) );
  AND U22131 ( .A(n22033), .B(n22034), .Z(n21815) );
  NANDN U22132 ( .A(n22035), .B(n22036), .Z(n22034) );
  OR U22133 ( .A(n22037), .B(n22038), .Z(n22036) );
  NAND U22134 ( .A(n22038), .B(n22037), .Z(n22033) );
  ANDN U22135 ( .B(B[223]), .A(n75), .Z(n21817) );
  XNOR U22136 ( .A(n21825), .B(n22039), .Z(n21818) );
  XNOR U22137 ( .A(n21824), .B(n21822), .Z(n22039) );
  AND U22138 ( .A(n22040), .B(n22041), .Z(n21822) );
  NANDN U22139 ( .A(n22042), .B(n22043), .Z(n22041) );
  NANDN U22140 ( .A(n22044), .B(n22045), .Z(n22043) );
  NANDN U22141 ( .A(n22045), .B(n22044), .Z(n22040) );
  ANDN U22142 ( .B(B[224]), .A(n76), .Z(n21824) );
  XNOR U22143 ( .A(n21832), .B(n22046), .Z(n21825) );
  XNOR U22144 ( .A(n21831), .B(n21829), .Z(n22046) );
  AND U22145 ( .A(n22047), .B(n22048), .Z(n21829) );
  NANDN U22146 ( .A(n22049), .B(n22050), .Z(n22048) );
  OR U22147 ( .A(n22051), .B(n22052), .Z(n22050) );
  NAND U22148 ( .A(n22052), .B(n22051), .Z(n22047) );
  ANDN U22149 ( .B(B[225]), .A(n77), .Z(n21831) );
  XNOR U22150 ( .A(n21839), .B(n22053), .Z(n21832) );
  XNOR U22151 ( .A(n21838), .B(n21836), .Z(n22053) );
  AND U22152 ( .A(n22054), .B(n22055), .Z(n21836) );
  NANDN U22153 ( .A(n22056), .B(n22057), .Z(n22055) );
  NANDN U22154 ( .A(n22058), .B(n22059), .Z(n22057) );
  NANDN U22155 ( .A(n22059), .B(n22058), .Z(n22054) );
  ANDN U22156 ( .B(B[226]), .A(n78), .Z(n21838) );
  XNOR U22157 ( .A(n21846), .B(n22060), .Z(n21839) );
  XNOR U22158 ( .A(n21845), .B(n21843), .Z(n22060) );
  AND U22159 ( .A(n22061), .B(n22062), .Z(n21843) );
  NANDN U22160 ( .A(n22063), .B(n22064), .Z(n22062) );
  OR U22161 ( .A(n22065), .B(n22066), .Z(n22064) );
  NAND U22162 ( .A(n22066), .B(n22065), .Z(n22061) );
  ANDN U22163 ( .B(B[227]), .A(n79), .Z(n21845) );
  XNOR U22164 ( .A(n21853), .B(n22067), .Z(n21846) );
  XNOR U22165 ( .A(n21852), .B(n21850), .Z(n22067) );
  AND U22166 ( .A(n22068), .B(n22069), .Z(n21850) );
  NANDN U22167 ( .A(n22070), .B(n22071), .Z(n22069) );
  NANDN U22168 ( .A(n22072), .B(n22073), .Z(n22071) );
  NANDN U22169 ( .A(n22073), .B(n22072), .Z(n22068) );
  ANDN U22170 ( .B(B[228]), .A(n80), .Z(n21852) );
  XNOR U22171 ( .A(n21860), .B(n22074), .Z(n21853) );
  XNOR U22172 ( .A(n21859), .B(n21857), .Z(n22074) );
  AND U22173 ( .A(n22075), .B(n22076), .Z(n21857) );
  NANDN U22174 ( .A(n22077), .B(n22078), .Z(n22076) );
  OR U22175 ( .A(n22079), .B(n22080), .Z(n22078) );
  NAND U22176 ( .A(n22080), .B(n22079), .Z(n22075) );
  ANDN U22177 ( .B(B[229]), .A(n81), .Z(n21859) );
  XNOR U22178 ( .A(n21867), .B(n22081), .Z(n21860) );
  XNOR U22179 ( .A(n21866), .B(n21864), .Z(n22081) );
  AND U22180 ( .A(n22082), .B(n22083), .Z(n21864) );
  NANDN U22181 ( .A(n22084), .B(n22085), .Z(n22083) );
  NAND U22182 ( .A(n22086), .B(n22087), .Z(n22085) );
  ANDN U22183 ( .B(B[230]), .A(n82), .Z(n21866) );
  XOR U22184 ( .A(n21873), .B(n22088), .Z(n21867) );
  XNOR U22185 ( .A(n21871), .B(n21874), .Z(n22088) );
  NAND U22186 ( .A(A[2]), .B(B[231]), .Z(n21874) );
  NANDN U22187 ( .A(n22089), .B(n22090), .Z(n21871) );
  AND U22188 ( .A(A[0]), .B(B[232]), .Z(n22090) );
  XNOR U22189 ( .A(n21876), .B(n22091), .Z(n21873) );
  NAND U22190 ( .A(A[0]), .B(B[233]), .Z(n22091) );
  NAND U22191 ( .A(B[232]), .B(A[1]), .Z(n21876) );
  NAND U22192 ( .A(n22092), .B(n22093), .Z(n330) );
  NANDN U22193 ( .A(n22094), .B(n22095), .Z(n22093) );
  OR U22194 ( .A(n22096), .B(n22097), .Z(n22095) );
  NAND U22195 ( .A(n22097), .B(n22096), .Z(n22092) );
  XOR U22196 ( .A(n332), .B(n331), .Z(\A1[230] ) );
  XOR U22197 ( .A(n22097), .B(n22098), .Z(n331) );
  XNOR U22198 ( .A(n22096), .B(n22094), .Z(n22098) );
  AND U22199 ( .A(n22099), .B(n22100), .Z(n22094) );
  NANDN U22200 ( .A(n22101), .B(n22102), .Z(n22100) );
  NANDN U22201 ( .A(n22103), .B(n22104), .Z(n22102) );
  NANDN U22202 ( .A(n22104), .B(n22103), .Z(n22099) );
  ANDN U22203 ( .B(B[201]), .A(n54), .Z(n22096) );
  XNOR U22204 ( .A(n21891), .B(n22105), .Z(n22097) );
  XNOR U22205 ( .A(n21890), .B(n21888), .Z(n22105) );
  AND U22206 ( .A(n22106), .B(n22107), .Z(n21888) );
  NANDN U22207 ( .A(n22108), .B(n22109), .Z(n22107) );
  OR U22208 ( .A(n22110), .B(n22111), .Z(n22109) );
  NAND U22209 ( .A(n22111), .B(n22110), .Z(n22106) );
  ANDN U22210 ( .B(B[202]), .A(n55), .Z(n21890) );
  XNOR U22211 ( .A(n21898), .B(n22112), .Z(n21891) );
  XNOR U22212 ( .A(n21897), .B(n21895), .Z(n22112) );
  AND U22213 ( .A(n22113), .B(n22114), .Z(n21895) );
  NANDN U22214 ( .A(n22115), .B(n22116), .Z(n22114) );
  NANDN U22215 ( .A(n22117), .B(n22118), .Z(n22116) );
  NANDN U22216 ( .A(n22118), .B(n22117), .Z(n22113) );
  ANDN U22217 ( .B(B[203]), .A(n56), .Z(n21897) );
  XNOR U22218 ( .A(n21905), .B(n22119), .Z(n21898) );
  XNOR U22219 ( .A(n21904), .B(n21902), .Z(n22119) );
  AND U22220 ( .A(n22120), .B(n22121), .Z(n21902) );
  NANDN U22221 ( .A(n22122), .B(n22123), .Z(n22121) );
  OR U22222 ( .A(n22124), .B(n22125), .Z(n22123) );
  NAND U22223 ( .A(n22125), .B(n22124), .Z(n22120) );
  ANDN U22224 ( .B(B[204]), .A(n57), .Z(n21904) );
  XNOR U22225 ( .A(n21912), .B(n22126), .Z(n21905) );
  XNOR U22226 ( .A(n21911), .B(n21909), .Z(n22126) );
  AND U22227 ( .A(n22127), .B(n22128), .Z(n21909) );
  NANDN U22228 ( .A(n22129), .B(n22130), .Z(n22128) );
  NANDN U22229 ( .A(n22131), .B(n22132), .Z(n22130) );
  NANDN U22230 ( .A(n22132), .B(n22131), .Z(n22127) );
  ANDN U22231 ( .B(B[205]), .A(n58), .Z(n21911) );
  XNOR U22232 ( .A(n21919), .B(n22133), .Z(n21912) );
  XNOR U22233 ( .A(n21918), .B(n21916), .Z(n22133) );
  AND U22234 ( .A(n22134), .B(n22135), .Z(n21916) );
  NANDN U22235 ( .A(n22136), .B(n22137), .Z(n22135) );
  OR U22236 ( .A(n22138), .B(n22139), .Z(n22137) );
  NAND U22237 ( .A(n22139), .B(n22138), .Z(n22134) );
  ANDN U22238 ( .B(B[206]), .A(n59), .Z(n21918) );
  XNOR U22239 ( .A(n21926), .B(n22140), .Z(n21919) );
  XNOR U22240 ( .A(n21925), .B(n21923), .Z(n22140) );
  AND U22241 ( .A(n22141), .B(n22142), .Z(n21923) );
  NANDN U22242 ( .A(n22143), .B(n22144), .Z(n22142) );
  NANDN U22243 ( .A(n22145), .B(n22146), .Z(n22144) );
  NANDN U22244 ( .A(n22146), .B(n22145), .Z(n22141) );
  ANDN U22245 ( .B(B[207]), .A(n60), .Z(n21925) );
  XNOR U22246 ( .A(n21933), .B(n22147), .Z(n21926) );
  XNOR U22247 ( .A(n21932), .B(n21930), .Z(n22147) );
  AND U22248 ( .A(n22148), .B(n22149), .Z(n21930) );
  NANDN U22249 ( .A(n22150), .B(n22151), .Z(n22149) );
  OR U22250 ( .A(n22152), .B(n22153), .Z(n22151) );
  NAND U22251 ( .A(n22153), .B(n22152), .Z(n22148) );
  ANDN U22252 ( .B(B[208]), .A(n61), .Z(n21932) );
  XNOR U22253 ( .A(n21940), .B(n22154), .Z(n21933) );
  XNOR U22254 ( .A(n21939), .B(n21937), .Z(n22154) );
  AND U22255 ( .A(n22155), .B(n22156), .Z(n21937) );
  NANDN U22256 ( .A(n22157), .B(n22158), .Z(n22156) );
  NANDN U22257 ( .A(n22159), .B(n22160), .Z(n22158) );
  NANDN U22258 ( .A(n22160), .B(n22159), .Z(n22155) );
  ANDN U22259 ( .B(B[209]), .A(n62), .Z(n21939) );
  XNOR U22260 ( .A(n21947), .B(n22161), .Z(n21940) );
  XNOR U22261 ( .A(n21946), .B(n21944), .Z(n22161) );
  AND U22262 ( .A(n22162), .B(n22163), .Z(n21944) );
  NANDN U22263 ( .A(n22164), .B(n22165), .Z(n22163) );
  OR U22264 ( .A(n22166), .B(n22167), .Z(n22165) );
  NAND U22265 ( .A(n22167), .B(n22166), .Z(n22162) );
  ANDN U22266 ( .B(B[210]), .A(n63), .Z(n21946) );
  XNOR U22267 ( .A(n21954), .B(n22168), .Z(n21947) );
  XNOR U22268 ( .A(n21953), .B(n21951), .Z(n22168) );
  AND U22269 ( .A(n22169), .B(n22170), .Z(n21951) );
  NANDN U22270 ( .A(n22171), .B(n22172), .Z(n22170) );
  NANDN U22271 ( .A(n22173), .B(n22174), .Z(n22172) );
  NANDN U22272 ( .A(n22174), .B(n22173), .Z(n22169) );
  ANDN U22273 ( .B(B[211]), .A(n64), .Z(n21953) );
  XNOR U22274 ( .A(n21961), .B(n22175), .Z(n21954) );
  XNOR U22275 ( .A(n21960), .B(n21958), .Z(n22175) );
  AND U22276 ( .A(n22176), .B(n22177), .Z(n21958) );
  NANDN U22277 ( .A(n22178), .B(n22179), .Z(n22177) );
  OR U22278 ( .A(n22180), .B(n22181), .Z(n22179) );
  NAND U22279 ( .A(n22181), .B(n22180), .Z(n22176) );
  ANDN U22280 ( .B(B[212]), .A(n65), .Z(n21960) );
  XNOR U22281 ( .A(n21968), .B(n22182), .Z(n21961) );
  XNOR U22282 ( .A(n21967), .B(n21965), .Z(n22182) );
  AND U22283 ( .A(n22183), .B(n22184), .Z(n21965) );
  NANDN U22284 ( .A(n22185), .B(n22186), .Z(n22184) );
  NANDN U22285 ( .A(n22187), .B(n22188), .Z(n22186) );
  NANDN U22286 ( .A(n22188), .B(n22187), .Z(n22183) );
  ANDN U22287 ( .B(B[213]), .A(n66), .Z(n21967) );
  XNOR U22288 ( .A(n21975), .B(n22189), .Z(n21968) );
  XNOR U22289 ( .A(n21974), .B(n21972), .Z(n22189) );
  AND U22290 ( .A(n22190), .B(n22191), .Z(n21972) );
  NANDN U22291 ( .A(n22192), .B(n22193), .Z(n22191) );
  OR U22292 ( .A(n22194), .B(n22195), .Z(n22193) );
  NAND U22293 ( .A(n22195), .B(n22194), .Z(n22190) );
  ANDN U22294 ( .B(B[214]), .A(n67), .Z(n21974) );
  XNOR U22295 ( .A(n21982), .B(n22196), .Z(n21975) );
  XNOR U22296 ( .A(n21981), .B(n21979), .Z(n22196) );
  AND U22297 ( .A(n22197), .B(n22198), .Z(n21979) );
  NANDN U22298 ( .A(n22199), .B(n22200), .Z(n22198) );
  NANDN U22299 ( .A(n22201), .B(n22202), .Z(n22200) );
  NANDN U22300 ( .A(n22202), .B(n22201), .Z(n22197) );
  ANDN U22301 ( .B(B[215]), .A(n68), .Z(n21981) );
  XNOR U22302 ( .A(n21989), .B(n22203), .Z(n21982) );
  XNOR U22303 ( .A(n21988), .B(n21986), .Z(n22203) );
  AND U22304 ( .A(n22204), .B(n22205), .Z(n21986) );
  NANDN U22305 ( .A(n22206), .B(n22207), .Z(n22205) );
  OR U22306 ( .A(n22208), .B(n22209), .Z(n22207) );
  NAND U22307 ( .A(n22209), .B(n22208), .Z(n22204) );
  ANDN U22308 ( .B(B[216]), .A(n69), .Z(n21988) );
  XNOR U22309 ( .A(n21996), .B(n22210), .Z(n21989) );
  XNOR U22310 ( .A(n21995), .B(n21993), .Z(n22210) );
  AND U22311 ( .A(n22211), .B(n22212), .Z(n21993) );
  NANDN U22312 ( .A(n22213), .B(n22214), .Z(n22212) );
  NANDN U22313 ( .A(n22215), .B(n22216), .Z(n22214) );
  NANDN U22314 ( .A(n22216), .B(n22215), .Z(n22211) );
  ANDN U22315 ( .B(B[217]), .A(n70), .Z(n21995) );
  XNOR U22316 ( .A(n22003), .B(n22217), .Z(n21996) );
  XNOR U22317 ( .A(n22002), .B(n22000), .Z(n22217) );
  AND U22318 ( .A(n22218), .B(n22219), .Z(n22000) );
  NANDN U22319 ( .A(n22220), .B(n22221), .Z(n22219) );
  OR U22320 ( .A(n22222), .B(n22223), .Z(n22221) );
  NAND U22321 ( .A(n22223), .B(n22222), .Z(n22218) );
  ANDN U22322 ( .B(B[218]), .A(n71), .Z(n22002) );
  XNOR U22323 ( .A(n22010), .B(n22224), .Z(n22003) );
  XNOR U22324 ( .A(n22009), .B(n22007), .Z(n22224) );
  AND U22325 ( .A(n22225), .B(n22226), .Z(n22007) );
  NANDN U22326 ( .A(n22227), .B(n22228), .Z(n22226) );
  NANDN U22327 ( .A(n22229), .B(n22230), .Z(n22228) );
  NANDN U22328 ( .A(n22230), .B(n22229), .Z(n22225) );
  ANDN U22329 ( .B(B[219]), .A(n72), .Z(n22009) );
  XNOR U22330 ( .A(n22017), .B(n22231), .Z(n22010) );
  XNOR U22331 ( .A(n22016), .B(n22014), .Z(n22231) );
  AND U22332 ( .A(n22232), .B(n22233), .Z(n22014) );
  NANDN U22333 ( .A(n22234), .B(n22235), .Z(n22233) );
  OR U22334 ( .A(n22236), .B(n22237), .Z(n22235) );
  NAND U22335 ( .A(n22237), .B(n22236), .Z(n22232) );
  ANDN U22336 ( .B(B[220]), .A(n73), .Z(n22016) );
  XNOR U22337 ( .A(n22024), .B(n22238), .Z(n22017) );
  XNOR U22338 ( .A(n22023), .B(n22021), .Z(n22238) );
  AND U22339 ( .A(n22239), .B(n22240), .Z(n22021) );
  NANDN U22340 ( .A(n22241), .B(n22242), .Z(n22240) );
  NANDN U22341 ( .A(n22243), .B(n22244), .Z(n22242) );
  NANDN U22342 ( .A(n22244), .B(n22243), .Z(n22239) );
  ANDN U22343 ( .B(B[221]), .A(n74), .Z(n22023) );
  XNOR U22344 ( .A(n22031), .B(n22245), .Z(n22024) );
  XNOR U22345 ( .A(n22030), .B(n22028), .Z(n22245) );
  AND U22346 ( .A(n22246), .B(n22247), .Z(n22028) );
  NANDN U22347 ( .A(n22248), .B(n22249), .Z(n22247) );
  OR U22348 ( .A(n22250), .B(n22251), .Z(n22249) );
  NAND U22349 ( .A(n22251), .B(n22250), .Z(n22246) );
  ANDN U22350 ( .B(B[222]), .A(n75), .Z(n22030) );
  XNOR U22351 ( .A(n22038), .B(n22252), .Z(n22031) );
  XNOR U22352 ( .A(n22037), .B(n22035), .Z(n22252) );
  AND U22353 ( .A(n22253), .B(n22254), .Z(n22035) );
  NANDN U22354 ( .A(n22255), .B(n22256), .Z(n22254) );
  NANDN U22355 ( .A(n22257), .B(n22258), .Z(n22256) );
  NANDN U22356 ( .A(n22258), .B(n22257), .Z(n22253) );
  ANDN U22357 ( .B(B[223]), .A(n76), .Z(n22037) );
  XNOR U22358 ( .A(n22045), .B(n22259), .Z(n22038) );
  XNOR U22359 ( .A(n22044), .B(n22042), .Z(n22259) );
  AND U22360 ( .A(n22260), .B(n22261), .Z(n22042) );
  NANDN U22361 ( .A(n22262), .B(n22263), .Z(n22261) );
  OR U22362 ( .A(n22264), .B(n22265), .Z(n22263) );
  NAND U22363 ( .A(n22265), .B(n22264), .Z(n22260) );
  ANDN U22364 ( .B(B[224]), .A(n77), .Z(n22044) );
  XNOR U22365 ( .A(n22052), .B(n22266), .Z(n22045) );
  XNOR U22366 ( .A(n22051), .B(n22049), .Z(n22266) );
  AND U22367 ( .A(n22267), .B(n22268), .Z(n22049) );
  NANDN U22368 ( .A(n22269), .B(n22270), .Z(n22268) );
  NANDN U22369 ( .A(n22271), .B(n22272), .Z(n22270) );
  NANDN U22370 ( .A(n22272), .B(n22271), .Z(n22267) );
  ANDN U22371 ( .B(B[225]), .A(n78), .Z(n22051) );
  XNOR U22372 ( .A(n22059), .B(n22273), .Z(n22052) );
  XNOR U22373 ( .A(n22058), .B(n22056), .Z(n22273) );
  AND U22374 ( .A(n22274), .B(n22275), .Z(n22056) );
  NANDN U22375 ( .A(n22276), .B(n22277), .Z(n22275) );
  OR U22376 ( .A(n22278), .B(n22279), .Z(n22277) );
  NAND U22377 ( .A(n22279), .B(n22278), .Z(n22274) );
  ANDN U22378 ( .B(B[226]), .A(n79), .Z(n22058) );
  XNOR U22379 ( .A(n22066), .B(n22280), .Z(n22059) );
  XNOR U22380 ( .A(n22065), .B(n22063), .Z(n22280) );
  AND U22381 ( .A(n22281), .B(n22282), .Z(n22063) );
  NANDN U22382 ( .A(n22283), .B(n22284), .Z(n22282) );
  NANDN U22383 ( .A(n22285), .B(n22286), .Z(n22284) );
  NANDN U22384 ( .A(n22286), .B(n22285), .Z(n22281) );
  ANDN U22385 ( .B(B[227]), .A(n80), .Z(n22065) );
  XNOR U22386 ( .A(n22073), .B(n22287), .Z(n22066) );
  XNOR U22387 ( .A(n22072), .B(n22070), .Z(n22287) );
  AND U22388 ( .A(n22288), .B(n22289), .Z(n22070) );
  NANDN U22389 ( .A(n22290), .B(n22291), .Z(n22289) );
  OR U22390 ( .A(n22292), .B(n22293), .Z(n22291) );
  NAND U22391 ( .A(n22293), .B(n22292), .Z(n22288) );
  ANDN U22392 ( .B(B[228]), .A(n81), .Z(n22072) );
  XNOR U22393 ( .A(n22080), .B(n22294), .Z(n22073) );
  XNOR U22394 ( .A(n22079), .B(n22077), .Z(n22294) );
  AND U22395 ( .A(n22295), .B(n22296), .Z(n22077) );
  NANDN U22396 ( .A(n22297), .B(n22298), .Z(n22296) );
  NAND U22397 ( .A(n22299), .B(n22300), .Z(n22298) );
  ANDN U22398 ( .B(B[229]), .A(n82), .Z(n22079) );
  XOR U22399 ( .A(n22086), .B(n22301), .Z(n22080) );
  XNOR U22400 ( .A(n22084), .B(n22087), .Z(n22301) );
  NAND U22401 ( .A(A[2]), .B(B[230]), .Z(n22087) );
  NANDN U22402 ( .A(n22302), .B(n22303), .Z(n22084) );
  AND U22403 ( .A(A[0]), .B(B[231]), .Z(n22303) );
  XNOR U22404 ( .A(n22089), .B(n22304), .Z(n22086) );
  NAND U22405 ( .A(A[0]), .B(B[232]), .Z(n22304) );
  NAND U22406 ( .A(B[231]), .B(A[1]), .Z(n22089) );
  NAND U22407 ( .A(n22305), .B(n22306), .Z(n332) );
  NANDN U22408 ( .A(n22307), .B(n22308), .Z(n22306) );
  OR U22409 ( .A(n22309), .B(n22310), .Z(n22308) );
  NAND U22410 ( .A(n22310), .B(n22309), .Z(n22305) );
  XOR U22411 ( .A(n20022), .B(n22311), .Z(\A1[22] ) );
  XNOR U22412 ( .A(n20021), .B(n20020), .Z(n22311) );
  NAND U22413 ( .A(n22312), .B(n22313), .Z(n20020) );
  NANDN U22414 ( .A(n22314), .B(n22315), .Z(n22313) );
  OR U22415 ( .A(n22316), .B(n22317), .Z(n22315) );
  NAND U22416 ( .A(n22317), .B(n22316), .Z(n22312) );
  ANDN U22417 ( .B(B[0]), .A(n61), .Z(n20021) );
  XNOR U22418 ( .A(n20029), .B(n22318), .Z(n20022) );
  XNOR U22419 ( .A(n20028), .B(n20026), .Z(n22318) );
  AND U22420 ( .A(n22319), .B(n22320), .Z(n20026) );
  NANDN U22421 ( .A(n22321), .B(n22322), .Z(n22320) );
  NANDN U22422 ( .A(n22323), .B(n22324), .Z(n22322) );
  NANDN U22423 ( .A(n22324), .B(n22323), .Z(n22319) );
  ANDN U22424 ( .B(B[1]), .A(n62), .Z(n20028) );
  XNOR U22425 ( .A(n20036), .B(n22325), .Z(n20029) );
  XNOR U22426 ( .A(n20035), .B(n20033), .Z(n22325) );
  AND U22427 ( .A(n22326), .B(n22327), .Z(n20033) );
  NANDN U22428 ( .A(n22328), .B(n22329), .Z(n22327) );
  OR U22429 ( .A(n22330), .B(n22331), .Z(n22329) );
  NAND U22430 ( .A(n22331), .B(n22330), .Z(n22326) );
  ANDN U22431 ( .B(B[2]), .A(n63), .Z(n20035) );
  XNOR U22432 ( .A(n20043), .B(n22332), .Z(n20036) );
  XNOR U22433 ( .A(n20042), .B(n20040), .Z(n22332) );
  AND U22434 ( .A(n22333), .B(n22334), .Z(n20040) );
  NANDN U22435 ( .A(n22335), .B(n22336), .Z(n22334) );
  NANDN U22436 ( .A(n22337), .B(n22338), .Z(n22336) );
  NANDN U22437 ( .A(n22338), .B(n22337), .Z(n22333) );
  ANDN U22438 ( .B(B[3]), .A(n64), .Z(n20042) );
  XNOR U22439 ( .A(n20050), .B(n22339), .Z(n20043) );
  XNOR U22440 ( .A(n20049), .B(n20047), .Z(n22339) );
  AND U22441 ( .A(n22340), .B(n22341), .Z(n20047) );
  NANDN U22442 ( .A(n22342), .B(n22343), .Z(n22341) );
  OR U22443 ( .A(n22344), .B(n22345), .Z(n22343) );
  NAND U22444 ( .A(n22345), .B(n22344), .Z(n22340) );
  ANDN U22445 ( .B(B[4]), .A(n65), .Z(n20049) );
  XNOR U22446 ( .A(n20057), .B(n22346), .Z(n20050) );
  XNOR U22447 ( .A(n20056), .B(n20054), .Z(n22346) );
  AND U22448 ( .A(n22347), .B(n22348), .Z(n20054) );
  NANDN U22449 ( .A(n22349), .B(n22350), .Z(n22348) );
  NANDN U22450 ( .A(n22351), .B(n22352), .Z(n22350) );
  NANDN U22451 ( .A(n22352), .B(n22351), .Z(n22347) );
  ANDN U22452 ( .B(B[5]), .A(n66), .Z(n20056) );
  XNOR U22453 ( .A(n20064), .B(n22353), .Z(n20057) );
  XNOR U22454 ( .A(n20063), .B(n20061), .Z(n22353) );
  AND U22455 ( .A(n22354), .B(n22355), .Z(n20061) );
  NANDN U22456 ( .A(n22356), .B(n22357), .Z(n22355) );
  OR U22457 ( .A(n22358), .B(n22359), .Z(n22357) );
  NAND U22458 ( .A(n22359), .B(n22358), .Z(n22354) );
  ANDN U22459 ( .B(B[6]), .A(n67), .Z(n20063) );
  XNOR U22460 ( .A(n20071), .B(n22360), .Z(n20064) );
  XNOR U22461 ( .A(n20070), .B(n20068), .Z(n22360) );
  AND U22462 ( .A(n22361), .B(n22362), .Z(n20068) );
  NANDN U22463 ( .A(n22363), .B(n22364), .Z(n22362) );
  NANDN U22464 ( .A(n22365), .B(n22366), .Z(n22364) );
  NANDN U22465 ( .A(n22366), .B(n22365), .Z(n22361) );
  ANDN U22466 ( .B(B[7]), .A(n68), .Z(n20070) );
  XNOR U22467 ( .A(n20078), .B(n22367), .Z(n20071) );
  XNOR U22468 ( .A(n20077), .B(n20075), .Z(n22367) );
  AND U22469 ( .A(n22368), .B(n22369), .Z(n20075) );
  NANDN U22470 ( .A(n22370), .B(n22371), .Z(n22369) );
  OR U22471 ( .A(n22372), .B(n22373), .Z(n22371) );
  NAND U22472 ( .A(n22373), .B(n22372), .Z(n22368) );
  ANDN U22473 ( .B(B[8]), .A(n69), .Z(n20077) );
  XNOR U22474 ( .A(n20085), .B(n22374), .Z(n20078) );
  XNOR U22475 ( .A(n20084), .B(n20082), .Z(n22374) );
  AND U22476 ( .A(n22375), .B(n22376), .Z(n20082) );
  NANDN U22477 ( .A(n22377), .B(n22378), .Z(n22376) );
  NANDN U22478 ( .A(n22379), .B(n22380), .Z(n22378) );
  NANDN U22479 ( .A(n22380), .B(n22379), .Z(n22375) );
  ANDN U22480 ( .B(B[9]), .A(n70), .Z(n20084) );
  XNOR U22481 ( .A(n20092), .B(n22381), .Z(n20085) );
  XNOR U22482 ( .A(n20091), .B(n20089), .Z(n22381) );
  AND U22483 ( .A(n22382), .B(n22383), .Z(n20089) );
  NANDN U22484 ( .A(n22384), .B(n22385), .Z(n22383) );
  OR U22485 ( .A(n22386), .B(n22387), .Z(n22385) );
  NAND U22486 ( .A(n22387), .B(n22386), .Z(n22382) );
  ANDN U22487 ( .B(B[10]), .A(n71), .Z(n20091) );
  XNOR U22488 ( .A(n20099), .B(n22388), .Z(n20092) );
  XNOR U22489 ( .A(n20098), .B(n20096), .Z(n22388) );
  AND U22490 ( .A(n22389), .B(n22390), .Z(n20096) );
  NANDN U22491 ( .A(n22391), .B(n22392), .Z(n22390) );
  NANDN U22492 ( .A(n22393), .B(n22394), .Z(n22392) );
  NANDN U22493 ( .A(n22394), .B(n22393), .Z(n22389) );
  ANDN U22494 ( .B(B[11]), .A(n72), .Z(n20098) );
  XNOR U22495 ( .A(n20106), .B(n22395), .Z(n20099) );
  XNOR U22496 ( .A(n20105), .B(n20103), .Z(n22395) );
  AND U22497 ( .A(n22396), .B(n22397), .Z(n20103) );
  NANDN U22498 ( .A(n22398), .B(n22399), .Z(n22397) );
  OR U22499 ( .A(n22400), .B(n22401), .Z(n22399) );
  NAND U22500 ( .A(n22401), .B(n22400), .Z(n22396) );
  ANDN U22501 ( .B(B[12]), .A(n73), .Z(n20105) );
  XNOR U22502 ( .A(n20113), .B(n22402), .Z(n20106) );
  XNOR U22503 ( .A(n20112), .B(n20110), .Z(n22402) );
  AND U22504 ( .A(n22403), .B(n22404), .Z(n20110) );
  NANDN U22505 ( .A(n22405), .B(n22406), .Z(n22404) );
  NANDN U22506 ( .A(n22407), .B(n22408), .Z(n22406) );
  NANDN U22507 ( .A(n22408), .B(n22407), .Z(n22403) );
  ANDN U22508 ( .B(B[13]), .A(n74), .Z(n20112) );
  XNOR U22509 ( .A(n20120), .B(n22409), .Z(n20113) );
  XNOR U22510 ( .A(n20119), .B(n20117), .Z(n22409) );
  AND U22511 ( .A(n22410), .B(n22411), .Z(n20117) );
  NANDN U22512 ( .A(n22412), .B(n22413), .Z(n22411) );
  OR U22513 ( .A(n22414), .B(n22415), .Z(n22413) );
  NAND U22514 ( .A(n22415), .B(n22414), .Z(n22410) );
  ANDN U22515 ( .B(B[14]), .A(n75), .Z(n20119) );
  XNOR U22516 ( .A(n20127), .B(n22416), .Z(n20120) );
  XNOR U22517 ( .A(n20126), .B(n20124), .Z(n22416) );
  AND U22518 ( .A(n22417), .B(n22418), .Z(n20124) );
  NANDN U22519 ( .A(n22419), .B(n22420), .Z(n22418) );
  NANDN U22520 ( .A(n22421), .B(n22422), .Z(n22420) );
  NANDN U22521 ( .A(n22422), .B(n22421), .Z(n22417) );
  ANDN U22522 ( .B(B[15]), .A(n76), .Z(n20126) );
  XNOR U22523 ( .A(n20134), .B(n22423), .Z(n20127) );
  XNOR U22524 ( .A(n20133), .B(n20131), .Z(n22423) );
  AND U22525 ( .A(n22424), .B(n22425), .Z(n20131) );
  NANDN U22526 ( .A(n22426), .B(n22427), .Z(n22425) );
  OR U22527 ( .A(n22428), .B(n22429), .Z(n22427) );
  NAND U22528 ( .A(n22429), .B(n22428), .Z(n22424) );
  ANDN U22529 ( .B(B[16]), .A(n77), .Z(n20133) );
  XNOR U22530 ( .A(n20141), .B(n22430), .Z(n20134) );
  XNOR U22531 ( .A(n20140), .B(n20138), .Z(n22430) );
  AND U22532 ( .A(n22431), .B(n22432), .Z(n20138) );
  NANDN U22533 ( .A(n22433), .B(n22434), .Z(n22432) );
  NANDN U22534 ( .A(n22435), .B(n22436), .Z(n22434) );
  NANDN U22535 ( .A(n22436), .B(n22435), .Z(n22431) );
  ANDN U22536 ( .B(B[17]), .A(n78), .Z(n20140) );
  XNOR U22537 ( .A(n20148), .B(n22437), .Z(n20141) );
  XNOR U22538 ( .A(n20147), .B(n20145), .Z(n22437) );
  AND U22539 ( .A(n22438), .B(n22439), .Z(n20145) );
  NANDN U22540 ( .A(n22440), .B(n22441), .Z(n22439) );
  OR U22541 ( .A(n22442), .B(n22443), .Z(n22441) );
  NAND U22542 ( .A(n22443), .B(n22442), .Z(n22438) );
  ANDN U22543 ( .B(B[18]), .A(n79), .Z(n20147) );
  XNOR U22544 ( .A(n20155), .B(n22444), .Z(n20148) );
  XNOR U22545 ( .A(n20154), .B(n20152), .Z(n22444) );
  AND U22546 ( .A(n22445), .B(n22446), .Z(n20152) );
  NANDN U22547 ( .A(n22447), .B(n22448), .Z(n22446) );
  NANDN U22548 ( .A(n22449), .B(n22450), .Z(n22448) );
  NANDN U22549 ( .A(n22450), .B(n22449), .Z(n22445) );
  ANDN U22550 ( .B(B[19]), .A(n80), .Z(n20154) );
  XNOR U22551 ( .A(n20162), .B(n22451), .Z(n20155) );
  XNOR U22552 ( .A(n20161), .B(n20159), .Z(n22451) );
  AND U22553 ( .A(n22452), .B(n22453), .Z(n20159) );
  NANDN U22554 ( .A(n22454), .B(n22455), .Z(n22453) );
  OR U22555 ( .A(n22456), .B(n22457), .Z(n22455) );
  NAND U22556 ( .A(n22457), .B(n22456), .Z(n22452) );
  ANDN U22557 ( .B(B[20]), .A(n81), .Z(n20161) );
  XNOR U22558 ( .A(n20169), .B(n22458), .Z(n20162) );
  XNOR U22559 ( .A(n20168), .B(n20166), .Z(n22458) );
  AND U22560 ( .A(n22459), .B(n22460), .Z(n20166) );
  NANDN U22561 ( .A(n22461), .B(n22462), .Z(n22460) );
  NAND U22562 ( .A(n22463), .B(n22464), .Z(n22462) );
  ANDN U22563 ( .B(B[21]), .A(n82), .Z(n20168) );
  XOR U22564 ( .A(n20175), .B(n22465), .Z(n20169) );
  XNOR U22565 ( .A(n20173), .B(n20176), .Z(n22465) );
  NAND U22566 ( .A(A[2]), .B(B[22]), .Z(n20176) );
  NANDN U22567 ( .A(n22466), .B(n22467), .Z(n20173) );
  AND U22568 ( .A(A[0]), .B(B[23]), .Z(n22467) );
  XNOR U22569 ( .A(n20178), .B(n22468), .Z(n20175) );
  NAND U22570 ( .A(A[0]), .B(B[24]), .Z(n22468) );
  NAND U22571 ( .A(B[23]), .B(A[1]), .Z(n20178) );
  XOR U22572 ( .A(n334), .B(n333), .Z(\A1[229] ) );
  XOR U22573 ( .A(n22310), .B(n22469), .Z(n333) );
  XNOR U22574 ( .A(n22309), .B(n22307), .Z(n22469) );
  AND U22575 ( .A(n22470), .B(n22471), .Z(n22307) );
  NANDN U22576 ( .A(n22472), .B(n22473), .Z(n22471) );
  NANDN U22577 ( .A(n22474), .B(n22475), .Z(n22473) );
  NANDN U22578 ( .A(n22475), .B(n22474), .Z(n22470) );
  ANDN U22579 ( .B(B[200]), .A(n54), .Z(n22309) );
  XNOR U22580 ( .A(n22104), .B(n22476), .Z(n22310) );
  XNOR U22581 ( .A(n22103), .B(n22101), .Z(n22476) );
  AND U22582 ( .A(n22477), .B(n22478), .Z(n22101) );
  NANDN U22583 ( .A(n22479), .B(n22480), .Z(n22478) );
  OR U22584 ( .A(n22481), .B(n22482), .Z(n22480) );
  NAND U22585 ( .A(n22482), .B(n22481), .Z(n22477) );
  ANDN U22586 ( .B(B[201]), .A(n55), .Z(n22103) );
  XNOR U22587 ( .A(n22111), .B(n22483), .Z(n22104) );
  XNOR U22588 ( .A(n22110), .B(n22108), .Z(n22483) );
  AND U22589 ( .A(n22484), .B(n22485), .Z(n22108) );
  NANDN U22590 ( .A(n22486), .B(n22487), .Z(n22485) );
  NANDN U22591 ( .A(n22488), .B(n22489), .Z(n22487) );
  NANDN U22592 ( .A(n22489), .B(n22488), .Z(n22484) );
  ANDN U22593 ( .B(B[202]), .A(n56), .Z(n22110) );
  XNOR U22594 ( .A(n22118), .B(n22490), .Z(n22111) );
  XNOR U22595 ( .A(n22117), .B(n22115), .Z(n22490) );
  AND U22596 ( .A(n22491), .B(n22492), .Z(n22115) );
  NANDN U22597 ( .A(n22493), .B(n22494), .Z(n22492) );
  OR U22598 ( .A(n22495), .B(n22496), .Z(n22494) );
  NAND U22599 ( .A(n22496), .B(n22495), .Z(n22491) );
  ANDN U22600 ( .B(B[203]), .A(n57), .Z(n22117) );
  XNOR U22601 ( .A(n22125), .B(n22497), .Z(n22118) );
  XNOR U22602 ( .A(n22124), .B(n22122), .Z(n22497) );
  AND U22603 ( .A(n22498), .B(n22499), .Z(n22122) );
  NANDN U22604 ( .A(n22500), .B(n22501), .Z(n22499) );
  NANDN U22605 ( .A(n22502), .B(n22503), .Z(n22501) );
  NANDN U22606 ( .A(n22503), .B(n22502), .Z(n22498) );
  ANDN U22607 ( .B(B[204]), .A(n58), .Z(n22124) );
  XNOR U22608 ( .A(n22132), .B(n22504), .Z(n22125) );
  XNOR U22609 ( .A(n22131), .B(n22129), .Z(n22504) );
  AND U22610 ( .A(n22505), .B(n22506), .Z(n22129) );
  NANDN U22611 ( .A(n22507), .B(n22508), .Z(n22506) );
  OR U22612 ( .A(n22509), .B(n22510), .Z(n22508) );
  NAND U22613 ( .A(n22510), .B(n22509), .Z(n22505) );
  ANDN U22614 ( .B(B[205]), .A(n59), .Z(n22131) );
  XNOR U22615 ( .A(n22139), .B(n22511), .Z(n22132) );
  XNOR U22616 ( .A(n22138), .B(n22136), .Z(n22511) );
  AND U22617 ( .A(n22512), .B(n22513), .Z(n22136) );
  NANDN U22618 ( .A(n22514), .B(n22515), .Z(n22513) );
  NANDN U22619 ( .A(n22516), .B(n22517), .Z(n22515) );
  NANDN U22620 ( .A(n22517), .B(n22516), .Z(n22512) );
  ANDN U22621 ( .B(B[206]), .A(n60), .Z(n22138) );
  XNOR U22622 ( .A(n22146), .B(n22518), .Z(n22139) );
  XNOR U22623 ( .A(n22145), .B(n22143), .Z(n22518) );
  AND U22624 ( .A(n22519), .B(n22520), .Z(n22143) );
  NANDN U22625 ( .A(n22521), .B(n22522), .Z(n22520) );
  OR U22626 ( .A(n22523), .B(n22524), .Z(n22522) );
  NAND U22627 ( .A(n22524), .B(n22523), .Z(n22519) );
  ANDN U22628 ( .B(B[207]), .A(n61), .Z(n22145) );
  XNOR U22629 ( .A(n22153), .B(n22525), .Z(n22146) );
  XNOR U22630 ( .A(n22152), .B(n22150), .Z(n22525) );
  AND U22631 ( .A(n22526), .B(n22527), .Z(n22150) );
  NANDN U22632 ( .A(n22528), .B(n22529), .Z(n22527) );
  NANDN U22633 ( .A(n22530), .B(n22531), .Z(n22529) );
  NANDN U22634 ( .A(n22531), .B(n22530), .Z(n22526) );
  ANDN U22635 ( .B(B[208]), .A(n62), .Z(n22152) );
  XNOR U22636 ( .A(n22160), .B(n22532), .Z(n22153) );
  XNOR U22637 ( .A(n22159), .B(n22157), .Z(n22532) );
  AND U22638 ( .A(n22533), .B(n22534), .Z(n22157) );
  NANDN U22639 ( .A(n22535), .B(n22536), .Z(n22534) );
  OR U22640 ( .A(n22537), .B(n22538), .Z(n22536) );
  NAND U22641 ( .A(n22538), .B(n22537), .Z(n22533) );
  ANDN U22642 ( .B(B[209]), .A(n63), .Z(n22159) );
  XNOR U22643 ( .A(n22167), .B(n22539), .Z(n22160) );
  XNOR U22644 ( .A(n22166), .B(n22164), .Z(n22539) );
  AND U22645 ( .A(n22540), .B(n22541), .Z(n22164) );
  NANDN U22646 ( .A(n22542), .B(n22543), .Z(n22541) );
  NANDN U22647 ( .A(n22544), .B(n22545), .Z(n22543) );
  NANDN U22648 ( .A(n22545), .B(n22544), .Z(n22540) );
  ANDN U22649 ( .B(B[210]), .A(n64), .Z(n22166) );
  XNOR U22650 ( .A(n22174), .B(n22546), .Z(n22167) );
  XNOR U22651 ( .A(n22173), .B(n22171), .Z(n22546) );
  AND U22652 ( .A(n22547), .B(n22548), .Z(n22171) );
  NANDN U22653 ( .A(n22549), .B(n22550), .Z(n22548) );
  OR U22654 ( .A(n22551), .B(n22552), .Z(n22550) );
  NAND U22655 ( .A(n22552), .B(n22551), .Z(n22547) );
  ANDN U22656 ( .B(B[211]), .A(n65), .Z(n22173) );
  XNOR U22657 ( .A(n22181), .B(n22553), .Z(n22174) );
  XNOR U22658 ( .A(n22180), .B(n22178), .Z(n22553) );
  AND U22659 ( .A(n22554), .B(n22555), .Z(n22178) );
  NANDN U22660 ( .A(n22556), .B(n22557), .Z(n22555) );
  NANDN U22661 ( .A(n22558), .B(n22559), .Z(n22557) );
  NANDN U22662 ( .A(n22559), .B(n22558), .Z(n22554) );
  ANDN U22663 ( .B(B[212]), .A(n66), .Z(n22180) );
  XNOR U22664 ( .A(n22188), .B(n22560), .Z(n22181) );
  XNOR U22665 ( .A(n22187), .B(n22185), .Z(n22560) );
  AND U22666 ( .A(n22561), .B(n22562), .Z(n22185) );
  NANDN U22667 ( .A(n22563), .B(n22564), .Z(n22562) );
  OR U22668 ( .A(n22565), .B(n22566), .Z(n22564) );
  NAND U22669 ( .A(n22566), .B(n22565), .Z(n22561) );
  ANDN U22670 ( .B(B[213]), .A(n67), .Z(n22187) );
  XNOR U22671 ( .A(n22195), .B(n22567), .Z(n22188) );
  XNOR U22672 ( .A(n22194), .B(n22192), .Z(n22567) );
  AND U22673 ( .A(n22568), .B(n22569), .Z(n22192) );
  NANDN U22674 ( .A(n22570), .B(n22571), .Z(n22569) );
  NANDN U22675 ( .A(n22572), .B(n22573), .Z(n22571) );
  NANDN U22676 ( .A(n22573), .B(n22572), .Z(n22568) );
  ANDN U22677 ( .B(B[214]), .A(n68), .Z(n22194) );
  XNOR U22678 ( .A(n22202), .B(n22574), .Z(n22195) );
  XNOR U22679 ( .A(n22201), .B(n22199), .Z(n22574) );
  AND U22680 ( .A(n22575), .B(n22576), .Z(n22199) );
  NANDN U22681 ( .A(n22577), .B(n22578), .Z(n22576) );
  OR U22682 ( .A(n22579), .B(n22580), .Z(n22578) );
  NAND U22683 ( .A(n22580), .B(n22579), .Z(n22575) );
  ANDN U22684 ( .B(B[215]), .A(n69), .Z(n22201) );
  XNOR U22685 ( .A(n22209), .B(n22581), .Z(n22202) );
  XNOR U22686 ( .A(n22208), .B(n22206), .Z(n22581) );
  AND U22687 ( .A(n22582), .B(n22583), .Z(n22206) );
  NANDN U22688 ( .A(n22584), .B(n22585), .Z(n22583) );
  NANDN U22689 ( .A(n22586), .B(n22587), .Z(n22585) );
  NANDN U22690 ( .A(n22587), .B(n22586), .Z(n22582) );
  ANDN U22691 ( .B(B[216]), .A(n70), .Z(n22208) );
  XNOR U22692 ( .A(n22216), .B(n22588), .Z(n22209) );
  XNOR U22693 ( .A(n22215), .B(n22213), .Z(n22588) );
  AND U22694 ( .A(n22589), .B(n22590), .Z(n22213) );
  NANDN U22695 ( .A(n22591), .B(n22592), .Z(n22590) );
  OR U22696 ( .A(n22593), .B(n22594), .Z(n22592) );
  NAND U22697 ( .A(n22594), .B(n22593), .Z(n22589) );
  ANDN U22698 ( .B(B[217]), .A(n71), .Z(n22215) );
  XNOR U22699 ( .A(n22223), .B(n22595), .Z(n22216) );
  XNOR U22700 ( .A(n22222), .B(n22220), .Z(n22595) );
  AND U22701 ( .A(n22596), .B(n22597), .Z(n22220) );
  NANDN U22702 ( .A(n22598), .B(n22599), .Z(n22597) );
  NANDN U22703 ( .A(n22600), .B(n22601), .Z(n22599) );
  NANDN U22704 ( .A(n22601), .B(n22600), .Z(n22596) );
  ANDN U22705 ( .B(B[218]), .A(n72), .Z(n22222) );
  XNOR U22706 ( .A(n22230), .B(n22602), .Z(n22223) );
  XNOR U22707 ( .A(n22229), .B(n22227), .Z(n22602) );
  AND U22708 ( .A(n22603), .B(n22604), .Z(n22227) );
  NANDN U22709 ( .A(n22605), .B(n22606), .Z(n22604) );
  OR U22710 ( .A(n22607), .B(n22608), .Z(n22606) );
  NAND U22711 ( .A(n22608), .B(n22607), .Z(n22603) );
  ANDN U22712 ( .B(B[219]), .A(n73), .Z(n22229) );
  XNOR U22713 ( .A(n22237), .B(n22609), .Z(n22230) );
  XNOR U22714 ( .A(n22236), .B(n22234), .Z(n22609) );
  AND U22715 ( .A(n22610), .B(n22611), .Z(n22234) );
  NANDN U22716 ( .A(n22612), .B(n22613), .Z(n22611) );
  NANDN U22717 ( .A(n22614), .B(n22615), .Z(n22613) );
  NANDN U22718 ( .A(n22615), .B(n22614), .Z(n22610) );
  ANDN U22719 ( .B(B[220]), .A(n74), .Z(n22236) );
  XNOR U22720 ( .A(n22244), .B(n22616), .Z(n22237) );
  XNOR U22721 ( .A(n22243), .B(n22241), .Z(n22616) );
  AND U22722 ( .A(n22617), .B(n22618), .Z(n22241) );
  NANDN U22723 ( .A(n22619), .B(n22620), .Z(n22618) );
  OR U22724 ( .A(n22621), .B(n22622), .Z(n22620) );
  NAND U22725 ( .A(n22622), .B(n22621), .Z(n22617) );
  ANDN U22726 ( .B(B[221]), .A(n75), .Z(n22243) );
  XNOR U22727 ( .A(n22251), .B(n22623), .Z(n22244) );
  XNOR U22728 ( .A(n22250), .B(n22248), .Z(n22623) );
  AND U22729 ( .A(n22624), .B(n22625), .Z(n22248) );
  NANDN U22730 ( .A(n22626), .B(n22627), .Z(n22625) );
  NANDN U22731 ( .A(n22628), .B(n22629), .Z(n22627) );
  NANDN U22732 ( .A(n22629), .B(n22628), .Z(n22624) );
  ANDN U22733 ( .B(B[222]), .A(n76), .Z(n22250) );
  XNOR U22734 ( .A(n22258), .B(n22630), .Z(n22251) );
  XNOR U22735 ( .A(n22257), .B(n22255), .Z(n22630) );
  AND U22736 ( .A(n22631), .B(n22632), .Z(n22255) );
  NANDN U22737 ( .A(n22633), .B(n22634), .Z(n22632) );
  OR U22738 ( .A(n22635), .B(n22636), .Z(n22634) );
  NAND U22739 ( .A(n22636), .B(n22635), .Z(n22631) );
  ANDN U22740 ( .B(B[223]), .A(n77), .Z(n22257) );
  XNOR U22741 ( .A(n22265), .B(n22637), .Z(n22258) );
  XNOR U22742 ( .A(n22264), .B(n22262), .Z(n22637) );
  AND U22743 ( .A(n22638), .B(n22639), .Z(n22262) );
  NANDN U22744 ( .A(n22640), .B(n22641), .Z(n22639) );
  NANDN U22745 ( .A(n22642), .B(n22643), .Z(n22641) );
  NANDN U22746 ( .A(n22643), .B(n22642), .Z(n22638) );
  ANDN U22747 ( .B(B[224]), .A(n78), .Z(n22264) );
  XNOR U22748 ( .A(n22272), .B(n22644), .Z(n22265) );
  XNOR U22749 ( .A(n22271), .B(n22269), .Z(n22644) );
  AND U22750 ( .A(n22645), .B(n22646), .Z(n22269) );
  NANDN U22751 ( .A(n22647), .B(n22648), .Z(n22646) );
  OR U22752 ( .A(n22649), .B(n22650), .Z(n22648) );
  NAND U22753 ( .A(n22650), .B(n22649), .Z(n22645) );
  ANDN U22754 ( .B(B[225]), .A(n79), .Z(n22271) );
  XNOR U22755 ( .A(n22279), .B(n22651), .Z(n22272) );
  XNOR U22756 ( .A(n22278), .B(n22276), .Z(n22651) );
  AND U22757 ( .A(n22652), .B(n22653), .Z(n22276) );
  NANDN U22758 ( .A(n22654), .B(n22655), .Z(n22653) );
  NANDN U22759 ( .A(n22656), .B(n22657), .Z(n22655) );
  NANDN U22760 ( .A(n22657), .B(n22656), .Z(n22652) );
  ANDN U22761 ( .B(B[226]), .A(n80), .Z(n22278) );
  XNOR U22762 ( .A(n22286), .B(n22658), .Z(n22279) );
  XNOR U22763 ( .A(n22285), .B(n22283), .Z(n22658) );
  AND U22764 ( .A(n22659), .B(n22660), .Z(n22283) );
  NANDN U22765 ( .A(n22661), .B(n22662), .Z(n22660) );
  OR U22766 ( .A(n22663), .B(n22664), .Z(n22662) );
  NAND U22767 ( .A(n22664), .B(n22663), .Z(n22659) );
  ANDN U22768 ( .B(B[227]), .A(n81), .Z(n22285) );
  XNOR U22769 ( .A(n22293), .B(n22665), .Z(n22286) );
  XNOR U22770 ( .A(n22292), .B(n22290), .Z(n22665) );
  AND U22771 ( .A(n22666), .B(n22667), .Z(n22290) );
  NANDN U22772 ( .A(n22668), .B(n22669), .Z(n22667) );
  NAND U22773 ( .A(n22670), .B(n22671), .Z(n22669) );
  ANDN U22774 ( .B(B[228]), .A(n82), .Z(n22292) );
  XOR U22775 ( .A(n22299), .B(n22672), .Z(n22293) );
  XNOR U22776 ( .A(n22297), .B(n22300), .Z(n22672) );
  NAND U22777 ( .A(A[2]), .B(B[229]), .Z(n22300) );
  NANDN U22778 ( .A(n22673), .B(n22674), .Z(n22297) );
  AND U22779 ( .A(A[0]), .B(B[230]), .Z(n22674) );
  XNOR U22780 ( .A(n22302), .B(n22675), .Z(n22299) );
  NAND U22781 ( .A(A[0]), .B(B[231]), .Z(n22675) );
  NAND U22782 ( .A(B[230]), .B(A[1]), .Z(n22302) );
  NAND U22783 ( .A(n22676), .B(n22677), .Z(n334) );
  NANDN U22784 ( .A(n22678), .B(n22679), .Z(n22677) );
  OR U22785 ( .A(n22680), .B(n22681), .Z(n22679) );
  NAND U22786 ( .A(n22681), .B(n22680), .Z(n22676) );
  XOR U22787 ( .A(n336), .B(n335), .Z(\A1[228] ) );
  XOR U22788 ( .A(n22681), .B(n22682), .Z(n335) );
  XNOR U22789 ( .A(n22680), .B(n22678), .Z(n22682) );
  AND U22790 ( .A(n22683), .B(n22684), .Z(n22678) );
  NANDN U22791 ( .A(n22685), .B(n22686), .Z(n22684) );
  NANDN U22792 ( .A(n22687), .B(n22688), .Z(n22686) );
  NANDN U22793 ( .A(n22688), .B(n22687), .Z(n22683) );
  ANDN U22794 ( .B(B[199]), .A(n54), .Z(n22680) );
  XNOR U22795 ( .A(n22475), .B(n22689), .Z(n22681) );
  XNOR U22796 ( .A(n22474), .B(n22472), .Z(n22689) );
  AND U22797 ( .A(n22690), .B(n22691), .Z(n22472) );
  NANDN U22798 ( .A(n22692), .B(n22693), .Z(n22691) );
  OR U22799 ( .A(n22694), .B(n22695), .Z(n22693) );
  NAND U22800 ( .A(n22695), .B(n22694), .Z(n22690) );
  ANDN U22801 ( .B(B[200]), .A(n55), .Z(n22474) );
  XNOR U22802 ( .A(n22482), .B(n22696), .Z(n22475) );
  XNOR U22803 ( .A(n22481), .B(n22479), .Z(n22696) );
  AND U22804 ( .A(n22697), .B(n22698), .Z(n22479) );
  NANDN U22805 ( .A(n22699), .B(n22700), .Z(n22698) );
  NANDN U22806 ( .A(n22701), .B(n22702), .Z(n22700) );
  NANDN U22807 ( .A(n22702), .B(n22701), .Z(n22697) );
  ANDN U22808 ( .B(B[201]), .A(n56), .Z(n22481) );
  XNOR U22809 ( .A(n22489), .B(n22703), .Z(n22482) );
  XNOR U22810 ( .A(n22488), .B(n22486), .Z(n22703) );
  AND U22811 ( .A(n22704), .B(n22705), .Z(n22486) );
  NANDN U22812 ( .A(n22706), .B(n22707), .Z(n22705) );
  OR U22813 ( .A(n22708), .B(n22709), .Z(n22707) );
  NAND U22814 ( .A(n22709), .B(n22708), .Z(n22704) );
  ANDN U22815 ( .B(B[202]), .A(n57), .Z(n22488) );
  XNOR U22816 ( .A(n22496), .B(n22710), .Z(n22489) );
  XNOR U22817 ( .A(n22495), .B(n22493), .Z(n22710) );
  AND U22818 ( .A(n22711), .B(n22712), .Z(n22493) );
  NANDN U22819 ( .A(n22713), .B(n22714), .Z(n22712) );
  NANDN U22820 ( .A(n22715), .B(n22716), .Z(n22714) );
  NANDN U22821 ( .A(n22716), .B(n22715), .Z(n22711) );
  ANDN U22822 ( .B(B[203]), .A(n58), .Z(n22495) );
  XNOR U22823 ( .A(n22503), .B(n22717), .Z(n22496) );
  XNOR U22824 ( .A(n22502), .B(n22500), .Z(n22717) );
  AND U22825 ( .A(n22718), .B(n22719), .Z(n22500) );
  NANDN U22826 ( .A(n22720), .B(n22721), .Z(n22719) );
  OR U22827 ( .A(n22722), .B(n22723), .Z(n22721) );
  NAND U22828 ( .A(n22723), .B(n22722), .Z(n22718) );
  ANDN U22829 ( .B(B[204]), .A(n59), .Z(n22502) );
  XNOR U22830 ( .A(n22510), .B(n22724), .Z(n22503) );
  XNOR U22831 ( .A(n22509), .B(n22507), .Z(n22724) );
  AND U22832 ( .A(n22725), .B(n22726), .Z(n22507) );
  NANDN U22833 ( .A(n22727), .B(n22728), .Z(n22726) );
  NANDN U22834 ( .A(n22729), .B(n22730), .Z(n22728) );
  NANDN U22835 ( .A(n22730), .B(n22729), .Z(n22725) );
  ANDN U22836 ( .B(B[205]), .A(n60), .Z(n22509) );
  XNOR U22837 ( .A(n22517), .B(n22731), .Z(n22510) );
  XNOR U22838 ( .A(n22516), .B(n22514), .Z(n22731) );
  AND U22839 ( .A(n22732), .B(n22733), .Z(n22514) );
  NANDN U22840 ( .A(n22734), .B(n22735), .Z(n22733) );
  OR U22841 ( .A(n22736), .B(n22737), .Z(n22735) );
  NAND U22842 ( .A(n22737), .B(n22736), .Z(n22732) );
  ANDN U22843 ( .B(B[206]), .A(n61), .Z(n22516) );
  XNOR U22844 ( .A(n22524), .B(n22738), .Z(n22517) );
  XNOR U22845 ( .A(n22523), .B(n22521), .Z(n22738) );
  AND U22846 ( .A(n22739), .B(n22740), .Z(n22521) );
  NANDN U22847 ( .A(n22741), .B(n22742), .Z(n22740) );
  NANDN U22848 ( .A(n22743), .B(n22744), .Z(n22742) );
  NANDN U22849 ( .A(n22744), .B(n22743), .Z(n22739) );
  ANDN U22850 ( .B(B[207]), .A(n62), .Z(n22523) );
  XNOR U22851 ( .A(n22531), .B(n22745), .Z(n22524) );
  XNOR U22852 ( .A(n22530), .B(n22528), .Z(n22745) );
  AND U22853 ( .A(n22746), .B(n22747), .Z(n22528) );
  NANDN U22854 ( .A(n22748), .B(n22749), .Z(n22747) );
  OR U22855 ( .A(n22750), .B(n22751), .Z(n22749) );
  NAND U22856 ( .A(n22751), .B(n22750), .Z(n22746) );
  ANDN U22857 ( .B(B[208]), .A(n63), .Z(n22530) );
  XNOR U22858 ( .A(n22538), .B(n22752), .Z(n22531) );
  XNOR U22859 ( .A(n22537), .B(n22535), .Z(n22752) );
  AND U22860 ( .A(n22753), .B(n22754), .Z(n22535) );
  NANDN U22861 ( .A(n22755), .B(n22756), .Z(n22754) );
  NANDN U22862 ( .A(n22757), .B(n22758), .Z(n22756) );
  NANDN U22863 ( .A(n22758), .B(n22757), .Z(n22753) );
  ANDN U22864 ( .B(B[209]), .A(n64), .Z(n22537) );
  XNOR U22865 ( .A(n22545), .B(n22759), .Z(n22538) );
  XNOR U22866 ( .A(n22544), .B(n22542), .Z(n22759) );
  AND U22867 ( .A(n22760), .B(n22761), .Z(n22542) );
  NANDN U22868 ( .A(n22762), .B(n22763), .Z(n22761) );
  OR U22869 ( .A(n22764), .B(n22765), .Z(n22763) );
  NAND U22870 ( .A(n22765), .B(n22764), .Z(n22760) );
  ANDN U22871 ( .B(B[210]), .A(n65), .Z(n22544) );
  XNOR U22872 ( .A(n22552), .B(n22766), .Z(n22545) );
  XNOR U22873 ( .A(n22551), .B(n22549), .Z(n22766) );
  AND U22874 ( .A(n22767), .B(n22768), .Z(n22549) );
  NANDN U22875 ( .A(n22769), .B(n22770), .Z(n22768) );
  NANDN U22876 ( .A(n22771), .B(n22772), .Z(n22770) );
  NANDN U22877 ( .A(n22772), .B(n22771), .Z(n22767) );
  ANDN U22878 ( .B(B[211]), .A(n66), .Z(n22551) );
  XNOR U22879 ( .A(n22559), .B(n22773), .Z(n22552) );
  XNOR U22880 ( .A(n22558), .B(n22556), .Z(n22773) );
  AND U22881 ( .A(n22774), .B(n22775), .Z(n22556) );
  NANDN U22882 ( .A(n22776), .B(n22777), .Z(n22775) );
  OR U22883 ( .A(n22778), .B(n22779), .Z(n22777) );
  NAND U22884 ( .A(n22779), .B(n22778), .Z(n22774) );
  ANDN U22885 ( .B(B[212]), .A(n67), .Z(n22558) );
  XNOR U22886 ( .A(n22566), .B(n22780), .Z(n22559) );
  XNOR U22887 ( .A(n22565), .B(n22563), .Z(n22780) );
  AND U22888 ( .A(n22781), .B(n22782), .Z(n22563) );
  NANDN U22889 ( .A(n22783), .B(n22784), .Z(n22782) );
  NANDN U22890 ( .A(n22785), .B(n22786), .Z(n22784) );
  NANDN U22891 ( .A(n22786), .B(n22785), .Z(n22781) );
  ANDN U22892 ( .B(B[213]), .A(n68), .Z(n22565) );
  XNOR U22893 ( .A(n22573), .B(n22787), .Z(n22566) );
  XNOR U22894 ( .A(n22572), .B(n22570), .Z(n22787) );
  AND U22895 ( .A(n22788), .B(n22789), .Z(n22570) );
  NANDN U22896 ( .A(n22790), .B(n22791), .Z(n22789) );
  OR U22897 ( .A(n22792), .B(n22793), .Z(n22791) );
  NAND U22898 ( .A(n22793), .B(n22792), .Z(n22788) );
  ANDN U22899 ( .B(B[214]), .A(n69), .Z(n22572) );
  XNOR U22900 ( .A(n22580), .B(n22794), .Z(n22573) );
  XNOR U22901 ( .A(n22579), .B(n22577), .Z(n22794) );
  AND U22902 ( .A(n22795), .B(n22796), .Z(n22577) );
  NANDN U22903 ( .A(n22797), .B(n22798), .Z(n22796) );
  NANDN U22904 ( .A(n22799), .B(n22800), .Z(n22798) );
  NANDN U22905 ( .A(n22800), .B(n22799), .Z(n22795) );
  ANDN U22906 ( .B(B[215]), .A(n70), .Z(n22579) );
  XNOR U22907 ( .A(n22587), .B(n22801), .Z(n22580) );
  XNOR U22908 ( .A(n22586), .B(n22584), .Z(n22801) );
  AND U22909 ( .A(n22802), .B(n22803), .Z(n22584) );
  NANDN U22910 ( .A(n22804), .B(n22805), .Z(n22803) );
  OR U22911 ( .A(n22806), .B(n22807), .Z(n22805) );
  NAND U22912 ( .A(n22807), .B(n22806), .Z(n22802) );
  ANDN U22913 ( .B(B[216]), .A(n71), .Z(n22586) );
  XNOR U22914 ( .A(n22594), .B(n22808), .Z(n22587) );
  XNOR U22915 ( .A(n22593), .B(n22591), .Z(n22808) );
  AND U22916 ( .A(n22809), .B(n22810), .Z(n22591) );
  NANDN U22917 ( .A(n22811), .B(n22812), .Z(n22810) );
  NANDN U22918 ( .A(n22813), .B(n22814), .Z(n22812) );
  NANDN U22919 ( .A(n22814), .B(n22813), .Z(n22809) );
  ANDN U22920 ( .B(B[217]), .A(n72), .Z(n22593) );
  XNOR U22921 ( .A(n22601), .B(n22815), .Z(n22594) );
  XNOR U22922 ( .A(n22600), .B(n22598), .Z(n22815) );
  AND U22923 ( .A(n22816), .B(n22817), .Z(n22598) );
  NANDN U22924 ( .A(n22818), .B(n22819), .Z(n22817) );
  OR U22925 ( .A(n22820), .B(n22821), .Z(n22819) );
  NAND U22926 ( .A(n22821), .B(n22820), .Z(n22816) );
  ANDN U22927 ( .B(B[218]), .A(n73), .Z(n22600) );
  XNOR U22928 ( .A(n22608), .B(n22822), .Z(n22601) );
  XNOR U22929 ( .A(n22607), .B(n22605), .Z(n22822) );
  AND U22930 ( .A(n22823), .B(n22824), .Z(n22605) );
  NANDN U22931 ( .A(n22825), .B(n22826), .Z(n22824) );
  NANDN U22932 ( .A(n22827), .B(n22828), .Z(n22826) );
  NANDN U22933 ( .A(n22828), .B(n22827), .Z(n22823) );
  ANDN U22934 ( .B(B[219]), .A(n74), .Z(n22607) );
  XNOR U22935 ( .A(n22615), .B(n22829), .Z(n22608) );
  XNOR U22936 ( .A(n22614), .B(n22612), .Z(n22829) );
  AND U22937 ( .A(n22830), .B(n22831), .Z(n22612) );
  NANDN U22938 ( .A(n22832), .B(n22833), .Z(n22831) );
  OR U22939 ( .A(n22834), .B(n22835), .Z(n22833) );
  NAND U22940 ( .A(n22835), .B(n22834), .Z(n22830) );
  ANDN U22941 ( .B(B[220]), .A(n75), .Z(n22614) );
  XNOR U22942 ( .A(n22622), .B(n22836), .Z(n22615) );
  XNOR U22943 ( .A(n22621), .B(n22619), .Z(n22836) );
  AND U22944 ( .A(n22837), .B(n22838), .Z(n22619) );
  NANDN U22945 ( .A(n22839), .B(n22840), .Z(n22838) );
  NANDN U22946 ( .A(n22841), .B(n22842), .Z(n22840) );
  NANDN U22947 ( .A(n22842), .B(n22841), .Z(n22837) );
  ANDN U22948 ( .B(B[221]), .A(n76), .Z(n22621) );
  XNOR U22949 ( .A(n22629), .B(n22843), .Z(n22622) );
  XNOR U22950 ( .A(n22628), .B(n22626), .Z(n22843) );
  AND U22951 ( .A(n22844), .B(n22845), .Z(n22626) );
  NANDN U22952 ( .A(n22846), .B(n22847), .Z(n22845) );
  OR U22953 ( .A(n22848), .B(n22849), .Z(n22847) );
  NAND U22954 ( .A(n22849), .B(n22848), .Z(n22844) );
  ANDN U22955 ( .B(B[222]), .A(n77), .Z(n22628) );
  XNOR U22956 ( .A(n22636), .B(n22850), .Z(n22629) );
  XNOR U22957 ( .A(n22635), .B(n22633), .Z(n22850) );
  AND U22958 ( .A(n22851), .B(n22852), .Z(n22633) );
  NANDN U22959 ( .A(n22853), .B(n22854), .Z(n22852) );
  NANDN U22960 ( .A(n22855), .B(n22856), .Z(n22854) );
  NANDN U22961 ( .A(n22856), .B(n22855), .Z(n22851) );
  ANDN U22962 ( .B(B[223]), .A(n78), .Z(n22635) );
  XNOR U22963 ( .A(n22643), .B(n22857), .Z(n22636) );
  XNOR U22964 ( .A(n22642), .B(n22640), .Z(n22857) );
  AND U22965 ( .A(n22858), .B(n22859), .Z(n22640) );
  NANDN U22966 ( .A(n22860), .B(n22861), .Z(n22859) );
  OR U22967 ( .A(n22862), .B(n22863), .Z(n22861) );
  NAND U22968 ( .A(n22863), .B(n22862), .Z(n22858) );
  ANDN U22969 ( .B(B[224]), .A(n79), .Z(n22642) );
  XNOR U22970 ( .A(n22650), .B(n22864), .Z(n22643) );
  XNOR U22971 ( .A(n22649), .B(n22647), .Z(n22864) );
  AND U22972 ( .A(n22865), .B(n22866), .Z(n22647) );
  NANDN U22973 ( .A(n22867), .B(n22868), .Z(n22866) );
  NANDN U22974 ( .A(n22869), .B(n22870), .Z(n22868) );
  NANDN U22975 ( .A(n22870), .B(n22869), .Z(n22865) );
  ANDN U22976 ( .B(B[225]), .A(n80), .Z(n22649) );
  XNOR U22977 ( .A(n22657), .B(n22871), .Z(n22650) );
  XNOR U22978 ( .A(n22656), .B(n22654), .Z(n22871) );
  AND U22979 ( .A(n22872), .B(n22873), .Z(n22654) );
  NANDN U22980 ( .A(n22874), .B(n22875), .Z(n22873) );
  OR U22981 ( .A(n22876), .B(n22877), .Z(n22875) );
  NAND U22982 ( .A(n22877), .B(n22876), .Z(n22872) );
  ANDN U22983 ( .B(B[226]), .A(n81), .Z(n22656) );
  XNOR U22984 ( .A(n22664), .B(n22878), .Z(n22657) );
  XNOR U22985 ( .A(n22663), .B(n22661), .Z(n22878) );
  AND U22986 ( .A(n22879), .B(n22880), .Z(n22661) );
  NANDN U22987 ( .A(n22881), .B(n22882), .Z(n22880) );
  NAND U22988 ( .A(n22883), .B(n22884), .Z(n22882) );
  ANDN U22989 ( .B(B[227]), .A(n82), .Z(n22663) );
  XOR U22990 ( .A(n22670), .B(n22885), .Z(n22664) );
  XNOR U22991 ( .A(n22668), .B(n22671), .Z(n22885) );
  NAND U22992 ( .A(A[2]), .B(B[228]), .Z(n22671) );
  NANDN U22993 ( .A(n22886), .B(n22887), .Z(n22668) );
  AND U22994 ( .A(A[0]), .B(B[229]), .Z(n22887) );
  XNOR U22995 ( .A(n22673), .B(n22888), .Z(n22670) );
  NAND U22996 ( .A(A[0]), .B(B[230]), .Z(n22888) );
  NAND U22997 ( .A(B[229]), .B(A[1]), .Z(n22673) );
  NAND U22998 ( .A(n22889), .B(n22890), .Z(n336) );
  NANDN U22999 ( .A(n22891), .B(n22892), .Z(n22890) );
  OR U23000 ( .A(n22893), .B(n22894), .Z(n22892) );
  NAND U23001 ( .A(n22894), .B(n22893), .Z(n22889) );
  XOR U23002 ( .A(n338), .B(n337), .Z(\A1[227] ) );
  XOR U23003 ( .A(n22894), .B(n22895), .Z(n337) );
  XNOR U23004 ( .A(n22893), .B(n22891), .Z(n22895) );
  AND U23005 ( .A(n22896), .B(n22897), .Z(n22891) );
  NANDN U23006 ( .A(n22898), .B(n22899), .Z(n22897) );
  NANDN U23007 ( .A(n22900), .B(n22901), .Z(n22899) );
  NANDN U23008 ( .A(n22901), .B(n22900), .Z(n22896) );
  ANDN U23009 ( .B(B[198]), .A(n54), .Z(n22893) );
  XNOR U23010 ( .A(n22688), .B(n22902), .Z(n22894) );
  XNOR U23011 ( .A(n22687), .B(n22685), .Z(n22902) );
  AND U23012 ( .A(n22903), .B(n22904), .Z(n22685) );
  NANDN U23013 ( .A(n22905), .B(n22906), .Z(n22904) );
  OR U23014 ( .A(n22907), .B(n22908), .Z(n22906) );
  NAND U23015 ( .A(n22908), .B(n22907), .Z(n22903) );
  ANDN U23016 ( .B(B[199]), .A(n55), .Z(n22687) );
  XNOR U23017 ( .A(n22695), .B(n22909), .Z(n22688) );
  XNOR U23018 ( .A(n22694), .B(n22692), .Z(n22909) );
  AND U23019 ( .A(n22910), .B(n22911), .Z(n22692) );
  NANDN U23020 ( .A(n22912), .B(n22913), .Z(n22911) );
  NANDN U23021 ( .A(n22914), .B(n22915), .Z(n22913) );
  NANDN U23022 ( .A(n22915), .B(n22914), .Z(n22910) );
  ANDN U23023 ( .B(B[200]), .A(n56), .Z(n22694) );
  XNOR U23024 ( .A(n22702), .B(n22916), .Z(n22695) );
  XNOR U23025 ( .A(n22701), .B(n22699), .Z(n22916) );
  AND U23026 ( .A(n22917), .B(n22918), .Z(n22699) );
  NANDN U23027 ( .A(n22919), .B(n22920), .Z(n22918) );
  OR U23028 ( .A(n22921), .B(n22922), .Z(n22920) );
  NAND U23029 ( .A(n22922), .B(n22921), .Z(n22917) );
  ANDN U23030 ( .B(B[201]), .A(n57), .Z(n22701) );
  XNOR U23031 ( .A(n22709), .B(n22923), .Z(n22702) );
  XNOR U23032 ( .A(n22708), .B(n22706), .Z(n22923) );
  AND U23033 ( .A(n22924), .B(n22925), .Z(n22706) );
  NANDN U23034 ( .A(n22926), .B(n22927), .Z(n22925) );
  NANDN U23035 ( .A(n22928), .B(n22929), .Z(n22927) );
  NANDN U23036 ( .A(n22929), .B(n22928), .Z(n22924) );
  ANDN U23037 ( .B(B[202]), .A(n58), .Z(n22708) );
  XNOR U23038 ( .A(n22716), .B(n22930), .Z(n22709) );
  XNOR U23039 ( .A(n22715), .B(n22713), .Z(n22930) );
  AND U23040 ( .A(n22931), .B(n22932), .Z(n22713) );
  NANDN U23041 ( .A(n22933), .B(n22934), .Z(n22932) );
  OR U23042 ( .A(n22935), .B(n22936), .Z(n22934) );
  NAND U23043 ( .A(n22936), .B(n22935), .Z(n22931) );
  ANDN U23044 ( .B(B[203]), .A(n59), .Z(n22715) );
  XNOR U23045 ( .A(n22723), .B(n22937), .Z(n22716) );
  XNOR U23046 ( .A(n22722), .B(n22720), .Z(n22937) );
  AND U23047 ( .A(n22938), .B(n22939), .Z(n22720) );
  NANDN U23048 ( .A(n22940), .B(n22941), .Z(n22939) );
  NANDN U23049 ( .A(n22942), .B(n22943), .Z(n22941) );
  NANDN U23050 ( .A(n22943), .B(n22942), .Z(n22938) );
  ANDN U23051 ( .B(B[204]), .A(n60), .Z(n22722) );
  XNOR U23052 ( .A(n22730), .B(n22944), .Z(n22723) );
  XNOR U23053 ( .A(n22729), .B(n22727), .Z(n22944) );
  AND U23054 ( .A(n22945), .B(n22946), .Z(n22727) );
  NANDN U23055 ( .A(n22947), .B(n22948), .Z(n22946) );
  OR U23056 ( .A(n22949), .B(n22950), .Z(n22948) );
  NAND U23057 ( .A(n22950), .B(n22949), .Z(n22945) );
  ANDN U23058 ( .B(B[205]), .A(n61), .Z(n22729) );
  XNOR U23059 ( .A(n22737), .B(n22951), .Z(n22730) );
  XNOR U23060 ( .A(n22736), .B(n22734), .Z(n22951) );
  AND U23061 ( .A(n22952), .B(n22953), .Z(n22734) );
  NANDN U23062 ( .A(n22954), .B(n22955), .Z(n22953) );
  NANDN U23063 ( .A(n22956), .B(n22957), .Z(n22955) );
  NANDN U23064 ( .A(n22957), .B(n22956), .Z(n22952) );
  ANDN U23065 ( .B(B[206]), .A(n62), .Z(n22736) );
  XNOR U23066 ( .A(n22744), .B(n22958), .Z(n22737) );
  XNOR U23067 ( .A(n22743), .B(n22741), .Z(n22958) );
  AND U23068 ( .A(n22959), .B(n22960), .Z(n22741) );
  NANDN U23069 ( .A(n22961), .B(n22962), .Z(n22960) );
  OR U23070 ( .A(n22963), .B(n22964), .Z(n22962) );
  NAND U23071 ( .A(n22964), .B(n22963), .Z(n22959) );
  ANDN U23072 ( .B(B[207]), .A(n63), .Z(n22743) );
  XNOR U23073 ( .A(n22751), .B(n22965), .Z(n22744) );
  XNOR U23074 ( .A(n22750), .B(n22748), .Z(n22965) );
  AND U23075 ( .A(n22966), .B(n22967), .Z(n22748) );
  NANDN U23076 ( .A(n22968), .B(n22969), .Z(n22967) );
  NANDN U23077 ( .A(n22970), .B(n22971), .Z(n22969) );
  NANDN U23078 ( .A(n22971), .B(n22970), .Z(n22966) );
  ANDN U23079 ( .B(B[208]), .A(n64), .Z(n22750) );
  XNOR U23080 ( .A(n22758), .B(n22972), .Z(n22751) );
  XNOR U23081 ( .A(n22757), .B(n22755), .Z(n22972) );
  AND U23082 ( .A(n22973), .B(n22974), .Z(n22755) );
  NANDN U23083 ( .A(n22975), .B(n22976), .Z(n22974) );
  OR U23084 ( .A(n22977), .B(n22978), .Z(n22976) );
  NAND U23085 ( .A(n22978), .B(n22977), .Z(n22973) );
  ANDN U23086 ( .B(B[209]), .A(n65), .Z(n22757) );
  XNOR U23087 ( .A(n22765), .B(n22979), .Z(n22758) );
  XNOR U23088 ( .A(n22764), .B(n22762), .Z(n22979) );
  AND U23089 ( .A(n22980), .B(n22981), .Z(n22762) );
  NANDN U23090 ( .A(n22982), .B(n22983), .Z(n22981) );
  NANDN U23091 ( .A(n22984), .B(n22985), .Z(n22983) );
  NANDN U23092 ( .A(n22985), .B(n22984), .Z(n22980) );
  ANDN U23093 ( .B(B[210]), .A(n66), .Z(n22764) );
  XNOR U23094 ( .A(n22772), .B(n22986), .Z(n22765) );
  XNOR U23095 ( .A(n22771), .B(n22769), .Z(n22986) );
  AND U23096 ( .A(n22987), .B(n22988), .Z(n22769) );
  NANDN U23097 ( .A(n22989), .B(n22990), .Z(n22988) );
  OR U23098 ( .A(n22991), .B(n22992), .Z(n22990) );
  NAND U23099 ( .A(n22992), .B(n22991), .Z(n22987) );
  ANDN U23100 ( .B(B[211]), .A(n67), .Z(n22771) );
  XNOR U23101 ( .A(n22779), .B(n22993), .Z(n22772) );
  XNOR U23102 ( .A(n22778), .B(n22776), .Z(n22993) );
  AND U23103 ( .A(n22994), .B(n22995), .Z(n22776) );
  NANDN U23104 ( .A(n22996), .B(n22997), .Z(n22995) );
  NANDN U23105 ( .A(n22998), .B(n22999), .Z(n22997) );
  NANDN U23106 ( .A(n22999), .B(n22998), .Z(n22994) );
  ANDN U23107 ( .B(B[212]), .A(n68), .Z(n22778) );
  XNOR U23108 ( .A(n22786), .B(n23000), .Z(n22779) );
  XNOR U23109 ( .A(n22785), .B(n22783), .Z(n23000) );
  AND U23110 ( .A(n23001), .B(n23002), .Z(n22783) );
  NANDN U23111 ( .A(n23003), .B(n23004), .Z(n23002) );
  OR U23112 ( .A(n23005), .B(n23006), .Z(n23004) );
  NAND U23113 ( .A(n23006), .B(n23005), .Z(n23001) );
  ANDN U23114 ( .B(B[213]), .A(n69), .Z(n22785) );
  XNOR U23115 ( .A(n22793), .B(n23007), .Z(n22786) );
  XNOR U23116 ( .A(n22792), .B(n22790), .Z(n23007) );
  AND U23117 ( .A(n23008), .B(n23009), .Z(n22790) );
  NANDN U23118 ( .A(n23010), .B(n23011), .Z(n23009) );
  NANDN U23119 ( .A(n23012), .B(n23013), .Z(n23011) );
  NANDN U23120 ( .A(n23013), .B(n23012), .Z(n23008) );
  ANDN U23121 ( .B(B[214]), .A(n70), .Z(n22792) );
  XNOR U23122 ( .A(n22800), .B(n23014), .Z(n22793) );
  XNOR U23123 ( .A(n22799), .B(n22797), .Z(n23014) );
  AND U23124 ( .A(n23015), .B(n23016), .Z(n22797) );
  NANDN U23125 ( .A(n23017), .B(n23018), .Z(n23016) );
  OR U23126 ( .A(n23019), .B(n23020), .Z(n23018) );
  NAND U23127 ( .A(n23020), .B(n23019), .Z(n23015) );
  ANDN U23128 ( .B(B[215]), .A(n71), .Z(n22799) );
  XNOR U23129 ( .A(n22807), .B(n23021), .Z(n22800) );
  XNOR U23130 ( .A(n22806), .B(n22804), .Z(n23021) );
  AND U23131 ( .A(n23022), .B(n23023), .Z(n22804) );
  NANDN U23132 ( .A(n23024), .B(n23025), .Z(n23023) );
  NANDN U23133 ( .A(n23026), .B(n23027), .Z(n23025) );
  NANDN U23134 ( .A(n23027), .B(n23026), .Z(n23022) );
  ANDN U23135 ( .B(B[216]), .A(n72), .Z(n22806) );
  XNOR U23136 ( .A(n22814), .B(n23028), .Z(n22807) );
  XNOR U23137 ( .A(n22813), .B(n22811), .Z(n23028) );
  AND U23138 ( .A(n23029), .B(n23030), .Z(n22811) );
  NANDN U23139 ( .A(n23031), .B(n23032), .Z(n23030) );
  OR U23140 ( .A(n23033), .B(n23034), .Z(n23032) );
  NAND U23141 ( .A(n23034), .B(n23033), .Z(n23029) );
  ANDN U23142 ( .B(B[217]), .A(n73), .Z(n22813) );
  XNOR U23143 ( .A(n22821), .B(n23035), .Z(n22814) );
  XNOR U23144 ( .A(n22820), .B(n22818), .Z(n23035) );
  AND U23145 ( .A(n23036), .B(n23037), .Z(n22818) );
  NANDN U23146 ( .A(n23038), .B(n23039), .Z(n23037) );
  NANDN U23147 ( .A(n23040), .B(n23041), .Z(n23039) );
  NANDN U23148 ( .A(n23041), .B(n23040), .Z(n23036) );
  ANDN U23149 ( .B(B[218]), .A(n74), .Z(n22820) );
  XNOR U23150 ( .A(n22828), .B(n23042), .Z(n22821) );
  XNOR U23151 ( .A(n22827), .B(n22825), .Z(n23042) );
  AND U23152 ( .A(n23043), .B(n23044), .Z(n22825) );
  NANDN U23153 ( .A(n23045), .B(n23046), .Z(n23044) );
  OR U23154 ( .A(n23047), .B(n23048), .Z(n23046) );
  NAND U23155 ( .A(n23048), .B(n23047), .Z(n23043) );
  ANDN U23156 ( .B(B[219]), .A(n75), .Z(n22827) );
  XNOR U23157 ( .A(n22835), .B(n23049), .Z(n22828) );
  XNOR U23158 ( .A(n22834), .B(n22832), .Z(n23049) );
  AND U23159 ( .A(n23050), .B(n23051), .Z(n22832) );
  NANDN U23160 ( .A(n23052), .B(n23053), .Z(n23051) );
  NANDN U23161 ( .A(n23054), .B(n23055), .Z(n23053) );
  NANDN U23162 ( .A(n23055), .B(n23054), .Z(n23050) );
  ANDN U23163 ( .B(B[220]), .A(n76), .Z(n22834) );
  XNOR U23164 ( .A(n22842), .B(n23056), .Z(n22835) );
  XNOR U23165 ( .A(n22841), .B(n22839), .Z(n23056) );
  AND U23166 ( .A(n23057), .B(n23058), .Z(n22839) );
  NANDN U23167 ( .A(n23059), .B(n23060), .Z(n23058) );
  OR U23168 ( .A(n23061), .B(n23062), .Z(n23060) );
  NAND U23169 ( .A(n23062), .B(n23061), .Z(n23057) );
  ANDN U23170 ( .B(B[221]), .A(n77), .Z(n22841) );
  XNOR U23171 ( .A(n22849), .B(n23063), .Z(n22842) );
  XNOR U23172 ( .A(n22848), .B(n22846), .Z(n23063) );
  AND U23173 ( .A(n23064), .B(n23065), .Z(n22846) );
  NANDN U23174 ( .A(n23066), .B(n23067), .Z(n23065) );
  NANDN U23175 ( .A(n23068), .B(n23069), .Z(n23067) );
  NANDN U23176 ( .A(n23069), .B(n23068), .Z(n23064) );
  ANDN U23177 ( .B(B[222]), .A(n78), .Z(n22848) );
  XNOR U23178 ( .A(n22856), .B(n23070), .Z(n22849) );
  XNOR U23179 ( .A(n22855), .B(n22853), .Z(n23070) );
  AND U23180 ( .A(n23071), .B(n23072), .Z(n22853) );
  NANDN U23181 ( .A(n23073), .B(n23074), .Z(n23072) );
  OR U23182 ( .A(n23075), .B(n23076), .Z(n23074) );
  NAND U23183 ( .A(n23076), .B(n23075), .Z(n23071) );
  ANDN U23184 ( .B(B[223]), .A(n79), .Z(n22855) );
  XNOR U23185 ( .A(n22863), .B(n23077), .Z(n22856) );
  XNOR U23186 ( .A(n22862), .B(n22860), .Z(n23077) );
  AND U23187 ( .A(n23078), .B(n23079), .Z(n22860) );
  NANDN U23188 ( .A(n23080), .B(n23081), .Z(n23079) );
  NANDN U23189 ( .A(n23082), .B(n23083), .Z(n23081) );
  NANDN U23190 ( .A(n23083), .B(n23082), .Z(n23078) );
  ANDN U23191 ( .B(B[224]), .A(n80), .Z(n22862) );
  XNOR U23192 ( .A(n22870), .B(n23084), .Z(n22863) );
  XNOR U23193 ( .A(n22869), .B(n22867), .Z(n23084) );
  AND U23194 ( .A(n23085), .B(n23086), .Z(n22867) );
  NANDN U23195 ( .A(n23087), .B(n23088), .Z(n23086) );
  OR U23196 ( .A(n23089), .B(n23090), .Z(n23088) );
  NAND U23197 ( .A(n23090), .B(n23089), .Z(n23085) );
  ANDN U23198 ( .B(B[225]), .A(n81), .Z(n22869) );
  XNOR U23199 ( .A(n22877), .B(n23091), .Z(n22870) );
  XNOR U23200 ( .A(n22876), .B(n22874), .Z(n23091) );
  AND U23201 ( .A(n23092), .B(n23093), .Z(n22874) );
  NANDN U23202 ( .A(n23094), .B(n23095), .Z(n23093) );
  NAND U23203 ( .A(n23096), .B(n23097), .Z(n23095) );
  ANDN U23204 ( .B(B[226]), .A(n82), .Z(n22876) );
  XOR U23205 ( .A(n22883), .B(n23098), .Z(n22877) );
  XNOR U23206 ( .A(n22881), .B(n22884), .Z(n23098) );
  NAND U23207 ( .A(A[2]), .B(B[227]), .Z(n22884) );
  NANDN U23208 ( .A(n23099), .B(n23100), .Z(n22881) );
  AND U23209 ( .A(A[0]), .B(B[228]), .Z(n23100) );
  XNOR U23210 ( .A(n22886), .B(n23101), .Z(n22883) );
  NAND U23211 ( .A(A[0]), .B(B[229]), .Z(n23101) );
  NAND U23212 ( .A(B[228]), .B(A[1]), .Z(n22886) );
  NAND U23213 ( .A(n23102), .B(n23103), .Z(n338) );
  NANDN U23214 ( .A(n23104), .B(n23105), .Z(n23103) );
  OR U23215 ( .A(n23106), .B(n23107), .Z(n23105) );
  NAND U23216 ( .A(n23107), .B(n23106), .Z(n23102) );
  XOR U23217 ( .A(n340), .B(n339), .Z(\A1[226] ) );
  XOR U23218 ( .A(n23107), .B(n23108), .Z(n339) );
  XNOR U23219 ( .A(n23106), .B(n23104), .Z(n23108) );
  AND U23220 ( .A(n23109), .B(n23110), .Z(n23104) );
  NANDN U23221 ( .A(n23111), .B(n23112), .Z(n23110) );
  NANDN U23222 ( .A(n23113), .B(n23114), .Z(n23112) );
  NANDN U23223 ( .A(n23114), .B(n23113), .Z(n23109) );
  ANDN U23224 ( .B(B[197]), .A(n54), .Z(n23106) );
  XNOR U23225 ( .A(n22901), .B(n23115), .Z(n23107) );
  XNOR U23226 ( .A(n22900), .B(n22898), .Z(n23115) );
  AND U23227 ( .A(n23116), .B(n23117), .Z(n22898) );
  NANDN U23228 ( .A(n23118), .B(n23119), .Z(n23117) );
  OR U23229 ( .A(n23120), .B(n23121), .Z(n23119) );
  NAND U23230 ( .A(n23121), .B(n23120), .Z(n23116) );
  ANDN U23231 ( .B(B[198]), .A(n55), .Z(n22900) );
  XNOR U23232 ( .A(n22908), .B(n23122), .Z(n22901) );
  XNOR U23233 ( .A(n22907), .B(n22905), .Z(n23122) );
  AND U23234 ( .A(n23123), .B(n23124), .Z(n22905) );
  NANDN U23235 ( .A(n23125), .B(n23126), .Z(n23124) );
  NANDN U23236 ( .A(n23127), .B(n23128), .Z(n23126) );
  NANDN U23237 ( .A(n23128), .B(n23127), .Z(n23123) );
  ANDN U23238 ( .B(B[199]), .A(n56), .Z(n22907) );
  XNOR U23239 ( .A(n22915), .B(n23129), .Z(n22908) );
  XNOR U23240 ( .A(n22914), .B(n22912), .Z(n23129) );
  AND U23241 ( .A(n23130), .B(n23131), .Z(n22912) );
  NANDN U23242 ( .A(n23132), .B(n23133), .Z(n23131) );
  OR U23243 ( .A(n23134), .B(n23135), .Z(n23133) );
  NAND U23244 ( .A(n23135), .B(n23134), .Z(n23130) );
  ANDN U23245 ( .B(B[200]), .A(n57), .Z(n22914) );
  XNOR U23246 ( .A(n22922), .B(n23136), .Z(n22915) );
  XNOR U23247 ( .A(n22921), .B(n22919), .Z(n23136) );
  AND U23248 ( .A(n23137), .B(n23138), .Z(n22919) );
  NANDN U23249 ( .A(n23139), .B(n23140), .Z(n23138) );
  NANDN U23250 ( .A(n23141), .B(n23142), .Z(n23140) );
  NANDN U23251 ( .A(n23142), .B(n23141), .Z(n23137) );
  ANDN U23252 ( .B(B[201]), .A(n58), .Z(n22921) );
  XNOR U23253 ( .A(n22929), .B(n23143), .Z(n22922) );
  XNOR U23254 ( .A(n22928), .B(n22926), .Z(n23143) );
  AND U23255 ( .A(n23144), .B(n23145), .Z(n22926) );
  NANDN U23256 ( .A(n23146), .B(n23147), .Z(n23145) );
  OR U23257 ( .A(n23148), .B(n23149), .Z(n23147) );
  NAND U23258 ( .A(n23149), .B(n23148), .Z(n23144) );
  ANDN U23259 ( .B(B[202]), .A(n59), .Z(n22928) );
  XNOR U23260 ( .A(n22936), .B(n23150), .Z(n22929) );
  XNOR U23261 ( .A(n22935), .B(n22933), .Z(n23150) );
  AND U23262 ( .A(n23151), .B(n23152), .Z(n22933) );
  NANDN U23263 ( .A(n23153), .B(n23154), .Z(n23152) );
  NANDN U23264 ( .A(n23155), .B(n23156), .Z(n23154) );
  NANDN U23265 ( .A(n23156), .B(n23155), .Z(n23151) );
  ANDN U23266 ( .B(B[203]), .A(n60), .Z(n22935) );
  XNOR U23267 ( .A(n22943), .B(n23157), .Z(n22936) );
  XNOR U23268 ( .A(n22942), .B(n22940), .Z(n23157) );
  AND U23269 ( .A(n23158), .B(n23159), .Z(n22940) );
  NANDN U23270 ( .A(n23160), .B(n23161), .Z(n23159) );
  OR U23271 ( .A(n23162), .B(n23163), .Z(n23161) );
  NAND U23272 ( .A(n23163), .B(n23162), .Z(n23158) );
  ANDN U23273 ( .B(B[204]), .A(n61), .Z(n22942) );
  XNOR U23274 ( .A(n22950), .B(n23164), .Z(n22943) );
  XNOR U23275 ( .A(n22949), .B(n22947), .Z(n23164) );
  AND U23276 ( .A(n23165), .B(n23166), .Z(n22947) );
  NANDN U23277 ( .A(n23167), .B(n23168), .Z(n23166) );
  NANDN U23278 ( .A(n23169), .B(n23170), .Z(n23168) );
  NANDN U23279 ( .A(n23170), .B(n23169), .Z(n23165) );
  ANDN U23280 ( .B(B[205]), .A(n62), .Z(n22949) );
  XNOR U23281 ( .A(n22957), .B(n23171), .Z(n22950) );
  XNOR U23282 ( .A(n22956), .B(n22954), .Z(n23171) );
  AND U23283 ( .A(n23172), .B(n23173), .Z(n22954) );
  NANDN U23284 ( .A(n23174), .B(n23175), .Z(n23173) );
  OR U23285 ( .A(n23176), .B(n23177), .Z(n23175) );
  NAND U23286 ( .A(n23177), .B(n23176), .Z(n23172) );
  ANDN U23287 ( .B(B[206]), .A(n63), .Z(n22956) );
  XNOR U23288 ( .A(n22964), .B(n23178), .Z(n22957) );
  XNOR U23289 ( .A(n22963), .B(n22961), .Z(n23178) );
  AND U23290 ( .A(n23179), .B(n23180), .Z(n22961) );
  NANDN U23291 ( .A(n23181), .B(n23182), .Z(n23180) );
  NANDN U23292 ( .A(n23183), .B(n23184), .Z(n23182) );
  NANDN U23293 ( .A(n23184), .B(n23183), .Z(n23179) );
  ANDN U23294 ( .B(B[207]), .A(n64), .Z(n22963) );
  XNOR U23295 ( .A(n22971), .B(n23185), .Z(n22964) );
  XNOR U23296 ( .A(n22970), .B(n22968), .Z(n23185) );
  AND U23297 ( .A(n23186), .B(n23187), .Z(n22968) );
  NANDN U23298 ( .A(n23188), .B(n23189), .Z(n23187) );
  OR U23299 ( .A(n23190), .B(n23191), .Z(n23189) );
  NAND U23300 ( .A(n23191), .B(n23190), .Z(n23186) );
  ANDN U23301 ( .B(B[208]), .A(n65), .Z(n22970) );
  XNOR U23302 ( .A(n22978), .B(n23192), .Z(n22971) );
  XNOR U23303 ( .A(n22977), .B(n22975), .Z(n23192) );
  AND U23304 ( .A(n23193), .B(n23194), .Z(n22975) );
  NANDN U23305 ( .A(n23195), .B(n23196), .Z(n23194) );
  NANDN U23306 ( .A(n23197), .B(n23198), .Z(n23196) );
  NANDN U23307 ( .A(n23198), .B(n23197), .Z(n23193) );
  ANDN U23308 ( .B(B[209]), .A(n66), .Z(n22977) );
  XNOR U23309 ( .A(n22985), .B(n23199), .Z(n22978) );
  XNOR U23310 ( .A(n22984), .B(n22982), .Z(n23199) );
  AND U23311 ( .A(n23200), .B(n23201), .Z(n22982) );
  NANDN U23312 ( .A(n23202), .B(n23203), .Z(n23201) );
  OR U23313 ( .A(n23204), .B(n23205), .Z(n23203) );
  NAND U23314 ( .A(n23205), .B(n23204), .Z(n23200) );
  ANDN U23315 ( .B(B[210]), .A(n67), .Z(n22984) );
  XNOR U23316 ( .A(n22992), .B(n23206), .Z(n22985) );
  XNOR U23317 ( .A(n22991), .B(n22989), .Z(n23206) );
  AND U23318 ( .A(n23207), .B(n23208), .Z(n22989) );
  NANDN U23319 ( .A(n23209), .B(n23210), .Z(n23208) );
  NANDN U23320 ( .A(n23211), .B(n23212), .Z(n23210) );
  NANDN U23321 ( .A(n23212), .B(n23211), .Z(n23207) );
  ANDN U23322 ( .B(B[211]), .A(n68), .Z(n22991) );
  XNOR U23323 ( .A(n22999), .B(n23213), .Z(n22992) );
  XNOR U23324 ( .A(n22998), .B(n22996), .Z(n23213) );
  AND U23325 ( .A(n23214), .B(n23215), .Z(n22996) );
  NANDN U23326 ( .A(n23216), .B(n23217), .Z(n23215) );
  OR U23327 ( .A(n23218), .B(n23219), .Z(n23217) );
  NAND U23328 ( .A(n23219), .B(n23218), .Z(n23214) );
  ANDN U23329 ( .B(B[212]), .A(n69), .Z(n22998) );
  XNOR U23330 ( .A(n23006), .B(n23220), .Z(n22999) );
  XNOR U23331 ( .A(n23005), .B(n23003), .Z(n23220) );
  AND U23332 ( .A(n23221), .B(n23222), .Z(n23003) );
  NANDN U23333 ( .A(n23223), .B(n23224), .Z(n23222) );
  NANDN U23334 ( .A(n23225), .B(n23226), .Z(n23224) );
  NANDN U23335 ( .A(n23226), .B(n23225), .Z(n23221) );
  ANDN U23336 ( .B(B[213]), .A(n70), .Z(n23005) );
  XNOR U23337 ( .A(n23013), .B(n23227), .Z(n23006) );
  XNOR U23338 ( .A(n23012), .B(n23010), .Z(n23227) );
  AND U23339 ( .A(n23228), .B(n23229), .Z(n23010) );
  NANDN U23340 ( .A(n23230), .B(n23231), .Z(n23229) );
  OR U23341 ( .A(n23232), .B(n23233), .Z(n23231) );
  NAND U23342 ( .A(n23233), .B(n23232), .Z(n23228) );
  ANDN U23343 ( .B(B[214]), .A(n71), .Z(n23012) );
  XNOR U23344 ( .A(n23020), .B(n23234), .Z(n23013) );
  XNOR U23345 ( .A(n23019), .B(n23017), .Z(n23234) );
  AND U23346 ( .A(n23235), .B(n23236), .Z(n23017) );
  NANDN U23347 ( .A(n23237), .B(n23238), .Z(n23236) );
  NANDN U23348 ( .A(n23239), .B(n23240), .Z(n23238) );
  NANDN U23349 ( .A(n23240), .B(n23239), .Z(n23235) );
  ANDN U23350 ( .B(B[215]), .A(n72), .Z(n23019) );
  XNOR U23351 ( .A(n23027), .B(n23241), .Z(n23020) );
  XNOR U23352 ( .A(n23026), .B(n23024), .Z(n23241) );
  AND U23353 ( .A(n23242), .B(n23243), .Z(n23024) );
  NANDN U23354 ( .A(n23244), .B(n23245), .Z(n23243) );
  OR U23355 ( .A(n23246), .B(n23247), .Z(n23245) );
  NAND U23356 ( .A(n23247), .B(n23246), .Z(n23242) );
  ANDN U23357 ( .B(B[216]), .A(n73), .Z(n23026) );
  XNOR U23358 ( .A(n23034), .B(n23248), .Z(n23027) );
  XNOR U23359 ( .A(n23033), .B(n23031), .Z(n23248) );
  AND U23360 ( .A(n23249), .B(n23250), .Z(n23031) );
  NANDN U23361 ( .A(n23251), .B(n23252), .Z(n23250) );
  NANDN U23362 ( .A(n23253), .B(n23254), .Z(n23252) );
  NANDN U23363 ( .A(n23254), .B(n23253), .Z(n23249) );
  ANDN U23364 ( .B(B[217]), .A(n74), .Z(n23033) );
  XNOR U23365 ( .A(n23041), .B(n23255), .Z(n23034) );
  XNOR U23366 ( .A(n23040), .B(n23038), .Z(n23255) );
  AND U23367 ( .A(n23256), .B(n23257), .Z(n23038) );
  NANDN U23368 ( .A(n23258), .B(n23259), .Z(n23257) );
  OR U23369 ( .A(n23260), .B(n23261), .Z(n23259) );
  NAND U23370 ( .A(n23261), .B(n23260), .Z(n23256) );
  ANDN U23371 ( .B(B[218]), .A(n75), .Z(n23040) );
  XNOR U23372 ( .A(n23048), .B(n23262), .Z(n23041) );
  XNOR U23373 ( .A(n23047), .B(n23045), .Z(n23262) );
  AND U23374 ( .A(n23263), .B(n23264), .Z(n23045) );
  NANDN U23375 ( .A(n23265), .B(n23266), .Z(n23264) );
  NANDN U23376 ( .A(n23267), .B(n23268), .Z(n23266) );
  NANDN U23377 ( .A(n23268), .B(n23267), .Z(n23263) );
  ANDN U23378 ( .B(B[219]), .A(n76), .Z(n23047) );
  XNOR U23379 ( .A(n23055), .B(n23269), .Z(n23048) );
  XNOR U23380 ( .A(n23054), .B(n23052), .Z(n23269) );
  AND U23381 ( .A(n23270), .B(n23271), .Z(n23052) );
  NANDN U23382 ( .A(n23272), .B(n23273), .Z(n23271) );
  OR U23383 ( .A(n23274), .B(n23275), .Z(n23273) );
  NAND U23384 ( .A(n23275), .B(n23274), .Z(n23270) );
  ANDN U23385 ( .B(B[220]), .A(n77), .Z(n23054) );
  XNOR U23386 ( .A(n23062), .B(n23276), .Z(n23055) );
  XNOR U23387 ( .A(n23061), .B(n23059), .Z(n23276) );
  AND U23388 ( .A(n23277), .B(n23278), .Z(n23059) );
  NANDN U23389 ( .A(n23279), .B(n23280), .Z(n23278) );
  NANDN U23390 ( .A(n23281), .B(n23282), .Z(n23280) );
  NANDN U23391 ( .A(n23282), .B(n23281), .Z(n23277) );
  ANDN U23392 ( .B(B[221]), .A(n78), .Z(n23061) );
  XNOR U23393 ( .A(n23069), .B(n23283), .Z(n23062) );
  XNOR U23394 ( .A(n23068), .B(n23066), .Z(n23283) );
  AND U23395 ( .A(n23284), .B(n23285), .Z(n23066) );
  NANDN U23396 ( .A(n23286), .B(n23287), .Z(n23285) );
  OR U23397 ( .A(n23288), .B(n23289), .Z(n23287) );
  NAND U23398 ( .A(n23289), .B(n23288), .Z(n23284) );
  ANDN U23399 ( .B(B[222]), .A(n79), .Z(n23068) );
  XNOR U23400 ( .A(n23076), .B(n23290), .Z(n23069) );
  XNOR U23401 ( .A(n23075), .B(n23073), .Z(n23290) );
  AND U23402 ( .A(n23291), .B(n23292), .Z(n23073) );
  NANDN U23403 ( .A(n23293), .B(n23294), .Z(n23292) );
  NANDN U23404 ( .A(n23295), .B(n23296), .Z(n23294) );
  NANDN U23405 ( .A(n23296), .B(n23295), .Z(n23291) );
  ANDN U23406 ( .B(B[223]), .A(n80), .Z(n23075) );
  XNOR U23407 ( .A(n23083), .B(n23297), .Z(n23076) );
  XNOR U23408 ( .A(n23082), .B(n23080), .Z(n23297) );
  AND U23409 ( .A(n23298), .B(n23299), .Z(n23080) );
  NANDN U23410 ( .A(n23300), .B(n23301), .Z(n23299) );
  OR U23411 ( .A(n23302), .B(n23303), .Z(n23301) );
  NAND U23412 ( .A(n23303), .B(n23302), .Z(n23298) );
  ANDN U23413 ( .B(B[224]), .A(n81), .Z(n23082) );
  XNOR U23414 ( .A(n23090), .B(n23304), .Z(n23083) );
  XNOR U23415 ( .A(n23089), .B(n23087), .Z(n23304) );
  AND U23416 ( .A(n23305), .B(n23306), .Z(n23087) );
  NANDN U23417 ( .A(n23307), .B(n23308), .Z(n23306) );
  NAND U23418 ( .A(n23309), .B(n23310), .Z(n23308) );
  ANDN U23419 ( .B(B[225]), .A(n82), .Z(n23089) );
  XOR U23420 ( .A(n23096), .B(n23311), .Z(n23090) );
  XNOR U23421 ( .A(n23094), .B(n23097), .Z(n23311) );
  NAND U23422 ( .A(A[2]), .B(B[226]), .Z(n23097) );
  NANDN U23423 ( .A(n23312), .B(n23313), .Z(n23094) );
  AND U23424 ( .A(A[0]), .B(B[227]), .Z(n23313) );
  XNOR U23425 ( .A(n23099), .B(n23314), .Z(n23096) );
  NAND U23426 ( .A(A[0]), .B(B[228]), .Z(n23314) );
  NAND U23427 ( .A(B[227]), .B(A[1]), .Z(n23099) );
  NAND U23428 ( .A(n23315), .B(n23316), .Z(n340) );
  NANDN U23429 ( .A(n23317), .B(n23318), .Z(n23316) );
  OR U23430 ( .A(n23319), .B(n23320), .Z(n23318) );
  NAND U23431 ( .A(n23320), .B(n23319), .Z(n23315) );
  XOR U23432 ( .A(n342), .B(n341), .Z(\A1[225] ) );
  XOR U23433 ( .A(n23320), .B(n23321), .Z(n341) );
  XNOR U23434 ( .A(n23319), .B(n23317), .Z(n23321) );
  AND U23435 ( .A(n23322), .B(n23323), .Z(n23317) );
  NANDN U23436 ( .A(n23324), .B(n23325), .Z(n23323) );
  NANDN U23437 ( .A(n23326), .B(n23327), .Z(n23325) );
  NANDN U23438 ( .A(n23327), .B(n23326), .Z(n23322) );
  ANDN U23439 ( .B(B[196]), .A(n54), .Z(n23319) );
  XNOR U23440 ( .A(n23114), .B(n23328), .Z(n23320) );
  XNOR U23441 ( .A(n23113), .B(n23111), .Z(n23328) );
  AND U23442 ( .A(n23329), .B(n23330), .Z(n23111) );
  NANDN U23443 ( .A(n23331), .B(n23332), .Z(n23330) );
  OR U23444 ( .A(n23333), .B(n23334), .Z(n23332) );
  NAND U23445 ( .A(n23334), .B(n23333), .Z(n23329) );
  ANDN U23446 ( .B(B[197]), .A(n55), .Z(n23113) );
  XNOR U23447 ( .A(n23121), .B(n23335), .Z(n23114) );
  XNOR U23448 ( .A(n23120), .B(n23118), .Z(n23335) );
  AND U23449 ( .A(n23336), .B(n23337), .Z(n23118) );
  NANDN U23450 ( .A(n23338), .B(n23339), .Z(n23337) );
  NANDN U23451 ( .A(n23340), .B(n23341), .Z(n23339) );
  NANDN U23452 ( .A(n23341), .B(n23340), .Z(n23336) );
  ANDN U23453 ( .B(B[198]), .A(n56), .Z(n23120) );
  XNOR U23454 ( .A(n23128), .B(n23342), .Z(n23121) );
  XNOR U23455 ( .A(n23127), .B(n23125), .Z(n23342) );
  AND U23456 ( .A(n23343), .B(n23344), .Z(n23125) );
  NANDN U23457 ( .A(n23345), .B(n23346), .Z(n23344) );
  OR U23458 ( .A(n23347), .B(n23348), .Z(n23346) );
  NAND U23459 ( .A(n23348), .B(n23347), .Z(n23343) );
  ANDN U23460 ( .B(B[199]), .A(n57), .Z(n23127) );
  XNOR U23461 ( .A(n23135), .B(n23349), .Z(n23128) );
  XNOR U23462 ( .A(n23134), .B(n23132), .Z(n23349) );
  AND U23463 ( .A(n23350), .B(n23351), .Z(n23132) );
  NANDN U23464 ( .A(n23352), .B(n23353), .Z(n23351) );
  NANDN U23465 ( .A(n23354), .B(n23355), .Z(n23353) );
  NANDN U23466 ( .A(n23355), .B(n23354), .Z(n23350) );
  ANDN U23467 ( .B(B[200]), .A(n58), .Z(n23134) );
  XNOR U23468 ( .A(n23142), .B(n23356), .Z(n23135) );
  XNOR U23469 ( .A(n23141), .B(n23139), .Z(n23356) );
  AND U23470 ( .A(n23357), .B(n23358), .Z(n23139) );
  NANDN U23471 ( .A(n23359), .B(n23360), .Z(n23358) );
  OR U23472 ( .A(n23361), .B(n23362), .Z(n23360) );
  NAND U23473 ( .A(n23362), .B(n23361), .Z(n23357) );
  ANDN U23474 ( .B(B[201]), .A(n59), .Z(n23141) );
  XNOR U23475 ( .A(n23149), .B(n23363), .Z(n23142) );
  XNOR U23476 ( .A(n23148), .B(n23146), .Z(n23363) );
  AND U23477 ( .A(n23364), .B(n23365), .Z(n23146) );
  NANDN U23478 ( .A(n23366), .B(n23367), .Z(n23365) );
  NANDN U23479 ( .A(n23368), .B(n23369), .Z(n23367) );
  NANDN U23480 ( .A(n23369), .B(n23368), .Z(n23364) );
  ANDN U23481 ( .B(B[202]), .A(n60), .Z(n23148) );
  XNOR U23482 ( .A(n23156), .B(n23370), .Z(n23149) );
  XNOR U23483 ( .A(n23155), .B(n23153), .Z(n23370) );
  AND U23484 ( .A(n23371), .B(n23372), .Z(n23153) );
  NANDN U23485 ( .A(n23373), .B(n23374), .Z(n23372) );
  OR U23486 ( .A(n23375), .B(n23376), .Z(n23374) );
  NAND U23487 ( .A(n23376), .B(n23375), .Z(n23371) );
  ANDN U23488 ( .B(B[203]), .A(n61), .Z(n23155) );
  XNOR U23489 ( .A(n23163), .B(n23377), .Z(n23156) );
  XNOR U23490 ( .A(n23162), .B(n23160), .Z(n23377) );
  AND U23491 ( .A(n23378), .B(n23379), .Z(n23160) );
  NANDN U23492 ( .A(n23380), .B(n23381), .Z(n23379) );
  NANDN U23493 ( .A(n23382), .B(n23383), .Z(n23381) );
  NANDN U23494 ( .A(n23383), .B(n23382), .Z(n23378) );
  ANDN U23495 ( .B(B[204]), .A(n62), .Z(n23162) );
  XNOR U23496 ( .A(n23170), .B(n23384), .Z(n23163) );
  XNOR U23497 ( .A(n23169), .B(n23167), .Z(n23384) );
  AND U23498 ( .A(n23385), .B(n23386), .Z(n23167) );
  NANDN U23499 ( .A(n23387), .B(n23388), .Z(n23386) );
  OR U23500 ( .A(n23389), .B(n23390), .Z(n23388) );
  NAND U23501 ( .A(n23390), .B(n23389), .Z(n23385) );
  ANDN U23502 ( .B(B[205]), .A(n63), .Z(n23169) );
  XNOR U23503 ( .A(n23177), .B(n23391), .Z(n23170) );
  XNOR U23504 ( .A(n23176), .B(n23174), .Z(n23391) );
  AND U23505 ( .A(n23392), .B(n23393), .Z(n23174) );
  NANDN U23506 ( .A(n23394), .B(n23395), .Z(n23393) );
  NANDN U23507 ( .A(n23396), .B(n23397), .Z(n23395) );
  NANDN U23508 ( .A(n23397), .B(n23396), .Z(n23392) );
  ANDN U23509 ( .B(B[206]), .A(n64), .Z(n23176) );
  XNOR U23510 ( .A(n23184), .B(n23398), .Z(n23177) );
  XNOR U23511 ( .A(n23183), .B(n23181), .Z(n23398) );
  AND U23512 ( .A(n23399), .B(n23400), .Z(n23181) );
  NANDN U23513 ( .A(n23401), .B(n23402), .Z(n23400) );
  OR U23514 ( .A(n23403), .B(n23404), .Z(n23402) );
  NAND U23515 ( .A(n23404), .B(n23403), .Z(n23399) );
  ANDN U23516 ( .B(B[207]), .A(n65), .Z(n23183) );
  XNOR U23517 ( .A(n23191), .B(n23405), .Z(n23184) );
  XNOR U23518 ( .A(n23190), .B(n23188), .Z(n23405) );
  AND U23519 ( .A(n23406), .B(n23407), .Z(n23188) );
  NANDN U23520 ( .A(n23408), .B(n23409), .Z(n23407) );
  NANDN U23521 ( .A(n23410), .B(n23411), .Z(n23409) );
  NANDN U23522 ( .A(n23411), .B(n23410), .Z(n23406) );
  ANDN U23523 ( .B(B[208]), .A(n66), .Z(n23190) );
  XNOR U23524 ( .A(n23198), .B(n23412), .Z(n23191) );
  XNOR U23525 ( .A(n23197), .B(n23195), .Z(n23412) );
  AND U23526 ( .A(n23413), .B(n23414), .Z(n23195) );
  NANDN U23527 ( .A(n23415), .B(n23416), .Z(n23414) );
  OR U23528 ( .A(n23417), .B(n23418), .Z(n23416) );
  NAND U23529 ( .A(n23418), .B(n23417), .Z(n23413) );
  ANDN U23530 ( .B(B[209]), .A(n67), .Z(n23197) );
  XNOR U23531 ( .A(n23205), .B(n23419), .Z(n23198) );
  XNOR U23532 ( .A(n23204), .B(n23202), .Z(n23419) );
  AND U23533 ( .A(n23420), .B(n23421), .Z(n23202) );
  NANDN U23534 ( .A(n23422), .B(n23423), .Z(n23421) );
  NANDN U23535 ( .A(n23424), .B(n23425), .Z(n23423) );
  NANDN U23536 ( .A(n23425), .B(n23424), .Z(n23420) );
  ANDN U23537 ( .B(B[210]), .A(n68), .Z(n23204) );
  XNOR U23538 ( .A(n23212), .B(n23426), .Z(n23205) );
  XNOR U23539 ( .A(n23211), .B(n23209), .Z(n23426) );
  AND U23540 ( .A(n23427), .B(n23428), .Z(n23209) );
  NANDN U23541 ( .A(n23429), .B(n23430), .Z(n23428) );
  OR U23542 ( .A(n23431), .B(n23432), .Z(n23430) );
  NAND U23543 ( .A(n23432), .B(n23431), .Z(n23427) );
  ANDN U23544 ( .B(B[211]), .A(n69), .Z(n23211) );
  XNOR U23545 ( .A(n23219), .B(n23433), .Z(n23212) );
  XNOR U23546 ( .A(n23218), .B(n23216), .Z(n23433) );
  AND U23547 ( .A(n23434), .B(n23435), .Z(n23216) );
  NANDN U23548 ( .A(n23436), .B(n23437), .Z(n23435) );
  NANDN U23549 ( .A(n23438), .B(n23439), .Z(n23437) );
  NANDN U23550 ( .A(n23439), .B(n23438), .Z(n23434) );
  ANDN U23551 ( .B(B[212]), .A(n70), .Z(n23218) );
  XNOR U23552 ( .A(n23226), .B(n23440), .Z(n23219) );
  XNOR U23553 ( .A(n23225), .B(n23223), .Z(n23440) );
  AND U23554 ( .A(n23441), .B(n23442), .Z(n23223) );
  NANDN U23555 ( .A(n23443), .B(n23444), .Z(n23442) );
  OR U23556 ( .A(n23445), .B(n23446), .Z(n23444) );
  NAND U23557 ( .A(n23446), .B(n23445), .Z(n23441) );
  ANDN U23558 ( .B(B[213]), .A(n71), .Z(n23225) );
  XNOR U23559 ( .A(n23233), .B(n23447), .Z(n23226) );
  XNOR U23560 ( .A(n23232), .B(n23230), .Z(n23447) );
  AND U23561 ( .A(n23448), .B(n23449), .Z(n23230) );
  NANDN U23562 ( .A(n23450), .B(n23451), .Z(n23449) );
  NANDN U23563 ( .A(n23452), .B(n23453), .Z(n23451) );
  NANDN U23564 ( .A(n23453), .B(n23452), .Z(n23448) );
  ANDN U23565 ( .B(B[214]), .A(n72), .Z(n23232) );
  XNOR U23566 ( .A(n23240), .B(n23454), .Z(n23233) );
  XNOR U23567 ( .A(n23239), .B(n23237), .Z(n23454) );
  AND U23568 ( .A(n23455), .B(n23456), .Z(n23237) );
  NANDN U23569 ( .A(n23457), .B(n23458), .Z(n23456) );
  OR U23570 ( .A(n23459), .B(n23460), .Z(n23458) );
  NAND U23571 ( .A(n23460), .B(n23459), .Z(n23455) );
  ANDN U23572 ( .B(B[215]), .A(n73), .Z(n23239) );
  XNOR U23573 ( .A(n23247), .B(n23461), .Z(n23240) );
  XNOR U23574 ( .A(n23246), .B(n23244), .Z(n23461) );
  AND U23575 ( .A(n23462), .B(n23463), .Z(n23244) );
  NANDN U23576 ( .A(n23464), .B(n23465), .Z(n23463) );
  NANDN U23577 ( .A(n23466), .B(n23467), .Z(n23465) );
  NANDN U23578 ( .A(n23467), .B(n23466), .Z(n23462) );
  ANDN U23579 ( .B(B[216]), .A(n74), .Z(n23246) );
  XNOR U23580 ( .A(n23254), .B(n23468), .Z(n23247) );
  XNOR U23581 ( .A(n23253), .B(n23251), .Z(n23468) );
  AND U23582 ( .A(n23469), .B(n23470), .Z(n23251) );
  NANDN U23583 ( .A(n23471), .B(n23472), .Z(n23470) );
  OR U23584 ( .A(n23473), .B(n23474), .Z(n23472) );
  NAND U23585 ( .A(n23474), .B(n23473), .Z(n23469) );
  ANDN U23586 ( .B(B[217]), .A(n75), .Z(n23253) );
  XNOR U23587 ( .A(n23261), .B(n23475), .Z(n23254) );
  XNOR U23588 ( .A(n23260), .B(n23258), .Z(n23475) );
  AND U23589 ( .A(n23476), .B(n23477), .Z(n23258) );
  NANDN U23590 ( .A(n23478), .B(n23479), .Z(n23477) );
  NANDN U23591 ( .A(n23480), .B(n23481), .Z(n23479) );
  NANDN U23592 ( .A(n23481), .B(n23480), .Z(n23476) );
  ANDN U23593 ( .B(B[218]), .A(n76), .Z(n23260) );
  XNOR U23594 ( .A(n23268), .B(n23482), .Z(n23261) );
  XNOR U23595 ( .A(n23267), .B(n23265), .Z(n23482) );
  AND U23596 ( .A(n23483), .B(n23484), .Z(n23265) );
  NANDN U23597 ( .A(n23485), .B(n23486), .Z(n23484) );
  OR U23598 ( .A(n23487), .B(n23488), .Z(n23486) );
  NAND U23599 ( .A(n23488), .B(n23487), .Z(n23483) );
  ANDN U23600 ( .B(B[219]), .A(n77), .Z(n23267) );
  XNOR U23601 ( .A(n23275), .B(n23489), .Z(n23268) );
  XNOR U23602 ( .A(n23274), .B(n23272), .Z(n23489) );
  AND U23603 ( .A(n23490), .B(n23491), .Z(n23272) );
  NANDN U23604 ( .A(n23492), .B(n23493), .Z(n23491) );
  NANDN U23605 ( .A(n23494), .B(n23495), .Z(n23493) );
  NANDN U23606 ( .A(n23495), .B(n23494), .Z(n23490) );
  ANDN U23607 ( .B(B[220]), .A(n78), .Z(n23274) );
  XNOR U23608 ( .A(n23282), .B(n23496), .Z(n23275) );
  XNOR U23609 ( .A(n23281), .B(n23279), .Z(n23496) );
  AND U23610 ( .A(n23497), .B(n23498), .Z(n23279) );
  NANDN U23611 ( .A(n23499), .B(n23500), .Z(n23498) );
  OR U23612 ( .A(n23501), .B(n23502), .Z(n23500) );
  NAND U23613 ( .A(n23502), .B(n23501), .Z(n23497) );
  ANDN U23614 ( .B(B[221]), .A(n79), .Z(n23281) );
  XNOR U23615 ( .A(n23289), .B(n23503), .Z(n23282) );
  XNOR U23616 ( .A(n23288), .B(n23286), .Z(n23503) );
  AND U23617 ( .A(n23504), .B(n23505), .Z(n23286) );
  NANDN U23618 ( .A(n23506), .B(n23507), .Z(n23505) );
  NANDN U23619 ( .A(n23508), .B(n23509), .Z(n23507) );
  NANDN U23620 ( .A(n23509), .B(n23508), .Z(n23504) );
  ANDN U23621 ( .B(B[222]), .A(n80), .Z(n23288) );
  XNOR U23622 ( .A(n23296), .B(n23510), .Z(n23289) );
  XNOR U23623 ( .A(n23295), .B(n23293), .Z(n23510) );
  AND U23624 ( .A(n23511), .B(n23512), .Z(n23293) );
  NANDN U23625 ( .A(n23513), .B(n23514), .Z(n23512) );
  OR U23626 ( .A(n23515), .B(n23516), .Z(n23514) );
  NAND U23627 ( .A(n23516), .B(n23515), .Z(n23511) );
  ANDN U23628 ( .B(B[223]), .A(n81), .Z(n23295) );
  XNOR U23629 ( .A(n23303), .B(n23517), .Z(n23296) );
  XNOR U23630 ( .A(n23302), .B(n23300), .Z(n23517) );
  AND U23631 ( .A(n23518), .B(n23519), .Z(n23300) );
  NANDN U23632 ( .A(n23520), .B(n23521), .Z(n23519) );
  NAND U23633 ( .A(n23522), .B(n23523), .Z(n23521) );
  ANDN U23634 ( .B(B[224]), .A(n82), .Z(n23302) );
  XOR U23635 ( .A(n23309), .B(n23524), .Z(n23303) );
  XNOR U23636 ( .A(n23307), .B(n23310), .Z(n23524) );
  NAND U23637 ( .A(A[2]), .B(B[225]), .Z(n23310) );
  NANDN U23638 ( .A(n23525), .B(n23526), .Z(n23307) );
  AND U23639 ( .A(A[0]), .B(B[226]), .Z(n23526) );
  XNOR U23640 ( .A(n23312), .B(n23527), .Z(n23309) );
  NAND U23641 ( .A(A[0]), .B(B[227]), .Z(n23527) );
  NAND U23642 ( .A(B[226]), .B(A[1]), .Z(n23312) );
  NAND U23643 ( .A(n23528), .B(n23529), .Z(n342) );
  NANDN U23644 ( .A(n23530), .B(n23531), .Z(n23529) );
  OR U23645 ( .A(n23532), .B(n23533), .Z(n23531) );
  NAND U23646 ( .A(n23533), .B(n23532), .Z(n23528) );
  XOR U23647 ( .A(n344), .B(n343), .Z(\A1[224] ) );
  XOR U23648 ( .A(n23533), .B(n23534), .Z(n343) );
  XNOR U23649 ( .A(n23532), .B(n23530), .Z(n23534) );
  AND U23650 ( .A(n23535), .B(n23536), .Z(n23530) );
  NANDN U23651 ( .A(n23537), .B(n23538), .Z(n23536) );
  NANDN U23652 ( .A(n23539), .B(n23540), .Z(n23538) );
  NANDN U23653 ( .A(n23540), .B(n23539), .Z(n23535) );
  ANDN U23654 ( .B(B[195]), .A(n54), .Z(n23532) );
  XNOR U23655 ( .A(n23327), .B(n23541), .Z(n23533) );
  XNOR U23656 ( .A(n23326), .B(n23324), .Z(n23541) );
  AND U23657 ( .A(n23542), .B(n23543), .Z(n23324) );
  NANDN U23658 ( .A(n23544), .B(n23545), .Z(n23543) );
  OR U23659 ( .A(n23546), .B(n23547), .Z(n23545) );
  NAND U23660 ( .A(n23547), .B(n23546), .Z(n23542) );
  ANDN U23661 ( .B(B[196]), .A(n55), .Z(n23326) );
  XNOR U23662 ( .A(n23334), .B(n23548), .Z(n23327) );
  XNOR U23663 ( .A(n23333), .B(n23331), .Z(n23548) );
  AND U23664 ( .A(n23549), .B(n23550), .Z(n23331) );
  NANDN U23665 ( .A(n23551), .B(n23552), .Z(n23550) );
  NANDN U23666 ( .A(n23553), .B(n23554), .Z(n23552) );
  NANDN U23667 ( .A(n23554), .B(n23553), .Z(n23549) );
  ANDN U23668 ( .B(B[197]), .A(n56), .Z(n23333) );
  XNOR U23669 ( .A(n23341), .B(n23555), .Z(n23334) );
  XNOR U23670 ( .A(n23340), .B(n23338), .Z(n23555) );
  AND U23671 ( .A(n23556), .B(n23557), .Z(n23338) );
  NANDN U23672 ( .A(n23558), .B(n23559), .Z(n23557) );
  OR U23673 ( .A(n23560), .B(n23561), .Z(n23559) );
  NAND U23674 ( .A(n23561), .B(n23560), .Z(n23556) );
  ANDN U23675 ( .B(B[198]), .A(n57), .Z(n23340) );
  XNOR U23676 ( .A(n23348), .B(n23562), .Z(n23341) );
  XNOR U23677 ( .A(n23347), .B(n23345), .Z(n23562) );
  AND U23678 ( .A(n23563), .B(n23564), .Z(n23345) );
  NANDN U23679 ( .A(n23565), .B(n23566), .Z(n23564) );
  NANDN U23680 ( .A(n23567), .B(n23568), .Z(n23566) );
  NANDN U23681 ( .A(n23568), .B(n23567), .Z(n23563) );
  ANDN U23682 ( .B(B[199]), .A(n58), .Z(n23347) );
  XNOR U23683 ( .A(n23355), .B(n23569), .Z(n23348) );
  XNOR U23684 ( .A(n23354), .B(n23352), .Z(n23569) );
  AND U23685 ( .A(n23570), .B(n23571), .Z(n23352) );
  NANDN U23686 ( .A(n23572), .B(n23573), .Z(n23571) );
  OR U23687 ( .A(n23574), .B(n23575), .Z(n23573) );
  NAND U23688 ( .A(n23575), .B(n23574), .Z(n23570) );
  ANDN U23689 ( .B(B[200]), .A(n59), .Z(n23354) );
  XNOR U23690 ( .A(n23362), .B(n23576), .Z(n23355) );
  XNOR U23691 ( .A(n23361), .B(n23359), .Z(n23576) );
  AND U23692 ( .A(n23577), .B(n23578), .Z(n23359) );
  NANDN U23693 ( .A(n23579), .B(n23580), .Z(n23578) );
  NANDN U23694 ( .A(n23581), .B(n23582), .Z(n23580) );
  NANDN U23695 ( .A(n23582), .B(n23581), .Z(n23577) );
  ANDN U23696 ( .B(B[201]), .A(n60), .Z(n23361) );
  XNOR U23697 ( .A(n23369), .B(n23583), .Z(n23362) );
  XNOR U23698 ( .A(n23368), .B(n23366), .Z(n23583) );
  AND U23699 ( .A(n23584), .B(n23585), .Z(n23366) );
  NANDN U23700 ( .A(n23586), .B(n23587), .Z(n23585) );
  OR U23701 ( .A(n23588), .B(n23589), .Z(n23587) );
  NAND U23702 ( .A(n23589), .B(n23588), .Z(n23584) );
  ANDN U23703 ( .B(B[202]), .A(n61), .Z(n23368) );
  XNOR U23704 ( .A(n23376), .B(n23590), .Z(n23369) );
  XNOR U23705 ( .A(n23375), .B(n23373), .Z(n23590) );
  AND U23706 ( .A(n23591), .B(n23592), .Z(n23373) );
  NANDN U23707 ( .A(n23593), .B(n23594), .Z(n23592) );
  NANDN U23708 ( .A(n23595), .B(n23596), .Z(n23594) );
  NANDN U23709 ( .A(n23596), .B(n23595), .Z(n23591) );
  ANDN U23710 ( .B(B[203]), .A(n62), .Z(n23375) );
  XNOR U23711 ( .A(n23383), .B(n23597), .Z(n23376) );
  XNOR U23712 ( .A(n23382), .B(n23380), .Z(n23597) );
  AND U23713 ( .A(n23598), .B(n23599), .Z(n23380) );
  NANDN U23714 ( .A(n23600), .B(n23601), .Z(n23599) );
  OR U23715 ( .A(n23602), .B(n23603), .Z(n23601) );
  NAND U23716 ( .A(n23603), .B(n23602), .Z(n23598) );
  ANDN U23717 ( .B(B[204]), .A(n63), .Z(n23382) );
  XNOR U23718 ( .A(n23390), .B(n23604), .Z(n23383) );
  XNOR U23719 ( .A(n23389), .B(n23387), .Z(n23604) );
  AND U23720 ( .A(n23605), .B(n23606), .Z(n23387) );
  NANDN U23721 ( .A(n23607), .B(n23608), .Z(n23606) );
  NANDN U23722 ( .A(n23609), .B(n23610), .Z(n23608) );
  NANDN U23723 ( .A(n23610), .B(n23609), .Z(n23605) );
  ANDN U23724 ( .B(B[205]), .A(n64), .Z(n23389) );
  XNOR U23725 ( .A(n23397), .B(n23611), .Z(n23390) );
  XNOR U23726 ( .A(n23396), .B(n23394), .Z(n23611) );
  AND U23727 ( .A(n23612), .B(n23613), .Z(n23394) );
  NANDN U23728 ( .A(n23614), .B(n23615), .Z(n23613) );
  OR U23729 ( .A(n23616), .B(n23617), .Z(n23615) );
  NAND U23730 ( .A(n23617), .B(n23616), .Z(n23612) );
  ANDN U23731 ( .B(B[206]), .A(n65), .Z(n23396) );
  XNOR U23732 ( .A(n23404), .B(n23618), .Z(n23397) );
  XNOR U23733 ( .A(n23403), .B(n23401), .Z(n23618) );
  AND U23734 ( .A(n23619), .B(n23620), .Z(n23401) );
  NANDN U23735 ( .A(n23621), .B(n23622), .Z(n23620) );
  NANDN U23736 ( .A(n23623), .B(n23624), .Z(n23622) );
  NANDN U23737 ( .A(n23624), .B(n23623), .Z(n23619) );
  ANDN U23738 ( .B(B[207]), .A(n66), .Z(n23403) );
  XNOR U23739 ( .A(n23411), .B(n23625), .Z(n23404) );
  XNOR U23740 ( .A(n23410), .B(n23408), .Z(n23625) );
  AND U23741 ( .A(n23626), .B(n23627), .Z(n23408) );
  NANDN U23742 ( .A(n23628), .B(n23629), .Z(n23627) );
  OR U23743 ( .A(n23630), .B(n23631), .Z(n23629) );
  NAND U23744 ( .A(n23631), .B(n23630), .Z(n23626) );
  ANDN U23745 ( .B(B[208]), .A(n67), .Z(n23410) );
  XNOR U23746 ( .A(n23418), .B(n23632), .Z(n23411) );
  XNOR U23747 ( .A(n23417), .B(n23415), .Z(n23632) );
  AND U23748 ( .A(n23633), .B(n23634), .Z(n23415) );
  NANDN U23749 ( .A(n23635), .B(n23636), .Z(n23634) );
  NANDN U23750 ( .A(n23637), .B(n23638), .Z(n23636) );
  NANDN U23751 ( .A(n23638), .B(n23637), .Z(n23633) );
  ANDN U23752 ( .B(B[209]), .A(n68), .Z(n23417) );
  XNOR U23753 ( .A(n23425), .B(n23639), .Z(n23418) );
  XNOR U23754 ( .A(n23424), .B(n23422), .Z(n23639) );
  AND U23755 ( .A(n23640), .B(n23641), .Z(n23422) );
  NANDN U23756 ( .A(n23642), .B(n23643), .Z(n23641) );
  OR U23757 ( .A(n23644), .B(n23645), .Z(n23643) );
  NAND U23758 ( .A(n23645), .B(n23644), .Z(n23640) );
  ANDN U23759 ( .B(B[210]), .A(n69), .Z(n23424) );
  XNOR U23760 ( .A(n23432), .B(n23646), .Z(n23425) );
  XNOR U23761 ( .A(n23431), .B(n23429), .Z(n23646) );
  AND U23762 ( .A(n23647), .B(n23648), .Z(n23429) );
  NANDN U23763 ( .A(n23649), .B(n23650), .Z(n23648) );
  NANDN U23764 ( .A(n23651), .B(n23652), .Z(n23650) );
  NANDN U23765 ( .A(n23652), .B(n23651), .Z(n23647) );
  ANDN U23766 ( .B(B[211]), .A(n70), .Z(n23431) );
  XNOR U23767 ( .A(n23439), .B(n23653), .Z(n23432) );
  XNOR U23768 ( .A(n23438), .B(n23436), .Z(n23653) );
  AND U23769 ( .A(n23654), .B(n23655), .Z(n23436) );
  NANDN U23770 ( .A(n23656), .B(n23657), .Z(n23655) );
  OR U23771 ( .A(n23658), .B(n23659), .Z(n23657) );
  NAND U23772 ( .A(n23659), .B(n23658), .Z(n23654) );
  ANDN U23773 ( .B(B[212]), .A(n71), .Z(n23438) );
  XNOR U23774 ( .A(n23446), .B(n23660), .Z(n23439) );
  XNOR U23775 ( .A(n23445), .B(n23443), .Z(n23660) );
  AND U23776 ( .A(n23661), .B(n23662), .Z(n23443) );
  NANDN U23777 ( .A(n23663), .B(n23664), .Z(n23662) );
  NANDN U23778 ( .A(n23665), .B(n23666), .Z(n23664) );
  NANDN U23779 ( .A(n23666), .B(n23665), .Z(n23661) );
  ANDN U23780 ( .B(B[213]), .A(n72), .Z(n23445) );
  XNOR U23781 ( .A(n23453), .B(n23667), .Z(n23446) );
  XNOR U23782 ( .A(n23452), .B(n23450), .Z(n23667) );
  AND U23783 ( .A(n23668), .B(n23669), .Z(n23450) );
  NANDN U23784 ( .A(n23670), .B(n23671), .Z(n23669) );
  OR U23785 ( .A(n23672), .B(n23673), .Z(n23671) );
  NAND U23786 ( .A(n23673), .B(n23672), .Z(n23668) );
  ANDN U23787 ( .B(B[214]), .A(n73), .Z(n23452) );
  XNOR U23788 ( .A(n23460), .B(n23674), .Z(n23453) );
  XNOR U23789 ( .A(n23459), .B(n23457), .Z(n23674) );
  AND U23790 ( .A(n23675), .B(n23676), .Z(n23457) );
  NANDN U23791 ( .A(n23677), .B(n23678), .Z(n23676) );
  NANDN U23792 ( .A(n23679), .B(n23680), .Z(n23678) );
  NANDN U23793 ( .A(n23680), .B(n23679), .Z(n23675) );
  ANDN U23794 ( .B(B[215]), .A(n74), .Z(n23459) );
  XNOR U23795 ( .A(n23467), .B(n23681), .Z(n23460) );
  XNOR U23796 ( .A(n23466), .B(n23464), .Z(n23681) );
  AND U23797 ( .A(n23682), .B(n23683), .Z(n23464) );
  NANDN U23798 ( .A(n23684), .B(n23685), .Z(n23683) );
  OR U23799 ( .A(n23686), .B(n23687), .Z(n23685) );
  NAND U23800 ( .A(n23687), .B(n23686), .Z(n23682) );
  ANDN U23801 ( .B(B[216]), .A(n75), .Z(n23466) );
  XNOR U23802 ( .A(n23474), .B(n23688), .Z(n23467) );
  XNOR U23803 ( .A(n23473), .B(n23471), .Z(n23688) );
  AND U23804 ( .A(n23689), .B(n23690), .Z(n23471) );
  NANDN U23805 ( .A(n23691), .B(n23692), .Z(n23690) );
  NANDN U23806 ( .A(n23693), .B(n23694), .Z(n23692) );
  NANDN U23807 ( .A(n23694), .B(n23693), .Z(n23689) );
  ANDN U23808 ( .B(B[217]), .A(n76), .Z(n23473) );
  XNOR U23809 ( .A(n23481), .B(n23695), .Z(n23474) );
  XNOR U23810 ( .A(n23480), .B(n23478), .Z(n23695) );
  AND U23811 ( .A(n23696), .B(n23697), .Z(n23478) );
  NANDN U23812 ( .A(n23698), .B(n23699), .Z(n23697) );
  OR U23813 ( .A(n23700), .B(n23701), .Z(n23699) );
  NAND U23814 ( .A(n23701), .B(n23700), .Z(n23696) );
  ANDN U23815 ( .B(B[218]), .A(n77), .Z(n23480) );
  XNOR U23816 ( .A(n23488), .B(n23702), .Z(n23481) );
  XNOR U23817 ( .A(n23487), .B(n23485), .Z(n23702) );
  AND U23818 ( .A(n23703), .B(n23704), .Z(n23485) );
  NANDN U23819 ( .A(n23705), .B(n23706), .Z(n23704) );
  NANDN U23820 ( .A(n23707), .B(n23708), .Z(n23706) );
  NANDN U23821 ( .A(n23708), .B(n23707), .Z(n23703) );
  ANDN U23822 ( .B(B[219]), .A(n78), .Z(n23487) );
  XNOR U23823 ( .A(n23495), .B(n23709), .Z(n23488) );
  XNOR U23824 ( .A(n23494), .B(n23492), .Z(n23709) );
  AND U23825 ( .A(n23710), .B(n23711), .Z(n23492) );
  NANDN U23826 ( .A(n23712), .B(n23713), .Z(n23711) );
  OR U23827 ( .A(n23714), .B(n23715), .Z(n23713) );
  NAND U23828 ( .A(n23715), .B(n23714), .Z(n23710) );
  ANDN U23829 ( .B(B[220]), .A(n79), .Z(n23494) );
  XNOR U23830 ( .A(n23502), .B(n23716), .Z(n23495) );
  XNOR U23831 ( .A(n23501), .B(n23499), .Z(n23716) );
  AND U23832 ( .A(n23717), .B(n23718), .Z(n23499) );
  NANDN U23833 ( .A(n23719), .B(n23720), .Z(n23718) );
  NANDN U23834 ( .A(n23721), .B(n23722), .Z(n23720) );
  NANDN U23835 ( .A(n23722), .B(n23721), .Z(n23717) );
  ANDN U23836 ( .B(B[221]), .A(n80), .Z(n23501) );
  XNOR U23837 ( .A(n23509), .B(n23723), .Z(n23502) );
  XNOR U23838 ( .A(n23508), .B(n23506), .Z(n23723) );
  AND U23839 ( .A(n23724), .B(n23725), .Z(n23506) );
  NANDN U23840 ( .A(n23726), .B(n23727), .Z(n23725) );
  OR U23841 ( .A(n23728), .B(n23729), .Z(n23727) );
  NAND U23842 ( .A(n23729), .B(n23728), .Z(n23724) );
  ANDN U23843 ( .B(B[222]), .A(n81), .Z(n23508) );
  XNOR U23844 ( .A(n23516), .B(n23730), .Z(n23509) );
  XNOR U23845 ( .A(n23515), .B(n23513), .Z(n23730) );
  AND U23846 ( .A(n23731), .B(n23732), .Z(n23513) );
  NANDN U23847 ( .A(n23733), .B(n23734), .Z(n23732) );
  NAND U23848 ( .A(n23735), .B(n23736), .Z(n23734) );
  ANDN U23849 ( .B(B[223]), .A(n82), .Z(n23515) );
  XOR U23850 ( .A(n23522), .B(n23737), .Z(n23516) );
  XNOR U23851 ( .A(n23520), .B(n23523), .Z(n23737) );
  NAND U23852 ( .A(A[2]), .B(B[224]), .Z(n23523) );
  NANDN U23853 ( .A(n23738), .B(n23739), .Z(n23520) );
  AND U23854 ( .A(A[0]), .B(B[225]), .Z(n23739) );
  XNOR U23855 ( .A(n23525), .B(n23740), .Z(n23522) );
  NAND U23856 ( .A(A[0]), .B(B[226]), .Z(n23740) );
  NAND U23857 ( .A(B[225]), .B(A[1]), .Z(n23525) );
  NAND U23858 ( .A(n23741), .B(n23742), .Z(n344) );
  NANDN U23859 ( .A(n23743), .B(n23744), .Z(n23742) );
  OR U23860 ( .A(n23745), .B(n23746), .Z(n23744) );
  NAND U23861 ( .A(n23746), .B(n23745), .Z(n23741) );
  XOR U23862 ( .A(n346), .B(n345), .Z(\A1[223] ) );
  XOR U23863 ( .A(n23746), .B(n23747), .Z(n345) );
  XNOR U23864 ( .A(n23745), .B(n23743), .Z(n23747) );
  AND U23865 ( .A(n23748), .B(n23749), .Z(n23743) );
  NANDN U23866 ( .A(n23750), .B(n23751), .Z(n23749) );
  NANDN U23867 ( .A(n23752), .B(n23753), .Z(n23751) );
  NANDN U23868 ( .A(n23753), .B(n23752), .Z(n23748) );
  ANDN U23869 ( .B(B[194]), .A(n54), .Z(n23745) );
  XNOR U23870 ( .A(n23540), .B(n23754), .Z(n23746) );
  XNOR U23871 ( .A(n23539), .B(n23537), .Z(n23754) );
  AND U23872 ( .A(n23755), .B(n23756), .Z(n23537) );
  NANDN U23873 ( .A(n23757), .B(n23758), .Z(n23756) );
  OR U23874 ( .A(n23759), .B(n23760), .Z(n23758) );
  NAND U23875 ( .A(n23760), .B(n23759), .Z(n23755) );
  ANDN U23876 ( .B(B[195]), .A(n55), .Z(n23539) );
  XNOR U23877 ( .A(n23547), .B(n23761), .Z(n23540) );
  XNOR U23878 ( .A(n23546), .B(n23544), .Z(n23761) );
  AND U23879 ( .A(n23762), .B(n23763), .Z(n23544) );
  NANDN U23880 ( .A(n23764), .B(n23765), .Z(n23763) );
  NANDN U23881 ( .A(n23766), .B(n23767), .Z(n23765) );
  NANDN U23882 ( .A(n23767), .B(n23766), .Z(n23762) );
  ANDN U23883 ( .B(B[196]), .A(n56), .Z(n23546) );
  XNOR U23884 ( .A(n23554), .B(n23768), .Z(n23547) );
  XNOR U23885 ( .A(n23553), .B(n23551), .Z(n23768) );
  AND U23886 ( .A(n23769), .B(n23770), .Z(n23551) );
  NANDN U23887 ( .A(n23771), .B(n23772), .Z(n23770) );
  OR U23888 ( .A(n23773), .B(n23774), .Z(n23772) );
  NAND U23889 ( .A(n23774), .B(n23773), .Z(n23769) );
  ANDN U23890 ( .B(B[197]), .A(n57), .Z(n23553) );
  XNOR U23891 ( .A(n23561), .B(n23775), .Z(n23554) );
  XNOR U23892 ( .A(n23560), .B(n23558), .Z(n23775) );
  AND U23893 ( .A(n23776), .B(n23777), .Z(n23558) );
  NANDN U23894 ( .A(n23778), .B(n23779), .Z(n23777) );
  NANDN U23895 ( .A(n23780), .B(n23781), .Z(n23779) );
  NANDN U23896 ( .A(n23781), .B(n23780), .Z(n23776) );
  ANDN U23897 ( .B(B[198]), .A(n58), .Z(n23560) );
  XNOR U23898 ( .A(n23568), .B(n23782), .Z(n23561) );
  XNOR U23899 ( .A(n23567), .B(n23565), .Z(n23782) );
  AND U23900 ( .A(n23783), .B(n23784), .Z(n23565) );
  NANDN U23901 ( .A(n23785), .B(n23786), .Z(n23784) );
  OR U23902 ( .A(n23787), .B(n23788), .Z(n23786) );
  NAND U23903 ( .A(n23788), .B(n23787), .Z(n23783) );
  ANDN U23904 ( .B(B[199]), .A(n59), .Z(n23567) );
  XNOR U23905 ( .A(n23575), .B(n23789), .Z(n23568) );
  XNOR U23906 ( .A(n23574), .B(n23572), .Z(n23789) );
  AND U23907 ( .A(n23790), .B(n23791), .Z(n23572) );
  NANDN U23908 ( .A(n23792), .B(n23793), .Z(n23791) );
  NANDN U23909 ( .A(n23794), .B(n23795), .Z(n23793) );
  NANDN U23910 ( .A(n23795), .B(n23794), .Z(n23790) );
  ANDN U23911 ( .B(B[200]), .A(n60), .Z(n23574) );
  XNOR U23912 ( .A(n23582), .B(n23796), .Z(n23575) );
  XNOR U23913 ( .A(n23581), .B(n23579), .Z(n23796) );
  AND U23914 ( .A(n23797), .B(n23798), .Z(n23579) );
  NANDN U23915 ( .A(n23799), .B(n23800), .Z(n23798) );
  OR U23916 ( .A(n23801), .B(n23802), .Z(n23800) );
  NAND U23917 ( .A(n23802), .B(n23801), .Z(n23797) );
  ANDN U23918 ( .B(B[201]), .A(n61), .Z(n23581) );
  XNOR U23919 ( .A(n23589), .B(n23803), .Z(n23582) );
  XNOR U23920 ( .A(n23588), .B(n23586), .Z(n23803) );
  AND U23921 ( .A(n23804), .B(n23805), .Z(n23586) );
  NANDN U23922 ( .A(n23806), .B(n23807), .Z(n23805) );
  NANDN U23923 ( .A(n23808), .B(n23809), .Z(n23807) );
  NANDN U23924 ( .A(n23809), .B(n23808), .Z(n23804) );
  ANDN U23925 ( .B(B[202]), .A(n62), .Z(n23588) );
  XNOR U23926 ( .A(n23596), .B(n23810), .Z(n23589) );
  XNOR U23927 ( .A(n23595), .B(n23593), .Z(n23810) );
  AND U23928 ( .A(n23811), .B(n23812), .Z(n23593) );
  NANDN U23929 ( .A(n23813), .B(n23814), .Z(n23812) );
  OR U23930 ( .A(n23815), .B(n23816), .Z(n23814) );
  NAND U23931 ( .A(n23816), .B(n23815), .Z(n23811) );
  ANDN U23932 ( .B(B[203]), .A(n63), .Z(n23595) );
  XNOR U23933 ( .A(n23603), .B(n23817), .Z(n23596) );
  XNOR U23934 ( .A(n23602), .B(n23600), .Z(n23817) );
  AND U23935 ( .A(n23818), .B(n23819), .Z(n23600) );
  NANDN U23936 ( .A(n23820), .B(n23821), .Z(n23819) );
  NANDN U23937 ( .A(n23822), .B(n23823), .Z(n23821) );
  NANDN U23938 ( .A(n23823), .B(n23822), .Z(n23818) );
  ANDN U23939 ( .B(B[204]), .A(n64), .Z(n23602) );
  XNOR U23940 ( .A(n23610), .B(n23824), .Z(n23603) );
  XNOR U23941 ( .A(n23609), .B(n23607), .Z(n23824) );
  AND U23942 ( .A(n23825), .B(n23826), .Z(n23607) );
  NANDN U23943 ( .A(n23827), .B(n23828), .Z(n23826) );
  OR U23944 ( .A(n23829), .B(n23830), .Z(n23828) );
  NAND U23945 ( .A(n23830), .B(n23829), .Z(n23825) );
  ANDN U23946 ( .B(B[205]), .A(n65), .Z(n23609) );
  XNOR U23947 ( .A(n23617), .B(n23831), .Z(n23610) );
  XNOR U23948 ( .A(n23616), .B(n23614), .Z(n23831) );
  AND U23949 ( .A(n23832), .B(n23833), .Z(n23614) );
  NANDN U23950 ( .A(n23834), .B(n23835), .Z(n23833) );
  NANDN U23951 ( .A(n23836), .B(n23837), .Z(n23835) );
  NANDN U23952 ( .A(n23837), .B(n23836), .Z(n23832) );
  ANDN U23953 ( .B(B[206]), .A(n66), .Z(n23616) );
  XNOR U23954 ( .A(n23624), .B(n23838), .Z(n23617) );
  XNOR U23955 ( .A(n23623), .B(n23621), .Z(n23838) );
  AND U23956 ( .A(n23839), .B(n23840), .Z(n23621) );
  NANDN U23957 ( .A(n23841), .B(n23842), .Z(n23840) );
  OR U23958 ( .A(n23843), .B(n23844), .Z(n23842) );
  NAND U23959 ( .A(n23844), .B(n23843), .Z(n23839) );
  ANDN U23960 ( .B(B[207]), .A(n67), .Z(n23623) );
  XNOR U23961 ( .A(n23631), .B(n23845), .Z(n23624) );
  XNOR U23962 ( .A(n23630), .B(n23628), .Z(n23845) );
  AND U23963 ( .A(n23846), .B(n23847), .Z(n23628) );
  NANDN U23964 ( .A(n23848), .B(n23849), .Z(n23847) );
  NANDN U23965 ( .A(n23850), .B(n23851), .Z(n23849) );
  NANDN U23966 ( .A(n23851), .B(n23850), .Z(n23846) );
  ANDN U23967 ( .B(B[208]), .A(n68), .Z(n23630) );
  XNOR U23968 ( .A(n23638), .B(n23852), .Z(n23631) );
  XNOR U23969 ( .A(n23637), .B(n23635), .Z(n23852) );
  AND U23970 ( .A(n23853), .B(n23854), .Z(n23635) );
  NANDN U23971 ( .A(n23855), .B(n23856), .Z(n23854) );
  OR U23972 ( .A(n23857), .B(n23858), .Z(n23856) );
  NAND U23973 ( .A(n23858), .B(n23857), .Z(n23853) );
  ANDN U23974 ( .B(B[209]), .A(n69), .Z(n23637) );
  XNOR U23975 ( .A(n23645), .B(n23859), .Z(n23638) );
  XNOR U23976 ( .A(n23644), .B(n23642), .Z(n23859) );
  AND U23977 ( .A(n23860), .B(n23861), .Z(n23642) );
  NANDN U23978 ( .A(n23862), .B(n23863), .Z(n23861) );
  NANDN U23979 ( .A(n23864), .B(n23865), .Z(n23863) );
  NANDN U23980 ( .A(n23865), .B(n23864), .Z(n23860) );
  ANDN U23981 ( .B(B[210]), .A(n70), .Z(n23644) );
  XNOR U23982 ( .A(n23652), .B(n23866), .Z(n23645) );
  XNOR U23983 ( .A(n23651), .B(n23649), .Z(n23866) );
  AND U23984 ( .A(n23867), .B(n23868), .Z(n23649) );
  NANDN U23985 ( .A(n23869), .B(n23870), .Z(n23868) );
  OR U23986 ( .A(n23871), .B(n23872), .Z(n23870) );
  NAND U23987 ( .A(n23872), .B(n23871), .Z(n23867) );
  ANDN U23988 ( .B(B[211]), .A(n71), .Z(n23651) );
  XNOR U23989 ( .A(n23659), .B(n23873), .Z(n23652) );
  XNOR U23990 ( .A(n23658), .B(n23656), .Z(n23873) );
  AND U23991 ( .A(n23874), .B(n23875), .Z(n23656) );
  NANDN U23992 ( .A(n23876), .B(n23877), .Z(n23875) );
  NANDN U23993 ( .A(n23878), .B(n23879), .Z(n23877) );
  NANDN U23994 ( .A(n23879), .B(n23878), .Z(n23874) );
  ANDN U23995 ( .B(B[212]), .A(n72), .Z(n23658) );
  XNOR U23996 ( .A(n23666), .B(n23880), .Z(n23659) );
  XNOR U23997 ( .A(n23665), .B(n23663), .Z(n23880) );
  AND U23998 ( .A(n23881), .B(n23882), .Z(n23663) );
  NANDN U23999 ( .A(n23883), .B(n23884), .Z(n23882) );
  OR U24000 ( .A(n23885), .B(n23886), .Z(n23884) );
  NAND U24001 ( .A(n23886), .B(n23885), .Z(n23881) );
  ANDN U24002 ( .B(B[213]), .A(n73), .Z(n23665) );
  XNOR U24003 ( .A(n23673), .B(n23887), .Z(n23666) );
  XNOR U24004 ( .A(n23672), .B(n23670), .Z(n23887) );
  AND U24005 ( .A(n23888), .B(n23889), .Z(n23670) );
  NANDN U24006 ( .A(n23890), .B(n23891), .Z(n23889) );
  NANDN U24007 ( .A(n23892), .B(n23893), .Z(n23891) );
  NANDN U24008 ( .A(n23893), .B(n23892), .Z(n23888) );
  ANDN U24009 ( .B(B[214]), .A(n74), .Z(n23672) );
  XNOR U24010 ( .A(n23680), .B(n23894), .Z(n23673) );
  XNOR U24011 ( .A(n23679), .B(n23677), .Z(n23894) );
  AND U24012 ( .A(n23895), .B(n23896), .Z(n23677) );
  NANDN U24013 ( .A(n23897), .B(n23898), .Z(n23896) );
  OR U24014 ( .A(n23899), .B(n23900), .Z(n23898) );
  NAND U24015 ( .A(n23900), .B(n23899), .Z(n23895) );
  ANDN U24016 ( .B(B[215]), .A(n75), .Z(n23679) );
  XNOR U24017 ( .A(n23687), .B(n23901), .Z(n23680) );
  XNOR U24018 ( .A(n23686), .B(n23684), .Z(n23901) );
  AND U24019 ( .A(n23902), .B(n23903), .Z(n23684) );
  NANDN U24020 ( .A(n23904), .B(n23905), .Z(n23903) );
  NANDN U24021 ( .A(n23906), .B(n23907), .Z(n23905) );
  NANDN U24022 ( .A(n23907), .B(n23906), .Z(n23902) );
  ANDN U24023 ( .B(B[216]), .A(n76), .Z(n23686) );
  XNOR U24024 ( .A(n23694), .B(n23908), .Z(n23687) );
  XNOR U24025 ( .A(n23693), .B(n23691), .Z(n23908) );
  AND U24026 ( .A(n23909), .B(n23910), .Z(n23691) );
  NANDN U24027 ( .A(n23911), .B(n23912), .Z(n23910) );
  OR U24028 ( .A(n23913), .B(n23914), .Z(n23912) );
  NAND U24029 ( .A(n23914), .B(n23913), .Z(n23909) );
  ANDN U24030 ( .B(B[217]), .A(n77), .Z(n23693) );
  XNOR U24031 ( .A(n23701), .B(n23915), .Z(n23694) );
  XNOR U24032 ( .A(n23700), .B(n23698), .Z(n23915) );
  AND U24033 ( .A(n23916), .B(n23917), .Z(n23698) );
  NANDN U24034 ( .A(n23918), .B(n23919), .Z(n23917) );
  NANDN U24035 ( .A(n23920), .B(n23921), .Z(n23919) );
  NANDN U24036 ( .A(n23921), .B(n23920), .Z(n23916) );
  ANDN U24037 ( .B(B[218]), .A(n78), .Z(n23700) );
  XNOR U24038 ( .A(n23708), .B(n23922), .Z(n23701) );
  XNOR U24039 ( .A(n23707), .B(n23705), .Z(n23922) );
  AND U24040 ( .A(n23923), .B(n23924), .Z(n23705) );
  NANDN U24041 ( .A(n23925), .B(n23926), .Z(n23924) );
  OR U24042 ( .A(n23927), .B(n23928), .Z(n23926) );
  NAND U24043 ( .A(n23928), .B(n23927), .Z(n23923) );
  ANDN U24044 ( .B(B[219]), .A(n79), .Z(n23707) );
  XNOR U24045 ( .A(n23715), .B(n23929), .Z(n23708) );
  XNOR U24046 ( .A(n23714), .B(n23712), .Z(n23929) );
  AND U24047 ( .A(n23930), .B(n23931), .Z(n23712) );
  NANDN U24048 ( .A(n23932), .B(n23933), .Z(n23931) );
  NANDN U24049 ( .A(n23934), .B(n23935), .Z(n23933) );
  NANDN U24050 ( .A(n23935), .B(n23934), .Z(n23930) );
  ANDN U24051 ( .B(B[220]), .A(n80), .Z(n23714) );
  XNOR U24052 ( .A(n23722), .B(n23936), .Z(n23715) );
  XNOR U24053 ( .A(n23721), .B(n23719), .Z(n23936) );
  AND U24054 ( .A(n23937), .B(n23938), .Z(n23719) );
  NANDN U24055 ( .A(n23939), .B(n23940), .Z(n23938) );
  OR U24056 ( .A(n23941), .B(n23942), .Z(n23940) );
  NAND U24057 ( .A(n23942), .B(n23941), .Z(n23937) );
  ANDN U24058 ( .B(B[221]), .A(n81), .Z(n23721) );
  XNOR U24059 ( .A(n23729), .B(n23943), .Z(n23722) );
  XNOR U24060 ( .A(n23728), .B(n23726), .Z(n23943) );
  AND U24061 ( .A(n23944), .B(n23945), .Z(n23726) );
  NANDN U24062 ( .A(n23946), .B(n23947), .Z(n23945) );
  NAND U24063 ( .A(n23948), .B(n23949), .Z(n23947) );
  ANDN U24064 ( .B(B[222]), .A(n82), .Z(n23728) );
  XOR U24065 ( .A(n23735), .B(n23950), .Z(n23729) );
  XNOR U24066 ( .A(n23733), .B(n23736), .Z(n23950) );
  NAND U24067 ( .A(A[2]), .B(B[223]), .Z(n23736) );
  NANDN U24068 ( .A(n23951), .B(n23952), .Z(n23733) );
  AND U24069 ( .A(A[0]), .B(B[224]), .Z(n23952) );
  XNOR U24070 ( .A(n23738), .B(n23953), .Z(n23735) );
  NAND U24071 ( .A(A[0]), .B(B[225]), .Z(n23953) );
  NAND U24072 ( .A(B[224]), .B(A[1]), .Z(n23738) );
  NAND U24073 ( .A(n23954), .B(n23955), .Z(n346) );
  NANDN U24074 ( .A(n23956), .B(n23957), .Z(n23955) );
  OR U24075 ( .A(n23958), .B(n23959), .Z(n23957) );
  NAND U24076 ( .A(n23959), .B(n23958), .Z(n23954) );
  XOR U24077 ( .A(n348), .B(n347), .Z(\A1[222] ) );
  XOR U24078 ( .A(n23959), .B(n23960), .Z(n347) );
  XNOR U24079 ( .A(n23958), .B(n23956), .Z(n23960) );
  AND U24080 ( .A(n23961), .B(n23962), .Z(n23956) );
  NANDN U24081 ( .A(n23963), .B(n23964), .Z(n23962) );
  NANDN U24082 ( .A(n23965), .B(n23966), .Z(n23964) );
  NANDN U24083 ( .A(n23966), .B(n23965), .Z(n23961) );
  ANDN U24084 ( .B(B[193]), .A(n54), .Z(n23958) );
  XNOR U24085 ( .A(n23753), .B(n23967), .Z(n23959) );
  XNOR U24086 ( .A(n23752), .B(n23750), .Z(n23967) );
  AND U24087 ( .A(n23968), .B(n23969), .Z(n23750) );
  NANDN U24088 ( .A(n23970), .B(n23971), .Z(n23969) );
  OR U24089 ( .A(n23972), .B(n23973), .Z(n23971) );
  NAND U24090 ( .A(n23973), .B(n23972), .Z(n23968) );
  ANDN U24091 ( .B(B[194]), .A(n55), .Z(n23752) );
  XNOR U24092 ( .A(n23760), .B(n23974), .Z(n23753) );
  XNOR U24093 ( .A(n23759), .B(n23757), .Z(n23974) );
  AND U24094 ( .A(n23975), .B(n23976), .Z(n23757) );
  NANDN U24095 ( .A(n23977), .B(n23978), .Z(n23976) );
  NANDN U24096 ( .A(n23979), .B(n23980), .Z(n23978) );
  NANDN U24097 ( .A(n23980), .B(n23979), .Z(n23975) );
  ANDN U24098 ( .B(B[195]), .A(n56), .Z(n23759) );
  XNOR U24099 ( .A(n23767), .B(n23981), .Z(n23760) );
  XNOR U24100 ( .A(n23766), .B(n23764), .Z(n23981) );
  AND U24101 ( .A(n23982), .B(n23983), .Z(n23764) );
  NANDN U24102 ( .A(n23984), .B(n23985), .Z(n23983) );
  OR U24103 ( .A(n23986), .B(n23987), .Z(n23985) );
  NAND U24104 ( .A(n23987), .B(n23986), .Z(n23982) );
  ANDN U24105 ( .B(B[196]), .A(n57), .Z(n23766) );
  XNOR U24106 ( .A(n23774), .B(n23988), .Z(n23767) );
  XNOR U24107 ( .A(n23773), .B(n23771), .Z(n23988) );
  AND U24108 ( .A(n23989), .B(n23990), .Z(n23771) );
  NANDN U24109 ( .A(n23991), .B(n23992), .Z(n23990) );
  NANDN U24110 ( .A(n23993), .B(n23994), .Z(n23992) );
  NANDN U24111 ( .A(n23994), .B(n23993), .Z(n23989) );
  ANDN U24112 ( .B(B[197]), .A(n58), .Z(n23773) );
  XNOR U24113 ( .A(n23781), .B(n23995), .Z(n23774) );
  XNOR U24114 ( .A(n23780), .B(n23778), .Z(n23995) );
  AND U24115 ( .A(n23996), .B(n23997), .Z(n23778) );
  NANDN U24116 ( .A(n23998), .B(n23999), .Z(n23997) );
  OR U24117 ( .A(n24000), .B(n24001), .Z(n23999) );
  NAND U24118 ( .A(n24001), .B(n24000), .Z(n23996) );
  ANDN U24119 ( .B(B[198]), .A(n59), .Z(n23780) );
  XNOR U24120 ( .A(n23788), .B(n24002), .Z(n23781) );
  XNOR U24121 ( .A(n23787), .B(n23785), .Z(n24002) );
  AND U24122 ( .A(n24003), .B(n24004), .Z(n23785) );
  NANDN U24123 ( .A(n24005), .B(n24006), .Z(n24004) );
  NANDN U24124 ( .A(n24007), .B(n24008), .Z(n24006) );
  NANDN U24125 ( .A(n24008), .B(n24007), .Z(n24003) );
  ANDN U24126 ( .B(B[199]), .A(n60), .Z(n23787) );
  XNOR U24127 ( .A(n23795), .B(n24009), .Z(n23788) );
  XNOR U24128 ( .A(n23794), .B(n23792), .Z(n24009) );
  AND U24129 ( .A(n24010), .B(n24011), .Z(n23792) );
  NANDN U24130 ( .A(n24012), .B(n24013), .Z(n24011) );
  OR U24131 ( .A(n24014), .B(n24015), .Z(n24013) );
  NAND U24132 ( .A(n24015), .B(n24014), .Z(n24010) );
  ANDN U24133 ( .B(B[200]), .A(n61), .Z(n23794) );
  XNOR U24134 ( .A(n23802), .B(n24016), .Z(n23795) );
  XNOR U24135 ( .A(n23801), .B(n23799), .Z(n24016) );
  AND U24136 ( .A(n24017), .B(n24018), .Z(n23799) );
  NANDN U24137 ( .A(n24019), .B(n24020), .Z(n24018) );
  NANDN U24138 ( .A(n24021), .B(n24022), .Z(n24020) );
  NANDN U24139 ( .A(n24022), .B(n24021), .Z(n24017) );
  ANDN U24140 ( .B(B[201]), .A(n62), .Z(n23801) );
  XNOR U24141 ( .A(n23809), .B(n24023), .Z(n23802) );
  XNOR U24142 ( .A(n23808), .B(n23806), .Z(n24023) );
  AND U24143 ( .A(n24024), .B(n24025), .Z(n23806) );
  NANDN U24144 ( .A(n24026), .B(n24027), .Z(n24025) );
  OR U24145 ( .A(n24028), .B(n24029), .Z(n24027) );
  NAND U24146 ( .A(n24029), .B(n24028), .Z(n24024) );
  ANDN U24147 ( .B(B[202]), .A(n63), .Z(n23808) );
  XNOR U24148 ( .A(n23816), .B(n24030), .Z(n23809) );
  XNOR U24149 ( .A(n23815), .B(n23813), .Z(n24030) );
  AND U24150 ( .A(n24031), .B(n24032), .Z(n23813) );
  NANDN U24151 ( .A(n24033), .B(n24034), .Z(n24032) );
  NANDN U24152 ( .A(n24035), .B(n24036), .Z(n24034) );
  NANDN U24153 ( .A(n24036), .B(n24035), .Z(n24031) );
  ANDN U24154 ( .B(B[203]), .A(n64), .Z(n23815) );
  XNOR U24155 ( .A(n23823), .B(n24037), .Z(n23816) );
  XNOR U24156 ( .A(n23822), .B(n23820), .Z(n24037) );
  AND U24157 ( .A(n24038), .B(n24039), .Z(n23820) );
  NANDN U24158 ( .A(n24040), .B(n24041), .Z(n24039) );
  OR U24159 ( .A(n24042), .B(n24043), .Z(n24041) );
  NAND U24160 ( .A(n24043), .B(n24042), .Z(n24038) );
  ANDN U24161 ( .B(B[204]), .A(n65), .Z(n23822) );
  XNOR U24162 ( .A(n23830), .B(n24044), .Z(n23823) );
  XNOR U24163 ( .A(n23829), .B(n23827), .Z(n24044) );
  AND U24164 ( .A(n24045), .B(n24046), .Z(n23827) );
  NANDN U24165 ( .A(n24047), .B(n24048), .Z(n24046) );
  NANDN U24166 ( .A(n24049), .B(n24050), .Z(n24048) );
  NANDN U24167 ( .A(n24050), .B(n24049), .Z(n24045) );
  ANDN U24168 ( .B(B[205]), .A(n66), .Z(n23829) );
  XNOR U24169 ( .A(n23837), .B(n24051), .Z(n23830) );
  XNOR U24170 ( .A(n23836), .B(n23834), .Z(n24051) );
  AND U24171 ( .A(n24052), .B(n24053), .Z(n23834) );
  NANDN U24172 ( .A(n24054), .B(n24055), .Z(n24053) );
  OR U24173 ( .A(n24056), .B(n24057), .Z(n24055) );
  NAND U24174 ( .A(n24057), .B(n24056), .Z(n24052) );
  ANDN U24175 ( .B(B[206]), .A(n67), .Z(n23836) );
  XNOR U24176 ( .A(n23844), .B(n24058), .Z(n23837) );
  XNOR U24177 ( .A(n23843), .B(n23841), .Z(n24058) );
  AND U24178 ( .A(n24059), .B(n24060), .Z(n23841) );
  NANDN U24179 ( .A(n24061), .B(n24062), .Z(n24060) );
  NANDN U24180 ( .A(n24063), .B(n24064), .Z(n24062) );
  NANDN U24181 ( .A(n24064), .B(n24063), .Z(n24059) );
  ANDN U24182 ( .B(B[207]), .A(n68), .Z(n23843) );
  XNOR U24183 ( .A(n23851), .B(n24065), .Z(n23844) );
  XNOR U24184 ( .A(n23850), .B(n23848), .Z(n24065) );
  AND U24185 ( .A(n24066), .B(n24067), .Z(n23848) );
  NANDN U24186 ( .A(n24068), .B(n24069), .Z(n24067) );
  OR U24187 ( .A(n24070), .B(n24071), .Z(n24069) );
  NAND U24188 ( .A(n24071), .B(n24070), .Z(n24066) );
  ANDN U24189 ( .B(B[208]), .A(n69), .Z(n23850) );
  XNOR U24190 ( .A(n23858), .B(n24072), .Z(n23851) );
  XNOR U24191 ( .A(n23857), .B(n23855), .Z(n24072) );
  AND U24192 ( .A(n24073), .B(n24074), .Z(n23855) );
  NANDN U24193 ( .A(n24075), .B(n24076), .Z(n24074) );
  NANDN U24194 ( .A(n24077), .B(n24078), .Z(n24076) );
  NANDN U24195 ( .A(n24078), .B(n24077), .Z(n24073) );
  ANDN U24196 ( .B(B[209]), .A(n70), .Z(n23857) );
  XNOR U24197 ( .A(n23865), .B(n24079), .Z(n23858) );
  XNOR U24198 ( .A(n23864), .B(n23862), .Z(n24079) );
  AND U24199 ( .A(n24080), .B(n24081), .Z(n23862) );
  NANDN U24200 ( .A(n24082), .B(n24083), .Z(n24081) );
  OR U24201 ( .A(n24084), .B(n24085), .Z(n24083) );
  NAND U24202 ( .A(n24085), .B(n24084), .Z(n24080) );
  ANDN U24203 ( .B(B[210]), .A(n71), .Z(n23864) );
  XNOR U24204 ( .A(n23872), .B(n24086), .Z(n23865) );
  XNOR U24205 ( .A(n23871), .B(n23869), .Z(n24086) );
  AND U24206 ( .A(n24087), .B(n24088), .Z(n23869) );
  NANDN U24207 ( .A(n24089), .B(n24090), .Z(n24088) );
  NANDN U24208 ( .A(n24091), .B(n24092), .Z(n24090) );
  NANDN U24209 ( .A(n24092), .B(n24091), .Z(n24087) );
  ANDN U24210 ( .B(B[211]), .A(n72), .Z(n23871) );
  XNOR U24211 ( .A(n23879), .B(n24093), .Z(n23872) );
  XNOR U24212 ( .A(n23878), .B(n23876), .Z(n24093) );
  AND U24213 ( .A(n24094), .B(n24095), .Z(n23876) );
  NANDN U24214 ( .A(n24096), .B(n24097), .Z(n24095) );
  OR U24215 ( .A(n24098), .B(n24099), .Z(n24097) );
  NAND U24216 ( .A(n24099), .B(n24098), .Z(n24094) );
  ANDN U24217 ( .B(B[212]), .A(n73), .Z(n23878) );
  XNOR U24218 ( .A(n23886), .B(n24100), .Z(n23879) );
  XNOR U24219 ( .A(n23885), .B(n23883), .Z(n24100) );
  AND U24220 ( .A(n24101), .B(n24102), .Z(n23883) );
  NANDN U24221 ( .A(n24103), .B(n24104), .Z(n24102) );
  NANDN U24222 ( .A(n24105), .B(n24106), .Z(n24104) );
  NANDN U24223 ( .A(n24106), .B(n24105), .Z(n24101) );
  ANDN U24224 ( .B(B[213]), .A(n74), .Z(n23885) );
  XNOR U24225 ( .A(n23893), .B(n24107), .Z(n23886) );
  XNOR U24226 ( .A(n23892), .B(n23890), .Z(n24107) );
  AND U24227 ( .A(n24108), .B(n24109), .Z(n23890) );
  NANDN U24228 ( .A(n24110), .B(n24111), .Z(n24109) );
  OR U24229 ( .A(n24112), .B(n24113), .Z(n24111) );
  NAND U24230 ( .A(n24113), .B(n24112), .Z(n24108) );
  ANDN U24231 ( .B(B[214]), .A(n75), .Z(n23892) );
  XNOR U24232 ( .A(n23900), .B(n24114), .Z(n23893) );
  XNOR U24233 ( .A(n23899), .B(n23897), .Z(n24114) );
  AND U24234 ( .A(n24115), .B(n24116), .Z(n23897) );
  NANDN U24235 ( .A(n24117), .B(n24118), .Z(n24116) );
  NANDN U24236 ( .A(n24119), .B(n24120), .Z(n24118) );
  NANDN U24237 ( .A(n24120), .B(n24119), .Z(n24115) );
  ANDN U24238 ( .B(B[215]), .A(n76), .Z(n23899) );
  XNOR U24239 ( .A(n23907), .B(n24121), .Z(n23900) );
  XNOR U24240 ( .A(n23906), .B(n23904), .Z(n24121) );
  AND U24241 ( .A(n24122), .B(n24123), .Z(n23904) );
  NANDN U24242 ( .A(n24124), .B(n24125), .Z(n24123) );
  OR U24243 ( .A(n24126), .B(n24127), .Z(n24125) );
  NAND U24244 ( .A(n24127), .B(n24126), .Z(n24122) );
  ANDN U24245 ( .B(B[216]), .A(n77), .Z(n23906) );
  XNOR U24246 ( .A(n23914), .B(n24128), .Z(n23907) );
  XNOR U24247 ( .A(n23913), .B(n23911), .Z(n24128) );
  AND U24248 ( .A(n24129), .B(n24130), .Z(n23911) );
  NANDN U24249 ( .A(n24131), .B(n24132), .Z(n24130) );
  NANDN U24250 ( .A(n24133), .B(n24134), .Z(n24132) );
  NANDN U24251 ( .A(n24134), .B(n24133), .Z(n24129) );
  ANDN U24252 ( .B(B[217]), .A(n78), .Z(n23913) );
  XNOR U24253 ( .A(n23921), .B(n24135), .Z(n23914) );
  XNOR U24254 ( .A(n23920), .B(n23918), .Z(n24135) );
  AND U24255 ( .A(n24136), .B(n24137), .Z(n23918) );
  NANDN U24256 ( .A(n24138), .B(n24139), .Z(n24137) );
  OR U24257 ( .A(n24140), .B(n24141), .Z(n24139) );
  NAND U24258 ( .A(n24141), .B(n24140), .Z(n24136) );
  ANDN U24259 ( .B(B[218]), .A(n79), .Z(n23920) );
  XNOR U24260 ( .A(n23928), .B(n24142), .Z(n23921) );
  XNOR U24261 ( .A(n23927), .B(n23925), .Z(n24142) );
  AND U24262 ( .A(n24143), .B(n24144), .Z(n23925) );
  NANDN U24263 ( .A(n24145), .B(n24146), .Z(n24144) );
  NANDN U24264 ( .A(n24147), .B(n24148), .Z(n24146) );
  NANDN U24265 ( .A(n24148), .B(n24147), .Z(n24143) );
  ANDN U24266 ( .B(B[219]), .A(n80), .Z(n23927) );
  XNOR U24267 ( .A(n23935), .B(n24149), .Z(n23928) );
  XNOR U24268 ( .A(n23934), .B(n23932), .Z(n24149) );
  AND U24269 ( .A(n24150), .B(n24151), .Z(n23932) );
  NANDN U24270 ( .A(n24152), .B(n24153), .Z(n24151) );
  OR U24271 ( .A(n24154), .B(n24155), .Z(n24153) );
  NAND U24272 ( .A(n24155), .B(n24154), .Z(n24150) );
  ANDN U24273 ( .B(B[220]), .A(n81), .Z(n23934) );
  XNOR U24274 ( .A(n23942), .B(n24156), .Z(n23935) );
  XNOR U24275 ( .A(n23941), .B(n23939), .Z(n24156) );
  AND U24276 ( .A(n24157), .B(n24158), .Z(n23939) );
  NANDN U24277 ( .A(n24159), .B(n24160), .Z(n24158) );
  NAND U24278 ( .A(n24161), .B(n24162), .Z(n24160) );
  ANDN U24279 ( .B(B[221]), .A(n82), .Z(n23941) );
  XOR U24280 ( .A(n23948), .B(n24163), .Z(n23942) );
  XNOR U24281 ( .A(n23946), .B(n23949), .Z(n24163) );
  NAND U24282 ( .A(A[2]), .B(B[222]), .Z(n23949) );
  NANDN U24283 ( .A(n24164), .B(n24165), .Z(n23946) );
  AND U24284 ( .A(A[0]), .B(B[223]), .Z(n24165) );
  XNOR U24285 ( .A(n23951), .B(n24166), .Z(n23948) );
  NAND U24286 ( .A(A[0]), .B(B[224]), .Z(n24166) );
  NAND U24287 ( .A(B[223]), .B(A[1]), .Z(n23951) );
  NAND U24288 ( .A(n24167), .B(n24168), .Z(n348) );
  NANDN U24289 ( .A(n24169), .B(n24170), .Z(n24168) );
  OR U24290 ( .A(n24171), .B(n24172), .Z(n24170) );
  NAND U24291 ( .A(n24172), .B(n24171), .Z(n24167) );
  XOR U24292 ( .A(n350), .B(n349), .Z(\A1[221] ) );
  XOR U24293 ( .A(n24172), .B(n24173), .Z(n349) );
  XNOR U24294 ( .A(n24171), .B(n24169), .Z(n24173) );
  AND U24295 ( .A(n24174), .B(n24175), .Z(n24169) );
  NANDN U24296 ( .A(n24176), .B(n24177), .Z(n24175) );
  NANDN U24297 ( .A(n24178), .B(n24179), .Z(n24177) );
  NANDN U24298 ( .A(n24179), .B(n24178), .Z(n24174) );
  ANDN U24299 ( .B(B[192]), .A(n54), .Z(n24171) );
  XNOR U24300 ( .A(n23966), .B(n24180), .Z(n24172) );
  XNOR U24301 ( .A(n23965), .B(n23963), .Z(n24180) );
  AND U24302 ( .A(n24181), .B(n24182), .Z(n23963) );
  NANDN U24303 ( .A(n24183), .B(n24184), .Z(n24182) );
  OR U24304 ( .A(n24185), .B(n24186), .Z(n24184) );
  NAND U24305 ( .A(n24186), .B(n24185), .Z(n24181) );
  ANDN U24306 ( .B(B[193]), .A(n55), .Z(n23965) );
  XNOR U24307 ( .A(n23973), .B(n24187), .Z(n23966) );
  XNOR U24308 ( .A(n23972), .B(n23970), .Z(n24187) );
  AND U24309 ( .A(n24188), .B(n24189), .Z(n23970) );
  NANDN U24310 ( .A(n24190), .B(n24191), .Z(n24189) );
  NANDN U24311 ( .A(n24192), .B(n24193), .Z(n24191) );
  NANDN U24312 ( .A(n24193), .B(n24192), .Z(n24188) );
  ANDN U24313 ( .B(B[194]), .A(n56), .Z(n23972) );
  XNOR U24314 ( .A(n23980), .B(n24194), .Z(n23973) );
  XNOR U24315 ( .A(n23979), .B(n23977), .Z(n24194) );
  AND U24316 ( .A(n24195), .B(n24196), .Z(n23977) );
  NANDN U24317 ( .A(n24197), .B(n24198), .Z(n24196) );
  OR U24318 ( .A(n24199), .B(n24200), .Z(n24198) );
  NAND U24319 ( .A(n24200), .B(n24199), .Z(n24195) );
  ANDN U24320 ( .B(B[195]), .A(n57), .Z(n23979) );
  XNOR U24321 ( .A(n23987), .B(n24201), .Z(n23980) );
  XNOR U24322 ( .A(n23986), .B(n23984), .Z(n24201) );
  AND U24323 ( .A(n24202), .B(n24203), .Z(n23984) );
  NANDN U24324 ( .A(n24204), .B(n24205), .Z(n24203) );
  NANDN U24325 ( .A(n24206), .B(n24207), .Z(n24205) );
  NANDN U24326 ( .A(n24207), .B(n24206), .Z(n24202) );
  ANDN U24327 ( .B(B[196]), .A(n58), .Z(n23986) );
  XNOR U24328 ( .A(n23994), .B(n24208), .Z(n23987) );
  XNOR U24329 ( .A(n23993), .B(n23991), .Z(n24208) );
  AND U24330 ( .A(n24209), .B(n24210), .Z(n23991) );
  NANDN U24331 ( .A(n24211), .B(n24212), .Z(n24210) );
  OR U24332 ( .A(n24213), .B(n24214), .Z(n24212) );
  NAND U24333 ( .A(n24214), .B(n24213), .Z(n24209) );
  ANDN U24334 ( .B(B[197]), .A(n59), .Z(n23993) );
  XNOR U24335 ( .A(n24001), .B(n24215), .Z(n23994) );
  XNOR U24336 ( .A(n24000), .B(n23998), .Z(n24215) );
  AND U24337 ( .A(n24216), .B(n24217), .Z(n23998) );
  NANDN U24338 ( .A(n24218), .B(n24219), .Z(n24217) );
  NANDN U24339 ( .A(n24220), .B(n24221), .Z(n24219) );
  NANDN U24340 ( .A(n24221), .B(n24220), .Z(n24216) );
  ANDN U24341 ( .B(B[198]), .A(n60), .Z(n24000) );
  XNOR U24342 ( .A(n24008), .B(n24222), .Z(n24001) );
  XNOR U24343 ( .A(n24007), .B(n24005), .Z(n24222) );
  AND U24344 ( .A(n24223), .B(n24224), .Z(n24005) );
  NANDN U24345 ( .A(n24225), .B(n24226), .Z(n24224) );
  OR U24346 ( .A(n24227), .B(n24228), .Z(n24226) );
  NAND U24347 ( .A(n24228), .B(n24227), .Z(n24223) );
  ANDN U24348 ( .B(B[199]), .A(n61), .Z(n24007) );
  XNOR U24349 ( .A(n24015), .B(n24229), .Z(n24008) );
  XNOR U24350 ( .A(n24014), .B(n24012), .Z(n24229) );
  AND U24351 ( .A(n24230), .B(n24231), .Z(n24012) );
  NANDN U24352 ( .A(n24232), .B(n24233), .Z(n24231) );
  NANDN U24353 ( .A(n24234), .B(n24235), .Z(n24233) );
  NANDN U24354 ( .A(n24235), .B(n24234), .Z(n24230) );
  ANDN U24355 ( .B(B[200]), .A(n62), .Z(n24014) );
  XNOR U24356 ( .A(n24022), .B(n24236), .Z(n24015) );
  XNOR U24357 ( .A(n24021), .B(n24019), .Z(n24236) );
  AND U24358 ( .A(n24237), .B(n24238), .Z(n24019) );
  NANDN U24359 ( .A(n24239), .B(n24240), .Z(n24238) );
  OR U24360 ( .A(n24241), .B(n24242), .Z(n24240) );
  NAND U24361 ( .A(n24242), .B(n24241), .Z(n24237) );
  ANDN U24362 ( .B(B[201]), .A(n63), .Z(n24021) );
  XNOR U24363 ( .A(n24029), .B(n24243), .Z(n24022) );
  XNOR U24364 ( .A(n24028), .B(n24026), .Z(n24243) );
  AND U24365 ( .A(n24244), .B(n24245), .Z(n24026) );
  NANDN U24366 ( .A(n24246), .B(n24247), .Z(n24245) );
  NANDN U24367 ( .A(n24248), .B(n24249), .Z(n24247) );
  NANDN U24368 ( .A(n24249), .B(n24248), .Z(n24244) );
  ANDN U24369 ( .B(B[202]), .A(n64), .Z(n24028) );
  XNOR U24370 ( .A(n24036), .B(n24250), .Z(n24029) );
  XNOR U24371 ( .A(n24035), .B(n24033), .Z(n24250) );
  AND U24372 ( .A(n24251), .B(n24252), .Z(n24033) );
  NANDN U24373 ( .A(n24253), .B(n24254), .Z(n24252) );
  OR U24374 ( .A(n24255), .B(n24256), .Z(n24254) );
  NAND U24375 ( .A(n24256), .B(n24255), .Z(n24251) );
  ANDN U24376 ( .B(B[203]), .A(n65), .Z(n24035) );
  XNOR U24377 ( .A(n24043), .B(n24257), .Z(n24036) );
  XNOR U24378 ( .A(n24042), .B(n24040), .Z(n24257) );
  AND U24379 ( .A(n24258), .B(n24259), .Z(n24040) );
  NANDN U24380 ( .A(n24260), .B(n24261), .Z(n24259) );
  NANDN U24381 ( .A(n24262), .B(n24263), .Z(n24261) );
  NANDN U24382 ( .A(n24263), .B(n24262), .Z(n24258) );
  ANDN U24383 ( .B(B[204]), .A(n66), .Z(n24042) );
  XNOR U24384 ( .A(n24050), .B(n24264), .Z(n24043) );
  XNOR U24385 ( .A(n24049), .B(n24047), .Z(n24264) );
  AND U24386 ( .A(n24265), .B(n24266), .Z(n24047) );
  NANDN U24387 ( .A(n24267), .B(n24268), .Z(n24266) );
  OR U24388 ( .A(n24269), .B(n24270), .Z(n24268) );
  NAND U24389 ( .A(n24270), .B(n24269), .Z(n24265) );
  ANDN U24390 ( .B(B[205]), .A(n67), .Z(n24049) );
  XNOR U24391 ( .A(n24057), .B(n24271), .Z(n24050) );
  XNOR U24392 ( .A(n24056), .B(n24054), .Z(n24271) );
  AND U24393 ( .A(n24272), .B(n24273), .Z(n24054) );
  NANDN U24394 ( .A(n24274), .B(n24275), .Z(n24273) );
  NANDN U24395 ( .A(n24276), .B(n24277), .Z(n24275) );
  NANDN U24396 ( .A(n24277), .B(n24276), .Z(n24272) );
  ANDN U24397 ( .B(B[206]), .A(n68), .Z(n24056) );
  XNOR U24398 ( .A(n24064), .B(n24278), .Z(n24057) );
  XNOR U24399 ( .A(n24063), .B(n24061), .Z(n24278) );
  AND U24400 ( .A(n24279), .B(n24280), .Z(n24061) );
  NANDN U24401 ( .A(n24281), .B(n24282), .Z(n24280) );
  OR U24402 ( .A(n24283), .B(n24284), .Z(n24282) );
  NAND U24403 ( .A(n24284), .B(n24283), .Z(n24279) );
  ANDN U24404 ( .B(B[207]), .A(n69), .Z(n24063) );
  XNOR U24405 ( .A(n24071), .B(n24285), .Z(n24064) );
  XNOR U24406 ( .A(n24070), .B(n24068), .Z(n24285) );
  AND U24407 ( .A(n24286), .B(n24287), .Z(n24068) );
  NANDN U24408 ( .A(n24288), .B(n24289), .Z(n24287) );
  NANDN U24409 ( .A(n24290), .B(n24291), .Z(n24289) );
  NANDN U24410 ( .A(n24291), .B(n24290), .Z(n24286) );
  ANDN U24411 ( .B(B[208]), .A(n70), .Z(n24070) );
  XNOR U24412 ( .A(n24078), .B(n24292), .Z(n24071) );
  XNOR U24413 ( .A(n24077), .B(n24075), .Z(n24292) );
  AND U24414 ( .A(n24293), .B(n24294), .Z(n24075) );
  NANDN U24415 ( .A(n24295), .B(n24296), .Z(n24294) );
  OR U24416 ( .A(n24297), .B(n24298), .Z(n24296) );
  NAND U24417 ( .A(n24298), .B(n24297), .Z(n24293) );
  ANDN U24418 ( .B(B[209]), .A(n71), .Z(n24077) );
  XNOR U24419 ( .A(n24085), .B(n24299), .Z(n24078) );
  XNOR U24420 ( .A(n24084), .B(n24082), .Z(n24299) );
  AND U24421 ( .A(n24300), .B(n24301), .Z(n24082) );
  NANDN U24422 ( .A(n24302), .B(n24303), .Z(n24301) );
  NANDN U24423 ( .A(n24304), .B(n24305), .Z(n24303) );
  NANDN U24424 ( .A(n24305), .B(n24304), .Z(n24300) );
  ANDN U24425 ( .B(B[210]), .A(n72), .Z(n24084) );
  XNOR U24426 ( .A(n24092), .B(n24306), .Z(n24085) );
  XNOR U24427 ( .A(n24091), .B(n24089), .Z(n24306) );
  AND U24428 ( .A(n24307), .B(n24308), .Z(n24089) );
  NANDN U24429 ( .A(n24309), .B(n24310), .Z(n24308) );
  OR U24430 ( .A(n24311), .B(n24312), .Z(n24310) );
  NAND U24431 ( .A(n24312), .B(n24311), .Z(n24307) );
  ANDN U24432 ( .B(B[211]), .A(n73), .Z(n24091) );
  XNOR U24433 ( .A(n24099), .B(n24313), .Z(n24092) );
  XNOR U24434 ( .A(n24098), .B(n24096), .Z(n24313) );
  AND U24435 ( .A(n24314), .B(n24315), .Z(n24096) );
  NANDN U24436 ( .A(n24316), .B(n24317), .Z(n24315) );
  NANDN U24437 ( .A(n24318), .B(n24319), .Z(n24317) );
  NANDN U24438 ( .A(n24319), .B(n24318), .Z(n24314) );
  ANDN U24439 ( .B(B[212]), .A(n74), .Z(n24098) );
  XNOR U24440 ( .A(n24106), .B(n24320), .Z(n24099) );
  XNOR U24441 ( .A(n24105), .B(n24103), .Z(n24320) );
  AND U24442 ( .A(n24321), .B(n24322), .Z(n24103) );
  NANDN U24443 ( .A(n24323), .B(n24324), .Z(n24322) );
  OR U24444 ( .A(n24325), .B(n24326), .Z(n24324) );
  NAND U24445 ( .A(n24326), .B(n24325), .Z(n24321) );
  ANDN U24446 ( .B(B[213]), .A(n75), .Z(n24105) );
  XNOR U24447 ( .A(n24113), .B(n24327), .Z(n24106) );
  XNOR U24448 ( .A(n24112), .B(n24110), .Z(n24327) );
  AND U24449 ( .A(n24328), .B(n24329), .Z(n24110) );
  NANDN U24450 ( .A(n24330), .B(n24331), .Z(n24329) );
  NANDN U24451 ( .A(n24332), .B(n24333), .Z(n24331) );
  NANDN U24452 ( .A(n24333), .B(n24332), .Z(n24328) );
  ANDN U24453 ( .B(B[214]), .A(n76), .Z(n24112) );
  XNOR U24454 ( .A(n24120), .B(n24334), .Z(n24113) );
  XNOR U24455 ( .A(n24119), .B(n24117), .Z(n24334) );
  AND U24456 ( .A(n24335), .B(n24336), .Z(n24117) );
  NANDN U24457 ( .A(n24337), .B(n24338), .Z(n24336) );
  OR U24458 ( .A(n24339), .B(n24340), .Z(n24338) );
  NAND U24459 ( .A(n24340), .B(n24339), .Z(n24335) );
  ANDN U24460 ( .B(B[215]), .A(n77), .Z(n24119) );
  XNOR U24461 ( .A(n24127), .B(n24341), .Z(n24120) );
  XNOR U24462 ( .A(n24126), .B(n24124), .Z(n24341) );
  AND U24463 ( .A(n24342), .B(n24343), .Z(n24124) );
  NANDN U24464 ( .A(n24344), .B(n24345), .Z(n24343) );
  NANDN U24465 ( .A(n24346), .B(n24347), .Z(n24345) );
  NANDN U24466 ( .A(n24347), .B(n24346), .Z(n24342) );
  ANDN U24467 ( .B(B[216]), .A(n78), .Z(n24126) );
  XNOR U24468 ( .A(n24134), .B(n24348), .Z(n24127) );
  XNOR U24469 ( .A(n24133), .B(n24131), .Z(n24348) );
  AND U24470 ( .A(n24349), .B(n24350), .Z(n24131) );
  NANDN U24471 ( .A(n24351), .B(n24352), .Z(n24350) );
  OR U24472 ( .A(n24353), .B(n24354), .Z(n24352) );
  NAND U24473 ( .A(n24354), .B(n24353), .Z(n24349) );
  ANDN U24474 ( .B(B[217]), .A(n79), .Z(n24133) );
  XNOR U24475 ( .A(n24141), .B(n24355), .Z(n24134) );
  XNOR U24476 ( .A(n24140), .B(n24138), .Z(n24355) );
  AND U24477 ( .A(n24356), .B(n24357), .Z(n24138) );
  NANDN U24478 ( .A(n24358), .B(n24359), .Z(n24357) );
  NANDN U24479 ( .A(n24360), .B(n24361), .Z(n24359) );
  NANDN U24480 ( .A(n24361), .B(n24360), .Z(n24356) );
  ANDN U24481 ( .B(B[218]), .A(n80), .Z(n24140) );
  XNOR U24482 ( .A(n24148), .B(n24362), .Z(n24141) );
  XNOR U24483 ( .A(n24147), .B(n24145), .Z(n24362) );
  AND U24484 ( .A(n24363), .B(n24364), .Z(n24145) );
  NANDN U24485 ( .A(n24365), .B(n24366), .Z(n24364) );
  OR U24486 ( .A(n24367), .B(n24368), .Z(n24366) );
  NAND U24487 ( .A(n24368), .B(n24367), .Z(n24363) );
  ANDN U24488 ( .B(B[219]), .A(n81), .Z(n24147) );
  XNOR U24489 ( .A(n24155), .B(n24369), .Z(n24148) );
  XNOR U24490 ( .A(n24154), .B(n24152), .Z(n24369) );
  AND U24491 ( .A(n24370), .B(n24371), .Z(n24152) );
  NANDN U24492 ( .A(n24372), .B(n24373), .Z(n24371) );
  NAND U24493 ( .A(n24374), .B(n24375), .Z(n24373) );
  ANDN U24494 ( .B(B[220]), .A(n82), .Z(n24154) );
  XOR U24495 ( .A(n24161), .B(n24376), .Z(n24155) );
  XNOR U24496 ( .A(n24159), .B(n24162), .Z(n24376) );
  NAND U24497 ( .A(A[2]), .B(B[221]), .Z(n24162) );
  NANDN U24498 ( .A(n24377), .B(n24378), .Z(n24159) );
  AND U24499 ( .A(A[0]), .B(B[222]), .Z(n24378) );
  XNOR U24500 ( .A(n24164), .B(n24379), .Z(n24161) );
  NAND U24501 ( .A(A[0]), .B(B[223]), .Z(n24379) );
  NAND U24502 ( .A(B[222]), .B(A[1]), .Z(n24164) );
  NAND U24503 ( .A(n24380), .B(n24381), .Z(n350) );
  NANDN U24504 ( .A(n24382), .B(n24383), .Z(n24381) );
  OR U24505 ( .A(n24384), .B(n24385), .Z(n24383) );
  NAND U24506 ( .A(n24385), .B(n24384), .Z(n24380) );
  XOR U24507 ( .A(n352), .B(n351), .Z(\A1[220] ) );
  XOR U24508 ( .A(n24385), .B(n24386), .Z(n351) );
  XNOR U24509 ( .A(n24384), .B(n24382), .Z(n24386) );
  AND U24510 ( .A(n24387), .B(n24388), .Z(n24382) );
  NANDN U24511 ( .A(n24389), .B(n24390), .Z(n24388) );
  NANDN U24512 ( .A(n24391), .B(n24392), .Z(n24390) );
  NANDN U24513 ( .A(n24392), .B(n24391), .Z(n24387) );
  ANDN U24514 ( .B(B[191]), .A(n54), .Z(n24384) );
  XNOR U24515 ( .A(n24179), .B(n24393), .Z(n24385) );
  XNOR U24516 ( .A(n24178), .B(n24176), .Z(n24393) );
  AND U24517 ( .A(n24394), .B(n24395), .Z(n24176) );
  NANDN U24518 ( .A(n24396), .B(n24397), .Z(n24395) );
  OR U24519 ( .A(n24398), .B(n24399), .Z(n24397) );
  NAND U24520 ( .A(n24399), .B(n24398), .Z(n24394) );
  ANDN U24521 ( .B(B[192]), .A(n55), .Z(n24178) );
  XNOR U24522 ( .A(n24186), .B(n24400), .Z(n24179) );
  XNOR U24523 ( .A(n24185), .B(n24183), .Z(n24400) );
  AND U24524 ( .A(n24401), .B(n24402), .Z(n24183) );
  NANDN U24525 ( .A(n24403), .B(n24404), .Z(n24402) );
  NANDN U24526 ( .A(n24405), .B(n24406), .Z(n24404) );
  NANDN U24527 ( .A(n24406), .B(n24405), .Z(n24401) );
  ANDN U24528 ( .B(B[193]), .A(n56), .Z(n24185) );
  XNOR U24529 ( .A(n24193), .B(n24407), .Z(n24186) );
  XNOR U24530 ( .A(n24192), .B(n24190), .Z(n24407) );
  AND U24531 ( .A(n24408), .B(n24409), .Z(n24190) );
  NANDN U24532 ( .A(n24410), .B(n24411), .Z(n24409) );
  OR U24533 ( .A(n24412), .B(n24413), .Z(n24411) );
  NAND U24534 ( .A(n24413), .B(n24412), .Z(n24408) );
  ANDN U24535 ( .B(B[194]), .A(n57), .Z(n24192) );
  XNOR U24536 ( .A(n24200), .B(n24414), .Z(n24193) );
  XNOR U24537 ( .A(n24199), .B(n24197), .Z(n24414) );
  AND U24538 ( .A(n24415), .B(n24416), .Z(n24197) );
  NANDN U24539 ( .A(n24417), .B(n24418), .Z(n24416) );
  NANDN U24540 ( .A(n24419), .B(n24420), .Z(n24418) );
  NANDN U24541 ( .A(n24420), .B(n24419), .Z(n24415) );
  ANDN U24542 ( .B(B[195]), .A(n58), .Z(n24199) );
  XNOR U24543 ( .A(n24207), .B(n24421), .Z(n24200) );
  XNOR U24544 ( .A(n24206), .B(n24204), .Z(n24421) );
  AND U24545 ( .A(n24422), .B(n24423), .Z(n24204) );
  NANDN U24546 ( .A(n24424), .B(n24425), .Z(n24423) );
  OR U24547 ( .A(n24426), .B(n24427), .Z(n24425) );
  NAND U24548 ( .A(n24427), .B(n24426), .Z(n24422) );
  ANDN U24549 ( .B(B[196]), .A(n59), .Z(n24206) );
  XNOR U24550 ( .A(n24214), .B(n24428), .Z(n24207) );
  XNOR U24551 ( .A(n24213), .B(n24211), .Z(n24428) );
  AND U24552 ( .A(n24429), .B(n24430), .Z(n24211) );
  NANDN U24553 ( .A(n24431), .B(n24432), .Z(n24430) );
  NANDN U24554 ( .A(n24433), .B(n24434), .Z(n24432) );
  NANDN U24555 ( .A(n24434), .B(n24433), .Z(n24429) );
  ANDN U24556 ( .B(B[197]), .A(n60), .Z(n24213) );
  XNOR U24557 ( .A(n24221), .B(n24435), .Z(n24214) );
  XNOR U24558 ( .A(n24220), .B(n24218), .Z(n24435) );
  AND U24559 ( .A(n24436), .B(n24437), .Z(n24218) );
  NANDN U24560 ( .A(n24438), .B(n24439), .Z(n24437) );
  OR U24561 ( .A(n24440), .B(n24441), .Z(n24439) );
  NAND U24562 ( .A(n24441), .B(n24440), .Z(n24436) );
  ANDN U24563 ( .B(B[198]), .A(n61), .Z(n24220) );
  XNOR U24564 ( .A(n24228), .B(n24442), .Z(n24221) );
  XNOR U24565 ( .A(n24227), .B(n24225), .Z(n24442) );
  AND U24566 ( .A(n24443), .B(n24444), .Z(n24225) );
  NANDN U24567 ( .A(n24445), .B(n24446), .Z(n24444) );
  NANDN U24568 ( .A(n24447), .B(n24448), .Z(n24446) );
  NANDN U24569 ( .A(n24448), .B(n24447), .Z(n24443) );
  ANDN U24570 ( .B(B[199]), .A(n62), .Z(n24227) );
  XNOR U24571 ( .A(n24235), .B(n24449), .Z(n24228) );
  XNOR U24572 ( .A(n24234), .B(n24232), .Z(n24449) );
  AND U24573 ( .A(n24450), .B(n24451), .Z(n24232) );
  NANDN U24574 ( .A(n24452), .B(n24453), .Z(n24451) );
  OR U24575 ( .A(n24454), .B(n24455), .Z(n24453) );
  NAND U24576 ( .A(n24455), .B(n24454), .Z(n24450) );
  ANDN U24577 ( .B(B[200]), .A(n63), .Z(n24234) );
  XNOR U24578 ( .A(n24242), .B(n24456), .Z(n24235) );
  XNOR U24579 ( .A(n24241), .B(n24239), .Z(n24456) );
  AND U24580 ( .A(n24457), .B(n24458), .Z(n24239) );
  NANDN U24581 ( .A(n24459), .B(n24460), .Z(n24458) );
  NANDN U24582 ( .A(n24461), .B(n24462), .Z(n24460) );
  NANDN U24583 ( .A(n24462), .B(n24461), .Z(n24457) );
  ANDN U24584 ( .B(B[201]), .A(n64), .Z(n24241) );
  XNOR U24585 ( .A(n24249), .B(n24463), .Z(n24242) );
  XNOR U24586 ( .A(n24248), .B(n24246), .Z(n24463) );
  AND U24587 ( .A(n24464), .B(n24465), .Z(n24246) );
  NANDN U24588 ( .A(n24466), .B(n24467), .Z(n24465) );
  OR U24589 ( .A(n24468), .B(n24469), .Z(n24467) );
  NAND U24590 ( .A(n24469), .B(n24468), .Z(n24464) );
  ANDN U24591 ( .B(B[202]), .A(n65), .Z(n24248) );
  XNOR U24592 ( .A(n24256), .B(n24470), .Z(n24249) );
  XNOR U24593 ( .A(n24255), .B(n24253), .Z(n24470) );
  AND U24594 ( .A(n24471), .B(n24472), .Z(n24253) );
  NANDN U24595 ( .A(n24473), .B(n24474), .Z(n24472) );
  NANDN U24596 ( .A(n24475), .B(n24476), .Z(n24474) );
  NANDN U24597 ( .A(n24476), .B(n24475), .Z(n24471) );
  ANDN U24598 ( .B(B[203]), .A(n66), .Z(n24255) );
  XNOR U24599 ( .A(n24263), .B(n24477), .Z(n24256) );
  XNOR U24600 ( .A(n24262), .B(n24260), .Z(n24477) );
  AND U24601 ( .A(n24478), .B(n24479), .Z(n24260) );
  NANDN U24602 ( .A(n24480), .B(n24481), .Z(n24479) );
  OR U24603 ( .A(n24482), .B(n24483), .Z(n24481) );
  NAND U24604 ( .A(n24483), .B(n24482), .Z(n24478) );
  ANDN U24605 ( .B(B[204]), .A(n67), .Z(n24262) );
  XNOR U24606 ( .A(n24270), .B(n24484), .Z(n24263) );
  XNOR U24607 ( .A(n24269), .B(n24267), .Z(n24484) );
  AND U24608 ( .A(n24485), .B(n24486), .Z(n24267) );
  NANDN U24609 ( .A(n24487), .B(n24488), .Z(n24486) );
  NANDN U24610 ( .A(n24489), .B(n24490), .Z(n24488) );
  NANDN U24611 ( .A(n24490), .B(n24489), .Z(n24485) );
  ANDN U24612 ( .B(B[205]), .A(n68), .Z(n24269) );
  XNOR U24613 ( .A(n24277), .B(n24491), .Z(n24270) );
  XNOR U24614 ( .A(n24276), .B(n24274), .Z(n24491) );
  AND U24615 ( .A(n24492), .B(n24493), .Z(n24274) );
  NANDN U24616 ( .A(n24494), .B(n24495), .Z(n24493) );
  OR U24617 ( .A(n24496), .B(n24497), .Z(n24495) );
  NAND U24618 ( .A(n24497), .B(n24496), .Z(n24492) );
  ANDN U24619 ( .B(B[206]), .A(n69), .Z(n24276) );
  XNOR U24620 ( .A(n24284), .B(n24498), .Z(n24277) );
  XNOR U24621 ( .A(n24283), .B(n24281), .Z(n24498) );
  AND U24622 ( .A(n24499), .B(n24500), .Z(n24281) );
  NANDN U24623 ( .A(n24501), .B(n24502), .Z(n24500) );
  NANDN U24624 ( .A(n24503), .B(n24504), .Z(n24502) );
  NANDN U24625 ( .A(n24504), .B(n24503), .Z(n24499) );
  ANDN U24626 ( .B(B[207]), .A(n70), .Z(n24283) );
  XNOR U24627 ( .A(n24291), .B(n24505), .Z(n24284) );
  XNOR U24628 ( .A(n24290), .B(n24288), .Z(n24505) );
  AND U24629 ( .A(n24506), .B(n24507), .Z(n24288) );
  NANDN U24630 ( .A(n24508), .B(n24509), .Z(n24507) );
  OR U24631 ( .A(n24510), .B(n24511), .Z(n24509) );
  NAND U24632 ( .A(n24511), .B(n24510), .Z(n24506) );
  ANDN U24633 ( .B(B[208]), .A(n71), .Z(n24290) );
  XNOR U24634 ( .A(n24298), .B(n24512), .Z(n24291) );
  XNOR U24635 ( .A(n24297), .B(n24295), .Z(n24512) );
  AND U24636 ( .A(n24513), .B(n24514), .Z(n24295) );
  NANDN U24637 ( .A(n24515), .B(n24516), .Z(n24514) );
  NANDN U24638 ( .A(n24517), .B(n24518), .Z(n24516) );
  NANDN U24639 ( .A(n24518), .B(n24517), .Z(n24513) );
  ANDN U24640 ( .B(B[209]), .A(n72), .Z(n24297) );
  XNOR U24641 ( .A(n24305), .B(n24519), .Z(n24298) );
  XNOR U24642 ( .A(n24304), .B(n24302), .Z(n24519) );
  AND U24643 ( .A(n24520), .B(n24521), .Z(n24302) );
  NANDN U24644 ( .A(n24522), .B(n24523), .Z(n24521) );
  OR U24645 ( .A(n24524), .B(n24525), .Z(n24523) );
  NAND U24646 ( .A(n24525), .B(n24524), .Z(n24520) );
  ANDN U24647 ( .B(B[210]), .A(n73), .Z(n24304) );
  XNOR U24648 ( .A(n24312), .B(n24526), .Z(n24305) );
  XNOR U24649 ( .A(n24311), .B(n24309), .Z(n24526) );
  AND U24650 ( .A(n24527), .B(n24528), .Z(n24309) );
  NANDN U24651 ( .A(n24529), .B(n24530), .Z(n24528) );
  NANDN U24652 ( .A(n24531), .B(n24532), .Z(n24530) );
  NANDN U24653 ( .A(n24532), .B(n24531), .Z(n24527) );
  ANDN U24654 ( .B(B[211]), .A(n74), .Z(n24311) );
  XNOR U24655 ( .A(n24319), .B(n24533), .Z(n24312) );
  XNOR U24656 ( .A(n24318), .B(n24316), .Z(n24533) );
  AND U24657 ( .A(n24534), .B(n24535), .Z(n24316) );
  NANDN U24658 ( .A(n24536), .B(n24537), .Z(n24535) );
  OR U24659 ( .A(n24538), .B(n24539), .Z(n24537) );
  NAND U24660 ( .A(n24539), .B(n24538), .Z(n24534) );
  ANDN U24661 ( .B(B[212]), .A(n75), .Z(n24318) );
  XNOR U24662 ( .A(n24326), .B(n24540), .Z(n24319) );
  XNOR U24663 ( .A(n24325), .B(n24323), .Z(n24540) );
  AND U24664 ( .A(n24541), .B(n24542), .Z(n24323) );
  NANDN U24665 ( .A(n24543), .B(n24544), .Z(n24542) );
  NANDN U24666 ( .A(n24545), .B(n24546), .Z(n24544) );
  NANDN U24667 ( .A(n24546), .B(n24545), .Z(n24541) );
  ANDN U24668 ( .B(B[213]), .A(n76), .Z(n24325) );
  XNOR U24669 ( .A(n24333), .B(n24547), .Z(n24326) );
  XNOR U24670 ( .A(n24332), .B(n24330), .Z(n24547) );
  AND U24671 ( .A(n24548), .B(n24549), .Z(n24330) );
  NANDN U24672 ( .A(n24550), .B(n24551), .Z(n24549) );
  OR U24673 ( .A(n24552), .B(n24553), .Z(n24551) );
  NAND U24674 ( .A(n24553), .B(n24552), .Z(n24548) );
  ANDN U24675 ( .B(B[214]), .A(n77), .Z(n24332) );
  XNOR U24676 ( .A(n24340), .B(n24554), .Z(n24333) );
  XNOR U24677 ( .A(n24339), .B(n24337), .Z(n24554) );
  AND U24678 ( .A(n24555), .B(n24556), .Z(n24337) );
  NANDN U24679 ( .A(n24557), .B(n24558), .Z(n24556) );
  NANDN U24680 ( .A(n24559), .B(n24560), .Z(n24558) );
  NANDN U24681 ( .A(n24560), .B(n24559), .Z(n24555) );
  ANDN U24682 ( .B(B[215]), .A(n78), .Z(n24339) );
  XNOR U24683 ( .A(n24347), .B(n24561), .Z(n24340) );
  XNOR U24684 ( .A(n24346), .B(n24344), .Z(n24561) );
  AND U24685 ( .A(n24562), .B(n24563), .Z(n24344) );
  NANDN U24686 ( .A(n24564), .B(n24565), .Z(n24563) );
  OR U24687 ( .A(n24566), .B(n24567), .Z(n24565) );
  NAND U24688 ( .A(n24567), .B(n24566), .Z(n24562) );
  ANDN U24689 ( .B(B[216]), .A(n79), .Z(n24346) );
  XNOR U24690 ( .A(n24354), .B(n24568), .Z(n24347) );
  XNOR U24691 ( .A(n24353), .B(n24351), .Z(n24568) );
  AND U24692 ( .A(n24569), .B(n24570), .Z(n24351) );
  NANDN U24693 ( .A(n24571), .B(n24572), .Z(n24570) );
  NANDN U24694 ( .A(n24573), .B(n24574), .Z(n24572) );
  NANDN U24695 ( .A(n24574), .B(n24573), .Z(n24569) );
  ANDN U24696 ( .B(B[217]), .A(n80), .Z(n24353) );
  XNOR U24697 ( .A(n24361), .B(n24575), .Z(n24354) );
  XNOR U24698 ( .A(n24360), .B(n24358), .Z(n24575) );
  AND U24699 ( .A(n24576), .B(n24577), .Z(n24358) );
  NANDN U24700 ( .A(n24578), .B(n24579), .Z(n24577) );
  OR U24701 ( .A(n24580), .B(n24581), .Z(n24579) );
  NAND U24702 ( .A(n24581), .B(n24580), .Z(n24576) );
  ANDN U24703 ( .B(B[218]), .A(n81), .Z(n24360) );
  XNOR U24704 ( .A(n24368), .B(n24582), .Z(n24361) );
  XNOR U24705 ( .A(n24367), .B(n24365), .Z(n24582) );
  AND U24706 ( .A(n24583), .B(n24584), .Z(n24365) );
  NANDN U24707 ( .A(n24585), .B(n24586), .Z(n24584) );
  NAND U24708 ( .A(n24587), .B(n24588), .Z(n24586) );
  ANDN U24709 ( .B(B[219]), .A(n82), .Z(n24367) );
  XOR U24710 ( .A(n24374), .B(n24589), .Z(n24368) );
  XNOR U24711 ( .A(n24372), .B(n24375), .Z(n24589) );
  NAND U24712 ( .A(A[2]), .B(B[220]), .Z(n24375) );
  NANDN U24713 ( .A(n24590), .B(n24591), .Z(n24372) );
  AND U24714 ( .A(A[0]), .B(B[221]), .Z(n24591) );
  XNOR U24715 ( .A(n24377), .B(n24592), .Z(n24374) );
  NAND U24716 ( .A(A[0]), .B(B[222]), .Z(n24592) );
  NAND U24717 ( .A(B[221]), .B(A[1]), .Z(n24377) );
  NAND U24718 ( .A(n24593), .B(n24594), .Z(n352) );
  NANDN U24719 ( .A(n24595), .B(n24596), .Z(n24594) );
  OR U24720 ( .A(n24597), .B(n24598), .Z(n24596) );
  NAND U24721 ( .A(n24598), .B(n24597), .Z(n24593) );
  XOR U24722 ( .A(n22317), .B(n24599), .Z(\A1[21] ) );
  XNOR U24723 ( .A(n22316), .B(n22314), .Z(n24599) );
  AND U24724 ( .A(n24600), .B(n24601), .Z(n22314) );
  NAND U24725 ( .A(n24602), .B(n24603), .Z(n24601) );
  NANDN U24726 ( .A(n24604), .B(n24605), .Z(n24602) );
  NANDN U24727 ( .A(n24605), .B(n24604), .Z(n24600) );
  ANDN U24728 ( .B(B[0]), .A(n62), .Z(n22316) );
  XNOR U24729 ( .A(n22324), .B(n24606), .Z(n22317) );
  XNOR U24730 ( .A(n22323), .B(n22321), .Z(n24606) );
  AND U24731 ( .A(n24607), .B(n24608), .Z(n22321) );
  NANDN U24732 ( .A(n24609), .B(n24610), .Z(n24608) );
  OR U24733 ( .A(n24611), .B(n24612), .Z(n24610) );
  NAND U24734 ( .A(n24612), .B(n24611), .Z(n24607) );
  ANDN U24735 ( .B(B[1]), .A(n63), .Z(n22323) );
  XNOR U24736 ( .A(n22331), .B(n24613), .Z(n22324) );
  XNOR U24737 ( .A(n22330), .B(n22328), .Z(n24613) );
  AND U24738 ( .A(n24614), .B(n24615), .Z(n22328) );
  NANDN U24739 ( .A(n24616), .B(n24617), .Z(n24615) );
  NANDN U24740 ( .A(n24618), .B(n24619), .Z(n24617) );
  NANDN U24741 ( .A(n24619), .B(n24618), .Z(n24614) );
  ANDN U24742 ( .B(B[2]), .A(n64), .Z(n22330) );
  XNOR U24743 ( .A(n22338), .B(n24620), .Z(n22331) );
  XNOR U24744 ( .A(n22337), .B(n22335), .Z(n24620) );
  AND U24745 ( .A(n24621), .B(n24622), .Z(n22335) );
  NANDN U24746 ( .A(n24623), .B(n24624), .Z(n24622) );
  OR U24747 ( .A(n24625), .B(n24626), .Z(n24624) );
  NAND U24748 ( .A(n24626), .B(n24625), .Z(n24621) );
  ANDN U24749 ( .B(B[3]), .A(n65), .Z(n22337) );
  XNOR U24750 ( .A(n22345), .B(n24627), .Z(n22338) );
  XNOR U24751 ( .A(n22344), .B(n22342), .Z(n24627) );
  AND U24752 ( .A(n24628), .B(n24629), .Z(n22342) );
  NANDN U24753 ( .A(n24630), .B(n24631), .Z(n24629) );
  NANDN U24754 ( .A(n24632), .B(n24633), .Z(n24631) );
  NANDN U24755 ( .A(n24633), .B(n24632), .Z(n24628) );
  ANDN U24756 ( .B(B[4]), .A(n66), .Z(n22344) );
  XNOR U24757 ( .A(n22352), .B(n24634), .Z(n22345) );
  XNOR U24758 ( .A(n22351), .B(n22349), .Z(n24634) );
  AND U24759 ( .A(n24635), .B(n24636), .Z(n22349) );
  NANDN U24760 ( .A(n24637), .B(n24638), .Z(n24636) );
  OR U24761 ( .A(n24639), .B(n24640), .Z(n24638) );
  NAND U24762 ( .A(n24640), .B(n24639), .Z(n24635) );
  ANDN U24763 ( .B(B[5]), .A(n67), .Z(n22351) );
  XNOR U24764 ( .A(n22359), .B(n24641), .Z(n22352) );
  XNOR U24765 ( .A(n22358), .B(n22356), .Z(n24641) );
  AND U24766 ( .A(n24642), .B(n24643), .Z(n22356) );
  NANDN U24767 ( .A(n24644), .B(n24645), .Z(n24643) );
  NANDN U24768 ( .A(n24646), .B(n24647), .Z(n24645) );
  NANDN U24769 ( .A(n24647), .B(n24646), .Z(n24642) );
  ANDN U24770 ( .B(B[6]), .A(n68), .Z(n22358) );
  XNOR U24771 ( .A(n22366), .B(n24648), .Z(n22359) );
  XNOR U24772 ( .A(n22365), .B(n22363), .Z(n24648) );
  AND U24773 ( .A(n24649), .B(n24650), .Z(n22363) );
  NANDN U24774 ( .A(n24651), .B(n24652), .Z(n24650) );
  OR U24775 ( .A(n24653), .B(n24654), .Z(n24652) );
  NAND U24776 ( .A(n24654), .B(n24653), .Z(n24649) );
  ANDN U24777 ( .B(B[7]), .A(n69), .Z(n22365) );
  XNOR U24778 ( .A(n22373), .B(n24655), .Z(n22366) );
  XNOR U24779 ( .A(n22372), .B(n22370), .Z(n24655) );
  AND U24780 ( .A(n24656), .B(n24657), .Z(n22370) );
  NANDN U24781 ( .A(n24658), .B(n24659), .Z(n24657) );
  NANDN U24782 ( .A(n24660), .B(n24661), .Z(n24659) );
  NANDN U24783 ( .A(n24661), .B(n24660), .Z(n24656) );
  ANDN U24784 ( .B(B[8]), .A(n70), .Z(n22372) );
  XNOR U24785 ( .A(n22380), .B(n24662), .Z(n22373) );
  XNOR U24786 ( .A(n22379), .B(n22377), .Z(n24662) );
  AND U24787 ( .A(n24663), .B(n24664), .Z(n22377) );
  NANDN U24788 ( .A(n24665), .B(n24666), .Z(n24664) );
  OR U24789 ( .A(n24667), .B(n24668), .Z(n24666) );
  NAND U24790 ( .A(n24668), .B(n24667), .Z(n24663) );
  ANDN U24791 ( .B(B[9]), .A(n71), .Z(n22379) );
  XNOR U24792 ( .A(n22387), .B(n24669), .Z(n22380) );
  XNOR U24793 ( .A(n22386), .B(n22384), .Z(n24669) );
  AND U24794 ( .A(n24670), .B(n24671), .Z(n22384) );
  NANDN U24795 ( .A(n24672), .B(n24673), .Z(n24671) );
  NANDN U24796 ( .A(n24674), .B(n24675), .Z(n24673) );
  NANDN U24797 ( .A(n24675), .B(n24674), .Z(n24670) );
  ANDN U24798 ( .B(B[10]), .A(n72), .Z(n22386) );
  XNOR U24799 ( .A(n22394), .B(n24676), .Z(n22387) );
  XNOR U24800 ( .A(n22393), .B(n22391), .Z(n24676) );
  AND U24801 ( .A(n24677), .B(n24678), .Z(n22391) );
  NANDN U24802 ( .A(n24679), .B(n24680), .Z(n24678) );
  OR U24803 ( .A(n24681), .B(n24682), .Z(n24680) );
  NAND U24804 ( .A(n24682), .B(n24681), .Z(n24677) );
  ANDN U24805 ( .B(B[11]), .A(n73), .Z(n22393) );
  XNOR U24806 ( .A(n22401), .B(n24683), .Z(n22394) );
  XNOR U24807 ( .A(n22400), .B(n22398), .Z(n24683) );
  AND U24808 ( .A(n24684), .B(n24685), .Z(n22398) );
  NANDN U24809 ( .A(n24686), .B(n24687), .Z(n24685) );
  NANDN U24810 ( .A(n24688), .B(n24689), .Z(n24687) );
  NANDN U24811 ( .A(n24689), .B(n24688), .Z(n24684) );
  ANDN U24812 ( .B(B[12]), .A(n74), .Z(n22400) );
  XNOR U24813 ( .A(n22408), .B(n24690), .Z(n22401) );
  XNOR U24814 ( .A(n22407), .B(n22405), .Z(n24690) );
  AND U24815 ( .A(n24691), .B(n24692), .Z(n22405) );
  NANDN U24816 ( .A(n24693), .B(n24694), .Z(n24692) );
  OR U24817 ( .A(n24695), .B(n24696), .Z(n24694) );
  NAND U24818 ( .A(n24696), .B(n24695), .Z(n24691) );
  ANDN U24819 ( .B(B[13]), .A(n75), .Z(n22407) );
  XNOR U24820 ( .A(n22415), .B(n24697), .Z(n22408) );
  XNOR U24821 ( .A(n22414), .B(n22412), .Z(n24697) );
  AND U24822 ( .A(n24698), .B(n24699), .Z(n22412) );
  NANDN U24823 ( .A(n24700), .B(n24701), .Z(n24699) );
  NANDN U24824 ( .A(n24702), .B(n24703), .Z(n24701) );
  NANDN U24825 ( .A(n24703), .B(n24702), .Z(n24698) );
  ANDN U24826 ( .B(B[14]), .A(n76), .Z(n22414) );
  XNOR U24827 ( .A(n22422), .B(n24704), .Z(n22415) );
  XNOR U24828 ( .A(n22421), .B(n22419), .Z(n24704) );
  AND U24829 ( .A(n24705), .B(n24706), .Z(n22419) );
  NANDN U24830 ( .A(n24707), .B(n24708), .Z(n24706) );
  OR U24831 ( .A(n24709), .B(n24710), .Z(n24708) );
  NAND U24832 ( .A(n24710), .B(n24709), .Z(n24705) );
  ANDN U24833 ( .B(B[15]), .A(n77), .Z(n22421) );
  XNOR U24834 ( .A(n22429), .B(n24711), .Z(n22422) );
  XNOR U24835 ( .A(n22428), .B(n22426), .Z(n24711) );
  AND U24836 ( .A(n24712), .B(n24713), .Z(n22426) );
  NANDN U24837 ( .A(n24714), .B(n24715), .Z(n24713) );
  NANDN U24838 ( .A(n24716), .B(n24717), .Z(n24715) );
  NANDN U24839 ( .A(n24717), .B(n24716), .Z(n24712) );
  ANDN U24840 ( .B(B[16]), .A(n78), .Z(n22428) );
  XNOR U24841 ( .A(n22436), .B(n24718), .Z(n22429) );
  XNOR U24842 ( .A(n22435), .B(n22433), .Z(n24718) );
  AND U24843 ( .A(n24719), .B(n24720), .Z(n22433) );
  NANDN U24844 ( .A(n24721), .B(n24722), .Z(n24720) );
  OR U24845 ( .A(n24723), .B(n24724), .Z(n24722) );
  NAND U24846 ( .A(n24724), .B(n24723), .Z(n24719) );
  ANDN U24847 ( .B(B[17]), .A(n79), .Z(n22435) );
  XNOR U24848 ( .A(n22443), .B(n24725), .Z(n22436) );
  XNOR U24849 ( .A(n22442), .B(n22440), .Z(n24725) );
  AND U24850 ( .A(n24726), .B(n24727), .Z(n22440) );
  NANDN U24851 ( .A(n24728), .B(n24729), .Z(n24727) );
  NANDN U24852 ( .A(n24730), .B(n24731), .Z(n24729) );
  NANDN U24853 ( .A(n24731), .B(n24730), .Z(n24726) );
  ANDN U24854 ( .B(B[18]), .A(n80), .Z(n22442) );
  XNOR U24855 ( .A(n22450), .B(n24732), .Z(n22443) );
  XNOR U24856 ( .A(n22449), .B(n22447), .Z(n24732) );
  AND U24857 ( .A(n24733), .B(n24734), .Z(n22447) );
  NANDN U24858 ( .A(n24735), .B(n24736), .Z(n24734) );
  OR U24859 ( .A(n24737), .B(n24738), .Z(n24736) );
  NAND U24860 ( .A(n24738), .B(n24737), .Z(n24733) );
  ANDN U24861 ( .B(B[19]), .A(n81), .Z(n22449) );
  XNOR U24862 ( .A(n22457), .B(n24739), .Z(n22450) );
  XNOR U24863 ( .A(n22456), .B(n22454), .Z(n24739) );
  AND U24864 ( .A(n24740), .B(n24741), .Z(n22454) );
  NANDN U24865 ( .A(n24742), .B(n24743), .Z(n24741) );
  NAND U24866 ( .A(n24744), .B(n24745), .Z(n24743) );
  ANDN U24867 ( .B(B[20]), .A(n82), .Z(n22456) );
  XOR U24868 ( .A(n22463), .B(n24746), .Z(n22457) );
  XNOR U24869 ( .A(n22461), .B(n22464), .Z(n24746) );
  NAND U24870 ( .A(A[2]), .B(B[21]), .Z(n22464) );
  NANDN U24871 ( .A(n24747), .B(n24748), .Z(n22461) );
  AND U24872 ( .A(A[0]), .B(B[22]), .Z(n24748) );
  XNOR U24873 ( .A(n22466), .B(n24749), .Z(n22463) );
  NAND U24874 ( .A(A[0]), .B(B[23]), .Z(n24749) );
  NAND U24875 ( .A(B[22]), .B(A[1]), .Z(n22466) );
  XOR U24876 ( .A(n354), .B(n353), .Z(\A1[219] ) );
  XOR U24877 ( .A(n24598), .B(n24750), .Z(n353) );
  XNOR U24878 ( .A(n24597), .B(n24595), .Z(n24750) );
  AND U24879 ( .A(n24751), .B(n24752), .Z(n24595) );
  NANDN U24880 ( .A(n24753), .B(n24754), .Z(n24752) );
  NANDN U24881 ( .A(n24755), .B(n24756), .Z(n24754) );
  NANDN U24882 ( .A(n24756), .B(n24755), .Z(n24751) );
  ANDN U24883 ( .B(B[190]), .A(n54), .Z(n24597) );
  XNOR U24884 ( .A(n24392), .B(n24757), .Z(n24598) );
  XNOR U24885 ( .A(n24391), .B(n24389), .Z(n24757) );
  AND U24886 ( .A(n24758), .B(n24759), .Z(n24389) );
  NANDN U24887 ( .A(n24760), .B(n24761), .Z(n24759) );
  OR U24888 ( .A(n24762), .B(n24763), .Z(n24761) );
  NAND U24889 ( .A(n24763), .B(n24762), .Z(n24758) );
  ANDN U24890 ( .B(B[191]), .A(n55), .Z(n24391) );
  XNOR U24891 ( .A(n24399), .B(n24764), .Z(n24392) );
  XNOR U24892 ( .A(n24398), .B(n24396), .Z(n24764) );
  AND U24893 ( .A(n24765), .B(n24766), .Z(n24396) );
  NANDN U24894 ( .A(n24767), .B(n24768), .Z(n24766) );
  NANDN U24895 ( .A(n24769), .B(n24770), .Z(n24768) );
  NANDN U24896 ( .A(n24770), .B(n24769), .Z(n24765) );
  ANDN U24897 ( .B(B[192]), .A(n56), .Z(n24398) );
  XNOR U24898 ( .A(n24406), .B(n24771), .Z(n24399) );
  XNOR U24899 ( .A(n24405), .B(n24403), .Z(n24771) );
  AND U24900 ( .A(n24772), .B(n24773), .Z(n24403) );
  NANDN U24901 ( .A(n24774), .B(n24775), .Z(n24773) );
  OR U24902 ( .A(n24776), .B(n24777), .Z(n24775) );
  NAND U24903 ( .A(n24777), .B(n24776), .Z(n24772) );
  ANDN U24904 ( .B(B[193]), .A(n57), .Z(n24405) );
  XNOR U24905 ( .A(n24413), .B(n24778), .Z(n24406) );
  XNOR U24906 ( .A(n24412), .B(n24410), .Z(n24778) );
  AND U24907 ( .A(n24779), .B(n24780), .Z(n24410) );
  NANDN U24908 ( .A(n24781), .B(n24782), .Z(n24780) );
  NANDN U24909 ( .A(n24783), .B(n24784), .Z(n24782) );
  NANDN U24910 ( .A(n24784), .B(n24783), .Z(n24779) );
  ANDN U24911 ( .B(B[194]), .A(n58), .Z(n24412) );
  XNOR U24912 ( .A(n24420), .B(n24785), .Z(n24413) );
  XNOR U24913 ( .A(n24419), .B(n24417), .Z(n24785) );
  AND U24914 ( .A(n24786), .B(n24787), .Z(n24417) );
  NANDN U24915 ( .A(n24788), .B(n24789), .Z(n24787) );
  OR U24916 ( .A(n24790), .B(n24791), .Z(n24789) );
  NAND U24917 ( .A(n24791), .B(n24790), .Z(n24786) );
  ANDN U24918 ( .B(B[195]), .A(n59), .Z(n24419) );
  XNOR U24919 ( .A(n24427), .B(n24792), .Z(n24420) );
  XNOR U24920 ( .A(n24426), .B(n24424), .Z(n24792) );
  AND U24921 ( .A(n24793), .B(n24794), .Z(n24424) );
  NANDN U24922 ( .A(n24795), .B(n24796), .Z(n24794) );
  NANDN U24923 ( .A(n24797), .B(n24798), .Z(n24796) );
  NANDN U24924 ( .A(n24798), .B(n24797), .Z(n24793) );
  ANDN U24925 ( .B(B[196]), .A(n60), .Z(n24426) );
  XNOR U24926 ( .A(n24434), .B(n24799), .Z(n24427) );
  XNOR U24927 ( .A(n24433), .B(n24431), .Z(n24799) );
  AND U24928 ( .A(n24800), .B(n24801), .Z(n24431) );
  NANDN U24929 ( .A(n24802), .B(n24803), .Z(n24801) );
  OR U24930 ( .A(n24804), .B(n24805), .Z(n24803) );
  NAND U24931 ( .A(n24805), .B(n24804), .Z(n24800) );
  ANDN U24932 ( .B(B[197]), .A(n61), .Z(n24433) );
  XNOR U24933 ( .A(n24441), .B(n24806), .Z(n24434) );
  XNOR U24934 ( .A(n24440), .B(n24438), .Z(n24806) );
  AND U24935 ( .A(n24807), .B(n24808), .Z(n24438) );
  NANDN U24936 ( .A(n24809), .B(n24810), .Z(n24808) );
  NANDN U24937 ( .A(n24811), .B(n24812), .Z(n24810) );
  NANDN U24938 ( .A(n24812), .B(n24811), .Z(n24807) );
  ANDN U24939 ( .B(B[198]), .A(n62), .Z(n24440) );
  XNOR U24940 ( .A(n24448), .B(n24813), .Z(n24441) );
  XNOR U24941 ( .A(n24447), .B(n24445), .Z(n24813) );
  AND U24942 ( .A(n24814), .B(n24815), .Z(n24445) );
  NANDN U24943 ( .A(n24816), .B(n24817), .Z(n24815) );
  OR U24944 ( .A(n24818), .B(n24819), .Z(n24817) );
  NAND U24945 ( .A(n24819), .B(n24818), .Z(n24814) );
  ANDN U24946 ( .B(B[199]), .A(n63), .Z(n24447) );
  XNOR U24947 ( .A(n24455), .B(n24820), .Z(n24448) );
  XNOR U24948 ( .A(n24454), .B(n24452), .Z(n24820) );
  AND U24949 ( .A(n24821), .B(n24822), .Z(n24452) );
  NANDN U24950 ( .A(n24823), .B(n24824), .Z(n24822) );
  NANDN U24951 ( .A(n24825), .B(n24826), .Z(n24824) );
  NANDN U24952 ( .A(n24826), .B(n24825), .Z(n24821) );
  ANDN U24953 ( .B(B[200]), .A(n64), .Z(n24454) );
  XNOR U24954 ( .A(n24462), .B(n24827), .Z(n24455) );
  XNOR U24955 ( .A(n24461), .B(n24459), .Z(n24827) );
  AND U24956 ( .A(n24828), .B(n24829), .Z(n24459) );
  NANDN U24957 ( .A(n24830), .B(n24831), .Z(n24829) );
  OR U24958 ( .A(n24832), .B(n24833), .Z(n24831) );
  NAND U24959 ( .A(n24833), .B(n24832), .Z(n24828) );
  ANDN U24960 ( .B(B[201]), .A(n65), .Z(n24461) );
  XNOR U24961 ( .A(n24469), .B(n24834), .Z(n24462) );
  XNOR U24962 ( .A(n24468), .B(n24466), .Z(n24834) );
  AND U24963 ( .A(n24835), .B(n24836), .Z(n24466) );
  NANDN U24964 ( .A(n24837), .B(n24838), .Z(n24836) );
  NANDN U24965 ( .A(n24839), .B(n24840), .Z(n24838) );
  NANDN U24966 ( .A(n24840), .B(n24839), .Z(n24835) );
  ANDN U24967 ( .B(B[202]), .A(n66), .Z(n24468) );
  XNOR U24968 ( .A(n24476), .B(n24841), .Z(n24469) );
  XNOR U24969 ( .A(n24475), .B(n24473), .Z(n24841) );
  AND U24970 ( .A(n24842), .B(n24843), .Z(n24473) );
  NANDN U24971 ( .A(n24844), .B(n24845), .Z(n24843) );
  OR U24972 ( .A(n24846), .B(n24847), .Z(n24845) );
  NAND U24973 ( .A(n24847), .B(n24846), .Z(n24842) );
  ANDN U24974 ( .B(B[203]), .A(n67), .Z(n24475) );
  XNOR U24975 ( .A(n24483), .B(n24848), .Z(n24476) );
  XNOR U24976 ( .A(n24482), .B(n24480), .Z(n24848) );
  AND U24977 ( .A(n24849), .B(n24850), .Z(n24480) );
  NANDN U24978 ( .A(n24851), .B(n24852), .Z(n24850) );
  NANDN U24979 ( .A(n24853), .B(n24854), .Z(n24852) );
  NANDN U24980 ( .A(n24854), .B(n24853), .Z(n24849) );
  ANDN U24981 ( .B(B[204]), .A(n68), .Z(n24482) );
  XNOR U24982 ( .A(n24490), .B(n24855), .Z(n24483) );
  XNOR U24983 ( .A(n24489), .B(n24487), .Z(n24855) );
  AND U24984 ( .A(n24856), .B(n24857), .Z(n24487) );
  NANDN U24985 ( .A(n24858), .B(n24859), .Z(n24857) );
  OR U24986 ( .A(n24860), .B(n24861), .Z(n24859) );
  NAND U24987 ( .A(n24861), .B(n24860), .Z(n24856) );
  ANDN U24988 ( .B(B[205]), .A(n69), .Z(n24489) );
  XNOR U24989 ( .A(n24497), .B(n24862), .Z(n24490) );
  XNOR U24990 ( .A(n24496), .B(n24494), .Z(n24862) );
  AND U24991 ( .A(n24863), .B(n24864), .Z(n24494) );
  NANDN U24992 ( .A(n24865), .B(n24866), .Z(n24864) );
  NANDN U24993 ( .A(n24867), .B(n24868), .Z(n24866) );
  NANDN U24994 ( .A(n24868), .B(n24867), .Z(n24863) );
  ANDN U24995 ( .B(B[206]), .A(n70), .Z(n24496) );
  XNOR U24996 ( .A(n24504), .B(n24869), .Z(n24497) );
  XNOR U24997 ( .A(n24503), .B(n24501), .Z(n24869) );
  AND U24998 ( .A(n24870), .B(n24871), .Z(n24501) );
  NANDN U24999 ( .A(n24872), .B(n24873), .Z(n24871) );
  OR U25000 ( .A(n24874), .B(n24875), .Z(n24873) );
  NAND U25001 ( .A(n24875), .B(n24874), .Z(n24870) );
  ANDN U25002 ( .B(B[207]), .A(n71), .Z(n24503) );
  XNOR U25003 ( .A(n24511), .B(n24876), .Z(n24504) );
  XNOR U25004 ( .A(n24510), .B(n24508), .Z(n24876) );
  AND U25005 ( .A(n24877), .B(n24878), .Z(n24508) );
  NANDN U25006 ( .A(n24879), .B(n24880), .Z(n24878) );
  NANDN U25007 ( .A(n24881), .B(n24882), .Z(n24880) );
  NANDN U25008 ( .A(n24882), .B(n24881), .Z(n24877) );
  ANDN U25009 ( .B(B[208]), .A(n72), .Z(n24510) );
  XNOR U25010 ( .A(n24518), .B(n24883), .Z(n24511) );
  XNOR U25011 ( .A(n24517), .B(n24515), .Z(n24883) );
  AND U25012 ( .A(n24884), .B(n24885), .Z(n24515) );
  NANDN U25013 ( .A(n24886), .B(n24887), .Z(n24885) );
  OR U25014 ( .A(n24888), .B(n24889), .Z(n24887) );
  NAND U25015 ( .A(n24889), .B(n24888), .Z(n24884) );
  ANDN U25016 ( .B(B[209]), .A(n73), .Z(n24517) );
  XNOR U25017 ( .A(n24525), .B(n24890), .Z(n24518) );
  XNOR U25018 ( .A(n24524), .B(n24522), .Z(n24890) );
  AND U25019 ( .A(n24891), .B(n24892), .Z(n24522) );
  NANDN U25020 ( .A(n24893), .B(n24894), .Z(n24892) );
  NANDN U25021 ( .A(n24895), .B(n24896), .Z(n24894) );
  NANDN U25022 ( .A(n24896), .B(n24895), .Z(n24891) );
  ANDN U25023 ( .B(B[210]), .A(n74), .Z(n24524) );
  XNOR U25024 ( .A(n24532), .B(n24897), .Z(n24525) );
  XNOR U25025 ( .A(n24531), .B(n24529), .Z(n24897) );
  AND U25026 ( .A(n24898), .B(n24899), .Z(n24529) );
  NANDN U25027 ( .A(n24900), .B(n24901), .Z(n24899) );
  OR U25028 ( .A(n24902), .B(n24903), .Z(n24901) );
  NAND U25029 ( .A(n24903), .B(n24902), .Z(n24898) );
  ANDN U25030 ( .B(B[211]), .A(n75), .Z(n24531) );
  XNOR U25031 ( .A(n24539), .B(n24904), .Z(n24532) );
  XNOR U25032 ( .A(n24538), .B(n24536), .Z(n24904) );
  AND U25033 ( .A(n24905), .B(n24906), .Z(n24536) );
  NANDN U25034 ( .A(n24907), .B(n24908), .Z(n24906) );
  NANDN U25035 ( .A(n24909), .B(n24910), .Z(n24908) );
  NANDN U25036 ( .A(n24910), .B(n24909), .Z(n24905) );
  ANDN U25037 ( .B(B[212]), .A(n76), .Z(n24538) );
  XNOR U25038 ( .A(n24546), .B(n24911), .Z(n24539) );
  XNOR U25039 ( .A(n24545), .B(n24543), .Z(n24911) );
  AND U25040 ( .A(n24912), .B(n24913), .Z(n24543) );
  NANDN U25041 ( .A(n24914), .B(n24915), .Z(n24913) );
  OR U25042 ( .A(n24916), .B(n24917), .Z(n24915) );
  NAND U25043 ( .A(n24917), .B(n24916), .Z(n24912) );
  ANDN U25044 ( .B(B[213]), .A(n77), .Z(n24545) );
  XNOR U25045 ( .A(n24553), .B(n24918), .Z(n24546) );
  XNOR U25046 ( .A(n24552), .B(n24550), .Z(n24918) );
  AND U25047 ( .A(n24919), .B(n24920), .Z(n24550) );
  NANDN U25048 ( .A(n24921), .B(n24922), .Z(n24920) );
  NANDN U25049 ( .A(n24923), .B(n24924), .Z(n24922) );
  NANDN U25050 ( .A(n24924), .B(n24923), .Z(n24919) );
  ANDN U25051 ( .B(B[214]), .A(n78), .Z(n24552) );
  XNOR U25052 ( .A(n24560), .B(n24925), .Z(n24553) );
  XNOR U25053 ( .A(n24559), .B(n24557), .Z(n24925) );
  AND U25054 ( .A(n24926), .B(n24927), .Z(n24557) );
  NANDN U25055 ( .A(n24928), .B(n24929), .Z(n24927) );
  OR U25056 ( .A(n24930), .B(n24931), .Z(n24929) );
  NAND U25057 ( .A(n24931), .B(n24930), .Z(n24926) );
  ANDN U25058 ( .B(B[215]), .A(n79), .Z(n24559) );
  XNOR U25059 ( .A(n24567), .B(n24932), .Z(n24560) );
  XNOR U25060 ( .A(n24566), .B(n24564), .Z(n24932) );
  AND U25061 ( .A(n24933), .B(n24934), .Z(n24564) );
  NANDN U25062 ( .A(n24935), .B(n24936), .Z(n24934) );
  NANDN U25063 ( .A(n24937), .B(n24938), .Z(n24936) );
  NANDN U25064 ( .A(n24938), .B(n24937), .Z(n24933) );
  ANDN U25065 ( .B(B[216]), .A(n80), .Z(n24566) );
  XNOR U25066 ( .A(n24574), .B(n24939), .Z(n24567) );
  XNOR U25067 ( .A(n24573), .B(n24571), .Z(n24939) );
  AND U25068 ( .A(n24940), .B(n24941), .Z(n24571) );
  NANDN U25069 ( .A(n24942), .B(n24943), .Z(n24941) );
  OR U25070 ( .A(n24944), .B(n24945), .Z(n24943) );
  NAND U25071 ( .A(n24945), .B(n24944), .Z(n24940) );
  ANDN U25072 ( .B(B[217]), .A(n81), .Z(n24573) );
  XNOR U25073 ( .A(n24581), .B(n24946), .Z(n24574) );
  XNOR U25074 ( .A(n24580), .B(n24578), .Z(n24946) );
  AND U25075 ( .A(n24947), .B(n24948), .Z(n24578) );
  NANDN U25076 ( .A(n24949), .B(n24950), .Z(n24948) );
  NAND U25077 ( .A(n24951), .B(n24952), .Z(n24950) );
  ANDN U25078 ( .B(B[218]), .A(n82), .Z(n24580) );
  XOR U25079 ( .A(n24587), .B(n24953), .Z(n24581) );
  XNOR U25080 ( .A(n24585), .B(n24588), .Z(n24953) );
  NAND U25081 ( .A(A[2]), .B(B[219]), .Z(n24588) );
  NANDN U25082 ( .A(n24954), .B(n24955), .Z(n24585) );
  AND U25083 ( .A(A[0]), .B(B[220]), .Z(n24955) );
  XNOR U25084 ( .A(n24590), .B(n24956), .Z(n24587) );
  NAND U25085 ( .A(A[0]), .B(B[221]), .Z(n24956) );
  NAND U25086 ( .A(B[220]), .B(A[1]), .Z(n24590) );
  NAND U25087 ( .A(n24957), .B(n24958), .Z(n354) );
  NANDN U25088 ( .A(n24959), .B(n24960), .Z(n24958) );
  OR U25089 ( .A(n24961), .B(n24962), .Z(n24960) );
  NAND U25090 ( .A(n24962), .B(n24961), .Z(n24957) );
  XOR U25091 ( .A(n356), .B(n355), .Z(\A1[218] ) );
  XOR U25092 ( .A(n24962), .B(n24963), .Z(n355) );
  XNOR U25093 ( .A(n24961), .B(n24959), .Z(n24963) );
  AND U25094 ( .A(n24964), .B(n24965), .Z(n24959) );
  NANDN U25095 ( .A(n24966), .B(n24967), .Z(n24965) );
  NANDN U25096 ( .A(n24968), .B(n24969), .Z(n24967) );
  NANDN U25097 ( .A(n24969), .B(n24968), .Z(n24964) );
  ANDN U25098 ( .B(B[189]), .A(n54), .Z(n24961) );
  XNOR U25099 ( .A(n24756), .B(n24970), .Z(n24962) );
  XNOR U25100 ( .A(n24755), .B(n24753), .Z(n24970) );
  AND U25101 ( .A(n24971), .B(n24972), .Z(n24753) );
  NANDN U25102 ( .A(n24973), .B(n24974), .Z(n24972) );
  OR U25103 ( .A(n24975), .B(n24976), .Z(n24974) );
  NAND U25104 ( .A(n24976), .B(n24975), .Z(n24971) );
  ANDN U25105 ( .B(B[190]), .A(n55), .Z(n24755) );
  XNOR U25106 ( .A(n24763), .B(n24977), .Z(n24756) );
  XNOR U25107 ( .A(n24762), .B(n24760), .Z(n24977) );
  AND U25108 ( .A(n24978), .B(n24979), .Z(n24760) );
  NANDN U25109 ( .A(n24980), .B(n24981), .Z(n24979) );
  NANDN U25110 ( .A(n24982), .B(n24983), .Z(n24981) );
  NANDN U25111 ( .A(n24983), .B(n24982), .Z(n24978) );
  ANDN U25112 ( .B(B[191]), .A(n56), .Z(n24762) );
  XNOR U25113 ( .A(n24770), .B(n24984), .Z(n24763) );
  XNOR U25114 ( .A(n24769), .B(n24767), .Z(n24984) );
  AND U25115 ( .A(n24985), .B(n24986), .Z(n24767) );
  NANDN U25116 ( .A(n24987), .B(n24988), .Z(n24986) );
  OR U25117 ( .A(n24989), .B(n24990), .Z(n24988) );
  NAND U25118 ( .A(n24990), .B(n24989), .Z(n24985) );
  ANDN U25119 ( .B(B[192]), .A(n57), .Z(n24769) );
  XNOR U25120 ( .A(n24777), .B(n24991), .Z(n24770) );
  XNOR U25121 ( .A(n24776), .B(n24774), .Z(n24991) );
  AND U25122 ( .A(n24992), .B(n24993), .Z(n24774) );
  NANDN U25123 ( .A(n24994), .B(n24995), .Z(n24993) );
  NANDN U25124 ( .A(n24996), .B(n24997), .Z(n24995) );
  NANDN U25125 ( .A(n24997), .B(n24996), .Z(n24992) );
  ANDN U25126 ( .B(B[193]), .A(n58), .Z(n24776) );
  XNOR U25127 ( .A(n24784), .B(n24998), .Z(n24777) );
  XNOR U25128 ( .A(n24783), .B(n24781), .Z(n24998) );
  AND U25129 ( .A(n24999), .B(n25000), .Z(n24781) );
  NANDN U25130 ( .A(n25001), .B(n25002), .Z(n25000) );
  OR U25131 ( .A(n25003), .B(n25004), .Z(n25002) );
  NAND U25132 ( .A(n25004), .B(n25003), .Z(n24999) );
  ANDN U25133 ( .B(B[194]), .A(n59), .Z(n24783) );
  XNOR U25134 ( .A(n24791), .B(n25005), .Z(n24784) );
  XNOR U25135 ( .A(n24790), .B(n24788), .Z(n25005) );
  AND U25136 ( .A(n25006), .B(n25007), .Z(n24788) );
  NANDN U25137 ( .A(n25008), .B(n25009), .Z(n25007) );
  NANDN U25138 ( .A(n25010), .B(n25011), .Z(n25009) );
  NANDN U25139 ( .A(n25011), .B(n25010), .Z(n25006) );
  ANDN U25140 ( .B(B[195]), .A(n60), .Z(n24790) );
  XNOR U25141 ( .A(n24798), .B(n25012), .Z(n24791) );
  XNOR U25142 ( .A(n24797), .B(n24795), .Z(n25012) );
  AND U25143 ( .A(n25013), .B(n25014), .Z(n24795) );
  NANDN U25144 ( .A(n25015), .B(n25016), .Z(n25014) );
  OR U25145 ( .A(n25017), .B(n25018), .Z(n25016) );
  NAND U25146 ( .A(n25018), .B(n25017), .Z(n25013) );
  ANDN U25147 ( .B(B[196]), .A(n61), .Z(n24797) );
  XNOR U25148 ( .A(n24805), .B(n25019), .Z(n24798) );
  XNOR U25149 ( .A(n24804), .B(n24802), .Z(n25019) );
  AND U25150 ( .A(n25020), .B(n25021), .Z(n24802) );
  NANDN U25151 ( .A(n25022), .B(n25023), .Z(n25021) );
  NANDN U25152 ( .A(n25024), .B(n25025), .Z(n25023) );
  NANDN U25153 ( .A(n25025), .B(n25024), .Z(n25020) );
  ANDN U25154 ( .B(B[197]), .A(n62), .Z(n24804) );
  XNOR U25155 ( .A(n24812), .B(n25026), .Z(n24805) );
  XNOR U25156 ( .A(n24811), .B(n24809), .Z(n25026) );
  AND U25157 ( .A(n25027), .B(n25028), .Z(n24809) );
  NANDN U25158 ( .A(n25029), .B(n25030), .Z(n25028) );
  OR U25159 ( .A(n25031), .B(n25032), .Z(n25030) );
  NAND U25160 ( .A(n25032), .B(n25031), .Z(n25027) );
  ANDN U25161 ( .B(B[198]), .A(n63), .Z(n24811) );
  XNOR U25162 ( .A(n24819), .B(n25033), .Z(n24812) );
  XNOR U25163 ( .A(n24818), .B(n24816), .Z(n25033) );
  AND U25164 ( .A(n25034), .B(n25035), .Z(n24816) );
  NANDN U25165 ( .A(n25036), .B(n25037), .Z(n25035) );
  NANDN U25166 ( .A(n25038), .B(n25039), .Z(n25037) );
  NANDN U25167 ( .A(n25039), .B(n25038), .Z(n25034) );
  ANDN U25168 ( .B(B[199]), .A(n64), .Z(n24818) );
  XNOR U25169 ( .A(n24826), .B(n25040), .Z(n24819) );
  XNOR U25170 ( .A(n24825), .B(n24823), .Z(n25040) );
  AND U25171 ( .A(n25041), .B(n25042), .Z(n24823) );
  NANDN U25172 ( .A(n25043), .B(n25044), .Z(n25042) );
  OR U25173 ( .A(n25045), .B(n25046), .Z(n25044) );
  NAND U25174 ( .A(n25046), .B(n25045), .Z(n25041) );
  ANDN U25175 ( .B(B[200]), .A(n65), .Z(n24825) );
  XNOR U25176 ( .A(n24833), .B(n25047), .Z(n24826) );
  XNOR U25177 ( .A(n24832), .B(n24830), .Z(n25047) );
  AND U25178 ( .A(n25048), .B(n25049), .Z(n24830) );
  NANDN U25179 ( .A(n25050), .B(n25051), .Z(n25049) );
  NANDN U25180 ( .A(n25052), .B(n25053), .Z(n25051) );
  NANDN U25181 ( .A(n25053), .B(n25052), .Z(n25048) );
  ANDN U25182 ( .B(B[201]), .A(n66), .Z(n24832) );
  XNOR U25183 ( .A(n24840), .B(n25054), .Z(n24833) );
  XNOR U25184 ( .A(n24839), .B(n24837), .Z(n25054) );
  AND U25185 ( .A(n25055), .B(n25056), .Z(n24837) );
  NANDN U25186 ( .A(n25057), .B(n25058), .Z(n25056) );
  OR U25187 ( .A(n25059), .B(n25060), .Z(n25058) );
  NAND U25188 ( .A(n25060), .B(n25059), .Z(n25055) );
  ANDN U25189 ( .B(B[202]), .A(n67), .Z(n24839) );
  XNOR U25190 ( .A(n24847), .B(n25061), .Z(n24840) );
  XNOR U25191 ( .A(n24846), .B(n24844), .Z(n25061) );
  AND U25192 ( .A(n25062), .B(n25063), .Z(n24844) );
  NANDN U25193 ( .A(n25064), .B(n25065), .Z(n25063) );
  NANDN U25194 ( .A(n25066), .B(n25067), .Z(n25065) );
  NANDN U25195 ( .A(n25067), .B(n25066), .Z(n25062) );
  ANDN U25196 ( .B(B[203]), .A(n68), .Z(n24846) );
  XNOR U25197 ( .A(n24854), .B(n25068), .Z(n24847) );
  XNOR U25198 ( .A(n24853), .B(n24851), .Z(n25068) );
  AND U25199 ( .A(n25069), .B(n25070), .Z(n24851) );
  NANDN U25200 ( .A(n25071), .B(n25072), .Z(n25070) );
  OR U25201 ( .A(n25073), .B(n25074), .Z(n25072) );
  NAND U25202 ( .A(n25074), .B(n25073), .Z(n25069) );
  ANDN U25203 ( .B(B[204]), .A(n69), .Z(n24853) );
  XNOR U25204 ( .A(n24861), .B(n25075), .Z(n24854) );
  XNOR U25205 ( .A(n24860), .B(n24858), .Z(n25075) );
  AND U25206 ( .A(n25076), .B(n25077), .Z(n24858) );
  NANDN U25207 ( .A(n25078), .B(n25079), .Z(n25077) );
  NANDN U25208 ( .A(n25080), .B(n25081), .Z(n25079) );
  NANDN U25209 ( .A(n25081), .B(n25080), .Z(n25076) );
  ANDN U25210 ( .B(B[205]), .A(n70), .Z(n24860) );
  XNOR U25211 ( .A(n24868), .B(n25082), .Z(n24861) );
  XNOR U25212 ( .A(n24867), .B(n24865), .Z(n25082) );
  AND U25213 ( .A(n25083), .B(n25084), .Z(n24865) );
  NANDN U25214 ( .A(n25085), .B(n25086), .Z(n25084) );
  OR U25215 ( .A(n25087), .B(n25088), .Z(n25086) );
  NAND U25216 ( .A(n25088), .B(n25087), .Z(n25083) );
  ANDN U25217 ( .B(B[206]), .A(n71), .Z(n24867) );
  XNOR U25218 ( .A(n24875), .B(n25089), .Z(n24868) );
  XNOR U25219 ( .A(n24874), .B(n24872), .Z(n25089) );
  AND U25220 ( .A(n25090), .B(n25091), .Z(n24872) );
  NANDN U25221 ( .A(n25092), .B(n25093), .Z(n25091) );
  NANDN U25222 ( .A(n25094), .B(n25095), .Z(n25093) );
  NANDN U25223 ( .A(n25095), .B(n25094), .Z(n25090) );
  ANDN U25224 ( .B(B[207]), .A(n72), .Z(n24874) );
  XNOR U25225 ( .A(n24882), .B(n25096), .Z(n24875) );
  XNOR U25226 ( .A(n24881), .B(n24879), .Z(n25096) );
  AND U25227 ( .A(n25097), .B(n25098), .Z(n24879) );
  NANDN U25228 ( .A(n25099), .B(n25100), .Z(n25098) );
  OR U25229 ( .A(n25101), .B(n25102), .Z(n25100) );
  NAND U25230 ( .A(n25102), .B(n25101), .Z(n25097) );
  ANDN U25231 ( .B(B[208]), .A(n73), .Z(n24881) );
  XNOR U25232 ( .A(n24889), .B(n25103), .Z(n24882) );
  XNOR U25233 ( .A(n24888), .B(n24886), .Z(n25103) );
  AND U25234 ( .A(n25104), .B(n25105), .Z(n24886) );
  NANDN U25235 ( .A(n25106), .B(n25107), .Z(n25105) );
  NANDN U25236 ( .A(n25108), .B(n25109), .Z(n25107) );
  NANDN U25237 ( .A(n25109), .B(n25108), .Z(n25104) );
  ANDN U25238 ( .B(B[209]), .A(n74), .Z(n24888) );
  XNOR U25239 ( .A(n24896), .B(n25110), .Z(n24889) );
  XNOR U25240 ( .A(n24895), .B(n24893), .Z(n25110) );
  AND U25241 ( .A(n25111), .B(n25112), .Z(n24893) );
  NANDN U25242 ( .A(n25113), .B(n25114), .Z(n25112) );
  OR U25243 ( .A(n25115), .B(n25116), .Z(n25114) );
  NAND U25244 ( .A(n25116), .B(n25115), .Z(n25111) );
  ANDN U25245 ( .B(B[210]), .A(n75), .Z(n24895) );
  XNOR U25246 ( .A(n24903), .B(n25117), .Z(n24896) );
  XNOR U25247 ( .A(n24902), .B(n24900), .Z(n25117) );
  AND U25248 ( .A(n25118), .B(n25119), .Z(n24900) );
  NANDN U25249 ( .A(n25120), .B(n25121), .Z(n25119) );
  NANDN U25250 ( .A(n25122), .B(n25123), .Z(n25121) );
  NANDN U25251 ( .A(n25123), .B(n25122), .Z(n25118) );
  ANDN U25252 ( .B(B[211]), .A(n76), .Z(n24902) );
  XNOR U25253 ( .A(n24910), .B(n25124), .Z(n24903) );
  XNOR U25254 ( .A(n24909), .B(n24907), .Z(n25124) );
  AND U25255 ( .A(n25125), .B(n25126), .Z(n24907) );
  NANDN U25256 ( .A(n25127), .B(n25128), .Z(n25126) );
  OR U25257 ( .A(n25129), .B(n25130), .Z(n25128) );
  NAND U25258 ( .A(n25130), .B(n25129), .Z(n25125) );
  ANDN U25259 ( .B(B[212]), .A(n77), .Z(n24909) );
  XNOR U25260 ( .A(n24917), .B(n25131), .Z(n24910) );
  XNOR U25261 ( .A(n24916), .B(n24914), .Z(n25131) );
  AND U25262 ( .A(n25132), .B(n25133), .Z(n24914) );
  NANDN U25263 ( .A(n25134), .B(n25135), .Z(n25133) );
  NANDN U25264 ( .A(n25136), .B(n25137), .Z(n25135) );
  NANDN U25265 ( .A(n25137), .B(n25136), .Z(n25132) );
  ANDN U25266 ( .B(B[213]), .A(n78), .Z(n24916) );
  XNOR U25267 ( .A(n24924), .B(n25138), .Z(n24917) );
  XNOR U25268 ( .A(n24923), .B(n24921), .Z(n25138) );
  AND U25269 ( .A(n25139), .B(n25140), .Z(n24921) );
  NANDN U25270 ( .A(n25141), .B(n25142), .Z(n25140) );
  OR U25271 ( .A(n25143), .B(n25144), .Z(n25142) );
  NAND U25272 ( .A(n25144), .B(n25143), .Z(n25139) );
  ANDN U25273 ( .B(B[214]), .A(n79), .Z(n24923) );
  XNOR U25274 ( .A(n24931), .B(n25145), .Z(n24924) );
  XNOR U25275 ( .A(n24930), .B(n24928), .Z(n25145) );
  AND U25276 ( .A(n25146), .B(n25147), .Z(n24928) );
  NANDN U25277 ( .A(n25148), .B(n25149), .Z(n25147) );
  NANDN U25278 ( .A(n25150), .B(n25151), .Z(n25149) );
  NANDN U25279 ( .A(n25151), .B(n25150), .Z(n25146) );
  ANDN U25280 ( .B(B[215]), .A(n80), .Z(n24930) );
  XNOR U25281 ( .A(n24938), .B(n25152), .Z(n24931) );
  XNOR U25282 ( .A(n24937), .B(n24935), .Z(n25152) );
  AND U25283 ( .A(n25153), .B(n25154), .Z(n24935) );
  NANDN U25284 ( .A(n25155), .B(n25156), .Z(n25154) );
  OR U25285 ( .A(n25157), .B(n25158), .Z(n25156) );
  NAND U25286 ( .A(n25158), .B(n25157), .Z(n25153) );
  ANDN U25287 ( .B(B[216]), .A(n81), .Z(n24937) );
  XNOR U25288 ( .A(n24945), .B(n25159), .Z(n24938) );
  XNOR U25289 ( .A(n24944), .B(n24942), .Z(n25159) );
  AND U25290 ( .A(n25160), .B(n25161), .Z(n24942) );
  NANDN U25291 ( .A(n25162), .B(n25163), .Z(n25161) );
  NAND U25292 ( .A(n25164), .B(n25165), .Z(n25163) );
  ANDN U25293 ( .B(B[217]), .A(n82), .Z(n24944) );
  XOR U25294 ( .A(n24951), .B(n25166), .Z(n24945) );
  XNOR U25295 ( .A(n24949), .B(n24952), .Z(n25166) );
  NAND U25296 ( .A(A[2]), .B(B[218]), .Z(n24952) );
  NANDN U25297 ( .A(n25167), .B(n25168), .Z(n24949) );
  AND U25298 ( .A(A[0]), .B(B[219]), .Z(n25168) );
  XNOR U25299 ( .A(n24954), .B(n25169), .Z(n24951) );
  NAND U25300 ( .A(A[0]), .B(B[220]), .Z(n25169) );
  NAND U25301 ( .A(B[219]), .B(A[1]), .Z(n24954) );
  NAND U25302 ( .A(n25170), .B(n25171), .Z(n356) );
  NANDN U25303 ( .A(n25172), .B(n25173), .Z(n25171) );
  OR U25304 ( .A(n25174), .B(n25175), .Z(n25173) );
  NAND U25305 ( .A(n25175), .B(n25174), .Z(n25170) );
  XOR U25306 ( .A(n358), .B(n357), .Z(\A1[217] ) );
  XOR U25307 ( .A(n25175), .B(n25176), .Z(n357) );
  XNOR U25308 ( .A(n25174), .B(n25172), .Z(n25176) );
  AND U25309 ( .A(n25177), .B(n25178), .Z(n25172) );
  NANDN U25310 ( .A(n25179), .B(n25180), .Z(n25178) );
  NANDN U25311 ( .A(n25181), .B(n25182), .Z(n25180) );
  NANDN U25312 ( .A(n25182), .B(n25181), .Z(n25177) );
  ANDN U25313 ( .B(B[188]), .A(n54), .Z(n25174) );
  XNOR U25314 ( .A(n24969), .B(n25183), .Z(n25175) );
  XNOR U25315 ( .A(n24968), .B(n24966), .Z(n25183) );
  AND U25316 ( .A(n25184), .B(n25185), .Z(n24966) );
  NANDN U25317 ( .A(n25186), .B(n25187), .Z(n25185) );
  OR U25318 ( .A(n25188), .B(n25189), .Z(n25187) );
  NAND U25319 ( .A(n25189), .B(n25188), .Z(n25184) );
  ANDN U25320 ( .B(B[189]), .A(n55), .Z(n24968) );
  XNOR U25321 ( .A(n24976), .B(n25190), .Z(n24969) );
  XNOR U25322 ( .A(n24975), .B(n24973), .Z(n25190) );
  AND U25323 ( .A(n25191), .B(n25192), .Z(n24973) );
  NANDN U25324 ( .A(n25193), .B(n25194), .Z(n25192) );
  NANDN U25325 ( .A(n25195), .B(n25196), .Z(n25194) );
  NANDN U25326 ( .A(n25196), .B(n25195), .Z(n25191) );
  ANDN U25327 ( .B(B[190]), .A(n56), .Z(n24975) );
  XNOR U25328 ( .A(n24983), .B(n25197), .Z(n24976) );
  XNOR U25329 ( .A(n24982), .B(n24980), .Z(n25197) );
  AND U25330 ( .A(n25198), .B(n25199), .Z(n24980) );
  NANDN U25331 ( .A(n25200), .B(n25201), .Z(n25199) );
  OR U25332 ( .A(n25202), .B(n25203), .Z(n25201) );
  NAND U25333 ( .A(n25203), .B(n25202), .Z(n25198) );
  ANDN U25334 ( .B(B[191]), .A(n57), .Z(n24982) );
  XNOR U25335 ( .A(n24990), .B(n25204), .Z(n24983) );
  XNOR U25336 ( .A(n24989), .B(n24987), .Z(n25204) );
  AND U25337 ( .A(n25205), .B(n25206), .Z(n24987) );
  NANDN U25338 ( .A(n25207), .B(n25208), .Z(n25206) );
  NANDN U25339 ( .A(n25209), .B(n25210), .Z(n25208) );
  NANDN U25340 ( .A(n25210), .B(n25209), .Z(n25205) );
  ANDN U25341 ( .B(B[192]), .A(n58), .Z(n24989) );
  XNOR U25342 ( .A(n24997), .B(n25211), .Z(n24990) );
  XNOR U25343 ( .A(n24996), .B(n24994), .Z(n25211) );
  AND U25344 ( .A(n25212), .B(n25213), .Z(n24994) );
  NANDN U25345 ( .A(n25214), .B(n25215), .Z(n25213) );
  OR U25346 ( .A(n25216), .B(n25217), .Z(n25215) );
  NAND U25347 ( .A(n25217), .B(n25216), .Z(n25212) );
  ANDN U25348 ( .B(B[193]), .A(n59), .Z(n24996) );
  XNOR U25349 ( .A(n25004), .B(n25218), .Z(n24997) );
  XNOR U25350 ( .A(n25003), .B(n25001), .Z(n25218) );
  AND U25351 ( .A(n25219), .B(n25220), .Z(n25001) );
  NANDN U25352 ( .A(n25221), .B(n25222), .Z(n25220) );
  NANDN U25353 ( .A(n25223), .B(n25224), .Z(n25222) );
  NANDN U25354 ( .A(n25224), .B(n25223), .Z(n25219) );
  ANDN U25355 ( .B(B[194]), .A(n60), .Z(n25003) );
  XNOR U25356 ( .A(n25011), .B(n25225), .Z(n25004) );
  XNOR U25357 ( .A(n25010), .B(n25008), .Z(n25225) );
  AND U25358 ( .A(n25226), .B(n25227), .Z(n25008) );
  NANDN U25359 ( .A(n25228), .B(n25229), .Z(n25227) );
  OR U25360 ( .A(n25230), .B(n25231), .Z(n25229) );
  NAND U25361 ( .A(n25231), .B(n25230), .Z(n25226) );
  ANDN U25362 ( .B(B[195]), .A(n61), .Z(n25010) );
  XNOR U25363 ( .A(n25018), .B(n25232), .Z(n25011) );
  XNOR U25364 ( .A(n25017), .B(n25015), .Z(n25232) );
  AND U25365 ( .A(n25233), .B(n25234), .Z(n25015) );
  NANDN U25366 ( .A(n25235), .B(n25236), .Z(n25234) );
  NANDN U25367 ( .A(n25237), .B(n25238), .Z(n25236) );
  NANDN U25368 ( .A(n25238), .B(n25237), .Z(n25233) );
  ANDN U25369 ( .B(B[196]), .A(n62), .Z(n25017) );
  XNOR U25370 ( .A(n25025), .B(n25239), .Z(n25018) );
  XNOR U25371 ( .A(n25024), .B(n25022), .Z(n25239) );
  AND U25372 ( .A(n25240), .B(n25241), .Z(n25022) );
  NANDN U25373 ( .A(n25242), .B(n25243), .Z(n25241) );
  OR U25374 ( .A(n25244), .B(n25245), .Z(n25243) );
  NAND U25375 ( .A(n25245), .B(n25244), .Z(n25240) );
  ANDN U25376 ( .B(B[197]), .A(n63), .Z(n25024) );
  XNOR U25377 ( .A(n25032), .B(n25246), .Z(n25025) );
  XNOR U25378 ( .A(n25031), .B(n25029), .Z(n25246) );
  AND U25379 ( .A(n25247), .B(n25248), .Z(n25029) );
  NANDN U25380 ( .A(n25249), .B(n25250), .Z(n25248) );
  NANDN U25381 ( .A(n25251), .B(n25252), .Z(n25250) );
  NANDN U25382 ( .A(n25252), .B(n25251), .Z(n25247) );
  ANDN U25383 ( .B(B[198]), .A(n64), .Z(n25031) );
  XNOR U25384 ( .A(n25039), .B(n25253), .Z(n25032) );
  XNOR U25385 ( .A(n25038), .B(n25036), .Z(n25253) );
  AND U25386 ( .A(n25254), .B(n25255), .Z(n25036) );
  NANDN U25387 ( .A(n25256), .B(n25257), .Z(n25255) );
  OR U25388 ( .A(n25258), .B(n25259), .Z(n25257) );
  NAND U25389 ( .A(n25259), .B(n25258), .Z(n25254) );
  ANDN U25390 ( .B(B[199]), .A(n65), .Z(n25038) );
  XNOR U25391 ( .A(n25046), .B(n25260), .Z(n25039) );
  XNOR U25392 ( .A(n25045), .B(n25043), .Z(n25260) );
  AND U25393 ( .A(n25261), .B(n25262), .Z(n25043) );
  NANDN U25394 ( .A(n25263), .B(n25264), .Z(n25262) );
  NANDN U25395 ( .A(n25265), .B(n25266), .Z(n25264) );
  NANDN U25396 ( .A(n25266), .B(n25265), .Z(n25261) );
  ANDN U25397 ( .B(B[200]), .A(n66), .Z(n25045) );
  XNOR U25398 ( .A(n25053), .B(n25267), .Z(n25046) );
  XNOR U25399 ( .A(n25052), .B(n25050), .Z(n25267) );
  AND U25400 ( .A(n25268), .B(n25269), .Z(n25050) );
  NANDN U25401 ( .A(n25270), .B(n25271), .Z(n25269) );
  OR U25402 ( .A(n25272), .B(n25273), .Z(n25271) );
  NAND U25403 ( .A(n25273), .B(n25272), .Z(n25268) );
  ANDN U25404 ( .B(B[201]), .A(n67), .Z(n25052) );
  XNOR U25405 ( .A(n25060), .B(n25274), .Z(n25053) );
  XNOR U25406 ( .A(n25059), .B(n25057), .Z(n25274) );
  AND U25407 ( .A(n25275), .B(n25276), .Z(n25057) );
  NANDN U25408 ( .A(n25277), .B(n25278), .Z(n25276) );
  NANDN U25409 ( .A(n25279), .B(n25280), .Z(n25278) );
  NANDN U25410 ( .A(n25280), .B(n25279), .Z(n25275) );
  ANDN U25411 ( .B(B[202]), .A(n68), .Z(n25059) );
  XNOR U25412 ( .A(n25067), .B(n25281), .Z(n25060) );
  XNOR U25413 ( .A(n25066), .B(n25064), .Z(n25281) );
  AND U25414 ( .A(n25282), .B(n25283), .Z(n25064) );
  NANDN U25415 ( .A(n25284), .B(n25285), .Z(n25283) );
  OR U25416 ( .A(n25286), .B(n25287), .Z(n25285) );
  NAND U25417 ( .A(n25287), .B(n25286), .Z(n25282) );
  ANDN U25418 ( .B(B[203]), .A(n69), .Z(n25066) );
  XNOR U25419 ( .A(n25074), .B(n25288), .Z(n25067) );
  XNOR U25420 ( .A(n25073), .B(n25071), .Z(n25288) );
  AND U25421 ( .A(n25289), .B(n25290), .Z(n25071) );
  NANDN U25422 ( .A(n25291), .B(n25292), .Z(n25290) );
  NANDN U25423 ( .A(n25293), .B(n25294), .Z(n25292) );
  NANDN U25424 ( .A(n25294), .B(n25293), .Z(n25289) );
  ANDN U25425 ( .B(B[204]), .A(n70), .Z(n25073) );
  XNOR U25426 ( .A(n25081), .B(n25295), .Z(n25074) );
  XNOR U25427 ( .A(n25080), .B(n25078), .Z(n25295) );
  AND U25428 ( .A(n25296), .B(n25297), .Z(n25078) );
  NANDN U25429 ( .A(n25298), .B(n25299), .Z(n25297) );
  OR U25430 ( .A(n25300), .B(n25301), .Z(n25299) );
  NAND U25431 ( .A(n25301), .B(n25300), .Z(n25296) );
  ANDN U25432 ( .B(B[205]), .A(n71), .Z(n25080) );
  XNOR U25433 ( .A(n25088), .B(n25302), .Z(n25081) );
  XNOR U25434 ( .A(n25087), .B(n25085), .Z(n25302) );
  AND U25435 ( .A(n25303), .B(n25304), .Z(n25085) );
  NANDN U25436 ( .A(n25305), .B(n25306), .Z(n25304) );
  NANDN U25437 ( .A(n25307), .B(n25308), .Z(n25306) );
  NANDN U25438 ( .A(n25308), .B(n25307), .Z(n25303) );
  ANDN U25439 ( .B(B[206]), .A(n72), .Z(n25087) );
  XNOR U25440 ( .A(n25095), .B(n25309), .Z(n25088) );
  XNOR U25441 ( .A(n25094), .B(n25092), .Z(n25309) );
  AND U25442 ( .A(n25310), .B(n25311), .Z(n25092) );
  NANDN U25443 ( .A(n25312), .B(n25313), .Z(n25311) );
  OR U25444 ( .A(n25314), .B(n25315), .Z(n25313) );
  NAND U25445 ( .A(n25315), .B(n25314), .Z(n25310) );
  ANDN U25446 ( .B(B[207]), .A(n73), .Z(n25094) );
  XNOR U25447 ( .A(n25102), .B(n25316), .Z(n25095) );
  XNOR U25448 ( .A(n25101), .B(n25099), .Z(n25316) );
  AND U25449 ( .A(n25317), .B(n25318), .Z(n25099) );
  NANDN U25450 ( .A(n25319), .B(n25320), .Z(n25318) );
  NANDN U25451 ( .A(n25321), .B(n25322), .Z(n25320) );
  NANDN U25452 ( .A(n25322), .B(n25321), .Z(n25317) );
  ANDN U25453 ( .B(B[208]), .A(n74), .Z(n25101) );
  XNOR U25454 ( .A(n25109), .B(n25323), .Z(n25102) );
  XNOR U25455 ( .A(n25108), .B(n25106), .Z(n25323) );
  AND U25456 ( .A(n25324), .B(n25325), .Z(n25106) );
  NANDN U25457 ( .A(n25326), .B(n25327), .Z(n25325) );
  OR U25458 ( .A(n25328), .B(n25329), .Z(n25327) );
  NAND U25459 ( .A(n25329), .B(n25328), .Z(n25324) );
  ANDN U25460 ( .B(B[209]), .A(n75), .Z(n25108) );
  XNOR U25461 ( .A(n25116), .B(n25330), .Z(n25109) );
  XNOR U25462 ( .A(n25115), .B(n25113), .Z(n25330) );
  AND U25463 ( .A(n25331), .B(n25332), .Z(n25113) );
  NANDN U25464 ( .A(n25333), .B(n25334), .Z(n25332) );
  NANDN U25465 ( .A(n25335), .B(n25336), .Z(n25334) );
  NANDN U25466 ( .A(n25336), .B(n25335), .Z(n25331) );
  ANDN U25467 ( .B(B[210]), .A(n76), .Z(n25115) );
  XNOR U25468 ( .A(n25123), .B(n25337), .Z(n25116) );
  XNOR U25469 ( .A(n25122), .B(n25120), .Z(n25337) );
  AND U25470 ( .A(n25338), .B(n25339), .Z(n25120) );
  NANDN U25471 ( .A(n25340), .B(n25341), .Z(n25339) );
  OR U25472 ( .A(n25342), .B(n25343), .Z(n25341) );
  NAND U25473 ( .A(n25343), .B(n25342), .Z(n25338) );
  ANDN U25474 ( .B(B[211]), .A(n77), .Z(n25122) );
  XNOR U25475 ( .A(n25130), .B(n25344), .Z(n25123) );
  XNOR U25476 ( .A(n25129), .B(n25127), .Z(n25344) );
  AND U25477 ( .A(n25345), .B(n25346), .Z(n25127) );
  NANDN U25478 ( .A(n25347), .B(n25348), .Z(n25346) );
  NANDN U25479 ( .A(n25349), .B(n25350), .Z(n25348) );
  NANDN U25480 ( .A(n25350), .B(n25349), .Z(n25345) );
  ANDN U25481 ( .B(B[212]), .A(n78), .Z(n25129) );
  XNOR U25482 ( .A(n25137), .B(n25351), .Z(n25130) );
  XNOR U25483 ( .A(n25136), .B(n25134), .Z(n25351) );
  AND U25484 ( .A(n25352), .B(n25353), .Z(n25134) );
  NANDN U25485 ( .A(n25354), .B(n25355), .Z(n25353) );
  OR U25486 ( .A(n25356), .B(n25357), .Z(n25355) );
  NAND U25487 ( .A(n25357), .B(n25356), .Z(n25352) );
  ANDN U25488 ( .B(B[213]), .A(n79), .Z(n25136) );
  XNOR U25489 ( .A(n25144), .B(n25358), .Z(n25137) );
  XNOR U25490 ( .A(n25143), .B(n25141), .Z(n25358) );
  AND U25491 ( .A(n25359), .B(n25360), .Z(n25141) );
  NANDN U25492 ( .A(n25361), .B(n25362), .Z(n25360) );
  NANDN U25493 ( .A(n25363), .B(n25364), .Z(n25362) );
  NANDN U25494 ( .A(n25364), .B(n25363), .Z(n25359) );
  ANDN U25495 ( .B(B[214]), .A(n80), .Z(n25143) );
  XNOR U25496 ( .A(n25151), .B(n25365), .Z(n25144) );
  XNOR U25497 ( .A(n25150), .B(n25148), .Z(n25365) );
  AND U25498 ( .A(n25366), .B(n25367), .Z(n25148) );
  NANDN U25499 ( .A(n25368), .B(n25369), .Z(n25367) );
  OR U25500 ( .A(n25370), .B(n25371), .Z(n25369) );
  NAND U25501 ( .A(n25371), .B(n25370), .Z(n25366) );
  ANDN U25502 ( .B(B[215]), .A(n81), .Z(n25150) );
  XNOR U25503 ( .A(n25158), .B(n25372), .Z(n25151) );
  XNOR U25504 ( .A(n25157), .B(n25155), .Z(n25372) );
  AND U25505 ( .A(n25373), .B(n25374), .Z(n25155) );
  NANDN U25506 ( .A(n25375), .B(n25376), .Z(n25374) );
  NAND U25507 ( .A(n25377), .B(n25378), .Z(n25376) );
  ANDN U25508 ( .B(B[216]), .A(n82), .Z(n25157) );
  XOR U25509 ( .A(n25164), .B(n25379), .Z(n25158) );
  XNOR U25510 ( .A(n25162), .B(n25165), .Z(n25379) );
  NAND U25511 ( .A(A[2]), .B(B[217]), .Z(n25165) );
  NANDN U25512 ( .A(n25380), .B(n25381), .Z(n25162) );
  AND U25513 ( .A(A[0]), .B(B[218]), .Z(n25381) );
  XNOR U25514 ( .A(n25167), .B(n25382), .Z(n25164) );
  NAND U25515 ( .A(A[0]), .B(B[219]), .Z(n25382) );
  NAND U25516 ( .A(B[218]), .B(A[1]), .Z(n25167) );
  NAND U25517 ( .A(n25383), .B(n25384), .Z(n358) );
  NANDN U25518 ( .A(n25385), .B(n25386), .Z(n25384) );
  OR U25519 ( .A(n25387), .B(n25388), .Z(n25386) );
  NAND U25520 ( .A(n25388), .B(n25387), .Z(n25383) );
  XOR U25521 ( .A(n360), .B(n359), .Z(\A1[216] ) );
  XOR U25522 ( .A(n25388), .B(n25389), .Z(n359) );
  XNOR U25523 ( .A(n25387), .B(n25385), .Z(n25389) );
  AND U25524 ( .A(n25390), .B(n25391), .Z(n25385) );
  NANDN U25525 ( .A(n25392), .B(n25393), .Z(n25391) );
  NANDN U25526 ( .A(n25394), .B(n25395), .Z(n25393) );
  NANDN U25527 ( .A(n25395), .B(n25394), .Z(n25390) );
  ANDN U25528 ( .B(B[187]), .A(n54), .Z(n25387) );
  XNOR U25529 ( .A(n25182), .B(n25396), .Z(n25388) );
  XNOR U25530 ( .A(n25181), .B(n25179), .Z(n25396) );
  AND U25531 ( .A(n25397), .B(n25398), .Z(n25179) );
  NANDN U25532 ( .A(n25399), .B(n25400), .Z(n25398) );
  OR U25533 ( .A(n25401), .B(n25402), .Z(n25400) );
  NAND U25534 ( .A(n25402), .B(n25401), .Z(n25397) );
  ANDN U25535 ( .B(B[188]), .A(n55), .Z(n25181) );
  XNOR U25536 ( .A(n25189), .B(n25403), .Z(n25182) );
  XNOR U25537 ( .A(n25188), .B(n25186), .Z(n25403) );
  AND U25538 ( .A(n25404), .B(n25405), .Z(n25186) );
  NANDN U25539 ( .A(n25406), .B(n25407), .Z(n25405) );
  NANDN U25540 ( .A(n25408), .B(n25409), .Z(n25407) );
  NANDN U25541 ( .A(n25409), .B(n25408), .Z(n25404) );
  ANDN U25542 ( .B(B[189]), .A(n56), .Z(n25188) );
  XNOR U25543 ( .A(n25196), .B(n25410), .Z(n25189) );
  XNOR U25544 ( .A(n25195), .B(n25193), .Z(n25410) );
  AND U25545 ( .A(n25411), .B(n25412), .Z(n25193) );
  NANDN U25546 ( .A(n25413), .B(n25414), .Z(n25412) );
  OR U25547 ( .A(n25415), .B(n25416), .Z(n25414) );
  NAND U25548 ( .A(n25416), .B(n25415), .Z(n25411) );
  ANDN U25549 ( .B(B[190]), .A(n57), .Z(n25195) );
  XNOR U25550 ( .A(n25203), .B(n25417), .Z(n25196) );
  XNOR U25551 ( .A(n25202), .B(n25200), .Z(n25417) );
  AND U25552 ( .A(n25418), .B(n25419), .Z(n25200) );
  NANDN U25553 ( .A(n25420), .B(n25421), .Z(n25419) );
  NANDN U25554 ( .A(n25422), .B(n25423), .Z(n25421) );
  NANDN U25555 ( .A(n25423), .B(n25422), .Z(n25418) );
  ANDN U25556 ( .B(B[191]), .A(n58), .Z(n25202) );
  XNOR U25557 ( .A(n25210), .B(n25424), .Z(n25203) );
  XNOR U25558 ( .A(n25209), .B(n25207), .Z(n25424) );
  AND U25559 ( .A(n25425), .B(n25426), .Z(n25207) );
  NANDN U25560 ( .A(n25427), .B(n25428), .Z(n25426) );
  OR U25561 ( .A(n25429), .B(n25430), .Z(n25428) );
  NAND U25562 ( .A(n25430), .B(n25429), .Z(n25425) );
  ANDN U25563 ( .B(B[192]), .A(n59), .Z(n25209) );
  XNOR U25564 ( .A(n25217), .B(n25431), .Z(n25210) );
  XNOR U25565 ( .A(n25216), .B(n25214), .Z(n25431) );
  AND U25566 ( .A(n25432), .B(n25433), .Z(n25214) );
  NANDN U25567 ( .A(n25434), .B(n25435), .Z(n25433) );
  NANDN U25568 ( .A(n25436), .B(n25437), .Z(n25435) );
  NANDN U25569 ( .A(n25437), .B(n25436), .Z(n25432) );
  ANDN U25570 ( .B(B[193]), .A(n60), .Z(n25216) );
  XNOR U25571 ( .A(n25224), .B(n25438), .Z(n25217) );
  XNOR U25572 ( .A(n25223), .B(n25221), .Z(n25438) );
  AND U25573 ( .A(n25439), .B(n25440), .Z(n25221) );
  NANDN U25574 ( .A(n25441), .B(n25442), .Z(n25440) );
  OR U25575 ( .A(n25443), .B(n25444), .Z(n25442) );
  NAND U25576 ( .A(n25444), .B(n25443), .Z(n25439) );
  ANDN U25577 ( .B(B[194]), .A(n61), .Z(n25223) );
  XNOR U25578 ( .A(n25231), .B(n25445), .Z(n25224) );
  XNOR U25579 ( .A(n25230), .B(n25228), .Z(n25445) );
  AND U25580 ( .A(n25446), .B(n25447), .Z(n25228) );
  NANDN U25581 ( .A(n25448), .B(n25449), .Z(n25447) );
  NANDN U25582 ( .A(n25450), .B(n25451), .Z(n25449) );
  NANDN U25583 ( .A(n25451), .B(n25450), .Z(n25446) );
  ANDN U25584 ( .B(B[195]), .A(n62), .Z(n25230) );
  XNOR U25585 ( .A(n25238), .B(n25452), .Z(n25231) );
  XNOR U25586 ( .A(n25237), .B(n25235), .Z(n25452) );
  AND U25587 ( .A(n25453), .B(n25454), .Z(n25235) );
  NANDN U25588 ( .A(n25455), .B(n25456), .Z(n25454) );
  OR U25589 ( .A(n25457), .B(n25458), .Z(n25456) );
  NAND U25590 ( .A(n25458), .B(n25457), .Z(n25453) );
  ANDN U25591 ( .B(B[196]), .A(n63), .Z(n25237) );
  XNOR U25592 ( .A(n25245), .B(n25459), .Z(n25238) );
  XNOR U25593 ( .A(n25244), .B(n25242), .Z(n25459) );
  AND U25594 ( .A(n25460), .B(n25461), .Z(n25242) );
  NANDN U25595 ( .A(n25462), .B(n25463), .Z(n25461) );
  NANDN U25596 ( .A(n25464), .B(n25465), .Z(n25463) );
  NANDN U25597 ( .A(n25465), .B(n25464), .Z(n25460) );
  ANDN U25598 ( .B(B[197]), .A(n64), .Z(n25244) );
  XNOR U25599 ( .A(n25252), .B(n25466), .Z(n25245) );
  XNOR U25600 ( .A(n25251), .B(n25249), .Z(n25466) );
  AND U25601 ( .A(n25467), .B(n25468), .Z(n25249) );
  NANDN U25602 ( .A(n25469), .B(n25470), .Z(n25468) );
  OR U25603 ( .A(n25471), .B(n25472), .Z(n25470) );
  NAND U25604 ( .A(n25472), .B(n25471), .Z(n25467) );
  ANDN U25605 ( .B(B[198]), .A(n65), .Z(n25251) );
  XNOR U25606 ( .A(n25259), .B(n25473), .Z(n25252) );
  XNOR U25607 ( .A(n25258), .B(n25256), .Z(n25473) );
  AND U25608 ( .A(n25474), .B(n25475), .Z(n25256) );
  NANDN U25609 ( .A(n25476), .B(n25477), .Z(n25475) );
  NANDN U25610 ( .A(n25478), .B(n25479), .Z(n25477) );
  NANDN U25611 ( .A(n25479), .B(n25478), .Z(n25474) );
  ANDN U25612 ( .B(B[199]), .A(n66), .Z(n25258) );
  XNOR U25613 ( .A(n25266), .B(n25480), .Z(n25259) );
  XNOR U25614 ( .A(n25265), .B(n25263), .Z(n25480) );
  AND U25615 ( .A(n25481), .B(n25482), .Z(n25263) );
  NANDN U25616 ( .A(n25483), .B(n25484), .Z(n25482) );
  OR U25617 ( .A(n25485), .B(n25486), .Z(n25484) );
  NAND U25618 ( .A(n25486), .B(n25485), .Z(n25481) );
  ANDN U25619 ( .B(B[200]), .A(n67), .Z(n25265) );
  XNOR U25620 ( .A(n25273), .B(n25487), .Z(n25266) );
  XNOR U25621 ( .A(n25272), .B(n25270), .Z(n25487) );
  AND U25622 ( .A(n25488), .B(n25489), .Z(n25270) );
  NANDN U25623 ( .A(n25490), .B(n25491), .Z(n25489) );
  NANDN U25624 ( .A(n25492), .B(n25493), .Z(n25491) );
  NANDN U25625 ( .A(n25493), .B(n25492), .Z(n25488) );
  ANDN U25626 ( .B(B[201]), .A(n68), .Z(n25272) );
  XNOR U25627 ( .A(n25280), .B(n25494), .Z(n25273) );
  XNOR U25628 ( .A(n25279), .B(n25277), .Z(n25494) );
  AND U25629 ( .A(n25495), .B(n25496), .Z(n25277) );
  NANDN U25630 ( .A(n25497), .B(n25498), .Z(n25496) );
  OR U25631 ( .A(n25499), .B(n25500), .Z(n25498) );
  NAND U25632 ( .A(n25500), .B(n25499), .Z(n25495) );
  ANDN U25633 ( .B(B[202]), .A(n69), .Z(n25279) );
  XNOR U25634 ( .A(n25287), .B(n25501), .Z(n25280) );
  XNOR U25635 ( .A(n25286), .B(n25284), .Z(n25501) );
  AND U25636 ( .A(n25502), .B(n25503), .Z(n25284) );
  NANDN U25637 ( .A(n25504), .B(n25505), .Z(n25503) );
  NANDN U25638 ( .A(n25506), .B(n25507), .Z(n25505) );
  NANDN U25639 ( .A(n25507), .B(n25506), .Z(n25502) );
  ANDN U25640 ( .B(B[203]), .A(n70), .Z(n25286) );
  XNOR U25641 ( .A(n25294), .B(n25508), .Z(n25287) );
  XNOR U25642 ( .A(n25293), .B(n25291), .Z(n25508) );
  AND U25643 ( .A(n25509), .B(n25510), .Z(n25291) );
  NANDN U25644 ( .A(n25511), .B(n25512), .Z(n25510) );
  OR U25645 ( .A(n25513), .B(n25514), .Z(n25512) );
  NAND U25646 ( .A(n25514), .B(n25513), .Z(n25509) );
  ANDN U25647 ( .B(B[204]), .A(n71), .Z(n25293) );
  XNOR U25648 ( .A(n25301), .B(n25515), .Z(n25294) );
  XNOR U25649 ( .A(n25300), .B(n25298), .Z(n25515) );
  AND U25650 ( .A(n25516), .B(n25517), .Z(n25298) );
  NANDN U25651 ( .A(n25518), .B(n25519), .Z(n25517) );
  NANDN U25652 ( .A(n25520), .B(n25521), .Z(n25519) );
  NANDN U25653 ( .A(n25521), .B(n25520), .Z(n25516) );
  ANDN U25654 ( .B(B[205]), .A(n72), .Z(n25300) );
  XNOR U25655 ( .A(n25308), .B(n25522), .Z(n25301) );
  XNOR U25656 ( .A(n25307), .B(n25305), .Z(n25522) );
  AND U25657 ( .A(n25523), .B(n25524), .Z(n25305) );
  NANDN U25658 ( .A(n25525), .B(n25526), .Z(n25524) );
  OR U25659 ( .A(n25527), .B(n25528), .Z(n25526) );
  NAND U25660 ( .A(n25528), .B(n25527), .Z(n25523) );
  ANDN U25661 ( .B(B[206]), .A(n73), .Z(n25307) );
  XNOR U25662 ( .A(n25315), .B(n25529), .Z(n25308) );
  XNOR U25663 ( .A(n25314), .B(n25312), .Z(n25529) );
  AND U25664 ( .A(n25530), .B(n25531), .Z(n25312) );
  NANDN U25665 ( .A(n25532), .B(n25533), .Z(n25531) );
  NANDN U25666 ( .A(n25534), .B(n25535), .Z(n25533) );
  NANDN U25667 ( .A(n25535), .B(n25534), .Z(n25530) );
  ANDN U25668 ( .B(B[207]), .A(n74), .Z(n25314) );
  XNOR U25669 ( .A(n25322), .B(n25536), .Z(n25315) );
  XNOR U25670 ( .A(n25321), .B(n25319), .Z(n25536) );
  AND U25671 ( .A(n25537), .B(n25538), .Z(n25319) );
  NANDN U25672 ( .A(n25539), .B(n25540), .Z(n25538) );
  OR U25673 ( .A(n25541), .B(n25542), .Z(n25540) );
  NAND U25674 ( .A(n25542), .B(n25541), .Z(n25537) );
  ANDN U25675 ( .B(B[208]), .A(n75), .Z(n25321) );
  XNOR U25676 ( .A(n25329), .B(n25543), .Z(n25322) );
  XNOR U25677 ( .A(n25328), .B(n25326), .Z(n25543) );
  AND U25678 ( .A(n25544), .B(n25545), .Z(n25326) );
  NANDN U25679 ( .A(n25546), .B(n25547), .Z(n25545) );
  NANDN U25680 ( .A(n25548), .B(n25549), .Z(n25547) );
  NANDN U25681 ( .A(n25549), .B(n25548), .Z(n25544) );
  ANDN U25682 ( .B(B[209]), .A(n76), .Z(n25328) );
  XNOR U25683 ( .A(n25336), .B(n25550), .Z(n25329) );
  XNOR U25684 ( .A(n25335), .B(n25333), .Z(n25550) );
  AND U25685 ( .A(n25551), .B(n25552), .Z(n25333) );
  NANDN U25686 ( .A(n25553), .B(n25554), .Z(n25552) );
  OR U25687 ( .A(n25555), .B(n25556), .Z(n25554) );
  NAND U25688 ( .A(n25556), .B(n25555), .Z(n25551) );
  ANDN U25689 ( .B(B[210]), .A(n77), .Z(n25335) );
  XNOR U25690 ( .A(n25343), .B(n25557), .Z(n25336) );
  XNOR U25691 ( .A(n25342), .B(n25340), .Z(n25557) );
  AND U25692 ( .A(n25558), .B(n25559), .Z(n25340) );
  NANDN U25693 ( .A(n25560), .B(n25561), .Z(n25559) );
  NANDN U25694 ( .A(n25562), .B(n25563), .Z(n25561) );
  NANDN U25695 ( .A(n25563), .B(n25562), .Z(n25558) );
  ANDN U25696 ( .B(B[211]), .A(n78), .Z(n25342) );
  XNOR U25697 ( .A(n25350), .B(n25564), .Z(n25343) );
  XNOR U25698 ( .A(n25349), .B(n25347), .Z(n25564) );
  AND U25699 ( .A(n25565), .B(n25566), .Z(n25347) );
  NANDN U25700 ( .A(n25567), .B(n25568), .Z(n25566) );
  OR U25701 ( .A(n25569), .B(n25570), .Z(n25568) );
  NAND U25702 ( .A(n25570), .B(n25569), .Z(n25565) );
  ANDN U25703 ( .B(B[212]), .A(n79), .Z(n25349) );
  XNOR U25704 ( .A(n25357), .B(n25571), .Z(n25350) );
  XNOR U25705 ( .A(n25356), .B(n25354), .Z(n25571) );
  AND U25706 ( .A(n25572), .B(n25573), .Z(n25354) );
  NANDN U25707 ( .A(n25574), .B(n25575), .Z(n25573) );
  NANDN U25708 ( .A(n25576), .B(n25577), .Z(n25575) );
  NANDN U25709 ( .A(n25577), .B(n25576), .Z(n25572) );
  ANDN U25710 ( .B(B[213]), .A(n80), .Z(n25356) );
  XNOR U25711 ( .A(n25364), .B(n25578), .Z(n25357) );
  XNOR U25712 ( .A(n25363), .B(n25361), .Z(n25578) );
  AND U25713 ( .A(n25579), .B(n25580), .Z(n25361) );
  NANDN U25714 ( .A(n25581), .B(n25582), .Z(n25580) );
  OR U25715 ( .A(n25583), .B(n25584), .Z(n25582) );
  NAND U25716 ( .A(n25584), .B(n25583), .Z(n25579) );
  ANDN U25717 ( .B(B[214]), .A(n81), .Z(n25363) );
  XNOR U25718 ( .A(n25371), .B(n25585), .Z(n25364) );
  XNOR U25719 ( .A(n25370), .B(n25368), .Z(n25585) );
  AND U25720 ( .A(n25586), .B(n25587), .Z(n25368) );
  NANDN U25721 ( .A(n25588), .B(n25589), .Z(n25587) );
  NAND U25722 ( .A(n25590), .B(n25591), .Z(n25589) );
  ANDN U25723 ( .B(B[215]), .A(n82), .Z(n25370) );
  XOR U25724 ( .A(n25377), .B(n25592), .Z(n25371) );
  XNOR U25725 ( .A(n25375), .B(n25378), .Z(n25592) );
  NAND U25726 ( .A(A[2]), .B(B[216]), .Z(n25378) );
  NANDN U25727 ( .A(n25593), .B(n25594), .Z(n25375) );
  AND U25728 ( .A(A[0]), .B(B[217]), .Z(n25594) );
  XNOR U25729 ( .A(n25380), .B(n25595), .Z(n25377) );
  NAND U25730 ( .A(A[0]), .B(B[218]), .Z(n25595) );
  NAND U25731 ( .A(B[217]), .B(A[1]), .Z(n25380) );
  NAND U25732 ( .A(n25596), .B(n25597), .Z(n360) );
  NANDN U25733 ( .A(n25598), .B(n25599), .Z(n25597) );
  OR U25734 ( .A(n25600), .B(n25601), .Z(n25599) );
  NAND U25735 ( .A(n25601), .B(n25600), .Z(n25596) );
  XOR U25736 ( .A(n362), .B(n361), .Z(\A1[215] ) );
  XOR U25737 ( .A(n25601), .B(n25602), .Z(n361) );
  XNOR U25738 ( .A(n25600), .B(n25598), .Z(n25602) );
  AND U25739 ( .A(n25603), .B(n25604), .Z(n25598) );
  NANDN U25740 ( .A(n25605), .B(n25606), .Z(n25604) );
  NANDN U25741 ( .A(n25607), .B(n25608), .Z(n25606) );
  NANDN U25742 ( .A(n25608), .B(n25607), .Z(n25603) );
  ANDN U25743 ( .B(B[186]), .A(n54), .Z(n25600) );
  XNOR U25744 ( .A(n25395), .B(n25609), .Z(n25601) );
  XNOR U25745 ( .A(n25394), .B(n25392), .Z(n25609) );
  AND U25746 ( .A(n25610), .B(n25611), .Z(n25392) );
  NANDN U25747 ( .A(n25612), .B(n25613), .Z(n25611) );
  OR U25748 ( .A(n25614), .B(n25615), .Z(n25613) );
  NAND U25749 ( .A(n25615), .B(n25614), .Z(n25610) );
  ANDN U25750 ( .B(B[187]), .A(n55), .Z(n25394) );
  XNOR U25751 ( .A(n25402), .B(n25616), .Z(n25395) );
  XNOR U25752 ( .A(n25401), .B(n25399), .Z(n25616) );
  AND U25753 ( .A(n25617), .B(n25618), .Z(n25399) );
  NANDN U25754 ( .A(n25619), .B(n25620), .Z(n25618) );
  NANDN U25755 ( .A(n25621), .B(n25622), .Z(n25620) );
  NANDN U25756 ( .A(n25622), .B(n25621), .Z(n25617) );
  ANDN U25757 ( .B(B[188]), .A(n56), .Z(n25401) );
  XNOR U25758 ( .A(n25409), .B(n25623), .Z(n25402) );
  XNOR U25759 ( .A(n25408), .B(n25406), .Z(n25623) );
  AND U25760 ( .A(n25624), .B(n25625), .Z(n25406) );
  NANDN U25761 ( .A(n25626), .B(n25627), .Z(n25625) );
  OR U25762 ( .A(n25628), .B(n25629), .Z(n25627) );
  NAND U25763 ( .A(n25629), .B(n25628), .Z(n25624) );
  ANDN U25764 ( .B(B[189]), .A(n57), .Z(n25408) );
  XNOR U25765 ( .A(n25416), .B(n25630), .Z(n25409) );
  XNOR U25766 ( .A(n25415), .B(n25413), .Z(n25630) );
  AND U25767 ( .A(n25631), .B(n25632), .Z(n25413) );
  NANDN U25768 ( .A(n25633), .B(n25634), .Z(n25632) );
  NANDN U25769 ( .A(n25635), .B(n25636), .Z(n25634) );
  NANDN U25770 ( .A(n25636), .B(n25635), .Z(n25631) );
  ANDN U25771 ( .B(B[190]), .A(n58), .Z(n25415) );
  XNOR U25772 ( .A(n25423), .B(n25637), .Z(n25416) );
  XNOR U25773 ( .A(n25422), .B(n25420), .Z(n25637) );
  AND U25774 ( .A(n25638), .B(n25639), .Z(n25420) );
  NANDN U25775 ( .A(n25640), .B(n25641), .Z(n25639) );
  OR U25776 ( .A(n25642), .B(n25643), .Z(n25641) );
  NAND U25777 ( .A(n25643), .B(n25642), .Z(n25638) );
  ANDN U25778 ( .B(B[191]), .A(n59), .Z(n25422) );
  XNOR U25779 ( .A(n25430), .B(n25644), .Z(n25423) );
  XNOR U25780 ( .A(n25429), .B(n25427), .Z(n25644) );
  AND U25781 ( .A(n25645), .B(n25646), .Z(n25427) );
  NANDN U25782 ( .A(n25647), .B(n25648), .Z(n25646) );
  NANDN U25783 ( .A(n25649), .B(n25650), .Z(n25648) );
  NANDN U25784 ( .A(n25650), .B(n25649), .Z(n25645) );
  ANDN U25785 ( .B(B[192]), .A(n60), .Z(n25429) );
  XNOR U25786 ( .A(n25437), .B(n25651), .Z(n25430) );
  XNOR U25787 ( .A(n25436), .B(n25434), .Z(n25651) );
  AND U25788 ( .A(n25652), .B(n25653), .Z(n25434) );
  NANDN U25789 ( .A(n25654), .B(n25655), .Z(n25653) );
  OR U25790 ( .A(n25656), .B(n25657), .Z(n25655) );
  NAND U25791 ( .A(n25657), .B(n25656), .Z(n25652) );
  ANDN U25792 ( .B(B[193]), .A(n61), .Z(n25436) );
  XNOR U25793 ( .A(n25444), .B(n25658), .Z(n25437) );
  XNOR U25794 ( .A(n25443), .B(n25441), .Z(n25658) );
  AND U25795 ( .A(n25659), .B(n25660), .Z(n25441) );
  NANDN U25796 ( .A(n25661), .B(n25662), .Z(n25660) );
  NANDN U25797 ( .A(n25663), .B(n25664), .Z(n25662) );
  NANDN U25798 ( .A(n25664), .B(n25663), .Z(n25659) );
  ANDN U25799 ( .B(B[194]), .A(n62), .Z(n25443) );
  XNOR U25800 ( .A(n25451), .B(n25665), .Z(n25444) );
  XNOR U25801 ( .A(n25450), .B(n25448), .Z(n25665) );
  AND U25802 ( .A(n25666), .B(n25667), .Z(n25448) );
  NANDN U25803 ( .A(n25668), .B(n25669), .Z(n25667) );
  OR U25804 ( .A(n25670), .B(n25671), .Z(n25669) );
  NAND U25805 ( .A(n25671), .B(n25670), .Z(n25666) );
  ANDN U25806 ( .B(B[195]), .A(n63), .Z(n25450) );
  XNOR U25807 ( .A(n25458), .B(n25672), .Z(n25451) );
  XNOR U25808 ( .A(n25457), .B(n25455), .Z(n25672) );
  AND U25809 ( .A(n25673), .B(n25674), .Z(n25455) );
  NANDN U25810 ( .A(n25675), .B(n25676), .Z(n25674) );
  NANDN U25811 ( .A(n25677), .B(n25678), .Z(n25676) );
  NANDN U25812 ( .A(n25678), .B(n25677), .Z(n25673) );
  ANDN U25813 ( .B(B[196]), .A(n64), .Z(n25457) );
  XNOR U25814 ( .A(n25465), .B(n25679), .Z(n25458) );
  XNOR U25815 ( .A(n25464), .B(n25462), .Z(n25679) );
  AND U25816 ( .A(n25680), .B(n25681), .Z(n25462) );
  NANDN U25817 ( .A(n25682), .B(n25683), .Z(n25681) );
  OR U25818 ( .A(n25684), .B(n25685), .Z(n25683) );
  NAND U25819 ( .A(n25685), .B(n25684), .Z(n25680) );
  ANDN U25820 ( .B(B[197]), .A(n65), .Z(n25464) );
  XNOR U25821 ( .A(n25472), .B(n25686), .Z(n25465) );
  XNOR U25822 ( .A(n25471), .B(n25469), .Z(n25686) );
  AND U25823 ( .A(n25687), .B(n25688), .Z(n25469) );
  NANDN U25824 ( .A(n25689), .B(n25690), .Z(n25688) );
  NANDN U25825 ( .A(n25691), .B(n25692), .Z(n25690) );
  NANDN U25826 ( .A(n25692), .B(n25691), .Z(n25687) );
  ANDN U25827 ( .B(B[198]), .A(n66), .Z(n25471) );
  XNOR U25828 ( .A(n25479), .B(n25693), .Z(n25472) );
  XNOR U25829 ( .A(n25478), .B(n25476), .Z(n25693) );
  AND U25830 ( .A(n25694), .B(n25695), .Z(n25476) );
  NANDN U25831 ( .A(n25696), .B(n25697), .Z(n25695) );
  OR U25832 ( .A(n25698), .B(n25699), .Z(n25697) );
  NAND U25833 ( .A(n25699), .B(n25698), .Z(n25694) );
  ANDN U25834 ( .B(B[199]), .A(n67), .Z(n25478) );
  XNOR U25835 ( .A(n25486), .B(n25700), .Z(n25479) );
  XNOR U25836 ( .A(n25485), .B(n25483), .Z(n25700) );
  AND U25837 ( .A(n25701), .B(n25702), .Z(n25483) );
  NANDN U25838 ( .A(n25703), .B(n25704), .Z(n25702) );
  NANDN U25839 ( .A(n25705), .B(n25706), .Z(n25704) );
  NANDN U25840 ( .A(n25706), .B(n25705), .Z(n25701) );
  ANDN U25841 ( .B(B[200]), .A(n68), .Z(n25485) );
  XNOR U25842 ( .A(n25493), .B(n25707), .Z(n25486) );
  XNOR U25843 ( .A(n25492), .B(n25490), .Z(n25707) );
  AND U25844 ( .A(n25708), .B(n25709), .Z(n25490) );
  NANDN U25845 ( .A(n25710), .B(n25711), .Z(n25709) );
  OR U25846 ( .A(n25712), .B(n25713), .Z(n25711) );
  NAND U25847 ( .A(n25713), .B(n25712), .Z(n25708) );
  ANDN U25848 ( .B(B[201]), .A(n69), .Z(n25492) );
  XNOR U25849 ( .A(n25500), .B(n25714), .Z(n25493) );
  XNOR U25850 ( .A(n25499), .B(n25497), .Z(n25714) );
  AND U25851 ( .A(n25715), .B(n25716), .Z(n25497) );
  NANDN U25852 ( .A(n25717), .B(n25718), .Z(n25716) );
  NANDN U25853 ( .A(n25719), .B(n25720), .Z(n25718) );
  NANDN U25854 ( .A(n25720), .B(n25719), .Z(n25715) );
  ANDN U25855 ( .B(B[202]), .A(n70), .Z(n25499) );
  XNOR U25856 ( .A(n25507), .B(n25721), .Z(n25500) );
  XNOR U25857 ( .A(n25506), .B(n25504), .Z(n25721) );
  AND U25858 ( .A(n25722), .B(n25723), .Z(n25504) );
  NANDN U25859 ( .A(n25724), .B(n25725), .Z(n25723) );
  OR U25860 ( .A(n25726), .B(n25727), .Z(n25725) );
  NAND U25861 ( .A(n25727), .B(n25726), .Z(n25722) );
  ANDN U25862 ( .B(B[203]), .A(n71), .Z(n25506) );
  XNOR U25863 ( .A(n25514), .B(n25728), .Z(n25507) );
  XNOR U25864 ( .A(n25513), .B(n25511), .Z(n25728) );
  AND U25865 ( .A(n25729), .B(n25730), .Z(n25511) );
  NANDN U25866 ( .A(n25731), .B(n25732), .Z(n25730) );
  NANDN U25867 ( .A(n25733), .B(n25734), .Z(n25732) );
  NANDN U25868 ( .A(n25734), .B(n25733), .Z(n25729) );
  ANDN U25869 ( .B(B[204]), .A(n72), .Z(n25513) );
  XNOR U25870 ( .A(n25521), .B(n25735), .Z(n25514) );
  XNOR U25871 ( .A(n25520), .B(n25518), .Z(n25735) );
  AND U25872 ( .A(n25736), .B(n25737), .Z(n25518) );
  NANDN U25873 ( .A(n25738), .B(n25739), .Z(n25737) );
  OR U25874 ( .A(n25740), .B(n25741), .Z(n25739) );
  NAND U25875 ( .A(n25741), .B(n25740), .Z(n25736) );
  ANDN U25876 ( .B(B[205]), .A(n73), .Z(n25520) );
  XNOR U25877 ( .A(n25528), .B(n25742), .Z(n25521) );
  XNOR U25878 ( .A(n25527), .B(n25525), .Z(n25742) );
  AND U25879 ( .A(n25743), .B(n25744), .Z(n25525) );
  NANDN U25880 ( .A(n25745), .B(n25746), .Z(n25744) );
  NANDN U25881 ( .A(n25747), .B(n25748), .Z(n25746) );
  NANDN U25882 ( .A(n25748), .B(n25747), .Z(n25743) );
  ANDN U25883 ( .B(B[206]), .A(n74), .Z(n25527) );
  XNOR U25884 ( .A(n25535), .B(n25749), .Z(n25528) );
  XNOR U25885 ( .A(n25534), .B(n25532), .Z(n25749) );
  AND U25886 ( .A(n25750), .B(n25751), .Z(n25532) );
  NANDN U25887 ( .A(n25752), .B(n25753), .Z(n25751) );
  OR U25888 ( .A(n25754), .B(n25755), .Z(n25753) );
  NAND U25889 ( .A(n25755), .B(n25754), .Z(n25750) );
  ANDN U25890 ( .B(B[207]), .A(n75), .Z(n25534) );
  XNOR U25891 ( .A(n25542), .B(n25756), .Z(n25535) );
  XNOR U25892 ( .A(n25541), .B(n25539), .Z(n25756) );
  AND U25893 ( .A(n25757), .B(n25758), .Z(n25539) );
  NANDN U25894 ( .A(n25759), .B(n25760), .Z(n25758) );
  NANDN U25895 ( .A(n25761), .B(n25762), .Z(n25760) );
  NANDN U25896 ( .A(n25762), .B(n25761), .Z(n25757) );
  ANDN U25897 ( .B(B[208]), .A(n76), .Z(n25541) );
  XNOR U25898 ( .A(n25549), .B(n25763), .Z(n25542) );
  XNOR U25899 ( .A(n25548), .B(n25546), .Z(n25763) );
  AND U25900 ( .A(n25764), .B(n25765), .Z(n25546) );
  NANDN U25901 ( .A(n25766), .B(n25767), .Z(n25765) );
  OR U25902 ( .A(n25768), .B(n25769), .Z(n25767) );
  NAND U25903 ( .A(n25769), .B(n25768), .Z(n25764) );
  ANDN U25904 ( .B(B[209]), .A(n77), .Z(n25548) );
  XNOR U25905 ( .A(n25556), .B(n25770), .Z(n25549) );
  XNOR U25906 ( .A(n25555), .B(n25553), .Z(n25770) );
  AND U25907 ( .A(n25771), .B(n25772), .Z(n25553) );
  NANDN U25908 ( .A(n25773), .B(n25774), .Z(n25772) );
  NANDN U25909 ( .A(n25775), .B(n25776), .Z(n25774) );
  NANDN U25910 ( .A(n25776), .B(n25775), .Z(n25771) );
  ANDN U25911 ( .B(B[210]), .A(n78), .Z(n25555) );
  XNOR U25912 ( .A(n25563), .B(n25777), .Z(n25556) );
  XNOR U25913 ( .A(n25562), .B(n25560), .Z(n25777) );
  AND U25914 ( .A(n25778), .B(n25779), .Z(n25560) );
  NANDN U25915 ( .A(n25780), .B(n25781), .Z(n25779) );
  OR U25916 ( .A(n25782), .B(n25783), .Z(n25781) );
  NAND U25917 ( .A(n25783), .B(n25782), .Z(n25778) );
  ANDN U25918 ( .B(B[211]), .A(n79), .Z(n25562) );
  XNOR U25919 ( .A(n25570), .B(n25784), .Z(n25563) );
  XNOR U25920 ( .A(n25569), .B(n25567), .Z(n25784) );
  AND U25921 ( .A(n25785), .B(n25786), .Z(n25567) );
  NANDN U25922 ( .A(n25787), .B(n25788), .Z(n25786) );
  NANDN U25923 ( .A(n25789), .B(n25790), .Z(n25788) );
  NANDN U25924 ( .A(n25790), .B(n25789), .Z(n25785) );
  ANDN U25925 ( .B(B[212]), .A(n80), .Z(n25569) );
  XNOR U25926 ( .A(n25577), .B(n25791), .Z(n25570) );
  XNOR U25927 ( .A(n25576), .B(n25574), .Z(n25791) );
  AND U25928 ( .A(n25792), .B(n25793), .Z(n25574) );
  NANDN U25929 ( .A(n25794), .B(n25795), .Z(n25793) );
  OR U25930 ( .A(n25796), .B(n25797), .Z(n25795) );
  NAND U25931 ( .A(n25797), .B(n25796), .Z(n25792) );
  ANDN U25932 ( .B(B[213]), .A(n81), .Z(n25576) );
  XNOR U25933 ( .A(n25584), .B(n25798), .Z(n25577) );
  XNOR U25934 ( .A(n25583), .B(n25581), .Z(n25798) );
  AND U25935 ( .A(n25799), .B(n25800), .Z(n25581) );
  NANDN U25936 ( .A(n25801), .B(n25802), .Z(n25800) );
  NAND U25937 ( .A(n25803), .B(n25804), .Z(n25802) );
  ANDN U25938 ( .B(B[214]), .A(n82), .Z(n25583) );
  XOR U25939 ( .A(n25590), .B(n25805), .Z(n25584) );
  XNOR U25940 ( .A(n25588), .B(n25591), .Z(n25805) );
  NAND U25941 ( .A(A[2]), .B(B[215]), .Z(n25591) );
  NANDN U25942 ( .A(n25806), .B(n25807), .Z(n25588) );
  AND U25943 ( .A(A[0]), .B(B[216]), .Z(n25807) );
  XNOR U25944 ( .A(n25593), .B(n25808), .Z(n25590) );
  NAND U25945 ( .A(A[0]), .B(B[217]), .Z(n25808) );
  NAND U25946 ( .A(B[216]), .B(A[1]), .Z(n25593) );
  NAND U25947 ( .A(n25809), .B(n25810), .Z(n362) );
  NANDN U25948 ( .A(n25811), .B(n25812), .Z(n25810) );
  OR U25949 ( .A(n25813), .B(n25814), .Z(n25812) );
  NAND U25950 ( .A(n25814), .B(n25813), .Z(n25809) );
  XOR U25951 ( .A(n364), .B(n363), .Z(\A1[214] ) );
  XOR U25952 ( .A(n25814), .B(n25815), .Z(n363) );
  XNOR U25953 ( .A(n25813), .B(n25811), .Z(n25815) );
  AND U25954 ( .A(n25816), .B(n25817), .Z(n25811) );
  NANDN U25955 ( .A(n25818), .B(n25819), .Z(n25817) );
  NANDN U25956 ( .A(n25820), .B(n25821), .Z(n25819) );
  NANDN U25957 ( .A(n25821), .B(n25820), .Z(n25816) );
  ANDN U25958 ( .B(B[185]), .A(n54), .Z(n25813) );
  XNOR U25959 ( .A(n25608), .B(n25822), .Z(n25814) );
  XNOR U25960 ( .A(n25607), .B(n25605), .Z(n25822) );
  AND U25961 ( .A(n25823), .B(n25824), .Z(n25605) );
  NANDN U25962 ( .A(n25825), .B(n25826), .Z(n25824) );
  OR U25963 ( .A(n25827), .B(n25828), .Z(n25826) );
  NAND U25964 ( .A(n25828), .B(n25827), .Z(n25823) );
  ANDN U25965 ( .B(B[186]), .A(n55), .Z(n25607) );
  XNOR U25966 ( .A(n25615), .B(n25829), .Z(n25608) );
  XNOR U25967 ( .A(n25614), .B(n25612), .Z(n25829) );
  AND U25968 ( .A(n25830), .B(n25831), .Z(n25612) );
  NANDN U25969 ( .A(n25832), .B(n25833), .Z(n25831) );
  NANDN U25970 ( .A(n25834), .B(n25835), .Z(n25833) );
  NANDN U25971 ( .A(n25835), .B(n25834), .Z(n25830) );
  ANDN U25972 ( .B(B[187]), .A(n56), .Z(n25614) );
  XNOR U25973 ( .A(n25622), .B(n25836), .Z(n25615) );
  XNOR U25974 ( .A(n25621), .B(n25619), .Z(n25836) );
  AND U25975 ( .A(n25837), .B(n25838), .Z(n25619) );
  NANDN U25976 ( .A(n25839), .B(n25840), .Z(n25838) );
  OR U25977 ( .A(n25841), .B(n25842), .Z(n25840) );
  NAND U25978 ( .A(n25842), .B(n25841), .Z(n25837) );
  ANDN U25979 ( .B(B[188]), .A(n57), .Z(n25621) );
  XNOR U25980 ( .A(n25629), .B(n25843), .Z(n25622) );
  XNOR U25981 ( .A(n25628), .B(n25626), .Z(n25843) );
  AND U25982 ( .A(n25844), .B(n25845), .Z(n25626) );
  NANDN U25983 ( .A(n25846), .B(n25847), .Z(n25845) );
  NANDN U25984 ( .A(n25848), .B(n25849), .Z(n25847) );
  NANDN U25985 ( .A(n25849), .B(n25848), .Z(n25844) );
  ANDN U25986 ( .B(B[189]), .A(n58), .Z(n25628) );
  XNOR U25987 ( .A(n25636), .B(n25850), .Z(n25629) );
  XNOR U25988 ( .A(n25635), .B(n25633), .Z(n25850) );
  AND U25989 ( .A(n25851), .B(n25852), .Z(n25633) );
  NANDN U25990 ( .A(n25853), .B(n25854), .Z(n25852) );
  OR U25991 ( .A(n25855), .B(n25856), .Z(n25854) );
  NAND U25992 ( .A(n25856), .B(n25855), .Z(n25851) );
  ANDN U25993 ( .B(B[190]), .A(n59), .Z(n25635) );
  XNOR U25994 ( .A(n25643), .B(n25857), .Z(n25636) );
  XNOR U25995 ( .A(n25642), .B(n25640), .Z(n25857) );
  AND U25996 ( .A(n25858), .B(n25859), .Z(n25640) );
  NANDN U25997 ( .A(n25860), .B(n25861), .Z(n25859) );
  NANDN U25998 ( .A(n25862), .B(n25863), .Z(n25861) );
  NANDN U25999 ( .A(n25863), .B(n25862), .Z(n25858) );
  ANDN U26000 ( .B(B[191]), .A(n60), .Z(n25642) );
  XNOR U26001 ( .A(n25650), .B(n25864), .Z(n25643) );
  XNOR U26002 ( .A(n25649), .B(n25647), .Z(n25864) );
  AND U26003 ( .A(n25865), .B(n25866), .Z(n25647) );
  NANDN U26004 ( .A(n25867), .B(n25868), .Z(n25866) );
  OR U26005 ( .A(n25869), .B(n25870), .Z(n25868) );
  NAND U26006 ( .A(n25870), .B(n25869), .Z(n25865) );
  ANDN U26007 ( .B(B[192]), .A(n61), .Z(n25649) );
  XNOR U26008 ( .A(n25657), .B(n25871), .Z(n25650) );
  XNOR U26009 ( .A(n25656), .B(n25654), .Z(n25871) );
  AND U26010 ( .A(n25872), .B(n25873), .Z(n25654) );
  NANDN U26011 ( .A(n25874), .B(n25875), .Z(n25873) );
  NANDN U26012 ( .A(n25876), .B(n25877), .Z(n25875) );
  NANDN U26013 ( .A(n25877), .B(n25876), .Z(n25872) );
  ANDN U26014 ( .B(B[193]), .A(n62), .Z(n25656) );
  XNOR U26015 ( .A(n25664), .B(n25878), .Z(n25657) );
  XNOR U26016 ( .A(n25663), .B(n25661), .Z(n25878) );
  AND U26017 ( .A(n25879), .B(n25880), .Z(n25661) );
  NANDN U26018 ( .A(n25881), .B(n25882), .Z(n25880) );
  OR U26019 ( .A(n25883), .B(n25884), .Z(n25882) );
  NAND U26020 ( .A(n25884), .B(n25883), .Z(n25879) );
  ANDN U26021 ( .B(B[194]), .A(n63), .Z(n25663) );
  XNOR U26022 ( .A(n25671), .B(n25885), .Z(n25664) );
  XNOR U26023 ( .A(n25670), .B(n25668), .Z(n25885) );
  AND U26024 ( .A(n25886), .B(n25887), .Z(n25668) );
  NANDN U26025 ( .A(n25888), .B(n25889), .Z(n25887) );
  NANDN U26026 ( .A(n25890), .B(n25891), .Z(n25889) );
  NANDN U26027 ( .A(n25891), .B(n25890), .Z(n25886) );
  ANDN U26028 ( .B(B[195]), .A(n64), .Z(n25670) );
  XNOR U26029 ( .A(n25678), .B(n25892), .Z(n25671) );
  XNOR U26030 ( .A(n25677), .B(n25675), .Z(n25892) );
  AND U26031 ( .A(n25893), .B(n25894), .Z(n25675) );
  NANDN U26032 ( .A(n25895), .B(n25896), .Z(n25894) );
  OR U26033 ( .A(n25897), .B(n25898), .Z(n25896) );
  NAND U26034 ( .A(n25898), .B(n25897), .Z(n25893) );
  ANDN U26035 ( .B(B[196]), .A(n65), .Z(n25677) );
  XNOR U26036 ( .A(n25685), .B(n25899), .Z(n25678) );
  XNOR U26037 ( .A(n25684), .B(n25682), .Z(n25899) );
  AND U26038 ( .A(n25900), .B(n25901), .Z(n25682) );
  NANDN U26039 ( .A(n25902), .B(n25903), .Z(n25901) );
  NANDN U26040 ( .A(n25904), .B(n25905), .Z(n25903) );
  NANDN U26041 ( .A(n25905), .B(n25904), .Z(n25900) );
  ANDN U26042 ( .B(B[197]), .A(n66), .Z(n25684) );
  XNOR U26043 ( .A(n25692), .B(n25906), .Z(n25685) );
  XNOR U26044 ( .A(n25691), .B(n25689), .Z(n25906) );
  AND U26045 ( .A(n25907), .B(n25908), .Z(n25689) );
  NANDN U26046 ( .A(n25909), .B(n25910), .Z(n25908) );
  OR U26047 ( .A(n25911), .B(n25912), .Z(n25910) );
  NAND U26048 ( .A(n25912), .B(n25911), .Z(n25907) );
  ANDN U26049 ( .B(B[198]), .A(n67), .Z(n25691) );
  XNOR U26050 ( .A(n25699), .B(n25913), .Z(n25692) );
  XNOR U26051 ( .A(n25698), .B(n25696), .Z(n25913) );
  AND U26052 ( .A(n25914), .B(n25915), .Z(n25696) );
  NANDN U26053 ( .A(n25916), .B(n25917), .Z(n25915) );
  NANDN U26054 ( .A(n25918), .B(n25919), .Z(n25917) );
  NANDN U26055 ( .A(n25919), .B(n25918), .Z(n25914) );
  ANDN U26056 ( .B(B[199]), .A(n68), .Z(n25698) );
  XNOR U26057 ( .A(n25706), .B(n25920), .Z(n25699) );
  XNOR U26058 ( .A(n25705), .B(n25703), .Z(n25920) );
  AND U26059 ( .A(n25921), .B(n25922), .Z(n25703) );
  NANDN U26060 ( .A(n25923), .B(n25924), .Z(n25922) );
  OR U26061 ( .A(n25925), .B(n25926), .Z(n25924) );
  NAND U26062 ( .A(n25926), .B(n25925), .Z(n25921) );
  ANDN U26063 ( .B(B[200]), .A(n69), .Z(n25705) );
  XNOR U26064 ( .A(n25713), .B(n25927), .Z(n25706) );
  XNOR U26065 ( .A(n25712), .B(n25710), .Z(n25927) );
  AND U26066 ( .A(n25928), .B(n25929), .Z(n25710) );
  NANDN U26067 ( .A(n25930), .B(n25931), .Z(n25929) );
  NANDN U26068 ( .A(n25932), .B(n25933), .Z(n25931) );
  NANDN U26069 ( .A(n25933), .B(n25932), .Z(n25928) );
  ANDN U26070 ( .B(B[201]), .A(n70), .Z(n25712) );
  XNOR U26071 ( .A(n25720), .B(n25934), .Z(n25713) );
  XNOR U26072 ( .A(n25719), .B(n25717), .Z(n25934) );
  AND U26073 ( .A(n25935), .B(n25936), .Z(n25717) );
  NANDN U26074 ( .A(n25937), .B(n25938), .Z(n25936) );
  OR U26075 ( .A(n25939), .B(n25940), .Z(n25938) );
  NAND U26076 ( .A(n25940), .B(n25939), .Z(n25935) );
  ANDN U26077 ( .B(B[202]), .A(n71), .Z(n25719) );
  XNOR U26078 ( .A(n25727), .B(n25941), .Z(n25720) );
  XNOR U26079 ( .A(n25726), .B(n25724), .Z(n25941) );
  AND U26080 ( .A(n25942), .B(n25943), .Z(n25724) );
  NANDN U26081 ( .A(n25944), .B(n25945), .Z(n25943) );
  NANDN U26082 ( .A(n25946), .B(n25947), .Z(n25945) );
  NANDN U26083 ( .A(n25947), .B(n25946), .Z(n25942) );
  ANDN U26084 ( .B(B[203]), .A(n72), .Z(n25726) );
  XNOR U26085 ( .A(n25734), .B(n25948), .Z(n25727) );
  XNOR U26086 ( .A(n25733), .B(n25731), .Z(n25948) );
  AND U26087 ( .A(n25949), .B(n25950), .Z(n25731) );
  NANDN U26088 ( .A(n25951), .B(n25952), .Z(n25950) );
  OR U26089 ( .A(n25953), .B(n25954), .Z(n25952) );
  NAND U26090 ( .A(n25954), .B(n25953), .Z(n25949) );
  ANDN U26091 ( .B(B[204]), .A(n73), .Z(n25733) );
  XNOR U26092 ( .A(n25741), .B(n25955), .Z(n25734) );
  XNOR U26093 ( .A(n25740), .B(n25738), .Z(n25955) );
  AND U26094 ( .A(n25956), .B(n25957), .Z(n25738) );
  NANDN U26095 ( .A(n25958), .B(n25959), .Z(n25957) );
  NANDN U26096 ( .A(n25960), .B(n25961), .Z(n25959) );
  NANDN U26097 ( .A(n25961), .B(n25960), .Z(n25956) );
  ANDN U26098 ( .B(B[205]), .A(n74), .Z(n25740) );
  XNOR U26099 ( .A(n25748), .B(n25962), .Z(n25741) );
  XNOR U26100 ( .A(n25747), .B(n25745), .Z(n25962) );
  AND U26101 ( .A(n25963), .B(n25964), .Z(n25745) );
  NANDN U26102 ( .A(n25965), .B(n25966), .Z(n25964) );
  OR U26103 ( .A(n25967), .B(n25968), .Z(n25966) );
  NAND U26104 ( .A(n25968), .B(n25967), .Z(n25963) );
  ANDN U26105 ( .B(B[206]), .A(n75), .Z(n25747) );
  XNOR U26106 ( .A(n25755), .B(n25969), .Z(n25748) );
  XNOR U26107 ( .A(n25754), .B(n25752), .Z(n25969) );
  AND U26108 ( .A(n25970), .B(n25971), .Z(n25752) );
  NANDN U26109 ( .A(n25972), .B(n25973), .Z(n25971) );
  NANDN U26110 ( .A(n25974), .B(n25975), .Z(n25973) );
  NANDN U26111 ( .A(n25975), .B(n25974), .Z(n25970) );
  ANDN U26112 ( .B(B[207]), .A(n76), .Z(n25754) );
  XNOR U26113 ( .A(n25762), .B(n25976), .Z(n25755) );
  XNOR U26114 ( .A(n25761), .B(n25759), .Z(n25976) );
  AND U26115 ( .A(n25977), .B(n25978), .Z(n25759) );
  NANDN U26116 ( .A(n25979), .B(n25980), .Z(n25978) );
  OR U26117 ( .A(n25981), .B(n25982), .Z(n25980) );
  NAND U26118 ( .A(n25982), .B(n25981), .Z(n25977) );
  ANDN U26119 ( .B(B[208]), .A(n77), .Z(n25761) );
  XNOR U26120 ( .A(n25769), .B(n25983), .Z(n25762) );
  XNOR U26121 ( .A(n25768), .B(n25766), .Z(n25983) );
  AND U26122 ( .A(n25984), .B(n25985), .Z(n25766) );
  NANDN U26123 ( .A(n25986), .B(n25987), .Z(n25985) );
  NANDN U26124 ( .A(n25988), .B(n25989), .Z(n25987) );
  NANDN U26125 ( .A(n25989), .B(n25988), .Z(n25984) );
  ANDN U26126 ( .B(B[209]), .A(n78), .Z(n25768) );
  XNOR U26127 ( .A(n25776), .B(n25990), .Z(n25769) );
  XNOR U26128 ( .A(n25775), .B(n25773), .Z(n25990) );
  AND U26129 ( .A(n25991), .B(n25992), .Z(n25773) );
  NANDN U26130 ( .A(n25993), .B(n25994), .Z(n25992) );
  OR U26131 ( .A(n25995), .B(n25996), .Z(n25994) );
  NAND U26132 ( .A(n25996), .B(n25995), .Z(n25991) );
  ANDN U26133 ( .B(B[210]), .A(n79), .Z(n25775) );
  XNOR U26134 ( .A(n25783), .B(n25997), .Z(n25776) );
  XNOR U26135 ( .A(n25782), .B(n25780), .Z(n25997) );
  AND U26136 ( .A(n25998), .B(n25999), .Z(n25780) );
  NANDN U26137 ( .A(n26000), .B(n26001), .Z(n25999) );
  NANDN U26138 ( .A(n26002), .B(n26003), .Z(n26001) );
  NANDN U26139 ( .A(n26003), .B(n26002), .Z(n25998) );
  ANDN U26140 ( .B(B[211]), .A(n80), .Z(n25782) );
  XNOR U26141 ( .A(n25790), .B(n26004), .Z(n25783) );
  XNOR U26142 ( .A(n25789), .B(n25787), .Z(n26004) );
  AND U26143 ( .A(n26005), .B(n26006), .Z(n25787) );
  NANDN U26144 ( .A(n26007), .B(n26008), .Z(n26006) );
  OR U26145 ( .A(n26009), .B(n26010), .Z(n26008) );
  NAND U26146 ( .A(n26010), .B(n26009), .Z(n26005) );
  ANDN U26147 ( .B(B[212]), .A(n81), .Z(n25789) );
  XNOR U26148 ( .A(n25797), .B(n26011), .Z(n25790) );
  XNOR U26149 ( .A(n25796), .B(n25794), .Z(n26011) );
  AND U26150 ( .A(n26012), .B(n26013), .Z(n25794) );
  NANDN U26151 ( .A(n26014), .B(n26015), .Z(n26013) );
  NAND U26152 ( .A(n26016), .B(n26017), .Z(n26015) );
  ANDN U26153 ( .B(B[213]), .A(n82), .Z(n25796) );
  XOR U26154 ( .A(n25803), .B(n26018), .Z(n25797) );
  XNOR U26155 ( .A(n25801), .B(n25804), .Z(n26018) );
  NAND U26156 ( .A(A[2]), .B(B[214]), .Z(n25804) );
  NANDN U26157 ( .A(n26019), .B(n26020), .Z(n25801) );
  AND U26158 ( .A(A[0]), .B(B[215]), .Z(n26020) );
  XNOR U26159 ( .A(n25806), .B(n26021), .Z(n25803) );
  NAND U26160 ( .A(A[0]), .B(B[216]), .Z(n26021) );
  NAND U26161 ( .A(B[215]), .B(A[1]), .Z(n25806) );
  NAND U26162 ( .A(n26022), .B(n26023), .Z(n364) );
  NANDN U26163 ( .A(n26024), .B(n26025), .Z(n26023) );
  OR U26164 ( .A(n26026), .B(n26027), .Z(n26025) );
  NAND U26165 ( .A(n26027), .B(n26026), .Z(n26022) );
  XOR U26166 ( .A(n366), .B(n365), .Z(\A1[213] ) );
  XOR U26167 ( .A(n26027), .B(n26028), .Z(n365) );
  XNOR U26168 ( .A(n26026), .B(n26024), .Z(n26028) );
  AND U26169 ( .A(n26029), .B(n26030), .Z(n26024) );
  NANDN U26170 ( .A(n26031), .B(n26032), .Z(n26030) );
  NANDN U26171 ( .A(n26033), .B(n26034), .Z(n26032) );
  NANDN U26172 ( .A(n26034), .B(n26033), .Z(n26029) );
  ANDN U26173 ( .B(B[184]), .A(n54), .Z(n26026) );
  XNOR U26174 ( .A(n25821), .B(n26035), .Z(n26027) );
  XNOR U26175 ( .A(n25820), .B(n25818), .Z(n26035) );
  AND U26176 ( .A(n26036), .B(n26037), .Z(n25818) );
  NANDN U26177 ( .A(n26038), .B(n26039), .Z(n26037) );
  OR U26178 ( .A(n26040), .B(n26041), .Z(n26039) );
  NAND U26179 ( .A(n26041), .B(n26040), .Z(n26036) );
  ANDN U26180 ( .B(B[185]), .A(n55), .Z(n25820) );
  XNOR U26181 ( .A(n25828), .B(n26042), .Z(n25821) );
  XNOR U26182 ( .A(n25827), .B(n25825), .Z(n26042) );
  AND U26183 ( .A(n26043), .B(n26044), .Z(n25825) );
  NANDN U26184 ( .A(n26045), .B(n26046), .Z(n26044) );
  NANDN U26185 ( .A(n26047), .B(n26048), .Z(n26046) );
  NANDN U26186 ( .A(n26048), .B(n26047), .Z(n26043) );
  ANDN U26187 ( .B(B[186]), .A(n56), .Z(n25827) );
  XNOR U26188 ( .A(n25835), .B(n26049), .Z(n25828) );
  XNOR U26189 ( .A(n25834), .B(n25832), .Z(n26049) );
  AND U26190 ( .A(n26050), .B(n26051), .Z(n25832) );
  NANDN U26191 ( .A(n26052), .B(n26053), .Z(n26051) );
  OR U26192 ( .A(n26054), .B(n26055), .Z(n26053) );
  NAND U26193 ( .A(n26055), .B(n26054), .Z(n26050) );
  ANDN U26194 ( .B(B[187]), .A(n57), .Z(n25834) );
  XNOR U26195 ( .A(n25842), .B(n26056), .Z(n25835) );
  XNOR U26196 ( .A(n25841), .B(n25839), .Z(n26056) );
  AND U26197 ( .A(n26057), .B(n26058), .Z(n25839) );
  NANDN U26198 ( .A(n26059), .B(n26060), .Z(n26058) );
  NANDN U26199 ( .A(n26061), .B(n26062), .Z(n26060) );
  NANDN U26200 ( .A(n26062), .B(n26061), .Z(n26057) );
  ANDN U26201 ( .B(B[188]), .A(n58), .Z(n25841) );
  XNOR U26202 ( .A(n25849), .B(n26063), .Z(n25842) );
  XNOR U26203 ( .A(n25848), .B(n25846), .Z(n26063) );
  AND U26204 ( .A(n26064), .B(n26065), .Z(n25846) );
  NANDN U26205 ( .A(n26066), .B(n26067), .Z(n26065) );
  OR U26206 ( .A(n26068), .B(n26069), .Z(n26067) );
  NAND U26207 ( .A(n26069), .B(n26068), .Z(n26064) );
  ANDN U26208 ( .B(B[189]), .A(n59), .Z(n25848) );
  XNOR U26209 ( .A(n25856), .B(n26070), .Z(n25849) );
  XNOR U26210 ( .A(n25855), .B(n25853), .Z(n26070) );
  AND U26211 ( .A(n26071), .B(n26072), .Z(n25853) );
  NANDN U26212 ( .A(n26073), .B(n26074), .Z(n26072) );
  NANDN U26213 ( .A(n26075), .B(n26076), .Z(n26074) );
  NANDN U26214 ( .A(n26076), .B(n26075), .Z(n26071) );
  ANDN U26215 ( .B(B[190]), .A(n60), .Z(n25855) );
  XNOR U26216 ( .A(n25863), .B(n26077), .Z(n25856) );
  XNOR U26217 ( .A(n25862), .B(n25860), .Z(n26077) );
  AND U26218 ( .A(n26078), .B(n26079), .Z(n25860) );
  NANDN U26219 ( .A(n26080), .B(n26081), .Z(n26079) );
  OR U26220 ( .A(n26082), .B(n26083), .Z(n26081) );
  NAND U26221 ( .A(n26083), .B(n26082), .Z(n26078) );
  ANDN U26222 ( .B(B[191]), .A(n61), .Z(n25862) );
  XNOR U26223 ( .A(n25870), .B(n26084), .Z(n25863) );
  XNOR U26224 ( .A(n25869), .B(n25867), .Z(n26084) );
  AND U26225 ( .A(n26085), .B(n26086), .Z(n25867) );
  NANDN U26226 ( .A(n26087), .B(n26088), .Z(n26086) );
  NANDN U26227 ( .A(n26089), .B(n26090), .Z(n26088) );
  NANDN U26228 ( .A(n26090), .B(n26089), .Z(n26085) );
  ANDN U26229 ( .B(B[192]), .A(n62), .Z(n25869) );
  XNOR U26230 ( .A(n25877), .B(n26091), .Z(n25870) );
  XNOR U26231 ( .A(n25876), .B(n25874), .Z(n26091) );
  AND U26232 ( .A(n26092), .B(n26093), .Z(n25874) );
  NANDN U26233 ( .A(n26094), .B(n26095), .Z(n26093) );
  OR U26234 ( .A(n26096), .B(n26097), .Z(n26095) );
  NAND U26235 ( .A(n26097), .B(n26096), .Z(n26092) );
  ANDN U26236 ( .B(B[193]), .A(n63), .Z(n25876) );
  XNOR U26237 ( .A(n25884), .B(n26098), .Z(n25877) );
  XNOR U26238 ( .A(n25883), .B(n25881), .Z(n26098) );
  AND U26239 ( .A(n26099), .B(n26100), .Z(n25881) );
  NANDN U26240 ( .A(n26101), .B(n26102), .Z(n26100) );
  NANDN U26241 ( .A(n26103), .B(n26104), .Z(n26102) );
  NANDN U26242 ( .A(n26104), .B(n26103), .Z(n26099) );
  ANDN U26243 ( .B(B[194]), .A(n64), .Z(n25883) );
  XNOR U26244 ( .A(n25891), .B(n26105), .Z(n25884) );
  XNOR U26245 ( .A(n25890), .B(n25888), .Z(n26105) );
  AND U26246 ( .A(n26106), .B(n26107), .Z(n25888) );
  NANDN U26247 ( .A(n26108), .B(n26109), .Z(n26107) );
  OR U26248 ( .A(n26110), .B(n26111), .Z(n26109) );
  NAND U26249 ( .A(n26111), .B(n26110), .Z(n26106) );
  ANDN U26250 ( .B(B[195]), .A(n65), .Z(n25890) );
  XNOR U26251 ( .A(n25898), .B(n26112), .Z(n25891) );
  XNOR U26252 ( .A(n25897), .B(n25895), .Z(n26112) );
  AND U26253 ( .A(n26113), .B(n26114), .Z(n25895) );
  NANDN U26254 ( .A(n26115), .B(n26116), .Z(n26114) );
  NANDN U26255 ( .A(n26117), .B(n26118), .Z(n26116) );
  NANDN U26256 ( .A(n26118), .B(n26117), .Z(n26113) );
  ANDN U26257 ( .B(B[196]), .A(n66), .Z(n25897) );
  XNOR U26258 ( .A(n25905), .B(n26119), .Z(n25898) );
  XNOR U26259 ( .A(n25904), .B(n25902), .Z(n26119) );
  AND U26260 ( .A(n26120), .B(n26121), .Z(n25902) );
  NANDN U26261 ( .A(n26122), .B(n26123), .Z(n26121) );
  OR U26262 ( .A(n26124), .B(n26125), .Z(n26123) );
  NAND U26263 ( .A(n26125), .B(n26124), .Z(n26120) );
  ANDN U26264 ( .B(B[197]), .A(n67), .Z(n25904) );
  XNOR U26265 ( .A(n25912), .B(n26126), .Z(n25905) );
  XNOR U26266 ( .A(n25911), .B(n25909), .Z(n26126) );
  AND U26267 ( .A(n26127), .B(n26128), .Z(n25909) );
  NANDN U26268 ( .A(n26129), .B(n26130), .Z(n26128) );
  NANDN U26269 ( .A(n26131), .B(n26132), .Z(n26130) );
  NANDN U26270 ( .A(n26132), .B(n26131), .Z(n26127) );
  ANDN U26271 ( .B(B[198]), .A(n68), .Z(n25911) );
  XNOR U26272 ( .A(n25919), .B(n26133), .Z(n25912) );
  XNOR U26273 ( .A(n25918), .B(n25916), .Z(n26133) );
  AND U26274 ( .A(n26134), .B(n26135), .Z(n25916) );
  NANDN U26275 ( .A(n26136), .B(n26137), .Z(n26135) );
  OR U26276 ( .A(n26138), .B(n26139), .Z(n26137) );
  NAND U26277 ( .A(n26139), .B(n26138), .Z(n26134) );
  ANDN U26278 ( .B(B[199]), .A(n69), .Z(n25918) );
  XNOR U26279 ( .A(n25926), .B(n26140), .Z(n25919) );
  XNOR U26280 ( .A(n25925), .B(n25923), .Z(n26140) );
  AND U26281 ( .A(n26141), .B(n26142), .Z(n25923) );
  NANDN U26282 ( .A(n26143), .B(n26144), .Z(n26142) );
  NANDN U26283 ( .A(n26145), .B(n26146), .Z(n26144) );
  NANDN U26284 ( .A(n26146), .B(n26145), .Z(n26141) );
  ANDN U26285 ( .B(B[200]), .A(n70), .Z(n25925) );
  XNOR U26286 ( .A(n25933), .B(n26147), .Z(n25926) );
  XNOR U26287 ( .A(n25932), .B(n25930), .Z(n26147) );
  AND U26288 ( .A(n26148), .B(n26149), .Z(n25930) );
  NANDN U26289 ( .A(n26150), .B(n26151), .Z(n26149) );
  OR U26290 ( .A(n26152), .B(n26153), .Z(n26151) );
  NAND U26291 ( .A(n26153), .B(n26152), .Z(n26148) );
  ANDN U26292 ( .B(B[201]), .A(n71), .Z(n25932) );
  XNOR U26293 ( .A(n25940), .B(n26154), .Z(n25933) );
  XNOR U26294 ( .A(n25939), .B(n25937), .Z(n26154) );
  AND U26295 ( .A(n26155), .B(n26156), .Z(n25937) );
  NANDN U26296 ( .A(n26157), .B(n26158), .Z(n26156) );
  NANDN U26297 ( .A(n26159), .B(n26160), .Z(n26158) );
  NANDN U26298 ( .A(n26160), .B(n26159), .Z(n26155) );
  ANDN U26299 ( .B(B[202]), .A(n72), .Z(n25939) );
  XNOR U26300 ( .A(n25947), .B(n26161), .Z(n25940) );
  XNOR U26301 ( .A(n25946), .B(n25944), .Z(n26161) );
  AND U26302 ( .A(n26162), .B(n26163), .Z(n25944) );
  NANDN U26303 ( .A(n26164), .B(n26165), .Z(n26163) );
  OR U26304 ( .A(n26166), .B(n26167), .Z(n26165) );
  NAND U26305 ( .A(n26167), .B(n26166), .Z(n26162) );
  ANDN U26306 ( .B(B[203]), .A(n73), .Z(n25946) );
  XNOR U26307 ( .A(n25954), .B(n26168), .Z(n25947) );
  XNOR U26308 ( .A(n25953), .B(n25951), .Z(n26168) );
  AND U26309 ( .A(n26169), .B(n26170), .Z(n25951) );
  NANDN U26310 ( .A(n26171), .B(n26172), .Z(n26170) );
  NANDN U26311 ( .A(n26173), .B(n26174), .Z(n26172) );
  NANDN U26312 ( .A(n26174), .B(n26173), .Z(n26169) );
  ANDN U26313 ( .B(B[204]), .A(n74), .Z(n25953) );
  XNOR U26314 ( .A(n25961), .B(n26175), .Z(n25954) );
  XNOR U26315 ( .A(n25960), .B(n25958), .Z(n26175) );
  AND U26316 ( .A(n26176), .B(n26177), .Z(n25958) );
  NANDN U26317 ( .A(n26178), .B(n26179), .Z(n26177) );
  OR U26318 ( .A(n26180), .B(n26181), .Z(n26179) );
  NAND U26319 ( .A(n26181), .B(n26180), .Z(n26176) );
  ANDN U26320 ( .B(B[205]), .A(n75), .Z(n25960) );
  XNOR U26321 ( .A(n25968), .B(n26182), .Z(n25961) );
  XNOR U26322 ( .A(n25967), .B(n25965), .Z(n26182) );
  AND U26323 ( .A(n26183), .B(n26184), .Z(n25965) );
  NANDN U26324 ( .A(n26185), .B(n26186), .Z(n26184) );
  NANDN U26325 ( .A(n26187), .B(n26188), .Z(n26186) );
  NANDN U26326 ( .A(n26188), .B(n26187), .Z(n26183) );
  ANDN U26327 ( .B(B[206]), .A(n76), .Z(n25967) );
  XNOR U26328 ( .A(n25975), .B(n26189), .Z(n25968) );
  XNOR U26329 ( .A(n25974), .B(n25972), .Z(n26189) );
  AND U26330 ( .A(n26190), .B(n26191), .Z(n25972) );
  NANDN U26331 ( .A(n26192), .B(n26193), .Z(n26191) );
  OR U26332 ( .A(n26194), .B(n26195), .Z(n26193) );
  NAND U26333 ( .A(n26195), .B(n26194), .Z(n26190) );
  ANDN U26334 ( .B(B[207]), .A(n77), .Z(n25974) );
  XNOR U26335 ( .A(n25982), .B(n26196), .Z(n25975) );
  XNOR U26336 ( .A(n25981), .B(n25979), .Z(n26196) );
  AND U26337 ( .A(n26197), .B(n26198), .Z(n25979) );
  NANDN U26338 ( .A(n26199), .B(n26200), .Z(n26198) );
  NANDN U26339 ( .A(n26201), .B(n26202), .Z(n26200) );
  NANDN U26340 ( .A(n26202), .B(n26201), .Z(n26197) );
  ANDN U26341 ( .B(B[208]), .A(n78), .Z(n25981) );
  XNOR U26342 ( .A(n25989), .B(n26203), .Z(n25982) );
  XNOR U26343 ( .A(n25988), .B(n25986), .Z(n26203) );
  AND U26344 ( .A(n26204), .B(n26205), .Z(n25986) );
  NANDN U26345 ( .A(n26206), .B(n26207), .Z(n26205) );
  OR U26346 ( .A(n26208), .B(n26209), .Z(n26207) );
  NAND U26347 ( .A(n26209), .B(n26208), .Z(n26204) );
  ANDN U26348 ( .B(B[209]), .A(n79), .Z(n25988) );
  XNOR U26349 ( .A(n25996), .B(n26210), .Z(n25989) );
  XNOR U26350 ( .A(n25995), .B(n25993), .Z(n26210) );
  AND U26351 ( .A(n26211), .B(n26212), .Z(n25993) );
  NANDN U26352 ( .A(n26213), .B(n26214), .Z(n26212) );
  NANDN U26353 ( .A(n26215), .B(n26216), .Z(n26214) );
  NANDN U26354 ( .A(n26216), .B(n26215), .Z(n26211) );
  ANDN U26355 ( .B(B[210]), .A(n80), .Z(n25995) );
  XNOR U26356 ( .A(n26003), .B(n26217), .Z(n25996) );
  XNOR U26357 ( .A(n26002), .B(n26000), .Z(n26217) );
  AND U26358 ( .A(n26218), .B(n26219), .Z(n26000) );
  NANDN U26359 ( .A(n26220), .B(n26221), .Z(n26219) );
  OR U26360 ( .A(n26222), .B(n26223), .Z(n26221) );
  NAND U26361 ( .A(n26223), .B(n26222), .Z(n26218) );
  ANDN U26362 ( .B(B[211]), .A(n81), .Z(n26002) );
  XNOR U26363 ( .A(n26010), .B(n26224), .Z(n26003) );
  XNOR U26364 ( .A(n26009), .B(n26007), .Z(n26224) );
  AND U26365 ( .A(n26225), .B(n26226), .Z(n26007) );
  NANDN U26366 ( .A(n26227), .B(n26228), .Z(n26226) );
  NAND U26367 ( .A(n26229), .B(n26230), .Z(n26228) );
  ANDN U26368 ( .B(B[212]), .A(n82), .Z(n26009) );
  XOR U26369 ( .A(n26016), .B(n26231), .Z(n26010) );
  XNOR U26370 ( .A(n26014), .B(n26017), .Z(n26231) );
  NAND U26371 ( .A(A[2]), .B(B[213]), .Z(n26017) );
  NANDN U26372 ( .A(n26232), .B(n26233), .Z(n26014) );
  AND U26373 ( .A(A[0]), .B(B[214]), .Z(n26233) );
  XNOR U26374 ( .A(n26019), .B(n26234), .Z(n26016) );
  NAND U26375 ( .A(A[0]), .B(B[215]), .Z(n26234) );
  NAND U26376 ( .A(B[214]), .B(A[1]), .Z(n26019) );
  NAND U26377 ( .A(n26235), .B(n26236), .Z(n366) );
  NANDN U26378 ( .A(n26237), .B(n26238), .Z(n26236) );
  OR U26379 ( .A(n26239), .B(n26240), .Z(n26238) );
  NAND U26380 ( .A(n26240), .B(n26239), .Z(n26235) );
  XOR U26381 ( .A(n368), .B(n367), .Z(\A1[212] ) );
  XOR U26382 ( .A(n26240), .B(n26241), .Z(n367) );
  XNOR U26383 ( .A(n26239), .B(n26237), .Z(n26241) );
  AND U26384 ( .A(n26242), .B(n26243), .Z(n26237) );
  NANDN U26385 ( .A(n26244), .B(n26245), .Z(n26243) );
  NANDN U26386 ( .A(n26246), .B(n26247), .Z(n26245) );
  NANDN U26387 ( .A(n26247), .B(n26246), .Z(n26242) );
  ANDN U26388 ( .B(B[183]), .A(n54), .Z(n26239) );
  XNOR U26389 ( .A(n26034), .B(n26248), .Z(n26240) );
  XNOR U26390 ( .A(n26033), .B(n26031), .Z(n26248) );
  AND U26391 ( .A(n26249), .B(n26250), .Z(n26031) );
  NANDN U26392 ( .A(n26251), .B(n26252), .Z(n26250) );
  OR U26393 ( .A(n26253), .B(n26254), .Z(n26252) );
  NAND U26394 ( .A(n26254), .B(n26253), .Z(n26249) );
  ANDN U26395 ( .B(B[184]), .A(n55), .Z(n26033) );
  XNOR U26396 ( .A(n26041), .B(n26255), .Z(n26034) );
  XNOR U26397 ( .A(n26040), .B(n26038), .Z(n26255) );
  AND U26398 ( .A(n26256), .B(n26257), .Z(n26038) );
  NANDN U26399 ( .A(n26258), .B(n26259), .Z(n26257) );
  NANDN U26400 ( .A(n26260), .B(n26261), .Z(n26259) );
  NANDN U26401 ( .A(n26261), .B(n26260), .Z(n26256) );
  ANDN U26402 ( .B(B[185]), .A(n56), .Z(n26040) );
  XNOR U26403 ( .A(n26048), .B(n26262), .Z(n26041) );
  XNOR U26404 ( .A(n26047), .B(n26045), .Z(n26262) );
  AND U26405 ( .A(n26263), .B(n26264), .Z(n26045) );
  NANDN U26406 ( .A(n26265), .B(n26266), .Z(n26264) );
  OR U26407 ( .A(n26267), .B(n26268), .Z(n26266) );
  NAND U26408 ( .A(n26268), .B(n26267), .Z(n26263) );
  ANDN U26409 ( .B(B[186]), .A(n57), .Z(n26047) );
  XNOR U26410 ( .A(n26055), .B(n26269), .Z(n26048) );
  XNOR U26411 ( .A(n26054), .B(n26052), .Z(n26269) );
  AND U26412 ( .A(n26270), .B(n26271), .Z(n26052) );
  NANDN U26413 ( .A(n26272), .B(n26273), .Z(n26271) );
  NANDN U26414 ( .A(n26274), .B(n26275), .Z(n26273) );
  NANDN U26415 ( .A(n26275), .B(n26274), .Z(n26270) );
  ANDN U26416 ( .B(B[187]), .A(n58), .Z(n26054) );
  XNOR U26417 ( .A(n26062), .B(n26276), .Z(n26055) );
  XNOR U26418 ( .A(n26061), .B(n26059), .Z(n26276) );
  AND U26419 ( .A(n26277), .B(n26278), .Z(n26059) );
  NANDN U26420 ( .A(n26279), .B(n26280), .Z(n26278) );
  OR U26421 ( .A(n26281), .B(n26282), .Z(n26280) );
  NAND U26422 ( .A(n26282), .B(n26281), .Z(n26277) );
  ANDN U26423 ( .B(B[188]), .A(n59), .Z(n26061) );
  XNOR U26424 ( .A(n26069), .B(n26283), .Z(n26062) );
  XNOR U26425 ( .A(n26068), .B(n26066), .Z(n26283) );
  AND U26426 ( .A(n26284), .B(n26285), .Z(n26066) );
  NANDN U26427 ( .A(n26286), .B(n26287), .Z(n26285) );
  NANDN U26428 ( .A(n26288), .B(n26289), .Z(n26287) );
  NANDN U26429 ( .A(n26289), .B(n26288), .Z(n26284) );
  ANDN U26430 ( .B(B[189]), .A(n60), .Z(n26068) );
  XNOR U26431 ( .A(n26076), .B(n26290), .Z(n26069) );
  XNOR U26432 ( .A(n26075), .B(n26073), .Z(n26290) );
  AND U26433 ( .A(n26291), .B(n26292), .Z(n26073) );
  NANDN U26434 ( .A(n26293), .B(n26294), .Z(n26292) );
  OR U26435 ( .A(n26295), .B(n26296), .Z(n26294) );
  NAND U26436 ( .A(n26296), .B(n26295), .Z(n26291) );
  ANDN U26437 ( .B(B[190]), .A(n61), .Z(n26075) );
  XNOR U26438 ( .A(n26083), .B(n26297), .Z(n26076) );
  XNOR U26439 ( .A(n26082), .B(n26080), .Z(n26297) );
  AND U26440 ( .A(n26298), .B(n26299), .Z(n26080) );
  NANDN U26441 ( .A(n26300), .B(n26301), .Z(n26299) );
  NANDN U26442 ( .A(n26302), .B(n26303), .Z(n26301) );
  NANDN U26443 ( .A(n26303), .B(n26302), .Z(n26298) );
  ANDN U26444 ( .B(B[191]), .A(n62), .Z(n26082) );
  XNOR U26445 ( .A(n26090), .B(n26304), .Z(n26083) );
  XNOR U26446 ( .A(n26089), .B(n26087), .Z(n26304) );
  AND U26447 ( .A(n26305), .B(n26306), .Z(n26087) );
  NANDN U26448 ( .A(n26307), .B(n26308), .Z(n26306) );
  OR U26449 ( .A(n26309), .B(n26310), .Z(n26308) );
  NAND U26450 ( .A(n26310), .B(n26309), .Z(n26305) );
  ANDN U26451 ( .B(B[192]), .A(n63), .Z(n26089) );
  XNOR U26452 ( .A(n26097), .B(n26311), .Z(n26090) );
  XNOR U26453 ( .A(n26096), .B(n26094), .Z(n26311) );
  AND U26454 ( .A(n26312), .B(n26313), .Z(n26094) );
  NANDN U26455 ( .A(n26314), .B(n26315), .Z(n26313) );
  NANDN U26456 ( .A(n26316), .B(n26317), .Z(n26315) );
  NANDN U26457 ( .A(n26317), .B(n26316), .Z(n26312) );
  ANDN U26458 ( .B(B[193]), .A(n64), .Z(n26096) );
  XNOR U26459 ( .A(n26104), .B(n26318), .Z(n26097) );
  XNOR U26460 ( .A(n26103), .B(n26101), .Z(n26318) );
  AND U26461 ( .A(n26319), .B(n26320), .Z(n26101) );
  NANDN U26462 ( .A(n26321), .B(n26322), .Z(n26320) );
  OR U26463 ( .A(n26323), .B(n26324), .Z(n26322) );
  NAND U26464 ( .A(n26324), .B(n26323), .Z(n26319) );
  ANDN U26465 ( .B(B[194]), .A(n65), .Z(n26103) );
  XNOR U26466 ( .A(n26111), .B(n26325), .Z(n26104) );
  XNOR U26467 ( .A(n26110), .B(n26108), .Z(n26325) );
  AND U26468 ( .A(n26326), .B(n26327), .Z(n26108) );
  NANDN U26469 ( .A(n26328), .B(n26329), .Z(n26327) );
  NANDN U26470 ( .A(n26330), .B(n26331), .Z(n26329) );
  NANDN U26471 ( .A(n26331), .B(n26330), .Z(n26326) );
  ANDN U26472 ( .B(B[195]), .A(n66), .Z(n26110) );
  XNOR U26473 ( .A(n26118), .B(n26332), .Z(n26111) );
  XNOR U26474 ( .A(n26117), .B(n26115), .Z(n26332) );
  AND U26475 ( .A(n26333), .B(n26334), .Z(n26115) );
  NANDN U26476 ( .A(n26335), .B(n26336), .Z(n26334) );
  OR U26477 ( .A(n26337), .B(n26338), .Z(n26336) );
  NAND U26478 ( .A(n26338), .B(n26337), .Z(n26333) );
  ANDN U26479 ( .B(B[196]), .A(n67), .Z(n26117) );
  XNOR U26480 ( .A(n26125), .B(n26339), .Z(n26118) );
  XNOR U26481 ( .A(n26124), .B(n26122), .Z(n26339) );
  AND U26482 ( .A(n26340), .B(n26341), .Z(n26122) );
  NANDN U26483 ( .A(n26342), .B(n26343), .Z(n26341) );
  NANDN U26484 ( .A(n26344), .B(n26345), .Z(n26343) );
  NANDN U26485 ( .A(n26345), .B(n26344), .Z(n26340) );
  ANDN U26486 ( .B(B[197]), .A(n68), .Z(n26124) );
  XNOR U26487 ( .A(n26132), .B(n26346), .Z(n26125) );
  XNOR U26488 ( .A(n26131), .B(n26129), .Z(n26346) );
  AND U26489 ( .A(n26347), .B(n26348), .Z(n26129) );
  NANDN U26490 ( .A(n26349), .B(n26350), .Z(n26348) );
  OR U26491 ( .A(n26351), .B(n26352), .Z(n26350) );
  NAND U26492 ( .A(n26352), .B(n26351), .Z(n26347) );
  ANDN U26493 ( .B(B[198]), .A(n69), .Z(n26131) );
  XNOR U26494 ( .A(n26139), .B(n26353), .Z(n26132) );
  XNOR U26495 ( .A(n26138), .B(n26136), .Z(n26353) );
  AND U26496 ( .A(n26354), .B(n26355), .Z(n26136) );
  NANDN U26497 ( .A(n26356), .B(n26357), .Z(n26355) );
  NANDN U26498 ( .A(n26358), .B(n26359), .Z(n26357) );
  NANDN U26499 ( .A(n26359), .B(n26358), .Z(n26354) );
  ANDN U26500 ( .B(B[199]), .A(n70), .Z(n26138) );
  XNOR U26501 ( .A(n26146), .B(n26360), .Z(n26139) );
  XNOR U26502 ( .A(n26145), .B(n26143), .Z(n26360) );
  AND U26503 ( .A(n26361), .B(n26362), .Z(n26143) );
  NANDN U26504 ( .A(n26363), .B(n26364), .Z(n26362) );
  OR U26505 ( .A(n26365), .B(n26366), .Z(n26364) );
  NAND U26506 ( .A(n26366), .B(n26365), .Z(n26361) );
  ANDN U26507 ( .B(B[200]), .A(n71), .Z(n26145) );
  XNOR U26508 ( .A(n26153), .B(n26367), .Z(n26146) );
  XNOR U26509 ( .A(n26152), .B(n26150), .Z(n26367) );
  AND U26510 ( .A(n26368), .B(n26369), .Z(n26150) );
  NANDN U26511 ( .A(n26370), .B(n26371), .Z(n26369) );
  NANDN U26512 ( .A(n26372), .B(n26373), .Z(n26371) );
  NANDN U26513 ( .A(n26373), .B(n26372), .Z(n26368) );
  ANDN U26514 ( .B(B[201]), .A(n72), .Z(n26152) );
  XNOR U26515 ( .A(n26160), .B(n26374), .Z(n26153) );
  XNOR U26516 ( .A(n26159), .B(n26157), .Z(n26374) );
  AND U26517 ( .A(n26375), .B(n26376), .Z(n26157) );
  NANDN U26518 ( .A(n26377), .B(n26378), .Z(n26376) );
  OR U26519 ( .A(n26379), .B(n26380), .Z(n26378) );
  NAND U26520 ( .A(n26380), .B(n26379), .Z(n26375) );
  ANDN U26521 ( .B(B[202]), .A(n73), .Z(n26159) );
  XNOR U26522 ( .A(n26167), .B(n26381), .Z(n26160) );
  XNOR U26523 ( .A(n26166), .B(n26164), .Z(n26381) );
  AND U26524 ( .A(n26382), .B(n26383), .Z(n26164) );
  NANDN U26525 ( .A(n26384), .B(n26385), .Z(n26383) );
  NANDN U26526 ( .A(n26386), .B(n26387), .Z(n26385) );
  NANDN U26527 ( .A(n26387), .B(n26386), .Z(n26382) );
  ANDN U26528 ( .B(B[203]), .A(n74), .Z(n26166) );
  XNOR U26529 ( .A(n26174), .B(n26388), .Z(n26167) );
  XNOR U26530 ( .A(n26173), .B(n26171), .Z(n26388) );
  AND U26531 ( .A(n26389), .B(n26390), .Z(n26171) );
  NANDN U26532 ( .A(n26391), .B(n26392), .Z(n26390) );
  OR U26533 ( .A(n26393), .B(n26394), .Z(n26392) );
  NAND U26534 ( .A(n26394), .B(n26393), .Z(n26389) );
  ANDN U26535 ( .B(B[204]), .A(n75), .Z(n26173) );
  XNOR U26536 ( .A(n26181), .B(n26395), .Z(n26174) );
  XNOR U26537 ( .A(n26180), .B(n26178), .Z(n26395) );
  AND U26538 ( .A(n26396), .B(n26397), .Z(n26178) );
  NANDN U26539 ( .A(n26398), .B(n26399), .Z(n26397) );
  NANDN U26540 ( .A(n26400), .B(n26401), .Z(n26399) );
  NANDN U26541 ( .A(n26401), .B(n26400), .Z(n26396) );
  ANDN U26542 ( .B(B[205]), .A(n76), .Z(n26180) );
  XNOR U26543 ( .A(n26188), .B(n26402), .Z(n26181) );
  XNOR U26544 ( .A(n26187), .B(n26185), .Z(n26402) );
  AND U26545 ( .A(n26403), .B(n26404), .Z(n26185) );
  NANDN U26546 ( .A(n26405), .B(n26406), .Z(n26404) );
  OR U26547 ( .A(n26407), .B(n26408), .Z(n26406) );
  NAND U26548 ( .A(n26408), .B(n26407), .Z(n26403) );
  ANDN U26549 ( .B(B[206]), .A(n77), .Z(n26187) );
  XNOR U26550 ( .A(n26195), .B(n26409), .Z(n26188) );
  XNOR U26551 ( .A(n26194), .B(n26192), .Z(n26409) );
  AND U26552 ( .A(n26410), .B(n26411), .Z(n26192) );
  NANDN U26553 ( .A(n26412), .B(n26413), .Z(n26411) );
  NANDN U26554 ( .A(n26414), .B(n26415), .Z(n26413) );
  NANDN U26555 ( .A(n26415), .B(n26414), .Z(n26410) );
  ANDN U26556 ( .B(B[207]), .A(n78), .Z(n26194) );
  XNOR U26557 ( .A(n26202), .B(n26416), .Z(n26195) );
  XNOR U26558 ( .A(n26201), .B(n26199), .Z(n26416) );
  AND U26559 ( .A(n26417), .B(n26418), .Z(n26199) );
  NANDN U26560 ( .A(n26419), .B(n26420), .Z(n26418) );
  OR U26561 ( .A(n26421), .B(n26422), .Z(n26420) );
  NAND U26562 ( .A(n26422), .B(n26421), .Z(n26417) );
  ANDN U26563 ( .B(B[208]), .A(n79), .Z(n26201) );
  XNOR U26564 ( .A(n26209), .B(n26423), .Z(n26202) );
  XNOR U26565 ( .A(n26208), .B(n26206), .Z(n26423) );
  AND U26566 ( .A(n26424), .B(n26425), .Z(n26206) );
  NANDN U26567 ( .A(n26426), .B(n26427), .Z(n26425) );
  NANDN U26568 ( .A(n26428), .B(n26429), .Z(n26427) );
  NANDN U26569 ( .A(n26429), .B(n26428), .Z(n26424) );
  ANDN U26570 ( .B(B[209]), .A(n80), .Z(n26208) );
  XNOR U26571 ( .A(n26216), .B(n26430), .Z(n26209) );
  XNOR U26572 ( .A(n26215), .B(n26213), .Z(n26430) );
  AND U26573 ( .A(n26431), .B(n26432), .Z(n26213) );
  NANDN U26574 ( .A(n26433), .B(n26434), .Z(n26432) );
  OR U26575 ( .A(n26435), .B(n26436), .Z(n26434) );
  NAND U26576 ( .A(n26436), .B(n26435), .Z(n26431) );
  ANDN U26577 ( .B(B[210]), .A(n81), .Z(n26215) );
  XNOR U26578 ( .A(n26223), .B(n26437), .Z(n26216) );
  XNOR U26579 ( .A(n26222), .B(n26220), .Z(n26437) );
  AND U26580 ( .A(n26438), .B(n26439), .Z(n26220) );
  NANDN U26581 ( .A(n26440), .B(n26441), .Z(n26439) );
  NAND U26582 ( .A(n26442), .B(n26443), .Z(n26441) );
  ANDN U26583 ( .B(B[211]), .A(n82), .Z(n26222) );
  XOR U26584 ( .A(n26229), .B(n26444), .Z(n26223) );
  XNOR U26585 ( .A(n26227), .B(n26230), .Z(n26444) );
  NAND U26586 ( .A(A[2]), .B(B[212]), .Z(n26230) );
  NANDN U26587 ( .A(n26445), .B(n26446), .Z(n26227) );
  AND U26588 ( .A(A[0]), .B(B[213]), .Z(n26446) );
  XNOR U26589 ( .A(n26232), .B(n26447), .Z(n26229) );
  NAND U26590 ( .A(A[0]), .B(B[214]), .Z(n26447) );
  NAND U26591 ( .A(B[213]), .B(A[1]), .Z(n26232) );
  NAND U26592 ( .A(n26448), .B(n26449), .Z(n368) );
  NANDN U26593 ( .A(n26450), .B(n26451), .Z(n26449) );
  OR U26594 ( .A(n26452), .B(n26453), .Z(n26451) );
  NAND U26595 ( .A(n26453), .B(n26452), .Z(n26448) );
  XOR U26596 ( .A(n370), .B(n369), .Z(\A1[211] ) );
  XOR U26597 ( .A(n26453), .B(n26454), .Z(n369) );
  XNOR U26598 ( .A(n26452), .B(n26450), .Z(n26454) );
  AND U26599 ( .A(n26455), .B(n26456), .Z(n26450) );
  NANDN U26600 ( .A(n26457), .B(n26458), .Z(n26456) );
  NANDN U26601 ( .A(n26459), .B(n26460), .Z(n26458) );
  NANDN U26602 ( .A(n26460), .B(n26459), .Z(n26455) );
  ANDN U26603 ( .B(B[182]), .A(n54), .Z(n26452) );
  XNOR U26604 ( .A(n26247), .B(n26461), .Z(n26453) );
  XNOR U26605 ( .A(n26246), .B(n26244), .Z(n26461) );
  AND U26606 ( .A(n26462), .B(n26463), .Z(n26244) );
  NANDN U26607 ( .A(n26464), .B(n26465), .Z(n26463) );
  OR U26608 ( .A(n26466), .B(n26467), .Z(n26465) );
  NAND U26609 ( .A(n26467), .B(n26466), .Z(n26462) );
  ANDN U26610 ( .B(B[183]), .A(n55), .Z(n26246) );
  XNOR U26611 ( .A(n26254), .B(n26468), .Z(n26247) );
  XNOR U26612 ( .A(n26253), .B(n26251), .Z(n26468) );
  AND U26613 ( .A(n26469), .B(n26470), .Z(n26251) );
  NANDN U26614 ( .A(n26471), .B(n26472), .Z(n26470) );
  NANDN U26615 ( .A(n26473), .B(n26474), .Z(n26472) );
  NANDN U26616 ( .A(n26474), .B(n26473), .Z(n26469) );
  ANDN U26617 ( .B(B[184]), .A(n56), .Z(n26253) );
  XNOR U26618 ( .A(n26261), .B(n26475), .Z(n26254) );
  XNOR U26619 ( .A(n26260), .B(n26258), .Z(n26475) );
  AND U26620 ( .A(n26476), .B(n26477), .Z(n26258) );
  NANDN U26621 ( .A(n26478), .B(n26479), .Z(n26477) );
  OR U26622 ( .A(n26480), .B(n26481), .Z(n26479) );
  NAND U26623 ( .A(n26481), .B(n26480), .Z(n26476) );
  ANDN U26624 ( .B(B[185]), .A(n57), .Z(n26260) );
  XNOR U26625 ( .A(n26268), .B(n26482), .Z(n26261) );
  XNOR U26626 ( .A(n26267), .B(n26265), .Z(n26482) );
  AND U26627 ( .A(n26483), .B(n26484), .Z(n26265) );
  NANDN U26628 ( .A(n26485), .B(n26486), .Z(n26484) );
  NANDN U26629 ( .A(n26487), .B(n26488), .Z(n26486) );
  NANDN U26630 ( .A(n26488), .B(n26487), .Z(n26483) );
  ANDN U26631 ( .B(B[186]), .A(n58), .Z(n26267) );
  XNOR U26632 ( .A(n26275), .B(n26489), .Z(n26268) );
  XNOR U26633 ( .A(n26274), .B(n26272), .Z(n26489) );
  AND U26634 ( .A(n26490), .B(n26491), .Z(n26272) );
  NANDN U26635 ( .A(n26492), .B(n26493), .Z(n26491) );
  OR U26636 ( .A(n26494), .B(n26495), .Z(n26493) );
  NAND U26637 ( .A(n26495), .B(n26494), .Z(n26490) );
  ANDN U26638 ( .B(B[187]), .A(n59), .Z(n26274) );
  XNOR U26639 ( .A(n26282), .B(n26496), .Z(n26275) );
  XNOR U26640 ( .A(n26281), .B(n26279), .Z(n26496) );
  AND U26641 ( .A(n26497), .B(n26498), .Z(n26279) );
  NANDN U26642 ( .A(n26499), .B(n26500), .Z(n26498) );
  NANDN U26643 ( .A(n26501), .B(n26502), .Z(n26500) );
  NANDN U26644 ( .A(n26502), .B(n26501), .Z(n26497) );
  ANDN U26645 ( .B(B[188]), .A(n60), .Z(n26281) );
  XNOR U26646 ( .A(n26289), .B(n26503), .Z(n26282) );
  XNOR U26647 ( .A(n26288), .B(n26286), .Z(n26503) );
  AND U26648 ( .A(n26504), .B(n26505), .Z(n26286) );
  NANDN U26649 ( .A(n26506), .B(n26507), .Z(n26505) );
  OR U26650 ( .A(n26508), .B(n26509), .Z(n26507) );
  NAND U26651 ( .A(n26509), .B(n26508), .Z(n26504) );
  ANDN U26652 ( .B(B[189]), .A(n61), .Z(n26288) );
  XNOR U26653 ( .A(n26296), .B(n26510), .Z(n26289) );
  XNOR U26654 ( .A(n26295), .B(n26293), .Z(n26510) );
  AND U26655 ( .A(n26511), .B(n26512), .Z(n26293) );
  NANDN U26656 ( .A(n26513), .B(n26514), .Z(n26512) );
  NANDN U26657 ( .A(n26515), .B(n26516), .Z(n26514) );
  NANDN U26658 ( .A(n26516), .B(n26515), .Z(n26511) );
  ANDN U26659 ( .B(B[190]), .A(n62), .Z(n26295) );
  XNOR U26660 ( .A(n26303), .B(n26517), .Z(n26296) );
  XNOR U26661 ( .A(n26302), .B(n26300), .Z(n26517) );
  AND U26662 ( .A(n26518), .B(n26519), .Z(n26300) );
  NANDN U26663 ( .A(n26520), .B(n26521), .Z(n26519) );
  OR U26664 ( .A(n26522), .B(n26523), .Z(n26521) );
  NAND U26665 ( .A(n26523), .B(n26522), .Z(n26518) );
  ANDN U26666 ( .B(B[191]), .A(n63), .Z(n26302) );
  XNOR U26667 ( .A(n26310), .B(n26524), .Z(n26303) );
  XNOR U26668 ( .A(n26309), .B(n26307), .Z(n26524) );
  AND U26669 ( .A(n26525), .B(n26526), .Z(n26307) );
  NANDN U26670 ( .A(n26527), .B(n26528), .Z(n26526) );
  NANDN U26671 ( .A(n26529), .B(n26530), .Z(n26528) );
  NANDN U26672 ( .A(n26530), .B(n26529), .Z(n26525) );
  ANDN U26673 ( .B(B[192]), .A(n64), .Z(n26309) );
  XNOR U26674 ( .A(n26317), .B(n26531), .Z(n26310) );
  XNOR U26675 ( .A(n26316), .B(n26314), .Z(n26531) );
  AND U26676 ( .A(n26532), .B(n26533), .Z(n26314) );
  NANDN U26677 ( .A(n26534), .B(n26535), .Z(n26533) );
  OR U26678 ( .A(n26536), .B(n26537), .Z(n26535) );
  NAND U26679 ( .A(n26537), .B(n26536), .Z(n26532) );
  ANDN U26680 ( .B(B[193]), .A(n65), .Z(n26316) );
  XNOR U26681 ( .A(n26324), .B(n26538), .Z(n26317) );
  XNOR U26682 ( .A(n26323), .B(n26321), .Z(n26538) );
  AND U26683 ( .A(n26539), .B(n26540), .Z(n26321) );
  NANDN U26684 ( .A(n26541), .B(n26542), .Z(n26540) );
  NANDN U26685 ( .A(n26543), .B(n26544), .Z(n26542) );
  NANDN U26686 ( .A(n26544), .B(n26543), .Z(n26539) );
  ANDN U26687 ( .B(B[194]), .A(n66), .Z(n26323) );
  XNOR U26688 ( .A(n26331), .B(n26545), .Z(n26324) );
  XNOR U26689 ( .A(n26330), .B(n26328), .Z(n26545) );
  AND U26690 ( .A(n26546), .B(n26547), .Z(n26328) );
  NANDN U26691 ( .A(n26548), .B(n26549), .Z(n26547) );
  OR U26692 ( .A(n26550), .B(n26551), .Z(n26549) );
  NAND U26693 ( .A(n26551), .B(n26550), .Z(n26546) );
  ANDN U26694 ( .B(B[195]), .A(n67), .Z(n26330) );
  XNOR U26695 ( .A(n26338), .B(n26552), .Z(n26331) );
  XNOR U26696 ( .A(n26337), .B(n26335), .Z(n26552) );
  AND U26697 ( .A(n26553), .B(n26554), .Z(n26335) );
  NANDN U26698 ( .A(n26555), .B(n26556), .Z(n26554) );
  NANDN U26699 ( .A(n26557), .B(n26558), .Z(n26556) );
  NANDN U26700 ( .A(n26558), .B(n26557), .Z(n26553) );
  ANDN U26701 ( .B(B[196]), .A(n68), .Z(n26337) );
  XNOR U26702 ( .A(n26345), .B(n26559), .Z(n26338) );
  XNOR U26703 ( .A(n26344), .B(n26342), .Z(n26559) );
  AND U26704 ( .A(n26560), .B(n26561), .Z(n26342) );
  NANDN U26705 ( .A(n26562), .B(n26563), .Z(n26561) );
  OR U26706 ( .A(n26564), .B(n26565), .Z(n26563) );
  NAND U26707 ( .A(n26565), .B(n26564), .Z(n26560) );
  ANDN U26708 ( .B(B[197]), .A(n69), .Z(n26344) );
  XNOR U26709 ( .A(n26352), .B(n26566), .Z(n26345) );
  XNOR U26710 ( .A(n26351), .B(n26349), .Z(n26566) );
  AND U26711 ( .A(n26567), .B(n26568), .Z(n26349) );
  NANDN U26712 ( .A(n26569), .B(n26570), .Z(n26568) );
  NANDN U26713 ( .A(n26571), .B(n26572), .Z(n26570) );
  NANDN U26714 ( .A(n26572), .B(n26571), .Z(n26567) );
  ANDN U26715 ( .B(B[198]), .A(n70), .Z(n26351) );
  XNOR U26716 ( .A(n26359), .B(n26573), .Z(n26352) );
  XNOR U26717 ( .A(n26358), .B(n26356), .Z(n26573) );
  AND U26718 ( .A(n26574), .B(n26575), .Z(n26356) );
  NANDN U26719 ( .A(n26576), .B(n26577), .Z(n26575) );
  OR U26720 ( .A(n26578), .B(n26579), .Z(n26577) );
  NAND U26721 ( .A(n26579), .B(n26578), .Z(n26574) );
  ANDN U26722 ( .B(B[199]), .A(n71), .Z(n26358) );
  XNOR U26723 ( .A(n26366), .B(n26580), .Z(n26359) );
  XNOR U26724 ( .A(n26365), .B(n26363), .Z(n26580) );
  AND U26725 ( .A(n26581), .B(n26582), .Z(n26363) );
  NANDN U26726 ( .A(n26583), .B(n26584), .Z(n26582) );
  NANDN U26727 ( .A(n26585), .B(n26586), .Z(n26584) );
  NANDN U26728 ( .A(n26586), .B(n26585), .Z(n26581) );
  ANDN U26729 ( .B(B[200]), .A(n72), .Z(n26365) );
  XNOR U26730 ( .A(n26373), .B(n26587), .Z(n26366) );
  XNOR U26731 ( .A(n26372), .B(n26370), .Z(n26587) );
  AND U26732 ( .A(n26588), .B(n26589), .Z(n26370) );
  NANDN U26733 ( .A(n26590), .B(n26591), .Z(n26589) );
  OR U26734 ( .A(n26592), .B(n26593), .Z(n26591) );
  NAND U26735 ( .A(n26593), .B(n26592), .Z(n26588) );
  ANDN U26736 ( .B(B[201]), .A(n73), .Z(n26372) );
  XNOR U26737 ( .A(n26380), .B(n26594), .Z(n26373) );
  XNOR U26738 ( .A(n26379), .B(n26377), .Z(n26594) );
  AND U26739 ( .A(n26595), .B(n26596), .Z(n26377) );
  NANDN U26740 ( .A(n26597), .B(n26598), .Z(n26596) );
  NANDN U26741 ( .A(n26599), .B(n26600), .Z(n26598) );
  NANDN U26742 ( .A(n26600), .B(n26599), .Z(n26595) );
  ANDN U26743 ( .B(B[202]), .A(n74), .Z(n26379) );
  XNOR U26744 ( .A(n26387), .B(n26601), .Z(n26380) );
  XNOR U26745 ( .A(n26386), .B(n26384), .Z(n26601) );
  AND U26746 ( .A(n26602), .B(n26603), .Z(n26384) );
  NANDN U26747 ( .A(n26604), .B(n26605), .Z(n26603) );
  OR U26748 ( .A(n26606), .B(n26607), .Z(n26605) );
  NAND U26749 ( .A(n26607), .B(n26606), .Z(n26602) );
  ANDN U26750 ( .B(B[203]), .A(n75), .Z(n26386) );
  XNOR U26751 ( .A(n26394), .B(n26608), .Z(n26387) );
  XNOR U26752 ( .A(n26393), .B(n26391), .Z(n26608) );
  AND U26753 ( .A(n26609), .B(n26610), .Z(n26391) );
  NANDN U26754 ( .A(n26611), .B(n26612), .Z(n26610) );
  NANDN U26755 ( .A(n26613), .B(n26614), .Z(n26612) );
  NANDN U26756 ( .A(n26614), .B(n26613), .Z(n26609) );
  ANDN U26757 ( .B(B[204]), .A(n76), .Z(n26393) );
  XNOR U26758 ( .A(n26401), .B(n26615), .Z(n26394) );
  XNOR U26759 ( .A(n26400), .B(n26398), .Z(n26615) );
  AND U26760 ( .A(n26616), .B(n26617), .Z(n26398) );
  NANDN U26761 ( .A(n26618), .B(n26619), .Z(n26617) );
  OR U26762 ( .A(n26620), .B(n26621), .Z(n26619) );
  NAND U26763 ( .A(n26621), .B(n26620), .Z(n26616) );
  ANDN U26764 ( .B(B[205]), .A(n77), .Z(n26400) );
  XNOR U26765 ( .A(n26408), .B(n26622), .Z(n26401) );
  XNOR U26766 ( .A(n26407), .B(n26405), .Z(n26622) );
  AND U26767 ( .A(n26623), .B(n26624), .Z(n26405) );
  NANDN U26768 ( .A(n26625), .B(n26626), .Z(n26624) );
  NANDN U26769 ( .A(n26627), .B(n26628), .Z(n26626) );
  NANDN U26770 ( .A(n26628), .B(n26627), .Z(n26623) );
  ANDN U26771 ( .B(B[206]), .A(n78), .Z(n26407) );
  XNOR U26772 ( .A(n26415), .B(n26629), .Z(n26408) );
  XNOR U26773 ( .A(n26414), .B(n26412), .Z(n26629) );
  AND U26774 ( .A(n26630), .B(n26631), .Z(n26412) );
  NANDN U26775 ( .A(n26632), .B(n26633), .Z(n26631) );
  OR U26776 ( .A(n26634), .B(n26635), .Z(n26633) );
  NAND U26777 ( .A(n26635), .B(n26634), .Z(n26630) );
  ANDN U26778 ( .B(B[207]), .A(n79), .Z(n26414) );
  XNOR U26779 ( .A(n26422), .B(n26636), .Z(n26415) );
  XNOR U26780 ( .A(n26421), .B(n26419), .Z(n26636) );
  AND U26781 ( .A(n26637), .B(n26638), .Z(n26419) );
  NANDN U26782 ( .A(n26639), .B(n26640), .Z(n26638) );
  NANDN U26783 ( .A(n26641), .B(n26642), .Z(n26640) );
  NANDN U26784 ( .A(n26642), .B(n26641), .Z(n26637) );
  ANDN U26785 ( .B(B[208]), .A(n80), .Z(n26421) );
  XNOR U26786 ( .A(n26429), .B(n26643), .Z(n26422) );
  XNOR U26787 ( .A(n26428), .B(n26426), .Z(n26643) );
  AND U26788 ( .A(n26644), .B(n26645), .Z(n26426) );
  NANDN U26789 ( .A(n26646), .B(n26647), .Z(n26645) );
  OR U26790 ( .A(n26648), .B(n26649), .Z(n26647) );
  NAND U26791 ( .A(n26649), .B(n26648), .Z(n26644) );
  ANDN U26792 ( .B(B[209]), .A(n81), .Z(n26428) );
  XNOR U26793 ( .A(n26436), .B(n26650), .Z(n26429) );
  XNOR U26794 ( .A(n26435), .B(n26433), .Z(n26650) );
  AND U26795 ( .A(n26651), .B(n26652), .Z(n26433) );
  NANDN U26796 ( .A(n26653), .B(n26654), .Z(n26652) );
  NAND U26797 ( .A(n26655), .B(n26656), .Z(n26654) );
  ANDN U26798 ( .B(B[210]), .A(n82), .Z(n26435) );
  XOR U26799 ( .A(n26442), .B(n26657), .Z(n26436) );
  XNOR U26800 ( .A(n26440), .B(n26443), .Z(n26657) );
  NAND U26801 ( .A(A[2]), .B(B[211]), .Z(n26443) );
  NANDN U26802 ( .A(n26658), .B(n26659), .Z(n26440) );
  AND U26803 ( .A(A[0]), .B(B[212]), .Z(n26659) );
  XNOR U26804 ( .A(n26445), .B(n26660), .Z(n26442) );
  NAND U26805 ( .A(A[0]), .B(B[213]), .Z(n26660) );
  NAND U26806 ( .A(B[212]), .B(A[1]), .Z(n26445) );
  NAND U26807 ( .A(n26661), .B(n26662), .Z(n370) );
  NANDN U26808 ( .A(n26663), .B(n26664), .Z(n26662) );
  OR U26809 ( .A(n26665), .B(n26666), .Z(n26664) );
  NAND U26810 ( .A(n26666), .B(n26665), .Z(n26661) );
  XOR U26811 ( .A(n372), .B(n371), .Z(\A1[210] ) );
  XOR U26812 ( .A(n26666), .B(n26667), .Z(n371) );
  XNOR U26813 ( .A(n26665), .B(n26663), .Z(n26667) );
  AND U26814 ( .A(n26668), .B(n26669), .Z(n26663) );
  NANDN U26815 ( .A(n26670), .B(n26671), .Z(n26669) );
  NANDN U26816 ( .A(n26672), .B(n26673), .Z(n26671) );
  NANDN U26817 ( .A(n26673), .B(n26672), .Z(n26668) );
  ANDN U26818 ( .B(B[181]), .A(n54), .Z(n26665) );
  XNOR U26819 ( .A(n26460), .B(n26674), .Z(n26666) );
  XNOR U26820 ( .A(n26459), .B(n26457), .Z(n26674) );
  AND U26821 ( .A(n26675), .B(n26676), .Z(n26457) );
  NANDN U26822 ( .A(n26677), .B(n26678), .Z(n26676) );
  OR U26823 ( .A(n26679), .B(n26680), .Z(n26678) );
  NAND U26824 ( .A(n26680), .B(n26679), .Z(n26675) );
  ANDN U26825 ( .B(B[182]), .A(n55), .Z(n26459) );
  XNOR U26826 ( .A(n26467), .B(n26681), .Z(n26460) );
  XNOR U26827 ( .A(n26466), .B(n26464), .Z(n26681) );
  AND U26828 ( .A(n26682), .B(n26683), .Z(n26464) );
  NANDN U26829 ( .A(n26684), .B(n26685), .Z(n26683) );
  NANDN U26830 ( .A(n26686), .B(n26687), .Z(n26685) );
  NANDN U26831 ( .A(n26687), .B(n26686), .Z(n26682) );
  ANDN U26832 ( .B(B[183]), .A(n56), .Z(n26466) );
  XNOR U26833 ( .A(n26474), .B(n26688), .Z(n26467) );
  XNOR U26834 ( .A(n26473), .B(n26471), .Z(n26688) );
  AND U26835 ( .A(n26689), .B(n26690), .Z(n26471) );
  NANDN U26836 ( .A(n26691), .B(n26692), .Z(n26690) );
  OR U26837 ( .A(n26693), .B(n26694), .Z(n26692) );
  NAND U26838 ( .A(n26694), .B(n26693), .Z(n26689) );
  ANDN U26839 ( .B(B[184]), .A(n57), .Z(n26473) );
  XNOR U26840 ( .A(n26481), .B(n26695), .Z(n26474) );
  XNOR U26841 ( .A(n26480), .B(n26478), .Z(n26695) );
  AND U26842 ( .A(n26696), .B(n26697), .Z(n26478) );
  NANDN U26843 ( .A(n26698), .B(n26699), .Z(n26697) );
  NANDN U26844 ( .A(n26700), .B(n26701), .Z(n26699) );
  NANDN U26845 ( .A(n26701), .B(n26700), .Z(n26696) );
  ANDN U26846 ( .B(B[185]), .A(n58), .Z(n26480) );
  XNOR U26847 ( .A(n26488), .B(n26702), .Z(n26481) );
  XNOR U26848 ( .A(n26487), .B(n26485), .Z(n26702) );
  AND U26849 ( .A(n26703), .B(n26704), .Z(n26485) );
  NANDN U26850 ( .A(n26705), .B(n26706), .Z(n26704) );
  OR U26851 ( .A(n26707), .B(n26708), .Z(n26706) );
  NAND U26852 ( .A(n26708), .B(n26707), .Z(n26703) );
  ANDN U26853 ( .B(B[186]), .A(n59), .Z(n26487) );
  XNOR U26854 ( .A(n26495), .B(n26709), .Z(n26488) );
  XNOR U26855 ( .A(n26494), .B(n26492), .Z(n26709) );
  AND U26856 ( .A(n26710), .B(n26711), .Z(n26492) );
  NANDN U26857 ( .A(n26712), .B(n26713), .Z(n26711) );
  NANDN U26858 ( .A(n26714), .B(n26715), .Z(n26713) );
  NANDN U26859 ( .A(n26715), .B(n26714), .Z(n26710) );
  ANDN U26860 ( .B(B[187]), .A(n60), .Z(n26494) );
  XNOR U26861 ( .A(n26502), .B(n26716), .Z(n26495) );
  XNOR U26862 ( .A(n26501), .B(n26499), .Z(n26716) );
  AND U26863 ( .A(n26717), .B(n26718), .Z(n26499) );
  NANDN U26864 ( .A(n26719), .B(n26720), .Z(n26718) );
  OR U26865 ( .A(n26721), .B(n26722), .Z(n26720) );
  NAND U26866 ( .A(n26722), .B(n26721), .Z(n26717) );
  ANDN U26867 ( .B(B[188]), .A(n61), .Z(n26501) );
  XNOR U26868 ( .A(n26509), .B(n26723), .Z(n26502) );
  XNOR U26869 ( .A(n26508), .B(n26506), .Z(n26723) );
  AND U26870 ( .A(n26724), .B(n26725), .Z(n26506) );
  NANDN U26871 ( .A(n26726), .B(n26727), .Z(n26725) );
  NANDN U26872 ( .A(n26728), .B(n26729), .Z(n26727) );
  NANDN U26873 ( .A(n26729), .B(n26728), .Z(n26724) );
  ANDN U26874 ( .B(B[189]), .A(n62), .Z(n26508) );
  XNOR U26875 ( .A(n26516), .B(n26730), .Z(n26509) );
  XNOR U26876 ( .A(n26515), .B(n26513), .Z(n26730) );
  AND U26877 ( .A(n26731), .B(n26732), .Z(n26513) );
  NANDN U26878 ( .A(n26733), .B(n26734), .Z(n26732) );
  OR U26879 ( .A(n26735), .B(n26736), .Z(n26734) );
  NAND U26880 ( .A(n26736), .B(n26735), .Z(n26731) );
  ANDN U26881 ( .B(B[190]), .A(n63), .Z(n26515) );
  XNOR U26882 ( .A(n26523), .B(n26737), .Z(n26516) );
  XNOR U26883 ( .A(n26522), .B(n26520), .Z(n26737) );
  AND U26884 ( .A(n26738), .B(n26739), .Z(n26520) );
  NANDN U26885 ( .A(n26740), .B(n26741), .Z(n26739) );
  NANDN U26886 ( .A(n26742), .B(n26743), .Z(n26741) );
  NANDN U26887 ( .A(n26743), .B(n26742), .Z(n26738) );
  ANDN U26888 ( .B(B[191]), .A(n64), .Z(n26522) );
  XNOR U26889 ( .A(n26530), .B(n26744), .Z(n26523) );
  XNOR U26890 ( .A(n26529), .B(n26527), .Z(n26744) );
  AND U26891 ( .A(n26745), .B(n26746), .Z(n26527) );
  NANDN U26892 ( .A(n26747), .B(n26748), .Z(n26746) );
  OR U26893 ( .A(n26749), .B(n26750), .Z(n26748) );
  NAND U26894 ( .A(n26750), .B(n26749), .Z(n26745) );
  ANDN U26895 ( .B(B[192]), .A(n65), .Z(n26529) );
  XNOR U26896 ( .A(n26537), .B(n26751), .Z(n26530) );
  XNOR U26897 ( .A(n26536), .B(n26534), .Z(n26751) );
  AND U26898 ( .A(n26752), .B(n26753), .Z(n26534) );
  NANDN U26899 ( .A(n26754), .B(n26755), .Z(n26753) );
  NANDN U26900 ( .A(n26756), .B(n26757), .Z(n26755) );
  NANDN U26901 ( .A(n26757), .B(n26756), .Z(n26752) );
  ANDN U26902 ( .B(B[193]), .A(n66), .Z(n26536) );
  XNOR U26903 ( .A(n26544), .B(n26758), .Z(n26537) );
  XNOR U26904 ( .A(n26543), .B(n26541), .Z(n26758) );
  AND U26905 ( .A(n26759), .B(n26760), .Z(n26541) );
  NANDN U26906 ( .A(n26761), .B(n26762), .Z(n26760) );
  OR U26907 ( .A(n26763), .B(n26764), .Z(n26762) );
  NAND U26908 ( .A(n26764), .B(n26763), .Z(n26759) );
  ANDN U26909 ( .B(B[194]), .A(n67), .Z(n26543) );
  XNOR U26910 ( .A(n26551), .B(n26765), .Z(n26544) );
  XNOR U26911 ( .A(n26550), .B(n26548), .Z(n26765) );
  AND U26912 ( .A(n26766), .B(n26767), .Z(n26548) );
  NANDN U26913 ( .A(n26768), .B(n26769), .Z(n26767) );
  NANDN U26914 ( .A(n26770), .B(n26771), .Z(n26769) );
  NANDN U26915 ( .A(n26771), .B(n26770), .Z(n26766) );
  ANDN U26916 ( .B(B[195]), .A(n68), .Z(n26550) );
  XNOR U26917 ( .A(n26558), .B(n26772), .Z(n26551) );
  XNOR U26918 ( .A(n26557), .B(n26555), .Z(n26772) );
  AND U26919 ( .A(n26773), .B(n26774), .Z(n26555) );
  NANDN U26920 ( .A(n26775), .B(n26776), .Z(n26774) );
  OR U26921 ( .A(n26777), .B(n26778), .Z(n26776) );
  NAND U26922 ( .A(n26778), .B(n26777), .Z(n26773) );
  ANDN U26923 ( .B(B[196]), .A(n69), .Z(n26557) );
  XNOR U26924 ( .A(n26565), .B(n26779), .Z(n26558) );
  XNOR U26925 ( .A(n26564), .B(n26562), .Z(n26779) );
  AND U26926 ( .A(n26780), .B(n26781), .Z(n26562) );
  NANDN U26927 ( .A(n26782), .B(n26783), .Z(n26781) );
  NANDN U26928 ( .A(n26784), .B(n26785), .Z(n26783) );
  NANDN U26929 ( .A(n26785), .B(n26784), .Z(n26780) );
  ANDN U26930 ( .B(B[197]), .A(n70), .Z(n26564) );
  XNOR U26931 ( .A(n26572), .B(n26786), .Z(n26565) );
  XNOR U26932 ( .A(n26571), .B(n26569), .Z(n26786) );
  AND U26933 ( .A(n26787), .B(n26788), .Z(n26569) );
  NANDN U26934 ( .A(n26789), .B(n26790), .Z(n26788) );
  OR U26935 ( .A(n26791), .B(n26792), .Z(n26790) );
  NAND U26936 ( .A(n26792), .B(n26791), .Z(n26787) );
  ANDN U26937 ( .B(B[198]), .A(n71), .Z(n26571) );
  XNOR U26938 ( .A(n26579), .B(n26793), .Z(n26572) );
  XNOR U26939 ( .A(n26578), .B(n26576), .Z(n26793) );
  AND U26940 ( .A(n26794), .B(n26795), .Z(n26576) );
  NANDN U26941 ( .A(n26796), .B(n26797), .Z(n26795) );
  NANDN U26942 ( .A(n26798), .B(n26799), .Z(n26797) );
  NANDN U26943 ( .A(n26799), .B(n26798), .Z(n26794) );
  ANDN U26944 ( .B(B[199]), .A(n72), .Z(n26578) );
  XNOR U26945 ( .A(n26586), .B(n26800), .Z(n26579) );
  XNOR U26946 ( .A(n26585), .B(n26583), .Z(n26800) );
  AND U26947 ( .A(n26801), .B(n26802), .Z(n26583) );
  NANDN U26948 ( .A(n26803), .B(n26804), .Z(n26802) );
  OR U26949 ( .A(n26805), .B(n26806), .Z(n26804) );
  NAND U26950 ( .A(n26806), .B(n26805), .Z(n26801) );
  ANDN U26951 ( .B(B[200]), .A(n73), .Z(n26585) );
  XNOR U26952 ( .A(n26593), .B(n26807), .Z(n26586) );
  XNOR U26953 ( .A(n26592), .B(n26590), .Z(n26807) );
  AND U26954 ( .A(n26808), .B(n26809), .Z(n26590) );
  NANDN U26955 ( .A(n26810), .B(n26811), .Z(n26809) );
  NANDN U26956 ( .A(n26812), .B(n26813), .Z(n26811) );
  NANDN U26957 ( .A(n26813), .B(n26812), .Z(n26808) );
  ANDN U26958 ( .B(B[201]), .A(n74), .Z(n26592) );
  XNOR U26959 ( .A(n26600), .B(n26814), .Z(n26593) );
  XNOR U26960 ( .A(n26599), .B(n26597), .Z(n26814) );
  AND U26961 ( .A(n26815), .B(n26816), .Z(n26597) );
  NANDN U26962 ( .A(n26817), .B(n26818), .Z(n26816) );
  OR U26963 ( .A(n26819), .B(n26820), .Z(n26818) );
  NAND U26964 ( .A(n26820), .B(n26819), .Z(n26815) );
  ANDN U26965 ( .B(B[202]), .A(n75), .Z(n26599) );
  XNOR U26966 ( .A(n26607), .B(n26821), .Z(n26600) );
  XNOR U26967 ( .A(n26606), .B(n26604), .Z(n26821) );
  AND U26968 ( .A(n26822), .B(n26823), .Z(n26604) );
  NANDN U26969 ( .A(n26824), .B(n26825), .Z(n26823) );
  NANDN U26970 ( .A(n26826), .B(n26827), .Z(n26825) );
  NANDN U26971 ( .A(n26827), .B(n26826), .Z(n26822) );
  ANDN U26972 ( .B(B[203]), .A(n76), .Z(n26606) );
  XNOR U26973 ( .A(n26614), .B(n26828), .Z(n26607) );
  XNOR U26974 ( .A(n26613), .B(n26611), .Z(n26828) );
  AND U26975 ( .A(n26829), .B(n26830), .Z(n26611) );
  NANDN U26976 ( .A(n26831), .B(n26832), .Z(n26830) );
  OR U26977 ( .A(n26833), .B(n26834), .Z(n26832) );
  NAND U26978 ( .A(n26834), .B(n26833), .Z(n26829) );
  ANDN U26979 ( .B(B[204]), .A(n77), .Z(n26613) );
  XNOR U26980 ( .A(n26621), .B(n26835), .Z(n26614) );
  XNOR U26981 ( .A(n26620), .B(n26618), .Z(n26835) );
  AND U26982 ( .A(n26836), .B(n26837), .Z(n26618) );
  NANDN U26983 ( .A(n26838), .B(n26839), .Z(n26837) );
  NANDN U26984 ( .A(n26840), .B(n26841), .Z(n26839) );
  NANDN U26985 ( .A(n26841), .B(n26840), .Z(n26836) );
  ANDN U26986 ( .B(B[205]), .A(n78), .Z(n26620) );
  XNOR U26987 ( .A(n26628), .B(n26842), .Z(n26621) );
  XNOR U26988 ( .A(n26627), .B(n26625), .Z(n26842) );
  AND U26989 ( .A(n26843), .B(n26844), .Z(n26625) );
  NANDN U26990 ( .A(n26845), .B(n26846), .Z(n26844) );
  OR U26991 ( .A(n26847), .B(n26848), .Z(n26846) );
  NAND U26992 ( .A(n26848), .B(n26847), .Z(n26843) );
  ANDN U26993 ( .B(B[206]), .A(n79), .Z(n26627) );
  XNOR U26994 ( .A(n26635), .B(n26849), .Z(n26628) );
  XNOR U26995 ( .A(n26634), .B(n26632), .Z(n26849) );
  AND U26996 ( .A(n26850), .B(n26851), .Z(n26632) );
  NANDN U26997 ( .A(n26852), .B(n26853), .Z(n26851) );
  NANDN U26998 ( .A(n26854), .B(n26855), .Z(n26853) );
  NANDN U26999 ( .A(n26855), .B(n26854), .Z(n26850) );
  ANDN U27000 ( .B(B[207]), .A(n80), .Z(n26634) );
  XNOR U27001 ( .A(n26642), .B(n26856), .Z(n26635) );
  XNOR U27002 ( .A(n26641), .B(n26639), .Z(n26856) );
  AND U27003 ( .A(n26857), .B(n26858), .Z(n26639) );
  NANDN U27004 ( .A(n26859), .B(n26860), .Z(n26858) );
  OR U27005 ( .A(n26861), .B(n26862), .Z(n26860) );
  NAND U27006 ( .A(n26862), .B(n26861), .Z(n26857) );
  ANDN U27007 ( .B(B[208]), .A(n81), .Z(n26641) );
  XNOR U27008 ( .A(n26649), .B(n26863), .Z(n26642) );
  XNOR U27009 ( .A(n26648), .B(n26646), .Z(n26863) );
  AND U27010 ( .A(n26864), .B(n26865), .Z(n26646) );
  NANDN U27011 ( .A(n26866), .B(n26867), .Z(n26865) );
  NAND U27012 ( .A(n26868), .B(n26869), .Z(n26867) );
  ANDN U27013 ( .B(B[209]), .A(n82), .Z(n26648) );
  XOR U27014 ( .A(n26655), .B(n26870), .Z(n26649) );
  XNOR U27015 ( .A(n26653), .B(n26656), .Z(n26870) );
  NAND U27016 ( .A(A[2]), .B(B[210]), .Z(n26656) );
  NANDN U27017 ( .A(n26871), .B(n26872), .Z(n26653) );
  AND U27018 ( .A(A[0]), .B(B[211]), .Z(n26872) );
  XNOR U27019 ( .A(n26658), .B(n26873), .Z(n26655) );
  NAND U27020 ( .A(A[0]), .B(B[212]), .Z(n26873) );
  NAND U27021 ( .A(B[211]), .B(A[1]), .Z(n26658) );
  NAND U27022 ( .A(n26874), .B(n26875), .Z(n372) );
  NANDN U27023 ( .A(n26876), .B(n26877), .Z(n26875) );
  OR U27024 ( .A(n26878), .B(n26879), .Z(n26877) );
  NAND U27025 ( .A(n26879), .B(n26878), .Z(n26874) );
  XOR U27026 ( .A(n24605), .B(n26880), .Z(\A1[20] ) );
  XNOR U27027 ( .A(n24604), .B(n24603), .Z(n26880) );
  NAND U27028 ( .A(n26881), .B(n26882), .Z(n24603) );
  NANDN U27029 ( .A(n26883), .B(n26884), .Z(n26882) );
  OR U27030 ( .A(n26885), .B(n26886), .Z(n26884) );
  NAND U27031 ( .A(n26886), .B(n26885), .Z(n26881) );
  ANDN U27032 ( .B(B[0]), .A(n63), .Z(n24604) );
  XNOR U27033 ( .A(n24612), .B(n26887), .Z(n24605) );
  XNOR U27034 ( .A(n24611), .B(n24609), .Z(n26887) );
  AND U27035 ( .A(n26888), .B(n26889), .Z(n24609) );
  NANDN U27036 ( .A(n26890), .B(n26891), .Z(n26889) );
  NANDN U27037 ( .A(n26892), .B(n26893), .Z(n26891) );
  NANDN U27038 ( .A(n26893), .B(n26892), .Z(n26888) );
  ANDN U27039 ( .B(B[1]), .A(n64), .Z(n24611) );
  XNOR U27040 ( .A(n24619), .B(n26894), .Z(n24612) );
  XNOR U27041 ( .A(n24618), .B(n24616), .Z(n26894) );
  AND U27042 ( .A(n26895), .B(n26896), .Z(n24616) );
  NANDN U27043 ( .A(n26897), .B(n26898), .Z(n26896) );
  OR U27044 ( .A(n26899), .B(n26900), .Z(n26898) );
  NAND U27045 ( .A(n26900), .B(n26899), .Z(n26895) );
  ANDN U27046 ( .B(B[2]), .A(n65), .Z(n24618) );
  XNOR U27047 ( .A(n24626), .B(n26901), .Z(n24619) );
  XNOR U27048 ( .A(n24625), .B(n24623), .Z(n26901) );
  AND U27049 ( .A(n26902), .B(n26903), .Z(n24623) );
  NANDN U27050 ( .A(n26904), .B(n26905), .Z(n26903) );
  NANDN U27051 ( .A(n26906), .B(n26907), .Z(n26905) );
  NANDN U27052 ( .A(n26907), .B(n26906), .Z(n26902) );
  ANDN U27053 ( .B(B[3]), .A(n66), .Z(n24625) );
  XNOR U27054 ( .A(n24633), .B(n26908), .Z(n24626) );
  XNOR U27055 ( .A(n24632), .B(n24630), .Z(n26908) );
  AND U27056 ( .A(n26909), .B(n26910), .Z(n24630) );
  NANDN U27057 ( .A(n26911), .B(n26912), .Z(n26910) );
  OR U27058 ( .A(n26913), .B(n26914), .Z(n26912) );
  NAND U27059 ( .A(n26914), .B(n26913), .Z(n26909) );
  ANDN U27060 ( .B(B[4]), .A(n67), .Z(n24632) );
  XNOR U27061 ( .A(n24640), .B(n26915), .Z(n24633) );
  XNOR U27062 ( .A(n24639), .B(n24637), .Z(n26915) );
  AND U27063 ( .A(n26916), .B(n26917), .Z(n24637) );
  NANDN U27064 ( .A(n26918), .B(n26919), .Z(n26917) );
  NANDN U27065 ( .A(n26920), .B(n26921), .Z(n26919) );
  NANDN U27066 ( .A(n26921), .B(n26920), .Z(n26916) );
  ANDN U27067 ( .B(B[5]), .A(n68), .Z(n24639) );
  XNOR U27068 ( .A(n24647), .B(n26922), .Z(n24640) );
  XNOR U27069 ( .A(n24646), .B(n24644), .Z(n26922) );
  AND U27070 ( .A(n26923), .B(n26924), .Z(n24644) );
  NANDN U27071 ( .A(n26925), .B(n26926), .Z(n26924) );
  OR U27072 ( .A(n26927), .B(n26928), .Z(n26926) );
  NAND U27073 ( .A(n26928), .B(n26927), .Z(n26923) );
  ANDN U27074 ( .B(B[6]), .A(n69), .Z(n24646) );
  XNOR U27075 ( .A(n24654), .B(n26929), .Z(n24647) );
  XNOR U27076 ( .A(n24653), .B(n24651), .Z(n26929) );
  AND U27077 ( .A(n26930), .B(n26931), .Z(n24651) );
  NANDN U27078 ( .A(n26932), .B(n26933), .Z(n26931) );
  NANDN U27079 ( .A(n26934), .B(n26935), .Z(n26933) );
  NANDN U27080 ( .A(n26935), .B(n26934), .Z(n26930) );
  ANDN U27081 ( .B(B[7]), .A(n70), .Z(n24653) );
  XNOR U27082 ( .A(n24661), .B(n26936), .Z(n24654) );
  XNOR U27083 ( .A(n24660), .B(n24658), .Z(n26936) );
  AND U27084 ( .A(n26937), .B(n26938), .Z(n24658) );
  NANDN U27085 ( .A(n26939), .B(n26940), .Z(n26938) );
  OR U27086 ( .A(n26941), .B(n26942), .Z(n26940) );
  NAND U27087 ( .A(n26942), .B(n26941), .Z(n26937) );
  ANDN U27088 ( .B(B[8]), .A(n71), .Z(n24660) );
  XNOR U27089 ( .A(n24668), .B(n26943), .Z(n24661) );
  XNOR U27090 ( .A(n24667), .B(n24665), .Z(n26943) );
  AND U27091 ( .A(n26944), .B(n26945), .Z(n24665) );
  NANDN U27092 ( .A(n26946), .B(n26947), .Z(n26945) );
  NANDN U27093 ( .A(n26948), .B(n26949), .Z(n26947) );
  NANDN U27094 ( .A(n26949), .B(n26948), .Z(n26944) );
  ANDN U27095 ( .B(B[9]), .A(n72), .Z(n24667) );
  XNOR U27096 ( .A(n24675), .B(n26950), .Z(n24668) );
  XNOR U27097 ( .A(n24674), .B(n24672), .Z(n26950) );
  AND U27098 ( .A(n26951), .B(n26952), .Z(n24672) );
  NANDN U27099 ( .A(n26953), .B(n26954), .Z(n26952) );
  OR U27100 ( .A(n26955), .B(n26956), .Z(n26954) );
  NAND U27101 ( .A(n26956), .B(n26955), .Z(n26951) );
  ANDN U27102 ( .B(B[10]), .A(n73), .Z(n24674) );
  XNOR U27103 ( .A(n24682), .B(n26957), .Z(n24675) );
  XNOR U27104 ( .A(n24681), .B(n24679), .Z(n26957) );
  AND U27105 ( .A(n26958), .B(n26959), .Z(n24679) );
  NANDN U27106 ( .A(n26960), .B(n26961), .Z(n26959) );
  NANDN U27107 ( .A(n26962), .B(n26963), .Z(n26961) );
  NANDN U27108 ( .A(n26963), .B(n26962), .Z(n26958) );
  ANDN U27109 ( .B(B[11]), .A(n74), .Z(n24681) );
  XNOR U27110 ( .A(n24689), .B(n26964), .Z(n24682) );
  XNOR U27111 ( .A(n24688), .B(n24686), .Z(n26964) );
  AND U27112 ( .A(n26965), .B(n26966), .Z(n24686) );
  NANDN U27113 ( .A(n26967), .B(n26968), .Z(n26966) );
  OR U27114 ( .A(n26969), .B(n26970), .Z(n26968) );
  NAND U27115 ( .A(n26970), .B(n26969), .Z(n26965) );
  ANDN U27116 ( .B(B[12]), .A(n75), .Z(n24688) );
  XNOR U27117 ( .A(n24696), .B(n26971), .Z(n24689) );
  XNOR U27118 ( .A(n24695), .B(n24693), .Z(n26971) );
  AND U27119 ( .A(n26972), .B(n26973), .Z(n24693) );
  NANDN U27120 ( .A(n26974), .B(n26975), .Z(n26973) );
  NANDN U27121 ( .A(n26976), .B(n26977), .Z(n26975) );
  NANDN U27122 ( .A(n26977), .B(n26976), .Z(n26972) );
  ANDN U27123 ( .B(B[13]), .A(n76), .Z(n24695) );
  XNOR U27124 ( .A(n24703), .B(n26978), .Z(n24696) );
  XNOR U27125 ( .A(n24702), .B(n24700), .Z(n26978) );
  AND U27126 ( .A(n26979), .B(n26980), .Z(n24700) );
  NANDN U27127 ( .A(n26981), .B(n26982), .Z(n26980) );
  OR U27128 ( .A(n26983), .B(n26984), .Z(n26982) );
  NAND U27129 ( .A(n26984), .B(n26983), .Z(n26979) );
  ANDN U27130 ( .B(B[14]), .A(n77), .Z(n24702) );
  XNOR U27131 ( .A(n24710), .B(n26985), .Z(n24703) );
  XNOR U27132 ( .A(n24709), .B(n24707), .Z(n26985) );
  AND U27133 ( .A(n26986), .B(n26987), .Z(n24707) );
  NANDN U27134 ( .A(n26988), .B(n26989), .Z(n26987) );
  NANDN U27135 ( .A(n26990), .B(n26991), .Z(n26989) );
  NANDN U27136 ( .A(n26991), .B(n26990), .Z(n26986) );
  ANDN U27137 ( .B(B[15]), .A(n78), .Z(n24709) );
  XNOR U27138 ( .A(n24717), .B(n26992), .Z(n24710) );
  XNOR U27139 ( .A(n24716), .B(n24714), .Z(n26992) );
  AND U27140 ( .A(n26993), .B(n26994), .Z(n24714) );
  NANDN U27141 ( .A(n26995), .B(n26996), .Z(n26994) );
  OR U27142 ( .A(n26997), .B(n26998), .Z(n26996) );
  NAND U27143 ( .A(n26998), .B(n26997), .Z(n26993) );
  ANDN U27144 ( .B(B[16]), .A(n79), .Z(n24716) );
  XNOR U27145 ( .A(n24724), .B(n26999), .Z(n24717) );
  XNOR U27146 ( .A(n24723), .B(n24721), .Z(n26999) );
  AND U27147 ( .A(n27000), .B(n27001), .Z(n24721) );
  NANDN U27148 ( .A(n27002), .B(n27003), .Z(n27001) );
  NANDN U27149 ( .A(n27004), .B(n27005), .Z(n27003) );
  NANDN U27150 ( .A(n27005), .B(n27004), .Z(n27000) );
  ANDN U27151 ( .B(B[17]), .A(n80), .Z(n24723) );
  XNOR U27152 ( .A(n24731), .B(n27006), .Z(n24724) );
  XNOR U27153 ( .A(n24730), .B(n24728), .Z(n27006) );
  AND U27154 ( .A(n27007), .B(n27008), .Z(n24728) );
  NANDN U27155 ( .A(n27009), .B(n27010), .Z(n27008) );
  OR U27156 ( .A(n27011), .B(n27012), .Z(n27010) );
  NAND U27157 ( .A(n27012), .B(n27011), .Z(n27007) );
  ANDN U27158 ( .B(B[18]), .A(n81), .Z(n24730) );
  XNOR U27159 ( .A(n24738), .B(n27013), .Z(n24731) );
  XNOR U27160 ( .A(n24737), .B(n24735), .Z(n27013) );
  AND U27161 ( .A(n27014), .B(n27015), .Z(n24735) );
  NANDN U27162 ( .A(n27016), .B(n27017), .Z(n27015) );
  NAND U27163 ( .A(n27018), .B(n27019), .Z(n27017) );
  ANDN U27164 ( .B(B[19]), .A(n82), .Z(n24737) );
  XOR U27165 ( .A(n24744), .B(n27020), .Z(n24738) );
  XNOR U27166 ( .A(n24742), .B(n24745), .Z(n27020) );
  NAND U27167 ( .A(A[2]), .B(B[20]), .Z(n24745) );
  NANDN U27168 ( .A(n27021), .B(n27022), .Z(n24742) );
  AND U27169 ( .A(A[0]), .B(B[21]), .Z(n27022) );
  XNOR U27170 ( .A(n24747), .B(n27023), .Z(n24744) );
  NAND U27171 ( .A(A[0]), .B(B[22]), .Z(n27023) );
  NAND U27172 ( .A(B[21]), .B(A[1]), .Z(n24747) );
  XOR U27173 ( .A(n374), .B(n373), .Z(\A1[209] ) );
  XOR U27174 ( .A(n26879), .B(n27024), .Z(n373) );
  XNOR U27175 ( .A(n26878), .B(n26876), .Z(n27024) );
  AND U27176 ( .A(n27025), .B(n27026), .Z(n26876) );
  NANDN U27177 ( .A(n27027), .B(n27028), .Z(n27026) );
  NANDN U27178 ( .A(n27029), .B(n27030), .Z(n27028) );
  NANDN U27179 ( .A(n27030), .B(n27029), .Z(n27025) );
  ANDN U27180 ( .B(B[180]), .A(n54), .Z(n26878) );
  XNOR U27181 ( .A(n26673), .B(n27031), .Z(n26879) );
  XNOR U27182 ( .A(n26672), .B(n26670), .Z(n27031) );
  AND U27183 ( .A(n27032), .B(n27033), .Z(n26670) );
  NANDN U27184 ( .A(n27034), .B(n27035), .Z(n27033) );
  OR U27185 ( .A(n27036), .B(n27037), .Z(n27035) );
  NAND U27186 ( .A(n27037), .B(n27036), .Z(n27032) );
  ANDN U27187 ( .B(B[181]), .A(n55), .Z(n26672) );
  XNOR U27188 ( .A(n26680), .B(n27038), .Z(n26673) );
  XNOR U27189 ( .A(n26679), .B(n26677), .Z(n27038) );
  AND U27190 ( .A(n27039), .B(n27040), .Z(n26677) );
  NANDN U27191 ( .A(n27041), .B(n27042), .Z(n27040) );
  NANDN U27192 ( .A(n27043), .B(n27044), .Z(n27042) );
  NANDN U27193 ( .A(n27044), .B(n27043), .Z(n27039) );
  ANDN U27194 ( .B(B[182]), .A(n56), .Z(n26679) );
  XNOR U27195 ( .A(n26687), .B(n27045), .Z(n26680) );
  XNOR U27196 ( .A(n26686), .B(n26684), .Z(n27045) );
  AND U27197 ( .A(n27046), .B(n27047), .Z(n26684) );
  NANDN U27198 ( .A(n27048), .B(n27049), .Z(n27047) );
  OR U27199 ( .A(n27050), .B(n27051), .Z(n27049) );
  NAND U27200 ( .A(n27051), .B(n27050), .Z(n27046) );
  ANDN U27201 ( .B(B[183]), .A(n57), .Z(n26686) );
  XNOR U27202 ( .A(n26694), .B(n27052), .Z(n26687) );
  XNOR U27203 ( .A(n26693), .B(n26691), .Z(n27052) );
  AND U27204 ( .A(n27053), .B(n27054), .Z(n26691) );
  NANDN U27205 ( .A(n27055), .B(n27056), .Z(n27054) );
  NANDN U27206 ( .A(n27057), .B(n27058), .Z(n27056) );
  NANDN U27207 ( .A(n27058), .B(n27057), .Z(n27053) );
  ANDN U27208 ( .B(B[184]), .A(n58), .Z(n26693) );
  XNOR U27209 ( .A(n26701), .B(n27059), .Z(n26694) );
  XNOR U27210 ( .A(n26700), .B(n26698), .Z(n27059) );
  AND U27211 ( .A(n27060), .B(n27061), .Z(n26698) );
  NANDN U27212 ( .A(n27062), .B(n27063), .Z(n27061) );
  OR U27213 ( .A(n27064), .B(n27065), .Z(n27063) );
  NAND U27214 ( .A(n27065), .B(n27064), .Z(n27060) );
  ANDN U27215 ( .B(B[185]), .A(n59), .Z(n26700) );
  XNOR U27216 ( .A(n26708), .B(n27066), .Z(n26701) );
  XNOR U27217 ( .A(n26707), .B(n26705), .Z(n27066) );
  AND U27218 ( .A(n27067), .B(n27068), .Z(n26705) );
  NANDN U27219 ( .A(n27069), .B(n27070), .Z(n27068) );
  NANDN U27220 ( .A(n27071), .B(n27072), .Z(n27070) );
  NANDN U27221 ( .A(n27072), .B(n27071), .Z(n27067) );
  ANDN U27222 ( .B(B[186]), .A(n60), .Z(n26707) );
  XNOR U27223 ( .A(n26715), .B(n27073), .Z(n26708) );
  XNOR U27224 ( .A(n26714), .B(n26712), .Z(n27073) );
  AND U27225 ( .A(n27074), .B(n27075), .Z(n26712) );
  NANDN U27226 ( .A(n27076), .B(n27077), .Z(n27075) );
  OR U27227 ( .A(n27078), .B(n27079), .Z(n27077) );
  NAND U27228 ( .A(n27079), .B(n27078), .Z(n27074) );
  ANDN U27229 ( .B(B[187]), .A(n61), .Z(n26714) );
  XNOR U27230 ( .A(n26722), .B(n27080), .Z(n26715) );
  XNOR U27231 ( .A(n26721), .B(n26719), .Z(n27080) );
  AND U27232 ( .A(n27081), .B(n27082), .Z(n26719) );
  NANDN U27233 ( .A(n27083), .B(n27084), .Z(n27082) );
  NANDN U27234 ( .A(n27085), .B(n27086), .Z(n27084) );
  NANDN U27235 ( .A(n27086), .B(n27085), .Z(n27081) );
  ANDN U27236 ( .B(B[188]), .A(n62), .Z(n26721) );
  XNOR U27237 ( .A(n26729), .B(n27087), .Z(n26722) );
  XNOR U27238 ( .A(n26728), .B(n26726), .Z(n27087) );
  AND U27239 ( .A(n27088), .B(n27089), .Z(n26726) );
  NANDN U27240 ( .A(n27090), .B(n27091), .Z(n27089) );
  OR U27241 ( .A(n27092), .B(n27093), .Z(n27091) );
  NAND U27242 ( .A(n27093), .B(n27092), .Z(n27088) );
  ANDN U27243 ( .B(B[189]), .A(n63), .Z(n26728) );
  XNOR U27244 ( .A(n26736), .B(n27094), .Z(n26729) );
  XNOR U27245 ( .A(n26735), .B(n26733), .Z(n27094) );
  AND U27246 ( .A(n27095), .B(n27096), .Z(n26733) );
  NANDN U27247 ( .A(n27097), .B(n27098), .Z(n27096) );
  NANDN U27248 ( .A(n27099), .B(n27100), .Z(n27098) );
  NANDN U27249 ( .A(n27100), .B(n27099), .Z(n27095) );
  ANDN U27250 ( .B(B[190]), .A(n64), .Z(n26735) );
  XNOR U27251 ( .A(n26743), .B(n27101), .Z(n26736) );
  XNOR U27252 ( .A(n26742), .B(n26740), .Z(n27101) );
  AND U27253 ( .A(n27102), .B(n27103), .Z(n26740) );
  NANDN U27254 ( .A(n27104), .B(n27105), .Z(n27103) );
  OR U27255 ( .A(n27106), .B(n27107), .Z(n27105) );
  NAND U27256 ( .A(n27107), .B(n27106), .Z(n27102) );
  ANDN U27257 ( .B(B[191]), .A(n65), .Z(n26742) );
  XNOR U27258 ( .A(n26750), .B(n27108), .Z(n26743) );
  XNOR U27259 ( .A(n26749), .B(n26747), .Z(n27108) );
  AND U27260 ( .A(n27109), .B(n27110), .Z(n26747) );
  NANDN U27261 ( .A(n27111), .B(n27112), .Z(n27110) );
  NANDN U27262 ( .A(n27113), .B(n27114), .Z(n27112) );
  NANDN U27263 ( .A(n27114), .B(n27113), .Z(n27109) );
  ANDN U27264 ( .B(B[192]), .A(n66), .Z(n26749) );
  XNOR U27265 ( .A(n26757), .B(n27115), .Z(n26750) );
  XNOR U27266 ( .A(n26756), .B(n26754), .Z(n27115) );
  AND U27267 ( .A(n27116), .B(n27117), .Z(n26754) );
  NANDN U27268 ( .A(n27118), .B(n27119), .Z(n27117) );
  OR U27269 ( .A(n27120), .B(n27121), .Z(n27119) );
  NAND U27270 ( .A(n27121), .B(n27120), .Z(n27116) );
  ANDN U27271 ( .B(B[193]), .A(n67), .Z(n26756) );
  XNOR U27272 ( .A(n26764), .B(n27122), .Z(n26757) );
  XNOR U27273 ( .A(n26763), .B(n26761), .Z(n27122) );
  AND U27274 ( .A(n27123), .B(n27124), .Z(n26761) );
  NANDN U27275 ( .A(n27125), .B(n27126), .Z(n27124) );
  NANDN U27276 ( .A(n27127), .B(n27128), .Z(n27126) );
  NANDN U27277 ( .A(n27128), .B(n27127), .Z(n27123) );
  ANDN U27278 ( .B(B[194]), .A(n68), .Z(n26763) );
  XNOR U27279 ( .A(n26771), .B(n27129), .Z(n26764) );
  XNOR U27280 ( .A(n26770), .B(n26768), .Z(n27129) );
  AND U27281 ( .A(n27130), .B(n27131), .Z(n26768) );
  NANDN U27282 ( .A(n27132), .B(n27133), .Z(n27131) );
  OR U27283 ( .A(n27134), .B(n27135), .Z(n27133) );
  NAND U27284 ( .A(n27135), .B(n27134), .Z(n27130) );
  ANDN U27285 ( .B(B[195]), .A(n69), .Z(n26770) );
  XNOR U27286 ( .A(n26778), .B(n27136), .Z(n26771) );
  XNOR U27287 ( .A(n26777), .B(n26775), .Z(n27136) );
  AND U27288 ( .A(n27137), .B(n27138), .Z(n26775) );
  NANDN U27289 ( .A(n27139), .B(n27140), .Z(n27138) );
  NANDN U27290 ( .A(n27141), .B(n27142), .Z(n27140) );
  NANDN U27291 ( .A(n27142), .B(n27141), .Z(n27137) );
  ANDN U27292 ( .B(B[196]), .A(n70), .Z(n26777) );
  XNOR U27293 ( .A(n26785), .B(n27143), .Z(n26778) );
  XNOR U27294 ( .A(n26784), .B(n26782), .Z(n27143) );
  AND U27295 ( .A(n27144), .B(n27145), .Z(n26782) );
  NANDN U27296 ( .A(n27146), .B(n27147), .Z(n27145) );
  OR U27297 ( .A(n27148), .B(n27149), .Z(n27147) );
  NAND U27298 ( .A(n27149), .B(n27148), .Z(n27144) );
  ANDN U27299 ( .B(B[197]), .A(n71), .Z(n26784) );
  XNOR U27300 ( .A(n26792), .B(n27150), .Z(n26785) );
  XNOR U27301 ( .A(n26791), .B(n26789), .Z(n27150) );
  AND U27302 ( .A(n27151), .B(n27152), .Z(n26789) );
  NANDN U27303 ( .A(n27153), .B(n27154), .Z(n27152) );
  NANDN U27304 ( .A(n27155), .B(n27156), .Z(n27154) );
  NANDN U27305 ( .A(n27156), .B(n27155), .Z(n27151) );
  ANDN U27306 ( .B(B[198]), .A(n72), .Z(n26791) );
  XNOR U27307 ( .A(n26799), .B(n27157), .Z(n26792) );
  XNOR U27308 ( .A(n26798), .B(n26796), .Z(n27157) );
  AND U27309 ( .A(n27158), .B(n27159), .Z(n26796) );
  NANDN U27310 ( .A(n27160), .B(n27161), .Z(n27159) );
  OR U27311 ( .A(n27162), .B(n27163), .Z(n27161) );
  NAND U27312 ( .A(n27163), .B(n27162), .Z(n27158) );
  ANDN U27313 ( .B(B[199]), .A(n73), .Z(n26798) );
  XNOR U27314 ( .A(n26806), .B(n27164), .Z(n26799) );
  XNOR U27315 ( .A(n26805), .B(n26803), .Z(n27164) );
  AND U27316 ( .A(n27165), .B(n27166), .Z(n26803) );
  NANDN U27317 ( .A(n27167), .B(n27168), .Z(n27166) );
  NANDN U27318 ( .A(n27169), .B(n27170), .Z(n27168) );
  NANDN U27319 ( .A(n27170), .B(n27169), .Z(n27165) );
  ANDN U27320 ( .B(B[200]), .A(n74), .Z(n26805) );
  XNOR U27321 ( .A(n26813), .B(n27171), .Z(n26806) );
  XNOR U27322 ( .A(n26812), .B(n26810), .Z(n27171) );
  AND U27323 ( .A(n27172), .B(n27173), .Z(n26810) );
  NANDN U27324 ( .A(n27174), .B(n27175), .Z(n27173) );
  OR U27325 ( .A(n27176), .B(n27177), .Z(n27175) );
  NAND U27326 ( .A(n27177), .B(n27176), .Z(n27172) );
  ANDN U27327 ( .B(B[201]), .A(n75), .Z(n26812) );
  XNOR U27328 ( .A(n26820), .B(n27178), .Z(n26813) );
  XNOR U27329 ( .A(n26819), .B(n26817), .Z(n27178) );
  AND U27330 ( .A(n27179), .B(n27180), .Z(n26817) );
  NANDN U27331 ( .A(n27181), .B(n27182), .Z(n27180) );
  NANDN U27332 ( .A(n27183), .B(n27184), .Z(n27182) );
  NANDN U27333 ( .A(n27184), .B(n27183), .Z(n27179) );
  ANDN U27334 ( .B(B[202]), .A(n76), .Z(n26819) );
  XNOR U27335 ( .A(n26827), .B(n27185), .Z(n26820) );
  XNOR U27336 ( .A(n26826), .B(n26824), .Z(n27185) );
  AND U27337 ( .A(n27186), .B(n27187), .Z(n26824) );
  NANDN U27338 ( .A(n27188), .B(n27189), .Z(n27187) );
  OR U27339 ( .A(n27190), .B(n27191), .Z(n27189) );
  NAND U27340 ( .A(n27191), .B(n27190), .Z(n27186) );
  ANDN U27341 ( .B(B[203]), .A(n77), .Z(n26826) );
  XNOR U27342 ( .A(n26834), .B(n27192), .Z(n26827) );
  XNOR U27343 ( .A(n26833), .B(n26831), .Z(n27192) );
  AND U27344 ( .A(n27193), .B(n27194), .Z(n26831) );
  NANDN U27345 ( .A(n27195), .B(n27196), .Z(n27194) );
  NANDN U27346 ( .A(n27197), .B(n27198), .Z(n27196) );
  NANDN U27347 ( .A(n27198), .B(n27197), .Z(n27193) );
  ANDN U27348 ( .B(B[204]), .A(n78), .Z(n26833) );
  XNOR U27349 ( .A(n26841), .B(n27199), .Z(n26834) );
  XNOR U27350 ( .A(n26840), .B(n26838), .Z(n27199) );
  AND U27351 ( .A(n27200), .B(n27201), .Z(n26838) );
  NANDN U27352 ( .A(n27202), .B(n27203), .Z(n27201) );
  OR U27353 ( .A(n27204), .B(n27205), .Z(n27203) );
  NAND U27354 ( .A(n27205), .B(n27204), .Z(n27200) );
  ANDN U27355 ( .B(B[205]), .A(n79), .Z(n26840) );
  XNOR U27356 ( .A(n26848), .B(n27206), .Z(n26841) );
  XNOR U27357 ( .A(n26847), .B(n26845), .Z(n27206) );
  AND U27358 ( .A(n27207), .B(n27208), .Z(n26845) );
  NANDN U27359 ( .A(n27209), .B(n27210), .Z(n27208) );
  NANDN U27360 ( .A(n27211), .B(n27212), .Z(n27210) );
  NANDN U27361 ( .A(n27212), .B(n27211), .Z(n27207) );
  ANDN U27362 ( .B(B[206]), .A(n80), .Z(n26847) );
  XNOR U27363 ( .A(n26855), .B(n27213), .Z(n26848) );
  XNOR U27364 ( .A(n26854), .B(n26852), .Z(n27213) );
  AND U27365 ( .A(n27214), .B(n27215), .Z(n26852) );
  NANDN U27366 ( .A(n27216), .B(n27217), .Z(n27215) );
  OR U27367 ( .A(n27218), .B(n27219), .Z(n27217) );
  NAND U27368 ( .A(n27219), .B(n27218), .Z(n27214) );
  ANDN U27369 ( .B(B[207]), .A(n81), .Z(n26854) );
  XNOR U27370 ( .A(n26862), .B(n27220), .Z(n26855) );
  XNOR U27371 ( .A(n26861), .B(n26859), .Z(n27220) );
  AND U27372 ( .A(n27221), .B(n27222), .Z(n26859) );
  NANDN U27373 ( .A(n27223), .B(n27224), .Z(n27222) );
  NAND U27374 ( .A(n27225), .B(n27226), .Z(n27224) );
  ANDN U27375 ( .B(B[208]), .A(n82), .Z(n26861) );
  XOR U27376 ( .A(n26868), .B(n27227), .Z(n26862) );
  XNOR U27377 ( .A(n26866), .B(n26869), .Z(n27227) );
  NAND U27378 ( .A(A[2]), .B(B[209]), .Z(n26869) );
  NANDN U27379 ( .A(n27228), .B(n27229), .Z(n26866) );
  AND U27380 ( .A(A[0]), .B(B[210]), .Z(n27229) );
  XNOR U27381 ( .A(n26871), .B(n27230), .Z(n26868) );
  NAND U27382 ( .A(A[0]), .B(B[211]), .Z(n27230) );
  NAND U27383 ( .A(B[210]), .B(A[1]), .Z(n26871) );
  NAND U27384 ( .A(n27231), .B(n27232), .Z(n374) );
  NANDN U27385 ( .A(n27233), .B(n27234), .Z(n27232) );
  OR U27386 ( .A(n27235), .B(n27236), .Z(n27234) );
  NAND U27387 ( .A(n27236), .B(n27235), .Z(n27231) );
  XOR U27388 ( .A(n376), .B(n375), .Z(\A1[208] ) );
  XOR U27389 ( .A(n27236), .B(n27237), .Z(n375) );
  XNOR U27390 ( .A(n27235), .B(n27233), .Z(n27237) );
  AND U27391 ( .A(n27238), .B(n27239), .Z(n27233) );
  NANDN U27392 ( .A(n27240), .B(n27241), .Z(n27239) );
  NANDN U27393 ( .A(n27242), .B(n27243), .Z(n27241) );
  NANDN U27394 ( .A(n27243), .B(n27242), .Z(n27238) );
  ANDN U27395 ( .B(B[179]), .A(n54), .Z(n27235) );
  XNOR U27396 ( .A(n27030), .B(n27244), .Z(n27236) );
  XNOR U27397 ( .A(n27029), .B(n27027), .Z(n27244) );
  AND U27398 ( .A(n27245), .B(n27246), .Z(n27027) );
  NANDN U27399 ( .A(n27247), .B(n27248), .Z(n27246) );
  OR U27400 ( .A(n27249), .B(n27250), .Z(n27248) );
  NAND U27401 ( .A(n27250), .B(n27249), .Z(n27245) );
  ANDN U27402 ( .B(B[180]), .A(n55), .Z(n27029) );
  XNOR U27403 ( .A(n27037), .B(n27251), .Z(n27030) );
  XNOR U27404 ( .A(n27036), .B(n27034), .Z(n27251) );
  AND U27405 ( .A(n27252), .B(n27253), .Z(n27034) );
  NANDN U27406 ( .A(n27254), .B(n27255), .Z(n27253) );
  NANDN U27407 ( .A(n27256), .B(n27257), .Z(n27255) );
  NANDN U27408 ( .A(n27257), .B(n27256), .Z(n27252) );
  ANDN U27409 ( .B(B[181]), .A(n56), .Z(n27036) );
  XNOR U27410 ( .A(n27044), .B(n27258), .Z(n27037) );
  XNOR U27411 ( .A(n27043), .B(n27041), .Z(n27258) );
  AND U27412 ( .A(n27259), .B(n27260), .Z(n27041) );
  NANDN U27413 ( .A(n27261), .B(n27262), .Z(n27260) );
  OR U27414 ( .A(n27263), .B(n27264), .Z(n27262) );
  NAND U27415 ( .A(n27264), .B(n27263), .Z(n27259) );
  ANDN U27416 ( .B(B[182]), .A(n57), .Z(n27043) );
  XNOR U27417 ( .A(n27051), .B(n27265), .Z(n27044) );
  XNOR U27418 ( .A(n27050), .B(n27048), .Z(n27265) );
  AND U27419 ( .A(n27266), .B(n27267), .Z(n27048) );
  NANDN U27420 ( .A(n27268), .B(n27269), .Z(n27267) );
  NANDN U27421 ( .A(n27270), .B(n27271), .Z(n27269) );
  NANDN U27422 ( .A(n27271), .B(n27270), .Z(n27266) );
  ANDN U27423 ( .B(B[183]), .A(n58), .Z(n27050) );
  XNOR U27424 ( .A(n27058), .B(n27272), .Z(n27051) );
  XNOR U27425 ( .A(n27057), .B(n27055), .Z(n27272) );
  AND U27426 ( .A(n27273), .B(n27274), .Z(n27055) );
  NANDN U27427 ( .A(n27275), .B(n27276), .Z(n27274) );
  OR U27428 ( .A(n27277), .B(n27278), .Z(n27276) );
  NAND U27429 ( .A(n27278), .B(n27277), .Z(n27273) );
  ANDN U27430 ( .B(B[184]), .A(n59), .Z(n27057) );
  XNOR U27431 ( .A(n27065), .B(n27279), .Z(n27058) );
  XNOR U27432 ( .A(n27064), .B(n27062), .Z(n27279) );
  AND U27433 ( .A(n27280), .B(n27281), .Z(n27062) );
  NANDN U27434 ( .A(n27282), .B(n27283), .Z(n27281) );
  NANDN U27435 ( .A(n27284), .B(n27285), .Z(n27283) );
  NANDN U27436 ( .A(n27285), .B(n27284), .Z(n27280) );
  ANDN U27437 ( .B(B[185]), .A(n60), .Z(n27064) );
  XNOR U27438 ( .A(n27072), .B(n27286), .Z(n27065) );
  XNOR U27439 ( .A(n27071), .B(n27069), .Z(n27286) );
  AND U27440 ( .A(n27287), .B(n27288), .Z(n27069) );
  NANDN U27441 ( .A(n27289), .B(n27290), .Z(n27288) );
  OR U27442 ( .A(n27291), .B(n27292), .Z(n27290) );
  NAND U27443 ( .A(n27292), .B(n27291), .Z(n27287) );
  ANDN U27444 ( .B(B[186]), .A(n61), .Z(n27071) );
  XNOR U27445 ( .A(n27079), .B(n27293), .Z(n27072) );
  XNOR U27446 ( .A(n27078), .B(n27076), .Z(n27293) );
  AND U27447 ( .A(n27294), .B(n27295), .Z(n27076) );
  NANDN U27448 ( .A(n27296), .B(n27297), .Z(n27295) );
  NANDN U27449 ( .A(n27298), .B(n27299), .Z(n27297) );
  NANDN U27450 ( .A(n27299), .B(n27298), .Z(n27294) );
  ANDN U27451 ( .B(B[187]), .A(n62), .Z(n27078) );
  XNOR U27452 ( .A(n27086), .B(n27300), .Z(n27079) );
  XNOR U27453 ( .A(n27085), .B(n27083), .Z(n27300) );
  AND U27454 ( .A(n27301), .B(n27302), .Z(n27083) );
  NANDN U27455 ( .A(n27303), .B(n27304), .Z(n27302) );
  OR U27456 ( .A(n27305), .B(n27306), .Z(n27304) );
  NAND U27457 ( .A(n27306), .B(n27305), .Z(n27301) );
  ANDN U27458 ( .B(B[188]), .A(n63), .Z(n27085) );
  XNOR U27459 ( .A(n27093), .B(n27307), .Z(n27086) );
  XNOR U27460 ( .A(n27092), .B(n27090), .Z(n27307) );
  AND U27461 ( .A(n27308), .B(n27309), .Z(n27090) );
  NANDN U27462 ( .A(n27310), .B(n27311), .Z(n27309) );
  NANDN U27463 ( .A(n27312), .B(n27313), .Z(n27311) );
  NANDN U27464 ( .A(n27313), .B(n27312), .Z(n27308) );
  ANDN U27465 ( .B(B[189]), .A(n64), .Z(n27092) );
  XNOR U27466 ( .A(n27100), .B(n27314), .Z(n27093) );
  XNOR U27467 ( .A(n27099), .B(n27097), .Z(n27314) );
  AND U27468 ( .A(n27315), .B(n27316), .Z(n27097) );
  NANDN U27469 ( .A(n27317), .B(n27318), .Z(n27316) );
  OR U27470 ( .A(n27319), .B(n27320), .Z(n27318) );
  NAND U27471 ( .A(n27320), .B(n27319), .Z(n27315) );
  ANDN U27472 ( .B(B[190]), .A(n65), .Z(n27099) );
  XNOR U27473 ( .A(n27107), .B(n27321), .Z(n27100) );
  XNOR U27474 ( .A(n27106), .B(n27104), .Z(n27321) );
  AND U27475 ( .A(n27322), .B(n27323), .Z(n27104) );
  NANDN U27476 ( .A(n27324), .B(n27325), .Z(n27323) );
  NANDN U27477 ( .A(n27326), .B(n27327), .Z(n27325) );
  NANDN U27478 ( .A(n27327), .B(n27326), .Z(n27322) );
  ANDN U27479 ( .B(B[191]), .A(n66), .Z(n27106) );
  XNOR U27480 ( .A(n27114), .B(n27328), .Z(n27107) );
  XNOR U27481 ( .A(n27113), .B(n27111), .Z(n27328) );
  AND U27482 ( .A(n27329), .B(n27330), .Z(n27111) );
  NANDN U27483 ( .A(n27331), .B(n27332), .Z(n27330) );
  OR U27484 ( .A(n27333), .B(n27334), .Z(n27332) );
  NAND U27485 ( .A(n27334), .B(n27333), .Z(n27329) );
  ANDN U27486 ( .B(B[192]), .A(n67), .Z(n27113) );
  XNOR U27487 ( .A(n27121), .B(n27335), .Z(n27114) );
  XNOR U27488 ( .A(n27120), .B(n27118), .Z(n27335) );
  AND U27489 ( .A(n27336), .B(n27337), .Z(n27118) );
  NANDN U27490 ( .A(n27338), .B(n27339), .Z(n27337) );
  NANDN U27491 ( .A(n27340), .B(n27341), .Z(n27339) );
  NANDN U27492 ( .A(n27341), .B(n27340), .Z(n27336) );
  ANDN U27493 ( .B(B[193]), .A(n68), .Z(n27120) );
  XNOR U27494 ( .A(n27128), .B(n27342), .Z(n27121) );
  XNOR U27495 ( .A(n27127), .B(n27125), .Z(n27342) );
  AND U27496 ( .A(n27343), .B(n27344), .Z(n27125) );
  NANDN U27497 ( .A(n27345), .B(n27346), .Z(n27344) );
  OR U27498 ( .A(n27347), .B(n27348), .Z(n27346) );
  NAND U27499 ( .A(n27348), .B(n27347), .Z(n27343) );
  ANDN U27500 ( .B(B[194]), .A(n69), .Z(n27127) );
  XNOR U27501 ( .A(n27135), .B(n27349), .Z(n27128) );
  XNOR U27502 ( .A(n27134), .B(n27132), .Z(n27349) );
  AND U27503 ( .A(n27350), .B(n27351), .Z(n27132) );
  NANDN U27504 ( .A(n27352), .B(n27353), .Z(n27351) );
  NANDN U27505 ( .A(n27354), .B(n27355), .Z(n27353) );
  NANDN U27506 ( .A(n27355), .B(n27354), .Z(n27350) );
  ANDN U27507 ( .B(B[195]), .A(n70), .Z(n27134) );
  XNOR U27508 ( .A(n27142), .B(n27356), .Z(n27135) );
  XNOR U27509 ( .A(n27141), .B(n27139), .Z(n27356) );
  AND U27510 ( .A(n27357), .B(n27358), .Z(n27139) );
  NANDN U27511 ( .A(n27359), .B(n27360), .Z(n27358) );
  OR U27512 ( .A(n27361), .B(n27362), .Z(n27360) );
  NAND U27513 ( .A(n27362), .B(n27361), .Z(n27357) );
  ANDN U27514 ( .B(B[196]), .A(n71), .Z(n27141) );
  XNOR U27515 ( .A(n27149), .B(n27363), .Z(n27142) );
  XNOR U27516 ( .A(n27148), .B(n27146), .Z(n27363) );
  AND U27517 ( .A(n27364), .B(n27365), .Z(n27146) );
  NANDN U27518 ( .A(n27366), .B(n27367), .Z(n27365) );
  NANDN U27519 ( .A(n27368), .B(n27369), .Z(n27367) );
  NANDN U27520 ( .A(n27369), .B(n27368), .Z(n27364) );
  ANDN U27521 ( .B(B[197]), .A(n72), .Z(n27148) );
  XNOR U27522 ( .A(n27156), .B(n27370), .Z(n27149) );
  XNOR U27523 ( .A(n27155), .B(n27153), .Z(n27370) );
  AND U27524 ( .A(n27371), .B(n27372), .Z(n27153) );
  NANDN U27525 ( .A(n27373), .B(n27374), .Z(n27372) );
  OR U27526 ( .A(n27375), .B(n27376), .Z(n27374) );
  NAND U27527 ( .A(n27376), .B(n27375), .Z(n27371) );
  ANDN U27528 ( .B(B[198]), .A(n73), .Z(n27155) );
  XNOR U27529 ( .A(n27163), .B(n27377), .Z(n27156) );
  XNOR U27530 ( .A(n27162), .B(n27160), .Z(n27377) );
  AND U27531 ( .A(n27378), .B(n27379), .Z(n27160) );
  NANDN U27532 ( .A(n27380), .B(n27381), .Z(n27379) );
  NANDN U27533 ( .A(n27382), .B(n27383), .Z(n27381) );
  NANDN U27534 ( .A(n27383), .B(n27382), .Z(n27378) );
  ANDN U27535 ( .B(B[199]), .A(n74), .Z(n27162) );
  XNOR U27536 ( .A(n27170), .B(n27384), .Z(n27163) );
  XNOR U27537 ( .A(n27169), .B(n27167), .Z(n27384) );
  AND U27538 ( .A(n27385), .B(n27386), .Z(n27167) );
  NANDN U27539 ( .A(n27387), .B(n27388), .Z(n27386) );
  OR U27540 ( .A(n27389), .B(n27390), .Z(n27388) );
  NAND U27541 ( .A(n27390), .B(n27389), .Z(n27385) );
  ANDN U27542 ( .B(B[200]), .A(n75), .Z(n27169) );
  XNOR U27543 ( .A(n27177), .B(n27391), .Z(n27170) );
  XNOR U27544 ( .A(n27176), .B(n27174), .Z(n27391) );
  AND U27545 ( .A(n27392), .B(n27393), .Z(n27174) );
  NANDN U27546 ( .A(n27394), .B(n27395), .Z(n27393) );
  NANDN U27547 ( .A(n27396), .B(n27397), .Z(n27395) );
  NANDN U27548 ( .A(n27397), .B(n27396), .Z(n27392) );
  ANDN U27549 ( .B(B[201]), .A(n76), .Z(n27176) );
  XNOR U27550 ( .A(n27184), .B(n27398), .Z(n27177) );
  XNOR U27551 ( .A(n27183), .B(n27181), .Z(n27398) );
  AND U27552 ( .A(n27399), .B(n27400), .Z(n27181) );
  NANDN U27553 ( .A(n27401), .B(n27402), .Z(n27400) );
  OR U27554 ( .A(n27403), .B(n27404), .Z(n27402) );
  NAND U27555 ( .A(n27404), .B(n27403), .Z(n27399) );
  ANDN U27556 ( .B(B[202]), .A(n77), .Z(n27183) );
  XNOR U27557 ( .A(n27191), .B(n27405), .Z(n27184) );
  XNOR U27558 ( .A(n27190), .B(n27188), .Z(n27405) );
  AND U27559 ( .A(n27406), .B(n27407), .Z(n27188) );
  NANDN U27560 ( .A(n27408), .B(n27409), .Z(n27407) );
  NANDN U27561 ( .A(n27410), .B(n27411), .Z(n27409) );
  NANDN U27562 ( .A(n27411), .B(n27410), .Z(n27406) );
  ANDN U27563 ( .B(B[203]), .A(n78), .Z(n27190) );
  XNOR U27564 ( .A(n27198), .B(n27412), .Z(n27191) );
  XNOR U27565 ( .A(n27197), .B(n27195), .Z(n27412) );
  AND U27566 ( .A(n27413), .B(n27414), .Z(n27195) );
  NANDN U27567 ( .A(n27415), .B(n27416), .Z(n27414) );
  OR U27568 ( .A(n27417), .B(n27418), .Z(n27416) );
  NAND U27569 ( .A(n27418), .B(n27417), .Z(n27413) );
  ANDN U27570 ( .B(B[204]), .A(n79), .Z(n27197) );
  XNOR U27571 ( .A(n27205), .B(n27419), .Z(n27198) );
  XNOR U27572 ( .A(n27204), .B(n27202), .Z(n27419) );
  AND U27573 ( .A(n27420), .B(n27421), .Z(n27202) );
  NANDN U27574 ( .A(n27422), .B(n27423), .Z(n27421) );
  NANDN U27575 ( .A(n27424), .B(n27425), .Z(n27423) );
  NANDN U27576 ( .A(n27425), .B(n27424), .Z(n27420) );
  ANDN U27577 ( .B(B[205]), .A(n80), .Z(n27204) );
  XNOR U27578 ( .A(n27212), .B(n27426), .Z(n27205) );
  XNOR U27579 ( .A(n27211), .B(n27209), .Z(n27426) );
  AND U27580 ( .A(n27427), .B(n27428), .Z(n27209) );
  NANDN U27581 ( .A(n27429), .B(n27430), .Z(n27428) );
  OR U27582 ( .A(n27431), .B(n27432), .Z(n27430) );
  NAND U27583 ( .A(n27432), .B(n27431), .Z(n27427) );
  ANDN U27584 ( .B(B[206]), .A(n81), .Z(n27211) );
  XNOR U27585 ( .A(n27219), .B(n27433), .Z(n27212) );
  XNOR U27586 ( .A(n27218), .B(n27216), .Z(n27433) );
  AND U27587 ( .A(n27434), .B(n27435), .Z(n27216) );
  NANDN U27588 ( .A(n27436), .B(n27437), .Z(n27435) );
  NAND U27589 ( .A(n27438), .B(n27439), .Z(n27437) );
  ANDN U27590 ( .B(B[207]), .A(n82), .Z(n27218) );
  XOR U27591 ( .A(n27225), .B(n27440), .Z(n27219) );
  XNOR U27592 ( .A(n27223), .B(n27226), .Z(n27440) );
  NAND U27593 ( .A(A[2]), .B(B[208]), .Z(n27226) );
  NANDN U27594 ( .A(n27441), .B(n27442), .Z(n27223) );
  AND U27595 ( .A(A[0]), .B(B[209]), .Z(n27442) );
  XNOR U27596 ( .A(n27228), .B(n27443), .Z(n27225) );
  NAND U27597 ( .A(A[0]), .B(B[210]), .Z(n27443) );
  NAND U27598 ( .A(B[209]), .B(A[1]), .Z(n27228) );
  NAND U27599 ( .A(n27444), .B(n27445), .Z(n376) );
  NANDN U27600 ( .A(n27446), .B(n27447), .Z(n27445) );
  OR U27601 ( .A(n27448), .B(n27449), .Z(n27447) );
  NAND U27602 ( .A(n27449), .B(n27448), .Z(n27444) );
  XOR U27603 ( .A(n378), .B(n377), .Z(\A1[207] ) );
  XOR U27604 ( .A(n27449), .B(n27450), .Z(n377) );
  XNOR U27605 ( .A(n27448), .B(n27446), .Z(n27450) );
  AND U27606 ( .A(n27451), .B(n27452), .Z(n27446) );
  NANDN U27607 ( .A(n27453), .B(n27454), .Z(n27452) );
  NANDN U27608 ( .A(n27455), .B(n27456), .Z(n27454) );
  NANDN U27609 ( .A(n27456), .B(n27455), .Z(n27451) );
  ANDN U27610 ( .B(B[178]), .A(n54), .Z(n27448) );
  XNOR U27611 ( .A(n27243), .B(n27457), .Z(n27449) );
  XNOR U27612 ( .A(n27242), .B(n27240), .Z(n27457) );
  AND U27613 ( .A(n27458), .B(n27459), .Z(n27240) );
  NANDN U27614 ( .A(n27460), .B(n27461), .Z(n27459) );
  OR U27615 ( .A(n27462), .B(n27463), .Z(n27461) );
  NAND U27616 ( .A(n27463), .B(n27462), .Z(n27458) );
  ANDN U27617 ( .B(B[179]), .A(n55), .Z(n27242) );
  XNOR U27618 ( .A(n27250), .B(n27464), .Z(n27243) );
  XNOR U27619 ( .A(n27249), .B(n27247), .Z(n27464) );
  AND U27620 ( .A(n27465), .B(n27466), .Z(n27247) );
  NANDN U27621 ( .A(n27467), .B(n27468), .Z(n27466) );
  NANDN U27622 ( .A(n27469), .B(n27470), .Z(n27468) );
  NANDN U27623 ( .A(n27470), .B(n27469), .Z(n27465) );
  ANDN U27624 ( .B(B[180]), .A(n56), .Z(n27249) );
  XNOR U27625 ( .A(n27257), .B(n27471), .Z(n27250) );
  XNOR U27626 ( .A(n27256), .B(n27254), .Z(n27471) );
  AND U27627 ( .A(n27472), .B(n27473), .Z(n27254) );
  NANDN U27628 ( .A(n27474), .B(n27475), .Z(n27473) );
  OR U27629 ( .A(n27476), .B(n27477), .Z(n27475) );
  NAND U27630 ( .A(n27477), .B(n27476), .Z(n27472) );
  ANDN U27631 ( .B(B[181]), .A(n57), .Z(n27256) );
  XNOR U27632 ( .A(n27264), .B(n27478), .Z(n27257) );
  XNOR U27633 ( .A(n27263), .B(n27261), .Z(n27478) );
  AND U27634 ( .A(n27479), .B(n27480), .Z(n27261) );
  NANDN U27635 ( .A(n27481), .B(n27482), .Z(n27480) );
  NANDN U27636 ( .A(n27483), .B(n27484), .Z(n27482) );
  NANDN U27637 ( .A(n27484), .B(n27483), .Z(n27479) );
  ANDN U27638 ( .B(B[182]), .A(n58), .Z(n27263) );
  XNOR U27639 ( .A(n27271), .B(n27485), .Z(n27264) );
  XNOR U27640 ( .A(n27270), .B(n27268), .Z(n27485) );
  AND U27641 ( .A(n27486), .B(n27487), .Z(n27268) );
  NANDN U27642 ( .A(n27488), .B(n27489), .Z(n27487) );
  OR U27643 ( .A(n27490), .B(n27491), .Z(n27489) );
  NAND U27644 ( .A(n27491), .B(n27490), .Z(n27486) );
  ANDN U27645 ( .B(B[183]), .A(n59), .Z(n27270) );
  XNOR U27646 ( .A(n27278), .B(n27492), .Z(n27271) );
  XNOR U27647 ( .A(n27277), .B(n27275), .Z(n27492) );
  AND U27648 ( .A(n27493), .B(n27494), .Z(n27275) );
  NANDN U27649 ( .A(n27495), .B(n27496), .Z(n27494) );
  NANDN U27650 ( .A(n27497), .B(n27498), .Z(n27496) );
  NANDN U27651 ( .A(n27498), .B(n27497), .Z(n27493) );
  ANDN U27652 ( .B(B[184]), .A(n60), .Z(n27277) );
  XNOR U27653 ( .A(n27285), .B(n27499), .Z(n27278) );
  XNOR U27654 ( .A(n27284), .B(n27282), .Z(n27499) );
  AND U27655 ( .A(n27500), .B(n27501), .Z(n27282) );
  NANDN U27656 ( .A(n27502), .B(n27503), .Z(n27501) );
  OR U27657 ( .A(n27504), .B(n27505), .Z(n27503) );
  NAND U27658 ( .A(n27505), .B(n27504), .Z(n27500) );
  ANDN U27659 ( .B(B[185]), .A(n61), .Z(n27284) );
  XNOR U27660 ( .A(n27292), .B(n27506), .Z(n27285) );
  XNOR U27661 ( .A(n27291), .B(n27289), .Z(n27506) );
  AND U27662 ( .A(n27507), .B(n27508), .Z(n27289) );
  NANDN U27663 ( .A(n27509), .B(n27510), .Z(n27508) );
  NANDN U27664 ( .A(n27511), .B(n27512), .Z(n27510) );
  NANDN U27665 ( .A(n27512), .B(n27511), .Z(n27507) );
  ANDN U27666 ( .B(B[186]), .A(n62), .Z(n27291) );
  XNOR U27667 ( .A(n27299), .B(n27513), .Z(n27292) );
  XNOR U27668 ( .A(n27298), .B(n27296), .Z(n27513) );
  AND U27669 ( .A(n27514), .B(n27515), .Z(n27296) );
  NANDN U27670 ( .A(n27516), .B(n27517), .Z(n27515) );
  OR U27671 ( .A(n27518), .B(n27519), .Z(n27517) );
  NAND U27672 ( .A(n27519), .B(n27518), .Z(n27514) );
  ANDN U27673 ( .B(B[187]), .A(n63), .Z(n27298) );
  XNOR U27674 ( .A(n27306), .B(n27520), .Z(n27299) );
  XNOR U27675 ( .A(n27305), .B(n27303), .Z(n27520) );
  AND U27676 ( .A(n27521), .B(n27522), .Z(n27303) );
  NANDN U27677 ( .A(n27523), .B(n27524), .Z(n27522) );
  NANDN U27678 ( .A(n27525), .B(n27526), .Z(n27524) );
  NANDN U27679 ( .A(n27526), .B(n27525), .Z(n27521) );
  ANDN U27680 ( .B(B[188]), .A(n64), .Z(n27305) );
  XNOR U27681 ( .A(n27313), .B(n27527), .Z(n27306) );
  XNOR U27682 ( .A(n27312), .B(n27310), .Z(n27527) );
  AND U27683 ( .A(n27528), .B(n27529), .Z(n27310) );
  NANDN U27684 ( .A(n27530), .B(n27531), .Z(n27529) );
  OR U27685 ( .A(n27532), .B(n27533), .Z(n27531) );
  NAND U27686 ( .A(n27533), .B(n27532), .Z(n27528) );
  ANDN U27687 ( .B(B[189]), .A(n65), .Z(n27312) );
  XNOR U27688 ( .A(n27320), .B(n27534), .Z(n27313) );
  XNOR U27689 ( .A(n27319), .B(n27317), .Z(n27534) );
  AND U27690 ( .A(n27535), .B(n27536), .Z(n27317) );
  NANDN U27691 ( .A(n27537), .B(n27538), .Z(n27536) );
  NANDN U27692 ( .A(n27539), .B(n27540), .Z(n27538) );
  NANDN U27693 ( .A(n27540), .B(n27539), .Z(n27535) );
  ANDN U27694 ( .B(B[190]), .A(n66), .Z(n27319) );
  XNOR U27695 ( .A(n27327), .B(n27541), .Z(n27320) );
  XNOR U27696 ( .A(n27326), .B(n27324), .Z(n27541) );
  AND U27697 ( .A(n27542), .B(n27543), .Z(n27324) );
  NANDN U27698 ( .A(n27544), .B(n27545), .Z(n27543) );
  OR U27699 ( .A(n27546), .B(n27547), .Z(n27545) );
  NAND U27700 ( .A(n27547), .B(n27546), .Z(n27542) );
  ANDN U27701 ( .B(B[191]), .A(n67), .Z(n27326) );
  XNOR U27702 ( .A(n27334), .B(n27548), .Z(n27327) );
  XNOR U27703 ( .A(n27333), .B(n27331), .Z(n27548) );
  AND U27704 ( .A(n27549), .B(n27550), .Z(n27331) );
  NANDN U27705 ( .A(n27551), .B(n27552), .Z(n27550) );
  NANDN U27706 ( .A(n27553), .B(n27554), .Z(n27552) );
  NANDN U27707 ( .A(n27554), .B(n27553), .Z(n27549) );
  ANDN U27708 ( .B(B[192]), .A(n68), .Z(n27333) );
  XNOR U27709 ( .A(n27341), .B(n27555), .Z(n27334) );
  XNOR U27710 ( .A(n27340), .B(n27338), .Z(n27555) );
  AND U27711 ( .A(n27556), .B(n27557), .Z(n27338) );
  NANDN U27712 ( .A(n27558), .B(n27559), .Z(n27557) );
  OR U27713 ( .A(n27560), .B(n27561), .Z(n27559) );
  NAND U27714 ( .A(n27561), .B(n27560), .Z(n27556) );
  ANDN U27715 ( .B(B[193]), .A(n69), .Z(n27340) );
  XNOR U27716 ( .A(n27348), .B(n27562), .Z(n27341) );
  XNOR U27717 ( .A(n27347), .B(n27345), .Z(n27562) );
  AND U27718 ( .A(n27563), .B(n27564), .Z(n27345) );
  NANDN U27719 ( .A(n27565), .B(n27566), .Z(n27564) );
  NANDN U27720 ( .A(n27567), .B(n27568), .Z(n27566) );
  NANDN U27721 ( .A(n27568), .B(n27567), .Z(n27563) );
  ANDN U27722 ( .B(B[194]), .A(n70), .Z(n27347) );
  XNOR U27723 ( .A(n27355), .B(n27569), .Z(n27348) );
  XNOR U27724 ( .A(n27354), .B(n27352), .Z(n27569) );
  AND U27725 ( .A(n27570), .B(n27571), .Z(n27352) );
  NANDN U27726 ( .A(n27572), .B(n27573), .Z(n27571) );
  OR U27727 ( .A(n27574), .B(n27575), .Z(n27573) );
  NAND U27728 ( .A(n27575), .B(n27574), .Z(n27570) );
  ANDN U27729 ( .B(B[195]), .A(n71), .Z(n27354) );
  XNOR U27730 ( .A(n27362), .B(n27576), .Z(n27355) );
  XNOR U27731 ( .A(n27361), .B(n27359), .Z(n27576) );
  AND U27732 ( .A(n27577), .B(n27578), .Z(n27359) );
  NANDN U27733 ( .A(n27579), .B(n27580), .Z(n27578) );
  NANDN U27734 ( .A(n27581), .B(n27582), .Z(n27580) );
  NANDN U27735 ( .A(n27582), .B(n27581), .Z(n27577) );
  ANDN U27736 ( .B(B[196]), .A(n72), .Z(n27361) );
  XNOR U27737 ( .A(n27369), .B(n27583), .Z(n27362) );
  XNOR U27738 ( .A(n27368), .B(n27366), .Z(n27583) );
  AND U27739 ( .A(n27584), .B(n27585), .Z(n27366) );
  NANDN U27740 ( .A(n27586), .B(n27587), .Z(n27585) );
  OR U27741 ( .A(n27588), .B(n27589), .Z(n27587) );
  NAND U27742 ( .A(n27589), .B(n27588), .Z(n27584) );
  ANDN U27743 ( .B(B[197]), .A(n73), .Z(n27368) );
  XNOR U27744 ( .A(n27376), .B(n27590), .Z(n27369) );
  XNOR U27745 ( .A(n27375), .B(n27373), .Z(n27590) );
  AND U27746 ( .A(n27591), .B(n27592), .Z(n27373) );
  NANDN U27747 ( .A(n27593), .B(n27594), .Z(n27592) );
  NANDN U27748 ( .A(n27595), .B(n27596), .Z(n27594) );
  NANDN U27749 ( .A(n27596), .B(n27595), .Z(n27591) );
  ANDN U27750 ( .B(B[198]), .A(n74), .Z(n27375) );
  XNOR U27751 ( .A(n27383), .B(n27597), .Z(n27376) );
  XNOR U27752 ( .A(n27382), .B(n27380), .Z(n27597) );
  AND U27753 ( .A(n27598), .B(n27599), .Z(n27380) );
  NANDN U27754 ( .A(n27600), .B(n27601), .Z(n27599) );
  OR U27755 ( .A(n27602), .B(n27603), .Z(n27601) );
  NAND U27756 ( .A(n27603), .B(n27602), .Z(n27598) );
  ANDN U27757 ( .B(B[199]), .A(n75), .Z(n27382) );
  XNOR U27758 ( .A(n27390), .B(n27604), .Z(n27383) );
  XNOR U27759 ( .A(n27389), .B(n27387), .Z(n27604) );
  AND U27760 ( .A(n27605), .B(n27606), .Z(n27387) );
  NANDN U27761 ( .A(n27607), .B(n27608), .Z(n27606) );
  NANDN U27762 ( .A(n27609), .B(n27610), .Z(n27608) );
  NANDN U27763 ( .A(n27610), .B(n27609), .Z(n27605) );
  ANDN U27764 ( .B(B[200]), .A(n76), .Z(n27389) );
  XNOR U27765 ( .A(n27397), .B(n27611), .Z(n27390) );
  XNOR U27766 ( .A(n27396), .B(n27394), .Z(n27611) );
  AND U27767 ( .A(n27612), .B(n27613), .Z(n27394) );
  NANDN U27768 ( .A(n27614), .B(n27615), .Z(n27613) );
  OR U27769 ( .A(n27616), .B(n27617), .Z(n27615) );
  NAND U27770 ( .A(n27617), .B(n27616), .Z(n27612) );
  ANDN U27771 ( .B(B[201]), .A(n77), .Z(n27396) );
  XNOR U27772 ( .A(n27404), .B(n27618), .Z(n27397) );
  XNOR U27773 ( .A(n27403), .B(n27401), .Z(n27618) );
  AND U27774 ( .A(n27619), .B(n27620), .Z(n27401) );
  NANDN U27775 ( .A(n27621), .B(n27622), .Z(n27620) );
  NANDN U27776 ( .A(n27623), .B(n27624), .Z(n27622) );
  NANDN U27777 ( .A(n27624), .B(n27623), .Z(n27619) );
  ANDN U27778 ( .B(B[202]), .A(n78), .Z(n27403) );
  XNOR U27779 ( .A(n27411), .B(n27625), .Z(n27404) );
  XNOR U27780 ( .A(n27410), .B(n27408), .Z(n27625) );
  AND U27781 ( .A(n27626), .B(n27627), .Z(n27408) );
  NANDN U27782 ( .A(n27628), .B(n27629), .Z(n27627) );
  OR U27783 ( .A(n27630), .B(n27631), .Z(n27629) );
  NAND U27784 ( .A(n27631), .B(n27630), .Z(n27626) );
  ANDN U27785 ( .B(B[203]), .A(n79), .Z(n27410) );
  XNOR U27786 ( .A(n27418), .B(n27632), .Z(n27411) );
  XNOR U27787 ( .A(n27417), .B(n27415), .Z(n27632) );
  AND U27788 ( .A(n27633), .B(n27634), .Z(n27415) );
  NANDN U27789 ( .A(n27635), .B(n27636), .Z(n27634) );
  NANDN U27790 ( .A(n27637), .B(n27638), .Z(n27636) );
  NANDN U27791 ( .A(n27638), .B(n27637), .Z(n27633) );
  ANDN U27792 ( .B(B[204]), .A(n80), .Z(n27417) );
  XNOR U27793 ( .A(n27425), .B(n27639), .Z(n27418) );
  XNOR U27794 ( .A(n27424), .B(n27422), .Z(n27639) );
  AND U27795 ( .A(n27640), .B(n27641), .Z(n27422) );
  NANDN U27796 ( .A(n27642), .B(n27643), .Z(n27641) );
  OR U27797 ( .A(n27644), .B(n27645), .Z(n27643) );
  NAND U27798 ( .A(n27645), .B(n27644), .Z(n27640) );
  ANDN U27799 ( .B(B[205]), .A(n81), .Z(n27424) );
  XNOR U27800 ( .A(n27432), .B(n27646), .Z(n27425) );
  XNOR U27801 ( .A(n27431), .B(n27429), .Z(n27646) );
  AND U27802 ( .A(n27647), .B(n27648), .Z(n27429) );
  NANDN U27803 ( .A(n27649), .B(n27650), .Z(n27648) );
  NAND U27804 ( .A(n27651), .B(n27652), .Z(n27650) );
  ANDN U27805 ( .B(B[206]), .A(n82), .Z(n27431) );
  XOR U27806 ( .A(n27438), .B(n27653), .Z(n27432) );
  XNOR U27807 ( .A(n27436), .B(n27439), .Z(n27653) );
  NAND U27808 ( .A(A[2]), .B(B[207]), .Z(n27439) );
  NANDN U27809 ( .A(n27654), .B(n27655), .Z(n27436) );
  AND U27810 ( .A(A[0]), .B(B[208]), .Z(n27655) );
  XNOR U27811 ( .A(n27441), .B(n27656), .Z(n27438) );
  NAND U27812 ( .A(A[0]), .B(B[209]), .Z(n27656) );
  NAND U27813 ( .A(B[208]), .B(A[1]), .Z(n27441) );
  NAND U27814 ( .A(n27657), .B(n27658), .Z(n378) );
  NANDN U27815 ( .A(n27659), .B(n27660), .Z(n27658) );
  OR U27816 ( .A(n27661), .B(n27662), .Z(n27660) );
  NAND U27817 ( .A(n27662), .B(n27661), .Z(n27657) );
  XOR U27818 ( .A(n380), .B(n379), .Z(\A1[206] ) );
  XOR U27819 ( .A(n27662), .B(n27663), .Z(n379) );
  XNOR U27820 ( .A(n27661), .B(n27659), .Z(n27663) );
  AND U27821 ( .A(n27664), .B(n27665), .Z(n27659) );
  NANDN U27822 ( .A(n27666), .B(n27667), .Z(n27665) );
  NANDN U27823 ( .A(n27668), .B(n27669), .Z(n27667) );
  NANDN U27824 ( .A(n27669), .B(n27668), .Z(n27664) );
  ANDN U27825 ( .B(B[177]), .A(n54), .Z(n27661) );
  XNOR U27826 ( .A(n27456), .B(n27670), .Z(n27662) );
  XNOR U27827 ( .A(n27455), .B(n27453), .Z(n27670) );
  AND U27828 ( .A(n27671), .B(n27672), .Z(n27453) );
  NANDN U27829 ( .A(n27673), .B(n27674), .Z(n27672) );
  OR U27830 ( .A(n27675), .B(n27676), .Z(n27674) );
  NAND U27831 ( .A(n27676), .B(n27675), .Z(n27671) );
  ANDN U27832 ( .B(B[178]), .A(n55), .Z(n27455) );
  XNOR U27833 ( .A(n27463), .B(n27677), .Z(n27456) );
  XNOR U27834 ( .A(n27462), .B(n27460), .Z(n27677) );
  AND U27835 ( .A(n27678), .B(n27679), .Z(n27460) );
  NANDN U27836 ( .A(n27680), .B(n27681), .Z(n27679) );
  NANDN U27837 ( .A(n27682), .B(n27683), .Z(n27681) );
  NANDN U27838 ( .A(n27683), .B(n27682), .Z(n27678) );
  ANDN U27839 ( .B(B[179]), .A(n56), .Z(n27462) );
  XNOR U27840 ( .A(n27470), .B(n27684), .Z(n27463) );
  XNOR U27841 ( .A(n27469), .B(n27467), .Z(n27684) );
  AND U27842 ( .A(n27685), .B(n27686), .Z(n27467) );
  NANDN U27843 ( .A(n27687), .B(n27688), .Z(n27686) );
  OR U27844 ( .A(n27689), .B(n27690), .Z(n27688) );
  NAND U27845 ( .A(n27690), .B(n27689), .Z(n27685) );
  ANDN U27846 ( .B(B[180]), .A(n57), .Z(n27469) );
  XNOR U27847 ( .A(n27477), .B(n27691), .Z(n27470) );
  XNOR U27848 ( .A(n27476), .B(n27474), .Z(n27691) );
  AND U27849 ( .A(n27692), .B(n27693), .Z(n27474) );
  NANDN U27850 ( .A(n27694), .B(n27695), .Z(n27693) );
  NANDN U27851 ( .A(n27696), .B(n27697), .Z(n27695) );
  NANDN U27852 ( .A(n27697), .B(n27696), .Z(n27692) );
  ANDN U27853 ( .B(B[181]), .A(n58), .Z(n27476) );
  XNOR U27854 ( .A(n27484), .B(n27698), .Z(n27477) );
  XNOR U27855 ( .A(n27483), .B(n27481), .Z(n27698) );
  AND U27856 ( .A(n27699), .B(n27700), .Z(n27481) );
  NANDN U27857 ( .A(n27701), .B(n27702), .Z(n27700) );
  OR U27858 ( .A(n27703), .B(n27704), .Z(n27702) );
  NAND U27859 ( .A(n27704), .B(n27703), .Z(n27699) );
  ANDN U27860 ( .B(B[182]), .A(n59), .Z(n27483) );
  XNOR U27861 ( .A(n27491), .B(n27705), .Z(n27484) );
  XNOR U27862 ( .A(n27490), .B(n27488), .Z(n27705) );
  AND U27863 ( .A(n27706), .B(n27707), .Z(n27488) );
  NANDN U27864 ( .A(n27708), .B(n27709), .Z(n27707) );
  NANDN U27865 ( .A(n27710), .B(n27711), .Z(n27709) );
  NANDN U27866 ( .A(n27711), .B(n27710), .Z(n27706) );
  ANDN U27867 ( .B(B[183]), .A(n60), .Z(n27490) );
  XNOR U27868 ( .A(n27498), .B(n27712), .Z(n27491) );
  XNOR U27869 ( .A(n27497), .B(n27495), .Z(n27712) );
  AND U27870 ( .A(n27713), .B(n27714), .Z(n27495) );
  NANDN U27871 ( .A(n27715), .B(n27716), .Z(n27714) );
  OR U27872 ( .A(n27717), .B(n27718), .Z(n27716) );
  NAND U27873 ( .A(n27718), .B(n27717), .Z(n27713) );
  ANDN U27874 ( .B(B[184]), .A(n61), .Z(n27497) );
  XNOR U27875 ( .A(n27505), .B(n27719), .Z(n27498) );
  XNOR U27876 ( .A(n27504), .B(n27502), .Z(n27719) );
  AND U27877 ( .A(n27720), .B(n27721), .Z(n27502) );
  NANDN U27878 ( .A(n27722), .B(n27723), .Z(n27721) );
  NANDN U27879 ( .A(n27724), .B(n27725), .Z(n27723) );
  NANDN U27880 ( .A(n27725), .B(n27724), .Z(n27720) );
  ANDN U27881 ( .B(B[185]), .A(n62), .Z(n27504) );
  XNOR U27882 ( .A(n27512), .B(n27726), .Z(n27505) );
  XNOR U27883 ( .A(n27511), .B(n27509), .Z(n27726) );
  AND U27884 ( .A(n27727), .B(n27728), .Z(n27509) );
  NANDN U27885 ( .A(n27729), .B(n27730), .Z(n27728) );
  OR U27886 ( .A(n27731), .B(n27732), .Z(n27730) );
  NAND U27887 ( .A(n27732), .B(n27731), .Z(n27727) );
  ANDN U27888 ( .B(B[186]), .A(n63), .Z(n27511) );
  XNOR U27889 ( .A(n27519), .B(n27733), .Z(n27512) );
  XNOR U27890 ( .A(n27518), .B(n27516), .Z(n27733) );
  AND U27891 ( .A(n27734), .B(n27735), .Z(n27516) );
  NANDN U27892 ( .A(n27736), .B(n27737), .Z(n27735) );
  NANDN U27893 ( .A(n27738), .B(n27739), .Z(n27737) );
  NANDN U27894 ( .A(n27739), .B(n27738), .Z(n27734) );
  ANDN U27895 ( .B(B[187]), .A(n64), .Z(n27518) );
  XNOR U27896 ( .A(n27526), .B(n27740), .Z(n27519) );
  XNOR U27897 ( .A(n27525), .B(n27523), .Z(n27740) );
  AND U27898 ( .A(n27741), .B(n27742), .Z(n27523) );
  NANDN U27899 ( .A(n27743), .B(n27744), .Z(n27742) );
  OR U27900 ( .A(n27745), .B(n27746), .Z(n27744) );
  NAND U27901 ( .A(n27746), .B(n27745), .Z(n27741) );
  ANDN U27902 ( .B(B[188]), .A(n65), .Z(n27525) );
  XNOR U27903 ( .A(n27533), .B(n27747), .Z(n27526) );
  XNOR U27904 ( .A(n27532), .B(n27530), .Z(n27747) );
  AND U27905 ( .A(n27748), .B(n27749), .Z(n27530) );
  NANDN U27906 ( .A(n27750), .B(n27751), .Z(n27749) );
  NANDN U27907 ( .A(n27752), .B(n27753), .Z(n27751) );
  NANDN U27908 ( .A(n27753), .B(n27752), .Z(n27748) );
  ANDN U27909 ( .B(B[189]), .A(n66), .Z(n27532) );
  XNOR U27910 ( .A(n27540), .B(n27754), .Z(n27533) );
  XNOR U27911 ( .A(n27539), .B(n27537), .Z(n27754) );
  AND U27912 ( .A(n27755), .B(n27756), .Z(n27537) );
  NANDN U27913 ( .A(n27757), .B(n27758), .Z(n27756) );
  OR U27914 ( .A(n27759), .B(n27760), .Z(n27758) );
  NAND U27915 ( .A(n27760), .B(n27759), .Z(n27755) );
  ANDN U27916 ( .B(B[190]), .A(n67), .Z(n27539) );
  XNOR U27917 ( .A(n27547), .B(n27761), .Z(n27540) );
  XNOR U27918 ( .A(n27546), .B(n27544), .Z(n27761) );
  AND U27919 ( .A(n27762), .B(n27763), .Z(n27544) );
  NANDN U27920 ( .A(n27764), .B(n27765), .Z(n27763) );
  NANDN U27921 ( .A(n27766), .B(n27767), .Z(n27765) );
  NANDN U27922 ( .A(n27767), .B(n27766), .Z(n27762) );
  ANDN U27923 ( .B(B[191]), .A(n68), .Z(n27546) );
  XNOR U27924 ( .A(n27554), .B(n27768), .Z(n27547) );
  XNOR U27925 ( .A(n27553), .B(n27551), .Z(n27768) );
  AND U27926 ( .A(n27769), .B(n27770), .Z(n27551) );
  NANDN U27927 ( .A(n27771), .B(n27772), .Z(n27770) );
  OR U27928 ( .A(n27773), .B(n27774), .Z(n27772) );
  NAND U27929 ( .A(n27774), .B(n27773), .Z(n27769) );
  ANDN U27930 ( .B(B[192]), .A(n69), .Z(n27553) );
  XNOR U27931 ( .A(n27561), .B(n27775), .Z(n27554) );
  XNOR U27932 ( .A(n27560), .B(n27558), .Z(n27775) );
  AND U27933 ( .A(n27776), .B(n27777), .Z(n27558) );
  NANDN U27934 ( .A(n27778), .B(n27779), .Z(n27777) );
  NANDN U27935 ( .A(n27780), .B(n27781), .Z(n27779) );
  NANDN U27936 ( .A(n27781), .B(n27780), .Z(n27776) );
  ANDN U27937 ( .B(B[193]), .A(n70), .Z(n27560) );
  XNOR U27938 ( .A(n27568), .B(n27782), .Z(n27561) );
  XNOR U27939 ( .A(n27567), .B(n27565), .Z(n27782) );
  AND U27940 ( .A(n27783), .B(n27784), .Z(n27565) );
  NANDN U27941 ( .A(n27785), .B(n27786), .Z(n27784) );
  OR U27942 ( .A(n27787), .B(n27788), .Z(n27786) );
  NAND U27943 ( .A(n27788), .B(n27787), .Z(n27783) );
  ANDN U27944 ( .B(B[194]), .A(n71), .Z(n27567) );
  XNOR U27945 ( .A(n27575), .B(n27789), .Z(n27568) );
  XNOR U27946 ( .A(n27574), .B(n27572), .Z(n27789) );
  AND U27947 ( .A(n27790), .B(n27791), .Z(n27572) );
  NANDN U27948 ( .A(n27792), .B(n27793), .Z(n27791) );
  NANDN U27949 ( .A(n27794), .B(n27795), .Z(n27793) );
  NANDN U27950 ( .A(n27795), .B(n27794), .Z(n27790) );
  ANDN U27951 ( .B(B[195]), .A(n72), .Z(n27574) );
  XNOR U27952 ( .A(n27582), .B(n27796), .Z(n27575) );
  XNOR U27953 ( .A(n27581), .B(n27579), .Z(n27796) );
  AND U27954 ( .A(n27797), .B(n27798), .Z(n27579) );
  NANDN U27955 ( .A(n27799), .B(n27800), .Z(n27798) );
  OR U27956 ( .A(n27801), .B(n27802), .Z(n27800) );
  NAND U27957 ( .A(n27802), .B(n27801), .Z(n27797) );
  ANDN U27958 ( .B(B[196]), .A(n73), .Z(n27581) );
  XNOR U27959 ( .A(n27589), .B(n27803), .Z(n27582) );
  XNOR U27960 ( .A(n27588), .B(n27586), .Z(n27803) );
  AND U27961 ( .A(n27804), .B(n27805), .Z(n27586) );
  NANDN U27962 ( .A(n27806), .B(n27807), .Z(n27805) );
  NANDN U27963 ( .A(n27808), .B(n27809), .Z(n27807) );
  NANDN U27964 ( .A(n27809), .B(n27808), .Z(n27804) );
  ANDN U27965 ( .B(B[197]), .A(n74), .Z(n27588) );
  XNOR U27966 ( .A(n27596), .B(n27810), .Z(n27589) );
  XNOR U27967 ( .A(n27595), .B(n27593), .Z(n27810) );
  AND U27968 ( .A(n27811), .B(n27812), .Z(n27593) );
  NANDN U27969 ( .A(n27813), .B(n27814), .Z(n27812) );
  OR U27970 ( .A(n27815), .B(n27816), .Z(n27814) );
  NAND U27971 ( .A(n27816), .B(n27815), .Z(n27811) );
  ANDN U27972 ( .B(B[198]), .A(n75), .Z(n27595) );
  XNOR U27973 ( .A(n27603), .B(n27817), .Z(n27596) );
  XNOR U27974 ( .A(n27602), .B(n27600), .Z(n27817) );
  AND U27975 ( .A(n27818), .B(n27819), .Z(n27600) );
  NANDN U27976 ( .A(n27820), .B(n27821), .Z(n27819) );
  NANDN U27977 ( .A(n27822), .B(n27823), .Z(n27821) );
  NANDN U27978 ( .A(n27823), .B(n27822), .Z(n27818) );
  ANDN U27979 ( .B(B[199]), .A(n76), .Z(n27602) );
  XNOR U27980 ( .A(n27610), .B(n27824), .Z(n27603) );
  XNOR U27981 ( .A(n27609), .B(n27607), .Z(n27824) );
  AND U27982 ( .A(n27825), .B(n27826), .Z(n27607) );
  NANDN U27983 ( .A(n27827), .B(n27828), .Z(n27826) );
  OR U27984 ( .A(n27829), .B(n27830), .Z(n27828) );
  NAND U27985 ( .A(n27830), .B(n27829), .Z(n27825) );
  ANDN U27986 ( .B(B[200]), .A(n77), .Z(n27609) );
  XNOR U27987 ( .A(n27617), .B(n27831), .Z(n27610) );
  XNOR U27988 ( .A(n27616), .B(n27614), .Z(n27831) );
  AND U27989 ( .A(n27832), .B(n27833), .Z(n27614) );
  NANDN U27990 ( .A(n27834), .B(n27835), .Z(n27833) );
  NANDN U27991 ( .A(n27836), .B(n27837), .Z(n27835) );
  NANDN U27992 ( .A(n27837), .B(n27836), .Z(n27832) );
  ANDN U27993 ( .B(B[201]), .A(n78), .Z(n27616) );
  XNOR U27994 ( .A(n27624), .B(n27838), .Z(n27617) );
  XNOR U27995 ( .A(n27623), .B(n27621), .Z(n27838) );
  AND U27996 ( .A(n27839), .B(n27840), .Z(n27621) );
  NANDN U27997 ( .A(n27841), .B(n27842), .Z(n27840) );
  OR U27998 ( .A(n27843), .B(n27844), .Z(n27842) );
  NAND U27999 ( .A(n27844), .B(n27843), .Z(n27839) );
  ANDN U28000 ( .B(B[202]), .A(n79), .Z(n27623) );
  XNOR U28001 ( .A(n27631), .B(n27845), .Z(n27624) );
  XNOR U28002 ( .A(n27630), .B(n27628), .Z(n27845) );
  AND U28003 ( .A(n27846), .B(n27847), .Z(n27628) );
  NANDN U28004 ( .A(n27848), .B(n27849), .Z(n27847) );
  NANDN U28005 ( .A(n27850), .B(n27851), .Z(n27849) );
  NANDN U28006 ( .A(n27851), .B(n27850), .Z(n27846) );
  ANDN U28007 ( .B(B[203]), .A(n80), .Z(n27630) );
  XNOR U28008 ( .A(n27638), .B(n27852), .Z(n27631) );
  XNOR U28009 ( .A(n27637), .B(n27635), .Z(n27852) );
  AND U28010 ( .A(n27853), .B(n27854), .Z(n27635) );
  NANDN U28011 ( .A(n27855), .B(n27856), .Z(n27854) );
  OR U28012 ( .A(n27857), .B(n27858), .Z(n27856) );
  NAND U28013 ( .A(n27858), .B(n27857), .Z(n27853) );
  ANDN U28014 ( .B(B[204]), .A(n81), .Z(n27637) );
  XNOR U28015 ( .A(n27645), .B(n27859), .Z(n27638) );
  XNOR U28016 ( .A(n27644), .B(n27642), .Z(n27859) );
  AND U28017 ( .A(n27860), .B(n27861), .Z(n27642) );
  NANDN U28018 ( .A(n27862), .B(n27863), .Z(n27861) );
  NAND U28019 ( .A(n27864), .B(n27865), .Z(n27863) );
  ANDN U28020 ( .B(B[205]), .A(n82), .Z(n27644) );
  XOR U28021 ( .A(n27651), .B(n27866), .Z(n27645) );
  XNOR U28022 ( .A(n27649), .B(n27652), .Z(n27866) );
  NAND U28023 ( .A(A[2]), .B(B[206]), .Z(n27652) );
  NANDN U28024 ( .A(n27867), .B(n27868), .Z(n27649) );
  AND U28025 ( .A(A[0]), .B(B[207]), .Z(n27868) );
  XNOR U28026 ( .A(n27654), .B(n27869), .Z(n27651) );
  NAND U28027 ( .A(A[0]), .B(B[208]), .Z(n27869) );
  NAND U28028 ( .A(B[207]), .B(A[1]), .Z(n27654) );
  NAND U28029 ( .A(n27870), .B(n27871), .Z(n380) );
  NANDN U28030 ( .A(n27872), .B(n27873), .Z(n27871) );
  OR U28031 ( .A(n27874), .B(n27875), .Z(n27873) );
  NAND U28032 ( .A(n27875), .B(n27874), .Z(n27870) );
  XOR U28033 ( .A(n382), .B(n381), .Z(\A1[205] ) );
  XOR U28034 ( .A(n27875), .B(n27876), .Z(n381) );
  XNOR U28035 ( .A(n27874), .B(n27872), .Z(n27876) );
  AND U28036 ( .A(n27877), .B(n27878), .Z(n27872) );
  NANDN U28037 ( .A(n27879), .B(n27880), .Z(n27878) );
  NANDN U28038 ( .A(n27881), .B(n27882), .Z(n27880) );
  NANDN U28039 ( .A(n27882), .B(n27881), .Z(n27877) );
  ANDN U28040 ( .B(B[176]), .A(n54), .Z(n27874) );
  XNOR U28041 ( .A(n27669), .B(n27883), .Z(n27875) );
  XNOR U28042 ( .A(n27668), .B(n27666), .Z(n27883) );
  AND U28043 ( .A(n27884), .B(n27885), .Z(n27666) );
  NANDN U28044 ( .A(n27886), .B(n27887), .Z(n27885) );
  OR U28045 ( .A(n27888), .B(n27889), .Z(n27887) );
  NAND U28046 ( .A(n27889), .B(n27888), .Z(n27884) );
  ANDN U28047 ( .B(B[177]), .A(n55), .Z(n27668) );
  XNOR U28048 ( .A(n27676), .B(n27890), .Z(n27669) );
  XNOR U28049 ( .A(n27675), .B(n27673), .Z(n27890) );
  AND U28050 ( .A(n27891), .B(n27892), .Z(n27673) );
  NANDN U28051 ( .A(n27893), .B(n27894), .Z(n27892) );
  NANDN U28052 ( .A(n27895), .B(n27896), .Z(n27894) );
  NANDN U28053 ( .A(n27896), .B(n27895), .Z(n27891) );
  ANDN U28054 ( .B(B[178]), .A(n56), .Z(n27675) );
  XNOR U28055 ( .A(n27683), .B(n27897), .Z(n27676) );
  XNOR U28056 ( .A(n27682), .B(n27680), .Z(n27897) );
  AND U28057 ( .A(n27898), .B(n27899), .Z(n27680) );
  NANDN U28058 ( .A(n27900), .B(n27901), .Z(n27899) );
  OR U28059 ( .A(n27902), .B(n27903), .Z(n27901) );
  NAND U28060 ( .A(n27903), .B(n27902), .Z(n27898) );
  ANDN U28061 ( .B(B[179]), .A(n57), .Z(n27682) );
  XNOR U28062 ( .A(n27690), .B(n27904), .Z(n27683) );
  XNOR U28063 ( .A(n27689), .B(n27687), .Z(n27904) );
  AND U28064 ( .A(n27905), .B(n27906), .Z(n27687) );
  NANDN U28065 ( .A(n27907), .B(n27908), .Z(n27906) );
  NANDN U28066 ( .A(n27909), .B(n27910), .Z(n27908) );
  NANDN U28067 ( .A(n27910), .B(n27909), .Z(n27905) );
  ANDN U28068 ( .B(B[180]), .A(n58), .Z(n27689) );
  XNOR U28069 ( .A(n27697), .B(n27911), .Z(n27690) );
  XNOR U28070 ( .A(n27696), .B(n27694), .Z(n27911) );
  AND U28071 ( .A(n27912), .B(n27913), .Z(n27694) );
  NANDN U28072 ( .A(n27914), .B(n27915), .Z(n27913) );
  OR U28073 ( .A(n27916), .B(n27917), .Z(n27915) );
  NAND U28074 ( .A(n27917), .B(n27916), .Z(n27912) );
  ANDN U28075 ( .B(B[181]), .A(n59), .Z(n27696) );
  XNOR U28076 ( .A(n27704), .B(n27918), .Z(n27697) );
  XNOR U28077 ( .A(n27703), .B(n27701), .Z(n27918) );
  AND U28078 ( .A(n27919), .B(n27920), .Z(n27701) );
  NANDN U28079 ( .A(n27921), .B(n27922), .Z(n27920) );
  NANDN U28080 ( .A(n27923), .B(n27924), .Z(n27922) );
  NANDN U28081 ( .A(n27924), .B(n27923), .Z(n27919) );
  ANDN U28082 ( .B(B[182]), .A(n60), .Z(n27703) );
  XNOR U28083 ( .A(n27711), .B(n27925), .Z(n27704) );
  XNOR U28084 ( .A(n27710), .B(n27708), .Z(n27925) );
  AND U28085 ( .A(n27926), .B(n27927), .Z(n27708) );
  NANDN U28086 ( .A(n27928), .B(n27929), .Z(n27927) );
  OR U28087 ( .A(n27930), .B(n27931), .Z(n27929) );
  NAND U28088 ( .A(n27931), .B(n27930), .Z(n27926) );
  ANDN U28089 ( .B(B[183]), .A(n61), .Z(n27710) );
  XNOR U28090 ( .A(n27718), .B(n27932), .Z(n27711) );
  XNOR U28091 ( .A(n27717), .B(n27715), .Z(n27932) );
  AND U28092 ( .A(n27933), .B(n27934), .Z(n27715) );
  NANDN U28093 ( .A(n27935), .B(n27936), .Z(n27934) );
  NANDN U28094 ( .A(n27937), .B(n27938), .Z(n27936) );
  NANDN U28095 ( .A(n27938), .B(n27937), .Z(n27933) );
  ANDN U28096 ( .B(B[184]), .A(n62), .Z(n27717) );
  XNOR U28097 ( .A(n27725), .B(n27939), .Z(n27718) );
  XNOR U28098 ( .A(n27724), .B(n27722), .Z(n27939) );
  AND U28099 ( .A(n27940), .B(n27941), .Z(n27722) );
  NANDN U28100 ( .A(n27942), .B(n27943), .Z(n27941) );
  OR U28101 ( .A(n27944), .B(n27945), .Z(n27943) );
  NAND U28102 ( .A(n27945), .B(n27944), .Z(n27940) );
  ANDN U28103 ( .B(B[185]), .A(n63), .Z(n27724) );
  XNOR U28104 ( .A(n27732), .B(n27946), .Z(n27725) );
  XNOR U28105 ( .A(n27731), .B(n27729), .Z(n27946) );
  AND U28106 ( .A(n27947), .B(n27948), .Z(n27729) );
  NANDN U28107 ( .A(n27949), .B(n27950), .Z(n27948) );
  NANDN U28108 ( .A(n27951), .B(n27952), .Z(n27950) );
  NANDN U28109 ( .A(n27952), .B(n27951), .Z(n27947) );
  ANDN U28110 ( .B(B[186]), .A(n64), .Z(n27731) );
  XNOR U28111 ( .A(n27739), .B(n27953), .Z(n27732) );
  XNOR U28112 ( .A(n27738), .B(n27736), .Z(n27953) );
  AND U28113 ( .A(n27954), .B(n27955), .Z(n27736) );
  NANDN U28114 ( .A(n27956), .B(n27957), .Z(n27955) );
  OR U28115 ( .A(n27958), .B(n27959), .Z(n27957) );
  NAND U28116 ( .A(n27959), .B(n27958), .Z(n27954) );
  ANDN U28117 ( .B(B[187]), .A(n65), .Z(n27738) );
  XNOR U28118 ( .A(n27746), .B(n27960), .Z(n27739) );
  XNOR U28119 ( .A(n27745), .B(n27743), .Z(n27960) );
  AND U28120 ( .A(n27961), .B(n27962), .Z(n27743) );
  NANDN U28121 ( .A(n27963), .B(n27964), .Z(n27962) );
  NANDN U28122 ( .A(n27965), .B(n27966), .Z(n27964) );
  NANDN U28123 ( .A(n27966), .B(n27965), .Z(n27961) );
  ANDN U28124 ( .B(B[188]), .A(n66), .Z(n27745) );
  XNOR U28125 ( .A(n27753), .B(n27967), .Z(n27746) );
  XNOR U28126 ( .A(n27752), .B(n27750), .Z(n27967) );
  AND U28127 ( .A(n27968), .B(n27969), .Z(n27750) );
  NANDN U28128 ( .A(n27970), .B(n27971), .Z(n27969) );
  OR U28129 ( .A(n27972), .B(n27973), .Z(n27971) );
  NAND U28130 ( .A(n27973), .B(n27972), .Z(n27968) );
  ANDN U28131 ( .B(B[189]), .A(n67), .Z(n27752) );
  XNOR U28132 ( .A(n27760), .B(n27974), .Z(n27753) );
  XNOR U28133 ( .A(n27759), .B(n27757), .Z(n27974) );
  AND U28134 ( .A(n27975), .B(n27976), .Z(n27757) );
  NANDN U28135 ( .A(n27977), .B(n27978), .Z(n27976) );
  NANDN U28136 ( .A(n27979), .B(n27980), .Z(n27978) );
  NANDN U28137 ( .A(n27980), .B(n27979), .Z(n27975) );
  ANDN U28138 ( .B(B[190]), .A(n68), .Z(n27759) );
  XNOR U28139 ( .A(n27767), .B(n27981), .Z(n27760) );
  XNOR U28140 ( .A(n27766), .B(n27764), .Z(n27981) );
  AND U28141 ( .A(n27982), .B(n27983), .Z(n27764) );
  NANDN U28142 ( .A(n27984), .B(n27985), .Z(n27983) );
  OR U28143 ( .A(n27986), .B(n27987), .Z(n27985) );
  NAND U28144 ( .A(n27987), .B(n27986), .Z(n27982) );
  ANDN U28145 ( .B(B[191]), .A(n69), .Z(n27766) );
  XNOR U28146 ( .A(n27774), .B(n27988), .Z(n27767) );
  XNOR U28147 ( .A(n27773), .B(n27771), .Z(n27988) );
  AND U28148 ( .A(n27989), .B(n27990), .Z(n27771) );
  NANDN U28149 ( .A(n27991), .B(n27992), .Z(n27990) );
  NANDN U28150 ( .A(n27993), .B(n27994), .Z(n27992) );
  NANDN U28151 ( .A(n27994), .B(n27993), .Z(n27989) );
  ANDN U28152 ( .B(B[192]), .A(n70), .Z(n27773) );
  XNOR U28153 ( .A(n27781), .B(n27995), .Z(n27774) );
  XNOR U28154 ( .A(n27780), .B(n27778), .Z(n27995) );
  AND U28155 ( .A(n27996), .B(n27997), .Z(n27778) );
  NANDN U28156 ( .A(n27998), .B(n27999), .Z(n27997) );
  OR U28157 ( .A(n28000), .B(n28001), .Z(n27999) );
  NAND U28158 ( .A(n28001), .B(n28000), .Z(n27996) );
  ANDN U28159 ( .B(B[193]), .A(n71), .Z(n27780) );
  XNOR U28160 ( .A(n27788), .B(n28002), .Z(n27781) );
  XNOR U28161 ( .A(n27787), .B(n27785), .Z(n28002) );
  AND U28162 ( .A(n28003), .B(n28004), .Z(n27785) );
  NANDN U28163 ( .A(n28005), .B(n28006), .Z(n28004) );
  NANDN U28164 ( .A(n28007), .B(n28008), .Z(n28006) );
  NANDN U28165 ( .A(n28008), .B(n28007), .Z(n28003) );
  ANDN U28166 ( .B(B[194]), .A(n72), .Z(n27787) );
  XNOR U28167 ( .A(n27795), .B(n28009), .Z(n27788) );
  XNOR U28168 ( .A(n27794), .B(n27792), .Z(n28009) );
  AND U28169 ( .A(n28010), .B(n28011), .Z(n27792) );
  NANDN U28170 ( .A(n28012), .B(n28013), .Z(n28011) );
  OR U28171 ( .A(n28014), .B(n28015), .Z(n28013) );
  NAND U28172 ( .A(n28015), .B(n28014), .Z(n28010) );
  ANDN U28173 ( .B(B[195]), .A(n73), .Z(n27794) );
  XNOR U28174 ( .A(n27802), .B(n28016), .Z(n27795) );
  XNOR U28175 ( .A(n27801), .B(n27799), .Z(n28016) );
  AND U28176 ( .A(n28017), .B(n28018), .Z(n27799) );
  NANDN U28177 ( .A(n28019), .B(n28020), .Z(n28018) );
  NANDN U28178 ( .A(n28021), .B(n28022), .Z(n28020) );
  NANDN U28179 ( .A(n28022), .B(n28021), .Z(n28017) );
  ANDN U28180 ( .B(B[196]), .A(n74), .Z(n27801) );
  XNOR U28181 ( .A(n27809), .B(n28023), .Z(n27802) );
  XNOR U28182 ( .A(n27808), .B(n27806), .Z(n28023) );
  AND U28183 ( .A(n28024), .B(n28025), .Z(n27806) );
  NANDN U28184 ( .A(n28026), .B(n28027), .Z(n28025) );
  OR U28185 ( .A(n28028), .B(n28029), .Z(n28027) );
  NAND U28186 ( .A(n28029), .B(n28028), .Z(n28024) );
  ANDN U28187 ( .B(B[197]), .A(n75), .Z(n27808) );
  XNOR U28188 ( .A(n27816), .B(n28030), .Z(n27809) );
  XNOR U28189 ( .A(n27815), .B(n27813), .Z(n28030) );
  AND U28190 ( .A(n28031), .B(n28032), .Z(n27813) );
  NANDN U28191 ( .A(n28033), .B(n28034), .Z(n28032) );
  NANDN U28192 ( .A(n28035), .B(n28036), .Z(n28034) );
  NANDN U28193 ( .A(n28036), .B(n28035), .Z(n28031) );
  ANDN U28194 ( .B(B[198]), .A(n76), .Z(n27815) );
  XNOR U28195 ( .A(n27823), .B(n28037), .Z(n27816) );
  XNOR U28196 ( .A(n27822), .B(n27820), .Z(n28037) );
  AND U28197 ( .A(n28038), .B(n28039), .Z(n27820) );
  NANDN U28198 ( .A(n28040), .B(n28041), .Z(n28039) );
  OR U28199 ( .A(n28042), .B(n28043), .Z(n28041) );
  NAND U28200 ( .A(n28043), .B(n28042), .Z(n28038) );
  ANDN U28201 ( .B(B[199]), .A(n77), .Z(n27822) );
  XNOR U28202 ( .A(n27830), .B(n28044), .Z(n27823) );
  XNOR U28203 ( .A(n27829), .B(n27827), .Z(n28044) );
  AND U28204 ( .A(n28045), .B(n28046), .Z(n27827) );
  NANDN U28205 ( .A(n28047), .B(n28048), .Z(n28046) );
  NANDN U28206 ( .A(n28049), .B(n28050), .Z(n28048) );
  NANDN U28207 ( .A(n28050), .B(n28049), .Z(n28045) );
  ANDN U28208 ( .B(B[200]), .A(n78), .Z(n27829) );
  XNOR U28209 ( .A(n27837), .B(n28051), .Z(n27830) );
  XNOR U28210 ( .A(n27836), .B(n27834), .Z(n28051) );
  AND U28211 ( .A(n28052), .B(n28053), .Z(n27834) );
  NANDN U28212 ( .A(n28054), .B(n28055), .Z(n28053) );
  OR U28213 ( .A(n28056), .B(n28057), .Z(n28055) );
  NAND U28214 ( .A(n28057), .B(n28056), .Z(n28052) );
  ANDN U28215 ( .B(B[201]), .A(n79), .Z(n27836) );
  XNOR U28216 ( .A(n27844), .B(n28058), .Z(n27837) );
  XNOR U28217 ( .A(n27843), .B(n27841), .Z(n28058) );
  AND U28218 ( .A(n28059), .B(n28060), .Z(n27841) );
  NANDN U28219 ( .A(n28061), .B(n28062), .Z(n28060) );
  NANDN U28220 ( .A(n28063), .B(n28064), .Z(n28062) );
  NANDN U28221 ( .A(n28064), .B(n28063), .Z(n28059) );
  ANDN U28222 ( .B(B[202]), .A(n80), .Z(n27843) );
  XNOR U28223 ( .A(n27851), .B(n28065), .Z(n27844) );
  XNOR U28224 ( .A(n27850), .B(n27848), .Z(n28065) );
  AND U28225 ( .A(n28066), .B(n28067), .Z(n27848) );
  NANDN U28226 ( .A(n28068), .B(n28069), .Z(n28067) );
  OR U28227 ( .A(n28070), .B(n28071), .Z(n28069) );
  NAND U28228 ( .A(n28071), .B(n28070), .Z(n28066) );
  ANDN U28229 ( .B(B[203]), .A(n81), .Z(n27850) );
  XNOR U28230 ( .A(n27858), .B(n28072), .Z(n27851) );
  XNOR U28231 ( .A(n27857), .B(n27855), .Z(n28072) );
  AND U28232 ( .A(n28073), .B(n28074), .Z(n27855) );
  NANDN U28233 ( .A(n28075), .B(n28076), .Z(n28074) );
  NAND U28234 ( .A(n28077), .B(n28078), .Z(n28076) );
  ANDN U28235 ( .B(B[204]), .A(n82), .Z(n27857) );
  XOR U28236 ( .A(n27864), .B(n28079), .Z(n27858) );
  XNOR U28237 ( .A(n27862), .B(n27865), .Z(n28079) );
  NAND U28238 ( .A(A[2]), .B(B[205]), .Z(n27865) );
  NANDN U28239 ( .A(n28080), .B(n28081), .Z(n27862) );
  AND U28240 ( .A(A[0]), .B(B[206]), .Z(n28081) );
  XNOR U28241 ( .A(n27867), .B(n28082), .Z(n27864) );
  NAND U28242 ( .A(A[0]), .B(B[207]), .Z(n28082) );
  NAND U28243 ( .A(B[206]), .B(A[1]), .Z(n27867) );
  NAND U28244 ( .A(n28083), .B(n28084), .Z(n382) );
  NANDN U28245 ( .A(n28085), .B(n28086), .Z(n28084) );
  OR U28246 ( .A(n28087), .B(n28088), .Z(n28086) );
  NAND U28247 ( .A(n28088), .B(n28087), .Z(n28083) );
  XOR U28248 ( .A(n384), .B(n383), .Z(\A1[204] ) );
  XOR U28249 ( .A(n28088), .B(n28089), .Z(n383) );
  XNOR U28250 ( .A(n28087), .B(n28085), .Z(n28089) );
  AND U28251 ( .A(n28090), .B(n28091), .Z(n28085) );
  NANDN U28252 ( .A(n28092), .B(n28093), .Z(n28091) );
  NANDN U28253 ( .A(n28094), .B(n28095), .Z(n28093) );
  NANDN U28254 ( .A(n28095), .B(n28094), .Z(n28090) );
  ANDN U28255 ( .B(B[175]), .A(n54), .Z(n28087) );
  XNOR U28256 ( .A(n27882), .B(n28096), .Z(n28088) );
  XNOR U28257 ( .A(n27881), .B(n27879), .Z(n28096) );
  AND U28258 ( .A(n28097), .B(n28098), .Z(n27879) );
  NANDN U28259 ( .A(n28099), .B(n28100), .Z(n28098) );
  OR U28260 ( .A(n28101), .B(n28102), .Z(n28100) );
  NAND U28261 ( .A(n28102), .B(n28101), .Z(n28097) );
  ANDN U28262 ( .B(B[176]), .A(n55), .Z(n27881) );
  XNOR U28263 ( .A(n27889), .B(n28103), .Z(n27882) );
  XNOR U28264 ( .A(n27888), .B(n27886), .Z(n28103) );
  AND U28265 ( .A(n28104), .B(n28105), .Z(n27886) );
  NANDN U28266 ( .A(n28106), .B(n28107), .Z(n28105) );
  NANDN U28267 ( .A(n28108), .B(n28109), .Z(n28107) );
  NANDN U28268 ( .A(n28109), .B(n28108), .Z(n28104) );
  ANDN U28269 ( .B(B[177]), .A(n56), .Z(n27888) );
  XNOR U28270 ( .A(n27896), .B(n28110), .Z(n27889) );
  XNOR U28271 ( .A(n27895), .B(n27893), .Z(n28110) );
  AND U28272 ( .A(n28111), .B(n28112), .Z(n27893) );
  NANDN U28273 ( .A(n28113), .B(n28114), .Z(n28112) );
  OR U28274 ( .A(n28115), .B(n28116), .Z(n28114) );
  NAND U28275 ( .A(n28116), .B(n28115), .Z(n28111) );
  ANDN U28276 ( .B(B[178]), .A(n57), .Z(n27895) );
  XNOR U28277 ( .A(n27903), .B(n28117), .Z(n27896) );
  XNOR U28278 ( .A(n27902), .B(n27900), .Z(n28117) );
  AND U28279 ( .A(n28118), .B(n28119), .Z(n27900) );
  NANDN U28280 ( .A(n28120), .B(n28121), .Z(n28119) );
  NANDN U28281 ( .A(n28122), .B(n28123), .Z(n28121) );
  NANDN U28282 ( .A(n28123), .B(n28122), .Z(n28118) );
  ANDN U28283 ( .B(B[179]), .A(n58), .Z(n27902) );
  XNOR U28284 ( .A(n27910), .B(n28124), .Z(n27903) );
  XNOR U28285 ( .A(n27909), .B(n27907), .Z(n28124) );
  AND U28286 ( .A(n28125), .B(n28126), .Z(n27907) );
  NANDN U28287 ( .A(n28127), .B(n28128), .Z(n28126) );
  OR U28288 ( .A(n28129), .B(n28130), .Z(n28128) );
  NAND U28289 ( .A(n28130), .B(n28129), .Z(n28125) );
  ANDN U28290 ( .B(B[180]), .A(n59), .Z(n27909) );
  XNOR U28291 ( .A(n27917), .B(n28131), .Z(n27910) );
  XNOR U28292 ( .A(n27916), .B(n27914), .Z(n28131) );
  AND U28293 ( .A(n28132), .B(n28133), .Z(n27914) );
  NANDN U28294 ( .A(n28134), .B(n28135), .Z(n28133) );
  NANDN U28295 ( .A(n28136), .B(n28137), .Z(n28135) );
  NANDN U28296 ( .A(n28137), .B(n28136), .Z(n28132) );
  ANDN U28297 ( .B(B[181]), .A(n60), .Z(n27916) );
  XNOR U28298 ( .A(n27924), .B(n28138), .Z(n27917) );
  XNOR U28299 ( .A(n27923), .B(n27921), .Z(n28138) );
  AND U28300 ( .A(n28139), .B(n28140), .Z(n27921) );
  NANDN U28301 ( .A(n28141), .B(n28142), .Z(n28140) );
  OR U28302 ( .A(n28143), .B(n28144), .Z(n28142) );
  NAND U28303 ( .A(n28144), .B(n28143), .Z(n28139) );
  ANDN U28304 ( .B(B[182]), .A(n61), .Z(n27923) );
  XNOR U28305 ( .A(n27931), .B(n28145), .Z(n27924) );
  XNOR U28306 ( .A(n27930), .B(n27928), .Z(n28145) );
  AND U28307 ( .A(n28146), .B(n28147), .Z(n27928) );
  NANDN U28308 ( .A(n28148), .B(n28149), .Z(n28147) );
  NANDN U28309 ( .A(n28150), .B(n28151), .Z(n28149) );
  NANDN U28310 ( .A(n28151), .B(n28150), .Z(n28146) );
  ANDN U28311 ( .B(B[183]), .A(n62), .Z(n27930) );
  XNOR U28312 ( .A(n27938), .B(n28152), .Z(n27931) );
  XNOR U28313 ( .A(n27937), .B(n27935), .Z(n28152) );
  AND U28314 ( .A(n28153), .B(n28154), .Z(n27935) );
  NANDN U28315 ( .A(n28155), .B(n28156), .Z(n28154) );
  OR U28316 ( .A(n28157), .B(n28158), .Z(n28156) );
  NAND U28317 ( .A(n28158), .B(n28157), .Z(n28153) );
  ANDN U28318 ( .B(B[184]), .A(n63), .Z(n27937) );
  XNOR U28319 ( .A(n27945), .B(n28159), .Z(n27938) );
  XNOR U28320 ( .A(n27944), .B(n27942), .Z(n28159) );
  AND U28321 ( .A(n28160), .B(n28161), .Z(n27942) );
  NANDN U28322 ( .A(n28162), .B(n28163), .Z(n28161) );
  NANDN U28323 ( .A(n28164), .B(n28165), .Z(n28163) );
  NANDN U28324 ( .A(n28165), .B(n28164), .Z(n28160) );
  ANDN U28325 ( .B(B[185]), .A(n64), .Z(n27944) );
  XNOR U28326 ( .A(n27952), .B(n28166), .Z(n27945) );
  XNOR U28327 ( .A(n27951), .B(n27949), .Z(n28166) );
  AND U28328 ( .A(n28167), .B(n28168), .Z(n27949) );
  NANDN U28329 ( .A(n28169), .B(n28170), .Z(n28168) );
  OR U28330 ( .A(n28171), .B(n28172), .Z(n28170) );
  NAND U28331 ( .A(n28172), .B(n28171), .Z(n28167) );
  ANDN U28332 ( .B(B[186]), .A(n65), .Z(n27951) );
  XNOR U28333 ( .A(n27959), .B(n28173), .Z(n27952) );
  XNOR U28334 ( .A(n27958), .B(n27956), .Z(n28173) );
  AND U28335 ( .A(n28174), .B(n28175), .Z(n27956) );
  NANDN U28336 ( .A(n28176), .B(n28177), .Z(n28175) );
  NANDN U28337 ( .A(n28178), .B(n28179), .Z(n28177) );
  NANDN U28338 ( .A(n28179), .B(n28178), .Z(n28174) );
  ANDN U28339 ( .B(B[187]), .A(n66), .Z(n27958) );
  XNOR U28340 ( .A(n27966), .B(n28180), .Z(n27959) );
  XNOR U28341 ( .A(n27965), .B(n27963), .Z(n28180) );
  AND U28342 ( .A(n28181), .B(n28182), .Z(n27963) );
  NANDN U28343 ( .A(n28183), .B(n28184), .Z(n28182) );
  OR U28344 ( .A(n28185), .B(n28186), .Z(n28184) );
  NAND U28345 ( .A(n28186), .B(n28185), .Z(n28181) );
  ANDN U28346 ( .B(B[188]), .A(n67), .Z(n27965) );
  XNOR U28347 ( .A(n27973), .B(n28187), .Z(n27966) );
  XNOR U28348 ( .A(n27972), .B(n27970), .Z(n28187) );
  AND U28349 ( .A(n28188), .B(n28189), .Z(n27970) );
  NANDN U28350 ( .A(n28190), .B(n28191), .Z(n28189) );
  NANDN U28351 ( .A(n28192), .B(n28193), .Z(n28191) );
  NANDN U28352 ( .A(n28193), .B(n28192), .Z(n28188) );
  ANDN U28353 ( .B(B[189]), .A(n68), .Z(n27972) );
  XNOR U28354 ( .A(n27980), .B(n28194), .Z(n27973) );
  XNOR U28355 ( .A(n27979), .B(n27977), .Z(n28194) );
  AND U28356 ( .A(n28195), .B(n28196), .Z(n27977) );
  NANDN U28357 ( .A(n28197), .B(n28198), .Z(n28196) );
  OR U28358 ( .A(n28199), .B(n28200), .Z(n28198) );
  NAND U28359 ( .A(n28200), .B(n28199), .Z(n28195) );
  ANDN U28360 ( .B(B[190]), .A(n69), .Z(n27979) );
  XNOR U28361 ( .A(n27987), .B(n28201), .Z(n27980) );
  XNOR U28362 ( .A(n27986), .B(n27984), .Z(n28201) );
  AND U28363 ( .A(n28202), .B(n28203), .Z(n27984) );
  NANDN U28364 ( .A(n28204), .B(n28205), .Z(n28203) );
  NANDN U28365 ( .A(n28206), .B(n28207), .Z(n28205) );
  NANDN U28366 ( .A(n28207), .B(n28206), .Z(n28202) );
  ANDN U28367 ( .B(B[191]), .A(n70), .Z(n27986) );
  XNOR U28368 ( .A(n27994), .B(n28208), .Z(n27987) );
  XNOR U28369 ( .A(n27993), .B(n27991), .Z(n28208) );
  AND U28370 ( .A(n28209), .B(n28210), .Z(n27991) );
  NANDN U28371 ( .A(n28211), .B(n28212), .Z(n28210) );
  OR U28372 ( .A(n28213), .B(n28214), .Z(n28212) );
  NAND U28373 ( .A(n28214), .B(n28213), .Z(n28209) );
  ANDN U28374 ( .B(B[192]), .A(n71), .Z(n27993) );
  XNOR U28375 ( .A(n28001), .B(n28215), .Z(n27994) );
  XNOR U28376 ( .A(n28000), .B(n27998), .Z(n28215) );
  AND U28377 ( .A(n28216), .B(n28217), .Z(n27998) );
  NANDN U28378 ( .A(n28218), .B(n28219), .Z(n28217) );
  NANDN U28379 ( .A(n28220), .B(n28221), .Z(n28219) );
  NANDN U28380 ( .A(n28221), .B(n28220), .Z(n28216) );
  ANDN U28381 ( .B(B[193]), .A(n72), .Z(n28000) );
  XNOR U28382 ( .A(n28008), .B(n28222), .Z(n28001) );
  XNOR U28383 ( .A(n28007), .B(n28005), .Z(n28222) );
  AND U28384 ( .A(n28223), .B(n28224), .Z(n28005) );
  NANDN U28385 ( .A(n28225), .B(n28226), .Z(n28224) );
  OR U28386 ( .A(n28227), .B(n28228), .Z(n28226) );
  NAND U28387 ( .A(n28228), .B(n28227), .Z(n28223) );
  ANDN U28388 ( .B(B[194]), .A(n73), .Z(n28007) );
  XNOR U28389 ( .A(n28015), .B(n28229), .Z(n28008) );
  XNOR U28390 ( .A(n28014), .B(n28012), .Z(n28229) );
  AND U28391 ( .A(n28230), .B(n28231), .Z(n28012) );
  NANDN U28392 ( .A(n28232), .B(n28233), .Z(n28231) );
  NANDN U28393 ( .A(n28234), .B(n28235), .Z(n28233) );
  NANDN U28394 ( .A(n28235), .B(n28234), .Z(n28230) );
  ANDN U28395 ( .B(B[195]), .A(n74), .Z(n28014) );
  XNOR U28396 ( .A(n28022), .B(n28236), .Z(n28015) );
  XNOR U28397 ( .A(n28021), .B(n28019), .Z(n28236) );
  AND U28398 ( .A(n28237), .B(n28238), .Z(n28019) );
  NANDN U28399 ( .A(n28239), .B(n28240), .Z(n28238) );
  OR U28400 ( .A(n28241), .B(n28242), .Z(n28240) );
  NAND U28401 ( .A(n28242), .B(n28241), .Z(n28237) );
  ANDN U28402 ( .B(B[196]), .A(n75), .Z(n28021) );
  XNOR U28403 ( .A(n28029), .B(n28243), .Z(n28022) );
  XNOR U28404 ( .A(n28028), .B(n28026), .Z(n28243) );
  AND U28405 ( .A(n28244), .B(n28245), .Z(n28026) );
  NANDN U28406 ( .A(n28246), .B(n28247), .Z(n28245) );
  NANDN U28407 ( .A(n28248), .B(n28249), .Z(n28247) );
  NANDN U28408 ( .A(n28249), .B(n28248), .Z(n28244) );
  ANDN U28409 ( .B(B[197]), .A(n76), .Z(n28028) );
  XNOR U28410 ( .A(n28036), .B(n28250), .Z(n28029) );
  XNOR U28411 ( .A(n28035), .B(n28033), .Z(n28250) );
  AND U28412 ( .A(n28251), .B(n28252), .Z(n28033) );
  NANDN U28413 ( .A(n28253), .B(n28254), .Z(n28252) );
  OR U28414 ( .A(n28255), .B(n28256), .Z(n28254) );
  NAND U28415 ( .A(n28256), .B(n28255), .Z(n28251) );
  ANDN U28416 ( .B(B[198]), .A(n77), .Z(n28035) );
  XNOR U28417 ( .A(n28043), .B(n28257), .Z(n28036) );
  XNOR U28418 ( .A(n28042), .B(n28040), .Z(n28257) );
  AND U28419 ( .A(n28258), .B(n28259), .Z(n28040) );
  NANDN U28420 ( .A(n28260), .B(n28261), .Z(n28259) );
  NANDN U28421 ( .A(n28262), .B(n28263), .Z(n28261) );
  NANDN U28422 ( .A(n28263), .B(n28262), .Z(n28258) );
  ANDN U28423 ( .B(B[199]), .A(n78), .Z(n28042) );
  XNOR U28424 ( .A(n28050), .B(n28264), .Z(n28043) );
  XNOR U28425 ( .A(n28049), .B(n28047), .Z(n28264) );
  AND U28426 ( .A(n28265), .B(n28266), .Z(n28047) );
  NANDN U28427 ( .A(n28267), .B(n28268), .Z(n28266) );
  OR U28428 ( .A(n28269), .B(n28270), .Z(n28268) );
  NAND U28429 ( .A(n28270), .B(n28269), .Z(n28265) );
  ANDN U28430 ( .B(B[200]), .A(n79), .Z(n28049) );
  XNOR U28431 ( .A(n28057), .B(n28271), .Z(n28050) );
  XNOR U28432 ( .A(n28056), .B(n28054), .Z(n28271) );
  AND U28433 ( .A(n28272), .B(n28273), .Z(n28054) );
  NANDN U28434 ( .A(n28274), .B(n28275), .Z(n28273) );
  NANDN U28435 ( .A(n28276), .B(n28277), .Z(n28275) );
  NANDN U28436 ( .A(n28277), .B(n28276), .Z(n28272) );
  ANDN U28437 ( .B(B[201]), .A(n80), .Z(n28056) );
  XNOR U28438 ( .A(n28064), .B(n28278), .Z(n28057) );
  XNOR U28439 ( .A(n28063), .B(n28061), .Z(n28278) );
  AND U28440 ( .A(n28279), .B(n28280), .Z(n28061) );
  NANDN U28441 ( .A(n28281), .B(n28282), .Z(n28280) );
  OR U28442 ( .A(n28283), .B(n28284), .Z(n28282) );
  NAND U28443 ( .A(n28284), .B(n28283), .Z(n28279) );
  ANDN U28444 ( .B(B[202]), .A(n81), .Z(n28063) );
  XNOR U28445 ( .A(n28071), .B(n28285), .Z(n28064) );
  XNOR U28446 ( .A(n28070), .B(n28068), .Z(n28285) );
  AND U28447 ( .A(n28286), .B(n28287), .Z(n28068) );
  NANDN U28448 ( .A(n28288), .B(n28289), .Z(n28287) );
  NAND U28449 ( .A(n28290), .B(n28291), .Z(n28289) );
  ANDN U28450 ( .B(B[203]), .A(n82), .Z(n28070) );
  XOR U28451 ( .A(n28077), .B(n28292), .Z(n28071) );
  XNOR U28452 ( .A(n28075), .B(n28078), .Z(n28292) );
  NAND U28453 ( .A(A[2]), .B(B[204]), .Z(n28078) );
  NANDN U28454 ( .A(n28293), .B(n28294), .Z(n28075) );
  AND U28455 ( .A(A[0]), .B(B[205]), .Z(n28294) );
  XNOR U28456 ( .A(n28080), .B(n28295), .Z(n28077) );
  NAND U28457 ( .A(A[0]), .B(B[206]), .Z(n28295) );
  NAND U28458 ( .A(B[205]), .B(A[1]), .Z(n28080) );
  NAND U28459 ( .A(n28296), .B(n28297), .Z(n384) );
  NANDN U28460 ( .A(n28298), .B(n28299), .Z(n28297) );
  OR U28461 ( .A(n28300), .B(n28301), .Z(n28299) );
  NAND U28462 ( .A(n28301), .B(n28300), .Z(n28296) );
  XOR U28463 ( .A(n386), .B(n385), .Z(\A1[203] ) );
  XOR U28464 ( .A(n28301), .B(n28302), .Z(n385) );
  XNOR U28465 ( .A(n28300), .B(n28298), .Z(n28302) );
  AND U28466 ( .A(n28303), .B(n28304), .Z(n28298) );
  NANDN U28467 ( .A(n28305), .B(n28306), .Z(n28304) );
  NANDN U28468 ( .A(n28307), .B(n28308), .Z(n28306) );
  NANDN U28469 ( .A(n28308), .B(n28307), .Z(n28303) );
  ANDN U28470 ( .B(B[174]), .A(n54), .Z(n28300) );
  XNOR U28471 ( .A(n28095), .B(n28309), .Z(n28301) );
  XNOR U28472 ( .A(n28094), .B(n28092), .Z(n28309) );
  AND U28473 ( .A(n28310), .B(n28311), .Z(n28092) );
  NANDN U28474 ( .A(n28312), .B(n28313), .Z(n28311) );
  OR U28475 ( .A(n28314), .B(n28315), .Z(n28313) );
  NAND U28476 ( .A(n28315), .B(n28314), .Z(n28310) );
  ANDN U28477 ( .B(B[175]), .A(n55), .Z(n28094) );
  XNOR U28478 ( .A(n28102), .B(n28316), .Z(n28095) );
  XNOR U28479 ( .A(n28101), .B(n28099), .Z(n28316) );
  AND U28480 ( .A(n28317), .B(n28318), .Z(n28099) );
  NANDN U28481 ( .A(n28319), .B(n28320), .Z(n28318) );
  NANDN U28482 ( .A(n28321), .B(n28322), .Z(n28320) );
  NANDN U28483 ( .A(n28322), .B(n28321), .Z(n28317) );
  ANDN U28484 ( .B(B[176]), .A(n56), .Z(n28101) );
  XNOR U28485 ( .A(n28109), .B(n28323), .Z(n28102) );
  XNOR U28486 ( .A(n28108), .B(n28106), .Z(n28323) );
  AND U28487 ( .A(n28324), .B(n28325), .Z(n28106) );
  NANDN U28488 ( .A(n28326), .B(n28327), .Z(n28325) );
  OR U28489 ( .A(n28328), .B(n28329), .Z(n28327) );
  NAND U28490 ( .A(n28329), .B(n28328), .Z(n28324) );
  ANDN U28491 ( .B(B[177]), .A(n57), .Z(n28108) );
  XNOR U28492 ( .A(n28116), .B(n28330), .Z(n28109) );
  XNOR U28493 ( .A(n28115), .B(n28113), .Z(n28330) );
  AND U28494 ( .A(n28331), .B(n28332), .Z(n28113) );
  NANDN U28495 ( .A(n28333), .B(n28334), .Z(n28332) );
  NANDN U28496 ( .A(n28335), .B(n28336), .Z(n28334) );
  NANDN U28497 ( .A(n28336), .B(n28335), .Z(n28331) );
  ANDN U28498 ( .B(B[178]), .A(n58), .Z(n28115) );
  XNOR U28499 ( .A(n28123), .B(n28337), .Z(n28116) );
  XNOR U28500 ( .A(n28122), .B(n28120), .Z(n28337) );
  AND U28501 ( .A(n28338), .B(n28339), .Z(n28120) );
  NANDN U28502 ( .A(n28340), .B(n28341), .Z(n28339) );
  OR U28503 ( .A(n28342), .B(n28343), .Z(n28341) );
  NAND U28504 ( .A(n28343), .B(n28342), .Z(n28338) );
  ANDN U28505 ( .B(B[179]), .A(n59), .Z(n28122) );
  XNOR U28506 ( .A(n28130), .B(n28344), .Z(n28123) );
  XNOR U28507 ( .A(n28129), .B(n28127), .Z(n28344) );
  AND U28508 ( .A(n28345), .B(n28346), .Z(n28127) );
  NANDN U28509 ( .A(n28347), .B(n28348), .Z(n28346) );
  NANDN U28510 ( .A(n28349), .B(n28350), .Z(n28348) );
  NANDN U28511 ( .A(n28350), .B(n28349), .Z(n28345) );
  ANDN U28512 ( .B(B[180]), .A(n60), .Z(n28129) );
  XNOR U28513 ( .A(n28137), .B(n28351), .Z(n28130) );
  XNOR U28514 ( .A(n28136), .B(n28134), .Z(n28351) );
  AND U28515 ( .A(n28352), .B(n28353), .Z(n28134) );
  NANDN U28516 ( .A(n28354), .B(n28355), .Z(n28353) );
  OR U28517 ( .A(n28356), .B(n28357), .Z(n28355) );
  NAND U28518 ( .A(n28357), .B(n28356), .Z(n28352) );
  ANDN U28519 ( .B(B[181]), .A(n61), .Z(n28136) );
  XNOR U28520 ( .A(n28144), .B(n28358), .Z(n28137) );
  XNOR U28521 ( .A(n28143), .B(n28141), .Z(n28358) );
  AND U28522 ( .A(n28359), .B(n28360), .Z(n28141) );
  NANDN U28523 ( .A(n28361), .B(n28362), .Z(n28360) );
  NANDN U28524 ( .A(n28363), .B(n28364), .Z(n28362) );
  NANDN U28525 ( .A(n28364), .B(n28363), .Z(n28359) );
  ANDN U28526 ( .B(B[182]), .A(n62), .Z(n28143) );
  XNOR U28527 ( .A(n28151), .B(n28365), .Z(n28144) );
  XNOR U28528 ( .A(n28150), .B(n28148), .Z(n28365) );
  AND U28529 ( .A(n28366), .B(n28367), .Z(n28148) );
  NANDN U28530 ( .A(n28368), .B(n28369), .Z(n28367) );
  OR U28531 ( .A(n28370), .B(n28371), .Z(n28369) );
  NAND U28532 ( .A(n28371), .B(n28370), .Z(n28366) );
  ANDN U28533 ( .B(B[183]), .A(n63), .Z(n28150) );
  XNOR U28534 ( .A(n28158), .B(n28372), .Z(n28151) );
  XNOR U28535 ( .A(n28157), .B(n28155), .Z(n28372) );
  AND U28536 ( .A(n28373), .B(n28374), .Z(n28155) );
  NANDN U28537 ( .A(n28375), .B(n28376), .Z(n28374) );
  NANDN U28538 ( .A(n28377), .B(n28378), .Z(n28376) );
  NANDN U28539 ( .A(n28378), .B(n28377), .Z(n28373) );
  ANDN U28540 ( .B(B[184]), .A(n64), .Z(n28157) );
  XNOR U28541 ( .A(n28165), .B(n28379), .Z(n28158) );
  XNOR U28542 ( .A(n28164), .B(n28162), .Z(n28379) );
  AND U28543 ( .A(n28380), .B(n28381), .Z(n28162) );
  NANDN U28544 ( .A(n28382), .B(n28383), .Z(n28381) );
  OR U28545 ( .A(n28384), .B(n28385), .Z(n28383) );
  NAND U28546 ( .A(n28385), .B(n28384), .Z(n28380) );
  ANDN U28547 ( .B(B[185]), .A(n65), .Z(n28164) );
  XNOR U28548 ( .A(n28172), .B(n28386), .Z(n28165) );
  XNOR U28549 ( .A(n28171), .B(n28169), .Z(n28386) );
  AND U28550 ( .A(n28387), .B(n28388), .Z(n28169) );
  NANDN U28551 ( .A(n28389), .B(n28390), .Z(n28388) );
  NANDN U28552 ( .A(n28391), .B(n28392), .Z(n28390) );
  NANDN U28553 ( .A(n28392), .B(n28391), .Z(n28387) );
  ANDN U28554 ( .B(B[186]), .A(n66), .Z(n28171) );
  XNOR U28555 ( .A(n28179), .B(n28393), .Z(n28172) );
  XNOR U28556 ( .A(n28178), .B(n28176), .Z(n28393) );
  AND U28557 ( .A(n28394), .B(n28395), .Z(n28176) );
  NANDN U28558 ( .A(n28396), .B(n28397), .Z(n28395) );
  OR U28559 ( .A(n28398), .B(n28399), .Z(n28397) );
  NAND U28560 ( .A(n28399), .B(n28398), .Z(n28394) );
  ANDN U28561 ( .B(B[187]), .A(n67), .Z(n28178) );
  XNOR U28562 ( .A(n28186), .B(n28400), .Z(n28179) );
  XNOR U28563 ( .A(n28185), .B(n28183), .Z(n28400) );
  AND U28564 ( .A(n28401), .B(n28402), .Z(n28183) );
  NANDN U28565 ( .A(n28403), .B(n28404), .Z(n28402) );
  NANDN U28566 ( .A(n28405), .B(n28406), .Z(n28404) );
  NANDN U28567 ( .A(n28406), .B(n28405), .Z(n28401) );
  ANDN U28568 ( .B(B[188]), .A(n68), .Z(n28185) );
  XNOR U28569 ( .A(n28193), .B(n28407), .Z(n28186) );
  XNOR U28570 ( .A(n28192), .B(n28190), .Z(n28407) );
  AND U28571 ( .A(n28408), .B(n28409), .Z(n28190) );
  NANDN U28572 ( .A(n28410), .B(n28411), .Z(n28409) );
  OR U28573 ( .A(n28412), .B(n28413), .Z(n28411) );
  NAND U28574 ( .A(n28413), .B(n28412), .Z(n28408) );
  ANDN U28575 ( .B(B[189]), .A(n69), .Z(n28192) );
  XNOR U28576 ( .A(n28200), .B(n28414), .Z(n28193) );
  XNOR U28577 ( .A(n28199), .B(n28197), .Z(n28414) );
  AND U28578 ( .A(n28415), .B(n28416), .Z(n28197) );
  NANDN U28579 ( .A(n28417), .B(n28418), .Z(n28416) );
  NANDN U28580 ( .A(n28419), .B(n28420), .Z(n28418) );
  NANDN U28581 ( .A(n28420), .B(n28419), .Z(n28415) );
  ANDN U28582 ( .B(B[190]), .A(n70), .Z(n28199) );
  XNOR U28583 ( .A(n28207), .B(n28421), .Z(n28200) );
  XNOR U28584 ( .A(n28206), .B(n28204), .Z(n28421) );
  AND U28585 ( .A(n28422), .B(n28423), .Z(n28204) );
  NANDN U28586 ( .A(n28424), .B(n28425), .Z(n28423) );
  OR U28587 ( .A(n28426), .B(n28427), .Z(n28425) );
  NAND U28588 ( .A(n28427), .B(n28426), .Z(n28422) );
  ANDN U28589 ( .B(B[191]), .A(n71), .Z(n28206) );
  XNOR U28590 ( .A(n28214), .B(n28428), .Z(n28207) );
  XNOR U28591 ( .A(n28213), .B(n28211), .Z(n28428) );
  AND U28592 ( .A(n28429), .B(n28430), .Z(n28211) );
  NANDN U28593 ( .A(n28431), .B(n28432), .Z(n28430) );
  NANDN U28594 ( .A(n28433), .B(n28434), .Z(n28432) );
  NANDN U28595 ( .A(n28434), .B(n28433), .Z(n28429) );
  ANDN U28596 ( .B(B[192]), .A(n72), .Z(n28213) );
  XNOR U28597 ( .A(n28221), .B(n28435), .Z(n28214) );
  XNOR U28598 ( .A(n28220), .B(n28218), .Z(n28435) );
  AND U28599 ( .A(n28436), .B(n28437), .Z(n28218) );
  NANDN U28600 ( .A(n28438), .B(n28439), .Z(n28437) );
  OR U28601 ( .A(n28440), .B(n28441), .Z(n28439) );
  NAND U28602 ( .A(n28441), .B(n28440), .Z(n28436) );
  ANDN U28603 ( .B(B[193]), .A(n73), .Z(n28220) );
  XNOR U28604 ( .A(n28228), .B(n28442), .Z(n28221) );
  XNOR U28605 ( .A(n28227), .B(n28225), .Z(n28442) );
  AND U28606 ( .A(n28443), .B(n28444), .Z(n28225) );
  NANDN U28607 ( .A(n28445), .B(n28446), .Z(n28444) );
  NANDN U28608 ( .A(n28447), .B(n28448), .Z(n28446) );
  NANDN U28609 ( .A(n28448), .B(n28447), .Z(n28443) );
  ANDN U28610 ( .B(B[194]), .A(n74), .Z(n28227) );
  XNOR U28611 ( .A(n28235), .B(n28449), .Z(n28228) );
  XNOR U28612 ( .A(n28234), .B(n28232), .Z(n28449) );
  AND U28613 ( .A(n28450), .B(n28451), .Z(n28232) );
  NANDN U28614 ( .A(n28452), .B(n28453), .Z(n28451) );
  OR U28615 ( .A(n28454), .B(n28455), .Z(n28453) );
  NAND U28616 ( .A(n28455), .B(n28454), .Z(n28450) );
  ANDN U28617 ( .B(B[195]), .A(n75), .Z(n28234) );
  XNOR U28618 ( .A(n28242), .B(n28456), .Z(n28235) );
  XNOR U28619 ( .A(n28241), .B(n28239), .Z(n28456) );
  AND U28620 ( .A(n28457), .B(n28458), .Z(n28239) );
  NANDN U28621 ( .A(n28459), .B(n28460), .Z(n28458) );
  NANDN U28622 ( .A(n28461), .B(n28462), .Z(n28460) );
  NANDN U28623 ( .A(n28462), .B(n28461), .Z(n28457) );
  ANDN U28624 ( .B(B[196]), .A(n76), .Z(n28241) );
  XNOR U28625 ( .A(n28249), .B(n28463), .Z(n28242) );
  XNOR U28626 ( .A(n28248), .B(n28246), .Z(n28463) );
  AND U28627 ( .A(n28464), .B(n28465), .Z(n28246) );
  NANDN U28628 ( .A(n28466), .B(n28467), .Z(n28465) );
  OR U28629 ( .A(n28468), .B(n28469), .Z(n28467) );
  NAND U28630 ( .A(n28469), .B(n28468), .Z(n28464) );
  ANDN U28631 ( .B(B[197]), .A(n77), .Z(n28248) );
  XNOR U28632 ( .A(n28256), .B(n28470), .Z(n28249) );
  XNOR U28633 ( .A(n28255), .B(n28253), .Z(n28470) );
  AND U28634 ( .A(n28471), .B(n28472), .Z(n28253) );
  NANDN U28635 ( .A(n28473), .B(n28474), .Z(n28472) );
  NANDN U28636 ( .A(n28475), .B(n28476), .Z(n28474) );
  NANDN U28637 ( .A(n28476), .B(n28475), .Z(n28471) );
  ANDN U28638 ( .B(B[198]), .A(n78), .Z(n28255) );
  XNOR U28639 ( .A(n28263), .B(n28477), .Z(n28256) );
  XNOR U28640 ( .A(n28262), .B(n28260), .Z(n28477) );
  AND U28641 ( .A(n28478), .B(n28479), .Z(n28260) );
  NANDN U28642 ( .A(n28480), .B(n28481), .Z(n28479) );
  OR U28643 ( .A(n28482), .B(n28483), .Z(n28481) );
  NAND U28644 ( .A(n28483), .B(n28482), .Z(n28478) );
  ANDN U28645 ( .B(B[199]), .A(n79), .Z(n28262) );
  XNOR U28646 ( .A(n28270), .B(n28484), .Z(n28263) );
  XNOR U28647 ( .A(n28269), .B(n28267), .Z(n28484) );
  AND U28648 ( .A(n28485), .B(n28486), .Z(n28267) );
  NANDN U28649 ( .A(n28487), .B(n28488), .Z(n28486) );
  NANDN U28650 ( .A(n28489), .B(n28490), .Z(n28488) );
  NANDN U28651 ( .A(n28490), .B(n28489), .Z(n28485) );
  ANDN U28652 ( .B(B[200]), .A(n80), .Z(n28269) );
  XNOR U28653 ( .A(n28277), .B(n28491), .Z(n28270) );
  XNOR U28654 ( .A(n28276), .B(n28274), .Z(n28491) );
  AND U28655 ( .A(n28492), .B(n28493), .Z(n28274) );
  NANDN U28656 ( .A(n28494), .B(n28495), .Z(n28493) );
  OR U28657 ( .A(n28496), .B(n28497), .Z(n28495) );
  NAND U28658 ( .A(n28497), .B(n28496), .Z(n28492) );
  ANDN U28659 ( .B(B[201]), .A(n81), .Z(n28276) );
  XNOR U28660 ( .A(n28284), .B(n28498), .Z(n28277) );
  XNOR U28661 ( .A(n28283), .B(n28281), .Z(n28498) );
  AND U28662 ( .A(n28499), .B(n28500), .Z(n28281) );
  NANDN U28663 ( .A(n28501), .B(n28502), .Z(n28500) );
  NAND U28664 ( .A(n28503), .B(n28504), .Z(n28502) );
  ANDN U28665 ( .B(B[202]), .A(n82), .Z(n28283) );
  XOR U28666 ( .A(n28290), .B(n28505), .Z(n28284) );
  XNOR U28667 ( .A(n28288), .B(n28291), .Z(n28505) );
  NAND U28668 ( .A(A[2]), .B(B[203]), .Z(n28291) );
  NANDN U28669 ( .A(n28506), .B(n28507), .Z(n28288) );
  AND U28670 ( .A(A[0]), .B(B[204]), .Z(n28507) );
  XNOR U28671 ( .A(n28293), .B(n28508), .Z(n28290) );
  NAND U28672 ( .A(A[0]), .B(B[205]), .Z(n28508) );
  NAND U28673 ( .A(B[204]), .B(A[1]), .Z(n28293) );
  NAND U28674 ( .A(n28509), .B(n28510), .Z(n386) );
  NANDN U28675 ( .A(n28511), .B(n28512), .Z(n28510) );
  OR U28676 ( .A(n28513), .B(n28514), .Z(n28512) );
  NAND U28677 ( .A(n28514), .B(n28513), .Z(n28509) );
  XOR U28678 ( .A(n388), .B(n387), .Z(\A1[202] ) );
  XOR U28679 ( .A(n28514), .B(n28515), .Z(n387) );
  XNOR U28680 ( .A(n28513), .B(n28511), .Z(n28515) );
  AND U28681 ( .A(n28516), .B(n28517), .Z(n28511) );
  NANDN U28682 ( .A(n28518), .B(n28519), .Z(n28517) );
  NANDN U28683 ( .A(n28520), .B(n28521), .Z(n28519) );
  NANDN U28684 ( .A(n28521), .B(n28520), .Z(n28516) );
  ANDN U28685 ( .B(B[173]), .A(n54), .Z(n28513) );
  XNOR U28686 ( .A(n28308), .B(n28522), .Z(n28514) );
  XNOR U28687 ( .A(n28307), .B(n28305), .Z(n28522) );
  AND U28688 ( .A(n28523), .B(n28524), .Z(n28305) );
  NANDN U28689 ( .A(n28525), .B(n28526), .Z(n28524) );
  OR U28690 ( .A(n28527), .B(n28528), .Z(n28526) );
  NAND U28691 ( .A(n28528), .B(n28527), .Z(n28523) );
  ANDN U28692 ( .B(B[174]), .A(n55), .Z(n28307) );
  XNOR U28693 ( .A(n28315), .B(n28529), .Z(n28308) );
  XNOR U28694 ( .A(n28314), .B(n28312), .Z(n28529) );
  AND U28695 ( .A(n28530), .B(n28531), .Z(n28312) );
  NANDN U28696 ( .A(n28532), .B(n28533), .Z(n28531) );
  NANDN U28697 ( .A(n28534), .B(n28535), .Z(n28533) );
  NANDN U28698 ( .A(n28535), .B(n28534), .Z(n28530) );
  ANDN U28699 ( .B(B[175]), .A(n56), .Z(n28314) );
  XNOR U28700 ( .A(n28322), .B(n28536), .Z(n28315) );
  XNOR U28701 ( .A(n28321), .B(n28319), .Z(n28536) );
  AND U28702 ( .A(n28537), .B(n28538), .Z(n28319) );
  NANDN U28703 ( .A(n28539), .B(n28540), .Z(n28538) );
  OR U28704 ( .A(n28541), .B(n28542), .Z(n28540) );
  NAND U28705 ( .A(n28542), .B(n28541), .Z(n28537) );
  ANDN U28706 ( .B(B[176]), .A(n57), .Z(n28321) );
  XNOR U28707 ( .A(n28329), .B(n28543), .Z(n28322) );
  XNOR U28708 ( .A(n28328), .B(n28326), .Z(n28543) );
  AND U28709 ( .A(n28544), .B(n28545), .Z(n28326) );
  NANDN U28710 ( .A(n28546), .B(n28547), .Z(n28545) );
  NANDN U28711 ( .A(n28548), .B(n28549), .Z(n28547) );
  NANDN U28712 ( .A(n28549), .B(n28548), .Z(n28544) );
  ANDN U28713 ( .B(B[177]), .A(n58), .Z(n28328) );
  XNOR U28714 ( .A(n28336), .B(n28550), .Z(n28329) );
  XNOR U28715 ( .A(n28335), .B(n28333), .Z(n28550) );
  AND U28716 ( .A(n28551), .B(n28552), .Z(n28333) );
  NANDN U28717 ( .A(n28553), .B(n28554), .Z(n28552) );
  OR U28718 ( .A(n28555), .B(n28556), .Z(n28554) );
  NAND U28719 ( .A(n28556), .B(n28555), .Z(n28551) );
  ANDN U28720 ( .B(B[178]), .A(n59), .Z(n28335) );
  XNOR U28721 ( .A(n28343), .B(n28557), .Z(n28336) );
  XNOR U28722 ( .A(n28342), .B(n28340), .Z(n28557) );
  AND U28723 ( .A(n28558), .B(n28559), .Z(n28340) );
  NANDN U28724 ( .A(n28560), .B(n28561), .Z(n28559) );
  NANDN U28725 ( .A(n28562), .B(n28563), .Z(n28561) );
  NANDN U28726 ( .A(n28563), .B(n28562), .Z(n28558) );
  ANDN U28727 ( .B(B[179]), .A(n60), .Z(n28342) );
  XNOR U28728 ( .A(n28350), .B(n28564), .Z(n28343) );
  XNOR U28729 ( .A(n28349), .B(n28347), .Z(n28564) );
  AND U28730 ( .A(n28565), .B(n28566), .Z(n28347) );
  NANDN U28731 ( .A(n28567), .B(n28568), .Z(n28566) );
  OR U28732 ( .A(n28569), .B(n28570), .Z(n28568) );
  NAND U28733 ( .A(n28570), .B(n28569), .Z(n28565) );
  ANDN U28734 ( .B(B[180]), .A(n61), .Z(n28349) );
  XNOR U28735 ( .A(n28357), .B(n28571), .Z(n28350) );
  XNOR U28736 ( .A(n28356), .B(n28354), .Z(n28571) );
  AND U28737 ( .A(n28572), .B(n28573), .Z(n28354) );
  NANDN U28738 ( .A(n28574), .B(n28575), .Z(n28573) );
  NANDN U28739 ( .A(n28576), .B(n28577), .Z(n28575) );
  NANDN U28740 ( .A(n28577), .B(n28576), .Z(n28572) );
  ANDN U28741 ( .B(B[181]), .A(n62), .Z(n28356) );
  XNOR U28742 ( .A(n28364), .B(n28578), .Z(n28357) );
  XNOR U28743 ( .A(n28363), .B(n28361), .Z(n28578) );
  AND U28744 ( .A(n28579), .B(n28580), .Z(n28361) );
  NANDN U28745 ( .A(n28581), .B(n28582), .Z(n28580) );
  OR U28746 ( .A(n28583), .B(n28584), .Z(n28582) );
  NAND U28747 ( .A(n28584), .B(n28583), .Z(n28579) );
  ANDN U28748 ( .B(B[182]), .A(n63), .Z(n28363) );
  XNOR U28749 ( .A(n28371), .B(n28585), .Z(n28364) );
  XNOR U28750 ( .A(n28370), .B(n28368), .Z(n28585) );
  AND U28751 ( .A(n28586), .B(n28587), .Z(n28368) );
  NANDN U28752 ( .A(n28588), .B(n28589), .Z(n28587) );
  NANDN U28753 ( .A(n28590), .B(n28591), .Z(n28589) );
  NANDN U28754 ( .A(n28591), .B(n28590), .Z(n28586) );
  ANDN U28755 ( .B(B[183]), .A(n64), .Z(n28370) );
  XNOR U28756 ( .A(n28378), .B(n28592), .Z(n28371) );
  XNOR U28757 ( .A(n28377), .B(n28375), .Z(n28592) );
  AND U28758 ( .A(n28593), .B(n28594), .Z(n28375) );
  NANDN U28759 ( .A(n28595), .B(n28596), .Z(n28594) );
  OR U28760 ( .A(n28597), .B(n28598), .Z(n28596) );
  NAND U28761 ( .A(n28598), .B(n28597), .Z(n28593) );
  ANDN U28762 ( .B(B[184]), .A(n65), .Z(n28377) );
  XNOR U28763 ( .A(n28385), .B(n28599), .Z(n28378) );
  XNOR U28764 ( .A(n28384), .B(n28382), .Z(n28599) );
  AND U28765 ( .A(n28600), .B(n28601), .Z(n28382) );
  NANDN U28766 ( .A(n28602), .B(n28603), .Z(n28601) );
  NANDN U28767 ( .A(n28604), .B(n28605), .Z(n28603) );
  NANDN U28768 ( .A(n28605), .B(n28604), .Z(n28600) );
  ANDN U28769 ( .B(B[185]), .A(n66), .Z(n28384) );
  XNOR U28770 ( .A(n28392), .B(n28606), .Z(n28385) );
  XNOR U28771 ( .A(n28391), .B(n28389), .Z(n28606) );
  AND U28772 ( .A(n28607), .B(n28608), .Z(n28389) );
  NANDN U28773 ( .A(n28609), .B(n28610), .Z(n28608) );
  OR U28774 ( .A(n28611), .B(n28612), .Z(n28610) );
  NAND U28775 ( .A(n28612), .B(n28611), .Z(n28607) );
  ANDN U28776 ( .B(B[186]), .A(n67), .Z(n28391) );
  XNOR U28777 ( .A(n28399), .B(n28613), .Z(n28392) );
  XNOR U28778 ( .A(n28398), .B(n28396), .Z(n28613) );
  AND U28779 ( .A(n28614), .B(n28615), .Z(n28396) );
  NANDN U28780 ( .A(n28616), .B(n28617), .Z(n28615) );
  NANDN U28781 ( .A(n28618), .B(n28619), .Z(n28617) );
  NANDN U28782 ( .A(n28619), .B(n28618), .Z(n28614) );
  ANDN U28783 ( .B(B[187]), .A(n68), .Z(n28398) );
  XNOR U28784 ( .A(n28406), .B(n28620), .Z(n28399) );
  XNOR U28785 ( .A(n28405), .B(n28403), .Z(n28620) );
  AND U28786 ( .A(n28621), .B(n28622), .Z(n28403) );
  NANDN U28787 ( .A(n28623), .B(n28624), .Z(n28622) );
  OR U28788 ( .A(n28625), .B(n28626), .Z(n28624) );
  NAND U28789 ( .A(n28626), .B(n28625), .Z(n28621) );
  ANDN U28790 ( .B(B[188]), .A(n69), .Z(n28405) );
  XNOR U28791 ( .A(n28413), .B(n28627), .Z(n28406) );
  XNOR U28792 ( .A(n28412), .B(n28410), .Z(n28627) );
  AND U28793 ( .A(n28628), .B(n28629), .Z(n28410) );
  NANDN U28794 ( .A(n28630), .B(n28631), .Z(n28629) );
  NANDN U28795 ( .A(n28632), .B(n28633), .Z(n28631) );
  NANDN U28796 ( .A(n28633), .B(n28632), .Z(n28628) );
  ANDN U28797 ( .B(B[189]), .A(n70), .Z(n28412) );
  XNOR U28798 ( .A(n28420), .B(n28634), .Z(n28413) );
  XNOR U28799 ( .A(n28419), .B(n28417), .Z(n28634) );
  AND U28800 ( .A(n28635), .B(n28636), .Z(n28417) );
  NANDN U28801 ( .A(n28637), .B(n28638), .Z(n28636) );
  OR U28802 ( .A(n28639), .B(n28640), .Z(n28638) );
  NAND U28803 ( .A(n28640), .B(n28639), .Z(n28635) );
  ANDN U28804 ( .B(B[190]), .A(n71), .Z(n28419) );
  XNOR U28805 ( .A(n28427), .B(n28641), .Z(n28420) );
  XNOR U28806 ( .A(n28426), .B(n28424), .Z(n28641) );
  AND U28807 ( .A(n28642), .B(n28643), .Z(n28424) );
  NANDN U28808 ( .A(n28644), .B(n28645), .Z(n28643) );
  NANDN U28809 ( .A(n28646), .B(n28647), .Z(n28645) );
  NANDN U28810 ( .A(n28647), .B(n28646), .Z(n28642) );
  ANDN U28811 ( .B(B[191]), .A(n72), .Z(n28426) );
  XNOR U28812 ( .A(n28434), .B(n28648), .Z(n28427) );
  XNOR U28813 ( .A(n28433), .B(n28431), .Z(n28648) );
  AND U28814 ( .A(n28649), .B(n28650), .Z(n28431) );
  NANDN U28815 ( .A(n28651), .B(n28652), .Z(n28650) );
  OR U28816 ( .A(n28653), .B(n28654), .Z(n28652) );
  NAND U28817 ( .A(n28654), .B(n28653), .Z(n28649) );
  ANDN U28818 ( .B(B[192]), .A(n73), .Z(n28433) );
  XNOR U28819 ( .A(n28441), .B(n28655), .Z(n28434) );
  XNOR U28820 ( .A(n28440), .B(n28438), .Z(n28655) );
  AND U28821 ( .A(n28656), .B(n28657), .Z(n28438) );
  NANDN U28822 ( .A(n28658), .B(n28659), .Z(n28657) );
  NANDN U28823 ( .A(n28660), .B(n28661), .Z(n28659) );
  NANDN U28824 ( .A(n28661), .B(n28660), .Z(n28656) );
  ANDN U28825 ( .B(B[193]), .A(n74), .Z(n28440) );
  XNOR U28826 ( .A(n28448), .B(n28662), .Z(n28441) );
  XNOR U28827 ( .A(n28447), .B(n28445), .Z(n28662) );
  AND U28828 ( .A(n28663), .B(n28664), .Z(n28445) );
  NANDN U28829 ( .A(n28665), .B(n28666), .Z(n28664) );
  OR U28830 ( .A(n28667), .B(n28668), .Z(n28666) );
  NAND U28831 ( .A(n28668), .B(n28667), .Z(n28663) );
  ANDN U28832 ( .B(B[194]), .A(n75), .Z(n28447) );
  XNOR U28833 ( .A(n28455), .B(n28669), .Z(n28448) );
  XNOR U28834 ( .A(n28454), .B(n28452), .Z(n28669) );
  AND U28835 ( .A(n28670), .B(n28671), .Z(n28452) );
  NANDN U28836 ( .A(n28672), .B(n28673), .Z(n28671) );
  NANDN U28837 ( .A(n28674), .B(n28675), .Z(n28673) );
  NANDN U28838 ( .A(n28675), .B(n28674), .Z(n28670) );
  ANDN U28839 ( .B(B[195]), .A(n76), .Z(n28454) );
  XNOR U28840 ( .A(n28462), .B(n28676), .Z(n28455) );
  XNOR U28841 ( .A(n28461), .B(n28459), .Z(n28676) );
  AND U28842 ( .A(n28677), .B(n28678), .Z(n28459) );
  NANDN U28843 ( .A(n28679), .B(n28680), .Z(n28678) );
  OR U28844 ( .A(n28681), .B(n28682), .Z(n28680) );
  NAND U28845 ( .A(n28682), .B(n28681), .Z(n28677) );
  ANDN U28846 ( .B(B[196]), .A(n77), .Z(n28461) );
  XNOR U28847 ( .A(n28469), .B(n28683), .Z(n28462) );
  XNOR U28848 ( .A(n28468), .B(n28466), .Z(n28683) );
  AND U28849 ( .A(n28684), .B(n28685), .Z(n28466) );
  NANDN U28850 ( .A(n28686), .B(n28687), .Z(n28685) );
  NANDN U28851 ( .A(n28688), .B(n28689), .Z(n28687) );
  NANDN U28852 ( .A(n28689), .B(n28688), .Z(n28684) );
  ANDN U28853 ( .B(B[197]), .A(n78), .Z(n28468) );
  XNOR U28854 ( .A(n28476), .B(n28690), .Z(n28469) );
  XNOR U28855 ( .A(n28475), .B(n28473), .Z(n28690) );
  AND U28856 ( .A(n28691), .B(n28692), .Z(n28473) );
  NANDN U28857 ( .A(n28693), .B(n28694), .Z(n28692) );
  OR U28858 ( .A(n28695), .B(n28696), .Z(n28694) );
  NAND U28859 ( .A(n28696), .B(n28695), .Z(n28691) );
  ANDN U28860 ( .B(B[198]), .A(n79), .Z(n28475) );
  XNOR U28861 ( .A(n28483), .B(n28697), .Z(n28476) );
  XNOR U28862 ( .A(n28482), .B(n28480), .Z(n28697) );
  AND U28863 ( .A(n28698), .B(n28699), .Z(n28480) );
  NANDN U28864 ( .A(n28700), .B(n28701), .Z(n28699) );
  NANDN U28865 ( .A(n28702), .B(n28703), .Z(n28701) );
  NANDN U28866 ( .A(n28703), .B(n28702), .Z(n28698) );
  ANDN U28867 ( .B(B[199]), .A(n80), .Z(n28482) );
  XNOR U28868 ( .A(n28490), .B(n28704), .Z(n28483) );
  XNOR U28869 ( .A(n28489), .B(n28487), .Z(n28704) );
  AND U28870 ( .A(n28705), .B(n28706), .Z(n28487) );
  NANDN U28871 ( .A(n28707), .B(n28708), .Z(n28706) );
  OR U28872 ( .A(n28709), .B(n28710), .Z(n28708) );
  NAND U28873 ( .A(n28710), .B(n28709), .Z(n28705) );
  ANDN U28874 ( .B(B[200]), .A(n81), .Z(n28489) );
  XNOR U28875 ( .A(n28497), .B(n28711), .Z(n28490) );
  XNOR U28876 ( .A(n28496), .B(n28494), .Z(n28711) );
  AND U28877 ( .A(n28712), .B(n28713), .Z(n28494) );
  NANDN U28878 ( .A(n28714), .B(n28715), .Z(n28713) );
  NAND U28879 ( .A(n28716), .B(n28717), .Z(n28715) );
  ANDN U28880 ( .B(B[201]), .A(n82), .Z(n28496) );
  XOR U28881 ( .A(n28503), .B(n28718), .Z(n28497) );
  XNOR U28882 ( .A(n28501), .B(n28504), .Z(n28718) );
  NAND U28883 ( .A(A[2]), .B(B[202]), .Z(n28504) );
  NANDN U28884 ( .A(n28719), .B(n28720), .Z(n28501) );
  AND U28885 ( .A(A[0]), .B(B[203]), .Z(n28720) );
  XNOR U28886 ( .A(n28506), .B(n28721), .Z(n28503) );
  NAND U28887 ( .A(A[0]), .B(B[204]), .Z(n28721) );
  NAND U28888 ( .A(B[203]), .B(A[1]), .Z(n28506) );
  NAND U28889 ( .A(n28722), .B(n28723), .Z(n388) );
  NANDN U28890 ( .A(n28724), .B(n28725), .Z(n28723) );
  OR U28891 ( .A(n28726), .B(n28727), .Z(n28725) );
  NAND U28892 ( .A(n28727), .B(n28726), .Z(n28722) );
  XOR U28893 ( .A(n390), .B(n389), .Z(\A1[201] ) );
  XOR U28894 ( .A(n28727), .B(n28728), .Z(n389) );
  XNOR U28895 ( .A(n28726), .B(n28724), .Z(n28728) );
  AND U28896 ( .A(n28729), .B(n28730), .Z(n28724) );
  NANDN U28897 ( .A(n28731), .B(n28732), .Z(n28730) );
  NANDN U28898 ( .A(n28733), .B(n28734), .Z(n28732) );
  NANDN U28899 ( .A(n28734), .B(n28733), .Z(n28729) );
  ANDN U28900 ( .B(B[172]), .A(n54), .Z(n28726) );
  XNOR U28901 ( .A(n28521), .B(n28735), .Z(n28727) );
  XNOR U28902 ( .A(n28520), .B(n28518), .Z(n28735) );
  AND U28903 ( .A(n28736), .B(n28737), .Z(n28518) );
  NANDN U28904 ( .A(n28738), .B(n28739), .Z(n28737) );
  OR U28905 ( .A(n28740), .B(n28741), .Z(n28739) );
  NAND U28906 ( .A(n28741), .B(n28740), .Z(n28736) );
  ANDN U28907 ( .B(B[173]), .A(n55), .Z(n28520) );
  XNOR U28908 ( .A(n28528), .B(n28742), .Z(n28521) );
  XNOR U28909 ( .A(n28527), .B(n28525), .Z(n28742) );
  AND U28910 ( .A(n28743), .B(n28744), .Z(n28525) );
  NANDN U28911 ( .A(n28745), .B(n28746), .Z(n28744) );
  NANDN U28912 ( .A(n28747), .B(n28748), .Z(n28746) );
  NANDN U28913 ( .A(n28748), .B(n28747), .Z(n28743) );
  ANDN U28914 ( .B(B[174]), .A(n56), .Z(n28527) );
  XNOR U28915 ( .A(n28535), .B(n28749), .Z(n28528) );
  XNOR U28916 ( .A(n28534), .B(n28532), .Z(n28749) );
  AND U28917 ( .A(n28750), .B(n28751), .Z(n28532) );
  NANDN U28918 ( .A(n28752), .B(n28753), .Z(n28751) );
  OR U28919 ( .A(n28754), .B(n28755), .Z(n28753) );
  NAND U28920 ( .A(n28755), .B(n28754), .Z(n28750) );
  ANDN U28921 ( .B(B[175]), .A(n57), .Z(n28534) );
  XNOR U28922 ( .A(n28542), .B(n28756), .Z(n28535) );
  XNOR U28923 ( .A(n28541), .B(n28539), .Z(n28756) );
  AND U28924 ( .A(n28757), .B(n28758), .Z(n28539) );
  NANDN U28925 ( .A(n28759), .B(n28760), .Z(n28758) );
  NANDN U28926 ( .A(n28761), .B(n28762), .Z(n28760) );
  NANDN U28927 ( .A(n28762), .B(n28761), .Z(n28757) );
  ANDN U28928 ( .B(B[176]), .A(n58), .Z(n28541) );
  XNOR U28929 ( .A(n28549), .B(n28763), .Z(n28542) );
  XNOR U28930 ( .A(n28548), .B(n28546), .Z(n28763) );
  AND U28931 ( .A(n28764), .B(n28765), .Z(n28546) );
  NANDN U28932 ( .A(n28766), .B(n28767), .Z(n28765) );
  OR U28933 ( .A(n28768), .B(n28769), .Z(n28767) );
  NAND U28934 ( .A(n28769), .B(n28768), .Z(n28764) );
  ANDN U28935 ( .B(B[177]), .A(n59), .Z(n28548) );
  XNOR U28936 ( .A(n28556), .B(n28770), .Z(n28549) );
  XNOR U28937 ( .A(n28555), .B(n28553), .Z(n28770) );
  AND U28938 ( .A(n28771), .B(n28772), .Z(n28553) );
  NANDN U28939 ( .A(n28773), .B(n28774), .Z(n28772) );
  NANDN U28940 ( .A(n28775), .B(n28776), .Z(n28774) );
  NANDN U28941 ( .A(n28776), .B(n28775), .Z(n28771) );
  ANDN U28942 ( .B(B[178]), .A(n60), .Z(n28555) );
  XNOR U28943 ( .A(n28563), .B(n28777), .Z(n28556) );
  XNOR U28944 ( .A(n28562), .B(n28560), .Z(n28777) );
  AND U28945 ( .A(n28778), .B(n28779), .Z(n28560) );
  NANDN U28946 ( .A(n28780), .B(n28781), .Z(n28779) );
  OR U28947 ( .A(n28782), .B(n28783), .Z(n28781) );
  NAND U28948 ( .A(n28783), .B(n28782), .Z(n28778) );
  ANDN U28949 ( .B(B[179]), .A(n61), .Z(n28562) );
  XNOR U28950 ( .A(n28570), .B(n28784), .Z(n28563) );
  XNOR U28951 ( .A(n28569), .B(n28567), .Z(n28784) );
  AND U28952 ( .A(n28785), .B(n28786), .Z(n28567) );
  NANDN U28953 ( .A(n28787), .B(n28788), .Z(n28786) );
  NANDN U28954 ( .A(n28789), .B(n28790), .Z(n28788) );
  NANDN U28955 ( .A(n28790), .B(n28789), .Z(n28785) );
  ANDN U28956 ( .B(B[180]), .A(n62), .Z(n28569) );
  XNOR U28957 ( .A(n28577), .B(n28791), .Z(n28570) );
  XNOR U28958 ( .A(n28576), .B(n28574), .Z(n28791) );
  AND U28959 ( .A(n28792), .B(n28793), .Z(n28574) );
  NANDN U28960 ( .A(n28794), .B(n28795), .Z(n28793) );
  OR U28961 ( .A(n28796), .B(n28797), .Z(n28795) );
  NAND U28962 ( .A(n28797), .B(n28796), .Z(n28792) );
  ANDN U28963 ( .B(B[181]), .A(n63), .Z(n28576) );
  XNOR U28964 ( .A(n28584), .B(n28798), .Z(n28577) );
  XNOR U28965 ( .A(n28583), .B(n28581), .Z(n28798) );
  AND U28966 ( .A(n28799), .B(n28800), .Z(n28581) );
  NANDN U28967 ( .A(n28801), .B(n28802), .Z(n28800) );
  NANDN U28968 ( .A(n28803), .B(n28804), .Z(n28802) );
  NANDN U28969 ( .A(n28804), .B(n28803), .Z(n28799) );
  ANDN U28970 ( .B(B[182]), .A(n64), .Z(n28583) );
  XNOR U28971 ( .A(n28591), .B(n28805), .Z(n28584) );
  XNOR U28972 ( .A(n28590), .B(n28588), .Z(n28805) );
  AND U28973 ( .A(n28806), .B(n28807), .Z(n28588) );
  NANDN U28974 ( .A(n28808), .B(n28809), .Z(n28807) );
  OR U28975 ( .A(n28810), .B(n28811), .Z(n28809) );
  NAND U28976 ( .A(n28811), .B(n28810), .Z(n28806) );
  ANDN U28977 ( .B(B[183]), .A(n65), .Z(n28590) );
  XNOR U28978 ( .A(n28598), .B(n28812), .Z(n28591) );
  XNOR U28979 ( .A(n28597), .B(n28595), .Z(n28812) );
  AND U28980 ( .A(n28813), .B(n28814), .Z(n28595) );
  NANDN U28981 ( .A(n28815), .B(n28816), .Z(n28814) );
  NANDN U28982 ( .A(n28817), .B(n28818), .Z(n28816) );
  NANDN U28983 ( .A(n28818), .B(n28817), .Z(n28813) );
  ANDN U28984 ( .B(B[184]), .A(n66), .Z(n28597) );
  XNOR U28985 ( .A(n28605), .B(n28819), .Z(n28598) );
  XNOR U28986 ( .A(n28604), .B(n28602), .Z(n28819) );
  AND U28987 ( .A(n28820), .B(n28821), .Z(n28602) );
  NANDN U28988 ( .A(n28822), .B(n28823), .Z(n28821) );
  OR U28989 ( .A(n28824), .B(n28825), .Z(n28823) );
  NAND U28990 ( .A(n28825), .B(n28824), .Z(n28820) );
  ANDN U28991 ( .B(B[185]), .A(n67), .Z(n28604) );
  XNOR U28992 ( .A(n28612), .B(n28826), .Z(n28605) );
  XNOR U28993 ( .A(n28611), .B(n28609), .Z(n28826) );
  AND U28994 ( .A(n28827), .B(n28828), .Z(n28609) );
  NANDN U28995 ( .A(n28829), .B(n28830), .Z(n28828) );
  NANDN U28996 ( .A(n28831), .B(n28832), .Z(n28830) );
  NANDN U28997 ( .A(n28832), .B(n28831), .Z(n28827) );
  ANDN U28998 ( .B(B[186]), .A(n68), .Z(n28611) );
  XNOR U28999 ( .A(n28619), .B(n28833), .Z(n28612) );
  XNOR U29000 ( .A(n28618), .B(n28616), .Z(n28833) );
  AND U29001 ( .A(n28834), .B(n28835), .Z(n28616) );
  NANDN U29002 ( .A(n28836), .B(n28837), .Z(n28835) );
  OR U29003 ( .A(n28838), .B(n28839), .Z(n28837) );
  NAND U29004 ( .A(n28839), .B(n28838), .Z(n28834) );
  ANDN U29005 ( .B(B[187]), .A(n69), .Z(n28618) );
  XNOR U29006 ( .A(n28626), .B(n28840), .Z(n28619) );
  XNOR U29007 ( .A(n28625), .B(n28623), .Z(n28840) );
  AND U29008 ( .A(n28841), .B(n28842), .Z(n28623) );
  NANDN U29009 ( .A(n28843), .B(n28844), .Z(n28842) );
  NANDN U29010 ( .A(n28845), .B(n28846), .Z(n28844) );
  NANDN U29011 ( .A(n28846), .B(n28845), .Z(n28841) );
  ANDN U29012 ( .B(B[188]), .A(n70), .Z(n28625) );
  XNOR U29013 ( .A(n28633), .B(n28847), .Z(n28626) );
  XNOR U29014 ( .A(n28632), .B(n28630), .Z(n28847) );
  AND U29015 ( .A(n28848), .B(n28849), .Z(n28630) );
  NANDN U29016 ( .A(n28850), .B(n28851), .Z(n28849) );
  OR U29017 ( .A(n28852), .B(n28853), .Z(n28851) );
  NAND U29018 ( .A(n28853), .B(n28852), .Z(n28848) );
  ANDN U29019 ( .B(B[189]), .A(n71), .Z(n28632) );
  XNOR U29020 ( .A(n28640), .B(n28854), .Z(n28633) );
  XNOR U29021 ( .A(n28639), .B(n28637), .Z(n28854) );
  AND U29022 ( .A(n28855), .B(n28856), .Z(n28637) );
  NANDN U29023 ( .A(n28857), .B(n28858), .Z(n28856) );
  NANDN U29024 ( .A(n28859), .B(n28860), .Z(n28858) );
  NANDN U29025 ( .A(n28860), .B(n28859), .Z(n28855) );
  ANDN U29026 ( .B(B[190]), .A(n72), .Z(n28639) );
  XNOR U29027 ( .A(n28647), .B(n28861), .Z(n28640) );
  XNOR U29028 ( .A(n28646), .B(n28644), .Z(n28861) );
  AND U29029 ( .A(n28862), .B(n28863), .Z(n28644) );
  NANDN U29030 ( .A(n28864), .B(n28865), .Z(n28863) );
  OR U29031 ( .A(n28866), .B(n28867), .Z(n28865) );
  NAND U29032 ( .A(n28867), .B(n28866), .Z(n28862) );
  ANDN U29033 ( .B(B[191]), .A(n73), .Z(n28646) );
  XNOR U29034 ( .A(n28654), .B(n28868), .Z(n28647) );
  XNOR U29035 ( .A(n28653), .B(n28651), .Z(n28868) );
  AND U29036 ( .A(n28869), .B(n28870), .Z(n28651) );
  NANDN U29037 ( .A(n28871), .B(n28872), .Z(n28870) );
  NANDN U29038 ( .A(n28873), .B(n28874), .Z(n28872) );
  NANDN U29039 ( .A(n28874), .B(n28873), .Z(n28869) );
  ANDN U29040 ( .B(B[192]), .A(n74), .Z(n28653) );
  XNOR U29041 ( .A(n28661), .B(n28875), .Z(n28654) );
  XNOR U29042 ( .A(n28660), .B(n28658), .Z(n28875) );
  AND U29043 ( .A(n28876), .B(n28877), .Z(n28658) );
  NANDN U29044 ( .A(n28878), .B(n28879), .Z(n28877) );
  OR U29045 ( .A(n28880), .B(n28881), .Z(n28879) );
  NAND U29046 ( .A(n28881), .B(n28880), .Z(n28876) );
  ANDN U29047 ( .B(B[193]), .A(n75), .Z(n28660) );
  XNOR U29048 ( .A(n28668), .B(n28882), .Z(n28661) );
  XNOR U29049 ( .A(n28667), .B(n28665), .Z(n28882) );
  AND U29050 ( .A(n28883), .B(n28884), .Z(n28665) );
  NANDN U29051 ( .A(n28885), .B(n28886), .Z(n28884) );
  NANDN U29052 ( .A(n28887), .B(n28888), .Z(n28886) );
  NANDN U29053 ( .A(n28888), .B(n28887), .Z(n28883) );
  ANDN U29054 ( .B(B[194]), .A(n76), .Z(n28667) );
  XNOR U29055 ( .A(n28675), .B(n28889), .Z(n28668) );
  XNOR U29056 ( .A(n28674), .B(n28672), .Z(n28889) );
  AND U29057 ( .A(n28890), .B(n28891), .Z(n28672) );
  NANDN U29058 ( .A(n28892), .B(n28893), .Z(n28891) );
  OR U29059 ( .A(n28894), .B(n28895), .Z(n28893) );
  NAND U29060 ( .A(n28895), .B(n28894), .Z(n28890) );
  ANDN U29061 ( .B(B[195]), .A(n77), .Z(n28674) );
  XNOR U29062 ( .A(n28682), .B(n28896), .Z(n28675) );
  XNOR U29063 ( .A(n28681), .B(n28679), .Z(n28896) );
  AND U29064 ( .A(n28897), .B(n28898), .Z(n28679) );
  NANDN U29065 ( .A(n28899), .B(n28900), .Z(n28898) );
  NANDN U29066 ( .A(n28901), .B(n28902), .Z(n28900) );
  NANDN U29067 ( .A(n28902), .B(n28901), .Z(n28897) );
  ANDN U29068 ( .B(B[196]), .A(n78), .Z(n28681) );
  XNOR U29069 ( .A(n28689), .B(n28903), .Z(n28682) );
  XNOR U29070 ( .A(n28688), .B(n28686), .Z(n28903) );
  AND U29071 ( .A(n28904), .B(n28905), .Z(n28686) );
  NANDN U29072 ( .A(n28906), .B(n28907), .Z(n28905) );
  OR U29073 ( .A(n28908), .B(n28909), .Z(n28907) );
  NAND U29074 ( .A(n28909), .B(n28908), .Z(n28904) );
  ANDN U29075 ( .B(B[197]), .A(n79), .Z(n28688) );
  XNOR U29076 ( .A(n28696), .B(n28910), .Z(n28689) );
  XNOR U29077 ( .A(n28695), .B(n28693), .Z(n28910) );
  AND U29078 ( .A(n28911), .B(n28912), .Z(n28693) );
  NANDN U29079 ( .A(n28913), .B(n28914), .Z(n28912) );
  NANDN U29080 ( .A(n28915), .B(n28916), .Z(n28914) );
  NANDN U29081 ( .A(n28916), .B(n28915), .Z(n28911) );
  ANDN U29082 ( .B(B[198]), .A(n80), .Z(n28695) );
  XNOR U29083 ( .A(n28703), .B(n28917), .Z(n28696) );
  XNOR U29084 ( .A(n28702), .B(n28700), .Z(n28917) );
  AND U29085 ( .A(n28918), .B(n28919), .Z(n28700) );
  NANDN U29086 ( .A(n28920), .B(n28921), .Z(n28919) );
  OR U29087 ( .A(n28922), .B(n28923), .Z(n28921) );
  NAND U29088 ( .A(n28923), .B(n28922), .Z(n28918) );
  ANDN U29089 ( .B(B[199]), .A(n81), .Z(n28702) );
  XNOR U29090 ( .A(n28710), .B(n28924), .Z(n28703) );
  XNOR U29091 ( .A(n28709), .B(n28707), .Z(n28924) );
  AND U29092 ( .A(n28925), .B(n28926), .Z(n28707) );
  NANDN U29093 ( .A(n28927), .B(n28928), .Z(n28926) );
  NAND U29094 ( .A(n28929), .B(n28930), .Z(n28928) );
  ANDN U29095 ( .B(B[200]), .A(n82), .Z(n28709) );
  XOR U29096 ( .A(n28716), .B(n28931), .Z(n28710) );
  XNOR U29097 ( .A(n28714), .B(n28717), .Z(n28931) );
  NAND U29098 ( .A(A[2]), .B(B[201]), .Z(n28717) );
  NANDN U29099 ( .A(n28932), .B(n28933), .Z(n28714) );
  AND U29100 ( .A(A[0]), .B(B[202]), .Z(n28933) );
  XNOR U29101 ( .A(n28719), .B(n28934), .Z(n28716) );
  NAND U29102 ( .A(A[0]), .B(B[203]), .Z(n28934) );
  NAND U29103 ( .A(B[202]), .B(A[1]), .Z(n28719) );
  NAND U29104 ( .A(n28935), .B(n28936), .Z(n390) );
  NANDN U29105 ( .A(n28937), .B(n28938), .Z(n28936) );
  OR U29106 ( .A(n28939), .B(n28940), .Z(n28938) );
  NAND U29107 ( .A(n28940), .B(n28939), .Z(n28935) );
  XOR U29108 ( .A(n392), .B(n391), .Z(\A1[200] ) );
  XOR U29109 ( .A(n28940), .B(n28941), .Z(n391) );
  XNOR U29110 ( .A(n28939), .B(n28937), .Z(n28941) );
  AND U29111 ( .A(n28942), .B(n28943), .Z(n28937) );
  NANDN U29112 ( .A(n28944), .B(n28945), .Z(n28943) );
  NANDN U29113 ( .A(n28946), .B(n28947), .Z(n28945) );
  NANDN U29114 ( .A(n28947), .B(n28946), .Z(n28942) );
  ANDN U29115 ( .B(B[171]), .A(n54), .Z(n28939) );
  XNOR U29116 ( .A(n28734), .B(n28948), .Z(n28940) );
  XNOR U29117 ( .A(n28733), .B(n28731), .Z(n28948) );
  AND U29118 ( .A(n28949), .B(n28950), .Z(n28731) );
  NANDN U29119 ( .A(n28951), .B(n28952), .Z(n28950) );
  OR U29120 ( .A(n28953), .B(n28954), .Z(n28952) );
  NAND U29121 ( .A(n28954), .B(n28953), .Z(n28949) );
  ANDN U29122 ( .B(B[172]), .A(n55), .Z(n28733) );
  XNOR U29123 ( .A(n28741), .B(n28955), .Z(n28734) );
  XNOR U29124 ( .A(n28740), .B(n28738), .Z(n28955) );
  AND U29125 ( .A(n28956), .B(n28957), .Z(n28738) );
  NANDN U29126 ( .A(n28958), .B(n28959), .Z(n28957) );
  NANDN U29127 ( .A(n28960), .B(n28961), .Z(n28959) );
  NANDN U29128 ( .A(n28961), .B(n28960), .Z(n28956) );
  ANDN U29129 ( .B(B[173]), .A(n56), .Z(n28740) );
  XNOR U29130 ( .A(n28748), .B(n28962), .Z(n28741) );
  XNOR U29131 ( .A(n28747), .B(n28745), .Z(n28962) );
  AND U29132 ( .A(n28963), .B(n28964), .Z(n28745) );
  NANDN U29133 ( .A(n28965), .B(n28966), .Z(n28964) );
  OR U29134 ( .A(n28967), .B(n28968), .Z(n28966) );
  NAND U29135 ( .A(n28968), .B(n28967), .Z(n28963) );
  ANDN U29136 ( .B(B[174]), .A(n57), .Z(n28747) );
  XNOR U29137 ( .A(n28755), .B(n28969), .Z(n28748) );
  XNOR U29138 ( .A(n28754), .B(n28752), .Z(n28969) );
  AND U29139 ( .A(n28970), .B(n28971), .Z(n28752) );
  NANDN U29140 ( .A(n28972), .B(n28973), .Z(n28971) );
  NANDN U29141 ( .A(n28974), .B(n28975), .Z(n28973) );
  NANDN U29142 ( .A(n28975), .B(n28974), .Z(n28970) );
  ANDN U29143 ( .B(B[175]), .A(n58), .Z(n28754) );
  XNOR U29144 ( .A(n28762), .B(n28976), .Z(n28755) );
  XNOR U29145 ( .A(n28761), .B(n28759), .Z(n28976) );
  AND U29146 ( .A(n28977), .B(n28978), .Z(n28759) );
  NANDN U29147 ( .A(n28979), .B(n28980), .Z(n28978) );
  OR U29148 ( .A(n28981), .B(n28982), .Z(n28980) );
  NAND U29149 ( .A(n28982), .B(n28981), .Z(n28977) );
  ANDN U29150 ( .B(B[176]), .A(n59), .Z(n28761) );
  XNOR U29151 ( .A(n28769), .B(n28983), .Z(n28762) );
  XNOR U29152 ( .A(n28768), .B(n28766), .Z(n28983) );
  AND U29153 ( .A(n28984), .B(n28985), .Z(n28766) );
  NANDN U29154 ( .A(n28986), .B(n28987), .Z(n28985) );
  NANDN U29155 ( .A(n28988), .B(n28989), .Z(n28987) );
  NANDN U29156 ( .A(n28989), .B(n28988), .Z(n28984) );
  ANDN U29157 ( .B(B[177]), .A(n60), .Z(n28768) );
  XNOR U29158 ( .A(n28776), .B(n28990), .Z(n28769) );
  XNOR U29159 ( .A(n28775), .B(n28773), .Z(n28990) );
  AND U29160 ( .A(n28991), .B(n28992), .Z(n28773) );
  NANDN U29161 ( .A(n28993), .B(n28994), .Z(n28992) );
  OR U29162 ( .A(n28995), .B(n28996), .Z(n28994) );
  NAND U29163 ( .A(n28996), .B(n28995), .Z(n28991) );
  ANDN U29164 ( .B(B[178]), .A(n61), .Z(n28775) );
  XNOR U29165 ( .A(n28783), .B(n28997), .Z(n28776) );
  XNOR U29166 ( .A(n28782), .B(n28780), .Z(n28997) );
  AND U29167 ( .A(n28998), .B(n28999), .Z(n28780) );
  NANDN U29168 ( .A(n29000), .B(n29001), .Z(n28999) );
  NANDN U29169 ( .A(n29002), .B(n29003), .Z(n29001) );
  NANDN U29170 ( .A(n29003), .B(n29002), .Z(n28998) );
  ANDN U29171 ( .B(B[179]), .A(n62), .Z(n28782) );
  XNOR U29172 ( .A(n28790), .B(n29004), .Z(n28783) );
  XNOR U29173 ( .A(n28789), .B(n28787), .Z(n29004) );
  AND U29174 ( .A(n29005), .B(n29006), .Z(n28787) );
  NANDN U29175 ( .A(n29007), .B(n29008), .Z(n29006) );
  OR U29176 ( .A(n29009), .B(n29010), .Z(n29008) );
  NAND U29177 ( .A(n29010), .B(n29009), .Z(n29005) );
  ANDN U29178 ( .B(B[180]), .A(n63), .Z(n28789) );
  XNOR U29179 ( .A(n28797), .B(n29011), .Z(n28790) );
  XNOR U29180 ( .A(n28796), .B(n28794), .Z(n29011) );
  AND U29181 ( .A(n29012), .B(n29013), .Z(n28794) );
  NANDN U29182 ( .A(n29014), .B(n29015), .Z(n29013) );
  NANDN U29183 ( .A(n29016), .B(n29017), .Z(n29015) );
  NANDN U29184 ( .A(n29017), .B(n29016), .Z(n29012) );
  ANDN U29185 ( .B(B[181]), .A(n64), .Z(n28796) );
  XNOR U29186 ( .A(n28804), .B(n29018), .Z(n28797) );
  XNOR U29187 ( .A(n28803), .B(n28801), .Z(n29018) );
  AND U29188 ( .A(n29019), .B(n29020), .Z(n28801) );
  NANDN U29189 ( .A(n29021), .B(n29022), .Z(n29020) );
  OR U29190 ( .A(n29023), .B(n29024), .Z(n29022) );
  NAND U29191 ( .A(n29024), .B(n29023), .Z(n29019) );
  ANDN U29192 ( .B(B[182]), .A(n65), .Z(n28803) );
  XNOR U29193 ( .A(n28811), .B(n29025), .Z(n28804) );
  XNOR U29194 ( .A(n28810), .B(n28808), .Z(n29025) );
  AND U29195 ( .A(n29026), .B(n29027), .Z(n28808) );
  NANDN U29196 ( .A(n29028), .B(n29029), .Z(n29027) );
  NANDN U29197 ( .A(n29030), .B(n29031), .Z(n29029) );
  NANDN U29198 ( .A(n29031), .B(n29030), .Z(n29026) );
  ANDN U29199 ( .B(B[183]), .A(n66), .Z(n28810) );
  XNOR U29200 ( .A(n28818), .B(n29032), .Z(n28811) );
  XNOR U29201 ( .A(n28817), .B(n28815), .Z(n29032) );
  AND U29202 ( .A(n29033), .B(n29034), .Z(n28815) );
  NANDN U29203 ( .A(n29035), .B(n29036), .Z(n29034) );
  OR U29204 ( .A(n29037), .B(n29038), .Z(n29036) );
  NAND U29205 ( .A(n29038), .B(n29037), .Z(n29033) );
  ANDN U29206 ( .B(B[184]), .A(n67), .Z(n28817) );
  XNOR U29207 ( .A(n28825), .B(n29039), .Z(n28818) );
  XNOR U29208 ( .A(n28824), .B(n28822), .Z(n29039) );
  AND U29209 ( .A(n29040), .B(n29041), .Z(n28822) );
  NANDN U29210 ( .A(n29042), .B(n29043), .Z(n29041) );
  NANDN U29211 ( .A(n29044), .B(n29045), .Z(n29043) );
  NANDN U29212 ( .A(n29045), .B(n29044), .Z(n29040) );
  ANDN U29213 ( .B(B[185]), .A(n68), .Z(n28824) );
  XNOR U29214 ( .A(n28832), .B(n29046), .Z(n28825) );
  XNOR U29215 ( .A(n28831), .B(n28829), .Z(n29046) );
  AND U29216 ( .A(n29047), .B(n29048), .Z(n28829) );
  NANDN U29217 ( .A(n29049), .B(n29050), .Z(n29048) );
  OR U29218 ( .A(n29051), .B(n29052), .Z(n29050) );
  NAND U29219 ( .A(n29052), .B(n29051), .Z(n29047) );
  ANDN U29220 ( .B(B[186]), .A(n69), .Z(n28831) );
  XNOR U29221 ( .A(n28839), .B(n29053), .Z(n28832) );
  XNOR U29222 ( .A(n28838), .B(n28836), .Z(n29053) );
  AND U29223 ( .A(n29054), .B(n29055), .Z(n28836) );
  NANDN U29224 ( .A(n29056), .B(n29057), .Z(n29055) );
  NANDN U29225 ( .A(n29058), .B(n29059), .Z(n29057) );
  NANDN U29226 ( .A(n29059), .B(n29058), .Z(n29054) );
  ANDN U29227 ( .B(B[187]), .A(n70), .Z(n28838) );
  XNOR U29228 ( .A(n28846), .B(n29060), .Z(n28839) );
  XNOR U29229 ( .A(n28845), .B(n28843), .Z(n29060) );
  AND U29230 ( .A(n29061), .B(n29062), .Z(n28843) );
  NANDN U29231 ( .A(n29063), .B(n29064), .Z(n29062) );
  OR U29232 ( .A(n29065), .B(n29066), .Z(n29064) );
  NAND U29233 ( .A(n29066), .B(n29065), .Z(n29061) );
  ANDN U29234 ( .B(B[188]), .A(n71), .Z(n28845) );
  XNOR U29235 ( .A(n28853), .B(n29067), .Z(n28846) );
  XNOR U29236 ( .A(n28852), .B(n28850), .Z(n29067) );
  AND U29237 ( .A(n29068), .B(n29069), .Z(n28850) );
  NANDN U29238 ( .A(n29070), .B(n29071), .Z(n29069) );
  NANDN U29239 ( .A(n29072), .B(n29073), .Z(n29071) );
  NANDN U29240 ( .A(n29073), .B(n29072), .Z(n29068) );
  ANDN U29241 ( .B(B[189]), .A(n72), .Z(n28852) );
  XNOR U29242 ( .A(n28860), .B(n29074), .Z(n28853) );
  XNOR U29243 ( .A(n28859), .B(n28857), .Z(n29074) );
  AND U29244 ( .A(n29075), .B(n29076), .Z(n28857) );
  NANDN U29245 ( .A(n29077), .B(n29078), .Z(n29076) );
  OR U29246 ( .A(n29079), .B(n29080), .Z(n29078) );
  NAND U29247 ( .A(n29080), .B(n29079), .Z(n29075) );
  ANDN U29248 ( .B(B[190]), .A(n73), .Z(n28859) );
  XNOR U29249 ( .A(n28867), .B(n29081), .Z(n28860) );
  XNOR U29250 ( .A(n28866), .B(n28864), .Z(n29081) );
  AND U29251 ( .A(n29082), .B(n29083), .Z(n28864) );
  NANDN U29252 ( .A(n29084), .B(n29085), .Z(n29083) );
  NANDN U29253 ( .A(n29086), .B(n29087), .Z(n29085) );
  NANDN U29254 ( .A(n29087), .B(n29086), .Z(n29082) );
  ANDN U29255 ( .B(B[191]), .A(n74), .Z(n28866) );
  XNOR U29256 ( .A(n28874), .B(n29088), .Z(n28867) );
  XNOR U29257 ( .A(n28873), .B(n28871), .Z(n29088) );
  AND U29258 ( .A(n29089), .B(n29090), .Z(n28871) );
  NANDN U29259 ( .A(n29091), .B(n29092), .Z(n29090) );
  OR U29260 ( .A(n29093), .B(n29094), .Z(n29092) );
  NAND U29261 ( .A(n29094), .B(n29093), .Z(n29089) );
  ANDN U29262 ( .B(B[192]), .A(n75), .Z(n28873) );
  XNOR U29263 ( .A(n28881), .B(n29095), .Z(n28874) );
  XNOR U29264 ( .A(n28880), .B(n28878), .Z(n29095) );
  AND U29265 ( .A(n29096), .B(n29097), .Z(n28878) );
  NANDN U29266 ( .A(n29098), .B(n29099), .Z(n29097) );
  NANDN U29267 ( .A(n29100), .B(n29101), .Z(n29099) );
  NANDN U29268 ( .A(n29101), .B(n29100), .Z(n29096) );
  ANDN U29269 ( .B(B[193]), .A(n76), .Z(n28880) );
  XNOR U29270 ( .A(n28888), .B(n29102), .Z(n28881) );
  XNOR U29271 ( .A(n28887), .B(n28885), .Z(n29102) );
  AND U29272 ( .A(n29103), .B(n29104), .Z(n28885) );
  NANDN U29273 ( .A(n29105), .B(n29106), .Z(n29104) );
  OR U29274 ( .A(n29107), .B(n29108), .Z(n29106) );
  NAND U29275 ( .A(n29108), .B(n29107), .Z(n29103) );
  ANDN U29276 ( .B(B[194]), .A(n77), .Z(n28887) );
  XNOR U29277 ( .A(n28895), .B(n29109), .Z(n28888) );
  XNOR U29278 ( .A(n28894), .B(n28892), .Z(n29109) );
  AND U29279 ( .A(n29110), .B(n29111), .Z(n28892) );
  NANDN U29280 ( .A(n29112), .B(n29113), .Z(n29111) );
  NANDN U29281 ( .A(n29114), .B(n29115), .Z(n29113) );
  NANDN U29282 ( .A(n29115), .B(n29114), .Z(n29110) );
  ANDN U29283 ( .B(B[195]), .A(n78), .Z(n28894) );
  XNOR U29284 ( .A(n28902), .B(n29116), .Z(n28895) );
  XNOR U29285 ( .A(n28901), .B(n28899), .Z(n29116) );
  AND U29286 ( .A(n29117), .B(n29118), .Z(n28899) );
  NANDN U29287 ( .A(n29119), .B(n29120), .Z(n29118) );
  OR U29288 ( .A(n29121), .B(n29122), .Z(n29120) );
  NAND U29289 ( .A(n29122), .B(n29121), .Z(n29117) );
  ANDN U29290 ( .B(B[196]), .A(n79), .Z(n28901) );
  XNOR U29291 ( .A(n28909), .B(n29123), .Z(n28902) );
  XNOR U29292 ( .A(n28908), .B(n28906), .Z(n29123) );
  AND U29293 ( .A(n29124), .B(n29125), .Z(n28906) );
  NANDN U29294 ( .A(n29126), .B(n29127), .Z(n29125) );
  NANDN U29295 ( .A(n29128), .B(n29129), .Z(n29127) );
  NANDN U29296 ( .A(n29129), .B(n29128), .Z(n29124) );
  ANDN U29297 ( .B(B[197]), .A(n80), .Z(n28908) );
  XNOR U29298 ( .A(n28916), .B(n29130), .Z(n28909) );
  XNOR U29299 ( .A(n28915), .B(n28913), .Z(n29130) );
  AND U29300 ( .A(n29131), .B(n29132), .Z(n28913) );
  NANDN U29301 ( .A(n29133), .B(n29134), .Z(n29132) );
  OR U29302 ( .A(n29135), .B(n29136), .Z(n29134) );
  NAND U29303 ( .A(n29136), .B(n29135), .Z(n29131) );
  ANDN U29304 ( .B(B[198]), .A(n81), .Z(n28915) );
  XNOR U29305 ( .A(n28923), .B(n29137), .Z(n28916) );
  XNOR U29306 ( .A(n28922), .B(n28920), .Z(n29137) );
  AND U29307 ( .A(n29138), .B(n29139), .Z(n28920) );
  NANDN U29308 ( .A(n29140), .B(n29141), .Z(n29139) );
  NAND U29309 ( .A(n29142), .B(n29143), .Z(n29141) );
  ANDN U29310 ( .B(B[199]), .A(n82), .Z(n28922) );
  XOR U29311 ( .A(n28929), .B(n29144), .Z(n28923) );
  XNOR U29312 ( .A(n28927), .B(n28930), .Z(n29144) );
  NAND U29313 ( .A(A[2]), .B(B[200]), .Z(n28930) );
  NANDN U29314 ( .A(n29145), .B(n29146), .Z(n28927) );
  AND U29315 ( .A(A[0]), .B(B[201]), .Z(n29146) );
  XNOR U29316 ( .A(n28932), .B(n29147), .Z(n28929) );
  NAND U29317 ( .A(A[0]), .B(B[202]), .Z(n29147) );
  NAND U29318 ( .A(B[201]), .B(A[1]), .Z(n28932) );
  NAND U29319 ( .A(n29148), .B(n29149), .Z(n392) );
  NANDN U29320 ( .A(n29150), .B(n29151), .Z(n29149) );
  OR U29321 ( .A(n29152), .B(n29153), .Z(n29151) );
  NAND U29322 ( .A(n29153), .B(n29152), .Z(n29148) );
  XOR U29323 ( .A(n29154), .B(n29155), .Z(\A1[1] ) );
  XNOR U29324 ( .A(n29156), .B(n29157), .Z(n29155) );
  XOR U29325 ( .A(n26886), .B(n29158), .Z(\A1[19] ) );
  XNOR U29326 ( .A(n26885), .B(n26883), .Z(n29158) );
  AND U29327 ( .A(n29159), .B(n29160), .Z(n26883) );
  NAND U29328 ( .A(n29161), .B(n29162), .Z(n29160) );
  NANDN U29329 ( .A(n29163), .B(n29164), .Z(n29161) );
  NANDN U29330 ( .A(n29164), .B(n29163), .Z(n29159) );
  ANDN U29331 ( .B(B[0]), .A(n64), .Z(n26885) );
  XNOR U29332 ( .A(n26893), .B(n29165), .Z(n26886) );
  XNOR U29333 ( .A(n26892), .B(n26890), .Z(n29165) );
  AND U29334 ( .A(n29166), .B(n29167), .Z(n26890) );
  NANDN U29335 ( .A(n29168), .B(n29169), .Z(n29167) );
  OR U29336 ( .A(n29170), .B(n29171), .Z(n29169) );
  NAND U29337 ( .A(n29171), .B(n29170), .Z(n29166) );
  ANDN U29338 ( .B(B[1]), .A(n65), .Z(n26892) );
  XNOR U29339 ( .A(n26900), .B(n29172), .Z(n26893) );
  XNOR U29340 ( .A(n26899), .B(n26897), .Z(n29172) );
  AND U29341 ( .A(n29173), .B(n29174), .Z(n26897) );
  NANDN U29342 ( .A(n29175), .B(n29176), .Z(n29174) );
  NANDN U29343 ( .A(n29177), .B(n29178), .Z(n29176) );
  NANDN U29344 ( .A(n29178), .B(n29177), .Z(n29173) );
  ANDN U29345 ( .B(B[2]), .A(n66), .Z(n26899) );
  XNOR U29346 ( .A(n26907), .B(n29179), .Z(n26900) );
  XNOR U29347 ( .A(n26906), .B(n26904), .Z(n29179) );
  AND U29348 ( .A(n29180), .B(n29181), .Z(n26904) );
  NANDN U29349 ( .A(n29182), .B(n29183), .Z(n29181) );
  OR U29350 ( .A(n29184), .B(n29185), .Z(n29183) );
  NAND U29351 ( .A(n29185), .B(n29184), .Z(n29180) );
  ANDN U29352 ( .B(B[3]), .A(n67), .Z(n26906) );
  XNOR U29353 ( .A(n26914), .B(n29186), .Z(n26907) );
  XNOR U29354 ( .A(n26913), .B(n26911), .Z(n29186) );
  AND U29355 ( .A(n29187), .B(n29188), .Z(n26911) );
  NANDN U29356 ( .A(n29189), .B(n29190), .Z(n29188) );
  NANDN U29357 ( .A(n29191), .B(n29192), .Z(n29190) );
  NANDN U29358 ( .A(n29192), .B(n29191), .Z(n29187) );
  ANDN U29359 ( .B(B[4]), .A(n68), .Z(n26913) );
  XNOR U29360 ( .A(n26921), .B(n29193), .Z(n26914) );
  XNOR U29361 ( .A(n26920), .B(n26918), .Z(n29193) );
  AND U29362 ( .A(n29194), .B(n29195), .Z(n26918) );
  NANDN U29363 ( .A(n29196), .B(n29197), .Z(n29195) );
  OR U29364 ( .A(n29198), .B(n29199), .Z(n29197) );
  NAND U29365 ( .A(n29199), .B(n29198), .Z(n29194) );
  ANDN U29366 ( .B(B[5]), .A(n69), .Z(n26920) );
  XNOR U29367 ( .A(n26928), .B(n29200), .Z(n26921) );
  XNOR U29368 ( .A(n26927), .B(n26925), .Z(n29200) );
  AND U29369 ( .A(n29201), .B(n29202), .Z(n26925) );
  NANDN U29370 ( .A(n29203), .B(n29204), .Z(n29202) );
  NANDN U29371 ( .A(n29205), .B(n29206), .Z(n29204) );
  NANDN U29372 ( .A(n29206), .B(n29205), .Z(n29201) );
  ANDN U29373 ( .B(B[6]), .A(n70), .Z(n26927) );
  XNOR U29374 ( .A(n26935), .B(n29207), .Z(n26928) );
  XNOR U29375 ( .A(n26934), .B(n26932), .Z(n29207) );
  AND U29376 ( .A(n29208), .B(n29209), .Z(n26932) );
  NANDN U29377 ( .A(n29210), .B(n29211), .Z(n29209) );
  OR U29378 ( .A(n29212), .B(n29213), .Z(n29211) );
  NAND U29379 ( .A(n29213), .B(n29212), .Z(n29208) );
  ANDN U29380 ( .B(B[7]), .A(n71), .Z(n26934) );
  XNOR U29381 ( .A(n26942), .B(n29214), .Z(n26935) );
  XNOR U29382 ( .A(n26941), .B(n26939), .Z(n29214) );
  AND U29383 ( .A(n29215), .B(n29216), .Z(n26939) );
  NANDN U29384 ( .A(n29217), .B(n29218), .Z(n29216) );
  NANDN U29385 ( .A(n29219), .B(n29220), .Z(n29218) );
  NANDN U29386 ( .A(n29220), .B(n29219), .Z(n29215) );
  ANDN U29387 ( .B(B[8]), .A(n72), .Z(n26941) );
  XNOR U29388 ( .A(n26949), .B(n29221), .Z(n26942) );
  XNOR U29389 ( .A(n26948), .B(n26946), .Z(n29221) );
  AND U29390 ( .A(n29222), .B(n29223), .Z(n26946) );
  NANDN U29391 ( .A(n29224), .B(n29225), .Z(n29223) );
  OR U29392 ( .A(n29226), .B(n29227), .Z(n29225) );
  NAND U29393 ( .A(n29227), .B(n29226), .Z(n29222) );
  ANDN U29394 ( .B(B[9]), .A(n73), .Z(n26948) );
  XNOR U29395 ( .A(n26956), .B(n29228), .Z(n26949) );
  XNOR U29396 ( .A(n26955), .B(n26953), .Z(n29228) );
  AND U29397 ( .A(n29229), .B(n29230), .Z(n26953) );
  NANDN U29398 ( .A(n29231), .B(n29232), .Z(n29230) );
  NANDN U29399 ( .A(n29233), .B(n29234), .Z(n29232) );
  NANDN U29400 ( .A(n29234), .B(n29233), .Z(n29229) );
  ANDN U29401 ( .B(B[10]), .A(n74), .Z(n26955) );
  XNOR U29402 ( .A(n26963), .B(n29235), .Z(n26956) );
  XNOR U29403 ( .A(n26962), .B(n26960), .Z(n29235) );
  AND U29404 ( .A(n29236), .B(n29237), .Z(n26960) );
  NANDN U29405 ( .A(n29238), .B(n29239), .Z(n29237) );
  OR U29406 ( .A(n29240), .B(n29241), .Z(n29239) );
  NAND U29407 ( .A(n29241), .B(n29240), .Z(n29236) );
  ANDN U29408 ( .B(B[11]), .A(n75), .Z(n26962) );
  XNOR U29409 ( .A(n26970), .B(n29242), .Z(n26963) );
  XNOR U29410 ( .A(n26969), .B(n26967), .Z(n29242) );
  AND U29411 ( .A(n29243), .B(n29244), .Z(n26967) );
  NANDN U29412 ( .A(n29245), .B(n29246), .Z(n29244) );
  NANDN U29413 ( .A(n29247), .B(n29248), .Z(n29246) );
  NANDN U29414 ( .A(n29248), .B(n29247), .Z(n29243) );
  ANDN U29415 ( .B(B[12]), .A(n76), .Z(n26969) );
  XNOR U29416 ( .A(n26977), .B(n29249), .Z(n26970) );
  XNOR U29417 ( .A(n26976), .B(n26974), .Z(n29249) );
  AND U29418 ( .A(n29250), .B(n29251), .Z(n26974) );
  NANDN U29419 ( .A(n29252), .B(n29253), .Z(n29251) );
  OR U29420 ( .A(n29254), .B(n29255), .Z(n29253) );
  NAND U29421 ( .A(n29255), .B(n29254), .Z(n29250) );
  ANDN U29422 ( .B(B[13]), .A(n77), .Z(n26976) );
  XNOR U29423 ( .A(n26984), .B(n29256), .Z(n26977) );
  XNOR U29424 ( .A(n26983), .B(n26981), .Z(n29256) );
  AND U29425 ( .A(n29257), .B(n29258), .Z(n26981) );
  NANDN U29426 ( .A(n29259), .B(n29260), .Z(n29258) );
  NANDN U29427 ( .A(n29261), .B(n29262), .Z(n29260) );
  NANDN U29428 ( .A(n29262), .B(n29261), .Z(n29257) );
  ANDN U29429 ( .B(B[14]), .A(n78), .Z(n26983) );
  XNOR U29430 ( .A(n26991), .B(n29263), .Z(n26984) );
  XNOR U29431 ( .A(n26990), .B(n26988), .Z(n29263) );
  AND U29432 ( .A(n29264), .B(n29265), .Z(n26988) );
  NANDN U29433 ( .A(n29266), .B(n29267), .Z(n29265) );
  OR U29434 ( .A(n29268), .B(n29269), .Z(n29267) );
  NAND U29435 ( .A(n29269), .B(n29268), .Z(n29264) );
  ANDN U29436 ( .B(B[15]), .A(n79), .Z(n26990) );
  XNOR U29437 ( .A(n26998), .B(n29270), .Z(n26991) );
  XNOR U29438 ( .A(n26997), .B(n26995), .Z(n29270) );
  AND U29439 ( .A(n29271), .B(n29272), .Z(n26995) );
  NANDN U29440 ( .A(n29273), .B(n29274), .Z(n29272) );
  NANDN U29441 ( .A(n29275), .B(n29276), .Z(n29274) );
  NANDN U29442 ( .A(n29276), .B(n29275), .Z(n29271) );
  ANDN U29443 ( .B(B[16]), .A(n80), .Z(n26997) );
  XNOR U29444 ( .A(n27005), .B(n29277), .Z(n26998) );
  XNOR U29445 ( .A(n27004), .B(n27002), .Z(n29277) );
  AND U29446 ( .A(n29278), .B(n29279), .Z(n27002) );
  NANDN U29447 ( .A(n29280), .B(n29281), .Z(n29279) );
  OR U29448 ( .A(n29282), .B(n29283), .Z(n29281) );
  NAND U29449 ( .A(n29283), .B(n29282), .Z(n29278) );
  ANDN U29450 ( .B(B[17]), .A(n81), .Z(n27004) );
  XNOR U29451 ( .A(n27012), .B(n29284), .Z(n27005) );
  XNOR U29452 ( .A(n27011), .B(n27009), .Z(n29284) );
  AND U29453 ( .A(n29285), .B(n29286), .Z(n27009) );
  NANDN U29454 ( .A(n29287), .B(n29288), .Z(n29286) );
  NAND U29455 ( .A(n29289), .B(n29290), .Z(n29288) );
  ANDN U29456 ( .B(B[18]), .A(n82), .Z(n27011) );
  XOR U29457 ( .A(n27018), .B(n29291), .Z(n27012) );
  XNOR U29458 ( .A(n27016), .B(n27019), .Z(n29291) );
  NAND U29459 ( .A(A[2]), .B(B[19]), .Z(n27019) );
  NANDN U29460 ( .A(n29292), .B(n29293), .Z(n27016) );
  AND U29461 ( .A(A[0]), .B(B[20]), .Z(n29293) );
  XNOR U29462 ( .A(n27021), .B(n29294), .Z(n27018) );
  NAND U29463 ( .A(A[0]), .B(B[21]), .Z(n29294) );
  NAND U29464 ( .A(B[20]), .B(A[1]), .Z(n27021) );
  XOR U29465 ( .A(n394), .B(n393), .Z(\A1[199] ) );
  XOR U29466 ( .A(n29153), .B(n29295), .Z(n393) );
  XNOR U29467 ( .A(n29152), .B(n29150), .Z(n29295) );
  AND U29468 ( .A(n29296), .B(n29297), .Z(n29150) );
  NANDN U29469 ( .A(n29298), .B(n29299), .Z(n29297) );
  NANDN U29470 ( .A(n29300), .B(n29301), .Z(n29299) );
  NANDN U29471 ( .A(n29301), .B(n29300), .Z(n29296) );
  ANDN U29472 ( .B(B[170]), .A(n54), .Z(n29152) );
  XNOR U29473 ( .A(n28947), .B(n29302), .Z(n29153) );
  XNOR U29474 ( .A(n28946), .B(n28944), .Z(n29302) );
  AND U29475 ( .A(n29303), .B(n29304), .Z(n28944) );
  NANDN U29476 ( .A(n29305), .B(n29306), .Z(n29304) );
  OR U29477 ( .A(n29307), .B(n29308), .Z(n29306) );
  NAND U29478 ( .A(n29308), .B(n29307), .Z(n29303) );
  ANDN U29479 ( .B(B[171]), .A(n55), .Z(n28946) );
  XNOR U29480 ( .A(n28954), .B(n29309), .Z(n28947) );
  XNOR U29481 ( .A(n28953), .B(n28951), .Z(n29309) );
  AND U29482 ( .A(n29310), .B(n29311), .Z(n28951) );
  NANDN U29483 ( .A(n29312), .B(n29313), .Z(n29311) );
  NANDN U29484 ( .A(n29314), .B(n29315), .Z(n29313) );
  NANDN U29485 ( .A(n29315), .B(n29314), .Z(n29310) );
  ANDN U29486 ( .B(B[172]), .A(n56), .Z(n28953) );
  XNOR U29487 ( .A(n28961), .B(n29316), .Z(n28954) );
  XNOR U29488 ( .A(n28960), .B(n28958), .Z(n29316) );
  AND U29489 ( .A(n29317), .B(n29318), .Z(n28958) );
  NANDN U29490 ( .A(n29319), .B(n29320), .Z(n29318) );
  OR U29491 ( .A(n29321), .B(n29322), .Z(n29320) );
  NAND U29492 ( .A(n29322), .B(n29321), .Z(n29317) );
  ANDN U29493 ( .B(B[173]), .A(n57), .Z(n28960) );
  XNOR U29494 ( .A(n28968), .B(n29323), .Z(n28961) );
  XNOR U29495 ( .A(n28967), .B(n28965), .Z(n29323) );
  AND U29496 ( .A(n29324), .B(n29325), .Z(n28965) );
  NANDN U29497 ( .A(n29326), .B(n29327), .Z(n29325) );
  NANDN U29498 ( .A(n29328), .B(n29329), .Z(n29327) );
  NANDN U29499 ( .A(n29329), .B(n29328), .Z(n29324) );
  ANDN U29500 ( .B(B[174]), .A(n58), .Z(n28967) );
  XNOR U29501 ( .A(n28975), .B(n29330), .Z(n28968) );
  XNOR U29502 ( .A(n28974), .B(n28972), .Z(n29330) );
  AND U29503 ( .A(n29331), .B(n29332), .Z(n28972) );
  NANDN U29504 ( .A(n29333), .B(n29334), .Z(n29332) );
  OR U29505 ( .A(n29335), .B(n29336), .Z(n29334) );
  NAND U29506 ( .A(n29336), .B(n29335), .Z(n29331) );
  ANDN U29507 ( .B(B[175]), .A(n59), .Z(n28974) );
  XNOR U29508 ( .A(n28982), .B(n29337), .Z(n28975) );
  XNOR U29509 ( .A(n28981), .B(n28979), .Z(n29337) );
  AND U29510 ( .A(n29338), .B(n29339), .Z(n28979) );
  NANDN U29511 ( .A(n29340), .B(n29341), .Z(n29339) );
  NANDN U29512 ( .A(n29342), .B(n29343), .Z(n29341) );
  NANDN U29513 ( .A(n29343), .B(n29342), .Z(n29338) );
  ANDN U29514 ( .B(B[176]), .A(n60), .Z(n28981) );
  XNOR U29515 ( .A(n28989), .B(n29344), .Z(n28982) );
  XNOR U29516 ( .A(n28988), .B(n28986), .Z(n29344) );
  AND U29517 ( .A(n29345), .B(n29346), .Z(n28986) );
  NANDN U29518 ( .A(n29347), .B(n29348), .Z(n29346) );
  OR U29519 ( .A(n29349), .B(n29350), .Z(n29348) );
  NAND U29520 ( .A(n29350), .B(n29349), .Z(n29345) );
  ANDN U29521 ( .B(B[177]), .A(n61), .Z(n28988) );
  XNOR U29522 ( .A(n28996), .B(n29351), .Z(n28989) );
  XNOR U29523 ( .A(n28995), .B(n28993), .Z(n29351) );
  AND U29524 ( .A(n29352), .B(n29353), .Z(n28993) );
  NANDN U29525 ( .A(n29354), .B(n29355), .Z(n29353) );
  NANDN U29526 ( .A(n29356), .B(n29357), .Z(n29355) );
  NANDN U29527 ( .A(n29357), .B(n29356), .Z(n29352) );
  ANDN U29528 ( .B(B[178]), .A(n62), .Z(n28995) );
  XNOR U29529 ( .A(n29003), .B(n29358), .Z(n28996) );
  XNOR U29530 ( .A(n29002), .B(n29000), .Z(n29358) );
  AND U29531 ( .A(n29359), .B(n29360), .Z(n29000) );
  NANDN U29532 ( .A(n29361), .B(n29362), .Z(n29360) );
  OR U29533 ( .A(n29363), .B(n29364), .Z(n29362) );
  NAND U29534 ( .A(n29364), .B(n29363), .Z(n29359) );
  ANDN U29535 ( .B(B[179]), .A(n63), .Z(n29002) );
  XNOR U29536 ( .A(n29010), .B(n29365), .Z(n29003) );
  XNOR U29537 ( .A(n29009), .B(n29007), .Z(n29365) );
  AND U29538 ( .A(n29366), .B(n29367), .Z(n29007) );
  NANDN U29539 ( .A(n29368), .B(n29369), .Z(n29367) );
  NANDN U29540 ( .A(n29370), .B(n29371), .Z(n29369) );
  NANDN U29541 ( .A(n29371), .B(n29370), .Z(n29366) );
  ANDN U29542 ( .B(B[180]), .A(n64), .Z(n29009) );
  XNOR U29543 ( .A(n29017), .B(n29372), .Z(n29010) );
  XNOR U29544 ( .A(n29016), .B(n29014), .Z(n29372) );
  AND U29545 ( .A(n29373), .B(n29374), .Z(n29014) );
  NANDN U29546 ( .A(n29375), .B(n29376), .Z(n29374) );
  OR U29547 ( .A(n29377), .B(n29378), .Z(n29376) );
  NAND U29548 ( .A(n29378), .B(n29377), .Z(n29373) );
  ANDN U29549 ( .B(B[181]), .A(n65), .Z(n29016) );
  XNOR U29550 ( .A(n29024), .B(n29379), .Z(n29017) );
  XNOR U29551 ( .A(n29023), .B(n29021), .Z(n29379) );
  AND U29552 ( .A(n29380), .B(n29381), .Z(n29021) );
  NANDN U29553 ( .A(n29382), .B(n29383), .Z(n29381) );
  NANDN U29554 ( .A(n29384), .B(n29385), .Z(n29383) );
  NANDN U29555 ( .A(n29385), .B(n29384), .Z(n29380) );
  ANDN U29556 ( .B(B[182]), .A(n66), .Z(n29023) );
  XNOR U29557 ( .A(n29031), .B(n29386), .Z(n29024) );
  XNOR U29558 ( .A(n29030), .B(n29028), .Z(n29386) );
  AND U29559 ( .A(n29387), .B(n29388), .Z(n29028) );
  NANDN U29560 ( .A(n29389), .B(n29390), .Z(n29388) );
  OR U29561 ( .A(n29391), .B(n29392), .Z(n29390) );
  NAND U29562 ( .A(n29392), .B(n29391), .Z(n29387) );
  ANDN U29563 ( .B(B[183]), .A(n67), .Z(n29030) );
  XNOR U29564 ( .A(n29038), .B(n29393), .Z(n29031) );
  XNOR U29565 ( .A(n29037), .B(n29035), .Z(n29393) );
  AND U29566 ( .A(n29394), .B(n29395), .Z(n29035) );
  NANDN U29567 ( .A(n29396), .B(n29397), .Z(n29395) );
  NANDN U29568 ( .A(n29398), .B(n29399), .Z(n29397) );
  NANDN U29569 ( .A(n29399), .B(n29398), .Z(n29394) );
  ANDN U29570 ( .B(B[184]), .A(n68), .Z(n29037) );
  XNOR U29571 ( .A(n29045), .B(n29400), .Z(n29038) );
  XNOR U29572 ( .A(n29044), .B(n29042), .Z(n29400) );
  AND U29573 ( .A(n29401), .B(n29402), .Z(n29042) );
  NANDN U29574 ( .A(n29403), .B(n29404), .Z(n29402) );
  OR U29575 ( .A(n29405), .B(n29406), .Z(n29404) );
  NAND U29576 ( .A(n29406), .B(n29405), .Z(n29401) );
  ANDN U29577 ( .B(B[185]), .A(n69), .Z(n29044) );
  XNOR U29578 ( .A(n29052), .B(n29407), .Z(n29045) );
  XNOR U29579 ( .A(n29051), .B(n29049), .Z(n29407) );
  AND U29580 ( .A(n29408), .B(n29409), .Z(n29049) );
  NANDN U29581 ( .A(n29410), .B(n29411), .Z(n29409) );
  NANDN U29582 ( .A(n29412), .B(n29413), .Z(n29411) );
  NANDN U29583 ( .A(n29413), .B(n29412), .Z(n29408) );
  ANDN U29584 ( .B(B[186]), .A(n70), .Z(n29051) );
  XNOR U29585 ( .A(n29059), .B(n29414), .Z(n29052) );
  XNOR U29586 ( .A(n29058), .B(n29056), .Z(n29414) );
  AND U29587 ( .A(n29415), .B(n29416), .Z(n29056) );
  NANDN U29588 ( .A(n29417), .B(n29418), .Z(n29416) );
  OR U29589 ( .A(n29419), .B(n29420), .Z(n29418) );
  NAND U29590 ( .A(n29420), .B(n29419), .Z(n29415) );
  ANDN U29591 ( .B(B[187]), .A(n71), .Z(n29058) );
  XNOR U29592 ( .A(n29066), .B(n29421), .Z(n29059) );
  XNOR U29593 ( .A(n29065), .B(n29063), .Z(n29421) );
  AND U29594 ( .A(n29422), .B(n29423), .Z(n29063) );
  NANDN U29595 ( .A(n29424), .B(n29425), .Z(n29423) );
  NANDN U29596 ( .A(n29426), .B(n29427), .Z(n29425) );
  NANDN U29597 ( .A(n29427), .B(n29426), .Z(n29422) );
  ANDN U29598 ( .B(B[188]), .A(n72), .Z(n29065) );
  XNOR U29599 ( .A(n29073), .B(n29428), .Z(n29066) );
  XNOR U29600 ( .A(n29072), .B(n29070), .Z(n29428) );
  AND U29601 ( .A(n29429), .B(n29430), .Z(n29070) );
  NANDN U29602 ( .A(n29431), .B(n29432), .Z(n29430) );
  OR U29603 ( .A(n29433), .B(n29434), .Z(n29432) );
  NAND U29604 ( .A(n29434), .B(n29433), .Z(n29429) );
  ANDN U29605 ( .B(B[189]), .A(n73), .Z(n29072) );
  XNOR U29606 ( .A(n29080), .B(n29435), .Z(n29073) );
  XNOR U29607 ( .A(n29079), .B(n29077), .Z(n29435) );
  AND U29608 ( .A(n29436), .B(n29437), .Z(n29077) );
  NANDN U29609 ( .A(n29438), .B(n29439), .Z(n29437) );
  NANDN U29610 ( .A(n29440), .B(n29441), .Z(n29439) );
  NANDN U29611 ( .A(n29441), .B(n29440), .Z(n29436) );
  ANDN U29612 ( .B(B[190]), .A(n74), .Z(n29079) );
  XNOR U29613 ( .A(n29087), .B(n29442), .Z(n29080) );
  XNOR U29614 ( .A(n29086), .B(n29084), .Z(n29442) );
  AND U29615 ( .A(n29443), .B(n29444), .Z(n29084) );
  NANDN U29616 ( .A(n29445), .B(n29446), .Z(n29444) );
  OR U29617 ( .A(n29447), .B(n29448), .Z(n29446) );
  NAND U29618 ( .A(n29448), .B(n29447), .Z(n29443) );
  ANDN U29619 ( .B(B[191]), .A(n75), .Z(n29086) );
  XNOR U29620 ( .A(n29094), .B(n29449), .Z(n29087) );
  XNOR U29621 ( .A(n29093), .B(n29091), .Z(n29449) );
  AND U29622 ( .A(n29450), .B(n29451), .Z(n29091) );
  NANDN U29623 ( .A(n29452), .B(n29453), .Z(n29451) );
  NANDN U29624 ( .A(n29454), .B(n29455), .Z(n29453) );
  NANDN U29625 ( .A(n29455), .B(n29454), .Z(n29450) );
  ANDN U29626 ( .B(B[192]), .A(n76), .Z(n29093) );
  XNOR U29627 ( .A(n29101), .B(n29456), .Z(n29094) );
  XNOR U29628 ( .A(n29100), .B(n29098), .Z(n29456) );
  AND U29629 ( .A(n29457), .B(n29458), .Z(n29098) );
  NANDN U29630 ( .A(n29459), .B(n29460), .Z(n29458) );
  OR U29631 ( .A(n29461), .B(n29462), .Z(n29460) );
  NAND U29632 ( .A(n29462), .B(n29461), .Z(n29457) );
  ANDN U29633 ( .B(B[193]), .A(n77), .Z(n29100) );
  XNOR U29634 ( .A(n29108), .B(n29463), .Z(n29101) );
  XNOR U29635 ( .A(n29107), .B(n29105), .Z(n29463) );
  AND U29636 ( .A(n29464), .B(n29465), .Z(n29105) );
  NANDN U29637 ( .A(n29466), .B(n29467), .Z(n29465) );
  NANDN U29638 ( .A(n29468), .B(n29469), .Z(n29467) );
  NANDN U29639 ( .A(n29469), .B(n29468), .Z(n29464) );
  ANDN U29640 ( .B(B[194]), .A(n78), .Z(n29107) );
  XNOR U29641 ( .A(n29115), .B(n29470), .Z(n29108) );
  XNOR U29642 ( .A(n29114), .B(n29112), .Z(n29470) );
  AND U29643 ( .A(n29471), .B(n29472), .Z(n29112) );
  NANDN U29644 ( .A(n29473), .B(n29474), .Z(n29472) );
  OR U29645 ( .A(n29475), .B(n29476), .Z(n29474) );
  NAND U29646 ( .A(n29476), .B(n29475), .Z(n29471) );
  ANDN U29647 ( .B(B[195]), .A(n79), .Z(n29114) );
  XNOR U29648 ( .A(n29122), .B(n29477), .Z(n29115) );
  XNOR U29649 ( .A(n29121), .B(n29119), .Z(n29477) );
  AND U29650 ( .A(n29478), .B(n29479), .Z(n29119) );
  NANDN U29651 ( .A(n29480), .B(n29481), .Z(n29479) );
  NANDN U29652 ( .A(n29482), .B(n29483), .Z(n29481) );
  NANDN U29653 ( .A(n29483), .B(n29482), .Z(n29478) );
  ANDN U29654 ( .B(B[196]), .A(n80), .Z(n29121) );
  XNOR U29655 ( .A(n29129), .B(n29484), .Z(n29122) );
  XNOR U29656 ( .A(n29128), .B(n29126), .Z(n29484) );
  AND U29657 ( .A(n29485), .B(n29486), .Z(n29126) );
  NANDN U29658 ( .A(n29487), .B(n29488), .Z(n29486) );
  OR U29659 ( .A(n29489), .B(n29490), .Z(n29488) );
  NAND U29660 ( .A(n29490), .B(n29489), .Z(n29485) );
  ANDN U29661 ( .B(B[197]), .A(n81), .Z(n29128) );
  XNOR U29662 ( .A(n29136), .B(n29491), .Z(n29129) );
  XNOR U29663 ( .A(n29135), .B(n29133), .Z(n29491) );
  AND U29664 ( .A(n29492), .B(n29493), .Z(n29133) );
  NANDN U29665 ( .A(n29494), .B(n29495), .Z(n29493) );
  NAND U29666 ( .A(n29496), .B(n29497), .Z(n29495) );
  ANDN U29667 ( .B(B[198]), .A(n82), .Z(n29135) );
  XOR U29668 ( .A(n29142), .B(n29498), .Z(n29136) );
  XNOR U29669 ( .A(n29140), .B(n29143), .Z(n29498) );
  NAND U29670 ( .A(A[2]), .B(B[199]), .Z(n29143) );
  NANDN U29671 ( .A(n29499), .B(n29500), .Z(n29140) );
  AND U29672 ( .A(A[0]), .B(B[200]), .Z(n29500) );
  XNOR U29673 ( .A(n29145), .B(n29501), .Z(n29142) );
  NAND U29674 ( .A(A[0]), .B(B[201]), .Z(n29501) );
  NAND U29675 ( .A(B[200]), .B(A[1]), .Z(n29145) );
  NAND U29676 ( .A(n29502), .B(n29503), .Z(n394) );
  NANDN U29677 ( .A(n29504), .B(n29505), .Z(n29503) );
  OR U29678 ( .A(n29506), .B(n29507), .Z(n29505) );
  NAND U29679 ( .A(n29507), .B(n29506), .Z(n29502) );
  XOR U29680 ( .A(n396), .B(n395), .Z(\A1[198] ) );
  XOR U29681 ( .A(n29507), .B(n29508), .Z(n395) );
  XNOR U29682 ( .A(n29506), .B(n29504), .Z(n29508) );
  AND U29683 ( .A(n29509), .B(n29510), .Z(n29504) );
  NANDN U29684 ( .A(n29511), .B(n29512), .Z(n29510) );
  NANDN U29685 ( .A(n29513), .B(n29514), .Z(n29512) );
  NANDN U29686 ( .A(n29514), .B(n29513), .Z(n29509) );
  ANDN U29687 ( .B(B[169]), .A(n54), .Z(n29506) );
  XNOR U29688 ( .A(n29301), .B(n29515), .Z(n29507) );
  XNOR U29689 ( .A(n29300), .B(n29298), .Z(n29515) );
  AND U29690 ( .A(n29516), .B(n29517), .Z(n29298) );
  NANDN U29691 ( .A(n29518), .B(n29519), .Z(n29517) );
  OR U29692 ( .A(n29520), .B(n29521), .Z(n29519) );
  NAND U29693 ( .A(n29521), .B(n29520), .Z(n29516) );
  ANDN U29694 ( .B(B[170]), .A(n55), .Z(n29300) );
  XNOR U29695 ( .A(n29308), .B(n29522), .Z(n29301) );
  XNOR U29696 ( .A(n29307), .B(n29305), .Z(n29522) );
  AND U29697 ( .A(n29523), .B(n29524), .Z(n29305) );
  NANDN U29698 ( .A(n29525), .B(n29526), .Z(n29524) );
  NANDN U29699 ( .A(n29527), .B(n29528), .Z(n29526) );
  NANDN U29700 ( .A(n29528), .B(n29527), .Z(n29523) );
  ANDN U29701 ( .B(B[171]), .A(n56), .Z(n29307) );
  XNOR U29702 ( .A(n29315), .B(n29529), .Z(n29308) );
  XNOR U29703 ( .A(n29314), .B(n29312), .Z(n29529) );
  AND U29704 ( .A(n29530), .B(n29531), .Z(n29312) );
  NANDN U29705 ( .A(n29532), .B(n29533), .Z(n29531) );
  OR U29706 ( .A(n29534), .B(n29535), .Z(n29533) );
  NAND U29707 ( .A(n29535), .B(n29534), .Z(n29530) );
  ANDN U29708 ( .B(B[172]), .A(n57), .Z(n29314) );
  XNOR U29709 ( .A(n29322), .B(n29536), .Z(n29315) );
  XNOR U29710 ( .A(n29321), .B(n29319), .Z(n29536) );
  AND U29711 ( .A(n29537), .B(n29538), .Z(n29319) );
  NANDN U29712 ( .A(n29539), .B(n29540), .Z(n29538) );
  NANDN U29713 ( .A(n29541), .B(n29542), .Z(n29540) );
  NANDN U29714 ( .A(n29542), .B(n29541), .Z(n29537) );
  ANDN U29715 ( .B(B[173]), .A(n58), .Z(n29321) );
  XNOR U29716 ( .A(n29329), .B(n29543), .Z(n29322) );
  XNOR U29717 ( .A(n29328), .B(n29326), .Z(n29543) );
  AND U29718 ( .A(n29544), .B(n29545), .Z(n29326) );
  NANDN U29719 ( .A(n29546), .B(n29547), .Z(n29545) );
  OR U29720 ( .A(n29548), .B(n29549), .Z(n29547) );
  NAND U29721 ( .A(n29549), .B(n29548), .Z(n29544) );
  ANDN U29722 ( .B(B[174]), .A(n59), .Z(n29328) );
  XNOR U29723 ( .A(n29336), .B(n29550), .Z(n29329) );
  XNOR U29724 ( .A(n29335), .B(n29333), .Z(n29550) );
  AND U29725 ( .A(n29551), .B(n29552), .Z(n29333) );
  NANDN U29726 ( .A(n29553), .B(n29554), .Z(n29552) );
  NANDN U29727 ( .A(n29555), .B(n29556), .Z(n29554) );
  NANDN U29728 ( .A(n29556), .B(n29555), .Z(n29551) );
  ANDN U29729 ( .B(B[175]), .A(n60), .Z(n29335) );
  XNOR U29730 ( .A(n29343), .B(n29557), .Z(n29336) );
  XNOR U29731 ( .A(n29342), .B(n29340), .Z(n29557) );
  AND U29732 ( .A(n29558), .B(n29559), .Z(n29340) );
  NANDN U29733 ( .A(n29560), .B(n29561), .Z(n29559) );
  OR U29734 ( .A(n29562), .B(n29563), .Z(n29561) );
  NAND U29735 ( .A(n29563), .B(n29562), .Z(n29558) );
  ANDN U29736 ( .B(B[176]), .A(n61), .Z(n29342) );
  XNOR U29737 ( .A(n29350), .B(n29564), .Z(n29343) );
  XNOR U29738 ( .A(n29349), .B(n29347), .Z(n29564) );
  AND U29739 ( .A(n29565), .B(n29566), .Z(n29347) );
  NANDN U29740 ( .A(n29567), .B(n29568), .Z(n29566) );
  NANDN U29741 ( .A(n29569), .B(n29570), .Z(n29568) );
  NANDN U29742 ( .A(n29570), .B(n29569), .Z(n29565) );
  ANDN U29743 ( .B(B[177]), .A(n62), .Z(n29349) );
  XNOR U29744 ( .A(n29357), .B(n29571), .Z(n29350) );
  XNOR U29745 ( .A(n29356), .B(n29354), .Z(n29571) );
  AND U29746 ( .A(n29572), .B(n29573), .Z(n29354) );
  NANDN U29747 ( .A(n29574), .B(n29575), .Z(n29573) );
  OR U29748 ( .A(n29576), .B(n29577), .Z(n29575) );
  NAND U29749 ( .A(n29577), .B(n29576), .Z(n29572) );
  ANDN U29750 ( .B(B[178]), .A(n63), .Z(n29356) );
  XNOR U29751 ( .A(n29364), .B(n29578), .Z(n29357) );
  XNOR U29752 ( .A(n29363), .B(n29361), .Z(n29578) );
  AND U29753 ( .A(n29579), .B(n29580), .Z(n29361) );
  NANDN U29754 ( .A(n29581), .B(n29582), .Z(n29580) );
  NANDN U29755 ( .A(n29583), .B(n29584), .Z(n29582) );
  NANDN U29756 ( .A(n29584), .B(n29583), .Z(n29579) );
  ANDN U29757 ( .B(B[179]), .A(n64), .Z(n29363) );
  XNOR U29758 ( .A(n29371), .B(n29585), .Z(n29364) );
  XNOR U29759 ( .A(n29370), .B(n29368), .Z(n29585) );
  AND U29760 ( .A(n29586), .B(n29587), .Z(n29368) );
  NANDN U29761 ( .A(n29588), .B(n29589), .Z(n29587) );
  OR U29762 ( .A(n29590), .B(n29591), .Z(n29589) );
  NAND U29763 ( .A(n29591), .B(n29590), .Z(n29586) );
  ANDN U29764 ( .B(B[180]), .A(n65), .Z(n29370) );
  XNOR U29765 ( .A(n29378), .B(n29592), .Z(n29371) );
  XNOR U29766 ( .A(n29377), .B(n29375), .Z(n29592) );
  AND U29767 ( .A(n29593), .B(n29594), .Z(n29375) );
  NANDN U29768 ( .A(n29595), .B(n29596), .Z(n29594) );
  NANDN U29769 ( .A(n29597), .B(n29598), .Z(n29596) );
  NANDN U29770 ( .A(n29598), .B(n29597), .Z(n29593) );
  ANDN U29771 ( .B(B[181]), .A(n66), .Z(n29377) );
  XNOR U29772 ( .A(n29385), .B(n29599), .Z(n29378) );
  XNOR U29773 ( .A(n29384), .B(n29382), .Z(n29599) );
  AND U29774 ( .A(n29600), .B(n29601), .Z(n29382) );
  NANDN U29775 ( .A(n29602), .B(n29603), .Z(n29601) );
  OR U29776 ( .A(n29604), .B(n29605), .Z(n29603) );
  NAND U29777 ( .A(n29605), .B(n29604), .Z(n29600) );
  ANDN U29778 ( .B(B[182]), .A(n67), .Z(n29384) );
  XNOR U29779 ( .A(n29392), .B(n29606), .Z(n29385) );
  XNOR U29780 ( .A(n29391), .B(n29389), .Z(n29606) );
  AND U29781 ( .A(n29607), .B(n29608), .Z(n29389) );
  NANDN U29782 ( .A(n29609), .B(n29610), .Z(n29608) );
  NANDN U29783 ( .A(n29611), .B(n29612), .Z(n29610) );
  NANDN U29784 ( .A(n29612), .B(n29611), .Z(n29607) );
  ANDN U29785 ( .B(B[183]), .A(n68), .Z(n29391) );
  XNOR U29786 ( .A(n29399), .B(n29613), .Z(n29392) );
  XNOR U29787 ( .A(n29398), .B(n29396), .Z(n29613) );
  AND U29788 ( .A(n29614), .B(n29615), .Z(n29396) );
  NANDN U29789 ( .A(n29616), .B(n29617), .Z(n29615) );
  OR U29790 ( .A(n29618), .B(n29619), .Z(n29617) );
  NAND U29791 ( .A(n29619), .B(n29618), .Z(n29614) );
  ANDN U29792 ( .B(B[184]), .A(n69), .Z(n29398) );
  XNOR U29793 ( .A(n29406), .B(n29620), .Z(n29399) );
  XNOR U29794 ( .A(n29405), .B(n29403), .Z(n29620) );
  AND U29795 ( .A(n29621), .B(n29622), .Z(n29403) );
  NANDN U29796 ( .A(n29623), .B(n29624), .Z(n29622) );
  NANDN U29797 ( .A(n29625), .B(n29626), .Z(n29624) );
  NANDN U29798 ( .A(n29626), .B(n29625), .Z(n29621) );
  ANDN U29799 ( .B(B[185]), .A(n70), .Z(n29405) );
  XNOR U29800 ( .A(n29413), .B(n29627), .Z(n29406) );
  XNOR U29801 ( .A(n29412), .B(n29410), .Z(n29627) );
  AND U29802 ( .A(n29628), .B(n29629), .Z(n29410) );
  NANDN U29803 ( .A(n29630), .B(n29631), .Z(n29629) );
  OR U29804 ( .A(n29632), .B(n29633), .Z(n29631) );
  NAND U29805 ( .A(n29633), .B(n29632), .Z(n29628) );
  ANDN U29806 ( .B(B[186]), .A(n71), .Z(n29412) );
  XNOR U29807 ( .A(n29420), .B(n29634), .Z(n29413) );
  XNOR U29808 ( .A(n29419), .B(n29417), .Z(n29634) );
  AND U29809 ( .A(n29635), .B(n29636), .Z(n29417) );
  NANDN U29810 ( .A(n29637), .B(n29638), .Z(n29636) );
  NANDN U29811 ( .A(n29639), .B(n29640), .Z(n29638) );
  NANDN U29812 ( .A(n29640), .B(n29639), .Z(n29635) );
  ANDN U29813 ( .B(B[187]), .A(n72), .Z(n29419) );
  XNOR U29814 ( .A(n29427), .B(n29641), .Z(n29420) );
  XNOR U29815 ( .A(n29426), .B(n29424), .Z(n29641) );
  AND U29816 ( .A(n29642), .B(n29643), .Z(n29424) );
  NANDN U29817 ( .A(n29644), .B(n29645), .Z(n29643) );
  OR U29818 ( .A(n29646), .B(n29647), .Z(n29645) );
  NAND U29819 ( .A(n29647), .B(n29646), .Z(n29642) );
  ANDN U29820 ( .B(B[188]), .A(n73), .Z(n29426) );
  XNOR U29821 ( .A(n29434), .B(n29648), .Z(n29427) );
  XNOR U29822 ( .A(n29433), .B(n29431), .Z(n29648) );
  AND U29823 ( .A(n29649), .B(n29650), .Z(n29431) );
  NANDN U29824 ( .A(n29651), .B(n29652), .Z(n29650) );
  NANDN U29825 ( .A(n29653), .B(n29654), .Z(n29652) );
  NANDN U29826 ( .A(n29654), .B(n29653), .Z(n29649) );
  ANDN U29827 ( .B(B[189]), .A(n74), .Z(n29433) );
  XNOR U29828 ( .A(n29441), .B(n29655), .Z(n29434) );
  XNOR U29829 ( .A(n29440), .B(n29438), .Z(n29655) );
  AND U29830 ( .A(n29656), .B(n29657), .Z(n29438) );
  NANDN U29831 ( .A(n29658), .B(n29659), .Z(n29657) );
  OR U29832 ( .A(n29660), .B(n29661), .Z(n29659) );
  NAND U29833 ( .A(n29661), .B(n29660), .Z(n29656) );
  ANDN U29834 ( .B(B[190]), .A(n75), .Z(n29440) );
  XNOR U29835 ( .A(n29448), .B(n29662), .Z(n29441) );
  XNOR U29836 ( .A(n29447), .B(n29445), .Z(n29662) );
  AND U29837 ( .A(n29663), .B(n29664), .Z(n29445) );
  NANDN U29838 ( .A(n29665), .B(n29666), .Z(n29664) );
  NANDN U29839 ( .A(n29667), .B(n29668), .Z(n29666) );
  NANDN U29840 ( .A(n29668), .B(n29667), .Z(n29663) );
  ANDN U29841 ( .B(B[191]), .A(n76), .Z(n29447) );
  XNOR U29842 ( .A(n29455), .B(n29669), .Z(n29448) );
  XNOR U29843 ( .A(n29454), .B(n29452), .Z(n29669) );
  AND U29844 ( .A(n29670), .B(n29671), .Z(n29452) );
  NANDN U29845 ( .A(n29672), .B(n29673), .Z(n29671) );
  OR U29846 ( .A(n29674), .B(n29675), .Z(n29673) );
  NAND U29847 ( .A(n29675), .B(n29674), .Z(n29670) );
  ANDN U29848 ( .B(B[192]), .A(n77), .Z(n29454) );
  XNOR U29849 ( .A(n29462), .B(n29676), .Z(n29455) );
  XNOR U29850 ( .A(n29461), .B(n29459), .Z(n29676) );
  AND U29851 ( .A(n29677), .B(n29678), .Z(n29459) );
  NANDN U29852 ( .A(n29679), .B(n29680), .Z(n29678) );
  NANDN U29853 ( .A(n29681), .B(n29682), .Z(n29680) );
  NANDN U29854 ( .A(n29682), .B(n29681), .Z(n29677) );
  ANDN U29855 ( .B(B[193]), .A(n78), .Z(n29461) );
  XNOR U29856 ( .A(n29469), .B(n29683), .Z(n29462) );
  XNOR U29857 ( .A(n29468), .B(n29466), .Z(n29683) );
  AND U29858 ( .A(n29684), .B(n29685), .Z(n29466) );
  NANDN U29859 ( .A(n29686), .B(n29687), .Z(n29685) );
  OR U29860 ( .A(n29688), .B(n29689), .Z(n29687) );
  NAND U29861 ( .A(n29689), .B(n29688), .Z(n29684) );
  ANDN U29862 ( .B(B[194]), .A(n79), .Z(n29468) );
  XNOR U29863 ( .A(n29476), .B(n29690), .Z(n29469) );
  XNOR U29864 ( .A(n29475), .B(n29473), .Z(n29690) );
  AND U29865 ( .A(n29691), .B(n29692), .Z(n29473) );
  NANDN U29866 ( .A(n29693), .B(n29694), .Z(n29692) );
  NANDN U29867 ( .A(n29695), .B(n29696), .Z(n29694) );
  NANDN U29868 ( .A(n29696), .B(n29695), .Z(n29691) );
  ANDN U29869 ( .B(B[195]), .A(n80), .Z(n29475) );
  XNOR U29870 ( .A(n29483), .B(n29697), .Z(n29476) );
  XNOR U29871 ( .A(n29482), .B(n29480), .Z(n29697) );
  AND U29872 ( .A(n29698), .B(n29699), .Z(n29480) );
  NANDN U29873 ( .A(n29700), .B(n29701), .Z(n29699) );
  OR U29874 ( .A(n29702), .B(n29703), .Z(n29701) );
  NAND U29875 ( .A(n29703), .B(n29702), .Z(n29698) );
  ANDN U29876 ( .B(B[196]), .A(n81), .Z(n29482) );
  XNOR U29877 ( .A(n29490), .B(n29704), .Z(n29483) );
  XNOR U29878 ( .A(n29489), .B(n29487), .Z(n29704) );
  AND U29879 ( .A(n29705), .B(n29706), .Z(n29487) );
  NANDN U29880 ( .A(n29707), .B(n29708), .Z(n29706) );
  NAND U29881 ( .A(n29709), .B(n29710), .Z(n29708) );
  ANDN U29882 ( .B(B[197]), .A(n82), .Z(n29489) );
  XOR U29883 ( .A(n29496), .B(n29711), .Z(n29490) );
  XNOR U29884 ( .A(n29494), .B(n29497), .Z(n29711) );
  NAND U29885 ( .A(A[2]), .B(B[198]), .Z(n29497) );
  NANDN U29886 ( .A(n29712), .B(n29713), .Z(n29494) );
  AND U29887 ( .A(A[0]), .B(B[199]), .Z(n29713) );
  XNOR U29888 ( .A(n29499), .B(n29714), .Z(n29496) );
  NAND U29889 ( .A(A[0]), .B(B[200]), .Z(n29714) );
  NAND U29890 ( .A(B[199]), .B(A[1]), .Z(n29499) );
  NAND U29891 ( .A(n29715), .B(n29716), .Z(n396) );
  NANDN U29892 ( .A(n29717), .B(n29718), .Z(n29716) );
  OR U29893 ( .A(n29719), .B(n29720), .Z(n29718) );
  NAND U29894 ( .A(n29720), .B(n29719), .Z(n29715) );
  XOR U29895 ( .A(n398), .B(n397), .Z(\A1[197] ) );
  XOR U29896 ( .A(n29720), .B(n29721), .Z(n397) );
  XNOR U29897 ( .A(n29719), .B(n29717), .Z(n29721) );
  AND U29898 ( .A(n29722), .B(n29723), .Z(n29717) );
  NANDN U29899 ( .A(n29724), .B(n29725), .Z(n29723) );
  NANDN U29900 ( .A(n29726), .B(n29727), .Z(n29725) );
  NANDN U29901 ( .A(n29727), .B(n29726), .Z(n29722) );
  ANDN U29902 ( .B(B[168]), .A(n54), .Z(n29719) );
  XNOR U29903 ( .A(n29514), .B(n29728), .Z(n29720) );
  XNOR U29904 ( .A(n29513), .B(n29511), .Z(n29728) );
  AND U29905 ( .A(n29729), .B(n29730), .Z(n29511) );
  NANDN U29906 ( .A(n29731), .B(n29732), .Z(n29730) );
  OR U29907 ( .A(n29733), .B(n29734), .Z(n29732) );
  NAND U29908 ( .A(n29734), .B(n29733), .Z(n29729) );
  ANDN U29909 ( .B(B[169]), .A(n55), .Z(n29513) );
  XNOR U29910 ( .A(n29521), .B(n29735), .Z(n29514) );
  XNOR U29911 ( .A(n29520), .B(n29518), .Z(n29735) );
  AND U29912 ( .A(n29736), .B(n29737), .Z(n29518) );
  NANDN U29913 ( .A(n29738), .B(n29739), .Z(n29737) );
  NANDN U29914 ( .A(n29740), .B(n29741), .Z(n29739) );
  NANDN U29915 ( .A(n29741), .B(n29740), .Z(n29736) );
  ANDN U29916 ( .B(B[170]), .A(n56), .Z(n29520) );
  XNOR U29917 ( .A(n29528), .B(n29742), .Z(n29521) );
  XNOR U29918 ( .A(n29527), .B(n29525), .Z(n29742) );
  AND U29919 ( .A(n29743), .B(n29744), .Z(n29525) );
  NANDN U29920 ( .A(n29745), .B(n29746), .Z(n29744) );
  OR U29921 ( .A(n29747), .B(n29748), .Z(n29746) );
  NAND U29922 ( .A(n29748), .B(n29747), .Z(n29743) );
  ANDN U29923 ( .B(B[171]), .A(n57), .Z(n29527) );
  XNOR U29924 ( .A(n29535), .B(n29749), .Z(n29528) );
  XNOR U29925 ( .A(n29534), .B(n29532), .Z(n29749) );
  AND U29926 ( .A(n29750), .B(n29751), .Z(n29532) );
  NANDN U29927 ( .A(n29752), .B(n29753), .Z(n29751) );
  NANDN U29928 ( .A(n29754), .B(n29755), .Z(n29753) );
  NANDN U29929 ( .A(n29755), .B(n29754), .Z(n29750) );
  ANDN U29930 ( .B(B[172]), .A(n58), .Z(n29534) );
  XNOR U29931 ( .A(n29542), .B(n29756), .Z(n29535) );
  XNOR U29932 ( .A(n29541), .B(n29539), .Z(n29756) );
  AND U29933 ( .A(n29757), .B(n29758), .Z(n29539) );
  NANDN U29934 ( .A(n29759), .B(n29760), .Z(n29758) );
  OR U29935 ( .A(n29761), .B(n29762), .Z(n29760) );
  NAND U29936 ( .A(n29762), .B(n29761), .Z(n29757) );
  ANDN U29937 ( .B(B[173]), .A(n59), .Z(n29541) );
  XNOR U29938 ( .A(n29549), .B(n29763), .Z(n29542) );
  XNOR U29939 ( .A(n29548), .B(n29546), .Z(n29763) );
  AND U29940 ( .A(n29764), .B(n29765), .Z(n29546) );
  NANDN U29941 ( .A(n29766), .B(n29767), .Z(n29765) );
  NANDN U29942 ( .A(n29768), .B(n29769), .Z(n29767) );
  NANDN U29943 ( .A(n29769), .B(n29768), .Z(n29764) );
  ANDN U29944 ( .B(B[174]), .A(n60), .Z(n29548) );
  XNOR U29945 ( .A(n29556), .B(n29770), .Z(n29549) );
  XNOR U29946 ( .A(n29555), .B(n29553), .Z(n29770) );
  AND U29947 ( .A(n29771), .B(n29772), .Z(n29553) );
  NANDN U29948 ( .A(n29773), .B(n29774), .Z(n29772) );
  OR U29949 ( .A(n29775), .B(n29776), .Z(n29774) );
  NAND U29950 ( .A(n29776), .B(n29775), .Z(n29771) );
  ANDN U29951 ( .B(B[175]), .A(n61), .Z(n29555) );
  XNOR U29952 ( .A(n29563), .B(n29777), .Z(n29556) );
  XNOR U29953 ( .A(n29562), .B(n29560), .Z(n29777) );
  AND U29954 ( .A(n29778), .B(n29779), .Z(n29560) );
  NANDN U29955 ( .A(n29780), .B(n29781), .Z(n29779) );
  NANDN U29956 ( .A(n29782), .B(n29783), .Z(n29781) );
  NANDN U29957 ( .A(n29783), .B(n29782), .Z(n29778) );
  ANDN U29958 ( .B(B[176]), .A(n62), .Z(n29562) );
  XNOR U29959 ( .A(n29570), .B(n29784), .Z(n29563) );
  XNOR U29960 ( .A(n29569), .B(n29567), .Z(n29784) );
  AND U29961 ( .A(n29785), .B(n29786), .Z(n29567) );
  NANDN U29962 ( .A(n29787), .B(n29788), .Z(n29786) );
  OR U29963 ( .A(n29789), .B(n29790), .Z(n29788) );
  NAND U29964 ( .A(n29790), .B(n29789), .Z(n29785) );
  ANDN U29965 ( .B(B[177]), .A(n63), .Z(n29569) );
  XNOR U29966 ( .A(n29577), .B(n29791), .Z(n29570) );
  XNOR U29967 ( .A(n29576), .B(n29574), .Z(n29791) );
  AND U29968 ( .A(n29792), .B(n29793), .Z(n29574) );
  NANDN U29969 ( .A(n29794), .B(n29795), .Z(n29793) );
  NANDN U29970 ( .A(n29796), .B(n29797), .Z(n29795) );
  NANDN U29971 ( .A(n29797), .B(n29796), .Z(n29792) );
  ANDN U29972 ( .B(B[178]), .A(n64), .Z(n29576) );
  XNOR U29973 ( .A(n29584), .B(n29798), .Z(n29577) );
  XNOR U29974 ( .A(n29583), .B(n29581), .Z(n29798) );
  AND U29975 ( .A(n29799), .B(n29800), .Z(n29581) );
  NANDN U29976 ( .A(n29801), .B(n29802), .Z(n29800) );
  OR U29977 ( .A(n29803), .B(n29804), .Z(n29802) );
  NAND U29978 ( .A(n29804), .B(n29803), .Z(n29799) );
  ANDN U29979 ( .B(B[179]), .A(n65), .Z(n29583) );
  XNOR U29980 ( .A(n29591), .B(n29805), .Z(n29584) );
  XNOR U29981 ( .A(n29590), .B(n29588), .Z(n29805) );
  AND U29982 ( .A(n29806), .B(n29807), .Z(n29588) );
  NANDN U29983 ( .A(n29808), .B(n29809), .Z(n29807) );
  NANDN U29984 ( .A(n29810), .B(n29811), .Z(n29809) );
  NANDN U29985 ( .A(n29811), .B(n29810), .Z(n29806) );
  ANDN U29986 ( .B(B[180]), .A(n66), .Z(n29590) );
  XNOR U29987 ( .A(n29598), .B(n29812), .Z(n29591) );
  XNOR U29988 ( .A(n29597), .B(n29595), .Z(n29812) );
  AND U29989 ( .A(n29813), .B(n29814), .Z(n29595) );
  NANDN U29990 ( .A(n29815), .B(n29816), .Z(n29814) );
  OR U29991 ( .A(n29817), .B(n29818), .Z(n29816) );
  NAND U29992 ( .A(n29818), .B(n29817), .Z(n29813) );
  ANDN U29993 ( .B(B[181]), .A(n67), .Z(n29597) );
  XNOR U29994 ( .A(n29605), .B(n29819), .Z(n29598) );
  XNOR U29995 ( .A(n29604), .B(n29602), .Z(n29819) );
  AND U29996 ( .A(n29820), .B(n29821), .Z(n29602) );
  NANDN U29997 ( .A(n29822), .B(n29823), .Z(n29821) );
  NANDN U29998 ( .A(n29824), .B(n29825), .Z(n29823) );
  NANDN U29999 ( .A(n29825), .B(n29824), .Z(n29820) );
  ANDN U30000 ( .B(B[182]), .A(n68), .Z(n29604) );
  XNOR U30001 ( .A(n29612), .B(n29826), .Z(n29605) );
  XNOR U30002 ( .A(n29611), .B(n29609), .Z(n29826) );
  AND U30003 ( .A(n29827), .B(n29828), .Z(n29609) );
  NANDN U30004 ( .A(n29829), .B(n29830), .Z(n29828) );
  OR U30005 ( .A(n29831), .B(n29832), .Z(n29830) );
  NAND U30006 ( .A(n29832), .B(n29831), .Z(n29827) );
  ANDN U30007 ( .B(B[183]), .A(n69), .Z(n29611) );
  XNOR U30008 ( .A(n29619), .B(n29833), .Z(n29612) );
  XNOR U30009 ( .A(n29618), .B(n29616), .Z(n29833) );
  AND U30010 ( .A(n29834), .B(n29835), .Z(n29616) );
  NANDN U30011 ( .A(n29836), .B(n29837), .Z(n29835) );
  NANDN U30012 ( .A(n29838), .B(n29839), .Z(n29837) );
  NANDN U30013 ( .A(n29839), .B(n29838), .Z(n29834) );
  ANDN U30014 ( .B(B[184]), .A(n70), .Z(n29618) );
  XNOR U30015 ( .A(n29626), .B(n29840), .Z(n29619) );
  XNOR U30016 ( .A(n29625), .B(n29623), .Z(n29840) );
  AND U30017 ( .A(n29841), .B(n29842), .Z(n29623) );
  NANDN U30018 ( .A(n29843), .B(n29844), .Z(n29842) );
  OR U30019 ( .A(n29845), .B(n29846), .Z(n29844) );
  NAND U30020 ( .A(n29846), .B(n29845), .Z(n29841) );
  ANDN U30021 ( .B(B[185]), .A(n71), .Z(n29625) );
  XNOR U30022 ( .A(n29633), .B(n29847), .Z(n29626) );
  XNOR U30023 ( .A(n29632), .B(n29630), .Z(n29847) );
  AND U30024 ( .A(n29848), .B(n29849), .Z(n29630) );
  NANDN U30025 ( .A(n29850), .B(n29851), .Z(n29849) );
  NANDN U30026 ( .A(n29852), .B(n29853), .Z(n29851) );
  NANDN U30027 ( .A(n29853), .B(n29852), .Z(n29848) );
  ANDN U30028 ( .B(B[186]), .A(n72), .Z(n29632) );
  XNOR U30029 ( .A(n29640), .B(n29854), .Z(n29633) );
  XNOR U30030 ( .A(n29639), .B(n29637), .Z(n29854) );
  AND U30031 ( .A(n29855), .B(n29856), .Z(n29637) );
  NANDN U30032 ( .A(n29857), .B(n29858), .Z(n29856) );
  OR U30033 ( .A(n29859), .B(n29860), .Z(n29858) );
  NAND U30034 ( .A(n29860), .B(n29859), .Z(n29855) );
  ANDN U30035 ( .B(B[187]), .A(n73), .Z(n29639) );
  XNOR U30036 ( .A(n29647), .B(n29861), .Z(n29640) );
  XNOR U30037 ( .A(n29646), .B(n29644), .Z(n29861) );
  AND U30038 ( .A(n29862), .B(n29863), .Z(n29644) );
  NANDN U30039 ( .A(n29864), .B(n29865), .Z(n29863) );
  NANDN U30040 ( .A(n29866), .B(n29867), .Z(n29865) );
  NANDN U30041 ( .A(n29867), .B(n29866), .Z(n29862) );
  ANDN U30042 ( .B(B[188]), .A(n74), .Z(n29646) );
  XNOR U30043 ( .A(n29654), .B(n29868), .Z(n29647) );
  XNOR U30044 ( .A(n29653), .B(n29651), .Z(n29868) );
  AND U30045 ( .A(n29869), .B(n29870), .Z(n29651) );
  NANDN U30046 ( .A(n29871), .B(n29872), .Z(n29870) );
  OR U30047 ( .A(n29873), .B(n29874), .Z(n29872) );
  NAND U30048 ( .A(n29874), .B(n29873), .Z(n29869) );
  ANDN U30049 ( .B(B[189]), .A(n75), .Z(n29653) );
  XNOR U30050 ( .A(n29661), .B(n29875), .Z(n29654) );
  XNOR U30051 ( .A(n29660), .B(n29658), .Z(n29875) );
  AND U30052 ( .A(n29876), .B(n29877), .Z(n29658) );
  NANDN U30053 ( .A(n29878), .B(n29879), .Z(n29877) );
  NANDN U30054 ( .A(n29880), .B(n29881), .Z(n29879) );
  NANDN U30055 ( .A(n29881), .B(n29880), .Z(n29876) );
  ANDN U30056 ( .B(B[190]), .A(n76), .Z(n29660) );
  XNOR U30057 ( .A(n29668), .B(n29882), .Z(n29661) );
  XNOR U30058 ( .A(n29667), .B(n29665), .Z(n29882) );
  AND U30059 ( .A(n29883), .B(n29884), .Z(n29665) );
  NANDN U30060 ( .A(n29885), .B(n29886), .Z(n29884) );
  OR U30061 ( .A(n29887), .B(n29888), .Z(n29886) );
  NAND U30062 ( .A(n29888), .B(n29887), .Z(n29883) );
  ANDN U30063 ( .B(B[191]), .A(n77), .Z(n29667) );
  XNOR U30064 ( .A(n29675), .B(n29889), .Z(n29668) );
  XNOR U30065 ( .A(n29674), .B(n29672), .Z(n29889) );
  AND U30066 ( .A(n29890), .B(n29891), .Z(n29672) );
  NANDN U30067 ( .A(n29892), .B(n29893), .Z(n29891) );
  NANDN U30068 ( .A(n29894), .B(n29895), .Z(n29893) );
  NANDN U30069 ( .A(n29895), .B(n29894), .Z(n29890) );
  ANDN U30070 ( .B(B[192]), .A(n78), .Z(n29674) );
  XNOR U30071 ( .A(n29682), .B(n29896), .Z(n29675) );
  XNOR U30072 ( .A(n29681), .B(n29679), .Z(n29896) );
  AND U30073 ( .A(n29897), .B(n29898), .Z(n29679) );
  NANDN U30074 ( .A(n29899), .B(n29900), .Z(n29898) );
  OR U30075 ( .A(n29901), .B(n29902), .Z(n29900) );
  NAND U30076 ( .A(n29902), .B(n29901), .Z(n29897) );
  ANDN U30077 ( .B(B[193]), .A(n79), .Z(n29681) );
  XNOR U30078 ( .A(n29689), .B(n29903), .Z(n29682) );
  XNOR U30079 ( .A(n29688), .B(n29686), .Z(n29903) );
  AND U30080 ( .A(n29904), .B(n29905), .Z(n29686) );
  NANDN U30081 ( .A(n29906), .B(n29907), .Z(n29905) );
  NANDN U30082 ( .A(n29908), .B(n29909), .Z(n29907) );
  NANDN U30083 ( .A(n29909), .B(n29908), .Z(n29904) );
  ANDN U30084 ( .B(B[194]), .A(n80), .Z(n29688) );
  XNOR U30085 ( .A(n29696), .B(n29910), .Z(n29689) );
  XNOR U30086 ( .A(n29695), .B(n29693), .Z(n29910) );
  AND U30087 ( .A(n29911), .B(n29912), .Z(n29693) );
  NANDN U30088 ( .A(n29913), .B(n29914), .Z(n29912) );
  OR U30089 ( .A(n29915), .B(n29916), .Z(n29914) );
  NAND U30090 ( .A(n29916), .B(n29915), .Z(n29911) );
  ANDN U30091 ( .B(B[195]), .A(n81), .Z(n29695) );
  XNOR U30092 ( .A(n29703), .B(n29917), .Z(n29696) );
  XNOR U30093 ( .A(n29702), .B(n29700), .Z(n29917) );
  AND U30094 ( .A(n29918), .B(n29919), .Z(n29700) );
  NANDN U30095 ( .A(n29920), .B(n29921), .Z(n29919) );
  NAND U30096 ( .A(n29922), .B(n29923), .Z(n29921) );
  ANDN U30097 ( .B(B[196]), .A(n82), .Z(n29702) );
  XOR U30098 ( .A(n29709), .B(n29924), .Z(n29703) );
  XNOR U30099 ( .A(n29707), .B(n29710), .Z(n29924) );
  NAND U30100 ( .A(A[2]), .B(B[197]), .Z(n29710) );
  NANDN U30101 ( .A(n29925), .B(n29926), .Z(n29707) );
  AND U30102 ( .A(A[0]), .B(B[198]), .Z(n29926) );
  XNOR U30103 ( .A(n29712), .B(n29927), .Z(n29709) );
  NAND U30104 ( .A(A[0]), .B(B[199]), .Z(n29927) );
  NAND U30105 ( .A(B[198]), .B(A[1]), .Z(n29712) );
  NAND U30106 ( .A(n29928), .B(n29929), .Z(n398) );
  NANDN U30107 ( .A(n29930), .B(n29931), .Z(n29929) );
  OR U30108 ( .A(n29932), .B(n29933), .Z(n29931) );
  NAND U30109 ( .A(n29933), .B(n29932), .Z(n29928) );
  XOR U30110 ( .A(n400), .B(n399), .Z(\A1[196] ) );
  XOR U30111 ( .A(n29933), .B(n29934), .Z(n399) );
  XNOR U30112 ( .A(n29932), .B(n29930), .Z(n29934) );
  AND U30113 ( .A(n29935), .B(n29936), .Z(n29930) );
  NANDN U30114 ( .A(n29937), .B(n29938), .Z(n29936) );
  NANDN U30115 ( .A(n29939), .B(n29940), .Z(n29938) );
  NANDN U30116 ( .A(n29940), .B(n29939), .Z(n29935) );
  ANDN U30117 ( .B(B[167]), .A(n54), .Z(n29932) );
  XNOR U30118 ( .A(n29727), .B(n29941), .Z(n29933) );
  XNOR U30119 ( .A(n29726), .B(n29724), .Z(n29941) );
  AND U30120 ( .A(n29942), .B(n29943), .Z(n29724) );
  NANDN U30121 ( .A(n29944), .B(n29945), .Z(n29943) );
  OR U30122 ( .A(n29946), .B(n29947), .Z(n29945) );
  NAND U30123 ( .A(n29947), .B(n29946), .Z(n29942) );
  ANDN U30124 ( .B(B[168]), .A(n55), .Z(n29726) );
  XNOR U30125 ( .A(n29734), .B(n29948), .Z(n29727) );
  XNOR U30126 ( .A(n29733), .B(n29731), .Z(n29948) );
  AND U30127 ( .A(n29949), .B(n29950), .Z(n29731) );
  NANDN U30128 ( .A(n29951), .B(n29952), .Z(n29950) );
  NANDN U30129 ( .A(n29953), .B(n29954), .Z(n29952) );
  NANDN U30130 ( .A(n29954), .B(n29953), .Z(n29949) );
  ANDN U30131 ( .B(B[169]), .A(n56), .Z(n29733) );
  XNOR U30132 ( .A(n29741), .B(n29955), .Z(n29734) );
  XNOR U30133 ( .A(n29740), .B(n29738), .Z(n29955) );
  AND U30134 ( .A(n29956), .B(n29957), .Z(n29738) );
  NANDN U30135 ( .A(n29958), .B(n29959), .Z(n29957) );
  OR U30136 ( .A(n29960), .B(n29961), .Z(n29959) );
  NAND U30137 ( .A(n29961), .B(n29960), .Z(n29956) );
  ANDN U30138 ( .B(B[170]), .A(n57), .Z(n29740) );
  XNOR U30139 ( .A(n29748), .B(n29962), .Z(n29741) );
  XNOR U30140 ( .A(n29747), .B(n29745), .Z(n29962) );
  AND U30141 ( .A(n29963), .B(n29964), .Z(n29745) );
  NANDN U30142 ( .A(n29965), .B(n29966), .Z(n29964) );
  NANDN U30143 ( .A(n29967), .B(n29968), .Z(n29966) );
  NANDN U30144 ( .A(n29968), .B(n29967), .Z(n29963) );
  ANDN U30145 ( .B(B[171]), .A(n58), .Z(n29747) );
  XNOR U30146 ( .A(n29755), .B(n29969), .Z(n29748) );
  XNOR U30147 ( .A(n29754), .B(n29752), .Z(n29969) );
  AND U30148 ( .A(n29970), .B(n29971), .Z(n29752) );
  NANDN U30149 ( .A(n29972), .B(n29973), .Z(n29971) );
  OR U30150 ( .A(n29974), .B(n29975), .Z(n29973) );
  NAND U30151 ( .A(n29975), .B(n29974), .Z(n29970) );
  ANDN U30152 ( .B(B[172]), .A(n59), .Z(n29754) );
  XNOR U30153 ( .A(n29762), .B(n29976), .Z(n29755) );
  XNOR U30154 ( .A(n29761), .B(n29759), .Z(n29976) );
  AND U30155 ( .A(n29977), .B(n29978), .Z(n29759) );
  NANDN U30156 ( .A(n29979), .B(n29980), .Z(n29978) );
  NANDN U30157 ( .A(n29981), .B(n29982), .Z(n29980) );
  NANDN U30158 ( .A(n29982), .B(n29981), .Z(n29977) );
  ANDN U30159 ( .B(B[173]), .A(n60), .Z(n29761) );
  XNOR U30160 ( .A(n29769), .B(n29983), .Z(n29762) );
  XNOR U30161 ( .A(n29768), .B(n29766), .Z(n29983) );
  AND U30162 ( .A(n29984), .B(n29985), .Z(n29766) );
  NANDN U30163 ( .A(n29986), .B(n29987), .Z(n29985) );
  OR U30164 ( .A(n29988), .B(n29989), .Z(n29987) );
  NAND U30165 ( .A(n29989), .B(n29988), .Z(n29984) );
  ANDN U30166 ( .B(B[174]), .A(n61), .Z(n29768) );
  XNOR U30167 ( .A(n29776), .B(n29990), .Z(n29769) );
  XNOR U30168 ( .A(n29775), .B(n29773), .Z(n29990) );
  AND U30169 ( .A(n29991), .B(n29992), .Z(n29773) );
  NANDN U30170 ( .A(n29993), .B(n29994), .Z(n29992) );
  NANDN U30171 ( .A(n29995), .B(n29996), .Z(n29994) );
  NANDN U30172 ( .A(n29996), .B(n29995), .Z(n29991) );
  ANDN U30173 ( .B(B[175]), .A(n62), .Z(n29775) );
  XNOR U30174 ( .A(n29783), .B(n29997), .Z(n29776) );
  XNOR U30175 ( .A(n29782), .B(n29780), .Z(n29997) );
  AND U30176 ( .A(n29998), .B(n29999), .Z(n29780) );
  NANDN U30177 ( .A(n30000), .B(n30001), .Z(n29999) );
  OR U30178 ( .A(n30002), .B(n30003), .Z(n30001) );
  NAND U30179 ( .A(n30003), .B(n30002), .Z(n29998) );
  ANDN U30180 ( .B(B[176]), .A(n63), .Z(n29782) );
  XNOR U30181 ( .A(n29790), .B(n30004), .Z(n29783) );
  XNOR U30182 ( .A(n29789), .B(n29787), .Z(n30004) );
  AND U30183 ( .A(n30005), .B(n30006), .Z(n29787) );
  NANDN U30184 ( .A(n30007), .B(n30008), .Z(n30006) );
  NANDN U30185 ( .A(n30009), .B(n30010), .Z(n30008) );
  NANDN U30186 ( .A(n30010), .B(n30009), .Z(n30005) );
  ANDN U30187 ( .B(B[177]), .A(n64), .Z(n29789) );
  XNOR U30188 ( .A(n29797), .B(n30011), .Z(n29790) );
  XNOR U30189 ( .A(n29796), .B(n29794), .Z(n30011) );
  AND U30190 ( .A(n30012), .B(n30013), .Z(n29794) );
  NANDN U30191 ( .A(n30014), .B(n30015), .Z(n30013) );
  OR U30192 ( .A(n30016), .B(n30017), .Z(n30015) );
  NAND U30193 ( .A(n30017), .B(n30016), .Z(n30012) );
  ANDN U30194 ( .B(B[178]), .A(n65), .Z(n29796) );
  XNOR U30195 ( .A(n29804), .B(n30018), .Z(n29797) );
  XNOR U30196 ( .A(n29803), .B(n29801), .Z(n30018) );
  AND U30197 ( .A(n30019), .B(n30020), .Z(n29801) );
  NANDN U30198 ( .A(n30021), .B(n30022), .Z(n30020) );
  NANDN U30199 ( .A(n30023), .B(n30024), .Z(n30022) );
  NANDN U30200 ( .A(n30024), .B(n30023), .Z(n30019) );
  ANDN U30201 ( .B(B[179]), .A(n66), .Z(n29803) );
  XNOR U30202 ( .A(n29811), .B(n30025), .Z(n29804) );
  XNOR U30203 ( .A(n29810), .B(n29808), .Z(n30025) );
  AND U30204 ( .A(n30026), .B(n30027), .Z(n29808) );
  NANDN U30205 ( .A(n30028), .B(n30029), .Z(n30027) );
  OR U30206 ( .A(n30030), .B(n30031), .Z(n30029) );
  NAND U30207 ( .A(n30031), .B(n30030), .Z(n30026) );
  ANDN U30208 ( .B(B[180]), .A(n67), .Z(n29810) );
  XNOR U30209 ( .A(n29818), .B(n30032), .Z(n29811) );
  XNOR U30210 ( .A(n29817), .B(n29815), .Z(n30032) );
  AND U30211 ( .A(n30033), .B(n30034), .Z(n29815) );
  NANDN U30212 ( .A(n30035), .B(n30036), .Z(n30034) );
  NANDN U30213 ( .A(n30037), .B(n30038), .Z(n30036) );
  NANDN U30214 ( .A(n30038), .B(n30037), .Z(n30033) );
  ANDN U30215 ( .B(B[181]), .A(n68), .Z(n29817) );
  XNOR U30216 ( .A(n29825), .B(n30039), .Z(n29818) );
  XNOR U30217 ( .A(n29824), .B(n29822), .Z(n30039) );
  AND U30218 ( .A(n30040), .B(n30041), .Z(n29822) );
  NANDN U30219 ( .A(n30042), .B(n30043), .Z(n30041) );
  OR U30220 ( .A(n30044), .B(n30045), .Z(n30043) );
  NAND U30221 ( .A(n30045), .B(n30044), .Z(n30040) );
  ANDN U30222 ( .B(B[182]), .A(n69), .Z(n29824) );
  XNOR U30223 ( .A(n29832), .B(n30046), .Z(n29825) );
  XNOR U30224 ( .A(n29831), .B(n29829), .Z(n30046) );
  AND U30225 ( .A(n30047), .B(n30048), .Z(n29829) );
  NANDN U30226 ( .A(n30049), .B(n30050), .Z(n30048) );
  NANDN U30227 ( .A(n30051), .B(n30052), .Z(n30050) );
  NANDN U30228 ( .A(n30052), .B(n30051), .Z(n30047) );
  ANDN U30229 ( .B(B[183]), .A(n70), .Z(n29831) );
  XNOR U30230 ( .A(n29839), .B(n30053), .Z(n29832) );
  XNOR U30231 ( .A(n29838), .B(n29836), .Z(n30053) );
  AND U30232 ( .A(n30054), .B(n30055), .Z(n29836) );
  NANDN U30233 ( .A(n30056), .B(n30057), .Z(n30055) );
  OR U30234 ( .A(n30058), .B(n30059), .Z(n30057) );
  NAND U30235 ( .A(n30059), .B(n30058), .Z(n30054) );
  ANDN U30236 ( .B(B[184]), .A(n71), .Z(n29838) );
  XNOR U30237 ( .A(n29846), .B(n30060), .Z(n29839) );
  XNOR U30238 ( .A(n29845), .B(n29843), .Z(n30060) );
  AND U30239 ( .A(n30061), .B(n30062), .Z(n29843) );
  NANDN U30240 ( .A(n30063), .B(n30064), .Z(n30062) );
  NANDN U30241 ( .A(n30065), .B(n30066), .Z(n30064) );
  NANDN U30242 ( .A(n30066), .B(n30065), .Z(n30061) );
  ANDN U30243 ( .B(B[185]), .A(n72), .Z(n29845) );
  XNOR U30244 ( .A(n29853), .B(n30067), .Z(n29846) );
  XNOR U30245 ( .A(n29852), .B(n29850), .Z(n30067) );
  AND U30246 ( .A(n30068), .B(n30069), .Z(n29850) );
  NANDN U30247 ( .A(n30070), .B(n30071), .Z(n30069) );
  OR U30248 ( .A(n30072), .B(n30073), .Z(n30071) );
  NAND U30249 ( .A(n30073), .B(n30072), .Z(n30068) );
  ANDN U30250 ( .B(B[186]), .A(n73), .Z(n29852) );
  XNOR U30251 ( .A(n29860), .B(n30074), .Z(n29853) );
  XNOR U30252 ( .A(n29859), .B(n29857), .Z(n30074) );
  AND U30253 ( .A(n30075), .B(n30076), .Z(n29857) );
  NANDN U30254 ( .A(n30077), .B(n30078), .Z(n30076) );
  NANDN U30255 ( .A(n30079), .B(n30080), .Z(n30078) );
  NANDN U30256 ( .A(n30080), .B(n30079), .Z(n30075) );
  ANDN U30257 ( .B(B[187]), .A(n74), .Z(n29859) );
  XNOR U30258 ( .A(n29867), .B(n30081), .Z(n29860) );
  XNOR U30259 ( .A(n29866), .B(n29864), .Z(n30081) );
  AND U30260 ( .A(n30082), .B(n30083), .Z(n29864) );
  NANDN U30261 ( .A(n30084), .B(n30085), .Z(n30083) );
  OR U30262 ( .A(n30086), .B(n30087), .Z(n30085) );
  NAND U30263 ( .A(n30087), .B(n30086), .Z(n30082) );
  ANDN U30264 ( .B(B[188]), .A(n75), .Z(n29866) );
  XNOR U30265 ( .A(n29874), .B(n30088), .Z(n29867) );
  XNOR U30266 ( .A(n29873), .B(n29871), .Z(n30088) );
  AND U30267 ( .A(n30089), .B(n30090), .Z(n29871) );
  NANDN U30268 ( .A(n30091), .B(n30092), .Z(n30090) );
  NANDN U30269 ( .A(n30093), .B(n30094), .Z(n30092) );
  NANDN U30270 ( .A(n30094), .B(n30093), .Z(n30089) );
  ANDN U30271 ( .B(B[189]), .A(n76), .Z(n29873) );
  XNOR U30272 ( .A(n29881), .B(n30095), .Z(n29874) );
  XNOR U30273 ( .A(n29880), .B(n29878), .Z(n30095) );
  AND U30274 ( .A(n30096), .B(n30097), .Z(n29878) );
  NANDN U30275 ( .A(n30098), .B(n30099), .Z(n30097) );
  OR U30276 ( .A(n30100), .B(n30101), .Z(n30099) );
  NAND U30277 ( .A(n30101), .B(n30100), .Z(n30096) );
  ANDN U30278 ( .B(B[190]), .A(n77), .Z(n29880) );
  XNOR U30279 ( .A(n29888), .B(n30102), .Z(n29881) );
  XNOR U30280 ( .A(n29887), .B(n29885), .Z(n30102) );
  AND U30281 ( .A(n30103), .B(n30104), .Z(n29885) );
  NANDN U30282 ( .A(n30105), .B(n30106), .Z(n30104) );
  NANDN U30283 ( .A(n30107), .B(n30108), .Z(n30106) );
  NANDN U30284 ( .A(n30108), .B(n30107), .Z(n30103) );
  ANDN U30285 ( .B(B[191]), .A(n78), .Z(n29887) );
  XNOR U30286 ( .A(n29895), .B(n30109), .Z(n29888) );
  XNOR U30287 ( .A(n29894), .B(n29892), .Z(n30109) );
  AND U30288 ( .A(n30110), .B(n30111), .Z(n29892) );
  NANDN U30289 ( .A(n30112), .B(n30113), .Z(n30111) );
  OR U30290 ( .A(n30114), .B(n30115), .Z(n30113) );
  NAND U30291 ( .A(n30115), .B(n30114), .Z(n30110) );
  ANDN U30292 ( .B(B[192]), .A(n79), .Z(n29894) );
  XNOR U30293 ( .A(n29902), .B(n30116), .Z(n29895) );
  XNOR U30294 ( .A(n29901), .B(n29899), .Z(n30116) );
  AND U30295 ( .A(n30117), .B(n30118), .Z(n29899) );
  NANDN U30296 ( .A(n30119), .B(n30120), .Z(n30118) );
  NANDN U30297 ( .A(n30121), .B(n30122), .Z(n30120) );
  NANDN U30298 ( .A(n30122), .B(n30121), .Z(n30117) );
  ANDN U30299 ( .B(B[193]), .A(n80), .Z(n29901) );
  XNOR U30300 ( .A(n29909), .B(n30123), .Z(n29902) );
  XNOR U30301 ( .A(n29908), .B(n29906), .Z(n30123) );
  AND U30302 ( .A(n30124), .B(n30125), .Z(n29906) );
  NANDN U30303 ( .A(n30126), .B(n30127), .Z(n30125) );
  OR U30304 ( .A(n30128), .B(n30129), .Z(n30127) );
  NAND U30305 ( .A(n30129), .B(n30128), .Z(n30124) );
  ANDN U30306 ( .B(B[194]), .A(n81), .Z(n29908) );
  XNOR U30307 ( .A(n29916), .B(n30130), .Z(n29909) );
  XNOR U30308 ( .A(n29915), .B(n29913), .Z(n30130) );
  AND U30309 ( .A(n30131), .B(n30132), .Z(n29913) );
  NANDN U30310 ( .A(n30133), .B(n30134), .Z(n30132) );
  NAND U30311 ( .A(n30135), .B(n30136), .Z(n30134) );
  ANDN U30312 ( .B(B[195]), .A(n82), .Z(n29915) );
  XOR U30313 ( .A(n29922), .B(n30137), .Z(n29916) );
  XNOR U30314 ( .A(n29920), .B(n29923), .Z(n30137) );
  NAND U30315 ( .A(A[2]), .B(B[196]), .Z(n29923) );
  NANDN U30316 ( .A(n30138), .B(n30139), .Z(n29920) );
  AND U30317 ( .A(A[0]), .B(B[197]), .Z(n30139) );
  XNOR U30318 ( .A(n29925), .B(n30140), .Z(n29922) );
  NAND U30319 ( .A(A[0]), .B(B[198]), .Z(n30140) );
  NAND U30320 ( .A(B[197]), .B(A[1]), .Z(n29925) );
  NAND U30321 ( .A(n30141), .B(n30142), .Z(n400) );
  NANDN U30322 ( .A(n30143), .B(n30144), .Z(n30142) );
  OR U30323 ( .A(n30145), .B(n30146), .Z(n30144) );
  NAND U30324 ( .A(n30146), .B(n30145), .Z(n30141) );
  XOR U30325 ( .A(n402), .B(n401), .Z(\A1[195] ) );
  XOR U30326 ( .A(n30146), .B(n30147), .Z(n401) );
  XNOR U30327 ( .A(n30145), .B(n30143), .Z(n30147) );
  AND U30328 ( .A(n30148), .B(n30149), .Z(n30143) );
  NANDN U30329 ( .A(n30150), .B(n30151), .Z(n30149) );
  NANDN U30330 ( .A(n30152), .B(n30153), .Z(n30151) );
  NANDN U30331 ( .A(n30153), .B(n30152), .Z(n30148) );
  ANDN U30332 ( .B(B[166]), .A(n54), .Z(n30145) );
  XNOR U30333 ( .A(n29940), .B(n30154), .Z(n30146) );
  XNOR U30334 ( .A(n29939), .B(n29937), .Z(n30154) );
  AND U30335 ( .A(n30155), .B(n30156), .Z(n29937) );
  NANDN U30336 ( .A(n30157), .B(n30158), .Z(n30156) );
  OR U30337 ( .A(n30159), .B(n30160), .Z(n30158) );
  NAND U30338 ( .A(n30160), .B(n30159), .Z(n30155) );
  ANDN U30339 ( .B(B[167]), .A(n55), .Z(n29939) );
  XNOR U30340 ( .A(n29947), .B(n30161), .Z(n29940) );
  XNOR U30341 ( .A(n29946), .B(n29944), .Z(n30161) );
  AND U30342 ( .A(n30162), .B(n30163), .Z(n29944) );
  NANDN U30343 ( .A(n30164), .B(n30165), .Z(n30163) );
  NANDN U30344 ( .A(n30166), .B(n30167), .Z(n30165) );
  NANDN U30345 ( .A(n30167), .B(n30166), .Z(n30162) );
  ANDN U30346 ( .B(B[168]), .A(n56), .Z(n29946) );
  XNOR U30347 ( .A(n29954), .B(n30168), .Z(n29947) );
  XNOR U30348 ( .A(n29953), .B(n29951), .Z(n30168) );
  AND U30349 ( .A(n30169), .B(n30170), .Z(n29951) );
  NANDN U30350 ( .A(n30171), .B(n30172), .Z(n30170) );
  OR U30351 ( .A(n30173), .B(n30174), .Z(n30172) );
  NAND U30352 ( .A(n30174), .B(n30173), .Z(n30169) );
  ANDN U30353 ( .B(B[169]), .A(n57), .Z(n29953) );
  XNOR U30354 ( .A(n29961), .B(n30175), .Z(n29954) );
  XNOR U30355 ( .A(n29960), .B(n29958), .Z(n30175) );
  AND U30356 ( .A(n30176), .B(n30177), .Z(n29958) );
  NANDN U30357 ( .A(n30178), .B(n30179), .Z(n30177) );
  NANDN U30358 ( .A(n30180), .B(n30181), .Z(n30179) );
  NANDN U30359 ( .A(n30181), .B(n30180), .Z(n30176) );
  ANDN U30360 ( .B(B[170]), .A(n58), .Z(n29960) );
  XNOR U30361 ( .A(n29968), .B(n30182), .Z(n29961) );
  XNOR U30362 ( .A(n29967), .B(n29965), .Z(n30182) );
  AND U30363 ( .A(n30183), .B(n30184), .Z(n29965) );
  NANDN U30364 ( .A(n30185), .B(n30186), .Z(n30184) );
  OR U30365 ( .A(n30187), .B(n30188), .Z(n30186) );
  NAND U30366 ( .A(n30188), .B(n30187), .Z(n30183) );
  ANDN U30367 ( .B(B[171]), .A(n59), .Z(n29967) );
  XNOR U30368 ( .A(n29975), .B(n30189), .Z(n29968) );
  XNOR U30369 ( .A(n29974), .B(n29972), .Z(n30189) );
  AND U30370 ( .A(n30190), .B(n30191), .Z(n29972) );
  NANDN U30371 ( .A(n30192), .B(n30193), .Z(n30191) );
  NANDN U30372 ( .A(n30194), .B(n30195), .Z(n30193) );
  NANDN U30373 ( .A(n30195), .B(n30194), .Z(n30190) );
  ANDN U30374 ( .B(B[172]), .A(n60), .Z(n29974) );
  XNOR U30375 ( .A(n29982), .B(n30196), .Z(n29975) );
  XNOR U30376 ( .A(n29981), .B(n29979), .Z(n30196) );
  AND U30377 ( .A(n30197), .B(n30198), .Z(n29979) );
  NANDN U30378 ( .A(n30199), .B(n30200), .Z(n30198) );
  OR U30379 ( .A(n30201), .B(n30202), .Z(n30200) );
  NAND U30380 ( .A(n30202), .B(n30201), .Z(n30197) );
  ANDN U30381 ( .B(B[173]), .A(n61), .Z(n29981) );
  XNOR U30382 ( .A(n29989), .B(n30203), .Z(n29982) );
  XNOR U30383 ( .A(n29988), .B(n29986), .Z(n30203) );
  AND U30384 ( .A(n30204), .B(n30205), .Z(n29986) );
  NANDN U30385 ( .A(n30206), .B(n30207), .Z(n30205) );
  NANDN U30386 ( .A(n30208), .B(n30209), .Z(n30207) );
  NANDN U30387 ( .A(n30209), .B(n30208), .Z(n30204) );
  ANDN U30388 ( .B(B[174]), .A(n62), .Z(n29988) );
  XNOR U30389 ( .A(n29996), .B(n30210), .Z(n29989) );
  XNOR U30390 ( .A(n29995), .B(n29993), .Z(n30210) );
  AND U30391 ( .A(n30211), .B(n30212), .Z(n29993) );
  NANDN U30392 ( .A(n30213), .B(n30214), .Z(n30212) );
  OR U30393 ( .A(n30215), .B(n30216), .Z(n30214) );
  NAND U30394 ( .A(n30216), .B(n30215), .Z(n30211) );
  ANDN U30395 ( .B(B[175]), .A(n63), .Z(n29995) );
  XNOR U30396 ( .A(n30003), .B(n30217), .Z(n29996) );
  XNOR U30397 ( .A(n30002), .B(n30000), .Z(n30217) );
  AND U30398 ( .A(n30218), .B(n30219), .Z(n30000) );
  NANDN U30399 ( .A(n30220), .B(n30221), .Z(n30219) );
  NANDN U30400 ( .A(n30222), .B(n30223), .Z(n30221) );
  NANDN U30401 ( .A(n30223), .B(n30222), .Z(n30218) );
  ANDN U30402 ( .B(B[176]), .A(n64), .Z(n30002) );
  XNOR U30403 ( .A(n30010), .B(n30224), .Z(n30003) );
  XNOR U30404 ( .A(n30009), .B(n30007), .Z(n30224) );
  AND U30405 ( .A(n30225), .B(n30226), .Z(n30007) );
  NANDN U30406 ( .A(n30227), .B(n30228), .Z(n30226) );
  OR U30407 ( .A(n30229), .B(n30230), .Z(n30228) );
  NAND U30408 ( .A(n30230), .B(n30229), .Z(n30225) );
  ANDN U30409 ( .B(B[177]), .A(n65), .Z(n30009) );
  XNOR U30410 ( .A(n30017), .B(n30231), .Z(n30010) );
  XNOR U30411 ( .A(n30016), .B(n30014), .Z(n30231) );
  AND U30412 ( .A(n30232), .B(n30233), .Z(n30014) );
  NANDN U30413 ( .A(n30234), .B(n30235), .Z(n30233) );
  NANDN U30414 ( .A(n30236), .B(n30237), .Z(n30235) );
  NANDN U30415 ( .A(n30237), .B(n30236), .Z(n30232) );
  ANDN U30416 ( .B(B[178]), .A(n66), .Z(n30016) );
  XNOR U30417 ( .A(n30024), .B(n30238), .Z(n30017) );
  XNOR U30418 ( .A(n30023), .B(n30021), .Z(n30238) );
  AND U30419 ( .A(n30239), .B(n30240), .Z(n30021) );
  NANDN U30420 ( .A(n30241), .B(n30242), .Z(n30240) );
  OR U30421 ( .A(n30243), .B(n30244), .Z(n30242) );
  NAND U30422 ( .A(n30244), .B(n30243), .Z(n30239) );
  ANDN U30423 ( .B(B[179]), .A(n67), .Z(n30023) );
  XNOR U30424 ( .A(n30031), .B(n30245), .Z(n30024) );
  XNOR U30425 ( .A(n30030), .B(n30028), .Z(n30245) );
  AND U30426 ( .A(n30246), .B(n30247), .Z(n30028) );
  NANDN U30427 ( .A(n30248), .B(n30249), .Z(n30247) );
  NANDN U30428 ( .A(n30250), .B(n30251), .Z(n30249) );
  NANDN U30429 ( .A(n30251), .B(n30250), .Z(n30246) );
  ANDN U30430 ( .B(B[180]), .A(n68), .Z(n30030) );
  XNOR U30431 ( .A(n30038), .B(n30252), .Z(n30031) );
  XNOR U30432 ( .A(n30037), .B(n30035), .Z(n30252) );
  AND U30433 ( .A(n30253), .B(n30254), .Z(n30035) );
  NANDN U30434 ( .A(n30255), .B(n30256), .Z(n30254) );
  OR U30435 ( .A(n30257), .B(n30258), .Z(n30256) );
  NAND U30436 ( .A(n30258), .B(n30257), .Z(n30253) );
  ANDN U30437 ( .B(B[181]), .A(n69), .Z(n30037) );
  XNOR U30438 ( .A(n30045), .B(n30259), .Z(n30038) );
  XNOR U30439 ( .A(n30044), .B(n30042), .Z(n30259) );
  AND U30440 ( .A(n30260), .B(n30261), .Z(n30042) );
  NANDN U30441 ( .A(n30262), .B(n30263), .Z(n30261) );
  NANDN U30442 ( .A(n30264), .B(n30265), .Z(n30263) );
  NANDN U30443 ( .A(n30265), .B(n30264), .Z(n30260) );
  ANDN U30444 ( .B(B[182]), .A(n70), .Z(n30044) );
  XNOR U30445 ( .A(n30052), .B(n30266), .Z(n30045) );
  XNOR U30446 ( .A(n30051), .B(n30049), .Z(n30266) );
  AND U30447 ( .A(n30267), .B(n30268), .Z(n30049) );
  NANDN U30448 ( .A(n30269), .B(n30270), .Z(n30268) );
  OR U30449 ( .A(n30271), .B(n30272), .Z(n30270) );
  NAND U30450 ( .A(n30272), .B(n30271), .Z(n30267) );
  ANDN U30451 ( .B(B[183]), .A(n71), .Z(n30051) );
  XNOR U30452 ( .A(n30059), .B(n30273), .Z(n30052) );
  XNOR U30453 ( .A(n30058), .B(n30056), .Z(n30273) );
  AND U30454 ( .A(n30274), .B(n30275), .Z(n30056) );
  NANDN U30455 ( .A(n30276), .B(n30277), .Z(n30275) );
  NANDN U30456 ( .A(n30278), .B(n30279), .Z(n30277) );
  NANDN U30457 ( .A(n30279), .B(n30278), .Z(n30274) );
  ANDN U30458 ( .B(B[184]), .A(n72), .Z(n30058) );
  XNOR U30459 ( .A(n30066), .B(n30280), .Z(n30059) );
  XNOR U30460 ( .A(n30065), .B(n30063), .Z(n30280) );
  AND U30461 ( .A(n30281), .B(n30282), .Z(n30063) );
  NANDN U30462 ( .A(n30283), .B(n30284), .Z(n30282) );
  OR U30463 ( .A(n30285), .B(n30286), .Z(n30284) );
  NAND U30464 ( .A(n30286), .B(n30285), .Z(n30281) );
  ANDN U30465 ( .B(B[185]), .A(n73), .Z(n30065) );
  XNOR U30466 ( .A(n30073), .B(n30287), .Z(n30066) );
  XNOR U30467 ( .A(n30072), .B(n30070), .Z(n30287) );
  AND U30468 ( .A(n30288), .B(n30289), .Z(n30070) );
  NANDN U30469 ( .A(n30290), .B(n30291), .Z(n30289) );
  NANDN U30470 ( .A(n30292), .B(n30293), .Z(n30291) );
  NANDN U30471 ( .A(n30293), .B(n30292), .Z(n30288) );
  ANDN U30472 ( .B(B[186]), .A(n74), .Z(n30072) );
  XNOR U30473 ( .A(n30080), .B(n30294), .Z(n30073) );
  XNOR U30474 ( .A(n30079), .B(n30077), .Z(n30294) );
  AND U30475 ( .A(n30295), .B(n30296), .Z(n30077) );
  NANDN U30476 ( .A(n30297), .B(n30298), .Z(n30296) );
  OR U30477 ( .A(n30299), .B(n30300), .Z(n30298) );
  NAND U30478 ( .A(n30300), .B(n30299), .Z(n30295) );
  ANDN U30479 ( .B(B[187]), .A(n75), .Z(n30079) );
  XNOR U30480 ( .A(n30087), .B(n30301), .Z(n30080) );
  XNOR U30481 ( .A(n30086), .B(n30084), .Z(n30301) );
  AND U30482 ( .A(n30302), .B(n30303), .Z(n30084) );
  NANDN U30483 ( .A(n30304), .B(n30305), .Z(n30303) );
  NANDN U30484 ( .A(n30306), .B(n30307), .Z(n30305) );
  NANDN U30485 ( .A(n30307), .B(n30306), .Z(n30302) );
  ANDN U30486 ( .B(B[188]), .A(n76), .Z(n30086) );
  XNOR U30487 ( .A(n30094), .B(n30308), .Z(n30087) );
  XNOR U30488 ( .A(n30093), .B(n30091), .Z(n30308) );
  AND U30489 ( .A(n30309), .B(n30310), .Z(n30091) );
  NANDN U30490 ( .A(n30311), .B(n30312), .Z(n30310) );
  OR U30491 ( .A(n30313), .B(n30314), .Z(n30312) );
  NAND U30492 ( .A(n30314), .B(n30313), .Z(n30309) );
  ANDN U30493 ( .B(B[189]), .A(n77), .Z(n30093) );
  XNOR U30494 ( .A(n30101), .B(n30315), .Z(n30094) );
  XNOR U30495 ( .A(n30100), .B(n30098), .Z(n30315) );
  AND U30496 ( .A(n30316), .B(n30317), .Z(n30098) );
  NANDN U30497 ( .A(n30318), .B(n30319), .Z(n30317) );
  NANDN U30498 ( .A(n30320), .B(n30321), .Z(n30319) );
  NANDN U30499 ( .A(n30321), .B(n30320), .Z(n30316) );
  ANDN U30500 ( .B(B[190]), .A(n78), .Z(n30100) );
  XNOR U30501 ( .A(n30108), .B(n30322), .Z(n30101) );
  XNOR U30502 ( .A(n30107), .B(n30105), .Z(n30322) );
  AND U30503 ( .A(n30323), .B(n30324), .Z(n30105) );
  NANDN U30504 ( .A(n30325), .B(n30326), .Z(n30324) );
  OR U30505 ( .A(n30327), .B(n30328), .Z(n30326) );
  NAND U30506 ( .A(n30328), .B(n30327), .Z(n30323) );
  ANDN U30507 ( .B(B[191]), .A(n79), .Z(n30107) );
  XNOR U30508 ( .A(n30115), .B(n30329), .Z(n30108) );
  XNOR U30509 ( .A(n30114), .B(n30112), .Z(n30329) );
  AND U30510 ( .A(n30330), .B(n30331), .Z(n30112) );
  NANDN U30511 ( .A(n30332), .B(n30333), .Z(n30331) );
  NANDN U30512 ( .A(n30334), .B(n30335), .Z(n30333) );
  NANDN U30513 ( .A(n30335), .B(n30334), .Z(n30330) );
  ANDN U30514 ( .B(B[192]), .A(n80), .Z(n30114) );
  XNOR U30515 ( .A(n30122), .B(n30336), .Z(n30115) );
  XNOR U30516 ( .A(n30121), .B(n30119), .Z(n30336) );
  AND U30517 ( .A(n30337), .B(n30338), .Z(n30119) );
  NANDN U30518 ( .A(n30339), .B(n30340), .Z(n30338) );
  OR U30519 ( .A(n30341), .B(n30342), .Z(n30340) );
  NAND U30520 ( .A(n30342), .B(n30341), .Z(n30337) );
  ANDN U30521 ( .B(B[193]), .A(n81), .Z(n30121) );
  XNOR U30522 ( .A(n30129), .B(n30343), .Z(n30122) );
  XNOR U30523 ( .A(n30128), .B(n30126), .Z(n30343) );
  AND U30524 ( .A(n30344), .B(n30345), .Z(n30126) );
  NANDN U30525 ( .A(n30346), .B(n30347), .Z(n30345) );
  NAND U30526 ( .A(n30348), .B(n30349), .Z(n30347) );
  ANDN U30527 ( .B(B[194]), .A(n82), .Z(n30128) );
  XOR U30528 ( .A(n30135), .B(n30350), .Z(n30129) );
  XNOR U30529 ( .A(n30133), .B(n30136), .Z(n30350) );
  NAND U30530 ( .A(A[2]), .B(B[195]), .Z(n30136) );
  NANDN U30531 ( .A(n30351), .B(n30352), .Z(n30133) );
  AND U30532 ( .A(A[0]), .B(B[196]), .Z(n30352) );
  XNOR U30533 ( .A(n30138), .B(n30353), .Z(n30135) );
  NAND U30534 ( .A(A[0]), .B(B[197]), .Z(n30353) );
  NAND U30535 ( .A(B[196]), .B(A[1]), .Z(n30138) );
  NAND U30536 ( .A(n30354), .B(n30355), .Z(n402) );
  NANDN U30537 ( .A(n30356), .B(n30357), .Z(n30355) );
  OR U30538 ( .A(n30358), .B(n30359), .Z(n30357) );
  NAND U30539 ( .A(n30359), .B(n30358), .Z(n30354) );
  XOR U30540 ( .A(n404), .B(n403), .Z(\A1[194] ) );
  XOR U30541 ( .A(n30359), .B(n30360), .Z(n403) );
  XNOR U30542 ( .A(n30358), .B(n30356), .Z(n30360) );
  AND U30543 ( .A(n30361), .B(n30362), .Z(n30356) );
  NANDN U30544 ( .A(n30363), .B(n30364), .Z(n30362) );
  NANDN U30545 ( .A(n30365), .B(n30366), .Z(n30364) );
  NANDN U30546 ( .A(n30366), .B(n30365), .Z(n30361) );
  ANDN U30547 ( .B(B[165]), .A(n54), .Z(n30358) );
  XNOR U30548 ( .A(n30153), .B(n30367), .Z(n30359) );
  XNOR U30549 ( .A(n30152), .B(n30150), .Z(n30367) );
  AND U30550 ( .A(n30368), .B(n30369), .Z(n30150) );
  NANDN U30551 ( .A(n30370), .B(n30371), .Z(n30369) );
  OR U30552 ( .A(n30372), .B(n30373), .Z(n30371) );
  NAND U30553 ( .A(n30373), .B(n30372), .Z(n30368) );
  ANDN U30554 ( .B(B[166]), .A(n55), .Z(n30152) );
  XNOR U30555 ( .A(n30160), .B(n30374), .Z(n30153) );
  XNOR U30556 ( .A(n30159), .B(n30157), .Z(n30374) );
  AND U30557 ( .A(n30375), .B(n30376), .Z(n30157) );
  NANDN U30558 ( .A(n30377), .B(n30378), .Z(n30376) );
  NANDN U30559 ( .A(n30379), .B(n30380), .Z(n30378) );
  NANDN U30560 ( .A(n30380), .B(n30379), .Z(n30375) );
  ANDN U30561 ( .B(B[167]), .A(n56), .Z(n30159) );
  XNOR U30562 ( .A(n30167), .B(n30381), .Z(n30160) );
  XNOR U30563 ( .A(n30166), .B(n30164), .Z(n30381) );
  AND U30564 ( .A(n30382), .B(n30383), .Z(n30164) );
  NANDN U30565 ( .A(n30384), .B(n30385), .Z(n30383) );
  OR U30566 ( .A(n30386), .B(n30387), .Z(n30385) );
  NAND U30567 ( .A(n30387), .B(n30386), .Z(n30382) );
  ANDN U30568 ( .B(B[168]), .A(n57), .Z(n30166) );
  XNOR U30569 ( .A(n30174), .B(n30388), .Z(n30167) );
  XNOR U30570 ( .A(n30173), .B(n30171), .Z(n30388) );
  AND U30571 ( .A(n30389), .B(n30390), .Z(n30171) );
  NANDN U30572 ( .A(n30391), .B(n30392), .Z(n30390) );
  NANDN U30573 ( .A(n30393), .B(n30394), .Z(n30392) );
  NANDN U30574 ( .A(n30394), .B(n30393), .Z(n30389) );
  ANDN U30575 ( .B(B[169]), .A(n58), .Z(n30173) );
  XNOR U30576 ( .A(n30181), .B(n30395), .Z(n30174) );
  XNOR U30577 ( .A(n30180), .B(n30178), .Z(n30395) );
  AND U30578 ( .A(n30396), .B(n30397), .Z(n30178) );
  NANDN U30579 ( .A(n30398), .B(n30399), .Z(n30397) );
  OR U30580 ( .A(n30400), .B(n30401), .Z(n30399) );
  NAND U30581 ( .A(n30401), .B(n30400), .Z(n30396) );
  ANDN U30582 ( .B(B[170]), .A(n59), .Z(n30180) );
  XNOR U30583 ( .A(n30188), .B(n30402), .Z(n30181) );
  XNOR U30584 ( .A(n30187), .B(n30185), .Z(n30402) );
  AND U30585 ( .A(n30403), .B(n30404), .Z(n30185) );
  NANDN U30586 ( .A(n30405), .B(n30406), .Z(n30404) );
  NANDN U30587 ( .A(n30407), .B(n30408), .Z(n30406) );
  NANDN U30588 ( .A(n30408), .B(n30407), .Z(n30403) );
  ANDN U30589 ( .B(B[171]), .A(n60), .Z(n30187) );
  XNOR U30590 ( .A(n30195), .B(n30409), .Z(n30188) );
  XNOR U30591 ( .A(n30194), .B(n30192), .Z(n30409) );
  AND U30592 ( .A(n30410), .B(n30411), .Z(n30192) );
  NANDN U30593 ( .A(n30412), .B(n30413), .Z(n30411) );
  OR U30594 ( .A(n30414), .B(n30415), .Z(n30413) );
  NAND U30595 ( .A(n30415), .B(n30414), .Z(n30410) );
  ANDN U30596 ( .B(B[172]), .A(n61), .Z(n30194) );
  XNOR U30597 ( .A(n30202), .B(n30416), .Z(n30195) );
  XNOR U30598 ( .A(n30201), .B(n30199), .Z(n30416) );
  AND U30599 ( .A(n30417), .B(n30418), .Z(n30199) );
  NANDN U30600 ( .A(n30419), .B(n30420), .Z(n30418) );
  NANDN U30601 ( .A(n30421), .B(n30422), .Z(n30420) );
  NANDN U30602 ( .A(n30422), .B(n30421), .Z(n30417) );
  ANDN U30603 ( .B(B[173]), .A(n62), .Z(n30201) );
  XNOR U30604 ( .A(n30209), .B(n30423), .Z(n30202) );
  XNOR U30605 ( .A(n30208), .B(n30206), .Z(n30423) );
  AND U30606 ( .A(n30424), .B(n30425), .Z(n30206) );
  NANDN U30607 ( .A(n30426), .B(n30427), .Z(n30425) );
  OR U30608 ( .A(n30428), .B(n30429), .Z(n30427) );
  NAND U30609 ( .A(n30429), .B(n30428), .Z(n30424) );
  ANDN U30610 ( .B(B[174]), .A(n63), .Z(n30208) );
  XNOR U30611 ( .A(n30216), .B(n30430), .Z(n30209) );
  XNOR U30612 ( .A(n30215), .B(n30213), .Z(n30430) );
  AND U30613 ( .A(n30431), .B(n30432), .Z(n30213) );
  NANDN U30614 ( .A(n30433), .B(n30434), .Z(n30432) );
  NANDN U30615 ( .A(n30435), .B(n30436), .Z(n30434) );
  NANDN U30616 ( .A(n30436), .B(n30435), .Z(n30431) );
  ANDN U30617 ( .B(B[175]), .A(n64), .Z(n30215) );
  XNOR U30618 ( .A(n30223), .B(n30437), .Z(n30216) );
  XNOR U30619 ( .A(n30222), .B(n30220), .Z(n30437) );
  AND U30620 ( .A(n30438), .B(n30439), .Z(n30220) );
  NANDN U30621 ( .A(n30440), .B(n30441), .Z(n30439) );
  OR U30622 ( .A(n30442), .B(n30443), .Z(n30441) );
  NAND U30623 ( .A(n30443), .B(n30442), .Z(n30438) );
  ANDN U30624 ( .B(B[176]), .A(n65), .Z(n30222) );
  XNOR U30625 ( .A(n30230), .B(n30444), .Z(n30223) );
  XNOR U30626 ( .A(n30229), .B(n30227), .Z(n30444) );
  AND U30627 ( .A(n30445), .B(n30446), .Z(n30227) );
  NANDN U30628 ( .A(n30447), .B(n30448), .Z(n30446) );
  NANDN U30629 ( .A(n30449), .B(n30450), .Z(n30448) );
  NANDN U30630 ( .A(n30450), .B(n30449), .Z(n30445) );
  ANDN U30631 ( .B(B[177]), .A(n66), .Z(n30229) );
  XNOR U30632 ( .A(n30237), .B(n30451), .Z(n30230) );
  XNOR U30633 ( .A(n30236), .B(n30234), .Z(n30451) );
  AND U30634 ( .A(n30452), .B(n30453), .Z(n30234) );
  NANDN U30635 ( .A(n30454), .B(n30455), .Z(n30453) );
  OR U30636 ( .A(n30456), .B(n30457), .Z(n30455) );
  NAND U30637 ( .A(n30457), .B(n30456), .Z(n30452) );
  ANDN U30638 ( .B(B[178]), .A(n67), .Z(n30236) );
  XNOR U30639 ( .A(n30244), .B(n30458), .Z(n30237) );
  XNOR U30640 ( .A(n30243), .B(n30241), .Z(n30458) );
  AND U30641 ( .A(n30459), .B(n30460), .Z(n30241) );
  NANDN U30642 ( .A(n30461), .B(n30462), .Z(n30460) );
  NANDN U30643 ( .A(n30463), .B(n30464), .Z(n30462) );
  NANDN U30644 ( .A(n30464), .B(n30463), .Z(n30459) );
  ANDN U30645 ( .B(B[179]), .A(n68), .Z(n30243) );
  XNOR U30646 ( .A(n30251), .B(n30465), .Z(n30244) );
  XNOR U30647 ( .A(n30250), .B(n30248), .Z(n30465) );
  AND U30648 ( .A(n30466), .B(n30467), .Z(n30248) );
  NANDN U30649 ( .A(n30468), .B(n30469), .Z(n30467) );
  OR U30650 ( .A(n30470), .B(n30471), .Z(n30469) );
  NAND U30651 ( .A(n30471), .B(n30470), .Z(n30466) );
  ANDN U30652 ( .B(B[180]), .A(n69), .Z(n30250) );
  XNOR U30653 ( .A(n30258), .B(n30472), .Z(n30251) );
  XNOR U30654 ( .A(n30257), .B(n30255), .Z(n30472) );
  AND U30655 ( .A(n30473), .B(n30474), .Z(n30255) );
  NANDN U30656 ( .A(n30475), .B(n30476), .Z(n30474) );
  NANDN U30657 ( .A(n30477), .B(n30478), .Z(n30476) );
  NANDN U30658 ( .A(n30478), .B(n30477), .Z(n30473) );
  ANDN U30659 ( .B(B[181]), .A(n70), .Z(n30257) );
  XNOR U30660 ( .A(n30265), .B(n30479), .Z(n30258) );
  XNOR U30661 ( .A(n30264), .B(n30262), .Z(n30479) );
  AND U30662 ( .A(n30480), .B(n30481), .Z(n30262) );
  NANDN U30663 ( .A(n30482), .B(n30483), .Z(n30481) );
  OR U30664 ( .A(n30484), .B(n30485), .Z(n30483) );
  NAND U30665 ( .A(n30485), .B(n30484), .Z(n30480) );
  ANDN U30666 ( .B(B[182]), .A(n71), .Z(n30264) );
  XNOR U30667 ( .A(n30272), .B(n30486), .Z(n30265) );
  XNOR U30668 ( .A(n30271), .B(n30269), .Z(n30486) );
  AND U30669 ( .A(n30487), .B(n30488), .Z(n30269) );
  NANDN U30670 ( .A(n30489), .B(n30490), .Z(n30488) );
  NANDN U30671 ( .A(n30491), .B(n30492), .Z(n30490) );
  NANDN U30672 ( .A(n30492), .B(n30491), .Z(n30487) );
  ANDN U30673 ( .B(B[183]), .A(n72), .Z(n30271) );
  XNOR U30674 ( .A(n30279), .B(n30493), .Z(n30272) );
  XNOR U30675 ( .A(n30278), .B(n30276), .Z(n30493) );
  AND U30676 ( .A(n30494), .B(n30495), .Z(n30276) );
  NANDN U30677 ( .A(n30496), .B(n30497), .Z(n30495) );
  OR U30678 ( .A(n30498), .B(n30499), .Z(n30497) );
  NAND U30679 ( .A(n30499), .B(n30498), .Z(n30494) );
  ANDN U30680 ( .B(B[184]), .A(n73), .Z(n30278) );
  XNOR U30681 ( .A(n30286), .B(n30500), .Z(n30279) );
  XNOR U30682 ( .A(n30285), .B(n30283), .Z(n30500) );
  AND U30683 ( .A(n30501), .B(n30502), .Z(n30283) );
  NANDN U30684 ( .A(n30503), .B(n30504), .Z(n30502) );
  NANDN U30685 ( .A(n30505), .B(n30506), .Z(n30504) );
  NANDN U30686 ( .A(n30506), .B(n30505), .Z(n30501) );
  ANDN U30687 ( .B(B[185]), .A(n74), .Z(n30285) );
  XNOR U30688 ( .A(n30293), .B(n30507), .Z(n30286) );
  XNOR U30689 ( .A(n30292), .B(n30290), .Z(n30507) );
  AND U30690 ( .A(n30508), .B(n30509), .Z(n30290) );
  NANDN U30691 ( .A(n30510), .B(n30511), .Z(n30509) );
  OR U30692 ( .A(n30512), .B(n30513), .Z(n30511) );
  NAND U30693 ( .A(n30513), .B(n30512), .Z(n30508) );
  ANDN U30694 ( .B(B[186]), .A(n75), .Z(n30292) );
  XNOR U30695 ( .A(n30300), .B(n30514), .Z(n30293) );
  XNOR U30696 ( .A(n30299), .B(n30297), .Z(n30514) );
  AND U30697 ( .A(n30515), .B(n30516), .Z(n30297) );
  NANDN U30698 ( .A(n30517), .B(n30518), .Z(n30516) );
  NANDN U30699 ( .A(n30519), .B(n30520), .Z(n30518) );
  NANDN U30700 ( .A(n30520), .B(n30519), .Z(n30515) );
  ANDN U30701 ( .B(B[187]), .A(n76), .Z(n30299) );
  XNOR U30702 ( .A(n30307), .B(n30521), .Z(n30300) );
  XNOR U30703 ( .A(n30306), .B(n30304), .Z(n30521) );
  AND U30704 ( .A(n30522), .B(n30523), .Z(n30304) );
  NANDN U30705 ( .A(n30524), .B(n30525), .Z(n30523) );
  OR U30706 ( .A(n30526), .B(n30527), .Z(n30525) );
  NAND U30707 ( .A(n30527), .B(n30526), .Z(n30522) );
  ANDN U30708 ( .B(B[188]), .A(n77), .Z(n30306) );
  XNOR U30709 ( .A(n30314), .B(n30528), .Z(n30307) );
  XNOR U30710 ( .A(n30313), .B(n30311), .Z(n30528) );
  AND U30711 ( .A(n30529), .B(n30530), .Z(n30311) );
  NANDN U30712 ( .A(n30531), .B(n30532), .Z(n30530) );
  NANDN U30713 ( .A(n30533), .B(n30534), .Z(n30532) );
  NANDN U30714 ( .A(n30534), .B(n30533), .Z(n30529) );
  ANDN U30715 ( .B(B[189]), .A(n78), .Z(n30313) );
  XNOR U30716 ( .A(n30321), .B(n30535), .Z(n30314) );
  XNOR U30717 ( .A(n30320), .B(n30318), .Z(n30535) );
  AND U30718 ( .A(n30536), .B(n30537), .Z(n30318) );
  NANDN U30719 ( .A(n30538), .B(n30539), .Z(n30537) );
  OR U30720 ( .A(n30540), .B(n30541), .Z(n30539) );
  NAND U30721 ( .A(n30541), .B(n30540), .Z(n30536) );
  ANDN U30722 ( .B(B[190]), .A(n79), .Z(n30320) );
  XNOR U30723 ( .A(n30328), .B(n30542), .Z(n30321) );
  XNOR U30724 ( .A(n30327), .B(n30325), .Z(n30542) );
  AND U30725 ( .A(n30543), .B(n30544), .Z(n30325) );
  NANDN U30726 ( .A(n30545), .B(n30546), .Z(n30544) );
  NANDN U30727 ( .A(n30547), .B(n30548), .Z(n30546) );
  NANDN U30728 ( .A(n30548), .B(n30547), .Z(n30543) );
  ANDN U30729 ( .B(B[191]), .A(n80), .Z(n30327) );
  XNOR U30730 ( .A(n30335), .B(n30549), .Z(n30328) );
  XNOR U30731 ( .A(n30334), .B(n30332), .Z(n30549) );
  AND U30732 ( .A(n30550), .B(n30551), .Z(n30332) );
  NANDN U30733 ( .A(n30552), .B(n30553), .Z(n30551) );
  OR U30734 ( .A(n30554), .B(n30555), .Z(n30553) );
  NAND U30735 ( .A(n30555), .B(n30554), .Z(n30550) );
  ANDN U30736 ( .B(B[192]), .A(n81), .Z(n30334) );
  XNOR U30737 ( .A(n30342), .B(n30556), .Z(n30335) );
  XNOR U30738 ( .A(n30341), .B(n30339), .Z(n30556) );
  AND U30739 ( .A(n30557), .B(n30558), .Z(n30339) );
  NANDN U30740 ( .A(n30559), .B(n30560), .Z(n30558) );
  NAND U30741 ( .A(n30561), .B(n30562), .Z(n30560) );
  ANDN U30742 ( .B(B[193]), .A(n82), .Z(n30341) );
  XOR U30743 ( .A(n30348), .B(n30563), .Z(n30342) );
  XNOR U30744 ( .A(n30346), .B(n30349), .Z(n30563) );
  NAND U30745 ( .A(A[2]), .B(B[194]), .Z(n30349) );
  NANDN U30746 ( .A(n30564), .B(n30565), .Z(n30346) );
  AND U30747 ( .A(A[0]), .B(B[195]), .Z(n30565) );
  XNOR U30748 ( .A(n30351), .B(n30566), .Z(n30348) );
  NAND U30749 ( .A(A[0]), .B(B[196]), .Z(n30566) );
  NAND U30750 ( .A(B[195]), .B(A[1]), .Z(n30351) );
  NAND U30751 ( .A(n30567), .B(n30568), .Z(n404) );
  NANDN U30752 ( .A(n30569), .B(n30570), .Z(n30568) );
  OR U30753 ( .A(n30571), .B(n30572), .Z(n30570) );
  NAND U30754 ( .A(n30572), .B(n30571), .Z(n30567) );
  XOR U30755 ( .A(n406), .B(n405), .Z(\A1[193] ) );
  XOR U30756 ( .A(n30572), .B(n30573), .Z(n405) );
  XNOR U30757 ( .A(n30571), .B(n30569), .Z(n30573) );
  AND U30758 ( .A(n30574), .B(n30575), .Z(n30569) );
  NANDN U30759 ( .A(n30576), .B(n30577), .Z(n30575) );
  NANDN U30760 ( .A(n30578), .B(n30579), .Z(n30577) );
  NANDN U30761 ( .A(n30579), .B(n30578), .Z(n30574) );
  ANDN U30762 ( .B(B[164]), .A(n54), .Z(n30571) );
  XNOR U30763 ( .A(n30366), .B(n30580), .Z(n30572) );
  XNOR U30764 ( .A(n30365), .B(n30363), .Z(n30580) );
  AND U30765 ( .A(n30581), .B(n30582), .Z(n30363) );
  NANDN U30766 ( .A(n30583), .B(n30584), .Z(n30582) );
  OR U30767 ( .A(n30585), .B(n30586), .Z(n30584) );
  NAND U30768 ( .A(n30586), .B(n30585), .Z(n30581) );
  ANDN U30769 ( .B(B[165]), .A(n55), .Z(n30365) );
  XNOR U30770 ( .A(n30373), .B(n30587), .Z(n30366) );
  XNOR U30771 ( .A(n30372), .B(n30370), .Z(n30587) );
  AND U30772 ( .A(n30588), .B(n30589), .Z(n30370) );
  NANDN U30773 ( .A(n30590), .B(n30591), .Z(n30589) );
  NANDN U30774 ( .A(n30592), .B(n30593), .Z(n30591) );
  NANDN U30775 ( .A(n30593), .B(n30592), .Z(n30588) );
  ANDN U30776 ( .B(B[166]), .A(n56), .Z(n30372) );
  XNOR U30777 ( .A(n30380), .B(n30594), .Z(n30373) );
  XNOR U30778 ( .A(n30379), .B(n30377), .Z(n30594) );
  AND U30779 ( .A(n30595), .B(n30596), .Z(n30377) );
  NANDN U30780 ( .A(n30597), .B(n30598), .Z(n30596) );
  OR U30781 ( .A(n30599), .B(n30600), .Z(n30598) );
  NAND U30782 ( .A(n30600), .B(n30599), .Z(n30595) );
  ANDN U30783 ( .B(B[167]), .A(n57), .Z(n30379) );
  XNOR U30784 ( .A(n30387), .B(n30601), .Z(n30380) );
  XNOR U30785 ( .A(n30386), .B(n30384), .Z(n30601) );
  AND U30786 ( .A(n30602), .B(n30603), .Z(n30384) );
  NANDN U30787 ( .A(n30604), .B(n30605), .Z(n30603) );
  NANDN U30788 ( .A(n30606), .B(n30607), .Z(n30605) );
  NANDN U30789 ( .A(n30607), .B(n30606), .Z(n30602) );
  ANDN U30790 ( .B(B[168]), .A(n58), .Z(n30386) );
  XNOR U30791 ( .A(n30394), .B(n30608), .Z(n30387) );
  XNOR U30792 ( .A(n30393), .B(n30391), .Z(n30608) );
  AND U30793 ( .A(n30609), .B(n30610), .Z(n30391) );
  NANDN U30794 ( .A(n30611), .B(n30612), .Z(n30610) );
  OR U30795 ( .A(n30613), .B(n30614), .Z(n30612) );
  NAND U30796 ( .A(n30614), .B(n30613), .Z(n30609) );
  ANDN U30797 ( .B(B[169]), .A(n59), .Z(n30393) );
  XNOR U30798 ( .A(n30401), .B(n30615), .Z(n30394) );
  XNOR U30799 ( .A(n30400), .B(n30398), .Z(n30615) );
  AND U30800 ( .A(n30616), .B(n30617), .Z(n30398) );
  NANDN U30801 ( .A(n30618), .B(n30619), .Z(n30617) );
  NANDN U30802 ( .A(n30620), .B(n30621), .Z(n30619) );
  NANDN U30803 ( .A(n30621), .B(n30620), .Z(n30616) );
  ANDN U30804 ( .B(B[170]), .A(n60), .Z(n30400) );
  XNOR U30805 ( .A(n30408), .B(n30622), .Z(n30401) );
  XNOR U30806 ( .A(n30407), .B(n30405), .Z(n30622) );
  AND U30807 ( .A(n30623), .B(n30624), .Z(n30405) );
  NANDN U30808 ( .A(n30625), .B(n30626), .Z(n30624) );
  OR U30809 ( .A(n30627), .B(n30628), .Z(n30626) );
  NAND U30810 ( .A(n30628), .B(n30627), .Z(n30623) );
  ANDN U30811 ( .B(B[171]), .A(n61), .Z(n30407) );
  XNOR U30812 ( .A(n30415), .B(n30629), .Z(n30408) );
  XNOR U30813 ( .A(n30414), .B(n30412), .Z(n30629) );
  AND U30814 ( .A(n30630), .B(n30631), .Z(n30412) );
  NANDN U30815 ( .A(n30632), .B(n30633), .Z(n30631) );
  NANDN U30816 ( .A(n30634), .B(n30635), .Z(n30633) );
  NANDN U30817 ( .A(n30635), .B(n30634), .Z(n30630) );
  ANDN U30818 ( .B(B[172]), .A(n62), .Z(n30414) );
  XNOR U30819 ( .A(n30422), .B(n30636), .Z(n30415) );
  XNOR U30820 ( .A(n30421), .B(n30419), .Z(n30636) );
  AND U30821 ( .A(n30637), .B(n30638), .Z(n30419) );
  NANDN U30822 ( .A(n30639), .B(n30640), .Z(n30638) );
  OR U30823 ( .A(n30641), .B(n30642), .Z(n30640) );
  NAND U30824 ( .A(n30642), .B(n30641), .Z(n30637) );
  ANDN U30825 ( .B(B[173]), .A(n63), .Z(n30421) );
  XNOR U30826 ( .A(n30429), .B(n30643), .Z(n30422) );
  XNOR U30827 ( .A(n30428), .B(n30426), .Z(n30643) );
  AND U30828 ( .A(n30644), .B(n30645), .Z(n30426) );
  NANDN U30829 ( .A(n30646), .B(n30647), .Z(n30645) );
  NANDN U30830 ( .A(n30648), .B(n30649), .Z(n30647) );
  NANDN U30831 ( .A(n30649), .B(n30648), .Z(n30644) );
  ANDN U30832 ( .B(B[174]), .A(n64), .Z(n30428) );
  XNOR U30833 ( .A(n30436), .B(n30650), .Z(n30429) );
  XNOR U30834 ( .A(n30435), .B(n30433), .Z(n30650) );
  AND U30835 ( .A(n30651), .B(n30652), .Z(n30433) );
  NANDN U30836 ( .A(n30653), .B(n30654), .Z(n30652) );
  OR U30837 ( .A(n30655), .B(n30656), .Z(n30654) );
  NAND U30838 ( .A(n30656), .B(n30655), .Z(n30651) );
  ANDN U30839 ( .B(B[175]), .A(n65), .Z(n30435) );
  XNOR U30840 ( .A(n30443), .B(n30657), .Z(n30436) );
  XNOR U30841 ( .A(n30442), .B(n30440), .Z(n30657) );
  AND U30842 ( .A(n30658), .B(n30659), .Z(n30440) );
  NANDN U30843 ( .A(n30660), .B(n30661), .Z(n30659) );
  NANDN U30844 ( .A(n30662), .B(n30663), .Z(n30661) );
  NANDN U30845 ( .A(n30663), .B(n30662), .Z(n30658) );
  ANDN U30846 ( .B(B[176]), .A(n66), .Z(n30442) );
  XNOR U30847 ( .A(n30450), .B(n30664), .Z(n30443) );
  XNOR U30848 ( .A(n30449), .B(n30447), .Z(n30664) );
  AND U30849 ( .A(n30665), .B(n30666), .Z(n30447) );
  NANDN U30850 ( .A(n30667), .B(n30668), .Z(n30666) );
  OR U30851 ( .A(n30669), .B(n30670), .Z(n30668) );
  NAND U30852 ( .A(n30670), .B(n30669), .Z(n30665) );
  ANDN U30853 ( .B(B[177]), .A(n67), .Z(n30449) );
  XNOR U30854 ( .A(n30457), .B(n30671), .Z(n30450) );
  XNOR U30855 ( .A(n30456), .B(n30454), .Z(n30671) );
  AND U30856 ( .A(n30672), .B(n30673), .Z(n30454) );
  NANDN U30857 ( .A(n30674), .B(n30675), .Z(n30673) );
  NANDN U30858 ( .A(n30676), .B(n30677), .Z(n30675) );
  NANDN U30859 ( .A(n30677), .B(n30676), .Z(n30672) );
  ANDN U30860 ( .B(B[178]), .A(n68), .Z(n30456) );
  XNOR U30861 ( .A(n30464), .B(n30678), .Z(n30457) );
  XNOR U30862 ( .A(n30463), .B(n30461), .Z(n30678) );
  AND U30863 ( .A(n30679), .B(n30680), .Z(n30461) );
  NANDN U30864 ( .A(n30681), .B(n30682), .Z(n30680) );
  OR U30865 ( .A(n30683), .B(n30684), .Z(n30682) );
  NAND U30866 ( .A(n30684), .B(n30683), .Z(n30679) );
  ANDN U30867 ( .B(B[179]), .A(n69), .Z(n30463) );
  XNOR U30868 ( .A(n30471), .B(n30685), .Z(n30464) );
  XNOR U30869 ( .A(n30470), .B(n30468), .Z(n30685) );
  AND U30870 ( .A(n30686), .B(n30687), .Z(n30468) );
  NANDN U30871 ( .A(n30688), .B(n30689), .Z(n30687) );
  NANDN U30872 ( .A(n30690), .B(n30691), .Z(n30689) );
  NANDN U30873 ( .A(n30691), .B(n30690), .Z(n30686) );
  ANDN U30874 ( .B(B[180]), .A(n70), .Z(n30470) );
  XNOR U30875 ( .A(n30478), .B(n30692), .Z(n30471) );
  XNOR U30876 ( .A(n30477), .B(n30475), .Z(n30692) );
  AND U30877 ( .A(n30693), .B(n30694), .Z(n30475) );
  NANDN U30878 ( .A(n30695), .B(n30696), .Z(n30694) );
  OR U30879 ( .A(n30697), .B(n30698), .Z(n30696) );
  NAND U30880 ( .A(n30698), .B(n30697), .Z(n30693) );
  ANDN U30881 ( .B(B[181]), .A(n71), .Z(n30477) );
  XNOR U30882 ( .A(n30485), .B(n30699), .Z(n30478) );
  XNOR U30883 ( .A(n30484), .B(n30482), .Z(n30699) );
  AND U30884 ( .A(n30700), .B(n30701), .Z(n30482) );
  NANDN U30885 ( .A(n30702), .B(n30703), .Z(n30701) );
  NANDN U30886 ( .A(n30704), .B(n30705), .Z(n30703) );
  NANDN U30887 ( .A(n30705), .B(n30704), .Z(n30700) );
  ANDN U30888 ( .B(B[182]), .A(n72), .Z(n30484) );
  XNOR U30889 ( .A(n30492), .B(n30706), .Z(n30485) );
  XNOR U30890 ( .A(n30491), .B(n30489), .Z(n30706) );
  AND U30891 ( .A(n30707), .B(n30708), .Z(n30489) );
  NANDN U30892 ( .A(n30709), .B(n30710), .Z(n30708) );
  OR U30893 ( .A(n30711), .B(n30712), .Z(n30710) );
  NAND U30894 ( .A(n30712), .B(n30711), .Z(n30707) );
  ANDN U30895 ( .B(B[183]), .A(n73), .Z(n30491) );
  XNOR U30896 ( .A(n30499), .B(n30713), .Z(n30492) );
  XNOR U30897 ( .A(n30498), .B(n30496), .Z(n30713) );
  AND U30898 ( .A(n30714), .B(n30715), .Z(n30496) );
  NANDN U30899 ( .A(n30716), .B(n30717), .Z(n30715) );
  NANDN U30900 ( .A(n30718), .B(n30719), .Z(n30717) );
  NANDN U30901 ( .A(n30719), .B(n30718), .Z(n30714) );
  ANDN U30902 ( .B(B[184]), .A(n74), .Z(n30498) );
  XNOR U30903 ( .A(n30506), .B(n30720), .Z(n30499) );
  XNOR U30904 ( .A(n30505), .B(n30503), .Z(n30720) );
  AND U30905 ( .A(n30721), .B(n30722), .Z(n30503) );
  NANDN U30906 ( .A(n30723), .B(n30724), .Z(n30722) );
  OR U30907 ( .A(n30725), .B(n30726), .Z(n30724) );
  NAND U30908 ( .A(n30726), .B(n30725), .Z(n30721) );
  ANDN U30909 ( .B(B[185]), .A(n75), .Z(n30505) );
  XNOR U30910 ( .A(n30513), .B(n30727), .Z(n30506) );
  XNOR U30911 ( .A(n30512), .B(n30510), .Z(n30727) );
  AND U30912 ( .A(n30728), .B(n30729), .Z(n30510) );
  NANDN U30913 ( .A(n30730), .B(n30731), .Z(n30729) );
  NANDN U30914 ( .A(n30732), .B(n30733), .Z(n30731) );
  NANDN U30915 ( .A(n30733), .B(n30732), .Z(n30728) );
  ANDN U30916 ( .B(B[186]), .A(n76), .Z(n30512) );
  XNOR U30917 ( .A(n30520), .B(n30734), .Z(n30513) );
  XNOR U30918 ( .A(n30519), .B(n30517), .Z(n30734) );
  AND U30919 ( .A(n30735), .B(n30736), .Z(n30517) );
  NANDN U30920 ( .A(n30737), .B(n30738), .Z(n30736) );
  OR U30921 ( .A(n30739), .B(n30740), .Z(n30738) );
  NAND U30922 ( .A(n30740), .B(n30739), .Z(n30735) );
  ANDN U30923 ( .B(B[187]), .A(n77), .Z(n30519) );
  XNOR U30924 ( .A(n30527), .B(n30741), .Z(n30520) );
  XNOR U30925 ( .A(n30526), .B(n30524), .Z(n30741) );
  AND U30926 ( .A(n30742), .B(n30743), .Z(n30524) );
  NANDN U30927 ( .A(n30744), .B(n30745), .Z(n30743) );
  NANDN U30928 ( .A(n30746), .B(n30747), .Z(n30745) );
  NANDN U30929 ( .A(n30747), .B(n30746), .Z(n30742) );
  ANDN U30930 ( .B(B[188]), .A(n78), .Z(n30526) );
  XNOR U30931 ( .A(n30534), .B(n30748), .Z(n30527) );
  XNOR U30932 ( .A(n30533), .B(n30531), .Z(n30748) );
  AND U30933 ( .A(n30749), .B(n30750), .Z(n30531) );
  NANDN U30934 ( .A(n30751), .B(n30752), .Z(n30750) );
  OR U30935 ( .A(n30753), .B(n30754), .Z(n30752) );
  NAND U30936 ( .A(n30754), .B(n30753), .Z(n30749) );
  ANDN U30937 ( .B(B[189]), .A(n79), .Z(n30533) );
  XNOR U30938 ( .A(n30541), .B(n30755), .Z(n30534) );
  XNOR U30939 ( .A(n30540), .B(n30538), .Z(n30755) );
  AND U30940 ( .A(n30756), .B(n30757), .Z(n30538) );
  NANDN U30941 ( .A(n30758), .B(n30759), .Z(n30757) );
  NANDN U30942 ( .A(n30760), .B(n30761), .Z(n30759) );
  NANDN U30943 ( .A(n30761), .B(n30760), .Z(n30756) );
  ANDN U30944 ( .B(B[190]), .A(n80), .Z(n30540) );
  XNOR U30945 ( .A(n30548), .B(n30762), .Z(n30541) );
  XNOR U30946 ( .A(n30547), .B(n30545), .Z(n30762) );
  AND U30947 ( .A(n30763), .B(n30764), .Z(n30545) );
  NANDN U30948 ( .A(n30765), .B(n30766), .Z(n30764) );
  OR U30949 ( .A(n30767), .B(n30768), .Z(n30766) );
  NAND U30950 ( .A(n30768), .B(n30767), .Z(n30763) );
  ANDN U30951 ( .B(B[191]), .A(n81), .Z(n30547) );
  XNOR U30952 ( .A(n30555), .B(n30769), .Z(n30548) );
  XNOR U30953 ( .A(n30554), .B(n30552), .Z(n30769) );
  AND U30954 ( .A(n30770), .B(n30771), .Z(n30552) );
  NANDN U30955 ( .A(n30772), .B(n30773), .Z(n30771) );
  NAND U30956 ( .A(n30774), .B(n30775), .Z(n30773) );
  ANDN U30957 ( .B(B[192]), .A(n82), .Z(n30554) );
  XOR U30958 ( .A(n30561), .B(n30776), .Z(n30555) );
  XNOR U30959 ( .A(n30559), .B(n30562), .Z(n30776) );
  NAND U30960 ( .A(A[2]), .B(B[193]), .Z(n30562) );
  NANDN U30961 ( .A(n30777), .B(n30778), .Z(n30559) );
  AND U30962 ( .A(A[0]), .B(B[194]), .Z(n30778) );
  XNOR U30963 ( .A(n30564), .B(n30779), .Z(n30561) );
  NAND U30964 ( .A(A[0]), .B(B[195]), .Z(n30779) );
  NAND U30965 ( .A(B[194]), .B(A[1]), .Z(n30564) );
  NAND U30966 ( .A(n30780), .B(n30781), .Z(n406) );
  NANDN U30967 ( .A(n30782), .B(n30783), .Z(n30781) );
  OR U30968 ( .A(n30784), .B(n30785), .Z(n30783) );
  NAND U30969 ( .A(n30785), .B(n30784), .Z(n30780) );
  XOR U30970 ( .A(n408), .B(n407), .Z(\A1[192] ) );
  XOR U30971 ( .A(n30785), .B(n30786), .Z(n407) );
  XNOR U30972 ( .A(n30784), .B(n30782), .Z(n30786) );
  AND U30973 ( .A(n30787), .B(n30788), .Z(n30782) );
  NANDN U30974 ( .A(n30789), .B(n30790), .Z(n30788) );
  NANDN U30975 ( .A(n30791), .B(n30792), .Z(n30790) );
  NANDN U30976 ( .A(n30792), .B(n30791), .Z(n30787) );
  ANDN U30977 ( .B(B[163]), .A(n54), .Z(n30784) );
  XNOR U30978 ( .A(n30579), .B(n30793), .Z(n30785) );
  XNOR U30979 ( .A(n30578), .B(n30576), .Z(n30793) );
  AND U30980 ( .A(n30794), .B(n30795), .Z(n30576) );
  NANDN U30981 ( .A(n30796), .B(n30797), .Z(n30795) );
  OR U30982 ( .A(n30798), .B(n30799), .Z(n30797) );
  NAND U30983 ( .A(n30799), .B(n30798), .Z(n30794) );
  ANDN U30984 ( .B(B[164]), .A(n55), .Z(n30578) );
  XNOR U30985 ( .A(n30586), .B(n30800), .Z(n30579) );
  XNOR U30986 ( .A(n30585), .B(n30583), .Z(n30800) );
  AND U30987 ( .A(n30801), .B(n30802), .Z(n30583) );
  NANDN U30988 ( .A(n30803), .B(n30804), .Z(n30802) );
  NANDN U30989 ( .A(n30805), .B(n30806), .Z(n30804) );
  NANDN U30990 ( .A(n30806), .B(n30805), .Z(n30801) );
  ANDN U30991 ( .B(B[165]), .A(n56), .Z(n30585) );
  XNOR U30992 ( .A(n30593), .B(n30807), .Z(n30586) );
  XNOR U30993 ( .A(n30592), .B(n30590), .Z(n30807) );
  AND U30994 ( .A(n30808), .B(n30809), .Z(n30590) );
  NANDN U30995 ( .A(n30810), .B(n30811), .Z(n30809) );
  OR U30996 ( .A(n30812), .B(n30813), .Z(n30811) );
  NAND U30997 ( .A(n30813), .B(n30812), .Z(n30808) );
  ANDN U30998 ( .B(B[166]), .A(n57), .Z(n30592) );
  XNOR U30999 ( .A(n30600), .B(n30814), .Z(n30593) );
  XNOR U31000 ( .A(n30599), .B(n30597), .Z(n30814) );
  AND U31001 ( .A(n30815), .B(n30816), .Z(n30597) );
  NANDN U31002 ( .A(n30817), .B(n30818), .Z(n30816) );
  NANDN U31003 ( .A(n30819), .B(n30820), .Z(n30818) );
  NANDN U31004 ( .A(n30820), .B(n30819), .Z(n30815) );
  ANDN U31005 ( .B(B[167]), .A(n58), .Z(n30599) );
  XNOR U31006 ( .A(n30607), .B(n30821), .Z(n30600) );
  XNOR U31007 ( .A(n30606), .B(n30604), .Z(n30821) );
  AND U31008 ( .A(n30822), .B(n30823), .Z(n30604) );
  NANDN U31009 ( .A(n30824), .B(n30825), .Z(n30823) );
  OR U31010 ( .A(n30826), .B(n30827), .Z(n30825) );
  NAND U31011 ( .A(n30827), .B(n30826), .Z(n30822) );
  ANDN U31012 ( .B(B[168]), .A(n59), .Z(n30606) );
  XNOR U31013 ( .A(n30614), .B(n30828), .Z(n30607) );
  XNOR U31014 ( .A(n30613), .B(n30611), .Z(n30828) );
  AND U31015 ( .A(n30829), .B(n30830), .Z(n30611) );
  NANDN U31016 ( .A(n30831), .B(n30832), .Z(n30830) );
  NANDN U31017 ( .A(n30833), .B(n30834), .Z(n30832) );
  NANDN U31018 ( .A(n30834), .B(n30833), .Z(n30829) );
  ANDN U31019 ( .B(B[169]), .A(n60), .Z(n30613) );
  XNOR U31020 ( .A(n30621), .B(n30835), .Z(n30614) );
  XNOR U31021 ( .A(n30620), .B(n30618), .Z(n30835) );
  AND U31022 ( .A(n30836), .B(n30837), .Z(n30618) );
  NANDN U31023 ( .A(n30838), .B(n30839), .Z(n30837) );
  OR U31024 ( .A(n30840), .B(n30841), .Z(n30839) );
  NAND U31025 ( .A(n30841), .B(n30840), .Z(n30836) );
  ANDN U31026 ( .B(B[170]), .A(n61), .Z(n30620) );
  XNOR U31027 ( .A(n30628), .B(n30842), .Z(n30621) );
  XNOR U31028 ( .A(n30627), .B(n30625), .Z(n30842) );
  AND U31029 ( .A(n30843), .B(n30844), .Z(n30625) );
  NANDN U31030 ( .A(n30845), .B(n30846), .Z(n30844) );
  NANDN U31031 ( .A(n30847), .B(n30848), .Z(n30846) );
  NANDN U31032 ( .A(n30848), .B(n30847), .Z(n30843) );
  ANDN U31033 ( .B(B[171]), .A(n62), .Z(n30627) );
  XNOR U31034 ( .A(n30635), .B(n30849), .Z(n30628) );
  XNOR U31035 ( .A(n30634), .B(n30632), .Z(n30849) );
  AND U31036 ( .A(n30850), .B(n30851), .Z(n30632) );
  NANDN U31037 ( .A(n30852), .B(n30853), .Z(n30851) );
  OR U31038 ( .A(n30854), .B(n30855), .Z(n30853) );
  NAND U31039 ( .A(n30855), .B(n30854), .Z(n30850) );
  ANDN U31040 ( .B(B[172]), .A(n63), .Z(n30634) );
  XNOR U31041 ( .A(n30642), .B(n30856), .Z(n30635) );
  XNOR U31042 ( .A(n30641), .B(n30639), .Z(n30856) );
  AND U31043 ( .A(n30857), .B(n30858), .Z(n30639) );
  NANDN U31044 ( .A(n30859), .B(n30860), .Z(n30858) );
  NANDN U31045 ( .A(n30861), .B(n30862), .Z(n30860) );
  NANDN U31046 ( .A(n30862), .B(n30861), .Z(n30857) );
  ANDN U31047 ( .B(B[173]), .A(n64), .Z(n30641) );
  XNOR U31048 ( .A(n30649), .B(n30863), .Z(n30642) );
  XNOR U31049 ( .A(n30648), .B(n30646), .Z(n30863) );
  AND U31050 ( .A(n30864), .B(n30865), .Z(n30646) );
  NANDN U31051 ( .A(n30866), .B(n30867), .Z(n30865) );
  OR U31052 ( .A(n30868), .B(n30869), .Z(n30867) );
  NAND U31053 ( .A(n30869), .B(n30868), .Z(n30864) );
  ANDN U31054 ( .B(B[174]), .A(n65), .Z(n30648) );
  XNOR U31055 ( .A(n30656), .B(n30870), .Z(n30649) );
  XNOR U31056 ( .A(n30655), .B(n30653), .Z(n30870) );
  AND U31057 ( .A(n30871), .B(n30872), .Z(n30653) );
  NANDN U31058 ( .A(n30873), .B(n30874), .Z(n30872) );
  NANDN U31059 ( .A(n30875), .B(n30876), .Z(n30874) );
  NANDN U31060 ( .A(n30876), .B(n30875), .Z(n30871) );
  ANDN U31061 ( .B(B[175]), .A(n66), .Z(n30655) );
  XNOR U31062 ( .A(n30663), .B(n30877), .Z(n30656) );
  XNOR U31063 ( .A(n30662), .B(n30660), .Z(n30877) );
  AND U31064 ( .A(n30878), .B(n30879), .Z(n30660) );
  NANDN U31065 ( .A(n30880), .B(n30881), .Z(n30879) );
  OR U31066 ( .A(n30882), .B(n30883), .Z(n30881) );
  NAND U31067 ( .A(n30883), .B(n30882), .Z(n30878) );
  ANDN U31068 ( .B(B[176]), .A(n67), .Z(n30662) );
  XNOR U31069 ( .A(n30670), .B(n30884), .Z(n30663) );
  XNOR U31070 ( .A(n30669), .B(n30667), .Z(n30884) );
  AND U31071 ( .A(n30885), .B(n30886), .Z(n30667) );
  NANDN U31072 ( .A(n30887), .B(n30888), .Z(n30886) );
  NANDN U31073 ( .A(n30889), .B(n30890), .Z(n30888) );
  NANDN U31074 ( .A(n30890), .B(n30889), .Z(n30885) );
  ANDN U31075 ( .B(B[177]), .A(n68), .Z(n30669) );
  XNOR U31076 ( .A(n30677), .B(n30891), .Z(n30670) );
  XNOR U31077 ( .A(n30676), .B(n30674), .Z(n30891) );
  AND U31078 ( .A(n30892), .B(n30893), .Z(n30674) );
  NANDN U31079 ( .A(n30894), .B(n30895), .Z(n30893) );
  OR U31080 ( .A(n30896), .B(n30897), .Z(n30895) );
  NAND U31081 ( .A(n30897), .B(n30896), .Z(n30892) );
  ANDN U31082 ( .B(B[178]), .A(n69), .Z(n30676) );
  XNOR U31083 ( .A(n30684), .B(n30898), .Z(n30677) );
  XNOR U31084 ( .A(n30683), .B(n30681), .Z(n30898) );
  AND U31085 ( .A(n30899), .B(n30900), .Z(n30681) );
  NANDN U31086 ( .A(n30901), .B(n30902), .Z(n30900) );
  NANDN U31087 ( .A(n30903), .B(n30904), .Z(n30902) );
  NANDN U31088 ( .A(n30904), .B(n30903), .Z(n30899) );
  ANDN U31089 ( .B(B[179]), .A(n70), .Z(n30683) );
  XNOR U31090 ( .A(n30691), .B(n30905), .Z(n30684) );
  XNOR U31091 ( .A(n30690), .B(n30688), .Z(n30905) );
  AND U31092 ( .A(n30906), .B(n30907), .Z(n30688) );
  NANDN U31093 ( .A(n30908), .B(n30909), .Z(n30907) );
  OR U31094 ( .A(n30910), .B(n30911), .Z(n30909) );
  NAND U31095 ( .A(n30911), .B(n30910), .Z(n30906) );
  ANDN U31096 ( .B(B[180]), .A(n71), .Z(n30690) );
  XNOR U31097 ( .A(n30698), .B(n30912), .Z(n30691) );
  XNOR U31098 ( .A(n30697), .B(n30695), .Z(n30912) );
  AND U31099 ( .A(n30913), .B(n30914), .Z(n30695) );
  NANDN U31100 ( .A(n30915), .B(n30916), .Z(n30914) );
  NANDN U31101 ( .A(n30917), .B(n30918), .Z(n30916) );
  NANDN U31102 ( .A(n30918), .B(n30917), .Z(n30913) );
  ANDN U31103 ( .B(B[181]), .A(n72), .Z(n30697) );
  XNOR U31104 ( .A(n30705), .B(n30919), .Z(n30698) );
  XNOR U31105 ( .A(n30704), .B(n30702), .Z(n30919) );
  AND U31106 ( .A(n30920), .B(n30921), .Z(n30702) );
  NANDN U31107 ( .A(n30922), .B(n30923), .Z(n30921) );
  OR U31108 ( .A(n30924), .B(n30925), .Z(n30923) );
  NAND U31109 ( .A(n30925), .B(n30924), .Z(n30920) );
  ANDN U31110 ( .B(B[182]), .A(n73), .Z(n30704) );
  XNOR U31111 ( .A(n30712), .B(n30926), .Z(n30705) );
  XNOR U31112 ( .A(n30711), .B(n30709), .Z(n30926) );
  AND U31113 ( .A(n30927), .B(n30928), .Z(n30709) );
  NANDN U31114 ( .A(n30929), .B(n30930), .Z(n30928) );
  NANDN U31115 ( .A(n30931), .B(n30932), .Z(n30930) );
  NANDN U31116 ( .A(n30932), .B(n30931), .Z(n30927) );
  ANDN U31117 ( .B(B[183]), .A(n74), .Z(n30711) );
  XNOR U31118 ( .A(n30719), .B(n30933), .Z(n30712) );
  XNOR U31119 ( .A(n30718), .B(n30716), .Z(n30933) );
  AND U31120 ( .A(n30934), .B(n30935), .Z(n30716) );
  NANDN U31121 ( .A(n30936), .B(n30937), .Z(n30935) );
  OR U31122 ( .A(n30938), .B(n30939), .Z(n30937) );
  NAND U31123 ( .A(n30939), .B(n30938), .Z(n30934) );
  ANDN U31124 ( .B(B[184]), .A(n75), .Z(n30718) );
  XNOR U31125 ( .A(n30726), .B(n30940), .Z(n30719) );
  XNOR U31126 ( .A(n30725), .B(n30723), .Z(n30940) );
  AND U31127 ( .A(n30941), .B(n30942), .Z(n30723) );
  NANDN U31128 ( .A(n30943), .B(n30944), .Z(n30942) );
  NANDN U31129 ( .A(n30945), .B(n30946), .Z(n30944) );
  NANDN U31130 ( .A(n30946), .B(n30945), .Z(n30941) );
  ANDN U31131 ( .B(B[185]), .A(n76), .Z(n30725) );
  XNOR U31132 ( .A(n30733), .B(n30947), .Z(n30726) );
  XNOR U31133 ( .A(n30732), .B(n30730), .Z(n30947) );
  AND U31134 ( .A(n30948), .B(n30949), .Z(n30730) );
  NANDN U31135 ( .A(n30950), .B(n30951), .Z(n30949) );
  OR U31136 ( .A(n30952), .B(n30953), .Z(n30951) );
  NAND U31137 ( .A(n30953), .B(n30952), .Z(n30948) );
  ANDN U31138 ( .B(B[186]), .A(n77), .Z(n30732) );
  XNOR U31139 ( .A(n30740), .B(n30954), .Z(n30733) );
  XNOR U31140 ( .A(n30739), .B(n30737), .Z(n30954) );
  AND U31141 ( .A(n30955), .B(n30956), .Z(n30737) );
  NANDN U31142 ( .A(n30957), .B(n30958), .Z(n30956) );
  NANDN U31143 ( .A(n30959), .B(n30960), .Z(n30958) );
  NANDN U31144 ( .A(n30960), .B(n30959), .Z(n30955) );
  ANDN U31145 ( .B(B[187]), .A(n78), .Z(n30739) );
  XNOR U31146 ( .A(n30747), .B(n30961), .Z(n30740) );
  XNOR U31147 ( .A(n30746), .B(n30744), .Z(n30961) );
  AND U31148 ( .A(n30962), .B(n30963), .Z(n30744) );
  NANDN U31149 ( .A(n30964), .B(n30965), .Z(n30963) );
  OR U31150 ( .A(n30966), .B(n30967), .Z(n30965) );
  NAND U31151 ( .A(n30967), .B(n30966), .Z(n30962) );
  ANDN U31152 ( .B(B[188]), .A(n79), .Z(n30746) );
  XNOR U31153 ( .A(n30754), .B(n30968), .Z(n30747) );
  XNOR U31154 ( .A(n30753), .B(n30751), .Z(n30968) );
  AND U31155 ( .A(n30969), .B(n30970), .Z(n30751) );
  NANDN U31156 ( .A(n30971), .B(n30972), .Z(n30970) );
  NANDN U31157 ( .A(n30973), .B(n30974), .Z(n30972) );
  NANDN U31158 ( .A(n30974), .B(n30973), .Z(n30969) );
  ANDN U31159 ( .B(B[189]), .A(n80), .Z(n30753) );
  XNOR U31160 ( .A(n30761), .B(n30975), .Z(n30754) );
  XNOR U31161 ( .A(n30760), .B(n30758), .Z(n30975) );
  AND U31162 ( .A(n30976), .B(n30977), .Z(n30758) );
  NANDN U31163 ( .A(n30978), .B(n30979), .Z(n30977) );
  OR U31164 ( .A(n30980), .B(n30981), .Z(n30979) );
  NAND U31165 ( .A(n30981), .B(n30980), .Z(n30976) );
  ANDN U31166 ( .B(B[190]), .A(n81), .Z(n30760) );
  XNOR U31167 ( .A(n30768), .B(n30982), .Z(n30761) );
  XNOR U31168 ( .A(n30767), .B(n30765), .Z(n30982) );
  AND U31169 ( .A(n30983), .B(n30984), .Z(n30765) );
  NANDN U31170 ( .A(n30985), .B(n30986), .Z(n30984) );
  NAND U31171 ( .A(n30987), .B(n30988), .Z(n30986) );
  ANDN U31172 ( .B(B[191]), .A(n82), .Z(n30767) );
  XOR U31173 ( .A(n30774), .B(n30989), .Z(n30768) );
  XNOR U31174 ( .A(n30772), .B(n30775), .Z(n30989) );
  NAND U31175 ( .A(A[2]), .B(B[192]), .Z(n30775) );
  NANDN U31176 ( .A(n30990), .B(n30991), .Z(n30772) );
  AND U31177 ( .A(A[0]), .B(B[193]), .Z(n30991) );
  XNOR U31178 ( .A(n30777), .B(n30992), .Z(n30774) );
  NAND U31179 ( .A(A[0]), .B(B[194]), .Z(n30992) );
  NAND U31180 ( .A(B[193]), .B(A[1]), .Z(n30777) );
  NAND U31181 ( .A(n30993), .B(n30994), .Z(n408) );
  NANDN U31182 ( .A(n30995), .B(n30996), .Z(n30994) );
  OR U31183 ( .A(n30997), .B(n30998), .Z(n30996) );
  NAND U31184 ( .A(n30998), .B(n30997), .Z(n30993) );
  XOR U31185 ( .A(n410), .B(n409), .Z(\A1[191] ) );
  XOR U31186 ( .A(n30998), .B(n30999), .Z(n409) );
  XNOR U31187 ( .A(n30997), .B(n30995), .Z(n30999) );
  AND U31188 ( .A(n31000), .B(n31001), .Z(n30995) );
  NANDN U31189 ( .A(n31002), .B(n31003), .Z(n31001) );
  NANDN U31190 ( .A(n31004), .B(n31005), .Z(n31003) );
  NANDN U31191 ( .A(n31005), .B(n31004), .Z(n31000) );
  ANDN U31192 ( .B(B[162]), .A(n54), .Z(n30997) );
  XNOR U31193 ( .A(n30792), .B(n31006), .Z(n30998) );
  XNOR U31194 ( .A(n30791), .B(n30789), .Z(n31006) );
  AND U31195 ( .A(n31007), .B(n31008), .Z(n30789) );
  NANDN U31196 ( .A(n31009), .B(n31010), .Z(n31008) );
  OR U31197 ( .A(n31011), .B(n31012), .Z(n31010) );
  NAND U31198 ( .A(n31012), .B(n31011), .Z(n31007) );
  ANDN U31199 ( .B(B[163]), .A(n55), .Z(n30791) );
  XNOR U31200 ( .A(n30799), .B(n31013), .Z(n30792) );
  XNOR U31201 ( .A(n30798), .B(n30796), .Z(n31013) );
  AND U31202 ( .A(n31014), .B(n31015), .Z(n30796) );
  NANDN U31203 ( .A(n31016), .B(n31017), .Z(n31015) );
  NANDN U31204 ( .A(n31018), .B(n31019), .Z(n31017) );
  NANDN U31205 ( .A(n31019), .B(n31018), .Z(n31014) );
  ANDN U31206 ( .B(B[164]), .A(n56), .Z(n30798) );
  XNOR U31207 ( .A(n30806), .B(n31020), .Z(n30799) );
  XNOR U31208 ( .A(n30805), .B(n30803), .Z(n31020) );
  AND U31209 ( .A(n31021), .B(n31022), .Z(n30803) );
  NANDN U31210 ( .A(n31023), .B(n31024), .Z(n31022) );
  OR U31211 ( .A(n31025), .B(n31026), .Z(n31024) );
  NAND U31212 ( .A(n31026), .B(n31025), .Z(n31021) );
  ANDN U31213 ( .B(B[165]), .A(n57), .Z(n30805) );
  XNOR U31214 ( .A(n30813), .B(n31027), .Z(n30806) );
  XNOR U31215 ( .A(n30812), .B(n30810), .Z(n31027) );
  AND U31216 ( .A(n31028), .B(n31029), .Z(n30810) );
  NANDN U31217 ( .A(n31030), .B(n31031), .Z(n31029) );
  NANDN U31218 ( .A(n31032), .B(n31033), .Z(n31031) );
  NANDN U31219 ( .A(n31033), .B(n31032), .Z(n31028) );
  ANDN U31220 ( .B(B[166]), .A(n58), .Z(n30812) );
  XNOR U31221 ( .A(n30820), .B(n31034), .Z(n30813) );
  XNOR U31222 ( .A(n30819), .B(n30817), .Z(n31034) );
  AND U31223 ( .A(n31035), .B(n31036), .Z(n30817) );
  NANDN U31224 ( .A(n31037), .B(n31038), .Z(n31036) );
  OR U31225 ( .A(n31039), .B(n31040), .Z(n31038) );
  NAND U31226 ( .A(n31040), .B(n31039), .Z(n31035) );
  ANDN U31227 ( .B(B[167]), .A(n59), .Z(n30819) );
  XNOR U31228 ( .A(n30827), .B(n31041), .Z(n30820) );
  XNOR U31229 ( .A(n30826), .B(n30824), .Z(n31041) );
  AND U31230 ( .A(n31042), .B(n31043), .Z(n30824) );
  NANDN U31231 ( .A(n31044), .B(n31045), .Z(n31043) );
  NANDN U31232 ( .A(n31046), .B(n31047), .Z(n31045) );
  NANDN U31233 ( .A(n31047), .B(n31046), .Z(n31042) );
  ANDN U31234 ( .B(B[168]), .A(n60), .Z(n30826) );
  XNOR U31235 ( .A(n30834), .B(n31048), .Z(n30827) );
  XNOR U31236 ( .A(n30833), .B(n30831), .Z(n31048) );
  AND U31237 ( .A(n31049), .B(n31050), .Z(n30831) );
  NANDN U31238 ( .A(n31051), .B(n31052), .Z(n31050) );
  OR U31239 ( .A(n31053), .B(n31054), .Z(n31052) );
  NAND U31240 ( .A(n31054), .B(n31053), .Z(n31049) );
  ANDN U31241 ( .B(B[169]), .A(n61), .Z(n30833) );
  XNOR U31242 ( .A(n30841), .B(n31055), .Z(n30834) );
  XNOR U31243 ( .A(n30840), .B(n30838), .Z(n31055) );
  AND U31244 ( .A(n31056), .B(n31057), .Z(n30838) );
  NANDN U31245 ( .A(n31058), .B(n31059), .Z(n31057) );
  NANDN U31246 ( .A(n31060), .B(n31061), .Z(n31059) );
  NANDN U31247 ( .A(n31061), .B(n31060), .Z(n31056) );
  ANDN U31248 ( .B(B[170]), .A(n62), .Z(n30840) );
  XNOR U31249 ( .A(n30848), .B(n31062), .Z(n30841) );
  XNOR U31250 ( .A(n30847), .B(n30845), .Z(n31062) );
  AND U31251 ( .A(n31063), .B(n31064), .Z(n30845) );
  NANDN U31252 ( .A(n31065), .B(n31066), .Z(n31064) );
  OR U31253 ( .A(n31067), .B(n31068), .Z(n31066) );
  NAND U31254 ( .A(n31068), .B(n31067), .Z(n31063) );
  ANDN U31255 ( .B(B[171]), .A(n63), .Z(n30847) );
  XNOR U31256 ( .A(n30855), .B(n31069), .Z(n30848) );
  XNOR U31257 ( .A(n30854), .B(n30852), .Z(n31069) );
  AND U31258 ( .A(n31070), .B(n31071), .Z(n30852) );
  NANDN U31259 ( .A(n31072), .B(n31073), .Z(n31071) );
  NANDN U31260 ( .A(n31074), .B(n31075), .Z(n31073) );
  NANDN U31261 ( .A(n31075), .B(n31074), .Z(n31070) );
  ANDN U31262 ( .B(B[172]), .A(n64), .Z(n30854) );
  XNOR U31263 ( .A(n30862), .B(n31076), .Z(n30855) );
  XNOR U31264 ( .A(n30861), .B(n30859), .Z(n31076) );
  AND U31265 ( .A(n31077), .B(n31078), .Z(n30859) );
  NANDN U31266 ( .A(n31079), .B(n31080), .Z(n31078) );
  OR U31267 ( .A(n31081), .B(n31082), .Z(n31080) );
  NAND U31268 ( .A(n31082), .B(n31081), .Z(n31077) );
  ANDN U31269 ( .B(B[173]), .A(n65), .Z(n30861) );
  XNOR U31270 ( .A(n30869), .B(n31083), .Z(n30862) );
  XNOR U31271 ( .A(n30868), .B(n30866), .Z(n31083) );
  AND U31272 ( .A(n31084), .B(n31085), .Z(n30866) );
  NANDN U31273 ( .A(n31086), .B(n31087), .Z(n31085) );
  NANDN U31274 ( .A(n31088), .B(n31089), .Z(n31087) );
  NANDN U31275 ( .A(n31089), .B(n31088), .Z(n31084) );
  ANDN U31276 ( .B(B[174]), .A(n66), .Z(n30868) );
  XNOR U31277 ( .A(n30876), .B(n31090), .Z(n30869) );
  XNOR U31278 ( .A(n30875), .B(n30873), .Z(n31090) );
  AND U31279 ( .A(n31091), .B(n31092), .Z(n30873) );
  NANDN U31280 ( .A(n31093), .B(n31094), .Z(n31092) );
  OR U31281 ( .A(n31095), .B(n31096), .Z(n31094) );
  NAND U31282 ( .A(n31096), .B(n31095), .Z(n31091) );
  ANDN U31283 ( .B(B[175]), .A(n67), .Z(n30875) );
  XNOR U31284 ( .A(n30883), .B(n31097), .Z(n30876) );
  XNOR U31285 ( .A(n30882), .B(n30880), .Z(n31097) );
  AND U31286 ( .A(n31098), .B(n31099), .Z(n30880) );
  NANDN U31287 ( .A(n31100), .B(n31101), .Z(n31099) );
  NANDN U31288 ( .A(n31102), .B(n31103), .Z(n31101) );
  NANDN U31289 ( .A(n31103), .B(n31102), .Z(n31098) );
  ANDN U31290 ( .B(B[176]), .A(n68), .Z(n30882) );
  XNOR U31291 ( .A(n30890), .B(n31104), .Z(n30883) );
  XNOR U31292 ( .A(n30889), .B(n30887), .Z(n31104) );
  AND U31293 ( .A(n31105), .B(n31106), .Z(n30887) );
  NANDN U31294 ( .A(n31107), .B(n31108), .Z(n31106) );
  OR U31295 ( .A(n31109), .B(n31110), .Z(n31108) );
  NAND U31296 ( .A(n31110), .B(n31109), .Z(n31105) );
  ANDN U31297 ( .B(B[177]), .A(n69), .Z(n30889) );
  XNOR U31298 ( .A(n30897), .B(n31111), .Z(n30890) );
  XNOR U31299 ( .A(n30896), .B(n30894), .Z(n31111) );
  AND U31300 ( .A(n31112), .B(n31113), .Z(n30894) );
  NANDN U31301 ( .A(n31114), .B(n31115), .Z(n31113) );
  NANDN U31302 ( .A(n31116), .B(n31117), .Z(n31115) );
  NANDN U31303 ( .A(n31117), .B(n31116), .Z(n31112) );
  ANDN U31304 ( .B(B[178]), .A(n70), .Z(n30896) );
  XNOR U31305 ( .A(n30904), .B(n31118), .Z(n30897) );
  XNOR U31306 ( .A(n30903), .B(n30901), .Z(n31118) );
  AND U31307 ( .A(n31119), .B(n31120), .Z(n30901) );
  NANDN U31308 ( .A(n31121), .B(n31122), .Z(n31120) );
  OR U31309 ( .A(n31123), .B(n31124), .Z(n31122) );
  NAND U31310 ( .A(n31124), .B(n31123), .Z(n31119) );
  ANDN U31311 ( .B(B[179]), .A(n71), .Z(n30903) );
  XNOR U31312 ( .A(n30911), .B(n31125), .Z(n30904) );
  XNOR U31313 ( .A(n30910), .B(n30908), .Z(n31125) );
  AND U31314 ( .A(n31126), .B(n31127), .Z(n30908) );
  NANDN U31315 ( .A(n31128), .B(n31129), .Z(n31127) );
  NANDN U31316 ( .A(n31130), .B(n31131), .Z(n31129) );
  NANDN U31317 ( .A(n31131), .B(n31130), .Z(n31126) );
  ANDN U31318 ( .B(B[180]), .A(n72), .Z(n30910) );
  XNOR U31319 ( .A(n30918), .B(n31132), .Z(n30911) );
  XNOR U31320 ( .A(n30917), .B(n30915), .Z(n31132) );
  AND U31321 ( .A(n31133), .B(n31134), .Z(n30915) );
  NANDN U31322 ( .A(n31135), .B(n31136), .Z(n31134) );
  OR U31323 ( .A(n31137), .B(n31138), .Z(n31136) );
  NAND U31324 ( .A(n31138), .B(n31137), .Z(n31133) );
  ANDN U31325 ( .B(B[181]), .A(n73), .Z(n30917) );
  XNOR U31326 ( .A(n30925), .B(n31139), .Z(n30918) );
  XNOR U31327 ( .A(n30924), .B(n30922), .Z(n31139) );
  AND U31328 ( .A(n31140), .B(n31141), .Z(n30922) );
  NANDN U31329 ( .A(n31142), .B(n31143), .Z(n31141) );
  NANDN U31330 ( .A(n31144), .B(n31145), .Z(n31143) );
  NANDN U31331 ( .A(n31145), .B(n31144), .Z(n31140) );
  ANDN U31332 ( .B(B[182]), .A(n74), .Z(n30924) );
  XNOR U31333 ( .A(n30932), .B(n31146), .Z(n30925) );
  XNOR U31334 ( .A(n30931), .B(n30929), .Z(n31146) );
  AND U31335 ( .A(n31147), .B(n31148), .Z(n30929) );
  NANDN U31336 ( .A(n31149), .B(n31150), .Z(n31148) );
  OR U31337 ( .A(n31151), .B(n31152), .Z(n31150) );
  NAND U31338 ( .A(n31152), .B(n31151), .Z(n31147) );
  ANDN U31339 ( .B(B[183]), .A(n75), .Z(n30931) );
  XNOR U31340 ( .A(n30939), .B(n31153), .Z(n30932) );
  XNOR U31341 ( .A(n30938), .B(n30936), .Z(n31153) );
  AND U31342 ( .A(n31154), .B(n31155), .Z(n30936) );
  NANDN U31343 ( .A(n31156), .B(n31157), .Z(n31155) );
  NANDN U31344 ( .A(n31158), .B(n31159), .Z(n31157) );
  NANDN U31345 ( .A(n31159), .B(n31158), .Z(n31154) );
  ANDN U31346 ( .B(B[184]), .A(n76), .Z(n30938) );
  XNOR U31347 ( .A(n30946), .B(n31160), .Z(n30939) );
  XNOR U31348 ( .A(n30945), .B(n30943), .Z(n31160) );
  AND U31349 ( .A(n31161), .B(n31162), .Z(n30943) );
  NANDN U31350 ( .A(n31163), .B(n31164), .Z(n31162) );
  OR U31351 ( .A(n31165), .B(n31166), .Z(n31164) );
  NAND U31352 ( .A(n31166), .B(n31165), .Z(n31161) );
  ANDN U31353 ( .B(B[185]), .A(n77), .Z(n30945) );
  XNOR U31354 ( .A(n30953), .B(n31167), .Z(n30946) );
  XNOR U31355 ( .A(n30952), .B(n30950), .Z(n31167) );
  AND U31356 ( .A(n31168), .B(n31169), .Z(n30950) );
  NANDN U31357 ( .A(n31170), .B(n31171), .Z(n31169) );
  NANDN U31358 ( .A(n31172), .B(n31173), .Z(n31171) );
  NANDN U31359 ( .A(n31173), .B(n31172), .Z(n31168) );
  ANDN U31360 ( .B(B[186]), .A(n78), .Z(n30952) );
  XNOR U31361 ( .A(n30960), .B(n31174), .Z(n30953) );
  XNOR U31362 ( .A(n30959), .B(n30957), .Z(n31174) );
  AND U31363 ( .A(n31175), .B(n31176), .Z(n30957) );
  NANDN U31364 ( .A(n31177), .B(n31178), .Z(n31176) );
  OR U31365 ( .A(n31179), .B(n31180), .Z(n31178) );
  NAND U31366 ( .A(n31180), .B(n31179), .Z(n31175) );
  ANDN U31367 ( .B(B[187]), .A(n79), .Z(n30959) );
  XNOR U31368 ( .A(n30967), .B(n31181), .Z(n30960) );
  XNOR U31369 ( .A(n30966), .B(n30964), .Z(n31181) );
  AND U31370 ( .A(n31182), .B(n31183), .Z(n30964) );
  NANDN U31371 ( .A(n31184), .B(n31185), .Z(n31183) );
  NANDN U31372 ( .A(n31186), .B(n31187), .Z(n31185) );
  NANDN U31373 ( .A(n31187), .B(n31186), .Z(n31182) );
  ANDN U31374 ( .B(B[188]), .A(n80), .Z(n30966) );
  XNOR U31375 ( .A(n30974), .B(n31188), .Z(n30967) );
  XNOR U31376 ( .A(n30973), .B(n30971), .Z(n31188) );
  AND U31377 ( .A(n31189), .B(n31190), .Z(n30971) );
  NANDN U31378 ( .A(n31191), .B(n31192), .Z(n31190) );
  OR U31379 ( .A(n31193), .B(n31194), .Z(n31192) );
  NAND U31380 ( .A(n31194), .B(n31193), .Z(n31189) );
  ANDN U31381 ( .B(B[189]), .A(n81), .Z(n30973) );
  XNOR U31382 ( .A(n30981), .B(n31195), .Z(n30974) );
  XNOR U31383 ( .A(n30980), .B(n30978), .Z(n31195) );
  AND U31384 ( .A(n31196), .B(n31197), .Z(n30978) );
  NANDN U31385 ( .A(n31198), .B(n31199), .Z(n31197) );
  NAND U31386 ( .A(n31200), .B(n31201), .Z(n31199) );
  ANDN U31387 ( .B(B[190]), .A(n82), .Z(n30980) );
  XOR U31388 ( .A(n30987), .B(n31202), .Z(n30981) );
  XNOR U31389 ( .A(n30985), .B(n30988), .Z(n31202) );
  NAND U31390 ( .A(A[2]), .B(B[191]), .Z(n30988) );
  NANDN U31391 ( .A(n31203), .B(n31204), .Z(n30985) );
  AND U31392 ( .A(A[0]), .B(B[192]), .Z(n31204) );
  XNOR U31393 ( .A(n30990), .B(n31205), .Z(n30987) );
  NAND U31394 ( .A(A[0]), .B(B[193]), .Z(n31205) );
  NAND U31395 ( .A(B[192]), .B(A[1]), .Z(n30990) );
  NAND U31396 ( .A(n31206), .B(n31207), .Z(n410) );
  NANDN U31397 ( .A(n31208), .B(n31209), .Z(n31207) );
  OR U31398 ( .A(n31210), .B(n31211), .Z(n31209) );
  NAND U31399 ( .A(n31211), .B(n31210), .Z(n31206) );
  XOR U31400 ( .A(n412), .B(n411), .Z(\A1[190] ) );
  XOR U31401 ( .A(n31211), .B(n31212), .Z(n411) );
  XNOR U31402 ( .A(n31210), .B(n31208), .Z(n31212) );
  AND U31403 ( .A(n31213), .B(n31214), .Z(n31208) );
  NANDN U31404 ( .A(n31215), .B(n31216), .Z(n31214) );
  NANDN U31405 ( .A(n31217), .B(n31218), .Z(n31216) );
  NANDN U31406 ( .A(n31218), .B(n31217), .Z(n31213) );
  ANDN U31407 ( .B(B[161]), .A(n54), .Z(n31210) );
  XNOR U31408 ( .A(n31005), .B(n31219), .Z(n31211) );
  XNOR U31409 ( .A(n31004), .B(n31002), .Z(n31219) );
  AND U31410 ( .A(n31220), .B(n31221), .Z(n31002) );
  NANDN U31411 ( .A(n31222), .B(n31223), .Z(n31221) );
  OR U31412 ( .A(n31224), .B(n31225), .Z(n31223) );
  NAND U31413 ( .A(n31225), .B(n31224), .Z(n31220) );
  ANDN U31414 ( .B(B[162]), .A(n55), .Z(n31004) );
  XNOR U31415 ( .A(n31012), .B(n31226), .Z(n31005) );
  XNOR U31416 ( .A(n31011), .B(n31009), .Z(n31226) );
  AND U31417 ( .A(n31227), .B(n31228), .Z(n31009) );
  NANDN U31418 ( .A(n31229), .B(n31230), .Z(n31228) );
  NANDN U31419 ( .A(n31231), .B(n31232), .Z(n31230) );
  NANDN U31420 ( .A(n31232), .B(n31231), .Z(n31227) );
  ANDN U31421 ( .B(B[163]), .A(n56), .Z(n31011) );
  XNOR U31422 ( .A(n31019), .B(n31233), .Z(n31012) );
  XNOR U31423 ( .A(n31018), .B(n31016), .Z(n31233) );
  AND U31424 ( .A(n31234), .B(n31235), .Z(n31016) );
  NANDN U31425 ( .A(n31236), .B(n31237), .Z(n31235) );
  OR U31426 ( .A(n31238), .B(n31239), .Z(n31237) );
  NAND U31427 ( .A(n31239), .B(n31238), .Z(n31234) );
  ANDN U31428 ( .B(B[164]), .A(n57), .Z(n31018) );
  XNOR U31429 ( .A(n31026), .B(n31240), .Z(n31019) );
  XNOR U31430 ( .A(n31025), .B(n31023), .Z(n31240) );
  AND U31431 ( .A(n31241), .B(n31242), .Z(n31023) );
  NANDN U31432 ( .A(n31243), .B(n31244), .Z(n31242) );
  NANDN U31433 ( .A(n31245), .B(n31246), .Z(n31244) );
  NANDN U31434 ( .A(n31246), .B(n31245), .Z(n31241) );
  ANDN U31435 ( .B(B[165]), .A(n58), .Z(n31025) );
  XNOR U31436 ( .A(n31033), .B(n31247), .Z(n31026) );
  XNOR U31437 ( .A(n31032), .B(n31030), .Z(n31247) );
  AND U31438 ( .A(n31248), .B(n31249), .Z(n31030) );
  NANDN U31439 ( .A(n31250), .B(n31251), .Z(n31249) );
  OR U31440 ( .A(n31252), .B(n31253), .Z(n31251) );
  NAND U31441 ( .A(n31253), .B(n31252), .Z(n31248) );
  ANDN U31442 ( .B(B[166]), .A(n59), .Z(n31032) );
  XNOR U31443 ( .A(n31040), .B(n31254), .Z(n31033) );
  XNOR U31444 ( .A(n31039), .B(n31037), .Z(n31254) );
  AND U31445 ( .A(n31255), .B(n31256), .Z(n31037) );
  NANDN U31446 ( .A(n31257), .B(n31258), .Z(n31256) );
  NANDN U31447 ( .A(n31259), .B(n31260), .Z(n31258) );
  NANDN U31448 ( .A(n31260), .B(n31259), .Z(n31255) );
  ANDN U31449 ( .B(B[167]), .A(n60), .Z(n31039) );
  XNOR U31450 ( .A(n31047), .B(n31261), .Z(n31040) );
  XNOR U31451 ( .A(n31046), .B(n31044), .Z(n31261) );
  AND U31452 ( .A(n31262), .B(n31263), .Z(n31044) );
  NANDN U31453 ( .A(n31264), .B(n31265), .Z(n31263) );
  OR U31454 ( .A(n31266), .B(n31267), .Z(n31265) );
  NAND U31455 ( .A(n31267), .B(n31266), .Z(n31262) );
  ANDN U31456 ( .B(B[168]), .A(n61), .Z(n31046) );
  XNOR U31457 ( .A(n31054), .B(n31268), .Z(n31047) );
  XNOR U31458 ( .A(n31053), .B(n31051), .Z(n31268) );
  AND U31459 ( .A(n31269), .B(n31270), .Z(n31051) );
  NANDN U31460 ( .A(n31271), .B(n31272), .Z(n31270) );
  NANDN U31461 ( .A(n31273), .B(n31274), .Z(n31272) );
  NANDN U31462 ( .A(n31274), .B(n31273), .Z(n31269) );
  ANDN U31463 ( .B(B[169]), .A(n62), .Z(n31053) );
  XNOR U31464 ( .A(n31061), .B(n31275), .Z(n31054) );
  XNOR U31465 ( .A(n31060), .B(n31058), .Z(n31275) );
  AND U31466 ( .A(n31276), .B(n31277), .Z(n31058) );
  NANDN U31467 ( .A(n31278), .B(n31279), .Z(n31277) );
  OR U31468 ( .A(n31280), .B(n31281), .Z(n31279) );
  NAND U31469 ( .A(n31281), .B(n31280), .Z(n31276) );
  ANDN U31470 ( .B(B[170]), .A(n63), .Z(n31060) );
  XNOR U31471 ( .A(n31068), .B(n31282), .Z(n31061) );
  XNOR U31472 ( .A(n31067), .B(n31065), .Z(n31282) );
  AND U31473 ( .A(n31283), .B(n31284), .Z(n31065) );
  NANDN U31474 ( .A(n31285), .B(n31286), .Z(n31284) );
  NANDN U31475 ( .A(n31287), .B(n31288), .Z(n31286) );
  NANDN U31476 ( .A(n31288), .B(n31287), .Z(n31283) );
  ANDN U31477 ( .B(B[171]), .A(n64), .Z(n31067) );
  XNOR U31478 ( .A(n31075), .B(n31289), .Z(n31068) );
  XNOR U31479 ( .A(n31074), .B(n31072), .Z(n31289) );
  AND U31480 ( .A(n31290), .B(n31291), .Z(n31072) );
  NANDN U31481 ( .A(n31292), .B(n31293), .Z(n31291) );
  OR U31482 ( .A(n31294), .B(n31295), .Z(n31293) );
  NAND U31483 ( .A(n31295), .B(n31294), .Z(n31290) );
  ANDN U31484 ( .B(B[172]), .A(n65), .Z(n31074) );
  XNOR U31485 ( .A(n31082), .B(n31296), .Z(n31075) );
  XNOR U31486 ( .A(n31081), .B(n31079), .Z(n31296) );
  AND U31487 ( .A(n31297), .B(n31298), .Z(n31079) );
  NANDN U31488 ( .A(n31299), .B(n31300), .Z(n31298) );
  NANDN U31489 ( .A(n31301), .B(n31302), .Z(n31300) );
  NANDN U31490 ( .A(n31302), .B(n31301), .Z(n31297) );
  ANDN U31491 ( .B(B[173]), .A(n66), .Z(n31081) );
  XNOR U31492 ( .A(n31089), .B(n31303), .Z(n31082) );
  XNOR U31493 ( .A(n31088), .B(n31086), .Z(n31303) );
  AND U31494 ( .A(n31304), .B(n31305), .Z(n31086) );
  NANDN U31495 ( .A(n31306), .B(n31307), .Z(n31305) );
  OR U31496 ( .A(n31308), .B(n31309), .Z(n31307) );
  NAND U31497 ( .A(n31309), .B(n31308), .Z(n31304) );
  ANDN U31498 ( .B(B[174]), .A(n67), .Z(n31088) );
  XNOR U31499 ( .A(n31096), .B(n31310), .Z(n31089) );
  XNOR U31500 ( .A(n31095), .B(n31093), .Z(n31310) );
  AND U31501 ( .A(n31311), .B(n31312), .Z(n31093) );
  NANDN U31502 ( .A(n31313), .B(n31314), .Z(n31312) );
  NANDN U31503 ( .A(n31315), .B(n31316), .Z(n31314) );
  NANDN U31504 ( .A(n31316), .B(n31315), .Z(n31311) );
  ANDN U31505 ( .B(B[175]), .A(n68), .Z(n31095) );
  XNOR U31506 ( .A(n31103), .B(n31317), .Z(n31096) );
  XNOR U31507 ( .A(n31102), .B(n31100), .Z(n31317) );
  AND U31508 ( .A(n31318), .B(n31319), .Z(n31100) );
  NANDN U31509 ( .A(n31320), .B(n31321), .Z(n31319) );
  OR U31510 ( .A(n31322), .B(n31323), .Z(n31321) );
  NAND U31511 ( .A(n31323), .B(n31322), .Z(n31318) );
  ANDN U31512 ( .B(B[176]), .A(n69), .Z(n31102) );
  XNOR U31513 ( .A(n31110), .B(n31324), .Z(n31103) );
  XNOR U31514 ( .A(n31109), .B(n31107), .Z(n31324) );
  AND U31515 ( .A(n31325), .B(n31326), .Z(n31107) );
  NANDN U31516 ( .A(n31327), .B(n31328), .Z(n31326) );
  NANDN U31517 ( .A(n31329), .B(n31330), .Z(n31328) );
  NANDN U31518 ( .A(n31330), .B(n31329), .Z(n31325) );
  ANDN U31519 ( .B(B[177]), .A(n70), .Z(n31109) );
  XNOR U31520 ( .A(n31117), .B(n31331), .Z(n31110) );
  XNOR U31521 ( .A(n31116), .B(n31114), .Z(n31331) );
  AND U31522 ( .A(n31332), .B(n31333), .Z(n31114) );
  NANDN U31523 ( .A(n31334), .B(n31335), .Z(n31333) );
  OR U31524 ( .A(n31336), .B(n31337), .Z(n31335) );
  NAND U31525 ( .A(n31337), .B(n31336), .Z(n31332) );
  ANDN U31526 ( .B(B[178]), .A(n71), .Z(n31116) );
  XNOR U31527 ( .A(n31124), .B(n31338), .Z(n31117) );
  XNOR U31528 ( .A(n31123), .B(n31121), .Z(n31338) );
  AND U31529 ( .A(n31339), .B(n31340), .Z(n31121) );
  NANDN U31530 ( .A(n31341), .B(n31342), .Z(n31340) );
  NANDN U31531 ( .A(n31343), .B(n31344), .Z(n31342) );
  NANDN U31532 ( .A(n31344), .B(n31343), .Z(n31339) );
  ANDN U31533 ( .B(B[179]), .A(n72), .Z(n31123) );
  XNOR U31534 ( .A(n31131), .B(n31345), .Z(n31124) );
  XNOR U31535 ( .A(n31130), .B(n31128), .Z(n31345) );
  AND U31536 ( .A(n31346), .B(n31347), .Z(n31128) );
  NANDN U31537 ( .A(n31348), .B(n31349), .Z(n31347) );
  OR U31538 ( .A(n31350), .B(n31351), .Z(n31349) );
  NAND U31539 ( .A(n31351), .B(n31350), .Z(n31346) );
  ANDN U31540 ( .B(B[180]), .A(n73), .Z(n31130) );
  XNOR U31541 ( .A(n31138), .B(n31352), .Z(n31131) );
  XNOR U31542 ( .A(n31137), .B(n31135), .Z(n31352) );
  AND U31543 ( .A(n31353), .B(n31354), .Z(n31135) );
  NANDN U31544 ( .A(n31355), .B(n31356), .Z(n31354) );
  NANDN U31545 ( .A(n31357), .B(n31358), .Z(n31356) );
  NANDN U31546 ( .A(n31358), .B(n31357), .Z(n31353) );
  ANDN U31547 ( .B(B[181]), .A(n74), .Z(n31137) );
  XNOR U31548 ( .A(n31145), .B(n31359), .Z(n31138) );
  XNOR U31549 ( .A(n31144), .B(n31142), .Z(n31359) );
  AND U31550 ( .A(n31360), .B(n31361), .Z(n31142) );
  NANDN U31551 ( .A(n31362), .B(n31363), .Z(n31361) );
  OR U31552 ( .A(n31364), .B(n31365), .Z(n31363) );
  NAND U31553 ( .A(n31365), .B(n31364), .Z(n31360) );
  ANDN U31554 ( .B(B[182]), .A(n75), .Z(n31144) );
  XNOR U31555 ( .A(n31152), .B(n31366), .Z(n31145) );
  XNOR U31556 ( .A(n31151), .B(n31149), .Z(n31366) );
  AND U31557 ( .A(n31367), .B(n31368), .Z(n31149) );
  NANDN U31558 ( .A(n31369), .B(n31370), .Z(n31368) );
  NANDN U31559 ( .A(n31371), .B(n31372), .Z(n31370) );
  NANDN U31560 ( .A(n31372), .B(n31371), .Z(n31367) );
  ANDN U31561 ( .B(B[183]), .A(n76), .Z(n31151) );
  XNOR U31562 ( .A(n31159), .B(n31373), .Z(n31152) );
  XNOR U31563 ( .A(n31158), .B(n31156), .Z(n31373) );
  AND U31564 ( .A(n31374), .B(n31375), .Z(n31156) );
  NANDN U31565 ( .A(n31376), .B(n31377), .Z(n31375) );
  OR U31566 ( .A(n31378), .B(n31379), .Z(n31377) );
  NAND U31567 ( .A(n31379), .B(n31378), .Z(n31374) );
  ANDN U31568 ( .B(B[184]), .A(n77), .Z(n31158) );
  XNOR U31569 ( .A(n31166), .B(n31380), .Z(n31159) );
  XNOR U31570 ( .A(n31165), .B(n31163), .Z(n31380) );
  AND U31571 ( .A(n31381), .B(n31382), .Z(n31163) );
  NANDN U31572 ( .A(n31383), .B(n31384), .Z(n31382) );
  NANDN U31573 ( .A(n31385), .B(n31386), .Z(n31384) );
  NANDN U31574 ( .A(n31386), .B(n31385), .Z(n31381) );
  ANDN U31575 ( .B(B[185]), .A(n78), .Z(n31165) );
  XNOR U31576 ( .A(n31173), .B(n31387), .Z(n31166) );
  XNOR U31577 ( .A(n31172), .B(n31170), .Z(n31387) );
  AND U31578 ( .A(n31388), .B(n31389), .Z(n31170) );
  NANDN U31579 ( .A(n31390), .B(n31391), .Z(n31389) );
  OR U31580 ( .A(n31392), .B(n31393), .Z(n31391) );
  NAND U31581 ( .A(n31393), .B(n31392), .Z(n31388) );
  ANDN U31582 ( .B(B[186]), .A(n79), .Z(n31172) );
  XNOR U31583 ( .A(n31180), .B(n31394), .Z(n31173) );
  XNOR U31584 ( .A(n31179), .B(n31177), .Z(n31394) );
  AND U31585 ( .A(n31395), .B(n31396), .Z(n31177) );
  NANDN U31586 ( .A(n31397), .B(n31398), .Z(n31396) );
  NANDN U31587 ( .A(n31399), .B(n31400), .Z(n31398) );
  NANDN U31588 ( .A(n31400), .B(n31399), .Z(n31395) );
  ANDN U31589 ( .B(B[187]), .A(n80), .Z(n31179) );
  XNOR U31590 ( .A(n31187), .B(n31401), .Z(n31180) );
  XNOR U31591 ( .A(n31186), .B(n31184), .Z(n31401) );
  AND U31592 ( .A(n31402), .B(n31403), .Z(n31184) );
  NANDN U31593 ( .A(n31404), .B(n31405), .Z(n31403) );
  OR U31594 ( .A(n31406), .B(n31407), .Z(n31405) );
  NAND U31595 ( .A(n31407), .B(n31406), .Z(n31402) );
  ANDN U31596 ( .B(B[188]), .A(n81), .Z(n31186) );
  XNOR U31597 ( .A(n31194), .B(n31408), .Z(n31187) );
  XNOR U31598 ( .A(n31193), .B(n31191), .Z(n31408) );
  AND U31599 ( .A(n31409), .B(n31410), .Z(n31191) );
  NANDN U31600 ( .A(n31411), .B(n31412), .Z(n31410) );
  NAND U31601 ( .A(n31413), .B(n31414), .Z(n31412) );
  ANDN U31602 ( .B(B[189]), .A(n82), .Z(n31193) );
  XOR U31603 ( .A(n31200), .B(n31415), .Z(n31194) );
  XNOR U31604 ( .A(n31198), .B(n31201), .Z(n31415) );
  NAND U31605 ( .A(A[2]), .B(B[190]), .Z(n31201) );
  NANDN U31606 ( .A(n31416), .B(n31417), .Z(n31198) );
  AND U31607 ( .A(A[0]), .B(B[191]), .Z(n31417) );
  XNOR U31608 ( .A(n31203), .B(n31418), .Z(n31200) );
  NAND U31609 ( .A(A[0]), .B(B[192]), .Z(n31418) );
  NAND U31610 ( .A(B[191]), .B(A[1]), .Z(n31203) );
  NAND U31611 ( .A(n31419), .B(n31420), .Z(n412) );
  NANDN U31612 ( .A(n31421), .B(n31422), .Z(n31420) );
  OR U31613 ( .A(n31423), .B(n31424), .Z(n31422) );
  NAND U31614 ( .A(n31424), .B(n31423), .Z(n31419) );
  XOR U31615 ( .A(n29164), .B(n31425), .Z(\A1[18] ) );
  XNOR U31616 ( .A(n29163), .B(n29162), .Z(n31425) );
  NAND U31617 ( .A(n31426), .B(n31427), .Z(n29162) );
  NANDN U31618 ( .A(n31428), .B(n31429), .Z(n31427) );
  OR U31619 ( .A(n31430), .B(n31431), .Z(n31429) );
  NAND U31620 ( .A(n31431), .B(n31430), .Z(n31426) );
  ANDN U31621 ( .B(B[0]), .A(n65), .Z(n29163) );
  XNOR U31622 ( .A(n29171), .B(n31432), .Z(n29164) );
  XNOR U31623 ( .A(n29170), .B(n29168), .Z(n31432) );
  AND U31624 ( .A(n31433), .B(n31434), .Z(n29168) );
  NANDN U31625 ( .A(n31435), .B(n31436), .Z(n31434) );
  NANDN U31626 ( .A(n31437), .B(n31438), .Z(n31436) );
  NANDN U31627 ( .A(n31438), .B(n31437), .Z(n31433) );
  ANDN U31628 ( .B(B[1]), .A(n66), .Z(n29170) );
  XNOR U31629 ( .A(n29178), .B(n31439), .Z(n29171) );
  XNOR U31630 ( .A(n29177), .B(n29175), .Z(n31439) );
  AND U31631 ( .A(n31440), .B(n31441), .Z(n29175) );
  NANDN U31632 ( .A(n31442), .B(n31443), .Z(n31441) );
  OR U31633 ( .A(n31444), .B(n31445), .Z(n31443) );
  NAND U31634 ( .A(n31445), .B(n31444), .Z(n31440) );
  ANDN U31635 ( .B(B[2]), .A(n67), .Z(n29177) );
  XNOR U31636 ( .A(n29185), .B(n31446), .Z(n29178) );
  XNOR U31637 ( .A(n29184), .B(n29182), .Z(n31446) );
  AND U31638 ( .A(n31447), .B(n31448), .Z(n29182) );
  NANDN U31639 ( .A(n31449), .B(n31450), .Z(n31448) );
  NANDN U31640 ( .A(n31451), .B(n31452), .Z(n31450) );
  NANDN U31641 ( .A(n31452), .B(n31451), .Z(n31447) );
  ANDN U31642 ( .B(B[3]), .A(n68), .Z(n29184) );
  XNOR U31643 ( .A(n29192), .B(n31453), .Z(n29185) );
  XNOR U31644 ( .A(n29191), .B(n29189), .Z(n31453) );
  AND U31645 ( .A(n31454), .B(n31455), .Z(n29189) );
  NANDN U31646 ( .A(n31456), .B(n31457), .Z(n31455) );
  OR U31647 ( .A(n31458), .B(n31459), .Z(n31457) );
  NAND U31648 ( .A(n31459), .B(n31458), .Z(n31454) );
  ANDN U31649 ( .B(B[4]), .A(n69), .Z(n29191) );
  XNOR U31650 ( .A(n29199), .B(n31460), .Z(n29192) );
  XNOR U31651 ( .A(n29198), .B(n29196), .Z(n31460) );
  AND U31652 ( .A(n31461), .B(n31462), .Z(n29196) );
  NANDN U31653 ( .A(n31463), .B(n31464), .Z(n31462) );
  NANDN U31654 ( .A(n31465), .B(n31466), .Z(n31464) );
  NANDN U31655 ( .A(n31466), .B(n31465), .Z(n31461) );
  ANDN U31656 ( .B(B[5]), .A(n70), .Z(n29198) );
  XNOR U31657 ( .A(n29206), .B(n31467), .Z(n29199) );
  XNOR U31658 ( .A(n29205), .B(n29203), .Z(n31467) );
  AND U31659 ( .A(n31468), .B(n31469), .Z(n29203) );
  NANDN U31660 ( .A(n31470), .B(n31471), .Z(n31469) );
  OR U31661 ( .A(n31472), .B(n31473), .Z(n31471) );
  NAND U31662 ( .A(n31473), .B(n31472), .Z(n31468) );
  ANDN U31663 ( .B(B[6]), .A(n71), .Z(n29205) );
  XNOR U31664 ( .A(n29213), .B(n31474), .Z(n29206) );
  XNOR U31665 ( .A(n29212), .B(n29210), .Z(n31474) );
  AND U31666 ( .A(n31475), .B(n31476), .Z(n29210) );
  NANDN U31667 ( .A(n31477), .B(n31478), .Z(n31476) );
  NANDN U31668 ( .A(n31479), .B(n31480), .Z(n31478) );
  NANDN U31669 ( .A(n31480), .B(n31479), .Z(n31475) );
  ANDN U31670 ( .B(B[7]), .A(n72), .Z(n29212) );
  XNOR U31671 ( .A(n29220), .B(n31481), .Z(n29213) );
  XNOR U31672 ( .A(n29219), .B(n29217), .Z(n31481) );
  AND U31673 ( .A(n31482), .B(n31483), .Z(n29217) );
  NANDN U31674 ( .A(n31484), .B(n31485), .Z(n31483) );
  OR U31675 ( .A(n31486), .B(n31487), .Z(n31485) );
  NAND U31676 ( .A(n31487), .B(n31486), .Z(n31482) );
  ANDN U31677 ( .B(B[8]), .A(n73), .Z(n29219) );
  XNOR U31678 ( .A(n29227), .B(n31488), .Z(n29220) );
  XNOR U31679 ( .A(n29226), .B(n29224), .Z(n31488) );
  AND U31680 ( .A(n31489), .B(n31490), .Z(n29224) );
  NANDN U31681 ( .A(n31491), .B(n31492), .Z(n31490) );
  NANDN U31682 ( .A(n31493), .B(n31494), .Z(n31492) );
  NANDN U31683 ( .A(n31494), .B(n31493), .Z(n31489) );
  ANDN U31684 ( .B(B[9]), .A(n74), .Z(n29226) );
  XNOR U31685 ( .A(n29234), .B(n31495), .Z(n29227) );
  XNOR U31686 ( .A(n29233), .B(n29231), .Z(n31495) );
  AND U31687 ( .A(n31496), .B(n31497), .Z(n29231) );
  NANDN U31688 ( .A(n31498), .B(n31499), .Z(n31497) );
  OR U31689 ( .A(n31500), .B(n31501), .Z(n31499) );
  NAND U31690 ( .A(n31501), .B(n31500), .Z(n31496) );
  ANDN U31691 ( .B(B[10]), .A(n75), .Z(n29233) );
  XNOR U31692 ( .A(n29241), .B(n31502), .Z(n29234) );
  XNOR U31693 ( .A(n29240), .B(n29238), .Z(n31502) );
  AND U31694 ( .A(n31503), .B(n31504), .Z(n29238) );
  NANDN U31695 ( .A(n31505), .B(n31506), .Z(n31504) );
  NANDN U31696 ( .A(n31507), .B(n31508), .Z(n31506) );
  NANDN U31697 ( .A(n31508), .B(n31507), .Z(n31503) );
  ANDN U31698 ( .B(B[11]), .A(n76), .Z(n29240) );
  XNOR U31699 ( .A(n29248), .B(n31509), .Z(n29241) );
  XNOR U31700 ( .A(n29247), .B(n29245), .Z(n31509) );
  AND U31701 ( .A(n31510), .B(n31511), .Z(n29245) );
  NANDN U31702 ( .A(n31512), .B(n31513), .Z(n31511) );
  OR U31703 ( .A(n31514), .B(n31515), .Z(n31513) );
  NAND U31704 ( .A(n31515), .B(n31514), .Z(n31510) );
  ANDN U31705 ( .B(B[12]), .A(n77), .Z(n29247) );
  XNOR U31706 ( .A(n29255), .B(n31516), .Z(n29248) );
  XNOR U31707 ( .A(n29254), .B(n29252), .Z(n31516) );
  AND U31708 ( .A(n31517), .B(n31518), .Z(n29252) );
  NANDN U31709 ( .A(n31519), .B(n31520), .Z(n31518) );
  NANDN U31710 ( .A(n31521), .B(n31522), .Z(n31520) );
  NANDN U31711 ( .A(n31522), .B(n31521), .Z(n31517) );
  ANDN U31712 ( .B(B[13]), .A(n78), .Z(n29254) );
  XNOR U31713 ( .A(n29262), .B(n31523), .Z(n29255) );
  XNOR U31714 ( .A(n29261), .B(n29259), .Z(n31523) );
  AND U31715 ( .A(n31524), .B(n31525), .Z(n29259) );
  NANDN U31716 ( .A(n31526), .B(n31527), .Z(n31525) );
  OR U31717 ( .A(n31528), .B(n31529), .Z(n31527) );
  NAND U31718 ( .A(n31529), .B(n31528), .Z(n31524) );
  ANDN U31719 ( .B(B[14]), .A(n79), .Z(n29261) );
  XNOR U31720 ( .A(n29269), .B(n31530), .Z(n29262) );
  XNOR U31721 ( .A(n29268), .B(n29266), .Z(n31530) );
  AND U31722 ( .A(n31531), .B(n31532), .Z(n29266) );
  NANDN U31723 ( .A(n31533), .B(n31534), .Z(n31532) );
  NANDN U31724 ( .A(n31535), .B(n31536), .Z(n31534) );
  NANDN U31725 ( .A(n31536), .B(n31535), .Z(n31531) );
  ANDN U31726 ( .B(B[15]), .A(n80), .Z(n29268) );
  XNOR U31727 ( .A(n29276), .B(n31537), .Z(n29269) );
  XNOR U31728 ( .A(n29275), .B(n29273), .Z(n31537) );
  AND U31729 ( .A(n31538), .B(n31539), .Z(n29273) );
  NANDN U31730 ( .A(n31540), .B(n31541), .Z(n31539) );
  OR U31731 ( .A(n31542), .B(n31543), .Z(n31541) );
  NAND U31732 ( .A(n31543), .B(n31542), .Z(n31538) );
  ANDN U31733 ( .B(B[16]), .A(n81), .Z(n29275) );
  XNOR U31734 ( .A(n29283), .B(n31544), .Z(n29276) );
  XNOR U31735 ( .A(n29282), .B(n29280), .Z(n31544) );
  AND U31736 ( .A(n31545), .B(n31546), .Z(n29280) );
  NANDN U31737 ( .A(n31547), .B(n31548), .Z(n31546) );
  NAND U31738 ( .A(n31549), .B(n31550), .Z(n31548) );
  ANDN U31739 ( .B(B[17]), .A(n82), .Z(n29282) );
  XOR U31740 ( .A(n29289), .B(n31551), .Z(n29283) );
  XNOR U31741 ( .A(n29287), .B(n29290), .Z(n31551) );
  NAND U31742 ( .A(A[2]), .B(B[18]), .Z(n29290) );
  NANDN U31743 ( .A(n31552), .B(n31553), .Z(n29287) );
  AND U31744 ( .A(A[0]), .B(B[19]), .Z(n31553) );
  XNOR U31745 ( .A(n29292), .B(n31554), .Z(n29289) );
  NAND U31746 ( .A(A[0]), .B(B[20]), .Z(n31554) );
  NAND U31747 ( .A(B[19]), .B(A[1]), .Z(n29292) );
  XOR U31748 ( .A(n414), .B(n413), .Z(\A1[189] ) );
  XOR U31749 ( .A(n31424), .B(n31555), .Z(n413) );
  XNOR U31750 ( .A(n31423), .B(n31421), .Z(n31555) );
  AND U31751 ( .A(n31556), .B(n31557), .Z(n31421) );
  NANDN U31752 ( .A(n31558), .B(n31559), .Z(n31557) );
  NANDN U31753 ( .A(n31560), .B(n31561), .Z(n31559) );
  NANDN U31754 ( .A(n31561), .B(n31560), .Z(n31556) );
  ANDN U31755 ( .B(B[160]), .A(n54), .Z(n31423) );
  XNOR U31756 ( .A(n31218), .B(n31562), .Z(n31424) );
  XNOR U31757 ( .A(n31217), .B(n31215), .Z(n31562) );
  AND U31758 ( .A(n31563), .B(n31564), .Z(n31215) );
  NANDN U31759 ( .A(n31565), .B(n31566), .Z(n31564) );
  OR U31760 ( .A(n31567), .B(n31568), .Z(n31566) );
  NAND U31761 ( .A(n31568), .B(n31567), .Z(n31563) );
  ANDN U31762 ( .B(B[161]), .A(n55), .Z(n31217) );
  XNOR U31763 ( .A(n31225), .B(n31569), .Z(n31218) );
  XNOR U31764 ( .A(n31224), .B(n31222), .Z(n31569) );
  AND U31765 ( .A(n31570), .B(n31571), .Z(n31222) );
  NANDN U31766 ( .A(n31572), .B(n31573), .Z(n31571) );
  NANDN U31767 ( .A(n31574), .B(n31575), .Z(n31573) );
  NANDN U31768 ( .A(n31575), .B(n31574), .Z(n31570) );
  ANDN U31769 ( .B(B[162]), .A(n56), .Z(n31224) );
  XNOR U31770 ( .A(n31232), .B(n31576), .Z(n31225) );
  XNOR U31771 ( .A(n31231), .B(n31229), .Z(n31576) );
  AND U31772 ( .A(n31577), .B(n31578), .Z(n31229) );
  NANDN U31773 ( .A(n31579), .B(n31580), .Z(n31578) );
  OR U31774 ( .A(n31581), .B(n31582), .Z(n31580) );
  NAND U31775 ( .A(n31582), .B(n31581), .Z(n31577) );
  ANDN U31776 ( .B(B[163]), .A(n57), .Z(n31231) );
  XNOR U31777 ( .A(n31239), .B(n31583), .Z(n31232) );
  XNOR U31778 ( .A(n31238), .B(n31236), .Z(n31583) );
  AND U31779 ( .A(n31584), .B(n31585), .Z(n31236) );
  NANDN U31780 ( .A(n31586), .B(n31587), .Z(n31585) );
  NANDN U31781 ( .A(n31588), .B(n31589), .Z(n31587) );
  NANDN U31782 ( .A(n31589), .B(n31588), .Z(n31584) );
  ANDN U31783 ( .B(B[164]), .A(n58), .Z(n31238) );
  XNOR U31784 ( .A(n31246), .B(n31590), .Z(n31239) );
  XNOR U31785 ( .A(n31245), .B(n31243), .Z(n31590) );
  AND U31786 ( .A(n31591), .B(n31592), .Z(n31243) );
  NANDN U31787 ( .A(n31593), .B(n31594), .Z(n31592) );
  OR U31788 ( .A(n31595), .B(n31596), .Z(n31594) );
  NAND U31789 ( .A(n31596), .B(n31595), .Z(n31591) );
  ANDN U31790 ( .B(B[165]), .A(n59), .Z(n31245) );
  XNOR U31791 ( .A(n31253), .B(n31597), .Z(n31246) );
  XNOR U31792 ( .A(n31252), .B(n31250), .Z(n31597) );
  AND U31793 ( .A(n31598), .B(n31599), .Z(n31250) );
  NANDN U31794 ( .A(n31600), .B(n31601), .Z(n31599) );
  NANDN U31795 ( .A(n31602), .B(n31603), .Z(n31601) );
  NANDN U31796 ( .A(n31603), .B(n31602), .Z(n31598) );
  ANDN U31797 ( .B(B[166]), .A(n60), .Z(n31252) );
  XNOR U31798 ( .A(n31260), .B(n31604), .Z(n31253) );
  XNOR U31799 ( .A(n31259), .B(n31257), .Z(n31604) );
  AND U31800 ( .A(n31605), .B(n31606), .Z(n31257) );
  NANDN U31801 ( .A(n31607), .B(n31608), .Z(n31606) );
  OR U31802 ( .A(n31609), .B(n31610), .Z(n31608) );
  NAND U31803 ( .A(n31610), .B(n31609), .Z(n31605) );
  ANDN U31804 ( .B(B[167]), .A(n61), .Z(n31259) );
  XNOR U31805 ( .A(n31267), .B(n31611), .Z(n31260) );
  XNOR U31806 ( .A(n31266), .B(n31264), .Z(n31611) );
  AND U31807 ( .A(n31612), .B(n31613), .Z(n31264) );
  NANDN U31808 ( .A(n31614), .B(n31615), .Z(n31613) );
  NANDN U31809 ( .A(n31616), .B(n31617), .Z(n31615) );
  NANDN U31810 ( .A(n31617), .B(n31616), .Z(n31612) );
  ANDN U31811 ( .B(B[168]), .A(n62), .Z(n31266) );
  XNOR U31812 ( .A(n31274), .B(n31618), .Z(n31267) );
  XNOR U31813 ( .A(n31273), .B(n31271), .Z(n31618) );
  AND U31814 ( .A(n31619), .B(n31620), .Z(n31271) );
  NANDN U31815 ( .A(n31621), .B(n31622), .Z(n31620) );
  OR U31816 ( .A(n31623), .B(n31624), .Z(n31622) );
  NAND U31817 ( .A(n31624), .B(n31623), .Z(n31619) );
  ANDN U31818 ( .B(B[169]), .A(n63), .Z(n31273) );
  XNOR U31819 ( .A(n31281), .B(n31625), .Z(n31274) );
  XNOR U31820 ( .A(n31280), .B(n31278), .Z(n31625) );
  AND U31821 ( .A(n31626), .B(n31627), .Z(n31278) );
  NANDN U31822 ( .A(n31628), .B(n31629), .Z(n31627) );
  NANDN U31823 ( .A(n31630), .B(n31631), .Z(n31629) );
  NANDN U31824 ( .A(n31631), .B(n31630), .Z(n31626) );
  ANDN U31825 ( .B(B[170]), .A(n64), .Z(n31280) );
  XNOR U31826 ( .A(n31288), .B(n31632), .Z(n31281) );
  XNOR U31827 ( .A(n31287), .B(n31285), .Z(n31632) );
  AND U31828 ( .A(n31633), .B(n31634), .Z(n31285) );
  NANDN U31829 ( .A(n31635), .B(n31636), .Z(n31634) );
  OR U31830 ( .A(n31637), .B(n31638), .Z(n31636) );
  NAND U31831 ( .A(n31638), .B(n31637), .Z(n31633) );
  ANDN U31832 ( .B(B[171]), .A(n65), .Z(n31287) );
  XNOR U31833 ( .A(n31295), .B(n31639), .Z(n31288) );
  XNOR U31834 ( .A(n31294), .B(n31292), .Z(n31639) );
  AND U31835 ( .A(n31640), .B(n31641), .Z(n31292) );
  NANDN U31836 ( .A(n31642), .B(n31643), .Z(n31641) );
  NANDN U31837 ( .A(n31644), .B(n31645), .Z(n31643) );
  NANDN U31838 ( .A(n31645), .B(n31644), .Z(n31640) );
  ANDN U31839 ( .B(B[172]), .A(n66), .Z(n31294) );
  XNOR U31840 ( .A(n31302), .B(n31646), .Z(n31295) );
  XNOR U31841 ( .A(n31301), .B(n31299), .Z(n31646) );
  AND U31842 ( .A(n31647), .B(n31648), .Z(n31299) );
  NANDN U31843 ( .A(n31649), .B(n31650), .Z(n31648) );
  OR U31844 ( .A(n31651), .B(n31652), .Z(n31650) );
  NAND U31845 ( .A(n31652), .B(n31651), .Z(n31647) );
  ANDN U31846 ( .B(B[173]), .A(n67), .Z(n31301) );
  XNOR U31847 ( .A(n31309), .B(n31653), .Z(n31302) );
  XNOR U31848 ( .A(n31308), .B(n31306), .Z(n31653) );
  AND U31849 ( .A(n31654), .B(n31655), .Z(n31306) );
  NANDN U31850 ( .A(n31656), .B(n31657), .Z(n31655) );
  NANDN U31851 ( .A(n31658), .B(n31659), .Z(n31657) );
  NANDN U31852 ( .A(n31659), .B(n31658), .Z(n31654) );
  ANDN U31853 ( .B(B[174]), .A(n68), .Z(n31308) );
  XNOR U31854 ( .A(n31316), .B(n31660), .Z(n31309) );
  XNOR U31855 ( .A(n31315), .B(n31313), .Z(n31660) );
  AND U31856 ( .A(n31661), .B(n31662), .Z(n31313) );
  NANDN U31857 ( .A(n31663), .B(n31664), .Z(n31662) );
  OR U31858 ( .A(n31665), .B(n31666), .Z(n31664) );
  NAND U31859 ( .A(n31666), .B(n31665), .Z(n31661) );
  ANDN U31860 ( .B(B[175]), .A(n69), .Z(n31315) );
  XNOR U31861 ( .A(n31323), .B(n31667), .Z(n31316) );
  XNOR U31862 ( .A(n31322), .B(n31320), .Z(n31667) );
  AND U31863 ( .A(n31668), .B(n31669), .Z(n31320) );
  NANDN U31864 ( .A(n31670), .B(n31671), .Z(n31669) );
  NANDN U31865 ( .A(n31672), .B(n31673), .Z(n31671) );
  NANDN U31866 ( .A(n31673), .B(n31672), .Z(n31668) );
  ANDN U31867 ( .B(B[176]), .A(n70), .Z(n31322) );
  XNOR U31868 ( .A(n31330), .B(n31674), .Z(n31323) );
  XNOR U31869 ( .A(n31329), .B(n31327), .Z(n31674) );
  AND U31870 ( .A(n31675), .B(n31676), .Z(n31327) );
  NANDN U31871 ( .A(n31677), .B(n31678), .Z(n31676) );
  OR U31872 ( .A(n31679), .B(n31680), .Z(n31678) );
  NAND U31873 ( .A(n31680), .B(n31679), .Z(n31675) );
  ANDN U31874 ( .B(B[177]), .A(n71), .Z(n31329) );
  XNOR U31875 ( .A(n31337), .B(n31681), .Z(n31330) );
  XNOR U31876 ( .A(n31336), .B(n31334), .Z(n31681) );
  AND U31877 ( .A(n31682), .B(n31683), .Z(n31334) );
  NANDN U31878 ( .A(n31684), .B(n31685), .Z(n31683) );
  NANDN U31879 ( .A(n31686), .B(n31687), .Z(n31685) );
  NANDN U31880 ( .A(n31687), .B(n31686), .Z(n31682) );
  ANDN U31881 ( .B(B[178]), .A(n72), .Z(n31336) );
  XNOR U31882 ( .A(n31344), .B(n31688), .Z(n31337) );
  XNOR U31883 ( .A(n31343), .B(n31341), .Z(n31688) );
  AND U31884 ( .A(n31689), .B(n31690), .Z(n31341) );
  NANDN U31885 ( .A(n31691), .B(n31692), .Z(n31690) );
  OR U31886 ( .A(n31693), .B(n31694), .Z(n31692) );
  NAND U31887 ( .A(n31694), .B(n31693), .Z(n31689) );
  ANDN U31888 ( .B(B[179]), .A(n73), .Z(n31343) );
  XNOR U31889 ( .A(n31351), .B(n31695), .Z(n31344) );
  XNOR U31890 ( .A(n31350), .B(n31348), .Z(n31695) );
  AND U31891 ( .A(n31696), .B(n31697), .Z(n31348) );
  NANDN U31892 ( .A(n31698), .B(n31699), .Z(n31697) );
  NANDN U31893 ( .A(n31700), .B(n31701), .Z(n31699) );
  NANDN U31894 ( .A(n31701), .B(n31700), .Z(n31696) );
  ANDN U31895 ( .B(B[180]), .A(n74), .Z(n31350) );
  XNOR U31896 ( .A(n31358), .B(n31702), .Z(n31351) );
  XNOR U31897 ( .A(n31357), .B(n31355), .Z(n31702) );
  AND U31898 ( .A(n31703), .B(n31704), .Z(n31355) );
  NANDN U31899 ( .A(n31705), .B(n31706), .Z(n31704) );
  OR U31900 ( .A(n31707), .B(n31708), .Z(n31706) );
  NAND U31901 ( .A(n31708), .B(n31707), .Z(n31703) );
  ANDN U31902 ( .B(B[181]), .A(n75), .Z(n31357) );
  XNOR U31903 ( .A(n31365), .B(n31709), .Z(n31358) );
  XNOR U31904 ( .A(n31364), .B(n31362), .Z(n31709) );
  AND U31905 ( .A(n31710), .B(n31711), .Z(n31362) );
  NANDN U31906 ( .A(n31712), .B(n31713), .Z(n31711) );
  NANDN U31907 ( .A(n31714), .B(n31715), .Z(n31713) );
  NANDN U31908 ( .A(n31715), .B(n31714), .Z(n31710) );
  ANDN U31909 ( .B(B[182]), .A(n76), .Z(n31364) );
  XNOR U31910 ( .A(n31372), .B(n31716), .Z(n31365) );
  XNOR U31911 ( .A(n31371), .B(n31369), .Z(n31716) );
  AND U31912 ( .A(n31717), .B(n31718), .Z(n31369) );
  NANDN U31913 ( .A(n31719), .B(n31720), .Z(n31718) );
  OR U31914 ( .A(n31721), .B(n31722), .Z(n31720) );
  NAND U31915 ( .A(n31722), .B(n31721), .Z(n31717) );
  ANDN U31916 ( .B(B[183]), .A(n77), .Z(n31371) );
  XNOR U31917 ( .A(n31379), .B(n31723), .Z(n31372) );
  XNOR U31918 ( .A(n31378), .B(n31376), .Z(n31723) );
  AND U31919 ( .A(n31724), .B(n31725), .Z(n31376) );
  NANDN U31920 ( .A(n31726), .B(n31727), .Z(n31725) );
  NANDN U31921 ( .A(n31728), .B(n31729), .Z(n31727) );
  NANDN U31922 ( .A(n31729), .B(n31728), .Z(n31724) );
  ANDN U31923 ( .B(B[184]), .A(n78), .Z(n31378) );
  XNOR U31924 ( .A(n31386), .B(n31730), .Z(n31379) );
  XNOR U31925 ( .A(n31385), .B(n31383), .Z(n31730) );
  AND U31926 ( .A(n31731), .B(n31732), .Z(n31383) );
  NANDN U31927 ( .A(n31733), .B(n31734), .Z(n31732) );
  OR U31928 ( .A(n31735), .B(n31736), .Z(n31734) );
  NAND U31929 ( .A(n31736), .B(n31735), .Z(n31731) );
  ANDN U31930 ( .B(B[185]), .A(n79), .Z(n31385) );
  XNOR U31931 ( .A(n31393), .B(n31737), .Z(n31386) );
  XNOR U31932 ( .A(n31392), .B(n31390), .Z(n31737) );
  AND U31933 ( .A(n31738), .B(n31739), .Z(n31390) );
  NANDN U31934 ( .A(n31740), .B(n31741), .Z(n31739) );
  NANDN U31935 ( .A(n31742), .B(n31743), .Z(n31741) );
  NANDN U31936 ( .A(n31743), .B(n31742), .Z(n31738) );
  ANDN U31937 ( .B(B[186]), .A(n80), .Z(n31392) );
  XNOR U31938 ( .A(n31400), .B(n31744), .Z(n31393) );
  XNOR U31939 ( .A(n31399), .B(n31397), .Z(n31744) );
  AND U31940 ( .A(n31745), .B(n31746), .Z(n31397) );
  NANDN U31941 ( .A(n31747), .B(n31748), .Z(n31746) );
  OR U31942 ( .A(n31749), .B(n31750), .Z(n31748) );
  NAND U31943 ( .A(n31750), .B(n31749), .Z(n31745) );
  ANDN U31944 ( .B(B[187]), .A(n81), .Z(n31399) );
  XNOR U31945 ( .A(n31407), .B(n31751), .Z(n31400) );
  XNOR U31946 ( .A(n31406), .B(n31404), .Z(n31751) );
  AND U31947 ( .A(n31752), .B(n31753), .Z(n31404) );
  NANDN U31948 ( .A(n31754), .B(n31755), .Z(n31753) );
  NAND U31949 ( .A(n31756), .B(n31757), .Z(n31755) );
  ANDN U31950 ( .B(B[188]), .A(n82), .Z(n31406) );
  XOR U31951 ( .A(n31413), .B(n31758), .Z(n31407) );
  XNOR U31952 ( .A(n31411), .B(n31414), .Z(n31758) );
  NAND U31953 ( .A(A[2]), .B(B[189]), .Z(n31414) );
  NANDN U31954 ( .A(n31759), .B(n31760), .Z(n31411) );
  AND U31955 ( .A(A[0]), .B(B[190]), .Z(n31760) );
  XNOR U31956 ( .A(n31416), .B(n31761), .Z(n31413) );
  NAND U31957 ( .A(A[0]), .B(B[191]), .Z(n31761) );
  NAND U31958 ( .A(B[190]), .B(A[1]), .Z(n31416) );
  NAND U31959 ( .A(n31762), .B(n31763), .Z(n414) );
  NANDN U31960 ( .A(n31764), .B(n31765), .Z(n31763) );
  OR U31961 ( .A(n31766), .B(n31767), .Z(n31765) );
  NAND U31962 ( .A(n31767), .B(n31766), .Z(n31762) );
  XOR U31963 ( .A(n416), .B(n415), .Z(\A1[188] ) );
  XOR U31964 ( .A(n31767), .B(n31768), .Z(n415) );
  XNOR U31965 ( .A(n31766), .B(n31764), .Z(n31768) );
  AND U31966 ( .A(n31769), .B(n31770), .Z(n31764) );
  NANDN U31967 ( .A(n31771), .B(n31772), .Z(n31770) );
  NANDN U31968 ( .A(n31773), .B(n31774), .Z(n31772) );
  NANDN U31969 ( .A(n31774), .B(n31773), .Z(n31769) );
  ANDN U31970 ( .B(B[159]), .A(n54), .Z(n31766) );
  XNOR U31971 ( .A(n31561), .B(n31775), .Z(n31767) );
  XNOR U31972 ( .A(n31560), .B(n31558), .Z(n31775) );
  AND U31973 ( .A(n31776), .B(n31777), .Z(n31558) );
  NANDN U31974 ( .A(n31778), .B(n31779), .Z(n31777) );
  OR U31975 ( .A(n31780), .B(n31781), .Z(n31779) );
  NAND U31976 ( .A(n31781), .B(n31780), .Z(n31776) );
  ANDN U31977 ( .B(B[160]), .A(n55), .Z(n31560) );
  XNOR U31978 ( .A(n31568), .B(n31782), .Z(n31561) );
  XNOR U31979 ( .A(n31567), .B(n31565), .Z(n31782) );
  AND U31980 ( .A(n31783), .B(n31784), .Z(n31565) );
  NANDN U31981 ( .A(n31785), .B(n31786), .Z(n31784) );
  NANDN U31982 ( .A(n31787), .B(n31788), .Z(n31786) );
  NANDN U31983 ( .A(n31788), .B(n31787), .Z(n31783) );
  ANDN U31984 ( .B(B[161]), .A(n56), .Z(n31567) );
  XNOR U31985 ( .A(n31575), .B(n31789), .Z(n31568) );
  XNOR U31986 ( .A(n31574), .B(n31572), .Z(n31789) );
  AND U31987 ( .A(n31790), .B(n31791), .Z(n31572) );
  NANDN U31988 ( .A(n31792), .B(n31793), .Z(n31791) );
  OR U31989 ( .A(n31794), .B(n31795), .Z(n31793) );
  NAND U31990 ( .A(n31795), .B(n31794), .Z(n31790) );
  ANDN U31991 ( .B(B[162]), .A(n57), .Z(n31574) );
  XNOR U31992 ( .A(n31582), .B(n31796), .Z(n31575) );
  XNOR U31993 ( .A(n31581), .B(n31579), .Z(n31796) );
  AND U31994 ( .A(n31797), .B(n31798), .Z(n31579) );
  NANDN U31995 ( .A(n31799), .B(n31800), .Z(n31798) );
  NANDN U31996 ( .A(n31801), .B(n31802), .Z(n31800) );
  NANDN U31997 ( .A(n31802), .B(n31801), .Z(n31797) );
  ANDN U31998 ( .B(B[163]), .A(n58), .Z(n31581) );
  XNOR U31999 ( .A(n31589), .B(n31803), .Z(n31582) );
  XNOR U32000 ( .A(n31588), .B(n31586), .Z(n31803) );
  AND U32001 ( .A(n31804), .B(n31805), .Z(n31586) );
  NANDN U32002 ( .A(n31806), .B(n31807), .Z(n31805) );
  OR U32003 ( .A(n31808), .B(n31809), .Z(n31807) );
  NAND U32004 ( .A(n31809), .B(n31808), .Z(n31804) );
  ANDN U32005 ( .B(B[164]), .A(n59), .Z(n31588) );
  XNOR U32006 ( .A(n31596), .B(n31810), .Z(n31589) );
  XNOR U32007 ( .A(n31595), .B(n31593), .Z(n31810) );
  AND U32008 ( .A(n31811), .B(n31812), .Z(n31593) );
  NANDN U32009 ( .A(n31813), .B(n31814), .Z(n31812) );
  NANDN U32010 ( .A(n31815), .B(n31816), .Z(n31814) );
  NANDN U32011 ( .A(n31816), .B(n31815), .Z(n31811) );
  ANDN U32012 ( .B(B[165]), .A(n60), .Z(n31595) );
  XNOR U32013 ( .A(n31603), .B(n31817), .Z(n31596) );
  XNOR U32014 ( .A(n31602), .B(n31600), .Z(n31817) );
  AND U32015 ( .A(n31818), .B(n31819), .Z(n31600) );
  NANDN U32016 ( .A(n31820), .B(n31821), .Z(n31819) );
  OR U32017 ( .A(n31822), .B(n31823), .Z(n31821) );
  NAND U32018 ( .A(n31823), .B(n31822), .Z(n31818) );
  ANDN U32019 ( .B(B[166]), .A(n61), .Z(n31602) );
  XNOR U32020 ( .A(n31610), .B(n31824), .Z(n31603) );
  XNOR U32021 ( .A(n31609), .B(n31607), .Z(n31824) );
  AND U32022 ( .A(n31825), .B(n31826), .Z(n31607) );
  NANDN U32023 ( .A(n31827), .B(n31828), .Z(n31826) );
  NANDN U32024 ( .A(n31829), .B(n31830), .Z(n31828) );
  NANDN U32025 ( .A(n31830), .B(n31829), .Z(n31825) );
  ANDN U32026 ( .B(B[167]), .A(n62), .Z(n31609) );
  XNOR U32027 ( .A(n31617), .B(n31831), .Z(n31610) );
  XNOR U32028 ( .A(n31616), .B(n31614), .Z(n31831) );
  AND U32029 ( .A(n31832), .B(n31833), .Z(n31614) );
  NANDN U32030 ( .A(n31834), .B(n31835), .Z(n31833) );
  OR U32031 ( .A(n31836), .B(n31837), .Z(n31835) );
  NAND U32032 ( .A(n31837), .B(n31836), .Z(n31832) );
  ANDN U32033 ( .B(B[168]), .A(n63), .Z(n31616) );
  XNOR U32034 ( .A(n31624), .B(n31838), .Z(n31617) );
  XNOR U32035 ( .A(n31623), .B(n31621), .Z(n31838) );
  AND U32036 ( .A(n31839), .B(n31840), .Z(n31621) );
  NANDN U32037 ( .A(n31841), .B(n31842), .Z(n31840) );
  NANDN U32038 ( .A(n31843), .B(n31844), .Z(n31842) );
  NANDN U32039 ( .A(n31844), .B(n31843), .Z(n31839) );
  ANDN U32040 ( .B(B[169]), .A(n64), .Z(n31623) );
  XNOR U32041 ( .A(n31631), .B(n31845), .Z(n31624) );
  XNOR U32042 ( .A(n31630), .B(n31628), .Z(n31845) );
  AND U32043 ( .A(n31846), .B(n31847), .Z(n31628) );
  NANDN U32044 ( .A(n31848), .B(n31849), .Z(n31847) );
  OR U32045 ( .A(n31850), .B(n31851), .Z(n31849) );
  NAND U32046 ( .A(n31851), .B(n31850), .Z(n31846) );
  ANDN U32047 ( .B(B[170]), .A(n65), .Z(n31630) );
  XNOR U32048 ( .A(n31638), .B(n31852), .Z(n31631) );
  XNOR U32049 ( .A(n31637), .B(n31635), .Z(n31852) );
  AND U32050 ( .A(n31853), .B(n31854), .Z(n31635) );
  NANDN U32051 ( .A(n31855), .B(n31856), .Z(n31854) );
  NANDN U32052 ( .A(n31857), .B(n31858), .Z(n31856) );
  NANDN U32053 ( .A(n31858), .B(n31857), .Z(n31853) );
  ANDN U32054 ( .B(B[171]), .A(n66), .Z(n31637) );
  XNOR U32055 ( .A(n31645), .B(n31859), .Z(n31638) );
  XNOR U32056 ( .A(n31644), .B(n31642), .Z(n31859) );
  AND U32057 ( .A(n31860), .B(n31861), .Z(n31642) );
  NANDN U32058 ( .A(n31862), .B(n31863), .Z(n31861) );
  OR U32059 ( .A(n31864), .B(n31865), .Z(n31863) );
  NAND U32060 ( .A(n31865), .B(n31864), .Z(n31860) );
  ANDN U32061 ( .B(B[172]), .A(n67), .Z(n31644) );
  XNOR U32062 ( .A(n31652), .B(n31866), .Z(n31645) );
  XNOR U32063 ( .A(n31651), .B(n31649), .Z(n31866) );
  AND U32064 ( .A(n31867), .B(n31868), .Z(n31649) );
  NANDN U32065 ( .A(n31869), .B(n31870), .Z(n31868) );
  NANDN U32066 ( .A(n31871), .B(n31872), .Z(n31870) );
  NANDN U32067 ( .A(n31872), .B(n31871), .Z(n31867) );
  ANDN U32068 ( .B(B[173]), .A(n68), .Z(n31651) );
  XNOR U32069 ( .A(n31659), .B(n31873), .Z(n31652) );
  XNOR U32070 ( .A(n31658), .B(n31656), .Z(n31873) );
  AND U32071 ( .A(n31874), .B(n31875), .Z(n31656) );
  NANDN U32072 ( .A(n31876), .B(n31877), .Z(n31875) );
  OR U32073 ( .A(n31878), .B(n31879), .Z(n31877) );
  NAND U32074 ( .A(n31879), .B(n31878), .Z(n31874) );
  ANDN U32075 ( .B(B[174]), .A(n69), .Z(n31658) );
  XNOR U32076 ( .A(n31666), .B(n31880), .Z(n31659) );
  XNOR U32077 ( .A(n31665), .B(n31663), .Z(n31880) );
  AND U32078 ( .A(n31881), .B(n31882), .Z(n31663) );
  NANDN U32079 ( .A(n31883), .B(n31884), .Z(n31882) );
  NANDN U32080 ( .A(n31885), .B(n31886), .Z(n31884) );
  NANDN U32081 ( .A(n31886), .B(n31885), .Z(n31881) );
  ANDN U32082 ( .B(B[175]), .A(n70), .Z(n31665) );
  XNOR U32083 ( .A(n31673), .B(n31887), .Z(n31666) );
  XNOR U32084 ( .A(n31672), .B(n31670), .Z(n31887) );
  AND U32085 ( .A(n31888), .B(n31889), .Z(n31670) );
  NANDN U32086 ( .A(n31890), .B(n31891), .Z(n31889) );
  OR U32087 ( .A(n31892), .B(n31893), .Z(n31891) );
  NAND U32088 ( .A(n31893), .B(n31892), .Z(n31888) );
  ANDN U32089 ( .B(B[176]), .A(n71), .Z(n31672) );
  XNOR U32090 ( .A(n31680), .B(n31894), .Z(n31673) );
  XNOR U32091 ( .A(n31679), .B(n31677), .Z(n31894) );
  AND U32092 ( .A(n31895), .B(n31896), .Z(n31677) );
  NANDN U32093 ( .A(n31897), .B(n31898), .Z(n31896) );
  NANDN U32094 ( .A(n31899), .B(n31900), .Z(n31898) );
  NANDN U32095 ( .A(n31900), .B(n31899), .Z(n31895) );
  ANDN U32096 ( .B(B[177]), .A(n72), .Z(n31679) );
  XNOR U32097 ( .A(n31687), .B(n31901), .Z(n31680) );
  XNOR U32098 ( .A(n31686), .B(n31684), .Z(n31901) );
  AND U32099 ( .A(n31902), .B(n31903), .Z(n31684) );
  NANDN U32100 ( .A(n31904), .B(n31905), .Z(n31903) );
  OR U32101 ( .A(n31906), .B(n31907), .Z(n31905) );
  NAND U32102 ( .A(n31907), .B(n31906), .Z(n31902) );
  ANDN U32103 ( .B(B[178]), .A(n73), .Z(n31686) );
  XNOR U32104 ( .A(n31694), .B(n31908), .Z(n31687) );
  XNOR U32105 ( .A(n31693), .B(n31691), .Z(n31908) );
  AND U32106 ( .A(n31909), .B(n31910), .Z(n31691) );
  NANDN U32107 ( .A(n31911), .B(n31912), .Z(n31910) );
  NANDN U32108 ( .A(n31913), .B(n31914), .Z(n31912) );
  NANDN U32109 ( .A(n31914), .B(n31913), .Z(n31909) );
  ANDN U32110 ( .B(B[179]), .A(n74), .Z(n31693) );
  XNOR U32111 ( .A(n31701), .B(n31915), .Z(n31694) );
  XNOR U32112 ( .A(n31700), .B(n31698), .Z(n31915) );
  AND U32113 ( .A(n31916), .B(n31917), .Z(n31698) );
  NANDN U32114 ( .A(n31918), .B(n31919), .Z(n31917) );
  OR U32115 ( .A(n31920), .B(n31921), .Z(n31919) );
  NAND U32116 ( .A(n31921), .B(n31920), .Z(n31916) );
  ANDN U32117 ( .B(B[180]), .A(n75), .Z(n31700) );
  XNOR U32118 ( .A(n31708), .B(n31922), .Z(n31701) );
  XNOR U32119 ( .A(n31707), .B(n31705), .Z(n31922) );
  AND U32120 ( .A(n31923), .B(n31924), .Z(n31705) );
  NANDN U32121 ( .A(n31925), .B(n31926), .Z(n31924) );
  NANDN U32122 ( .A(n31927), .B(n31928), .Z(n31926) );
  NANDN U32123 ( .A(n31928), .B(n31927), .Z(n31923) );
  ANDN U32124 ( .B(B[181]), .A(n76), .Z(n31707) );
  XNOR U32125 ( .A(n31715), .B(n31929), .Z(n31708) );
  XNOR U32126 ( .A(n31714), .B(n31712), .Z(n31929) );
  AND U32127 ( .A(n31930), .B(n31931), .Z(n31712) );
  NANDN U32128 ( .A(n31932), .B(n31933), .Z(n31931) );
  OR U32129 ( .A(n31934), .B(n31935), .Z(n31933) );
  NAND U32130 ( .A(n31935), .B(n31934), .Z(n31930) );
  ANDN U32131 ( .B(B[182]), .A(n77), .Z(n31714) );
  XNOR U32132 ( .A(n31722), .B(n31936), .Z(n31715) );
  XNOR U32133 ( .A(n31721), .B(n31719), .Z(n31936) );
  AND U32134 ( .A(n31937), .B(n31938), .Z(n31719) );
  NANDN U32135 ( .A(n31939), .B(n31940), .Z(n31938) );
  NANDN U32136 ( .A(n31941), .B(n31942), .Z(n31940) );
  NANDN U32137 ( .A(n31942), .B(n31941), .Z(n31937) );
  ANDN U32138 ( .B(B[183]), .A(n78), .Z(n31721) );
  XNOR U32139 ( .A(n31729), .B(n31943), .Z(n31722) );
  XNOR U32140 ( .A(n31728), .B(n31726), .Z(n31943) );
  AND U32141 ( .A(n31944), .B(n31945), .Z(n31726) );
  NANDN U32142 ( .A(n31946), .B(n31947), .Z(n31945) );
  OR U32143 ( .A(n31948), .B(n31949), .Z(n31947) );
  NAND U32144 ( .A(n31949), .B(n31948), .Z(n31944) );
  ANDN U32145 ( .B(B[184]), .A(n79), .Z(n31728) );
  XNOR U32146 ( .A(n31736), .B(n31950), .Z(n31729) );
  XNOR U32147 ( .A(n31735), .B(n31733), .Z(n31950) );
  AND U32148 ( .A(n31951), .B(n31952), .Z(n31733) );
  NANDN U32149 ( .A(n31953), .B(n31954), .Z(n31952) );
  NANDN U32150 ( .A(n31955), .B(n31956), .Z(n31954) );
  NANDN U32151 ( .A(n31956), .B(n31955), .Z(n31951) );
  ANDN U32152 ( .B(B[185]), .A(n80), .Z(n31735) );
  XNOR U32153 ( .A(n31743), .B(n31957), .Z(n31736) );
  XNOR U32154 ( .A(n31742), .B(n31740), .Z(n31957) );
  AND U32155 ( .A(n31958), .B(n31959), .Z(n31740) );
  NANDN U32156 ( .A(n31960), .B(n31961), .Z(n31959) );
  OR U32157 ( .A(n31962), .B(n31963), .Z(n31961) );
  NAND U32158 ( .A(n31963), .B(n31962), .Z(n31958) );
  ANDN U32159 ( .B(B[186]), .A(n81), .Z(n31742) );
  XNOR U32160 ( .A(n31750), .B(n31964), .Z(n31743) );
  XNOR U32161 ( .A(n31749), .B(n31747), .Z(n31964) );
  AND U32162 ( .A(n31965), .B(n31966), .Z(n31747) );
  NANDN U32163 ( .A(n31967), .B(n31968), .Z(n31966) );
  NAND U32164 ( .A(n31969), .B(n31970), .Z(n31968) );
  ANDN U32165 ( .B(B[187]), .A(n82), .Z(n31749) );
  XOR U32166 ( .A(n31756), .B(n31971), .Z(n31750) );
  XNOR U32167 ( .A(n31754), .B(n31757), .Z(n31971) );
  NAND U32168 ( .A(A[2]), .B(B[188]), .Z(n31757) );
  NANDN U32169 ( .A(n31972), .B(n31973), .Z(n31754) );
  AND U32170 ( .A(A[0]), .B(B[189]), .Z(n31973) );
  XNOR U32171 ( .A(n31759), .B(n31974), .Z(n31756) );
  NAND U32172 ( .A(A[0]), .B(B[190]), .Z(n31974) );
  NAND U32173 ( .A(B[189]), .B(A[1]), .Z(n31759) );
  NAND U32174 ( .A(n31975), .B(n31976), .Z(n416) );
  NANDN U32175 ( .A(n31977), .B(n31978), .Z(n31976) );
  OR U32176 ( .A(n31979), .B(n31980), .Z(n31978) );
  NAND U32177 ( .A(n31980), .B(n31979), .Z(n31975) );
  XOR U32178 ( .A(n418), .B(n417), .Z(\A1[187] ) );
  XOR U32179 ( .A(n31980), .B(n31981), .Z(n417) );
  XNOR U32180 ( .A(n31979), .B(n31977), .Z(n31981) );
  AND U32181 ( .A(n31982), .B(n31983), .Z(n31977) );
  NANDN U32182 ( .A(n31984), .B(n31985), .Z(n31983) );
  NANDN U32183 ( .A(n31986), .B(n31987), .Z(n31985) );
  NANDN U32184 ( .A(n31987), .B(n31986), .Z(n31982) );
  ANDN U32185 ( .B(B[158]), .A(n54), .Z(n31979) );
  XNOR U32186 ( .A(n31774), .B(n31988), .Z(n31980) );
  XNOR U32187 ( .A(n31773), .B(n31771), .Z(n31988) );
  AND U32188 ( .A(n31989), .B(n31990), .Z(n31771) );
  NANDN U32189 ( .A(n31991), .B(n31992), .Z(n31990) );
  OR U32190 ( .A(n31993), .B(n31994), .Z(n31992) );
  NAND U32191 ( .A(n31994), .B(n31993), .Z(n31989) );
  ANDN U32192 ( .B(B[159]), .A(n55), .Z(n31773) );
  XNOR U32193 ( .A(n31781), .B(n31995), .Z(n31774) );
  XNOR U32194 ( .A(n31780), .B(n31778), .Z(n31995) );
  AND U32195 ( .A(n31996), .B(n31997), .Z(n31778) );
  NANDN U32196 ( .A(n31998), .B(n31999), .Z(n31997) );
  NANDN U32197 ( .A(n32000), .B(n32001), .Z(n31999) );
  NANDN U32198 ( .A(n32001), .B(n32000), .Z(n31996) );
  ANDN U32199 ( .B(B[160]), .A(n56), .Z(n31780) );
  XNOR U32200 ( .A(n31788), .B(n32002), .Z(n31781) );
  XNOR U32201 ( .A(n31787), .B(n31785), .Z(n32002) );
  AND U32202 ( .A(n32003), .B(n32004), .Z(n31785) );
  NANDN U32203 ( .A(n32005), .B(n32006), .Z(n32004) );
  OR U32204 ( .A(n32007), .B(n32008), .Z(n32006) );
  NAND U32205 ( .A(n32008), .B(n32007), .Z(n32003) );
  ANDN U32206 ( .B(B[161]), .A(n57), .Z(n31787) );
  XNOR U32207 ( .A(n31795), .B(n32009), .Z(n31788) );
  XNOR U32208 ( .A(n31794), .B(n31792), .Z(n32009) );
  AND U32209 ( .A(n32010), .B(n32011), .Z(n31792) );
  NANDN U32210 ( .A(n32012), .B(n32013), .Z(n32011) );
  NANDN U32211 ( .A(n32014), .B(n32015), .Z(n32013) );
  NANDN U32212 ( .A(n32015), .B(n32014), .Z(n32010) );
  ANDN U32213 ( .B(B[162]), .A(n58), .Z(n31794) );
  XNOR U32214 ( .A(n31802), .B(n32016), .Z(n31795) );
  XNOR U32215 ( .A(n31801), .B(n31799), .Z(n32016) );
  AND U32216 ( .A(n32017), .B(n32018), .Z(n31799) );
  NANDN U32217 ( .A(n32019), .B(n32020), .Z(n32018) );
  OR U32218 ( .A(n32021), .B(n32022), .Z(n32020) );
  NAND U32219 ( .A(n32022), .B(n32021), .Z(n32017) );
  ANDN U32220 ( .B(B[163]), .A(n59), .Z(n31801) );
  XNOR U32221 ( .A(n31809), .B(n32023), .Z(n31802) );
  XNOR U32222 ( .A(n31808), .B(n31806), .Z(n32023) );
  AND U32223 ( .A(n32024), .B(n32025), .Z(n31806) );
  NANDN U32224 ( .A(n32026), .B(n32027), .Z(n32025) );
  NANDN U32225 ( .A(n32028), .B(n32029), .Z(n32027) );
  NANDN U32226 ( .A(n32029), .B(n32028), .Z(n32024) );
  ANDN U32227 ( .B(B[164]), .A(n60), .Z(n31808) );
  XNOR U32228 ( .A(n31816), .B(n32030), .Z(n31809) );
  XNOR U32229 ( .A(n31815), .B(n31813), .Z(n32030) );
  AND U32230 ( .A(n32031), .B(n32032), .Z(n31813) );
  NANDN U32231 ( .A(n32033), .B(n32034), .Z(n32032) );
  OR U32232 ( .A(n32035), .B(n32036), .Z(n32034) );
  NAND U32233 ( .A(n32036), .B(n32035), .Z(n32031) );
  ANDN U32234 ( .B(B[165]), .A(n61), .Z(n31815) );
  XNOR U32235 ( .A(n31823), .B(n32037), .Z(n31816) );
  XNOR U32236 ( .A(n31822), .B(n31820), .Z(n32037) );
  AND U32237 ( .A(n32038), .B(n32039), .Z(n31820) );
  NANDN U32238 ( .A(n32040), .B(n32041), .Z(n32039) );
  NANDN U32239 ( .A(n32042), .B(n32043), .Z(n32041) );
  NANDN U32240 ( .A(n32043), .B(n32042), .Z(n32038) );
  ANDN U32241 ( .B(B[166]), .A(n62), .Z(n31822) );
  XNOR U32242 ( .A(n31830), .B(n32044), .Z(n31823) );
  XNOR U32243 ( .A(n31829), .B(n31827), .Z(n32044) );
  AND U32244 ( .A(n32045), .B(n32046), .Z(n31827) );
  NANDN U32245 ( .A(n32047), .B(n32048), .Z(n32046) );
  OR U32246 ( .A(n32049), .B(n32050), .Z(n32048) );
  NAND U32247 ( .A(n32050), .B(n32049), .Z(n32045) );
  ANDN U32248 ( .B(B[167]), .A(n63), .Z(n31829) );
  XNOR U32249 ( .A(n31837), .B(n32051), .Z(n31830) );
  XNOR U32250 ( .A(n31836), .B(n31834), .Z(n32051) );
  AND U32251 ( .A(n32052), .B(n32053), .Z(n31834) );
  NANDN U32252 ( .A(n32054), .B(n32055), .Z(n32053) );
  NANDN U32253 ( .A(n32056), .B(n32057), .Z(n32055) );
  NANDN U32254 ( .A(n32057), .B(n32056), .Z(n32052) );
  ANDN U32255 ( .B(B[168]), .A(n64), .Z(n31836) );
  XNOR U32256 ( .A(n31844), .B(n32058), .Z(n31837) );
  XNOR U32257 ( .A(n31843), .B(n31841), .Z(n32058) );
  AND U32258 ( .A(n32059), .B(n32060), .Z(n31841) );
  NANDN U32259 ( .A(n32061), .B(n32062), .Z(n32060) );
  OR U32260 ( .A(n32063), .B(n32064), .Z(n32062) );
  NAND U32261 ( .A(n32064), .B(n32063), .Z(n32059) );
  ANDN U32262 ( .B(B[169]), .A(n65), .Z(n31843) );
  XNOR U32263 ( .A(n31851), .B(n32065), .Z(n31844) );
  XNOR U32264 ( .A(n31850), .B(n31848), .Z(n32065) );
  AND U32265 ( .A(n32066), .B(n32067), .Z(n31848) );
  NANDN U32266 ( .A(n32068), .B(n32069), .Z(n32067) );
  NANDN U32267 ( .A(n32070), .B(n32071), .Z(n32069) );
  NANDN U32268 ( .A(n32071), .B(n32070), .Z(n32066) );
  ANDN U32269 ( .B(B[170]), .A(n66), .Z(n31850) );
  XNOR U32270 ( .A(n31858), .B(n32072), .Z(n31851) );
  XNOR U32271 ( .A(n31857), .B(n31855), .Z(n32072) );
  AND U32272 ( .A(n32073), .B(n32074), .Z(n31855) );
  NANDN U32273 ( .A(n32075), .B(n32076), .Z(n32074) );
  OR U32274 ( .A(n32077), .B(n32078), .Z(n32076) );
  NAND U32275 ( .A(n32078), .B(n32077), .Z(n32073) );
  ANDN U32276 ( .B(B[171]), .A(n67), .Z(n31857) );
  XNOR U32277 ( .A(n31865), .B(n32079), .Z(n31858) );
  XNOR U32278 ( .A(n31864), .B(n31862), .Z(n32079) );
  AND U32279 ( .A(n32080), .B(n32081), .Z(n31862) );
  NANDN U32280 ( .A(n32082), .B(n32083), .Z(n32081) );
  NANDN U32281 ( .A(n32084), .B(n32085), .Z(n32083) );
  NANDN U32282 ( .A(n32085), .B(n32084), .Z(n32080) );
  ANDN U32283 ( .B(B[172]), .A(n68), .Z(n31864) );
  XNOR U32284 ( .A(n31872), .B(n32086), .Z(n31865) );
  XNOR U32285 ( .A(n31871), .B(n31869), .Z(n32086) );
  AND U32286 ( .A(n32087), .B(n32088), .Z(n31869) );
  NANDN U32287 ( .A(n32089), .B(n32090), .Z(n32088) );
  OR U32288 ( .A(n32091), .B(n32092), .Z(n32090) );
  NAND U32289 ( .A(n32092), .B(n32091), .Z(n32087) );
  ANDN U32290 ( .B(B[173]), .A(n69), .Z(n31871) );
  XNOR U32291 ( .A(n31879), .B(n32093), .Z(n31872) );
  XNOR U32292 ( .A(n31878), .B(n31876), .Z(n32093) );
  AND U32293 ( .A(n32094), .B(n32095), .Z(n31876) );
  NANDN U32294 ( .A(n32096), .B(n32097), .Z(n32095) );
  NANDN U32295 ( .A(n32098), .B(n32099), .Z(n32097) );
  NANDN U32296 ( .A(n32099), .B(n32098), .Z(n32094) );
  ANDN U32297 ( .B(B[174]), .A(n70), .Z(n31878) );
  XNOR U32298 ( .A(n31886), .B(n32100), .Z(n31879) );
  XNOR U32299 ( .A(n31885), .B(n31883), .Z(n32100) );
  AND U32300 ( .A(n32101), .B(n32102), .Z(n31883) );
  NANDN U32301 ( .A(n32103), .B(n32104), .Z(n32102) );
  OR U32302 ( .A(n32105), .B(n32106), .Z(n32104) );
  NAND U32303 ( .A(n32106), .B(n32105), .Z(n32101) );
  ANDN U32304 ( .B(B[175]), .A(n71), .Z(n31885) );
  XNOR U32305 ( .A(n31893), .B(n32107), .Z(n31886) );
  XNOR U32306 ( .A(n31892), .B(n31890), .Z(n32107) );
  AND U32307 ( .A(n32108), .B(n32109), .Z(n31890) );
  NANDN U32308 ( .A(n32110), .B(n32111), .Z(n32109) );
  NANDN U32309 ( .A(n32112), .B(n32113), .Z(n32111) );
  NANDN U32310 ( .A(n32113), .B(n32112), .Z(n32108) );
  ANDN U32311 ( .B(B[176]), .A(n72), .Z(n31892) );
  XNOR U32312 ( .A(n31900), .B(n32114), .Z(n31893) );
  XNOR U32313 ( .A(n31899), .B(n31897), .Z(n32114) );
  AND U32314 ( .A(n32115), .B(n32116), .Z(n31897) );
  NANDN U32315 ( .A(n32117), .B(n32118), .Z(n32116) );
  OR U32316 ( .A(n32119), .B(n32120), .Z(n32118) );
  NAND U32317 ( .A(n32120), .B(n32119), .Z(n32115) );
  ANDN U32318 ( .B(B[177]), .A(n73), .Z(n31899) );
  XNOR U32319 ( .A(n31907), .B(n32121), .Z(n31900) );
  XNOR U32320 ( .A(n31906), .B(n31904), .Z(n32121) );
  AND U32321 ( .A(n32122), .B(n32123), .Z(n31904) );
  NANDN U32322 ( .A(n32124), .B(n32125), .Z(n32123) );
  NANDN U32323 ( .A(n32126), .B(n32127), .Z(n32125) );
  NANDN U32324 ( .A(n32127), .B(n32126), .Z(n32122) );
  ANDN U32325 ( .B(B[178]), .A(n74), .Z(n31906) );
  XNOR U32326 ( .A(n31914), .B(n32128), .Z(n31907) );
  XNOR U32327 ( .A(n31913), .B(n31911), .Z(n32128) );
  AND U32328 ( .A(n32129), .B(n32130), .Z(n31911) );
  NANDN U32329 ( .A(n32131), .B(n32132), .Z(n32130) );
  OR U32330 ( .A(n32133), .B(n32134), .Z(n32132) );
  NAND U32331 ( .A(n32134), .B(n32133), .Z(n32129) );
  ANDN U32332 ( .B(B[179]), .A(n75), .Z(n31913) );
  XNOR U32333 ( .A(n31921), .B(n32135), .Z(n31914) );
  XNOR U32334 ( .A(n31920), .B(n31918), .Z(n32135) );
  AND U32335 ( .A(n32136), .B(n32137), .Z(n31918) );
  NANDN U32336 ( .A(n32138), .B(n32139), .Z(n32137) );
  NANDN U32337 ( .A(n32140), .B(n32141), .Z(n32139) );
  NANDN U32338 ( .A(n32141), .B(n32140), .Z(n32136) );
  ANDN U32339 ( .B(B[180]), .A(n76), .Z(n31920) );
  XNOR U32340 ( .A(n31928), .B(n32142), .Z(n31921) );
  XNOR U32341 ( .A(n31927), .B(n31925), .Z(n32142) );
  AND U32342 ( .A(n32143), .B(n32144), .Z(n31925) );
  NANDN U32343 ( .A(n32145), .B(n32146), .Z(n32144) );
  OR U32344 ( .A(n32147), .B(n32148), .Z(n32146) );
  NAND U32345 ( .A(n32148), .B(n32147), .Z(n32143) );
  ANDN U32346 ( .B(B[181]), .A(n77), .Z(n31927) );
  XNOR U32347 ( .A(n31935), .B(n32149), .Z(n31928) );
  XNOR U32348 ( .A(n31934), .B(n31932), .Z(n32149) );
  AND U32349 ( .A(n32150), .B(n32151), .Z(n31932) );
  NANDN U32350 ( .A(n32152), .B(n32153), .Z(n32151) );
  NANDN U32351 ( .A(n32154), .B(n32155), .Z(n32153) );
  NANDN U32352 ( .A(n32155), .B(n32154), .Z(n32150) );
  ANDN U32353 ( .B(B[182]), .A(n78), .Z(n31934) );
  XNOR U32354 ( .A(n31942), .B(n32156), .Z(n31935) );
  XNOR U32355 ( .A(n31941), .B(n31939), .Z(n32156) );
  AND U32356 ( .A(n32157), .B(n32158), .Z(n31939) );
  NANDN U32357 ( .A(n32159), .B(n32160), .Z(n32158) );
  OR U32358 ( .A(n32161), .B(n32162), .Z(n32160) );
  NAND U32359 ( .A(n32162), .B(n32161), .Z(n32157) );
  ANDN U32360 ( .B(B[183]), .A(n79), .Z(n31941) );
  XNOR U32361 ( .A(n31949), .B(n32163), .Z(n31942) );
  XNOR U32362 ( .A(n31948), .B(n31946), .Z(n32163) );
  AND U32363 ( .A(n32164), .B(n32165), .Z(n31946) );
  NANDN U32364 ( .A(n32166), .B(n32167), .Z(n32165) );
  NANDN U32365 ( .A(n32168), .B(n32169), .Z(n32167) );
  NANDN U32366 ( .A(n32169), .B(n32168), .Z(n32164) );
  ANDN U32367 ( .B(B[184]), .A(n80), .Z(n31948) );
  XNOR U32368 ( .A(n31956), .B(n32170), .Z(n31949) );
  XNOR U32369 ( .A(n31955), .B(n31953), .Z(n32170) );
  AND U32370 ( .A(n32171), .B(n32172), .Z(n31953) );
  NANDN U32371 ( .A(n32173), .B(n32174), .Z(n32172) );
  OR U32372 ( .A(n32175), .B(n32176), .Z(n32174) );
  NAND U32373 ( .A(n32176), .B(n32175), .Z(n32171) );
  ANDN U32374 ( .B(B[185]), .A(n81), .Z(n31955) );
  XNOR U32375 ( .A(n31963), .B(n32177), .Z(n31956) );
  XNOR U32376 ( .A(n31962), .B(n31960), .Z(n32177) );
  AND U32377 ( .A(n32178), .B(n32179), .Z(n31960) );
  NANDN U32378 ( .A(n32180), .B(n32181), .Z(n32179) );
  NAND U32379 ( .A(n32182), .B(n32183), .Z(n32181) );
  ANDN U32380 ( .B(B[186]), .A(n82), .Z(n31962) );
  XOR U32381 ( .A(n31969), .B(n32184), .Z(n31963) );
  XNOR U32382 ( .A(n31967), .B(n31970), .Z(n32184) );
  NAND U32383 ( .A(A[2]), .B(B[187]), .Z(n31970) );
  NANDN U32384 ( .A(n32185), .B(n32186), .Z(n31967) );
  AND U32385 ( .A(A[0]), .B(B[188]), .Z(n32186) );
  XNOR U32386 ( .A(n31972), .B(n32187), .Z(n31969) );
  NAND U32387 ( .A(A[0]), .B(B[189]), .Z(n32187) );
  NAND U32388 ( .A(B[188]), .B(A[1]), .Z(n31972) );
  NAND U32389 ( .A(n32188), .B(n32189), .Z(n418) );
  NANDN U32390 ( .A(n32190), .B(n32191), .Z(n32189) );
  OR U32391 ( .A(n32192), .B(n32193), .Z(n32191) );
  NAND U32392 ( .A(n32193), .B(n32192), .Z(n32188) );
  XOR U32393 ( .A(n420), .B(n419), .Z(\A1[186] ) );
  XOR U32394 ( .A(n32193), .B(n32194), .Z(n419) );
  XNOR U32395 ( .A(n32192), .B(n32190), .Z(n32194) );
  AND U32396 ( .A(n32195), .B(n32196), .Z(n32190) );
  NANDN U32397 ( .A(n32197), .B(n32198), .Z(n32196) );
  NANDN U32398 ( .A(n32199), .B(n32200), .Z(n32198) );
  NANDN U32399 ( .A(n32200), .B(n32199), .Z(n32195) );
  ANDN U32400 ( .B(B[157]), .A(n54), .Z(n32192) );
  XNOR U32401 ( .A(n31987), .B(n32201), .Z(n32193) );
  XNOR U32402 ( .A(n31986), .B(n31984), .Z(n32201) );
  AND U32403 ( .A(n32202), .B(n32203), .Z(n31984) );
  NANDN U32404 ( .A(n32204), .B(n32205), .Z(n32203) );
  OR U32405 ( .A(n32206), .B(n32207), .Z(n32205) );
  NAND U32406 ( .A(n32207), .B(n32206), .Z(n32202) );
  ANDN U32407 ( .B(B[158]), .A(n55), .Z(n31986) );
  XNOR U32408 ( .A(n31994), .B(n32208), .Z(n31987) );
  XNOR U32409 ( .A(n31993), .B(n31991), .Z(n32208) );
  AND U32410 ( .A(n32209), .B(n32210), .Z(n31991) );
  NANDN U32411 ( .A(n32211), .B(n32212), .Z(n32210) );
  NANDN U32412 ( .A(n32213), .B(n32214), .Z(n32212) );
  NANDN U32413 ( .A(n32214), .B(n32213), .Z(n32209) );
  ANDN U32414 ( .B(B[159]), .A(n56), .Z(n31993) );
  XNOR U32415 ( .A(n32001), .B(n32215), .Z(n31994) );
  XNOR U32416 ( .A(n32000), .B(n31998), .Z(n32215) );
  AND U32417 ( .A(n32216), .B(n32217), .Z(n31998) );
  NANDN U32418 ( .A(n32218), .B(n32219), .Z(n32217) );
  OR U32419 ( .A(n32220), .B(n32221), .Z(n32219) );
  NAND U32420 ( .A(n32221), .B(n32220), .Z(n32216) );
  ANDN U32421 ( .B(B[160]), .A(n57), .Z(n32000) );
  XNOR U32422 ( .A(n32008), .B(n32222), .Z(n32001) );
  XNOR U32423 ( .A(n32007), .B(n32005), .Z(n32222) );
  AND U32424 ( .A(n32223), .B(n32224), .Z(n32005) );
  NANDN U32425 ( .A(n32225), .B(n32226), .Z(n32224) );
  NANDN U32426 ( .A(n32227), .B(n32228), .Z(n32226) );
  NANDN U32427 ( .A(n32228), .B(n32227), .Z(n32223) );
  ANDN U32428 ( .B(B[161]), .A(n58), .Z(n32007) );
  XNOR U32429 ( .A(n32015), .B(n32229), .Z(n32008) );
  XNOR U32430 ( .A(n32014), .B(n32012), .Z(n32229) );
  AND U32431 ( .A(n32230), .B(n32231), .Z(n32012) );
  NANDN U32432 ( .A(n32232), .B(n32233), .Z(n32231) );
  OR U32433 ( .A(n32234), .B(n32235), .Z(n32233) );
  NAND U32434 ( .A(n32235), .B(n32234), .Z(n32230) );
  ANDN U32435 ( .B(B[162]), .A(n59), .Z(n32014) );
  XNOR U32436 ( .A(n32022), .B(n32236), .Z(n32015) );
  XNOR U32437 ( .A(n32021), .B(n32019), .Z(n32236) );
  AND U32438 ( .A(n32237), .B(n32238), .Z(n32019) );
  NANDN U32439 ( .A(n32239), .B(n32240), .Z(n32238) );
  NANDN U32440 ( .A(n32241), .B(n32242), .Z(n32240) );
  NANDN U32441 ( .A(n32242), .B(n32241), .Z(n32237) );
  ANDN U32442 ( .B(B[163]), .A(n60), .Z(n32021) );
  XNOR U32443 ( .A(n32029), .B(n32243), .Z(n32022) );
  XNOR U32444 ( .A(n32028), .B(n32026), .Z(n32243) );
  AND U32445 ( .A(n32244), .B(n32245), .Z(n32026) );
  NANDN U32446 ( .A(n32246), .B(n32247), .Z(n32245) );
  OR U32447 ( .A(n32248), .B(n32249), .Z(n32247) );
  NAND U32448 ( .A(n32249), .B(n32248), .Z(n32244) );
  ANDN U32449 ( .B(B[164]), .A(n61), .Z(n32028) );
  XNOR U32450 ( .A(n32036), .B(n32250), .Z(n32029) );
  XNOR U32451 ( .A(n32035), .B(n32033), .Z(n32250) );
  AND U32452 ( .A(n32251), .B(n32252), .Z(n32033) );
  NANDN U32453 ( .A(n32253), .B(n32254), .Z(n32252) );
  NANDN U32454 ( .A(n32255), .B(n32256), .Z(n32254) );
  NANDN U32455 ( .A(n32256), .B(n32255), .Z(n32251) );
  ANDN U32456 ( .B(B[165]), .A(n62), .Z(n32035) );
  XNOR U32457 ( .A(n32043), .B(n32257), .Z(n32036) );
  XNOR U32458 ( .A(n32042), .B(n32040), .Z(n32257) );
  AND U32459 ( .A(n32258), .B(n32259), .Z(n32040) );
  NANDN U32460 ( .A(n32260), .B(n32261), .Z(n32259) );
  OR U32461 ( .A(n32262), .B(n32263), .Z(n32261) );
  NAND U32462 ( .A(n32263), .B(n32262), .Z(n32258) );
  ANDN U32463 ( .B(B[166]), .A(n63), .Z(n32042) );
  XNOR U32464 ( .A(n32050), .B(n32264), .Z(n32043) );
  XNOR U32465 ( .A(n32049), .B(n32047), .Z(n32264) );
  AND U32466 ( .A(n32265), .B(n32266), .Z(n32047) );
  NANDN U32467 ( .A(n32267), .B(n32268), .Z(n32266) );
  NANDN U32468 ( .A(n32269), .B(n32270), .Z(n32268) );
  NANDN U32469 ( .A(n32270), .B(n32269), .Z(n32265) );
  ANDN U32470 ( .B(B[167]), .A(n64), .Z(n32049) );
  XNOR U32471 ( .A(n32057), .B(n32271), .Z(n32050) );
  XNOR U32472 ( .A(n32056), .B(n32054), .Z(n32271) );
  AND U32473 ( .A(n32272), .B(n32273), .Z(n32054) );
  NANDN U32474 ( .A(n32274), .B(n32275), .Z(n32273) );
  OR U32475 ( .A(n32276), .B(n32277), .Z(n32275) );
  NAND U32476 ( .A(n32277), .B(n32276), .Z(n32272) );
  ANDN U32477 ( .B(B[168]), .A(n65), .Z(n32056) );
  XNOR U32478 ( .A(n32064), .B(n32278), .Z(n32057) );
  XNOR U32479 ( .A(n32063), .B(n32061), .Z(n32278) );
  AND U32480 ( .A(n32279), .B(n32280), .Z(n32061) );
  NANDN U32481 ( .A(n32281), .B(n32282), .Z(n32280) );
  NANDN U32482 ( .A(n32283), .B(n32284), .Z(n32282) );
  NANDN U32483 ( .A(n32284), .B(n32283), .Z(n32279) );
  ANDN U32484 ( .B(B[169]), .A(n66), .Z(n32063) );
  XNOR U32485 ( .A(n32071), .B(n32285), .Z(n32064) );
  XNOR U32486 ( .A(n32070), .B(n32068), .Z(n32285) );
  AND U32487 ( .A(n32286), .B(n32287), .Z(n32068) );
  NANDN U32488 ( .A(n32288), .B(n32289), .Z(n32287) );
  OR U32489 ( .A(n32290), .B(n32291), .Z(n32289) );
  NAND U32490 ( .A(n32291), .B(n32290), .Z(n32286) );
  ANDN U32491 ( .B(B[170]), .A(n67), .Z(n32070) );
  XNOR U32492 ( .A(n32078), .B(n32292), .Z(n32071) );
  XNOR U32493 ( .A(n32077), .B(n32075), .Z(n32292) );
  AND U32494 ( .A(n32293), .B(n32294), .Z(n32075) );
  NANDN U32495 ( .A(n32295), .B(n32296), .Z(n32294) );
  NANDN U32496 ( .A(n32297), .B(n32298), .Z(n32296) );
  NANDN U32497 ( .A(n32298), .B(n32297), .Z(n32293) );
  ANDN U32498 ( .B(B[171]), .A(n68), .Z(n32077) );
  XNOR U32499 ( .A(n32085), .B(n32299), .Z(n32078) );
  XNOR U32500 ( .A(n32084), .B(n32082), .Z(n32299) );
  AND U32501 ( .A(n32300), .B(n32301), .Z(n32082) );
  NANDN U32502 ( .A(n32302), .B(n32303), .Z(n32301) );
  OR U32503 ( .A(n32304), .B(n32305), .Z(n32303) );
  NAND U32504 ( .A(n32305), .B(n32304), .Z(n32300) );
  ANDN U32505 ( .B(B[172]), .A(n69), .Z(n32084) );
  XNOR U32506 ( .A(n32092), .B(n32306), .Z(n32085) );
  XNOR U32507 ( .A(n32091), .B(n32089), .Z(n32306) );
  AND U32508 ( .A(n32307), .B(n32308), .Z(n32089) );
  NANDN U32509 ( .A(n32309), .B(n32310), .Z(n32308) );
  NANDN U32510 ( .A(n32311), .B(n32312), .Z(n32310) );
  NANDN U32511 ( .A(n32312), .B(n32311), .Z(n32307) );
  ANDN U32512 ( .B(B[173]), .A(n70), .Z(n32091) );
  XNOR U32513 ( .A(n32099), .B(n32313), .Z(n32092) );
  XNOR U32514 ( .A(n32098), .B(n32096), .Z(n32313) );
  AND U32515 ( .A(n32314), .B(n32315), .Z(n32096) );
  NANDN U32516 ( .A(n32316), .B(n32317), .Z(n32315) );
  OR U32517 ( .A(n32318), .B(n32319), .Z(n32317) );
  NAND U32518 ( .A(n32319), .B(n32318), .Z(n32314) );
  ANDN U32519 ( .B(B[174]), .A(n71), .Z(n32098) );
  XNOR U32520 ( .A(n32106), .B(n32320), .Z(n32099) );
  XNOR U32521 ( .A(n32105), .B(n32103), .Z(n32320) );
  AND U32522 ( .A(n32321), .B(n32322), .Z(n32103) );
  NANDN U32523 ( .A(n32323), .B(n32324), .Z(n32322) );
  NANDN U32524 ( .A(n32325), .B(n32326), .Z(n32324) );
  NANDN U32525 ( .A(n32326), .B(n32325), .Z(n32321) );
  ANDN U32526 ( .B(B[175]), .A(n72), .Z(n32105) );
  XNOR U32527 ( .A(n32113), .B(n32327), .Z(n32106) );
  XNOR U32528 ( .A(n32112), .B(n32110), .Z(n32327) );
  AND U32529 ( .A(n32328), .B(n32329), .Z(n32110) );
  NANDN U32530 ( .A(n32330), .B(n32331), .Z(n32329) );
  OR U32531 ( .A(n32332), .B(n32333), .Z(n32331) );
  NAND U32532 ( .A(n32333), .B(n32332), .Z(n32328) );
  ANDN U32533 ( .B(B[176]), .A(n73), .Z(n32112) );
  XNOR U32534 ( .A(n32120), .B(n32334), .Z(n32113) );
  XNOR U32535 ( .A(n32119), .B(n32117), .Z(n32334) );
  AND U32536 ( .A(n32335), .B(n32336), .Z(n32117) );
  NANDN U32537 ( .A(n32337), .B(n32338), .Z(n32336) );
  NANDN U32538 ( .A(n32339), .B(n32340), .Z(n32338) );
  NANDN U32539 ( .A(n32340), .B(n32339), .Z(n32335) );
  ANDN U32540 ( .B(B[177]), .A(n74), .Z(n32119) );
  XNOR U32541 ( .A(n32127), .B(n32341), .Z(n32120) );
  XNOR U32542 ( .A(n32126), .B(n32124), .Z(n32341) );
  AND U32543 ( .A(n32342), .B(n32343), .Z(n32124) );
  NANDN U32544 ( .A(n32344), .B(n32345), .Z(n32343) );
  OR U32545 ( .A(n32346), .B(n32347), .Z(n32345) );
  NAND U32546 ( .A(n32347), .B(n32346), .Z(n32342) );
  ANDN U32547 ( .B(B[178]), .A(n75), .Z(n32126) );
  XNOR U32548 ( .A(n32134), .B(n32348), .Z(n32127) );
  XNOR U32549 ( .A(n32133), .B(n32131), .Z(n32348) );
  AND U32550 ( .A(n32349), .B(n32350), .Z(n32131) );
  NANDN U32551 ( .A(n32351), .B(n32352), .Z(n32350) );
  NANDN U32552 ( .A(n32353), .B(n32354), .Z(n32352) );
  NANDN U32553 ( .A(n32354), .B(n32353), .Z(n32349) );
  ANDN U32554 ( .B(B[179]), .A(n76), .Z(n32133) );
  XNOR U32555 ( .A(n32141), .B(n32355), .Z(n32134) );
  XNOR U32556 ( .A(n32140), .B(n32138), .Z(n32355) );
  AND U32557 ( .A(n32356), .B(n32357), .Z(n32138) );
  NANDN U32558 ( .A(n32358), .B(n32359), .Z(n32357) );
  OR U32559 ( .A(n32360), .B(n32361), .Z(n32359) );
  NAND U32560 ( .A(n32361), .B(n32360), .Z(n32356) );
  ANDN U32561 ( .B(B[180]), .A(n77), .Z(n32140) );
  XNOR U32562 ( .A(n32148), .B(n32362), .Z(n32141) );
  XNOR U32563 ( .A(n32147), .B(n32145), .Z(n32362) );
  AND U32564 ( .A(n32363), .B(n32364), .Z(n32145) );
  NANDN U32565 ( .A(n32365), .B(n32366), .Z(n32364) );
  NANDN U32566 ( .A(n32367), .B(n32368), .Z(n32366) );
  NANDN U32567 ( .A(n32368), .B(n32367), .Z(n32363) );
  ANDN U32568 ( .B(B[181]), .A(n78), .Z(n32147) );
  XNOR U32569 ( .A(n32155), .B(n32369), .Z(n32148) );
  XNOR U32570 ( .A(n32154), .B(n32152), .Z(n32369) );
  AND U32571 ( .A(n32370), .B(n32371), .Z(n32152) );
  NANDN U32572 ( .A(n32372), .B(n32373), .Z(n32371) );
  OR U32573 ( .A(n32374), .B(n32375), .Z(n32373) );
  NAND U32574 ( .A(n32375), .B(n32374), .Z(n32370) );
  ANDN U32575 ( .B(B[182]), .A(n79), .Z(n32154) );
  XNOR U32576 ( .A(n32162), .B(n32376), .Z(n32155) );
  XNOR U32577 ( .A(n32161), .B(n32159), .Z(n32376) );
  AND U32578 ( .A(n32377), .B(n32378), .Z(n32159) );
  NANDN U32579 ( .A(n32379), .B(n32380), .Z(n32378) );
  NANDN U32580 ( .A(n32381), .B(n32382), .Z(n32380) );
  NANDN U32581 ( .A(n32382), .B(n32381), .Z(n32377) );
  ANDN U32582 ( .B(B[183]), .A(n80), .Z(n32161) );
  XNOR U32583 ( .A(n32169), .B(n32383), .Z(n32162) );
  XNOR U32584 ( .A(n32168), .B(n32166), .Z(n32383) );
  AND U32585 ( .A(n32384), .B(n32385), .Z(n32166) );
  NANDN U32586 ( .A(n32386), .B(n32387), .Z(n32385) );
  OR U32587 ( .A(n32388), .B(n32389), .Z(n32387) );
  NAND U32588 ( .A(n32389), .B(n32388), .Z(n32384) );
  ANDN U32589 ( .B(B[184]), .A(n81), .Z(n32168) );
  XNOR U32590 ( .A(n32176), .B(n32390), .Z(n32169) );
  XNOR U32591 ( .A(n32175), .B(n32173), .Z(n32390) );
  AND U32592 ( .A(n32391), .B(n32392), .Z(n32173) );
  NANDN U32593 ( .A(n32393), .B(n32394), .Z(n32392) );
  NAND U32594 ( .A(n32395), .B(n32396), .Z(n32394) );
  ANDN U32595 ( .B(B[185]), .A(n82), .Z(n32175) );
  XOR U32596 ( .A(n32182), .B(n32397), .Z(n32176) );
  XNOR U32597 ( .A(n32180), .B(n32183), .Z(n32397) );
  NAND U32598 ( .A(A[2]), .B(B[186]), .Z(n32183) );
  NANDN U32599 ( .A(n32398), .B(n32399), .Z(n32180) );
  AND U32600 ( .A(A[0]), .B(B[187]), .Z(n32399) );
  XNOR U32601 ( .A(n32185), .B(n32400), .Z(n32182) );
  NAND U32602 ( .A(A[0]), .B(B[188]), .Z(n32400) );
  NAND U32603 ( .A(B[187]), .B(A[1]), .Z(n32185) );
  NAND U32604 ( .A(n32401), .B(n32402), .Z(n420) );
  NANDN U32605 ( .A(n32403), .B(n32404), .Z(n32402) );
  OR U32606 ( .A(n32405), .B(n32406), .Z(n32404) );
  NAND U32607 ( .A(n32406), .B(n32405), .Z(n32401) );
  XOR U32608 ( .A(n422), .B(n421), .Z(\A1[185] ) );
  XOR U32609 ( .A(n32406), .B(n32407), .Z(n421) );
  XNOR U32610 ( .A(n32405), .B(n32403), .Z(n32407) );
  AND U32611 ( .A(n32408), .B(n32409), .Z(n32403) );
  NANDN U32612 ( .A(n32410), .B(n32411), .Z(n32409) );
  NANDN U32613 ( .A(n32412), .B(n32413), .Z(n32411) );
  NANDN U32614 ( .A(n32413), .B(n32412), .Z(n32408) );
  ANDN U32615 ( .B(B[156]), .A(n54), .Z(n32405) );
  XNOR U32616 ( .A(n32200), .B(n32414), .Z(n32406) );
  XNOR U32617 ( .A(n32199), .B(n32197), .Z(n32414) );
  AND U32618 ( .A(n32415), .B(n32416), .Z(n32197) );
  NANDN U32619 ( .A(n32417), .B(n32418), .Z(n32416) );
  OR U32620 ( .A(n32419), .B(n32420), .Z(n32418) );
  NAND U32621 ( .A(n32420), .B(n32419), .Z(n32415) );
  ANDN U32622 ( .B(B[157]), .A(n55), .Z(n32199) );
  XNOR U32623 ( .A(n32207), .B(n32421), .Z(n32200) );
  XNOR U32624 ( .A(n32206), .B(n32204), .Z(n32421) );
  AND U32625 ( .A(n32422), .B(n32423), .Z(n32204) );
  NANDN U32626 ( .A(n32424), .B(n32425), .Z(n32423) );
  NANDN U32627 ( .A(n32426), .B(n32427), .Z(n32425) );
  NANDN U32628 ( .A(n32427), .B(n32426), .Z(n32422) );
  ANDN U32629 ( .B(B[158]), .A(n56), .Z(n32206) );
  XNOR U32630 ( .A(n32214), .B(n32428), .Z(n32207) );
  XNOR U32631 ( .A(n32213), .B(n32211), .Z(n32428) );
  AND U32632 ( .A(n32429), .B(n32430), .Z(n32211) );
  NANDN U32633 ( .A(n32431), .B(n32432), .Z(n32430) );
  OR U32634 ( .A(n32433), .B(n32434), .Z(n32432) );
  NAND U32635 ( .A(n32434), .B(n32433), .Z(n32429) );
  ANDN U32636 ( .B(B[159]), .A(n57), .Z(n32213) );
  XNOR U32637 ( .A(n32221), .B(n32435), .Z(n32214) );
  XNOR U32638 ( .A(n32220), .B(n32218), .Z(n32435) );
  AND U32639 ( .A(n32436), .B(n32437), .Z(n32218) );
  NANDN U32640 ( .A(n32438), .B(n32439), .Z(n32437) );
  NANDN U32641 ( .A(n32440), .B(n32441), .Z(n32439) );
  NANDN U32642 ( .A(n32441), .B(n32440), .Z(n32436) );
  ANDN U32643 ( .B(B[160]), .A(n58), .Z(n32220) );
  XNOR U32644 ( .A(n32228), .B(n32442), .Z(n32221) );
  XNOR U32645 ( .A(n32227), .B(n32225), .Z(n32442) );
  AND U32646 ( .A(n32443), .B(n32444), .Z(n32225) );
  NANDN U32647 ( .A(n32445), .B(n32446), .Z(n32444) );
  OR U32648 ( .A(n32447), .B(n32448), .Z(n32446) );
  NAND U32649 ( .A(n32448), .B(n32447), .Z(n32443) );
  ANDN U32650 ( .B(B[161]), .A(n59), .Z(n32227) );
  XNOR U32651 ( .A(n32235), .B(n32449), .Z(n32228) );
  XNOR U32652 ( .A(n32234), .B(n32232), .Z(n32449) );
  AND U32653 ( .A(n32450), .B(n32451), .Z(n32232) );
  NANDN U32654 ( .A(n32452), .B(n32453), .Z(n32451) );
  NANDN U32655 ( .A(n32454), .B(n32455), .Z(n32453) );
  NANDN U32656 ( .A(n32455), .B(n32454), .Z(n32450) );
  ANDN U32657 ( .B(B[162]), .A(n60), .Z(n32234) );
  XNOR U32658 ( .A(n32242), .B(n32456), .Z(n32235) );
  XNOR U32659 ( .A(n32241), .B(n32239), .Z(n32456) );
  AND U32660 ( .A(n32457), .B(n32458), .Z(n32239) );
  NANDN U32661 ( .A(n32459), .B(n32460), .Z(n32458) );
  OR U32662 ( .A(n32461), .B(n32462), .Z(n32460) );
  NAND U32663 ( .A(n32462), .B(n32461), .Z(n32457) );
  ANDN U32664 ( .B(B[163]), .A(n61), .Z(n32241) );
  XNOR U32665 ( .A(n32249), .B(n32463), .Z(n32242) );
  XNOR U32666 ( .A(n32248), .B(n32246), .Z(n32463) );
  AND U32667 ( .A(n32464), .B(n32465), .Z(n32246) );
  NANDN U32668 ( .A(n32466), .B(n32467), .Z(n32465) );
  NANDN U32669 ( .A(n32468), .B(n32469), .Z(n32467) );
  NANDN U32670 ( .A(n32469), .B(n32468), .Z(n32464) );
  ANDN U32671 ( .B(B[164]), .A(n62), .Z(n32248) );
  XNOR U32672 ( .A(n32256), .B(n32470), .Z(n32249) );
  XNOR U32673 ( .A(n32255), .B(n32253), .Z(n32470) );
  AND U32674 ( .A(n32471), .B(n32472), .Z(n32253) );
  NANDN U32675 ( .A(n32473), .B(n32474), .Z(n32472) );
  OR U32676 ( .A(n32475), .B(n32476), .Z(n32474) );
  NAND U32677 ( .A(n32476), .B(n32475), .Z(n32471) );
  ANDN U32678 ( .B(B[165]), .A(n63), .Z(n32255) );
  XNOR U32679 ( .A(n32263), .B(n32477), .Z(n32256) );
  XNOR U32680 ( .A(n32262), .B(n32260), .Z(n32477) );
  AND U32681 ( .A(n32478), .B(n32479), .Z(n32260) );
  NANDN U32682 ( .A(n32480), .B(n32481), .Z(n32479) );
  NANDN U32683 ( .A(n32482), .B(n32483), .Z(n32481) );
  NANDN U32684 ( .A(n32483), .B(n32482), .Z(n32478) );
  ANDN U32685 ( .B(B[166]), .A(n64), .Z(n32262) );
  XNOR U32686 ( .A(n32270), .B(n32484), .Z(n32263) );
  XNOR U32687 ( .A(n32269), .B(n32267), .Z(n32484) );
  AND U32688 ( .A(n32485), .B(n32486), .Z(n32267) );
  NANDN U32689 ( .A(n32487), .B(n32488), .Z(n32486) );
  OR U32690 ( .A(n32489), .B(n32490), .Z(n32488) );
  NAND U32691 ( .A(n32490), .B(n32489), .Z(n32485) );
  ANDN U32692 ( .B(B[167]), .A(n65), .Z(n32269) );
  XNOR U32693 ( .A(n32277), .B(n32491), .Z(n32270) );
  XNOR U32694 ( .A(n32276), .B(n32274), .Z(n32491) );
  AND U32695 ( .A(n32492), .B(n32493), .Z(n32274) );
  NANDN U32696 ( .A(n32494), .B(n32495), .Z(n32493) );
  NANDN U32697 ( .A(n32496), .B(n32497), .Z(n32495) );
  NANDN U32698 ( .A(n32497), .B(n32496), .Z(n32492) );
  ANDN U32699 ( .B(B[168]), .A(n66), .Z(n32276) );
  XNOR U32700 ( .A(n32284), .B(n32498), .Z(n32277) );
  XNOR U32701 ( .A(n32283), .B(n32281), .Z(n32498) );
  AND U32702 ( .A(n32499), .B(n32500), .Z(n32281) );
  NANDN U32703 ( .A(n32501), .B(n32502), .Z(n32500) );
  OR U32704 ( .A(n32503), .B(n32504), .Z(n32502) );
  NAND U32705 ( .A(n32504), .B(n32503), .Z(n32499) );
  ANDN U32706 ( .B(B[169]), .A(n67), .Z(n32283) );
  XNOR U32707 ( .A(n32291), .B(n32505), .Z(n32284) );
  XNOR U32708 ( .A(n32290), .B(n32288), .Z(n32505) );
  AND U32709 ( .A(n32506), .B(n32507), .Z(n32288) );
  NANDN U32710 ( .A(n32508), .B(n32509), .Z(n32507) );
  NANDN U32711 ( .A(n32510), .B(n32511), .Z(n32509) );
  NANDN U32712 ( .A(n32511), .B(n32510), .Z(n32506) );
  ANDN U32713 ( .B(B[170]), .A(n68), .Z(n32290) );
  XNOR U32714 ( .A(n32298), .B(n32512), .Z(n32291) );
  XNOR U32715 ( .A(n32297), .B(n32295), .Z(n32512) );
  AND U32716 ( .A(n32513), .B(n32514), .Z(n32295) );
  NANDN U32717 ( .A(n32515), .B(n32516), .Z(n32514) );
  OR U32718 ( .A(n32517), .B(n32518), .Z(n32516) );
  NAND U32719 ( .A(n32518), .B(n32517), .Z(n32513) );
  ANDN U32720 ( .B(B[171]), .A(n69), .Z(n32297) );
  XNOR U32721 ( .A(n32305), .B(n32519), .Z(n32298) );
  XNOR U32722 ( .A(n32304), .B(n32302), .Z(n32519) );
  AND U32723 ( .A(n32520), .B(n32521), .Z(n32302) );
  NANDN U32724 ( .A(n32522), .B(n32523), .Z(n32521) );
  NANDN U32725 ( .A(n32524), .B(n32525), .Z(n32523) );
  NANDN U32726 ( .A(n32525), .B(n32524), .Z(n32520) );
  ANDN U32727 ( .B(B[172]), .A(n70), .Z(n32304) );
  XNOR U32728 ( .A(n32312), .B(n32526), .Z(n32305) );
  XNOR U32729 ( .A(n32311), .B(n32309), .Z(n32526) );
  AND U32730 ( .A(n32527), .B(n32528), .Z(n32309) );
  NANDN U32731 ( .A(n32529), .B(n32530), .Z(n32528) );
  OR U32732 ( .A(n32531), .B(n32532), .Z(n32530) );
  NAND U32733 ( .A(n32532), .B(n32531), .Z(n32527) );
  ANDN U32734 ( .B(B[173]), .A(n71), .Z(n32311) );
  XNOR U32735 ( .A(n32319), .B(n32533), .Z(n32312) );
  XNOR U32736 ( .A(n32318), .B(n32316), .Z(n32533) );
  AND U32737 ( .A(n32534), .B(n32535), .Z(n32316) );
  NANDN U32738 ( .A(n32536), .B(n32537), .Z(n32535) );
  NANDN U32739 ( .A(n32538), .B(n32539), .Z(n32537) );
  NANDN U32740 ( .A(n32539), .B(n32538), .Z(n32534) );
  ANDN U32741 ( .B(B[174]), .A(n72), .Z(n32318) );
  XNOR U32742 ( .A(n32326), .B(n32540), .Z(n32319) );
  XNOR U32743 ( .A(n32325), .B(n32323), .Z(n32540) );
  AND U32744 ( .A(n32541), .B(n32542), .Z(n32323) );
  NANDN U32745 ( .A(n32543), .B(n32544), .Z(n32542) );
  OR U32746 ( .A(n32545), .B(n32546), .Z(n32544) );
  NAND U32747 ( .A(n32546), .B(n32545), .Z(n32541) );
  ANDN U32748 ( .B(B[175]), .A(n73), .Z(n32325) );
  XNOR U32749 ( .A(n32333), .B(n32547), .Z(n32326) );
  XNOR U32750 ( .A(n32332), .B(n32330), .Z(n32547) );
  AND U32751 ( .A(n32548), .B(n32549), .Z(n32330) );
  NANDN U32752 ( .A(n32550), .B(n32551), .Z(n32549) );
  NANDN U32753 ( .A(n32552), .B(n32553), .Z(n32551) );
  NANDN U32754 ( .A(n32553), .B(n32552), .Z(n32548) );
  ANDN U32755 ( .B(B[176]), .A(n74), .Z(n32332) );
  XNOR U32756 ( .A(n32340), .B(n32554), .Z(n32333) );
  XNOR U32757 ( .A(n32339), .B(n32337), .Z(n32554) );
  AND U32758 ( .A(n32555), .B(n32556), .Z(n32337) );
  NANDN U32759 ( .A(n32557), .B(n32558), .Z(n32556) );
  OR U32760 ( .A(n32559), .B(n32560), .Z(n32558) );
  NAND U32761 ( .A(n32560), .B(n32559), .Z(n32555) );
  ANDN U32762 ( .B(B[177]), .A(n75), .Z(n32339) );
  XNOR U32763 ( .A(n32347), .B(n32561), .Z(n32340) );
  XNOR U32764 ( .A(n32346), .B(n32344), .Z(n32561) );
  AND U32765 ( .A(n32562), .B(n32563), .Z(n32344) );
  NANDN U32766 ( .A(n32564), .B(n32565), .Z(n32563) );
  NANDN U32767 ( .A(n32566), .B(n32567), .Z(n32565) );
  NANDN U32768 ( .A(n32567), .B(n32566), .Z(n32562) );
  ANDN U32769 ( .B(B[178]), .A(n76), .Z(n32346) );
  XNOR U32770 ( .A(n32354), .B(n32568), .Z(n32347) );
  XNOR U32771 ( .A(n32353), .B(n32351), .Z(n32568) );
  AND U32772 ( .A(n32569), .B(n32570), .Z(n32351) );
  NANDN U32773 ( .A(n32571), .B(n32572), .Z(n32570) );
  OR U32774 ( .A(n32573), .B(n32574), .Z(n32572) );
  NAND U32775 ( .A(n32574), .B(n32573), .Z(n32569) );
  ANDN U32776 ( .B(B[179]), .A(n77), .Z(n32353) );
  XNOR U32777 ( .A(n32361), .B(n32575), .Z(n32354) );
  XNOR U32778 ( .A(n32360), .B(n32358), .Z(n32575) );
  AND U32779 ( .A(n32576), .B(n32577), .Z(n32358) );
  NANDN U32780 ( .A(n32578), .B(n32579), .Z(n32577) );
  NANDN U32781 ( .A(n32580), .B(n32581), .Z(n32579) );
  NANDN U32782 ( .A(n32581), .B(n32580), .Z(n32576) );
  ANDN U32783 ( .B(B[180]), .A(n78), .Z(n32360) );
  XNOR U32784 ( .A(n32368), .B(n32582), .Z(n32361) );
  XNOR U32785 ( .A(n32367), .B(n32365), .Z(n32582) );
  AND U32786 ( .A(n32583), .B(n32584), .Z(n32365) );
  NANDN U32787 ( .A(n32585), .B(n32586), .Z(n32584) );
  OR U32788 ( .A(n32587), .B(n32588), .Z(n32586) );
  NAND U32789 ( .A(n32588), .B(n32587), .Z(n32583) );
  ANDN U32790 ( .B(B[181]), .A(n79), .Z(n32367) );
  XNOR U32791 ( .A(n32375), .B(n32589), .Z(n32368) );
  XNOR U32792 ( .A(n32374), .B(n32372), .Z(n32589) );
  AND U32793 ( .A(n32590), .B(n32591), .Z(n32372) );
  NANDN U32794 ( .A(n32592), .B(n32593), .Z(n32591) );
  NANDN U32795 ( .A(n32594), .B(n32595), .Z(n32593) );
  NANDN U32796 ( .A(n32595), .B(n32594), .Z(n32590) );
  ANDN U32797 ( .B(B[182]), .A(n80), .Z(n32374) );
  XNOR U32798 ( .A(n32382), .B(n32596), .Z(n32375) );
  XNOR U32799 ( .A(n32381), .B(n32379), .Z(n32596) );
  AND U32800 ( .A(n32597), .B(n32598), .Z(n32379) );
  NANDN U32801 ( .A(n32599), .B(n32600), .Z(n32598) );
  OR U32802 ( .A(n32601), .B(n32602), .Z(n32600) );
  NAND U32803 ( .A(n32602), .B(n32601), .Z(n32597) );
  ANDN U32804 ( .B(B[183]), .A(n81), .Z(n32381) );
  XNOR U32805 ( .A(n32389), .B(n32603), .Z(n32382) );
  XNOR U32806 ( .A(n32388), .B(n32386), .Z(n32603) );
  AND U32807 ( .A(n32604), .B(n32605), .Z(n32386) );
  NANDN U32808 ( .A(n32606), .B(n32607), .Z(n32605) );
  NAND U32809 ( .A(n32608), .B(n32609), .Z(n32607) );
  ANDN U32810 ( .B(B[184]), .A(n82), .Z(n32388) );
  XOR U32811 ( .A(n32395), .B(n32610), .Z(n32389) );
  XNOR U32812 ( .A(n32393), .B(n32396), .Z(n32610) );
  NAND U32813 ( .A(A[2]), .B(B[185]), .Z(n32396) );
  NANDN U32814 ( .A(n32611), .B(n32612), .Z(n32393) );
  AND U32815 ( .A(A[0]), .B(B[186]), .Z(n32612) );
  XNOR U32816 ( .A(n32398), .B(n32613), .Z(n32395) );
  NAND U32817 ( .A(A[0]), .B(B[187]), .Z(n32613) );
  NAND U32818 ( .A(B[186]), .B(A[1]), .Z(n32398) );
  NAND U32819 ( .A(n32614), .B(n32615), .Z(n422) );
  NANDN U32820 ( .A(n32616), .B(n32617), .Z(n32615) );
  OR U32821 ( .A(n32618), .B(n32619), .Z(n32617) );
  NAND U32822 ( .A(n32619), .B(n32618), .Z(n32614) );
  XOR U32823 ( .A(n424), .B(n423), .Z(\A1[184] ) );
  XOR U32824 ( .A(n32619), .B(n32620), .Z(n423) );
  XNOR U32825 ( .A(n32618), .B(n32616), .Z(n32620) );
  AND U32826 ( .A(n32621), .B(n32622), .Z(n32616) );
  NANDN U32827 ( .A(n32623), .B(n32624), .Z(n32622) );
  NANDN U32828 ( .A(n32625), .B(n32626), .Z(n32624) );
  NANDN U32829 ( .A(n32626), .B(n32625), .Z(n32621) );
  ANDN U32830 ( .B(B[155]), .A(n54), .Z(n32618) );
  XNOR U32831 ( .A(n32413), .B(n32627), .Z(n32619) );
  XNOR U32832 ( .A(n32412), .B(n32410), .Z(n32627) );
  AND U32833 ( .A(n32628), .B(n32629), .Z(n32410) );
  NANDN U32834 ( .A(n32630), .B(n32631), .Z(n32629) );
  OR U32835 ( .A(n32632), .B(n32633), .Z(n32631) );
  NAND U32836 ( .A(n32633), .B(n32632), .Z(n32628) );
  ANDN U32837 ( .B(B[156]), .A(n55), .Z(n32412) );
  XNOR U32838 ( .A(n32420), .B(n32634), .Z(n32413) );
  XNOR U32839 ( .A(n32419), .B(n32417), .Z(n32634) );
  AND U32840 ( .A(n32635), .B(n32636), .Z(n32417) );
  NANDN U32841 ( .A(n32637), .B(n32638), .Z(n32636) );
  NANDN U32842 ( .A(n32639), .B(n32640), .Z(n32638) );
  NANDN U32843 ( .A(n32640), .B(n32639), .Z(n32635) );
  ANDN U32844 ( .B(B[157]), .A(n56), .Z(n32419) );
  XNOR U32845 ( .A(n32427), .B(n32641), .Z(n32420) );
  XNOR U32846 ( .A(n32426), .B(n32424), .Z(n32641) );
  AND U32847 ( .A(n32642), .B(n32643), .Z(n32424) );
  NANDN U32848 ( .A(n32644), .B(n32645), .Z(n32643) );
  OR U32849 ( .A(n32646), .B(n32647), .Z(n32645) );
  NAND U32850 ( .A(n32647), .B(n32646), .Z(n32642) );
  ANDN U32851 ( .B(B[158]), .A(n57), .Z(n32426) );
  XNOR U32852 ( .A(n32434), .B(n32648), .Z(n32427) );
  XNOR U32853 ( .A(n32433), .B(n32431), .Z(n32648) );
  AND U32854 ( .A(n32649), .B(n32650), .Z(n32431) );
  NANDN U32855 ( .A(n32651), .B(n32652), .Z(n32650) );
  NANDN U32856 ( .A(n32653), .B(n32654), .Z(n32652) );
  NANDN U32857 ( .A(n32654), .B(n32653), .Z(n32649) );
  ANDN U32858 ( .B(B[159]), .A(n58), .Z(n32433) );
  XNOR U32859 ( .A(n32441), .B(n32655), .Z(n32434) );
  XNOR U32860 ( .A(n32440), .B(n32438), .Z(n32655) );
  AND U32861 ( .A(n32656), .B(n32657), .Z(n32438) );
  NANDN U32862 ( .A(n32658), .B(n32659), .Z(n32657) );
  OR U32863 ( .A(n32660), .B(n32661), .Z(n32659) );
  NAND U32864 ( .A(n32661), .B(n32660), .Z(n32656) );
  ANDN U32865 ( .B(B[160]), .A(n59), .Z(n32440) );
  XNOR U32866 ( .A(n32448), .B(n32662), .Z(n32441) );
  XNOR U32867 ( .A(n32447), .B(n32445), .Z(n32662) );
  AND U32868 ( .A(n32663), .B(n32664), .Z(n32445) );
  NANDN U32869 ( .A(n32665), .B(n32666), .Z(n32664) );
  NANDN U32870 ( .A(n32667), .B(n32668), .Z(n32666) );
  NANDN U32871 ( .A(n32668), .B(n32667), .Z(n32663) );
  ANDN U32872 ( .B(B[161]), .A(n60), .Z(n32447) );
  XNOR U32873 ( .A(n32455), .B(n32669), .Z(n32448) );
  XNOR U32874 ( .A(n32454), .B(n32452), .Z(n32669) );
  AND U32875 ( .A(n32670), .B(n32671), .Z(n32452) );
  NANDN U32876 ( .A(n32672), .B(n32673), .Z(n32671) );
  OR U32877 ( .A(n32674), .B(n32675), .Z(n32673) );
  NAND U32878 ( .A(n32675), .B(n32674), .Z(n32670) );
  ANDN U32879 ( .B(B[162]), .A(n61), .Z(n32454) );
  XNOR U32880 ( .A(n32462), .B(n32676), .Z(n32455) );
  XNOR U32881 ( .A(n32461), .B(n32459), .Z(n32676) );
  AND U32882 ( .A(n32677), .B(n32678), .Z(n32459) );
  NANDN U32883 ( .A(n32679), .B(n32680), .Z(n32678) );
  NANDN U32884 ( .A(n32681), .B(n32682), .Z(n32680) );
  NANDN U32885 ( .A(n32682), .B(n32681), .Z(n32677) );
  ANDN U32886 ( .B(B[163]), .A(n62), .Z(n32461) );
  XNOR U32887 ( .A(n32469), .B(n32683), .Z(n32462) );
  XNOR U32888 ( .A(n32468), .B(n32466), .Z(n32683) );
  AND U32889 ( .A(n32684), .B(n32685), .Z(n32466) );
  NANDN U32890 ( .A(n32686), .B(n32687), .Z(n32685) );
  OR U32891 ( .A(n32688), .B(n32689), .Z(n32687) );
  NAND U32892 ( .A(n32689), .B(n32688), .Z(n32684) );
  ANDN U32893 ( .B(B[164]), .A(n63), .Z(n32468) );
  XNOR U32894 ( .A(n32476), .B(n32690), .Z(n32469) );
  XNOR U32895 ( .A(n32475), .B(n32473), .Z(n32690) );
  AND U32896 ( .A(n32691), .B(n32692), .Z(n32473) );
  NANDN U32897 ( .A(n32693), .B(n32694), .Z(n32692) );
  NANDN U32898 ( .A(n32695), .B(n32696), .Z(n32694) );
  NANDN U32899 ( .A(n32696), .B(n32695), .Z(n32691) );
  ANDN U32900 ( .B(B[165]), .A(n64), .Z(n32475) );
  XNOR U32901 ( .A(n32483), .B(n32697), .Z(n32476) );
  XNOR U32902 ( .A(n32482), .B(n32480), .Z(n32697) );
  AND U32903 ( .A(n32698), .B(n32699), .Z(n32480) );
  NANDN U32904 ( .A(n32700), .B(n32701), .Z(n32699) );
  OR U32905 ( .A(n32702), .B(n32703), .Z(n32701) );
  NAND U32906 ( .A(n32703), .B(n32702), .Z(n32698) );
  ANDN U32907 ( .B(B[166]), .A(n65), .Z(n32482) );
  XNOR U32908 ( .A(n32490), .B(n32704), .Z(n32483) );
  XNOR U32909 ( .A(n32489), .B(n32487), .Z(n32704) );
  AND U32910 ( .A(n32705), .B(n32706), .Z(n32487) );
  NANDN U32911 ( .A(n32707), .B(n32708), .Z(n32706) );
  NANDN U32912 ( .A(n32709), .B(n32710), .Z(n32708) );
  NANDN U32913 ( .A(n32710), .B(n32709), .Z(n32705) );
  ANDN U32914 ( .B(B[167]), .A(n66), .Z(n32489) );
  XNOR U32915 ( .A(n32497), .B(n32711), .Z(n32490) );
  XNOR U32916 ( .A(n32496), .B(n32494), .Z(n32711) );
  AND U32917 ( .A(n32712), .B(n32713), .Z(n32494) );
  NANDN U32918 ( .A(n32714), .B(n32715), .Z(n32713) );
  OR U32919 ( .A(n32716), .B(n32717), .Z(n32715) );
  NAND U32920 ( .A(n32717), .B(n32716), .Z(n32712) );
  ANDN U32921 ( .B(B[168]), .A(n67), .Z(n32496) );
  XNOR U32922 ( .A(n32504), .B(n32718), .Z(n32497) );
  XNOR U32923 ( .A(n32503), .B(n32501), .Z(n32718) );
  AND U32924 ( .A(n32719), .B(n32720), .Z(n32501) );
  NANDN U32925 ( .A(n32721), .B(n32722), .Z(n32720) );
  NANDN U32926 ( .A(n32723), .B(n32724), .Z(n32722) );
  NANDN U32927 ( .A(n32724), .B(n32723), .Z(n32719) );
  ANDN U32928 ( .B(B[169]), .A(n68), .Z(n32503) );
  XNOR U32929 ( .A(n32511), .B(n32725), .Z(n32504) );
  XNOR U32930 ( .A(n32510), .B(n32508), .Z(n32725) );
  AND U32931 ( .A(n32726), .B(n32727), .Z(n32508) );
  NANDN U32932 ( .A(n32728), .B(n32729), .Z(n32727) );
  OR U32933 ( .A(n32730), .B(n32731), .Z(n32729) );
  NAND U32934 ( .A(n32731), .B(n32730), .Z(n32726) );
  ANDN U32935 ( .B(B[170]), .A(n69), .Z(n32510) );
  XNOR U32936 ( .A(n32518), .B(n32732), .Z(n32511) );
  XNOR U32937 ( .A(n32517), .B(n32515), .Z(n32732) );
  AND U32938 ( .A(n32733), .B(n32734), .Z(n32515) );
  NANDN U32939 ( .A(n32735), .B(n32736), .Z(n32734) );
  NANDN U32940 ( .A(n32737), .B(n32738), .Z(n32736) );
  NANDN U32941 ( .A(n32738), .B(n32737), .Z(n32733) );
  ANDN U32942 ( .B(B[171]), .A(n70), .Z(n32517) );
  XNOR U32943 ( .A(n32525), .B(n32739), .Z(n32518) );
  XNOR U32944 ( .A(n32524), .B(n32522), .Z(n32739) );
  AND U32945 ( .A(n32740), .B(n32741), .Z(n32522) );
  NANDN U32946 ( .A(n32742), .B(n32743), .Z(n32741) );
  OR U32947 ( .A(n32744), .B(n32745), .Z(n32743) );
  NAND U32948 ( .A(n32745), .B(n32744), .Z(n32740) );
  ANDN U32949 ( .B(B[172]), .A(n71), .Z(n32524) );
  XNOR U32950 ( .A(n32532), .B(n32746), .Z(n32525) );
  XNOR U32951 ( .A(n32531), .B(n32529), .Z(n32746) );
  AND U32952 ( .A(n32747), .B(n32748), .Z(n32529) );
  NANDN U32953 ( .A(n32749), .B(n32750), .Z(n32748) );
  NANDN U32954 ( .A(n32751), .B(n32752), .Z(n32750) );
  NANDN U32955 ( .A(n32752), .B(n32751), .Z(n32747) );
  ANDN U32956 ( .B(B[173]), .A(n72), .Z(n32531) );
  XNOR U32957 ( .A(n32539), .B(n32753), .Z(n32532) );
  XNOR U32958 ( .A(n32538), .B(n32536), .Z(n32753) );
  AND U32959 ( .A(n32754), .B(n32755), .Z(n32536) );
  NANDN U32960 ( .A(n32756), .B(n32757), .Z(n32755) );
  OR U32961 ( .A(n32758), .B(n32759), .Z(n32757) );
  NAND U32962 ( .A(n32759), .B(n32758), .Z(n32754) );
  ANDN U32963 ( .B(B[174]), .A(n73), .Z(n32538) );
  XNOR U32964 ( .A(n32546), .B(n32760), .Z(n32539) );
  XNOR U32965 ( .A(n32545), .B(n32543), .Z(n32760) );
  AND U32966 ( .A(n32761), .B(n32762), .Z(n32543) );
  NANDN U32967 ( .A(n32763), .B(n32764), .Z(n32762) );
  NANDN U32968 ( .A(n32765), .B(n32766), .Z(n32764) );
  NANDN U32969 ( .A(n32766), .B(n32765), .Z(n32761) );
  ANDN U32970 ( .B(B[175]), .A(n74), .Z(n32545) );
  XNOR U32971 ( .A(n32553), .B(n32767), .Z(n32546) );
  XNOR U32972 ( .A(n32552), .B(n32550), .Z(n32767) );
  AND U32973 ( .A(n32768), .B(n32769), .Z(n32550) );
  NANDN U32974 ( .A(n32770), .B(n32771), .Z(n32769) );
  OR U32975 ( .A(n32772), .B(n32773), .Z(n32771) );
  NAND U32976 ( .A(n32773), .B(n32772), .Z(n32768) );
  ANDN U32977 ( .B(B[176]), .A(n75), .Z(n32552) );
  XNOR U32978 ( .A(n32560), .B(n32774), .Z(n32553) );
  XNOR U32979 ( .A(n32559), .B(n32557), .Z(n32774) );
  AND U32980 ( .A(n32775), .B(n32776), .Z(n32557) );
  NANDN U32981 ( .A(n32777), .B(n32778), .Z(n32776) );
  NANDN U32982 ( .A(n32779), .B(n32780), .Z(n32778) );
  NANDN U32983 ( .A(n32780), .B(n32779), .Z(n32775) );
  ANDN U32984 ( .B(B[177]), .A(n76), .Z(n32559) );
  XNOR U32985 ( .A(n32567), .B(n32781), .Z(n32560) );
  XNOR U32986 ( .A(n32566), .B(n32564), .Z(n32781) );
  AND U32987 ( .A(n32782), .B(n32783), .Z(n32564) );
  NANDN U32988 ( .A(n32784), .B(n32785), .Z(n32783) );
  OR U32989 ( .A(n32786), .B(n32787), .Z(n32785) );
  NAND U32990 ( .A(n32787), .B(n32786), .Z(n32782) );
  ANDN U32991 ( .B(B[178]), .A(n77), .Z(n32566) );
  XNOR U32992 ( .A(n32574), .B(n32788), .Z(n32567) );
  XNOR U32993 ( .A(n32573), .B(n32571), .Z(n32788) );
  AND U32994 ( .A(n32789), .B(n32790), .Z(n32571) );
  NANDN U32995 ( .A(n32791), .B(n32792), .Z(n32790) );
  NANDN U32996 ( .A(n32793), .B(n32794), .Z(n32792) );
  NANDN U32997 ( .A(n32794), .B(n32793), .Z(n32789) );
  ANDN U32998 ( .B(B[179]), .A(n78), .Z(n32573) );
  XNOR U32999 ( .A(n32581), .B(n32795), .Z(n32574) );
  XNOR U33000 ( .A(n32580), .B(n32578), .Z(n32795) );
  AND U33001 ( .A(n32796), .B(n32797), .Z(n32578) );
  NANDN U33002 ( .A(n32798), .B(n32799), .Z(n32797) );
  OR U33003 ( .A(n32800), .B(n32801), .Z(n32799) );
  NAND U33004 ( .A(n32801), .B(n32800), .Z(n32796) );
  ANDN U33005 ( .B(B[180]), .A(n79), .Z(n32580) );
  XNOR U33006 ( .A(n32588), .B(n32802), .Z(n32581) );
  XNOR U33007 ( .A(n32587), .B(n32585), .Z(n32802) );
  AND U33008 ( .A(n32803), .B(n32804), .Z(n32585) );
  NANDN U33009 ( .A(n32805), .B(n32806), .Z(n32804) );
  NANDN U33010 ( .A(n32807), .B(n32808), .Z(n32806) );
  NANDN U33011 ( .A(n32808), .B(n32807), .Z(n32803) );
  ANDN U33012 ( .B(B[181]), .A(n80), .Z(n32587) );
  XNOR U33013 ( .A(n32595), .B(n32809), .Z(n32588) );
  XNOR U33014 ( .A(n32594), .B(n32592), .Z(n32809) );
  AND U33015 ( .A(n32810), .B(n32811), .Z(n32592) );
  NANDN U33016 ( .A(n32812), .B(n32813), .Z(n32811) );
  OR U33017 ( .A(n32814), .B(n32815), .Z(n32813) );
  NAND U33018 ( .A(n32815), .B(n32814), .Z(n32810) );
  ANDN U33019 ( .B(B[182]), .A(n81), .Z(n32594) );
  XNOR U33020 ( .A(n32602), .B(n32816), .Z(n32595) );
  XNOR U33021 ( .A(n32601), .B(n32599), .Z(n32816) );
  AND U33022 ( .A(n32817), .B(n32818), .Z(n32599) );
  NANDN U33023 ( .A(n32819), .B(n32820), .Z(n32818) );
  NAND U33024 ( .A(n32821), .B(n32822), .Z(n32820) );
  ANDN U33025 ( .B(B[183]), .A(n82), .Z(n32601) );
  XOR U33026 ( .A(n32608), .B(n32823), .Z(n32602) );
  XNOR U33027 ( .A(n32606), .B(n32609), .Z(n32823) );
  NAND U33028 ( .A(A[2]), .B(B[184]), .Z(n32609) );
  NANDN U33029 ( .A(n32824), .B(n32825), .Z(n32606) );
  AND U33030 ( .A(A[0]), .B(B[185]), .Z(n32825) );
  XNOR U33031 ( .A(n32611), .B(n32826), .Z(n32608) );
  NAND U33032 ( .A(A[0]), .B(B[186]), .Z(n32826) );
  NAND U33033 ( .A(B[185]), .B(A[1]), .Z(n32611) );
  NAND U33034 ( .A(n32827), .B(n32828), .Z(n424) );
  NANDN U33035 ( .A(n32829), .B(n32830), .Z(n32828) );
  OR U33036 ( .A(n32831), .B(n32832), .Z(n32830) );
  NAND U33037 ( .A(n32832), .B(n32831), .Z(n32827) );
  XOR U33038 ( .A(n426), .B(n425), .Z(\A1[183] ) );
  XOR U33039 ( .A(n32832), .B(n32833), .Z(n425) );
  XNOR U33040 ( .A(n32831), .B(n32829), .Z(n32833) );
  AND U33041 ( .A(n32834), .B(n32835), .Z(n32829) );
  NANDN U33042 ( .A(n32836), .B(n32837), .Z(n32835) );
  NANDN U33043 ( .A(n32838), .B(n32839), .Z(n32837) );
  NANDN U33044 ( .A(n32839), .B(n32838), .Z(n32834) );
  ANDN U33045 ( .B(B[154]), .A(n54), .Z(n32831) );
  XNOR U33046 ( .A(n32626), .B(n32840), .Z(n32832) );
  XNOR U33047 ( .A(n32625), .B(n32623), .Z(n32840) );
  AND U33048 ( .A(n32841), .B(n32842), .Z(n32623) );
  NANDN U33049 ( .A(n32843), .B(n32844), .Z(n32842) );
  OR U33050 ( .A(n32845), .B(n32846), .Z(n32844) );
  NAND U33051 ( .A(n32846), .B(n32845), .Z(n32841) );
  ANDN U33052 ( .B(B[155]), .A(n55), .Z(n32625) );
  XNOR U33053 ( .A(n32633), .B(n32847), .Z(n32626) );
  XNOR U33054 ( .A(n32632), .B(n32630), .Z(n32847) );
  AND U33055 ( .A(n32848), .B(n32849), .Z(n32630) );
  NANDN U33056 ( .A(n32850), .B(n32851), .Z(n32849) );
  NANDN U33057 ( .A(n32852), .B(n32853), .Z(n32851) );
  NANDN U33058 ( .A(n32853), .B(n32852), .Z(n32848) );
  ANDN U33059 ( .B(B[156]), .A(n56), .Z(n32632) );
  XNOR U33060 ( .A(n32640), .B(n32854), .Z(n32633) );
  XNOR U33061 ( .A(n32639), .B(n32637), .Z(n32854) );
  AND U33062 ( .A(n32855), .B(n32856), .Z(n32637) );
  NANDN U33063 ( .A(n32857), .B(n32858), .Z(n32856) );
  OR U33064 ( .A(n32859), .B(n32860), .Z(n32858) );
  NAND U33065 ( .A(n32860), .B(n32859), .Z(n32855) );
  ANDN U33066 ( .B(B[157]), .A(n57), .Z(n32639) );
  XNOR U33067 ( .A(n32647), .B(n32861), .Z(n32640) );
  XNOR U33068 ( .A(n32646), .B(n32644), .Z(n32861) );
  AND U33069 ( .A(n32862), .B(n32863), .Z(n32644) );
  NANDN U33070 ( .A(n32864), .B(n32865), .Z(n32863) );
  NANDN U33071 ( .A(n32866), .B(n32867), .Z(n32865) );
  NANDN U33072 ( .A(n32867), .B(n32866), .Z(n32862) );
  ANDN U33073 ( .B(B[158]), .A(n58), .Z(n32646) );
  XNOR U33074 ( .A(n32654), .B(n32868), .Z(n32647) );
  XNOR U33075 ( .A(n32653), .B(n32651), .Z(n32868) );
  AND U33076 ( .A(n32869), .B(n32870), .Z(n32651) );
  NANDN U33077 ( .A(n32871), .B(n32872), .Z(n32870) );
  OR U33078 ( .A(n32873), .B(n32874), .Z(n32872) );
  NAND U33079 ( .A(n32874), .B(n32873), .Z(n32869) );
  ANDN U33080 ( .B(B[159]), .A(n59), .Z(n32653) );
  XNOR U33081 ( .A(n32661), .B(n32875), .Z(n32654) );
  XNOR U33082 ( .A(n32660), .B(n32658), .Z(n32875) );
  AND U33083 ( .A(n32876), .B(n32877), .Z(n32658) );
  NANDN U33084 ( .A(n32878), .B(n32879), .Z(n32877) );
  NANDN U33085 ( .A(n32880), .B(n32881), .Z(n32879) );
  NANDN U33086 ( .A(n32881), .B(n32880), .Z(n32876) );
  ANDN U33087 ( .B(B[160]), .A(n60), .Z(n32660) );
  XNOR U33088 ( .A(n32668), .B(n32882), .Z(n32661) );
  XNOR U33089 ( .A(n32667), .B(n32665), .Z(n32882) );
  AND U33090 ( .A(n32883), .B(n32884), .Z(n32665) );
  NANDN U33091 ( .A(n32885), .B(n32886), .Z(n32884) );
  OR U33092 ( .A(n32887), .B(n32888), .Z(n32886) );
  NAND U33093 ( .A(n32888), .B(n32887), .Z(n32883) );
  ANDN U33094 ( .B(B[161]), .A(n61), .Z(n32667) );
  XNOR U33095 ( .A(n32675), .B(n32889), .Z(n32668) );
  XNOR U33096 ( .A(n32674), .B(n32672), .Z(n32889) );
  AND U33097 ( .A(n32890), .B(n32891), .Z(n32672) );
  NANDN U33098 ( .A(n32892), .B(n32893), .Z(n32891) );
  NANDN U33099 ( .A(n32894), .B(n32895), .Z(n32893) );
  NANDN U33100 ( .A(n32895), .B(n32894), .Z(n32890) );
  ANDN U33101 ( .B(B[162]), .A(n62), .Z(n32674) );
  XNOR U33102 ( .A(n32682), .B(n32896), .Z(n32675) );
  XNOR U33103 ( .A(n32681), .B(n32679), .Z(n32896) );
  AND U33104 ( .A(n32897), .B(n32898), .Z(n32679) );
  NANDN U33105 ( .A(n32899), .B(n32900), .Z(n32898) );
  OR U33106 ( .A(n32901), .B(n32902), .Z(n32900) );
  NAND U33107 ( .A(n32902), .B(n32901), .Z(n32897) );
  ANDN U33108 ( .B(B[163]), .A(n63), .Z(n32681) );
  XNOR U33109 ( .A(n32689), .B(n32903), .Z(n32682) );
  XNOR U33110 ( .A(n32688), .B(n32686), .Z(n32903) );
  AND U33111 ( .A(n32904), .B(n32905), .Z(n32686) );
  NANDN U33112 ( .A(n32906), .B(n32907), .Z(n32905) );
  NANDN U33113 ( .A(n32908), .B(n32909), .Z(n32907) );
  NANDN U33114 ( .A(n32909), .B(n32908), .Z(n32904) );
  ANDN U33115 ( .B(B[164]), .A(n64), .Z(n32688) );
  XNOR U33116 ( .A(n32696), .B(n32910), .Z(n32689) );
  XNOR U33117 ( .A(n32695), .B(n32693), .Z(n32910) );
  AND U33118 ( .A(n32911), .B(n32912), .Z(n32693) );
  NANDN U33119 ( .A(n32913), .B(n32914), .Z(n32912) );
  OR U33120 ( .A(n32915), .B(n32916), .Z(n32914) );
  NAND U33121 ( .A(n32916), .B(n32915), .Z(n32911) );
  ANDN U33122 ( .B(B[165]), .A(n65), .Z(n32695) );
  XNOR U33123 ( .A(n32703), .B(n32917), .Z(n32696) );
  XNOR U33124 ( .A(n32702), .B(n32700), .Z(n32917) );
  AND U33125 ( .A(n32918), .B(n32919), .Z(n32700) );
  NANDN U33126 ( .A(n32920), .B(n32921), .Z(n32919) );
  NANDN U33127 ( .A(n32922), .B(n32923), .Z(n32921) );
  NANDN U33128 ( .A(n32923), .B(n32922), .Z(n32918) );
  ANDN U33129 ( .B(B[166]), .A(n66), .Z(n32702) );
  XNOR U33130 ( .A(n32710), .B(n32924), .Z(n32703) );
  XNOR U33131 ( .A(n32709), .B(n32707), .Z(n32924) );
  AND U33132 ( .A(n32925), .B(n32926), .Z(n32707) );
  NANDN U33133 ( .A(n32927), .B(n32928), .Z(n32926) );
  OR U33134 ( .A(n32929), .B(n32930), .Z(n32928) );
  NAND U33135 ( .A(n32930), .B(n32929), .Z(n32925) );
  ANDN U33136 ( .B(B[167]), .A(n67), .Z(n32709) );
  XNOR U33137 ( .A(n32717), .B(n32931), .Z(n32710) );
  XNOR U33138 ( .A(n32716), .B(n32714), .Z(n32931) );
  AND U33139 ( .A(n32932), .B(n32933), .Z(n32714) );
  NANDN U33140 ( .A(n32934), .B(n32935), .Z(n32933) );
  NANDN U33141 ( .A(n32936), .B(n32937), .Z(n32935) );
  NANDN U33142 ( .A(n32937), .B(n32936), .Z(n32932) );
  ANDN U33143 ( .B(B[168]), .A(n68), .Z(n32716) );
  XNOR U33144 ( .A(n32724), .B(n32938), .Z(n32717) );
  XNOR U33145 ( .A(n32723), .B(n32721), .Z(n32938) );
  AND U33146 ( .A(n32939), .B(n32940), .Z(n32721) );
  NANDN U33147 ( .A(n32941), .B(n32942), .Z(n32940) );
  OR U33148 ( .A(n32943), .B(n32944), .Z(n32942) );
  NAND U33149 ( .A(n32944), .B(n32943), .Z(n32939) );
  ANDN U33150 ( .B(B[169]), .A(n69), .Z(n32723) );
  XNOR U33151 ( .A(n32731), .B(n32945), .Z(n32724) );
  XNOR U33152 ( .A(n32730), .B(n32728), .Z(n32945) );
  AND U33153 ( .A(n32946), .B(n32947), .Z(n32728) );
  NANDN U33154 ( .A(n32948), .B(n32949), .Z(n32947) );
  NANDN U33155 ( .A(n32950), .B(n32951), .Z(n32949) );
  NANDN U33156 ( .A(n32951), .B(n32950), .Z(n32946) );
  ANDN U33157 ( .B(B[170]), .A(n70), .Z(n32730) );
  XNOR U33158 ( .A(n32738), .B(n32952), .Z(n32731) );
  XNOR U33159 ( .A(n32737), .B(n32735), .Z(n32952) );
  AND U33160 ( .A(n32953), .B(n32954), .Z(n32735) );
  NANDN U33161 ( .A(n32955), .B(n32956), .Z(n32954) );
  OR U33162 ( .A(n32957), .B(n32958), .Z(n32956) );
  NAND U33163 ( .A(n32958), .B(n32957), .Z(n32953) );
  ANDN U33164 ( .B(B[171]), .A(n71), .Z(n32737) );
  XNOR U33165 ( .A(n32745), .B(n32959), .Z(n32738) );
  XNOR U33166 ( .A(n32744), .B(n32742), .Z(n32959) );
  AND U33167 ( .A(n32960), .B(n32961), .Z(n32742) );
  NANDN U33168 ( .A(n32962), .B(n32963), .Z(n32961) );
  NANDN U33169 ( .A(n32964), .B(n32965), .Z(n32963) );
  NANDN U33170 ( .A(n32965), .B(n32964), .Z(n32960) );
  ANDN U33171 ( .B(B[172]), .A(n72), .Z(n32744) );
  XNOR U33172 ( .A(n32752), .B(n32966), .Z(n32745) );
  XNOR U33173 ( .A(n32751), .B(n32749), .Z(n32966) );
  AND U33174 ( .A(n32967), .B(n32968), .Z(n32749) );
  NANDN U33175 ( .A(n32969), .B(n32970), .Z(n32968) );
  OR U33176 ( .A(n32971), .B(n32972), .Z(n32970) );
  NAND U33177 ( .A(n32972), .B(n32971), .Z(n32967) );
  ANDN U33178 ( .B(B[173]), .A(n73), .Z(n32751) );
  XNOR U33179 ( .A(n32759), .B(n32973), .Z(n32752) );
  XNOR U33180 ( .A(n32758), .B(n32756), .Z(n32973) );
  AND U33181 ( .A(n32974), .B(n32975), .Z(n32756) );
  NANDN U33182 ( .A(n32976), .B(n32977), .Z(n32975) );
  NANDN U33183 ( .A(n32978), .B(n32979), .Z(n32977) );
  NANDN U33184 ( .A(n32979), .B(n32978), .Z(n32974) );
  ANDN U33185 ( .B(B[174]), .A(n74), .Z(n32758) );
  XNOR U33186 ( .A(n32766), .B(n32980), .Z(n32759) );
  XNOR U33187 ( .A(n32765), .B(n32763), .Z(n32980) );
  AND U33188 ( .A(n32981), .B(n32982), .Z(n32763) );
  NANDN U33189 ( .A(n32983), .B(n32984), .Z(n32982) );
  OR U33190 ( .A(n32985), .B(n32986), .Z(n32984) );
  NAND U33191 ( .A(n32986), .B(n32985), .Z(n32981) );
  ANDN U33192 ( .B(B[175]), .A(n75), .Z(n32765) );
  XNOR U33193 ( .A(n32773), .B(n32987), .Z(n32766) );
  XNOR U33194 ( .A(n32772), .B(n32770), .Z(n32987) );
  AND U33195 ( .A(n32988), .B(n32989), .Z(n32770) );
  NANDN U33196 ( .A(n32990), .B(n32991), .Z(n32989) );
  NANDN U33197 ( .A(n32992), .B(n32993), .Z(n32991) );
  NANDN U33198 ( .A(n32993), .B(n32992), .Z(n32988) );
  ANDN U33199 ( .B(B[176]), .A(n76), .Z(n32772) );
  XNOR U33200 ( .A(n32780), .B(n32994), .Z(n32773) );
  XNOR U33201 ( .A(n32779), .B(n32777), .Z(n32994) );
  AND U33202 ( .A(n32995), .B(n32996), .Z(n32777) );
  NANDN U33203 ( .A(n32997), .B(n32998), .Z(n32996) );
  OR U33204 ( .A(n32999), .B(n33000), .Z(n32998) );
  NAND U33205 ( .A(n33000), .B(n32999), .Z(n32995) );
  ANDN U33206 ( .B(B[177]), .A(n77), .Z(n32779) );
  XNOR U33207 ( .A(n32787), .B(n33001), .Z(n32780) );
  XNOR U33208 ( .A(n32786), .B(n32784), .Z(n33001) );
  AND U33209 ( .A(n33002), .B(n33003), .Z(n32784) );
  NANDN U33210 ( .A(n33004), .B(n33005), .Z(n33003) );
  NANDN U33211 ( .A(n33006), .B(n33007), .Z(n33005) );
  NANDN U33212 ( .A(n33007), .B(n33006), .Z(n33002) );
  ANDN U33213 ( .B(B[178]), .A(n78), .Z(n32786) );
  XNOR U33214 ( .A(n32794), .B(n33008), .Z(n32787) );
  XNOR U33215 ( .A(n32793), .B(n32791), .Z(n33008) );
  AND U33216 ( .A(n33009), .B(n33010), .Z(n32791) );
  NANDN U33217 ( .A(n33011), .B(n33012), .Z(n33010) );
  OR U33218 ( .A(n33013), .B(n33014), .Z(n33012) );
  NAND U33219 ( .A(n33014), .B(n33013), .Z(n33009) );
  ANDN U33220 ( .B(B[179]), .A(n79), .Z(n32793) );
  XNOR U33221 ( .A(n32801), .B(n33015), .Z(n32794) );
  XNOR U33222 ( .A(n32800), .B(n32798), .Z(n33015) );
  AND U33223 ( .A(n33016), .B(n33017), .Z(n32798) );
  NANDN U33224 ( .A(n33018), .B(n33019), .Z(n33017) );
  NANDN U33225 ( .A(n33020), .B(n33021), .Z(n33019) );
  NANDN U33226 ( .A(n33021), .B(n33020), .Z(n33016) );
  ANDN U33227 ( .B(B[180]), .A(n80), .Z(n32800) );
  XNOR U33228 ( .A(n32808), .B(n33022), .Z(n32801) );
  XNOR U33229 ( .A(n32807), .B(n32805), .Z(n33022) );
  AND U33230 ( .A(n33023), .B(n33024), .Z(n32805) );
  NANDN U33231 ( .A(n33025), .B(n33026), .Z(n33024) );
  OR U33232 ( .A(n33027), .B(n33028), .Z(n33026) );
  NAND U33233 ( .A(n33028), .B(n33027), .Z(n33023) );
  ANDN U33234 ( .B(B[181]), .A(n81), .Z(n32807) );
  XNOR U33235 ( .A(n32815), .B(n33029), .Z(n32808) );
  XNOR U33236 ( .A(n32814), .B(n32812), .Z(n33029) );
  AND U33237 ( .A(n33030), .B(n33031), .Z(n32812) );
  NANDN U33238 ( .A(n33032), .B(n33033), .Z(n33031) );
  NAND U33239 ( .A(n33034), .B(n33035), .Z(n33033) );
  ANDN U33240 ( .B(B[182]), .A(n82), .Z(n32814) );
  XOR U33241 ( .A(n32821), .B(n33036), .Z(n32815) );
  XNOR U33242 ( .A(n32819), .B(n32822), .Z(n33036) );
  NAND U33243 ( .A(A[2]), .B(B[183]), .Z(n32822) );
  NANDN U33244 ( .A(n33037), .B(n33038), .Z(n32819) );
  AND U33245 ( .A(A[0]), .B(B[184]), .Z(n33038) );
  XNOR U33246 ( .A(n32824), .B(n33039), .Z(n32821) );
  NAND U33247 ( .A(A[0]), .B(B[185]), .Z(n33039) );
  NAND U33248 ( .A(B[184]), .B(A[1]), .Z(n32824) );
  NAND U33249 ( .A(n33040), .B(n33041), .Z(n426) );
  NANDN U33250 ( .A(n33042), .B(n33043), .Z(n33041) );
  OR U33251 ( .A(n33044), .B(n33045), .Z(n33043) );
  NAND U33252 ( .A(n33045), .B(n33044), .Z(n33040) );
  XOR U33253 ( .A(n428), .B(n427), .Z(\A1[182] ) );
  XOR U33254 ( .A(n33045), .B(n33046), .Z(n427) );
  XNOR U33255 ( .A(n33044), .B(n33042), .Z(n33046) );
  AND U33256 ( .A(n33047), .B(n33048), .Z(n33042) );
  NANDN U33257 ( .A(n33049), .B(n33050), .Z(n33048) );
  NANDN U33258 ( .A(n33051), .B(n33052), .Z(n33050) );
  NANDN U33259 ( .A(n33052), .B(n33051), .Z(n33047) );
  ANDN U33260 ( .B(B[153]), .A(n54), .Z(n33044) );
  XNOR U33261 ( .A(n32839), .B(n33053), .Z(n33045) );
  XNOR U33262 ( .A(n32838), .B(n32836), .Z(n33053) );
  AND U33263 ( .A(n33054), .B(n33055), .Z(n32836) );
  NANDN U33264 ( .A(n33056), .B(n33057), .Z(n33055) );
  OR U33265 ( .A(n33058), .B(n33059), .Z(n33057) );
  NAND U33266 ( .A(n33059), .B(n33058), .Z(n33054) );
  ANDN U33267 ( .B(B[154]), .A(n55), .Z(n32838) );
  XNOR U33268 ( .A(n32846), .B(n33060), .Z(n32839) );
  XNOR U33269 ( .A(n32845), .B(n32843), .Z(n33060) );
  AND U33270 ( .A(n33061), .B(n33062), .Z(n32843) );
  NANDN U33271 ( .A(n33063), .B(n33064), .Z(n33062) );
  NANDN U33272 ( .A(n33065), .B(n33066), .Z(n33064) );
  NANDN U33273 ( .A(n33066), .B(n33065), .Z(n33061) );
  ANDN U33274 ( .B(B[155]), .A(n56), .Z(n32845) );
  XNOR U33275 ( .A(n32853), .B(n33067), .Z(n32846) );
  XNOR U33276 ( .A(n32852), .B(n32850), .Z(n33067) );
  AND U33277 ( .A(n33068), .B(n33069), .Z(n32850) );
  NANDN U33278 ( .A(n33070), .B(n33071), .Z(n33069) );
  OR U33279 ( .A(n33072), .B(n33073), .Z(n33071) );
  NAND U33280 ( .A(n33073), .B(n33072), .Z(n33068) );
  ANDN U33281 ( .B(B[156]), .A(n57), .Z(n32852) );
  XNOR U33282 ( .A(n32860), .B(n33074), .Z(n32853) );
  XNOR U33283 ( .A(n32859), .B(n32857), .Z(n33074) );
  AND U33284 ( .A(n33075), .B(n33076), .Z(n32857) );
  NANDN U33285 ( .A(n33077), .B(n33078), .Z(n33076) );
  NANDN U33286 ( .A(n33079), .B(n33080), .Z(n33078) );
  NANDN U33287 ( .A(n33080), .B(n33079), .Z(n33075) );
  ANDN U33288 ( .B(B[157]), .A(n58), .Z(n32859) );
  XNOR U33289 ( .A(n32867), .B(n33081), .Z(n32860) );
  XNOR U33290 ( .A(n32866), .B(n32864), .Z(n33081) );
  AND U33291 ( .A(n33082), .B(n33083), .Z(n32864) );
  NANDN U33292 ( .A(n33084), .B(n33085), .Z(n33083) );
  OR U33293 ( .A(n33086), .B(n33087), .Z(n33085) );
  NAND U33294 ( .A(n33087), .B(n33086), .Z(n33082) );
  ANDN U33295 ( .B(B[158]), .A(n59), .Z(n32866) );
  XNOR U33296 ( .A(n32874), .B(n33088), .Z(n32867) );
  XNOR U33297 ( .A(n32873), .B(n32871), .Z(n33088) );
  AND U33298 ( .A(n33089), .B(n33090), .Z(n32871) );
  NANDN U33299 ( .A(n33091), .B(n33092), .Z(n33090) );
  NANDN U33300 ( .A(n33093), .B(n33094), .Z(n33092) );
  NANDN U33301 ( .A(n33094), .B(n33093), .Z(n33089) );
  ANDN U33302 ( .B(B[159]), .A(n60), .Z(n32873) );
  XNOR U33303 ( .A(n32881), .B(n33095), .Z(n32874) );
  XNOR U33304 ( .A(n32880), .B(n32878), .Z(n33095) );
  AND U33305 ( .A(n33096), .B(n33097), .Z(n32878) );
  NANDN U33306 ( .A(n33098), .B(n33099), .Z(n33097) );
  OR U33307 ( .A(n33100), .B(n33101), .Z(n33099) );
  NAND U33308 ( .A(n33101), .B(n33100), .Z(n33096) );
  ANDN U33309 ( .B(B[160]), .A(n61), .Z(n32880) );
  XNOR U33310 ( .A(n32888), .B(n33102), .Z(n32881) );
  XNOR U33311 ( .A(n32887), .B(n32885), .Z(n33102) );
  AND U33312 ( .A(n33103), .B(n33104), .Z(n32885) );
  NANDN U33313 ( .A(n33105), .B(n33106), .Z(n33104) );
  NANDN U33314 ( .A(n33107), .B(n33108), .Z(n33106) );
  NANDN U33315 ( .A(n33108), .B(n33107), .Z(n33103) );
  ANDN U33316 ( .B(B[161]), .A(n62), .Z(n32887) );
  XNOR U33317 ( .A(n32895), .B(n33109), .Z(n32888) );
  XNOR U33318 ( .A(n32894), .B(n32892), .Z(n33109) );
  AND U33319 ( .A(n33110), .B(n33111), .Z(n32892) );
  NANDN U33320 ( .A(n33112), .B(n33113), .Z(n33111) );
  OR U33321 ( .A(n33114), .B(n33115), .Z(n33113) );
  NAND U33322 ( .A(n33115), .B(n33114), .Z(n33110) );
  ANDN U33323 ( .B(B[162]), .A(n63), .Z(n32894) );
  XNOR U33324 ( .A(n32902), .B(n33116), .Z(n32895) );
  XNOR U33325 ( .A(n32901), .B(n32899), .Z(n33116) );
  AND U33326 ( .A(n33117), .B(n33118), .Z(n32899) );
  NANDN U33327 ( .A(n33119), .B(n33120), .Z(n33118) );
  NANDN U33328 ( .A(n33121), .B(n33122), .Z(n33120) );
  NANDN U33329 ( .A(n33122), .B(n33121), .Z(n33117) );
  ANDN U33330 ( .B(B[163]), .A(n64), .Z(n32901) );
  XNOR U33331 ( .A(n32909), .B(n33123), .Z(n32902) );
  XNOR U33332 ( .A(n32908), .B(n32906), .Z(n33123) );
  AND U33333 ( .A(n33124), .B(n33125), .Z(n32906) );
  NANDN U33334 ( .A(n33126), .B(n33127), .Z(n33125) );
  OR U33335 ( .A(n33128), .B(n33129), .Z(n33127) );
  NAND U33336 ( .A(n33129), .B(n33128), .Z(n33124) );
  ANDN U33337 ( .B(B[164]), .A(n65), .Z(n32908) );
  XNOR U33338 ( .A(n32916), .B(n33130), .Z(n32909) );
  XNOR U33339 ( .A(n32915), .B(n32913), .Z(n33130) );
  AND U33340 ( .A(n33131), .B(n33132), .Z(n32913) );
  NANDN U33341 ( .A(n33133), .B(n33134), .Z(n33132) );
  NANDN U33342 ( .A(n33135), .B(n33136), .Z(n33134) );
  NANDN U33343 ( .A(n33136), .B(n33135), .Z(n33131) );
  ANDN U33344 ( .B(B[165]), .A(n66), .Z(n32915) );
  XNOR U33345 ( .A(n32923), .B(n33137), .Z(n32916) );
  XNOR U33346 ( .A(n32922), .B(n32920), .Z(n33137) );
  AND U33347 ( .A(n33138), .B(n33139), .Z(n32920) );
  NANDN U33348 ( .A(n33140), .B(n33141), .Z(n33139) );
  OR U33349 ( .A(n33142), .B(n33143), .Z(n33141) );
  NAND U33350 ( .A(n33143), .B(n33142), .Z(n33138) );
  ANDN U33351 ( .B(B[166]), .A(n67), .Z(n32922) );
  XNOR U33352 ( .A(n32930), .B(n33144), .Z(n32923) );
  XNOR U33353 ( .A(n32929), .B(n32927), .Z(n33144) );
  AND U33354 ( .A(n33145), .B(n33146), .Z(n32927) );
  NANDN U33355 ( .A(n33147), .B(n33148), .Z(n33146) );
  NANDN U33356 ( .A(n33149), .B(n33150), .Z(n33148) );
  NANDN U33357 ( .A(n33150), .B(n33149), .Z(n33145) );
  ANDN U33358 ( .B(B[167]), .A(n68), .Z(n32929) );
  XNOR U33359 ( .A(n32937), .B(n33151), .Z(n32930) );
  XNOR U33360 ( .A(n32936), .B(n32934), .Z(n33151) );
  AND U33361 ( .A(n33152), .B(n33153), .Z(n32934) );
  NANDN U33362 ( .A(n33154), .B(n33155), .Z(n33153) );
  OR U33363 ( .A(n33156), .B(n33157), .Z(n33155) );
  NAND U33364 ( .A(n33157), .B(n33156), .Z(n33152) );
  ANDN U33365 ( .B(B[168]), .A(n69), .Z(n32936) );
  XNOR U33366 ( .A(n32944), .B(n33158), .Z(n32937) );
  XNOR U33367 ( .A(n32943), .B(n32941), .Z(n33158) );
  AND U33368 ( .A(n33159), .B(n33160), .Z(n32941) );
  NANDN U33369 ( .A(n33161), .B(n33162), .Z(n33160) );
  NANDN U33370 ( .A(n33163), .B(n33164), .Z(n33162) );
  NANDN U33371 ( .A(n33164), .B(n33163), .Z(n33159) );
  ANDN U33372 ( .B(B[169]), .A(n70), .Z(n32943) );
  XNOR U33373 ( .A(n32951), .B(n33165), .Z(n32944) );
  XNOR U33374 ( .A(n32950), .B(n32948), .Z(n33165) );
  AND U33375 ( .A(n33166), .B(n33167), .Z(n32948) );
  NANDN U33376 ( .A(n33168), .B(n33169), .Z(n33167) );
  OR U33377 ( .A(n33170), .B(n33171), .Z(n33169) );
  NAND U33378 ( .A(n33171), .B(n33170), .Z(n33166) );
  ANDN U33379 ( .B(B[170]), .A(n71), .Z(n32950) );
  XNOR U33380 ( .A(n32958), .B(n33172), .Z(n32951) );
  XNOR U33381 ( .A(n32957), .B(n32955), .Z(n33172) );
  AND U33382 ( .A(n33173), .B(n33174), .Z(n32955) );
  NANDN U33383 ( .A(n33175), .B(n33176), .Z(n33174) );
  NANDN U33384 ( .A(n33177), .B(n33178), .Z(n33176) );
  NANDN U33385 ( .A(n33178), .B(n33177), .Z(n33173) );
  ANDN U33386 ( .B(B[171]), .A(n72), .Z(n32957) );
  XNOR U33387 ( .A(n32965), .B(n33179), .Z(n32958) );
  XNOR U33388 ( .A(n32964), .B(n32962), .Z(n33179) );
  AND U33389 ( .A(n33180), .B(n33181), .Z(n32962) );
  NANDN U33390 ( .A(n33182), .B(n33183), .Z(n33181) );
  OR U33391 ( .A(n33184), .B(n33185), .Z(n33183) );
  NAND U33392 ( .A(n33185), .B(n33184), .Z(n33180) );
  ANDN U33393 ( .B(B[172]), .A(n73), .Z(n32964) );
  XNOR U33394 ( .A(n32972), .B(n33186), .Z(n32965) );
  XNOR U33395 ( .A(n32971), .B(n32969), .Z(n33186) );
  AND U33396 ( .A(n33187), .B(n33188), .Z(n32969) );
  NANDN U33397 ( .A(n33189), .B(n33190), .Z(n33188) );
  NANDN U33398 ( .A(n33191), .B(n33192), .Z(n33190) );
  NANDN U33399 ( .A(n33192), .B(n33191), .Z(n33187) );
  ANDN U33400 ( .B(B[173]), .A(n74), .Z(n32971) );
  XNOR U33401 ( .A(n32979), .B(n33193), .Z(n32972) );
  XNOR U33402 ( .A(n32978), .B(n32976), .Z(n33193) );
  AND U33403 ( .A(n33194), .B(n33195), .Z(n32976) );
  NANDN U33404 ( .A(n33196), .B(n33197), .Z(n33195) );
  OR U33405 ( .A(n33198), .B(n33199), .Z(n33197) );
  NAND U33406 ( .A(n33199), .B(n33198), .Z(n33194) );
  ANDN U33407 ( .B(B[174]), .A(n75), .Z(n32978) );
  XNOR U33408 ( .A(n32986), .B(n33200), .Z(n32979) );
  XNOR U33409 ( .A(n32985), .B(n32983), .Z(n33200) );
  AND U33410 ( .A(n33201), .B(n33202), .Z(n32983) );
  NANDN U33411 ( .A(n33203), .B(n33204), .Z(n33202) );
  NANDN U33412 ( .A(n33205), .B(n33206), .Z(n33204) );
  NANDN U33413 ( .A(n33206), .B(n33205), .Z(n33201) );
  ANDN U33414 ( .B(B[175]), .A(n76), .Z(n32985) );
  XNOR U33415 ( .A(n32993), .B(n33207), .Z(n32986) );
  XNOR U33416 ( .A(n32992), .B(n32990), .Z(n33207) );
  AND U33417 ( .A(n33208), .B(n33209), .Z(n32990) );
  NANDN U33418 ( .A(n33210), .B(n33211), .Z(n33209) );
  OR U33419 ( .A(n33212), .B(n33213), .Z(n33211) );
  NAND U33420 ( .A(n33213), .B(n33212), .Z(n33208) );
  ANDN U33421 ( .B(B[176]), .A(n77), .Z(n32992) );
  XNOR U33422 ( .A(n33000), .B(n33214), .Z(n32993) );
  XNOR U33423 ( .A(n32999), .B(n32997), .Z(n33214) );
  AND U33424 ( .A(n33215), .B(n33216), .Z(n32997) );
  NANDN U33425 ( .A(n33217), .B(n33218), .Z(n33216) );
  NANDN U33426 ( .A(n33219), .B(n33220), .Z(n33218) );
  NANDN U33427 ( .A(n33220), .B(n33219), .Z(n33215) );
  ANDN U33428 ( .B(B[177]), .A(n78), .Z(n32999) );
  XNOR U33429 ( .A(n33007), .B(n33221), .Z(n33000) );
  XNOR U33430 ( .A(n33006), .B(n33004), .Z(n33221) );
  AND U33431 ( .A(n33222), .B(n33223), .Z(n33004) );
  NANDN U33432 ( .A(n33224), .B(n33225), .Z(n33223) );
  OR U33433 ( .A(n33226), .B(n33227), .Z(n33225) );
  NAND U33434 ( .A(n33227), .B(n33226), .Z(n33222) );
  ANDN U33435 ( .B(B[178]), .A(n79), .Z(n33006) );
  XNOR U33436 ( .A(n33014), .B(n33228), .Z(n33007) );
  XNOR U33437 ( .A(n33013), .B(n33011), .Z(n33228) );
  AND U33438 ( .A(n33229), .B(n33230), .Z(n33011) );
  NANDN U33439 ( .A(n33231), .B(n33232), .Z(n33230) );
  NANDN U33440 ( .A(n33233), .B(n33234), .Z(n33232) );
  NANDN U33441 ( .A(n33234), .B(n33233), .Z(n33229) );
  ANDN U33442 ( .B(B[179]), .A(n80), .Z(n33013) );
  XNOR U33443 ( .A(n33021), .B(n33235), .Z(n33014) );
  XNOR U33444 ( .A(n33020), .B(n33018), .Z(n33235) );
  AND U33445 ( .A(n33236), .B(n33237), .Z(n33018) );
  NANDN U33446 ( .A(n33238), .B(n33239), .Z(n33237) );
  OR U33447 ( .A(n33240), .B(n33241), .Z(n33239) );
  NAND U33448 ( .A(n33241), .B(n33240), .Z(n33236) );
  ANDN U33449 ( .B(B[180]), .A(n81), .Z(n33020) );
  XNOR U33450 ( .A(n33028), .B(n33242), .Z(n33021) );
  XNOR U33451 ( .A(n33027), .B(n33025), .Z(n33242) );
  AND U33452 ( .A(n33243), .B(n33244), .Z(n33025) );
  NANDN U33453 ( .A(n33245), .B(n33246), .Z(n33244) );
  NAND U33454 ( .A(n33247), .B(n33248), .Z(n33246) );
  ANDN U33455 ( .B(B[181]), .A(n82), .Z(n33027) );
  XOR U33456 ( .A(n33034), .B(n33249), .Z(n33028) );
  XNOR U33457 ( .A(n33032), .B(n33035), .Z(n33249) );
  NAND U33458 ( .A(A[2]), .B(B[182]), .Z(n33035) );
  NANDN U33459 ( .A(n33250), .B(n33251), .Z(n33032) );
  AND U33460 ( .A(A[0]), .B(B[183]), .Z(n33251) );
  XNOR U33461 ( .A(n33037), .B(n33252), .Z(n33034) );
  NAND U33462 ( .A(A[0]), .B(B[184]), .Z(n33252) );
  NAND U33463 ( .A(B[183]), .B(A[1]), .Z(n33037) );
  NAND U33464 ( .A(n33253), .B(n33254), .Z(n428) );
  NANDN U33465 ( .A(n33255), .B(n33256), .Z(n33254) );
  OR U33466 ( .A(n33257), .B(n33258), .Z(n33256) );
  NAND U33467 ( .A(n33258), .B(n33257), .Z(n33253) );
  XOR U33468 ( .A(n430), .B(n429), .Z(\A1[181] ) );
  XOR U33469 ( .A(n33258), .B(n33259), .Z(n429) );
  XNOR U33470 ( .A(n33257), .B(n33255), .Z(n33259) );
  AND U33471 ( .A(n33260), .B(n33261), .Z(n33255) );
  NANDN U33472 ( .A(n33262), .B(n33263), .Z(n33261) );
  NANDN U33473 ( .A(n33264), .B(n33265), .Z(n33263) );
  NANDN U33474 ( .A(n33265), .B(n33264), .Z(n33260) );
  ANDN U33475 ( .B(B[152]), .A(n54), .Z(n33257) );
  XNOR U33476 ( .A(n33052), .B(n33266), .Z(n33258) );
  XNOR U33477 ( .A(n33051), .B(n33049), .Z(n33266) );
  AND U33478 ( .A(n33267), .B(n33268), .Z(n33049) );
  NANDN U33479 ( .A(n33269), .B(n33270), .Z(n33268) );
  OR U33480 ( .A(n33271), .B(n33272), .Z(n33270) );
  NAND U33481 ( .A(n33272), .B(n33271), .Z(n33267) );
  ANDN U33482 ( .B(B[153]), .A(n55), .Z(n33051) );
  XNOR U33483 ( .A(n33059), .B(n33273), .Z(n33052) );
  XNOR U33484 ( .A(n33058), .B(n33056), .Z(n33273) );
  AND U33485 ( .A(n33274), .B(n33275), .Z(n33056) );
  NANDN U33486 ( .A(n33276), .B(n33277), .Z(n33275) );
  NANDN U33487 ( .A(n33278), .B(n33279), .Z(n33277) );
  NANDN U33488 ( .A(n33279), .B(n33278), .Z(n33274) );
  ANDN U33489 ( .B(B[154]), .A(n56), .Z(n33058) );
  XNOR U33490 ( .A(n33066), .B(n33280), .Z(n33059) );
  XNOR U33491 ( .A(n33065), .B(n33063), .Z(n33280) );
  AND U33492 ( .A(n33281), .B(n33282), .Z(n33063) );
  NANDN U33493 ( .A(n33283), .B(n33284), .Z(n33282) );
  OR U33494 ( .A(n33285), .B(n33286), .Z(n33284) );
  NAND U33495 ( .A(n33286), .B(n33285), .Z(n33281) );
  ANDN U33496 ( .B(B[155]), .A(n57), .Z(n33065) );
  XNOR U33497 ( .A(n33073), .B(n33287), .Z(n33066) );
  XNOR U33498 ( .A(n33072), .B(n33070), .Z(n33287) );
  AND U33499 ( .A(n33288), .B(n33289), .Z(n33070) );
  NANDN U33500 ( .A(n33290), .B(n33291), .Z(n33289) );
  NANDN U33501 ( .A(n33292), .B(n33293), .Z(n33291) );
  NANDN U33502 ( .A(n33293), .B(n33292), .Z(n33288) );
  ANDN U33503 ( .B(B[156]), .A(n58), .Z(n33072) );
  XNOR U33504 ( .A(n33080), .B(n33294), .Z(n33073) );
  XNOR U33505 ( .A(n33079), .B(n33077), .Z(n33294) );
  AND U33506 ( .A(n33295), .B(n33296), .Z(n33077) );
  NANDN U33507 ( .A(n33297), .B(n33298), .Z(n33296) );
  OR U33508 ( .A(n33299), .B(n33300), .Z(n33298) );
  NAND U33509 ( .A(n33300), .B(n33299), .Z(n33295) );
  ANDN U33510 ( .B(B[157]), .A(n59), .Z(n33079) );
  XNOR U33511 ( .A(n33087), .B(n33301), .Z(n33080) );
  XNOR U33512 ( .A(n33086), .B(n33084), .Z(n33301) );
  AND U33513 ( .A(n33302), .B(n33303), .Z(n33084) );
  NANDN U33514 ( .A(n33304), .B(n33305), .Z(n33303) );
  NANDN U33515 ( .A(n33306), .B(n33307), .Z(n33305) );
  NANDN U33516 ( .A(n33307), .B(n33306), .Z(n33302) );
  ANDN U33517 ( .B(B[158]), .A(n60), .Z(n33086) );
  XNOR U33518 ( .A(n33094), .B(n33308), .Z(n33087) );
  XNOR U33519 ( .A(n33093), .B(n33091), .Z(n33308) );
  AND U33520 ( .A(n33309), .B(n33310), .Z(n33091) );
  NANDN U33521 ( .A(n33311), .B(n33312), .Z(n33310) );
  OR U33522 ( .A(n33313), .B(n33314), .Z(n33312) );
  NAND U33523 ( .A(n33314), .B(n33313), .Z(n33309) );
  ANDN U33524 ( .B(B[159]), .A(n61), .Z(n33093) );
  XNOR U33525 ( .A(n33101), .B(n33315), .Z(n33094) );
  XNOR U33526 ( .A(n33100), .B(n33098), .Z(n33315) );
  AND U33527 ( .A(n33316), .B(n33317), .Z(n33098) );
  NANDN U33528 ( .A(n33318), .B(n33319), .Z(n33317) );
  NANDN U33529 ( .A(n33320), .B(n33321), .Z(n33319) );
  NANDN U33530 ( .A(n33321), .B(n33320), .Z(n33316) );
  ANDN U33531 ( .B(B[160]), .A(n62), .Z(n33100) );
  XNOR U33532 ( .A(n33108), .B(n33322), .Z(n33101) );
  XNOR U33533 ( .A(n33107), .B(n33105), .Z(n33322) );
  AND U33534 ( .A(n33323), .B(n33324), .Z(n33105) );
  NANDN U33535 ( .A(n33325), .B(n33326), .Z(n33324) );
  OR U33536 ( .A(n33327), .B(n33328), .Z(n33326) );
  NAND U33537 ( .A(n33328), .B(n33327), .Z(n33323) );
  ANDN U33538 ( .B(B[161]), .A(n63), .Z(n33107) );
  XNOR U33539 ( .A(n33115), .B(n33329), .Z(n33108) );
  XNOR U33540 ( .A(n33114), .B(n33112), .Z(n33329) );
  AND U33541 ( .A(n33330), .B(n33331), .Z(n33112) );
  NANDN U33542 ( .A(n33332), .B(n33333), .Z(n33331) );
  NANDN U33543 ( .A(n33334), .B(n33335), .Z(n33333) );
  NANDN U33544 ( .A(n33335), .B(n33334), .Z(n33330) );
  ANDN U33545 ( .B(B[162]), .A(n64), .Z(n33114) );
  XNOR U33546 ( .A(n33122), .B(n33336), .Z(n33115) );
  XNOR U33547 ( .A(n33121), .B(n33119), .Z(n33336) );
  AND U33548 ( .A(n33337), .B(n33338), .Z(n33119) );
  NANDN U33549 ( .A(n33339), .B(n33340), .Z(n33338) );
  OR U33550 ( .A(n33341), .B(n33342), .Z(n33340) );
  NAND U33551 ( .A(n33342), .B(n33341), .Z(n33337) );
  ANDN U33552 ( .B(B[163]), .A(n65), .Z(n33121) );
  XNOR U33553 ( .A(n33129), .B(n33343), .Z(n33122) );
  XNOR U33554 ( .A(n33128), .B(n33126), .Z(n33343) );
  AND U33555 ( .A(n33344), .B(n33345), .Z(n33126) );
  NANDN U33556 ( .A(n33346), .B(n33347), .Z(n33345) );
  NANDN U33557 ( .A(n33348), .B(n33349), .Z(n33347) );
  NANDN U33558 ( .A(n33349), .B(n33348), .Z(n33344) );
  ANDN U33559 ( .B(B[164]), .A(n66), .Z(n33128) );
  XNOR U33560 ( .A(n33136), .B(n33350), .Z(n33129) );
  XNOR U33561 ( .A(n33135), .B(n33133), .Z(n33350) );
  AND U33562 ( .A(n33351), .B(n33352), .Z(n33133) );
  NANDN U33563 ( .A(n33353), .B(n33354), .Z(n33352) );
  OR U33564 ( .A(n33355), .B(n33356), .Z(n33354) );
  NAND U33565 ( .A(n33356), .B(n33355), .Z(n33351) );
  ANDN U33566 ( .B(B[165]), .A(n67), .Z(n33135) );
  XNOR U33567 ( .A(n33143), .B(n33357), .Z(n33136) );
  XNOR U33568 ( .A(n33142), .B(n33140), .Z(n33357) );
  AND U33569 ( .A(n33358), .B(n33359), .Z(n33140) );
  NANDN U33570 ( .A(n33360), .B(n33361), .Z(n33359) );
  NANDN U33571 ( .A(n33362), .B(n33363), .Z(n33361) );
  NANDN U33572 ( .A(n33363), .B(n33362), .Z(n33358) );
  ANDN U33573 ( .B(B[166]), .A(n68), .Z(n33142) );
  XNOR U33574 ( .A(n33150), .B(n33364), .Z(n33143) );
  XNOR U33575 ( .A(n33149), .B(n33147), .Z(n33364) );
  AND U33576 ( .A(n33365), .B(n33366), .Z(n33147) );
  NANDN U33577 ( .A(n33367), .B(n33368), .Z(n33366) );
  OR U33578 ( .A(n33369), .B(n33370), .Z(n33368) );
  NAND U33579 ( .A(n33370), .B(n33369), .Z(n33365) );
  ANDN U33580 ( .B(B[167]), .A(n69), .Z(n33149) );
  XNOR U33581 ( .A(n33157), .B(n33371), .Z(n33150) );
  XNOR U33582 ( .A(n33156), .B(n33154), .Z(n33371) );
  AND U33583 ( .A(n33372), .B(n33373), .Z(n33154) );
  NANDN U33584 ( .A(n33374), .B(n33375), .Z(n33373) );
  NANDN U33585 ( .A(n33376), .B(n33377), .Z(n33375) );
  NANDN U33586 ( .A(n33377), .B(n33376), .Z(n33372) );
  ANDN U33587 ( .B(B[168]), .A(n70), .Z(n33156) );
  XNOR U33588 ( .A(n33164), .B(n33378), .Z(n33157) );
  XNOR U33589 ( .A(n33163), .B(n33161), .Z(n33378) );
  AND U33590 ( .A(n33379), .B(n33380), .Z(n33161) );
  NANDN U33591 ( .A(n33381), .B(n33382), .Z(n33380) );
  OR U33592 ( .A(n33383), .B(n33384), .Z(n33382) );
  NAND U33593 ( .A(n33384), .B(n33383), .Z(n33379) );
  ANDN U33594 ( .B(B[169]), .A(n71), .Z(n33163) );
  XNOR U33595 ( .A(n33171), .B(n33385), .Z(n33164) );
  XNOR U33596 ( .A(n33170), .B(n33168), .Z(n33385) );
  AND U33597 ( .A(n33386), .B(n33387), .Z(n33168) );
  NANDN U33598 ( .A(n33388), .B(n33389), .Z(n33387) );
  NANDN U33599 ( .A(n33390), .B(n33391), .Z(n33389) );
  NANDN U33600 ( .A(n33391), .B(n33390), .Z(n33386) );
  ANDN U33601 ( .B(B[170]), .A(n72), .Z(n33170) );
  XNOR U33602 ( .A(n33178), .B(n33392), .Z(n33171) );
  XNOR U33603 ( .A(n33177), .B(n33175), .Z(n33392) );
  AND U33604 ( .A(n33393), .B(n33394), .Z(n33175) );
  NANDN U33605 ( .A(n33395), .B(n33396), .Z(n33394) );
  OR U33606 ( .A(n33397), .B(n33398), .Z(n33396) );
  NAND U33607 ( .A(n33398), .B(n33397), .Z(n33393) );
  ANDN U33608 ( .B(B[171]), .A(n73), .Z(n33177) );
  XNOR U33609 ( .A(n33185), .B(n33399), .Z(n33178) );
  XNOR U33610 ( .A(n33184), .B(n33182), .Z(n33399) );
  AND U33611 ( .A(n33400), .B(n33401), .Z(n33182) );
  NANDN U33612 ( .A(n33402), .B(n33403), .Z(n33401) );
  NANDN U33613 ( .A(n33404), .B(n33405), .Z(n33403) );
  NANDN U33614 ( .A(n33405), .B(n33404), .Z(n33400) );
  ANDN U33615 ( .B(B[172]), .A(n74), .Z(n33184) );
  XNOR U33616 ( .A(n33192), .B(n33406), .Z(n33185) );
  XNOR U33617 ( .A(n33191), .B(n33189), .Z(n33406) );
  AND U33618 ( .A(n33407), .B(n33408), .Z(n33189) );
  NANDN U33619 ( .A(n33409), .B(n33410), .Z(n33408) );
  OR U33620 ( .A(n33411), .B(n33412), .Z(n33410) );
  NAND U33621 ( .A(n33412), .B(n33411), .Z(n33407) );
  ANDN U33622 ( .B(B[173]), .A(n75), .Z(n33191) );
  XNOR U33623 ( .A(n33199), .B(n33413), .Z(n33192) );
  XNOR U33624 ( .A(n33198), .B(n33196), .Z(n33413) );
  AND U33625 ( .A(n33414), .B(n33415), .Z(n33196) );
  NANDN U33626 ( .A(n33416), .B(n33417), .Z(n33415) );
  NANDN U33627 ( .A(n33418), .B(n33419), .Z(n33417) );
  NANDN U33628 ( .A(n33419), .B(n33418), .Z(n33414) );
  ANDN U33629 ( .B(B[174]), .A(n76), .Z(n33198) );
  XNOR U33630 ( .A(n33206), .B(n33420), .Z(n33199) );
  XNOR U33631 ( .A(n33205), .B(n33203), .Z(n33420) );
  AND U33632 ( .A(n33421), .B(n33422), .Z(n33203) );
  NANDN U33633 ( .A(n33423), .B(n33424), .Z(n33422) );
  OR U33634 ( .A(n33425), .B(n33426), .Z(n33424) );
  NAND U33635 ( .A(n33426), .B(n33425), .Z(n33421) );
  ANDN U33636 ( .B(B[175]), .A(n77), .Z(n33205) );
  XNOR U33637 ( .A(n33213), .B(n33427), .Z(n33206) );
  XNOR U33638 ( .A(n33212), .B(n33210), .Z(n33427) );
  AND U33639 ( .A(n33428), .B(n33429), .Z(n33210) );
  NANDN U33640 ( .A(n33430), .B(n33431), .Z(n33429) );
  NANDN U33641 ( .A(n33432), .B(n33433), .Z(n33431) );
  NANDN U33642 ( .A(n33433), .B(n33432), .Z(n33428) );
  ANDN U33643 ( .B(B[176]), .A(n78), .Z(n33212) );
  XNOR U33644 ( .A(n33220), .B(n33434), .Z(n33213) );
  XNOR U33645 ( .A(n33219), .B(n33217), .Z(n33434) );
  AND U33646 ( .A(n33435), .B(n33436), .Z(n33217) );
  NANDN U33647 ( .A(n33437), .B(n33438), .Z(n33436) );
  OR U33648 ( .A(n33439), .B(n33440), .Z(n33438) );
  NAND U33649 ( .A(n33440), .B(n33439), .Z(n33435) );
  ANDN U33650 ( .B(B[177]), .A(n79), .Z(n33219) );
  XNOR U33651 ( .A(n33227), .B(n33441), .Z(n33220) );
  XNOR U33652 ( .A(n33226), .B(n33224), .Z(n33441) );
  AND U33653 ( .A(n33442), .B(n33443), .Z(n33224) );
  NANDN U33654 ( .A(n33444), .B(n33445), .Z(n33443) );
  NANDN U33655 ( .A(n33446), .B(n33447), .Z(n33445) );
  NANDN U33656 ( .A(n33447), .B(n33446), .Z(n33442) );
  ANDN U33657 ( .B(B[178]), .A(n80), .Z(n33226) );
  XNOR U33658 ( .A(n33234), .B(n33448), .Z(n33227) );
  XNOR U33659 ( .A(n33233), .B(n33231), .Z(n33448) );
  AND U33660 ( .A(n33449), .B(n33450), .Z(n33231) );
  NANDN U33661 ( .A(n33451), .B(n33452), .Z(n33450) );
  OR U33662 ( .A(n33453), .B(n33454), .Z(n33452) );
  NAND U33663 ( .A(n33454), .B(n33453), .Z(n33449) );
  ANDN U33664 ( .B(B[179]), .A(n81), .Z(n33233) );
  XNOR U33665 ( .A(n33241), .B(n33455), .Z(n33234) );
  XNOR U33666 ( .A(n33240), .B(n33238), .Z(n33455) );
  AND U33667 ( .A(n33456), .B(n33457), .Z(n33238) );
  NANDN U33668 ( .A(n33458), .B(n33459), .Z(n33457) );
  NAND U33669 ( .A(n33460), .B(n33461), .Z(n33459) );
  ANDN U33670 ( .B(B[180]), .A(n82), .Z(n33240) );
  XOR U33671 ( .A(n33247), .B(n33462), .Z(n33241) );
  XNOR U33672 ( .A(n33245), .B(n33248), .Z(n33462) );
  NAND U33673 ( .A(A[2]), .B(B[181]), .Z(n33248) );
  NANDN U33674 ( .A(n33463), .B(n33464), .Z(n33245) );
  AND U33675 ( .A(A[0]), .B(B[182]), .Z(n33464) );
  XNOR U33676 ( .A(n33250), .B(n33465), .Z(n33247) );
  NAND U33677 ( .A(A[0]), .B(B[183]), .Z(n33465) );
  NAND U33678 ( .A(B[182]), .B(A[1]), .Z(n33250) );
  NAND U33679 ( .A(n33466), .B(n33467), .Z(n430) );
  NANDN U33680 ( .A(n33468), .B(n33469), .Z(n33467) );
  OR U33681 ( .A(n33470), .B(n33471), .Z(n33469) );
  NAND U33682 ( .A(n33471), .B(n33470), .Z(n33466) );
  XOR U33683 ( .A(n432), .B(n431), .Z(\A1[180] ) );
  XOR U33684 ( .A(n33471), .B(n33472), .Z(n431) );
  XNOR U33685 ( .A(n33470), .B(n33468), .Z(n33472) );
  AND U33686 ( .A(n33473), .B(n33474), .Z(n33468) );
  NANDN U33687 ( .A(n33475), .B(n33476), .Z(n33474) );
  NANDN U33688 ( .A(n33477), .B(n33478), .Z(n33476) );
  NANDN U33689 ( .A(n33478), .B(n33477), .Z(n33473) );
  ANDN U33690 ( .B(B[151]), .A(n54), .Z(n33470) );
  XNOR U33691 ( .A(n33265), .B(n33479), .Z(n33471) );
  XNOR U33692 ( .A(n33264), .B(n33262), .Z(n33479) );
  AND U33693 ( .A(n33480), .B(n33481), .Z(n33262) );
  NANDN U33694 ( .A(n33482), .B(n33483), .Z(n33481) );
  OR U33695 ( .A(n33484), .B(n33485), .Z(n33483) );
  NAND U33696 ( .A(n33485), .B(n33484), .Z(n33480) );
  ANDN U33697 ( .B(B[152]), .A(n55), .Z(n33264) );
  XNOR U33698 ( .A(n33272), .B(n33486), .Z(n33265) );
  XNOR U33699 ( .A(n33271), .B(n33269), .Z(n33486) );
  AND U33700 ( .A(n33487), .B(n33488), .Z(n33269) );
  NANDN U33701 ( .A(n33489), .B(n33490), .Z(n33488) );
  NANDN U33702 ( .A(n33491), .B(n33492), .Z(n33490) );
  NANDN U33703 ( .A(n33492), .B(n33491), .Z(n33487) );
  ANDN U33704 ( .B(B[153]), .A(n56), .Z(n33271) );
  XNOR U33705 ( .A(n33279), .B(n33493), .Z(n33272) );
  XNOR U33706 ( .A(n33278), .B(n33276), .Z(n33493) );
  AND U33707 ( .A(n33494), .B(n33495), .Z(n33276) );
  NANDN U33708 ( .A(n33496), .B(n33497), .Z(n33495) );
  OR U33709 ( .A(n33498), .B(n33499), .Z(n33497) );
  NAND U33710 ( .A(n33499), .B(n33498), .Z(n33494) );
  ANDN U33711 ( .B(B[154]), .A(n57), .Z(n33278) );
  XNOR U33712 ( .A(n33286), .B(n33500), .Z(n33279) );
  XNOR U33713 ( .A(n33285), .B(n33283), .Z(n33500) );
  AND U33714 ( .A(n33501), .B(n33502), .Z(n33283) );
  NANDN U33715 ( .A(n33503), .B(n33504), .Z(n33502) );
  NANDN U33716 ( .A(n33505), .B(n33506), .Z(n33504) );
  NANDN U33717 ( .A(n33506), .B(n33505), .Z(n33501) );
  ANDN U33718 ( .B(B[155]), .A(n58), .Z(n33285) );
  XNOR U33719 ( .A(n33293), .B(n33507), .Z(n33286) );
  XNOR U33720 ( .A(n33292), .B(n33290), .Z(n33507) );
  AND U33721 ( .A(n33508), .B(n33509), .Z(n33290) );
  NANDN U33722 ( .A(n33510), .B(n33511), .Z(n33509) );
  OR U33723 ( .A(n33512), .B(n33513), .Z(n33511) );
  NAND U33724 ( .A(n33513), .B(n33512), .Z(n33508) );
  ANDN U33725 ( .B(B[156]), .A(n59), .Z(n33292) );
  XNOR U33726 ( .A(n33300), .B(n33514), .Z(n33293) );
  XNOR U33727 ( .A(n33299), .B(n33297), .Z(n33514) );
  AND U33728 ( .A(n33515), .B(n33516), .Z(n33297) );
  NANDN U33729 ( .A(n33517), .B(n33518), .Z(n33516) );
  NANDN U33730 ( .A(n33519), .B(n33520), .Z(n33518) );
  NANDN U33731 ( .A(n33520), .B(n33519), .Z(n33515) );
  ANDN U33732 ( .B(B[157]), .A(n60), .Z(n33299) );
  XNOR U33733 ( .A(n33307), .B(n33521), .Z(n33300) );
  XNOR U33734 ( .A(n33306), .B(n33304), .Z(n33521) );
  AND U33735 ( .A(n33522), .B(n33523), .Z(n33304) );
  NANDN U33736 ( .A(n33524), .B(n33525), .Z(n33523) );
  OR U33737 ( .A(n33526), .B(n33527), .Z(n33525) );
  NAND U33738 ( .A(n33527), .B(n33526), .Z(n33522) );
  ANDN U33739 ( .B(B[158]), .A(n61), .Z(n33306) );
  XNOR U33740 ( .A(n33314), .B(n33528), .Z(n33307) );
  XNOR U33741 ( .A(n33313), .B(n33311), .Z(n33528) );
  AND U33742 ( .A(n33529), .B(n33530), .Z(n33311) );
  NANDN U33743 ( .A(n33531), .B(n33532), .Z(n33530) );
  NANDN U33744 ( .A(n33533), .B(n33534), .Z(n33532) );
  NANDN U33745 ( .A(n33534), .B(n33533), .Z(n33529) );
  ANDN U33746 ( .B(B[159]), .A(n62), .Z(n33313) );
  XNOR U33747 ( .A(n33321), .B(n33535), .Z(n33314) );
  XNOR U33748 ( .A(n33320), .B(n33318), .Z(n33535) );
  AND U33749 ( .A(n33536), .B(n33537), .Z(n33318) );
  NANDN U33750 ( .A(n33538), .B(n33539), .Z(n33537) );
  OR U33751 ( .A(n33540), .B(n33541), .Z(n33539) );
  NAND U33752 ( .A(n33541), .B(n33540), .Z(n33536) );
  ANDN U33753 ( .B(B[160]), .A(n63), .Z(n33320) );
  XNOR U33754 ( .A(n33328), .B(n33542), .Z(n33321) );
  XNOR U33755 ( .A(n33327), .B(n33325), .Z(n33542) );
  AND U33756 ( .A(n33543), .B(n33544), .Z(n33325) );
  NANDN U33757 ( .A(n33545), .B(n33546), .Z(n33544) );
  NANDN U33758 ( .A(n33547), .B(n33548), .Z(n33546) );
  NANDN U33759 ( .A(n33548), .B(n33547), .Z(n33543) );
  ANDN U33760 ( .B(B[161]), .A(n64), .Z(n33327) );
  XNOR U33761 ( .A(n33335), .B(n33549), .Z(n33328) );
  XNOR U33762 ( .A(n33334), .B(n33332), .Z(n33549) );
  AND U33763 ( .A(n33550), .B(n33551), .Z(n33332) );
  NANDN U33764 ( .A(n33552), .B(n33553), .Z(n33551) );
  OR U33765 ( .A(n33554), .B(n33555), .Z(n33553) );
  NAND U33766 ( .A(n33555), .B(n33554), .Z(n33550) );
  ANDN U33767 ( .B(B[162]), .A(n65), .Z(n33334) );
  XNOR U33768 ( .A(n33342), .B(n33556), .Z(n33335) );
  XNOR U33769 ( .A(n33341), .B(n33339), .Z(n33556) );
  AND U33770 ( .A(n33557), .B(n33558), .Z(n33339) );
  NANDN U33771 ( .A(n33559), .B(n33560), .Z(n33558) );
  NANDN U33772 ( .A(n33561), .B(n33562), .Z(n33560) );
  NANDN U33773 ( .A(n33562), .B(n33561), .Z(n33557) );
  ANDN U33774 ( .B(B[163]), .A(n66), .Z(n33341) );
  XNOR U33775 ( .A(n33349), .B(n33563), .Z(n33342) );
  XNOR U33776 ( .A(n33348), .B(n33346), .Z(n33563) );
  AND U33777 ( .A(n33564), .B(n33565), .Z(n33346) );
  NANDN U33778 ( .A(n33566), .B(n33567), .Z(n33565) );
  OR U33779 ( .A(n33568), .B(n33569), .Z(n33567) );
  NAND U33780 ( .A(n33569), .B(n33568), .Z(n33564) );
  ANDN U33781 ( .B(B[164]), .A(n67), .Z(n33348) );
  XNOR U33782 ( .A(n33356), .B(n33570), .Z(n33349) );
  XNOR U33783 ( .A(n33355), .B(n33353), .Z(n33570) );
  AND U33784 ( .A(n33571), .B(n33572), .Z(n33353) );
  NANDN U33785 ( .A(n33573), .B(n33574), .Z(n33572) );
  NANDN U33786 ( .A(n33575), .B(n33576), .Z(n33574) );
  NANDN U33787 ( .A(n33576), .B(n33575), .Z(n33571) );
  ANDN U33788 ( .B(B[165]), .A(n68), .Z(n33355) );
  XNOR U33789 ( .A(n33363), .B(n33577), .Z(n33356) );
  XNOR U33790 ( .A(n33362), .B(n33360), .Z(n33577) );
  AND U33791 ( .A(n33578), .B(n33579), .Z(n33360) );
  NANDN U33792 ( .A(n33580), .B(n33581), .Z(n33579) );
  OR U33793 ( .A(n33582), .B(n33583), .Z(n33581) );
  NAND U33794 ( .A(n33583), .B(n33582), .Z(n33578) );
  ANDN U33795 ( .B(B[166]), .A(n69), .Z(n33362) );
  XNOR U33796 ( .A(n33370), .B(n33584), .Z(n33363) );
  XNOR U33797 ( .A(n33369), .B(n33367), .Z(n33584) );
  AND U33798 ( .A(n33585), .B(n33586), .Z(n33367) );
  NANDN U33799 ( .A(n33587), .B(n33588), .Z(n33586) );
  NANDN U33800 ( .A(n33589), .B(n33590), .Z(n33588) );
  NANDN U33801 ( .A(n33590), .B(n33589), .Z(n33585) );
  ANDN U33802 ( .B(B[167]), .A(n70), .Z(n33369) );
  XNOR U33803 ( .A(n33377), .B(n33591), .Z(n33370) );
  XNOR U33804 ( .A(n33376), .B(n33374), .Z(n33591) );
  AND U33805 ( .A(n33592), .B(n33593), .Z(n33374) );
  NANDN U33806 ( .A(n33594), .B(n33595), .Z(n33593) );
  OR U33807 ( .A(n33596), .B(n33597), .Z(n33595) );
  NAND U33808 ( .A(n33597), .B(n33596), .Z(n33592) );
  ANDN U33809 ( .B(B[168]), .A(n71), .Z(n33376) );
  XNOR U33810 ( .A(n33384), .B(n33598), .Z(n33377) );
  XNOR U33811 ( .A(n33383), .B(n33381), .Z(n33598) );
  AND U33812 ( .A(n33599), .B(n33600), .Z(n33381) );
  NANDN U33813 ( .A(n33601), .B(n33602), .Z(n33600) );
  NANDN U33814 ( .A(n33603), .B(n33604), .Z(n33602) );
  NANDN U33815 ( .A(n33604), .B(n33603), .Z(n33599) );
  ANDN U33816 ( .B(B[169]), .A(n72), .Z(n33383) );
  XNOR U33817 ( .A(n33391), .B(n33605), .Z(n33384) );
  XNOR U33818 ( .A(n33390), .B(n33388), .Z(n33605) );
  AND U33819 ( .A(n33606), .B(n33607), .Z(n33388) );
  NANDN U33820 ( .A(n33608), .B(n33609), .Z(n33607) );
  OR U33821 ( .A(n33610), .B(n33611), .Z(n33609) );
  NAND U33822 ( .A(n33611), .B(n33610), .Z(n33606) );
  ANDN U33823 ( .B(B[170]), .A(n73), .Z(n33390) );
  XNOR U33824 ( .A(n33398), .B(n33612), .Z(n33391) );
  XNOR U33825 ( .A(n33397), .B(n33395), .Z(n33612) );
  AND U33826 ( .A(n33613), .B(n33614), .Z(n33395) );
  NANDN U33827 ( .A(n33615), .B(n33616), .Z(n33614) );
  NANDN U33828 ( .A(n33617), .B(n33618), .Z(n33616) );
  NANDN U33829 ( .A(n33618), .B(n33617), .Z(n33613) );
  ANDN U33830 ( .B(B[171]), .A(n74), .Z(n33397) );
  XNOR U33831 ( .A(n33405), .B(n33619), .Z(n33398) );
  XNOR U33832 ( .A(n33404), .B(n33402), .Z(n33619) );
  AND U33833 ( .A(n33620), .B(n33621), .Z(n33402) );
  NANDN U33834 ( .A(n33622), .B(n33623), .Z(n33621) );
  OR U33835 ( .A(n33624), .B(n33625), .Z(n33623) );
  NAND U33836 ( .A(n33625), .B(n33624), .Z(n33620) );
  ANDN U33837 ( .B(B[172]), .A(n75), .Z(n33404) );
  XNOR U33838 ( .A(n33412), .B(n33626), .Z(n33405) );
  XNOR U33839 ( .A(n33411), .B(n33409), .Z(n33626) );
  AND U33840 ( .A(n33627), .B(n33628), .Z(n33409) );
  NANDN U33841 ( .A(n33629), .B(n33630), .Z(n33628) );
  NANDN U33842 ( .A(n33631), .B(n33632), .Z(n33630) );
  NANDN U33843 ( .A(n33632), .B(n33631), .Z(n33627) );
  ANDN U33844 ( .B(B[173]), .A(n76), .Z(n33411) );
  XNOR U33845 ( .A(n33419), .B(n33633), .Z(n33412) );
  XNOR U33846 ( .A(n33418), .B(n33416), .Z(n33633) );
  AND U33847 ( .A(n33634), .B(n33635), .Z(n33416) );
  NANDN U33848 ( .A(n33636), .B(n33637), .Z(n33635) );
  OR U33849 ( .A(n33638), .B(n33639), .Z(n33637) );
  NAND U33850 ( .A(n33639), .B(n33638), .Z(n33634) );
  ANDN U33851 ( .B(B[174]), .A(n77), .Z(n33418) );
  XNOR U33852 ( .A(n33426), .B(n33640), .Z(n33419) );
  XNOR U33853 ( .A(n33425), .B(n33423), .Z(n33640) );
  AND U33854 ( .A(n33641), .B(n33642), .Z(n33423) );
  NANDN U33855 ( .A(n33643), .B(n33644), .Z(n33642) );
  NANDN U33856 ( .A(n33645), .B(n33646), .Z(n33644) );
  NANDN U33857 ( .A(n33646), .B(n33645), .Z(n33641) );
  ANDN U33858 ( .B(B[175]), .A(n78), .Z(n33425) );
  XNOR U33859 ( .A(n33433), .B(n33647), .Z(n33426) );
  XNOR U33860 ( .A(n33432), .B(n33430), .Z(n33647) );
  AND U33861 ( .A(n33648), .B(n33649), .Z(n33430) );
  NANDN U33862 ( .A(n33650), .B(n33651), .Z(n33649) );
  OR U33863 ( .A(n33652), .B(n33653), .Z(n33651) );
  NAND U33864 ( .A(n33653), .B(n33652), .Z(n33648) );
  ANDN U33865 ( .B(B[176]), .A(n79), .Z(n33432) );
  XNOR U33866 ( .A(n33440), .B(n33654), .Z(n33433) );
  XNOR U33867 ( .A(n33439), .B(n33437), .Z(n33654) );
  AND U33868 ( .A(n33655), .B(n33656), .Z(n33437) );
  NANDN U33869 ( .A(n33657), .B(n33658), .Z(n33656) );
  NANDN U33870 ( .A(n33659), .B(n33660), .Z(n33658) );
  NANDN U33871 ( .A(n33660), .B(n33659), .Z(n33655) );
  ANDN U33872 ( .B(B[177]), .A(n80), .Z(n33439) );
  XNOR U33873 ( .A(n33447), .B(n33661), .Z(n33440) );
  XNOR U33874 ( .A(n33446), .B(n33444), .Z(n33661) );
  AND U33875 ( .A(n33662), .B(n33663), .Z(n33444) );
  NANDN U33876 ( .A(n33664), .B(n33665), .Z(n33663) );
  OR U33877 ( .A(n33666), .B(n33667), .Z(n33665) );
  NAND U33878 ( .A(n33667), .B(n33666), .Z(n33662) );
  ANDN U33879 ( .B(B[178]), .A(n81), .Z(n33446) );
  XNOR U33880 ( .A(n33454), .B(n33668), .Z(n33447) );
  XNOR U33881 ( .A(n33453), .B(n33451), .Z(n33668) );
  AND U33882 ( .A(n33669), .B(n33670), .Z(n33451) );
  NANDN U33883 ( .A(n33671), .B(n33672), .Z(n33670) );
  NAND U33884 ( .A(n33673), .B(n33674), .Z(n33672) );
  ANDN U33885 ( .B(B[179]), .A(n82), .Z(n33453) );
  XOR U33886 ( .A(n33460), .B(n33675), .Z(n33454) );
  XNOR U33887 ( .A(n33458), .B(n33461), .Z(n33675) );
  NAND U33888 ( .A(A[2]), .B(B[180]), .Z(n33461) );
  NANDN U33889 ( .A(n33676), .B(n33677), .Z(n33458) );
  AND U33890 ( .A(A[0]), .B(B[181]), .Z(n33677) );
  XNOR U33891 ( .A(n33463), .B(n33678), .Z(n33460) );
  NAND U33892 ( .A(A[0]), .B(B[182]), .Z(n33678) );
  NAND U33893 ( .A(B[181]), .B(A[1]), .Z(n33463) );
  NAND U33894 ( .A(n33679), .B(n33680), .Z(n432) );
  NANDN U33895 ( .A(n33681), .B(n33682), .Z(n33680) );
  OR U33896 ( .A(n33683), .B(n33684), .Z(n33682) );
  NAND U33897 ( .A(n33684), .B(n33683), .Z(n33679) );
  XOR U33898 ( .A(n31431), .B(n33685), .Z(\A1[17] ) );
  XNOR U33899 ( .A(n31430), .B(n31428), .Z(n33685) );
  AND U33900 ( .A(n33686), .B(n33687), .Z(n31428) );
  NAND U33901 ( .A(n33688), .B(n33689), .Z(n33687) );
  NANDN U33902 ( .A(n33690), .B(n33691), .Z(n33688) );
  NANDN U33903 ( .A(n33691), .B(n33690), .Z(n33686) );
  ANDN U33904 ( .B(B[0]), .A(n66), .Z(n31430) );
  XNOR U33905 ( .A(n31438), .B(n33692), .Z(n31431) );
  XNOR U33906 ( .A(n31437), .B(n31435), .Z(n33692) );
  AND U33907 ( .A(n33693), .B(n33694), .Z(n31435) );
  NANDN U33908 ( .A(n33695), .B(n33696), .Z(n33694) );
  OR U33909 ( .A(n33697), .B(n33698), .Z(n33696) );
  NAND U33910 ( .A(n33698), .B(n33697), .Z(n33693) );
  ANDN U33911 ( .B(B[1]), .A(n67), .Z(n31437) );
  XNOR U33912 ( .A(n31445), .B(n33699), .Z(n31438) );
  XNOR U33913 ( .A(n31444), .B(n31442), .Z(n33699) );
  AND U33914 ( .A(n33700), .B(n33701), .Z(n31442) );
  NANDN U33915 ( .A(n33702), .B(n33703), .Z(n33701) );
  NANDN U33916 ( .A(n33704), .B(n33705), .Z(n33703) );
  NANDN U33917 ( .A(n33705), .B(n33704), .Z(n33700) );
  ANDN U33918 ( .B(B[2]), .A(n68), .Z(n31444) );
  XNOR U33919 ( .A(n31452), .B(n33706), .Z(n31445) );
  XNOR U33920 ( .A(n31451), .B(n31449), .Z(n33706) );
  AND U33921 ( .A(n33707), .B(n33708), .Z(n31449) );
  NANDN U33922 ( .A(n33709), .B(n33710), .Z(n33708) );
  OR U33923 ( .A(n33711), .B(n33712), .Z(n33710) );
  NAND U33924 ( .A(n33712), .B(n33711), .Z(n33707) );
  ANDN U33925 ( .B(B[3]), .A(n69), .Z(n31451) );
  XNOR U33926 ( .A(n31459), .B(n33713), .Z(n31452) );
  XNOR U33927 ( .A(n31458), .B(n31456), .Z(n33713) );
  AND U33928 ( .A(n33714), .B(n33715), .Z(n31456) );
  NANDN U33929 ( .A(n33716), .B(n33717), .Z(n33715) );
  NANDN U33930 ( .A(n33718), .B(n33719), .Z(n33717) );
  NANDN U33931 ( .A(n33719), .B(n33718), .Z(n33714) );
  ANDN U33932 ( .B(B[4]), .A(n70), .Z(n31458) );
  XNOR U33933 ( .A(n31466), .B(n33720), .Z(n31459) );
  XNOR U33934 ( .A(n31465), .B(n31463), .Z(n33720) );
  AND U33935 ( .A(n33721), .B(n33722), .Z(n31463) );
  NANDN U33936 ( .A(n33723), .B(n33724), .Z(n33722) );
  OR U33937 ( .A(n33725), .B(n33726), .Z(n33724) );
  NAND U33938 ( .A(n33726), .B(n33725), .Z(n33721) );
  ANDN U33939 ( .B(B[5]), .A(n71), .Z(n31465) );
  XNOR U33940 ( .A(n31473), .B(n33727), .Z(n31466) );
  XNOR U33941 ( .A(n31472), .B(n31470), .Z(n33727) );
  AND U33942 ( .A(n33728), .B(n33729), .Z(n31470) );
  NANDN U33943 ( .A(n33730), .B(n33731), .Z(n33729) );
  NANDN U33944 ( .A(n33732), .B(n33733), .Z(n33731) );
  NANDN U33945 ( .A(n33733), .B(n33732), .Z(n33728) );
  ANDN U33946 ( .B(B[6]), .A(n72), .Z(n31472) );
  XNOR U33947 ( .A(n31480), .B(n33734), .Z(n31473) );
  XNOR U33948 ( .A(n31479), .B(n31477), .Z(n33734) );
  AND U33949 ( .A(n33735), .B(n33736), .Z(n31477) );
  NANDN U33950 ( .A(n33737), .B(n33738), .Z(n33736) );
  OR U33951 ( .A(n33739), .B(n33740), .Z(n33738) );
  NAND U33952 ( .A(n33740), .B(n33739), .Z(n33735) );
  ANDN U33953 ( .B(B[7]), .A(n73), .Z(n31479) );
  XNOR U33954 ( .A(n31487), .B(n33741), .Z(n31480) );
  XNOR U33955 ( .A(n31486), .B(n31484), .Z(n33741) );
  AND U33956 ( .A(n33742), .B(n33743), .Z(n31484) );
  NANDN U33957 ( .A(n33744), .B(n33745), .Z(n33743) );
  NANDN U33958 ( .A(n33746), .B(n33747), .Z(n33745) );
  NANDN U33959 ( .A(n33747), .B(n33746), .Z(n33742) );
  ANDN U33960 ( .B(B[8]), .A(n74), .Z(n31486) );
  XNOR U33961 ( .A(n31494), .B(n33748), .Z(n31487) );
  XNOR U33962 ( .A(n31493), .B(n31491), .Z(n33748) );
  AND U33963 ( .A(n33749), .B(n33750), .Z(n31491) );
  NANDN U33964 ( .A(n33751), .B(n33752), .Z(n33750) );
  OR U33965 ( .A(n33753), .B(n33754), .Z(n33752) );
  NAND U33966 ( .A(n33754), .B(n33753), .Z(n33749) );
  ANDN U33967 ( .B(B[9]), .A(n75), .Z(n31493) );
  XNOR U33968 ( .A(n31501), .B(n33755), .Z(n31494) );
  XNOR U33969 ( .A(n31500), .B(n31498), .Z(n33755) );
  AND U33970 ( .A(n33756), .B(n33757), .Z(n31498) );
  NANDN U33971 ( .A(n33758), .B(n33759), .Z(n33757) );
  NANDN U33972 ( .A(n33760), .B(n33761), .Z(n33759) );
  NANDN U33973 ( .A(n33761), .B(n33760), .Z(n33756) );
  ANDN U33974 ( .B(B[10]), .A(n76), .Z(n31500) );
  XNOR U33975 ( .A(n31508), .B(n33762), .Z(n31501) );
  XNOR U33976 ( .A(n31507), .B(n31505), .Z(n33762) );
  AND U33977 ( .A(n33763), .B(n33764), .Z(n31505) );
  NANDN U33978 ( .A(n33765), .B(n33766), .Z(n33764) );
  OR U33979 ( .A(n33767), .B(n33768), .Z(n33766) );
  NAND U33980 ( .A(n33768), .B(n33767), .Z(n33763) );
  ANDN U33981 ( .B(B[11]), .A(n77), .Z(n31507) );
  XNOR U33982 ( .A(n31515), .B(n33769), .Z(n31508) );
  XNOR U33983 ( .A(n31514), .B(n31512), .Z(n33769) );
  AND U33984 ( .A(n33770), .B(n33771), .Z(n31512) );
  NANDN U33985 ( .A(n33772), .B(n33773), .Z(n33771) );
  NANDN U33986 ( .A(n33774), .B(n33775), .Z(n33773) );
  NANDN U33987 ( .A(n33775), .B(n33774), .Z(n33770) );
  ANDN U33988 ( .B(B[12]), .A(n78), .Z(n31514) );
  XNOR U33989 ( .A(n31522), .B(n33776), .Z(n31515) );
  XNOR U33990 ( .A(n31521), .B(n31519), .Z(n33776) );
  AND U33991 ( .A(n33777), .B(n33778), .Z(n31519) );
  NANDN U33992 ( .A(n33779), .B(n33780), .Z(n33778) );
  OR U33993 ( .A(n33781), .B(n33782), .Z(n33780) );
  NAND U33994 ( .A(n33782), .B(n33781), .Z(n33777) );
  ANDN U33995 ( .B(B[13]), .A(n79), .Z(n31521) );
  XNOR U33996 ( .A(n31529), .B(n33783), .Z(n31522) );
  XNOR U33997 ( .A(n31528), .B(n31526), .Z(n33783) );
  AND U33998 ( .A(n33784), .B(n33785), .Z(n31526) );
  NANDN U33999 ( .A(n33786), .B(n33787), .Z(n33785) );
  NANDN U34000 ( .A(n33788), .B(n33789), .Z(n33787) );
  NANDN U34001 ( .A(n33789), .B(n33788), .Z(n33784) );
  ANDN U34002 ( .B(B[14]), .A(n80), .Z(n31528) );
  XNOR U34003 ( .A(n31536), .B(n33790), .Z(n31529) );
  XNOR U34004 ( .A(n31535), .B(n31533), .Z(n33790) );
  AND U34005 ( .A(n33791), .B(n33792), .Z(n31533) );
  NANDN U34006 ( .A(n33793), .B(n33794), .Z(n33792) );
  OR U34007 ( .A(n33795), .B(n33796), .Z(n33794) );
  NAND U34008 ( .A(n33796), .B(n33795), .Z(n33791) );
  ANDN U34009 ( .B(B[15]), .A(n81), .Z(n31535) );
  XNOR U34010 ( .A(n31543), .B(n33797), .Z(n31536) );
  XNOR U34011 ( .A(n31542), .B(n31540), .Z(n33797) );
  AND U34012 ( .A(n33798), .B(n33799), .Z(n31540) );
  NANDN U34013 ( .A(n33800), .B(n33801), .Z(n33799) );
  NAND U34014 ( .A(n33802), .B(n33803), .Z(n33801) );
  ANDN U34015 ( .B(B[16]), .A(n82), .Z(n31542) );
  XOR U34016 ( .A(n31549), .B(n33804), .Z(n31543) );
  XNOR U34017 ( .A(n31547), .B(n31550), .Z(n33804) );
  NAND U34018 ( .A(A[2]), .B(B[17]), .Z(n31550) );
  NANDN U34019 ( .A(n33805), .B(n33806), .Z(n31547) );
  AND U34020 ( .A(A[0]), .B(B[18]), .Z(n33806) );
  XNOR U34021 ( .A(n31552), .B(n33807), .Z(n31549) );
  NAND U34022 ( .A(A[0]), .B(B[19]), .Z(n33807) );
  NAND U34023 ( .A(B[18]), .B(A[1]), .Z(n31552) );
  XOR U34024 ( .A(n434), .B(n433), .Z(\A1[179] ) );
  XOR U34025 ( .A(n33684), .B(n33808), .Z(n433) );
  XNOR U34026 ( .A(n33683), .B(n33681), .Z(n33808) );
  AND U34027 ( .A(n33809), .B(n33810), .Z(n33681) );
  NANDN U34028 ( .A(n33811), .B(n33812), .Z(n33810) );
  NANDN U34029 ( .A(n33813), .B(n33814), .Z(n33812) );
  NANDN U34030 ( .A(n33814), .B(n33813), .Z(n33809) );
  ANDN U34031 ( .B(B[150]), .A(n54), .Z(n33683) );
  XNOR U34032 ( .A(n33478), .B(n33815), .Z(n33684) );
  XNOR U34033 ( .A(n33477), .B(n33475), .Z(n33815) );
  AND U34034 ( .A(n33816), .B(n33817), .Z(n33475) );
  NANDN U34035 ( .A(n33818), .B(n33819), .Z(n33817) );
  OR U34036 ( .A(n33820), .B(n33821), .Z(n33819) );
  NAND U34037 ( .A(n33821), .B(n33820), .Z(n33816) );
  ANDN U34038 ( .B(B[151]), .A(n55), .Z(n33477) );
  XNOR U34039 ( .A(n33485), .B(n33822), .Z(n33478) );
  XNOR U34040 ( .A(n33484), .B(n33482), .Z(n33822) );
  AND U34041 ( .A(n33823), .B(n33824), .Z(n33482) );
  NANDN U34042 ( .A(n33825), .B(n33826), .Z(n33824) );
  NANDN U34043 ( .A(n33827), .B(n33828), .Z(n33826) );
  NANDN U34044 ( .A(n33828), .B(n33827), .Z(n33823) );
  ANDN U34045 ( .B(B[152]), .A(n56), .Z(n33484) );
  XNOR U34046 ( .A(n33492), .B(n33829), .Z(n33485) );
  XNOR U34047 ( .A(n33491), .B(n33489), .Z(n33829) );
  AND U34048 ( .A(n33830), .B(n33831), .Z(n33489) );
  NANDN U34049 ( .A(n33832), .B(n33833), .Z(n33831) );
  OR U34050 ( .A(n33834), .B(n33835), .Z(n33833) );
  NAND U34051 ( .A(n33835), .B(n33834), .Z(n33830) );
  ANDN U34052 ( .B(B[153]), .A(n57), .Z(n33491) );
  XNOR U34053 ( .A(n33499), .B(n33836), .Z(n33492) );
  XNOR U34054 ( .A(n33498), .B(n33496), .Z(n33836) );
  AND U34055 ( .A(n33837), .B(n33838), .Z(n33496) );
  NANDN U34056 ( .A(n33839), .B(n33840), .Z(n33838) );
  NANDN U34057 ( .A(n33841), .B(n33842), .Z(n33840) );
  NANDN U34058 ( .A(n33842), .B(n33841), .Z(n33837) );
  ANDN U34059 ( .B(B[154]), .A(n58), .Z(n33498) );
  XNOR U34060 ( .A(n33506), .B(n33843), .Z(n33499) );
  XNOR U34061 ( .A(n33505), .B(n33503), .Z(n33843) );
  AND U34062 ( .A(n33844), .B(n33845), .Z(n33503) );
  NANDN U34063 ( .A(n33846), .B(n33847), .Z(n33845) );
  OR U34064 ( .A(n33848), .B(n33849), .Z(n33847) );
  NAND U34065 ( .A(n33849), .B(n33848), .Z(n33844) );
  ANDN U34066 ( .B(B[155]), .A(n59), .Z(n33505) );
  XNOR U34067 ( .A(n33513), .B(n33850), .Z(n33506) );
  XNOR U34068 ( .A(n33512), .B(n33510), .Z(n33850) );
  AND U34069 ( .A(n33851), .B(n33852), .Z(n33510) );
  NANDN U34070 ( .A(n33853), .B(n33854), .Z(n33852) );
  NANDN U34071 ( .A(n33855), .B(n33856), .Z(n33854) );
  NANDN U34072 ( .A(n33856), .B(n33855), .Z(n33851) );
  ANDN U34073 ( .B(B[156]), .A(n60), .Z(n33512) );
  XNOR U34074 ( .A(n33520), .B(n33857), .Z(n33513) );
  XNOR U34075 ( .A(n33519), .B(n33517), .Z(n33857) );
  AND U34076 ( .A(n33858), .B(n33859), .Z(n33517) );
  NANDN U34077 ( .A(n33860), .B(n33861), .Z(n33859) );
  OR U34078 ( .A(n33862), .B(n33863), .Z(n33861) );
  NAND U34079 ( .A(n33863), .B(n33862), .Z(n33858) );
  ANDN U34080 ( .B(B[157]), .A(n61), .Z(n33519) );
  XNOR U34081 ( .A(n33527), .B(n33864), .Z(n33520) );
  XNOR U34082 ( .A(n33526), .B(n33524), .Z(n33864) );
  AND U34083 ( .A(n33865), .B(n33866), .Z(n33524) );
  NANDN U34084 ( .A(n33867), .B(n33868), .Z(n33866) );
  NANDN U34085 ( .A(n33869), .B(n33870), .Z(n33868) );
  NANDN U34086 ( .A(n33870), .B(n33869), .Z(n33865) );
  ANDN U34087 ( .B(B[158]), .A(n62), .Z(n33526) );
  XNOR U34088 ( .A(n33534), .B(n33871), .Z(n33527) );
  XNOR U34089 ( .A(n33533), .B(n33531), .Z(n33871) );
  AND U34090 ( .A(n33872), .B(n33873), .Z(n33531) );
  NANDN U34091 ( .A(n33874), .B(n33875), .Z(n33873) );
  OR U34092 ( .A(n33876), .B(n33877), .Z(n33875) );
  NAND U34093 ( .A(n33877), .B(n33876), .Z(n33872) );
  ANDN U34094 ( .B(B[159]), .A(n63), .Z(n33533) );
  XNOR U34095 ( .A(n33541), .B(n33878), .Z(n33534) );
  XNOR U34096 ( .A(n33540), .B(n33538), .Z(n33878) );
  AND U34097 ( .A(n33879), .B(n33880), .Z(n33538) );
  NANDN U34098 ( .A(n33881), .B(n33882), .Z(n33880) );
  NANDN U34099 ( .A(n33883), .B(n33884), .Z(n33882) );
  NANDN U34100 ( .A(n33884), .B(n33883), .Z(n33879) );
  ANDN U34101 ( .B(B[160]), .A(n64), .Z(n33540) );
  XNOR U34102 ( .A(n33548), .B(n33885), .Z(n33541) );
  XNOR U34103 ( .A(n33547), .B(n33545), .Z(n33885) );
  AND U34104 ( .A(n33886), .B(n33887), .Z(n33545) );
  NANDN U34105 ( .A(n33888), .B(n33889), .Z(n33887) );
  OR U34106 ( .A(n33890), .B(n33891), .Z(n33889) );
  NAND U34107 ( .A(n33891), .B(n33890), .Z(n33886) );
  ANDN U34108 ( .B(B[161]), .A(n65), .Z(n33547) );
  XNOR U34109 ( .A(n33555), .B(n33892), .Z(n33548) );
  XNOR U34110 ( .A(n33554), .B(n33552), .Z(n33892) );
  AND U34111 ( .A(n33893), .B(n33894), .Z(n33552) );
  NANDN U34112 ( .A(n33895), .B(n33896), .Z(n33894) );
  NANDN U34113 ( .A(n33897), .B(n33898), .Z(n33896) );
  NANDN U34114 ( .A(n33898), .B(n33897), .Z(n33893) );
  ANDN U34115 ( .B(B[162]), .A(n66), .Z(n33554) );
  XNOR U34116 ( .A(n33562), .B(n33899), .Z(n33555) );
  XNOR U34117 ( .A(n33561), .B(n33559), .Z(n33899) );
  AND U34118 ( .A(n33900), .B(n33901), .Z(n33559) );
  NANDN U34119 ( .A(n33902), .B(n33903), .Z(n33901) );
  OR U34120 ( .A(n33904), .B(n33905), .Z(n33903) );
  NAND U34121 ( .A(n33905), .B(n33904), .Z(n33900) );
  ANDN U34122 ( .B(B[163]), .A(n67), .Z(n33561) );
  XNOR U34123 ( .A(n33569), .B(n33906), .Z(n33562) );
  XNOR U34124 ( .A(n33568), .B(n33566), .Z(n33906) );
  AND U34125 ( .A(n33907), .B(n33908), .Z(n33566) );
  NANDN U34126 ( .A(n33909), .B(n33910), .Z(n33908) );
  NANDN U34127 ( .A(n33911), .B(n33912), .Z(n33910) );
  NANDN U34128 ( .A(n33912), .B(n33911), .Z(n33907) );
  ANDN U34129 ( .B(B[164]), .A(n68), .Z(n33568) );
  XNOR U34130 ( .A(n33576), .B(n33913), .Z(n33569) );
  XNOR U34131 ( .A(n33575), .B(n33573), .Z(n33913) );
  AND U34132 ( .A(n33914), .B(n33915), .Z(n33573) );
  NANDN U34133 ( .A(n33916), .B(n33917), .Z(n33915) );
  OR U34134 ( .A(n33918), .B(n33919), .Z(n33917) );
  NAND U34135 ( .A(n33919), .B(n33918), .Z(n33914) );
  ANDN U34136 ( .B(B[165]), .A(n69), .Z(n33575) );
  XNOR U34137 ( .A(n33583), .B(n33920), .Z(n33576) );
  XNOR U34138 ( .A(n33582), .B(n33580), .Z(n33920) );
  AND U34139 ( .A(n33921), .B(n33922), .Z(n33580) );
  NANDN U34140 ( .A(n33923), .B(n33924), .Z(n33922) );
  NANDN U34141 ( .A(n33925), .B(n33926), .Z(n33924) );
  NANDN U34142 ( .A(n33926), .B(n33925), .Z(n33921) );
  ANDN U34143 ( .B(B[166]), .A(n70), .Z(n33582) );
  XNOR U34144 ( .A(n33590), .B(n33927), .Z(n33583) );
  XNOR U34145 ( .A(n33589), .B(n33587), .Z(n33927) );
  AND U34146 ( .A(n33928), .B(n33929), .Z(n33587) );
  NANDN U34147 ( .A(n33930), .B(n33931), .Z(n33929) );
  OR U34148 ( .A(n33932), .B(n33933), .Z(n33931) );
  NAND U34149 ( .A(n33933), .B(n33932), .Z(n33928) );
  ANDN U34150 ( .B(B[167]), .A(n71), .Z(n33589) );
  XNOR U34151 ( .A(n33597), .B(n33934), .Z(n33590) );
  XNOR U34152 ( .A(n33596), .B(n33594), .Z(n33934) );
  AND U34153 ( .A(n33935), .B(n33936), .Z(n33594) );
  NANDN U34154 ( .A(n33937), .B(n33938), .Z(n33936) );
  NANDN U34155 ( .A(n33939), .B(n33940), .Z(n33938) );
  NANDN U34156 ( .A(n33940), .B(n33939), .Z(n33935) );
  ANDN U34157 ( .B(B[168]), .A(n72), .Z(n33596) );
  XNOR U34158 ( .A(n33604), .B(n33941), .Z(n33597) );
  XNOR U34159 ( .A(n33603), .B(n33601), .Z(n33941) );
  AND U34160 ( .A(n33942), .B(n33943), .Z(n33601) );
  NANDN U34161 ( .A(n33944), .B(n33945), .Z(n33943) );
  OR U34162 ( .A(n33946), .B(n33947), .Z(n33945) );
  NAND U34163 ( .A(n33947), .B(n33946), .Z(n33942) );
  ANDN U34164 ( .B(B[169]), .A(n73), .Z(n33603) );
  XNOR U34165 ( .A(n33611), .B(n33948), .Z(n33604) );
  XNOR U34166 ( .A(n33610), .B(n33608), .Z(n33948) );
  AND U34167 ( .A(n33949), .B(n33950), .Z(n33608) );
  NANDN U34168 ( .A(n33951), .B(n33952), .Z(n33950) );
  NANDN U34169 ( .A(n33953), .B(n33954), .Z(n33952) );
  NANDN U34170 ( .A(n33954), .B(n33953), .Z(n33949) );
  ANDN U34171 ( .B(B[170]), .A(n74), .Z(n33610) );
  XNOR U34172 ( .A(n33618), .B(n33955), .Z(n33611) );
  XNOR U34173 ( .A(n33617), .B(n33615), .Z(n33955) );
  AND U34174 ( .A(n33956), .B(n33957), .Z(n33615) );
  NANDN U34175 ( .A(n33958), .B(n33959), .Z(n33957) );
  OR U34176 ( .A(n33960), .B(n33961), .Z(n33959) );
  NAND U34177 ( .A(n33961), .B(n33960), .Z(n33956) );
  ANDN U34178 ( .B(B[171]), .A(n75), .Z(n33617) );
  XNOR U34179 ( .A(n33625), .B(n33962), .Z(n33618) );
  XNOR U34180 ( .A(n33624), .B(n33622), .Z(n33962) );
  AND U34181 ( .A(n33963), .B(n33964), .Z(n33622) );
  NANDN U34182 ( .A(n33965), .B(n33966), .Z(n33964) );
  NANDN U34183 ( .A(n33967), .B(n33968), .Z(n33966) );
  NANDN U34184 ( .A(n33968), .B(n33967), .Z(n33963) );
  ANDN U34185 ( .B(B[172]), .A(n76), .Z(n33624) );
  XNOR U34186 ( .A(n33632), .B(n33969), .Z(n33625) );
  XNOR U34187 ( .A(n33631), .B(n33629), .Z(n33969) );
  AND U34188 ( .A(n33970), .B(n33971), .Z(n33629) );
  NANDN U34189 ( .A(n33972), .B(n33973), .Z(n33971) );
  OR U34190 ( .A(n33974), .B(n33975), .Z(n33973) );
  NAND U34191 ( .A(n33975), .B(n33974), .Z(n33970) );
  ANDN U34192 ( .B(B[173]), .A(n77), .Z(n33631) );
  XNOR U34193 ( .A(n33639), .B(n33976), .Z(n33632) );
  XNOR U34194 ( .A(n33638), .B(n33636), .Z(n33976) );
  AND U34195 ( .A(n33977), .B(n33978), .Z(n33636) );
  NANDN U34196 ( .A(n33979), .B(n33980), .Z(n33978) );
  NANDN U34197 ( .A(n33981), .B(n33982), .Z(n33980) );
  NANDN U34198 ( .A(n33982), .B(n33981), .Z(n33977) );
  ANDN U34199 ( .B(B[174]), .A(n78), .Z(n33638) );
  XNOR U34200 ( .A(n33646), .B(n33983), .Z(n33639) );
  XNOR U34201 ( .A(n33645), .B(n33643), .Z(n33983) );
  AND U34202 ( .A(n33984), .B(n33985), .Z(n33643) );
  NANDN U34203 ( .A(n33986), .B(n33987), .Z(n33985) );
  OR U34204 ( .A(n33988), .B(n33989), .Z(n33987) );
  NAND U34205 ( .A(n33989), .B(n33988), .Z(n33984) );
  ANDN U34206 ( .B(B[175]), .A(n79), .Z(n33645) );
  XNOR U34207 ( .A(n33653), .B(n33990), .Z(n33646) );
  XNOR U34208 ( .A(n33652), .B(n33650), .Z(n33990) );
  AND U34209 ( .A(n33991), .B(n33992), .Z(n33650) );
  NANDN U34210 ( .A(n33993), .B(n33994), .Z(n33992) );
  NANDN U34211 ( .A(n33995), .B(n33996), .Z(n33994) );
  NANDN U34212 ( .A(n33996), .B(n33995), .Z(n33991) );
  ANDN U34213 ( .B(B[176]), .A(n80), .Z(n33652) );
  XNOR U34214 ( .A(n33660), .B(n33997), .Z(n33653) );
  XNOR U34215 ( .A(n33659), .B(n33657), .Z(n33997) );
  AND U34216 ( .A(n33998), .B(n33999), .Z(n33657) );
  NANDN U34217 ( .A(n34000), .B(n34001), .Z(n33999) );
  OR U34218 ( .A(n34002), .B(n34003), .Z(n34001) );
  NAND U34219 ( .A(n34003), .B(n34002), .Z(n33998) );
  ANDN U34220 ( .B(B[177]), .A(n81), .Z(n33659) );
  XNOR U34221 ( .A(n33667), .B(n34004), .Z(n33660) );
  XNOR U34222 ( .A(n33666), .B(n33664), .Z(n34004) );
  AND U34223 ( .A(n34005), .B(n34006), .Z(n33664) );
  NANDN U34224 ( .A(n34007), .B(n34008), .Z(n34006) );
  NAND U34225 ( .A(n34009), .B(n34010), .Z(n34008) );
  ANDN U34226 ( .B(B[178]), .A(n82), .Z(n33666) );
  XOR U34227 ( .A(n33673), .B(n34011), .Z(n33667) );
  XNOR U34228 ( .A(n33671), .B(n33674), .Z(n34011) );
  NAND U34229 ( .A(A[2]), .B(B[179]), .Z(n33674) );
  NANDN U34230 ( .A(n34012), .B(n34013), .Z(n33671) );
  AND U34231 ( .A(A[0]), .B(B[180]), .Z(n34013) );
  XNOR U34232 ( .A(n33676), .B(n34014), .Z(n33673) );
  NAND U34233 ( .A(A[0]), .B(B[181]), .Z(n34014) );
  NAND U34234 ( .A(B[180]), .B(A[1]), .Z(n33676) );
  NAND U34235 ( .A(n34015), .B(n34016), .Z(n434) );
  NANDN U34236 ( .A(n34017), .B(n34018), .Z(n34016) );
  OR U34237 ( .A(n34019), .B(n34020), .Z(n34018) );
  NAND U34238 ( .A(n34020), .B(n34019), .Z(n34015) );
  XOR U34239 ( .A(n436), .B(n435), .Z(\A1[178] ) );
  XOR U34240 ( .A(n34020), .B(n34021), .Z(n435) );
  XNOR U34241 ( .A(n34019), .B(n34017), .Z(n34021) );
  AND U34242 ( .A(n34022), .B(n34023), .Z(n34017) );
  NANDN U34243 ( .A(n34024), .B(n34025), .Z(n34023) );
  NANDN U34244 ( .A(n34026), .B(n34027), .Z(n34025) );
  NANDN U34245 ( .A(n34027), .B(n34026), .Z(n34022) );
  ANDN U34246 ( .B(B[149]), .A(n54), .Z(n34019) );
  XNOR U34247 ( .A(n33814), .B(n34028), .Z(n34020) );
  XNOR U34248 ( .A(n33813), .B(n33811), .Z(n34028) );
  AND U34249 ( .A(n34029), .B(n34030), .Z(n33811) );
  NANDN U34250 ( .A(n34031), .B(n34032), .Z(n34030) );
  OR U34251 ( .A(n34033), .B(n34034), .Z(n34032) );
  NAND U34252 ( .A(n34034), .B(n34033), .Z(n34029) );
  ANDN U34253 ( .B(B[150]), .A(n55), .Z(n33813) );
  XNOR U34254 ( .A(n33821), .B(n34035), .Z(n33814) );
  XNOR U34255 ( .A(n33820), .B(n33818), .Z(n34035) );
  AND U34256 ( .A(n34036), .B(n34037), .Z(n33818) );
  NANDN U34257 ( .A(n34038), .B(n34039), .Z(n34037) );
  NANDN U34258 ( .A(n34040), .B(n34041), .Z(n34039) );
  NANDN U34259 ( .A(n34041), .B(n34040), .Z(n34036) );
  ANDN U34260 ( .B(B[151]), .A(n56), .Z(n33820) );
  XNOR U34261 ( .A(n33828), .B(n34042), .Z(n33821) );
  XNOR U34262 ( .A(n33827), .B(n33825), .Z(n34042) );
  AND U34263 ( .A(n34043), .B(n34044), .Z(n33825) );
  NANDN U34264 ( .A(n34045), .B(n34046), .Z(n34044) );
  OR U34265 ( .A(n34047), .B(n34048), .Z(n34046) );
  NAND U34266 ( .A(n34048), .B(n34047), .Z(n34043) );
  ANDN U34267 ( .B(B[152]), .A(n57), .Z(n33827) );
  XNOR U34268 ( .A(n33835), .B(n34049), .Z(n33828) );
  XNOR U34269 ( .A(n33834), .B(n33832), .Z(n34049) );
  AND U34270 ( .A(n34050), .B(n34051), .Z(n33832) );
  NANDN U34271 ( .A(n34052), .B(n34053), .Z(n34051) );
  NANDN U34272 ( .A(n34054), .B(n34055), .Z(n34053) );
  NANDN U34273 ( .A(n34055), .B(n34054), .Z(n34050) );
  ANDN U34274 ( .B(B[153]), .A(n58), .Z(n33834) );
  XNOR U34275 ( .A(n33842), .B(n34056), .Z(n33835) );
  XNOR U34276 ( .A(n33841), .B(n33839), .Z(n34056) );
  AND U34277 ( .A(n34057), .B(n34058), .Z(n33839) );
  NANDN U34278 ( .A(n34059), .B(n34060), .Z(n34058) );
  OR U34279 ( .A(n34061), .B(n34062), .Z(n34060) );
  NAND U34280 ( .A(n34062), .B(n34061), .Z(n34057) );
  ANDN U34281 ( .B(B[154]), .A(n59), .Z(n33841) );
  XNOR U34282 ( .A(n33849), .B(n34063), .Z(n33842) );
  XNOR U34283 ( .A(n33848), .B(n33846), .Z(n34063) );
  AND U34284 ( .A(n34064), .B(n34065), .Z(n33846) );
  NANDN U34285 ( .A(n34066), .B(n34067), .Z(n34065) );
  NANDN U34286 ( .A(n34068), .B(n34069), .Z(n34067) );
  NANDN U34287 ( .A(n34069), .B(n34068), .Z(n34064) );
  ANDN U34288 ( .B(B[155]), .A(n60), .Z(n33848) );
  XNOR U34289 ( .A(n33856), .B(n34070), .Z(n33849) );
  XNOR U34290 ( .A(n33855), .B(n33853), .Z(n34070) );
  AND U34291 ( .A(n34071), .B(n34072), .Z(n33853) );
  NANDN U34292 ( .A(n34073), .B(n34074), .Z(n34072) );
  OR U34293 ( .A(n34075), .B(n34076), .Z(n34074) );
  NAND U34294 ( .A(n34076), .B(n34075), .Z(n34071) );
  ANDN U34295 ( .B(B[156]), .A(n61), .Z(n33855) );
  XNOR U34296 ( .A(n33863), .B(n34077), .Z(n33856) );
  XNOR U34297 ( .A(n33862), .B(n33860), .Z(n34077) );
  AND U34298 ( .A(n34078), .B(n34079), .Z(n33860) );
  NANDN U34299 ( .A(n34080), .B(n34081), .Z(n34079) );
  NANDN U34300 ( .A(n34082), .B(n34083), .Z(n34081) );
  NANDN U34301 ( .A(n34083), .B(n34082), .Z(n34078) );
  ANDN U34302 ( .B(B[157]), .A(n62), .Z(n33862) );
  XNOR U34303 ( .A(n33870), .B(n34084), .Z(n33863) );
  XNOR U34304 ( .A(n33869), .B(n33867), .Z(n34084) );
  AND U34305 ( .A(n34085), .B(n34086), .Z(n33867) );
  NANDN U34306 ( .A(n34087), .B(n34088), .Z(n34086) );
  OR U34307 ( .A(n34089), .B(n34090), .Z(n34088) );
  NAND U34308 ( .A(n34090), .B(n34089), .Z(n34085) );
  ANDN U34309 ( .B(B[158]), .A(n63), .Z(n33869) );
  XNOR U34310 ( .A(n33877), .B(n34091), .Z(n33870) );
  XNOR U34311 ( .A(n33876), .B(n33874), .Z(n34091) );
  AND U34312 ( .A(n34092), .B(n34093), .Z(n33874) );
  NANDN U34313 ( .A(n34094), .B(n34095), .Z(n34093) );
  NANDN U34314 ( .A(n34096), .B(n34097), .Z(n34095) );
  NANDN U34315 ( .A(n34097), .B(n34096), .Z(n34092) );
  ANDN U34316 ( .B(B[159]), .A(n64), .Z(n33876) );
  XNOR U34317 ( .A(n33884), .B(n34098), .Z(n33877) );
  XNOR U34318 ( .A(n33883), .B(n33881), .Z(n34098) );
  AND U34319 ( .A(n34099), .B(n34100), .Z(n33881) );
  NANDN U34320 ( .A(n34101), .B(n34102), .Z(n34100) );
  OR U34321 ( .A(n34103), .B(n34104), .Z(n34102) );
  NAND U34322 ( .A(n34104), .B(n34103), .Z(n34099) );
  ANDN U34323 ( .B(B[160]), .A(n65), .Z(n33883) );
  XNOR U34324 ( .A(n33891), .B(n34105), .Z(n33884) );
  XNOR U34325 ( .A(n33890), .B(n33888), .Z(n34105) );
  AND U34326 ( .A(n34106), .B(n34107), .Z(n33888) );
  NANDN U34327 ( .A(n34108), .B(n34109), .Z(n34107) );
  NANDN U34328 ( .A(n34110), .B(n34111), .Z(n34109) );
  NANDN U34329 ( .A(n34111), .B(n34110), .Z(n34106) );
  ANDN U34330 ( .B(B[161]), .A(n66), .Z(n33890) );
  XNOR U34331 ( .A(n33898), .B(n34112), .Z(n33891) );
  XNOR U34332 ( .A(n33897), .B(n33895), .Z(n34112) );
  AND U34333 ( .A(n34113), .B(n34114), .Z(n33895) );
  NANDN U34334 ( .A(n34115), .B(n34116), .Z(n34114) );
  OR U34335 ( .A(n34117), .B(n34118), .Z(n34116) );
  NAND U34336 ( .A(n34118), .B(n34117), .Z(n34113) );
  ANDN U34337 ( .B(B[162]), .A(n67), .Z(n33897) );
  XNOR U34338 ( .A(n33905), .B(n34119), .Z(n33898) );
  XNOR U34339 ( .A(n33904), .B(n33902), .Z(n34119) );
  AND U34340 ( .A(n34120), .B(n34121), .Z(n33902) );
  NANDN U34341 ( .A(n34122), .B(n34123), .Z(n34121) );
  NANDN U34342 ( .A(n34124), .B(n34125), .Z(n34123) );
  NANDN U34343 ( .A(n34125), .B(n34124), .Z(n34120) );
  ANDN U34344 ( .B(B[163]), .A(n68), .Z(n33904) );
  XNOR U34345 ( .A(n33912), .B(n34126), .Z(n33905) );
  XNOR U34346 ( .A(n33911), .B(n33909), .Z(n34126) );
  AND U34347 ( .A(n34127), .B(n34128), .Z(n33909) );
  NANDN U34348 ( .A(n34129), .B(n34130), .Z(n34128) );
  OR U34349 ( .A(n34131), .B(n34132), .Z(n34130) );
  NAND U34350 ( .A(n34132), .B(n34131), .Z(n34127) );
  ANDN U34351 ( .B(B[164]), .A(n69), .Z(n33911) );
  XNOR U34352 ( .A(n33919), .B(n34133), .Z(n33912) );
  XNOR U34353 ( .A(n33918), .B(n33916), .Z(n34133) );
  AND U34354 ( .A(n34134), .B(n34135), .Z(n33916) );
  NANDN U34355 ( .A(n34136), .B(n34137), .Z(n34135) );
  NANDN U34356 ( .A(n34138), .B(n34139), .Z(n34137) );
  NANDN U34357 ( .A(n34139), .B(n34138), .Z(n34134) );
  ANDN U34358 ( .B(B[165]), .A(n70), .Z(n33918) );
  XNOR U34359 ( .A(n33926), .B(n34140), .Z(n33919) );
  XNOR U34360 ( .A(n33925), .B(n33923), .Z(n34140) );
  AND U34361 ( .A(n34141), .B(n34142), .Z(n33923) );
  NANDN U34362 ( .A(n34143), .B(n34144), .Z(n34142) );
  OR U34363 ( .A(n34145), .B(n34146), .Z(n34144) );
  NAND U34364 ( .A(n34146), .B(n34145), .Z(n34141) );
  ANDN U34365 ( .B(B[166]), .A(n71), .Z(n33925) );
  XNOR U34366 ( .A(n33933), .B(n34147), .Z(n33926) );
  XNOR U34367 ( .A(n33932), .B(n33930), .Z(n34147) );
  AND U34368 ( .A(n34148), .B(n34149), .Z(n33930) );
  NANDN U34369 ( .A(n34150), .B(n34151), .Z(n34149) );
  NANDN U34370 ( .A(n34152), .B(n34153), .Z(n34151) );
  NANDN U34371 ( .A(n34153), .B(n34152), .Z(n34148) );
  ANDN U34372 ( .B(B[167]), .A(n72), .Z(n33932) );
  XNOR U34373 ( .A(n33940), .B(n34154), .Z(n33933) );
  XNOR U34374 ( .A(n33939), .B(n33937), .Z(n34154) );
  AND U34375 ( .A(n34155), .B(n34156), .Z(n33937) );
  NANDN U34376 ( .A(n34157), .B(n34158), .Z(n34156) );
  OR U34377 ( .A(n34159), .B(n34160), .Z(n34158) );
  NAND U34378 ( .A(n34160), .B(n34159), .Z(n34155) );
  ANDN U34379 ( .B(B[168]), .A(n73), .Z(n33939) );
  XNOR U34380 ( .A(n33947), .B(n34161), .Z(n33940) );
  XNOR U34381 ( .A(n33946), .B(n33944), .Z(n34161) );
  AND U34382 ( .A(n34162), .B(n34163), .Z(n33944) );
  NANDN U34383 ( .A(n34164), .B(n34165), .Z(n34163) );
  NANDN U34384 ( .A(n34166), .B(n34167), .Z(n34165) );
  NANDN U34385 ( .A(n34167), .B(n34166), .Z(n34162) );
  ANDN U34386 ( .B(B[169]), .A(n74), .Z(n33946) );
  XNOR U34387 ( .A(n33954), .B(n34168), .Z(n33947) );
  XNOR U34388 ( .A(n33953), .B(n33951), .Z(n34168) );
  AND U34389 ( .A(n34169), .B(n34170), .Z(n33951) );
  NANDN U34390 ( .A(n34171), .B(n34172), .Z(n34170) );
  OR U34391 ( .A(n34173), .B(n34174), .Z(n34172) );
  NAND U34392 ( .A(n34174), .B(n34173), .Z(n34169) );
  ANDN U34393 ( .B(B[170]), .A(n75), .Z(n33953) );
  XNOR U34394 ( .A(n33961), .B(n34175), .Z(n33954) );
  XNOR U34395 ( .A(n33960), .B(n33958), .Z(n34175) );
  AND U34396 ( .A(n34176), .B(n34177), .Z(n33958) );
  NANDN U34397 ( .A(n34178), .B(n34179), .Z(n34177) );
  NANDN U34398 ( .A(n34180), .B(n34181), .Z(n34179) );
  NANDN U34399 ( .A(n34181), .B(n34180), .Z(n34176) );
  ANDN U34400 ( .B(B[171]), .A(n76), .Z(n33960) );
  XNOR U34401 ( .A(n33968), .B(n34182), .Z(n33961) );
  XNOR U34402 ( .A(n33967), .B(n33965), .Z(n34182) );
  AND U34403 ( .A(n34183), .B(n34184), .Z(n33965) );
  NANDN U34404 ( .A(n34185), .B(n34186), .Z(n34184) );
  OR U34405 ( .A(n34187), .B(n34188), .Z(n34186) );
  NAND U34406 ( .A(n34188), .B(n34187), .Z(n34183) );
  ANDN U34407 ( .B(B[172]), .A(n77), .Z(n33967) );
  XNOR U34408 ( .A(n33975), .B(n34189), .Z(n33968) );
  XNOR U34409 ( .A(n33974), .B(n33972), .Z(n34189) );
  AND U34410 ( .A(n34190), .B(n34191), .Z(n33972) );
  NANDN U34411 ( .A(n34192), .B(n34193), .Z(n34191) );
  NANDN U34412 ( .A(n34194), .B(n34195), .Z(n34193) );
  NANDN U34413 ( .A(n34195), .B(n34194), .Z(n34190) );
  ANDN U34414 ( .B(B[173]), .A(n78), .Z(n33974) );
  XNOR U34415 ( .A(n33982), .B(n34196), .Z(n33975) );
  XNOR U34416 ( .A(n33981), .B(n33979), .Z(n34196) );
  AND U34417 ( .A(n34197), .B(n34198), .Z(n33979) );
  NANDN U34418 ( .A(n34199), .B(n34200), .Z(n34198) );
  OR U34419 ( .A(n34201), .B(n34202), .Z(n34200) );
  NAND U34420 ( .A(n34202), .B(n34201), .Z(n34197) );
  ANDN U34421 ( .B(B[174]), .A(n79), .Z(n33981) );
  XNOR U34422 ( .A(n33989), .B(n34203), .Z(n33982) );
  XNOR U34423 ( .A(n33988), .B(n33986), .Z(n34203) );
  AND U34424 ( .A(n34204), .B(n34205), .Z(n33986) );
  NANDN U34425 ( .A(n34206), .B(n34207), .Z(n34205) );
  NANDN U34426 ( .A(n34208), .B(n34209), .Z(n34207) );
  NANDN U34427 ( .A(n34209), .B(n34208), .Z(n34204) );
  ANDN U34428 ( .B(B[175]), .A(n80), .Z(n33988) );
  XNOR U34429 ( .A(n33996), .B(n34210), .Z(n33989) );
  XNOR U34430 ( .A(n33995), .B(n33993), .Z(n34210) );
  AND U34431 ( .A(n34211), .B(n34212), .Z(n33993) );
  NANDN U34432 ( .A(n34213), .B(n34214), .Z(n34212) );
  OR U34433 ( .A(n34215), .B(n34216), .Z(n34214) );
  NAND U34434 ( .A(n34216), .B(n34215), .Z(n34211) );
  ANDN U34435 ( .B(B[176]), .A(n81), .Z(n33995) );
  XNOR U34436 ( .A(n34003), .B(n34217), .Z(n33996) );
  XNOR U34437 ( .A(n34002), .B(n34000), .Z(n34217) );
  AND U34438 ( .A(n34218), .B(n34219), .Z(n34000) );
  NANDN U34439 ( .A(n34220), .B(n34221), .Z(n34219) );
  NAND U34440 ( .A(n34222), .B(n34223), .Z(n34221) );
  ANDN U34441 ( .B(B[177]), .A(n82), .Z(n34002) );
  XOR U34442 ( .A(n34009), .B(n34224), .Z(n34003) );
  XNOR U34443 ( .A(n34007), .B(n34010), .Z(n34224) );
  NAND U34444 ( .A(A[2]), .B(B[178]), .Z(n34010) );
  NANDN U34445 ( .A(n34225), .B(n34226), .Z(n34007) );
  AND U34446 ( .A(A[0]), .B(B[179]), .Z(n34226) );
  XNOR U34447 ( .A(n34012), .B(n34227), .Z(n34009) );
  NAND U34448 ( .A(A[0]), .B(B[180]), .Z(n34227) );
  NAND U34449 ( .A(B[179]), .B(A[1]), .Z(n34012) );
  NAND U34450 ( .A(n34228), .B(n34229), .Z(n436) );
  NANDN U34451 ( .A(n34230), .B(n34231), .Z(n34229) );
  OR U34452 ( .A(n34232), .B(n34233), .Z(n34231) );
  NAND U34453 ( .A(n34233), .B(n34232), .Z(n34228) );
  XOR U34454 ( .A(n438), .B(n437), .Z(\A1[177] ) );
  XOR U34455 ( .A(n34233), .B(n34234), .Z(n437) );
  XNOR U34456 ( .A(n34232), .B(n34230), .Z(n34234) );
  AND U34457 ( .A(n34235), .B(n34236), .Z(n34230) );
  NANDN U34458 ( .A(n34237), .B(n34238), .Z(n34236) );
  NANDN U34459 ( .A(n34239), .B(n34240), .Z(n34238) );
  NANDN U34460 ( .A(n34240), .B(n34239), .Z(n34235) );
  ANDN U34461 ( .B(B[148]), .A(n54), .Z(n34232) );
  XNOR U34462 ( .A(n34027), .B(n34241), .Z(n34233) );
  XNOR U34463 ( .A(n34026), .B(n34024), .Z(n34241) );
  AND U34464 ( .A(n34242), .B(n34243), .Z(n34024) );
  NANDN U34465 ( .A(n34244), .B(n34245), .Z(n34243) );
  OR U34466 ( .A(n34246), .B(n34247), .Z(n34245) );
  NAND U34467 ( .A(n34247), .B(n34246), .Z(n34242) );
  ANDN U34468 ( .B(B[149]), .A(n55), .Z(n34026) );
  XNOR U34469 ( .A(n34034), .B(n34248), .Z(n34027) );
  XNOR U34470 ( .A(n34033), .B(n34031), .Z(n34248) );
  AND U34471 ( .A(n34249), .B(n34250), .Z(n34031) );
  NANDN U34472 ( .A(n34251), .B(n34252), .Z(n34250) );
  NANDN U34473 ( .A(n34253), .B(n34254), .Z(n34252) );
  NANDN U34474 ( .A(n34254), .B(n34253), .Z(n34249) );
  ANDN U34475 ( .B(B[150]), .A(n56), .Z(n34033) );
  XNOR U34476 ( .A(n34041), .B(n34255), .Z(n34034) );
  XNOR U34477 ( .A(n34040), .B(n34038), .Z(n34255) );
  AND U34478 ( .A(n34256), .B(n34257), .Z(n34038) );
  NANDN U34479 ( .A(n34258), .B(n34259), .Z(n34257) );
  OR U34480 ( .A(n34260), .B(n34261), .Z(n34259) );
  NAND U34481 ( .A(n34261), .B(n34260), .Z(n34256) );
  ANDN U34482 ( .B(B[151]), .A(n57), .Z(n34040) );
  XNOR U34483 ( .A(n34048), .B(n34262), .Z(n34041) );
  XNOR U34484 ( .A(n34047), .B(n34045), .Z(n34262) );
  AND U34485 ( .A(n34263), .B(n34264), .Z(n34045) );
  NANDN U34486 ( .A(n34265), .B(n34266), .Z(n34264) );
  NANDN U34487 ( .A(n34267), .B(n34268), .Z(n34266) );
  NANDN U34488 ( .A(n34268), .B(n34267), .Z(n34263) );
  ANDN U34489 ( .B(B[152]), .A(n58), .Z(n34047) );
  XNOR U34490 ( .A(n34055), .B(n34269), .Z(n34048) );
  XNOR U34491 ( .A(n34054), .B(n34052), .Z(n34269) );
  AND U34492 ( .A(n34270), .B(n34271), .Z(n34052) );
  NANDN U34493 ( .A(n34272), .B(n34273), .Z(n34271) );
  OR U34494 ( .A(n34274), .B(n34275), .Z(n34273) );
  NAND U34495 ( .A(n34275), .B(n34274), .Z(n34270) );
  ANDN U34496 ( .B(B[153]), .A(n59), .Z(n34054) );
  XNOR U34497 ( .A(n34062), .B(n34276), .Z(n34055) );
  XNOR U34498 ( .A(n34061), .B(n34059), .Z(n34276) );
  AND U34499 ( .A(n34277), .B(n34278), .Z(n34059) );
  NANDN U34500 ( .A(n34279), .B(n34280), .Z(n34278) );
  NANDN U34501 ( .A(n34281), .B(n34282), .Z(n34280) );
  NANDN U34502 ( .A(n34282), .B(n34281), .Z(n34277) );
  ANDN U34503 ( .B(B[154]), .A(n60), .Z(n34061) );
  XNOR U34504 ( .A(n34069), .B(n34283), .Z(n34062) );
  XNOR U34505 ( .A(n34068), .B(n34066), .Z(n34283) );
  AND U34506 ( .A(n34284), .B(n34285), .Z(n34066) );
  NANDN U34507 ( .A(n34286), .B(n34287), .Z(n34285) );
  OR U34508 ( .A(n34288), .B(n34289), .Z(n34287) );
  NAND U34509 ( .A(n34289), .B(n34288), .Z(n34284) );
  ANDN U34510 ( .B(B[155]), .A(n61), .Z(n34068) );
  XNOR U34511 ( .A(n34076), .B(n34290), .Z(n34069) );
  XNOR U34512 ( .A(n34075), .B(n34073), .Z(n34290) );
  AND U34513 ( .A(n34291), .B(n34292), .Z(n34073) );
  NANDN U34514 ( .A(n34293), .B(n34294), .Z(n34292) );
  NANDN U34515 ( .A(n34295), .B(n34296), .Z(n34294) );
  NANDN U34516 ( .A(n34296), .B(n34295), .Z(n34291) );
  ANDN U34517 ( .B(B[156]), .A(n62), .Z(n34075) );
  XNOR U34518 ( .A(n34083), .B(n34297), .Z(n34076) );
  XNOR U34519 ( .A(n34082), .B(n34080), .Z(n34297) );
  AND U34520 ( .A(n34298), .B(n34299), .Z(n34080) );
  NANDN U34521 ( .A(n34300), .B(n34301), .Z(n34299) );
  OR U34522 ( .A(n34302), .B(n34303), .Z(n34301) );
  NAND U34523 ( .A(n34303), .B(n34302), .Z(n34298) );
  ANDN U34524 ( .B(B[157]), .A(n63), .Z(n34082) );
  XNOR U34525 ( .A(n34090), .B(n34304), .Z(n34083) );
  XNOR U34526 ( .A(n34089), .B(n34087), .Z(n34304) );
  AND U34527 ( .A(n34305), .B(n34306), .Z(n34087) );
  NANDN U34528 ( .A(n34307), .B(n34308), .Z(n34306) );
  NANDN U34529 ( .A(n34309), .B(n34310), .Z(n34308) );
  NANDN U34530 ( .A(n34310), .B(n34309), .Z(n34305) );
  ANDN U34531 ( .B(B[158]), .A(n64), .Z(n34089) );
  XNOR U34532 ( .A(n34097), .B(n34311), .Z(n34090) );
  XNOR U34533 ( .A(n34096), .B(n34094), .Z(n34311) );
  AND U34534 ( .A(n34312), .B(n34313), .Z(n34094) );
  NANDN U34535 ( .A(n34314), .B(n34315), .Z(n34313) );
  OR U34536 ( .A(n34316), .B(n34317), .Z(n34315) );
  NAND U34537 ( .A(n34317), .B(n34316), .Z(n34312) );
  ANDN U34538 ( .B(B[159]), .A(n65), .Z(n34096) );
  XNOR U34539 ( .A(n34104), .B(n34318), .Z(n34097) );
  XNOR U34540 ( .A(n34103), .B(n34101), .Z(n34318) );
  AND U34541 ( .A(n34319), .B(n34320), .Z(n34101) );
  NANDN U34542 ( .A(n34321), .B(n34322), .Z(n34320) );
  NANDN U34543 ( .A(n34323), .B(n34324), .Z(n34322) );
  NANDN U34544 ( .A(n34324), .B(n34323), .Z(n34319) );
  ANDN U34545 ( .B(B[160]), .A(n66), .Z(n34103) );
  XNOR U34546 ( .A(n34111), .B(n34325), .Z(n34104) );
  XNOR U34547 ( .A(n34110), .B(n34108), .Z(n34325) );
  AND U34548 ( .A(n34326), .B(n34327), .Z(n34108) );
  NANDN U34549 ( .A(n34328), .B(n34329), .Z(n34327) );
  OR U34550 ( .A(n34330), .B(n34331), .Z(n34329) );
  NAND U34551 ( .A(n34331), .B(n34330), .Z(n34326) );
  ANDN U34552 ( .B(B[161]), .A(n67), .Z(n34110) );
  XNOR U34553 ( .A(n34118), .B(n34332), .Z(n34111) );
  XNOR U34554 ( .A(n34117), .B(n34115), .Z(n34332) );
  AND U34555 ( .A(n34333), .B(n34334), .Z(n34115) );
  NANDN U34556 ( .A(n34335), .B(n34336), .Z(n34334) );
  NANDN U34557 ( .A(n34337), .B(n34338), .Z(n34336) );
  NANDN U34558 ( .A(n34338), .B(n34337), .Z(n34333) );
  ANDN U34559 ( .B(B[162]), .A(n68), .Z(n34117) );
  XNOR U34560 ( .A(n34125), .B(n34339), .Z(n34118) );
  XNOR U34561 ( .A(n34124), .B(n34122), .Z(n34339) );
  AND U34562 ( .A(n34340), .B(n34341), .Z(n34122) );
  NANDN U34563 ( .A(n34342), .B(n34343), .Z(n34341) );
  OR U34564 ( .A(n34344), .B(n34345), .Z(n34343) );
  NAND U34565 ( .A(n34345), .B(n34344), .Z(n34340) );
  ANDN U34566 ( .B(B[163]), .A(n69), .Z(n34124) );
  XNOR U34567 ( .A(n34132), .B(n34346), .Z(n34125) );
  XNOR U34568 ( .A(n34131), .B(n34129), .Z(n34346) );
  AND U34569 ( .A(n34347), .B(n34348), .Z(n34129) );
  NANDN U34570 ( .A(n34349), .B(n34350), .Z(n34348) );
  NANDN U34571 ( .A(n34351), .B(n34352), .Z(n34350) );
  NANDN U34572 ( .A(n34352), .B(n34351), .Z(n34347) );
  ANDN U34573 ( .B(B[164]), .A(n70), .Z(n34131) );
  XNOR U34574 ( .A(n34139), .B(n34353), .Z(n34132) );
  XNOR U34575 ( .A(n34138), .B(n34136), .Z(n34353) );
  AND U34576 ( .A(n34354), .B(n34355), .Z(n34136) );
  NANDN U34577 ( .A(n34356), .B(n34357), .Z(n34355) );
  OR U34578 ( .A(n34358), .B(n34359), .Z(n34357) );
  NAND U34579 ( .A(n34359), .B(n34358), .Z(n34354) );
  ANDN U34580 ( .B(B[165]), .A(n71), .Z(n34138) );
  XNOR U34581 ( .A(n34146), .B(n34360), .Z(n34139) );
  XNOR U34582 ( .A(n34145), .B(n34143), .Z(n34360) );
  AND U34583 ( .A(n34361), .B(n34362), .Z(n34143) );
  NANDN U34584 ( .A(n34363), .B(n34364), .Z(n34362) );
  NANDN U34585 ( .A(n34365), .B(n34366), .Z(n34364) );
  NANDN U34586 ( .A(n34366), .B(n34365), .Z(n34361) );
  ANDN U34587 ( .B(B[166]), .A(n72), .Z(n34145) );
  XNOR U34588 ( .A(n34153), .B(n34367), .Z(n34146) );
  XNOR U34589 ( .A(n34152), .B(n34150), .Z(n34367) );
  AND U34590 ( .A(n34368), .B(n34369), .Z(n34150) );
  NANDN U34591 ( .A(n34370), .B(n34371), .Z(n34369) );
  OR U34592 ( .A(n34372), .B(n34373), .Z(n34371) );
  NAND U34593 ( .A(n34373), .B(n34372), .Z(n34368) );
  ANDN U34594 ( .B(B[167]), .A(n73), .Z(n34152) );
  XNOR U34595 ( .A(n34160), .B(n34374), .Z(n34153) );
  XNOR U34596 ( .A(n34159), .B(n34157), .Z(n34374) );
  AND U34597 ( .A(n34375), .B(n34376), .Z(n34157) );
  NANDN U34598 ( .A(n34377), .B(n34378), .Z(n34376) );
  NANDN U34599 ( .A(n34379), .B(n34380), .Z(n34378) );
  NANDN U34600 ( .A(n34380), .B(n34379), .Z(n34375) );
  ANDN U34601 ( .B(B[168]), .A(n74), .Z(n34159) );
  XNOR U34602 ( .A(n34167), .B(n34381), .Z(n34160) );
  XNOR U34603 ( .A(n34166), .B(n34164), .Z(n34381) );
  AND U34604 ( .A(n34382), .B(n34383), .Z(n34164) );
  NANDN U34605 ( .A(n34384), .B(n34385), .Z(n34383) );
  OR U34606 ( .A(n34386), .B(n34387), .Z(n34385) );
  NAND U34607 ( .A(n34387), .B(n34386), .Z(n34382) );
  ANDN U34608 ( .B(B[169]), .A(n75), .Z(n34166) );
  XNOR U34609 ( .A(n34174), .B(n34388), .Z(n34167) );
  XNOR U34610 ( .A(n34173), .B(n34171), .Z(n34388) );
  AND U34611 ( .A(n34389), .B(n34390), .Z(n34171) );
  NANDN U34612 ( .A(n34391), .B(n34392), .Z(n34390) );
  NANDN U34613 ( .A(n34393), .B(n34394), .Z(n34392) );
  NANDN U34614 ( .A(n34394), .B(n34393), .Z(n34389) );
  ANDN U34615 ( .B(B[170]), .A(n76), .Z(n34173) );
  XNOR U34616 ( .A(n34181), .B(n34395), .Z(n34174) );
  XNOR U34617 ( .A(n34180), .B(n34178), .Z(n34395) );
  AND U34618 ( .A(n34396), .B(n34397), .Z(n34178) );
  NANDN U34619 ( .A(n34398), .B(n34399), .Z(n34397) );
  OR U34620 ( .A(n34400), .B(n34401), .Z(n34399) );
  NAND U34621 ( .A(n34401), .B(n34400), .Z(n34396) );
  ANDN U34622 ( .B(B[171]), .A(n77), .Z(n34180) );
  XNOR U34623 ( .A(n34188), .B(n34402), .Z(n34181) );
  XNOR U34624 ( .A(n34187), .B(n34185), .Z(n34402) );
  AND U34625 ( .A(n34403), .B(n34404), .Z(n34185) );
  NANDN U34626 ( .A(n34405), .B(n34406), .Z(n34404) );
  NANDN U34627 ( .A(n34407), .B(n34408), .Z(n34406) );
  NANDN U34628 ( .A(n34408), .B(n34407), .Z(n34403) );
  ANDN U34629 ( .B(B[172]), .A(n78), .Z(n34187) );
  XNOR U34630 ( .A(n34195), .B(n34409), .Z(n34188) );
  XNOR U34631 ( .A(n34194), .B(n34192), .Z(n34409) );
  AND U34632 ( .A(n34410), .B(n34411), .Z(n34192) );
  NANDN U34633 ( .A(n34412), .B(n34413), .Z(n34411) );
  OR U34634 ( .A(n34414), .B(n34415), .Z(n34413) );
  NAND U34635 ( .A(n34415), .B(n34414), .Z(n34410) );
  ANDN U34636 ( .B(B[173]), .A(n79), .Z(n34194) );
  XNOR U34637 ( .A(n34202), .B(n34416), .Z(n34195) );
  XNOR U34638 ( .A(n34201), .B(n34199), .Z(n34416) );
  AND U34639 ( .A(n34417), .B(n34418), .Z(n34199) );
  NANDN U34640 ( .A(n34419), .B(n34420), .Z(n34418) );
  NANDN U34641 ( .A(n34421), .B(n34422), .Z(n34420) );
  NANDN U34642 ( .A(n34422), .B(n34421), .Z(n34417) );
  ANDN U34643 ( .B(B[174]), .A(n80), .Z(n34201) );
  XNOR U34644 ( .A(n34209), .B(n34423), .Z(n34202) );
  XNOR U34645 ( .A(n34208), .B(n34206), .Z(n34423) );
  AND U34646 ( .A(n34424), .B(n34425), .Z(n34206) );
  NANDN U34647 ( .A(n34426), .B(n34427), .Z(n34425) );
  OR U34648 ( .A(n34428), .B(n34429), .Z(n34427) );
  NAND U34649 ( .A(n34429), .B(n34428), .Z(n34424) );
  ANDN U34650 ( .B(B[175]), .A(n81), .Z(n34208) );
  XNOR U34651 ( .A(n34216), .B(n34430), .Z(n34209) );
  XNOR U34652 ( .A(n34215), .B(n34213), .Z(n34430) );
  AND U34653 ( .A(n34431), .B(n34432), .Z(n34213) );
  NANDN U34654 ( .A(n34433), .B(n34434), .Z(n34432) );
  NAND U34655 ( .A(n34435), .B(n34436), .Z(n34434) );
  ANDN U34656 ( .B(B[176]), .A(n82), .Z(n34215) );
  XOR U34657 ( .A(n34222), .B(n34437), .Z(n34216) );
  XNOR U34658 ( .A(n34220), .B(n34223), .Z(n34437) );
  NAND U34659 ( .A(A[2]), .B(B[177]), .Z(n34223) );
  NANDN U34660 ( .A(n34438), .B(n34439), .Z(n34220) );
  AND U34661 ( .A(A[0]), .B(B[178]), .Z(n34439) );
  XNOR U34662 ( .A(n34225), .B(n34440), .Z(n34222) );
  NAND U34663 ( .A(A[0]), .B(B[179]), .Z(n34440) );
  NAND U34664 ( .A(B[178]), .B(A[1]), .Z(n34225) );
  NAND U34665 ( .A(n34441), .B(n34442), .Z(n438) );
  NANDN U34666 ( .A(n34443), .B(n34444), .Z(n34442) );
  OR U34667 ( .A(n34445), .B(n34446), .Z(n34444) );
  NAND U34668 ( .A(n34446), .B(n34445), .Z(n34441) );
  XOR U34669 ( .A(n440), .B(n439), .Z(\A1[176] ) );
  XOR U34670 ( .A(n34446), .B(n34447), .Z(n439) );
  XNOR U34671 ( .A(n34445), .B(n34443), .Z(n34447) );
  AND U34672 ( .A(n34448), .B(n34449), .Z(n34443) );
  NANDN U34673 ( .A(n34450), .B(n34451), .Z(n34449) );
  NANDN U34674 ( .A(n34452), .B(n34453), .Z(n34451) );
  NANDN U34675 ( .A(n34453), .B(n34452), .Z(n34448) );
  ANDN U34676 ( .B(B[147]), .A(n54), .Z(n34445) );
  XNOR U34677 ( .A(n34240), .B(n34454), .Z(n34446) );
  XNOR U34678 ( .A(n34239), .B(n34237), .Z(n34454) );
  AND U34679 ( .A(n34455), .B(n34456), .Z(n34237) );
  NANDN U34680 ( .A(n34457), .B(n34458), .Z(n34456) );
  OR U34681 ( .A(n34459), .B(n34460), .Z(n34458) );
  NAND U34682 ( .A(n34460), .B(n34459), .Z(n34455) );
  ANDN U34683 ( .B(B[148]), .A(n55), .Z(n34239) );
  XNOR U34684 ( .A(n34247), .B(n34461), .Z(n34240) );
  XNOR U34685 ( .A(n34246), .B(n34244), .Z(n34461) );
  AND U34686 ( .A(n34462), .B(n34463), .Z(n34244) );
  NANDN U34687 ( .A(n34464), .B(n34465), .Z(n34463) );
  NANDN U34688 ( .A(n34466), .B(n34467), .Z(n34465) );
  NANDN U34689 ( .A(n34467), .B(n34466), .Z(n34462) );
  ANDN U34690 ( .B(B[149]), .A(n56), .Z(n34246) );
  XNOR U34691 ( .A(n34254), .B(n34468), .Z(n34247) );
  XNOR U34692 ( .A(n34253), .B(n34251), .Z(n34468) );
  AND U34693 ( .A(n34469), .B(n34470), .Z(n34251) );
  NANDN U34694 ( .A(n34471), .B(n34472), .Z(n34470) );
  OR U34695 ( .A(n34473), .B(n34474), .Z(n34472) );
  NAND U34696 ( .A(n34474), .B(n34473), .Z(n34469) );
  ANDN U34697 ( .B(B[150]), .A(n57), .Z(n34253) );
  XNOR U34698 ( .A(n34261), .B(n34475), .Z(n34254) );
  XNOR U34699 ( .A(n34260), .B(n34258), .Z(n34475) );
  AND U34700 ( .A(n34476), .B(n34477), .Z(n34258) );
  NANDN U34701 ( .A(n34478), .B(n34479), .Z(n34477) );
  NANDN U34702 ( .A(n34480), .B(n34481), .Z(n34479) );
  NANDN U34703 ( .A(n34481), .B(n34480), .Z(n34476) );
  ANDN U34704 ( .B(B[151]), .A(n58), .Z(n34260) );
  XNOR U34705 ( .A(n34268), .B(n34482), .Z(n34261) );
  XNOR U34706 ( .A(n34267), .B(n34265), .Z(n34482) );
  AND U34707 ( .A(n34483), .B(n34484), .Z(n34265) );
  NANDN U34708 ( .A(n34485), .B(n34486), .Z(n34484) );
  OR U34709 ( .A(n34487), .B(n34488), .Z(n34486) );
  NAND U34710 ( .A(n34488), .B(n34487), .Z(n34483) );
  ANDN U34711 ( .B(B[152]), .A(n59), .Z(n34267) );
  XNOR U34712 ( .A(n34275), .B(n34489), .Z(n34268) );
  XNOR U34713 ( .A(n34274), .B(n34272), .Z(n34489) );
  AND U34714 ( .A(n34490), .B(n34491), .Z(n34272) );
  NANDN U34715 ( .A(n34492), .B(n34493), .Z(n34491) );
  NANDN U34716 ( .A(n34494), .B(n34495), .Z(n34493) );
  NANDN U34717 ( .A(n34495), .B(n34494), .Z(n34490) );
  ANDN U34718 ( .B(B[153]), .A(n60), .Z(n34274) );
  XNOR U34719 ( .A(n34282), .B(n34496), .Z(n34275) );
  XNOR U34720 ( .A(n34281), .B(n34279), .Z(n34496) );
  AND U34721 ( .A(n34497), .B(n34498), .Z(n34279) );
  NANDN U34722 ( .A(n34499), .B(n34500), .Z(n34498) );
  OR U34723 ( .A(n34501), .B(n34502), .Z(n34500) );
  NAND U34724 ( .A(n34502), .B(n34501), .Z(n34497) );
  ANDN U34725 ( .B(B[154]), .A(n61), .Z(n34281) );
  XNOR U34726 ( .A(n34289), .B(n34503), .Z(n34282) );
  XNOR U34727 ( .A(n34288), .B(n34286), .Z(n34503) );
  AND U34728 ( .A(n34504), .B(n34505), .Z(n34286) );
  NANDN U34729 ( .A(n34506), .B(n34507), .Z(n34505) );
  NANDN U34730 ( .A(n34508), .B(n34509), .Z(n34507) );
  NANDN U34731 ( .A(n34509), .B(n34508), .Z(n34504) );
  ANDN U34732 ( .B(B[155]), .A(n62), .Z(n34288) );
  XNOR U34733 ( .A(n34296), .B(n34510), .Z(n34289) );
  XNOR U34734 ( .A(n34295), .B(n34293), .Z(n34510) );
  AND U34735 ( .A(n34511), .B(n34512), .Z(n34293) );
  NANDN U34736 ( .A(n34513), .B(n34514), .Z(n34512) );
  OR U34737 ( .A(n34515), .B(n34516), .Z(n34514) );
  NAND U34738 ( .A(n34516), .B(n34515), .Z(n34511) );
  ANDN U34739 ( .B(B[156]), .A(n63), .Z(n34295) );
  XNOR U34740 ( .A(n34303), .B(n34517), .Z(n34296) );
  XNOR U34741 ( .A(n34302), .B(n34300), .Z(n34517) );
  AND U34742 ( .A(n34518), .B(n34519), .Z(n34300) );
  NANDN U34743 ( .A(n34520), .B(n34521), .Z(n34519) );
  NANDN U34744 ( .A(n34522), .B(n34523), .Z(n34521) );
  NANDN U34745 ( .A(n34523), .B(n34522), .Z(n34518) );
  ANDN U34746 ( .B(B[157]), .A(n64), .Z(n34302) );
  XNOR U34747 ( .A(n34310), .B(n34524), .Z(n34303) );
  XNOR U34748 ( .A(n34309), .B(n34307), .Z(n34524) );
  AND U34749 ( .A(n34525), .B(n34526), .Z(n34307) );
  NANDN U34750 ( .A(n34527), .B(n34528), .Z(n34526) );
  OR U34751 ( .A(n34529), .B(n34530), .Z(n34528) );
  NAND U34752 ( .A(n34530), .B(n34529), .Z(n34525) );
  ANDN U34753 ( .B(B[158]), .A(n65), .Z(n34309) );
  XNOR U34754 ( .A(n34317), .B(n34531), .Z(n34310) );
  XNOR U34755 ( .A(n34316), .B(n34314), .Z(n34531) );
  AND U34756 ( .A(n34532), .B(n34533), .Z(n34314) );
  NANDN U34757 ( .A(n34534), .B(n34535), .Z(n34533) );
  NANDN U34758 ( .A(n34536), .B(n34537), .Z(n34535) );
  NANDN U34759 ( .A(n34537), .B(n34536), .Z(n34532) );
  ANDN U34760 ( .B(B[159]), .A(n66), .Z(n34316) );
  XNOR U34761 ( .A(n34324), .B(n34538), .Z(n34317) );
  XNOR U34762 ( .A(n34323), .B(n34321), .Z(n34538) );
  AND U34763 ( .A(n34539), .B(n34540), .Z(n34321) );
  NANDN U34764 ( .A(n34541), .B(n34542), .Z(n34540) );
  OR U34765 ( .A(n34543), .B(n34544), .Z(n34542) );
  NAND U34766 ( .A(n34544), .B(n34543), .Z(n34539) );
  ANDN U34767 ( .B(B[160]), .A(n67), .Z(n34323) );
  XNOR U34768 ( .A(n34331), .B(n34545), .Z(n34324) );
  XNOR U34769 ( .A(n34330), .B(n34328), .Z(n34545) );
  AND U34770 ( .A(n34546), .B(n34547), .Z(n34328) );
  NANDN U34771 ( .A(n34548), .B(n34549), .Z(n34547) );
  NANDN U34772 ( .A(n34550), .B(n34551), .Z(n34549) );
  NANDN U34773 ( .A(n34551), .B(n34550), .Z(n34546) );
  ANDN U34774 ( .B(B[161]), .A(n68), .Z(n34330) );
  XNOR U34775 ( .A(n34338), .B(n34552), .Z(n34331) );
  XNOR U34776 ( .A(n34337), .B(n34335), .Z(n34552) );
  AND U34777 ( .A(n34553), .B(n34554), .Z(n34335) );
  NANDN U34778 ( .A(n34555), .B(n34556), .Z(n34554) );
  OR U34779 ( .A(n34557), .B(n34558), .Z(n34556) );
  NAND U34780 ( .A(n34558), .B(n34557), .Z(n34553) );
  ANDN U34781 ( .B(B[162]), .A(n69), .Z(n34337) );
  XNOR U34782 ( .A(n34345), .B(n34559), .Z(n34338) );
  XNOR U34783 ( .A(n34344), .B(n34342), .Z(n34559) );
  AND U34784 ( .A(n34560), .B(n34561), .Z(n34342) );
  NANDN U34785 ( .A(n34562), .B(n34563), .Z(n34561) );
  NANDN U34786 ( .A(n34564), .B(n34565), .Z(n34563) );
  NANDN U34787 ( .A(n34565), .B(n34564), .Z(n34560) );
  ANDN U34788 ( .B(B[163]), .A(n70), .Z(n34344) );
  XNOR U34789 ( .A(n34352), .B(n34566), .Z(n34345) );
  XNOR U34790 ( .A(n34351), .B(n34349), .Z(n34566) );
  AND U34791 ( .A(n34567), .B(n34568), .Z(n34349) );
  NANDN U34792 ( .A(n34569), .B(n34570), .Z(n34568) );
  OR U34793 ( .A(n34571), .B(n34572), .Z(n34570) );
  NAND U34794 ( .A(n34572), .B(n34571), .Z(n34567) );
  ANDN U34795 ( .B(B[164]), .A(n71), .Z(n34351) );
  XNOR U34796 ( .A(n34359), .B(n34573), .Z(n34352) );
  XNOR U34797 ( .A(n34358), .B(n34356), .Z(n34573) );
  AND U34798 ( .A(n34574), .B(n34575), .Z(n34356) );
  NANDN U34799 ( .A(n34576), .B(n34577), .Z(n34575) );
  NANDN U34800 ( .A(n34578), .B(n34579), .Z(n34577) );
  NANDN U34801 ( .A(n34579), .B(n34578), .Z(n34574) );
  ANDN U34802 ( .B(B[165]), .A(n72), .Z(n34358) );
  XNOR U34803 ( .A(n34366), .B(n34580), .Z(n34359) );
  XNOR U34804 ( .A(n34365), .B(n34363), .Z(n34580) );
  AND U34805 ( .A(n34581), .B(n34582), .Z(n34363) );
  NANDN U34806 ( .A(n34583), .B(n34584), .Z(n34582) );
  OR U34807 ( .A(n34585), .B(n34586), .Z(n34584) );
  NAND U34808 ( .A(n34586), .B(n34585), .Z(n34581) );
  ANDN U34809 ( .B(B[166]), .A(n73), .Z(n34365) );
  XNOR U34810 ( .A(n34373), .B(n34587), .Z(n34366) );
  XNOR U34811 ( .A(n34372), .B(n34370), .Z(n34587) );
  AND U34812 ( .A(n34588), .B(n34589), .Z(n34370) );
  NANDN U34813 ( .A(n34590), .B(n34591), .Z(n34589) );
  NANDN U34814 ( .A(n34592), .B(n34593), .Z(n34591) );
  NANDN U34815 ( .A(n34593), .B(n34592), .Z(n34588) );
  ANDN U34816 ( .B(B[167]), .A(n74), .Z(n34372) );
  XNOR U34817 ( .A(n34380), .B(n34594), .Z(n34373) );
  XNOR U34818 ( .A(n34379), .B(n34377), .Z(n34594) );
  AND U34819 ( .A(n34595), .B(n34596), .Z(n34377) );
  NANDN U34820 ( .A(n34597), .B(n34598), .Z(n34596) );
  OR U34821 ( .A(n34599), .B(n34600), .Z(n34598) );
  NAND U34822 ( .A(n34600), .B(n34599), .Z(n34595) );
  ANDN U34823 ( .B(B[168]), .A(n75), .Z(n34379) );
  XNOR U34824 ( .A(n34387), .B(n34601), .Z(n34380) );
  XNOR U34825 ( .A(n34386), .B(n34384), .Z(n34601) );
  AND U34826 ( .A(n34602), .B(n34603), .Z(n34384) );
  NANDN U34827 ( .A(n34604), .B(n34605), .Z(n34603) );
  NANDN U34828 ( .A(n34606), .B(n34607), .Z(n34605) );
  NANDN U34829 ( .A(n34607), .B(n34606), .Z(n34602) );
  ANDN U34830 ( .B(B[169]), .A(n76), .Z(n34386) );
  XNOR U34831 ( .A(n34394), .B(n34608), .Z(n34387) );
  XNOR U34832 ( .A(n34393), .B(n34391), .Z(n34608) );
  AND U34833 ( .A(n34609), .B(n34610), .Z(n34391) );
  NANDN U34834 ( .A(n34611), .B(n34612), .Z(n34610) );
  OR U34835 ( .A(n34613), .B(n34614), .Z(n34612) );
  NAND U34836 ( .A(n34614), .B(n34613), .Z(n34609) );
  ANDN U34837 ( .B(B[170]), .A(n77), .Z(n34393) );
  XNOR U34838 ( .A(n34401), .B(n34615), .Z(n34394) );
  XNOR U34839 ( .A(n34400), .B(n34398), .Z(n34615) );
  AND U34840 ( .A(n34616), .B(n34617), .Z(n34398) );
  NANDN U34841 ( .A(n34618), .B(n34619), .Z(n34617) );
  NANDN U34842 ( .A(n34620), .B(n34621), .Z(n34619) );
  NANDN U34843 ( .A(n34621), .B(n34620), .Z(n34616) );
  ANDN U34844 ( .B(B[171]), .A(n78), .Z(n34400) );
  XNOR U34845 ( .A(n34408), .B(n34622), .Z(n34401) );
  XNOR U34846 ( .A(n34407), .B(n34405), .Z(n34622) );
  AND U34847 ( .A(n34623), .B(n34624), .Z(n34405) );
  NANDN U34848 ( .A(n34625), .B(n34626), .Z(n34624) );
  OR U34849 ( .A(n34627), .B(n34628), .Z(n34626) );
  NAND U34850 ( .A(n34628), .B(n34627), .Z(n34623) );
  ANDN U34851 ( .B(B[172]), .A(n79), .Z(n34407) );
  XNOR U34852 ( .A(n34415), .B(n34629), .Z(n34408) );
  XNOR U34853 ( .A(n34414), .B(n34412), .Z(n34629) );
  AND U34854 ( .A(n34630), .B(n34631), .Z(n34412) );
  NANDN U34855 ( .A(n34632), .B(n34633), .Z(n34631) );
  NANDN U34856 ( .A(n34634), .B(n34635), .Z(n34633) );
  NANDN U34857 ( .A(n34635), .B(n34634), .Z(n34630) );
  ANDN U34858 ( .B(B[173]), .A(n80), .Z(n34414) );
  XNOR U34859 ( .A(n34422), .B(n34636), .Z(n34415) );
  XNOR U34860 ( .A(n34421), .B(n34419), .Z(n34636) );
  AND U34861 ( .A(n34637), .B(n34638), .Z(n34419) );
  NANDN U34862 ( .A(n34639), .B(n34640), .Z(n34638) );
  OR U34863 ( .A(n34641), .B(n34642), .Z(n34640) );
  NAND U34864 ( .A(n34642), .B(n34641), .Z(n34637) );
  ANDN U34865 ( .B(B[174]), .A(n81), .Z(n34421) );
  XNOR U34866 ( .A(n34429), .B(n34643), .Z(n34422) );
  XNOR U34867 ( .A(n34428), .B(n34426), .Z(n34643) );
  AND U34868 ( .A(n34644), .B(n34645), .Z(n34426) );
  NANDN U34869 ( .A(n34646), .B(n34647), .Z(n34645) );
  NAND U34870 ( .A(n34648), .B(n34649), .Z(n34647) );
  ANDN U34871 ( .B(B[175]), .A(n82), .Z(n34428) );
  XOR U34872 ( .A(n34435), .B(n34650), .Z(n34429) );
  XNOR U34873 ( .A(n34433), .B(n34436), .Z(n34650) );
  NAND U34874 ( .A(A[2]), .B(B[176]), .Z(n34436) );
  NANDN U34875 ( .A(n34651), .B(n34652), .Z(n34433) );
  AND U34876 ( .A(A[0]), .B(B[177]), .Z(n34652) );
  XNOR U34877 ( .A(n34438), .B(n34653), .Z(n34435) );
  NAND U34878 ( .A(A[0]), .B(B[178]), .Z(n34653) );
  NAND U34879 ( .A(B[177]), .B(A[1]), .Z(n34438) );
  NAND U34880 ( .A(n34654), .B(n34655), .Z(n440) );
  NANDN U34881 ( .A(n34656), .B(n34657), .Z(n34655) );
  OR U34882 ( .A(n34658), .B(n34659), .Z(n34657) );
  NAND U34883 ( .A(n34659), .B(n34658), .Z(n34654) );
  XOR U34884 ( .A(n442), .B(n441), .Z(\A1[175] ) );
  XOR U34885 ( .A(n34659), .B(n34660), .Z(n441) );
  XNOR U34886 ( .A(n34658), .B(n34656), .Z(n34660) );
  AND U34887 ( .A(n34661), .B(n34662), .Z(n34656) );
  NANDN U34888 ( .A(n34663), .B(n34664), .Z(n34662) );
  NANDN U34889 ( .A(n34665), .B(n34666), .Z(n34664) );
  NANDN U34890 ( .A(n34666), .B(n34665), .Z(n34661) );
  ANDN U34891 ( .B(B[146]), .A(n54), .Z(n34658) );
  XNOR U34892 ( .A(n34453), .B(n34667), .Z(n34659) );
  XNOR U34893 ( .A(n34452), .B(n34450), .Z(n34667) );
  AND U34894 ( .A(n34668), .B(n34669), .Z(n34450) );
  NANDN U34895 ( .A(n34670), .B(n34671), .Z(n34669) );
  OR U34896 ( .A(n34672), .B(n34673), .Z(n34671) );
  NAND U34897 ( .A(n34673), .B(n34672), .Z(n34668) );
  ANDN U34898 ( .B(B[147]), .A(n55), .Z(n34452) );
  XNOR U34899 ( .A(n34460), .B(n34674), .Z(n34453) );
  XNOR U34900 ( .A(n34459), .B(n34457), .Z(n34674) );
  AND U34901 ( .A(n34675), .B(n34676), .Z(n34457) );
  NANDN U34902 ( .A(n34677), .B(n34678), .Z(n34676) );
  NANDN U34903 ( .A(n34679), .B(n34680), .Z(n34678) );
  NANDN U34904 ( .A(n34680), .B(n34679), .Z(n34675) );
  ANDN U34905 ( .B(B[148]), .A(n56), .Z(n34459) );
  XNOR U34906 ( .A(n34467), .B(n34681), .Z(n34460) );
  XNOR U34907 ( .A(n34466), .B(n34464), .Z(n34681) );
  AND U34908 ( .A(n34682), .B(n34683), .Z(n34464) );
  NANDN U34909 ( .A(n34684), .B(n34685), .Z(n34683) );
  OR U34910 ( .A(n34686), .B(n34687), .Z(n34685) );
  NAND U34911 ( .A(n34687), .B(n34686), .Z(n34682) );
  ANDN U34912 ( .B(B[149]), .A(n57), .Z(n34466) );
  XNOR U34913 ( .A(n34474), .B(n34688), .Z(n34467) );
  XNOR U34914 ( .A(n34473), .B(n34471), .Z(n34688) );
  AND U34915 ( .A(n34689), .B(n34690), .Z(n34471) );
  NANDN U34916 ( .A(n34691), .B(n34692), .Z(n34690) );
  NANDN U34917 ( .A(n34693), .B(n34694), .Z(n34692) );
  NANDN U34918 ( .A(n34694), .B(n34693), .Z(n34689) );
  ANDN U34919 ( .B(B[150]), .A(n58), .Z(n34473) );
  XNOR U34920 ( .A(n34481), .B(n34695), .Z(n34474) );
  XNOR U34921 ( .A(n34480), .B(n34478), .Z(n34695) );
  AND U34922 ( .A(n34696), .B(n34697), .Z(n34478) );
  NANDN U34923 ( .A(n34698), .B(n34699), .Z(n34697) );
  OR U34924 ( .A(n34700), .B(n34701), .Z(n34699) );
  NAND U34925 ( .A(n34701), .B(n34700), .Z(n34696) );
  ANDN U34926 ( .B(B[151]), .A(n59), .Z(n34480) );
  XNOR U34927 ( .A(n34488), .B(n34702), .Z(n34481) );
  XNOR U34928 ( .A(n34487), .B(n34485), .Z(n34702) );
  AND U34929 ( .A(n34703), .B(n34704), .Z(n34485) );
  NANDN U34930 ( .A(n34705), .B(n34706), .Z(n34704) );
  NANDN U34931 ( .A(n34707), .B(n34708), .Z(n34706) );
  NANDN U34932 ( .A(n34708), .B(n34707), .Z(n34703) );
  ANDN U34933 ( .B(B[152]), .A(n60), .Z(n34487) );
  XNOR U34934 ( .A(n34495), .B(n34709), .Z(n34488) );
  XNOR U34935 ( .A(n34494), .B(n34492), .Z(n34709) );
  AND U34936 ( .A(n34710), .B(n34711), .Z(n34492) );
  NANDN U34937 ( .A(n34712), .B(n34713), .Z(n34711) );
  OR U34938 ( .A(n34714), .B(n34715), .Z(n34713) );
  NAND U34939 ( .A(n34715), .B(n34714), .Z(n34710) );
  ANDN U34940 ( .B(B[153]), .A(n61), .Z(n34494) );
  XNOR U34941 ( .A(n34502), .B(n34716), .Z(n34495) );
  XNOR U34942 ( .A(n34501), .B(n34499), .Z(n34716) );
  AND U34943 ( .A(n34717), .B(n34718), .Z(n34499) );
  NANDN U34944 ( .A(n34719), .B(n34720), .Z(n34718) );
  NANDN U34945 ( .A(n34721), .B(n34722), .Z(n34720) );
  NANDN U34946 ( .A(n34722), .B(n34721), .Z(n34717) );
  ANDN U34947 ( .B(B[154]), .A(n62), .Z(n34501) );
  XNOR U34948 ( .A(n34509), .B(n34723), .Z(n34502) );
  XNOR U34949 ( .A(n34508), .B(n34506), .Z(n34723) );
  AND U34950 ( .A(n34724), .B(n34725), .Z(n34506) );
  NANDN U34951 ( .A(n34726), .B(n34727), .Z(n34725) );
  OR U34952 ( .A(n34728), .B(n34729), .Z(n34727) );
  NAND U34953 ( .A(n34729), .B(n34728), .Z(n34724) );
  ANDN U34954 ( .B(B[155]), .A(n63), .Z(n34508) );
  XNOR U34955 ( .A(n34516), .B(n34730), .Z(n34509) );
  XNOR U34956 ( .A(n34515), .B(n34513), .Z(n34730) );
  AND U34957 ( .A(n34731), .B(n34732), .Z(n34513) );
  NANDN U34958 ( .A(n34733), .B(n34734), .Z(n34732) );
  NANDN U34959 ( .A(n34735), .B(n34736), .Z(n34734) );
  NANDN U34960 ( .A(n34736), .B(n34735), .Z(n34731) );
  ANDN U34961 ( .B(B[156]), .A(n64), .Z(n34515) );
  XNOR U34962 ( .A(n34523), .B(n34737), .Z(n34516) );
  XNOR U34963 ( .A(n34522), .B(n34520), .Z(n34737) );
  AND U34964 ( .A(n34738), .B(n34739), .Z(n34520) );
  NANDN U34965 ( .A(n34740), .B(n34741), .Z(n34739) );
  OR U34966 ( .A(n34742), .B(n34743), .Z(n34741) );
  NAND U34967 ( .A(n34743), .B(n34742), .Z(n34738) );
  ANDN U34968 ( .B(B[157]), .A(n65), .Z(n34522) );
  XNOR U34969 ( .A(n34530), .B(n34744), .Z(n34523) );
  XNOR U34970 ( .A(n34529), .B(n34527), .Z(n34744) );
  AND U34971 ( .A(n34745), .B(n34746), .Z(n34527) );
  NANDN U34972 ( .A(n34747), .B(n34748), .Z(n34746) );
  NANDN U34973 ( .A(n34749), .B(n34750), .Z(n34748) );
  NANDN U34974 ( .A(n34750), .B(n34749), .Z(n34745) );
  ANDN U34975 ( .B(B[158]), .A(n66), .Z(n34529) );
  XNOR U34976 ( .A(n34537), .B(n34751), .Z(n34530) );
  XNOR U34977 ( .A(n34536), .B(n34534), .Z(n34751) );
  AND U34978 ( .A(n34752), .B(n34753), .Z(n34534) );
  NANDN U34979 ( .A(n34754), .B(n34755), .Z(n34753) );
  OR U34980 ( .A(n34756), .B(n34757), .Z(n34755) );
  NAND U34981 ( .A(n34757), .B(n34756), .Z(n34752) );
  ANDN U34982 ( .B(B[159]), .A(n67), .Z(n34536) );
  XNOR U34983 ( .A(n34544), .B(n34758), .Z(n34537) );
  XNOR U34984 ( .A(n34543), .B(n34541), .Z(n34758) );
  AND U34985 ( .A(n34759), .B(n34760), .Z(n34541) );
  NANDN U34986 ( .A(n34761), .B(n34762), .Z(n34760) );
  NANDN U34987 ( .A(n34763), .B(n34764), .Z(n34762) );
  NANDN U34988 ( .A(n34764), .B(n34763), .Z(n34759) );
  ANDN U34989 ( .B(B[160]), .A(n68), .Z(n34543) );
  XNOR U34990 ( .A(n34551), .B(n34765), .Z(n34544) );
  XNOR U34991 ( .A(n34550), .B(n34548), .Z(n34765) );
  AND U34992 ( .A(n34766), .B(n34767), .Z(n34548) );
  NANDN U34993 ( .A(n34768), .B(n34769), .Z(n34767) );
  OR U34994 ( .A(n34770), .B(n34771), .Z(n34769) );
  NAND U34995 ( .A(n34771), .B(n34770), .Z(n34766) );
  ANDN U34996 ( .B(B[161]), .A(n69), .Z(n34550) );
  XNOR U34997 ( .A(n34558), .B(n34772), .Z(n34551) );
  XNOR U34998 ( .A(n34557), .B(n34555), .Z(n34772) );
  AND U34999 ( .A(n34773), .B(n34774), .Z(n34555) );
  NANDN U35000 ( .A(n34775), .B(n34776), .Z(n34774) );
  NANDN U35001 ( .A(n34777), .B(n34778), .Z(n34776) );
  NANDN U35002 ( .A(n34778), .B(n34777), .Z(n34773) );
  ANDN U35003 ( .B(B[162]), .A(n70), .Z(n34557) );
  XNOR U35004 ( .A(n34565), .B(n34779), .Z(n34558) );
  XNOR U35005 ( .A(n34564), .B(n34562), .Z(n34779) );
  AND U35006 ( .A(n34780), .B(n34781), .Z(n34562) );
  NANDN U35007 ( .A(n34782), .B(n34783), .Z(n34781) );
  OR U35008 ( .A(n34784), .B(n34785), .Z(n34783) );
  NAND U35009 ( .A(n34785), .B(n34784), .Z(n34780) );
  ANDN U35010 ( .B(B[163]), .A(n71), .Z(n34564) );
  XNOR U35011 ( .A(n34572), .B(n34786), .Z(n34565) );
  XNOR U35012 ( .A(n34571), .B(n34569), .Z(n34786) );
  AND U35013 ( .A(n34787), .B(n34788), .Z(n34569) );
  NANDN U35014 ( .A(n34789), .B(n34790), .Z(n34788) );
  NANDN U35015 ( .A(n34791), .B(n34792), .Z(n34790) );
  NANDN U35016 ( .A(n34792), .B(n34791), .Z(n34787) );
  ANDN U35017 ( .B(B[164]), .A(n72), .Z(n34571) );
  XNOR U35018 ( .A(n34579), .B(n34793), .Z(n34572) );
  XNOR U35019 ( .A(n34578), .B(n34576), .Z(n34793) );
  AND U35020 ( .A(n34794), .B(n34795), .Z(n34576) );
  NANDN U35021 ( .A(n34796), .B(n34797), .Z(n34795) );
  OR U35022 ( .A(n34798), .B(n34799), .Z(n34797) );
  NAND U35023 ( .A(n34799), .B(n34798), .Z(n34794) );
  ANDN U35024 ( .B(B[165]), .A(n73), .Z(n34578) );
  XNOR U35025 ( .A(n34586), .B(n34800), .Z(n34579) );
  XNOR U35026 ( .A(n34585), .B(n34583), .Z(n34800) );
  AND U35027 ( .A(n34801), .B(n34802), .Z(n34583) );
  NANDN U35028 ( .A(n34803), .B(n34804), .Z(n34802) );
  NANDN U35029 ( .A(n34805), .B(n34806), .Z(n34804) );
  NANDN U35030 ( .A(n34806), .B(n34805), .Z(n34801) );
  ANDN U35031 ( .B(B[166]), .A(n74), .Z(n34585) );
  XNOR U35032 ( .A(n34593), .B(n34807), .Z(n34586) );
  XNOR U35033 ( .A(n34592), .B(n34590), .Z(n34807) );
  AND U35034 ( .A(n34808), .B(n34809), .Z(n34590) );
  NANDN U35035 ( .A(n34810), .B(n34811), .Z(n34809) );
  OR U35036 ( .A(n34812), .B(n34813), .Z(n34811) );
  NAND U35037 ( .A(n34813), .B(n34812), .Z(n34808) );
  ANDN U35038 ( .B(B[167]), .A(n75), .Z(n34592) );
  XNOR U35039 ( .A(n34600), .B(n34814), .Z(n34593) );
  XNOR U35040 ( .A(n34599), .B(n34597), .Z(n34814) );
  AND U35041 ( .A(n34815), .B(n34816), .Z(n34597) );
  NANDN U35042 ( .A(n34817), .B(n34818), .Z(n34816) );
  NANDN U35043 ( .A(n34819), .B(n34820), .Z(n34818) );
  NANDN U35044 ( .A(n34820), .B(n34819), .Z(n34815) );
  ANDN U35045 ( .B(B[168]), .A(n76), .Z(n34599) );
  XNOR U35046 ( .A(n34607), .B(n34821), .Z(n34600) );
  XNOR U35047 ( .A(n34606), .B(n34604), .Z(n34821) );
  AND U35048 ( .A(n34822), .B(n34823), .Z(n34604) );
  NANDN U35049 ( .A(n34824), .B(n34825), .Z(n34823) );
  OR U35050 ( .A(n34826), .B(n34827), .Z(n34825) );
  NAND U35051 ( .A(n34827), .B(n34826), .Z(n34822) );
  ANDN U35052 ( .B(B[169]), .A(n77), .Z(n34606) );
  XNOR U35053 ( .A(n34614), .B(n34828), .Z(n34607) );
  XNOR U35054 ( .A(n34613), .B(n34611), .Z(n34828) );
  AND U35055 ( .A(n34829), .B(n34830), .Z(n34611) );
  NANDN U35056 ( .A(n34831), .B(n34832), .Z(n34830) );
  NANDN U35057 ( .A(n34833), .B(n34834), .Z(n34832) );
  NANDN U35058 ( .A(n34834), .B(n34833), .Z(n34829) );
  ANDN U35059 ( .B(B[170]), .A(n78), .Z(n34613) );
  XNOR U35060 ( .A(n34621), .B(n34835), .Z(n34614) );
  XNOR U35061 ( .A(n34620), .B(n34618), .Z(n34835) );
  AND U35062 ( .A(n34836), .B(n34837), .Z(n34618) );
  NANDN U35063 ( .A(n34838), .B(n34839), .Z(n34837) );
  OR U35064 ( .A(n34840), .B(n34841), .Z(n34839) );
  NAND U35065 ( .A(n34841), .B(n34840), .Z(n34836) );
  ANDN U35066 ( .B(B[171]), .A(n79), .Z(n34620) );
  XNOR U35067 ( .A(n34628), .B(n34842), .Z(n34621) );
  XNOR U35068 ( .A(n34627), .B(n34625), .Z(n34842) );
  AND U35069 ( .A(n34843), .B(n34844), .Z(n34625) );
  NANDN U35070 ( .A(n34845), .B(n34846), .Z(n34844) );
  NANDN U35071 ( .A(n34847), .B(n34848), .Z(n34846) );
  NANDN U35072 ( .A(n34848), .B(n34847), .Z(n34843) );
  ANDN U35073 ( .B(B[172]), .A(n80), .Z(n34627) );
  XNOR U35074 ( .A(n34635), .B(n34849), .Z(n34628) );
  XNOR U35075 ( .A(n34634), .B(n34632), .Z(n34849) );
  AND U35076 ( .A(n34850), .B(n34851), .Z(n34632) );
  NANDN U35077 ( .A(n34852), .B(n34853), .Z(n34851) );
  OR U35078 ( .A(n34854), .B(n34855), .Z(n34853) );
  NAND U35079 ( .A(n34855), .B(n34854), .Z(n34850) );
  ANDN U35080 ( .B(B[173]), .A(n81), .Z(n34634) );
  XNOR U35081 ( .A(n34642), .B(n34856), .Z(n34635) );
  XNOR U35082 ( .A(n34641), .B(n34639), .Z(n34856) );
  AND U35083 ( .A(n34857), .B(n34858), .Z(n34639) );
  NANDN U35084 ( .A(n34859), .B(n34860), .Z(n34858) );
  NAND U35085 ( .A(n34861), .B(n34862), .Z(n34860) );
  ANDN U35086 ( .B(B[174]), .A(n82), .Z(n34641) );
  XOR U35087 ( .A(n34648), .B(n34863), .Z(n34642) );
  XNOR U35088 ( .A(n34646), .B(n34649), .Z(n34863) );
  NAND U35089 ( .A(A[2]), .B(B[175]), .Z(n34649) );
  NANDN U35090 ( .A(n34864), .B(n34865), .Z(n34646) );
  AND U35091 ( .A(A[0]), .B(B[176]), .Z(n34865) );
  XNOR U35092 ( .A(n34651), .B(n34866), .Z(n34648) );
  NAND U35093 ( .A(A[0]), .B(B[177]), .Z(n34866) );
  NAND U35094 ( .A(B[176]), .B(A[1]), .Z(n34651) );
  NAND U35095 ( .A(n34867), .B(n34868), .Z(n442) );
  NANDN U35096 ( .A(n34869), .B(n34870), .Z(n34868) );
  OR U35097 ( .A(n34871), .B(n34872), .Z(n34870) );
  NAND U35098 ( .A(n34872), .B(n34871), .Z(n34867) );
  XOR U35099 ( .A(n444), .B(n443), .Z(\A1[174] ) );
  XOR U35100 ( .A(n34872), .B(n34873), .Z(n443) );
  XNOR U35101 ( .A(n34871), .B(n34869), .Z(n34873) );
  AND U35102 ( .A(n34874), .B(n34875), .Z(n34869) );
  NANDN U35103 ( .A(n34876), .B(n34877), .Z(n34875) );
  NANDN U35104 ( .A(n34878), .B(n34879), .Z(n34877) );
  NANDN U35105 ( .A(n34879), .B(n34878), .Z(n34874) );
  ANDN U35106 ( .B(B[145]), .A(n54), .Z(n34871) );
  XNOR U35107 ( .A(n34666), .B(n34880), .Z(n34872) );
  XNOR U35108 ( .A(n34665), .B(n34663), .Z(n34880) );
  AND U35109 ( .A(n34881), .B(n34882), .Z(n34663) );
  NANDN U35110 ( .A(n34883), .B(n34884), .Z(n34882) );
  OR U35111 ( .A(n34885), .B(n34886), .Z(n34884) );
  NAND U35112 ( .A(n34886), .B(n34885), .Z(n34881) );
  ANDN U35113 ( .B(B[146]), .A(n55), .Z(n34665) );
  XNOR U35114 ( .A(n34673), .B(n34887), .Z(n34666) );
  XNOR U35115 ( .A(n34672), .B(n34670), .Z(n34887) );
  AND U35116 ( .A(n34888), .B(n34889), .Z(n34670) );
  NANDN U35117 ( .A(n34890), .B(n34891), .Z(n34889) );
  NANDN U35118 ( .A(n34892), .B(n34893), .Z(n34891) );
  NANDN U35119 ( .A(n34893), .B(n34892), .Z(n34888) );
  ANDN U35120 ( .B(B[147]), .A(n56), .Z(n34672) );
  XNOR U35121 ( .A(n34680), .B(n34894), .Z(n34673) );
  XNOR U35122 ( .A(n34679), .B(n34677), .Z(n34894) );
  AND U35123 ( .A(n34895), .B(n34896), .Z(n34677) );
  NANDN U35124 ( .A(n34897), .B(n34898), .Z(n34896) );
  OR U35125 ( .A(n34899), .B(n34900), .Z(n34898) );
  NAND U35126 ( .A(n34900), .B(n34899), .Z(n34895) );
  ANDN U35127 ( .B(B[148]), .A(n57), .Z(n34679) );
  XNOR U35128 ( .A(n34687), .B(n34901), .Z(n34680) );
  XNOR U35129 ( .A(n34686), .B(n34684), .Z(n34901) );
  AND U35130 ( .A(n34902), .B(n34903), .Z(n34684) );
  NANDN U35131 ( .A(n34904), .B(n34905), .Z(n34903) );
  NANDN U35132 ( .A(n34906), .B(n34907), .Z(n34905) );
  NANDN U35133 ( .A(n34907), .B(n34906), .Z(n34902) );
  ANDN U35134 ( .B(B[149]), .A(n58), .Z(n34686) );
  XNOR U35135 ( .A(n34694), .B(n34908), .Z(n34687) );
  XNOR U35136 ( .A(n34693), .B(n34691), .Z(n34908) );
  AND U35137 ( .A(n34909), .B(n34910), .Z(n34691) );
  NANDN U35138 ( .A(n34911), .B(n34912), .Z(n34910) );
  OR U35139 ( .A(n34913), .B(n34914), .Z(n34912) );
  NAND U35140 ( .A(n34914), .B(n34913), .Z(n34909) );
  ANDN U35141 ( .B(B[150]), .A(n59), .Z(n34693) );
  XNOR U35142 ( .A(n34701), .B(n34915), .Z(n34694) );
  XNOR U35143 ( .A(n34700), .B(n34698), .Z(n34915) );
  AND U35144 ( .A(n34916), .B(n34917), .Z(n34698) );
  NANDN U35145 ( .A(n34918), .B(n34919), .Z(n34917) );
  NANDN U35146 ( .A(n34920), .B(n34921), .Z(n34919) );
  NANDN U35147 ( .A(n34921), .B(n34920), .Z(n34916) );
  ANDN U35148 ( .B(B[151]), .A(n60), .Z(n34700) );
  XNOR U35149 ( .A(n34708), .B(n34922), .Z(n34701) );
  XNOR U35150 ( .A(n34707), .B(n34705), .Z(n34922) );
  AND U35151 ( .A(n34923), .B(n34924), .Z(n34705) );
  NANDN U35152 ( .A(n34925), .B(n34926), .Z(n34924) );
  OR U35153 ( .A(n34927), .B(n34928), .Z(n34926) );
  NAND U35154 ( .A(n34928), .B(n34927), .Z(n34923) );
  ANDN U35155 ( .B(B[152]), .A(n61), .Z(n34707) );
  XNOR U35156 ( .A(n34715), .B(n34929), .Z(n34708) );
  XNOR U35157 ( .A(n34714), .B(n34712), .Z(n34929) );
  AND U35158 ( .A(n34930), .B(n34931), .Z(n34712) );
  NANDN U35159 ( .A(n34932), .B(n34933), .Z(n34931) );
  NANDN U35160 ( .A(n34934), .B(n34935), .Z(n34933) );
  NANDN U35161 ( .A(n34935), .B(n34934), .Z(n34930) );
  ANDN U35162 ( .B(B[153]), .A(n62), .Z(n34714) );
  XNOR U35163 ( .A(n34722), .B(n34936), .Z(n34715) );
  XNOR U35164 ( .A(n34721), .B(n34719), .Z(n34936) );
  AND U35165 ( .A(n34937), .B(n34938), .Z(n34719) );
  NANDN U35166 ( .A(n34939), .B(n34940), .Z(n34938) );
  OR U35167 ( .A(n34941), .B(n34942), .Z(n34940) );
  NAND U35168 ( .A(n34942), .B(n34941), .Z(n34937) );
  ANDN U35169 ( .B(B[154]), .A(n63), .Z(n34721) );
  XNOR U35170 ( .A(n34729), .B(n34943), .Z(n34722) );
  XNOR U35171 ( .A(n34728), .B(n34726), .Z(n34943) );
  AND U35172 ( .A(n34944), .B(n34945), .Z(n34726) );
  NANDN U35173 ( .A(n34946), .B(n34947), .Z(n34945) );
  NANDN U35174 ( .A(n34948), .B(n34949), .Z(n34947) );
  NANDN U35175 ( .A(n34949), .B(n34948), .Z(n34944) );
  ANDN U35176 ( .B(B[155]), .A(n64), .Z(n34728) );
  XNOR U35177 ( .A(n34736), .B(n34950), .Z(n34729) );
  XNOR U35178 ( .A(n34735), .B(n34733), .Z(n34950) );
  AND U35179 ( .A(n34951), .B(n34952), .Z(n34733) );
  NANDN U35180 ( .A(n34953), .B(n34954), .Z(n34952) );
  OR U35181 ( .A(n34955), .B(n34956), .Z(n34954) );
  NAND U35182 ( .A(n34956), .B(n34955), .Z(n34951) );
  ANDN U35183 ( .B(B[156]), .A(n65), .Z(n34735) );
  XNOR U35184 ( .A(n34743), .B(n34957), .Z(n34736) );
  XNOR U35185 ( .A(n34742), .B(n34740), .Z(n34957) );
  AND U35186 ( .A(n34958), .B(n34959), .Z(n34740) );
  NANDN U35187 ( .A(n34960), .B(n34961), .Z(n34959) );
  NANDN U35188 ( .A(n34962), .B(n34963), .Z(n34961) );
  NANDN U35189 ( .A(n34963), .B(n34962), .Z(n34958) );
  ANDN U35190 ( .B(B[157]), .A(n66), .Z(n34742) );
  XNOR U35191 ( .A(n34750), .B(n34964), .Z(n34743) );
  XNOR U35192 ( .A(n34749), .B(n34747), .Z(n34964) );
  AND U35193 ( .A(n34965), .B(n34966), .Z(n34747) );
  NANDN U35194 ( .A(n34967), .B(n34968), .Z(n34966) );
  OR U35195 ( .A(n34969), .B(n34970), .Z(n34968) );
  NAND U35196 ( .A(n34970), .B(n34969), .Z(n34965) );
  ANDN U35197 ( .B(B[158]), .A(n67), .Z(n34749) );
  XNOR U35198 ( .A(n34757), .B(n34971), .Z(n34750) );
  XNOR U35199 ( .A(n34756), .B(n34754), .Z(n34971) );
  AND U35200 ( .A(n34972), .B(n34973), .Z(n34754) );
  NANDN U35201 ( .A(n34974), .B(n34975), .Z(n34973) );
  NANDN U35202 ( .A(n34976), .B(n34977), .Z(n34975) );
  NANDN U35203 ( .A(n34977), .B(n34976), .Z(n34972) );
  ANDN U35204 ( .B(B[159]), .A(n68), .Z(n34756) );
  XNOR U35205 ( .A(n34764), .B(n34978), .Z(n34757) );
  XNOR U35206 ( .A(n34763), .B(n34761), .Z(n34978) );
  AND U35207 ( .A(n34979), .B(n34980), .Z(n34761) );
  NANDN U35208 ( .A(n34981), .B(n34982), .Z(n34980) );
  OR U35209 ( .A(n34983), .B(n34984), .Z(n34982) );
  NAND U35210 ( .A(n34984), .B(n34983), .Z(n34979) );
  ANDN U35211 ( .B(B[160]), .A(n69), .Z(n34763) );
  XNOR U35212 ( .A(n34771), .B(n34985), .Z(n34764) );
  XNOR U35213 ( .A(n34770), .B(n34768), .Z(n34985) );
  AND U35214 ( .A(n34986), .B(n34987), .Z(n34768) );
  NANDN U35215 ( .A(n34988), .B(n34989), .Z(n34987) );
  NANDN U35216 ( .A(n34990), .B(n34991), .Z(n34989) );
  NANDN U35217 ( .A(n34991), .B(n34990), .Z(n34986) );
  ANDN U35218 ( .B(B[161]), .A(n70), .Z(n34770) );
  XNOR U35219 ( .A(n34778), .B(n34992), .Z(n34771) );
  XNOR U35220 ( .A(n34777), .B(n34775), .Z(n34992) );
  AND U35221 ( .A(n34993), .B(n34994), .Z(n34775) );
  NANDN U35222 ( .A(n34995), .B(n34996), .Z(n34994) );
  OR U35223 ( .A(n34997), .B(n34998), .Z(n34996) );
  NAND U35224 ( .A(n34998), .B(n34997), .Z(n34993) );
  ANDN U35225 ( .B(B[162]), .A(n71), .Z(n34777) );
  XNOR U35226 ( .A(n34785), .B(n34999), .Z(n34778) );
  XNOR U35227 ( .A(n34784), .B(n34782), .Z(n34999) );
  AND U35228 ( .A(n35000), .B(n35001), .Z(n34782) );
  NANDN U35229 ( .A(n35002), .B(n35003), .Z(n35001) );
  NANDN U35230 ( .A(n35004), .B(n35005), .Z(n35003) );
  NANDN U35231 ( .A(n35005), .B(n35004), .Z(n35000) );
  ANDN U35232 ( .B(B[163]), .A(n72), .Z(n34784) );
  XNOR U35233 ( .A(n34792), .B(n35006), .Z(n34785) );
  XNOR U35234 ( .A(n34791), .B(n34789), .Z(n35006) );
  AND U35235 ( .A(n35007), .B(n35008), .Z(n34789) );
  NANDN U35236 ( .A(n35009), .B(n35010), .Z(n35008) );
  OR U35237 ( .A(n35011), .B(n35012), .Z(n35010) );
  NAND U35238 ( .A(n35012), .B(n35011), .Z(n35007) );
  ANDN U35239 ( .B(B[164]), .A(n73), .Z(n34791) );
  XNOR U35240 ( .A(n34799), .B(n35013), .Z(n34792) );
  XNOR U35241 ( .A(n34798), .B(n34796), .Z(n35013) );
  AND U35242 ( .A(n35014), .B(n35015), .Z(n34796) );
  NANDN U35243 ( .A(n35016), .B(n35017), .Z(n35015) );
  NANDN U35244 ( .A(n35018), .B(n35019), .Z(n35017) );
  NANDN U35245 ( .A(n35019), .B(n35018), .Z(n35014) );
  ANDN U35246 ( .B(B[165]), .A(n74), .Z(n34798) );
  XNOR U35247 ( .A(n34806), .B(n35020), .Z(n34799) );
  XNOR U35248 ( .A(n34805), .B(n34803), .Z(n35020) );
  AND U35249 ( .A(n35021), .B(n35022), .Z(n34803) );
  NANDN U35250 ( .A(n35023), .B(n35024), .Z(n35022) );
  OR U35251 ( .A(n35025), .B(n35026), .Z(n35024) );
  NAND U35252 ( .A(n35026), .B(n35025), .Z(n35021) );
  ANDN U35253 ( .B(B[166]), .A(n75), .Z(n34805) );
  XNOR U35254 ( .A(n34813), .B(n35027), .Z(n34806) );
  XNOR U35255 ( .A(n34812), .B(n34810), .Z(n35027) );
  AND U35256 ( .A(n35028), .B(n35029), .Z(n34810) );
  NANDN U35257 ( .A(n35030), .B(n35031), .Z(n35029) );
  NANDN U35258 ( .A(n35032), .B(n35033), .Z(n35031) );
  NANDN U35259 ( .A(n35033), .B(n35032), .Z(n35028) );
  ANDN U35260 ( .B(B[167]), .A(n76), .Z(n34812) );
  XNOR U35261 ( .A(n34820), .B(n35034), .Z(n34813) );
  XNOR U35262 ( .A(n34819), .B(n34817), .Z(n35034) );
  AND U35263 ( .A(n35035), .B(n35036), .Z(n34817) );
  NANDN U35264 ( .A(n35037), .B(n35038), .Z(n35036) );
  OR U35265 ( .A(n35039), .B(n35040), .Z(n35038) );
  NAND U35266 ( .A(n35040), .B(n35039), .Z(n35035) );
  ANDN U35267 ( .B(B[168]), .A(n77), .Z(n34819) );
  XNOR U35268 ( .A(n34827), .B(n35041), .Z(n34820) );
  XNOR U35269 ( .A(n34826), .B(n34824), .Z(n35041) );
  AND U35270 ( .A(n35042), .B(n35043), .Z(n34824) );
  NANDN U35271 ( .A(n35044), .B(n35045), .Z(n35043) );
  NANDN U35272 ( .A(n35046), .B(n35047), .Z(n35045) );
  NANDN U35273 ( .A(n35047), .B(n35046), .Z(n35042) );
  ANDN U35274 ( .B(B[169]), .A(n78), .Z(n34826) );
  XNOR U35275 ( .A(n34834), .B(n35048), .Z(n34827) );
  XNOR U35276 ( .A(n34833), .B(n34831), .Z(n35048) );
  AND U35277 ( .A(n35049), .B(n35050), .Z(n34831) );
  NANDN U35278 ( .A(n35051), .B(n35052), .Z(n35050) );
  OR U35279 ( .A(n35053), .B(n35054), .Z(n35052) );
  NAND U35280 ( .A(n35054), .B(n35053), .Z(n35049) );
  ANDN U35281 ( .B(B[170]), .A(n79), .Z(n34833) );
  XNOR U35282 ( .A(n34841), .B(n35055), .Z(n34834) );
  XNOR U35283 ( .A(n34840), .B(n34838), .Z(n35055) );
  AND U35284 ( .A(n35056), .B(n35057), .Z(n34838) );
  NANDN U35285 ( .A(n35058), .B(n35059), .Z(n35057) );
  NANDN U35286 ( .A(n35060), .B(n35061), .Z(n35059) );
  NANDN U35287 ( .A(n35061), .B(n35060), .Z(n35056) );
  ANDN U35288 ( .B(B[171]), .A(n80), .Z(n34840) );
  XNOR U35289 ( .A(n34848), .B(n35062), .Z(n34841) );
  XNOR U35290 ( .A(n34847), .B(n34845), .Z(n35062) );
  AND U35291 ( .A(n35063), .B(n35064), .Z(n34845) );
  NANDN U35292 ( .A(n35065), .B(n35066), .Z(n35064) );
  OR U35293 ( .A(n35067), .B(n35068), .Z(n35066) );
  NAND U35294 ( .A(n35068), .B(n35067), .Z(n35063) );
  ANDN U35295 ( .B(B[172]), .A(n81), .Z(n34847) );
  XNOR U35296 ( .A(n34855), .B(n35069), .Z(n34848) );
  XNOR U35297 ( .A(n34854), .B(n34852), .Z(n35069) );
  AND U35298 ( .A(n35070), .B(n35071), .Z(n34852) );
  NANDN U35299 ( .A(n35072), .B(n35073), .Z(n35071) );
  NAND U35300 ( .A(n35074), .B(n35075), .Z(n35073) );
  ANDN U35301 ( .B(B[173]), .A(n82), .Z(n34854) );
  XOR U35302 ( .A(n34861), .B(n35076), .Z(n34855) );
  XNOR U35303 ( .A(n34859), .B(n34862), .Z(n35076) );
  NAND U35304 ( .A(A[2]), .B(B[174]), .Z(n34862) );
  NANDN U35305 ( .A(n35077), .B(n35078), .Z(n34859) );
  AND U35306 ( .A(A[0]), .B(B[175]), .Z(n35078) );
  XNOR U35307 ( .A(n34864), .B(n35079), .Z(n34861) );
  NAND U35308 ( .A(A[0]), .B(B[176]), .Z(n35079) );
  NAND U35309 ( .A(B[175]), .B(A[1]), .Z(n34864) );
  NAND U35310 ( .A(n35080), .B(n35081), .Z(n444) );
  NANDN U35311 ( .A(n35082), .B(n35083), .Z(n35081) );
  OR U35312 ( .A(n35084), .B(n35085), .Z(n35083) );
  NAND U35313 ( .A(n35085), .B(n35084), .Z(n35080) );
  XOR U35314 ( .A(n446), .B(n445), .Z(\A1[173] ) );
  XOR U35315 ( .A(n35085), .B(n35086), .Z(n445) );
  XNOR U35316 ( .A(n35084), .B(n35082), .Z(n35086) );
  AND U35317 ( .A(n35087), .B(n35088), .Z(n35082) );
  NANDN U35318 ( .A(n35089), .B(n35090), .Z(n35088) );
  NANDN U35319 ( .A(n35091), .B(n35092), .Z(n35090) );
  NANDN U35320 ( .A(n35092), .B(n35091), .Z(n35087) );
  ANDN U35321 ( .B(B[144]), .A(n54), .Z(n35084) );
  XNOR U35322 ( .A(n34879), .B(n35093), .Z(n35085) );
  XNOR U35323 ( .A(n34878), .B(n34876), .Z(n35093) );
  AND U35324 ( .A(n35094), .B(n35095), .Z(n34876) );
  NANDN U35325 ( .A(n35096), .B(n35097), .Z(n35095) );
  OR U35326 ( .A(n35098), .B(n35099), .Z(n35097) );
  NAND U35327 ( .A(n35099), .B(n35098), .Z(n35094) );
  ANDN U35328 ( .B(B[145]), .A(n55), .Z(n34878) );
  XNOR U35329 ( .A(n34886), .B(n35100), .Z(n34879) );
  XNOR U35330 ( .A(n34885), .B(n34883), .Z(n35100) );
  AND U35331 ( .A(n35101), .B(n35102), .Z(n34883) );
  NANDN U35332 ( .A(n35103), .B(n35104), .Z(n35102) );
  NANDN U35333 ( .A(n35105), .B(n35106), .Z(n35104) );
  NANDN U35334 ( .A(n35106), .B(n35105), .Z(n35101) );
  ANDN U35335 ( .B(B[146]), .A(n56), .Z(n34885) );
  XNOR U35336 ( .A(n34893), .B(n35107), .Z(n34886) );
  XNOR U35337 ( .A(n34892), .B(n34890), .Z(n35107) );
  AND U35338 ( .A(n35108), .B(n35109), .Z(n34890) );
  NANDN U35339 ( .A(n35110), .B(n35111), .Z(n35109) );
  OR U35340 ( .A(n35112), .B(n35113), .Z(n35111) );
  NAND U35341 ( .A(n35113), .B(n35112), .Z(n35108) );
  ANDN U35342 ( .B(B[147]), .A(n57), .Z(n34892) );
  XNOR U35343 ( .A(n34900), .B(n35114), .Z(n34893) );
  XNOR U35344 ( .A(n34899), .B(n34897), .Z(n35114) );
  AND U35345 ( .A(n35115), .B(n35116), .Z(n34897) );
  NANDN U35346 ( .A(n35117), .B(n35118), .Z(n35116) );
  NANDN U35347 ( .A(n35119), .B(n35120), .Z(n35118) );
  NANDN U35348 ( .A(n35120), .B(n35119), .Z(n35115) );
  ANDN U35349 ( .B(B[148]), .A(n58), .Z(n34899) );
  XNOR U35350 ( .A(n34907), .B(n35121), .Z(n34900) );
  XNOR U35351 ( .A(n34906), .B(n34904), .Z(n35121) );
  AND U35352 ( .A(n35122), .B(n35123), .Z(n34904) );
  NANDN U35353 ( .A(n35124), .B(n35125), .Z(n35123) );
  OR U35354 ( .A(n35126), .B(n35127), .Z(n35125) );
  NAND U35355 ( .A(n35127), .B(n35126), .Z(n35122) );
  ANDN U35356 ( .B(B[149]), .A(n59), .Z(n34906) );
  XNOR U35357 ( .A(n34914), .B(n35128), .Z(n34907) );
  XNOR U35358 ( .A(n34913), .B(n34911), .Z(n35128) );
  AND U35359 ( .A(n35129), .B(n35130), .Z(n34911) );
  NANDN U35360 ( .A(n35131), .B(n35132), .Z(n35130) );
  NANDN U35361 ( .A(n35133), .B(n35134), .Z(n35132) );
  NANDN U35362 ( .A(n35134), .B(n35133), .Z(n35129) );
  ANDN U35363 ( .B(B[150]), .A(n60), .Z(n34913) );
  XNOR U35364 ( .A(n34921), .B(n35135), .Z(n34914) );
  XNOR U35365 ( .A(n34920), .B(n34918), .Z(n35135) );
  AND U35366 ( .A(n35136), .B(n35137), .Z(n34918) );
  NANDN U35367 ( .A(n35138), .B(n35139), .Z(n35137) );
  OR U35368 ( .A(n35140), .B(n35141), .Z(n35139) );
  NAND U35369 ( .A(n35141), .B(n35140), .Z(n35136) );
  ANDN U35370 ( .B(B[151]), .A(n61), .Z(n34920) );
  XNOR U35371 ( .A(n34928), .B(n35142), .Z(n34921) );
  XNOR U35372 ( .A(n34927), .B(n34925), .Z(n35142) );
  AND U35373 ( .A(n35143), .B(n35144), .Z(n34925) );
  NANDN U35374 ( .A(n35145), .B(n35146), .Z(n35144) );
  NANDN U35375 ( .A(n35147), .B(n35148), .Z(n35146) );
  NANDN U35376 ( .A(n35148), .B(n35147), .Z(n35143) );
  ANDN U35377 ( .B(B[152]), .A(n62), .Z(n34927) );
  XNOR U35378 ( .A(n34935), .B(n35149), .Z(n34928) );
  XNOR U35379 ( .A(n34934), .B(n34932), .Z(n35149) );
  AND U35380 ( .A(n35150), .B(n35151), .Z(n34932) );
  NANDN U35381 ( .A(n35152), .B(n35153), .Z(n35151) );
  OR U35382 ( .A(n35154), .B(n35155), .Z(n35153) );
  NAND U35383 ( .A(n35155), .B(n35154), .Z(n35150) );
  ANDN U35384 ( .B(B[153]), .A(n63), .Z(n34934) );
  XNOR U35385 ( .A(n34942), .B(n35156), .Z(n34935) );
  XNOR U35386 ( .A(n34941), .B(n34939), .Z(n35156) );
  AND U35387 ( .A(n35157), .B(n35158), .Z(n34939) );
  NANDN U35388 ( .A(n35159), .B(n35160), .Z(n35158) );
  NANDN U35389 ( .A(n35161), .B(n35162), .Z(n35160) );
  NANDN U35390 ( .A(n35162), .B(n35161), .Z(n35157) );
  ANDN U35391 ( .B(B[154]), .A(n64), .Z(n34941) );
  XNOR U35392 ( .A(n34949), .B(n35163), .Z(n34942) );
  XNOR U35393 ( .A(n34948), .B(n34946), .Z(n35163) );
  AND U35394 ( .A(n35164), .B(n35165), .Z(n34946) );
  NANDN U35395 ( .A(n35166), .B(n35167), .Z(n35165) );
  OR U35396 ( .A(n35168), .B(n35169), .Z(n35167) );
  NAND U35397 ( .A(n35169), .B(n35168), .Z(n35164) );
  ANDN U35398 ( .B(B[155]), .A(n65), .Z(n34948) );
  XNOR U35399 ( .A(n34956), .B(n35170), .Z(n34949) );
  XNOR U35400 ( .A(n34955), .B(n34953), .Z(n35170) );
  AND U35401 ( .A(n35171), .B(n35172), .Z(n34953) );
  NANDN U35402 ( .A(n35173), .B(n35174), .Z(n35172) );
  NANDN U35403 ( .A(n35175), .B(n35176), .Z(n35174) );
  NANDN U35404 ( .A(n35176), .B(n35175), .Z(n35171) );
  ANDN U35405 ( .B(B[156]), .A(n66), .Z(n34955) );
  XNOR U35406 ( .A(n34963), .B(n35177), .Z(n34956) );
  XNOR U35407 ( .A(n34962), .B(n34960), .Z(n35177) );
  AND U35408 ( .A(n35178), .B(n35179), .Z(n34960) );
  NANDN U35409 ( .A(n35180), .B(n35181), .Z(n35179) );
  OR U35410 ( .A(n35182), .B(n35183), .Z(n35181) );
  NAND U35411 ( .A(n35183), .B(n35182), .Z(n35178) );
  ANDN U35412 ( .B(B[157]), .A(n67), .Z(n34962) );
  XNOR U35413 ( .A(n34970), .B(n35184), .Z(n34963) );
  XNOR U35414 ( .A(n34969), .B(n34967), .Z(n35184) );
  AND U35415 ( .A(n35185), .B(n35186), .Z(n34967) );
  NANDN U35416 ( .A(n35187), .B(n35188), .Z(n35186) );
  NANDN U35417 ( .A(n35189), .B(n35190), .Z(n35188) );
  NANDN U35418 ( .A(n35190), .B(n35189), .Z(n35185) );
  ANDN U35419 ( .B(B[158]), .A(n68), .Z(n34969) );
  XNOR U35420 ( .A(n34977), .B(n35191), .Z(n34970) );
  XNOR U35421 ( .A(n34976), .B(n34974), .Z(n35191) );
  AND U35422 ( .A(n35192), .B(n35193), .Z(n34974) );
  NANDN U35423 ( .A(n35194), .B(n35195), .Z(n35193) );
  OR U35424 ( .A(n35196), .B(n35197), .Z(n35195) );
  NAND U35425 ( .A(n35197), .B(n35196), .Z(n35192) );
  ANDN U35426 ( .B(B[159]), .A(n69), .Z(n34976) );
  XNOR U35427 ( .A(n34984), .B(n35198), .Z(n34977) );
  XNOR U35428 ( .A(n34983), .B(n34981), .Z(n35198) );
  AND U35429 ( .A(n35199), .B(n35200), .Z(n34981) );
  NANDN U35430 ( .A(n35201), .B(n35202), .Z(n35200) );
  NANDN U35431 ( .A(n35203), .B(n35204), .Z(n35202) );
  NANDN U35432 ( .A(n35204), .B(n35203), .Z(n35199) );
  ANDN U35433 ( .B(B[160]), .A(n70), .Z(n34983) );
  XNOR U35434 ( .A(n34991), .B(n35205), .Z(n34984) );
  XNOR U35435 ( .A(n34990), .B(n34988), .Z(n35205) );
  AND U35436 ( .A(n35206), .B(n35207), .Z(n34988) );
  NANDN U35437 ( .A(n35208), .B(n35209), .Z(n35207) );
  OR U35438 ( .A(n35210), .B(n35211), .Z(n35209) );
  NAND U35439 ( .A(n35211), .B(n35210), .Z(n35206) );
  ANDN U35440 ( .B(B[161]), .A(n71), .Z(n34990) );
  XNOR U35441 ( .A(n34998), .B(n35212), .Z(n34991) );
  XNOR U35442 ( .A(n34997), .B(n34995), .Z(n35212) );
  AND U35443 ( .A(n35213), .B(n35214), .Z(n34995) );
  NANDN U35444 ( .A(n35215), .B(n35216), .Z(n35214) );
  NANDN U35445 ( .A(n35217), .B(n35218), .Z(n35216) );
  NANDN U35446 ( .A(n35218), .B(n35217), .Z(n35213) );
  ANDN U35447 ( .B(B[162]), .A(n72), .Z(n34997) );
  XNOR U35448 ( .A(n35005), .B(n35219), .Z(n34998) );
  XNOR U35449 ( .A(n35004), .B(n35002), .Z(n35219) );
  AND U35450 ( .A(n35220), .B(n35221), .Z(n35002) );
  NANDN U35451 ( .A(n35222), .B(n35223), .Z(n35221) );
  OR U35452 ( .A(n35224), .B(n35225), .Z(n35223) );
  NAND U35453 ( .A(n35225), .B(n35224), .Z(n35220) );
  ANDN U35454 ( .B(B[163]), .A(n73), .Z(n35004) );
  XNOR U35455 ( .A(n35012), .B(n35226), .Z(n35005) );
  XNOR U35456 ( .A(n35011), .B(n35009), .Z(n35226) );
  AND U35457 ( .A(n35227), .B(n35228), .Z(n35009) );
  NANDN U35458 ( .A(n35229), .B(n35230), .Z(n35228) );
  NANDN U35459 ( .A(n35231), .B(n35232), .Z(n35230) );
  NANDN U35460 ( .A(n35232), .B(n35231), .Z(n35227) );
  ANDN U35461 ( .B(B[164]), .A(n74), .Z(n35011) );
  XNOR U35462 ( .A(n35019), .B(n35233), .Z(n35012) );
  XNOR U35463 ( .A(n35018), .B(n35016), .Z(n35233) );
  AND U35464 ( .A(n35234), .B(n35235), .Z(n35016) );
  NANDN U35465 ( .A(n35236), .B(n35237), .Z(n35235) );
  OR U35466 ( .A(n35238), .B(n35239), .Z(n35237) );
  NAND U35467 ( .A(n35239), .B(n35238), .Z(n35234) );
  ANDN U35468 ( .B(B[165]), .A(n75), .Z(n35018) );
  XNOR U35469 ( .A(n35026), .B(n35240), .Z(n35019) );
  XNOR U35470 ( .A(n35025), .B(n35023), .Z(n35240) );
  AND U35471 ( .A(n35241), .B(n35242), .Z(n35023) );
  NANDN U35472 ( .A(n35243), .B(n35244), .Z(n35242) );
  NANDN U35473 ( .A(n35245), .B(n35246), .Z(n35244) );
  NANDN U35474 ( .A(n35246), .B(n35245), .Z(n35241) );
  ANDN U35475 ( .B(B[166]), .A(n76), .Z(n35025) );
  XNOR U35476 ( .A(n35033), .B(n35247), .Z(n35026) );
  XNOR U35477 ( .A(n35032), .B(n35030), .Z(n35247) );
  AND U35478 ( .A(n35248), .B(n35249), .Z(n35030) );
  NANDN U35479 ( .A(n35250), .B(n35251), .Z(n35249) );
  OR U35480 ( .A(n35252), .B(n35253), .Z(n35251) );
  NAND U35481 ( .A(n35253), .B(n35252), .Z(n35248) );
  ANDN U35482 ( .B(B[167]), .A(n77), .Z(n35032) );
  XNOR U35483 ( .A(n35040), .B(n35254), .Z(n35033) );
  XNOR U35484 ( .A(n35039), .B(n35037), .Z(n35254) );
  AND U35485 ( .A(n35255), .B(n35256), .Z(n35037) );
  NANDN U35486 ( .A(n35257), .B(n35258), .Z(n35256) );
  NANDN U35487 ( .A(n35259), .B(n35260), .Z(n35258) );
  NANDN U35488 ( .A(n35260), .B(n35259), .Z(n35255) );
  ANDN U35489 ( .B(B[168]), .A(n78), .Z(n35039) );
  XNOR U35490 ( .A(n35047), .B(n35261), .Z(n35040) );
  XNOR U35491 ( .A(n35046), .B(n35044), .Z(n35261) );
  AND U35492 ( .A(n35262), .B(n35263), .Z(n35044) );
  NANDN U35493 ( .A(n35264), .B(n35265), .Z(n35263) );
  OR U35494 ( .A(n35266), .B(n35267), .Z(n35265) );
  NAND U35495 ( .A(n35267), .B(n35266), .Z(n35262) );
  ANDN U35496 ( .B(B[169]), .A(n79), .Z(n35046) );
  XNOR U35497 ( .A(n35054), .B(n35268), .Z(n35047) );
  XNOR U35498 ( .A(n35053), .B(n35051), .Z(n35268) );
  AND U35499 ( .A(n35269), .B(n35270), .Z(n35051) );
  NANDN U35500 ( .A(n35271), .B(n35272), .Z(n35270) );
  NANDN U35501 ( .A(n35273), .B(n35274), .Z(n35272) );
  NANDN U35502 ( .A(n35274), .B(n35273), .Z(n35269) );
  ANDN U35503 ( .B(B[170]), .A(n80), .Z(n35053) );
  XNOR U35504 ( .A(n35061), .B(n35275), .Z(n35054) );
  XNOR U35505 ( .A(n35060), .B(n35058), .Z(n35275) );
  AND U35506 ( .A(n35276), .B(n35277), .Z(n35058) );
  NANDN U35507 ( .A(n35278), .B(n35279), .Z(n35277) );
  OR U35508 ( .A(n35280), .B(n35281), .Z(n35279) );
  NAND U35509 ( .A(n35281), .B(n35280), .Z(n35276) );
  ANDN U35510 ( .B(B[171]), .A(n81), .Z(n35060) );
  XNOR U35511 ( .A(n35068), .B(n35282), .Z(n35061) );
  XNOR U35512 ( .A(n35067), .B(n35065), .Z(n35282) );
  AND U35513 ( .A(n35283), .B(n35284), .Z(n35065) );
  NANDN U35514 ( .A(n35285), .B(n35286), .Z(n35284) );
  NAND U35515 ( .A(n35287), .B(n35288), .Z(n35286) );
  ANDN U35516 ( .B(B[172]), .A(n82), .Z(n35067) );
  XOR U35517 ( .A(n35074), .B(n35289), .Z(n35068) );
  XNOR U35518 ( .A(n35072), .B(n35075), .Z(n35289) );
  NAND U35519 ( .A(A[2]), .B(B[173]), .Z(n35075) );
  NANDN U35520 ( .A(n35290), .B(n35291), .Z(n35072) );
  AND U35521 ( .A(A[0]), .B(B[174]), .Z(n35291) );
  XNOR U35522 ( .A(n35077), .B(n35292), .Z(n35074) );
  NAND U35523 ( .A(A[0]), .B(B[175]), .Z(n35292) );
  NAND U35524 ( .A(B[174]), .B(A[1]), .Z(n35077) );
  NAND U35525 ( .A(n35293), .B(n35294), .Z(n446) );
  NANDN U35526 ( .A(n35295), .B(n35296), .Z(n35294) );
  OR U35527 ( .A(n35297), .B(n35298), .Z(n35296) );
  NAND U35528 ( .A(n35298), .B(n35297), .Z(n35293) );
  XOR U35529 ( .A(n448), .B(n447), .Z(\A1[172] ) );
  XOR U35530 ( .A(n35298), .B(n35299), .Z(n447) );
  XNOR U35531 ( .A(n35297), .B(n35295), .Z(n35299) );
  AND U35532 ( .A(n35300), .B(n35301), .Z(n35295) );
  NANDN U35533 ( .A(n35302), .B(n35303), .Z(n35301) );
  NANDN U35534 ( .A(n35304), .B(n35305), .Z(n35303) );
  NANDN U35535 ( .A(n35305), .B(n35304), .Z(n35300) );
  ANDN U35536 ( .B(B[143]), .A(n54), .Z(n35297) );
  XNOR U35537 ( .A(n35092), .B(n35306), .Z(n35298) );
  XNOR U35538 ( .A(n35091), .B(n35089), .Z(n35306) );
  AND U35539 ( .A(n35307), .B(n35308), .Z(n35089) );
  NANDN U35540 ( .A(n35309), .B(n35310), .Z(n35308) );
  OR U35541 ( .A(n35311), .B(n35312), .Z(n35310) );
  NAND U35542 ( .A(n35312), .B(n35311), .Z(n35307) );
  ANDN U35543 ( .B(B[144]), .A(n55), .Z(n35091) );
  XNOR U35544 ( .A(n35099), .B(n35313), .Z(n35092) );
  XNOR U35545 ( .A(n35098), .B(n35096), .Z(n35313) );
  AND U35546 ( .A(n35314), .B(n35315), .Z(n35096) );
  NANDN U35547 ( .A(n35316), .B(n35317), .Z(n35315) );
  NANDN U35548 ( .A(n35318), .B(n35319), .Z(n35317) );
  NANDN U35549 ( .A(n35319), .B(n35318), .Z(n35314) );
  ANDN U35550 ( .B(B[145]), .A(n56), .Z(n35098) );
  XNOR U35551 ( .A(n35106), .B(n35320), .Z(n35099) );
  XNOR U35552 ( .A(n35105), .B(n35103), .Z(n35320) );
  AND U35553 ( .A(n35321), .B(n35322), .Z(n35103) );
  NANDN U35554 ( .A(n35323), .B(n35324), .Z(n35322) );
  OR U35555 ( .A(n35325), .B(n35326), .Z(n35324) );
  NAND U35556 ( .A(n35326), .B(n35325), .Z(n35321) );
  ANDN U35557 ( .B(B[146]), .A(n57), .Z(n35105) );
  XNOR U35558 ( .A(n35113), .B(n35327), .Z(n35106) );
  XNOR U35559 ( .A(n35112), .B(n35110), .Z(n35327) );
  AND U35560 ( .A(n35328), .B(n35329), .Z(n35110) );
  NANDN U35561 ( .A(n35330), .B(n35331), .Z(n35329) );
  NANDN U35562 ( .A(n35332), .B(n35333), .Z(n35331) );
  NANDN U35563 ( .A(n35333), .B(n35332), .Z(n35328) );
  ANDN U35564 ( .B(B[147]), .A(n58), .Z(n35112) );
  XNOR U35565 ( .A(n35120), .B(n35334), .Z(n35113) );
  XNOR U35566 ( .A(n35119), .B(n35117), .Z(n35334) );
  AND U35567 ( .A(n35335), .B(n35336), .Z(n35117) );
  NANDN U35568 ( .A(n35337), .B(n35338), .Z(n35336) );
  OR U35569 ( .A(n35339), .B(n35340), .Z(n35338) );
  NAND U35570 ( .A(n35340), .B(n35339), .Z(n35335) );
  ANDN U35571 ( .B(B[148]), .A(n59), .Z(n35119) );
  XNOR U35572 ( .A(n35127), .B(n35341), .Z(n35120) );
  XNOR U35573 ( .A(n35126), .B(n35124), .Z(n35341) );
  AND U35574 ( .A(n35342), .B(n35343), .Z(n35124) );
  NANDN U35575 ( .A(n35344), .B(n35345), .Z(n35343) );
  NANDN U35576 ( .A(n35346), .B(n35347), .Z(n35345) );
  NANDN U35577 ( .A(n35347), .B(n35346), .Z(n35342) );
  ANDN U35578 ( .B(B[149]), .A(n60), .Z(n35126) );
  XNOR U35579 ( .A(n35134), .B(n35348), .Z(n35127) );
  XNOR U35580 ( .A(n35133), .B(n35131), .Z(n35348) );
  AND U35581 ( .A(n35349), .B(n35350), .Z(n35131) );
  NANDN U35582 ( .A(n35351), .B(n35352), .Z(n35350) );
  OR U35583 ( .A(n35353), .B(n35354), .Z(n35352) );
  NAND U35584 ( .A(n35354), .B(n35353), .Z(n35349) );
  ANDN U35585 ( .B(B[150]), .A(n61), .Z(n35133) );
  XNOR U35586 ( .A(n35141), .B(n35355), .Z(n35134) );
  XNOR U35587 ( .A(n35140), .B(n35138), .Z(n35355) );
  AND U35588 ( .A(n35356), .B(n35357), .Z(n35138) );
  NANDN U35589 ( .A(n35358), .B(n35359), .Z(n35357) );
  NANDN U35590 ( .A(n35360), .B(n35361), .Z(n35359) );
  NANDN U35591 ( .A(n35361), .B(n35360), .Z(n35356) );
  ANDN U35592 ( .B(B[151]), .A(n62), .Z(n35140) );
  XNOR U35593 ( .A(n35148), .B(n35362), .Z(n35141) );
  XNOR U35594 ( .A(n35147), .B(n35145), .Z(n35362) );
  AND U35595 ( .A(n35363), .B(n35364), .Z(n35145) );
  NANDN U35596 ( .A(n35365), .B(n35366), .Z(n35364) );
  OR U35597 ( .A(n35367), .B(n35368), .Z(n35366) );
  NAND U35598 ( .A(n35368), .B(n35367), .Z(n35363) );
  ANDN U35599 ( .B(B[152]), .A(n63), .Z(n35147) );
  XNOR U35600 ( .A(n35155), .B(n35369), .Z(n35148) );
  XNOR U35601 ( .A(n35154), .B(n35152), .Z(n35369) );
  AND U35602 ( .A(n35370), .B(n35371), .Z(n35152) );
  NANDN U35603 ( .A(n35372), .B(n35373), .Z(n35371) );
  NANDN U35604 ( .A(n35374), .B(n35375), .Z(n35373) );
  NANDN U35605 ( .A(n35375), .B(n35374), .Z(n35370) );
  ANDN U35606 ( .B(B[153]), .A(n64), .Z(n35154) );
  XNOR U35607 ( .A(n35162), .B(n35376), .Z(n35155) );
  XNOR U35608 ( .A(n35161), .B(n35159), .Z(n35376) );
  AND U35609 ( .A(n35377), .B(n35378), .Z(n35159) );
  NANDN U35610 ( .A(n35379), .B(n35380), .Z(n35378) );
  OR U35611 ( .A(n35381), .B(n35382), .Z(n35380) );
  NAND U35612 ( .A(n35382), .B(n35381), .Z(n35377) );
  ANDN U35613 ( .B(B[154]), .A(n65), .Z(n35161) );
  XNOR U35614 ( .A(n35169), .B(n35383), .Z(n35162) );
  XNOR U35615 ( .A(n35168), .B(n35166), .Z(n35383) );
  AND U35616 ( .A(n35384), .B(n35385), .Z(n35166) );
  NANDN U35617 ( .A(n35386), .B(n35387), .Z(n35385) );
  NANDN U35618 ( .A(n35388), .B(n35389), .Z(n35387) );
  NANDN U35619 ( .A(n35389), .B(n35388), .Z(n35384) );
  ANDN U35620 ( .B(B[155]), .A(n66), .Z(n35168) );
  XNOR U35621 ( .A(n35176), .B(n35390), .Z(n35169) );
  XNOR U35622 ( .A(n35175), .B(n35173), .Z(n35390) );
  AND U35623 ( .A(n35391), .B(n35392), .Z(n35173) );
  NANDN U35624 ( .A(n35393), .B(n35394), .Z(n35392) );
  OR U35625 ( .A(n35395), .B(n35396), .Z(n35394) );
  NAND U35626 ( .A(n35396), .B(n35395), .Z(n35391) );
  ANDN U35627 ( .B(B[156]), .A(n67), .Z(n35175) );
  XNOR U35628 ( .A(n35183), .B(n35397), .Z(n35176) );
  XNOR U35629 ( .A(n35182), .B(n35180), .Z(n35397) );
  AND U35630 ( .A(n35398), .B(n35399), .Z(n35180) );
  NANDN U35631 ( .A(n35400), .B(n35401), .Z(n35399) );
  NANDN U35632 ( .A(n35402), .B(n35403), .Z(n35401) );
  NANDN U35633 ( .A(n35403), .B(n35402), .Z(n35398) );
  ANDN U35634 ( .B(B[157]), .A(n68), .Z(n35182) );
  XNOR U35635 ( .A(n35190), .B(n35404), .Z(n35183) );
  XNOR U35636 ( .A(n35189), .B(n35187), .Z(n35404) );
  AND U35637 ( .A(n35405), .B(n35406), .Z(n35187) );
  NANDN U35638 ( .A(n35407), .B(n35408), .Z(n35406) );
  OR U35639 ( .A(n35409), .B(n35410), .Z(n35408) );
  NAND U35640 ( .A(n35410), .B(n35409), .Z(n35405) );
  ANDN U35641 ( .B(B[158]), .A(n69), .Z(n35189) );
  XNOR U35642 ( .A(n35197), .B(n35411), .Z(n35190) );
  XNOR U35643 ( .A(n35196), .B(n35194), .Z(n35411) );
  AND U35644 ( .A(n35412), .B(n35413), .Z(n35194) );
  NANDN U35645 ( .A(n35414), .B(n35415), .Z(n35413) );
  NANDN U35646 ( .A(n35416), .B(n35417), .Z(n35415) );
  NANDN U35647 ( .A(n35417), .B(n35416), .Z(n35412) );
  ANDN U35648 ( .B(B[159]), .A(n70), .Z(n35196) );
  XNOR U35649 ( .A(n35204), .B(n35418), .Z(n35197) );
  XNOR U35650 ( .A(n35203), .B(n35201), .Z(n35418) );
  AND U35651 ( .A(n35419), .B(n35420), .Z(n35201) );
  NANDN U35652 ( .A(n35421), .B(n35422), .Z(n35420) );
  OR U35653 ( .A(n35423), .B(n35424), .Z(n35422) );
  NAND U35654 ( .A(n35424), .B(n35423), .Z(n35419) );
  ANDN U35655 ( .B(B[160]), .A(n71), .Z(n35203) );
  XNOR U35656 ( .A(n35211), .B(n35425), .Z(n35204) );
  XNOR U35657 ( .A(n35210), .B(n35208), .Z(n35425) );
  AND U35658 ( .A(n35426), .B(n35427), .Z(n35208) );
  NANDN U35659 ( .A(n35428), .B(n35429), .Z(n35427) );
  NANDN U35660 ( .A(n35430), .B(n35431), .Z(n35429) );
  NANDN U35661 ( .A(n35431), .B(n35430), .Z(n35426) );
  ANDN U35662 ( .B(B[161]), .A(n72), .Z(n35210) );
  XNOR U35663 ( .A(n35218), .B(n35432), .Z(n35211) );
  XNOR U35664 ( .A(n35217), .B(n35215), .Z(n35432) );
  AND U35665 ( .A(n35433), .B(n35434), .Z(n35215) );
  NANDN U35666 ( .A(n35435), .B(n35436), .Z(n35434) );
  OR U35667 ( .A(n35437), .B(n35438), .Z(n35436) );
  NAND U35668 ( .A(n35438), .B(n35437), .Z(n35433) );
  ANDN U35669 ( .B(B[162]), .A(n73), .Z(n35217) );
  XNOR U35670 ( .A(n35225), .B(n35439), .Z(n35218) );
  XNOR U35671 ( .A(n35224), .B(n35222), .Z(n35439) );
  AND U35672 ( .A(n35440), .B(n35441), .Z(n35222) );
  NANDN U35673 ( .A(n35442), .B(n35443), .Z(n35441) );
  NANDN U35674 ( .A(n35444), .B(n35445), .Z(n35443) );
  NANDN U35675 ( .A(n35445), .B(n35444), .Z(n35440) );
  ANDN U35676 ( .B(B[163]), .A(n74), .Z(n35224) );
  XNOR U35677 ( .A(n35232), .B(n35446), .Z(n35225) );
  XNOR U35678 ( .A(n35231), .B(n35229), .Z(n35446) );
  AND U35679 ( .A(n35447), .B(n35448), .Z(n35229) );
  NANDN U35680 ( .A(n35449), .B(n35450), .Z(n35448) );
  OR U35681 ( .A(n35451), .B(n35452), .Z(n35450) );
  NAND U35682 ( .A(n35452), .B(n35451), .Z(n35447) );
  ANDN U35683 ( .B(B[164]), .A(n75), .Z(n35231) );
  XNOR U35684 ( .A(n35239), .B(n35453), .Z(n35232) );
  XNOR U35685 ( .A(n35238), .B(n35236), .Z(n35453) );
  AND U35686 ( .A(n35454), .B(n35455), .Z(n35236) );
  NANDN U35687 ( .A(n35456), .B(n35457), .Z(n35455) );
  NANDN U35688 ( .A(n35458), .B(n35459), .Z(n35457) );
  NANDN U35689 ( .A(n35459), .B(n35458), .Z(n35454) );
  ANDN U35690 ( .B(B[165]), .A(n76), .Z(n35238) );
  XNOR U35691 ( .A(n35246), .B(n35460), .Z(n35239) );
  XNOR U35692 ( .A(n35245), .B(n35243), .Z(n35460) );
  AND U35693 ( .A(n35461), .B(n35462), .Z(n35243) );
  NANDN U35694 ( .A(n35463), .B(n35464), .Z(n35462) );
  OR U35695 ( .A(n35465), .B(n35466), .Z(n35464) );
  NAND U35696 ( .A(n35466), .B(n35465), .Z(n35461) );
  ANDN U35697 ( .B(B[166]), .A(n77), .Z(n35245) );
  XNOR U35698 ( .A(n35253), .B(n35467), .Z(n35246) );
  XNOR U35699 ( .A(n35252), .B(n35250), .Z(n35467) );
  AND U35700 ( .A(n35468), .B(n35469), .Z(n35250) );
  NANDN U35701 ( .A(n35470), .B(n35471), .Z(n35469) );
  NANDN U35702 ( .A(n35472), .B(n35473), .Z(n35471) );
  NANDN U35703 ( .A(n35473), .B(n35472), .Z(n35468) );
  ANDN U35704 ( .B(B[167]), .A(n78), .Z(n35252) );
  XNOR U35705 ( .A(n35260), .B(n35474), .Z(n35253) );
  XNOR U35706 ( .A(n35259), .B(n35257), .Z(n35474) );
  AND U35707 ( .A(n35475), .B(n35476), .Z(n35257) );
  NANDN U35708 ( .A(n35477), .B(n35478), .Z(n35476) );
  OR U35709 ( .A(n35479), .B(n35480), .Z(n35478) );
  NAND U35710 ( .A(n35480), .B(n35479), .Z(n35475) );
  ANDN U35711 ( .B(B[168]), .A(n79), .Z(n35259) );
  XNOR U35712 ( .A(n35267), .B(n35481), .Z(n35260) );
  XNOR U35713 ( .A(n35266), .B(n35264), .Z(n35481) );
  AND U35714 ( .A(n35482), .B(n35483), .Z(n35264) );
  NANDN U35715 ( .A(n35484), .B(n35485), .Z(n35483) );
  NANDN U35716 ( .A(n35486), .B(n35487), .Z(n35485) );
  NANDN U35717 ( .A(n35487), .B(n35486), .Z(n35482) );
  ANDN U35718 ( .B(B[169]), .A(n80), .Z(n35266) );
  XNOR U35719 ( .A(n35274), .B(n35488), .Z(n35267) );
  XNOR U35720 ( .A(n35273), .B(n35271), .Z(n35488) );
  AND U35721 ( .A(n35489), .B(n35490), .Z(n35271) );
  NANDN U35722 ( .A(n35491), .B(n35492), .Z(n35490) );
  OR U35723 ( .A(n35493), .B(n35494), .Z(n35492) );
  NAND U35724 ( .A(n35494), .B(n35493), .Z(n35489) );
  ANDN U35725 ( .B(B[170]), .A(n81), .Z(n35273) );
  XNOR U35726 ( .A(n35281), .B(n35495), .Z(n35274) );
  XNOR U35727 ( .A(n35280), .B(n35278), .Z(n35495) );
  AND U35728 ( .A(n35496), .B(n35497), .Z(n35278) );
  NANDN U35729 ( .A(n35498), .B(n35499), .Z(n35497) );
  NAND U35730 ( .A(n35500), .B(n35501), .Z(n35499) );
  ANDN U35731 ( .B(B[171]), .A(n82), .Z(n35280) );
  XOR U35732 ( .A(n35287), .B(n35502), .Z(n35281) );
  XNOR U35733 ( .A(n35285), .B(n35288), .Z(n35502) );
  NAND U35734 ( .A(A[2]), .B(B[172]), .Z(n35288) );
  NANDN U35735 ( .A(n35503), .B(n35504), .Z(n35285) );
  AND U35736 ( .A(A[0]), .B(B[173]), .Z(n35504) );
  XNOR U35737 ( .A(n35290), .B(n35505), .Z(n35287) );
  NAND U35738 ( .A(A[0]), .B(B[174]), .Z(n35505) );
  NAND U35739 ( .A(B[173]), .B(A[1]), .Z(n35290) );
  NAND U35740 ( .A(n35506), .B(n35507), .Z(n448) );
  NANDN U35741 ( .A(n35508), .B(n35509), .Z(n35507) );
  OR U35742 ( .A(n35510), .B(n35511), .Z(n35509) );
  NAND U35743 ( .A(n35511), .B(n35510), .Z(n35506) );
  XOR U35744 ( .A(n450), .B(n449), .Z(\A1[171] ) );
  XOR U35745 ( .A(n35511), .B(n35512), .Z(n449) );
  XNOR U35746 ( .A(n35510), .B(n35508), .Z(n35512) );
  AND U35747 ( .A(n35513), .B(n35514), .Z(n35508) );
  NANDN U35748 ( .A(n35515), .B(n35516), .Z(n35514) );
  NANDN U35749 ( .A(n35517), .B(n35518), .Z(n35516) );
  NANDN U35750 ( .A(n35518), .B(n35517), .Z(n35513) );
  ANDN U35751 ( .B(B[142]), .A(n54), .Z(n35510) );
  XNOR U35752 ( .A(n35305), .B(n35519), .Z(n35511) );
  XNOR U35753 ( .A(n35304), .B(n35302), .Z(n35519) );
  AND U35754 ( .A(n35520), .B(n35521), .Z(n35302) );
  NANDN U35755 ( .A(n35522), .B(n35523), .Z(n35521) );
  OR U35756 ( .A(n35524), .B(n35525), .Z(n35523) );
  NAND U35757 ( .A(n35525), .B(n35524), .Z(n35520) );
  ANDN U35758 ( .B(B[143]), .A(n55), .Z(n35304) );
  XNOR U35759 ( .A(n35312), .B(n35526), .Z(n35305) );
  XNOR U35760 ( .A(n35311), .B(n35309), .Z(n35526) );
  AND U35761 ( .A(n35527), .B(n35528), .Z(n35309) );
  NANDN U35762 ( .A(n35529), .B(n35530), .Z(n35528) );
  NANDN U35763 ( .A(n35531), .B(n35532), .Z(n35530) );
  NANDN U35764 ( .A(n35532), .B(n35531), .Z(n35527) );
  ANDN U35765 ( .B(B[144]), .A(n56), .Z(n35311) );
  XNOR U35766 ( .A(n35319), .B(n35533), .Z(n35312) );
  XNOR U35767 ( .A(n35318), .B(n35316), .Z(n35533) );
  AND U35768 ( .A(n35534), .B(n35535), .Z(n35316) );
  NANDN U35769 ( .A(n35536), .B(n35537), .Z(n35535) );
  OR U35770 ( .A(n35538), .B(n35539), .Z(n35537) );
  NAND U35771 ( .A(n35539), .B(n35538), .Z(n35534) );
  ANDN U35772 ( .B(B[145]), .A(n57), .Z(n35318) );
  XNOR U35773 ( .A(n35326), .B(n35540), .Z(n35319) );
  XNOR U35774 ( .A(n35325), .B(n35323), .Z(n35540) );
  AND U35775 ( .A(n35541), .B(n35542), .Z(n35323) );
  NANDN U35776 ( .A(n35543), .B(n35544), .Z(n35542) );
  NANDN U35777 ( .A(n35545), .B(n35546), .Z(n35544) );
  NANDN U35778 ( .A(n35546), .B(n35545), .Z(n35541) );
  ANDN U35779 ( .B(B[146]), .A(n58), .Z(n35325) );
  XNOR U35780 ( .A(n35333), .B(n35547), .Z(n35326) );
  XNOR U35781 ( .A(n35332), .B(n35330), .Z(n35547) );
  AND U35782 ( .A(n35548), .B(n35549), .Z(n35330) );
  NANDN U35783 ( .A(n35550), .B(n35551), .Z(n35549) );
  OR U35784 ( .A(n35552), .B(n35553), .Z(n35551) );
  NAND U35785 ( .A(n35553), .B(n35552), .Z(n35548) );
  ANDN U35786 ( .B(B[147]), .A(n59), .Z(n35332) );
  XNOR U35787 ( .A(n35340), .B(n35554), .Z(n35333) );
  XNOR U35788 ( .A(n35339), .B(n35337), .Z(n35554) );
  AND U35789 ( .A(n35555), .B(n35556), .Z(n35337) );
  NANDN U35790 ( .A(n35557), .B(n35558), .Z(n35556) );
  NANDN U35791 ( .A(n35559), .B(n35560), .Z(n35558) );
  NANDN U35792 ( .A(n35560), .B(n35559), .Z(n35555) );
  ANDN U35793 ( .B(B[148]), .A(n60), .Z(n35339) );
  XNOR U35794 ( .A(n35347), .B(n35561), .Z(n35340) );
  XNOR U35795 ( .A(n35346), .B(n35344), .Z(n35561) );
  AND U35796 ( .A(n35562), .B(n35563), .Z(n35344) );
  NANDN U35797 ( .A(n35564), .B(n35565), .Z(n35563) );
  OR U35798 ( .A(n35566), .B(n35567), .Z(n35565) );
  NAND U35799 ( .A(n35567), .B(n35566), .Z(n35562) );
  ANDN U35800 ( .B(B[149]), .A(n61), .Z(n35346) );
  XNOR U35801 ( .A(n35354), .B(n35568), .Z(n35347) );
  XNOR U35802 ( .A(n35353), .B(n35351), .Z(n35568) );
  AND U35803 ( .A(n35569), .B(n35570), .Z(n35351) );
  NANDN U35804 ( .A(n35571), .B(n35572), .Z(n35570) );
  NANDN U35805 ( .A(n35573), .B(n35574), .Z(n35572) );
  NANDN U35806 ( .A(n35574), .B(n35573), .Z(n35569) );
  ANDN U35807 ( .B(B[150]), .A(n62), .Z(n35353) );
  XNOR U35808 ( .A(n35361), .B(n35575), .Z(n35354) );
  XNOR U35809 ( .A(n35360), .B(n35358), .Z(n35575) );
  AND U35810 ( .A(n35576), .B(n35577), .Z(n35358) );
  NANDN U35811 ( .A(n35578), .B(n35579), .Z(n35577) );
  OR U35812 ( .A(n35580), .B(n35581), .Z(n35579) );
  NAND U35813 ( .A(n35581), .B(n35580), .Z(n35576) );
  ANDN U35814 ( .B(B[151]), .A(n63), .Z(n35360) );
  XNOR U35815 ( .A(n35368), .B(n35582), .Z(n35361) );
  XNOR U35816 ( .A(n35367), .B(n35365), .Z(n35582) );
  AND U35817 ( .A(n35583), .B(n35584), .Z(n35365) );
  NANDN U35818 ( .A(n35585), .B(n35586), .Z(n35584) );
  NANDN U35819 ( .A(n35587), .B(n35588), .Z(n35586) );
  NANDN U35820 ( .A(n35588), .B(n35587), .Z(n35583) );
  ANDN U35821 ( .B(B[152]), .A(n64), .Z(n35367) );
  XNOR U35822 ( .A(n35375), .B(n35589), .Z(n35368) );
  XNOR U35823 ( .A(n35374), .B(n35372), .Z(n35589) );
  AND U35824 ( .A(n35590), .B(n35591), .Z(n35372) );
  NANDN U35825 ( .A(n35592), .B(n35593), .Z(n35591) );
  OR U35826 ( .A(n35594), .B(n35595), .Z(n35593) );
  NAND U35827 ( .A(n35595), .B(n35594), .Z(n35590) );
  ANDN U35828 ( .B(B[153]), .A(n65), .Z(n35374) );
  XNOR U35829 ( .A(n35382), .B(n35596), .Z(n35375) );
  XNOR U35830 ( .A(n35381), .B(n35379), .Z(n35596) );
  AND U35831 ( .A(n35597), .B(n35598), .Z(n35379) );
  NANDN U35832 ( .A(n35599), .B(n35600), .Z(n35598) );
  NANDN U35833 ( .A(n35601), .B(n35602), .Z(n35600) );
  NANDN U35834 ( .A(n35602), .B(n35601), .Z(n35597) );
  ANDN U35835 ( .B(B[154]), .A(n66), .Z(n35381) );
  XNOR U35836 ( .A(n35389), .B(n35603), .Z(n35382) );
  XNOR U35837 ( .A(n35388), .B(n35386), .Z(n35603) );
  AND U35838 ( .A(n35604), .B(n35605), .Z(n35386) );
  NANDN U35839 ( .A(n35606), .B(n35607), .Z(n35605) );
  OR U35840 ( .A(n35608), .B(n35609), .Z(n35607) );
  NAND U35841 ( .A(n35609), .B(n35608), .Z(n35604) );
  ANDN U35842 ( .B(B[155]), .A(n67), .Z(n35388) );
  XNOR U35843 ( .A(n35396), .B(n35610), .Z(n35389) );
  XNOR U35844 ( .A(n35395), .B(n35393), .Z(n35610) );
  AND U35845 ( .A(n35611), .B(n35612), .Z(n35393) );
  NANDN U35846 ( .A(n35613), .B(n35614), .Z(n35612) );
  NANDN U35847 ( .A(n35615), .B(n35616), .Z(n35614) );
  NANDN U35848 ( .A(n35616), .B(n35615), .Z(n35611) );
  ANDN U35849 ( .B(B[156]), .A(n68), .Z(n35395) );
  XNOR U35850 ( .A(n35403), .B(n35617), .Z(n35396) );
  XNOR U35851 ( .A(n35402), .B(n35400), .Z(n35617) );
  AND U35852 ( .A(n35618), .B(n35619), .Z(n35400) );
  NANDN U35853 ( .A(n35620), .B(n35621), .Z(n35619) );
  OR U35854 ( .A(n35622), .B(n35623), .Z(n35621) );
  NAND U35855 ( .A(n35623), .B(n35622), .Z(n35618) );
  ANDN U35856 ( .B(B[157]), .A(n69), .Z(n35402) );
  XNOR U35857 ( .A(n35410), .B(n35624), .Z(n35403) );
  XNOR U35858 ( .A(n35409), .B(n35407), .Z(n35624) );
  AND U35859 ( .A(n35625), .B(n35626), .Z(n35407) );
  NANDN U35860 ( .A(n35627), .B(n35628), .Z(n35626) );
  NANDN U35861 ( .A(n35629), .B(n35630), .Z(n35628) );
  NANDN U35862 ( .A(n35630), .B(n35629), .Z(n35625) );
  ANDN U35863 ( .B(B[158]), .A(n70), .Z(n35409) );
  XNOR U35864 ( .A(n35417), .B(n35631), .Z(n35410) );
  XNOR U35865 ( .A(n35416), .B(n35414), .Z(n35631) );
  AND U35866 ( .A(n35632), .B(n35633), .Z(n35414) );
  NANDN U35867 ( .A(n35634), .B(n35635), .Z(n35633) );
  OR U35868 ( .A(n35636), .B(n35637), .Z(n35635) );
  NAND U35869 ( .A(n35637), .B(n35636), .Z(n35632) );
  ANDN U35870 ( .B(B[159]), .A(n71), .Z(n35416) );
  XNOR U35871 ( .A(n35424), .B(n35638), .Z(n35417) );
  XNOR U35872 ( .A(n35423), .B(n35421), .Z(n35638) );
  AND U35873 ( .A(n35639), .B(n35640), .Z(n35421) );
  NANDN U35874 ( .A(n35641), .B(n35642), .Z(n35640) );
  NANDN U35875 ( .A(n35643), .B(n35644), .Z(n35642) );
  NANDN U35876 ( .A(n35644), .B(n35643), .Z(n35639) );
  ANDN U35877 ( .B(B[160]), .A(n72), .Z(n35423) );
  XNOR U35878 ( .A(n35431), .B(n35645), .Z(n35424) );
  XNOR U35879 ( .A(n35430), .B(n35428), .Z(n35645) );
  AND U35880 ( .A(n35646), .B(n35647), .Z(n35428) );
  NANDN U35881 ( .A(n35648), .B(n35649), .Z(n35647) );
  OR U35882 ( .A(n35650), .B(n35651), .Z(n35649) );
  NAND U35883 ( .A(n35651), .B(n35650), .Z(n35646) );
  ANDN U35884 ( .B(B[161]), .A(n73), .Z(n35430) );
  XNOR U35885 ( .A(n35438), .B(n35652), .Z(n35431) );
  XNOR U35886 ( .A(n35437), .B(n35435), .Z(n35652) );
  AND U35887 ( .A(n35653), .B(n35654), .Z(n35435) );
  NANDN U35888 ( .A(n35655), .B(n35656), .Z(n35654) );
  NANDN U35889 ( .A(n35657), .B(n35658), .Z(n35656) );
  NANDN U35890 ( .A(n35658), .B(n35657), .Z(n35653) );
  ANDN U35891 ( .B(B[162]), .A(n74), .Z(n35437) );
  XNOR U35892 ( .A(n35445), .B(n35659), .Z(n35438) );
  XNOR U35893 ( .A(n35444), .B(n35442), .Z(n35659) );
  AND U35894 ( .A(n35660), .B(n35661), .Z(n35442) );
  NANDN U35895 ( .A(n35662), .B(n35663), .Z(n35661) );
  OR U35896 ( .A(n35664), .B(n35665), .Z(n35663) );
  NAND U35897 ( .A(n35665), .B(n35664), .Z(n35660) );
  ANDN U35898 ( .B(B[163]), .A(n75), .Z(n35444) );
  XNOR U35899 ( .A(n35452), .B(n35666), .Z(n35445) );
  XNOR U35900 ( .A(n35451), .B(n35449), .Z(n35666) );
  AND U35901 ( .A(n35667), .B(n35668), .Z(n35449) );
  NANDN U35902 ( .A(n35669), .B(n35670), .Z(n35668) );
  NANDN U35903 ( .A(n35671), .B(n35672), .Z(n35670) );
  NANDN U35904 ( .A(n35672), .B(n35671), .Z(n35667) );
  ANDN U35905 ( .B(B[164]), .A(n76), .Z(n35451) );
  XNOR U35906 ( .A(n35459), .B(n35673), .Z(n35452) );
  XNOR U35907 ( .A(n35458), .B(n35456), .Z(n35673) );
  AND U35908 ( .A(n35674), .B(n35675), .Z(n35456) );
  NANDN U35909 ( .A(n35676), .B(n35677), .Z(n35675) );
  OR U35910 ( .A(n35678), .B(n35679), .Z(n35677) );
  NAND U35911 ( .A(n35679), .B(n35678), .Z(n35674) );
  ANDN U35912 ( .B(B[165]), .A(n77), .Z(n35458) );
  XNOR U35913 ( .A(n35466), .B(n35680), .Z(n35459) );
  XNOR U35914 ( .A(n35465), .B(n35463), .Z(n35680) );
  AND U35915 ( .A(n35681), .B(n35682), .Z(n35463) );
  NANDN U35916 ( .A(n35683), .B(n35684), .Z(n35682) );
  NANDN U35917 ( .A(n35685), .B(n35686), .Z(n35684) );
  NANDN U35918 ( .A(n35686), .B(n35685), .Z(n35681) );
  ANDN U35919 ( .B(B[166]), .A(n78), .Z(n35465) );
  XNOR U35920 ( .A(n35473), .B(n35687), .Z(n35466) );
  XNOR U35921 ( .A(n35472), .B(n35470), .Z(n35687) );
  AND U35922 ( .A(n35688), .B(n35689), .Z(n35470) );
  NANDN U35923 ( .A(n35690), .B(n35691), .Z(n35689) );
  OR U35924 ( .A(n35692), .B(n35693), .Z(n35691) );
  NAND U35925 ( .A(n35693), .B(n35692), .Z(n35688) );
  ANDN U35926 ( .B(B[167]), .A(n79), .Z(n35472) );
  XNOR U35927 ( .A(n35480), .B(n35694), .Z(n35473) );
  XNOR U35928 ( .A(n35479), .B(n35477), .Z(n35694) );
  AND U35929 ( .A(n35695), .B(n35696), .Z(n35477) );
  NANDN U35930 ( .A(n35697), .B(n35698), .Z(n35696) );
  NANDN U35931 ( .A(n35699), .B(n35700), .Z(n35698) );
  NANDN U35932 ( .A(n35700), .B(n35699), .Z(n35695) );
  ANDN U35933 ( .B(B[168]), .A(n80), .Z(n35479) );
  XNOR U35934 ( .A(n35487), .B(n35701), .Z(n35480) );
  XNOR U35935 ( .A(n35486), .B(n35484), .Z(n35701) );
  AND U35936 ( .A(n35702), .B(n35703), .Z(n35484) );
  NANDN U35937 ( .A(n35704), .B(n35705), .Z(n35703) );
  OR U35938 ( .A(n35706), .B(n35707), .Z(n35705) );
  NAND U35939 ( .A(n35707), .B(n35706), .Z(n35702) );
  ANDN U35940 ( .B(B[169]), .A(n81), .Z(n35486) );
  XNOR U35941 ( .A(n35494), .B(n35708), .Z(n35487) );
  XNOR U35942 ( .A(n35493), .B(n35491), .Z(n35708) );
  AND U35943 ( .A(n35709), .B(n35710), .Z(n35491) );
  NANDN U35944 ( .A(n35711), .B(n35712), .Z(n35710) );
  NAND U35945 ( .A(n35713), .B(n35714), .Z(n35712) );
  ANDN U35946 ( .B(B[170]), .A(n82), .Z(n35493) );
  XOR U35947 ( .A(n35500), .B(n35715), .Z(n35494) );
  XNOR U35948 ( .A(n35498), .B(n35501), .Z(n35715) );
  NAND U35949 ( .A(A[2]), .B(B[171]), .Z(n35501) );
  NANDN U35950 ( .A(n35716), .B(n35717), .Z(n35498) );
  AND U35951 ( .A(A[0]), .B(B[172]), .Z(n35717) );
  XNOR U35952 ( .A(n35503), .B(n35718), .Z(n35500) );
  NAND U35953 ( .A(A[0]), .B(B[173]), .Z(n35718) );
  NAND U35954 ( .A(B[172]), .B(A[1]), .Z(n35503) );
  NAND U35955 ( .A(n35719), .B(n35720), .Z(n450) );
  NANDN U35956 ( .A(n35721), .B(n35722), .Z(n35720) );
  OR U35957 ( .A(n35723), .B(n35724), .Z(n35722) );
  NAND U35958 ( .A(n35724), .B(n35723), .Z(n35719) );
  XOR U35959 ( .A(n452), .B(n451), .Z(\A1[170] ) );
  XOR U35960 ( .A(n35724), .B(n35725), .Z(n451) );
  XNOR U35961 ( .A(n35723), .B(n35721), .Z(n35725) );
  AND U35962 ( .A(n35726), .B(n35727), .Z(n35721) );
  NANDN U35963 ( .A(n35728), .B(n35729), .Z(n35727) );
  NANDN U35964 ( .A(n35730), .B(n35731), .Z(n35729) );
  NANDN U35965 ( .A(n35731), .B(n35730), .Z(n35726) );
  ANDN U35966 ( .B(B[141]), .A(n54), .Z(n35723) );
  XNOR U35967 ( .A(n35518), .B(n35732), .Z(n35724) );
  XNOR U35968 ( .A(n35517), .B(n35515), .Z(n35732) );
  AND U35969 ( .A(n35733), .B(n35734), .Z(n35515) );
  NANDN U35970 ( .A(n35735), .B(n35736), .Z(n35734) );
  OR U35971 ( .A(n35737), .B(n35738), .Z(n35736) );
  NAND U35972 ( .A(n35738), .B(n35737), .Z(n35733) );
  ANDN U35973 ( .B(B[142]), .A(n55), .Z(n35517) );
  XNOR U35974 ( .A(n35525), .B(n35739), .Z(n35518) );
  XNOR U35975 ( .A(n35524), .B(n35522), .Z(n35739) );
  AND U35976 ( .A(n35740), .B(n35741), .Z(n35522) );
  NANDN U35977 ( .A(n35742), .B(n35743), .Z(n35741) );
  NANDN U35978 ( .A(n35744), .B(n35745), .Z(n35743) );
  NANDN U35979 ( .A(n35745), .B(n35744), .Z(n35740) );
  ANDN U35980 ( .B(B[143]), .A(n56), .Z(n35524) );
  XNOR U35981 ( .A(n35532), .B(n35746), .Z(n35525) );
  XNOR U35982 ( .A(n35531), .B(n35529), .Z(n35746) );
  AND U35983 ( .A(n35747), .B(n35748), .Z(n35529) );
  NANDN U35984 ( .A(n35749), .B(n35750), .Z(n35748) );
  OR U35985 ( .A(n35751), .B(n35752), .Z(n35750) );
  NAND U35986 ( .A(n35752), .B(n35751), .Z(n35747) );
  ANDN U35987 ( .B(B[144]), .A(n57), .Z(n35531) );
  XNOR U35988 ( .A(n35539), .B(n35753), .Z(n35532) );
  XNOR U35989 ( .A(n35538), .B(n35536), .Z(n35753) );
  AND U35990 ( .A(n35754), .B(n35755), .Z(n35536) );
  NANDN U35991 ( .A(n35756), .B(n35757), .Z(n35755) );
  NANDN U35992 ( .A(n35758), .B(n35759), .Z(n35757) );
  NANDN U35993 ( .A(n35759), .B(n35758), .Z(n35754) );
  ANDN U35994 ( .B(B[145]), .A(n58), .Z(n35538) );
  XNOR U35995 ( .A(n35546), .B(n35760), .Z(n35539) );
  XNOR U35996 ( .A(n35545), .B(n35543), .Z(n35760) );
  AND U35997 ( .A(n35761), .B(n35762), .Z(n35543) );
  NANDN U35998 ( .A(n35763), .B(n35764), .Z(n35762) );
  OR U35999 ( .A(n35765), .B(n35766), .Z(n35764) );
  NAND U36000 ( .A(n35766), .B(n35765), .Z(n35761) );
  ANDN U36001 ( .B(B[146]), .A(n59), .Z(n35545) );
  XNOR U36002 ( .A(n35553), .B(n35767), .Z(n35546) );
  XNOR U36003 ( .A(n35552), .B(n35550), .Z(n35767) );
  AND U36004 ( .A(n35768), .B(n35769), .Z(n35550) );
  NANDN U36005 ( .A(n35770), .B(n35771), .Z(n35769) );
  NANDN U36006 ( .A(n35772), .B(n35773), .Z(n35771) );
  NANDN U36007 ( .A(n35773), .B(n35772), .Z(n35768) );
  ANDN U36008 ( .B(B[147]), .A(n60), .Z(n35552) );
  XNOR U36009 ( .A(n35560), .B(n35774), .Z(n35553) );
  XNOR U36010 ( .A(n35559), .B(n35557), .Z(n35774) );
  AND U36011 ( .A(n35775), .B(n35776), .Z(n35557) );
  NANDN U36012 ( .A(n35777), .B(n35778), .Z(n35776) );
  OR U36013 ( .A(n35779), .B(n35780), .Z(n35778) );
  NAND U36014 ( .A(n35780), .B(n35779), .Z(n35775) );
  ANDN U36015 ( .B(B[148]), .A(n61), .Z(n35559) );
  XNOR U36016 ( .A(n35567), .B(n35781), .Z(n35560) );
  XNOR U36017 ( .A(n35566), .B(n35564), .Z(n35781) );
  AND U36018 ( .A(n35782), .B(n35783), .Z(n35564) );
  NANDN U36019 ( .A(n35784), .B(n35785), .Z(n35783) );
  NANDN U36020 ( .A(n35786), .B(n35787), .Z(n35785) );
  NANDN U36021 ( .A(n35787), .B(n35786), .Z(n35782) );
  ANDN U36022 ( .B(B[149]), .A(n62), .Z(n35566) );
  XNOR U36023 ( .A(n35574), .B(n35788), .Z(n35567) );
  XNOR U36024 ( .A(n35573), .B(n35571), .Z(n35788) );
  AND U36025 ( .A(n35789), .B(n35790), .Z(n35571) );
  NANDN U36026 ( .A(n35791), .B(n35792), .Z(n35790) );
  OR U36027 ( .A(n35793), .B(n35794), .Z(n35792) );
  NAND U36028 ( .A(n35794), .B(n35793), .Z(n35789) );
  ANDN U36029 ( .B(B[150]), .A(n63), .Z(n35573) );
  XNOR U36030 ( .A(n35581), .B(n35795), .Z(n35574) );
  XNOR U36031 ( .A(n35580), .B(n35578), .Z(n35795) );
  AND U36032 ( .A(n35796), .B(n35797), .Z(n35578) );
  NANDN U36033 ( .A(n35798), .B(n35799), .Z(n35797) );
  NANDN U36034 ( .A(n35800), .B(n35801), .Z(n35799) );
  NANDN U36035 ( .A(n35801), .B(n35800), .Z(n35796) );
  ANDN U36036 ( .B(B[151]), .A(n64), .Z(n35580) );
  XNOR U36037 ( .A(n35588), .B(n35802), .Z(n35581) );
  XNOR U36038 ( .A(n35587), .B(n35585), .Z(n35802) );
  AND U36039 ( .A(n35803), .B(n35804), .Z(n35585) );
  NANDN U36040 ( .A(n35805), .B(n35806), .Z(n35804) );
  OR U36041 ( .A(n35807), .B(n35808), .Z(n35806) );
  NAND U36042 ( .A(n35808), .B(n35807), .Z(n35803) );
  ANDN U36043 ( .B(B[152]), .A(n65), .Z(n35587) );
  XNOR U36044 ( .A(n35595), .B(n35809), .Z(n35588) );
  XNOR U36045 ( .A(n35594), .B(n35592), .Z(n35809) );
  AND U36046 ( .A(n35810), .B(n35811), .Z(n35592) );
  NANDN U36047 ( .A(n35812), .B(n35813), .Z(n35811) );
  NANDN U36048 ( .A(n35814), .B(n35815), .Z(n35813) );
  NANDN U36049 ( .A(n35815), .B(n35814), .Z(n35810) );
  ANDN U36050 ( .B(B[153]), .A(n66), .Z(n35594) );
  XNOR U36051 ( .A(n35602), .B(n35816), .Z(n35595) );
  XNOR U36052 ( .A(n35601), .B(n35599), .Z(n35816) );
  AND U36053 ( .A(n35817), .B(n35818), .Z(n35599) );
  NANDN U36054 ( .A(n35819), .B(n35820), .Z(n35818) );
  OR U36055 ( .A(n35821), .B(n35822), .Z(n35820) );
  NAND U36056 ( .A(n35822), .B(n35821), .Z(n35817) );
  ANDN U36057 ( .B(B[154]), .A(n67), .Z(n35601) );
  XNOR U36058 ( .A(n35609), .B(n35823), .Z(n35602) );
  XNOR U36059 ( .A(n35608), .B(n35606), .Z(n35823) );
  AND U36060 ( .A(n35824), .B(n35825), .Z(n35606) );
  NANDN U36061 ( .A(n35826), .B(n35827), .Z(n35825) );
  NANDN U36062 ( .A(n35828), .B(n35829), .Z(n35827) );
  NANDN U36063 ( .A(n35829), .B(n35828), .Z(n35824) );
  ANDN U36064 ( .B(B[155]), .A(n68), .Z(n35608) );
  XNOR U36065 ( .A(n35616), .B(n35830), .Z(n35609) );
  XNOR U36066 ( .A(n35615), .B(n35613), .Z(n35830) );
  AND U36067 ( .A(n35831), .B(n35832), .Z(n35613) );
  NANDN U36068 ( .A(n35833), .B(n35834), .Z(n35832) );
  OR U36069 ( .A(n35835), .B(n35836), .Z(n35834) );
  NAND U36070 ( .A(n35836), .B(n35835), .Z(n35831) );
  ANDN U36071 ( .B(B[156]), .A(n69), .Z(n35615) );
  XNOR U36072 ( .A(n35623), .B(n35837), .Z(n35616) );
  XNOR U36073 ( .A(n35622), .B(n35620), .Z(n35837) );
  AND U36074 ( .A(n35838), .B(n35839), .Z(n35620) );
  NANDN U36075 ( .A(n35840), .B(n35841), .Z(n35839) );
  NANDN U36076 ( .A(n35842), .B(n35843), .Z(n35841) );
  NANDN U36077 ( .A(n35843), .B(n35842), .Z(n35838) );
  ANDN U36078 ( .B(B[157]), .A(n70), .Z(n35622) );
  XNOR U36079 ( .A(n35630), .B(n35844), .Z(n35623) );
  XNOR U36080 ( .A(n35629), .B(n35627), .Z(n35844) );
  AND U36081 ( .A(n35845), .B(n35846), .Z(n35627) );
  NANDN U36082 ( .A(n35847), .B(n35848), .Z(n35846) );
  OR U36083 ( .A(n35849), .B(n35850), .Z(n35848) );
  NAND U36084 ( .A(n35850), .B(n35849), .Z(n35845) );
  ANDN U36085 ( .B(B[158]), .A(n71), .Z(n35629) );
  XNOR U36086 ( .A(n35637), .B(n35851), .Z(n35630) );
  XNOR U36087 ( .A(n35636), .B(n35634), .Z(n35851) );
  AND U36088 ( .A(n35852), .B(n35853), .Z(n35634) );
  NANDN U36089 ( .A(n35854), .B(n35855), .Z(n35853) );
  NANDN U36090 ( .A(n35856), .B(n35857), .Z(n35855) );
  NANDN U36091 ( .A(n35857), .B(n35856), .Z(n35852) );
  ANDN U36092 ( .B(B[159]), .A(n72), .Z(n35636) );
  XNOR U36093 ( .A(n35644), .B(n35858), .Z(n35637) );
  XNOR U36094 ( .A(n35643), .B(n35641), .Z(n35858) );
  AND U36095 ( .A(n35859), .B(n35860), .Z(n35641) );
  NANDN U36096 ( .A(n35861), .B(n35862), .Z(n35860) );
  OR U36097 ( .A(n35863), .B(n35864), .Z(n35862) );
  NAND U36098 ( .A(n35864), .B(n35863), .Z(n35859) );
  ANDN U36099 ( .B(B[160]), .A(n73), .Z(n35643) );
  XNOR U36100 ( .A(n35651), .B(n35865), .Z(n35644) );
  XNOR U36101 ( .A(n35650), .B(n35648), .Z(n35865) );
  AND U36102 ( .A(n35866), .B(n35867), .Z(n35648) );
  NANDN U36103 ( .A(n35868), .B(n35869), .Z(n35867) );
  NANDN U36104 ( .A(n35870), .B(n35871), .Z(n35869) );
  NANDN U36105 ( .A(n35871), .B(n35870), .Z(n35866) );
  ANDN U36106 ( .B(B[161]), .A(n74), .Z(n35650) );
  XNOR U36107 ( .A(n35658), .B(n35872), .Z(n35651) );
  XNOR U36108 ( .A(n35657), .B(n35655), .Z(n35872) );
  AND U36109 ( .A(n35873), .B(n35874), .Z(n35655) );
  NANDN U36110 ( .A(n35875), .B(n35876), .Z(n35874) );
  OR U36111 ( .A(n35877), .B(n35878), .Z(n35876) );
  NAND U36112 ( .A(n35878), .B(n35877), .Z(n35873) );
  ANDN U36113 ( .B(B[162]), .A(n75), .Z(n35657) );
  XNOR U36114 ( .A(n35665), .B(n35879), .Z(n35658) );
  XNOR U36115 ( .A(n35664), .B(n35662), .Z(n35879) );
  AND U36116 ( .A(n35880), .B(n35881), .Z(n35662) );
  NANDN U36117 ( .A(n35882), .B(n35883), .Z(n35881) );
  NANDN U36118 ( .A(n35884), .B(n35885), .Z(n35883) );
  NANDN U36119 ( .A(n35885), .B(n35884), .Z(n35880) );
  ANDN U36120 ( .B(B[163]), .A(n76), .Z(n35664) );
  XNOR U36121 ( .A(n35672), .B(n35886), .Z(n35665) );
  XNOR U36122 ( .A(n35671), .B(n35669), .Z(n35886) );
  AND U36123 ( .A(n35887), .B(n35888), .Z(n35669) );
  NANDN U36124 ( .A(n35889), .B(n35890), .Z(n35888) );
  OR U36125 ( .A(n35891), .B(n35892), .Z(n35890) );
  NAND U36126 ( .A(n35892), .B(n35891), .Z(n35887) );
  ANDN U36127 ( .B(B[164]), .A(n77), .Z(n35671) );
  XNOR U36128 ( .A(n35679), .B(n35893), .Z(n35672) );
  XNOR U36129 ( .A(n35678), .B(n35676), .Z(n35893) );
  AND U36130 ( .A(n35894), .B(n35895), .Z(n35676) );
  NANDN U36131 ( .A(n35896), .B(n35897), .Z(n35895) );
  NANDN U36132 ( .A(n35898), .B(n35899), .Z(n35897) );
  NANDN U36133 ( .A(n35899), .B(n35898), .Z(n35894) );
  ANDN U36134 ( .B(B[165]), .A(n78), .Z(n35678) );
  XNOR U36135 ( .A(n35686), .B(n35900), .Z(n35679) );
  XNOR U36136 ( .A(n35685), .B(n35683), .Z(n35900) );
  AND U36137 ( .A(n35901), .B(n35902), .Z(n35683) );
  NANDN U36138 ( .A(n35903), .B(n35904), .Z(n35902) );
  OR U36139 ( .A(n35905), .B(n35906), .Z(n35904) );
  NAND U36140 ( .A(n35906), .B(n35905), .Z(n35901) );
  ANDN U36141 ( .B(B[166]), .A(n79), .Z(n35685) );
  XNOR U36142 ( .A(n35693), .B(n35907), .Z(n35686) );
  XNOR U36143 ( .A(n35692), .B(n35690), .Z(n35907) );
  AND U36144 ( .A(n35908), .B(n35909), .Z(n35690) );
  NANDN U36145 ( .A(n35910), .B(n35911), .Z(n35909) );
  NANDN U36146 ( .A(n35912), .B(n35913), .Z(n35911) );
  NANDN U36147 ( .A(n35913), .B(n35912), .Z(n35908) );
  ANDN U36148 ( .B(B[167]), .A(n80), .Z(n35692) );
  XNOR U36149 ( .A(n35700), .B(n35914), .Z(n35693) );
  XNOR U36150 ( .A(n35699), .B(n35697), .Z(n35914) );
  AND U36151 ( .A(n35915), .B(n35916), .Z(n35697) );
  NANDN U36152 ( .A(n35917), .B(n35918), .Z(n35916) );
  OR U36153 ( .A(n35919), .B(n35920), .Z(n35918) );
  NAND U36154 ( .A(n35920), .B(n35919), .Z(n35915) );
  ANDN U36155 ( .B(B[168]), .A(n81), .Z(n35699) );
  XNOR U36156 ( .A(n35707), .B(n35921), .Z(n35700) );
  XNOR U36157 ( .A(n35706), .B(n35704), .Z(n35921) );
  AND U36158 ( .A(n35922), .B(n35923), .Z(n35704) );
  NANDN U36159 ( .A(n35924), .B(n35925), .Z(n35923) );
  NAND U36160 ( .A(n35926), .B(n35927), .Z(n35925) );
  ANDN U36161 ( .B(B[169]), .A(n82), .Z(n35706) );
  XOR U36162 ( .A(n35713), .B(n35928), .Z(n35707) );
  XNOR U36163 ( .A(n35711), .B(n35714), .Z(n35928) );
  NAND U36164 ( .A(A[2]), .B(B[170]), .Z(n35714) );
  NANDN U36165 ( .A(n35929), .B(n35930), .Z(n35711) );
  AND U36166 ( .A(A[0]), .B(B[171]), .Z(n35930) );
  XNOR U36167 ( .A(n35716), .B(n35931), .Z(n35713) );
  NAND U36168 ( .A(A[0]), .B(B[172]), .Z(n35931) );
  NAND U36169 ( .A(B[171]), .B(A[1]), .Z(n35716) );
  NAND U36170 ( .A(n35932), .B(n35933), .Z(n452) );
  NANDN U36171 ( .A(n35934), .B(n35935), .Z(n35933) );
  OR U36172 ( .A(n35936), .B(n35937), .Z(n35935) );
  NAND U36173 ( .A(n35937), .B(n35936), .Z(n35932) );
  XOR U36174 ( .A(n33691), .B(n35938), .Z(\A1[16] ) );
  XNOR U36175 ( .A(n33690), .B(n33689), .Z(n35938) );
  NAND U36176 ( .A(n35939), .B(n35940), .Z(n33689) );
  NANDN U36177 ( .A(n35941), .B(n35942), .Z(n35940) );
  OR U36178 ( .A(n35943), .B(n35944), .Z(n35942) );
  NAND U36179 ( .A(n35944), .B(n35943), .Z(n35939) );
  ANDN U36180 ( .B(B[0]), .A(n67), .Z(n33690) );
  XNOR U36181 ( .A(n33698), .B(n35945), .Z(n33691) );
  XNOR U36182 ( .A(n33697), .B(n33695), .Z(n35945) );
  AND U36183 ( .A(n35946), .B(n35947), .Z(n33695) );
  NANDN U36184 ( .A(n35948), .B(n35949), .Z(n35947) );
  NANDN U36185 ( .A(n35950), .B(n35951), .Z(n35949) );
  NANDN U36186 ( .A(n35951), .B(n35950), .Z(n35946) );
  ANDN U36187 ( .B(B[1]), .A(n68), .Z(n33697) );
  XNOR U36188 ( .A(n33705), .B(n35952), .Z(n33698) );
  XNOR U36189 ( .A(n33704), .B(n33702), .Z(n35952) );
  AND U36190 ( .A(n35953), .B(n35954), .Z(n33702) );
  NANDN U36191 ( .A(n35955), .B(n35956), .Z(n35954) );
  OR U36192 ( .A(n35957), .B(n35958), .Z(n35956) );
  NAND U36193 ( .A(n35958), .B(n35957), .Z(n35953) );
  ANDN U36194 ( .B(B[2]), .A(n69), .Z(n33704) );
  XNOR U36195 ( .A(n33712), .B(n35959), .Z(n33705) );
  XNOR U36196 ( .A(n33711), .B(n33709), .Z(n35959) );
  AND U36197 ( .A(n35960), .B(n35961), .Z(n33709) );
  NANDN U36198 ( .A(n35962), .B(n35963), .Z(n35961) );
  NANDN U36199 ( .A(n35964), .B(n35965), .Z(n35963) );
  NANDN U36200 ( .A(n35965), .B(n35964), .Z(n35960) );
  ANDN U36201 ( .B(B[3]), .A(n70), .Z(n33711) );
  XNOR U36202 ( .A(n33719), .B(n35966), .Z(n33712) );
  XNOR U36203 ( .A(n33718), .B(n33716), .Z(n35966) );
  AND U36204 ( .A(n35967), .B(n35968), .Z(n33716) );
  NANDN U36205 ( .A(n35969), .B(n35970), .Z(n35968) );
  OR U36206 ( .A(n35971), .B(n35972), .Z(n35970) );
  NAND U36207 ( .A(n35972), .B(n35971), .Z(n35967) );
  ANDN U36208 ( .B(B[4]), .A(n71), .Z(n33718) );
  XNOR U36209 ( .A(n33726), .B(n35973), .Z(n33719) );
  XNOR U36210 ( .A(n33725), .B(n33723), .Z(n35973) );
  AND U36211 ( .A(n35974), .B(n35975), .Z(n33723) );
  NANDN U36212 ( .A(n35976), .B(n35977), .Z(n35975) );
  NANDN U36213 ( .A(n35978), .B(n35979), .Z(n35977) );
  NANDN U36214 ( .A(n35979), .B(n35978), .Z(n35974) );
  ANDN U36215 ( .B(B[5]), .A(n72), .Z(n33725) );
  XNOR U36216 ( .A(n33733), .B(n35980), .Z(n33726) );
  XNOR U36217 ( .A(n33732), .B(n33730), .Z(n35980) );
  AND U36218 ( .A(n35981), .B(n35982), .Z(n33730) );
  NANDN U36219 ( .A(n35983), .B(n35984), .Z(n35982) );
  OR U36220 ( .A(n35985), .B(n35986), .Z(n35984) );
  NAND U36221 ( .A(n35986), .B(n35985), .Z(n35981) );
  ANDN U36222 ( .B(B[6]), .A(n73), .Z(n33732) );
  XNOR U36223 ( .A(n33740), .B(n35987), .Z(n33733) );
  XNOR U36224 ( .A(n33739), .B(n33737), .Z(n35987) );
  AND U36225 ( .A(n35988), .B(n35989), .Z(n33737) );
  NANDN U36226 ( .A(n35990), .B(n35991), .Z(n35989) );
  NANDN U36227 ( .A(n35992), .B(n35993), .Z(n35991) );
  NANDN U36228 ( .A(n35993), .B(n35992), .Z(n35988) );
  ANDN U36229 ( .B(B[7]), .A(n74), .Z(n33739) );
  XNOR U36230 ( .A(n33747), .B(n35994), .Z(n33740) );
  XNOR U36231 ( .A(n33746), .B(n33744), .Z(n35994) );
  AND U36232 ( .A(n35995), .B(n35996), .Z(n33744) );
  NANDN U36233 ( .A(n35997), .B(n35998), .Z(n35996) );
  OR U36234 ( .A(n35999), .B(n36000), .Z(n35998) );
  NAND U36235 ( .A(n36000), .B(n35999), .Z(n35995) );
  ANDN U36236 ( .B(B[8]), .A(n75), .Z(n33746) );
  XNOR U36237 ( .A(n33754), .B(n36001), .Z(n33747) );
  XNOR U36238 ( .A(n33753), .B(n33751), .Z(n36001) );
  AND U36239 ( .A(n36002), .B(n36003), .Z(n33751) );
  NANDN U36240 ( .A(n36004), .B(n36005), .Z(n36003) );
  NANDN U36241 ( .A(n36006), .B(n36007), .Z(n36005) );
  NANDN U36242 ( .A(n36007), .B(n36006), .Z(n36002) );
  ANDN U36243 ( .B(B[9]), .A(n76), .Z(n33753) );
  XNOR U36244 ( .A(n33761), .B(n36008), .Z(n33754) );
  XNOR U36245 ( .A(n33760), .B(n33758), .Z(n36008) );
  AND U36246 ( .A(n36009), .B(n36010), .Z(n33758) );
  NANDN U36247 ( .A(n36011), .B(n36012), .Z(n36010) );
  OR U36248 ( .A(n36013), .B(n36014), .Z(n36012) );
  NAND U36249 ( .A(n36014), .B(n36013), .Z(n36009) );
  ANDN U36250 ( .B(B[10]), .A(n77), .Z(n33760) );
  XNOR U36251 ( .A(n33768), .B(n36015), .Z(n33761) );
  XNOR U36252 ( .A(n33767), .B(n33765), .Z(n36015) );
  AND U36253 ( .A(n36016), .B(n36017), .Z(n33765) );
  NANDN U36254 ( .A(n36018), .B(n36019), .Z(n36017) );
  NANDN U36255 ( .A(n36020), .B(n36021), .Z(n36019) );
  NANDN U36256 ( .A(n36021), .B(n36020), .Z(n36016) );
  ANDN U36257 ( .B(B[11]), .A(n78), .Z(n33767) );
  XNOR U36258 ( .A(n33775), .B(n36022), .Z(n33768) );
  XNOR U36259 ( .A(n33774), .B(n33772), .Z(n36022) );
  AND U36260 ( .A(n36023), .B(n36024), .Z(n33772) );
  NANDN U36261 ( .A(n36025), .B(n36026), .Z(n36024) );
  OR U36262 ( .A(n36027), .B(n36028), .Z(n36026) );
  NAND U36263 ( .A(n36028), .B(n36027), .Z(n36023) );
  ANDN U36264 ( .B(B[12]), .A(n79), .Z(n33774) );
  XNOR U36265 ( .A(n33782), .B(n36029), .Z(n33775) );
  XNOR U36266 ( .A(n33781), .B(n33779), .Z(n36029) );
  AND U36267 ( .A(n36030), .B(n36031), .Z(n33779) );
  NANDN U36268 ( .A(n36032), .B(n36033), .Z(n36031) );
  NANDN U36269 ( .A(n36034), .B(n36035), .Z(n36033) );
  NANDN U36270 ( .A(n36035), .B(n36034), .Z(n36030) );
  ANDN U36271 ( .B(B[13]), .A(n80), .Z(n33781) );
  XNOR U36272 ( .A(n33789), .B(n36036), .Z(n33782) );
  XNOR U36273 ( .A(n33788), .B(n33786), .Z(n36036) );
  AND U36274 ( .A(n36037), .B(n36038), .Z(n33786) );
  NANDN U36275 ( .A(n36039), .B(n36040), .Z(n36038) );
  OR U36276 ( .A(n36041), .B(n36042), .Z(n36040) );
  NAND U36277 ( .A(n36042), .B(n36041), .Z(n36037) );
  ANDN U36278 ( .B(B[14]), .A(n81), .Z(n33788) );
  XNOR U36279 ( .A(n33796), .B(n36043), .Z(n33789) );
  XNOR U36280 ( .A(n33795), .B(n33793), .Z(n36043) );
  AND U36281 ( .A(n36044), .B(n36045), .Z(n33793) );
  NANDN U36282 ( .A(n36046), .B(n36047), .Z(n36045) );
  NAND U36283 ( .A(n36048), .B(n36049), .Z(n36047) );
  ANDN U36284 ( .B(B[15]), .A(n82), .Z(n33795) );
  XOR U36285 ( .A(n33802), .B(n36050), .Z(n33796) );
  XNOR U36286 ( .A(n33800), .B(n33803), .Z(n36050) );
  NAND U36287 ( .A(A[2]), .B(B[16]), .Z(n33803) );
  NANDN U36288 ( .A(n36051), .B(n36052), .Z(n33800) );
  AND U36289 ( .A(A[0]), .B(B[17]), .Z(n36052) );
  XNOR U36290 ( .A(n33805), .B(n36053), .Z(n33802) );
  NAND U36291 ( .A(A[0]), .B(B[18]), .Z(n36053) );
  NAND U36292 ( .A(B[17]), .B(A[1]), .Z(n33805) );
  XOR U36293 ( .A(n454), .B(n453), .Z(\A1[169] ) );
  XOR U36294 ( .A(n35937), .B(n36054), .Z(n453) );
  XNOR U36295 ( .A(n35936), .B(n35934), .Z(n36054) );
  AND U36296 ( .A(n36055), .B(n36056), .Z(n35934) );
  NANDN U36297 ( .A(n36057), .B(n36058), .Z(n36056) );
  NANDN U36298 ( .A(n36059), .B(n36060), .Z(n36058) );
  NANDN U36299 ( .A(n36060), .B(n36059), .Z(n36055) );
  ANDN U36300 ( .B(B[140]), .A(n54), .Z(n35936) );
  XNOR U36301 ( .A(n35731), .B(n36061), .Z(n35937) );
  XNOR U36302 ( .A(n35730), .B(n35728), .Z(n36061) );
  AND U36303 ( .A(n36062), .B(n36063), .Z(n35728) );
  NANDN U36304 ( .A(n36064), .B(n36065), .Z(n36063) );
  OR U36305 ( .A(n36066), .B(n36067), .Z(n36065) );
  NAND U36306 ( .A(n36067), .B(n36066), .Z(n36062) );
  ANDN U36307 ( .B(B[141]), .A(n55), .Z(n35730) );
  XNOR U36308 ( .A(n35738), .B(n36068), .Z(n35731) );
  XNOR U36309 ( .A(n35737), .B(n35735), .Z(n36068) );
  AND U36310 ( .A(n36069), .B(n36070), .Z(n35735) );
  NANDN U36311 ( .A(n36071), .B(n36072), .Z(n36070) );
  NANDN U36312 ( .A(n36073), .B(n36074), .Z(n36072) );
  NANDN U36313 ( .A(n36074), .B(n36073), .Z(n36069) );
  ANDN U36314 ( .B(B[142]), .A(n56), .Z(n35737) );
  XNOR U36315 ( .A(n35745), .B(n36075), .Z(n35738) );
  XNOR U36316 ( .A(n35744), .B(n35742), .Z(n36075) );
  AND U36317 ( .A(n36076), .B(n36077), .Z(n35742) );
  NANDN U36318 ( .A(n36078), .B(n36079), .Z(n36077) );
  OR U36319 ( .A(n36080), .B(n36081), .Z(n36079) );
  NAND U36320 ( .A(n36081), .B(n36080), .Z(n36076) );
  ANDN U36321 ( .B(B[143]), .A(n57), .Z(n35744) );
  XNOR U36322 ( .A(n35752), .B(n36082), .Z(n35745) );
  XNOR U36323 ( .A(n35751), .B(n35749), .Z(n36082) );
  AND U36324 ( .A(n36083), .B(n36084), .Z(n35749) );
  NANDN U36325 ( .A(n36085), .B(n36086), .Z(n36084) );
  NANDN U36326 ( .A(n36087), .B(n36088), .Z(n36086) );
  NANDN U36327 ( .A(n36088), .B(n36087), .Z(n36083) );
  ANDN U36328 ( .B(B[144]), .A(n58), .Z(n35751) );
  XNOR U36329 ( .A(n35759), .B(n36089), .Z(n35752) );
  XNOR U36330 ( .A(n35758), .B(n35756), .Z(n36089) );
  AND U36331 ( .A(n36090), .B(n36091), .Z(n35756) );
  NANDN U36332 ( .A(n36092), .B(n36093), .Z(n36091) );
  OR U36333 ( .A(n36094), .B(n36095), .Z(n36093) );
  NAND U36334 ( .A(n36095), .B(n36094), .Z(n36090) );
  ANDN U36335 ( .B(B[145]), .A(n59), .Z(n35758) );
  XNOR U36336 ( .A(n35766), .B(n36096), .Z(n35759) );
  XNOR U36337 ( .A(n35765), .B(n35763), .Z(n36096) );
  AND U36338 ( .A(n36097), .B(n36098), .Z(n35763) );
  NANDN U36339 ( .A(n36099), .B(n36100), .Z(n36098) );
  NANDN U36340 ( .A(n36101), .B(n36102), .Z(n36100) );
  NANDN U36341 ( .A(n36102), .B(n36101), .Z(n36097) );
  ANDN U36342 ( .B(B[146]), .A(n60), .Z(n35765) );
  XNOR U36343 ( .A(n35773), .B(n36103), .Z(n35766) );
  XNOR U36344 ( .A(n35772), .B(n35770), .Z(n36103) );
  AND U36345 ( .A(n36104), .B(n36105), .Z(n35770) );
  NANDN U36346 ( .A(n36106), .B(n36107), .Z(n36105) );
  OR U36347 ( .A(n36108), .B(n36109), .Z(n36107) );
  NAND U36348 ( .A(n36109), .B(n36108), .Z(n36104) );
  ANDN U36349 ( .B(B[147]), .A(n61), .Z(n35772) );
  XNOR U36350 ( .A(n35780), .B(n36110), .Z(n35773) );
  XNOR U36351 ( .A(n35779), .B(n35777), .Z(n36110) );
  AND U36352 ( .A(n36111), .B(n36112), .Z(n35777) );
  NANDN U36353 ( .A(n36113), .B(n36114), .Z(n36112) );
  NANDN U36354 ( .A(n36115), .B(n36116), .Z(n36114) );
  NANDN U36355 ( .A(n36116), .B(n36115), .Z(n36111) );
  ANDN U36356 ( .B(B[148]), .A(n62), .Z(n35779) );
  XNOR U36357 ( .A(n35787), .B(n36117), .Z(n35780) );
  XNOR U36358 ( .A(n35786), .B(n35784), .Z(n36117) );
  AND U36359 ( .A(n36118), .B(n36119), .Z(n35784) );
  NANDN U36360 ( .A(n36120), .B(n36121), .Z(n36119) );
  OR U36361 ( .A(n36122), .B(n36123), .Z(n36121) );
  NAND U36362 ( .A(n36123), .B(n36122), .Z(n36118) );
  ANDN U36363 ( .B(B[149]), .A(n63), .Z(n35786) );
  XNOR U36364 ( .A(n35794), .B(n36124), .Z(n35787) );
  XNOR U36365 ( .A(n35793), .B(n35791), .Z(n36124) );
  AND U36366 ( .A(n36125), .B(n36126), .Z(n35791) );
  NANDN U36367 ( .A(n36127), .B(n36128), .Z(n36126) );
  NANDN U36368 ( .A(n36129), .B(n36130), .Z(n36128) );
  NANDN U36369 ( .A(n36130), .B(n36129), .Z(n36125) );
  ANDN U36370 ( .B(B[150]), .A(n64), .Z(n35793) );
  XNOR U36371 ( .A(n35801), .B(n36131), .Z(n35794) );
  XNOR U36372 ( .A(n35800), .B(n35798), .Z(n36131) );
  AND U36373 ( .A(n36132), .B(n36133), .Z(n35798) );
  NANDN U36374 ( .A(n36134), .B(n36135), .Z(n36133) );
  OR U36375 ( .A(n36136), .B(n36137), .Z(n36135) );
  NAND U36376 ( .A(n36137), .B(n36136), .Z(n36132) );
  ANDN U36377 ( .B(B[151]), .A(n65), .Z(n35800) );
  XNOR U36378 ( .A(n35808), .B(n36138), .Z(n35801) );
  XNOR U36379 ( .A(n35807), .B(n35805), .Z(n36138) );
  AND U36380 ( .A(n36139), .B(n36140), .Z(n35805) );
  NANDN U36381 ( .A(n36141), .B(n36142), .Z(n36140) );
  NANDN U36382 ( .A(n36143), .B(n36144), .Z(n36142) );
  NANDN U36383 ( .A(n36144), .B(n36143), .Z(n36139) );
  ANDN U36384 ( .B(B[152]), .A(n66), .Z(n35807) );
  XNOR U36385 ( .A(n35815), .B(n36145), .Z(n35808) );
  XNOR U36386 ( .A(n35814), .B(n35812), .Z(n36145) );
  AND U36387 ( .A(n36146), .B(n36147), .Z(n35812) );
  NANDN U36388 ( .A(n36148), .B(n36149), .Z(n36147) );
  OR U36389 ( .A(n36150), .B(n36151), .Z(n36149) );
  NAND U36390 ( .A(n36151), .B(n36150), .Z(n36146) );
  ANDN U36391 ( .B(B[153]), .A(n67), .Z(n35814) );
  XNOR U36392 ( .A(n35822), .B(n36152), .Z(n35815) );
  XNOR U36393 ( .A(n35821), .B(n35819), .Z(n36152) );
  AND U36394 ( .A(n36153), .B(n36154), .Z(n35819) );
  NANDN U36395 ( .A(n36155), .B(n36156), .Z(n36154) );
  NANDN U36396 ( .A(n36157), .B(n36158), .Z(n36156) );
  NANDN U36397 ( .A(n36158), .B(n36157), .Z(n36153) );
  ANDN U36398 ( .B(B[154]), .A(n68), .Z(n35821) );
  XNOR U36399 ( .A(n35829), .B(n36159), .Z(n35822) );
  XNOR U36400 ( .A(n35828), .B(n35826), .Z(n36159) );
  AND U36401 ( .A(n36160), .B(n36161), .Z(n35826) );
  NANDN U36402 ( .A(n36162), .B(n36163), .Z(n36161) );
  OR U36403 ( .A(n36164), .B(n36165), .Z(n36163) );
  NAND U36404 ( .A(n36165), .B(n36164), .Z(n36160) );
  ANDN U36405 ( .B(B[155]), .A(n69), .Z(n35828) );
  XNOR U36406 ( .A(n35836), .B(n36166), .Z(n35829) );
  XNOR U36407 ( .A(n35835), .B(n35833), .Z(n36166) );
  AND U36408 ( .A(n36167), .B(n36168), .Z(n35833) );
  NANDN U36409 ( .A(n36169), .B(n36170), .Z(n36168) );
  NANDN U36410 ( .A(n36171), .B(n36172), .Z(n36170) );
  NANDN U36411 ( .A(n36172), .B(n36171), .Z(n36167) );
  ANDN U36412 ( .B(B[156]), .A(n70), .Z(n35835) );
  XNOR U36413 ( .A(n35843), .B(n36173), .Z(n35836) );
  XNOR U36414 ( .A(n35842), .B(n35840), .Z(n36173) );
  AND U36415 ( .A(n36174), .B(n36175), .Z(n35840) );
  NANDN U36416 ( .A(n36176), .B(n36177), .Z(n36175) );
  OR U36417 ( .A(n36178), .B(n36179), .Z(n36177) );
  NAND U36418 ( .A(n36179), .B(n36178), .Z(n36174) );
  ANDN U36419 ( .B(B[157]), .A(n71), .Z(n35842) );
  XNOR U36420 ( .A(n35850), .B(n36180), .Z(n35843) );
  XNOR U36421 ( .A(n35849), .B(n35847), .Z(n36180) );
  AND U36422 ( .A(n36181), .B(n36182), .Z(n35847) );
  NANDN U36423 ( .A(n36183), .B(n36184), .Z(n36182) );
  NANDN U36424 ( .A(n36185), .B(n36186), .Z(n36184) );
  NANDN U36425 ( .A(n36186), .B(n36185), .Z(n36181) );
  ANDN U36426 ( .B(B[158]), .A(n72), .Z(n35849) );
  XNOR U36427 ( .A(n35857), .B(n36187), .Z(n35850) );
  XNOR U36428 ( .A(n35856), .B(n35854), .Z(n36187) );
  AND U36429 ( .A(n36188), .B(n36189), .Z(n35854) );
  NANDN U36430 ( .A(n36190), .B(n36191), .Z(n36189) );
  OR U36431 ( .A(n36192), .B(n36193), .Z(n36191) );
  NAND U36432 ( .A(n36193), .B(n36192), .Z(n36188) );
  ANDN U36433 ( .B(B[159]), .A(n73), .Z(n35856) );
  XNOR U36434 ( .A(n35864), .B(n36194), .Z(n35857) );
  XNOR U36435 ( .A(n35863), .B(n35861), .Z(n36194) );
  AND U36436 ( .A(n36195), .B(n36196), .Z(n35861) );
  NANDN U36437 ( .A(n36197), .B(n36198), .Z(n36196) );
  NANDN U36438 ( .A(n36199), .B(n36200), .Z(n36198) );
  NANDN U36439 ( .A(n36200), .B(n36199), .Z(n36195) );
  ANDN U36440 ( .B(B[160]), .A(n74), .Z(n35863) );
  XNOR U36441 ( .A(n35871), .B(n36201), .Z(n35864) );
  XNOR U36442 ( .A(n35870), .B(n35868), .Z(n36201) );
  AND U36443 ( .A(n36202), .B(n36203), .Z(n35868) );
  NANDN U36444 ( .A(n36204), .B(n36205), .Z(n36203) );
  OR U36445 ( .A(n36206), .B(n36207), .Z(n36205) );
  NAND U36446 ( .A(n36207), .B(n36206), .Z(n36202) );
  ANDN U36447 ( .B(B[161]), .A(n75), .Z(n35870) );
  XNOR U36448 ( .A(n35878), .B(n36208), .Z(n35871) );
  XNOR U36449 ( .A(n35877), .B(n35875), .Z(n36208) );
  AND U36450 ( .A(n36209), .B(n36210), .Z(n35875) );
  NANDN U36451 ( .A(n36211), .B(n36212), .Z(n36210) );
  NANDN U36452 ( .A(n36213), .B(n36214), .Z(n36212) );
  NANDN U36453 ( .A(n36214), .B(n36213), .Z(n36209) );
  ANDN U36454 ( .B(B[162]), .A(n76), .Z(n35877) );
  XNOR U36455 ( .A(n35885), .B(n36215), .Z(n35878) );
  XNOR U36456 ( .A(n35884), .B(n35882), .Z(n36215) );
  AND U36457 ( .A(n36216), .B(n36217), .Z(n35882) );
  NANDN U36458 ( .A(n36218), .B(n36219), .Z(n36217) );
  OR U36459 ( .A(n36220), .B(n36221), .Z(n36219) );
  NAND U36460 ( .A(n36221), .B(n36220), .Z(n36216) );
  ANDN U36461 ( .B(B[163]), .A(n77), .Z(n35884) );
  XNOR U36462 ( .A(n35892), .B(n36222), .Z(n35885) );
  XNOR U36463 ( .A(n35891), .B(n35889), .Z(n36222) );
  AND U36464 ( .A(n36223), .B(n36224), .Z(n35889) );
  NANDN U36465 ( .A(n36225), .B(n36226), .Z(n36224) );
  NANDN U36466 ( .A(n36227), .B(n36228), .Z(n36226) );
  NANDN U36467 ( .A(n36228), .B(n36227), .Z(n36223) );
  ANDN U36468 ( .B(B[164]), .A(n78), .Z(n35891) );
  XNOR U36469 ( .A(n35899), .B(n36229), .Z(n35892) );
  XNOR U36470 ( .A(n35898), .B(n35896), .Z(n36229) );
  AND U36471 ( .A(n36230), .B(n36231), .Z(n35896) );
  NANDN U36472 ( .A(n36232), .B(n36233), .Z(n36231) );
  OR U36473 ( .A(n36234), .B(n36235), .Z(n36233) );
  NAND U36474 ( .A(n36235), .B(n36234), .Z(n36230) );
  ANDN U36475 ( .B(B[165]), .A(n79), .Z(n35898) );
  XNOR U36476 ( .A(n35906), .B(n36236), .Z(n35899) );
  XNOR U36477 ( .A(n35905), .B(n35903), .Z(n36236) );
  AND U36478 ( .A(n36237), .B(n36238), .Z(n35903) );
  NANDN U36479 ( .A(n36239), .B(n36240), .Z(n36238) );
  NANDN U36480 ( .A(n36241), .B(n36242), .Z(n36240) );
  NANDN U36481 ( .A(n36242), .B(n36241), .Z(n36237) );
  ANDN U36482 ( .B(B[166]), .A(n80), .Z(n35905) );
  XNOR U36483 ( .A(n35913), .B(n36243), .Z(n35906) );
  XNOR U36484 ( .A(n35912), .B(n35910), .Z(n36243) );
  AND U36485 ( .A(n36244), .B(n36245), .Z(n35910) );
  NANDN U36486 ( .A(n36246), .B(n36247), .Z(n36245) );
  OR U36487 ( .A(n36248), .B(n36249), .Z(n36247) );
  NAND U36488 ( .A(n36249), .B(n36248), .Z(n36244) );
  ANDN U36489 ( .B(B[167]), .A(n81), .Z(n35912) );
  XNOR U36490 ( .A(n35920), .B(n36250), .Z(n35913) );
  XNOR U36491 ( .A(n35919), .B(n35917), .Z(n36250) );
  AND U36492 ( .A(n36251), .B(n36252), .Z(n35917) );
  NANDN U36493 ( .A(n36253), .B(n36254), .Z(n36252) );
  NAND U36494 ( .A(n36255), .B(n36256), .Z(n36254) );
  ANDN U36495 ( .B(B[168]), .A(n82), .Z(n35919) );
  XOR U36496 ( .A(n35926), .B(n36257), .Z(n35920) );
  XNOR U36497 ( .A(n35924), .B(n35927), .Z(n36257) );
  NAND U36498 ( .A(A[2]), .B(B[169]), .Z(n35927) );
  NANDN U36499 ( .A(n36258), .B(n36259), .Z(n35924) );
  AND U36500 ( .A(A[0]), .B(B[170]), .Z(n36259) );
  XNOR U36501 ( .A(n35929), .B(n36260), .Z(n35926) );
  NAND U36502 ( .A(A[0]), .B(B[171]), .Z(n36260) );
  NAND U36503 ( .A(B[170]), .B(A[1]), .Z(n35929) );
  NAND U36504 ( .A(n36261), .B(n36262), .Z(n454) );
  NANDN U36505 ( .A(n36263), .B(n36264), .Z(n36262) );
  OR U36506 ( .A(n36265), .B(n36266), .Z(n36264) );
  NAND U36507 ( .A(n36266), .B(n36265), .Z(n36261) );
  XOR U36508 ( .A(n456), .B(n455), .Z(\A1[168] ) );
  XOR U36509 ( .A(n36266), .B(n36267), .Z(n455) );
  XNOR U36510 ( .A(n36265), .B(n36263), .Z(n36267) );
  AND U36511 ( .A(n36268), .B(n36269), .Z(n36263) );
  NANDN U36512 ( .A(n36270), .B(n36271), .Z(n36269) );
  NANDN U36513 ( .A(n36272), .B(n36273), .Z(n36271) );
  NANDN U36514 ( .A(n36273), .B(n36272), .Z(n36268) );
  ANDN U36515 ( .B(B[139]), .A(n54), .Z(n36265) );
  XNOR U36516 ( .A(n36060), .B(n36274), .Z(n36266) );
  XNOR U36517 ( .A(n36059), .B(n36057), .Z(n36274) );
  AND U36518 ( .A(n36275), .B(n36276), .Z(n36057) );
  NANDN U36519 ( .A(n36277), .B(n36278), .Z(n36276) );
  OR U36520 ( .A(n36279), .B(n36280), .Z(n36278) );
  NAND U36521 ( .A(n36280), .B(n36279), .Z(n36275) );
  ANDN U36522 ( .B(B[140]), .A(n55), .Z(n36059) );
  XNOR U36523 ( .A(n36067), .B(n36281), .Z(n36060) );
  XNOR U36524 ( .A(n36066), .B(n36064), .Z(n36281) );
  AND U36525 ( .A(n36282), .B(n36283), .Z(n36064) );
  NANDN U36526 ( .A(n36284), .B(n36285), .Z(n36283) );
  NANDN U36527 ( .A(n36286), .B(n36287), .Z(n36285) );
  NANDN U36528 ( .A(n36287), .B(n36286), .Z(n36282) );
  ANDN U36529 ( .B(B[141]), .A(n56), .Z(n36066) );
  XNOR U36530 ( .A(n36074), .B(n36288), .Z(n36067) );
  XNOR U36531 ( .A(n36073), .B(n36071), .Z(n36288) );
  AND U36532 ( .A(n36289), .B(n36290), .Z(n36071) );
  NANDN U36533 ( .A(n36291), .B(n36292), .Z(n36290) );
  OR U36534 ( .A(n36293), .B(n36294), .Z(n36292) );
  NAND U36535 ( .A(n36294), .B(n36293), .Z(n36289) );
  ANDN U36536 ( .B(B[142]), .A(n57), .Z(n36073) );
  XNOR U36537 ( .A(n36081), .B(n36295), .Z(n36074) );
  XNOR U36538 ( .A(n36080), .B(n36078), .Z(n36295) );
  AND U36539 ( .A(n36296), .B(n36297), .Z(n36078) );
  NANDN U36540 ( .A(n36298), .B(n36299), .Z(n36297) );
  NANDN U36541 ( .A(n36300), .B(n36301), .Z(n36299) );
  NANDN U36542 ( .A(n36301), .B(n36300), .Z(n36296) );
  ANDN U36543 ( .B(B[143]), .A(n58), .Z(n36080) );
  XNOR U36544 ( .A(n36088), .B(n36302), .Z(n36081) );
  XNOR U36545 ( .A(n36087), .B(n36085), .Z(n36302) );
  AND U36546 ( .A(n36303), .B(n36304), .Z(n36085) );
  NANDN U36547 ( .A(n36305), .B(n36306), .Z(n36304) );
  OR U36548 ( .A(n36307), .B(n36308), .Z(n36306) );
  NAND U36549 ( .A(n36308), .B(n36307), .Z(n36303) );
  ANDN U36550 ( .B(B[144]), .A(n59), .Z(n36087) );
  XNOR U36551 ( .A(n36095), .B(n36309), .Z(n36088) );
  XNOR U36552 ( .A(n36094), .B(n36092), .Z(n36309) );
  AND U36553 ( .A(n36310), .B(n36311), .Z(n36092) );
  NANDN U36554 ( .A(n36312), .B(n36313), .Z(n36311) );
  NANDN U36555 ( .A(n36314), .B(n36315), .Z(n36313) );
  NANDN U36556 ( .A(n36315), .B(n36314), .Z(n36310) );
  ANDN U36557 ( .B(B[145]), .A(n60), .Z(n36094) );
  XNOR U36558 ( .A(n36102), .B(n36316), .Z(n36095) );
  XNOR U36559 ( .A(n36101), .B(n36099), .Z(n36316) );
  AND U36560 ( .A(n36317), .B(n36318), .Z(n36099) );
  NANDN U36561 ( .A(n36319), .B(n36320), .Z(n36318) );
  OR U36562 ( .A(n36321), .B(n36322), .Z(n36320) );
  NAND U36563 ( .A(n36322), .B(n36321), .Z(n36317) );
  ANDN U36564 ( .B(B[146]), .A(n61), .Z(n36101) );
  XNOR U36565 ( .A(n36109), .B(n36323), .Z(n36102) );
  XNOR U36566 ( .A(n36108), .B(n36106), .Z(n36323) );
  AND U36567 ( .A(n36324), .B(n36325), .Z(n36106) );
  NANDN U36568 ( .A(n36326), .B(n36327), .Z(n36325) );
  NANDN U36569 ( .A(n36328), .B(n36329), .Z(n36327) );
  NANDN U36570 ( .A(n36329), .B(n36328), .Z(n36324) );
  ANDN U36571 ( .B(B[147]), .A(n62), .Z(n36108) );
  XNOR U36572 ( .A(n36116), .B(n36330), .Z(n36109) );
  XNOR U36573 ( .A(n36115), .B(n36113), .Z(n36330) );
  AND U36574 ( .A(n36331), .B(n36332), .Z(n36113) );
  NANDN U36575 ( .A(n36333), .B(n36334), .Z(n36332) );
  OR U36576 ( .A(n36335), .B(n36336), .Z(n36334) );
  NAND U36577 ( .A(n36336), .B(n36335), .Z(n36331) );
  ANDN U36578 ( .B(B[148]), .A(n63), .Z(n36115) );
  XNOR U36579 ( .A(n36123), .B(n36337), .Z(n36116) );
  XNOR U36580 ( .A(n36122), .B(n36120), .Z(n36337) );
  AND U36581 ( .A(n36338), .B(n36339), .Z(n36120) );
  NANDN U36582 ( .A(n36340), .B(n36341), .Z(n36339) );
  NANDN U36583 ( .A(n36342), .B(n36343), .Z(n36341) );
  NANDN U36584 ( .A(n36343), .B(n36342), .Z(n36338) );
  ANDN U36585 ( .B(B[149]), .A(n64), .Z(n36122) );
  XNOR U36586 ( .A(n36130), .B(n36344), .Z(n36123) );
  XNOR U36587 ( .A(n36129), .B(n36127), .Z(n36344) );
  AND U36588 ( .A(n36345), .B(n36346), .Z(n36127) );
  NANDN U36589 ( .A(n36347), .B(n36348), .Z(n36346) );
  OR U36590 ( .A(n36349), .B(n36350), .Z(n36348) );
  NAND U36591 ( .A(n36350), .B(n36349), .Z(n36345) );
  ANDN U36592 ( .B(B[150]), .A(n65), .Z(n36129) );
  XNOR U36593 ( .A(n36137), .B(n36351), .Z(n36130) );
  XNOR U36594 ( .A(n36136), .B(n36134), .Z(n36351) );
  AND U36595 ( .A(n36352), .B(n36353), .Z(n36134) );
  NANDN U36596 ( .A(n36354), .B(n36355), .Z(n36353) );
  NANDN U36597 ( .A(n36356), .B(n36357), .Z(n36355) );
  NANDN U36598 ( .A(n36357), .B(n36356), .Z(n36352) );
  ANDN U36599 ( .B(B[151]), .A(n66), .Z(n36136) );
  XNOR U36600 ( .A(n36144), .B(n36358), .Z(n36137) );
  XNOR U36601 ( .A(n36143), .B(n36141), .Z(n36358) );
  AND U36602 ( .A(n36359), .B(n36360), .Z(n36141) );
  NANDN U36603 ( .A(n36361), .B(n36362), .Z(n36360) );
  OR U36604 ( .A(n36363), .B(n36364), .Z(n36362) );
  NAND U36605 ( .A(n36364), .B(n36363), .Z(n36359) );
  ANDN U36606 ( .B(B[152]), .A(n67), .Z(n36143) );
  XNOR U36607 ( .A(n36151), .B(n36365), .Z(n36144) );
  XNOR U36608 ( .A(n36150), .B(n36148), .Z(n36365) );
  AND U36609 ( .A(n36366), .B(n36367), .Z(n36148) );
  NANDN U36610 ( .A(n36368), .B(n36369), .Z(n36367) );
  NANDN U36611 ( .A(n36370), .B(n36371), .Z(n36369) );
  NANDN U36612 ( .A(n36371), .B(n36370), .Z(n36366) );
  ANDN U36613 ( .B(B[153]), .A(n68), .Z(n36150) );
  XNOR U36614 ( .A(n36158), .B(n36372), .Z(n36151) );
  XNOR U36615 ( .A(n36157), .B(n36155), .Z(n36372) );
  AND U36616 ( .A(n36373), .B(n36374), .Z(n36155) );
  NANDN U36617 ( .A(n36375), .B(n36376), .Z(n36374) );
  OR U36618 ( .A(n36377), .B(n36378), .Z(n36376) );
  NAND U36619 ( .A(n36378), .B(n36377), .Z(n36373) );
  ANDN U36620 ( .B(B[154]), .A(n69), .Z(n36157) );
  XNOR U36621 ( .A(n36165), .B(n36379), .Z(n36158) );
  XNOR U36622 ( .A(n36164), .B(n36162), .Z(n36379) );
  AND U36623 ( .A(n36380), .B(n36381), .Z(n36162) );
  NANDN U36624 ( .A(n36382), .B(n36383), .Z(n36381) );
  NANDN U36625 ( .A(n36384), .B(n36385), .Z(n36383) );
  NANDN U36626 ( .A(n36385), .B(n36384), .Z(n36380) );
  ANDN U36627 ( .B(B[155]), .A(n70), .Z(n36164) );
  XNOR U36628 ( .A(n36172), .B(n36386), .Z(n36165) );
  XNOR U36629 ( .A(n36171), .B(n36169), .Z(n36386) );
  AND U36630 ( .A(n36387), .B(n36388), .Z(n36169) );
  NANDN U36631 ( .A(n36389), .B(n36390), .Z(n36388) );
  OR U36632 ( .A(n36391), .B(n36392), .Z(n36390) );
  NAND U36633 ( .A(n36392), .B(n36391), .Z(n36387) );
  ANDN U36634 ( .B(B[156]), .A(n71), .Z(n36171) );
  XNOR U36635 ( .A(n36179), .B(n36393), .Z(n36172) );
  XNOR U36636 ( .A(n36178), .B(n36176), .Z(n36393) );
  AND U36637 ( .A(n36394), .B(n36395), .Z(n36176) );
  NANDN U36638 ( .A(n36396), .B(n36397), .Z(n36395) );
  NANDN U36639 ( .A(n36398), .B(n36399), .Z(n36397) );
  NANDN U36640 ( .A(n36399), .B(n36398), .Z(n36394) );
  ANDN U36641 ( .B(B[157]), .A(n72), .Z(n36178) );
  XNOR U36642 ( .A(n36186), .B(n36400), .Z(n36179) );
  XNOR U36643 ( .A(n36185), .B(n36183), .Z(n36400) );
  AND U36644 ( .A(n36401), .B(n36402), .Z(n36183) );
  NANDN U36645 ( .A(n36403), .B(n36404), .Z(n36402) );
  OR U36646 ( .A(n36405), .B(n36406), .Z(n36404) );
  NAND U36647 ( .A(n36406), .B(n36405), .Z(n36401) );
  ANDN U36648 ( .B(B[158]), .A(n73), .Z(n36185) );
  XNOR U36649 ( .A(n36193), .B(n36407), .Z(n36186) );
  XNOR U36650 ( .A(n36192), .B(n36190), .Z(n36407) );
  AND U36651 ( .A(n36408), .B(n36409), .Z(n36190) );
  NANDN U36652 ( .A(n36410), .B(n36411), .Z(n36409) );
  NANDN U36653 ( .A(n36412), .B(n36413), .Z(n36411) );
  NANDN U36654 ( .A(n36413), .B(n36412), .Z(n36408) );
  ANDN U36655 ( .B(B[159]), .A(n74), .Z(n36192) );
  XNOR U36656 ( .A(n36200), .B(n36414), .Z(n36193) );
  XNOR U36657 ( .A(n36199), .B(n36197), .Z(n36414) );
  AND U36658 ( .A(n36415), .B(n36416), .Z(n36197) );
  NANDN U36659 ( .A(n36417), .B(n36418), .Z(n36416) );
  OR U36660 ( .A(n36419), .B(n36420), .Z(n36418) );
  NAND U36661 ( .A(n36420), .B(n36419), .Z(n36415) );
  ANDN U36662 ( .B(B[160]), .A(n75), .Z(n36199) );
  XNOR U36663 ( .A(n36207), .B(n36421), .Z(n36200) );
  XNOR U36664 ( .A(n36206), .B(n36204), .Z(n36421) );
  AND U36665 ( .A(n36422), .B(n36423), .Z(n36204) );
  NANDN U36666 ( .A(n36424), .B(n36425), .Z(n36423) );
  NANDN U36667 ( .A(n36426), .B(n36427), .Z(n36425) );
  NANDN U36668 ( .A(n36427), .B(n36426), .Z(n36422) );
  ANDN U36669 ( .B(B[161]), .A(n76), .Z(n36206) );
  XNOR U36670 ( .A(n36214), .B(n36428), .Z(n36207) );
  XNOR U36671 ( .A(n36213), .B(n36211), .Z(n36428) );
  AND U36672 ( .A(n36429), .B(n36430), .Z(n36211) );
  NANDN U36673 ( .A(n36431), .B(n36432), .Z(n36430) );
  OR U36674 ( .A(n36433), .B(n36434), .Z(n36432) );
  NAND U36675 ( .A(n36434), .B(n36433), .Z(n36429) );
  ANDN U36676 ( .B(B[162]), .A(n77), .Z(n36213) );
  XNOR U36677 ( .A(n36221), .B(n36435), .Z(n36214) );
  XNOR U36678 ( .A(n36220), .B(n36218), .Z(n36435) );
  AND U36679 ( .A(n36436), .B(n36437), .Z(n36218) );
  NANDN U36680 ( .A(n36438), .B(n36439), .Z(n36437) );
  NANDN U36681 ( .A(n36440), .B(n36441), .Z(n36439) );
  NANDN U36682 ( .A(n36441), .B(n36440), .Z(n36436) );
  ANDN U36683 ( .B(B[163]), .A(n78), .Z(n36220) );
  XNOR U36684 ( .A(n36228), .B(n36442), .Z(n36221) );
  XNOR U36685 ( .A(n36227), .B(n36225), .Z(n36442) );
  AND U36686 ( .A(n36443), .B(n36444), .Z(n36225) );
  NANDN U36687 ( .A(n36445), .B(n36446), .Z(n36444) );
  OR U36688 ( .A(n36447), .B(n36448), .Z(n36446) );
  NAND U36689 ( .A(n36448), .B(n36447), .Z(n36443) );
  ANDN U36690 ( .B(B[164]), .A(n79), .Z(n36227) );
  XNOR U36691 ( .A(n36235), .B(n36449), .Z(n36228) );
  XNOR U36692 ( .A(n36234), .B(n36232), .Z(n36449) );
  AND U36693 ( .A(n36450), .B(n36451), .Z(n36232) );
  NANDN U36694 ( .A(n36452), .B(n36453), .Z(n36451) );
  NANDN U36695 ( .A(n36454), .B(n36455), .Z(n36453) );
  NANDN U36696 ( .A(n36455), .B(n36454), .Z(n36450) );
  ANDN U36697 ( .B(B[165]), .A(n80), .Z(n36234) );
  XNOR U36698 ( .A(n36242), .B(n36456), .Z(n36235) );
  XNOR U36699 ( .A(n36241), .B(n36239), .Z(n36456) );
  AND U36700 ( .A(n36457), .B(n36458), .Z(n36239) );
  NANDN U36701 ( .A(n36459), .B(n36460), .Z(n36458) );
  OR U36702 ( .A(n36461), .B(n36462), .Z(n36460) );
  NAND U36703 ( .A(n36462), .B(n36461), .Z(n36457) );
  ANDN U36704 ( .B(B[166]), .A(n81), .Z(n36241) );
  XNOR U36705 ( .A(n36249), .B(n36463), .Z(n36242) );
  XNOR U36706 ( .A(n36248), .B(n36246), .Z(n36463) );
  AND U36707 ( .A(n36464), .B(n36465), .Z(n36246) );
  NANDN U36708 ( .A(n36466), .B(n36467), .Z(n36465) );
  NAND U36709 ( .A(n36468), .B(n36469), .Z(n36467) );
  ANDN U36710 ( .B(B[167]), .A(n82), .Z(n36248) );
  XOR U36711 ( .A(n36255), .B(n36470), .Z(n36249) );
  XNOR U36712 ( .A(n36253), .B(n36256), .Z(n36470) );
  NAND U36713 ( .A(A[2]), .B(B[168]), .Z(n36256) );
  NANDN U36714 ( .A(n36471), .B(n36472), .Z(n36253) );
  AND U36715 ( .A(A[0]), .B(B[169]), .Z(n36472) );
  XNOR U36716 ( .A(n36258), .B(n36473), .Z(n36255) );
  NAND U36717 ( .A(A[0]), .B(B[170]), .Z(n36473) );
  NAND U36718 ( .A(B[169]), .B(A[1]), .Z(n36258) );
  NAND U36719 ( .A(n36474), .B(n36475), .Z(n456) );
  NANDN U36720 ( .A(n36476), .B(n36477), .Z(n36475) );
  OR U36721 ( .A(n36478), .B(n36479), .Z(n36477) );
  NAND U36722 ( .A(n36479), .B(n36478), .Z(n36474) );
  XOR U36723 ( .A(n458), .B(n457), .Z(\A1[167] ) );
  XOR U36724 ( .A(n36479), .B(n36480), .Z(n457) );
  XNOR U36725 ( .A(n36478), .B(n36476), .Z(n36480) );
  AND U36726 ( .A(n36481), .B(n36482), .Z(n36476) );
  NANDN U36727 ( .A(n36483), .B(n36484), .Z(n36482) );
  NANDN U36728 ( .A(n36485), .B(n36486), .Z(n36484) );
  NANDN U36729 ( .A(n36486), .B(n36485), .Z(n36481) );
  ANDN U36730 ( .B(B[138]), .A(n54), .Z(n36478) );
  XNOR U36731 ( .A(n36273), .B(n36487), .Z(n36479) );
  XNOR U36732 ( .A(n36272), .B(n36270), .Z(n36487) );
  AND U36733 ( .A(n36488), .B(n36489), .Z(n36270) );
  NANDN U36734 ( .A(n36490), .B(n36491), .Z(n36489) );
  OR U36735 ( .A(n36492), .B(n36493), .Z(n36491) );
  NAND U36736 ( .A(n36493), .B(n36492), .Z(n36488) );
  ANDN U36737 ( .B(B[139]), .A(n55), .Z(n36272) );
  XNOR U36738 ( .A(n36280), .B(n36494), .Z(n36273) );
  XNOR U36739 ( .A(n36279), .B(n36277), .Z(n36494) );
  AND U36740 ( .A(n36495), .B(n36496), .Z(n36277) );
  NANDN U36741 ( .A(n36497), .B(n36498), .Z(n36496) );
  NANDN U36742 ( .A(n36499), .B(n36500), .Z(n36498) );
  NANDN U36743 ( .A(n36500), .B(n36499), .Z(n36495) );
  ANDN U36744 ( .B(B[140]), .A(n56), .Z(n36279) );
  XNOR U36745 ( .A(n36287), .B(n36501), .Z(n36280) );
  XNOR U36746 ( .A(n36286), .B(n36284), .Z(n36501) );
  AND U36747 ( .A(n36502), .B(n36503), .Z(n36284) );
  NANDN U36748 ( .A(n36504), .B(n36505), .Z(n36503) );
  OR U36749 ( .A(n36506), .B(n36507), .Z(n36505) );
  NAND U36750 ( .A(n36507), .B(n36506), .Z(n36502) );
  ANDN U36751 ( .B(B[141]), .A(n57), .Z(n36286) );
  XNOR U36752 ( .A(n36294), .B(n36508), .Z(n36287) );
  XNOR U36753 ( .A(n36293), .B(n36291), .Z(n36508) );
  AND U36754 ( .A(n36509), .B(n36510), .Z(n36291) );
  NANDN U36755 ( .A(n36511), .B(n36512), .Z(n36510) );
  NANDN U36756 ( .A(n36513), .B(n36514), .Z(n36512) );
  NANDN U36757 ( .A(n36514), .B(n36513), .Z(n36509) );
  ANDN U36758 ( .B(B[142]), .A(n58), .Z(n36293) );
  XNOR U36759 ( .A(n36301), .B(n36515), .Z(n36294) );
  XNOR U36760 ( .A(n36300), .B(n36298), .Z(n36515) );
  AND U36761 ( .A(n36516), .B(n36517), .Z(n36298) );
  NANDN U36762 ( .A(n36518), .B(n36519), .Z(n36517) );
  OR U36763 ( .A(n36520), .B(n36521), .Z(n36519) );
  NAND U36764 ( .A(n36521), .B(n36520), .Z(n36516) );
  ANDN U36765 ( .B(B[143]), .A(n59), .Z(n36300) );
  XNOR U36766 ( .A(n36308), .B(n36522), .Z(n36301) );
  XNOR U36767 ( .A(n36307), .B(n36305), .Z(n36522) );
  AND U36768 ( .A(n36523), .B(n36524), .Z(n36305) );
  NANDN U36769 ( .A(n36525), .B(n36526), .Z(n36524) );
  NANDN U36770 ( .A(n36527), .B(n36528), .Z(n36526) );
  NANDN U36771 ( .A(n36528), .B(n36527), .Z(n36523) );
  ANDN U36772 ( .B(B[144]), .A(n60), .Z(n36307) );
  XNOR U36773 ( .A(n36315), .B(n36529), .Z(n36308) );
  XNOR U36774 ( .A(n36314), .B(n36312), .Z(n36529) );
  AND U36775 ( .A(n36530), .B(n36531), .Z(n36312) );
  NANDN U36776 ( .A(n36532), .B(n36533), .Z(n36531) );
  OR U36777 ( .A(n36534), .B(n36535), .Z(n36533) );
  NAND U36778 ( .A(n36535), .B(n36534), .Z(n36530) );
  ANDN U36779 ( .B(B[145]), .A(n61), .Z(n36314) );
  XNOR U36780 ( .A(n36322), .B(n36536), .Z(n36315) );
  XNOR U36781 ( .A(n36321), .B(n36319), .Z(n36536) );
  AND U36782 ( .A(n36537), .B(n36538), .Z(n36319) );
  NANDN U36783 ( .A(n36539), .B(n36540), .Z(n36538) );
  NANDN U36784 ( .A(n36541), .B(n36542), .Z(n36540) );
  NANDN U36785 ( .A(n36542), .B(n36541), .Z(n36537) );
  ANDN U36786 ( .B(B[146]), .A(n62), .Z(n36321) );
  XNOR U36787 ( .A(n36329), .B(n36543), .Z(n36322) );
  XNOR U36788 ( .A(n36328), .B(n36326), .Z(n36543) );
  AND U36789 ( .A(n36544), .B(n36545), .Z(n36326) );
  NANDN U36790 ( .A(n36546), .B(n36547), .Z(n36545) );
  OR U36791 ( .A(n36548), .B(n36549), .Z(n36547) );
  NAND U36792 ( .A(n36549), .B(n36548), .Z(n36544) );
  ANDN U36793 ( .B(B[147]), .A(n63), .Z(n36328) );
  XNOR U36794 ( .A(n36336), .B(n36550), .Z(n36329) );
  XNOR U36795 ( .A(n36335), .B(n36333), .Z(n36550) );
  AND U36796 ( .A(n36551), .B(n36552), .Z(n36333) );
  NANDN U36797 ( .A(n36553), .B(n36554), .Z(n36552) );
  NANDN U36798 ( .A(n36555), .B(n36556), .Z(n36554) );
  NANDN U36799 ( .A(n36556), .B(n36555), .Z(n36551) );
  ANDN U36800 ( .B(B[148]), .A(n64), .Z(n36335) );
  XNOR U36801 ( .A(n36343), .B(n36557), .Z(n36336) );
  XNOR U36802 ( .A(n36342), .B(n36340), .Z(n36557) );
  AND U36803 ( .A(n36558), .B(n36559), .Z(n36340) );
  NANDN U36804 ( .A(n36560), .B(n36561), .Z(n36559) );
  OR U36805 ( .A(n36562), .B(n36563), .Z(n36561) );
  NAND U36806 ( .A(n36563), .B(n36562), .Z(n36558) );
  ANDN U36807 ( .B(B[149]), .A(n65), .Z(n36342) );
  XNOR U36808 ( .A(n36350), .B(n36564), .Z(n36343) );
  XNOR U36809 ( .A(n36349), .B(n36347), .Z(n36564) );
  AND U36810 ( .A(n36565), .B(n36566), .Z(n36347) );
  NANDN U36811 ( .A(n36567), .B(n36568), .Z(n36566) );
  NANDN U36812 ( .A(n36569), .B(n36570), .Z(n36568) );
  NANDN U36813 ( .A(n36570), .B(n36569), .Z(n36565) );
  ANDN U36814 ( .B(B[150]), .A(n66), .Z(n36349) );
  XNOR U36815 ( .A(n36357), .B(n36571), .Z(n36350) );
  XNOR U36816 ( .A(n36356), .B(n36354), .Z(n36571) );
  AND U36817 ( .A(n36572), .B(n36573), .Z(n36354) );
  NANDN U36818 ( .A(n36574), .B(n36575), .Z(n36573) );
  OR U36819 ( .A(n36576), .B(n36577), .Z(n36575) );
  NAND U36820 ( .A(n36577), .B(n36576), .Z(n36572) );
  ANDN U36821 ( .B(B[151]), .A(n67), .Z(n36356) );
  XNOR U36822 ( .A(n36364), .B(n36578), .Z(n36357) );
  XNOR U36823 ( .A(n36363), .B(n36361), .Z(n36578) );
  AND U36824 ( .A(n36579), .B(n36580), .Z(n36361) );
  NANDN U36825 ( .A(n36581), .B(n36582), .Z(n36580) );
  NANDN U36826 ( .A(n36583), .B(n36584), .Z(n36582) );
  NANDN U36827 ( .A(n36584), .B(n36583), .Z(n36579) );
  ANDN U36828 ( .B(B[152]), .A(n68), .Z(n36363) );
  XNOR U36829 ( .A(n36371), .B(n36585), .Z(n36364) );
  XNOR U36830 ( .A(n36370), .B(n36368), .Z(n36585) );
  AND U36831 ( .A(n36586), .B(n36587), .Z(n36368) );
  NANDN U36832 ( .A(n36588), .B(n36589), .Z(n36587) );
  OR U36833 ( .A(n36590), .B(n36591), .Z(n36589) );
  NAND U36834 ( .A(n36591), .B(n36590), .Z(n36586) );
  ANDN U36835 ( .B(B[153]), .A(n69), .Z(n36370) );
  XNOR U36836 ( .A(n36378), .B(n36592), .Z(n36371) );
  XNOR U36837 ( .A(n36377), .B(n36375), .Z(n36592) );
  AND U36838 ( .A(n36593), .B(n36594), .Z(n36375) );
  NANDN U36839 ( .A(n36595), .B(n36596), .Z(n36594) );
  NANDN U36840 ( .A(n36597), .B(n36598), .Z(n36596) );
  NANDN U36841 ( .A(n36598), .B(n36597), .Z(n36593) );
  ANDN U36842 ( .B(B[154]), .A(n70), .Z(n36377) );
  XNOR U36843 ( .A(n36385), .B(n36599), .Z(n36378) );
  XNOR U36844 ( .A(n36384), .B(n36382), .Z(n36599) );
  AND U36845 ( .A(n36600), .B(n36601), .Z(n36382) );
  NANDN U36846 ( .A(n36602), .B(n36603), .Z(n36601) );
  OR U36847 ( .A(n36604), .B(n36605), .Z(n36603) );
  NAND U36848 ( .A(n36605), .B(n36604), .Z(n36600) );
  ANDN U36849 ( .B(B[155]), .A(n71), .Z(n36384) );
  XNOR U36850 ( .A(n36392), .B(n36606), .Z(n36385) );
  XNOR U36851 ( .A(n36391), .B(n36389), .Z(n36606) );
  AND U36852 ( .A(n36607), .B(n36608), .Z(n36389) );
  NANDN U36853 ( .A(n36609), .B(n36610), .Z(n36608) );
  NANDN U36854 ( .A(n36611), .B(n36612), .Z(n36610) );
  NANDN U36855 ( .A(n36612), .B(n36611), .Z(n36607) );
  ANDN U36856 ( .B(B[156]), .A(n72), .Z(n36391) );
  XNOR U36857 ( .A(n36399), .B(n36613), .Z(n36392) );
  XNOR U36858 ( .A(n36398), .B(n36396), .Z(n36613) );
  AND U36859 ( .A(n36614), .B(n36615), .Z(n36396) );
  NANDN U36860 ( .A(n36616), .B(n36617), .Z(n36615) );
  OR U36861 ( .A(n36618), .B(n36619), .Z(n36617) );
  NAND U36862 ( .A(n36619), .B(n36618), .Z(n36614) );
  ANDN U36863 ( .B(B[157]), .A(n73), .Z(n36398) );
  XNOR U36864 ( .A(n36406), .B(n36620), .Z(n36399) );
  XNOR U36865 ( .A(n36405), .B(n36403), .Z(n36620) );
  AND U36866 ( .A(n36621), .B(n36622), .Z(n36403) );
  NANDN U36867 ( .A(n36623), .B(n36624), .Z(n36622) );
  NANDN U36868 ( .A(n36625), .B(n36626), .Z(n36624) );
  NANDN U36869 ( .A(n36626), .B(n36625), .Z(n36621) );
  ANDN U36870 ( .B(B[158]), .A(n74), .Z(n36405) );
  XNOR U36871 ( .A(n36413), .B(n36627), .Z(n36406) );
  XNOR U36872 ( .A(n36412), .B(n36410), .Z(n36627) );
  AND U36873 ( .A(n36628), .B(n36629), .Z(n36410) );
  NANDN U36874 ( .A(n36630), .B(n36631), .Z(n36629) );
  OR U36875 ( .A(n36632), .B(n36633), .Z(n36631) );
  NAND U36876 ( .A(n36633), .B(n36632), .Z(n36628) );
  ANDN U36877 ( .B(B[159]), .A(n75), .Z(n36412) );
  XNOR U36878 ( .A(n36420), .B(n36634), .Z(n36413) );
  XNOR U36879 ( .A(n36419), .B(n36417), .Z(n36634) );
  AND U36880 ( .A(n36635), .B(n36636), .Z(n36417) );
  NANDN U36881 ( .A(n36637), .B(n36638), .Z(n36636) );
  NANDN U36882 ( .A(n36639), .B(n36640), .Z(n36638) );
  NANDN U36883 ( .A(n36640), .B(n36639), .Z(n36635) );
  ANDN U36884 ( .B(B[160]), .A(n76), .Z(n36419) );
  XNOR U36885 ( .A(n36427), .B(n36641), .Z(n36420) );
  XNOR U36886 ( .A(n36426), .B(n36424), .Z(n36641) );
  AND U36887 ( .A(n36642), .B(n36643), .Z(n36424) );
  NANDN U36888 ( .A(n36644), .B(n36645), .Z(n36643) );
  OR U36889 ( .A(n36646), .B(n36647), .Z(n36645) );
  NAND U36890 ( .A(n36647), .B(n36646), .Z(n36642) );
  ANDN U36891 ( .B(B[161]), .A(n77), .Z(n36426) );
  XNOR U36892 ( .A(n36434), .B(n36648), .Z(n36427) );
  XNOR U36893 ( .A(n36433), .B(n36431), .Z(n36648) );
  AND U36894 ( .A(n36649), .B(n36650), .Z(n36431) );
  NANDN U36895 ( .A(n36651), .B(n36652), .Z(n36650) );
  NANDN U36896 ( .A(n36653), .B(n36654), .Z(n36652) );
  NANDN U36897 ( .A(n36654), .B(n36653), .Z(n36649) );
  ANDN U36898 ( .B(B[162]), .A(n78), .Z(n36433) );
  XNOR U36899 ( .A(n36441), .B(n36655), .Z(n36434) );
  XNOR U36900 ( .A(n36440), .B(n36438), .Z(n36655) );
  AND U36901 ( .A(n36656), .B(n36657), .Z(n36438) );
  NANDN U36902 ( .A(n36658), .B(n36659), .Z(n36657) );
  OR U36903 ( .A(n36660), .B(n36661), .Z(n36659) );
  NAND U36904 ( .A(n36661), .B(n36660), .Z(n36656) );
  ANDN U36905 ( .B(B[163]), .A(n79), .Z(n36440) );
  XNOR U36906 ( .A(n36448), .B(n36662), .Z(n36441) );
  XNOR U36907 ( .A(n36447), .B(n36445), .Z(n36662) );
  AND U36908 ( .A(n36663), .B(n36664), .Z(n36445) );
  NANDN U36909 ( .A(n36665), .B(n36666), .Z(n36664) );
  NANDN U36910 ( .A(n36667), .B(n36668), .Z(n36666) );
  NANDN U36911 ( .A(n36668), .B(n36667), .Z(n36663) );
  ANDN U36912 ( .B(B[164]), .A(n80), .Z(n36447) );
  XNOR U36913 ( .A(n36455), .B(n36669), .Z(n36448) );
  XNOR U36914 ( .A(n36454), .B(n36452), .Z(n36669) );
  AND U36915 ( .A(n36670), .B(n36671), .Z(n36452) );
  NANDN U36916 ( .A(n36672), .B(n36673), .Z(n36671) );
  OR U36917 ( .A(n36674), .B(n36675), .Z(n36673) );
  NAND U36918 ( .A(n36675), .B(n36674), .Z(n36670) );
  ANDN U36919 ( .B(B[165]), .A(n81), .Z(n36454) );
  XNOR U36920 ( .A(n36462), .B(n36676), .Z(n36455) );
  XNOR U36921 ( .A(n36461), .B(n36459), .Z(n36676) );
  AND U36922 ( .A(n36677), .B(n36678), .Z(n36459) );
  NANDN U36923 ( .A(n36679), .B(n36680), .Z(n36678) );
  NAND U36924 ( .A(n36681), .B(n36682), .Z(n36680) );
  ANDN U36925 ( .B(B[166]), .A(n82), .Z(n36461) );
  XOR U36926 ( .A(n36468), .B(n36683), .Z(n36462) );
  XNOR U36927 ( .A(n36466), .B(n36469), .Z(n36683) );
  NAND U36928 ( .A(A[2]), .B(B[167]), .Z(n36469) );
  NANDN U36929 ( .A(n36684), .B(n36685), .Z(n36466) );
  AND U36930 ( .A(A[0]), .B(B[168]), .Z(n36685) );
  XNOR U36931 ( .A(n36471), .B(n36686), .Z(n36468) );
  NAND U36932 ( .A(A[0]), .B(B[169]), .Z(n36686) );
  NAND U36933 ( .A(B[168]), .B(A[1]), .Z(n36471) );
  NAND U36934 ( .A(n36687), .B(n36688), .Z(n458) );
  NANDN U36935 ( .A(n36689), .B(n36690), .Z(n36688) );
  OR U36936 ( .A(n36691), .B(n36692), .Z(n36690) );
  NAND U36937 ( .A(n36692), .B(n36691), .Z(n36687) );
  XOR U36938 ( .A(n460), .B(n459), .Z(\A1[166] ) );
  XOR U36939 ( .A(n36692), .B(n36693), .Z(n459) );
  XNOR U36940 ( .A(n36691), .B(n36689), .Z(n36693) );
  AND U36941 ( .A(n36694), .B(n36695), .Z(n36689) );
  NANDN U36942 ( .A(n36696), .B(n36697), .Z(n36695) );
  NANDN U36943 ( .A(n36698), .B(n36699), .Z(n36697) );
  NANDN U36944 ( .A(n36699), .B(n36698), .Z(n36694) );
  ANDN U36945 ( .B(B[137]), .A(n54), .Z(n36691) );
  XNOR U36946 ( .A(n36486), .B(n36700), .Z(n36692) );
  XNOR U36947 ( .A(n36485), .B(n36483), .Z(n36700) );
  AND U36948 ( .A(n36701), .B(n36702), .Z(n36483) );
  NANDN U36949 ( .A(n36703), .B(n36704), .Z(n36702) );
  OR U36950 ( .A(n36705), .B(n36706), .Z(n36704) );
  NAND U36951 ( .A(n36706), .B(n36705), .Z(n36701) );
  ANDN U36952 ( .B(B[138]), .A(n55), .Z(n36485) );
  XNOR U36953 ( .A(n36493), .B(n36707), .Z(n36486) );
  XNOR U36954 ( .A(n36492), .B(n36490), .Z(n36707) );
  AND U36955 ( .A(n36708), .B(n36709), .Z(n36490) );
  NANDN U36956 ( .A(n36710), .B(n36711), .Z(n36709) );
  NANDN U36957 ( .A(n36712), .B(n36713), .Z(n36711) );
  NANDN U36958 ( .A(n36713), .B(n36712), .Z(n36708) );
  ANDN U36959 ( .B(B[139]), .A(n56), .Z(n36492) );
  XNOR U36960 ( .A(n36500), .B(n36714), .Z(n36493) );
  XNOR U36961 ( .A(n36499), .B(n36497), .Z(n36714) );
  AND U36962 ( .A(n36715), .B(n36716), .Z(n36497) );
  NANDN U36963 ( .A(n36717), .B(n36718), .Z(n36716) );
  OR U36964 ( .A(n36719), .B(n36720), .Z(n36718) );
  NAND U36965 ( .A(n36720), .B(n36719), .Z(n36715) );
  ANDN U36966 ( .B(B[140]), .A(n57), .Z(n36499) );
  XNOR U36967 ( .A(n36507), .B(n36721), .Z(n36500) );
  XNOR U36968 ( .A(n36506), .B(n36504), .Z(n36721) );
  AND U36969 ( .A(n36722), .B(n36723), .Z(n36504) );
  NANDN U36970 ( .A(n36724), .B(n36725), .Z(n36723) );
  NANDN U36971 ( .A(n36726), .B(n36727), .Z(n36725) );
  NANDN U36972 ( .A(n36727), .B(n36726), .Z(n36722) );
  ANDN U36973 ( .B(B[141]), .A(n58), .Z(n36506) );
  XNOR U36974 ( .A(n36514), .B(n36728), .Z(n36507) );
  XNOR U36975 ( .A(n36513), .B(n36511), .Z(n36728) );
  AND U36976 ( .A(n36729), .B(n36730), .Z(n36511) );
  NANDN U36977 ( .A(n36731), .B(n36732), .Z(n36730) );
  OR U36978 ( .A(n36733), .B(n36734), .Z(n36732) );
  NAND U36979 ( .A(n36734), .B(n36733), .Z(n36729) );
  ANDN U36980 ( .B(B[142]), .A(n59), .Z(n36513) );
  XNOR U36981 ( .A(n36521), .B(n36735), .Z(n36514) );
  XNOR U36982 ( .A(n36520), .B(n36518), .Z(n36735) );
  AND U36983 ( .A(n36736), .B(n36737), .Z(n36518) );
  NANDN U36984 ( .A(n36738), .B(n36739), .Z(n36737) );
  NANDN U36985 ( .A(n36740), .B(n36741), .Z(n36739) );
  NANDN U36986 ( .A(n36741), .B(n36740), .Z(n36736) );
  ANDN U36987 ( .B(B[143]), .A(n60), .Z(n36520) );
  XNOR U36988 ( .A(n36528), .B(n36742), .Z(n36521) );
  XNOR U36989 ( .A(n36527), .B(n36525), .Z(n36742) );
  AND U36990 ( .A(n36743), .B(n36744), .Z(n36525) );
  NANDN U36991 ( .A(n36745), .B(n36746), .Z(n36744) );
  OR U36992 ( .A(n36747), .B(n36748), .Z(n36746) );
  NAND U36993 ( .A(n36748), .B(n36747), .Z(n36743) );
  ANDN U36994 ( .B(B[144]), .A(n61), .Z(n36527) );
  XNOR U36995 ( .A(n36535), .B(n36749), .Z(n36528) );
  XNOR U36996 ( .A(n36534), .B(n36532), .Z(n36749) );
  AND U36997 ( .A(n36750), .B(n36751), .Z(n36532) );
  NANDN U36998 ( .A(n36752), .B(n36753), .Z(n36751) );
  NANDN U36999 ( .A(n36754), .B(n36755), .Z(n36753) );
  NANDN U37000 ( .A(n36755), .B(n36754), .Z(n36750) );
  ANDN U37001 ( .B(B[145]), .A(n62), .Z(n36534) );
  XNOR U37002 ( .A(n36542), .B(n36756), .Z(n36535) );
  XNOR U37003 ( .A(n36541), .B(n36539), .Z(n36756) );
  AND U37004 ( .A(n36757), .B(n36758), .Z(n36539) );
  NANDN U37005 ( .A(n36759), .B(n36760), .Z(n36758) );
  OR U37006 ( .A(n36761), .B(n36762), .Z(n36760) );
  NAND U37007 ( .A(n36762), .B(n36761), .Z(n36757) );
  ANDN U37008 ( .B(B[146]), .A(n63), .Z(n36541) );
  XNOR U37009 ( .A(n36549), .B(n36763), .Z(n36542) );
  XNOR U37010 ( .A(n36548), .B(n36546), .Z(n36763) );
  AND U37011 ( .A(n36764), .B(n36765), .Z(n36546) );
  NANDN U37012 ( .A(n36766), .B(n36767), .Z(n36765) );
  NANDN U37013 ( .A(n36768), .B(n36769), .Z(n36767) );
  NANDN U37014 ( .A(n36769), .B(n36768), .Z(n36764) );
  ANDN U37015 ( .B(B[147]), .A(n64), .Z(n36548) );
  XNOR U37016 ( .A(n36556), .B(n36770), .Z(n36549) );
  XNOR U37017 ( .A(n36555), .B(n36553), .Z(n36770) );
  AND U37018 ( .A(n36771), .B(n36772), .Z(n36553) );
  NANDN U37019 ( .A(n36773), .B(n36774), .Z(n36772) );
  OR U37020 ( .A(n36775), .B(n36776), .Z(n36774) );
  NAND U37021 ( .A(n36776), .B(n36775), .Z(n36771) );
  ANDN U37022 ( .B(B[148]), .A(n65), .Z(n36555) );
  XNOR U37023 ( .A(n36563), .B(n36777), .Z(n36556) );
  XNOR U37024 ( .A(n36562), .B(n36560), .Z(n36777) );
  AND U37025 ( .A(n36778), .B(n36779), .Z(n36560) );
  NANDN U37026 ( .A(n36780), .B(n36781), .Z(n36779) );
  NANDN U37027 ( .A(n36782), .B(n36783), .Z(n36781) );
  NANDN U37028 ( .A(n36783), .B(n36782), .Z(n36778) );
  ANDN U37029 ( .B(B[149]), .A(n66), .Z(n36562) );
  XNOR U37030 ( .A(n36570), .B(n36784), .Z(n36563) );
  XNOR U37031 ( .A(n36569), .B(n36567), .Z(n36784) );
  AND U37032 ( .A(n36785), .B(n36786), .Z(n36567) );
  NANDN U37033 ( .A(n36787), .B(n36788), .Z(n36786) );
  OR U37034 ( .A(n36789), .B(n36790), .Z(n36788) );
  NAND U37035 ( .A(n36790), .B(n36789), .Z(n36785) );
  ANDN U37036 ( .B(B[150]), .A(n67), .Z(n36569) );
  XNOR U37037 ( .A(n36577), .B(n36791), .Z(n36570) );
  XNOR U37038 ( .A(n36576), .B(n36574), .Z(n36791) );
  AND U37039 ( .A(n36792), .B(n36793), .Z(n36574) );
  NANDN U37040 ( .A(n36794), .B(n36795), .Z(n36793) );
  NANDN U37041 ( .A(n36796), .B(n36797), .Z(n36795) );
  NANDN U37042 ( .A(n36797), .B(n36796), .Z(n36792) );
  ANDN U37043 ( .B(B[151]), .A(n68), .Z(n36576) );
  XNOR U37044 ( .A(n36584), .B(n36798), .Z(n36577) );
  XNOR U37045 ( .A(n36583), .B(n36581), .Z(n36798) );
  AND U37046 ( .A(n36799), .B(n36800), .Z(n36581) );
  NANDN U37047 ( .A(n36801), .B(n36802), .Z(n36800) );
  OR U37048 ( .A(n36803), .B(n36804), .Z(n36802) );
  NAND U37049 ( .A(n36804), .B(n36803), .Z(n36799) );
  ANDN U37050 ( .B(B[152]), .A(n69), .Z(n36583) );
  XNOR U37051 ( .A(n36591), .B(n36805), .Z(n36584) );
  XNOR U37052 ( .A(n36590), .B(n36588), .Z(n36805) );
  AND U37053 ( .A(n36806), .B(n36807), .Z(n36588) );
  NANDN U37054 ( .A(n36808), .B(n36809), .Z(n36807) );
  NANDN U37055 ( .A(n36810), .B(n36811), .Z(n36809) );
  NANDN U37056 ( .A(n36811), .B(n36810), .Z(n36806) );
  ANDN U37057 ( .B(B[153]), .A(n70), .Z(n36590) );
  XNOR U37058 ( .A(n36598), .B(n36812), .Z(n36591) );
  XNOR U37059 ( .A(n36597), .B(n36595), .Z(n36812) );
  AND U37060 ( .A(n36813), .B(n36814), .Z(n36595) );
  NANDN U37061 ( .A(n36815), .B(n36816), .Z(n36814) );
  OR U37062 ( .A(n36817), .B(n36818), .Z(n36816) );
  NAND U37063 ( .A(n36818), .B(n36817), .Z(n36813) );
  ANDN U37064 ( .B(B[154]), .A(n71), .Z(n36597) );
  XNOR U37065 ( .A(n36605), .B(n36819), .Z(n36598) );
  XNOR U37066 ( .A(n36604), .B(n36602), .Z(n36819) );
  AND U37067 ( .A(n36820), .B(n36821), .Z(n36602) );
  NANDN U37068 ( .A(n36822), .B(n36823), .Z(n36821) );
  NANDN U37069 ( .A(n36824), .B(n36825), .Z(n36823) );
  NANDN U37070 ( .A(n36825), .B(n36824), .Z(n36820) );
  ANDN U37071 ( .B(B[155]), .A(n72), .Z(n36604) );
  XNOR U37072 ( .A(n36612), .B(n36826), .Z(n36605) );
  XNOR U37073 ( .A(n36611), .B(n36609), .Z(n36826) );
  AND U37074 ( .A(n36827), .B(n36828), .Z(n36609) );
  NANDN U37075 ( .A(n36829), .B(n36830), .Z(n36828) );
  OR U37076 ( .A(n36831), .B(n36832), .Z(n36830) );
  NAND U37077 ( .A(n36832), .B(n36831), .Z(n36827) );
  ANDN U37078 ( .B(B[156]), .A(n73), .Z(n36611) );
  XNOR U37079 ( .A(n36619), .B(n36833), .Z(n36612) );
  XNOR U37080 ( .A(n36618), .B(n36616), .Z(n36833) );
  AND U37081 ( .A(n36834), .B(n36835), .Z(n36616) );
  NANDN U37082 ( .A(n36836), .B(n36837), .Z(n36835) );
  NANDN U37083 ( .A(n36838), .B(n36839), .Z(n36837) );
  NANDN U37084 ( .A(n36839), .B(n36838), .Z(n36834) );
  ANDN U37085 ( .B(B[157]), .A(n74), .Z(n36618) );
  XNOR U37086 ( .A(n36626), .B(n36840), .Z(n36619) );
  XNOR U37087 ( .A(n36625), .B(n36623), .Z(n36840) );
  AND U37088 ( .A(n36841), .B(n36842), .Z(n36623) );
  NANDN U37089 ( .A(n36843), .B(n36844), .Z(n36842) );
  OR U37090 ( .A(n36845), .B(n36846), .Z(n36844) );
  NAND U37091 ( .A(n36846), .B(n36845), .Z(n36841) );
  ANDN U37092 ( .B(B[158]), .A(n75), .Z(n36625) );
  XNOR U37093 ( .A(n36633), .B(n36847), .Z(n36626) );
  XNOR U37094 ( .A(n36632), .B(n36630), .Z(n36847) );
  AND U37095 ( .A(n36848), .B(n36849), .Z(n36630) );
  NANDN U37096 ( .A(n36850), .B(n36851), .Z(n36849) );
  NANDN U37097 ( .A(n36852), .B(n36853), .Z(n36851) );
  NANDN U37098 ( .A(n36853), .B(n36852), .Z(n36848) );
  ANDN U37099 ( .B(B[159]), .A(n76), .Z(n36632) );
  XNOR U37100 ( .A(n36640), .B(n36854), .Z(n36633) );
  XNOR U37101 ( .A(n36639), .B(n36637), .Z(n36854) );
  AND U37102 ( .A(n36855), .B(n36856), .Z(n36637) );
  NANDN U37103 ( .A(n36857), .B(n36858), .Z(n36856) );
  OR U37104 ( .A(n36859), .B(n36860), .Z(n36858) );
  NAND U37105 ( .A(n36860), .B(n36859), .Z(n36855) );
  ANDN U37106 ( .B(B[160]), .A(n77), .Z(n36639) );
  XNOR U37107 ( .A(n36647), .B(n36861), .Z(n36640) );
  XNOR U37108 ( .A(n36646), .B(n36644), .Z(n36861) );
  AND U37109 ( .A(n36862), .B(n36863), .Z(n36644) );
  NANDN U37110 ( .A(n36864), .B(n36865), .Z(n36863) );
  NANDN U37111 ( .A(n36866), .B(n36867), .Z(n36865) );
  NANDN U37112 ( .A(n36867), .B(n36866), .Z(n36862) );
  ANDN U37113 ( .B(B[161]), .A(n78), .Z(n36646) );
  XNOR U37114 ( .A(n36654), .B(n36868), .Z(n36647) );
  XNOR U37115 ( .A(n36653), .B(n36651), .Z(n36868) );
  AND U37116 ( .A(n36869), .B(n36870), .Z(n36651) );
  NANDN U37117 ( .A(n36871), .B(n36872), .Z(n36870) );
  OR U37118 ( .A(n36873), .B(n36874), .Z(n36872) );
  NAND U37119 ( .A(n36874), .B(n36873), .Z(n36869) );
  ANDN U37120 ( .B(B[162]), .A(n79), .Z(n36653) );
  XNOR U37121 ( .A(n36661), .B(n36875), .Z(n36654) );
  XNOR U37122 ( .A(n36660), .B(n36658), .Z(n36875) );
  AND U37123 ( .A(n36876), .B(n36877), .Z(n36658) );
  NANDN U37124 ( .A(n36878), .B(n36879), .Z(n36877) );
  NANDN U37125 ( .A(n36880), .B(n36881), .Z(n36879) );
  NANDN U37126 ( .A(n36881), .B(n36880), .Z(n36876) );
  ANDN U37127 ( .B(B[163]), .A(n80), .Z(n36660) );
  XNOR U37128 ( .A(n36668), .B(n36882), .Z(n36661) );
  XNOR U37129 ( .A(n36667), .B(n36665), .Z(n36882) );
  AND U37130 ( .A(n36883), .B(n36884), .Z(n36665) );
  NANDN U37131 ( .A(n36885), .B(n36886), .Z(n36884) );
  OR U37132 ( .A(n36887), .B(n36888), .Z(n36886) );
  NAND U37133 ( .A(n36888), .B(n36887), .Z(n36883) );
  ANDN U37134 ( .B(B[164]), .A(n81), .Z(n36667) );
  XNOR U37135 ( .A(n36675), .B(n36889), .Z(n36668) );
  XNOR U37136 ( .A(n36674), .B(n36672), .Z(n36889) );
  AND U37137 ( .A(n36890), .B(n36891), .Z(n36672) );
  NANDN U37138 ( .A(n36892), .B(n36893), .Z(n36891) );
  NAND U37139 ( .A(n36894), .B(n36895), .Z(n36893) );
  ANDN U37140 ( .B(B[165]), .A(n82), .Z(n36674) );
  XOR U37141 ( .A(n36681), .B(n36896), .Z(n36675) );
  XNOR U37142 ( .A(n36679), .B(n36682), .Z(n36896) );
  NAND U37143 ( .A(A[2]), .B(B[166]), .Z(n36682) );
  NANDN U37144 ( .A(n36897), .B(n36898), .Z(n36679) );
  AND U37145 ( .A(A[0]), .B(B[167]), .Z(n36898) );
  XNOR U37146 ( .A(n36684), .B(n36899), .Z(n36681) );
  NAND U37147 ( .A(A[0]), .B(B[168]), .Z(n36899) );
  NAND U37148 ( .A(B[167]), .B(A[1]), .Z(n36684) );
  NAND U37149 ( .A(n36900), .B(n36901), .Z(n460) );
  NANDN U37150 ( .A(n36902), .B(n36903), .Z(n36901) );
  OR U37151 ( .A(n36904), .B(n36905), .Z(n36903) );
  NAND U37152 ( .A(n36905), .B(n36904), .Z(n36900) );
  XOR U37153 ( .A(n462), .B(n461), .Z(\A1[165] ) );
  XOR U37154 ( .A(n36905), .B(n36906), .Z(n461) );
  XNOR U37155 ( .A(n36904), .B(n36902), .Z(n36906) );
  AND U37156 ( .A(n36907), .B(n36908), .Z(n36902) );
  NANDN U37157 ( .A(n36909), .B(n36910), .Z(n36908) );
  NANDN U37158 ( .A(n36911), .B(n36912), .Z(n36910) );
  NANDN U37159 ( .A(n36912), .B(n36911), .Z(n36907) );
  ANDN U37160 ( .B(B[136]), .A(n54), .Z(n36904) );
  XNOR U37161 ( .A(n36699), .B(n36913), .Z(n36905) );
  XNOR U37162 ( .A(n36698), .B(n36696), .Z(n36913) );
  AND U37163 ( .A(n36914), .B(n36915), .Z(n36696) );
  NANDN U37164 ( .A(n36916), .B(n36917), .Z(n36915) );
  OR U37165 ( .A(n36918), .B(n36919), .Z(n36917) );
  NAND U37166 ( .A(n36919), .B(n36918), .Z(n36914) );
  ANDN U37167 ( .B(B[137]), .A(n55), .Z(n36698) );
  XNOR U37168 ( .A(n36706), .B(n36920), .Z(n36699) );
  XNOR U37169 ( .A(n36705), .B(n36703), .Z(n36920) );
  AND U37170 ( .A(n36921), .B(n36922), .Z(n36703) );
  NANDN U37171 ( .A(n36923), .B(n36924), .Z(n36922) );
  NANDN U37172 ( .A(n36925), .B(n36926), .Z(n36924) );
  NANDN U37173 ( .A(n36926), .B(n36925), .Z(n36921) );
  ANDN U37174 ( .B(B[138]), .A(n56), .Z(n36705) );
  XNOR U37175 ( .A(n36713), .B(n36927), .Z(n36706) );
  XNOR U37176 ( .A(n36712), .B(n36710), .Z(n36927) );
  AND U37177 ( .A(n36928), .B(n36929), .Z(n36710) );
  NANDN U37178 ( .A(n36930), .B(n36931), .Z(n36929) );
  OR U37179 ( .A(n36932), .B(n36933), .Z(n36931) );
  NAND U37180 ( .A(n36933), .B(n36932), .Z(n36928) );
  ANDN U37181 ( .B(B[139]), .A(n57), .Z(n36712) );
  XNOR U37182 ( .A(n36720), .B(n36934), .Z(n36713) );
  XNOR U37183 ( .A(n36719), .B(n36717), .Z(n36934) );
  AND U37184 ( .A(n36935), .B(n36936), .Z(n36717) );
  NANDN U37185 ( .A(n36937), .B(n36938), .Z(n36936) );
  NANDN U37186 ( .A(n36939), .B(n36940), .Z(n36938) );
  NANDN U37187 ( .A(n36940), .B(n36939), .Z(n36935) );
  ANDN U37188 ( .B(B[140]), .A(n58), .Z(n36719) );
  XNOR U37189 ( .A(n36727), .B(n36941), .Z(n36720) );
  XNOR U37190 ( .A(n36726), .B(n36724), .Z(n36941) );
  AND U37191 ( .A(n36942), .B(n36943), .Z(n36724) );
  NANDN U37192 ( .A(n36944), .B(n36945), .Z(n36943) );
  OR U37193 ( .A(n36946), .B(n36947), .Z(n36945) );
  NAND U37194 ( .A(n36947), .B(n36946), .Z(n36942) );
  ANDN U37195 ( .B(B[141]), .A(n59), .Z(n36726) );
  XNOR U37196 ( .A(n36734), .B(n36948), .Z(n36727) );
  XNOR U37197 ( .A(n36733), .B(n36731), .Z(n36948) );
  AND U37198 ( .A(n36949), .B(n36950), .Z(n36731) );
  NANDN U37199 ( .A(n36951), .B(n36952), .Z(n36950) );
  NANDN U37200 ( .A(n36953), .B(n36954), .Z(n36952) );
  NANDN U37201 ( .A(n36954), .B(n36953), .Z(n36949) );
  ANDN U37202 ( .B(B[142]), .A(n60), .Z(n36733) );
  XNOR U37203 ( .A(n36741), .B(n36955), .Z(n36734) );
  XNOR U37204 ( .A(n36740), .B(n36738), .Z(n36955) );
  AND U37205 ( .A(n36956), .B(n36957), .Z(n36738) );
  NANDN U37206 ( .A(n36958), .B(n36959), .Z(n36957) );
  OR U37207 ( .A(n36960), .B(n36961), .Z(n36959) );
  NAND U37208 ( .A(n36961), .B(n36960), .Z(n36956) );
  ANDN U37209 ( .B(B[143]), .A(n61), .Z(n36740) );
  XNOR U37210 ( .A(n36748), .B(n36962), .Z(n36741) );
  XNOR U37211 ( .A(n36747), .B(n36745), .Z(n36962) );
  AND U37212 ( .A(n36963), .B(n36964), .Z(n36745) );
  NANDN U37213 ( .A(n36965), .B(n36966), .Z(n36964) );
  NANDN U37214 ( .A(n36967), .B(n36968), .Z(n36966) );
  NANDN U37215 ( .A(n36968), .B(n36967), .Z(n36963) );
  ANDN U37216 ( .B(B[144]), .A(n62), .Z(n36747) );
  XNOR U37217 ( .A(n36755), .B(n36969), .Z(n36748) );
  XNOR U37218 ( .A(n36754), .B(n36752), .Z(n36969) );
  AND U37219 ( .A(n36970), .B(n36971), .Z(n36752) );
  NANDN U37220 ( .A(n36972), .B(n36973), .Z(n36971) );
  OR U37221 ( .A(n36974), .B(n36975), .Z(n36973) );
  NAND U37222 ( .A(n36975), .B(n36974), .Z(n36970) );
  ANDN U37223 ( .B(B[145]), .A(n63), .Z(n36754) );
  XNOR U37224 ( .A(n36762), .B(n36976), .Z(n36755) );
  XNOR U37225 ( .A(n36761), .B(n36759), .Z(n36976) );
  AND U37226 ( .A(n36977), .B(n36978), .Z(n36759) );
  NANDN U37227 ( .A(n36979), .B(n36980), .Z(n36978) );
  NANDN U37228 ( .A(n36981), .B(n36982), .Z(n36980) );
  NANDN U37229 ( .A(n36982), .B(n36981), .Z(n36977) );
  ANDN U37230 ( .B(B[146]), .A(n64), .Z(n36761) );
  XNOR U37231 ( .A(n36769), .B(n36983), .Z(n36762) );
  XNOR U37232 ( .A(n36768), .B(n36766), .Z(n36983) );
  AND U37233 ( .A(n36984), .B(n36985), .Z(n36766) );
  NANDN U37234 ( .A(n36986), .B(n36987), .Z(n36985) );
  OR U37235 ( .A(n36988), .B(n36989), .Z(n36987) );
  NAND U37236 ( .A(n36989), .B(n36988), .Z(n36984) );
  ANDN U37237 ( .B(B[147]), .A(n65), .Z(n36768) );
  XNOR U37238 ( .A(n36776), .B(n36990), .Z(n36769) );
  XNOR U37239 ( .A(n36775), .B(n36773), .Z(n36990) );
  AND U37240 ( .A(n36991), .B(n36992), .Z(n36773) );
  NANDN U37241 ( .A(n36993), .B(n36994), .Z(n36992) );
  NANDN U37242 ( .A(n36995), .B(n36996), .Z(n36994) );
  NANDN U37243 ( .A(n36996), .B(n36995), .Z(n36991) );
  ANDN U37244 ( .B(B[148]), .A(n66), .Z(n36775) );
  XNOR U37245 ( .A(n36783), .B(n36997), .Z(n36776) );
  XNOR U37246 ( .A(n36782), .B(n36780), .Z(n36997) );
  AND U37247 ( .A(n36998), .B(n36999), .Z(n36780) );
  NANDN U37248 ( .A(n37000), .B(n37001), .Z(n36999) );
  OR U37249 ( .A(n37002), .B(n37003), .Z(n37001) );
  NAND U37250 ( .A(n37003), .B(n37002), .Z(n36998) );
  ANDN U37251 ( .B(B[149]), .A(n67), .Z(n36782) );
  XNOR U37252 ( .A(n36790), .B(n37004), .Z(n36783) );
  XNOR U37253 ( .A(n36789), .B(n36787), .Z(n37004) );
  AND U37254 ( .A(n37005), .B(n37006), .Z(n36787) );
  NANDN U37255 ( .A(n37007), .B(n37008), .Z(n37006) );
  NANDN U37256 ( .A(n37009), .B(n37010), .Z(n37008) );
  NANDN U37257 ( .A(n37010), .B(n37009), .Z(n37005) );
  ANDN U37258 ( .B(B[150]), .A(n68), .Z(n36789) );
  XNOR U37259 ( .A(n36797), .B(n37011), .Z(n36790) );
  XNOR U37260 ( .A(n36796), .B(n36794), .Z(n37011) );
  AND U37261 ( .A(n37012), .B(n37013), .Z(n36794) );
  NANDN U37262 ( .A(n37014), .B(n37015), .Z(n37013) );
  OR U37263 ( .A(n37016), .B(n37017), .Z(n37015) );
  NAND U37264 ( .A(n37017), .B(n37016), .Z(n37012) );
  ANDN U37265 ( .B(B[151]), .A(n69), .Z(n36796) );
  XNOR U37266 ( .A(n36804), .B(n37018), .Z(n36797) );
  XNOR U37267 ( .A(n36803), .B(n36801), .Z(n37018) );
  AND U37268 ( .A(n37019), .B(n37020), .Z(n36801) );
  NANDN U37269 ( .A(n37021), .B(n37022), .Z(n37020) );
  NANDN U37270 ( .A(n37023), .B(n37024), .Z(n37022) );
  NANDN U37271 ( .A(n37024), .B(n37023), .Z(n37019) );
  ANDN U37272 ( .B(B[152]), .A(n70), .Z(n36803) );
  XNOR U37273 ( .A(n36811), .B(n37025), .Z(n36804) );
  XNOR U37274 ( .A(n36810), .B(n36808), .Z(n37025) );
  AND U37275 ( .A(n37026), .B(n37027), .Z(n36808) );
  NANDN U37276 ( .A(n37028), .B(n37029), .Z(n37027) );
  OR U37277 ( .A(n37030), .B(n37031), .Z(n37029) );
  NAND U37278 ( .A(n37031), .B(n37030), .Z(n37026) );
  ANDN U37279 ( .B(B[153]), .A(n71), .Z(n36810) );
  XNOR U37280 ( .A(n36818), .B(n37032), .Z(n36811) );
  XNOR U37281 ( .A(n36817), .B(n36815), .Z(n37032) );
  AND U37282 ( .A(n37033), .B(n37034), .Z(n36815) );
  NANDN U37283 ( .A(n37035), .B(n37036), .Z(n37034) );
  NANDN U37284 ( .A(n37037), .B(n37038), .Z(n37036) );
  NANDN U37285 ( .A(n37038), .B(n37037), .Z(n37033) );
  ANDN U37286 ( .B(B[154]), .A(n72), .Z(n36817) );
  XNOR U37287 ( .A(n36825), .B(n37039), .Z(n36818) );
  XNOR U37288 ( .A(n36824), .B(n36822), .Z(n37039) );
  AND U37289 ( .A(n37040), .B(n37041), .Z(n36822) );
  NANDN U37290 ( .A(n37042), .B(n37043), .Z(n37041) );
  OR U37291 ( .A(n37044), .B(n37045), .Z(n37043) );
  NAND U37292 ( .A(n37045), .B(n37044), .Z(n37040) );
  ANDN U37293 ( .B(B[155]), .A(n73), .Z(n36824) );
  XNOR U37294 ( .A(n36832), .B(n37046), .Z(n36825) );
  XNOR U37295 ( .A(n36831), .B(n36829), .Z(n37046) );
  AND U37296 ( .A(n37047), .B(n37048), .Z(n36829) );
  NANDN U37297 ( .A(n37049), .B(n37050), .Z(n37048) );
  NANDN U37298 ( .A(n37051), .B(n37052), .Z(n37050) );
  NANDN U37299 ( .A(n37052), .B(n37051), .Z(n37047) );
  ANDN U37300 ( .B(B[156]), .A(n74), .Z(n36831) );
  XNOR U37301 ( .A(n36839), .B(n37053), .Z(n36832) );
  XNOR U37302 ( .A(n36838), .B(n36836), .Z(n37053) );
  AND U37303 ( .A(n37054), .B(n37055), .Z(n36836) );
  NANDN U37304 ( .A(n37056), .B(n37057), .Z(n37055) );
  OR U37305 ( .A(n37058), .B(n37059), .Z(n37057) );
  NAND U37306 ( .A(n37059), .B(n37058), .Z(n37054) );
  ANDN U37307 ( .B(B[157]), .A(n75), .Z(n36838) );
  XNOR U37308 ( .A(n36846), .B(n37060), .Z(n36839) );
  XNOR U37309 ( .A(n36845), .B(n36843), .Z(n37060) );
  AND U37310 ( .A(n37061), .B(n37062), .Z(n36843) );
  NANDN U37311 ( .A(n37063), .B(n37064), .Z(n37062) );
  NANDN U37312 ( .A(n37065), .B(n37066), .Z(n37064) );
  NANDN U37313 ( .A(n37066), .B(n37065), .Z(n37061) );
  ANDN U37314 ( .B(B[158]), .A(n76), .Z(n36845) );
  XNOR U37315 ( .A(n36853), .B(n37067), .Z(n36846) );
  XNOR U37316 ( .A(n36852), .B(n36850), .Z(n37067) );
  AND U37317 ( .A(n37068), .B(n37069), .Z(n36850) );
  NANDN U37318 ( .A(n37070), .B(n37071), .Z(n37069) );
  OR U37319 ( .A(n37072), .B(n37073), .Z(n37071) );
  NAND U37320 ( .A(n37073), .B(n37072), .Z(n37068) );
  ANDN U37321 ( .B(B[159]), .A(n77), .Z(n36852) );
  XNOR U37322 ( .A(n36860), .B(n37074), .Z(n36853) );
  XNOR U37323 ( .A(n36859), .B(n36857), .Z(n37074) );
  AND U37324 ( .A(n37075), .B(n37076), .Z(n36857) );
  NANDN U37325 ( .A(n37077), .B(n37078), .Z(n37076) );
  NANDN U37326 ( .A(n37079), .B(n37080), .Z(n37078) );
  NANDN U37327 ( .A(n37080), .B(n37079), .Z(n37075) );
  ANDN U37328 ( .B(B[160]), .A(n78), .Z(n36859) );
  XNOR U37329 ( .A(n36867), .B(n37081), .Z(n36860) );
  XNOR U37330 ( .A(n36866), .B(n36864), .Z(n37081) );
  AND U37331 ( .A(n37082), .B(n37083), .Z(n36864) );
  NANDN U37332 ( .A(n37084), .B(n37085), .Z(n37083) );
  OR U37333 ( .A(n37086), .B(n37087), .Z(n37085) );
  NAND U37334 ( .A(n37087), .B(n37086), .Z(n37082) );
  ANDN U37335 ( .B(B[161]), .A(n79), .Z(n36866) );
  XNOR U37336 ( .A(n36874), .B(n37088), .Z(n36867) );
  XNOR U37337 ( .A(n36873), .B(n36871), .Z(n37088) );
  AND U37338 ( .A(n37089), .B(n37090), .Z(n36871) );
  NANDN U37339 ( .A(n37091), .B(n37092), .Z(n37090) );
  NANDN U37340 ( .A(n37093), .B(n37094), .Z(n37092) );
  NANDN U37341 ( .A(n37094), .B(n37093), .Z(n37089) );
  ANDN U37342 ( .B(B[162]), .A(n80), .Z(n36873) );
  XNOR U37343 ( .A(n36881), .B(n37095), .Z(n36874) );
  XNOR U37344 ( .A(n36880), .B(n36878), .Z(n37095) );
  AND U37345 ( .A(n37096), .B(n37097), .Z(n36878) );
  NANDN U37346 ( .A(n37098), .B(n37099), .Z(n37097) );
  OR U37347 ( .A(n37100), .B(n37101), .Z(n37099) );
  NAND U37348 ( .A(n37101), .B(n37100), .Z(n37096) );
  ANDN U37349 ( .B(B[163]), .A(n81), .Z(n36880) );
  XNOR U37350 ( .A(n36888), .B(n37102), .Z(n36881) );
  XNOR U37351 ( .A(n36887), .B(n36885), .Z(n37102) );
  AND U37352 ( .A(n37103), .B(n37104), .Z(n36885) );
  NANDN U37353 ( .A(n37105), .B(n37106), .Z(n37104) );
  NAND U37354 ( .A(n37107), .B(n37108), .Z(n37106) );
  ANDN U37355 ( .B(B[164]), .A(n82), .Z(n36887) );
  XOR U37356 ( .A(n36894), .B(n37109), .Z(n36888) );
  XNOR U37357 ( .A(n36892), .B(n36895), .Z(n37109) );
  NAND U37358 ( .A(A[2]), .B(B[165]), .Z(n36895) );
  NANDN U37359 ( .A(n37110), .B(n37111), .Z(n36892) );
  AND U37360 ( .A(A[0]), .B(B[166]), .Z(n37111) );
  XNOR U37361 ( .A(n36897), .B(n37112), .Z(n36894) );
  NAND U37362 ( .A(A[0]), .B(B[167]), .Z(n37112) );
  NAND U37363 ( .A(B[166]), .B(A[1]), .Z(n36897) );
  NAND U37364 ( .A(n37113), .B(n37114), .Z(n462) );
  NANDN U37365 ( .A(n37115), .B(n37116), .Z(n37114) );
  OR U37366 ( .A(n37117), .B(n37118), .Z(n37116) );
  NAND U37367 ( .A(n37118), .B(n37117), .Z(n37113) );
  XOR U37368 ( .A(n464), .B(n463), .Z(\A1[164] ) );
  XOR U37369 ( .A(n37118), .B(n37119), .Z(n463) );
  XNOR U37370 ( .A(n37117), .B(n37115), .Z(n37119) );
  AND U37371 ( .A(n37120), .B(n37121), .Z(n37115) );
  NANDN U37372 ( .A(n37122), .B(n37123), .Z(n37121) );
  NANDN U37373 ( .A(n37124), .B(n37125), .Z(n37123) );
  NANDN U37374 ( .A(n37125), .B(n37124), .Z(n37120) );
  ANDN U37375 ( .B(B[135]), .A(n54), .Z(n37117) );
  XNOR U37376 ( .A(n36912), .B(n37126), .Z(n37118) );
  XNOR U37377 ( .A(n36911), .B(n36909), .Z(n37126) );
  AND U37378 ( .A(n37127), .B(n37128), .Z(n36909) );
  NANDN U37379 ( .A(n37129), .B(n37130), .Z(n37128) );
  OR U37380 ( .A(n37131), .B(n37132), .Z(n37130) );
  NAND U37381 ( .A(n37132), .B(n37131), .Z(n37127) );
  ANDN U37382 ( .B(B[136]), .A(n55), .Z(n36911) );
  XNOR U37383 ( .A(n36919), .B(n37133), .Z(n36912) );
  XNOR U37384 ( .A(n36918), .B(n36916), .Z(n37133) );
  AND U37385 ( .A(n37134), .B(n37135), .Z(n36916) );
  NANDN U37386 ( .A(n37136), .B(n37137), .Z(n37135) );
  NANDN U37387 ( .A(n37138), .B(n37139), .Z(n37137) );
  NANDN U37388 ( .A(n37139), .B(n37138), .Z(n37134) );
  ANDN U37389 ( .B(B[137]), .A(n56), .Z(n36918) );
  XNOR U37390 ( .A(n36926), .B(n37140), .Z(n36919) );
  XNOR U37391 ( .A(n36925), .B(n36923), .Z(n37140) );
  AND U37392 ( .A(n37141), .B(n37142), .Z(n36923) );
  NANDN U37393 ( .A(n37143), .B(n37144), .Z(n37142) );
  OR U37394 ( .A(n37145), .B(n37146), .Z(n37144) );
  NAND U37395 ( .A(n37146), .B(n37145), .Z(n37141) );
  ANDN U37396 ( .B(B[138]), .A(n57), .Z(n36925) );
  XNOR U37397 ( .A(n36933), .B(n37147), .Z(n36926) );
  XNOR U37398 ( .A(n36932), .B(n36930), .Z(n37147) );
  AND U37399 ( .A(n37148), .B(n37149), .Z(n36930) );
  NANDN U37400 ( .A(n37150), .B(n37151), .Z(n37149) );
  NANDN U37401 ( .A(n37152), .B(n37153), .Z(n37151) );
  NANDN U37402 ( .A(n37153), .B(n37152), .Z(n37148) );
  ANDN U37403 ( .B(B[139]), .A(n58), .Z(n36932) );
  XNOR U37404 ( .A(n36940), .B(n37154), .Z(n36933) );
  XNOR U37405 ( .A(n36939), .B(n36937), .Z(n37154) );
  AND U37406 ( .A(n37155), .B(n37156), .Z(n36937) );
  NANDN U37407 ( .A(n37157), .B(n37158), .Z(n37156) );
  OR U37408 ( .A(n37159), .B(n37160), .Z(n37158) );
  NAND U37409 ( .A(n37160), .B(n37159), .Z(n37155) );
  ANDN U37410 ( .B(B[140]), .A(n59), .Z(n36939) );
  XNOR U37411 ( .A(n36947), .B(n37161), .Z(n36940) );
  XNOR U37412 ( .A(n36946), .B(n36944), .Z(n37161) );
  AND U37413 ( .A(n37162), .B(n37163), .Z(n36944) );
  NANDN U37414 ( .A(n37164), .B(n37165), .Z(n37163) );
  NANDN U37415 ( .A(n37166), .B(n37167), .Z(n37165) );
  NANDN U37416 ( .A(n37167), .B(n37166), .Z(n37162) );
  ANDN U37417 ( .B(B[141]), .A(n60), .Z(n36946) );
  XNOR U37418 ( .A(n36954), .B(n37168), .Z(n36947) );
  XNOR U37419 ( .A(n36953), .B(n36951), .Z(n37168) );
  AND U37420 ( .A(n37169), .B(n37170), .Z(n36951) );
  NANDN U37421 ( .A(n37171), .B(n37172), .Z(n37170) );
  OR U37422 ( .A(n37173), .B(n37174), .Z(n37172) );
  NAND U37423 ( .A(n37174), .B(n37173), .Z(n37169) );
  ANDN U37424 ( .B(B[142]), .A(n61), .Z(n36953) );
  XNOR U37425 ( .A(n36961), .B(n37175), .Z(n36954) );
  XNOR U37426 ( .A(n36960), .B(n36958), .Z(n37175) );
  AND U37427 ( .A(n37176), .B(n37177), .Z(n36958) );
  NANDN U37428 ( .A(n37178), .B(n37179), .Z(n37177) );
  NANDN U37429 ( .A(n37180), .B(n37181), .Z(n37179) );
  NANDN U37430 ( .A(n37181), .B(n37180), .Z(n37176) );
  ANDN U37431 ( .B(B[143]), .A(n62), .Z(n36960) );
  XNOR U37432 ( .A(n36968), .B(n37182), .Z(n36961) );
  XNOR U37433 ( .A(n36967), .B(n36965), .Z(n37182) );
  AND U37434 ( .A(n37183), .B(n37184), .Z(n36965) );
  NANDN U37435 ( .A(n37185), .B(n37186), .Z(n37184) );
  OR U37436 ( .A(n37187), .B(n37188), .Z(n37186) );
  NAND U37437 ( .A(n37188), .B(n37187), .Z(n37183) );
  ANDN U37438 ( .B(B[144]), .A(n63), .Z(n36967) );
  XNOR U37439 ( .A(n36975), .B(n37189), .Z(n36968) );
  XNOR U37440 ( .A(n36974), .B(n36972), .Z(n37189) );
  AND U37441 ( .A(n37190), .B(n37191), .Z(n36972) );
  NANDN U37442 ( .A(n37192), .B(n37193), .Z(n37191) );
  NANDN U37443 ( .A(n37194), .B(n37195), .Z(n37193) );
  NANDN U37444 ( .A(n37195), .B(n37194), .Z(n37190) );
  ANDN U37445 ( .B(B[145]), .A(n64), .Z(n36974) );
  XNOR U37446 ( .A(n36982), .B(n37196), .Z(n36975) );
  XNOR U37447 ( .A(n36981), .B(n36979), .Z(n37196) );
  AND U37448 ( .A(n37197), .B(n37198), .Z(n36979) );
  NANDN U37449 ( .A(n37199), .B(n37200), .Z(n37198) );
  OR U37450 ( .A(n37201), .B(n37202), .Z(n37200) );
  NAND U37451 ( .A(n37202), .B(n37201), .Z(n37197) );
  ANDN U37452 ( .B(B[146]), .A(n65), .Z(n36981) );
  XNOR U37453 ( .A(n36989), .B(n37203), .Z(n36982) );
  XNOR U37454 ( .A(n36988), .B(n36986), .Z(n37203) );
  AND U37455 ( .A(n37204), .B(n37205), .Z(n36986) );
  NANDN U37456 ( .A(n37206), .B(n37207), .Z(n37205) );
  NANDN U37457 ( .A(n37208), .B(n37209), .Z(n37207) );
  NANDN U37458 ( .A(n37209), .B(n37208), .Z(n37204) );
  ANDN U37459 ( .B(B[147]), .A(n66), .Z(n36988) );
  XNOR U37460 ( .A(n36996), .B(n37210), .Z(n36989) );
  XNOR U37461 ( .A(n36995), .B(n36993), .Z(n37210) );
  AND U37462 ( .A(n37211), .B(n37212), .Z(n36993) );
  NANDN U37463 ( .A(n37213), .B(n37214), .Z(n37212) );
  OR U37464 ( .A(n37215), .B(n37216), .Z(n37214) );
  NAND U37465 ( .A(n37216), .B(n37215), .Z(n37211) );
  ANDN U37466 ( .B(B[148]), .A(n67), .Z(n36995) );
  XNOR U37467 ( .A(n37003), .B(n37217), .Z(n36996) );
  XNOR U37468 ( .A(n37002), .B(n37000), .Z(n37217) );
  AND U37469 ( .A(n37218), .B(n37219), .Z(n37000) );
  NANDN U37470 ( .A(n37220), .B(n37221), .Z(n37219) );
  NANDN U37471 ( .A(n37222), .B(n37223), .Z(n37221) );
  NANDN U37472 ( .A(n37223), .B(n37222), .Z(n37218) );
  ANDN U37473 ( .B(B[149]), .A(n68), .Z(n37002) );
  XNOR U37474 ( .A(n37010), .B(n37224), .Z(n37003) );
  XNOR U37475 ( .A(n37009), .B(n37007), .Z(n37224) );
  AND U37476 ( .A(n37225), .B(n37226), .Z(n37007) );
  NANDN U37477 ( .A(n37227), .B(n37228), .Z(n37226) );
  OR U37478 ( .A(n37229), .B(n37230), .Z(n37228) );
  NAND U37479 ( .A(n37230), .B(n37229), .Z(n37225) );
  ANDN U37480 ( .B(B[150]), .A(n69), .Z(n37009) );
  XNOR U37481 ( .A(n37017), .B(n37231), .Z(n37010) );
  XNOR U37482 ( .A(n37016), .B(n37014), .Z(n37231) );
  AND U37483 ( .A(n37232), .B(n37233), .Z(n37014) );
  NANDN U37484 ( .A(n37234), .B(n37235), .Z(n37233) );
  NANDN U37485 ( .A(n37236), .B(n37237), .Z(n37235) );
  NANDN U37486 ( .A(n37237), .B(n37236), .Z(n37232) );
  ANDN U37487 ( .B(B[151]), .A(n70), .Z(n37016) );
  XNOR U37488 ( .A(n37024), .B(n37238), .Z(n37017) );
  XNOR U37489 ( .A(n37023), .B(n37021), .Z(n37238) );
  AND U37490 ( .A(n37239), .B(n37240), .Z(n37021) );
  NANDN U37491 ( .A(n37241), .B(n37242), .Z(n37240) );
  OR U37492 ( .A(n37243), .B(n37244), .Z(n37242) );
  NAND U37493 ( .A(n37244), .B(n37243), .Z(n37239) );
  ANDN U37494 ( .B(B[152]), .A(n71), .Z(n37023) );
  XNOR U37495 ( .A(n37031), .B(n37245), .Z(n37024) );
  XNOR U37496 ( .A(n37030), .B(n37028), .Z(n37245) );
  AND U37497 ( .A(n37246), .B(n37247), .Z(n37028) );
  NANDN U37498 ( .A(n37248), .B(n37249), .Z(n37247) );
  NANDN U37499 ( .A(n37250), .B(n37251), .Z(n37249) );
  NANDN U37500 ( .A(n37251), .B(n37250), .Z(n37246) );
  ANDN U37501 ( .B(B[153]), .A(n72), .Z(n37030) );
  XNOR U37502 ( .A(n37038), .B(n37252), .Z(n37031) );
  XNOR U37503 ( .A(n37037), .B(n37035), .Z(n37252) );
  AND U37504 ( .A(n37253), .B(n37254), .Z(n37035) );
  NANDN U37505 ( .A(n37255), .B(n37256), .Z(n37254) );
  OR U37506 ( .A(n37257), .B(n37258), .Z(n37256) );
  NAND U37507 ( .A(n37258), .B(n37257), .Z(n37253) );
  ANDN U37508 ( .B(B[154]), .A(n73), .Z(n37037) );
  XNOR U37509 ( .A(n37045), .B(n37259), .Z(n37038) );
  XNOR U37510 ( .A(n37044), .B(n37042), .Z(n37259) );
  AND U37511 ( .A(n37260), .B(n37261), .Z(n37042) );
  NANDN U37512 ( .A(n37262), .B(n37263), .Z(n37261) );
  NANDN U37513 ( .A(n37264), .B(n37265), .Z(n37263) );
  NANDN U37514 ( .A(n37265), .B(n37264), .Z(n37260) );
  ANDN U37515 ( .B(B[155]), .A(n74), .Z(n37044) );
  XNOR U37516 ( .A(n37052), .B(n37266), .Z(n37045) );
  XNOR U37517 ( .A(n37051), .B(n37049), .Z(n37266) );
  AND U37518 ( .A(n37267), .B(n37268), .Z(n37049) );
  NANDN U37519 ( .A(n37269), .B(n37270), .Z(n37268) );
  OR U37520 ( .A(n37271), .B(n37272), .Z(n37270) );
  NAND U37521 ( .A(n37272), .B(n37271), .Z(n37267) );
  ANDN U37522 ( .B(B[156]), .A(n75), .Z(n37051) );
  XNOR U37523 ( .A(n37059), .B(n37273), .Z(n37052) );
  XNOR U37524 ( .A(n37058), .B(n37056), .Z(n37273) );
  AND U37525 ( .A(n37274), .B(n37275), .Z(n37056) );
  NANDN U37526 ( .A(n37276), .B(n37277), .Z(n37275) );
  NANDN U37527 ( .A(n37278), .B(n37279), .Z(n37277) );
  NANDN U37528 ( .A(n37279), .B(n37278), .Z(n37274) );
  ANDN U37529 ( .B(B[157]), .A(n76), .Z(n37058) );
  XNOR U37530 ( .A(n37066), .B(n37280), .Z(n37059) );
  XNOR U37531 ( .A(n37065), .B(n37063), .Z(n37280) );
  AND U37532 ( .A(n37281), .B(n37282), .Z(n37063) );
  NANDN U37533 ( .A(n37283), .B(n37284), .Z(n37282) );
  OR U37534 ( .A(n37285), .B(n37286), .Z(n37284) );
  NAND U37535 ( .A(n37286), .B(n37285), .Z(n37281) );
  ANDN U37536 ( .B(B[158]), .A(n77), .Z(n37065) );
  XNOR U37537 ( .A(n37073), .B(n37287), .Z(n37066) );
  XNOR U37538 ( .A(n37072), .B(n37070), .Z(n37287) );
  AND U37539 ( .A(n37288), .B(n37289), .Z(n37070) );
  NANDN U37540 ( .A(n37290), .B(n37291), .Z(n37289) );
  NANDN U37541 ( .A(n37292), .B(n37293), .Z(n37291) );
  NANDN U37542 ( .A(n37293), .B(n37292), .Z(n37288) );
  ANDN U37543 ( .B(B[159]), .A(n78), .Z(n37072) );
  XNOR U37544 ( .A(n37080), .B(n37294), .Z(n37073) );
  XNOR U37545 ( .A(n37079), .B(n37077), .Z(n37294) );
  AND U37546 ( .A(n37295), .B(n37296), .Z(n37077) );
  NANDN U37547 ( .A(n37297), .B(n37298), .Z(n37296) );
  OR U37548 ( .A(n37299), .B(n37300), .Z(n37298) );
  NAND U37549 ( .A(n37300), .B(n37299), .Z(n37295) );
  ANDN U37550 ( .B(B[160]), .A(n79), .Z(n37079) );
  XNOR U37551 ( .A(n37087), .B(n37301), .Z(n37080) );
  XNOR U37552 ( .A(n37086), .B(n37084), .Z(n37301) );
  AND U37553 ( .A(n37302), .B(n37303), .Z(n37084) );
  NANDN U37554 ( .A(n37304), .B(n37305), .Z(n37303) );
  NANDN U37555 ( .A(n37306), .B(n37307), .Z(n37305) );
  NANDN U37556 ( .A(n37307), .B(n37306), .Z(n37302) );
  ANDN U37557 ( .B(B[161]), .A(n80), .Z(n37086) );
  XNOR U37558 ( .A(n37094), .B(n37308), .Z(n37087) );
  XNOR U37559 ( .A(n37093), .B(n37091), .Z(n37308) );
  AND U37560 ( .A(n37309), .B(n37310), .Z(n37091) );
  NANDN U37561 ( .A(n37311), .B(n37312), .Z(n37310) );
  OR U37562 ( .A(n37313), .B(n37314), .Z(n37312) );
  NAND U37563 ( .A(n37314), .B(n37313), .Z(n37309) );
  ANDN U37564 ( .B(B[162]), .A(n81), .Z(n37093) );
  XNOR U37565 ( .A(n37101), .B(n37315), .Z(n37094) );
  XNOR U37566 ( .A(n37100), .B(n37098), .Z(n37315) );
  AND U37567 ( .A(n37316), .B(n37317), .Z(n37098) );
  NANDN U37568 ( .A(n37318), .B(n37319), .Z(n37317) );
  NAND U37569 ( .A(n37320), .B(n37321), .Z(n37319) );
  ANDN U37570 ( .B(B[163]), .A(n82), .Z(n37100) );
  XOR U37571 ( .A(n37107), .B(n37322), .Z(n37101) );
  XNOR U37572 ( .A(n37105), .B(n37108), .Z(n37322) );
  NAND U37573 ( .A(A[2]), .B(B[164]), .Z(n37108) );
  NANDN U37574 ( .A(n37323), .B(n37324), .Z(n37105) );
  AND U37575 ( .A(A[0]), .B(B[165]), .Z(n37324) );
  XNOR U37576 ( .A(n37110), .B(n37325), .Z(n37107) );
  NAND U37577 ( .A(A[0]), .B(B[166]), .Z(n37325) );
  NAND U37578 ( .A(B[165]), .B(A[1]), .Z(n37110) );
  NAND U37579 ( .A(n37326), .B(n37327), .Z(n464) );
  NANDN U37580 ( .A(n37328), .B(n37329), .Z(n37327) );
  OR U37581 ( .A(n37330), .B(n37331), .Z(n37329) );
  NAND U37582 ( .A(n37331), .B(n37330), .Z(n37326) );
  XOR U37583 ( .A(n466), .B(n465), .Z(\A1[163] ) );
  XOR U37584 ( .A(n37331), .B(n37332), .Z(n465) );
  XNOR U37585 ( .A(n37330), .B(n37328), .Z(n37332) );
  AND U37586 ( .A(n37333), .B(n37334), .Z(n37328) );
  NANDN U37587 ( .A(n37335), .B(n37336), .Z(n37334) );
  NANDN U37588 ( .A(n37337), .B(n37338), .Z(n37336) );
  NANDN U37589 ( .A(n37338), .B(n37337), .Z(n37333) );
  ANDN U37590 ( .B(B[134]), .A(n54), .Z(n37330) );
  XNOR U37591 ( .A(n37125), .B(n37339), .Z(n37331) );
  XNOR U37592 ( .A(n37124), .B(n37122), .Z(n37339) );
  AND U37593 ( .A(n37340), .B(n37341), .Z(n37122) );
  NANDN U37594 ( .A(n37342), .B(n37343), .Z(n37341) );
  OR U37595 ( .A(n37344), .B(n37345), .Z(n37343) );
  NAND U37596 ( .A(n37345), .B(n37344), .Z(n37340) );
  ANDN U37597 ( .B(B[135]), .A(n55), .Z(n37124) );
  XNOR U37598 ( .A(n37132), .B(n37346), .Z(n37125) );
  XNOR U37599 ( .A(n37131), .B(n37129), .Z(n37346) );
  AND U37600 ( .A(n37347), .B(n37348), .Z(n37129) );
  NANDN U37601 ( .A(n37349), .B(n37350), .Z(n37348) );
  NANDN U37602 ( .A(n37351), .B(n37352), .Z(n37350) );
  NANDN U37603 ( .A(n37352), .B(n37351), .Z(n37347) );
  ANDN U37604 ( .B(B[136]), .A(n56), .Z(n37131) );
  XNOR U37605 ( .A(n37139), .B(n37353), .Z(n37132) );
  XNOR U37606 ( .A(n37138), .B(n37136), .Z(n37353) );
  AND U37607 ( .A(n37354), .B(n37355), .Z(n37136) );
  NANDN U37608 ( .A(n37356), .B(n37357), .Z(n37355) );
  OR U37609 ( .A(n37358), .B(n37359), .Z(n37357) );
  NAND U37610 ( .A(n37359), .B(n37358), .Z(n37354) );
  ANDN U37611 ( .B(B[137]), .A(n57), .Z(n37138) );
  XNOR U37612 ( .A(n37146), .B(n37360), .Z(n37139) );
  XNOR U37613 ( .A(n37145), .B(n37143), .Z(n37360) );
  AND U37614 ( .A(n37361), .B(n37362), .Z(n37143) );
  NANDN U37615 ( .A(n37363), .B(n37364), .Z(n37362) );
  NANDN U37616 ( .A(n37365), .B(n37366), .Z(n37364) );
  NANDN U37617 ( .A(n37366), .B(n37365), .Z(n37361) );
  ANDN U37618 ( .B(B[138]), .A(n58), .Z(n37145) );
  XNOR U37619 ( .A(n37153), .B(n37367), .Z(n37146) );
  XNOR U37620 ( .A(n37152), .B(n37150), .Z(n37367) );
  AND U37621 ( .A(n37368), .B(n37369), .Z(n37150) );
  NANDN U37622 ( .A(n37370), .B(n37371), .Z(n37369) );
  OR U37623 ( .A(n37372), .B(n37373), .Z(n37371) );
  NAND U37624 ( .A(n37373), .B(n37372), .Z(n37368) );
  ANDN U37625 ( .B(B[139]), .A(n59), .Z(n37152) );
  XNOR U37626 ( .A(n37160), .B(n37374), .Z(n37153) );
  XNOR U37627 ( .A(n37159), .B(n37157), .Z(n37374) );
  AND U37628 ( .A(n37375), .B(n37376), .Z(n37157) );
  NANDN U37629 ( .A(n37377), .B(n37378), .Z(n37376) );
  NANDN U37630 ( .A(n37379), .B(n37380), .Z(n37378) );
  NANDN U37631 ( .A(n37380), .B(n37379), .Z(n37375) );
  ANDN U37632 ( .B(B[140]), .A(n60), .Z(n37159) );
  XNOR U37633 ( .A(n37167), .B(n37381), .Z(n37160) );
  XNOR U37634 ( .A(n37166), .B(n37164), .Z(n37381) );
  AND U37635 ( .A(n37382), .B(n37383), .Z(n37164) );
  NANDN U37636 ( .A(n37384), .B(n37385), .Z(n37383) );
  OR U37637 ( .A(n37386), .B(n37387), .Z(n37385) );
  NAND U37638 ( .A(n37387), .B(n37386), .Z(n37382) );
  ANDN U37639 ( .B(B[141]), .A(n61), .Z(n37166) );
  XNOR U37640 ( .A(n37174), .B(n37388), .Z(n37167) );
  XNOR U37641 ( .A(n37173), .B(n37171), .Z(n37388) );
  AND U37642 ( .A(n37389), .B(n37390), .Z(n37171) );
  NANDN U37643 ( .A(n37391), .B(n37392), .Z(n37390) );
  NANDN U37644 ( .A(n37393), .B(n37394), .Z(n37392) );
  NANDN U37645 ( .A(n37394), .B(n37393), .Z(n37389) );
  ANDN U37646 ( .B(B[142]), .A(n62), .Z(n37173) );
  XNOR U37647 ( .A(n37181), .B(n37395), .Z(n37174) );
  XNOR U37648 ( .A(n37180), .B(n37178), .Z(n37395) );
  AND U37649 ( .A(n37396), .B(n37397), .Z(n37178) );
  NANDN U37650 ( .A(n37398), .B(n37399), .Z(n37397) );
  OR U37651 ( .A(n37400), .B(n37401), .Z(n37399) );
  NAND U37652 ( .A(n37401), .B(n37400), .Z(n37396) );
  ANDN U37653 ( .B(B[143]), .A(n63), .Z(n37180) );
  XNOR U37654 ( .A(n37188), .B(n37402), .Z(n37181) );
  XNOR U37655 ( .A(n37187), .B(n37185), .Z(n37402) );
  AND U37656 ( .A(n37403), .B(n37404), .Z(n37185) );
  NANDN U37657 ( .A(n37405), .B(n37406), .Z(n37404) );
  NANDN U37658 ( .A(n37407), .B(n37408), .Z(n37406) );
  NANDN U37659 ( .A(n37408), .B(n37407), .Z(n37403) );
  ANDN U37660 ( .B(B[144]), .A(n64), .Z(n37187) );
  XNOR U37661 ( .A(n37195), .B(n37409), .Z(n37188) );
  XNOR U37662 ( .A(n37194), .B(n37192), .Z(n37409) );
  AND U37663 ( .A(n37410), .B(n37411), .Z(n37192) );
  NANDN U37664 ( .A(n37412), .B(n37413), .Z(n37411) );
  OR U37665 ( .A(n37414), .B(n37415), .Z(n37413) );
  NAND U37666 ( .A(n37415), .B(n37414), .Z(n37410) );
  ANDN U37667 ( .B(B[145]), .A(n65), .Z(n37194) );
  XNOR U37668 ( .A(n37202), .B(n37416), .Z(n37195) );
  XNOR U37669 ( .A(n37201), .B(n37199), .Z(n37416) );
  AND U37670 ( .A(n37417), .B(n37418), .Z(n37199) );
  NANDN U37671 ( .A(n37419), .B(n37420), .Z(n37418) );
  NANDN U37672 ( .A(n37421), .B(n37422), .Z(n37420) );
  NANDN U37673 ( .A(n37422), .B(n37421), .Z(n37417) );
  ANDN U37674 ( .B(B[146]), .A(n66), .Z(n37201) );
  XNOR U37675 ( .A(n37209), .B(n37423), .Z(n37202) );
  XNOR U37676 ( .A(n37208), .B(n37206), .Z(n37423) );
  AND U37677 ( .A(n37424), .B(n37425), .Z(n37206) );
  NANDN U37678 ( .A(n37426), .B(n37427), .Z(n37425) );
  OR U37679 ( .A(n37428), .B(n37429), .Z(n37427) );
  NAND U37680 ( .A(n37429), .B(n37428), .Z(n37424) );
  ANDN U37681 ( .B(B[147]), .A(n67), .Z(n37208) );
  XNOR U37682 ( .A(n37216), .B(n37430), .Z(n37209) );
  XNOR U37683 ( .A(n37215), .B(n37213), .Z(n37430) );
  AND U37684 ( .A(n37431), .B(n37432), .Z(n37213) );
  NANDN U37685 ( .A(n37433), .B(n37434), .Z(n37432) );
  NANDN U37686 ( .A(n37435), .B(n37436), .Z(n37434) );
  NANDN U37687 ( .A(n37436), .B(n37435), .Z(n37431) );
  ANDN U37688 ( .B(B[148]), .A(n68), .Z(n37215) );
  XNOR U37689 ( .A(n37223), .B(n37437), .Z(n37216) );
  XNOR U37690 ( .A(n37222), .B(n37220), .Z(n37437) );
  AND U37691 ( .A(n37438), .B(n37439), .Z(n37220) );
  NANDN U37692 ( .A(n37440), .B(n37441), .Z(n37439) );
  OR U37693 ( .A(n37442), .B(n37443), .Z(n37441) );
  NAND U37694 ( .A(n37443), .B(n37442), .Z(n37438) );
  ANDN U37695 ( .B(B[149]), .A(n69), .Z(n37222) );
  XNOR U37696 ( .A(n37230), .B(n37444), .Z(n37223) );
  XNOR U37697 ( .A(n37229), .B(n37227), .Z(n37444) );
  AND U37698 ( .A(n37445), .B(n37446), .Z(n37227) );
  NANDN U37699 ( .A(n37447), .B(n37448), .Z(n37446) );
  NANDN U37700 ( .A(n37449), .B(n37450), .Z(n37448) );
  NANDN U37701 ( .A(n37450), .B(n37449), .Z(n37445) );
  ANDN U37702 ( .B(B[150]), .A(n70), .Z(n37229) );
  XNOR U37703 ( .A(n37237), .B(n37451), .Z(n37230) );
  XNOR U37704 ( .A(n37236), .B(n37234), .Z(n37451) );
  AND U37705 ( .A(n37452), .B(n37453), .Z(n37234) );
  NANDN U37706 ( .A(n37454), .B(n37455), .Z(n37453) );
  OR U37707 ( .A(n37456), .B(n37457), .Z(n37455) );
  NAND U37708 ( .A(n37457), .B(n37456), .Z(n37452) );
  ANDN U37709 ( .B(B[151]), .A(n71), .Z(n37236) );
  XNOR U37710 ( .A(n37244), .B(n37458), .Z(n37237) );
  XNOR U37711 ( .A(n37243), .B(n37241), .Z(n37458) );
  AND U37712 ( .A(n37459), .B(n37460), .Z(n37241) );
  NANDN U37713 ( .A(n37461), .B(n37462), .Z(n37460) );
  NANDN U37714 ( .A(n37463), .B(n37464), .Z(n37462) );
  NANDN U37715 ( .A(n37464), .B(n37463), .Z(n37459) );
  ANDN U37716 ( .B(B[152]), .A(n72), .Z(n37243) );
  XNOR U37717 ( .A(n37251), .B(n37465), .Z(n37244) );
  XNOR U37718 ( .A(n37250), .B(n37248), .Z(n37465) );
  AND U37719 ( .A(n37466), .B(n37467), .Z(n37248) );
  NANDN U37720 ( .A(n37468), .B(n37469), .Z(n37467) );
  OR U37721 ( .A(n37470), .B(n37471), .Z(n37469) );
  NAND U37722 ( .A(n37471), .B(n37470), .Z(n37466) );
  ANDN U37723 ( .B(B[153]), .A(n73), .Z(n37250) );
  XNOR U37724 ( .A(n37258), .B(n37472), .Z(n37251) );
  XNOR U37725 ( .A(n37257), .B(n37255), .Z(n37472) );
  AND U37726 ( .A(n37473), .B(n37474), .Z(n37255) );
  NANDN U37727 ( .A(n37475), .B(n37476), .Z(n37474) );
  NANDN U37728 ( .A(n37477), .B(n37478), .Z(n37476) );
  NANDN U37729 ( .A(n37478), .B(n37477), .Z(n37473) );
  ANDN U37730 ( .B(B[154]), .A(n74), .Z(n37257) );
  XNOR U37731 ( .A(n37265), .B(n37479), .Z(n37258) );
  XNOR U37732 ( .A(n37264), .B(n37262), .Z(n37479) );
  AND U37733 ( .A(n37480), .B(n37481), .Z(n37262) );
  NANDN U37734 ( .A(n37482), .B(n37483), .Z(n37481) );
  OR U37735 ( .A(n37484), .B(n37485), .Z(n37483) );
  NAND U37736 ( .A(n37485), .B(n37484), .Z(n37480) );
  ANDN U37737 ( .B(B[155]), .A(n75), .Z(n37264) );
  XNOR U37738 ( .A(n37272), .B(n37486), .Z(n37265) );
  XNOR U37739 ( .A(n37271), .B(n37269), .Z(n37486) );
  AND U37740 ( .A(n37487), .B(n37488), .Z(n37269) );
  NANDN U37741 ( .A(n37489), .B(n37490), .Z(n37488) );
  NANDN U37742 ( .A(n37491), .B(n37492), .Z(n37490) );
  NANDN U37743 ( .A(n37492), .B(n37491), .Z(n37487) );
  ANDN U37744 ( .B(B[156]), .A(n76), .Z(n37271) );
  XNOR U37745 ( .A(n37279), .B(n37493), .Z(n37272) );
  XNOR U37746 ( .A(n37278), .B(n37276), .Z(n37493) );
  AND U37747 ( .A(n37494), .B(n37495), .Z(n37276) );
  NANDN U37748 ( .A(n37496), .B(n37497), .Z(n37495) );
  OR U37749 ( .A(n37498), .B(n37499), .Z(n37497) );
  NAND U37750 ( .A(n37499), .B(n37498), .Z(n37494) );
  ANDN U37751 ( .B(B[157]), .A(n77), .Z(n37278) );
  XNOR U37752 ( .A(n37286), .B(n37500), .Z(n37279) );
  XNOR U37753 ( .A(n37285), .B(n37283), .Z(n37500) );
  AND U37754 ( .A(n37501), .B(n37502), .Z(n37283) );
  NANDN U37755 ( .A(n37503), .B(n37504), .Z(n37502) );
  NANDN U37756 ( .A(n37505), .B(n37506), .Z(n37504) );
  NANDN U37757 ( .A(n37506), .B(n37505), .Z(n37501) );
  ANDN U37758 ( .B(B[158]), .A(n78), .Z(n37285) );
  XNOR U37759 ( .A(n37293), .B(n37507), .Z(n37286) );
  XNOR U37760 ( .A(n37292), .B(n37290), .Z(n37507) );
  AND U37761 ( .A(n37508), .B(n37509), .Z(n37290) );
  NANDN U37762 ( .A(n37510), .B(n37511), .Z(n37509) );
  OR U37763 ( .A(n37512), .B(n37513), .Z(n37511) );
  NAND U37764 ( .A(n37513), .B(n37512), .Z(n37508) );
  ANDN U37765 ( .B(B[159]), .A(n79), .Z(n37292) );
  XNOR U37766 ( .A(n37300), .B(n37514), .Z(n37293) );
  XNOR U37767 ( .A(n37299), .B(n37297), .Z(n37514) );
  AND U37768 ( .A(n37515), .B(n37516), .Z(n37297) );
  NANDN U37769 ( .A(n37517), .B(n37518), .Z(n37516) );
  NANDN U37770 ( .A(n37519), .B(n37520), .Z(n37518) );
  NANDN U37771 ( .A(n37520), .B(n37519), .Z(n37515) );
  ANDN U37772 ( .B(B[160]), .A(n80), .Z(n37299) );
  XNOR U37773 ( .A(n37307), .B(n37521), .Z(n37300) );
  XNOR U37774 ( .A(n37306), .B(n37304), .Z(n37521) );
  AND U37775 ( .A(n37522), .B(n37523), .Z(n37304) );
  NANDN U37776 ( .A(n37524), .B(n37525), .Z(n37523) );
  OR U37777 ( .A(n37526), .B(n37527), .Z(n37525) );
  NAND U37778 ( .A(n37527), .B(n37526), .Z(n37522) );
  ANDN U37779 ( .B(B[161]), .A(n81), .Z(n37306) );
  XNOR U37780 ( .A(n37314), .B(n37528), .Z(n37307) );
  XNOR U37781 ( .A(n37313), .B(n37311), .Z(n37528) );
  AND U37782 ( .A(n37529), .B(n37530), .Z(n37311) );
  NANDN U37783 ( .A(n37531), .B(n37532), .Z(n37530) );
  NAND U37784 ( .A(n37533), .B(n37534), .Z(n37532) );
  ANDN U37785 ( .B(B[162]), .A(n82), .Z(n37313) );
  XOR U37786 ( .A(n37320), .B(n37535), .Z(n37314) );
  XNOR U37787 ( .A(n37318), .B(n37321), .Z(n37535) );
  NAND U37788 ( .A(A[2]), .B(B[163]), .Z(n37321) );
  NANDN U37789 ( .A(n37536), .B(n37537), .Z(n37318) );
  AND U37790 ( .A(A[0]), .B(B[164]), .Z(n37537) );
  XNOR U37791 ( .A(n37323), .B(n37538), .Z(n37320) );
  NAND U37792 ( .A(A[0]), .B(B[165]), .Z(n37538) );
  NAND U37793 ( .A(B[164]), .B(A[1]), .Z(n37323) );
  NAND U37794 ( .A(n37539), .B(n37540), .Z(n466) );
  NANDN U37795 ( .A(n37541), .B(n37542), .Z(n37540) );
  OR U37796 ( .A(n37543), .B(n37544), .Z(n37542) );
  NAND U37797 ( .A(n37544), .B(n37543), .Z(n37539) );
  XOR U37798 ( .A(n468), .B(n467), .Z(\A1[162] ) );
  XOR U37799 ( .A(n37544), .B(n37545), .Z(n467) );
  XNOR U37800 ( .A(n37543), .B(n37541), .Z(n37545) );
  AND U37801 ( .A(n37546), .B(n37547), .Z(n37541) );
  NANDN U37802 ( .A(n37548), .B(n37549), .Z(n37547) );
  NANDN U37803 ( .A(n37550), .B(n37551), .Z(n37549) );
  NANDN U37804 ( .A(n37551), .B(n37550), .Z(n37546) );
  ANDN U37805 ( .B(B[133]), .A(n54), .Z(n37543) );
  XNOR U37806 ( .A(n37338), .B(n37552), .Z(n37544) );
  XNOR U37807 ( .A(n37337), .B(n37335), .Z(n37552) );
  AND U37808 ( .A(n37553), .B(n37554), .Z(n37335) );
  NANDN U37809 ( .A(n37555), .B(n37556), .Z(n37554) );
  OR U37810 ( .A(n37557), .B(n37558), .Z(n37556) );
  NAND U37811 ( .A(n37558), .B(n37557), .Z(n37553) );
  ANDN U37812 ( .B(B[134]), .A(n55), .Z(n37337) );
  XNOR U37813 ( .A(n37345), .B(n37559), .Z(n37338) );
  XNOR U37814 ( .A(n37344), .B(n37342), .Z(n37559) );
  AND U37815 ( .A(n37560), .B(n37561), .Z(n37342) );
  NANDN U37816 ( .A(n37562), .B(n37563), .Z(n37561) );
  NANDN U37817 ( .A(n37564), .B(n37565), .Z(n37563) );
  NANDN U37818 ( .A(n37565), .B(n37564), .Z(n37560) );
  ANDN U37819 ( .B(B[135]), .A(n56), .Z(n37344) );
  XNOR U37820 ( .A(n37352), .B(n37566), .Z(n37345) );
  XNOR U37821 ( .A(n37351), .B(n37349), .Z(n37566) );
  AND U37822 ( .A(n37567), .B(n37568), .Z(n37349) );
  NANDN U37823 ( .A(n37569), .B(n37570), .Z(n37568) );
  OR U37824 ( .A(n37571), .B(n37572), .Z(n37570) );
  NAND U37825 ( .A(n37572), .B(n37571), .Z(n37567) );
  ANDN U37826 ( .B(B[136]), .A(n57), .Z(n37351) );
  XNOR U37827 ( .A(n37359), .B(n37573), .Z(n37352) );
  XNOR U37828 ( .A(n37358), .B(n37356), .Z(n37573) );
  AND U37829 ( .A(n37574), .B(n37575), .Z(n37356) );
  NANDN U37830 ( .A(n37576), .B(n37577), .Z(n37575) );
  NANDN U37831 ( .A(n37578), .B(n37579), .Z(n37577) );
  NANDN U37832 ( .A(n37579), .B(n37578), .Z(n37574) );
  ANDN U37833 ( .B(B[137]), .A(n58), .Z(n37358) );
  XNOR U37834 ( .A(n37366), .B(n37580), .Z(n37359) );
  XNOR U37835 ( .A(n37365), .B(n37363), .Z(n37580) );
  AND U37836 ( .A(n37581), .B(n37582), .Z(n37363) );
  NANDN U37837 ( .A(n37583), .B(n37584), .Z(n37582) );
  OR U37838 ( .A(n37585), .B(n37586), .Z(n37584) );
  NAND U37839 ( .A(n37586), .B(n37585), .Z(n37581) );
  ANDN U37840 ( .B(B[138]), .A(n59), .Z(n37365) );
  XNOR U37841 ( .A(n37373), .B(n37587), .Z(n37366) );
  XNOR U37842 ( .A(n37372), .B(n37370), .Z(n37587) );
  AND U37843 ( .A(n37588), .B(n37589), .Z(n37370) );
  NANDN U37844 ( .A(n37590), .B(n37591), .Z(n37589) );
  NANDN U37845 ( .A(n37592), .B(n37593), .Z(n37591) );
  NANDN U37846 ( .A(n37593), .B(n37592), .Z(n37588) );
  ANDN U37847 ( .B(B[139]), .A(n60), .Z(n37372) );
  XNOR U37848 ( .A(n37380), .B(n37594), .Z(n37373) );
  XNOR U37849 ( .A(n37379), .B(n37377), .Z(n37594) );
  AND U37850 ( .A(n37595), .B(n37596), .Z(n37377) );
  NANDN U37851 ( .A(n37597), .B(n37598), .Z(n37596) );
  OR U37852 ( .A(n37599), .B(n37600), .Z(n37598) );
  NAND U37853 ( .A(n37600), .B(n37599), .Z(n37595) );
  ANDN U37854 ( .B(B[140]), .A(n61), .Z(n37379) );
  XNOR U37855 ( .A(n37387), .B(n37601), .Z(n37380) );
  XNOR U37856 ( .A(n37386), .B(n37384), .Z(n37601) );
  AND U37857 ( .A(n37602), .B(n37603), .Z(n37384) );
  NANDN U37858 ( .A(n37604), .B(n37605), .Z(n37603) );
  NANDN U37859 ( .A(n37606), .B(n37607), .Z(n37605) );
  NANDN U37860 ( .A(n37607), .B(n37606), .Z(n37602) );
  ANDN U37861 ( .B(B[141]), .A(n62), .Z(n37386) );
  XNOR U37862 ( .A(n37394), .B(n37608), .Z(n37387) );
  XNOR U37863 ( .A(n37393), .B(n37391), .Z(n37608) );
  AND U37864 ( .A(n37609), .B(n37610), .Z(n37391) );
  NANDN U37865 ( .A(n37611), .B(n37612), .Z(n37610) );
  OR U37866 ( .A(n37613), .B(n37614), .Z(n37612) );
  NAND U37867 ( .A(n37614), .B(n37613), .Z(n37609) );
  ANDN U37868 ( .B(B[142]), .A(n63), .Z(n37393) );
  XNOR U37869 ( .A(n37401), .B(n37615), .Z(n37394) );
  XNOR U37870 ( .A(n37400), .B(n37398), .Z(n37615) );
  AND U37871 ( .A(n37616), .B(n37617), .Z(n37398) );
  NANDN U37872 ( .A(n37618), .B(n37619), .Z(n37617) );
  NANDN U37873 ( .A(n37620), .B(n37621), .Z(n37619) );
  NANDN U37874 ( .A(n37621), .B(n37620), .Z(n37616) );
  ANDN U37875 ( .B(B[143]), .A(n64), .Z(n37400) );
  XNOR U37876 ( .A(n37408), .B(n37622), .Z(n37401) );
  XNOR U37877 ( .A(n37407), .B(n37405), .Z(n37622) );
  AND U37878 ( .A(n37623), .B(n37624), .Z(n37405) );
  NANDN U37879 ( .A(n37625), .B(n37626), .Z(n37624) );
  OR U37880 ( .A(n37627), .B(n37628), .Z(n37626) );
  NAND U37881 ( .A(n37628), .B(n37627), .Z(n37623) );
  ANDN U37882 ( .B(B[144]), .A(n65), .Z(n37407) );
  XNOR U37883 ( .A(n37415), .B(n37629), .Z(n37408) );
  XNOR U37884 ( .A(n37414), .B(n37412), .Z(n37629) );
  AND U37885 ( .A(n37630), .B(n37631), .Z(n37412) );
  NANDN U37886 ( .A(n37632), .B(n37633), .Z(n37631) );
  NANDN U37887 ( .A(n37634), .B(n37635), .Z(n37633) );
  NANDN U37888 ( .A(n37635), .B(n37634), .Z(n37630) );
  ANDN U37889 ( .B(B[145]), .A(n66), .Z(n37414) );
  XNOR U37890 ( .A(n37422), .B(n37636), .Z(n37415) );
  XNOR U37891 ( .A(n37421), .B(n37419), .Z(n37636) );
  AND U37892 ( .A(n37637), .B(n37638), .Z(n37419) );
  NANDN U37893 ( .A(n37639), .B(n37640), .Z(n37638) );
  OR U37894 ( .A(n37641), .B(n37642), .Z(n37640) );
  NAND U37895 ( .A(n37642), .B(n37641), .Z(n37637) );
  ANDN U37896 ( .B(B[146]), .A(n67), .Z(n37421) );
  XNOR U37897 ( .A(n37429), .B(n37643), .Z(n37422) );
  XNOR U37898 ( .A(n37428), .B(n37426), .Z(n37643) );
  AND U37899 ( .A(n37644), .B(n37645), .Z(n37426) );
  NANDN U37900 ( .A(n37646), .B(n37647), .Z(n37645) );
  NANDN U37901 ( .A(n37648), .B(n37649), .Z(n37647) );
  NANDN U37902 ( .A(n37649), .B(n37648), .Z(n37644) );
  ANDN U37903 ( .B(B[147]), .A(n68), .Z(n37428) );
  XNOR U37904 ( .A(n37436), .B(n37650), .Z(n37429) );
  XNOR U37905 ( .A(n37435), .B(n37433), .Z(n37650) );
  AND U37906 ( .A(n37651), .B(n37652), .Z(n37433) );
  NANDN U37907 ( .A(n37653), .B(n37654), .Z(n37652) );
  OR U37908 ( .A(n37655), .B(n37656), .Z(n37654) );
  NAND U37909 ( .A(n37656), .B(n37655), .Z(n37651) );
  ANDN U37910 ( .B(B[148]), .A(n69), .Z(n37435) );
  XNOR U37911 ( .A(n37443), .B(n37657), .Z(n37436) );
  XNOR U37912 ( .A(n37442), .B(n37440), .Z(n37657) );
  AND U37913 ( .A(n37658), .B(n37659), .Z(n37440) );
  NANDN U37914 ( .A(n37660), .B(n37661), .Z(n37659) );
  NANDN U37915 ( .A(n37662), .B(n37663), .Z(n37661) );
  NANDN U37916 ( .A(n37663), .B(n37662), .Z(n37658) );
  ANDN U37917 ( .B(B[149]), .A(n70), .Z(n37442) );
  XNOR U37918 ( .A(n37450), .B(n37664), .Z(n37443) );
  XNOR U37919 ( .A(n37449), .B(n37447), .Z(n37664) );
  AND U37920 ( .A(n37665), .B(n37666), .Z(n37447) );
  NANDN U37921 ( .A(n37667), .B(n37668), .Z(n37666) );
  OR U37922 ( .A(n37669), .B(n37670), .Z(n37668) );
  NAND U37923 ( .A(n37670), .B(n37669), .Z(n37665) );
  ANDN U37924 ( .B(B[150]), .A(n71), .Z(n37449) );
  XNOR U37925 ( .A(n37457), .B(n37671), .Z(n37450) );
  XNOR U37926 ( .A(n37456), .B(n37454), .Z(n37671) );
  AND U37927 ( .A(n37672), .B(n37673), .Z(n37454) );
  NANDN U37928 ( .A(n37674), .B(n37675), .Z(n37673) );
  NANDN U37929 ( .A(n37676), .B(n37677), .Z(n37675) );
  NANDN U37930 ( .A(n37677), .B(n37676), .Z(n37672) );
  ANDN U37931 ( .B(B[151]), .A(n72), .Z(n37456) );
  XNOR U37932 ( .A(n37464), .B(n37678), .Z(n37457) );
  XNOR U37933 ( .A(n37463), .B(n37461), .Z(n37678) );
  AND U37934 ( .A(n37679), .B(n37680), .Z(n37461) );
  NANDN U37935 ( .A(n37681), .B(n37682), .Z(n37680) );
  OR U37936 ( .A(n37683), .B(n37684), .Z(n37682) );
  NAND U37937 ( .A(n37684), .B(n37683), .Z(n37679) );
  ANDN U37938 ( .B(B[152]), .A(n73), .Z(n37463) );
  XNOR U37939 ( .A(n37471), .B(n37685), .Z(n37464) );
  XNOR U37940 ( .A(n37470), .B(n37468), .Z(n37685) );
  AND U37941 ( .A(n37686), .B(n37687), .Z(n37468) );
  NANDN U37942 ( .A(n37688), .B(n37689), .Z(n37687) );
  NANDN U37943 ( .A(n37690), .B(n37691), .Z(n37689) );
  NANDN U37944 ( .A(n37691), .B(n37690), .Z(n37686) );
  ANDN U37945 ( .B(B[153]), .A(n74), .Z(n37470) );
  XNOR U37946 ( .A(n37478), .B(n37692), .Z(n37471) );
  XNOR U37947 ( .A(n37477), .B(n37475), .Z(n37692) );
  AND U37948 ( .A(n37693), .B(n37694), .Z(n37475) );
  NANDN U37949 ( .A(n37695), .B(n37696), .Z(n37694) );
  OR U37950 ( .A(n37697), .B(n37698), .Z(n37696) );
  NAND U37951 ( .A(n37698), .B(n37697), .Z(n37693) );
  ANDN U37952 ( .B(B[154]), .A(n75), .Z(n37477) );
  XNOR U37953 ( .A(n37485), .B(n37699), .Z(n37478) );
  XNOR U37954 ( .A(n37484), .B(n37482), .Z(n37699) );
  AND U37955 ( .A(n37700), .B(n37701), .Z(n37482) );
  NANDN U37956 ( .A(n37702), .B(n37703), .Z(n37701) );
  NANDN U37957 ( .A(n37704), .B(n37705), .Z(n37703) );
  NANDN U37958 ( .A(n37705), .B(n37704), .Z(n37700) );
  ANDN U37959 ( .B(B[155]), .A(n76), .Z(n37484) );
  XNOR U37960 ( .A(n37492), .B(n37706), .Z(n37485) );
  XNOR U37961 ( .A(n37491), .B(n37489), .Z(n37706) );
  AND U37962 ( .A(n37707), .B(n37708), .Z(n37489) );
  NANDN U37963 ( .A(n37709), .B(n37710), .Z(n37708) );
  OR U37964 ( .A(n37711), .B(n37712), .Z(n37710) );
  NAND U37965 ( .A(n37712), .B(n37711), .Z(n37707) );
  ANDN U37966 ( .B(B[156]), .A(n77), .Z(n37491) );
  XNOR U37967 ( .A(n37499), .B(n37713), .Z(n37492) );
  XNOR U37968 ( .A(n37498), .B(n37496), .Z(n37713) );
  AND U37969 ( .A(n37714), .B(n37715), .Z(n37496) );
  NANDN U37970 ( .A(n37716), .B(n37717), .Z(n37715) );
  NANDN U37971 ( .A(n37718), .B(n37719), .Z(n37717) );
  NANDN U37972 ( .A(n37719), .B(n37718), .Z(n37714) );
  ANDN U37973 ( .B(B[157]), .A(n78), .Z(n37498) );
  XNOR U37974 ( .A(n37506), .B(n37720), .Z(n37499) );
  XNOR U37975 ( .A(n37505), .B(n37503), .Z(n37720) );
  AND U37976 ( .A(n37721), .B(n37722), .Z(n37503) );
  NANDN U37977 ( .A(n37723), .B(n37724), .Z(n37722) );
  OR U37978 ( .A(n37725), .B(n37726), .Z(n37724) );
  NAND U37979 ( .A(n37726), .B(n37725), .Z(n37721) );
  ANDN U37980 ( .B(B[158]), .A(n79), .Z(n37505) );
  XNOR U37981 ( .A(n37513), .B(n37727), .Z(n37506) );
  XNOR U37982 ( .A(n37512), .B(n37510), .Z(n37727) );
  AND U37983 ( .A(n37728), .B(n37729), .Z(n37510) );
  NANDN U37984 ( .A(n37730), .B(n37731), .Z(n37729) );
  NANDN U37985 ( .A(n37732), .B(n37733), .Z(n37731) );
  NANDN U37986 ( .A(n37733), .B(n37732), .Z(n37728) );
  ANDN U37987 ( .B(B[159]), .A(n80), .Z(n37512) );
  XNOR U37988 ( .A(n37520), .B(n37734), .Z(n37513) );
  XNOR U37989 ( .A(n37519), .B(n37517), .Z(n37734) );
  AND U37990 ( .A(n37735), .B(n37736), .Z(n37517) );
  NANDN U37991 ( .A(n37737), .B(n37738), .Z(n37736) );
  OR U37992 ( .A(n37739), .B(n37740), .Z(n37738) );
  NAND U37993 ( .A(n37740), .B(n37739), .Z(n37735) );
  ANDN U37994 ( .B(B[160]), .A(n81), .Z(n37519) );
  XNOR U37995 ( .A(n37527), .B(n37741), .Z(n37520) );
  XNOR U37996 ( .A(n37526), .B(n37524), .Z(n37741) );
  AND U37997 ( .A(n37742), .B(n37743), .Z(n37524) );
  NANDN U37998 ( .A(n37744), .B(n37745), .Z(n37743) );
  NAND U37999 ( .A(n37746), .B(n37747), .Z(n37745) );
  ANDN U38000 ( .B(B[161]), .A(n82), .Z(n37526) );
  XOR U38001 ( .A(n37533), .B(n37748), .Z(n37527) );
  XNOR U38002 ( .A(n37531), .B(n37534), .Z(n37748) );
  NAND U38003 ( .A(A[2]), .B(B[162]), .Z(n37534) );
  NANDN U38004 ( .A(n37749), .B(n37750), .Z(n37531) );
  AND U38005 ( .A(A[0]), .B(B[163]), .Z(n37750) );
  XNOR U38006 ( .A(n37536), .B(n37751), .Z(n37533) );
  NAND U38007 ( .A(A[0]), .B(B[164]), .Z(n37751) );
  NAND U38008 ( .A(B[163]), .B(A[1]), .Z(n37536) );
  NAND U38009 ( .A(n37752), .B(n37753), .Z(n468) );
  NANDN U38010 ( .A(n37754), .B(n37755), .Z(n37753) );
  OR U38011 ( .A(n37756), .B(n37757), .Z(n37755) );
  NAND U38012 ( .A(n37757), .B(n37756), .Z(n37752) );
  XOR U38013 ( .A(n470), .B(n469), .Z(\A1[161] ) );
  XOR U38014 ( .A(n37757), .B(n37758), .Z(n469) );
  XNOR U38015 ( .A(n37756), .B(n37754), .Z(n37758) );
  AND U38016 ( .A(n37759), .B(n37760), .Z(n37754) );
  NANDN U38017 ( .A(n37761), .B(n37762), .Z(n37760) );
  NANDN U38018 ( .A(n37763), .B(n37764), .Z(n37762) );
  NANDN U38019 ( .A(n37764), .B(n37763), .Z(n37759) );
  ANDN U38020 ( .B(B[132]), .A(n54), .Z(n37756) );
  XNOR U38021 ( .A(n37551), .B(n37765), .Z(n37757) );
  XNOR U38022 ( .A(n37550), .B(n37548), .Z(n37765) );
  AND U38023 ( .A(n37766), .B(n37767), .Z(n37548) );
  NANDN U38024 ( .A(n37768), .B(n37769), .Z(n37767) );
  OR U38025 ( .A(n37770), .B(n37771), .Z(n37769) );
  NAND U38026 ( .A(n37771), .B(n37770), .Z(n37766) );
  ANDN U38027 ( .B(B[133]), .A(n55), .Z(n37550) );
  XNOR U38028 ( .A(n37558), .B(n37772), .Z(n37551) );
  XNOR U38029 ( .A(n37557), .B(n37555), .Z(n37772) );
  AND U38030 ( .A(n37773), .B(n37774), .Z(n37555) );
  NANDN U38031 ( .A(n37775), .B(n37776), .Z(n37774) );
  NANDN U38032 ( .A(n37777), .B(n37778), .Z(n37776) );
  NANDN U38033 ( .A(n37778), .B(n37777), .Z(n37773) );
  ANDN U38034 ( .B(B[134]), .A(n56), .Z(n37557) );
  XNOR U38035 ( .A(n37565), .B(n37779), .Z(n37558) );
  XNOR U38036 ( .A(n37564), .B(n37562), .Z(n37779) );
  AND U38037 ( .A(n37780), .B(n37781), .Z(n37562) );
  NANDN U38038 ( .A(n37782), .B(n37783), .Z(n37781) );
  OR U38039 ( .A(n37784), .B(n37785), .Z(n37783) );
  NAND U38040 ( .A(n37785), .B(n37784), .Z(n37780) );
  ANDN U38041 ( .B(B[135]), .A(n57), .Z(n37564) );
  XNOR U38042 ( .A(n37572), .B(n37786), .Z(n37565) );
  XNOR U38043 ( .A(n37571), .B(n37569), .Z(n37786) );
  AND U38044 ( .A(n37787), .B(n37788), .Z(n37569) );
  NANDN U38045 ( .A(n37789), .B(n37790), .Z(n37788) );
  NANDN U38046 ( .A(n37791), .B(n37792), .Z(n37790) );
  NANDN U38047 ( .A(n37792), .B(n37791), .Z(n37787) );
  ANDN U38048 ( .B(B[136]), .A(n58), .Z(n37571) );
  XNOR U38049 ( .A(n37579), .B(n37793), .Z(n37572) );
  XNOR U38050 ( .A(n37578), .B(n37576), .Z(n37793) );
  AND U38051 ( .A(n37794), .B(n37795), .Z(n37576) );
  NANDN U38052 ( .A(n37796), .B(n37797), .Z(n37795) );
  OR U38053 ( .A(n37798), .B(n37799), .Z(n37797) );
  NAND U38054 ( .A(n37799), .B(n37798), .Z(n37794) );
  ANDN U38055 ( .B(B[137]), .A(n59), .Z(n37578) );
  XNOR U38056 ( .A(n37586), .B(n37800), .Z(n37579) );
  XNOR U38057 ( .A(n37585), .B(n37583), .Z(n37800) );
  AND U38058 ( .A(n37801), .B(n37802), .Z(n37583) );
  NANDN U38059 ( .A(n37803), .B(n37804), .Z(n37802) );
  NANDN U38060 ( .A(n37805), .B(n37806), .Z(n37804) );
  NANDN U38061 ( .A(n37806), .B(n37805), .Z(n37801) );
  ANDN U38062 ( .B(B[138]), .A(n60), .Z(n37585) );
  XNOR U38063 ( .A(n37593), .B(n37807), .Z(n37586) );
  XNOR U38064 ( .A(n37592), .B(n37590), .Z(n37807) );
  AND U38065 ( .A(n37808), .B(n37809), .Z(n37590) );
  NANDN U38066 ( .A(n37810), .B(n37811), .Z(n37809) );
  OR U38067 ( .A(n37812), .B(n37813), .Z(n37811) );
  NAND U38068 ( .A(n37813), .B(n37812), .Z(n37808) );
  ANDN U38069 ( .B(B[139]), .A(n61), .Z(n37592) );
  XNOR U38070 ( .A(n37600), .B(n37814), .Z(n37593) );
  XNOR U38071 ( .A(n37599), .B(n37597), .Z(n37814) );
  AND U38072 ( .A(n37815), .B(n37816), .Z(n37597) );
  NANDN U38073 ( .A(n37817), .B(n37818), .Z(n37816) );
  NANDN U38074 ( .A(n37819), .B(n37820), .Z(n37818) );
  NANDN U38075 ( .A(n37820), .B(n37819), .Z(n37815) );
  ANDN U38076 ( .B(B[140]), .A(n62), .Z(n37599) );
  XNOR U38077 ( .A(n37607), .B(n37821), .Z(n37600) );
  XNOR U38078 ( .A(n37606), .B(n37604), .Z(n37821) );
  AND U38079 ( .A(n37822), .B(n37823), .Z(n37604) );
  NANDN U38080 ( .A(n37824), .B(n37825), .Z(n37823) );
  OR U38081 ( .A(n37826), .B(n37827), .Z(n37825) );
  NAND U38082 ( .A(n37827), .B(n37826), .Z(n37822) );
  ANDN U38083 ( .B(B[141]), .A(n63), .Z(n37606) );
  XNOR U38084 ( .A(n37614), .B(n37828), .Z(n37607) );
  XNOR U38085 ( .A(n37613), .B(n37611), .Z(n37828) );
  AND U38086 ( .A(n37829), .B(n37830), .Z(n37611) );
  NANDN U38087 ( .A(n37831), .B(n37832), .Z(n37830) );
  NANDN U38088 ( .A(n37833), .B(n37834), .Z(n37832) );
  NANDN U38089 ( .A(n37834), .B(n37833), .Z(n37829) );
  ANDN U38090 ( .B(B[142]), .A(n64), .Z(n37613) );
  XNOR U38091 ( .A(n37621), .B(n37835), .Z(n37614) );
  XNOR U38092 ( .A(n37620), .B(n37618), .Z(n37835) );
  AND U38093 ( .A(n37836), .B(n37837), .Z(n37618) );
  NANDN U38094 ( .A(n37838), .B(n37839), .Z(n37837) );
  OR U38095 ( .A(n37840), .B(n37841), .Z(n37839) );
  NAND U38096 ( .A(n37841), .B(n37840), .Z(n37836) );
  ANDN U38097 ( .B(B[143]), .A(n65), .Z(n37620) );
  XNOR U38098 ( .A(n37628), .B(n37842), .Z(n37621) );
  XNOR U38099 ( .A(n37627), .B(n37625), .Z(n37842) );
  AND U38100 ( .A(n37843), .B(n37844), .Z(n37625) );
  NANDN U38101 ( .A(n37845), .B(n37846), .Z(n37844) );
  NANDN U38102 ( .A(n37847), .B(n37848), .Z(n37846) );
  NANDN U38103 ( .A(n37848), .B(n37847), .Z(n37843) );
  ANDN U38104 ( .B(B[144]), .A(n66), .Z(n37627) );
  XNOR U38105 ( .A(n37635), .B(n37849), .Z(n37628) );
  XNOR U38106 ( .A(n37634), .B(n37632), .Z(n37849) );
  AND U38107 ( .A(n37850), .B(n37851), .Z(n37632) );
  NANDN U38108 ( .A(n37852), .B(n37853), .Z(n37851) );
  OR U38109 ( .A(n37854), .B(n37855), .Z(n37853) );
  NAND U38110 ( .A(n37855), .B(n37854), .Z(n37850) );
  ANDN U38111 ( .B(B[145]), .A(n67), .Z(n37634) );
  XNOR U38112 ( .A(n37642), .B(n37856), .Z(n37635) );
  XNOR U38113 ( .A(n37641), .B(n37639), .Z(n37856) );
  AND U38114 ( .A(n37857), .B(n37858), .Z(n37639) );
  NANDN U38115 ( .A(n37859), .B(n37860), .Z(n37858) );
  NANDN U38116 ( .A(n37861), .B(n37862), .Z(n37860) );
  NANDN U38117 ( .A(n37862), .B(n37861), .Z(n37857) );
  ANDN U38118 ( .B(B[146]), .A(n68), .Z(n37641) );
  XNOR U38119 ( .A(n37649), .B(n37863), .Z(n37642) );
  XNOR U38120 ( .A(n37648), .B(n37646), .Z(n37863) );
  AND U38121 ( .A(n37864), .B(n37865), .Z(n37646) );
  NANDN U38122 ( .A(n37866), .B(n37867), .Z(n37865) );
  OR U38123 ( .A(n37868), .B(n37869), .Z(n37867) );
  NAND U38124 ( .A(n37869), .B(n37868), .Z(n37864) );
  ANDN U38125 ( .B(B[147]), .A(n69), .Z(n37648) );
  XNOR U38126 ( .A(n37656), .B(n37870), .Z(n37649) );
  XNOR U38127 ( .A(n37655), .B(n37653), .Z(n37870) );
  AND U38128 ( .A(n37871), .B(n37872), .Z(n37653) );
  NANDN U38129 ( .A(n37873), .B(n37874), .Z(n37872) );
  NANDN U38130 ( .A(n37875), .B(n37876), .Z(n37874) );
  NANDN U38131 ( .A(n37876), .B(n37875), .Z(n37871) );
  ANDN U38132 ( .B(B[148]), .A(n70), .Z(n37655) );
  XNOR U38133 ( .A(n37663), .B(n37877), .Z(n37656) );
  XNOR U38134 ( .A(n37662), .B(n37660), .Z(n37877) );
  AND U38135 ( .A(n37878), .B(n37879), .Z(n37660) );
  NANDN U38136 ( .A(n37880), .B(n37881), .Z(n37879) );
  OR U38137 ( .A(n37882), .B(n37883), .Z(n37881) );
  NAND U38138 ( .A(n37883), .B(n37882), .Z(n37878) );
  ANDN U38139 ( .B(B[149]), .A(n71), .Z(n37662) );
  XNOR U38140 ( .A(n37670), .B(n37884), .Z(n37663) );
  XNOR U38141 ( .A(n37669), .B(n37667), .Z(n37884) );
  AND U38142 ( .A(n37885), .B(n37886), .Z(n37667) );
  NANDN U38143 ( .A(n37887), .B(n37888), .Z(n37886) );
  NANDN U38144 ( .A(n37889), .B(n37890), .Z(n37888) );
  NANDN U38145 ( .A(n37890), .B(n37889), .Z(n37885) );
  ANDN U38146 ( .B(B[150]), .A(n72), .Z(n37669) );
  XNOR U38147 ( .A(n37677), .B(n37891), .Z(n37670) );
  XNOR U38148 ( .A(n37676), .B(n37674), .Z(n37891) );
  AND U38149 ( .A(n37892), .B(n37893), .Z(n37674) );
  NANDN U38150 ( .A(n37894), .B(n37895), .Z(n37893) );
  OR U38151 ( .A(n37896), .B(n37897), .Z(n37895) );
  NAND U38152 ( .A(n37897), .B(n37896), .Z(n37892) );
  ANDN U38153 ( .B(B[151]), .A(n73), .Z(n37676) );
  XNOR U38154 ( .A(n37684), .B(n37898), .Z(n37677) );
  XNOR U38155 ( .A(n37683), .B(n37681), .Z(n37898) );
  AND U38156 ( .A(n37899), .B(n37900), .Z(n37681) );
  NANDN U38157 ( .A(n37901), .B(n37902), .Z(n37900) );
  NANDN U38158 ( .A(n37903), .B(n37904), .Z(n37902) );
  NANDN U38159 ( .A(n37904), .B(n37903), .Z(n37899) );
  ANDN U38160 ( .B(B[152]), .A(n74), .Z(n37683) );
  XNOR U38161 ( .A(n37691), .B(n37905), .Z(n37684) );
  XNOR U38162 ( .A(n37690), .B(n37688), .Z(n37905) );
  AND U38163 ( .A(n37906), .B(n37907), .Z(n37688) );
  NANDN U38164 ( .A(n37908), .B(n37909), .Z(n37907) );
  OR U38165 ( .A(n37910), .B(n37911), .Z(n37909) );
  NAND U38166 ( .A(n37911), .B(n37910), .Z(n37906) );
  ANDN U38167 ( .B(B[153]), .A(n75), .Z(n37690) );
  XNOR U38168 ( .A(n37698), .B(n37912), .Z(n37691) );
  XNOR U38169 ( .A(n37697), .B(n37695), .Z(n37912) );
  AND U38170 ( .A(n37913), .B(n37914), .Z(n37695) );
  NANDN U38171 ( .A(n37915), .B(n37916), .Z(n37914) );
  NANDN U38172 ( .A(n37917), .B(n37918), .Z(n37916) );
  NANDN U38173 ( .A(n37918), .B(n37917), .Z(n37913) );
  ANDN U38174 ( .B(B[154]), .A(n76), .Z(n37697) );
  XNOR U38175 ( .A(n37705), .B(n37919), .Z(n37698) );
  XNOR U38176 ( .A(n37704), .B(n37702), .Z(n37919) );
  AND U38177 ( .A(n37920), .B(n37921), .Z(n37702) );
  NANDN U38178 ( .A(n37922), .B(n37923), .Z(n37921) );
  OR U38179 ( .A(n37924), .B(n37925), .Z(n37923) );
  NAND U38180 ( .A(n37925), .B(n37924), .Z(n37920) );
  ANDN U38181 ( .B(B[155]), .A(n77), .Z(n37704) );
  XNOR U38182 ( .A(n37712), .B(n37926), .Z(n37705) );
  XNOR U38183 ( .A(n37711), .B(n37709), .Z(n37926) );
  AND U38184 ( .A(n37927), .B(n37928), .Z(n37709) );
  NANDN U38185 ( .A(n37929), .B(n37930), .Z(n37928) );
  NANDN U38186 ( .A(n37931), .B(n37932), .Z(n37930) );
  NANDN U38187 ( .A(n37932), .B(n37931), .Z(n37927) );
  ANDN U38188 ( .B(B[156]), .A(n78), .Z(n37711) );
  XNOR U38189 ( .A(n37719), .B(n37933), .Z(n37712) );
  XNOR U38190 ( .A(n37718), .B(n37716), .Z(n37933) );
  AND U38191 ( .A(n37934), .B(n37935), .Z(n37716) );
  NANDN U38192 ( .A(n37936), .B(n37937), .Z(n37935) );
  OR U38193 ( .A(n37938), .B(n37939), .Z(n37937) );
  NAND U38194 ( .A(n37939), .B(n37938), .Z(n37934) );
  ANDN U38195 ( .B(B[157]), .A(n79), .Z(n37718) );
  XNOR U38196 ( .A(n37726), .B(n37940), .Z(n37719) );
  XNOR U38197 ( .A(n37725), .B(n37723), .Z(n37940) );
  AND U38198 ( .A(n37941), .B(n37942), .Z(n37723) );
  NANDN U38199 ( .A(n37943), .B(n37944), .Z(n37942) );
  NANDN U38200 ( .A(n37945), .B(n37946), .Z(n37944) );
  NANDN U38201 ( .A(n37946), .B(n37945), .Z(n37941) );
  ANDN U38202 ( .B(B[158]), .A(n80), .Z(n37725) );
  XNOR U38203 ( .A(n37733), .B(n37947), .Z(n37726) );
  XNOR U38204 ( .A(n37732), .B(n37730), .Z(n37947) );
  AND U38205 ( .A(n37948), .B(n37949), .Z(n37730) );
  NANDN U38206 ( .A(n37950), .B(n37951), .Z(n37949) );
  OR U38207 ( .A(n37952), .B(n37953), .Z(n37951) );
  NAND U38208 ( .A(n37953), .B(n37952), .Z(n37948) );
  ANDN U38209 ( .B(B[159]), .A(n81), .Z(n37732) );
  XNOR U38210 ( .A(n37740), .B(n37954), .Z(n37733) );
  XNOR U38211 ( .A(n37739), .B(n37737), .Z(n37954) );
  AND U38212 ( .A(n37955), .B(n37956), .Z(n37737) );
  NANDN U38213 ( .A(n37957), .B(n37958), .Z(n37956) );
  NAND U38214 ( .A(n37959), .B(n37960), .Z(n37958) );
  ANDN U38215 ( .B(B[160]), .A(n82), .Z(n37739) );
  XOR U38216 ( .A(n37746), .B(n37961), .Z(n37740) );
  XNOR U38217 ( .A(n37744), .B(n37747), .Z(n37961) );
  NAND U38218 ( .A(A[2]), .B(B[161]), .Z(n37747) );
  NANDN U38219 ( .A(n37962), .B(n37963), .Z(n37744) );
  AND U38220 ( .A(A[0]), .B(B[162]), .Z(n37963) );
  XNOR U38221 ( .A(n37749), .B(n37964), .Z(n37746) );
  NAND U38222 ( .A(A[0]), .B(B[163]), .Z(n37964) );
  NAND U38223 ( .A(B[162]), .B(A[1]), .Z(n37749) );
  NAND U38224 ( .A(n37965), .B(n37966), .Z(n470) );
  NANDN U38225 ( .A(n37967), .B(n37968), .Z(n37966) );
  OR U38226 ( .A(n37969), .B(n37970), .Z(n37968) );
  NAND U38227 ( .A(n37970), .B(n37969), .Z(n37965) );
  XOR U38228 ( .A(n472), .B(n471), .Z(\A1[160] ) );
  XOR U38229 ( .A(n37970), .B(n37971), .Z(n471) );
  XNOR U38230 ( .A(n37969), .B(n37967), .Z(n37971) );
  AND U38231 ( .A(n37972), .B(n37973), .Z(n37967) );
  NANDN U38232 ( .A(n37974), .B(n37975), .Z(n37973) );
  NANDN U38233 ( .A(n37976), .B(n37977), .Z(n37975) );
  NANDN U38234 ( .A(n37977), .B(n37976), .Z(n37972) );
  ANDN U38235 ( .B(B[131]), .A(n54), .Z(n37969) );
  XNOR U38236 ( .A(n37764), .B(n37978), .Z(n37970) );
  XNOR U38237 ( .A(n37763), .B(n37761), .Z(n37978) );
  AND U38238 ( .A(n37979), .B(n37980), .Z(n37761) );
  NANDN U38239 ( .A(n37981), .B(n37982), .Z(n37980) );
  OR U38240 ( .A(n37983), .B(n37984), .Z(n37982) );
  NAND U38241 ( .A(n37984), .B(n37983), .Z(n37979) );
  ANDN U38242 ( .B(B[132]), .A(n55), .Z(n37763) );
  XNOR U38243 ( .A(n37771), .B(n37985), .Z(n37764) );
  XNOR U38244 ( .A(n37770), .B(n37768), .Z(n37985) );
  AND U38245 ( .A(n37986), .B(n37987), .Z(n37768) );
  NANDN U38246 ( .A(n37988), .B(n37989), .Z(n37987) );
  NANDN U38247 ( .A(n37990), .B(n37991), .Z(n37989) );
  NANDN U38248 ( .A(n37991), .B(n37990), .Z(n37986) );
  ANDN U38249 ( .B(B[133]), .A(n56), .Z(n37770) );
  XNOR U38250 ( .A(n37778), .B(n37992), .Z(n37771) );
  XNOR U38251 ( .A(n37777), .B(n37775), .Z(n37992) );
  AND U38252 ( .A(n37993), .B(n37994), .Z(n37775) );
  NANDN U38253 ( .A(n37995), .B(n37996), .Z(n37994) );
  OR U38254 ( .A(n37997), .B(n37998), .Z(n37996) );
  NAND U38255 ( .A(n37998), .B(n37997), .Z(n37993) );
  ANDN U38256 ( .B(B[134]), .A(n57), .Z(n37777) );
  XNOR U38257 ( .A(n37785), .B(n37999), .Z(n37778) );
  XNOR U38258 ( .A(n37784), .B(n37782), .Z(n37999) );
  AND U38259 ( .A(n38000), .B(n38001), .Z(n37782) );
  NANDN U38260 ( .A(n38002), .B(n38003), .Z(n38001) );
  NANDN U38261 ( .A(n38004), .B(n38005), .Z(n38003) );
  NANDN U38262 ( .A(n38005), .B(n38004), .Z(n38000) );
  ANDN U38263 ( .B(B[135]), .A(n58), .Z(n37784) );
  XNOR U38264 ( .A(n37792), .B(n38006), .Z(n37785) );
  XNOR U38265 ( .A(n37791), .B(n37789), .Z(n38006) );
  AND U38266 ( .A(n38007), .B(n38008), .Z(n37789) );
  NANDN U38267 ( .A(n38009), .B(n38010), .Z(n38008) );
  OR U38268 ( .A(n38011), .B(n38012), .Z(n38010) );
  NAND U38269 ( .A(n38012), .B(n38011), .Z(n38007) );
  ANDN U38270 ( .B(B[136]), .A(n59), .Z(n37791) );
  XNOR U38271 ( .A(n37799), .B(n38013), .Z(n37792) );
  XNOR U38272 ( .A(n37798), .B(n37796), .Z(n38013) );
  AND U38273 ( .A(n38014), .B(n38015), .Z(n37796) );
  NANDN U38274 ( .A(n38016), .B(n38017), .Z(n38015) );
  NANDN U38275 ( .A(n38018), .B(n38019), .Z(n38017) );
  NANDN U38276 ( .A(n38019), .B(n38018), .Z(n38014) );
  ANDN U38277 ( .B(B[137]), .A(n60), .Z(n37798) );
  XNOR U38278 ( .A(n37806), .B(n38020), .Z(n37799) );
  XNOR U38279 ( .A(n37805), .B(n37803), .Z(n38020) );
  AND U38280 ( .A(n38021), .B(n38022), .Z(n37803) );
  NANDN U38281 ( .A(n38023), .B(n38024), .Z(n38022) );
  OR U38282 ( .A(n38025), .B(n38026), .Z(n38024) );
  NAND U38283 ( .A(n38026), .B(n38025), .Z(n38021) );
  ANDN U38284 ( .B(B[138]), .A(n61), .Z(n37805) );
  XNOR U38285 ( .A(n37813), .B(n38027), .Z(n37806) );
  XNOR U38286 ( .A(n37812), .B(n37810), .Z(n38027) );
  AND U38287 ( .A(n38028), .B(n38029), .Z(n37810) );
  NANDN U38288 ( .A(n38030), .B(n38031), .Z(n38029) );
  NANDN U38289 ( .A(n38032), .B(n38033), .Z(n38031) );
  NANDN U38290 ( .A(n38033), .B(n38032), .Z(n38028) );
  ANDN U38291 ( .B(B[139]), .A(n62), .Z(n37812) );
  XNOR U38292 ( .A(n37820), .B(n38034), .Z(n37813) );
  XNOR U38293 ( .A(n37819), .B(n37817), .Z(n38034) );
  AND U38294 ( .A(n38035), .B(n38036), .Z(n37817) );
  NANDN U38295 ( .A(n38037), .B(n38038), .Z(n38036) );
  OR U38296 ( .A(n38039), .B(n38040), .Z(n38038) );
  NAND U38297 ( .A(n38040), .B(n38039), .Z(n38035) );
  ANDN U38298 ( .B(B[140]), .A(n63), .Z(n37819) );
  XNOR U38299 ( .A(n37827), .B(n38041), .Z(n37820) );
  XNOR U38300 ( .A(n37826), .B(n37824), .Z(n38041) );
  AND U38301 ( .A(n38042), .B(n38043), .Z(n37824) );
  NANDN U38302 ( .A(n38044), .B(n38045), .Z(n38043) );
  NANDN U38303 ( .A(n38046), .B(n38047), .Z(n38045) );
  NANDN U38304 ( .A(n38047), .B(n38046), .Z(n38042) );
  ANDN U38305 ( .B(B[141]), .A(n64), .Z(n37826) );
  XNOR U38306 ( .A(n37834), .B(n38048), .Z(n37827) );
  XNOR U38307 ( .A(n37833), .B(n37831), .Z(n38048) );
  AND U38308 ( .A(n38049), .B(n38050), .Z(n37831) );
  NANDN U38309 ( .A(n38051), .B(n38052), .Z(n38050) );
  OR U38310 ( .A(n38053), .B(n38054), .Z(n38052) );
  NAND U38311 ( .A(n38054), .B(n38053), .Z(n38049) );
  ANDN U38312 ( .B(B[142]), .A(n65), .Z(n37833) );
  XNOR U38313 ( .A(n37841), .B(n38055), .Z(n37834) );
  XNOR U38314 ( .A(n37840), .B(n37838), .Z(n38055) );
  AND U38315 ( .A(n38056), .B(n38057), .Z(n37838) );
  NANDN U38316 ( .A(n38058), .B(n38059), .Z(n38057) );
  NANDN U38317 ( .A(n38060), .B(n38061), .Z(n38059) );
  NANDN U38318 ( .A(n38061), .B(n38060), .Z(n38056) );
  ANDN U38319 ( .B(B[143]), .A(n66), .Z(n37840) );
  XNOR U38320 ( .A(n37848), .B(n38062), .Z(n37841) );
  XNOR U38321 ( .A(n37847), .B(n37845), .Z(n38062) );
  AND U38322 ( .A(n38063), .B(n38064), .Z(n37845) );
  NANDN U38323 ( .A(n38065), .B(n38066), .Z(n38064) );
  OR U38324 ( .A(n38067), .B(n38068), .Z(n38066) );
  NAND U38325 ( .A(n38068), .B(n38067), .Z(n38063) );
  ANDN U38326 ( .B(B[144]), .A(n67), .Z(n37847) );
  XNOR U38327 ( .A(n37855), .B(n38069), .Z(n37848) );
  XNOR U38328 ( .A(n37854), .B(n37852), .Z(n38069) );
  AND U38329 ( .A(n38070), .B(n38071), .Z(n37852) );
  NANDN U38330 ( .A(n38072), .B(n38073), .Z(n38071) );
  NANDN U38331 ( .A(n38074), .B(n38075), .Z(n38073) );
  NANDN U38332 ( .A(n38075), .B(n38074), .Z(n38070) );
  ANDN U38333 ( .B(B[145]), .A(n68), .Z(n37854) );
  XNOR U38334 ( .A(n37862), .B(n38076), .Z(n37855) );
  XNOR U38335 ( .A(n37861), .B(n37859), .Z(n38076) );
  AND U38336 ( .A(n38077), .B(n38078), .Z(n37859) );
  NANDN U38337 ( .A(n38079), .B(n38080), .Z(n38078) );
  OR U38338 ( .A(n38081), .B(n38082), .Z(n38080) );
  NAND U38339 ( .A(n38082), .B(n38081), .Z(n38077) );
  ANDN U38340 ( .B(B[146]), .A(n69), .Z(n37861) );
  XNOR U38341 ( .A(n37869), .B(n38083), .Z(n37862) );
  XNOR U38342 ( .A(n37868), .B(n37866), .Z(n38083) );
  AND U38343 ( .A(n38084), .B(n38085), .Z(n37866) );
  NANDN U38344 ( .A(n38086), .B(n38087), .Z(n38085) );
  NANDN U38345 ( .A(n38088), .B(n38089), .Z(n38087) );
  NANDN U38346 ( .A(n38089), .B(n38088), .Z(n38084) );
  ANDN U38347 ( .B(B[147]), .A(n70), .Z(n37868) );
  XNOR U38348 ( .A(n37876), .B(n38090), .Z(n37869) );
  XNOR U38349 ( .A(n37875), .B(n37873), .Z(n38090) );
  AND U38350 ( .A(n38091), .B(n38092), .Z(n37873) );
  NANDN U38351 ( .A(n38093), .B(n38094), .Z(n38092) );
  OR U38352 ( .A(n38095), .B(n38096), .Z(n38094) );
  NAND U38353 ( .A(n38096), .B(n38095), .Z(n38091) );
  ANDN U38354 ( .B(B[148]), .A(n71), .Z(n37875) );
  XNOR U38355 ( .A(n37883), .B(n38097), .Z(n37876) );
  XNOR U38356 ( .A(n37882), .B(n37880), .Z(n38097) );
  AND U38357 ( .A(n38098), .B(n38099), .Z(n37880) );
  NANDN U38358 ( .A(n38100), .B(n38101), .Z(n38099) );
  NANDN U38359 ( .A(n38102), .B(n38103), .Z(n38101) );
  NANDN U38360 ( .A(n38103), .B(n38102), .Z(n38098) );
  ANDN U38361 ( .B(B[149]), .A(n72), .Z(n37882) );
  XNOR U38362 ( .A(n37890), .B(n38104), .Z(n37883) );
  XNOR U38363 ( .A(n37889), .B(n37887), .Z(n38104) );
  AND U38364 ( .A(n38105), .B(n38106), .Z(n37887) );
  NANDN U38365 ( .A(n38107), .B(n38108), .Z(n38106) );
  OR U38366 ( .A(n38109), .B(n38110), .Z(n38108) );
  NAND U38367 ( .A(n38110), .B(n38109), .Z(n38105) );
  ANDN U38368 ( .B(B[150]), .A(n73), .Z(n37889) );
  XNOR U38369 ( .A(n37897), .B(n38111), .Z(n37890) );
  XNOR U38370 ( .A(n37896), .B(n37894), .Z(n38111) );
  AND U38371 ( .A(n38112), .B(n38113), .Z(n37894) );
  NANDN U38372 ( .A(n38114), .B(n38115), .Z(n38113) );
  NANDN U38373 ( .A(n38116), .B(n38117), .Z(n38115) );
  NANDN U38374 ( .A(n38117), .B(n38116), .Z(n38112) );
  ANDN U38375 ( .B(B[151]), .A(n74), .Z(n37896) );
  XNOR U38376 ( .A(n37904), .B(n38118), .Z(n37897) );
  XNOR U38377 ( .A(n37903), .B(n37901), .Z(n38118) );
  AND U38378 ( .A(n38119), .B(n38120), .Z(n37901) );
  NANDN U38379 ( .A(n38121), .B(n38122), .Z(n38120) );
  OR U38380 ( .A(n38123), .B(n38124), .Z(n38122) );
  NAND U38381 ( .A(n38124), .B(n38123), .Z(n38119) );
  ANDN U38382 ( .B(B[152]), .A(n75), .Z(n37903) );
  XNOR U38383 ( .A(n37911), .B(n38125), .Z(n37904) );
  XNOR U38384 ( .A(n37910), .B(n37908), .Z(n38125) );
  AND U38385 ( .A(n38126), .B(n38127), .Z(n37908) );
  NANDN U38386 ( .A(n38128), .B(n38129), .Z(n38127) );
  NANDN U38387 ( .A(n38130), .B(n38131), .Z(n38129) );
  NANDN U38388 ( .A(n38131), .B(n38130), .Z(n38126) );
  ANDN U38389 ( .B(B[153]), .A(n76), .Z(n37910) );
  XNOR U38390 ( .A(n37918), .B(n38132), .Z(n37911) );
  XNOR U38391 ( .A(n37917), .B(n37915), .Z(n38132) );
  AND U38392 ( .A(n38133), .B(n38134), .Z(n37915) );
  NANDN U38393 ( .A(n38135), .B(n38136), .Z(n38134) );
  OR U38394 ( .A(n38137), .B(n38138), .Z(n38136) );
  NAND U38395 ( .A(n38138), .B(n38137), .Z(n38133) );
  ANDN U38396 ( .B(B[154]), .A(n77), .Z(n37917) );
  XNOR U38397 ( .A(n37925), .B(n38139), .Z(n37918) );
  XNOR U38398 ( .A(n37924), .B(n37922), .Z(n38139) );
  AND U38399 ( .A(n38140), .B(n38141), .Z(n37922) );
  NANDN U38400 ( .A(n38142), .B(n38143), .Z(n38141) );
  NANDN U38401 ( .A(n38144), .B(n38145), .Z(n38143) );
  NANDN U38402 ( .A(n38145), .B(n38144), .Z(n38140) );
  ANDN U38403 ( .B(B[155]), .A(n78), .Z(n37924) );
  XNOR U38404 ( .A(n37932), .B(n38146), .Z(n37925) );
  XNOR U38405 ( .A(n37931), .B(n37929), .Z(n38146) );
  AND U38406 ( .A(n38147), .B(n38148), .Z(n37929) );
  NANDN U38407 ( .A(n38149), .B(n38150), .Z(n38148) );
  OR U38408 ( .A(n38151), .B(n38152), .Z(n38150) );
  NAND U38409 ( .A(n38152), .B(n38151), .Z(n38147) );
  ANDN U38410 ( .B(B[156]), .A(n79), .Z(n37931) );
  XNOR U38411 ( .A(n37939), .B(n38153), .Z(n37932) );
  XNOR U38412 ( .A(n37938), .B(n37936), .Z(n38153) );
  AND U38413 ( .A(n38154), .B(n38155), .Z(n37936) );
  NANDN U38414 ( .A(n38156), .B(n38157), .Z(n38155) );
  NANDN U38415 ( .A(n38158), .B(n38159), .Z(n38157) );
  NANDN U38416 ( .A(n38159), .B(n38158), .Z(n38154) );
  ANDN U38417 ( .B(B[157]), .A(n80), .Z(n37938) );
  XNOR U38418 ( .A(n37946), .B(n38160), .Z(n37939) );
  XNOR U38419 ( .A(n37945), .B(n37943), .Z(n38160) );
  AND U38420 ( .A(n38161), .B(n38162), .Z(n37943) );
  NANDN U38421 ( .A(n38163), .B(n38164), .Z(n38162) );
  OR U38422 ( .A(n38165), .B(n38166), .Z(n38164) );
  NAND U38423 ( .A(n38166), .B(n38165), .Z(n38161) );
  ANDN U38424 ( .B(B[158]), .A(n81), .Z(n37945) );
  XNOR U38425 ( .A(n37953), .B(n38167), .Z(n37946) );
  XNOR U38426 ( .A(n37952), .B(n37950), .Z(n38167) );
  AND U38427 ( .A(n38168), .B(n38169), .Z(n37950) );
  NANDN U38428 ( .A(n38170), .B(n38171), .Z(n38169) );
  NAND U38429 ( .A(n38172), .B(n38173), .Z(n38171) );
  ANDN U38430 ( .B(B[159]), .A(n82), .Z(n37952) );
  XOR U38431 ( .A(n37959), .B(n38174), .Z(n37953) );
  XNOR U38432 ( .A(n37957), .B(n37960), .Z(n38174) );
  NAND U38433 ( .A(A[2]), .B(B[160]), .Z(n37960) );
  NANDN U38434 ( .A(n38175), .B(n38176), .Z(n37957) );
  AND U38435 ( .A(A[0]), .B(B[161]), .Z(n38176) );
  XNOR U38436 ( .A(n37962), .B(n38177), .Z(n37959) );
  NAND U38437 ( .A(A[0]), .B(B[162]), .Z(n38177) );
  NAND U38438 ( .A(B[161]), .B(A[1]), .Z(n37962) );
  NAND U38439 ( .A(n38178), .B(n38179), .Z(n472) );
  NANDN U38440 ( .A(n38180), .B(n38181), .Z(n38179) );
  OR U38441 ( .A(n38182), .B(n38183), .Z(n38181) );
  NAND U38442 ( .A(n38183), .B(n38182), .Z(n38178) );
  XOR U38443 ( .A(n35944), .B(n38184), .Z(\A1[15] ) );
  XNOR U38444 ( .A(n35943), .B(n35941), .Z(n38184) );
  AND U38445 ( .A(n38185), .B(n38186), .Z(n35941) );
  NAND U38446 ( .A(n38187), .B(n38188), .Z(n38186) );
  NANDN U38447 ( .A(n38189), .B(n38190), .Z(n38187) );
  NANDN U38448 ( .A(n38190), .B(n38189), .Z(n38185) );
  ANDN U38449 ( .B(B[0]), .A(n68), .Z(n35943) );
  XNOR U38450 ( .A(n35951), .B(n38191), .Z(n35944) );
  XNOR U38451 ( .A(n35950), .B(n35948), .Z(n38191) );
  AND U38452 ( .A(n38192), .B(n38193), .Z(n35948) );
  NANDN U38453 ( .A(n38194), .B(n38195), .Z(n38193) );
  OR U38454 ( .A(n38196), .B(n38197), .Z(n38195) );
  NAND U38455 ( .A(n38197), .B(n38196), .Z(n38192) );
  ANDN U38456 ( .B(B[1]), .A(n69), .Z(n35950) );
  XNOR U38457 ( .A(n35958), .B(n38198), .Z(n35951) );
  XNOR U38458 ( .A(n35957), .B(n35955), .Z(n38198) );
  AND U38459 ( .A(n38199), .B(n38200), .Z(n35955) );
  NANDN U38460 ( .A(n38201), .B(n38202), .Z(n38200) );
  NANDN U38461 ( .A(n38203), .B(n38204), .Z(n38202) );
  NANDN U38462 ( .A(n38204), .B(n38203), .Z(n38199) );
  ANDN U38463 ( .B(B[2]), .A(n70), .Z(n35957) );
  XNOR U38464 ( .A(n35965), .B(n38205), .Z(n35958) );
  XNOR U38465 ( .A(n35964), .B(n35962), .Z(n38205) );
  AND U38466 ( .A(n38206), .B(n38207), .Z(n35962) );
  NANDN U38467 ( .A(n38208), .B(n38209), .Z(n38207) );
  OR U38468 ( .A(n38210), .B(n38211), .Z(n38209) );
  NAND U38469 ( .A(n38211), .B(n38210), .Z(n38206) );
  ANDN U38470 ( .B(B[3]), .A(n71), .Z(n35964) );
  XNOR U38471 ( .A(n35972), .B(n38212), .Z(n35965) );
  XNOR U38472 ( .A(n35971), .B(n35969), .Z(n38212) );
  AND U38473 ( .A(n38213), .B(n38214), .Z(n35969) );
  NANDN U38474 ( .A(n38215), .B(n38216), .Z(n38214) );
  NANDN U38475 ( .A(n38217), .B(n38218), .Z(n38216) );
  NANDN U38476 ( .A(n38218), .B(n38217), .Z(n38213) );
  ANDN U38477 ( .B(B[4]), .A(n72), .Z(n35971) );
  XNOR U38478 ( .A(n35979), .B(n38219), .Z(n35972) );
  XNOR U38479 ( .A(n35978), .B(n35976), .Z(n38219) );
  AND U38480 ( .A(n38220), .B(n38221), .Z(n35976) );
  NANDN U38481 ( .A(n38222), .B(n38223), .Z(n38221) );
  OR U38482 ( .A(n38224), .B(n38225), .Z(n38223) );
  NAND U38483 ( .A(n38225), .B(n38224), .Z(n38220) );
  ANDN U38484 ( .B(B[5]), .A(n73), .Z(n35978) );
  XNOR U38485 ( .A(n35986), .B(n38226), .Z(n35979) );
  XNOR U38486 ( .A(n35985), .B(n35983), .Z(n38226) );
  AND U38487 ( .A(n38227), .B(n38228), .Z(n35983) );
  NANDN U38488 ( .A(n38229), .B(n38230), .Z(n38228) );
  NANDN U38489 ( .A(n38231), .B(n38232), .Z(n38230) );
  NANDN U38490 ( .A(n38232), .B(n38231), .Z(n38227) );
  ANDN U38491 ( .B(B[6]), .A(n74), .Z(n35985) );
  XNOR U38492 ( .A(n35993), .B(n38233), .Z(n35986) );
  XNOR U38493 ( .A(n35992), .B(n35990), .Z(n38233) );
  AND U38494 ( .A(n38234), .B(n38235), .Z(n35990) );
  NANDN U38495 ( .A(n38236), .B(n38237), .Z(n38235) );
  OR U38496 ( .A(n38238), .B(n38239), .Z(n38237) );
  NAND U38497 ( .A(n38239), .B(n38238), .Z(n38234) );
  ANDN U38498 ( .B(B[7]), .A(n75), .Z(n35992) );
  XNOR U38499 ( .A(n36000), .B(n38240), .Z(n35993) );
  XNOR U38500 ( .A(n35999), .B(n35997), .Z(n38240) );
  AND U38501 ( .A(n38241), .B(n38242), .Z(n35997) );
  NANDN U38502 ( .A(n38243), .B(n38244), .Z(n38242) );
  NANDN U38503 ( .A(n38245), .B(n38246), .Z(n38244) );
  NANDN U38504 ( .A(n38246), .B(n38245), .Z(n38241) );
  ANDN U38505 ( .B(B[8]), .A(n76), .Z(n35999) );
  XNOR U38506 ( .A(n36007), .B(n38247), .Z(n36000) );
  XNOR U38507 ( .A(n36006), .B(n36004), .Z(n38247) );
  AND U38508 ( .A(n38248), .B(n38249), .Z(n36004) );
  NANDN U38509 ( .A(n38250), .B(n38251), .Z(n38249) );
  OR U38510 ( .A(n38252), .B(n38253), .Z(n38251) );
  NAND U38511 ( .A(n38253), .B(n38252), .Z(n38248) );
  ANDN U38512 ( .B(B[9]), .A(n77), .Z(n36006) );
  XNOR U38513 ( .A(n36014), .B(n38254), .Z(n36007) );
  XNOR U38514 ( .A(n36013), .B(n36011), .Z(n38254) );
  AND U38515 ( .A(n38255), .B(n38256), .Z(n36011) );
  NANDN U38516 ( .A(n38257), .B(n38258), .Z(n38256) );
  NANDN U38517 ( .A(n38259), .B(n38260), .Z(n38258) );
  NANDN U38518 ( .A(n38260), .B(n38259), .Z(n38255) );
  ANDN U38519 ( .B(B[10]), .A(n78), .Z(n36013) );
  XNOR U38520 ( .A(n36021), .B(n38261), .Z(n36014) );
  XNOR U38521 ( .A(n36020), .B(n36018), .Z(n38261) );
  AND U38522 ( .A(n38262), .B(n38263), .Z(n36018) );
  NANDN U38523 ( .A(n38264), .B(n38265), .Z(n38263) );
  OR U38524 ( .A(n38266), .B(n38267), .Z(n38265) );
  NAND U38525 ( .A(n38267), .B(n38266), .Z(n38262) );
  ANDN U38526 ( .B(B[11]), .A(n79), .Z(n36020) );
  XNOR U38527 ( .A(n36028), .B(n38268), .Z(n36021) );
  XNOR U38528 ( .A(n36027), .B(n36025), .Z(n38268) );
  AND U38529 ( .A(n38269), .B(n38270), .Z(n36025) );
  NANDN U38530 ( .A(n38271), .B(n38272), .Z(n38270) );
  NANDN U38531 ( .A(n38273), .B(n38274), .Z(n38272) );
  NANDN U38532 ( .A(n38274), .B(n38273), .Z(n38269) );
  ANDN U38533 ( .B(B[12]), .A(n80), .Z(n36027) );
  XNOR U38534 ( .A(n36035), .B(n38275), .Z(n36028) );
  XNOR U38535 ( .A(n36034), .B(n36032), .Z(n38275) );
  AND U38536 ( .A(n38276), .B(n38277), .Z(n36032) );
  NANDN U38537 ( .A(n38278), .B(n38279), .Z(n38277) );
  OR U38538 ( .A(n38280), .B(n38281), .Z(n38279) );
  NAND U38539 ( .A(n38281), .B(n38280), .Z(n38276) );
  ANDN U38540 ( .B(B[13]), .A(n81), .Z(n36034) );
  XNOR U38541 ( .A(n36042), .B(n38282), .Z(n36035) );
  XNOR U38542 ( .A(n36041), .B(n36039), .Z(n38282) );
  AND U38543 ( .A(n38283), .B(n38284), .Z(n36039) );
  NANDN U38544 ( .A(n38285), .B(n38286), .Z(n38284) );
  NAND U38545 ( .A(n38287), .B(n38288), .Z(n38286) );
  ANDN U38546 ( .B(B[14]), .A(n82), .Z(n36041) );
  XOR U38547 ( .A(n36048), .B(n38289), .Z(n36042) );
  XNOR U38548 ( .A(n36046), .B(n36049), .Z(n38289) );
  NAND U38549 ( .A(A[2]), .B(B[15]), .Z(n36049) );
  NANDN U38550 ( .A(n38290), .B(n38291), .Z(n36046) );
  AND U38551 ( .A(A[0]), .B(B[16]), .Z(n38291) );
  XNOR U38552 ( .A(n36051), .B(n38292), .Z(n36048) );
  NAND U38553 ( .A(A[0]), .B(B[17]), .Z(n38292) );
  NAND U38554 ( .A(B[16]), .B(A[1]), .Z(n36051) );
  XOR U38555 ( .A(n474), .B(n473), .Z(\A1[159] ) );
  XOR U38556 ( .A(n38183), .B(n38293), .Z(n473) );
  XNOR U38557 ( .A(n38182), .B(n38180), .Z(n38293) );
  AND U38558 ( .A(n38294), .B(n38295), .Z(n38180) );
  NANDN U38559 ( .A(n38296), .B(n38297), .Z(n38295) );
  NANDN U38560 ( .A(n38298), .B(n38299), .Z(n38297) );
  NANDN U38561 ( .A(n38299), .B(n38298), .Z(n38294) );
  ANDN U38562 ( .B(B[130]), .A(n54), .Z(n38182) );
  XNOR U38563 ( .A(n37977), .B(n38300), .Z(n38183) );
  XNOR U38564 ( .A(n37976), .B(n37974), .Z(n38300) );
  AND U38565 ( .A(n38301), .B(n38302), .Z(n37974) );
  NANDN U38566 ( .A(n38303), .B(n38304), .Z(n38302) );
  OR U38567 ( .A(n38305), .B(n38306), .Z(n38304) );
  NAND U38568 ( .A(n38306), .B(n38305), .Z(n38301) );
  ANDN U38569 ( .B(B[131]), .A(n55), .Z(n37976) );
  XNOR U38570 ( .A(n37984), .B(n38307), .Z(n37977) );
  XNOR U38571 ( .A(n37983), .B(n37981), .Z(n38307) );
  AND U38572 ( .A(n38308), .B(n38309), .Z(n37981) );
  NANDN U38573 ( .A(n38310), .B(n38311), .Z(n38309) );
  NANDN U38574 ( .A(n38312), .B(n38313), .Z(n38311) );
  NANDN U38575 ( .A(n38313), .B(n38312), .Z(n38308) );
  ANDN U38576 ( .B(B[132]), .A(n56), .Z(n37983) );
  XNOR U38577 ( .A(n37991), .B(n38314), .Z(n37984) );
  XNOR U38578 ( .A(n37990), .B(n37988), .Z(n38314) );
  AND U38579 ( .A(n38315), .B(n38316), .Z(n37988) );
  NANDN U38580 ( .A(n38317), .B(n38318), .Z(n38316) );
  OR U38581 ( .A(n38319), .B(n38320), .Z(n38318) );
  NAND U38582 ( .A(n38320), .B(n38319), .Z(n38315) );
  ANDN U38583 ( .B(B[133]), .A(n57), .Z(n37990) );
  XNOR U38584 ( .A(n37998), .B(n38321), .Z(n37991) );
  XNOR U38585 ( .A(n37997), .B(n37995), .Z(n38321) );
  AND U38586 ( .A(n38322), .B(n38323), .Z(n37995) );
  NANDN U38587 ( .A(n38324), .B(n38325), .Z(n38323) );
  NANDN U38588 ( .A(n38326), .B(n38327), .Z(n38325) );
  NANDN U38589 ( .A(n38327), .B(n38326), .Z(n38322) );
  ANDN U38590 ( .B(B[134]), .A(n58), .Z(n37997) );
  XNOR U38591 ( .A(n38005), .B(n38328), .Z(n37998) );
  XNOR U38592 ( .A(n38004), .B(n38002), .Z(n38328) );
  AND U38593 ( .A(n38329), .B(n38330), .Z(n38002) );
  NANDN U38594 ( .A(n38331), .B(n38332), .Z(n38330) );
  OR U38595 ( .A(n38333), .B(n38334), .Z(n38332) );
  NAND U38596 ( .A(n38334), .B(n38333), .Z(n38329) );
  ANDN U38597 ( .B(B[135]), .A(n59), .Z(n38004) );
  XNOR U38598 ( .A(n38012), .B(n38335), .Z(n38005) );
  XNOR U38599 ( .A(n38011), .B(n38009), .Z(n38335) );
  AND U38600 ( .A(n38336), .B(n38337), .Z(n38009) );
  NANDN U38601 ( .A(n38338), .B(n38339), .Z(n38337) );
  NANDN U38602 ( .A(n38340), .B(n38341), .Z(n38339) );
  NANDN U38603 ( .A(n38341), .B(n38340), .Z(n38336) );
  ANDN U38604 ( .B(B[136]), .A(n60), .Z(n38011) );
  XNOR U38605 ( .A(n38019), .B(n38342), .Z(n38012) );
  XNOR U38606 ( .A(n38018), .B(n38016), .Z(n38342) );
  AND U38607 ( .A(n38343), .B(n38344), .Z(n38016) );
  NANDN U38608 ( .A(n38345), .B(n38346), .Z(n38344) );
  OR U38609 ( .A(n38347), .B(n38348), .Z(n38346) );
  NAND U38610 ( .A(n38348), .B(n38347), .Z(n38343) );
  ANDN U38611 ( .B(B[137]), .A(n61), .Z(n38018) );
  XNOR U38612 ( .A(n38026), .B(n38349), .Z(n38019) );
  XNOR U38613 ( .A(n38025), .B(n38023), .Z(n38349) );
  AND U38614 ( .A(n38350), .B(n38351), .Z(n38023) );
  NANDN U38615 ( .A(n38352), .B(n38353), .Z(n38351) );
  NANDN U38616 ( .A(n38354), .B(n38355), .Z(n38353) );
  NANDN U38617 ( .A(n38355), .B(n38354), .Z(n38350) );
  ANDN U38618 ( .B(B[138]), .A(n62), .Z(n38025) );
  XNOR U38619 ( .A(n38033), .B(n38356), .Z(n38026) );
  XNOR U38620 ( .A(n38032), .B(n38030), .Z(n38356) );
  AND U38621 ( .A(n38357), .B(n38358), .Z(n38030) );
  NANDN U38622 ( .A(n38359), .B(n38360), .Z(n38358) );
  OR U38623 ( .A(n38361), .B(n38362), .Z(n38360) );
  NAND U38624 ( .A(n38362), .B(n38361), .Z(n38357) );
  ANDN U38625 ( .B(B[139]), .A(n63), .Z(n38032) );
  XNOR U38626 ( .A(n38040), .B(n38363), .Z(n38033) );
  XNOR U38627 ( .A(n38039), .B(n38037), .Z(n38363) );
  AND U38628 ( .A(n38364), .B(n38365), .Z(n38037) );
  NANDN U38629 ( .A(n38366), .B(n38367), .Z(n38365) );
  NANDN U38630 ( .A(n38368), .B(n38369), .Z(n38367) );
  NANDN U38631 ( .A(n38369), .B(n38368), .Z(n38364) );
  ANDN U38632 ( .B(B[140]), .A(n64), .Z(n38039) );
  XNOR U38633 ( .A(n38047), .B(n38370), .Z(n38040) );
  XNOR U38634 ( .A(n38046), .B(n38044), .Z(n38370) );
  AND U38635 ( .A(n38371), .B(n38372), .Z(n38044) );
  NANDN U38636 ( .A(n38373), .B(n38374), .Z(n38372) );
  OR U38637 ( .A(n38375), .B(n38376), .Z(n38374) );
  NAND U38638 ( .A(n38376), .B(n38375), .Z(n38371) );
  ANDN U38639 ( .B(B[141]), .A(n65), .Z(n38046) );
  XNOR U38640 ( .A(n38054), .B(n38377), .Z(n38047) );
  XNOR U38641 ( .A(n38053), .B(n38051), .Z(n38377) );
  AND U38642 ( .A(n38378), .B(n38379), .Z(n38051) );
  NANDN U38643 ( .A(n38380), .B(n38381), .Z(n38379) );
  NANDN U38644 ( .A(n38382), .B(n38383), .Z(n38381) );
  NANDN U38645 ( .A(n38383), .B(n38382), .Z(n38378) );
  ANDN U38646 ( .B(B[142]), .A(n66), .Z(n38053) );
  XNOR U38647 ( .A(n38061), .B(n38384), .Z(n38054) );
  XNOR U38648 ( .A(n38060), .B(n38058), .Z(n38384) );
  AND U38649 ( .A(n38385), .B(n38386), .Z(n38058) );
  NANDN U38650 ( .A(n38387), .B(n38388), .Z(n38386) );
  OR U38651 ( .A(n38389), .B(n38390), .Z(n38388) );
  NAND U38652 ( .A(n38390), .B(n38389), .Z(n38385) );
  ANDN U38653 ( .B(B[143]), .A(n67), .Z(n38060) );
  XNOR U38654 ( .A(n38068), .B(n38391), .Z(n38061) );
  XNOR U38655 ( .A(n38067), .B(n38065), .Z(n38391) );
  AND U38656 ( .A(n38392), .B(n38393), .Z(n38065) );
  NANDN U38657 ( .A(n38394), .B(n38395), .Z(n38393) );
  NANDN U38658 ( .A(n38396), .B(n38397), .Z(n38395) );
  NANDN U38659 ( .A(n38397), .B(n38396), .Z(n38392) );
  ANDN U38660 ( .B(B[144]), .A(n68), .Z(n38067) );
  XNOR U38661 ( .A(n38075), .B(n38398), .Z(n38068) );
  XNOR U38662 ( .A(n38074), .B(n38072), .Z(n38398) );
  AND U38663 ( .A(n38399), .B(n38400), .Z(n38072) );
  NANDN U38664 ( .A(n38401), .B(n38402), .Z(n38400) );
  OR U38665 ( .A(n38403), .B(n38404), .Z(n38402) );
  NAND U38666 ( .A(n38404), .B(n38403), .Z(n38399) );
  ANDN U38667 ( .B(B[145]), .A(n69), .Z(n38074) );
  XNOR U38668 ( .A(n38082), .B(n38405), .Z(n38075) );
  XNOR U38669 ( .A(n38081), .B(n38079), .Z(n38405) );
  AND U38670 ( .A(n38406), .B(n38407), .Z(n38079) );
  NANDN U38671 ( .A(n38408), .B(n38409), .Z(n38407) );
  NANDN U38672 ( .A(n38410), .B(n38411), .Z(n38409) );
  NANDN U38673 ( .A(n38411), .B(n38410), .Z(n38406) );
  ANDN U38674 ( .B(B[146]), .A(n70), .Z(n38081) );
  XNOR U38675 ( .A(n38089), .B(n38412), .Z(n38082) );
  XNOR U38676 ( .A(n38088), .B(n38086), .Z(n38412) );
  AND U38677 ( .A(n38413), .B(n38414), .Z(n38086) );
  NANDN U38678 ( .A(n38415), .B(n38416), .Z(n38414) );
  OR U38679 ( .A(n38417), .B(n38418), .Z(n38416) );
  NAND U38680 ( .A(n38418), .B(n38417), .Z(n38413) );
  ANDN U38681 ( .B(B[147]), .A(n71), .Z(n38088) );
  XNOR U38682 ( .A(n38096), .B(n38419), .Z(n38089) );
  XNOR U38683 ( .A(n38095), .B(n38093), .Z(n38419) );
  AND U38684 ( .A(n38420), .B(n38421), .Z(n38093) );
  NANDN U38685 ( .A(n38422), .B(n38423), .Z(n38421) );
  NANDN U38686 ( .A(n38424), .B(n38425), .Z(n38423) );
  NANDN U38687 ( .A(n38425), .B(n38424), .Z(n38420) );
  ANDN U38688 ( .B(B[148]), .A(n72), .Z(n38095) );
  XNOR U38689 ( .A(n38103), .B(n38426), .Z(n38096) );
  XNOR U38690 ( .A(n38102), .B(n38100), .Z(n38426) );
  AND U38691 ( .A(n38427), .B(n38428), .Z(n38100) );
  NANDN U38692 ( .A(n38429), .B(n38430), .Z(n38428) );
  OR U38693 ( .A(n38431), .B(n38432), .Z(n38430) );
  NAND U38694 ( .A(n38432), .B(n38431), .Z(n38427) );
  ANDN U38695 ( .B(B[149]), .A(n73), .Z(n38102) );
  XNOR U38696 ( .A(n38110), .B(n38433), .Z(n38103) );
  XNOR U38697 ( .A(n38109), .B(n38107), .Z(n38433) );
  AND U38698 ( .A(n38434), .B(n38435), .Z(n38107) );
  NANDN U38699 ( .A(n38436), .B(n38437), .Z(n38435) );
  NANDN U38700 ( .A(n38438), .B(n38439), .Z(n38437) );
  NANDN U38701 ( .A(n38439), .B(n38438), .Z(n38434) );
  ANDN U38702 ( .B(B[150]), .A(n74), .Z(n38109) );
  XNOR U38703 ( .A(n38117), .B(n38440), .Z(n38110) );
  XNOR U38704 ( .A(n38116), .B(n38114), .Z(n38440) );
  AND U38705 ( .A(n38441), .B(n38442), .Z(n38114) );
  NANDN U38706 ( .A(n38443), .B(n38444), .Z(n38442) );
  OR U38707 ( .A(n38445), .B(n38446), .Z(n38444) );
  NAND U38708 ( .A(n38446), .B(n38445), .Z(n38441) );
  ANDN U38709 ( .B(B[151]), .A(n75), .Z(n38116) );
  XNOR U38710 ( .A(n38124), .B(n38447), .Z(n38117) );
  XNOR U38711 ( .A(n38123), .B(n38121), .Z(n38447) );
  AND U38712 ( .A(n38448), .B(n38449), .Z(n38121) );
  NANDN U38713 ( .A(n38450), .B(n38451), .Z(n38449) );
  NANDN U38714 ( .A(n38452), .B(n38453), .Z(n38451) );
  NANDN U38715 ( .A(n38453), .B(n38452), .Z(n38448) );
  ANDN U38716 ( .B(B[152]), .A(n76), .Z(n38123) );
  XNOR U38717 ( .A(n38131), .B(n38454), .Z(n38124) );
  XNOR U38718 ( .A(n38130), .B(n38128), .Z(n38454) );
  AND U38719 ( .A(n38455), .B(n38456), .Z(n38128) );
  NANDN U38720 ( .A(n38457), .B(n38458), .Z(n38456) );
  OR U38721 ( .A(n38459), .B(n38460), .Z(n38458) );
  NAND U38722 ( .A(n38460), .B(n38459), .Z(n38455) );
  ANDN U38723 ( .B(B[153]), .A(n77), .Z(n38130) );
  XNOR U38724 ( .A(n38138), .B(n38461), .Z(n38131) );
  XNOR U38725 ( .A(n38137), .B(n38135), .Z(n38461) );
  AND U38726 ( .A(n38462), .B(n38463), .Z(n38135) );
  NANDN U38727 ( .A(n38464), .B(n38465), .Z(n38463) );
  NANDN U38728 ( .A(n38466), .B(n38467), .Z(n38465) );
  NANDN U38729 ( .A(n38467), .B(n38466), .Z(n38462) );
  ANDN U38730 ( .B(B[154]), .A(n78), .Z(n38137) );
  XNOR U38731 ( .A(n38145), .B(n38468), .Z(n38138) );
  XNOR U38732 ( .A(n38144), .B(n38142), .Z(n38468) );
  AND U38733 ( .A(n38469), .B(n38470), .Z(n38142) );
  NANDN U38734 ( .A(n38471), .B(n38472), .Z(n38470) );
  OR U38735 ( .A(n38473), .B(n38474), .Z(n38472) );
  NAND U38736 ( .A(n38474), .B(n38473), .Z(n38469) );
  ANDN U38737 ( .B(B[155]), .A(n79), .Z(n38144) );
  XNOR U38738 ( .A(n38152), .B(n38475), .Z(n38145) );
  XNOR U38739 ( .A(n38151), .B(n38149), .Z(n38475) );
  AND U38740 ( .A(n38476), .B(n38477), .Z(n38149) );
  NANDN U38741 ( .A(n38478), .B(n38479), .Z(n38477) );
  NANDN U38742 ( .A(n38480), .B(n38481), .Z(n38479) );
  NANDN U38743 ( .A(n38481), .B(n38480), .Z(n38476) );
  ANDN U38744 ( .B(B[156]), .A(n80), .Z(n38151) );
  XNOR U38745 ( .A(n38159), .B(n38482), .Z(n38152) );
  XNOR U38746 ( .A(n38158), .B(n38156), .Z(n38482) );
  AND U38747 ( .A(n38483), .B(n38484), .Z(n38156) );
  NANDN U38748 ( .A(n38485), .B(n38486), .Z(n38484) );
  OR U38749 ( .A(n38487), .B(n38488), .Z(n38486) );
  NAND U38750 ( .A(n38488), .B(n38487), .Z(n38483) );
  ANDN U38751 ( .B(B[157]), .A(n81), .Z(n38158) );
  XNOR U38752 ( .A(n38166), .B(n38489), .Z(n38159) );
  XNOR U38753 ( .A(n38165), .B(n38163), .Z(n38489) );
  AND U38754 ( .A(n38490), .B(n38491), .Z(n38163) );
  NANDN U38755 ( .A(n38492), .B(n38493), .Z(n38491) );
  NAND U38756 ( .A(n38494), .B(n38495), .Z(n38493) );
  ANDN U38757 ( .B(B[158]), .A(n82), .Z(n38165) );
  XOR U38758 ( .A(n38172), .B(n38496), .Z(n38166) );
  XNOR U38759 ( .A(n38170), .B(n38173), .Z(n38496) );
  NAND U38760 ( .A(A[2]), .B(B[159]), .Z(n38173) );
  NANDN U38761 ( .A(n38497), .B(n38498), .Z(n38170) );
  AND U38762 ( .A(A[0]), .B(B[160]), .Z(n38498) );
  XNOR U38763 ( .A(n38175), .B(n38499), .Z(n38172) );
  NAND U38764 ( .A(A[0]), .B(B[161]), .Z(n38499) );
  NAND U38765 ( .A(B[160]), .B(A[1]), .Z(n38175) );
  NAND U38766 ( .A(n38500), .B(n38501), .Z(n474) );
  NANDN U38767 ( .A(n38502), .B(n38503), .Z(n38501) );
  OR U38768 ( .A(n38504), .B(n38505), .Z(n38503) );
  NAND U38769 ( .A(n38505), .B(n38504), .Z(n38500) );
  XOR U38770 ( .A(n476), .B(n475), .Z(\A1[158] ) );
  XOR U38771 ( .A(n38505), .B(n38506), .Z(n475) );
  XNOR U38772 ( .A(n38504), .B(n38502), .Z(n38506) );
  AND U38773 ( .A(n38507), .B(n38508), .Z(n38502) );
  NANDN U38774 ( .A(n38509), .B(n38510), .Z(n38508) );
  NANDN U38775 ( .A(n38511), .B(n38512), .Z(n38510) );
  NANDN U38776 ( .A(n38512), .B(n38511), .Z(n38507) );
  ANDN U38777 ( .B(B[129]), .A(n54), .Z(n38504) );
  XNOR U38778 ( .A(n38299), .B(n38513), .Z(n38505) );
  XNOR U38779 ( .A(n38298), .B(n38296), .Z(n38513) );
  AND U38780 ( .A(n38514), .B(n38515), .Z(n38296) );
  NANDN U38781 ( .A(n38516), .B(n38517), .Z(n38515) );
  OR U38782 ( .A(n38518), .B(n38519), .Z(n38517) );
  NAND U38783 ( .A(n38519), .B(n38518), .Z(n38514) );
  ANDN U38784 ( .B(B[130]), .A(n55), .Z(n38298) );
  XNOR U38785 ( .A(n38306), .B(n38520), .Z(n38299) );
  XNOR U38786 ( .A(n38305), .B(n38303), .Z(n38520) );
  AND U38787 ( .A(n38521), .B(n38522), .Z(n38303) );
  NANDN U38788 ( .A(n38523), .B(n38524), .Z(n38522) );
  NANDN U38789 ( .A(n38525), .B(n38526), .Z(n38524) );
  NANDN U38790 ( .A(n38526), .B(n38525), .Z(n38521) );
  ANDN U38791 ( .B(B[131]), .A(n56), .Z(n38305) );
  XNOR U38792 ( .A(n38313), .B(n38527), .Z(n38306) );
  XNOR U38793 ( .A(n38312), .B(n38310), .Z(n38527) );
  AND U38794 ( .A(n38528), .B(n38529), .Z(n38310) );
  NANDN U38795 ( .A(n38530), .B(n38531), .Z(n38529) );
  OR U38796 ( .A(n38532), .B(n38533), .Z(n38531) );
  NAND U38797 ( .A(n38533), .B(n38532), .Z(n38528) );
  ANDN U38798 ( .B(B[132]), .A(n57), .Z(n38312) );
  XNOR U38799 ( .A(n38320), .B(n38534), .Z(n38313) );
  XNOR U38800 ( .A(n38319), .B(n38317), .Z(n38534) );
  AND U38801 ( .A(n38535), .B(n38536), .Z(n38317) );
  NANDN U38802 ( .A(n38537), .B(n38538), .Z(n38536) );
  NANDN U38803 ( .A(n38539), .B(n38540), .Z(n38538) );
  NANDN U38804 ( .A(n38540), .B(n38539), .Z(n38535) );
  ANDN U38805 ( .B(B[133]), .A(n58), .Z(n38319) );
  XNOR U38806 ( .A(n38327), .B(n38541), .Z(n38320) );
  XNOR U38807 ( .A(n38326), .B(n38324), .Z(n38541) );
  AND U38808 ( .A(n38542), .B(n38543), .Z(n38324) );
  NANDN U38809 ( .A(n38544), .B(n38545), .Z(n38543) );
  OR U38810 ( .A(n38546), .B(n38547), .Z(n38545) );
  NAND U38811 ( .A(n38547), .B(n38546), .Z(n38542) );
  ANDN U38812 ( .B(B[134]), .A(n59), .Z(n38326) );
  XNOR U38813 ( .A(n38334), .B(n38548), .Z(n38327) );
  XNOR U38814 ( .A(n38333), .B(n38331), .Z(n38548) );
  AND U38815 ( .A(n38549), .B(n38550), .Z(n38331) );
  NANDN U38816 ( .A(n38551), .B(n38552), .Z(n38550) );
  NANDN U38817 ( .A(n38553), .B(n38554), .Z(n38552) );
  NANDN U38818 ( .A(n38554), .B(n38553), .Z(n38549) );
  ANDN U38819 ( .B(B[135]), .A(n60), .Z(n38333) );
  XNOR U38820 ( .A(n38341), .B(n38555), .Z(n38334) );
  XNOR U38821 ( .A(n38340), .B(n38338), .Z(n38555) );
  AND U38822 ( .A(n38556), .B(n38557), .Z(n38338) );
  NANDN U38823 ( .A(n38558), .B(n38559), .Z(n38557) );
  OR U38824 ( .A(n38560), .B(n38561), .Z(n38559) );
  NAND U38825 ( .A(n38561), .B(n38560), .Z(n38556) );
  ANDN U38826 ( .B(B[136]), .A(n61), .Z(n38340) );
  XNOR U38827 ( .A(n38348), .B(n38562), .Z(n38341) );
  XNOR U38828 ( .A(n38347), .B(n38345), .Z(n38562) );
  AND U38829 ( .A(n38563), .B(n38564), .Z(n38345) );
  NANDN U38830 ( .A(n38565), .B(n38566), .Z(n38564) );
  NANDN U38831 ( .A(n38567), .B(n38568), .Z(n38566) );
  NANDN U38832 ( .A(n38568), .B(n38567), .Z(n38563) );
  ANDN U38833 ( .B(B[137]), .A(n62), .Z(n38347) );
  XNOR U38834 ( .A(n38355), .B(n38569), .Z(n38348) );
  XNOR U38835 ( .A(n38354), .B(n38352), .Z(n38569) );
  AND U38836 ( .A(n38570), .B(n38571), .Z(n38352) );
  NANDN U38837 ( .A(n38572), .B(n38573), .Z(n38571) );
  OR U38838 ( .A(n38574), .B(n38575), .Z(n38573) );
  NAND U38839 ( .A(n38575), .B(n38574), .Z(n38570) );
  ANDN U38840 ( .B(B[138]), .A(n63), .Z(n38354) );
  XNOR U38841 ( .A(n38362), .B(n38576), .Z(n38355) );
  XNOR U38842 ( .A(n38361), .B(n38359), .Z(n38576) );
  AND U38843 ( .A(n38577), .B(n38578), .Z(n38359) );
  NANDN U38844 ( .A(n38579), .B(n38580), .Z(n38578) );
  NANDN U38845 ( .A(n38581), .B(n38582), .Z(n38580) );
  NANDN U38846 ( .A(n38582), .B(n38581), .Z(n38577) );
  ANDN U38847 ( .B(B[139]), .A(n64), .Z(n38361) );
  XNOR U38848 ( .A(n38369), .B(n38583), .Z(n38362) );
  XNOR U38849 ( .A(n38368), .B(n38366), .Z(n38583) );
  AND U38850 ( .A(n38584), .B(n38585), .Z(n38366) );
  NANDN U38851 ( .A(n38586), .B(n38587), .Z(n38585) );
  OR U38852 ( .A(n38588), .B(n38589), .Z(n38587) );
  NAND U38853 ( .A(n38589), .B(n38588), .Z(n38584) );
  ANDN U38854 ( .B(B[140]), .A(n65), .Z(n38368) );
  XNOR U38855 ( .A(n38376), .B(n38590), .Z(n38369) );
  XNOR U38856 ( .A(n38375), .B(n38373), .Z(n38590) );
  AND U38857 ( .A(n38591), .B(n38592), .Z(n38373) );
  NANDN U38858 ( .A(n38593), .B(n38594), .Z(n38592) );
  NANDN U38859 ( .A(n38595), .B(n38596), .Z(n38594) );
  NANDN U38860 ( .A(n38596), .B(n38595), .Z(n38591) );
  ANDN U38861 ( .B(B[141]), .A(n66), .Z(n38375) );
  XNOR U38862 ( .A(n38383), .B(n38597), .Z(n38376) );
  XNOR U38863 ( .A(n38382), .B(n38380), .Z(n38597) );
  AND U38864 ( .A(n38598), .B(n38599), .Z(n38380) );
  NANDN U38865 ( .A(n38600), .B(n38601), .Z(n38599) );
  OR U38866 ( .A(n38602), .B(n38603), .Z(n38601) );
  NAND U38867 ( .A(n38603), .B(n38602), .Z(n38598) );
  ANDN U38868 ( .B(B[142]), .A(n67), .Z(n38382) );
  XNOR U38869 ( .A(n38390), .B(n38604), .Z(n38383) );
  XNOR U38870 ( .A(n38389), .B(n38387), .Z(n38604) );
  AND U38871 ( .A(n38605), .B(n38606), .Z(n38387) );
  NANDN U38872 ( .A(n38607), .B(n38608), .Z(n38606) );
  NANDN U38873 ( .A(n38609), .B(n38610), .Z(n38608) );
  NANDN U38874 ( .A(n38610), .B(n38609), .Z(n38605) );
  ANDN U38875 ( .B(B[143]), .A(n68), .Z(n38389) );
  XNOR U38876 ( .A(n38397), .B(n38611), .Z(n38390) );
  XNOR U38877 ( .A(n38396), .B(n38394), .Z(n38611) );
  AND U38878 ( .A(n38612), .B(n38613), .Z(n38394) );
  NANDN U38879 ( .A(n38614), .B(n38615), .Z(n38613) );
  OR U38880 ( .A(n38616), .B(n38617), .Z(n38615) );
  NAND U38881 ( .A(n38617), .B(n38616), .Z(n38612) );
  ANDN U38882 ( .B(B[144]), .A(n69), .Z(n38396) );
  XNOR U38883 ( .A(n38404), .B(n38618), .Z(n38397) );
  XNOR U38884 ( .A(n38403), .B(n38401), .Z(n38618) );
  AND U38885 ( .A(n38619), .B(n38620), .Z(n38401) );
  NANDN U38886 ( .A(n38621), .B(n38622), .Z(n38620) );
  NANDN U38887 ( .A(n38623), .B(n38624), .Z(n38622) );
  NANDN U38888 ( .A(n38624), .B(n38623), .Z(n38619) );
  ANDN U38889 ( .B(B[145]), .A(n70), .Z(n38403) );
  XNOR U38890 ( .A(n38411), .B(n38625), .Z(n38404) );
  XNOR U38891 ( .A(n38410), .B(n38408), .Z(n38625) );
  AND U38892 ( .A(n38626), .B(n38627), .Z(n38408) );
  NANDN U38893 ( .A(n38628), .B(n38629), .Z(n38627) );
  OR U38894 ( .A(n38630), .B(n38631), .Z(n38629) );
  NAND U38895 ( .A(n38631), .B(n38630), .Z(n38626) );
  ANDN U38896 ( .B(B[146]), .A(n71), .Z(n38410) );
  XNOR U38897 ( .A(n38418), .B(n38632), .Z(n38411) );
  XNOR U38898 ( .A(n38417), .B(n38415), .Z(n38632) );
  AND U38899 ( .A(n38633), .B(n38634), .Z(n38415) );
  NANDN U38900 ( .A(n38635), .B(n38636), .Z(n38634) );
  NANDN U38901 ( .A(n38637), .B(n38638), .Z(n38636) );
  NANDN U38902 ( .A(n38638), .B(n38637), .Z(n38633) );
  ANDN U38903 ( .B(B[147]), .A(n72), .Z(n38417) );
  XNOR U38904 ( .A(n38425), .B(n38639), .Z(n38418) );
  XNOR U38905 ( .A(n38424), .B(n38422), .Z(n38639) );
  AND U38906 ( .A(n38640), .B(n38641), .Z(n38422) );
  NANDN U38907 ( .A(n38642), .B(n38643), .Z(n38641) );
  OR U38908 ( .A(n38644), .B(n38645), .Z(n38643) );
  NAND U38909 ( .A(n38645), .B(n38644), .Z(n38640) );
  ANDN U38910 ( .B(B[148]), .A(n73), .Z(n38424) );
  XNOR U38911 ( .A(n38432), .B(n38646), .Z(n38425) );
  XNOR U38912 ( .A(n38431), .B(n38429), .Z(n38646) );
  AND U38913 ( .A(n38647), .B(n38648), .Z(n38429) );
  NANDN U38914 ( .A(n38649), .B(n38650), .Z(n38648) );
  NANDN U38915 ( .A(n38651), .B(n38652), .Z(n38650) );
  NANDN U38916 ( .A(n38652), .B(n38651), .Z(n38647) );
  ANDN U38917 ( .B(B[149]), .A(n74), .Z(n38431) );
  XNOR U38918 ( .A(n38439), .B(n38653), .Z(n38432) );
  XNOR U38919 ( .A(n38438), .B(n38436), .Z(n38653) );
  AND U38920 ( .A(n38654), .B(n38655), .Z(n38436) );
  NANDN U38921 ( .A(n38656), .B(n38657), .Z(n38655) );
  OR U38922 ( .A(n38658), .B(n38659), .Z(n38657) );
  NAND U38923 ( .A(n38659), .B(n38658), .Z(n38654) );
  ANDN U38924 ( .B(B[150]), .A(n75), .Z(n38438) );
  XNOR U38925 ( .A(n38446), .B(n38660), .Z(n38439) );
  XNOR U38926 ( .A(n38445), .B(n38443), .Z(n38660) );
  AND U38927 ( .A(n38661), .B(n38662), .Z(n38443) );
  NANDN U38928 ( .A(n38663), .B(n38664), .Z(n38662) );
  NANDN U38929 ( .A(n38665), .B(n38666), .Z(n38664) );
  NANDN U38930 ( .A(n38666), .B(n38665), .Z(n38661) );
  ANDN U38931 ( .B(B[151]), .A(n76), .Z(n38445) );
  XNOR U38932 ( .A(n38453), .B(n38667), .Z(n38446) );
  XNOR U38933 ( .A(n38452), .B(n38450), .Z(n38667) );
  AND U38934 ( .A(n38668), .B(n38669), .Z(n38450) );
  NANDN U38935 ( .A(n38670), .B(n38671), .Z(n38669) );
  OR U38936 ( .A(n38672), .B(n38673), .Z(n38671) );
  NAND U38937 ( .A(n38673), .B(n38672), .Z(n38668) );
  ANDN U38938 ( .B(B[152]), .A(n77), .Z(n38452) );
  XNOR U38939 ( .A(n38460), .B(n38674), .Z(n38453) );
  XNOR U38940 ( .A(n38459), .B(n38457), .Z(n38674) );
  AND U38941 ( .A(n38675), .B(n38676), .Z(n38457) );
  NANDN U38942 ( .A(n38677), .B(n38678), .Z(n38676) );
  NANDN U38943 ( .A(n38679), .B(n38680), .Z(n38678) );
  NANDN U38944 ( .A(n38680), .B(n38679), .Z(n38675) );
  ANDN U38945 ( .B(B[153]), .A(n78), .Z(n38459) );
  XNOR U38946 ( .A(n38467), .B(n38681), .Z(n38460) );
  XNOR U38947 ( .A(n38466), .B(n38464), .Z(n38681) );
  AND U38948 ( .A(n38682), .B(n38683), .Z(n38464) );
  NANDN U38949 ( .A(n38684), .B(n38685), .Z(n38683) );
  OR U38950 ( .A(n38686), .B(n38687), .Z(n38685) );
  NAND U38951 ( .A(n38687), .B(n38686), .Z(n38682) );
  ANDN U38952 ( .B(B[154]), .A(n79), .Z(n38466) );
  XNOR U38953 ( .A(n38474), .B(n38688), .Z(n38467) );
  XNOR U38954 ( .A(n38473), .B(n38471), .Z(n38688) );
  AND U38955 ( .A(n38689), .B(n38690), .Z(n38471) );
  NANDN U38956 ( .A(n38691), .B(n38692), .Z(n38690) );
  NANDN U38957 ( .A(n38693), .B(n38694), .Z(n38692) );
  NANDN U38958 ( .A(n38694), .B(n38693), .Z(n38689) );
  ANDN U38959 ( .B(B[155]), .A(n80), .Z(n38473) );
  XNOR U38960 ( .A(n38481), .B(n38695), .Z(n38474) );
  XNOR U38961 ( .A(n38480), .B(n38478), .Z(n38695) );
  AND U38962 ( .A(n38696), .B(n38697), .Z(n38478) );
  NANDN U38963 ( .A(n38698), .B(n38699), .Z(n38697) );
  OR U38964 ( .A(n38700), .B(n38701), .Z(n38699) );
  NAND U38965 ( .A(n38701), .B(n38700), .Z(n38696) );
  ANDN U38966 ( .B(B[156]), .A(n81), .Z(n38480) );
  XNOR U38967 ( .A(n38488), .B(n38702), .Z(n38481) );
  XNOR U38968 ( .A(n38487), .B(n38485), .Z(n38702) );
  AND U38969 ( .A(n38703), .B(n38704), .Z(n38485) );
  NANDN U38970 ( .A(n38705), .B(n38706), .Z(n38704) );
  NAND U38971 ( .A(n38707), .B(n38708), .Z(n38706) );
  ANDN U38972 ( .B(B[157]), .A(n82), .Z(n38487) );
  XOR U38973 ( .A(n38494), .B(n38709), .Z(n38488) );
  XNOR U38974 ( .A(n38492), .B(n38495), .Z(n38709) );
  NAND U38975 ( .A(A[2]), .B(B[158]), .Z(n38495) );
  NANDN U38976 ( .A(n38710), .B(n38711), .Z(n38492) );
  AND U38977 ( .A(A[0]), .B(B[159]), .Z(n38711) );
  XNOR U38978 ( .A(n38497), .B(n38712), .Z(n38494) );
  NAND U38979 ( .A(A[0]), .B(B[160]), .Z(n38712) );
  NAND U38980 ( .A(B[159]), .B(A[1]), .Z(n38497) );
  NAND U38981 ( .A(n38713), .B(n38714), .Z(n476) );
  NANDN U38982 ( .A(n38715), .B(n38716), .Z(n38714) );
  OR U38983 ( .A(n38717), .B(n38718), .Z(n38716) );
  NAND U38984 ( .A(n38718), .B(n38717), .Z(n38713) );
  XOR U38985 ( .A(n478), .B(n477), .Z(\A1[157] ) );
  XOR U38986 ( .A(n38718), .B(n38719), .Z(n477) );
  XNOR U38987 ( .A(n38717), .B(n38715), .Z(n38719) );
  AND U38988 ( .A(n38720), .B(n38721), .Z(n38715) );
  NANDN U38989 ( .A(n38722), .B(n38723), .Z(n38721) );
  NANDN U38990 ( .A(n38724), .B(n38725), .Z(n38723) );
  NANDN U38991 ( .A(n38725), .B(n38724), .Z(n38720) );
  ANDN U38992 ( .B(B[128]), .A(n54), .Z(n38717) );
  XNOR U38993 ( .A(n38512), .B(n38726), .Z(n38718) );
  XNOR U38994 ( .A(n38511), .B(n38509), .Z(n38726) );
  AND U38995 ( .A(n38727), .B(n38728), .Z(n38509) );
  NANDN U38996 ( .A(n38729), .B(n38730), .Z(n38728) );
  OR U38997 ( .A(n38731), .B(n38732), .Z(n38730) );
  NAND U38998 ( .A(n38732), .B(n38731), .Z(n38727) );
  ANDN U38999 ( .B(B[129]), .A(n55), .Z(n38511) );
  XNOR U39000 ( .A(n38519), .B(n38733), .Z(n38512) );
  XNOR U39001 ( .A(n38518), .B(n38516), .Z(n38733) );
  AND U39002 ( .A(n38734), .B(n38735), .Z(n38516) );
  NANDN U39003 ( .A(n38736), .B(n38737), .Z(n38735) );
  NANDN U39004 ( .A(n38738), .B(n38739), .Z(n38737) );
  NANDN U39005 ( .A(n38739), .B(n38738), .Z(n38734) );
  ANDN U39006 ( .B(B[130]), .A(n56), .Z(n38518) );
  XNOR U39007 ( .A(n38526), .B(n38740), .Z(n38519) );
  XNOR U39008 ( .A(n38525), .B(n38523), .Z(n38740) );
  AND U39009 ( .A(n38741), .B(n38742), .Z(n38523) );
  NANDN U39010 ( .A(n38743), .B(n38744), .Z(n38742) );
  OR U39011 ( .A(n38745), .B(n38746), .Z(n38744) );
  NAND U39012 ( .A(n38746), .B(n38745), .Z(n38741) );
  ANDN U39013 ( .B(B[131]), .A(n57), .Z(n38525) );
  XNOR U39014 ( .A(n38533), .B(n38747), .Z(n38526) );
  XNOR U39015 ( .A(n38532), .B(n38530), .Z(n38747) );
  AND U39016 ( .A(n38748), .B(n38749), .Z(n38530) );
  NANDN U39017 ( .A(n38750), .B(n38751), .Z(n38749) );
  NANDN U39018 ( .A(n38752), .B(n38753), .Z(n38751) );
  NANDN U39019 ( .A(n38753), .B(n38752), .Z(n38748) );
  ANDN U39020 ( .B(B[132]), .A(n58), .Z(n38532) );
  XNOR U39021 ( .A(n38540), .B(n38754), .Z(n38533) );
  XNOR U39022 ( .A(n38539), .B(n38537), .Z(n38754) );
  AND U39023 ( .A(n38755), .B(n38756), .Z(n38537) );
  NANDN U39024 ( .A(n38757), .B(n38758), .Z(n38756) );
  OR U39025 ( .A(n38759), .B(n38760), .Z(n38758) );
  NAND U39026 ( .A(n38760), .B(n38759), .Z(n38755) );
  ANDN U39027 ( .B(B[133]), .A(n59), .Z(n38539) );
  XNOR U39028 ( .A(n38547), .B(n38761), .Z(n38540) );
  XNOR U39029 ( .A(n38546), .B(n38544), .Z(n38761) );
  AND U39030 ( .A(n38762), .B(n38763), .Z(n38544) );
  NANDN U39031 ( .A(n38764), .B(n38765), .Z(n38763) );
  NANDN U39032 ( .A(n38766), .B(n38767), .Z(n38765) );
  NANDN U39033 ( .A(n38767), .B(n38766), .Z(n38762) );
  ANDN U39034 ( .B(B[134]), .A(n60), .Z(n38546) );
  XNOR U39035 ( .A(n38554), .B(n38768), .Z(n38547) );
  XNOR U39036 ( .A(n38553), .B(n38551), .Z(n38768) );
  AND U39037 ( .A(n38769), .B(n38770), .Z(n38551) );
  NANDN U39038 ( .A(n38771), .B(n38772), .Z(n38770) );
  OR U39039 ( .A(n38773), .B(n38774), .Z(n38772) );
  NAND U39040 ( .A(n38774), .B(n38773), .Z(n38769) );
  ANDN U39041 ( .B(B[135]), .A(n61), .Z(n38553) );
  XNOR U39042 ( .A(n38561), .B(n38775), .Z(n38554) );
  XNOR U39043 ( .A(n38560), .B(n38558), .Z(n38775) );
  AND U39044 ( .A(n38776), .B(n38777), .Z(n38558) );
  NANDN U39045 ( .A(n38778), .B(n38779), .Z(n38777) );
  NANDN U39046 ( .A(n38780), .B(n38781), .Z(n38779) );
  NANDN U39047 ( .A(n38781), .B(n38780), .Z(n38776) );
  ANDN U39048 ( .B(B[136]), .A(n62), .Z(n38560) );
  XNOR U39049 ( .A(n38568), .B(n38782), .Z(n38561) );
  XNOR U39050 ( .A(n38567), .B(n38565), .Z(n38782) );
  AND U39051 ( .A(n38783), .B(n38784), .Z(n38565) );
  NANDN U39052 ( .A(n38785), .B(n38786), .Z(n38784) );
  OR U39053 ( .A(n38787), .B(n38788), .Z(n38786) );
  NAND U39054 ( .A(n38788), .B(n38787), .Z(n38783) );
  ANDN U39055 ( .B(B[137]), .A(n63), .Z(n38567) );
  XNOR U39056 ( .A(n38575), .B(n38789), .Z(n38568) );
  XNOR U39057 ( .A(n38574), .B(n38572), .Z(n38789) );
  AND U39058 ( .A(n38790), .B(n38791), .Z(n38572) );
  NANDN U39059 ( .A(n38792), .B(n38793), .Z(n38791) );
  NANDN U39060 ( .A(n38794), .B(n38795), .Z(n38793) );
  NANDN U39061 ( .A(n38795), .B(n38794), .Z(n38790) );
  ANDN U39062 ( .B(B[138]), .A(n64), .Z(n38574) );
  XNOR U39063 ( .A(n38582), .B(n38796), .Z(n38575) );
  XNOR U39064 ( .A(n38581), .B(n38579), .Z(n38796) );
  AND U39065 ( .A(n38797), .B(n38798), .Z(n38579) );
  NANDN U39066 ( .A(n38799), .B(n38800), .Z(n38798) );
  OR U39067 ( .A(n38801), .B(n38802), .Z(n38800) );
  NAND U39068 ( .A(n38802), .B(n38801), .Z(n38797) );
  ANDN U39069 ( .B(B[139]), .A(n65), .Z(n38581) );
  XNOR U39070 ( .A(n38589), .B(n38803), .Z(n38582) );
  XNOR U39071 ( .A(n38588), .B(n38586), .Z(n38803) );
  AND U39072 ( .A(n38804), .B(n38805), .Z(n38586) );
  NANDN U39073 ( .A(n38806), .B(n38807), .Z(n38805) );
  NANDN U39074 ( .A(n38808), .B(n38809), .Z(n38807) );
  NANDN U39075 ( .A(n38809), .B(n38808), .Z(n38804) );
  ANDN U39076 ( .B(B[140]), .A(n66), .Z(n38588) );
  XNOR U39077 ( .A(n38596), .B(n38810), .Z(n38589) );
  XNOR U39078 ( .A(n38595), .B(n38593), .Z(n38810) );
  AND U39079 ( .A(n38811), .B(n38812), .Z(n38593) );
  NANDN U39080 ( .A(n38813), .B(n38814), .Z(n38812) );
  OR U39081 ( .A(n38815), .B(n38816), .Z(n38814) );
  NAND U39082 ( .A(n38816), .B(n38815), .Z(n38811) );
  ANDN U39083 ( .B(B[141]), .A(n67), .Z(n38595) );
  XNOR U39084 ( .A(n38603), .B(n38817), .Z(n38596) );
  XNOR U39085 ( .A(n38602), .B(n38600), .Z(n38817) );
  AND U39086 ( .A(n38818), .B(n38819), .Z(n38600) );
  NANDN U39087 ( .A(n38820), .B(n38821), .Z(n38819) );
  NANDN U39088 ( .A(n38822), .B(n38823), .Z(n38821) );
  NANDN U39089 ( .A(n38823), .B(n38822), .Z(n38818) );
  ANDN U39090 ( .B(B[142]), .A(n68), .Z(n38602) );
  XNOR U39091 ( .A(n38610), .B(n38824), .Z(n38603) );
  XNOR U39092 ( .A(n38609), .B(n38607), .Z(n38824) );
  AND U39093 ( .A(n38825), .B(n38826), .Z(n38607) );
  NANDN U39094 ( .A(n38827), .B(n38828), .Z(n38826) );
  OR U39095 ( .A(n38829), .B(n38830), .Z(n38828) );
  NAND U39096 ( .A(n38830), .B(n38829), .Z(n38825) );
  ANDN U39097 ( .B(B[143]), .A(n69), .Z(n38609) );
  XNOR U39098 ( .A(n38617), .B(n38831), .Z(n38610) );
  XNOR U39099 ( .A(n38616), .B(n38614), .Z(n38831) );
  AND U39100 ( .A(n38832), .B(n38833), .Z(n38614) );
  NANDN U39101 ( .A(n38834), .B(n38835), .Z(n38833) );
  NANDN U39102 ( .A(n38836), .B(n38837), .Z(n38835) );
  NANDN U39103 ( .A(n38837), .B(n38836), .Z(n38832) );
  ANDN U39104 ( .B(B[144]), .A(n70), .Z(n38616) );
  XNOR U39105 ( .A(n38624), .B(n38838), .Z(n38617) );
  XNOR U39106 ( .A(n38623), .B(n38621), .Z(n38838) );
  AND U39107 ( .A(n38839), .B(n38840), .Z(n38621) );
  NANDN U39108 ( .A(n38841), .B(n38842), .Z(n38840) );
  OR U39109 ( .A(n38843), .B(n38844), .Z(n38842) );
  NAND U39110 ( .A(n38844), .B(n38843), .Z(n38839) );
  ANDN U39111 ( .B(B[145]), .A(n71), .Z(n38623) );
  XNOR U39112 ( .A(n38631), .B(n38845), .Z(n38624) );
  XNOR U39113 ( .A(n38630), .B(n38628), .Z(n38845) );
  AND U39114 ( .A(n38846), .B(n38847), .Z(n38628) );
  NANDN U39115 ( .A(n38848), .B(n38849), .Z(n38847) );
  NANDN U39116 ( .A(n38850), .B(n38851), .Z(n38849) );
  NANDN U39117 ( .A(n38851), .B(n38850), .Z(n38846) );
  ANDN U39118 ( .B(B[146]), .A(n72), .Z(n38630) );
  XNOR U39119 ( .A(n38638), .B(n38852), .Z(n38631) );
  XNOR U39120 ( .A(n38637), .B(n38635), .Z(n38852) );
  AND U39121 ( .A(n38853), .B(n38854), .Z(n38635) );
  NANDN U39122 ( .A(n38855), .B(n38856), .Z(n38854) );
  OR U39123 ( .A(n38857), .B(n38858), .Z(n38856) );
  NAND U39124 ( .A(n38858), .B(n38857), .Z(n38853) );
  ANDN U39125 ( .B(B[147]), .A(n73), .Z(n38637) );
  XNOR U39126 ( .A(n38645), .B(n38859), .Z(n38638) );
  XNOR U39127 ( .A(n38644), .B(n38642), .Z(n38859) );
  AND U39128 ( .A(n38860), .B(n38861), .Z(n38642) );
  NANDN U39129 ( .A(n38862), .B(n38863), .Z(n38861) );
  NANDN U39130 ( .A(n38864), .B(n38865), .Z(n38863) );
  NANDN U39131 ( .A(n38865), .B(n38864), .Z(n38860) );
  ANDN U39132 ( .B(B[148]), .A(n74), .Z(n38644) );
  XNOR U39133 ( .A(n38652), .B(n38866), .Z(n38645) );
  XNOR U39134 ( .A(n38651), .B(n38649), .Z(n38866) );
  AND U39135 ( .A(n38867), .B(n38868), .Z(n38649) );
  NANDN U39136 ( .A(n38869), .B(n38870), .Z(n38868) );
  OR U39137 ( .A(n38871), .B(n38872), .Z(n38870) );
  NAND U39138 ( .A(n38872), .B(n38871), .Z(n38867) );
  ANDN U39139 ( .B(B[149]), .A(n75), .Z(n38651) );
  XNOR U39140 ( .A(n38659), .B(n38873), .Z(n38652) );
  XNOR U39141 ( .A(n38658), .B(n38656), .Z(n38873) );
  AND U39142 ( .A(n38874), .B(n38875), .Z(n38656) );
  NANDN U39143 ( .A(n38876), .B(n38877), .Z(n38875) );
  NANDN U39144 ( .A(n38878), .B(n38879), .Z(n38877) );
  NANDN U39145 ( .A(n38879), .B(n38878), .Z(n38874) );
  ANDN U39146 ( .B(B[150]), .A(n76), .Z(n38658) );
  XNOR U39147 ( .A(n38666), .B(n38880), .Z(n38659) );
  XNOR U39148 ( .A(n38665), .B(n38663), .Z(n38880) );
  AND U39149 ( .A(n38881), .B(n38882), .Z(n38663) );
  NANDN U39150 ( .A(n38883), .B(n38884), .Z(n38882) );
  OR U39151 ( .A(n38885), .B(n38886), .Z(n38884) );
  NAND U39152 ( .A(n38886), .B(n38885), .Z(n38881) );
  ANDN U39153 ( .B(B[151]), .A(n77), .Z(n38665) );
  XNOR U39154 ( .A(n38673), .B(n38887), .Z(n38666) );
  XNOR U39155 ( .A(n38672), .B(n38670), .Z(n38887) );
  AND U39156 ( .A(n38888), .B(n38889), .Z(n38670) );
  NANDN U39157 ( .A(n38890), .B(n38891), .Z(n38889) );
  NANDN U39158 ( .A(n38892), .B(n38893), .Z(n38891) );
  NANDN U39159 ( .A(n38893), .B(n38892), .Z(n38888) );
  ANDN U39160 ( .B(B[152]), .A(n78), .Z(n38672) );
  XNOR U39161 ( .A(n38680), .B(n38894), .Z(n38673) );
  XNOR U39162 ( .A(n38679), .B(n38677), .Z(n38894) );
  AND U39163 ( .A(n38895), .B(n38896), .Z(n38677) );
  NANDN U39164 ( .A(n38897), .B(n38898), .Z(n38896) );
  OR U39165 ( .A(n38899), .B(n38900), .Z(n38898) );
  NAND U39166 ( .A(n38900), .B(n38899), .Z(n38895) );
  ANDN U39167 ( .B(B[153]), .A(n79), .Z(n38679) );
  XNOR U39168 ( .A(n38687), .B(n38901), .Z(n38680) );
  XNOR U39169 ( .A(n38686), .B(n38684), .Z(n38901) );
  AND U39170 ( .A(n38902), .B(n38903), .Z(n38684) );
  NANDN U39171 ( .A(n38904), .B(n38905), .Z(n38903) );
  NANDN U39172 ( .A(n38906), .B(n38907), .Z(n38905) );
  NANDN U39173 ( .A(n38907), .B(n38906), .Z(n38902) );
  ANDN U39174 ( .B(B[154]), .A(n80), .Z(n38686) );
  XNOR U39175 ( .A(n38694), .B(n38908), .Z(n38687) );
  XNOR U39176 ( .A(n38693), .B(n38691), .Z(n38908) );
  AND U39177 ( .A(n38909), .B(n38910), .Z(n38691) );
  NANDN U39178 ( .A(n38911), .B(n38912), .Z(n38910) );
  OR U39179 ( .A(n38913), .B(n38914), .Z(n38912) );
  NAND U39180 ( .A(n38914), .B(n38913), .Z(n38909) );
  ANDN U39181 ( .B(B[155]), .A(n81), .Z(n38693) );
  XNOR U39182 ( .A(n38701), .B(n38915), .Z(n38694) );
  XNOR U39183 ( .A(n38700), .B(n38698), .Z(n38915) );
  AND U39184 ( .A(n38916), .B(n38917), .Z(n38698) );
  NANDN U39185 ( .A(n38918), .B(n38919), .Z(n38917) );
  NAND U39186 ( .A(n38920), .B(n38921), .Z(n38919) );
  ANDN U39187 ( .B(B[156]), .A(n82), .Z(n38700) );
  XOR U39188 ( .A(n38707), .B(n38922), .Z(n38701) );
  XNOR U39189 ( .A(n38705), .B(n38708), .Z(n38922) );
  NAND U39190 ( .A(A[2]), .B(B[157]), .Z(n38708) );
  NANDN U39191 ( .A(n38923), .B(n38924), .Z(n38705) );
  AND U39192 ( .A(A[0]), .B(B[158]), .Z(n38924) );
  XNOR U39193 ( .A(n38710), .B(n38925), .Z(n38707) );
  NAND U39194 ( .A(A[0]), .B(B[159]), .Z(n38925) );
  NAND U39195 ( .A(B[158]), .B(A[1]), .Z(n38710) );
  NAND U39196 ( .A(n38926), .B(n38927), .Z(n478) );
  NANDN U39197 ( .A(n38928), .B(n38929), .Z(n38927) );
  OR U39198 ( .A(n38930), .B(n38931), .Z(n38929) );
  NAND U39199 ( .A(n38931), .B(n38930), .Z(n38926) );
  XOR U39200 ( .A(n480), .B(n479), .Z(\A1[156] ) );
  XOR U39201 ( .A(n38931), .B(n38932), .Z(n479) );
  XNOR U39202 ( .A(n38930), .B(n38928), .Z(n38932) );
  AND U39203 ( .A(n38933), .B(n38934), .Z(n38928) );
  NANDN U39204 ( .A(n38935), .B(n38936), .Z(n38934) );
  NANDN U39205 ( .A(n38937), .B(n38938), .Z(n38936) );
  NANDN U39206 ( .A(n38938), .B(n38937), .Z(n38933) );
  ANDN U39207 ( .B(B[127]), .A(n54), .Z(n38930) );
  XNOR U39208 ( .A(n38725), .B(n38939), .Z(n38931) );
  XNOR U39209 ( .A(n38724), .B(n38722), .Z(n38939) );
  AND U39210 ( .A(n38940), .B(n38941), .Z(n38722) );
  NANDN U39211 ( .A(n38942), .B(n38943), .Z(n38941) );
  OR U39212 ( .A(n38944), .B(n38945), .Z(n38943) );
  NAND U39213 ( .A(n38945), .B(n38944), .Z(n38940) );
  ANDN U39214 ( .B(B[128]), .A(n55), .Z(n38724) );
  XNOR U39215 ( .A(n38732), .B(n38946), .Z(n38725) );
  XNOR U39216 ( .A(n38731), .B(n38729), .Z(n38946) );
  AND U39217 ( .A(n38947), .B(n38948), .Z(n38729) );
  NANDN U39218 ( .A(n38949), .B(n38950), .Z(n38948) );
  NANDN U39219 ( .A(n38951), .B(n38952), .Z(n38950) );
  NANDN U39220 ( .A(n38952), .B(n38951), .Z(n38947) );
  ANDN U39221 ( .B(B[129]), .A(n56), .Z(n38731) );
  XNOR U39222 ( .A(n38739), .B(n38953), .Z(n38732) );
  XNOR U39223 ( .A(n38738), .B(n38736), .Z(n38953) );
  AND U39224 ( .A(n38954), .B(n38955), .Z(n38736) );
  NANDN U39225 ( .A(n38956), .B(n38957), .Z(n38955) );
  OR U39226 ( .A(n38958), .B(n38959), .Z(n38957) );
  NAND U39227 ( .A(n38959), .B(n38958), .Z(n38954) );
  ANDN U39228 ( .B(B[130]), .A(n57), .Z(n38738) );
  XNOR U39229 ( .A(n38746), .B(n38960), .Z(n38739) );
  XNOR U39230 ( .A(n38745), .B(n38743), .Z(n38960) );
  AND U39231 ( .A(n38961), .B(n38962), .Z(n38743) );
  NANDN U39232 ( .A(n38963), .B(n38964), .Z(n38962) );
  NANDN U39233 ( .A(n38965), .B(n38966), .Z(n38964) );
  NANDN U39234 ( .A(n38966), .B(n38965), .Z(n38961) );
  ANDN U39235 ( .B(B[131]), .A(n58), .Z(n38745) );
  XNOR U39236 ( .A(n38753), .B(n38967), .Z(n38746) );
  XNOR U39237 ( .A(n38752), .B(n38750), .Z(n38967) );
  AND U39238 ( .A(n38968), .B(n38969), .Z(n38750) );
  NANDN U39239 ( .A(n38970), .B(n38971), .Z(n38969) );
  OR U39240 ( .A(n38972), .B(n38973), .Z(n38971) );
  NAND U39241 ( .A(n38973), .B(n38972), .Z(n38968) );
  ANDN U39242 ( .B(B[132]), .A(n59), .Z(n38752) );
  XNOR U39243 ( .A(n38760), .B(n38974), .Z(n38753) );
  XNOR U39244 ( .A(n38759), .B(n38757), .Z(n38974) );
  AND U39245 ( .A(n38975), .B(n38976), .Z(n38757) );
  NANDN U39246 ( .A(n38977), .B(n38978), .Z(n38976) );
  NANDN U39247 ( .A(n38979), .B(n38980), .Z(n38978) );
  NANDN U39248 ( .A(n38980), .B(n38979), .Z(n38975) );
  ANDN U39249 ( .B(B[133]), .A(n60), .Z(n38759) );
  XNOR U39250 ( .A(n38767), .B(n38981), .Z(n38760) );
  XNOR U39251 ( .A(n38766), .B(n38764), .Z(n38981) );
  AND U39252 ( .A(n38982), .B(n38983), .Z(n38764) );
  NANDN U39253 ( .A(n38984), .B(n38985), .Z(n38983) );
  OR U39254 ( .A(n38986), .B(n38987), .Z(n38985) );
  NAND U39255 ( .A(n38987), .B(n38986), .Z(n38982) );
  ANDN U39256 ( .B(B[134]), .A(n61), .Z(n38766) );
  XNOR U39257 ( .A(n38774), .B(n38988), .Z(n38767) );
  XNOR U39258 ( .A(n38773), .B(n38771), .Z(n38988) );
  AND U39259 ( .A(n38989), .B(n38990), .Z(n38771) );
  NANDN U39260 ( .A(n38991), .B(n38992), .Z(n38990) );
  NANDN U39261 ( .A(n38993), .B(n38994), .Z(n38992) );
  NANDN U39262 ( .A(n38994), .B(n38993), .Z(n38989) );
  ANDN U39263 ( .B(B[135]), .A(n62), .Z(n38773) );
  XNOR U39264 ( .A(n38781), .B(n38995), .Z(n38774) );
  XNOR U39265 ( .A(n38780), .B(n38778), .Z(n38995) );
  AND U39266 ( .A(n38996), .B(n38997), .Z(n38778) );
  NANDN U39267 ( .A(n38998), .B(n38999), .Z(n38997) );
  OR U39268 ( .A(n39000), .B(n39001), .Z(n38999) );
  NAND U39269 ( .A(n39001), .B(n39000), .Z(n38996) );
  ANDN U39270 ( .B(B[136]), .A(n63), .Z(n38780) );
  XNOR U39271 ( .A(n38788), .B(n39002), .Z(n38781) );
  XNOR U39272 ( .A(n38787), .B(n38785), .Z(n39002) );
  AND U39273 ( .A(n39003), .B(n39004), .Z(n38785) );
  NANDN U39274 ( .A(n39005), .B(n39006), .Z(n39004) );
  NANDN U39275 ( .A(n39007), .B(n39008), .Z(n39006) );
  NANDN U39276 ( .A(n39008), .B(n39007), .Z(n39003) );
  ANDN U39277 ( .B(B[137]), .A(n64), .Z(n38787) );
  XNOR U39278 ( .A(n38795), .B(n39009), .Z(n38788) );
  XNOR U39279 ( .A(n38794), .B(n38792), .Z(n39009) );
  AND U39280 ( .A(n39010), .B(n39011), .Z(n38792) );
  NANDN U39281 ( .A(n39012), .B(n39013), .Z(n39011) );
  OR U39282 ( .A(n39014), .B(n39015), .Z(n39013) );
  NAND U39283 ( .A(n39015), .B(n39014), .Z(n39010) );
  ANDN U39284 ( .B(B[138]), .A(n65), .Z(n38794) );
  XNOR U39285 ( .A(n38802), .B(n39016), .Z(n38795) );
  XNOR U39286 ( .A(n38801), .B(n38799), .Z(n39016) );
  AND U39287 ( .A(n39017), .B(n39018), .Z(n38799) );
  NANDN U39288 ( .A(n39019), .B(n39020), .Z(n39018) );
  NANDN U39289 ( .A(n39021), .B(n39022), .Z(n39020) );
  NANDN U39290 ( .A(n39022), .B(n39021), .Z(n39017) );
  ANDN U39291 ( .B(B[139]), .A(n66), .Z(n38801) );
  XNOR U39292 ( .A(n38809), .B(n39023), .Z(n38802) );
  XNOR U39293 ( .A(n38808), .B(n38806), .Z(n39023) );
  AND U39294 ( .A(n39024), .B(n39025), .Z(n38806) );
  NANDN U39295 ( .A(n39026), .B(n39027), .Z(n39025) );
  OR U39296 ( .A(n39028), .B(n39029), .Z(n39027) );
  NAND U39297 ( .A(n39029), .B(n39028), .Z(n39024) );
  ANDN U39298 ( .B(B[140]), .A(n67), .Z(n38808) );
  XNOR U39299 ( .A(n38816), .B(n39030), .Z(n38809) );
  XNOR U39300 ( .A(n38815), .B(n38813), .Z(n39030) );
  AND U39301 ( .A(n39031), .B(n39032), .Z(n38813) );
  NANDN U39302 ( .A(n39033), .B(n39034), .Z(n39032) );
  NANDN U39303 ( .A(n39035), .B(n39036), .Z(n39034) );
  NANDN U39304 ( .A(n39036), .B(n39035), .Z(n39031) );
  ANDN U39305 ( .B(B[141]), .A(n68), .Z(n38815) );
  XNOR U39306 ( .A(n38823), .B(n39037), .Z(n38816) );
  XNOR U39307 ( .A(n38822), .B(n38820), .Z(n39037) );
  AND U39308 ( .A(n39038), .B(n39039), .Z(n38820) );
  NANDN U39309 ( .A(n39040), .B(n39041), .Z(n39039) );
  OR U39310 ( .A(n39042), .B(n39043), .Z(n39041) );
  NAND U39311 ( .A(n39043), .B(n39042), .Z(n39038) );
  ANDN U39312 ( .B(B[142]), .A(n69), .Z(n38822) );
  XNOR U39313 ( .A(n38830), .B(n39044), .Z(n38823) );
  XNOR U39314 ( .A(n38829), .B(n38827), .Z(n39044) );
  AND U39315 ( .A(n39045), .B(n39046), .Z(n38827) );
  NANDN U39316 ( .A(n39047), .B(n39048), .Z(n39046) );
  NANDN U39317 ( .A(n39049), .B(n39050), .Z(n39048) );
  NANDN U39318 ( .A(n39050), .B(n39049), .Z(n39045) );
  ANDN U39319 ( .B(B[143]), .A(n70), .Z(n38829) );
  XNOR U39320 ( .A(n38837), .B(n39051), .Z(n38830) );
  XNOR U39321 ( .A(n38836), .B(n38834), .Z(n39051) );
  AND U39322 ( .A(n39052), .B(n39053), .Z(n38834) );
  NANDN U39323 ( .A(n39054), .B(n39055), .Z(n39053) );
  OR U39324 ( .A(n39056), .B(n39057), .Z(n39055) );
  NAND U39325 ( .A(n39057), .B(n39056), .Z(n39052) );
  ANDN U39326 ( .B(B[144]), .A(n71), .Z(n38836) );
  XNOR U39327 ( .A(n38844), .B(n39058), .Z(n38837) );
  XNOR U39328 ( .A(n38843), .B(n38841), .Z(n39058) );
  AND U39329 ( .A(n39059), .B(n39060), .Z(n38841) );
  NANDN U39330 ( .A(n39061), .B(n39062), .Z(n39060) );
  NANDN U39331 ( .A(n39063), .B(n39064), .Z(n39062) );
  NANDN U39332 ( .A(n39064), .B(n39063), .Z(n39059) );
  ANDN U39333 ( .B(B[145]), .A(n72), .Z(n38843) );
  XNOR U39334 ( .A(n38851), .B(n39065), .Z(n38844) );
  XNOR U39335 ( .A(n38850), .B(n38848), .Z(n39065) );
  AND U39336 ( .A(n39066), .B(n39067), .Z(n38848) );
  NANDN U39337 ( .A(n39068), .B(n39069), .Z(n39067) );
  OR U39338 ( .A(n39070), .B(n39071), .Z(n39069) );
  NAND U39339 ( .A(n39071), .B(n39070), .Z(n39066) );
  ANDN U39340 ( .B(B[146]), .A(n73), .Z(n38850) );
  XNOR U39341 ( .A(n38858), .B(n39072), .Z(n38851) );
  XNOR U39342 ( .A(n38857), .B(n38855), .Z(n39072) );
  AND U39343 ( .A(n39073), .B(n39074), .Z(n38855) );
  NANDN U39344 ( .A(n39075), .B(n39076), .Z(n39074) );
  NANDN U39345 ( .A(n39077), .B(n39078), .Z(n39076) );
  NANDN U39346 ( .A(n39078), .B(n39077), .Z(n39073) );
  ANDN U39347 ( .B(B[147]), .A(n74), .Z(n38857) );
  XNOR U39348 ( .A(n38865), .B(n39079), .Z(n38858) );
  XNOR U39349 ( .A(n38864), .B(n38862), .Z(n39079) );
  AND U39350 ( .A(n39080), .B(n39081), .Z(n38862) );
  NANDN U39351 ( .A(n39082), .B(n39083), .Z(n39081) );
  OR U39352 ( .A(n39084), .B(n39085), .Z(n39083) );
  NAND U39353 ( .A(n39085), .B(n39084), .Z(n39080) );
  ANDN U39354 ( .B(B[148]), .A(n75), .Z(n38864) );
  XNOR U39355 ( .A(n38872), .B(n39086), .Z(n38865) );
  XNOR U39356 ( .A(n38871), .B(n38869), .Z(n39086) );
  AND U39357 ( .A(n39087), .B(n39088), .Z(n38869) );
  NANDN U39358 ( .A(n39089), .B(n39090), .Z(n39088) );
  NANDN U39359 ( .A(n39091), .B(n39092), .Z(n39090) );
  NANDN U39360 ( .A(n39092), .B(n39091), .Z(n39087) );
  ANDN U39361 ( .B(B[149]), .A(n76), .Z(n38871) );
  XNOR U39362 ( .A(n38879), .B(n39093), .Z(n38872) );
  XNOR U39363 ( .A(n38878), .B(n38876), .Z(n39093) );
  AND U39364 ( .A(n39094), .B(n39095), .Z(n38876) );
  NANDN U39365 ( .A(n39096), .B(n39097), .Z(n39095) );
  OR U39366 ( .A(n39098), .B(n39099), .Z(n39097) );
  NAND U39367 ( .A(n39099), .B(n39098), .Z(n39094) );
  ANDN U39368 ( .B(B[150]), .A(n77), .Z(n38878) );
  XNOR U39369 ( .A(n38886), .B(n39100), .Z(n38879) );
  XNOR U39370 ( .A(n38885), .B(n38883), .Z(n39100) );
  AND U39371 ( .A(n39101), .B(n39102), .Z(n38883) );
  NANDN U39372 ( .A(n39103), .B(n39104), .Z(n39102) );
  NANDN U39373 ( .A(n39105), .B(n39106), .Z(n39104) );
  NANDN U39374 ( .A(n39106), .B(n39105), .Z(n39101) );
  ANDN U39375 ( .B(B[151]), .A(n78), .Z(n38885) );
  XNOR U39376 ( .A(n38893), .B(n39107), .Z(n38886) );
  XNOR U39377 ( .A(n38892), .B(n38890), .Z(n39107) );
  AND U39378 ( .A(n39108), .B(n39109), .Z(n38890) );
  NANDN U39379 ( .A(n39110), .B(n39111), .Z(n39109) );
  OR U39380 ( .A(n39112), .B(n39113), .Z(n39111) );
  NAND U39381 ( .A(n39113), .B(n39112), .Z(n39108) );
  ANDN U39382 ( .B(B[152]), .A(n79), .Z(n38892) );
  XNOR U39383 ( .A(n38900), .B(n39114), .Z(n38893) );
  XNOR U39384 ( .A(n38899), .B(n38897), .Z(n39114) );
  AND U39385 ( .A(n39115), .B(n39116), .Z(n38897) );
  NANDN U39386 ( .A(n39117), .B(n39118), .Z(n39116) );
  NANDN U39387 ( .A(n39119), .B(n39120), .Z(n39118) );
  NANDN U39388 ( .A(n39120), .B(n39119), .Z(n39115) );
  ANDN U39389 ( .B(B[153]), .A(n80), .Z(n38899) );
  XNOR U39390 ( .A(n38907), .B(n39121), .Z(n38900) );
  XNOR U39391 ( .A(n38906), .B(n38904), .Z(n39121) );
  AND U39392 ( .A(n39122), .B(n39123), .Z(n38904) );
  NANDN U39393 ( .A(n39124), .B(n39125), .Z(n39123) );
  OR U39394 ( .A(n39126), .B(n39127), .Z(n39125) );
  NAND U39395 ( .A(n39127), .B(n39126), .Z(n39122) );
  ANDN U39396 ( .B(B[154]), .A(n81), .Z(n38906) );
  XNOR U39397 ( .A(n38914), .B(n39128), .Z(n38907) );
  XNOR U39398 ( .A(n38913), .B(n38911), .Z(n39128) );
  AND U39399 ( .A(n39129), .B(n39130), .Z(n38911) );
  NANDN U39400 ( .A(n39131), .B(n39132), .Z(n39130) );
  NAND U39401 ( .A(n39133), .B(n39134), .Z(n39132) );
  ANDN U39402 ( .B(B[155]), .A(n82), .Z(n38913) );
  XOR U39403 ( .A(n38920), .B(n39135), .Z(n38914) );
  XNOR U39404 ( .A(n38918), .B(n38921), .Z(n39135) );
  NAND U39405 ( .A(A[2]), .B(B[156]), .Z(n38921) );
  NANDN U39406 ( .A(n39136), .B(n39137), .Z(n38918) );
  AND U39407 ( .A(A[0]), .B(B[157]), .Z(n39137) );
  XNOR U39408 ( .A(n38923), .B(n39138), .Z(n38920) );
  NAND U39409 ( .A(A[0]), .B(B[158]), .Z(n39138) );
  NAND U39410 ( .A(B[157]), .B(A[1]), .Z(n38923) );
  NAND U39411 ( .A(n39139), .B(n39140), .Z(n480) );
  NANDN U39412 ( .A(n39141), .B(n39142), .Z(n39140) );
  OR U39413 ( .A(n39143), .B(n39144), .Z(n39142) );
  NAND U39414 ( .A(n39144), .B(n39143), .Z(n39139) );
  XOR U39415 ( .A(n482), .B(n481), .Z(\A1[155] ) );
  XOR U39416 ( .A(n39144), .B(n39145), .Z(n481) );
  XNOR U39417 ( .A(n39143), .B(n39141), .Z(n39145) );
  AND U39418 ( .A(n39146), .B(n39147), .Z(n39141) );
  NANDN U39419 ( .A(n39148), .B(n39149), .Z(n39147) );
  NANDN U39420 ( .A(n39150), .B(n39151), .Z(n39149) );
  NANDN U39421 ( .A(n39151), .B(n39150), .Z(n39146) );
  ANDN U39422 ( .B(B[126]), .A(n54), .Z(n39143) );
  XNOR U39423 ( .A(n38938), .B(n39152), .Z(n39144) );
  XNOR U39424 ( .A(n38937), .B(n38935), .Z(n39152) );
  AND U39425 ( .A(n39153), .B(n39154), .Z(n38935) );
  NANDN U39426 ( .A(n39155), .B(n39156), .Z(n39154) );
  OR U39427 ( .A(n39157), .B(n39158), .Z(n39156) );
  NAND U39428 ( .A(n39158), .B(n39157), .Z(n39153) );
  ANDN U39429 ( .B(B[127]), .A(n55), .Z(n38937) );
  XNOR U39430 ( .A(n38945), .B(n39159), .Z(n38938) );
  XNOR U39431 ( .A(n38944), .B(n38942), .Z(n39159) );
  AND U39432 ( .A(n39160), .B(n39161), .Z(n38942) );
  NANDN U39433 ( .A(n39162), .B(n39163), .Z(n39161) );
  NANDN U39434 ( .A(n39164), .B(n39165), .Z(n39163) );
  NANDN U39435 ( .A(n39165), .B(n39164), .Z(n39160) );
  ANDN U39436 ( .B(B[128]), .A(n56), .Z(n38944) );
  XNOR U39437 ( .A(n38952), .B(n39166), .Z(n38945) );
  XNOR U39438 ( .A(n38951), .B(n38949), .Z(n39166) );
  AND U39439 ( .A(n39167), .B(n39168), .Z(n38949) );
  NANDN U39440 ( .A(n39169), .B(n39170), .Z(n39168) );
  OR U39441 ( .A(n39171), .B(n39172), .Z(n39170) );
  NAND U39442 ( .A(n39172), .B(n39171), .Z(n39167) );
  ANDN U39443 ( .B(B[129]), .A(n57), .Z(n38951) );
  XNOR U39444 ( .A(n38959), .B(n39173), .Z(n38952) );
  XNOR U39445 ( .A(n38958), .B(n38956), .Z(n39173) );
  AND U39446 ( .A(n39174), .B(n39175), .Z(n38956) );
  NANDN U39447 ( .A(n39176), .B(n39177), .Z(n39175) );
  NANDN U39448 ( .A(n39178), .B(n39179), .Z(n39177) );
  NANDN U39449 ( .A(n39179), .B(n39178), .Z(n39174) );
  ANDN U39450 ( .B(B[130]), .A(n58), .Z(n38958) );
  XNOR U39451 ( .A(n38966), .B(n39180), .Z(n38959) );
  XNOR U39452 ( .A(n38965), .B(n38963), .Z(n39180) );
  AND U39453 ( .A(n39181), .B(n39182), .Z(n38963) );
  NANDN U39454 ( .A(n39183), .B(n39184), .Z(n39182) );
  OR U39455 ( .A(n39185), .B(n39186), .Z(n39184) );
  NAND U39456 ( .A(n39186), .B(n39185), .Z(n39181) );
  ANDN U39457 ( .B(B[131]), .A(n59), .Z(n38965) );
  XNOR U39458 ( .A(n38973), .B(n39187), .Z(n38966) );
  XNOR U39459 ( .A(n38972), .B(n38970), .Z(n39187) );
  AND U39460 ( .A(n39188), .B(n39189), .Z(n38970) );
  NANDN U39461 ( .A(n39190), .B(n39191), .Z(n39189) );
  NANDN U39462 ( .A(n39192), .B(n39193), .Z(n39191) );
  NANDN U39463 ( .A(n39193), .B(n39192), .Z(n39188) );
  ANDN U39464 ( .B(B[132]), .A(n60), .Z(n38972) );
  XNOR U39465 ( .A(n38980), .B(n39194), .Z(n38973) );
  XNOR U39466 ( .A(n38979), .B(n38977), .Z(n39194) );
  AND U39467 ( .A(n39195), .B(n39196), .Z(n38977) );
  NANDN U39468 ( .A(n39197), .B(n39198), .Z(n39196) );
  OR U39469 ( .A(n39199), .B(n39200), .Z(n39198) );
  NAND U39470 ( .A(n39200), .B(n39199), .Z(n39195) );
  ANDN U39471 ( .B(B[133]), .A(n61), .Z(n38979) );
  XNOR U39472 ( .A(n38987), .B(n39201), .Z(n38980) );
  XNOR U39473 ( .A(n38986), .B(n38984), .Z(n39201) );
  AND U39474 ( .A(n39202), .B(n39203), .Z(n38984) );
  NANDN U39475 ( .A(n39204), .B(n39205), .Z(n39203) );
  NANDN U39476 ( .A(n39206), .B(n39207), .Z(n39205) );
  NANDN U39477 ( .A(n39207), .B(n39206), .Z(n39202) );
  ANDN U39478 ( .B(B[134]), .A(n62), .Z(n38986) );
  XNOR U39479 ( .A(n38994), .B(n39208), .Z(n38987) );
  XNOR U39480 ( .A(n38993), .B(n38991), .Z(n39208) );
  AND U39481 ( .A(n39209), .B(n39210), .Z(n38991) );
  NANDN U39482 ( .A(n39211), .B(n39212), .Z(n39210) );
  OR U39483 ( .A(n39213), .B(n39214), .Z(n39212) );
  NAND U39484 ( .A(n39214), .B(n39213), .Z(n39209) );
  ANDN U39485 ( .B(B[135]), .A(n63), .Z(n38993) );
  XNOR U39486 ( .A(n39001), .B(n39215), .Z(n38994) );
  XNOR U39487 ( .A(n39000), .B(n38998), .Z(n39215) );
  AND U39488 ( .A(n39216), .B(n39217), .Z(n38998) );
  NANDN U39489 ( .A(n39218), .B(n39219), .Z(n39217) );
  NANDN U39490 ( .A(n39220), .B(n39221), .Z(n39219) );
  NANDN U39491 ( .A(n39221), .B(n39220), .Z(n39216) );
  ANDN U39492 ( .B(B[136]), .A(n64), .Z(n39000) );
  XNOR U39493 ( .A(n39008), .B(n39222), .Z(n39001) );
  XNOR U39494 ( .A(n39007), .B(n39005), .Z(n39222) );
  AND U39495 ( .A(n39223), .B(n39224), .Z(n39005) );
  NANDN U39496 ( .A(n39225), .B(n39226), .Z(n39224) );
  OR U39497 ( .A(n39227), .B(n39228), .Z(n39226) );
  NAND U39498 ( .A(n39228), .B(n39227), .Z(n39223) );
  ANDN U39499 ( .B(B[137]), .A(n65), .Z(n39007) );
  XNOR U39500 ( .A(n39015), .B(n39229), .Z(n39008) );
  XNOR U39501 ( .A(n39014), .B(n39012), .Z(n39229) );
  AND U39502 ( .A(n39230), .B(n39231), .Z(n39012) );
  NANDN U39503 ( .A(n39232), .B(n39233), .Z(n39231) );
  NANDN U39504 ( .A(n39234), .B(n39235), .Z(n39233) );
  NANDN U39505 ( .A(n39235), .B(n39234), .Z(n39230) );
  ANDN U39506 ( .B(B[138]), .A(n66), .Z(n39014) );
  XNOR U39507 ( .A(n39022), .B(n39236), .Z(n39015) );
  XNOR U39508 ( .A(n39021), .B(n39019), .Z(n39236) );
  AND U39509 ( .A(n39237), .B(n39238), .Z(n39019) );
  NANDN U39510 ( .A(n39239), .B(n39240), .Z(n39238) );
  OR U39511 ( .A(n39241), .B(n39242), .Z(n39240) );
  NAND U39512 ( .A(n39242), .B(n39241), .Z(n39237) );
  ANDN U39513 ( .B(B[139]), .A(n67), .Z(n39021) );
  XNOR U39514 ( .A(n39029), .B(n39243), .Z(n39022) );
  XNOR U39515 ( .A(n39028), .B(n39026), .Z(n39243) );
  AND U39516 ( .A(n39244), .B(n39245), .Z(n39026) );
  NANDN U39517 ( .A(n39246), .B(n39247), .Z(n39245) );
  NANDN U39518 ( .A(n39248), .B(n39249), .Z(n39247) );
  NANDN U39519 ( .A(n39249), .B(n39248), .Z(n39244) );
  ANDN U39520 ( .B(B[140]), .A(n68), .Z(n39028) );
  XNOR U39521 ( .A(n39036), .B(n39250), .Z(n39029) );
  XNOR U39522 ( .A(n39035), .B(n39033), .Z(n39250) );
  AND U39523 ( .A(n39251), .B(n39252), .Z(n39033) );
  NANDN U39524 ( .A(n39253), .B(n39254), .Z(n39252) );
  OR U39525 ( .A(n39255), .B(n39256), .Z(n39254) );
  NAND U39526 ( .A(n39256), .B(n39255), .Z(n39251) );
  ANDN U39527 ( .B(B[141]), .A(n69), .Z(n39035) );
  XNOR U39528 ( .A(n39043), .B(n39257), .Z(n39036) );
  XNOR U39529 ( .A(n39042), .B(n39040), .Z(n39257) );
  AND U39530 ( .A(n39258), .B(n39259), .Z(n39040) );
  NANDN U39531 ( .A(n39260), .B(n39261), .Z(n39259) );
  NANDN U39532 ( .A(n39262), .B(n39263), .Z(n39261) );
  NANDN U39533 ( .A(n39263), .B(n39262), .Z(n39258) );
  ANDN U39534 ( .B(B[142]), .A(n70), .Z(n39042) );
  XNOR U39535 ( .A(n39050), .B(n39264), .Z(n39043) );
  XNOR U39536 ( .A(n39049), .B(n39047), .Z(n39264) );
  AND U39537 ( .A(n39265), .B(n39266), .Z(n39047) );
  NANDN U39538 ( .A(n39267), .B(n39268), .Z(n39266) );
  OR U39539 ( .A(n39269), .B(n39270), .Z(n39268) );
  NAND U39540 ( .A(n39270), .B(n39269), .Z(n39265) );
  ANDN U39541 ( .B(B[143]), .A(n71), .Z(n39049) );
  XNOR U39542 ( .A(n39057), .B(n39271), .Z(n39050) );
  XNOR U39543 ( .A(n39056), .B(n39054), .Z(n39271) );
  AND U39544 ( .A(n39272), .B(n39273), .Z(n39054) );
  NANDN U39545 ( .A(n39274), .B(n39275), .Z(n39273) );
  NANDN U39546 ( .A(n39276), .B(n39277), .Z(n39275) );
  NANDN U39547 ( .A(n39277), .B(n39276), .Z(n39272) );
  ANDN U39548 ( .B(B[144]), .A(n72), .Z(n39056) );
  XNOR U39549 ( .A(n39064), .B(n39278), .Z(n39057) );
  XNOR U39550 ( .A(n39063), .B(n39061), .Z(n39278) );
  AND U39551 ( .A(n39279), .B(n39280), .Z(n39061) );
  NANDN U39552 ( .A(n39281), .B(n39282), .Z(n39280) );
  OR U39553 ( .A(n39283), .B(n39284), .Z(n39282) );
  NAND U39554 ( .A(n39284), .B(n39283), .Z(n39279) );
  ANDN U39555 ( .B(B[145]), .A(n73), .Z(n39063) );
  XNOR U39556 ( .A(n39071), .B(n39285), .Z(n39064) );
  XNOR U39557 ( .A(n39070), .B(n39068), .Z(n39285) );
  AND U39558 ( .A(n39286), .B(n39287), .Z(n39068) );
  NANDN U39559 ( .A(n39288), .B(n39289), .Z(n39287) );
  NANDN U39560 ( .A(n39290), .B(n39291), .Z(n39289) );
  NANDN U39561 ( .A(n39291), .B(n39290), .Z(n39286) );
  ANDN U39562 ( .B(B[146]), .A(n74), .Z(n39070) );
  XNOR U39563 ( .A(n39078), .B(n39292), .Z(n39071) );
  XNOR U39564 ( .A(n39077), .B(n39075), .Z(n39292) );
  AND U39565 ( .A(n39293), .B(n39294), .Z(n39075) );
  NANDN U39566 ( .A(n39295), .B(n39296), .Z(n39294) );
  OR U39567 ( .A(n39297), .B(n39298), .Z(n39296) );
  NAND U39568 ( .A(n39298), .B(n39297), .Z(n39293) );
  ANDN U39569 ( .B(B[147]), .A(n75), .Z(n39077) );
  XNOR U39570 ( .A(n39085), .B(n39299), .Z(n39078) );
  XNOR U39571 ( .A(n39084), .B(n39082), .Z(n39299) );
  AND U39572 ( .A(n39300), .B(n39301), .Z(n39082) );
  NANDN U39573 ( .A(n39302), .B(n39303), .Z(n39301) );
  NANDN U39574 ( .A(n39304), .B(n39305), .Z(n39303) );
  NANDN U39575 ( .A(n39305), .B(n39304), .Z(n39300) );
  ANDN U39576 ( .B(B[148]), .A(n76), .Z(n39084) );
  XNOR U39577 ( .A(n39092), .B(n39306), .Z(n39085) );
  XNOR U39578 ( .A(n39091), .B(n39089), .Z(n39306) );
  AND U39579 ( .A(n39307), .B(n39308), .Z(n39089) );
  NANDN U39580 ( .A(n39309), .B(n39310), .Z(n39308) );
  OR U39581 ( .A(n39311), .B(n39312), .Z(n39310) );
  NAND U39582 ( .A(n39312), .B(n39311), .Z(n39307) );
  ANDN U39583 ( .B(B[149]), .A(n77), .Z(n39091) );
  XNOR U39584 ( .A(n39099), .B(n39313), .Z(n39092) );
  XNOR U39585 ( .A(n39098), .B(n39096), .Z(n39313) );
  AND U39586 ( .A(n39314), .B(n39315), .Z(n39096) );
  NANDN U39587 ( .A(n39316), .B(n39317), .Z(n39315) );
  NANDN U39588 ( .A(n39318), .B(n39319), .Z(n39317) );
  NANDN U39589 ( .A(n39319), .B(n39318), .Z(n39314) );
  ANDN U39590 ( .B(B[150]), .A(n78), .Z(n39098) );
  XNOR U39591 ( .A(n39106), .B(n39320), .Z(n39099) );
  XNOR U39592 ( .A(n39105), .B(n39103), .Z(n39320) );
  AND U39593 ( .A(n39321), .B(n39322), .Z(n39103) );
  NANDN U39594 ( .A(n39323), .B(n39324), .Z(n39322) );
  OR U39595 ( .A(n39325), .B(n39326), .Z(n39324) );
  NAND U39596 ( .A(n39326), .B(n39325), .Z(n39321) );
  ANDN U39597 ( .B(B[151]), .A(n79), .Z(n39105) );
  XNOR U39598 ( .A(n39113), .B(n39327), .Z(n39106) );
  XNOR U39599 ( .A(n39112), .B(n39110), .Z(n39327) );
  AND U39600 ( .A(n39328), .B(n39329), .Z(n39110) );
  NANDN U39601 ( .A(n39330), .B(n39331), .Z(n39329) );
  NANDN U39602 ( .A(n39332), .B(n39333), .Z(n39331) );
  NANDN U39603 ( .A(n39333), .B(n39332), .Z(n39328) );
  ANDN U39604 ( .B(B[152]), .A(n80), .Z(n39112) );
  XNOR U39605 ( .A(n39120), .B(n39334), .Z(n39113) );
  XNOR U39606 ( .A(n39119), .B(n39117), .Z(n39334) );
  AND U39607 ( .A(n39335), .B(n39336), .Z(n39117) );
  NANDN U39608 ( .A(n39337), .B(n39338), .Z(n39336) );
  OR U39609 ( .A(n39339), .B(n39340), .Z(n39338) );
  NAND U39610 ( .A(n39340), .B(n39339), .Z(n39335) );
  ANDN U39611 ( .B(B[153]), .A(n81), .Z(n39119) );
  XNOR U39612 ( .A(n39127), .B(n39341), .Z(n39120) );
  XNOR U39613 ( .A(n39126), .B(n39124), .Z(n39341) );
  AND U39614 ( .A(n39342), .B(n39343), .Z(n39124) );
  NANDN U39615 ( .A(n39344), .B(n39345), .Z(n39343) );
  NAND U39616 ( .A(n39346), .B(n39347), .Z(n39345) );
  ANDN U39617 ( .B(B[154]), .A(n82), .Z(n39126) );
  XOR U39618 ( .A(n39133), .B(n39348), .Z(n39127) );
  XNOR U39619 ( .A(n39131), .B(n39134), .Z(n39348) );
  NAND U39620 ( .A(A[2]), .B(B[155]), .Z(n39134) );
  NANDN U39621 ( .A(n39349), .B(n39350), .Z(n39131) );
  AND U39622 ( .A(A[0]), .B(B[156]), .Z(n39350) );
  XNOR U39623 ( .A(n39136), .B(n39351), .Z(n39133) );
  NAND U39624 ( .A(A[0]), .B(B[157]), .Z(n39351) );
  NAND U39625 ( .A(B[156]), .B(A[1]), .Z(n39136) );
  NAND U39626 ( .A(n39352), .B(n39353), .Z(n482) );
  NANDN U39627 ( .A(n39354), .B(n39355), .Z(n39353) );
  OR U39628 ( .A(n39356), .B(n39357), .Z(n39355) );
  NAND U39629 ( .A(n39357), .B(n39356), .Z(n39352) );
  XOR U39630 ( .A(n484), .B(n483), .Z(\A1[154] ) );
  XOR U39631 ( .A(n39357), .B(n39358), .Z(n483) );
  XNOR U39632 ( .A(n39356), .B(n39354), .Z(n39358) );
  AND U39633 ( .A(n39359), .B(n39360), .Z(n39354) );
  NANDN U39634 ( .A(n39361), .B(n39362), .Z(n39360) );
  NANDN U39635 ( .A(n39363), .B(n39364), .Z(n39362) );
  NANDN U39636 ( .A(n39364), .B(n39363), .Z(n39359) );
  ANDN U39637 ( .B(B[125]), .A(n54), .Z(n39356) );
  XNOR U39638 ( .A(n39151), .B(n39365), .Z(n39357) );
  XNOR U39639 ( .A(n39150), .B(n39148), .Z(n39365) );
  AND U39640 ( .A(n39366), .B(n39367), .Z(n39148) );
  NANDN U39641 ( .A(n39368), .B(n39369), .Z(n39367) );
  OR U39642 ( .A(n39370), .B(n39371), .Z(n39369) );
  NAND U39643 ( .A(n39371), .B(n39370), .Z(n39366) );
  ANDN U39644 ( .B(B[126]), .A(n55), .Z(n39150) );
  XNOR U39645 ( .A(n39158), .B(n39372), .Z(n39151) );
  XNOR U39646 ( .A(n39157), .B(n39155), .Z(n39372) );
  AND U39647 ( .A(n39373), .B(n39374), .Z(n39155) );
  NANDN U39648 ( .A(n39375), .B(n39376), .Z(n39374) );
  NANDN U39649 ( .A(n39377), .B(n39378), .Z(n39376) );
  NANDN U39650 ( .A(n39378), .B(n39377), .Z(n39373) );
  ANDN U39651 ( .B(B[127]), .A(n56), .Z(n39157) );
  XNOR U39652 ( .A(n39165), .B(n39379), .Z(n39158) );
  XNOR U39653 ( .A(n39164), .B(n39162), .Z(n39379) );
  AND U39654 ( .A(n39380), .B(n39381), .Z(n39162) );
  NANDN U39655 ( .A(n39382), .B(n39383), .Z(n39381) );
  OR U39656 ( .A(n39384), .B(n39385), .Z(n39383) );
  NAND U39657 ( .A(n39385), .B(n39384), .Z(n39380) );
  ANDN U39658 ( .B(B[128]), .A(n57), .Z(n39164) );
  XNOR U39659 ( .A(n39172), .B(n39386), .Z(n39165) );
  XNOR U39660 ( .A(n39171), .B(n39169), .Z(n39386) );
  AND U39661 ( .A(n39387), .B(n39388), .Z(n39169) );
  NANDN U39662 ( .A(n39389), .B(n39390), .Z(n39388) );
  NANDN U39663 ( .A(n39391), .B(n39392), .Z(n39390) );
  NANDN U39664 ( .A(n39392), .B(n39391), .Z(n39387) );
  ANDN U39665 ( .B(B[129]), .A(n58), .Z(n39171) );
  XNOR U39666 ( .A(n39179), .B(n39393), .Z(n39172) );
  XNOR U39667 ( .A(n39178), .B(n39176), .Z(n39393) );
  AND U39668 ( .A(n39394), .B(n39395), .Z(n39176) );
  NANDN U39669 ( .A(n39396), .B(n39397), .Z(n39395) );
  OR U39670 ( .A(n39398), .B(n39399), .Z(n39397) );
  NAND U39671 ( .A(n39399), .B(n39398), .Z(n39394) );
  ANDN U39672 ( .B(B[130]), .A(n59), .Z(n39178) );
  XNOR U39673 ( .A(n39186), .B(n39400), .Z(n39179) );
  XNOR U39674 ( .A(n39185), .B(n39183), .Z(n39400) );
  AND U39675 ( .A(n39401), .B(n39402), .Z(n39183) );
  NANDN U39676 ( .A(n39403), .B(n39404), .Z(n39402) );
  NANDN U39677 ( .A(n39405), .B(n39406), .Z(n39404) );
  NANDN U39678 ( .A(n39406), .B(n39405), .Z(n39401) );
  ANDN U39679 ( .B(B[131]), .A(n60), .Z(n39185) );
  XNOR U39680 ( .A(n39193), .B(n39407), .Z(n39186) );
  XNOR U39681 ( .A(n39192), .B(n39190), .Z(n39407) );
  AND U39682 ( .A(n39408), .B(n39409), .Z(n39190) );
  NANDN U39683 ( .A(n39410), .B(n39411), .Z(n39409) );
  OR U39684 ( .A(n39412), .B(n39413), .Z(n39411) );
  NAND U39685 ( .A(n39413), .B(n39412), .Z(n39408) );
  ANDN U39686 ( .B(B[132]), .A(n61), .Z(n39192) );
  XNOR U39687 ( .A(n39200), .B(n39414), .Z(n39193) );
  XNOR U39688 ( .A(n39199), .B(n39197), .Z(n39414) );
  AND U39689 ( .A(n39415), .B(n39416), .Z(n39197) );
  NANDN U39690 ( .A(n39417), .B(n39418), .Z(n39416) );
  NANDN U39691 ( .A(n39419), .B(n39420), .Z(n39418) );
  NANDN U39692 ( .A(n39420), .B(n39419), .Z(n39415) );
  ANDN U39693 ( .B(B[133]), .A(n62), .Z(n39199) );
  XNOR U39694 ( .A(n39207), .B(n39421), .Z(n39200) );
  XNOR U39695 ( .A(n39206), .B(n39204), .Z(n39421) );
  AND U39696 ( .A(n39422), .B(n39423), .Z(n39204) );
  NANDN U39697 ( .A(n39424), .B(n39425), .Z(n39423) );
  OR U39698 ( .A(n39426), .B(n39427), .Z(n39425) );
  NAND U39699 ( .A(n39427), .B(n39426), .Z(n39422) );
  ANDN U39700 ( .B(B[134]), .A(n63), .Z(n39206) );
  XNOR U39701 ( .A(n39214), .B(n39428), .Z(n39207) );
  XNOR U39702 ( .A(n39213), .B(n39211), .Z(n39428) );
  AND U39703 ( .A(n39429), .B(n39430), .Z(n39211) );
  NANDN U39704 ( .A(n39431), .B(n39432), .Z(n39430) );
  NANDN U39705 ( .A(n39433), .B(n39434), .Z(n39432) );
  NANDN U39706 ( .A(n39434), .B(n39433), .Z(n39429) );
  ANDN U39707 ( .B(B[135]), .A(n64), .Z(n39213) );
  XNOR U39708 ( .A(n39221), .B(n39435), .Z(n39214) );
  XNOR U39709 ( .A(n39220), .B(n39218), .Z(n39435) );
  AND U39710 ( .A(n39436), .B(n39437), .Z(n39218) );
  NANDN U39711 ( .A(n39438), .B(n39439), .Z(n39437) );
  OR U39712 ( .A(n39440), .B(n39441), .Z(n39439) );
  NAND U39713 ( .A(n39441), .B(n39440), .Z(n39436) );
  ANDN U39714 ( .B(B[136]), .A(n65), .Z(n39220) );
  XNOR U39715 ( .A(n39228), .B(n39442), .Z(n39221) );
  XNOR U39716 ( .A(n39227), .B(n39225), .Z(n39442) );
  AND U39717 ( .A(n39443), .B(n39444), .Z(n39225) );
  NANDN U39718 ( .A(n39445), .B(n39446), .Z(n39444) );
  NANDN U39719 ( .A(n39447), .B(n39448), .Z(n39446) );
  NANDN U39720 ( .A(n39448), .B(n39447), .Z(n39443) );
  ANDN U39721 ( .B(B[137]), .A(n66), .Z(n39227) );
  XNOR U39722 ( .A(n39235), .B(n39449), .Z(n39228) );
  XNOR U39723 ( .A(n39234), .B(n39232), .Z(n39449) );
  AND U39724 ( .A(n39450), .B(n39451), .Z(n39232) );
  NANDN U39725 ( .A(n39452), .B(n39453), .Z(n39451) );
  OR U39726 ( .A(n39454), .B(n39455), .Z(n39453) );
  NAND U39727 ( .A(n39455), .B(n39454), .Z(n39450) );
  ANDN U39728 ( .B(B[138]), .A(n67), .Z(n39234) );
  XNOR U39729 ( .A(n39242), .B(n39456), .Z(n39235) );
  XNOR U39730 ( .A(n39241), .B(n39239), .Z(n39456) );
  AND U39731 ( .A(n39457), .B(n39458), .Z(n39239) );
  NANDN U39732 ( .A(n39459), .B(n39460), .Z(n39458) );
  NANDN U39733 ( .A(n39461), .B(n39462), .Z(n39460) );
  NANDN U39734 ( .A(n39462), .B(n39461), .Z(n39457) );
  ANDN U39735 ( .B(B[139]), .A(n68), .Z(n39241) );
  XNOR U39736 ( .A(n39249), .B(n39463), .Z(n39242) );
  XNOR U39737 ( .A(n39248), .B(n39246), .Z(n39463) );
  AND U39738 ( .A(n39464), .B(n39465), .Z(n39246) );
  NANDN U39739 ( .A(n39466), .B(n39467), .Z(n39465) );
  OR U39740 ( .A(n39468), .B(n39469), .Z(n39467) );
  NAND U39741 ( .A(n39469), .B(n39468), .Z(n39464) );
  ANDN U39742 ( .B(B[140]), .A(n69), .Z(n39248) );
  XNOR U39743 ( .A(n39256), .B(n39470), .Z(n39249) );
  XNOR U39744 ( .A(n39255), .B(n39253), .Z(n39470) );
  AND U39745 ( .A(n39471), .B(n39472), .Z(n39253) );
  NANDN U39746 ( .A(n39473), .B(n39474), .Z(n39472) );
  NANDN U39747 ( .A(n39475), .B(n39476), .Z(n39474) );
  NANDN U39748 ( .A(n39476), .B(n39475), .Z(n39471) );
  ANDN U39749 ( .B(B[141]), .A(n70), .Z(n39255) );
  XNOR U39750 ( .A(n39263), .B(n39477), .Z(n39256) );
  XNOR U39751 ( .A(n39262), .B(n39260), .Z(n39477) );
  AND U39752 ( .A(n39478), .B(n39479), .Z(n39260) );
  NANDN U39753 ( .A(n39480), .B(n39481), .Z(n39479) );
  OR U39754 ( .A(n39482), .B(n39483), .Z(n39481) );
  NAND U39755 ( .A(n39483), .B(n39482), .Z(n39478) );
  ANDN U39756 ( .B(B[142]), .A(n71), .Z(n39262) );
  XNOR U39757 ( .A(n39270), .B(n39484), .Z(n39263) );
  XNOR U39758 ( .A(n39269), .B(n39267), .Z(n39484) );
  AND U39759 ( .A(n39485), .B(n39486), .Z(n39267) );
  NANDN U39760 ( .A(n39487), .B(n39488), .Z(n39486) );
  NANDN U39761 ( .A(n39489), .B(n39490), .Z(n39488) );
  NANDN U39762 ( .A(n39490), .B(n39489), .Z(n39485) );
  ANDN U39763 ( .B(B[143]), .A(n72), .Z(n39269) );
  XNOR U39764 ( .A(n39277), .B(n39491), .Z(n39270) );
  XNOR U39765 ( .A(n39276), .B(n39274), .Z(n39491) );
  AND U39766 ( .A(n39492), .B(n39493), .Z(n39274) );
  NANDN U39767 ( .A(n39494), .B(n39495), .Z(n39493) );
  OR U39768 ( .A(n39496), .B(n39497), .Z(n39495) );
  NAND U39769 ( .A(n39497), .B(n39496), .Z(n39492) );
  ANDN U39770 ( .B(B[144]), .A(n73), .Z(n39276) );
  XNOR U39771 ( .A(n39284), .B(n39498), .Z(n39277) );
  XNOR U39772 ( .A(n39283), .B(n39281), .Z(n39498) );
  AND U39773 ( .A(n39499), .B(n39500), .Z(n39281) );
  NANDN U39774 ( .A(n39501), .B(n39502), .Z(n39500) );
  NANDN U39775 ( .A(n39503), .B(n39504), .Z(n39502) );
  NANDN U39776 ( .A(n39504), .B(n39503), .Z(n39499) );
  ANDN U39777 ( .B(B[145]), .A(n74), .Z(n39283) );
  XNOR U39778 ( .A(n39291), .B(n39505), .Z(n39284) );
  XNOR U39779 ( .A(n39290), .B(n39288), .Z(n39505) );
  AND U39780 ( .A(n39506), .B(n39507), .Z(n39288) );
  NANDN U39781 ( .A(n39508), .B(n39509), .Z(n39507) );
  OR U39782 ( .A(n39510), .B(n39511), .Z(n39509) );
  NAND U39783 ( .A(n39511), .B(n39510), .Z(n39506) );
  ANDN U39784 ( .B(B[146]), .A(n75), .Z(n39290) );
  XNOR U39785 ( .A(n39298), .B(n39512), .Z(n39291) );
  XNOR U39786 ( .A(n39297), .B(n39295), .Z(n39512) );
  AND U39787 ( .A(n39513), .B(n39514), .Z(n39295) );
  NANDN U39788 ( .A(n39515), .B(n39516), .Z(n39514) );
  NANDN U39789 ( .A(n39517), .B(n39518), .Z(n39516) );
  NANDN U39790 ( .A(n39518), .B(n39517), .Z(n39513) );
  ANDN U39791 ( .B(B[147]), .A(n76), .Z(n39297) );
  XNOR U39792 ( .A(n39305), .B(n39519), .Z(n39298) );
  XNOR U39793 ( .A(n39304), .B(n39302), .Z(n39519) );
  AND U39794 ( .A(n39520), .B(n39521), .Z(n39302) );
  NANDN U39795 ( .A(n39522), .B(n39523), .Z(n39521) );
  OR U39796 ( .A(n39524), .B(n39525), .Z(n39523) );
  NAND U39797 ( .A(n39525), .B(n39524), .Z(n39520) );
  ANDN U39798 ( .B(B[148]), .A(n77), .Z(n39304) );
  XNOR U39799 ( .A(n39312), .B(n39526), .Z(n39305) );
  XNOR U39800 ( .A(n39311), .B(n39309), .Z(n39526) );
  AND U39801 ( .A(n39527), .B(n39528), .Z(n39309) );
  NANDN U39802 ( .A(n39529), .B(n39530), .Z(n39528) );
  NANDN U39803 ( .A(n39531), .B(n39532), .Z(n39530) );
  NANDN U39804 ( .A(n39532), .B(n39531), .Z(n39527) );
  ANDN U39805 ( .B(B[149]), .A(n78), .Z(n39311) );
  XNOR U39806 ( .A(n39319), .B(n39533), .Z(n39312) );
  XNOR U39807 ( .A(n39318), .B(n39316), .Z(n39533) );
  AND U39808 ( .A(n39534), .B(n39535), .Z(n39316) );
  NANDN U39809 ( .A(n39536), .B(n39537), .Z(n39535) );
  OR U39810 ( .A(n39538), .B(n39539), .Z(n39537) );
  NAND U39811 ( .A(n39539), .B(n39538), .Z(n39534) );
  ANDN U39812 ( .B(B[150]), .A(n79), .Z(n39318) );
  XNOR U39813 ( .A(n39326), .B(n39540), .Z(n39319) );
  XNOR U39814 ( .A(n39325), .B(n39323), .Z(n39540) );
  AND U39815 ( .A(n39541), .B(n39542), .Z(n39323) );
  NANDN U39816 ( .A(n39543), .B(n39544), .Z(n39542) );
  NANDN U39817 ( .A(n39545), .B(n39546), .Z(n39544) );
  NANDN U39818 ( .A(n39546), .B(n39545), .Z(n39541) );
  ANDN U39819 ( .B(B[151]), .A(n80), .Z(n39325) );
  XNOR U39820 ( .A(n39333), .B(n39547), .Z(n39326) );
  XNOR U39821 ( .A(n39332), .B(n39330), .Z(n39547) );
  AND U39822 ( .A(n39548), .B(n39549), .Z(n39330) );
  NANDN U39823 ( .A(n39550), .B(n39551), .Z(n39549) );
  OR U39824 ( .A(n39552), .B(n39553), .Z(n39551) );
  NAND U39825 ( .A(n39553), .B(n39552), .Z(n39548) );
  ANDN U39826 ( .B(B[152]), .A(n81), .Z(n39332) );
  XNOR U39827 ( .A(n39340), .B(n39554), .Z(n39333) );
  XNOR U39828 ( .A(n39339), .B(n39337), .Z(n39554) );
  AND U39829 ( .A(n39555), .B(n39556), .Z(n39337) );
  NANDN U39830 ( .A(n39557), .B(n39558), .Z(n39556) );
  NAND U39831 ( .A(n39559), .B(n39560), .Z(n39558) );
  ANDN U39832 ( .B(B[153]), .A(n82), .Z(n39339) );
  XOR U39833 ( .A(n39346), .B(n39561), .Z(n39340) );
  XNOR U39834 ( .A(n39344), .B(n39347), .Z(n39561) );
  NAND U39835 ( .A(A[2]), .B(B[154]), .Z(n39347) );
  NANDN U39836 ( .A(n39562), .B(n39563), .Z(n39344) );
  AND U39837 ( .A(A[0]), .B(B[155]), .Z(n39563) );
  XNOR U39838 ( .A(n39349), .B(n39564), .Z(n39346) );
  NAND U39839 ( .A(A[0]), .B(B[156]), .Z(n39564) );
  NAND U39840 ( .A(B[155]), .B(A[1]), .Z(n39349) );
  NAND U39841 ( .A(n39565), .B(n39566), .Z(n484) );
  NANDN U39842 ( .A(n39567), .B(n39568), .Z(n39566) );
  OR U39843 ( .A(n39569), .B(n39570), .Z(n39568) );
  NAND U39844 ( .A(n39570), .B(n39569), .Z(n39565) );
  XOR U39845 ( .A(n486), .B(n485), .Z(\A1[153] ) );
  XOR U39846 ( .A(n39570), .B(n39571), .Z(n485) );
  XNOR U39847 ( .A(n39569), .B(n39567), .Z(n39571) );
  AND U39848 ( .A(n39572), .B(n39573), .Z(n39567) );
  NANDN U39849 ( .A(n39574), .B(n39575), .Z(n39573) );
  NANDN U39850 ( .A(n39576), .B(n39577), .Z(n39575) );
  NANDN U39851 ( .A(n39577), .B(n39576), .Z(n39572) );
  ANDN U39852 ( .B(B[124]), .A(n54), .Z(n39569) );
  XNOR U39853 ( .A(n39364), .B(n39578), .Z(n39570) );
  XNOR U39854 ( .A(n39363), .B(n39361), .Z(n39578) );
  AND U39855 ( .A(n39579), .B(n39580), .Z(n39361) );
  NANDN U39856 ( .A(n39581), .B(n39582), .Z(n39580) );
  OR U39857 ( .A(n39583), .B(n39584), .Z(n39582) );
  NAND U39858 ( .A(n39584), .B(n39583), .Z(n39579) );
  ANDN U39859 ( .B(B[125]), .A(n55), .Z(n39363) );
  XNOR U39860 ( .A(n39371), .B(n39585), .Z(n39364) );
  XNOR U39861 ( .A(n39370), .B(n39368), .Z(n39585) );
  AND U39862 ( .A(n39586), .B(n39587), .Z(n39368) );
  NANDN U39863 ( .A(n39588), .B(n39589), .Z(n39587) );
  NANDN U39864 ( .A(n39590), .B(n39591), .Z(n39589) );
  NANDN U39865 ( .A(n39591), .B(n39590), .Z(n39586) );
  ANDN U39866 ( .B(B[126]), .A(n56), .Z(n39370) );
  XNOR U39867 ( .A(n39378), .B(n39592), .Z(n39371) );
  XNOR U39868 ( .A(n39377), .B(n39375), .Z(n39592) );
  AND U39869 ( .A(n39593), .B(n39594), .Z(n39375) );
  NANDN U39870 ( .A(n39595), .B(n39596), .Z(n39594) );
  OR U39871 ( .A(n39597), .B(n39598), .Z(n39596) );
  NAND U39872 ( .A(n39598), .B(n39597), .Z(n39593) );
  ANDN U39873 ( .B(B[127]), .A(n57), .Z(n39377) );
  XNOR U39874 ( .A(n39385), .B(n39599), .Z(n39378) );
  XNOR U39875 ( .A(n39384), .B(n39382), .Z(n39599) );
  AND U39876 ( .A(n39600), .B(n39601), .Z(n39382) );
  NANDN U39877 ( .A(n39602), .B(n39603), .Z(n39601) );
  NANDN U39878 ( .A(n39604), .B(n39605), .Z(n39603) );
  NANDN U39879 ( .A(n39605), .B(n39604), .Z(n39600) );
  ANDN U39880 ( .B(B[128]), .A(n58), .Z(n39384) );
  XNOR U39881 ( .A(n39392), .B(n39606), .Z(n39385) );
  XNOR U39882 ( .A(n39391), .B(n39389), .Z(n39606) );
  AND U39883 ( .A(n39607), .B(n39608), .Z(n39389) );
  NANDN U39884 ( .A(n39609), .B(n39610), .Z(n39608) );
  OR U39885 ( .A(n39611), .B(n39612), .Z(n39610) );
  NAND U39886 ( .A(n39612), .B(n39611), .Z(n39607) );
  ANDN U39887 ( .B(B[129]), .A(n59), .Z(n39391) );
  XNOR U39888 ( .A(n39399), .B(n39613), .Z(n39392) );
  XNOR U39889 ( .A(n39398), .B(n39396), .Z(n39613) );
  AND U39890 ( .A(n39614), .B(n39615), .Z(n39396) );
  NANDN U39891 ( .A(n39616), .B(n39617), .Z(n39615) );
  NANDN U39892 ( .A(n39618), .B(n39619), .Z(n39617) );
  NANDN U39893 ( .A(n39619), .B(n39618), .Z(n39614) );
  ANDN U39894 ( .B(B[130]), .A(n60), .Z(n39398) );
  XNOR U39895 ( .A(n39406), .B(n39620), .Z(n39399) );
  XNOR U39896 ( .A(n39405), .B(n39403), .Z(n39620) );
  AND U39897 ( .A(n39621), .B(n39622), .Z(n39403) );
  NANDN U39898 ( .A(n39623), .B(n39624), .Z(n39622) );
  OR U39899 ( .A(n39625), .B(n39626), .Z(n39624) );
  NAND U39900 ( .A(n39626), .B(n39625), .Z(n39621) );
  ANDN U39901 ( .B(B[131]), .A(n61), .Z(n39405) );
  XNOR U39902 ( .A(n39413), .B(n39627), .Z(n39406) );
  XNOR U39903 ( .A(n39412), .B(n39410), .Z(n39627) );
  AND U39904 ( .A(n39628), .B(n39629), .Z(n39410) );
  NANDN U39905 ( .A(n39630), .B(n39631), .Z(n39629) );
  NANDN U39906 ( .A(n39632), .B(n39633), .Z(n39631) );
  NANDN U39907 ( .A(n39633), .B(n39632), .Z(n39628) );
  ANDN U39908 ( .B(B[132]), .A(n62), .Z(n39412) );
  XNOR U39909 ( .A(n39420), .B(n39634), .Z(n39413) );
  XNOR U39910 ( .A(n39419), .B(n39417), .Z(n39634) );
  AND U39911 ( .A(n39635), .B(n39636), .Z(n39417) );
  NANDN U39912 ( .A(n39637), .B(n39638), .Z(n39636) );
  OR U39913 ( .A(n39639), .B(n39640), .Z(n39638) );
  NAND U39914 ( .A(n39640), .B(n39639), .Z(n39635) );
  ANDN U39915 ( .B(B[133]), .A(n63), .Z(n39419) );
  XNOR U39916 ( .A(n39427), .B(n39641), .Z(n39420) );
  XNOR U39917 ( .A(n39426), .B(n39424), .Z(n39641) );
  AND U39918 ( .A(n39642), .B(n39643), .Z(n39424) );
  NANDN U39919 ( .A(n39644), .B(n39645), .Z(n39643) );
  NANDN U39920 ( .A(n39646), .B(n39647), .Z(n39645) );
  NANDN U39921 ( .A(n39647), .B(n39646), .Z(n39642) );
  ANDN U39922 ( .B(B[134]), .A(n64), .Z(n39426) );
  XNOR U39923 ( .A(n39434), .B(n39648), .Z(n39427) );
  XNOR U39924 ( .A(n39433), .B(n39431), .Z(n39648) );
  AND U39925 ( .A(n39649), .B(n39650), .Z(n39431) );
  NANDN U39926 ( .A(n39651), .B(n39652), .Z(n39650) );
  OR U39927 ( .A(n39653), .B(n39654), .Z(n39652) );
  NAND U39928 ( .A(n39654), .B(n39653), .Z(n39649) );
  ANDN U39929 ( .B(B[135]), .A(n65), .Z(n39433) );
  XNOR U39930 ( .A(n39441), .B(n39655), .Z(n39434) );
  XNOR U39931 ( .A(n39440), .B(n39438), .Z(n39655) );
  AND U39932 ( .A(n39656), .B(n39657), .Z(n39438) );
  NANDN U39933 ( .A(n39658), .B(n39659), .Z(n39657) );
  NANDN U39934 ( .A(n39660), .B(n39661), .Z(n39659) );
  NANDN U39935 ( .A(n39661), .B(n39660), .Z(n39656) );
  ANDN U39936 ( .B(B[136]), .A(n66), .Z(n39440) );
  XNOR U39937 ( .A(n39448), .B(n39662), .Z(n39441) );
  XNOR U39938 ( .A(n39447), .B(n39445), .Z(n39662) );
  AND U39939 ( .A(n39663), .B(n39664), .Z(n39445) );
  NANDN U39940 ( .A(n39665), .B(n39666), .Z(n39664) );
  OR U39941 ( .A(n39667), .B(n39668), .Z(n39666) );
  NAND U39942 ( .A(n39668), .B(n39667), .Z(n39663) );
  ANDN U39943 ( .B(B[137]), .A(n67), .Z(n39447) );
  XNOR U39944 ( .A(n39455), .B(n39669), .Z(n39448) );
  XNOR U39945 ( .A(n39454), .B(n39452), .Z(n39669) );
  AND U39946 ( .A(n39670), .B(n39671), .Z(n39452) );
  NANDN U39947 ( .A(n39672), .B(n39673), .Z(n39671) );
  NANDN U39948 ( .A(n39674), .B(n39675), .Z(n39673) );
  NANDN U39949 ( .A(n39675), .B(n39674), .Z(n39670) );
  ANDN U39950 ( .B(B[138]), .A(n68), .Z(n39454) );
  XNOR U39951 ( .A(n39462), .B(n39676), .Z(n39455) );
  XNOR U39952 ( .A(n39461), .B(n39459), .Z(n39676) );
  AND U39953 ( .A(n39677), .B(n39678), .Z(n39459) );
  NANDN U39954 ( .A(n39679), .B(n39680), .Z(n39678) );
  OR U39955 ( .A(n39681), .B(n39682), .Z(n39680) );
  NAND U39956 ( .A(n39682), .B(n39681), .Z(n39677) );
  ANDN U39957 ( .B(B[139]), .A(n69), .Z(n39461) );
  XNOR U39958 ( .A(n39469), .B(n39683), .Z(n39462) );
  XNOR U39959 ( .A(n39468), .B(n39466), .Z(n39683) );
  AND U39960 ( .A(n39684), .B(n39685), .Z(n39466) );
  NANDN U39961 ( .A(n39686), .B(n39687), .Z(n39685) );
  NANDN U39962 ( .A(n39688), .B(n39689), .Z(n39687) );
  NANDN U39963 ( .A(n39689), .B(n39688), .Z(n39684) );
  ANDN U39964 ( .B(B[140]), .A(n70), .Z(n39468) );
  XNOR U39965 ( .A(n39476), .B(n39690), .Z(n39469) );
  XNOR U39966 ( .A(n39475), .B(n39473), .Z(n39690) );
  AND U39967 ( .A(n39691), .B(n39692), .Z(n39473) );
  NANDN U39968 ( .A(n39693), .B(n39694), .Z(n39692) );
  OR U39969 ( .A(n39695), .B(n39696), .Z(n39694) );
  NAND U39970 ( .A(n39696), .B(n39695), .Z(n39691) );
  ANDN U39971 ( .B(B[141]), .A(n71), .Z(n39475) );
  XNOR U39972 ( .A(n39483), .B(n39697), .Z(n39476) );
  XNOR U39973 ( .A(n39482), .B(n39480), .Z(n39697) );
  AND U39974 ( .A(n39698), .B(n39699), .Z(n39480) );
  NANDN U39975 ( .A(n39700), .B(n39701), .Z(n39699) );
  NANDN U39976 ( .A(n39702), .B(n39703), .Z(n39701) );
  NANDN U39977 ( .A(n39703), .B(n39702), .Z(n39698) );
  ANDN U39978 ( .B(B[142]), .A(n72), .Z(n39482) );
  XNOR U39979 ( .A(n39490), .B(n39704), .Z(n39483) );
  XNOR U39980 ( .A(n39489), .B(n39487), .Z(n39704) );
  AND U39981 ( .A(n39705), .B(n39706), .Z(n39487) );
  NANDN U39982 ( .A(n39707), .B(n39708), .Z(n39706) );
  OR U39983 ( .A(n39709), .B(n39710), .Z(n39708) );
  NAND U39984 ( .A(n39710), .B(n39709), .Z(n39705) );
  ANDN U39985 ( .B(B[143]), .A(n73), .Z(n39489) );
  XNOR U39986 ( .A(n39497), .B(n39711), .Z(n39490) );
  XNOR U39987 ( .A(n39496), .B(n39494), .Z(n39711) );
  AND U39988 ( .A(n39712), .B(n39713), .Z(n39494) );
  NANDN U39989 ( .A(n39714), .B(n39715), .Z(n39713) );
  NANDN U39990 ( .A(n39716), .B(n39717), .Z(n39715) );
  NANDN U39991 ( .A(n39717), .B(n39716), .Z(n39712) );
  ANDN U39992 ( .B(B[144]), .A(n74), .Z(n39496) );
  XNOR U39993 ( .A(n39504), .B(n39718), .Z(n39497) );
  XNOR U39994 ( .A(n39503), .B(n39501), .Z(n39718) );
  AND U39995 ( .A(n39719), .B(n39720), .Z(n39501) );
  NANDN U39996 ( .A(n39721), .B(n39722), .Z(n39720) );
  OR U39997 ( .A(n39723), .B(n39724), .Z(n39722) );
  NAND U39998 ( .A(n39724), .B(n39723), .Z(n39719) );
  ANDN U39999 ( .B(B[145]), .A(n75), .Z(n39503) );
  XNOR U40000 ( .A(n39511), .B(n39725), .Z(n39504) );
  XNOR U40001 ( .A(n39510), .B(n39508), .Z(n39725) );
  AND U40002 ( .A(n39726), .B(n39727), .Z(n39508) );
  NANDN U40003 ( .A(n39728), .B(n39729), .Z(n39727) );
  NANDN U40004 ( .A(n39730), .B(n39731), .Z(n39729) );
  NANDN U40005 ( .A(n39731), .B(n39730), .Z(n39726) );
  ANDN U40006 ( .B(B[146]), .A(n76), .Z(n39510) );
  XNOR U40007 ( .A(n39518), .B(n39732), .Z(n39511) );
  XNOR U40008 ( .A(n39517), .B(n39515), .Z(n39732) );
  AND U40009 ( .A(n39733), .B(n39734), .Z(n39515) );
  NANDN U40010 ( .A(n39735), .B(n39736), .Z(n39734) );
  OR U40011 ( .A(n39737), .B(n39738), .Z(n39736) );
  NAND U40012 ( .A(n39738), .B(n39737), .Z(n39733) );
  ANDN U40013 ( .B(B[147]), .A(n77), .Z(n39517) );
  XNOR U40014 ( .A(n39525), .B(n39739), .Z(n39518) );
  XNOR U40015 ( .A(n39524), .B(n39522), .Z(n39739) );
  AND U40016 ( .A(n39740), .B(n39741), .Z(n39522) );
  NANDN U40017 ( .A(n39742), .B(n39743), .Z(n39741) );
  NANDN U40018 ( .A(n39744), .B(n39745), .Z(n39743) );
  NANDN U40019 ( .A(n39745), .B(n39744), .Z(n39740) );
  ANDN U40020 ( .B(B[148]), .A(n78), .Z(n39524) );
  XNOR U40021 ( .A(n39532), .B(n39746), .Z(n39525) );
  XNOR U40022 ( .A(n39531), .B(n39529), .Z(n39746) );
  AND U40023 ( .A(n39747), .B(n39748), .Z(n39529) );
  NANDN U40024 ( .A(n39749), .B(n39750), .Z(n39748) );
  OR U40025 ( .A(n39751), .B(n39752), .Z(n39750) );
  NAND U40026 ( .A(n39752), .B(n39751), .Z(n39747) );
  ANDN U40027 ( .B(B[149]), .A(n79), .Z(n39531) );
  XNOR U40028 ( .A(n39539), .B(n39753), .Z(n39532) );
  XNOR U40029 ( .A(n39538), .B(n39536), .Z(n39753) );
  AND U40030 ( .A(n39754), .B(n39755), .Z(n39536) );
  NANDN U40031 ( .A(n39756), .B(n39757), .Z(n39755) );
  NANDN U40032 ( .A(n39758), .B(n39759), .Z(n39757) );
  NANDN U40033 ( .A(n39759), .B(n39758), .Z(n39754) );
  ANDN U40034 ( .B(B[150]), .A(n80), .Z(n39538) );
  XNOR U40035 ( .A(n39546), .B(n39760), .Z(n39539) );
  XNOR U40036 ( .A(n39545), .B(n39543), .Z(n39760) );
  AND U40037 ( .A(n39761), .B(n39762), .Z(n39543) );
  NANDN U40038 ( .A(n39763), .B(n39764), .Z(n39762) );
  OR U40039 ( .A(n39765), .B(n39766), .Z(n39764) );
  NAND U40040 ( .A(n39766), .B(n39765), .Z(n39761) );
  ANDN U40041 ( .B(B[151]), .A(n81), .Z(n39545) );
  XNOR U40042 ( .A(n39553), .B(n39767), .Z(n39546) );
  XNOR U40043 ( .A(n39552), .B(n39550), .Z(n39767) );
  AND U40044 ( .A(n39768), .B(n39769), .Z(n39550) );
  NANDN U40045 ( .A(n39770), .B(n39771), .Z(n39769) );
  NAND U40046 ( .A(n39772), .B(n39773), .Z(n39771) );
  ANDN U40047 ( .B(B[152]), .A(n82), .Z(n39552) );
  XOR U40048 ( .A(n39559), .B(n39774), .Z(n39553) );
  XNOR U40049 ( .A(n39557), .B(n39560), .Z(n39774) );
  NAND U40050 ( .A(A[2]), .B(B[153]), .Z(n39560) );
  NANDN U40051 ( .A(n39775), .B(n39776), .Z(n39557) );
  AND U40052 ( .A(A[0]), .B(B[154]), .Z(n39776) );
  XNOR U40053 ( .A(n39562), .B(n39777), .Z(n39559) );
  NAND U40054 ( .A(A[0]), .B(B[155]), .Z(n39777) );
  NAND U40055 ( .A(B[154]), .B(A[1]), .Z(n39562) );
  NAND U40056 ( .A(n39778), .B(n39779), .Z(n486) );
  NANDN U40057 ( .A(n39780), .B(n39781), .Z(n39779) );
  OR U40058 ( .A(n39782), .B(n39783), .Z(n39781) );
  NAND U40059 ( .A(n39783), .B(n39782), .Z(n39778) );
  XOR U40060 ( .A(n488), .B(n487), .Z(\A1[152] ) );
  XOR U40061 ( .A(n39783), .B(n39784), .Z(n487) );
  XNOR U40062 ( .A(n39782), .B(n39780), .Z(n39784) );
  AND U40063 ( .A(n39785), .B(n39786), .Z(n39780) );
  NANDN U40064 ( .A(n39787), .B(n39788), .Z(n39786) );
  NANDN U40065 ( .A(n39789), .B(n39790), .Z(n39788) );
  NANDN U40066 ( .A(n39790), .B(n39789), .Z(n39785) );
  ANDN U40067 ( .B(B[123]), .A(n54), .Z(n39782) );
  XNOR U40068 ( .A(n39577), .B(n39791), .Z(n39783) );
  XNOR U40069 ( .A(n39576), .B(n39574), .Z(n39791) );
  AND U40070 ( .A(n39792), .B(n39793), .Z(n39574) );
  NANDN U40071 ( .A(n39794), .B(n39795), .Z(n39793) );
  OR U40072 ( .A(n39796), .B(n39797), .Z(n39795) );
  NAND U40073 ( .A(n39797), .B(n39796), .Z(n39792) );
  ANDN U40074 ( .B(B[124]), .A(n55), .Z(n39576) );
  XNOR U40075 ( .A(n39584), .B(n39798), .Z(n39577) );
  XNOR U40076 ( .A(n39583), .B(n39581), .Z(n39798) );
  AND U40077 ( .A(n39799), .B(n39800), .Z(n39581) );
  NANDN U40078 ( .A(n39801), .B(n39802), .Z(n39800) );
  NANDN U40079 ( .A(n39803), .B(n39804), .Z(n39802) );
  NANDN U40080 ( .A(n39804), .B(n39803), .Z(n39799) );
  ANDN U40081 ( .B(B[125]), .A(n56), .Z(n39583) );
  XNOR U40082 ( .A(n39591), .B(n39805), .Z(n39584) );
  XNOR U40083 ( .A(n39590), .B(n39588), .Z(n39805) );
  AND U40084 ( .A(n39806), .B(n39807), .Z(n39588) );
  NANDN U40085 ( .A(n39808), .B(n39809), .Z(n39807) );
  OR U40086 ( .A(n39810), .B(n39811), .Z(n39809) );
  NAND U40087 ( .A(n39811), .B(n39810), .Z(n39806) );
  ANDN U40088 ( .B(B[126]), .A(n57), .Z(n39590) );
  XNOR U40089 ( .A(n39598), .B(n39812), .Z(n39591) );
  XNOR U40090 ( .A(n39597), .B(n39595), .Z(n39812) );
  AND U40091 ( .A(n39813), .B(n39814), .Z(n39595) );
  NANDN U40092 ( .A(n39815), .B(n39816), .Z(n39814) );
  NANDN U40093 ( .A(n39817), .B(n39818), .Z(n39816) );
  NANDN U40094 ( .A(n39818), .B(n39817), .Z(n39813) );
  ANDN U40095 ( .B(B[127]), .A(n58), .Z(n39597) );
  XNOR U40096 ( .A(n39605), .B(n39819), .Z(n39598) );
  XNOR U40097 ( .A(n39604), .B(n39602), .Z(n39819) );
  AND U40098 ( .A(n39820), .B(n39821), .Z(n39602) );
  NANDN U40099 ( .A(n39822), .B(n39823), .Z(n39821) );
  OR U40100 ( .A(n39824), .B(n39825), .Z(n39823) );
  NAND U40101 ( .A(n39825), .B(n39824), .Z(n39820) );
  ANDN U40102 ( .B(B[128]), .A(n59), .Z(n39604) );
  XNOR U40103 ( .A(n39612), .B(n39826), .Z(n39605) );
  XNOR U40104 ( .A(n39611), .B(n39609), .Z(n39826) );
  AND U40105 ( .A(n39827), .B(n39828), .Z(n39609) );
  NANDN U40106 ( .A(n39829), .B(n39830), .Z(n39828) );
  NANDN U40107 ( .A(n39831), .B(n39832), .Z(n39830) );
  NANDN U40108 ( .A(n39832), .B(n39831), .Z(n39827) );
  ANDN U40109 ( .B(B[129]), .A(n60), .Z(n39611) );
  XNOR U40110 ( .A(n39619), .B(n39833), .Z(n39612) );
  XNOR U40111 ( .A(n39618), .B(n39616), .Z(n39833) );
  AND U40112 ( .A(n39834), .B(n39835), .Z(n39616) );
  NANDN U40113 ( .A(n39836), .B(n39837), .Z(n39835) );
  OR U40114 ( .A(n39838), .B(n39839), .Z(n39837) );
  NAND U40115 ( .A(n39839), .B(n39838), .Z(n39834) );
  ANDN U40116 ( .B(B[130]), .A(n61), .Z(n39618) );
  XNOR U40117 ( .A(n39626), .B(n39840), .Z(n39619) );
  XNOR U40118 ( .A(n39625), .B(n39623), .Z(n39840) );
  AND U40119 ( .A(n39841), .B(n39842), .Z(n39623) );
  NANDN U40120 ( .A(n39843), .B(n39844), .Z(n39842) );
  NANDN U40121 ( .A(n39845), .B(n39846), .Z(n39844) );
  NANDN U40122 ( .A(n39846), .B(n39845), .Z(n39841) );
  ANDN U40123 ( .B(B[131]), .A(n62), .Z(n39625) );
  XNOR U40124 ( .A(n39633), .B(n39847), .Z(n39626) );
  XNOR U40125 ( .A(n39632), .B(n39630), .Z(n39847) );
  AND U40126 ( .A(n39848), .B(n39849), .Z(n39630) );
  NANDN U40127 ( .A(n39850), .B(n39851), .Z(n39849) );
  OR U40128 ( .A(n39852), .B(n39853), .Z(n39851) );
  NAND U40129 ( .A(n39853), .B(n39852), .Z(n39848) );
  ANDN U40130 ( .B(B[132]), .A(n63), .Z(n39632) );
  XNOR U40131 ( .A(n39640), .B(n39854), .Z(n39633) );
  XNOR U40132 ( .A(n39639), .B(n39637), .Z(n39854) );
  AND U40133 ( .A(n39855), .B(n39856), .Z(n39637) );
  NANDN U40134 ( .A(n39857), .B(n39858), .Z(n39856) );
  NANDN U40135 ( .A(n39859), .B(n39860), .Z(n39858) );
  NANDN U40136 ( .A(n39860), .B(n39859), .Z(n39855) );
  ANDN U40137 ( .B(B[133]), .A(n64), .Z(n39639) );
  XNOR U40138 ( .A(n39647), .B(n39861), .Z(n39640) );
  XNOR U40139 ( .A(n39646), .B(n39644), .Z(n39861) );
  AND U40140 ( .A(n39862), .B(n39863), .Z(n39644) );
  NANDN U40141 ( .A(n39864), .B(n39865), .Z(n39863) );
  OR U40142 ( .A(n39866), .B(n39867), .Z(n39865) );
  NAND U40143 ( .A(n39867), .B(n39866), .Z(n39862) );
  ANDN U40144 ( .B(B[134]), .A(n65), .Z(n39646) );
  XNOR U40145 ( .A(n39654), .B(n39868), .Z(n39647) );
  XNOR U40146 ( .A(n39653), .B(n39651), .Z(n39868) );
  AND U40147 ( .A(n39869), .B(n39870), .Z(n39651) );
  NANDN U40148 ( .A(n39871), .B(n39872), .Z(n39870) );
  NANDN U40149 ( .A(n39873), .B(n39874), .Z(n39872) );
  NANDN U40150 ( .A(n39874), .B(n39873), .Z(n39869) );
  ANDN U40151 ( .B(B[135]), .A(n66), .Z(n39653) );
  XNOR U40152 ( .A(n39661), .B(n39875), .Z(n39654) );
  XNOR U40153 ( .A(n39660), .B(n39658), .Z(n39875) );
  AND U40154 ( .A(n39876), .B(n39877), .Z(n39658) );
  NANDN U40155 ( .A(n39878), .B(n39879), .Z(n39877) );
  OR U40156 ( .A(n39880), .B(n39881), .Z(n39879) );
  NAND U40157 ( .A(n39881), .B(n39880), .Z(n39876) );
  ANDN U40158 ( .B(B[136]), .A(n67), .Z(n39660) );
  XNOR U40159 ( .A(n39668), .B(n39882), .Z(n39661) );
  XNOR U40160 ( .A(n39667), .B(n39665), .Z(n39882) );
  AND U40161 ( .A(n39883), .B(n39884), .Z(n39665) );
  NANDN U40162 ( .A(n39885), .B(n39886), .Z(n39884) );
  NANDN U40163 ( .A(n39887), .B(n39888), .Z(n39886) );
  NANDN U40164 ( .A(n39888), .B(n39887), .Z(n39883) );
  ANDN U40165 ( .B(B[137]), .A(n68), .Z(n39667) );
  XNOR U40166 ( .A(n39675), .B(n39889), .Z(n39668) );
  XNOR U40167 ( .A(n39674), .B(n39672), .Z(n39889) );
  AND U40168 ( .A(n39890), .B(n39891), .Z(n39672) );
  NANDN U40169 ( .A(n39892), .B(n39893), .Z(n39891) );
  OR U40170 ( .A(n39894), .B(n39895), .Z(n39893) );
  NAND U40171 ( .A(n39895), .B(n39894), .Z(n39890) );
  ANDN U40172 ( .B(B[138]), .A(n69), .Z(n39674) );
  XNOR U40173 ( .A(n39682), .B(n39896), .Z(n39675) );
  XNOR U40174 ( .A(n39681), .B(n39679), .Z(n39896) );
  AND U40175 ( .A(n39897), .B(n39898), .Z(n39679) );
  NANDN U40176 ( .A(n39899), .B(n39900), .Z(n39898) );
  NANDN U40177 ( .A(n39901), .B(n39902), .Z(n39900) );
  NANDN U40178 ( .A(n39902), .B(n39901), .Z(n39897) );
  ANDN U40179 ( .B(B[139]), .A(n70), .Z(n39681) );
  XNOR U40180 ( .A(n39689), .B(n39903), .Z(n39682) );
  XNOR U40181 ( .A(n39688), .B(n39686), .Z(n39903) );
  AND U40182 ( .A(n39904), .B(n39905), .Z(n39686) );
  NANDN U40183 ( .A(n39906), .B(n39907), .Z(n39905) );
  OR U40184 ( .A(n39908), .B(n39909), .Z(n39907) );
  NAND U40185 ( .A(n39909), .B(n39908), .Z(n39904) );
  ANDN U40186 ( .B(B[140]), .A(n71), .Z(n39688) );
  XNOR U40187 ( .A(n39696), .B(n39910), .Z(n39689) );
  XNOR U40188 ( .A(n39695), .B(n39693), .Z(n39910) );
  AND U40189 ( .A(n39911), .B(n39912), .Z(n39693) );
  NANDN U40190 ( .A(n39913), .B(n39914), .Z(n39912) );
  NANDN U40191 ( .A(n39915), .B(n39916), .Z(n39914) );
  NANDN U40192 ( .A(n39916), .B(n39915), .Z(n39911) );
  ANDN U40193 ( .B(B[141]), .A(n72), .Z(n39695) );
  XNOR U40194 ( .A(n39703), .B(n39917), .Z(n39696) );
  XNOR U40195 ( .A(n39702), .B(n39700), .Z(n39917) );
  AND U40196 ( .A(n39918), .B(n39919), .Z(n39700) );
  NANDN U40197 ( .A(n39920), .B(n39921), .Z(n39919) );
  OR U40198 ( .A(n39922), .B(n39923), .Z(n39921) );
  NAND U40199 ( .A(n39923), .B(n39922), .Z(n39918) );
  ANDN U40200 ( .B(B[142]), .A(n73), .Z(n39702) );
  XNOR U40201 ( .A(n39710), .B(n39924), .Z(n39703) );
  XNOR U40202 ( .A(n39709), .B(n39707), .Z(n39924) );
  AND U40203 ( .A(n39925), .B(n39926), .Z(n39707) );
  NANDN U40204 ( .A(n39927), .B(n39928), .Z(n39926) );
  NANDN U40205 ( .A(n39929), .B(n39930), .Z(n39928) );
  NANDN U40206 ( .A(n39930), .B(n39929), .Z(n39925) );
  ANDN U40207 ( .B(B[143]), .A(n74), .Z(n39709) );
  XNOR U40208 ( .A(n39717), .B(n39931), .Z(n39710) );
  XNOR U40209 ( .A(n39716), .B(n39714), .Z(n39931) );
  AND U40210 ( .A(n39932), .B(n39933), .Z(n39714) );
  NANDN U40211 ( .A(n39934), .B(n39935), .Z(n39933) );
  OR U40212 ( .A(n39936), .B(n39937), .Z(n39935) );
  NAND U40213 ( .A(n39937), .B(n39936), .Z(n39932) );
  ANDN U40214 ( .B(B[144]), .A(n75), .Z(n39716) );
  XNOR U40215 ( .A(n39724), .B(n39938), .Z(n39717) );
  XNOR U40216 ( .A(n39723), .B(n39721), .Z(n39938) );
  AND U40217 ( .A(n39939), .B(n39940), .Z(n39721) );
  NANDN U40218 ( .A(n39941), .B(n39942), .Z(n39940) );
  NANDN U40219 ( .A(n39943), .B(n39944), .Z(n39942) );
  NANDN U40220 ( .A(n39944), .B(n39943), .Z(n39939) );
  ANDN U40221 ( .B(B[145]), .A(n76), .Z(n39723) );
  XNOR U40222 ( .A(n39731), .B(n39945), .Z(n39724) );
  XNOR U40223 ( .A(n39730), .B(n39728), .Z(n39945) );
  AND U40224 ( .A(n39946), .B(n39947), .Z(n39728) );
  NANDN U40225 ( .A(n39948), .B(n39949), .Z(n39947) );
  OR U40226 ( .A(n39950), .B(n39951), .Z(n39949) );
  NAND U40227 ( .A(n39951), .B(n39950), .Z(n39946) );
  ANDN U40228 ( .B(B[146]), .A(n77), .Z(n39730) );
  XNOR U40229 ( .A(n39738), .B(n39952), .Z(n39731) );
  XNOR U40230 ( .A(n39737), .B(n39735), .Z(n39952) );
  AND U40231 ( .A(n39953), .B(n39954), .Z(n39735) );
  NANDN U40232 ( .A(n39955), .B(n39956), .Z(n39954) );
  NANDN U40233 ( .A(n39957), .B(n39958), .Z(n39956) );
  NANDN U40234 ( .A(n39958), .B(n39957), .Z(n39953) );
  ANDN U40235 ( .B(B[147]), .A(n78), .Z(n39737) );
  XNOR U40236 ( .A(n39745), .B(n39959), .Z(n39738) );
  XNOR U40237 ( .A(n39744), .B(n39742), .Z(n39959) );
  AND U40238 ( .A(n39960), .B(n39961), .Z(n39742) );
  NANDN U40239 ( .A(n39962), .B(n39963), .Z(n39961) );
  OR U40240 ( .A(n39964), .B(n39965), .Z(n39963) );
  NAND U40241 ( .A(n39965), .B(n39964), .Z(n39960) );
  ANDN U40242 ( .B(B[148]), .A(n79), .Z(n39744) );
  XNOR U40243 ( .A(n39752), .B(n39966), .Z(n39745) );
  XNOR U40244 ( .A(n39751), .B(n39749), .Z(n39966) );
  AND U40245 ( .A(n39967), .B(n39968), .Z(n39749) );
  NANDN U40246 ( .A(n39969), .B(n39970), .Z(n39968) );
  NANDN U40247 ( .A(n39971), .B(n39972), .Z(n39970) );
  NANDN U40248 ( .A(n39972), .B(n39971), .Z(n39967) );
  ANDN U40249 ( .B(B[149]), .A(n80), .Z(n39751) );
  XNOR U40250 ( .A(n39759), .B(n39973), .Z(n39752) );
  XNOR U40251 ( .A(n39758), .B(n39756), .Z(n39973) );
  AND U40252 ( .A(n39974), .B(n39975), .Z(n39756) );
  NANDN U40253 ( .A(n39976), .B(n39977), .Z(n39975) );
  OR U40254 ( .A(n39978), .B(n39979), .Z(n39977) );
  NAND U40255 ( .A(n39979), .B(n39978), .Z(n39974) );
  ANDN U40256 ( .B(B[150]), .A(n81), .Z(n39758) );
  XNOR U40257 ( .A(n39766), .B(n39980), .Z(n39759) );
  XNOR U40258 ( .A(n39765), .B(n39763), .Z(n39980) );
  AND U40259 ( .A(n39981), .B(n39982), .Z(n39763) );
  NANDN U40260 ( .A(n39983), .B(n39984), .Z(n39982) );
  NAND U40261 ( .A(n39985), .B(n39986), .Z(n39984) );
  ANDN U40262 ( .B(B[151]), .A(n82), .Z(n39765) );
  XOR U40263 ( .A(n39772), .B(n39987), .Z(n39766) );
  XNOR U40264 ( .A(n39770), .B(n39773), .Z(n39987) );
  NAND U40265 ( .A(A[2]), .B(B[152]), .Z(n39773) );
  NANDN U40266 ( .A(n39988), .B(n39989), .Z(n39770) );
  AND U40267 ( .A(A[0]), .B(B[153]), .Z(n39989) );
  XNOR U40268 ( .A(n39775), .B(n39990), .Z(n39772) );
  NAND U40269 ( .A(A[0]), .B(B[154]), .Z(n39990) );
  NAND U40270 ( .A(B[153]), .B(A[1]), .Z(n39775) );
  NAND U40271 ( .A(n39991), .B(n39992), .Z(n488) );
  NANDN U40272 ( .A(n39993), .B(n39994), .Z(n39992) );
  OR U40273 ( .A(n39995), .B(n39996), .Z(n39994) );
  NAND U40274 ( .A(n39996), .B(n39995), .Z(n39991) );
  XOR U40275 ( .A(n490), .B(n489), .Z(\A1[151] ) );
  XOR U40276 ( .A(n39996), .B(n39997), .Z(n489) );
  XNOR U40277 ( .A(n39995), .B(n39993), .Z(n39997) );
  AND U40278 ( .A(n39998), .B(n39999), .Z(n39993) );
  NANDN U40279 ( .A(n40000), .B(n40001), .Z(n39999) );
  NANDN U40280 ( .A(n40002), .B(n40003), .Z(n40001) );
  NANDN U40281 ( .A(n40003), .B(n40002), .Z(n39998) );
  ANDN U40282 ( .B(B[122]), .A(n54), .Z(n39995) );
  XNOR U40283 ( .A(n39790), .B(n40004), .Z(n39996) );
  XNOR U40284 ( .A(n39789), .B(n39787), .Z(n40004) );
  AND U40285 ( .A(n40005), .B(n40006), .Z(n39787) );
  NANDN U40286 ( .A(n40007), .B(n40008), .Z(n40006) );
  OR U40287 ( .A(n40009), .B(n40010), .Z(n40008) );
  NAND U40288 ( .A(n40010), .B(n40009), .Z(n40005) );
  ANDN U40289 ( .B(B[123]), .A(n55), .Z(n39789) );
  XNOR U40290 ( .A(n39797), .B(n40011), .Z(n39790) );
  XNOR U40291 ( .A(n39796), .B(n39794), .Z(n40011) );
  AND U40292 ( .A(n40012), .B(n40013), .Z(n39794) );
  NANDN U40293 ( .A(n40014), .B(n40015), .Z(n40013) );
  NANDN U40294 ( .A(n40016), .B(n40017), .Z(n40015) );
  NANDN U40295 ( .A(n40017), .B(n40016), .Z(n40012) );
  ANDN U40296 ( .B(B[124]), .A(n56), .Z(n39796) );
  XNOR U40297 ( .A(n39804), .B(n40018), .Z(n39797) );
  XNOR U40298 ( .A(n39803), .B(n39801), .Z(n40018) );
  AND U40299 ( .A(n40019), .B(n40020), .Z(n39801) );
  NANDN U40300 ( .A(n40021), .B(n40022), .Z(n40020) );
  OR U40301 ( .A(n40023), .B(n40024), .Z(n40022) );
  NAND U40302 ( .A(n40024), .B(n40023), .Z(n40019) );
  ANDN U40303 ( .B(B[125]), .A(n57), .Z(n39803) );
  XNOR U40304 ( .A(n39811), .B(n40025), .Z(n39804) );
  XNOR U40305 ( .A(n39810), .B(n39808), .Z(n40025) );
  AND U40306 ( .A(n40026), .B(n40027), .Z(n39808) );
  NANDN U40307 ( .A(n40028), .B(n40029), .Z(n40027) );
  NANDN U40308 ( .A(n40030), .B(n40031), .Z(n40029) );
  NANDN U40309 ( .A(n40031), .B(n40030), .Z(n40026) );
  ANDN U40310 ( .B(B[126]), .A(n58), .Z(n39810) );
  XNOR U40311 ( .A(n39818), .B(n40032), .Z(n39811) );
  XNOR U40312 ( .A(n39817), .B(n39815), .Z(n40032) );
  AND U40313 ( .A(n40033), .B(n40034), .Z(n39815) );
  NANDN U40314 ( .A(n40035), .B(n40036), .Z(n40034) );
  OR U40315 ( .A(n40037), .B(n40038), .Z(n40036) );
  NAND U40316 ( .A(n40038), .B(n40037), .Z(n40033) );
  ANDN U40317 ( .B(B[127]), .A(n59), .Z(n39817) );
  XNOR U40318 ( .A(n39825), .B(n40039), .Z(n39818) );
  XNOR U40319 ( .A(n39824), .B(n39822), .Z(n40039) );
  AND U40320 ( .A(n40040), .B(n40041), .Z(n39822) );
  NANDN U40321 ( .A(n40042), .B(n40043), .Z(n40041) );
  NANDN U40322 ( .A(n40044), .B(n40045), .Z(n40043) );
  NANDN U40323 ( .A(n40045), .B(n40044), .Z(n40040) );
  ANDN U40324 ( .B(B[128]), .A(n60), .Z(n39824) );
  XNOR U40325 ( .A(n39832), .B(n40046), .Z(n39825) );
  XNOR U40326 ( .A(n39831), .B(n39829), .Z(n40046) );
  AND U40327 ( .A(n40047), .B(n40048), .Z(n39829) );
  NANDN U40328 ( .A(n40049), .B(n40050), .Z(n40048) );
  OR U40329 ( .A(n40051), .B(n40052), .Z(n40050) );
  NAND U40330 ( .A(n40052), .B(n40051), .Z(n40047) );
  ANDN U40331 ( .B(B[129]), .A(n61), .Z(n39831) );
  XNOR U40332 ( .A(n39839), .B(n40053), .Z(n39832) );
  XNOR U40333 ( .A(n39838), .B(n39836), .Z(n40053) );
  AND U40334 ( .A(n40054), .B(n40055), .Z(n39836) );
  NANDN U40335 ( .A(n40056), .B(n40057), .Z(n40055) );
  NANDN U40336 ( .A(n40058), .B(n40059), .Z(n40057) );
  NANDN U40337 ( .A(n40059), .B(n40058), .Z(n40054) );
  ANDN U40338 ( .B(B[130]), .A(n62), .Z(n39838) );
  XNOR U40339 ( .A(n39846), .B(n40060), .Z(n39839) );
  XNOR U40340 ( .A(n39845), .B(n39843), .Z(n40060) );
  AND U40341 ( .A(n40061), .B(n40062), .Z(n39843) );
  NANDN U40342 ( .A(n40063), .B(n40064), .Z(n40062) );
  OR U40343 ( .A(n40065), .B(n40066), .Z(n40064) );
  NAND U40344 ( .A(n40066), .B(n40065), .Z(n40061) );
  ANDN U40345 ( .B(B[131]), .A(n63), .Z(n39845) );
  XNOR U40346 ( .A(n39853), .B(n40067), .Z(n39846) );
  XNOR U40347 ( .A(n39852), .B(n39850), .Z(n40067) );
  AND U40348 ( .A(n40068), .B(n40069), .Z(n39850) );
  NANDN U40349 ( .A(n40070), .B(n40071), .Z(n40069) );
  NANDN U40350 ( .A(n40072), .B(n40073), .Z(n40071) );
  NANDN U40351 ( .A(n40073), .B(n40072), .Z(n40068) );
  ANDN U40352 ( .B(B[132]), .A(n64), .Z(n39852) );
  XNOR U40353 ( .A(n39860), .B(n40074), .Z(n39853) );
  XNOR U40354 ( .A(n39859), .B(n39857), .Z(n40074) );
  AND U40355 ( .A(n40075), .B(n40076), .Z(n39857) );
  NANDN U40356 ( .A(n40077), .B(n40078), .Z(n40076) );
  OR U40357 ( .A(n40079), .B(n40080), .Z(n40078) );
  NAND U40358 ( .A(n40080), .B(n40079), .Z(n40075) );
  ANDN U40359 ( .B(B[133]), .A(n65), .Z(n39859) );
  XNOR U40360 ( .A(n39867), .B(n40081), .Z(n39860) );
  XNOR U40361 ( .A(n39866), .B(n39864), .Z(n40081) );
  AND U40362 ( .A(n40082), .B(n40083), .Z(n39864) );
  NANDN U40363 ( .A(n40084), .B(n40085), .Z(n40083) );
  NANDN U40364 ( .A(n40086), .B(n40087), .Z(n40085) );
  NANDN U40365 ( .A(n40087), .B(n40086), .Z(n40082) );
  ANDN U40366 ( .B(B[134]), .A(n66), .Z(n39866) );
  XNOR U40367 ( .A(n39874), .B(n40088), .Z(n39867) );
  XNOR U40368 ( .A(n39873), .B(n39871), .Z(n40088) );
  AND U40369 ( .A(n40089), .B(n40090), .Z(n39871) );
  NANDN U40370 ( .A(n40091), .B(n40092), .Z(n40090) );
  OR U40371 ( .A(n40093), .B(n40094), .Z(n40092) );
  NAND U40372 ( .A(n40094), .B(n40093), .Z(n40089) );
  ANDN U40373 ( .B(B[135]), .A(n67), .Z(n39873) );
  XNOR U40374 ( .A(n39881), .B(n40095), .Z(n39874) );
  XNOR U40375 ( .A(n39880), .B(n39878), .Z(n40095) );
  AND U40376 ( .A(n40096), .B(n40097), .Z(n39878) );
  NANDN U40377 ( .A(n40098), .B(n40099), .Z(n40097) );
  NANDN U40378 ( .A(n40100), .B(n40101), .Z(n40099) );
  NANDN U40379 ( .A(n40101), .B(n40100), .Z(n40096) );
  ANDN U40380 ( .B(B[136]), .A(n68), .Z(n39880) );
  XNOR U40381 ( .A(n39888), .B(n40102), .Z(n39881) );
  XNOR U40382 ( .A(n39887), .B(n39885), .Z(n40102) );
  AND U40383 ( .A(n40103), .B(n40104), .Z(n39885) );
  NANDN U40384 ( .A(n40105), .B(n40106), .Z(n40104) );
  OR U40385 ( .A(n40107), .B(n40108), .Z(n40106) );
  NAND U40386 ( .A(n40108), .B(n40107), .Z(n40103) );
  ANDN U40387 ( .B(B[137]), .A(n69), .Z(n39887) );
  XNOR U40388 ( .A(n39895), .B(n40109), .Z(n39888) );
  XNOR U40389 ( .A(n39894), .B(n39892), .Z(n40109) );
  AND U40390 ( .A(n40110), .B(n40111), .Z(n39892) );
  NANDN U40391 ( .A(n40112), .B(n40113), .Z(n40111) );
  NANDN U40392 ( .A(n40114), .B(n40115), .Z(n40113) );
  NANDN U40393 ( .A(n40115), .B(n40114), .Z(n40110) );
  ANDN U40394 ( .B(B[138]), .A(n70), .Z(n39894) );
  XNOR U40395 ( .A(n39902), .B(n40116), .Z(n39895) );
  XNOR U40396 ( .A(n39901), .B(n39899), .Z(n40116) );
  AND U40397 ( .A(n40117), .B(n40118), .Z(n39899) );
  NANDN U40398 ( .A(n40119), .B(n40120), .Z(n40118) );
  OR U40399 ( .A(n40121), .B(n40122), .Z(n40120) );
  NAND U40400 ( .A(n40122), .B(n40121), .Z(n40117) );
  ANDN U40401 ( .B(B[139]), .A(n71), .Z(n39901) );
  XNOR U40402 ( .A(n39909), .B(n40123), .Z(n39902) );
  XNOR U40403 ( .A(n39908), .B(n39906), .Z(n40123) );
  AND U40404 ( .A(n40124), .B(n40125), .Z(n39906) );
  NANDN U40405 ( .A(n40126), .B(n40127), .Z(n40125) );
  NANDN U40406 ( .A(n40128), .B(n40129), .Z(n40127) );
  NANDN U40407 ( .A(n40129), .B(n40128), .Z(n40124) );
  ANDN U40408 ( .B(B[140]), .A(n72), .Z(n39908) );
  XNOR U40409 ( .A(n39916), .B(n40130), .Z(n39909) );
  XNOR U40410 ( .A(n39915), .B(n39913), .Z(n40130) );
  AND U40411 ( .A(n40131), .B(n40132), .Z(n39913) );
  NANDN U40412 ( .A(n40133), .B(n40134), .Z(n40132) );
  OR U40413 ( .A(n40135), .B(n40136), .Z(n40134) );
  NAND U40414 ( .A(n40136), .B(n40135), .Z(n40131) );
  ANDN U40415 ( .B(B[141]), .A(n73), .Z(n39915) );
  XNOR U40416 ( .A(n39923), .B(n40137), .Z(n39916) );
  XNOR U40417 ( .A(n39922), .B(n39920), .Z(n40137) );
  AND U40418 ( .A(n40138), .B(n40139), .Z(n39920) );
  NANDN U40419 ( .A(n40140), .B(n40141), .Z(n40139) );
  NANDN U40420 ( .A(n40142), .B(n40143), .Z(n40141) );
  NANDN U40421 ( .A(n40143), .B(n40142), .Z(n40138) );
  ANDN U40422 ( .B(B[142]), .A(n74), .Z(n39922) );
  XNOR U40423 ( .A(n39930), .B(n40144), .Z(n39923) );
  XNOR U40424 ( .A(n39929), .B(n39927), .Z(n40144) );
  AND U40425 ( .A(n40145), .B(n40146), .Z(n39927) );
  NANDN U40426 ( .A(n40147), .B(n40148), .Z(n40146) );
  OR U40427 ( .A(n40149), .B(n40150), .Z(n40148) );
  NAND U40428 ( .A(n40150), .B(n40149), .Z(n40145) );
  ANDN U40429 ( .B(B[143]), .A(n75), .Z(n39929) );
  XNOR U40430 ( .A(n39937), .B(n40151), .Z(n39930) );
  XNOR U40431 ( .A(n39936), .B(n39934), .Z(n40151) );
  AND U40432 ( .A(n40152), .B(n40153), .Z(n39934) );
  NANDN U40433 ( .A(n40154), .B(n40155), .Z(n40153) );
  NANDN U40434 ( .A(n40156), .B(n40157), .Z(n40155) );
  NANDN U40435 ( .A(n40157), .B(n40156), .Z(n40152) );
  ANDN U40436 ( .B(B[144]), .A(n76), .Z(n39936) );
  XNOR U40437 ( .A(n39944), .B(n40158), .Z(n39937) );
  XNOR U40438 ( .A(n39943), .B(n39941), .Z(n40158) );
  AND U40439 ( .A(n40159), .B(n40160), .Z(n39941) );
  NANDN U40440 ( .A(n40161), .B(n40162), .Z(n40160) );
  OR U40441 ( .A(n40163), .B(n40164), .Z(n40162) );
  NAND U40442 ( .A(n40164), .B(n40163), .Z(n40159) );
  ANDN U40443 ( .B(B[145]), .A(n77), .Z(n39943) );
  XNOR U40444 ( .A(n39951), .B(n40165), .Z(n39944) );
  XNOR U40445 ( .A(n39950), .B(n39948), .Z(n40165) );
  AND U40446 ( .A(n40166), .B(n40167), .Z(n39948) );
  NANDN U40447 ( .A(n40168), .B(n40169), .Z(n40167) );
  NANDN U40448 ( .A(n40170), .B(n40171), .Z(n40169) );
  NANDN U40449 ( .A(n40171), .B(n40170), .Z(n40166) );
  ANDN U40450 ( .B(B[146]), .A(n78), .Z(n39950) );
  XNOR U40451 ( .A(n39958), .B(n40172), .Z(n39951) );
  XNOR U40452 ( .A(n39957), .B(n39955), .Z(n40172) );
  AND U40453 ( .A(n40173), .B(n40174), .Z(n39955) );
  NANDN U40454 ( .A(n40175), .B(n40176), .Z(n40174) );
  OR U40455 ( .A(n40177), .B(n40178), .Z(n40176) );
  NAND U40456 ( .A(n40178), .B(n40177), .Z(n40173) );
  ANDN U40457 ( .B(B[147]), .A(n79), .Z(n39957) );
  XNOR U40458 ( .A(n39965), .B(n40179), .Z(n39958) );
  XNOR U40459 ( .A(n39964), .B(n39962), .Z(n40179) );
  AND U40460 ( .A(n40180), .B(n40181), .Z(n39962) );
  NANDN U40461 ( .A(n40182), .B(n40183), .Z(n40181) );
  NANDN U40462 ( .A(n40184), .B(n40185), .Z(n40183) );
  NANDN U40463 ( .A(n40185), .B(n40184), .Z(n40180) );
  ANDN U40464 ( .B(B[148]), .A(n80), .Z(n39964) );
  XNOR U40465 ( .A(n39972), .B(n40186), .Z(n39965) );
  XNOR U40466 ( .A(n39971), .B(n39969), .Z(n40186) );
  AND U40467 ( .A(n40187), .B(n40188), .Z(n39969) );
  NANDN U40468 ( .A(n40189), .B(n40190), .Z(n40188) );
  OR U40469 ( .A(n40191), .B(n40192), .Z(n40190) );
  NAND U40470 ( .A(n40192), .B(n40191), .Z(n40187) );
  ANDN U40471 ( .B(B[149]), .A(n81), .Z(n39971) );
  XNOR U40472 ( .A(n39979), .B(n40193), .Z(n39972) );
  XNOR U40473 ( .A(n39978), .B(n39976), .Z(n40193) );
  AND U40474 ( .A(n40194), .B(n40195), .Z(n39976) );
  NANDN U40475 ( .A(n40196), .B(n40197), .Z(n40195) );
  NAND U40476 ( .A(n40198), .B(n40199), .Z(n40197) );
  ANDN U40477 ( .B(B[150]), .A(n82), .Z(n39978) );
  XOR U40478 ( .A(n39985), .B(n40200), .Z(n39979) );
  XNOR U40479 ( .A(n39983), .B(n39986), .Z(n40200) );
  NAND U40480 ( .A(A[2]), .B(B[151]), .Z(n39986) );
  NANDN U40481 ( .A(n40201), .B(n40202), .Z(n39983) );
  AND U40482 ( .A(A[0]), .B(B[152]), .Z(n40202) );
  XNOR U40483 ( .A(n39988), .B(n40203), .Z(n39985) );
  NAND U40484 ( .A(A[0]), .B(B[153]), .Z(n40203) );
  NAND U40485 ( .A(B[152]), .B(A[1]), .Z(n39988) );
  NAND U40486 ( .A(n40204), .B(n40205), .Z(n490) );
  NANDN U40487 ( .A(n40206), .B(n40207), .Z(n40205) );
  OR U40488 ( .A(n40208), .B(n40209), .Z(n40207) );
  NAND U40489 ( .A(n40209), .B(n40208), .Z(n40204) );
  XOR U40490 ( .A(n492), .B(n491), .Z(\A1[150] ) );
  XOR U40491 ( .A(n40209), .B(n40210), .Z(n491) );
  XNOR U40492 ( .A(n40208), .B(n40206), .Z(n40210) );
  AND U40493 ( .A(n40211), .B(n40212), .Z(n40206) );
  NANDN U40494 ( .A(n40213), .B(n40214), .Z(n40212) );
  NANDN U40495 ( .A(n40215), .B(n40216), .Z(n40214) );
  NANDN U40496 ( .A(n40216), .B(n40215), .Z(n40211) );
  ANDN U40497 ( .B(B[121]), .A(n54), .Z(n40208) );
  XNOR U40498 ( .A(n40003), .B(n40217), .Z(n40209) );
  XNOR U40499 ( .A(n40002), .B(n40000), .Z(n40217) );
  AND U40500 ( .A(n40218), .B(n40219), .Z(n40000) );
  NANDN U40501 ( .A(n40220), .B(n40221), .Z(n40219) );
  OR U40502 ( .A(n40222), .B(n40223), .Z(n40221) );
  NAND U40503 ( .A(n40223), .B(n40222), .Z(n40218) );
  ANDN U40504 ( .B(B[122]), .A(n55), .Z(n40002) );
  XNOR U40505 ( .A(n40010), .B(n40224), .Z(n40003) );
  XNOR U40506 ( .A(n40009), .B(n40007), .Z(n40224) );
  AND U40507 ( .A(n40225), .B(n40226), .Z(n40007) );
  NANDN U40508 ( .A(n40227), .B(n40228), .Z(n40226) );
  NANDN U40509 ( .A(n40229), .B(n40230), .Z(n40228) );
  NANDN U40510 ( .A(n40230), .B(n40229), .Z(n40225) );
  ANDN U40511 ( .B(B[123]), .A(n56), .Z(n40009) );
  XNOR U40512 ( .A(n40017), .B(n40231), .Z(n40010) );
  XNOR U40513 ( .A(n40016), .B(n40014), .Z(n40231) );
  AND U40514 ( .A(n40232), .B(n40233), .Z(n40014) );
  NANDN U40515 ( .A(n40234), .B(n40235), .Z(n40233) );
  OR U40516 ( .A(n40236), .B(n40237), .Z(n40235) );
  NAND U40517 ( .A(n40237), .B(n40236), .Z(n40232) );
  ANDN U40518 ( .B(B[124]), .A(n57), .Z(n40016) );
  XNOR U40519 ( .A(n40024), .B(n40238), .Z(n40017) );
  XNOR U40520 ( .A(n40023), .B(n40021), .Z(n40238) );
  AND U40521 ( .A(n40239), .B(n40240), .Z(n40021) );
  NANDN U40522 ( .A(n40241), .B(n40242), .Z(n40240) );
  NANDN U40523 ( .A(n40243), .B(n40244), .Z(n40242) );
  NANDN U40524 ( .A(n40244), .B(n40243), .Z(n40239) );
  ANDN U40525 ( .B(B[125]), .A(n58), .Z(n40023) );
  XNOR U40526 ( .A(n40031), .B(n40245), .Z(n40024) );
  XNOR U40527 ( .A(n40030), .B(n40028), .Z(n40245) );
  AND U40528 ( .A(n40246), .B(n40247), .Z(n40028) );
  NANDN U40529 ( .A(n40248), .B(n40249), .Z(n40247) );
  OR U40530 ( .A(n40250), .B(n40251), .Z(n40249) );
  NAND U40531 ( .A(n40251), .B(n40250), .Z(n40246) );
  ANDN U40532 ( .B(B[126]), .A(n59), .Z(n40030) );
  XNOR U40533 ( .A(n40038), .B(n40252), .Z(n40031) );
  XNOR U40534 ( .A(n40037), .B(n40035), .Z(n40252) );
  AND U40535 ( .A(n40253), .B(n40254), .Z(n40035) );
  NANDN U40536 ( .A(n40255), .B(n40256), .Z(n40254) );
  NANDN U40537 ( .A(n40257), .B(n40258), .Z(n40256) );
  NANDN U40538 ( .A(n40258), .B(n40257), .Z(n40253) );
  ANDN U40539 ( .B(B[127]), .A(n60), .Z(n40037) );
  XNOR U40540 ( .A(n40045), .B(n40259), .Z(n40038) );
  XNOR U40541 ( .A(n40044), .B(n40042), .Z(n40259) );
  AND U40542 ( .A(n40260), .B(n40261), .Z(n40042) );
  NANDN U40543 ( .A(n40262), .B(n40263), .Z(n40261) );
  OR U40544 ( .A(n40264), .B(n40265), .Z(n40263) );
  NAND U40545 ( .A(n40265), .B(n40264), .Z(n40260) );
  ANDN U40546 ( .B(B[128]), .A(n61), .Z(n40044) );
  XNOR U40547 ( .A(n40052), .B(n40266), .Z(n40045) );
  XNOR U40548 ( .A(n40051), .B(n40049), .Z(n40266) );
  AND U40549 ( .A(n40267), .B(n40268), .Z(n40049) );
  NANDN U40550 ( .A(n40269), .B(n40270), .Z(n40268) );
  NANDN U40551 ( .A(n40271), .B(n40272), .Z(n40270) );
  NANDN U40552 ( .A(n40272), .B(n40271), .Z(n40267) );
  ANDN U40553 ( .B(B[129]), .A(n62), .Z(n40051) );
  XNOR U40554 ( .A(n40059), .B(n40273), .Z(n40052) );
  XNOR U40555 ( .A(n40058), .B(n40056), .Z(n40273) );
  AND U40556 ( .A(n40274), .B(n40275), .Z(n40056) );
  NANDN U40557 ( .A(n40276), .B(n40277), .Z(n40275) );
  OR U40558 ( .A(n40278), .B(n40279), .Z(n40277) );
  NAND U40559 ( .A(n40279), .B(n40278), .Z(n40274) );
  ANDN U40560 ( .B(B[130]), .A(n63), .Z(n40058) );
  XNOR U40561 ( .A(n40066), .B(n40280), .Z(n40059) );
  XNOR U40562 ( .A(n40065), .B(n40063), .Z(n40280) );
  AND U40563 ( .A(n40281), .B(n40282), .Z(n40063) );
  NANDN U40564 ( .A(n40283), .B(n40284), .Z(n40282) );
  NANDN U40565 ( .A(n40285), .B(n40286), .Z(n40284) );
  NANDN U40566 ( .A(n40286), .B(n40285), .Z(n40281) );
  ANDN U40567 ( .B(B[131]), .A(n64), .Z(n40065) );
  XNOR U40568 ( .A(n40073), .B(n40287), .Z(n40066) );
  XNOR U40569 ( .A(n40072), .B(n40070), .Z(n40287) );
  AND U40570 ( .A(n40288), .B(n40289), .Z(n40070) );
  NANDN U40571 ( .A(n40290), .B(n40291), .Z(n40289) );
  OR U40572 ( .A(n40292), .B(n40293), .Z(n40291) );
  NAND U40573 ( .A(n40293), .B(n40292), .Z(n40288) );
  ANDN U40574 ( .B(B[132]), .A(n65), .Z(n40072) );
  XNOR U40575 ( .A(n40080), .B(n40294), .Z(n40073) );
  XNOR U40576 ( .A(n40079), .B(n40077), .Z(n40294) );
  AND U40577 ( .A(n40295), .B(n40296), .Z(n40077) );
  NANDN U40578 ( .A(n40297), .B(n40298), .Z(n40296) );
  NANDN U40579 ( .A(n40299), .B(n40300), .Z(n40298) );
  NANDN U40580 ( .A(n40300), .B(n40299), .Z(n40295) );
  ANDN U40581 ( .B(B[133]), .A(n66), .Z(n40079) );
  XNOR U40582 ( .A(n40087), .B(n40301), .Z(n40080) );
  XNOR U40583 ( .A(n40086), .B(n40084), .Z(n40301) );
  AND U40584 ( .A(n40302), .B(n40303), .Z(n40084) );
  NANDN U40585 ( .A(n40304), .B(n40305), .Z(n40303) );
  OR U40586 ( .A(n40306), .B(n40307), .Z(n40305) );
  NAND U40587 ( .A(n40307), .B(n40306), .Z(n40302) );
  ANDN U40588 ( .B(B[134]), .A(n67), .Z(n40086) );
  XNOR U40589 ( .A(n40094), .B(n40308), .Z(n40087) );
  XNOR U40590 ( .A(n40093), .B(n40091), .Z(n40308) );
  AND U40591 ( .A(n40309), .B(n40310), .Z(n40091) );
  NANDN U40592 ( .A(n40311), .B(n40312), .Z(n40310) );
  NANDN U40593 ( .A(n40313), .B(n40314), .Z(n40312) );
  NANDN U40594 ( .A(n40314), .B(n40313), .Z(n40309) );
  ANDN U40595 ( .B(B[135]), .A(n68), .Z(n40093) );
  XNOR U40596 ( .A(n40101), .B(n40315), .Z(n40094) );
  XNOR U40597 ( .A(n40100), .B(n40098), .Z(n40315) );
  AND U40598 ( .A(n40316), .B(n40317), .Z(n40098) );
  NANDN U40599 ( .A(n40318), .B(n40319), .Z(n40317) );
  OR U40600 ( .A(n40320), .B(n40321), .Z(n40319) );
  NAND U40601 ( .A(n40321), .B(n40320), .Z(n40316) );
  ANDN U40602 ( .B(B[136]), .A(n69), .Z(n40100) );
  XNOR U40603 ( .A(n40108), .B(n40322), .Z(n40101) );
  XNOR U40604 ( .A(n40107), .B(n40105), .Z(n40322) );
  AND U40605 ( .A(n40323), .B(n40324), .Z(n40105) );
  NANDN U40606 ( .A(n40325), .B(n40326), .Z(n40324) );
  NANDN U40607 ( .A(n40327), .B(n40328), .Z(n40326) );
  NANDN U40608 ( .A(n40328), .B(n40327), .Z(n40323) );
  ANDN U40609 ( .B(B[137]), .A(n70), .Z(n40107) );
  XNOR U40610 ( .A(n40115), .B(n40329), .Z(n40108) );
  XNOR U40611 ( .A(n40114), .B(n40112), .Z(n40329) );
  AND U40612 ( .A(n40330), .B(n40331), .Z(n40112) );
  NANDN U40613 ( .A(n40332), .B(n40333), .Z(n40331) );
  OR U40614 ( .A(n40334), .B(n40335), .Z(n40333) );
  NAND U40615 ( .A(n40335), .B(n40334), .Z(n40330) );
  ANDN U40616 ( .B(B[138]), .A(n71), .Z(n40114) );
  XNOR U40617 ( .A(n40122), .B(n40336), .Z(n40115) );
  XNOR U40618 ( .A(n40121), .B(n40119), .Z(n40336) );
  AND U40619 ( .A(n40337), .B(n40338), .Z(n40119) );
  NANDN U40620 ( .A(n40339), .B(n40340), .Z(n40338) );
  NANDN U40621 ( .A(n40341), .B(n40342), .Z(n40340) );
  NANDN U40622 ( .A(n40342), .B(n40341), .Z(n40337) );
  ANDN U40623 ( .B(B[139]), .A(n72), .Z(n40121) );
  XNOR U40624 ( .A(n40129), .B(n40343), .Z(n40122) );
  XNOR U40625 ( .A(n40128), .B(n40126), .Z(n40343) );
  AND U40626 ( .A(n40344), .B(n40345), .Z(n40126) );
  NANDN U40627 ( .A(n40346), .B(n40347), .Z(n40345) );
  OR U40628 ( .A(n40348), .B(n40349), .Z(n40347) );
  NAND U40629 ( .A(n40349), .B(n40348), .Z(n40344) );
  ANDN U40630 ( .B(B[140]), .A(n73), .Z(n40128) );
  XNOR U40631 ( .A(n40136), .B(n40350), .Z(n40129) );
  XNOR U40632 ( .A(n40135), .B(n40133), .Z(n40350) );
  AND U40633 ( .A(n40351), .B(n40352), .Z(n40133) );
  NANDN U40634 ( .A(n40353), .B(n40354), .Z(n40352) );
  NANDN U40635 ( .A(n40355), .B(n40356), .Z(n40354) );
  NANDN U40636 ( .A(n40356), .B(n40355), .Z(n40351) );
  ANDN U40637 ( .B(B[141]), .A(n74), .Z(n40135) );
  XNOR U40638 ( .A(n40143), .B(n40357), .Z(n40136) );
  XNOR U40639 ( .A(n40142), .B(n40140), .Z(n40357) );
  AND U40640 ( .A(n40358), .B(n40359), .Z(n40140) );
  NANDN U40641 ( .A(n40360), .B(n40361), .Z(n40359) );
  OR U40642 ( .A(n40362), .B(n40363), .Z(n40361) );
  NAND U40643 ( .A(n40363), .B(n40362), .Z(n40358) );
  ANDN U40644 ( .B(B[142]), .A(n75), .Z(n40142) );
  XNOR U40645 ( .A(n40150), .B(n40364), .Z(n40143) );
  XNOR U40646 ( .A(n40149), .B(n40147), .Z(n40364) );
  AND U40647 ( .A(n40365), .B(n40366), .Z(n40147) );
  NANDN U40648 ( .A(n40367), .B(n40368), .Z(n40366) );
  NANDN U40649 ( .A(n40369), .B(n40370), .Z(n40368) );
  NANDN U40650 ( .A(n40370), .B(n40369), .Z(n40365) );
  ANDN U40651 ( .B(B[143]), .A(n76), .Z(n40149) );
  XNOR U40652 ( .A(n40157), .B(n40371), .Z(n40150) );
  XNOR U40653 ( .A(n40156), .B(n40154), .Z(n40371) );
  AND U40654 ( .A(n40372), .B(n40373), .Z(n40154) );
  NANDN U40655 ( .A(n40374), .B(n40375), .Z(n40373) );
  OR U40656 ( .A(n40376), .B(n40377), .Z(n40375) );
  NAND U40657 ( .A(n40377), .B(n40376), .Z(n40372) );
  ANDN U40658 ( .B(B[144]), .A(n77), .Z(n40156) );
  XNOR U40659 ( .A(n40164), .B(n40378), .Z(n40157) );
  XNOR U40660 ( .A(n40163), .B(n40161), .Z(n40378) );
  AND U40661 ( .A(n40379), .B(n40380), .Z(n40161) );
  NANDN U40662 ( .A(n40381), .B(n40382), .Z(n40380) );
  NANDN U40663 ( .A(n40383), .B(n40384), .Z(n40382) );
  NANDN U40664 ( .A(n40384), .B(n40383), .Z(n40379) );
  ANDN U40665 ( .B(B[145]), .A(n78), .Z(n40163) );
  XNOR U40666 ( .A(n40171), .B(n40385), .Z(n40164) );
  XNOR U40667 ( .A(n40170), .B(n40168), .Z(n40385) );
  AND U40668 ( .A(n40386), .B(n40387), .Z(n40168) );
  NANDN U40669 ( .A(n40388), .B(n40389), .Z(n40387) );
  OR U40670 ( .A(n40390), .B(n40391), .Z(n40389) );
  NAND U40671 ( .A(n40391), .B(n40390), .Z(n40386) );
  ANDN U40672 ( .B(B[146]), .A(n79), .Z(n40170) );
  XNOR U40673 ( .A(n40178), .B(n40392), .Z(n40171) );
  XNOR U40674 ( .A(n40177), .B(n40175), .Z(n40392) );
  AND U40675 ( .A(n40393), .B(n40394), .Z(n40175) );
  NANDN U40676 ( .A(n40395), .B(n40396), .Z(n40394) );
  NANDN U40677 ( .A(n40397), .B(n40398), .Z(n40396) );
  NANDN U40678 ( .A(n40398), .B(n40397), .Z(n40393) );
  ANDN U40679 ( .B(B[147]), .A(n80), .Z(n40177) );
  XNOR U40680 ( .A(n40185), .B(n40399), .Z(n40178) );
  XNOR U40681 ( .A(n40184), .B(n40182), .Z(n40399) );
  AND U40682 ( .A(n40400), .B(n40401), .Z(n40182) );
  NANDN U40683 ( .A(n40402), .B(n40403), .Z(n40401) );
  OR U40684 ( .A(n40404), .B(n40405), .Z(n40403) );
  NAND U40685 ( .A(n40405), .B(n40404), .Z(n40400) );
  ANDN U40686 ( .B(B[148]), .A(n81), .Z(n40184) );
  XNOR U40687 ( .A(n40192), .B(n40406), .Z(n40185) );
  XNOR U40688 ( .A(n40191), .B(n40189), .Z(n40406) );
  AND U40689 ( .A(n40407), .B(n40408), .Z(n40189) );
  NANDN U40690 ( .A(n40409), .B(n40410), .Z(n40408) );
  NAND U40691 ( .A(n40411), .B(n40412), .Z(n40410) );
  ANDN U40692 ( .B(B[149]), .A(n82), .Z(n40191) );
  XOR U40693 ( .A(n40198), .B(n40413), .Z(n40192) );
  XNOR U40694 ( .A(n40196), .B(n40199), .Z(n40413) );
  NAND U40695 ( .A(A[2]), .B(B[150]), .Z(n40199) );
  NANDN U40696 ( .A(n40414), .B(n40415), .Z(n40196) );
  AND U40697 ( .A(A[0]), .B(B[151]), .Z(n40415) );
  XNOR U40698 ( .A(n40201), .B(n40416), .Z(n40198) );
  NAND U40699 ( .A(A[0]), .B(B[152]), .Z(n40416) );
  NAND U40700 ( .A(B[151]), .B(A[1]), .Z(n40201) );
  NAND U40701 ( .A(n40417), .B(n40418), .Z(n492) );
  NANDN U40702 ( .A(n40419), .B(n40420), .Z(n40418) );
  OR U40703 ( .A(n40421), .B(n40422), .Z(n40420) );
  NAND U40704 ( .A(n40422), .B(n40421), .Z(n40417) );
  XOR U40705 ( .A(n38190), .B(n40423), .Z(\A1[14] ) );
  XNOR U40706 ( .A(n38189), .B(n38188), .Z(n40423) );
  NAND U40707 ( .A(n40424), .B(n40425), .Z(n38188) );
  NANDN U40708 ( .A(n40426), .B(n40427), .Z(n40425) );
  OR U40709 ( .A(n40428), .B(n40429), .Z(n40427) );
  NAND U40710 ( .A(n40429), .B(n40428), .Z(n40424) );
  ANDN U40711 ( .B(B[0]), .A(n69), .Z(n38189) );
  XNOR U40712 ( .A(n38197), .B(n40430), .Z(n38190) );
  XNOR U40713 ( .A(n38196), .B(n38194), .Z(n40430) );
  AND U40714 ( .A(n40431), .B(n40432), .Z(n38194) );
  NANDN U40715 ( .A(n40433), .B(n40434), .Z(n40432) );
  NANDN U40716 ( .A(n40435), .B(n40436), .Z(n40434) );
  NANDN U40717 ( .A(n40436), .B(n40435), .Z(n40431) );
  ANDN U40718 ( .B(B[1]), .A(n70), .Z(n38196) );
  XNOR U40719 ( .A(n38204), .B(n40437), .Z(n38197) );
  XNOR U40720 ( .A(n38203), .B(n38201), .Z(n40437) );
  AND U40721 ( .A(n40438), .B(n40439), .Z(n38201) );
  NANDN U40722 ( .A(n40440), .B(n40441), .Z(n40439) );
  OR U40723 ( .A(n40442), .B(n40443), .Z(n40441) );
  NAND U40724 ( .A(n40443), .B(n40442), .Z(n40438) );
  ANDN U40725 ( .B(B[2]), .A(n71), .Z(n38203) );
  XNOR U40726 ( .A(n38211), .B(n40444), .Z(n38204) );
  XNOR U40727 ( .A(n38210), .B(n38208), .Z(n40444) );
  AND U40728 ( .A(n40445), .B(n40446), .Z(n38208) );
  NANDN U40729 ( .A(n40447), .B(n40448), .Z(n40446) );
  NANDN U40730 ( .A(n40449), .B(n40450), .Z(n40448) );
  NANDN U40731 ( .A(n40450), .B(n40449), .Z(n40445) );
  ANDN U40732 ( .B(B[3]), .A(n72), .Z(n38210) );
  XNOR U40733 ( .A(n38218), .B(n40451), .Z(n38211) );
  XNOR U40734 ( .A(n38217), .B(n38215), .Z(n40451) );
  AND U40735 ( .A(n40452), .B(n40453), .Z(n38215) );
  NANDN U40736 ( .A(n40454), .B(n40455), .Z(n40453) );
  OR U40737 ( .A(n40456), .B(n40457), .Z(n40455) );
  NAND U40738 ( .A(n40457), .B(n40456), .Z(n40452) );
  ANDN U40739 ( .B(B[4]), .A(n73), .Z(n38217) );
  XNOR U40740 ( .A(n38225), .B(n40458), .Z(n38218) );
  XNOR U40741 ( .A(n38224), .B(n38222), .Z(n40458) );
  AND U40742 ( .A(n40459), .B(n40460), .Z(n38222) );
  NANDN U40743 ( .A(n40461), .B(n40462), .Z(n40460) );
  NANDN U40744 ( .A(n40463), .B(n40464), .Z(n40462) );
  NANDN U40745 ( .A(n40464), .B(n40463), .Z(n40459) );
  ANDN U40746 ( .B(B[5]), .A(n74), .Z(n38224) );
  XNOR U40747 ( .A(n38232), .B(n40465), .Z(n38225) );
  XNOR U40748 ( .A(n38231), .B(n38229), .Z(n40465) );
  AND U40749 ( .A(n40466), .B(n40467), .Z(n38229) );
  NANDN U40750 ( .A(n40468), .B(n40469), .Z(n40467) );
  OR U40751 ( .A(n40470), .B(n40471), .Z(n40469) );
  NAND U40752 ( .A(n40471), .B(n40470), .Z(n40466) );
  ANDN U40753 ( .B(B[6]), .A(n75), .Z(n38231) );
  XNOR U40754 ( .A(n38239), .B(n40472), .Z(n38232) );
  XNOR U40755 ( .A(n38238), .B(n38236), .Z(n40472) );
  AND U40756 ( .A(n40473), .B(n40474), .Z(n38236) );
  NANDN U40757 ( .A(n40475), .B(n40476), .Z(n40474) );
  NANDN U40758 ( .A(n40477), .B(n40478), .Z(n40476) );
  NANDN U40759 ( .A(n40478), .B(n40477), .Z(n40473) );
  ANDN U40760 ( .B(B[7]), .A(n76), .Z(n38238) );
  XNOR U40761 ( .A(n38246), .B(n40479), .Z(n38239) );
  XNOR U40762 ( .A(n38245), .B(n38243), .Z(n40479) );
  AND U40763 ( .A(n40480), .B(n40481), .Z(n38243) );
  NANDN U40764 ( .A(n40482), .B(n40483), .Z(n40481) );
  OR U40765 ( .A(n40484), .B(n40485), .Z(n40483) );
  NAND U40766 ( .A(n40485), .B(n40484), .Z(n40480) );
  ANDN U40767 ( .B(B[8]), .A(n77), .Z(n38245) );
  XNOR U40768 ( .A(n38253), .B(n40486), .Z(n38246) );
  XNOR U40769 ( .A(n38252), .B(n38250), .Z(n40486) );
  AND U40770 ( .A(n40487), .B(n40488), .Z(n38250) );
  NANDN U40771 ( .A(n40489), .B(n40490), .Z(n40488) );
  NANDN U40772 ( .A(n40491), .B(n40492), .Z(n40490) );
  NANDN U40773 ( .A(n40492), .B(n40491), .Z(n40487) );
  ANDN U40774 ( .B(B[9]), .A(n78), .Z(n38252) );
  XNOR U40775 ( .A(n38260), .B(n40493), .Z(n38253) );
  XNOR U40776 ( .A(n38259), .B(n38257), .Z(n40493) );
  AND U40777 ( .A(n40494), .B(n40495), .Z(n38257) );
  NANDN U40778 ( .A(n40496), .B(n40497), .Z(n40495) );
  OR U40779 ( .A(n40498), .B(n40499), .Z(n40497) );
  NAND U40780 ( .A(n40499), .B(n40498), .Z(n40494) );
  ANDN U40781 ( .B(B[10]), .A(n79), .Z(n38259) );
  XNOR U40782 ( .A(n38267), .B(n40500), .Z(n38260) );
  XNOR U40783 ( .A(n38266), .B(n38264), .Z(n40500) );
  AND U40784 ( .A(n40501), .B(n40502), .Z(n38264) );
  NANDN U40785 ( .A(n40503), .B(n40504), .Z(n40502) );
  NANDN U40786 ( .A(n40505), .B(n40506), .Z(n40504) );
  NANDN U40787 ( .A(n40506), .B(n40505), .Z(n40501) );
  ANDN U40788 ( .B(B[11]), .A(n80), .Z(n38266) );
  XNOR U40789 ( .A(n38274), .B(n40507), .Z(n38267) );
  XNOR U40790 ( .A(n38273), .B(n38271), .Z(n40507) );
  AND U40791 ( .A(n40508), .B(n40509), .Z(n38271) );
  NANDN U40792 ( .A(n40510), .B(n40511), .Z(n40509) );
  OR U40793 ( .A(n40512), .B(n40513), .Z(n40511) );
  NAND U40794 ( .A(n40513), .B(n40512), .Z(n40508) );
  ANDN U40795 ( .B(B[12]), .A(n81), .Z(n38273) );
  XNOR U40796 ( .A(n38281), .B(n40514), .Z(n38274) );
  XNOR U40797 ( .A(n38280), .B(n38278), .Z(n40514) );
  AND U40798 ( .A(n40515), .B(n40516), .Z(n38278) );
  NANDN U40799 ( .A(n40517), .B(n40518), .Z(n40516) );
  NAND U40800 ( .A(n40519), .B(n40520), .Z(n40518) );
  ANDN U40801 ( .B(B[13]), .A(n82), .Z(n38280) );
  XOR U40802 ( .A(n38287), .B(n40521), .Z(n38281) );
  XNOR U40803 ( .A(n38285), .B(n38288), .Z(n40521) );
  NAND U40804 ( .A(A[2]), .B(B[14]), .Z(n38288) );
  NANDN U40805 ( .A(n40522), .B(n40523), .Z(n38285) );
  AND U40806 ( .A(A[0]), .B(B[15]), .Z(n40523) );
  XNOR U40807 ( .A(n38290), .B(n40524), .Z(n38287) );
  NAND U40808 ( .A(A[0]), .B(B[16]), .Z(n40524) );
  NAND U40809 ( .A(B[15]), .B(A[1]), .Z(n38290) );
  XOR U40810 ( .A(n494), .B(n493), .Z(\A1[149] ) );
  XOR U40811 ( .A(n40422), .B(n40525), .Z(n493) );
  XNOR U40812 ( .A(n40421), .B(n40419), .Z(n40525) );
  AND U40813 ( .A(n40526), .B(n40527), .Z(n40419) );
  NANDN U40814 ( .A(n40528), .B(n40529), .Z(n40527) );
  NANDN U40815 ( .A(n40530), .B(n40531), .Z(n40529) );
  NANDN U40816 ( .A(n40531), .B(n40530), .Z(n40526) );
  ANDN U40817 ( .B(B[120]), .A(n54), .Z(n40421) );
  XNOR U40818 ( .A(n40216), .B(n40532), .Z(n40422) );
  XNOR U40819 ( .A(n40215), .B(n40213), .Z(n40532) );
  AND U40820 ( .A(n40533), .B(n40534), .Z(n40213) );
  NANDN U40821 ( .A(n40535), .B(n40536), .Z(n40534) );
  OR U40822 ( .A(n40537), .B(n40538), .Z(n40536) );
  NAND U40823 ( .A(n40538), .B(n40537), .Z(n40533) );
  ANDN U40824 ( .B(B[121]), .A(n55), .Z(n40215) );
  XNOR U40825 ( .A(n40223), .B(n40539), .Z(n40216) );
  XNOR U40826 ( .A(n40222), .B(n40220), .Z(n40539) );
  AND U40827 ( .A(n40540), .B(n40541), .Z(n40220) );
  NANDN U40828 ( .A(n40542), .B(n40543), .Z(n40541) );
  NANDN U40829 ( .A(n40544), .B(n40545), .Z(n40543) );
  NANDN U40830 ( .A(n40545), .B(n40544), .Z(n40540) );
  ANDN U40831 ( .B(B[122]), .A(n56), .Z(n40222) );
  XNOR U40832 ( .A(n40230), .B(n40546), .Z(n40223) );
  XNOR U40833 ( .A(n40229), .B(n40227), .Z(n40546) );
  AND U40834 ( .A(n40547), .B(n40548), .Z(n40227) );
  NANDN U40835 ( .A(n40549), .B(n40550), .Z(n40548) );
  OR U40836 ( .A(n40551), .B(n40552), .Z(n40550) );
  NAND U40837 ( .A(n40552), .B(n40551), .Z(n40547) );
  ANDN U40838 ( .B(B[123]), .A(n57), .Z(n40229) );
  XNOR U40839 ( .A(n40237), .B(n40553), .Z(n40230) );
  XNOR U40840 ( .A(n40236), .B(n40234), .Z(n40553) );
  AND U40841 ( .A(n40554), .B(n40555), .Z(n40234) );
  NANDN U40842 ( .A(n40556), .B(n40557), .Z(n40555) );
  NANDN U40843 ( .A(n40558), .B(n40559), .Z(n40557) );
  NANDN U40844 ( .A(n40559), .B(n40558), .Z(n40554) );
  ANDN U40845 ( .B(B[124]), .A(n58), .Z(n40236) );
  XNOR U40846 ( .A(n40244), .B(n40560), .Z(n40237) );
  XNOR U40847 ( .A(n40243), .B(n40241), .Z(n40560) );
  AND U40848 ( .A(n40561), .B(n40562), .Z(n40241) );
  NANDN U40849 ( .A(n40563), .B(n40564), .Z(n40562) );
  OR U40850 ( .A(n40565), .B(n40566), .Z(n40564) );
  NAND U40851 ( .A(n40566), .B(n40565), .Z(n40561) );
  ANDN U40852 ( .B(B[125]), .A(n59), .Z(n40243) );
  XNOR U40853 ( .A(n40251), .B(n40567), .Z(n40244) );
  XNOR U40854 ( .A(n40250), .B(n40248), .Z(n40567) );
  AND U40855 ( .A(n40568), .B(n40569), .Z(n40248) );
  NANDN U40856 ( .A(n40570), .B(n40571), .Z(n40569) );
  NANDN U40857 ( .A(n40572), .B(n40573), .Z(n40571) );
  NANDN U40858 ( .A(n40573), .B(n40572), .Z(n40568) );
  ANDN U40859 ( .B(B[126]), .A(n60), .Z(n40250) );
  XNOR U40860 ( .A(n40258), .B(n40574), .Z(n40251) );
  XNOR U40861 ( .A(n40257), .B(n40255), .Z(n40574) );
  AND U40862 ( .A(n40575), .B(n40576), .Z(n40255) );
  NANDN U40863 ( .A(n40577), .B(n40578), .Z(n40576) );
  OR U40864 ( .A(n40579), .B(n40580), .Z(n40578) );
  NAND U40865 ( .A(n40580), .B(n40579), .Z(n40575) );
  ANDN U40866 ( .B(B[127]), .A(n61), .Z(n40257) );
  XNOR U40867 ( .A(n40265), .B(n40581), .Z(n40258) );
  XNOR U40868 ( .A(n40264), .B(n40262), .Z(n40581) );
  AND U40869 ( .A(n40582), .B(n40583), .Z(n40262) );
  NANDN U40870 ( .A(n40584), .B(n40585), .Z(n40583) );
  NANDN U40871 ( .A(n40586), .B(n40587), .Z(n40585) );
  NANDN U40872 ( .A(n40587), .B(n40586), .Z(n40582) );
  ANDN U40873 ( .B(B[128]), .A(n62), .Z(n40264) );
  XNOR U40874 ( .A(n40272), .B(n40588), .Z(n40265) );
  XNOR U40875 ( .A(n40271), .B(n40269), .Z(n40588) );
  AND U40876 ( .A(n40589), .B(n40590), .Z(n40269) );
  NANDN U40877 ( .A(n40591), .B(n40592), .Z(n40590) );
  OR U40878 ( .A(n40593), .B(n40594), .Z(n40592) );
  NAND U40879 ( .A(n40594), .B(n40593), .Z(n40589) );
  ANDN U40880 ( .B(B[129]), .A(n63), .Z(n40271) );
  XNOR U40881 ( .A(n40279), .B(n40595), .Z(n40272) );
  XNOR U40882 ( .A(n40278), .B(n40276), .Z(n40595) );
  AND U40883 ( .A(n40596), .B(n40597), .Z(n40276) );
  NANDN U40884 ( .A(n40598), .B(n40599), .Z(n40597) );
  NANDN U40885 ( .A(n40600), .B(n40601), .Z(n40599) );
  NANDN U40886 ( .A(n40601), .B(n40600), .Z(n40596) );
  ANDN U40887 ( .B(B[130]), .A(n64), .Z(n40278) );
  XNOR U40888 ( .A(n40286), .B(n40602), .Z(n40279) );
  XNOR U40889 ( .A(n40285), .B(n40283), .Z(n40602) );
  AND U40890 ( .A(n40603), .B(n40604), .Z(n40283) );
  NANDN U40891 ( .A(n40605), .B(n40606), .Z(n40604) );
  OR U40892 ( .A(n40607), .B(n40608), .Z(n40606) );
  NAND U40893 ( .A(n40608), .B(n40607), .Z(n40603) );
  ANDN U40894 ( .B(B[131]), .A(n65), .Z(n40285) );
  XNOR U40895 ( .A(n40293), .B(n40609), .Z(n40286) );
  XNOR U40896 ( .A(n40292), .B(n40290), .Z(n40609) );
  AND U40897 ( .A(n40610), .B(n40611), .Z(n40290) );
  NANDN U40898 ( .A(n40612), .B(n40613), .Z(n40611) );
  NANDN U40899 ( .A(n40614), .B(n40615), .Z(n40613) );
  NANDN U40900 ( .A(n40615), .B(n40614), .Z(n40610) );
  ANDN U40901 ( .B(B[132]), .A(n66), .Z(n40292) );
  XNOR U40902 ( .A(n40300), .B(n40616), .Z(n40293) );
  XNOR U40903 ( .A(n40299), .B(n40297), .Z(n40616) );
  AND U40904 ( .A(n40617), .B(n40618), .Z(n40297) );
  NANDN U40905 ( .A(n40619), .B(n40620), .Z(n40618) );
  OR U40906 ( .A(n40621), .B(n40622), .Z(n40620) );
  NAND U40907 ( .A(n40622), .B(n40621), .Z(n40617) );
  ANDN U40908 ( .B(B[133]), .A(n67), .Z(n40299) );
  XNOR U40909 ( .A(n40307), .B(n40623), .Z(n40300) );
  XNOR U40910 ( .A(n40306), .B(n40304), .Z(n40623) );
  AND U40911 ( .A(n40624), .B(n40625), .Z(n40304) );
  NANDN U40912 ( .A(n40626), .B(n40627), .Z(n40625) );
  NANDN U40913 ( .A(n40628), .B(n40629), .Z(n40627) );
  NANDN U40914 ( .A(n40629), .B(n40628), .Z(n40624) );
  ANDN U40915 ( .B(B[134]), .A(n68), .Z(n40306) );
  XNOR U40916 ( .A(n40314), .B(n40630), .Z(n40307) );
  XNOR U40917 ( .A(n40313), .B(n40311), .Z(n40630) );
  AND U40918 ( .A(n40631), .B(n40632), .Z(n40311) );
  NANDN U40919 ( .A(n40633), .B(n40634), .Z(n40632) );
  OR U40920 ( .A(n40635), .B(n40636), .Z(n40634) );
  NAND U40921 ( .A(n40636), .B(n40635), .Z(n40631) );
  ANDN U40922 ( .B(B[135]), .A(n69), .Z(n40313) );
  XNOR U40923 ( .A(n40321), .B(n40637), .Z(n40314) );
  XNOR U40924 ( .A(n40320), .B(n40318), .Z(n40637) );
  AND U40925 ( .A(n40638), .B(n40639), .Z(n40318) );
  NANDN U40926 ( .A(n40640), .B(n40641), .Z(n40639) );
  NANDN U40927 ( .A(n40642), .B(n40643), .Z(n40641) );
  NANDN U40928 ( .A(n40643), .B(n40642), .Z(n40638) );
  ANDN U40929 ( .B(B[136]), .A(n70), .Z(n40320) );
  XNOR U40930 ( .A(n40328), .B(n40644), .Z(n40321) );
  XNOR U40931 ( .A(n40327), .B(n40325), .Z(n40644) );
  AND U40932 ( .A(n40645), .B(n40646), .Z(n40325) );
  NANDN U40933 ( .A(n40647), .B(n40648), .Z(n40646) );
  OR U40934 ( .A(n40649), .B(n40650), .Z(n40648) );
  NAND U40935 ( .A(n40650), .B(n40649), .Z(n40645) );
  ANDN U40936 ( .B(B[137]), .A(n71), .Z(n40327) );
  XNOR U40937 ( .A(n40335), .B(n40651), .Z(n40328) );
  XNOR U40938 ( .A(n40334), .B(n40332), .Z(n40651) );
  AND U40939 ( .A(n40652), .B(n40653), .Z(n40332) );
  NANDN U40940 ( .A(n40654), .B(n40655), .Z(n40653) );
  NANDN U40941 ( .A(n40656), .B(n40657), .Z(n40655) );
  NANDN U40942 ( .A(n40657), .B(n40656), .Z(n40652) );
  ANDN U40943 ( .B(B[138]), .A(n72), .Z(n40334) );
  XNOR U40944 ( .A(n40342), .B(n40658), .Z(n40335) );
  XNOR U40945 ( .A(n40341), .B(n40339), .Z(n40658) );
  AND U40946 ( .A(n40659), .B(n40660), .Z(n40339) );
  NANDN U40947 ( .A(n40661), .B(n40662), .Z(n40660) );
  OR U40948 ( .A(n40663), .B(n40664), .Z(n40662) );
  NAND U40949 ( .A(n40664), .B(n40663), .Z(n40659) );
  ANDN U40950 ( .B(B[139]), .A(n73), .Z(n40341) );
  XNOR U40951 ( .A(n40349), .B(n40665), .Z(n40342) );
  XNOR U40952 ( .A(n40348), .B(n40346), .Z(n40665) );
  AND U40953 ( .A(n40666), .B(n40667), .Z(n40346) );
  NANDN U40954 ( .A(n40668), .B(n40669), .Z(n40667) );
  NANDN U40955 ( .A(n40670), .B(n40671), .Z(n40669) );
  NANDN U40956 ( .A(n40671), .B(n40670), .Z(n40666) );
  ANDN U40957 ( .B(B[140]), .A(n74), .Z(n40348) );
  XNOR U40958 ( .A(n40356), .B(n40672), .Z(n40349) );
  XNOR U40959 ( .A(n40355), .B(n40353), .Z(n40672) );
  AND U40960 ( .A(n40673), .B(n40674), .Z(n40353) );
  NANDN U40961 ( .A(n40675), .B(n40676), .Z(n40674) );
  OR U40962 ( .A(n40677), .B(n40678), .Z(n40676) );
  NAND U40963 ( .A(n40678), .B(n40677), .Z(n40673) );
  ANDN U40964 ( .B(B[141]), .A(n75), .Z(n40355) );
  XNOR U40965 ( .A(n40363), .B(n40679), .Z(n40356) );
  XNOR U40966 ( .A(n40362), .B(n40360), .Z(n40679) );
  AND U40967 ( .A(n40680), .B(n40681), .Z(n40360) );
  NANDN U40968 ( .A(n40682), .B(n40683), .Z(n40681) );
  NANDN U40969 ( .A(n40684), .B(n40685), .Z(n40683) );
  NANDN U40970 ( .A(n40685), .B(n40684), .Z(n40680) );
  ANDN U40971 ( .B(B[142]), .A(n76), .Z(n40362) );
  XNOR U40972 ( .A(n40370), .B(n40686), .Z(n40363) );
  XNOR U40973 ( .A(n40369), .B(n40367), .Z(n40686) );
  AND U40974 ( .A(n40687), .B(n40688), .Z(n40367) );
  NANDN U40975 ( .A(n40689), .B(n40690), .Z(n40688) );
  OR U40976 ( .A(n40691), .B(n40692), .Z(n40690) );
  NAND U40977 ( .A(n40692), .B(n40691), .Z(n40687) );
  ANDN U40978 ( .B(B[143]), .A(n77), .Z(n40369) );
  XNOR U40979 ( .A(n40377), .B(n40693), .Z(n40370) );
  XNOR U40980 ( .A(n40376), .B(n40374), .Z(n40693) );
  AND U40981 ( .A(n40694), .B(n40695), .Z(n40374) );
  NANDN U40982 ( .A(n40696), .B(n40697), .Z(n40695) );
  NANDN U40983 ( .A(n40698), .B(n40699), .Z(n40697) );
  NANDN U40984 ( .A(n40699), .B(n40698), .Z(n40694) );
  ANDN U40985 ( .B(B[144]), .A(n78), .Z(n40376) );
  XNOR U40986 ( .A(n40384), .B(n40700), .Z(n40377) );
  XNOR U40987 ( .A(n40383), .B(n40381), .Z(n40700) );
  AND U40988 ( .A(n40701), .B(n40702), .Z(n40381) );
  NANDN U40989 ( .A(n40703), .B(n40704), .Z(n40702) );
  OR U40990 ( .A(n40705), .B(n40706), .Z(n40704) );
  NAND U40991 ( .A(n40706), .B(n40705), .Z(n40701) );
  ANDN U40992 ( .B(B[145]), .A(n79), .Z(n40383) );
  XNOR U40993 ( .A(n40391), .B(n40707), .Z(n40384) );
  XNOR U40994 ( .A(n40390), .B(n40388), .Z(n40707) );
  AND U40995 ( .A(n40708), .B(n40709), .Z(n40388) );
  NANDN U40996 ( .A(n40710), .B(n40711), .Z(n40709) );
  NANDN U40997 ( .A(n40712), .B(n40713), .Z(n40711) );
  NANDN U40998 ( .A(n40713), .B(n40712), .Z(n40708) );
  ANDN U40999 ( .B(B[146]), .A(n80), .Z(n40390) );
  XNOR U41000 ( .A(n40398), .B(n40714), .Z(n40391) );
  XNOR U41001 ( .A(n40397), .B(n40395), .Z(n40714) );
  AND U41002 ( .A(n40715), .B(n40716), .Z(n40395) );
  NANDN U41003 ( .A(n40717), .B(n40718), .Z(n40716) );
  OR U41004 ( .A(n40719), .B(n40720), .Z(n40718) );
  NAND U41005 ( .A(n40720), .B(n40719), .Z(n40715) );
  ANDN U41006 ( .B(B[147]), .A(n81), .Z(n40397) );
  XNOR U41007 ( .A(n40405), .B(n40721), .Z(n40398) );
  XNOR U41008 ( .A(n40404), .B(n40402), .Z(n40721) );
  AND U41009 ( .A(n40722), .B(n40723), .Z(n40402) );
  NANDN U41010 ( .A(n40724), .B(n40725), .Z(n40723) );
  NAND U41011 ( .A(n40726), .B(n40727), .Z(n40725) );
  ANDN U41012 ( .B(B[148]), .A(n82), .Z(n40404) );
  XOR U41013 ( .A(n40411), .B(n40728), .Z(n40405) );
  XNOR U41014 ( .A(n40409), .B(n40412), .Z(n40728) );
  NAND U41015 ( .A(A[2]), .B(B[149]), .Z(n40412) );
  NANDN U41016 ( .A(n40729), .B(n40730), .Z(n40409) );
  AND U41017 ( .A(A[0]), .B(B[150]), .Z(n40730) );
  XNOR U41018 ( .A(n40414), .B(n40731), .Z(n40411) );
  NAND U41019 ( .A(A[0]), .B(B[151]), .Z(n40731) );
  NAND U41020 ( .A(B[150]), .B(A[1]), .Z(n40414) );
  NAND U41021 ( .A(n40732), .B(n40733), .Z(n494) );
  NANDN U41022 ( .A(n40734), .B(n40735), .Z(n40733) );
  OR U41023 ( .A(n40736), .B(n40737), .Z(n40735) );
  NAND U41024 ( .A(n40737), .B(n40736), .Z(n40732) );
  XOR U41025 ( .A(n496), .B(n495), .Z(\A1[148] ) );
  XOR U41026 ( .A(n40737), .B(n40738), .Z(n495) );
  XNOR U41027 ( .A(n40736), .B(n40734), .Z(n40738) );
  AND U41028 ( .A(n40739), .B(n40740), .Z(n40734) );
  NANDN U41029 ( .A(n40741), .B(n40742), .Z(n40740) );
  NANDN U41030 ( .A(n40743), .B(n40744), .Z(n40742) );
  NANDN U41031 ( .A(n40744), .B(n40743), .Z(n40739) );
  ANDN U41032 ( .B(B[119]), .A(n54), .Z(n40736) );
  XNOR U41033 ( .A(n40531), .B(n40745), .Z(n40737) );
  XNOR U41034 ( .A(n40530), .B(n40528), .Z(n40745) );
  AND U41035 ( .A(n40746), .B(n40747), .Z(n40528) );
  NANDN U41036 ( .A(n40748), .B(n40749), .Z(n40747) );
  OR U41037 ( .A(n40750), .B(n40751), .Z(n40749) );
  NAND U41038 ( .A(n40751), .B(n40750), .Z(n40746) );
  ANDN U41039 ( .B(B[120]), .A(n55), .Z(n40530) );
  XNOR U41040 ( .A(n40538), .B(n40752), .Z(n40531) );
  XNOR U41041 ( .A(n40537), .B(n40535), .Z(n40752) );
  AND U41042 ( .A(n40753), .B(n40754), .Z(n40535) );
  NANDN U41043 ( .A(n40755), .B(n40756), .Z(n40754) );
  NANDN U41044 ( .A(n40757), .B(n40758), .Z(n40756) );
  NANDN U41045 ( .A(n40758), .B(n40757), .Z(n40753) );
  ANDN U41046 ( .B(B[121]), .A(n56), .Z(n40537) );
  XNOR U41047 ( .A(n40545), .B(n40759), .Z(n40538) );
  XNOR U41048 ( .A(n40544), .B(n40542), .Z(n40759) );
  AND U41049 ( .A(n40760), .B(n40761), .Z(n40542) );
  NANDN U41050 ( .A(n40762), .B(n40763), .Z(n40761) );
  OR U41051 ( .A(n40764), .B(n40765), .Z(n40763) );
  NAND U41052 ( .A(n40765), .B(n40764), .Z(n40760) );
  ANDN U41053 ( .B(B[122]), .A(n57), .Z(n40544) );
  XNOR U41054 ( .A(n40552), .B(n40766), .Z(n40545) );
  XNOR U41055 ( .A(n40551), .B(n40549), .Z(n40766) );
  AND U41056 ( .A(n40767), .B(n40768), .Z(n40549) );
  NANDN U41057 ( .A(n40769), .B(n40770), .Z(n40768) );
  NANDN U41058 ( .A(n40771), .B(n40772), .Z(n40770) );
  NANDN U41059 ( .A(n40772), .B(n40771), .Z(n40767) );
  ANDN U41060 ( .B(B[123]), .A(n58), .Z(n40551) );
  XNOR U41061 ( .A(n40559), .B(n40773), .Z(n40552) );
  XNOR U41062 ( .A(n40558), .B(n40556), .Z(n40773) );
  AND U41063 ( .A(n40774), .B(n40775), .Z(n40556) );
  NANDN U41064 ( .A(n40776), .B(n40777), .Z(n40775) );
  OR U41065 ( .A(n40778), .B(n40779), .Z(n40777) );
  NAND U41066 ( .A(n40779), .B(n40778), .Z(n40774) );
  ANDN U41067 ( .B(B[124]), .A(n59), .Z(n40558) );
  XNOR U41068 ( .A(n40566), .B(n40780), .Z(n40559) );
  XNOR U41069 ( .A(n40565), .B(n40563), .Z(n40780) );
  AND U41070 ( .A(n40781), .B(n40782), .Z(n40563) );
  NANDN U41071 ( .A(n40783), .B(n40784), .Z(n40782) );
  NANDN U41072 ( .A(n40785), .B(n40786), .Z(n40784) );
  NANDN U41073 ( .A(n40786), .B(n40785), .Z(n40781) );
  ANDN U41074 ( .B(B[125]), .A(n60), .Z(n40565) );
  XNOR U41075 ( .A(n40573), .B(n40787), .Z(n40566) );
  XNOR U41076 ( .A(n40572), .B(n40570), .Z(n40787) );
  AND U41077 ( .A(n40788), .B(n40789), .Z(n40570) );
  NANDN U41078 ( .A(n40790), .B(n40791), .Z(n40789) );
  OR U41079 ( .A(n40792), .B(n40793), .Z(n40791) );
  NAND U41080 ( .A(n40793), .B(n40792), .Z(n40788) );
  ANDN U41081 ( .B(B[126]), .A(n61), .Z(n40572) );
  XNOR U41082 ( .A(n40580), .B(n40794), .Z(n40573) );
  XNOR U41083 ( .A(n40579), .B(n40577), .Z(n40794) );
  AND U41084 ( .A(n40795), .B(n40796), .Z(n40577) );
  NANDN U41085 ( .A(n40797), .B(n40798), .Z(n40796) );
  NANDN U41086 ( .A(n40799), .B(n40800), .Z(n40798) );
  NANDN U41087 ( .A(n40800), .B(n40799), .Z(n40795) );
  ANDN U41088 ( .B(B[127]), .A(n62), .Z(n40579) );
  XNOR U41089 ( .A(n40587), .B(n40801), .Z(n40580) );
  XNOR U41090 ( .A(n40586), .B(n40584), .Z(n40801) );
  AND U41091 ( .A(n40802), .B(n40803), .Z(n40584) );
  NANDN U41092 ( .A(n40804), .B(n40805), .Z(n40803) );
  OR U41093 ( .A(n40806), .B(n40807), .Z(n40805) );
  NAND U41094 ( .A(n40807), .B(n40806), .Z(n40802) );
  ANDN U41095 ( .B(B[128]), .A(n63), .Z(n40586) );
  XNOR U41096 ( .A(n40594), .B(n40808), .Z(n40587) );
  XNOR U41097 ( .A(n40593), .B(n40591), .Z(n40808) );
  AND U41098 ( .A(n40809), .B(n40810), .Z(n40591) );
  NANDN U41099 ( .A(n40811), .B(n40812), .Z(n40810) );
  NANDN U41100 ( .A(n40813), .B(n40814), .Z(n40812) );
  NANDN U41101 ( .A(n40814), .B(n40813), .Z(n40809) );
  ANDN U41102 ( .B(B[129]), .A(n64), .Z(n40593) );
  XNOR U41103 ( .A(n40601), .B(n40815), .Z(n40594) );
  XNOR U41104 ( .A(n40600), .B(n40598), .Z(n40815) );
  AND U41105 ( .A(n40816), .B(n40817), .Z(n40598) );
  NANDN U41106 ( .A(n40818), .B(n40819), .Z(n40817) );
  OR U41107 ( .A(n40820), .B(n40821), .Z(n40819) );
  NAND U41108 ( .A(n40821), .B(n40820), .Z(n40816) );
  ANDN U41109 ( .B(B[130]), .A(n65), .Z(n40600) );
  XNOR U41110 ( .A(n40608), .B(n40822), .Z(n40601) );
  XNOR U41111 ( .A(n40607), .B(n40605), .Z(n40822) );
  AND U41112 ( .A(n40823), .B(n40824), .Z(n40605) );
  NANDN U41113 ( .A(n40825), .B(n40826), .Z(n40824) );
  NANDN U41114 ( .A(n40827), .B(n40828), .Z(n40826) );
  NANDN U41115 ( .A(n40828), .B(n40827), .Z(n40823) );
  ANDN U41116 ( .B(B[131]), .A(n66), .Z(n40607) );
  XNOR U41117 ( .A(n40615), .B(n40829), .Z(n40608) );
  XNOR U41118 ( .A(n40614), .B(n40612), .Z(n40829) );
  AND U41119 ( .A(n40830), .B(n40831), .Z(n40612) );
  NANDN U41120 ( .A(n40832), .B(n40833), .Z(n40831) );
  OR U41121 ( .A(n40834), .B(n40835), .Z(n40833) );
  NAND U41122 ( .A(n40835), .B(n40834), .Z(n40830) );
  ANDN U41123 ( .B(B[132]), .A(n67), .Z(n40614) );
  XNOR U41124 ( .A(n40622), .B(n40836), .Z(n40615) );
  XNOR U41125 ( .A(n40621), .B(n40619), .Z(n40836) );
  AND U41126 ( .A(n40837), .B(n40838), .Z(n40619) );
  NANDN U41127 ( .A(n40839), .B(n40840), .Z(n40838) );
  NANDN U41128 ( .A(n40841), .B(n40842), .Z(n40840) );
  NANDN U41129 ( .A(n40842), .B(n40841), .Z(n40837) );
  ANDN U41130 ( .B(B[133]), .A(n68), .Z(n40621) );
  XNOR U41131 ( .A(n40629), .B(n40843), .Z(n40622) );
  XNOR U41132 ( .A(n40628), .B(n40626), .Z(n40843) );
  AND U41133 ( .A(n40844), .B(n40845), .Z(n40626) );
  NANDN U41134 ( .A(n40846), .B(n40847), .Z(n40845) );
  OR U41135 ( .A(n40848), .B(n40849), .Z(n40847) );
  NAND U41136 ( .A(n40849), .B(n40848), .Z(n40844) );
  ANDN U41137 ( .B(B[134]), .A(n69), .Z(n40628) );
  XNOR U41138 ( .A(n40636), .B(n40850), .Z(n40629) );
  XNOR U41139 ( .A(n40635), .B(n40633), .Z(n40850) );
  AND U41140 ( .A(n40851), .B(n40852), .Z(n40633) );
  NANDN U41141 ( .A(n40853), .B(n40854), .Z(n40852) );
  NANDN U41142 ( .A(n40855), .B(n40856), .Z(n40854) );
  NANDN U41143 ( .A(n40856), .B(n40855), .Z(n40851) );
  ANDN U41144 ( .B(B[135]), .A(n70), .Z(n40635) );
  XNOR U41145 ( .A(n40643), .B(n40857), .Z(n40636) );
  XNOR U41146 ( .A(n40642), .B(n40640), .Z(n40857) );
  AND U41147 ( .A(n40858), .B(n40859), .Z(n40640) );
  NANDN U41148 ( .A(n40860), .B(n40861), .Z(n40859) );
  OR U41149 ( .A(n40862), .B(n40863), .Z(n40861) );
  NAND U41150 ( .A(n40863), .B(n40862), .Z(n40858) );
  ANDN U41151 ( .B(B[136]), .A(n71), .Z(n40642) );
  XNOR U41152 ( .A(n40650), .B(n40864), .Z(n40643) );
  XNOR U41153 ( .A(n40649), .B(n40647), .Z(n40864) );
  AND U41154 ( .A(n40865), .B(n40866), .Z(n40647) );
  NANDN U41155 ( .A(n40867), .B(n40868), .Z(n40866) );
  NANDN U41156 ( .A(n40869), .B(n40870), .Z(n40868) );
  NANDN U41157 ( .A(n40870), .B(n40869), .Z(n40865) );
  ANDN U41158 ( .B(B[137]), .A(n72), .Z(n40649) );
  XNOR U41159 ( .A(n40657), .B(n40871), .Z(n40650) );
  XNOR U41160 ( .A(n40656), .B(n40654), .Z(n40871) );
  AND U41161 ( .A(n40872), .B(n40873), .Z(n40654) );
  NANDN U41162 ( .A(n40874), .B(n40875), .Z(n40873) );
  OR U41163 ( .A(n40876), .B(n40877), .Z(n40875) );
  NAND U41164 ( .A(n40877), .B(n40876), .Z(n40872) );
  ANDN U41165 ( .B(B[138]), .A(n73), .Z(n40656) );
  XNOR U41166 ( .A(n40664), .B(n40878), .Z(n40657) );
  XNOR U41167 ( .A(n40663), .B(n40661), .Z(n40878) );
  AND U41168 ( .A(n40879), .B(n40880), .Z(n40661) );
  NANDN U41169 ( .A(n40881), .B(n40882), .Z(n40880) );
  NANDN U41170 ( .A(n40883), .B(n40884), .Z(n40882) );
  NANDN U41171 ( .A(n40884), .B(n40883), .Z(n40879) );
  ANDN U41172 ( .B(B[139]), .A(n74), .Z(n40663) );
  XNOR U41173 ( .A(n40671), .B(n40885), .Z(n40664) );
  XNOR U41174 ( .A(n40670), .B(n40668), .Z(n40885) );
  AND U41175 ( .A(n40886), .B(n40887), .Z(n40668) );
  NANDN U41176 ( .A(n40888), .B(n40889), .Z(n40887) );
  OR U41177 ( .A(n40890), .B(n40891), .Z(n40889) );
  NAND U41178 ( .A(n40891), .B(n40890), .Z(n40886) );
  ANDN U41179 ( .B(B[140]), .A(n75), .Z(n40670) );
  XNOR U41180 ( .A(n40678), .B(n40892), .Z(n40671) );
  XNOR U41181 ( .A(n40677), .B(n40675), .Z(n40892) );
  AND U41182 ( .A(n40893), .B(n40894), .Z(n40675) );
  NANDN U41183 ( .A(n40895), .B(n40896), .Z(n40894) );
  NANDN U41184 ( .A(n40897), .B(n40898), .Z(n40896) );
  NANDN U41185 ( .A(n40898), .B(n40897), .Z(n40893) );
  ANDN U41186 ( .B(B[141]), .A(n76), .Z(n40677) );
  XNOR U41187 ( .A(n40685), .B(n40899), .Z(n40678) );
  XNOR U41188 ( .A(n40684), .B(n40682), .Z(n40899) );
  AND U41189 ( .A(n40900), .B(n40901), .Z(n40682) );
  NANDN U41190 ( .A(n40902), .B(n40903), .Z(n40901) );
  OR U41191 ( .A(n40904), .B(n40905), .Z(n40903) );
  NAND U41192 ( .A(n40905), .B(n40904), .Z(n40900) );
  ANDN U41193 ( .B(B[142]), .A(n77), .Z(n40684) );
  XNOR U41194 ( .A(n40692), .B(n40906), .Z(n40685) );
  XNOR U41195 ( .A(n40691), .B(n40689), .Z(n40906) );
  AND U41196 ( .A(n40907), .B(n40908), .Z(n40689) );
  NANDN U41197 ( .A(n40909), .B(n40910), .Z(n40908) );
  NANDN U41198 ( .A(n40911), .B(n40912), .Z(n40910) );
  NANDN U41199 ( .A(n40912), .B(n40911), .Z(n40907) );
  ANDN U41200 ( .B(B[143]), .A(n78), .Z(n40691) );
  XNOR U41201 ( .A(n40699), .B(n40913), .Z(n40692) );
  XNOR U41202 ( .A(n40698), .B(n40696), .Z(n40913) );
  AND U41203 ( .A(n40914), .B(n40915), .Z(n40696) );
  NANDN U41204 ( .A(n40916), .B(n40917), .Z(n40915) );
  OR U41205 ( .A(n40918), .B(n40919), .Z(n40917) );
  NAND U41206 ( .A(n40919), .B(n40918), .Z(n40914) );
  ANDN U41207 ( .B(B[144]), .A(n79), .Z(n40698) );
  XNOR U41208 ( .A(n40706), .B(n40920), .Z(n40699) );
  XNOR U41209 ( .A(n40705), .B(n40703), .Z(n40920) );
  AND U41210 ( .A(n40921), .B(n40922), .Z(n40703) );
  NANDN U41211 ( .A(n40923), .B(n40924), .Z(n40922) );
  NANDN U41212 ( .A(n40925), .B(n40926), .Z(n40924) );
  NANDN U41213 ( .A(n40926), .B(n40925), .Z(n40921) );
  ANDN U41214 ( .B(B[145]), .A(n80), .Z(n40705) );
  XNOR U41215 ( .A(n40713), .B(n40927), .Z(n40706) );
  XNOR U41216 ( .A(n40712), .B(n40710), .Z(n40927) );
  AND U41217 ( .A(n40928), .B(n40929), .Z(n40710) );
  NANDN U41218 ( .A(n40930), .B(n40931), .Z(n40929) );
  OR U41219 ( .A(n40932), .B(n40933), .Z(n40931) );
  NAND U41220 ( .A(n40933), .B(n40932), .Z(n40928) );
  ANDN U41221 ( .B(B[146]), .A(n81), .Z(n40712) );
  XNOR U41222 ( .A(n40720), .B(n40934), .Z(n40713) );
  XNOR U41223 ( .A(n40719), .B(n40717), .Z(n40934) );
  AND U41224 ( .A(n40935), .B(n40936), .Z(n40717) );
  NANDN U41225 ( .A(n40937), .B(n40938), .Z(n40936) );
  NAND U41226 ( .A(n40939), .B(n40940), .Z(n40938) );
  ANDN U41227 ( .B(B[147]), .A(n82), .Z(n40719) );
  XOR U41228 ( .A(n40726), .B(n40941), .Z(n40720) );
  XNOR U41229 ( .A(n40724), .B(n40727), .Z(n40941) );
  NAND U41230 ( .A(A[2]), .B(B[148]), .Z(n40727) );
  NANDN U41231 ( .A(n40942), .B(n40943), .Z(n40724) );
  AND U41232 ( .A(A[0]), .B(B[149]), .Z(n40943) );
  XNOR U41233 ( .A(n40729), .B(n40944), .Z(n40726) );
  NAND U41234 ( .A(A[0]), .B(B[150]), .Z(n40944) );
  NAND U41235 ( .A(B[149]), .B(A[1]), .Z(n40729) );
  NAND U41236 ( .A(n40945), .B(n40946), .Z(n496) );
  NANDN U41237 ( .A(n40947), .B(n40948), .Z(n40946) );
  OR U41238 ( .A(n40949), .B(n40950), .Z(n40948) );
  NAND U41239 ( .A(n40950), .B(n40949), .Z(n40945) );
  XOR U41240 ( .A(n498), .B(n497), .Z(\A1[147] ) );
  XOR U41241 ( .A(n40950), .B(n40951), .Z(n497) );
  XNOR U41242 ( .A(n40949), .B(n40947), .Z(n40951) );
  AND U41243 ( .A(n40952), .B(n40953), .Z(n40947) );
  NANDN U41244 ( .A(n40954), .B(n40955), .Z(n40953) );
  NANDN U41245 ( .A(n40956), .B(n40957), .Z(n40955) );
  NANDN U41246 ( .A(n40957), .B(n40956), .Z(n40952) );
  ANDN U41247 ( .B(B[118]), .A(n54), .Z(n40949) );
  XNOR U41248 ( .A(n40744), .B(n40958), .Z(n40950) );
  XNOR U41249 ( .A(n40743), .B(n40741), .Z(n40958) );
  AND U41250 ( .A(n40959), .B(n40960), .Z(n40741) );
  NANDN U41251 ( .A(n40961), .B(n40962), .Z(n40960) );
  OR U41252 ( .A(n40963), .B(n40964), .Z(n40962) );
  NAND U41253 ( .A(n40964), .B(n40963), .Z(n40959) );
  ANDN U41254 ( .B(B[119]), .A(n55), .Z(n40743) );
  XNOR U41255 ( .A(n40751), .B(n40965), .Z(n40744) );
  XNOR U41256 ( .A(n40750), .B(n40748), .Z(n40965) );
  AND U41257 ( .A(n40966), .B(n40967), .Z(n40748) );
  NANDN U41258 ( .A(n40968), .B(n40969), .Z(n40967) );
  NANDN U41259 ( .A(n40970), .B(n40971), .Z(n40969) );
  NANDN U41260 ( .A(n40971), .B(n40970), .Z(n40966) );
  ANDN U41261 ( .B(B[120]), .A(n56), .Z(n40750) );
  XNOR U41262 ( .A(n40758), .B(n40972), .Z(n40751) );
  XNOR U41263 ( .A(n40757), .B(n40755), .Z(n40972) );
  AND U41264 ( .A(n40973), .B(n40974), .Z(n40755) );
  NANDN U41265 ( .A(n40975), .B(n40976), .Z(n40974) );
  OR U41266 ( .A(n40977), .B(n40978), .Z(n40976) );
  NAND U41267 ( .A(n40978), .B(n40977), .Z(n40973) );
  ANDN U41268 ( .B(B[121]), .A(n57), .Z(n40757) );
  XNOR U41269 ( .A(n40765), .B(n40979), .Z(n40758) );
  XNOR U41270 ( .A(n40764), .B(n40762), .Z(n40979) );
  AND U41271 ( .A(n40980), .B(n40981), .Z(n40762) );
  NANDN U41272 ( .A(n40982), .B(n40983), .Z(n40981) );
  NANDN U41273 ( .A(n40984), .B(n40985), .Z(n40983) );
  NANDN U41274 ( .A(n40985), .B(n40984), .Z(n40980) );
  ANDN U41275 ( .B(B[122]), .A(n58), .Z(n40764) );
  XNOR U41276 ( .A(n40772), .B(n40986), .Z(n40765) );
  XNOR U41277 ( .A(n40771), .B(n40769), .Z(n40986) );
  AND U41278 ( .A(n40987), .B(n40988), .Z(n40769) );
  NANDN U41279 ( .A(n40989), .B(n40990), .Z(n40988) );
  OR U41280 ( .A(n40991), .B(n40992), .Z(n40990) );
  NAND U41281 ( .A(n40992), .B(n40991), .Z(n40987) );
  ANDN U41282 ( .B(B[123]), .A(n59), .Z(n40771) );
  XNOR U41283 ( .A(n40779), .B(n40993), .Z(n40772) );
  XNOR U41284 ( .A(n40778), .B(n40776), .Z(n40993) );
  AND U41285 ( .A(n40994), .B(n40995), .Z(n40776) );
  NANDN U41286 ( .A(n40996), .B(n40997), .Z(n40995) );
  NANDN U41287 ( .A(n40998), .B(n40999), .Z(n40997) );
  NANDN U41288 ( .A(n40999), .B(n40998), .Z(n40994) );
  ANDN U41289 ( .B(B[124]), .A(n60), .Z(n40778) );
  XNOR U41290 ( .A(n40786), .B(n41000), .Z(n40779) );
  XNOR U41291 ( .A(n40785), .B(n40783), .Z(n41000) );
  AND U41292 ( .A(n41001), .B(n41002), .Z(n40783) );
  NANDN U41293 ( .A(n41003), .B(n41004), .Z(n41002) );
  OR U41294 ( .A(n41005), .B(n41006), .Z(n41004) );
  NAND U41295 ( .A(n41006), .B(n41005), .Z(n41001) );
  ANDN U41296 ( .B(B[125]), .A(n61), .Z(n40785) );
  XNOR U41297 ( .A(n40793), .B(n41007), .Z(n40786) );
  XNOR U41298 ( .A(n40792), .B(n40790), .Z(n41007) );
  AND U41299 ( .A(n41008), .B(n41009), .Z(n40790) );
  NANDN U41300 ( .A(n41010), .B(n41011), .Z(n41009) );
  NANDN U41301 ( .A(n41012), .B(n41013), .Z(n41011) );
  NANDN U41302 ( .A(n41013), .B(n41012), .Z(n41008) );
  ANDN U41303 ( .B(B[126]), .A(n62), .Z(n40792) );
  XNOR U41304 ( .A(n40800), .B(n41014), .Z(n40793) );
  XNOR U41305 ( .A(n40799), .B(n40797), .Z(n41014) );
  AND U41306 ( .A(n41015), .B(n41016), .Z(n40797) );
  NANDN U41307 ( .A(n41017), .B(n41018), .Z(n41016) );
  OR U41308 ( .A(n41019), .B(n41020), .Z(n41018) );
  NAND U41309 ( .A(n41020), .B(n41019), .Z(n41015) );
  ANDN U41310 ( .B(B[127]), .A(n63), .Z(n40799) );
  XNOR U41311 ( .A(n40807), .B(n41021), .Z(n40800) );
  XNOR U41312 ( .A(n40806), .B(n40804), .Z(n41021) );
  AND U41313 ( .A(n41022), .B(n41023), .Z(n40804) );
  NANDN U41314 ( .A(n41024), .B(n41025), .Z(n41023) );
  NANDN U41315 ( .A(n41026), .B(n41027), .Z(n41025) );
  NANDN U41316 ( .A(n41027), .B(n41026), .Z(n41022) );
  ANDN U41317 ( .B(B[128]), .A(n64), .Z(n40806) );
  XNOR U41318 ( .A(n40814), .B(n41028), .Z(n40807) );
  XNOR U41319 ( .A(n40813), .B(n40811), .Z(n41028) );
  AND U41320 ( .A(n41029), .B(n41030), .Z(n40811) );
  NANDN U41321 ( .A(n41031), .B(n41032), .Z(n41030) );
  OR U41322 ( .A(n41033), .B(n41034), .Z(n41032) );
  NAND U41323 ( .A(n41034), .B(n41033), .Z(n41029) );
  ANDN U41324 ( .B(B[129]), .A(n65), .Z(n40813) );
  XNOR U41325 ( .A(n40821), .B(n41035), .Z(n40814) );
  XNOR U41326 ( .A(n40820), .B(n40818), .Z(n41035) );
  AND U41327 ( .A(n41036), .B(n41037), .Z(n40818) );
  NANDN U41328 ( .A(n41038), .B(n41039), .Z(n41037) );
  NANDN U41329 ( .A(n41040), .B(n41041), .Z(n41039) );
  NANDN U41330 ( .A(n41041), .B(n41040), .Z(n41036) );
  ANDN U41331 ( .B(B[130]), .A(n66), .Z(n40820) );
  XNOR U41332 ( .A(n40828), .B(n41042), .Z(n40821) );
  XNOR U41333 ( .A(n40827), .B(n40825), .Z(n41042) );
  AND U41334 ( .A(n41043), .B(n41044), .Z(n40825) );
  NANDN U41335 ( .A(n41045), .B(n41046), .Z(n41044) );
  OR U41336 ( .A(n41047), .B(n41048), .Z(n41046) );
  NAND U41337 ( .A(n41048), .B(n41047), .Z(n41043) );
  ANDN U41338 ( .B(B[131]), .A(n67), .Z(n40827) );
  XNOR U41339 ( .A(n40835), .B(n41049), .Z(n40828) );
  XNOR U41340 ( .A(n40834), .B(n40832), .Z(n41049) );
  AND U41341 ( .A(n41050), .B(n41051), .Z(n40832) );
  NANDN U41342 ( .A(n41052), .B(n41053), .Z(n41051) );
  NANDN U41343 ( .A(n41054), .B(n41055), .Z(n41053) );
  NANDN U41344 ( .A(n41055), .B(n41054), .Z(n41050) );
  ANDN U41345 ( .B(B[132]), .A(n68), .Z(n40834) );
  XNOR U41346 ( .A(n40842), .B(n41056), .Z(n40835) );
  XNOR U41347 ( .A(n40841), .B(n40839), .Z(n41056) );
  AND U41348 ( .A(n41057), .B(n41058), .Z(n40839) );
  NANDN U41349 ( .A(n41059), .B(n41060), .Z(n41058) );
  OR U41350 ( .A(n41061), .B(n41062), .Z(n41060) );
  NAND U41351 ( .A(n41062), .B(n41061), .Z(n41057) );
  ANDN U41352 ( .B(B[133]), .A(n69), .Z(n40841) );
  XNOR U41353 ( .A(n40849), .B(n41063), .Z(n40842) );
  XNOR U41354 ( .A(n40848), .B(n40846), .Z(n41063) );
  AND U41355 ( .A(n41064), .B(n41065), .Z(n40846) );
  NANDN U41356 ( .A(n41066), .B(n41067), .Z(n41065) );
  NANDN U41357 ( .A(n41068), .B(n41069), .Z(n41067) );
  NANDN U41358 ( .A(n41069), .B(n41068), .Z(n41064) );
  ANDN U41359 ( .B(B[134]), .A(n70), .Z(n40848) );
  XNOR U41360 ( .A(n40856), .B(n41070), .Z(n40849) );
  XNOR U41361 ( .A(n40855), .B(n40853), .Z(n41070) );
  AND U41362 ( .A(n41071), .B(n41072), .Z(n40853) );
  NANDN U41363 ( .A(n41073), .B(n41074), .Z(n41072) );
  OR U41364 ( .A(n41075), .B(n41076), .Z(n41074) );
  NAND U41365 ( .A(n41076), .B(n41075), .Z(n41071) );
  ANDN U41366 ( .B(B[135]), .A(n71), .Z(n40855) );
  XNOR U41367 ( .A(n40863), .B(n41077), .Z(n40856) );
  XNOR U41368 ( .A(n40862), .B(n40860), .Z(n41077) );
  AND U41369 ( .A(n41078), .B(n41079), .Z(n40860) );
  NANDN U41370 ( .A(n41080), .B(n41081), .Z(n41079) );
  NANDN U41371 ( .A(n41082), .B(n41083), .Z(n41081) );
  NANDN U41372 ( .A(n41083), .B(n41082), .Z(n41078) );
  ANDN U41373 ( .B(B[136]), .A(n72), .Z(n40862) );
  XNOR U41374 ( .A(n40870), .B(n41084), .Z(n40863) );
  XNOR U41375 ( .A(n40869), .B(n40867), .Z(n41084) );
  AND U41376 ( .A(n41085), .B(n41086), .Z(n40867) );
  NANDN U41377 ( .A(n41087), .B(n41088), .Z(n41086) );
  OR U41378 ( .A(n41089), .B(n41090), .Z(n41088) );
  NAND U41379 ( .A(n41090), .B(n41089), .Z(n41085) );
  ANDN U41380 ( .B(B[137]), .A(n73), .Z(n40869) );
  XNOR U41381 ( .A(n40877), .B(n41091), .Z(n40870) );
  XNOR U41382 ( .A(n40876), .B(n40874), .Z(n41091) );
  AND U41383 ( .A(n41092), .B(n41093), .Z(n40874) );
  NANDN U41384 ( .A(n41094), .B(n41095), .Z(n41093) );
  NANDN U41385 ( .A(n41096), .B(n41097), .Z(n41095) );
  NANDN U41386 ( .A(n41097), .B(n41096), .Z(n41092) );
  ANDN U41387 ( .B(B[138]), .A(n74), .Z(n40876) );
  XNOR U41388 ( .A(n40884), .B(n41098), .Z(n40877) );
  XNOR U41389 ( .A(n40883), .B(n40881), .Z(n41098) );
  AND U41390 ( .A(n41099), .B(n41100), .Z(n40881) );
  NANDN U41391 ( .A(n41101), .B(n41102), .Z(n41100) );
  OR U41392 ( .A(n41103), .B(n41104), .Z(n41102) );
  NAND U41393 ( .A(n41104), .B(n41103), .Z(n41099) );
  ANDN U41394 ( .B(B[139]), .A(n75), .Z(n40883) );
  XNOR U41395 ( .A(n40891), .B(n41105), .Z(n40884) );
  XNOR U41396 ( .A(n40890), .B(n40888), .Z(n41105) );
  AND U41397 ( .A(n41106), .B(n41107), .Z(n40888) );
  NANDN U41398 ( .A(n41108), .B(n41109), .Z(n41107) );
  NANDN U41399 ( .A(n41110), .B(n41111), .Z(n41109) );
  NANDN U41400 ( .A(n41111), .B(n41110), .Z(n41106) );
  ANDN U41401 ( .B(B[140]), .A(n76), .Z(n40890) );
  XNOR U41402 ( .A(n40898), .B(n41112), .Z(n40891) );
  XNOR U41403 ( .A(n40897), .B(n40895), .Z(n41112) );
  AND U41404 ( .A(n41113), .B(n41114), .Z(n40895) );
  NANDN U41405 ( .A(n41115), .B(n41116), .Z(n41114) );
  OR U41406 ( .A(n41117), .B(n41118), .Z(n41116) );
  NAND U41407 ( .A(n41118), .B(n41117), .Z(n41113) );
  ANDN U41408 ( .B(B[141]), .A(n77), .Z(n40897) );
  XNOR U41409 ( .A(n40905), .B(n41119), .Z(n40898) );
  XNOR U41410 ( .A(n40904), .B(n40902), .Z(n41119) );
  AND U41411 ( .A(n41120), .B(n41121), .Z(n40902) );
  NANDN U41412 ( .A(n41122), .B(n41123), .Z(n41121) );
  NANDN U41413 ( .A(n41124), .B(n41125), .Z(n41123) );
  NANDN U41414 ( .A(n41125), .B(n41124), .Z(n41120) );
  ANDN U41415 ( .B(B[142]), .A(n78), .Z(n40904) );
  XNOR U41416 ( .A(n40912), .B(n41126), .Z(n40905) );
  XNOR U41417 ( .A(n40911), .B(n40909), .Z(n41126) );
  AND U41418 ( .A(n41127), .B(n41128), .Z(n40909) );
  NANDN U41419 ( .A(n41129), .B(n41130), .Z(n41128) );
  OR U41420 ( .A(n41131), .B(n41132), .Z(n41130) );
  NAND U41421 ( .A(n41132), .B(n41131), .Z(n41127) );
  ANDN U41422 ( .B(B[143]), .A(n79), .Z(n40911) );
  XNOR U41423 ( .A(n40919), .B(n41133), .Z(n40912) );
  XNOR U41424 ( .A(n40918), .B(n40916), .Z(n41133) );
  AND U41425 ( .A(n41134), .B(n41135), .Z(n40916) );
  NANDN U41426 ( .A(n41136), .B(n41137), .Z(n41135) );
  NANDN U41427 ( .A(n41138), .B(n41139), .Z(n41137) );
  NANDN U41428 ( .A(n41139), .B(n41138), .Z(n41134) );
  ANDN U41429 ( .B(B[144]), .A(n80), .Z(n40918) );
  XNOR U41430 ( .A(n40926), .B(n41140), .Z(n40919) );
  XNOR U41431 ( .A(n40925), .B(n40923), .Z(n41140) );
  AND U41432 ( .A(n41141), .B(n41142), .Z(n40923) );
  NANDN U41433 ( .A(n41143), .B(n41144), .Z(n41142) );
  OR U41434 ( .A(n41145), .B(n41146), .Z(n41144) );
  NAND U41435 ( .A(n41146), .B(n41145), .Z(n41141) );
  ANDN U41436 ( .B(B[145]), .A(n81), .Z(n40925) );
  XNOR U41437 ( .A(n40933), .B(n41147), .Z(n40926) );
  XNOR U41438 ( .A(n40932), .B(n40930), .Z(n41147) );
  AND U41439 ( .A(n41148), .B(n41149), .Z(n40930) );
  NANDN U41440 ( .A(n41150), .B(n41151), .Z(n41149) );
  NAND U41441 ( .A(n41152), .B(n41153), .Z(n41151) );
  ANDN U41442 ( .B(B[146]), .A(n82), .Z(n40932) );
  XOR U41443 ( .A(n40939), .B(n41154), .Z(n40933) );
  XNOR U41444 ( .A(n40937), .B(n40940), .Z(n41154) );
  NAND U41445 ( .A(A[2]), .B(B[147]), .Z(n40940) );
  NANDN U41446 ( .A(n41155), .B(n41156), .Z(n40937) );
  AND U41447 ( .A(A[0]), .B(B[148]), .Z(n41156) );
  XNOR U41448 ( .A(n40942), .B(n41157), .Z(n40939) );
  NAND U41449 ( .A(A[0]), .B(B[149]), .Z(n41157) );
  NAND U41450 ( .A(B[148]), .B(A[1]), .Z(n40942) );
  NAND U41451 ( .A(n41158), .B(n41159), .Z(n498) );
  NANDN U41452 ( .A(n41160), .B(n41161), .Z(n41159) );
  OR U41453 ( .A(n41162), .B(n41163), .Z(n41161) );
  NAND U41454 ( .A(n41163), .B(n41162), .Z(n41158) );
  XOR U41455 ( .A(n500), .B(n499), .Z(\A1[146] ) );
  XOR U41456 ( .A(n41163), .B(n41164), .Z(n499) );
  XNOR U41457 ( .A(n41162), .B(n41160), .Z(n41164) );
  AND U41458 ( .A(n41165), .B(n41166), .Z(n41160) );
  NANDN U41459 ( .A(n41167), .B(n41168), .Z(n41166) );
  NANDN U41460 ( .A(n41169), .B(n41170), .Z(n41168) );
  NANDN U41461 ( .A(n41170), .B(n41169), .Z(n41165) );
  ANDN U41462 ( .B(B[117]), .A(n54), .Z(n41162) );
  XNOR U41463 ( .A(n40957), .B(n41171), .Z(n41163) );
  XNOR U41464 ( .A(n40956), .B(n40954), .Z(n41171) );
  AND U41465 ( .A(n41172), .B(n41173), .Z(n40954) );
  NANDN U41466 ( .A(n41174), .B(n41175), .Z(n41173) );
  OR U41467 ( .A(n41176), .B(n41177), .Z(n41175) );
  NAND U41468 ( .A(n41177), .B(n41176), .Z(n41172) );
  ANDN U41469 ( .B(B[118]), .A(n55), .Z(n40956) );
  XNOR U41470 ( .A(n40964), .B(n41178), .Z(n40957) );
  XNOR U41471 ( .A(n40963), .B(n40961), .Z(n41178) );
  AND U41472 ( .A(n41179), .B(n41180), .Z(n40961) );
  NANDN U41473 ( .A(n41181), .B(n41182), .Z(n41180) );
  NANDN U41474 ( .A(n41183), .B(n41184), .Z(n41182) );
  NANDN U41475 ( .A(n41184), .B(n41183), .Z(n41179) );
  ANDN U41476 ( .B(B[119]), .A(n56), .Z(n40963) );
  XNOR U41477 ( .A(n40971), .B(n41185), .Z(n40964) );
  XNOR U41478 ( .A(n40970), .B(n40968), .Z(n41185) );
  AND U41479 ( .A(n41186), .B(n41187), .Z(n40968) );
  NANDN U41480 ( .A(n41188), .B(n41189), .Z(n41187) );
  OR U41481 ( .A(n41190), .B(n41191), .Z(n41189) );
  NAND U41482 ( .A(n41191), .B(n41190), .Z(n41186) );
  ANDN U41483 ( .B(B[120]), .A(n57), .Z(n40970) );
  XNOR U41484 ( .A(n40978), .B(n41192), .Z(n40971) );
  XNOR U41485 ( .A(n40977), .B(n40975), .Z(n41192) );
  AND U41486 ( .A(n41193), .B(n41194), .Z(n40975) );
  NANDN U41487 ( .A(n41195), .B(n41196), .Z(n41194) );
  NANDN U41488 ( .A(n41197), .B(n41198), .Z(n41196) );
  NANDN U41489 ( .A(n41198), .B(n41197), .Z(n41193) );
  ANDN U41490 ( .B(B[121]), .A(n58), .Z(n40977) );
  XNOR U41491 ( .A(n40985), .B(n41199), .Z(n40978) );
  XNOR U41492 ( .A(n40984), .B(n40982), .Z(n41199) );
  AND U41493 ( .A(n41200), .B(n41201), .Z(n40982) );
  NANDN U41494 ( .A(n41202), .B(n41203), .Z(n41201) );
  OR U41495 ( .A(n41204), .B(n41205), .Z(n41203) );
  NAND U41496 ( .A(n41205), .B(n41204), .Z(n41200) );
  ANDN U41497 ( .B(B[122]), .A(n59), .Z(n40984) );
  XNOR U41498 ( .A(n40992), .B(n41206), .Z(n40985) );
  XNOR U41499 ( .A(n40991), .B(n40989), .Z(n41206) );
  AND U41500 ( .A(n41207), .B(n41208), .Z(n40989) );
  NANDN U41501 ( .A(n41209), .B(n41210), .Z(n41208) );
  NANDN U41502 ( .A(n41211), .B(n41212), .Z(n41210) );
  NANDN U41503 ( .A(n41212), .B(n41211), .Z(n41207) );
  ANDN U41504 ( .B(B[123]), .A(n60), .Z(n40991) );
  XNOR U41505 ( .A(n40999), .B(n41213), .Z(n40992) );
  XNOR U41506 ( .A(n40998), .B(n40996), .Z(n41213) );
  AND U41507 ( .A(n41214), .B(n41215), .Z(n40996) );
  NANDN U41508 ( .A(n41216), .B(n41217), .Z(n41215) );
  OR U41509 ( .A(n41218), .B(n41219), .Z(n41217) );
  NAND U41510 ( .A(n41219), .B(n41218), .Z(n41214) );
  ANDN U41511 ( .B(B[124]), .A(n61), .Z(n40998) );
  XNOR U41512 ( .A(n41006), .B(n41220), .Z(n40999) );
  XNOR U41513 ( .A(n41005), .B(n41003), .Z(n41220) );
  AND U41514 ( .A(n41221), .B(n41222), .Z(n41003) );
  NANDN U41515 ( .A(n41223), .B(n41224), .Z(n41222) );
  NANDN U41516 ( .A(n41225), .B(n41226), .Z(n41224) );
  NANDN U41517 ( .A(n41226), .B(n41225), .Z(n41221) );
  ANDN U41518 ( .B(B[125]), .A(n62), .Z(n41005) );
  XNOR U41519 ( .A(n41013), .B(n41227), .Z(n41006) );
  XNOR U41520 ( .A(n41012), .B(n41010), .Z(n41227) );
  AND U41521 ( .A(n41228), .B(n41229), .Z(n41010) );
  NANDN U41522 ( .A(n41230), .B(n41231), .Z(n41229) );
  OR U41523 ( .A(n41232), .B(n41233), .Z(n41231) );
  NAND U41524 ( .A(n41233), .B(n41232), .Z(n41228) );
  ANDN U41525 ( .B(B[126]), .A(n63), .Z(n41012) );
  XNOR U41526 ( .A(n41020), .B(n41234), .Z(n41013) );
  XNOR U41527 ( .A(n41019), .B(n41017), .Z(n41234) );
  AND U41528 ( .A(n41235), .B(n41236), .Z(n41017) );
  NANDN U41529 ( .A(n41237), .B(n41238), .Z(n41236) );
  NANDN U41530 ( .A(n41239), .B(n41240), .Z(n41238) );
  NANDN U41531 ( .A(n41240), .B(n41239), .Z(n41235) );
  ANDN U41532 ( .B(B[127]), .A(n64), .Z(n41019) );
  XNOR U41533 ( .A(n41027), .B(n41241), .Z(n41020) );
  XNOR U41534 ( .A(n41026), .B(n41024), .Z(n41241) );
  AND U41535 ( .A(n41242), .B(n41243), .Z(n41024) );
  NANDN U41536 ( .A(n41244), .B(n41245), .Z(n41243) );
  OR U41537 ( .A(n41246), .B(n41247), .Z(n41245) );
  NAND U41538 ( .A(n41247), .B(n41246), .Z(n41242) );
  ANDN U41539 ( .B(B[128]), .A(n65), .Z(n41026) );
  XNOR U41540 ( .A(n41034), .B(n41248), .Z(n41027) );
  XNOR U41541 ( .A(n41033), .B(n41031), .Z(n41248) );
  AND U41542 ( .A(n41249), .B(n41250), .Z(n41031) );
  NANDN U41543 ( .A(n41251), .B(n41252), .Z(n41250) );
  NANDN U41544 ( .A(n41253), .B(n41254), .Z(n41252) );
  NANDN U41545 ( .A(n41254), .B(n41253), .Z(n41249) );
  ANDN U41546 ( .B(B[129]), .A(n66), .Z(n41033) );
  XNOR U41547 ( .A(n41041), .B(n41255), .Z(n41034) );
  XNOR U41548 ( .A(n41040), .B(n41038), .Z(n41255) );
  AND U41549 ( .A(n41256), .B(n41257), .Z(n41038) );
  NANDN U41550 ( .A(n41258), .B(n41259), .Z(n41257) );
  OR U41551 ( .A(n41260), .B(n41261), .Z(n41259) );
  NAND U41552 ( .A(n41261), .B(n41260), .Z(n41256) );
  ANDN U41553 ( .B(B[130]), .A(n67), .Z(n41040) );
  XNOR U41554 ( .A(n41048), .B(n41262), .Z(n41041) );
  XNOR U41555 ( .A(n41047), .B(n41045), .Z(n41262) );
  AND U41556 ( .A(n41263), .B(n41264), .Z(n41045) );
  NANDN U41557 ( .A(n41265), .B(n41266), .Z(n41264) );
  NANDN U41558 ( .A(n41267), .B(n41268), .Z(n41266) );
  NANDN U41559 ( .A(n41268), .B(n41267), .Z(n41263) );
  ANDN U41560 ( .B(B[131]), .A(n68), .Z(n41047) );
  XNOR U41561 ( .A(n41055), .B(n41269), .Z(n41048) );
  XNOR U41562 ( .A(n41054), .B(n41052), .Z(n41269) );
  AND U41563 ( .A(n41270), .B(n41271), .Z(n41052) );
  NANDN U41564 ( .A(n41272), .B(n41273), .Z(n41271) );
  OR U41565 ( .A(n41274), .B(n41275), .Z(n41273) );
  NAND U41566 ( .A(n41275), .B(n41274), .Z(n41270) );
  ANDN U41567 ( .B(B[132]), .A(n69), .Z(n41054) );
  XNOR U41568 ( .A(n41062), .B(n41276), .Z(n41055) );
  XNOR U41569 ( .A(n41061), .B(n41059), .Z(n41276) );
  AND U41570 ( .A(n41277), .B(n41278), .Z(n41059) );
  NANDN U41571 ( .A(n41279), .B(n41280), .Z(n41278) );
  NANDN U41572 ( .A(n41281), .B(n41282), .Z(n41280) );
  NANDN U41573 ( .A(n41282), .B(n41281), .Z(n41277) );
  ANDN U41574 ( .B(B[133]), .A(n70), .Z(n41061) );
  XNOR U41575 ( .A(n41069), .B(n41283), .Z(n41062) );
  XNOR U41576 ( .A(n41068), .B(n41066), .Z(n41283) );
  AND U41577 ( .A(n41284), .B(n41285), .Z(n41066) );
  NANDN U41578 ( .A(n41286), .B(n41287), .Z(n41285) );
  OR U41579 ( .A(n41288), .B(n41289), .Z(n41287) );
  NAND U41580 ( .A(n41289), .B(n41288), .Z(n41284) );
  ANDN U41581 ( .B(B[134]), .A(n71), .Z(n41068) );
  XNOR U41582 ( .A(n41076), .B(n41290), .Z(n41069) );
  XNOR U41583 ( .A(n41075), .B(n41073), .Z(n41290) );
  AND U41584 ( .A(n41291), .B(n41292), .Z(n41073) );
  NANDN U41585 ( .A(n41293), .B(n41294), .Z(n41292) );
  NANDN U41586 ( .A(n41295), .B(n41296), .Z(n41294) );
  NANDN U41587 ( .A(n41296), .B(n41295), .Z(n41291) );
  ANDN U41588 ( .B(B[135]), .A(n72), .Z(n41075) );
  XNOR U41589 ( .A(n41083), .B(n41297), .Z(n41076) );
  XNOR U41590 ( .A(n41082), .B(n41080), .Z(n41297) );
  AND U41591 ( .A(n41298), .B(n41299), .Z(n41080) );
  NANDN U41592 ( .A(n41300), .B(n41301), .Z(n41299) );
  OR U41593 ( .A(n41302), .B(n41303), .Z(n41301) );
  NAND U41594 ( .A(n41303), .B(n41302), .Z(n41298) );
  ANDN U41595 ( .B(B[136]), .A(n73), .Z(n41082) );
  XNOR U41596 ( .A(n41090), .B(n41304), .Z(n41083) );
  XNOR U41597 ( .A(n41089), .B(n41087), .Z(n41304) );
  AND U41598 ( .A(n41305), .B(n41306), .Z(n41087) );
  NANDN U41599 ( .A(n41307), .B(n41308), .Z(n41306) );
  NANDN U41600 ( .A(n41309), .B(n41310), .Z(n41308) );
  NANDN U41601 ( .A(n41310), .B(n41309), .Z(n41305) );
  ANDN U41602 ( .B(B[137]), .A(n74), .Z(n41089) );
  XNOR U41603 ( .A(n41097), .B(n41311), .Z(n41090) );
  XNOR U41604 ( .A(n41096), .B(n41094), .Z(n41311) );
  AND U41605 ( .A(n41312), .B(n41313), .Z(n41094) );
  NANDN U41606 ( .A(n41314), .B(n41315), .Z(n41313) );
  OR U41607 ( .A(n41316), .B(n41317), .Z(n41315) );
  NAND U41608 ( .A(n41317), .B(n41316), .Z(n41312) );
  ANDN U41609 ( .B(B[138]), .A(n75), .Z(n41096) );
  XNOR U41610 ( .A(n41104), .B(n41318), .Z(n41097) );
  XNOR U41611 ( .A(n41103), .B(n41101), .Z(n41318) );
  AND U41612 ( .A(n41319), .B(n41320), .Z(n41101) );
  NANDN U41613 ( .A(n41321), .B(n41322), .Z(n41320) );
  NANDN U41614 ( .A(n41323), .B(n41324), .Z(n41322) );
  NANDN U41615 ( .A(n41324), .B(n41323), .Z(n41319) );
  ANDN U41616 ( .B(B[139]), .A(n76), .Z(n41103) );
  XNOR U41617 ( .A(n41111), .B(n41325), .Z(n41104) );
  XNOR U41618 ( .A(n41110), .B(n41108), .Z(n41325) );
  AND U41619 ( .A(n41326), .B(n41327), .Z(n41108) );
  NANDN U41620 ( .A(n41328), .B(n41329), .Z(n41327) );
  OR U41621 ( .A(n41330), .B(n41331), .Z(n41329) );
  NAND U41622 ( .A(n41331), .B(n41330), .Z(n41326) );
  ANDN U41623 ( .B(B[140]), .A(n77), .Z(n41110) );
  XNOR U41624 ( .A(n41118), .B(n41332), .Z(n41111) );
  XNOR U41625 ( .A(n41117), .B(n41115), .Z(n41332) );
  AND U41626 ( .A(n41333), .B(n41334), .Z(n41115) );
  NANDN U41627 ( .A(n41335), .B(n41336), .Z(n41334) );
  NANDN U41628 ( .A(n41337), .B(n41338), .Z(n41336) );
  NANDN U41629 ( .A(n41338), .B(n41337), .Z(n41333) );
  ANDN U41630 ( .B(B[141]), .A(n78), .Z(n41117) );
  XNOR U41631 ( .A(n41125), .B(n41339), .Z(n41118) );
  XNOR U41632 ( .A(n41124), .B(n41122), .Z(n41339) );
  AND U41633 ( .A(n41340), .B(n41341), .Z(n41122) );
  NANDN U41634 ( .A(n41342), .B(n41343), .Z(n41341) );
  OR U41635 ( .A(n41344), .B(n41345), .Z(n41343) );
  NAND U41636 ( .A(n41345), .B(n41344), .Z(n41340) );
  ANDN U41637 ( .B(B[142]), .A(n79), .Z(n41124) );
  XNOR U41638 ( .A(n41132), .B(n41346), .Z(n41125) );
  XNOR U41639 ( .A(n41131), .B(n41129), .Z(n41346) );
  AND U41640 ( .A(n41347), .B(n41348), .Z(n41129) );
  NANDN U41641 ( .A(n41349), .B(n41350), .Z(n41348) );
  NANDN U41642 ( .A(n41351), .B(n41352), .Z(n41350) );
  NANDN U41643 ( .A(n41352), .B(n41351), .Z(n41347) );
  ANDN U41644 ( .B(B[143]), .A(n80), .Z(n41131) );
  XNOR U41645 ( .A(n41139), .B(n41353), .Z(n41132) );
  XNOR U41646 ( .A(n41138), .B(n41136), .Z(n41353) );
  AND U41647 ( .A(n41354), .B(n41355), .Z(n41136) );
  NANDN U41648 ( .A(n41356), .B(n41357), .Z(n41355) );
  OR U41649 ( .A(n41358), .B(n41359), .Z(n41357) );
  NAND U41650 ( .A(n41359), .B(n41358), .Z(n41354) );
  ANDN U41651 ( .B(B[144]), .A(n81), .Z(n41138) );
  XNOR U41652 ( .A(n41146), .B(n41360), .Z(n41139) );
  XNOR U41653 ( .A(n41145), .B(n41143), .Z(n41360) );
  AND U41654 ( .A(n41361), .B(n41362), .Z(n41143) );
  NANDN U41655 ( .A(n41363), .B(n41364), .Z(n41362) );
  NAND U41656 ( .A(n41365), .B(n41366), .Z(n41364) );
  ANDN U41657 ( .B(B[145]), .A(n82), .Z(n41145) );
  XOR U41658 ( .A(n41152), .B(n41367), .Z(n41146) );
  XNOR U41659 ( .A(n41150), .B(n41153), .Z(n41367) );
  NAND U41660 ( .A(A[2]), .B(B[146]), .Z(n41153) );
  NANDN U41661 ( .A(n41368), .B(n41369), .Z(n41150) );
  AND U41662 ( .A(A[0]), .B(B[147]), .Z(n41369) );
  XNOR U41663 ( .A(n41155), .B(n41370), .Z(n41152) );
  NAND U41664 ( .A(A[0]), .B(B[148]), .Z(n41370) );
  NAND U41665 ( .A(B[147]), .B(A[1]), .Z(n41155) );
  NAND U41666 ( .A(n41371), .B(n41372), .Z(n500) );
  NANDN U41667 ( .A(n41373), .B(n41374), .Z(n41372) );
  OR U41668 ( .A(n41375), .B(n41376), .Z(n41374) );
  NAND U41669 ( .A(n41376), .B(n41375), .Z(n41371) );
  XOR U41670 ( .A(n502), .B(n501), .Z(\A1[145] ) );
  XOR U41671 ( .A(n41376), .B(n41377), .Z(n501) );
  XNOR U41672 ( .A(n41375), .B(n41373), .Z(n41377) );
  AND U41673 ( .A(n41378), .B(n41379), .Z(n41373) );
  NANDN U41674 ( .A(n41380), .B(n41381), .Z(n41379) );
  NANDN U41675 ( .A(n41382), .B(n41383), .Z(n41381) );
  NANDN U41676 ( .A(n41383), .B(n41382), .Z(n41378) );
  ANDN U41677 ( .B(B[116]), .A(n54), .Z(n41375) );
  XNOR U41678 ( .A(n41170), .B(n41384), .Z(n41376) );
  XNOR U41679 ( .A(n41169), .B(n41167), .Z(n41384) );
  AND U41680 ( .A(n41385), .B(n41386), .Z(n41167) );
  NANDN U41681 ( .A(n41387), .B(n41388), .Z(n41386) );
  OR U41682 ( .A(n41389), .B(n41390), .Z(n41388) );
  NAND U41683 ( .A(n41390), .B(n41389), .Z(n41385) );
  ANDN U41684 ( .B(B[117]), .A(n55), .Z(n41169) );
  XNOR U41685 ( .A(n41177), .B(n41391), .Z(n41170) );
  XNOR U41686 ( .A(n41176), .B(n41174), .Z(n41391) );
  AND U41687 ( .A(n41392), .B(n41393), .Z(n41174) );
  NANDN U41688 ( .A(n41394), .B(n41395), .Z(n41393) );
  NANDN U41689 ( .A(n41396), .B(n41397), .Z(n41395) );
  NANDN U41690 ( .A(n41397), .B(n41396), .Z(n41392) );
  ANDN U41691 ( .B(B[118]), .A(n56), .Z(n41176) );
  XNOR U41692 ( .A(n41184), .B(n41398), .Z(n41177) );
  XNOR U41693 ( .A(n41183), .B(n41181), .Z(n41398) );
  AND U41694 ( .A(n41399), .B(n41400), .Z(n41181) );
  NANDN U41695 ( .A(n41401), .B(n41402), .Z(n41400) );
  OR U41696 ( .A(n41403), .B(n41404), .Z(n41402) );
  NAND U41697 ( .A(n41404), .B(n41403), .Z(n41399) );
  ANDN U41698 ( .B(B[119]), .A(n57), .Z(n41183) );
  XNOR U41699 ( .A(n41191), .B(n41405), .Z(n41184) );
  XNOR U41700 ( .A(n41190), .B(n41188), .Z(n41405) );
  AND U41701 ( .A(n41406), .B(n41407), .Z(n41188) );
  NANDN U41702 ( .A(n41408), .B(n41409), .Z(n41407) );
  NANDN U41703 ( .A(n41410), .B(n41411), .Z(n41409) );
  NANDN U41704 ( .A(n41411), .B(n41410), .Z(n41406) );
  ANDN U41705 ( .B(B[120]), .A(n58), .Z(n41190) );
  XNOR U41706 ( .A(n41198), .B(n41412), .Z(n41191) );
  XNOR U41707 ( .A(n41197), .B(n41195), .Z(n41412) );
  AND U41708 ( .A(n41413), .B(n41414), .Z(n41195) );
  NANDN U41709 ( .A(n41415), .B(n41416), .Z(n41414) );
  OR U41710 ( .A(n41417), .B(n41418), .Z(n41416) );
  NAND U41711 ( .A(n41418), .B(n41417), .Z(n41413) );
  ANDN U41712 ( .B(B[121]), .A(n59), .Z(n41197) );
  XNOR U41713 ( .A(n41205), .B(n41419), .Z(n41198) );
  XNOR U41714 ( .A(n41204), .B(n41202), .Z(n41419) );
  AND U41715 ( .A(n41420), .B(n41421), .Z(n41202) );
  NANDN U41716 ( .A(n41422), .B(n41423), .Z(n41421) );
  NANDN U41717 ( .A(n41424), .B(n41425), .Z(n41423) );
  NANDN U41718 ( .A(n41425), .B(n41424), .Z(n41420) );
  ANDN U41719 ( .B(B[122]), .A(n60), .Z(n41204) );
  XNOR U41720 ( .A(n41212), .B(n41426), .Z(n41205) );
  XNOR U41721 ( .A(n41211), .B(n41209), .Z(n41426) );
  AND U41722 ( .A(n41427), .B(n41428), .Z(n41209) );
  NANDN U41723 ( .A(n41429), .B(n41430), .Z(n41428) );
  OR U41724 ( .A(n41431), .B(n41432), .Z(n41430) );
  NAND U41725 ( .A(n41432), .B(n41431), .Z(n41427) );
  ANDN U41726 ( .B(B[123]), .A(n61), .Z(n41211) );
  XNOR U41727 ( .A(n41219), .B(n41433), .Z(n41212) );
  XNOR U41728 ( .A(n41218), .B(n41216), .Z(n41433) );
  AND U41729 ( .A(n41434), .B(n41435), .Z(n41216) );
  NANDN U41730 ( .A(n41436), .B(n41437), .Z(n41435) );
  NANDN U41731 ( .A(n41438), .B(n41439), .Z(n41437) );
  NANDN U41732 ( .A(n41439), .B(n41438), .Z(n41434) );
  ANDN U41733 ( .B(B[124]), .A(n62), .Z(n41218) );
  XNOR U41734 ( .A(n41226), .B(n41440), .Z(n41219) );
  XNOR U41735 ( .A(n41225), .B(n41223), .Z(n41440) );
  AND U41736 ( .A(n41441), .B(n41442), .Z(n41223) );
  NANDN U41737 ( .A(n41443), .B(n41444), .Z(n41442) );
  OR U41738 ( .A(n41445), .B(n41446), .Z(n41444) );
  NAND U41739 ( .A(n41446), .B(n41445), .Z(n41441) );
  ANDN U41740 ( .B(B[125]), .A(n63), .Z(n41225) );
  XNOR U41741 ( .A(n41233), .B(n41447), .Z(n41226) );
  XNOR U41742 ( .A(n41232), .B(n41230), .Z(n41447) );
  AND U41743 ( .A(n41448), .B(n41449), .Z(n41230) );
  NANDN U41744 ( .A(n41450), .B(n41451), .Z(n41449) );
  NANDN U41745 ( .A(n41452), .B(n41453), .Z(n41451) );
  NANDN U41746 ( .A(n41453), .B(n41452), .Z(n41448) );
  ANDN U41747 ( .B(B[126]), .A(n64), .Z(n41232) );
  XNOR U41748 ( .A(n41240), .B(n41454), .Z(n41233) );
  XNOR U41749 ( .A(n41239), .B(n41237), .Z(n41454) );
  AND U41750 ( .A(n41455), .B(n41456), .Z(n41237) );
  NANDN U41751 ( .A(n41457), .B(n41458), .Z(n41456) );
  OR U41752 ( .A(n41459), .B(n41460), .Z(n41458) );
  NAND U41753 ( .A(n41460), .B(n41459), .Z(n41455) );
  ANDN U41754 ( .B(B[127]), .A(n65), .Z(n41239) );
  XNOR U41755 ( .A(n41247), .B(n41461), .Z(n41240) );
  XNOR U41756 ( .A(n41246), .B(n41244), .Z(n41461) );
  AND U41757 ( .A(n41462), .B(n41463), .Z(n41244) );
  NANDN U41758 ( .A(n41464), .B(n41465), .Z(n41463) );
  NANDN U41759 ( .A(n41466), .B(n41467), .Z(n41465) );
  NANDN U41760 ( .A(n41467), .B(n41466), .Z(n41462) );
  ANDN U41761 ( .B(B[128]), .A(n66), .Z(n41246) );
  XNOR U41762 ( .A(n41254), .B(n41468), .Z(n41247) );
  XNOR U41763 ( .A(n41253), .B(n41251), .Z(n41468) );
  AND U41764 ( .A(n41469), .B(n41470), .Z(n41251) );
  NANDN U41765 ( .A(n41471), .B(n41472), .Z(n41470) );
  OR U41766 ( .A(n41473), .B(n41474), .Z(n41472) );
  NAND U41767 ( .A(n41474), .B(n41473), .Z(n41469) );
  ANDN U41768 ( .B(B[129]), .A(n67), .Z(n41253) );
  XNOR U41769 ( .A(n41261), .B(n41475), .Z(n41254) );
  XNOR U41770 ( .A(n41260), .B(n41258), .Z(n41475) );
  AND U41771 ( .A(n41476), .B(n41477), .Z(n41258) );
  NANDN U41772 ( .A(n41478), .B(n41479), .Z(n41477) );
  NANDN U41773 ( .A(n41480), .B(n41481), .Z(n41479) );
  NANDN U41774 ( .A(n41481), .B(n41480), .Z(n41476) );
  ANDN U41775 ( .B(B[130]), .A(n68), .Z(n41260) );
  XNOR U41776 ( .A(n41268), .B(n41482), .Z(n41261) );
  XNOR U41777 ( .A(n41267), .B(n41265), .Z(n41482) );
  AND U41778 ( .A(n41483), .B(n41484), .Z(n41265) );
  NANDN U41779 ( .A(n41485), .B(n41486), .Z(n41484) );
  OR U41780 ( .A(n41487), .B(n41488), .Z(n41486) );
  NAND U41781 ( .A(n41488), .B(n41487), .Z(n41483) );
  ANDN U41782 ( .B(B[131]), .A(n69), .Z(n41267) );
  XNOR U41783 ( .A(n41275), .B(n41489), .Z(n41268) );
  XNOR U41784 ( .A(n41274), .B(n41272), .Z(n41489) );
  AND U41785 ( .A(n41490), .B(n41491), .Z(n41272) );
  NANDN U41786 ( .A(n41492), .B(n41493), .Z(n41491) );
  NANDN U41787 ( .A(n41494), .B(n41495), .Z(n41493) );
  NANDN U41788 ( .A(n41495), .B(n41494), .Z(n41490) );
  ANDN U41789 ( .B(B[132]), .A(n70), .Z(n41274) );
  XNOR U41790 ( .A(n41282), .B(n41496), .Z(n41275) );
  XNOR U41791 ( .A(n41281), .B(n41279), .Z(n41496) );
  AND U41792 ( .A(n41497), .B(n41498), .Z(n41279) );
  NANDN U41793 ( .A(n41499), .B(n41500), .Z(n41498) );
  OR U41794 ( .A(n41501), .B(n41502), .Z(n41500) );
  NAND U41795 ( .A(n41502), .B(n41501), .Z(n41497) );
  ANDN U41796 ( .B(B[133]), .A(n71), .Z(n41281) );
  XNOR U41797 ( .A(n41289), .B(n41503), .Z(n41282) );
  XNOR U41798 ( .A(n41288), .B(n41286), .Z(n41503) );
  AND U41799 ( .A(n41504), .B(n41505), .Z(n41286) );
  NANDN U41800 ( .A(n41506), .B(n41507), .Z(n41505) );
  NANDN U41801 ( .A(n41508), .B(n41509), .Z(n41507) );
  NANDN U41802 ( .A(n41509), .B(n41508), .Z(n41504) );
  ANDN U41803 ( .B(B[134]), .A(n72), .Z(n41288) );
  XNOR U41804 ( .A(n41296), .B(n41510), .Z(n41289) );
  XNOR U41805 ( .A(n41295), .B(n41293), .Z(n41510) );
  AND U41806 ( .A(n41511), .B(n41512), .Z(n41293) );
  NANDN U41807 ( .A(n41513), .B(n41514), .Z(n41512) );
  OR U41808 ( .A(n41515), .B(n41516), .Z(n41514) );
  NAND U41809 ( .A(n41516), .B(n41515), .Z(n41511) );
  ANDN U41810 ( .B(B[135]), .A(n73), .Z(n41295) );
  XNOR U41811 ( .A(n41303), .B(n41517), .Z(n41296) );
  XNOR U41812 ( .A(n41302), .B(n41300), .Z(n41517) );
  AND U41813 ( .A(n41518), .B(n41519), .Z(n41300) );
  NANDN U41814 ( .A(n41520), .B(n41521), .Z(n41519) );
  NANDN U41815 ( .A(n41522), .B(n41523), .Z(n41521) );
  NANDN U41816 ( .A(n41523), .B(n41522), .Z(n41518) );
  ANDN U41817 ( .B(B[136]), .A(n74), .Z(n41302) );
  XNOR U41818 ( .A(n41310), .B(n41524), .Z(n41303) );
  XNOR U41819 ( .A(n41309), .B(n41307), .Z(n41524) );
  AND U41820 ( .A(n41525), .B(n41526), .Z(n41307) );
  NANDN U41821 ( .A(n41527), .B(n41528), .Z(n41526) );
  OR U41822 ( .A(n41529), .B(n41530), .Z(n41528) );
  NAND U41823 ( .A(n41530), .B(n41529), .Z(n41525) );
  ANDN U41824 ( .B(B[137]), .A(n75), .Z(n41309) );
  XNOR U41825 ( .A(n41317), .B(n41531), .Z(n41310) );
  XNOR U41826 ( .A(n41316), .B(n41314), .Z(n41531) );
  AND U41827 ( .A(n41532), .B(n41533), .Z(n41314) );
  NANDN U41828 ( .A(n41534), .B(n41535), .Z(n41533) );
  NANDN U41829 ( .A(n41536), .B(n41537), .Z(n41535) );
  NANDN U41830 ( .A(n41537), .B(n41536), .Z(n41532) );
  ANDN U41831 ( .B(B[138]), .A(n76), .Z(n41316) );
  XNOR U41832 ( .A(n41324), .B(n41538), .Z(n41317) );
  XNOR U41833 ( .A(n41323), .B(n41321), .Z(n41538) );
  AND U41834 ( .A(n41539), .B(n41540), .Z(n41321) );
  NANDN U41835 ( .A(n41541), .B(n41542), .Z(n41540) );
  OR U41836 ( .A(n41543), .B(n41544), .Z(n41542) );
  NAND U41837 ( .A(n41544), .B(n41543), .Z(n41539) );
  ANDN U41838 ( .B(B[139]), .A(n77), .Z(n41323) );
  XNOR U41839 ( .A(n41331), .B(n41545), .Z(n41324) );
  XNOR U41840 ( .A(n41330), .B(n41328), .Z(n41545) );
  AND U41841 ( .A(n41546), .B(n41547), .Z(n41328) );
  NANDN U41842 ( .A(n41548), .B(n41549), .Z(n41547) );
  NANDN U41843 ( .A(n41550), .B(n41551), .Z(n41549) );
  NANDN U41844 ( .A(n41551), .B(n41550), .Z(n41546) );
  ANDN U41845 ( .B(B[140]), .A(n78), .Z(n41330) );
  XNOR U41846 ( .A(n41338), .B(n41552), .Z(n41331) );
  XNOR U41847 ( .A(n41337), .B(n41335), .Z(n41552) );
  AND U41848 ( .A(n41553), .B(n41554), .Z(n41335) );
  NANDN U41849 ( .A(n41555), .B(n41556), .Z(n41554) );
  OR U41850 ( .A(n41557), .B(n41558), .Z(n41556) );
  NAND U41851 ( .A(n41558), .B(n41557), .Z(n41553) );
  ANDN U41852 ( .B(B[141]), .A(n79), .Z(n41337) );
  XNOR U41853 ( .A(n41345), .B(n41559), .Z(n41338) );
  XNOR U41854 ( .A(n41344), .B(n41342), .Z(n41559) );
  AND U41855 ( .A(n41560), .B(n41561), .Z(n41342) );
  NANDN U41856 ( .A(n41562), .B(n41563), .Z(n41561) );
  NANDN U41857 ( .A(n41564), .B(n41565), .Z(n41563) );
  NANDN U41858 ( .A(n41565), .B(n41564), .Z(n41560) );
  ANDN U41859 ( .B(B[142]), .A(n80), .Z(n41344) );
  XNOR U41860 ( .A(n41352), .B(n41566), .Z(n41345) );
  XNOR U41861 ( .A(n41351), .B(n41349), .Z(n41566) );
  AND U41862 ( .A(n41567), .B(n41568), .Z(n41349) );
  NANDN U41863 ( .A(n41569), .B(n41570), .Z(n41568) );
  OR U41864 ( .A(n41571), .B(n41572), .Z(n41570) );
  NAND U41865 ( .A(n41572), .B(n41571), .Z(n41567) );
  ANDN U41866 ( .B(B[143]), .A(n81), .Z(n41351) );
  XNOR U41867 ( .A(n41359), .B(n41573), .Z(n41352) );
  XNOR U41868 ( .A(n41358), .B(n41356), .Z(n41573) );
  AND U41869 ( .A(n41574), .B(n41575), .Z(n41356) );
  NANDN U41870 ( .A(n41576), .B(n41577), .Z(n41575) );
  NAND U41871 ( .A(n41578), .B(n41579), .Z(n41577) );
  ANDN U41872 ( .B(B[144]), .A(n82), .Z(n41358) );
  XOR U41873 ( .A(n41365), .B(n41580), .Z(n41359) );
  XNOR U41874 ( .A(n41363), .B(n41366), .Z(n41580) );
  NAND U41875 ( .A(A[2]), .B(B[145]), .Z(n41366) );
  NANDN U41876 ( .A(n41581), .B(n41582), .Z(n41363) );
  AND U41877 ( .A(A[0]), .B(B[146]), .Z(n41582) );
  XNOR U41878 ( .A(n41368), .B(n41583), .Z(n41365) );
  NAND U41879 ( .A(A[0]), .B(B[147]), .Z(n41583) );
  NAND U41880 ( .A(B[146]), .B(A[1]), .Z(n41368) );
  NAND U41881 ( .A(n41584), .B(n41585), .Z(n502) );
  NANDN U41882 ( .A(n41586), .B(n41587), .Z(n41585) );
  OR U41883 ( .A(n41588), .B(n41589), .Z(n41587) );
  NAND U41884 ( .A(n41589), .B(n41588), .Z(n41584) );
  XOR U41885 ( .A(n504), .B(n503), .Z(\A1[144] ) );
  XOR U41886 ( .A(n41589), .B(n41590), .Z(n503) );
  XNOR U41887 ( .A(n41588), .B(n41586), .Z(n41590) );
  AND U41888 ( .A(n41591), .B(n41592), .Z(n41586) );
  NANDN U41889 ( .A(n41593), .B(n41594), .Z(n41592) );
  NANDN U41890 ( .A(n41595), .B(n41596), .Z(n41594) );
  NANDN U41891 ( .A(n41596), .B(n41595), .Z(n41591) );
  ANDN U41892 ( .B(B[115]), .A(n54), .Z(n41588) );
  XNOR U41893 ( .A(n41383), .B(n41597), .Z(n41589) );
  XNOR U41894 ( .A(n41382), .B(n41380), .Z(n41597) );
  AND U41895 ( .A(n41598), .B(n41599), .Z(n41380) );
  NANDN U41896 ( .A(n41600), .B(n41601), .Z(n41599) );
  OR U41897 ( .A(n41602), .B(n41603), .Z(n41601) );
  NAND U41898 ( .A(n41603), .B(n41602), .Z(n41598) );
  ANDN U41899 ( .B(B[116]), .A(n55), .Z(n41382) );
  XNOR U41900 ( .A(n41390), .B(n41604), .Z(n41383) );
  XNOR U41901 ( .A(n41389), .B(n41387), .Z(n41604) );
  AND U41902 ( .A(n41605), .B(n41606), .Z(n41387) );
  NANDN U41903 ( .A(n41607), .B(n41608), .Z(n41606) );
  NANDN U41904 ( .A(n41609), .B(n41610), .Z(n41608) );
  NANDN U41905 ( .A(n41610), .B(n41609), .Z(n41605) );
  ANDN U41906 ( .B(B[117]), .A(n56), .Z(n41389) );
  XNOR U41907 ( .A(n41397), .B(n41611), .Z(n41390) );
  XNOR U41908 ( .A(n41396), .B(n41394), .Z(n41611) );
  AND U41909 ( .A(n41612), .B(n41613), .Z(n41394) );
  NANDN U41910 ( .A(n41614), .B(n41615), .Z(n41613) );
  OR U41911 ( .A(n41616), .B(n41617), .Z(n41615) );
  NAND U41912 ( .A(n41617), .B(n41616), .Z(n41612) );
  ANDN U41913 ( .B(B[118]), .A(n57), .Z(n41396) );
  XNOR U41914 ( .A(n41404), .B(n41618), .Z(n41397) );
  XNOR U41915 ( .A(n41403), .B(n41401), .Z(n41618) );
  AND U41916 ( .A(n41619), .B(n41620), .Z(n41401) );
  NANDN U41917 ( .A(n41621), .B(n41622), .Z(n41620) );
  NANDN U41918 ( .A(n41623), .B(n41624), .Z(n41622) );
  NANDN U41919 ( .A(n41624), .B(n41623), .Z(n41619) );
  ANDN U41920 ( .B(B[119]), .A(n58), .Z(n41403) );
  XNOR U41921 ( .A(n41411), .B(n41625), .Z(n41404) );
  XNOR U41922 ( .A(n41410), .B(n41408), .Z(n41625) );
  AND U41923 ( .A(n41626), .B(n41627), .Z(n41408) );
  NANDN U41924 ( .A(n41628), .B(n41629), .Z(n41627) );
  OR U41925 ( .A(n41630), .B(n41631), .Z(n41629) );
  NAND U41926 ( .A(n41631), .B(n41630), .Z(n41626) );
  ANDN U41927 ( .B(B[120]), .A(n59), .Z(n41410) );
  XNOR U41928 ( .A(n41418), .B(n41632), .Z(n41411) );
  XNOR U41929 ( .A(n41417), .B(n41415), .Z(n41632) );
  AND U41930 ( .A(n41633), .B(n41634), .Z(n41415) );
  NANDN U41931 ( .A(n41635), .B(n41636), .Z(n41634) );
  NANDN U41932 ( .A(n41637), .B(n41638), .Z(n41636) );
  NANDN U41933 ( .A(n41638), .B(n41637), .Z(n41633) );
  ANDN U41934 ( .B(B[121]), .A(n60), .Z(n41417) );
  XNOR U41935 ( .A(n41425), .B(n41639), .Z(n41418) );
  XNOR U41936 ( .A(n41424), .B(n41422), .Z(n41639) );
  AND U41937 ( .A(n41640), .B(n41641), .Z(n41422) );
  NANDN U41938 ( .A(n41642), .B(n41643), .Z(n41641) );
  OR U41939 ( .A(n41644), .B(n41645), .Z(n41643) );
  NAND U41940 ( .A(n41645), .B(n41644), .Z(n41640) );
  ANDN U41941 ( .B(B[122]), .A(n61), .Z(n41424) );
  XNOR U41942 ( .A(n41432), .B(n41646), .Z(n41425) );
  XNOR U41943 ( .A(n41431), .B(n41429), .Z(n41646) );
  AND U41944 ( .A(n41647), .B(n41648), .Z(n41429) );
  NANDN U41945 ( .A(n41649), .B(n41650), .Z(n41648) );
  NANDN U41946 ( .A(n41651), .B(n41652), .Z(n41650) );
  NANDN U41947 ( .A(n41652), .B(n41651), .Z(n41647) );
  ANDN U41948 ( .B(B[123]), .A(n62), .Z(n41431) );
  XNOR U41949 ( .A(n41439), .B(n41653), .Z(n41432) );
  XNOR U41950 ( .A(n41438), .B(n41436), .Z(n41653) );
  AND U41951 ( .A(n41654), .B(n41655), .Z(n41436) );
  NANDN U41952 ( .A(n41656), .B(n41657), .Z(n41655) );
  OR U41953 ( .A(n41658), .B(n41659), .Z(n41657) );
  NAND U41954 ( .A(n41659), .B(n41658), .Z(n41654) );
  ANDN U41955 ( .B(B[124]), .A(n63), .Z(n41438) );
  XNOR U41956 ( .A(n41446), .B(n41660), .Z(n41439) );
  XNOR U41957 ( .A(n41445), .B(n41443), .Z(n41660) );
  AND U41958 ( .A(n41661), .B(n41662), .Z(n41443) );
  NANDN U41959 ( .A(n41663), .B(n41664), .Z(n41662) );
  NANDN U41960 ( .A(n41665), .B(n41666), .Z(n41664) );
  NANDN U41961 ( .A(n41666), .B(n41665), .Z(n41661) );
  ANDN U41962 ( .B(B[125]), .A(n64), .Z(n41445) );
  XNOR U41963 ( .A(n41453), .B(n41667), .Z(n41446) );
  XNOR U41964 ( .A(n41452), .B(n41450), .Z(n41667) );
  AND U41965 ( .A(n41668), .B(n41669), .Z(n41450) );
  NANDN U41966 ( .A(n41670), .B(n41671), .Z(n41669) );
  OR U41967 ( .A(n41672), .B(n41673), .Z(n41671) );
  NAND U41968 ( .A(n41673), .B(n41672), .Z(n41668) );
  ANDN U41969 ( .B(B[126]), .A(n65), .Z(n41452) );
  XNOR U41970 ( .A(n41460), .B(n41674), .Z(n41453) );
  XNOR U41971 ( .A(n41459), .B(n41457), .Z(n41674) );
  AND U41972 ( .A(n41675), .B(n41676), .Z(n41457) );
  NANDN U41973 ( .A(n41677), .B(n41678), .Z(n41676) );
  NANDN U41974 ( .A(n41679), .B(n41680), .Z(n41678) );
  NANDN U41975 ( .A(n41680), .B(n41679), .Z(n41675) );
  ANDN U41976 ( .B(B[127]), .A(n66), .Z(n41459) );
  XNOR U41977 ( .A(n41467), .B(n41681), .Z(n41460) );
  XNOR U41978 ( .A(n41466), .B(n41464), .Z(n41681) );
  AND U41979 ( .A(n41682), .B(n41683), .Z(n41464) );
  NANDN U41980 ( .A(n41684), .B(n41685), .Z(n41683) );
  OR U41981 ( .A(n41686), .B(n41687), .Z(n41685) );
  NAND U41982 ( .A(n41687), .B(n41686), .Z(n41682) );
  ANDN U41983 ( .B(B[128]), .A(n67), .Z(n41466) );
  XNOR U41984 ( .A(n41474), .B(n41688), .Z(n41467) );
  XNOR U41985 ( .A(n41473), .B(n41471), .Z(n41688) );
  AND U41986 ( .A(n41689), .B(n41690), .Z(n41471) );
  NANDN U41987 ( .A(n41691), .B(n41692), .Z(n41690) );
  NANDN U41988 ( .A(n41693), .B(n41694), .Z(n41692) );
  NANDN U41989 ( .A(n41694), .B(n41693), .Z(n41689) );
  ANDN U41990 ( .B(B[129]), .A(n68), .Z(n41473) );
  XNOR U41991 ( .A(n41481), .B(n41695), .Z(n41474) );
  XNOR U41992 ( .A(n41480), .B(n41478), .Z(n41695) );
  AND U41993 ( .A(n41696), .B(n41697), .Z(n41478) );
  NANDN U41994 ( .A(n41698), .B(n41699), .Z(n41697) );
  OR U41995 ( .A(n41700), .B(n41701), .Z(n41699) );
  NAND U41996 ( .A(n41701), .B(n41700), .Z(n41696) );
  ANDN U41997 ( .B(B[130]), .A(n69), .Z(n41480) );
  XNOR U41998 ( .A(n41488), .B(n41702), .Z(n41481) );
  XNOR U41999 ( .A(n41487), .B(n41485), .Z(n41702) );
  AND U42000 ( .A(n41703), .B(n41704), .Z(n41485) );
  NANDN U42001 ( .A(n41705), .B(n41706), .Z(n41704) );
  NANDN U42002 ( .A(n41707), .B(n41708), .Z(n41706) );
  NANDN U42003 ( .A(n41708), .B(n41707), .Z(n41703) );
  ANDN U42004 ( .B(B[131]), .A(n70), .Z(n41487) );
  XNOR U42005 ( .A(n41495), .B(n41709), .Z(n41488) );
  XNOR U42006 ( .A(n41494), .B(n41492), .Z(n41709) );
  AND U42007 ( .A(n41710), .B(n41711), .Z(n41492) );
  NANDN U42008 ( .A(n41712), .B(n41713), .Z(n41711) );
  OR U42009 ( .A(n41714), .B(n41715), .Z(n41713) );
  NAND U42010 ( .A(n41715), .B(n41714), .Z(n41710) );
  ANDN U42011 ( .B(B[132]), .A(n71), .Z(n41494) );
  XNOR U42012 ( .A(n41502), .B(n41716), .Z(n41495) );
  XNOR U42013 ( .A(n41501), .B(n41499), .Z(n41716) );
  AND U42014 ( .A(n41717), .B(n41718), .Z(n41499) );
  NANDN U42015 ( .A(n41719), .B(n41720), .Z(n41718) );
  NANDN U42016 ( .A(n41721), .B(n41722), .Z(n41720) );
  NANDN U42017 ( .A(n41722), .B(n41721), .Z(n41717) );
  ANDN U42018 ( .B(B[133]), .A(n72), .Z(n41501) );
  XNOR U42019 ( .A(n41509), .B(n41723), .Z(n41502) );
  XNOR U42020 ( .A(n41508), .B(n41506), .Z(n41723) );
  AND U42021 ( .A(n41724), .B(n41725), .Z(n41506) );
  NANDN U42022 ( .A(n41726), .B(n41727), .Z(n41725) );
  OR U42023 ( .A(n41728), .B(n41729), .Z(n41727) );
  NAND U42024 ( .A(n41729), .B(n41728), .Z(n41724) );
  ANDN U42025 ( .B(B[134]), .A(n73), .Z(n41508) );
  XNOR U42026 ( .A(n41516), .B(n41730), .Z(n41509) );
  XNOR U42027 ( .A(n41515), .B(n41513), .Z(n41730) );
  AND U42028 ( .A(n41731), .B(n41732), .Z(n41513) );
  NANDN U42029 ( .A(n41733), .B(n41734), .Z(n41732) );
  NANDN U42030 ( .A(n41735), .B(n41736), .Z(n41734) );
  NANDN U42031 ( .A(n41736), .B(n41735), .Z(n41731) );
  ANDN U42032 ( .B(B[135]), .A(n74), .Z(n41515) );
  XNOR U42033 ( .A(n41523), .B(n41737), .Z(n41516) );
  XNOR U42034 ( .A(n41522), .B(n41520), .Z(n41737) );
  AND U42035 ( .A(n41738), .B(n41739), .Z(n41520) );
  NANDN U42036 ( .A(n41740), .B(n41741), .Z(n41739) );
  OR U42037 ( .A(n41742), .B(n41743), .Z(n41741) );
  NAND U42038 ( .A(n41743), .B(n41742), .Z(n41738) );
  ANDN U42039 ( .B(B[136]), .A(n75), .Z(n41522) );
  XNOR U42040 ( .A(n41530), .B(n41744), .Z(n41523) );
  XNOR U42041 ( .A(n41529), .B(n41527), .Z(n41744) );
  AND U42042 ( .A(n41745), .B(n41746), .Z(n41527) );
  NANDN U42043 ( .A(n41747), .B(n41748), .Z(n41746) );
  NANDN U42044 ( .A(n41749), .B(n41750), .Z(n41748) );
  NANDN U42045 ( .A(n41750), .B(n41749), .Z(n41745) );
  ANDN U42046 ( .B(B[137]), .A(n76), .Z(n41529) );
  XNOR U42047 ( .A(n41537), .B(n41751), .Z(n41530) );
  XNOR U42048 ( .A(n41536), .B(n41534), .Z(n41751) );
  AND U42049 ( .A(n41752), .B(n41753), .Z(n41534) );
  NANDN U42050 ( .A(n41754), .B(n41755), .Z(n41753) );
  OR U42051 ( .A(n41756), .B(n41757), .Z(n41755) );
  NAND U42052 ( .A(n41757), .B(n41756), .Z(n41752) );
  ANDN U42053 ( .B(B[138]), .A(n77), .Z(n41536) );
  XNOR U42054 ( .A(n41544), .B(n41758), .Z(n41537) );
  XNOR U42055 ( .A(n41543), .B(n41541), .Z(n41758) );
  AND U42056 ( .A(n41759), .B(n41760), .Z(n41541) );
  NANDN U42057 ( .A(n41761), .B(n41762), .Z(n41760) );
  NANDN U42058 ( .A(n41763), .B(n41764), .Z(n41762) );
  NANDN U42059 ( .A(n41764), .B(n41763), .Z(n41759) );
  ANDN U42060 ( .B(B[139]), .A(n78), .Z(n41543) );
  XNOR U42061 ( .A(n41551), .B(n41765), .Z(n41544) );
  XNOR U42062 ( .A(n41550), .B(n41548), .Z(n41765) );
  AND U42063 ( .A(n41766), .B(n41767), .Z(n41548) );
  NANDN U42064 ( .A(n41768), .B(n41769), .Z(n41767) );
  OR U42065 ( .A(n41770), .B(n41771), .Z(n41769) );
  NAND U42066 ( .A(n41771), .B(n41770), .Z(n41766) );
  ANDN U42067 ( .B(B[140]), .A(n79), .Z(n41550) );
  XNOR U42068 ( .A(n41558), .B(n41772), .Z(n41551) );
  XNOR U42069 ( .A(n41557), .B(n41555), .Z(n41772) );
  AND U42070 ( .A(n41773), .B(n41774), .Z(n41555) );
  NANDN U42071 ( .A(n41775), .B(n41776), .Z(n41774) );
  NANDN U42072 ( .A(n41777), .B(n41778), .Z(n41776) );
  NANDN U42073 ( .A(n41778), .B(n41777), .Z(n41773) );
  ANDN U42074 ( .B(B[141]), .A(n80), .Z(n41557) );
  XNOR U42075 ( .A(n41565), .B(n41779), .Z(n41558) );
  XNOR U42076 ( .A(n41564), .B(n41562), .Z(n41779) );
  AND U42077 ( .A(n41780), .B(n41781), .Z(n41562) );
  NANDN U42078 ( .A(n41782), .B(n41783), .Z(n41781) );
  OR U42079 ( .A(n41784), .B(n41785), .Z(n41783) );
  NAND U42080 ( .A(n41785), .B(n41784), .Z(n41780) );
  ANDN U42081 ( .B(B[142]), .A(n81), .Z(n41564) );
  XNOR U42082 ( .A(n41572), .B(n41786), .Z(n41565) );
  XNOR U42083 ( .A(n41571), .B(n41569), .Z(n41786) );
  AND U42084 ( .A(n41787), .B(n41788), .Z(n41569) );
  NANDN U42085 ( .A(n41789), .B(n41790), .Z(n41788) );
  NAND U42086 ( .A(n41791), .B(n41792), .Z(n41790) );
  ANDN U42087 ( .B(B[143]), .A(n82), .Z(n41571) );
  XOR U42088 ( .A(n41578), .B(n41793), .Z(n41572) );
  XNOR U42089 ( .A(n41576), .B(n41579), .Z(n41793) );
  NAND U42090 ( .A(A[2]), .B(B[144]), .Z(n41579) );
  NANDN U42091 ( .A(n41794), .B(n41795), .Z(n41576) );
  AND U42092 ( .A(A[0]), .B(B[145]), .Z(n41795) );
  XNOR U42093 ( .A(n41581), .B(n41796), .Z(n41578) );
  NAND U42094 ( .A(A[0]), .B(B[146]), .Z(n41796) );
  NAND U42095 ( .A(B[145]), .B(A[1]), .Z(n41581) );
  NAND U42096 ( .A(n41797), .B(n41798), .Z(n504) );
  NANDN U42097 ( .A(n41799), .B(n41800), .Z(n41798) );
  OR U42098 ( .A(n41801), .B(n41802), .Z(n41800) );
  NAND U42099 ( .A(n41802), .B(n41801), .Z(n41797) );
  XOR U42100 ( .A(n506), .B(n505), .Z(\A1[143] ) );
  XOR U42101 ( .A(n41802), .B(n41803), .Z(n505) );
  XNOR U42102 ( .A(n41801), .B(n41799), .Z(n41803) );
  AND U42103 ( .A(n41804), .B(n41805), .Z(n41799) );
  NANDN U42104 ( .A(n41806), .B(n41807), .Z(n41805) );
  NANDN U42105 ( .A(n41808), .B(n41809), .Z(n41807) );
  NANDN U42106 ( .A(n41809), .B(n41808), .Z(n41804) );
  ANDN U42107 ( .B(B[114]), .A(n54), .Z(n41801) );
  XNOR U42108 ( .A(n41596), .B(n41810), .Z(n41802) );
  XNOR U42109 ( .A(n41595), .B(n41593), .Z(n41810) );
  AND U42110 ( .A(n41811), .B(n41812), .Z(n41593) );
  NANDN U42111 ( .A(n41813), .B(n41814), .Z(n41812) );
  OR U42112 ( .A(n41815), .B(n41816), .Z(n41814) );
  NAND U42113 ( .A(n41816), .B(n41815), .Z(n41811) );
  ANDN U42114 ( .B(B[115]), .A(n55), .Z(n41595) );
  XNOR U42115 ( .A(n41603), .B(n41817), .Z(n41596) );
  XNOR U42116 ( .A(n41602), .B(n41600), .Z(n41817) );
  AND U42117 ( .A(n41818), .B(n41819), .Z(n41600) );
  NANDN U42118 ( .A(n41820), .B(n41821), .Z(n41819) );
  NANDN U42119 ( .A(n41822), .B(n41823), .Z(n41821) );
  NANDN U42120 ( .A(n41823), .B(n41822), .Z(n41818) );
  ANDN U42121 ( .B(B[116]), .A(n56), .Z(n41602) );
  XNOR U42122 ( .A(n41610), .B(n41824), .Z(n41603) );
  XNOR U42123 ( .A(n41609), .B(n41607), .Z(n41824) );
  AND U42124 ( .A(n41825), .B(n41826), .Z(n41607) );
  NANDN U42125 ( .A(n41827), .B(n41828), .Z(n41826) );
  OR U42126 ( .A(n41829), .B(n41830), .Z(n41828) );
  NAND U42127 ( .A(n41830), .B(n41829), .Z(n41825) );
  ANDN U42128 ( .B(B[117]), .A(n57), .Z(n41609) );
  XNOR U42129 ( .A(n41617), .B(n41831), .Z(n41610) );
  XNOR U42130 ( .A(n41616), .B(n41614), .Z(n41831) );
  AND U42131 ( .A(n41832), .B(n41833), .Z(n41614) );
  NANDN U42132 ( .A(n41834), .B(n41835), .Z(n41833) );
  NANDN U42133 ( .A(n41836), .B(n41837), .Z(n41835) );
  NANDN U42134 ( .A(n41837), .B(n41836), .Z(n41832) );
  ANDN U42135 ( .B(B[118]), .A(n58), .Z(n41616) );
  XNOR U42136 ( .A(n41624), .B(n41838), .Z(n41617) );
  XNOR U42137 ( .A(n41623), .B(n41621), .Z(n41838) );
  AND U42138 ( .A(n41839), .B(n41840), .Z(n41621) );
  NANDN U42139 ( .A(n41841), .B(n41842), .Z(n41840) );
  OR U42140 ( .A(n41843), .B(n41844), .Z(n41842) );
  NAND U42141 ( .A(n41844), .B(n41843), .Z(n41839) );
  ANDN U42142 ( .B(B[119]), .A(n59), .Z(n41623) );
  XNOR U42143 ( .A(n41631), .B(n41845), .Z(n41624) );
  XNOR U42144 ( .A(n41630), .B(n41628), .Z(n41845) );
  AND U42145 ( .A(n41846), .B(n41847), .Z(n41628) );
  NANDN U42146 ( .A(n41848), .B(n41849), .Z(n41847) );
  NANDN U42147 ( .A(n41850), .B(n41851), .Z(n41849) );
  NANDN U42148 ( .A(n41851), .B(n41850), .Z(n41846) );
  ANDN U42149 ( .B(B[120]), .A(n60), .Z(n41630) );
  XNOR U42150 ( .A(n41638), .B(n41852), .Z(n41631) );
  XNOR U42151 ( .A(n41637), .B(n41635), .Z(n41852) );
  AND U42152 ( .A(n41853), .B(n41854), .Z(n41635) );
  NANDN U42153 ( .A(n41855), .B(n41856), .Z(n41854) );
  OR U42154 ( .A(n41857), .B(n41858), .Z(n41856) );
  NAND U42155 ( .A(n41858), .B(n41857), .Z(n41853) );
  ANDN U42156 ( .B(B[121]), .A(n61), .Z(n41637) );
  XNOR U42157 ( .A(n41645), .B(n41859), .Z(n41638) );
  XNOR U42158 ( .A(n41644), .B(n41642), .Z(n41859) );
  AND U42159 ( .A(n41860), .B(n41861), .Z(n41642) );
  NANDN U42160 ( .A(n41862), .B(n41863), .Z(n41861) );
  NANDN U42161 ( .A(n41864), .B(n41865), .Z(n41863) );
  NANDN U42162 ( .A(n41865), .B(n41864), .Z(n41860) );
  ANDN U42163 ( .B(B[122]), .A(n62), .Z(n41644) );
  XNOR U42164 ( .A(n41652), .B(n41866), .Z(n41645) );
  XNOR U42165 ( .A(n41651), .B(n41649), .Z(n41866) );
  AND U42166 ( .A(n41867), .B(n41868), .Z(n41649) );
  NANDN U42167 ( .A(n41869), .B(n41870), .Z(n41868) );
  OR U42168 ( .A(n41871), .B(n41872), .Z(n41870) );
  NAND U42169 ( .A(n41872), .B(n41871), .Z(n41867) );
  ANDN U42170 ( .B(B[123]), .A(n63), .Z(n41651) );
  XNOR U42171 ( .A(n41659), .B(n41873), .Z(n41652) );
  XNOR U42172 ( .A(n41658), .B(n41656), .Z(n41873) );
  AND U42173 ( .A(n41874), .B(n41875), .Z(n41656) );
  NANDN U42174 ( .A(n41876), .B(n41877), .Z(n41875) );
  NANDN U42175 ( .A(n41878), .B(n41879), .Z(n41877) );
  NANDN U42176 ( .A(n41879), .B(n41878), .Z(n41874) );
  ANDN U42177 ( .B(B[124]), .A(n64), .Z(n41658) );
  XNOR U42178 ( .A(n41666), .B(n41880), .Z(n41659) );
  XNOR U42179 ( .A(n41665), .B(n41663), .Z(n41880) );
  AND U42180 ( .A(n41881), .B(n41882), .Z(n41663) );
  NANDN U42181 ( .A(n41883), .B(n41884), .Z(n41882) );
  OR U42182 ( .A(n41885), .B(n41886), .Z(n41884) );
  NAND U42183 ( .A(n41886), .B(n41885), .Z(n41881) );
  ANDN U42184 ( .B(B[125]), .A(n65), .Z(n41665) );
  XNOR U42185 ( .A(n41673), .B(n41887), .Z(n41666) );
  XNOR U42186 ( .A(n41672), .B(n41670), .Z(n41887) );
  AND U42187 ( .A(n41888), .B(n41889), .Z(n41670) );
  NANDN U42188 ( .A(n41890), .B(n41891), .Z(n41889) );
  NANDN U42189 ( .A(n41892), .B(n41893), .Z(n41891) );
  NANDN U42190 ( .A(n41893), .B(n41892), .Z(n41888) );
  ANDN U42191 ( .B(B[126]), .A(n66), .Z(n41672) );
  XNOR U42192 ( .A(n41680), .B(n41894), .Z(n41673) );
  XNOR U42193 ( .A(n41679), .B(n41677), .Z(n41894) );
  AND U42194 ( .A(n41895), .B(n41896), .Z(n41677) );
  NANDN U42195 ( .A(n41897), .B(n41898), .Z(n41896) );
  OR U42196 ( .A(n41899), .B(n41900), .Z(n41898) );
  NAND U42197 ( .A(n41900), .B(n41899), .Z(n41895) );
  ANDN U42198 ( .B(B[127]), .A(n67), .Z(n41679) );
  XNOR U42199 ( .A(n41687), .B(n41901), .Z(n41680) );
  XNOR U42200 ( .A(n41686), .B(n41684), .Z(n41901) );
  AND U42201 ( .A(n41902), .B(n41903), .Z(n41684) );
  NANDN U42202 ( .A(n41904), .B(n41905), .Z(n41903) );
  NANDN U42203 ( .A(n41906), .B(n41907), .Z(n41905) );
  NANDN U42204 ( .A(n41907), .B(n41906), .Z(n41902) );
  ANDN U42205 ( .B(B[128]), .A(n68), .Z(n41686) );
  XNOR U42206 ( .A(n41694), .B(n41908), .Z(n41687) );
  XNOR U42207 ( .A(n41693), .B(n41691), .Z(n41908) );
  AND U42208 ( .A(n41909), .B(n41910), .Z(n41691) );
  NANDN U42209 ( .A(n41911), .B(n41912), .Z(n41910) );
  OR U42210 ( .A(n41913), .B(n41914), .Z(n41912) );
  NAND U42211 ( .A(n41914), .B(n41913), .Z(n41909) );
  ANDN U42212 ( .B(B[129]), .A(n69), .Z(n41693) );
  XNOR U42213 ( .A(n41701), .B(n41915), .Z(n41694) );
  XNOR U42214 ( .A(n41700), .B(n41698), .Z(n41915) );
  AND U42215 ( .A(n41916), .B(n41917), .Z(n41698) );
  NANDN U42216 ( .A(n41918), .B(n41919), .Z(n41917) );
  NANDN U42217 ( .A(n41920), .B(n41921), .Z(n41919) );
  NANDN U42218 ( .A(n41921), .B(n41920), .Z(n41916) );
  ANDN U42219 ( .B(B[130]), .A(n70), .Z(n41700) );
  XNOR U42220 ( .A(n41708), .B(n41922), .Z(n41701) );
  XNOR U42221 ( .A(n41707), .B(n41705), .Z(n41922) );
  AND U42222 ( .A(n41923), .B(n41924), .Z(n41705) );
  NANDN U42223 ( .A(n41925), .B(n41926), .Z(n41924) );
  OR U42224 ( .A(n41927), .B(n41928), .Z(n41926) );
  NAND U42225 ( .A(n41928), .B(n41927), .Z(n41923) );
  ANDN U42226 ( .B(B[131]), .A(n71), .Z(n41707) );
  XNOR U42227 ( .A(n41715), .B(n41929), .Z(n41708) );
  XNOR U42228 ( .A(n41714), .B(n41712), .Z(n41929) );
  AND U42229 ( .A(n41930), .B(n41931), .Z(n41712) );
  NANDN U42230 ( .A(n41932), .B(n41933), .Z(n41931) );
  NANDN U42231 ( .A(n41934), .B(n41935), .Z(n41933) );
  NANDN U42232 ( .A(n41935), .B(n41934), .Z(n41930) );
  ANDN U42233 ( .B(B[132]), .A(n72), .Z(n41714) );
  XNOR U42234 ( .A(n41722), .B(n41936), .Z(n41715) );
  XNOR U42235 ( .A(n41721), .B(n41719), .Z(n41936) );
  AND U42236 ( .A(n41937), .B(n41938), .Z(n41719) );
  NANDN U42237 ( .A(n41939), .B(n41940), .Z(n41938) );
  OR U42238 ( .A(n41941), .B(n41942), .Z(n41940) );
  NAND U42239 ( .A(n41942), .B(n41941), .Z(n41937) );
  ANDN U42240 ( .B(B[133]), .A(n73), .Z(n41721) );
  XNOR U42241 ( .A(n41729), .B(n41943), .Z(n41722) );
  XNOR U42242 ( .A(n41728), .B(n41726), .Z(n41943) );
  AND U42243 ( .A(n41944), .B(n41945), .Z(n41726) );
  NANDN U42244 ( .A(n41946), .B(n41947), .Z(n41945) );
  NANDN U42245 ( .A(n41948), .B(n41949), .Z(n41947) );
  NANDN U42246 ( .A(n41949), .B(n41948), .Z(n41944) );
  ANDN U42247 ( .B(B[134]), .A(n74), .Z(n41728) );
  XNOR U42248 ( .A(n41736), .B(n41950), .Z(n41729) );
  XNOR U42249 ( .A(n41735), .B(n41733), .Z(n41950) );
  AND U42250 ( .A(n41951), .B(n41952), .Z(n41733) );
  NANDN U42251 ( .A(n41953), .B(n41954), .Z(n41952) );
  OR U42252 ( .A(n41955), .B(n41956), .Z(n41954) );
  NAND U42253 ( .A(n41956), .B(n41955), .Z(n41951) );
  ANDN U42254 ( .B(B[135]), .A(n75), .Z(n41735) );
  XNOR U42255 ( .A(n41743), .B(n41957), .Z(n41736) );
  XNOR U42256 ( .A(n41742), .B(n41740), .Z(n41957) );
  AND U42257 ( .A(n41958), .B(n41959), .Z(n41740) );
  NANDN U42258 ( .A(n41960), .B(n41961), .Z(n41959) );
  NANDN U42259 ( .A(n41962), .B(n41963), .Z(n41961) );
  NANDN U42260 ( .A(n41963), .B(n41962), .Z(n41958) );
  ANDN U42261 ( .B(B[136]), .A(n76), .Z(n41742) );
  XNOR U42262 ( .A(n41750), .B(n41964), .Z(n41743) );
  XNOR U42263 ( .A(n41749), .B(n41747), .Z(n41964) );
  AND U42264 ( .A(n41965), .B(n41966), .Z(n41747) );
  NANDN U42265 ( .A(n41967), .B(n41968), .Z(n41966) );
  OR U42266 ( .A(n41969), .B(n41970), .Z(n41968) );
  NAND U42267 ( .A(n41970), .B(n41969), .Z(n41965) );
  ANDN U42268 ( .B(B[137]), .A(n77), .Z(n41749) );
  XNOR U42269 ( .A(n41757), .B(n41971), .Z(n41750) );
  XNOR U42270 ( .A(n41756), .B(n41754), .Z(n41971) );
  AND U42271 ( .A(n41972), .B(n41973), .Z(n41754) );
  NANDN U42272 ( .A(n41974), .B(n41975), .Z(n41973) );
  NANDN U42273 ( .A(n41976), .B(n41977), .Z(n41975) );
  NANDN U42274 ( .A(n41977), .B(n41976), .Z(n41972) );
  ANDN U42275 ( .B(B[138]), .A(n78), .Z(n41756) );
  XNOR U42276 ( .A(n41764), .B(n41978), .Z(n41757) );
  XNOR U42277 ( .A(n41763), .B(n41761), .Z(n41978) );
  AND U42278 ( .A(n41979), .B(n41980), .Z(n41761) );
  NANDN U42279 ( .A(n41981), .B(n41982), .Z(n41980) );
  OR U42280 ( .A(n41983), .B(n41984), .Z(n41982) );
  NAND U42281 ( .A(n41984), .B(n41983), .Z(n41979) );
  ANDN U42282 ( .B(B[139]), .A(n79), .Z(n41763) );
  XNOR U42283 ( .A(n41771), .B(n41985), .Z(n41764) );
  XNOR U42284 ( .A(n41770), .B(n41768), .Z(n41985) );
  AND U42285 ( .A(n41986), .B(n41987), .Z(n41768) );
  NANDN U42286 ( .A(n41988), .B(n41989), .Z(n41987) );
  NANDN U42287 ( .A(n41990), .B(n41991), .Z(n41989) );
  NANDN U42288 ( .A(n41991), .B(n41990), .Z(n41986) );
  ANDN U42289 ( .B(B[140]), .A(n80), .Z(n41770) );
  XNOR U42290 ( .A(n41778), .B(n41992), .Z(n41771) );
  XNOR U42291 ( .A(n41777), .B(n41775), .Z(n41992) );
  AND U42292 ( .A(n41993), .B(n41994), .Z(n41775) );
  NANDN U42293 ( .A(n41995), .B(n41996), .Z(n41994) );
  OR U42294 ( .A(n41997), .B(n41998), .Z(n41996) );
  NAND U42295 ( .A(n41998), .B(n41997), .Z(n41993) );
  ANDN U42296 ( .B(B[141]), .A(n81), .Z(n41777) );
  XNOR U42297 ( .A(n41785), .B(n41999), .Z(n41778) );
  XNOR U42298 ( .A(n41784), .B(n41782), .Z(n41999) );
  AND U42299 ( .A(n42000), .B(n42001), .Z(n41782) );
  NANDN U42300 ( .A(n42002), .B(n42003), .Z(n42001) );
  NAND U42301 ( .A(n42004), .B(n42005), .Z(n42003) );
  ANDN U42302 ( .B(B[142]), .A(n82), .Z(n41784) );
  XOR U42303 ( .A(n41791), .B(n42006), .Z(n41785) );
  XNOR U42304 ( .A(n41789), .B(n41792), .Z(n42006) );
  NAND U42305 ( .A(A[2]), .B(B[143]), .Z(n41792) );
  NANDN U42306 ( .A(n42007), .B(n42008), .Z(n41789) );
  AND U42307 ( .A(A[0]), .B(B[144]), .Z(n42008) );
  XNOR U42308 ( .A(n41794), .B(n42009), .Z(n41791) );
  NAND U42309 ( .A(A[0]), .B(B[145]), .Z(n42009) );
  NAND U42310 ( .A(B[144]), .B(A[1]), .Z(n41794) );
  NAND U42311 ( .A(n42010), .B(n42011), .Z(n506) );
  NANDN U42312 ( .A(n42012), .B(n42013), .Z(n42011) );
  OR U42313 ( .A(n42014), .B(n42015), .Z(n42013) );
  NAND U42314 ( .A(n42015), .B(n42014), .Z(n42010) );
  XOR U42315 ( .A(n508), .B(n507), .Z(\A1[142] ) );
  XOR U42316 ( .A(n42015), .B(n42016), .Z(n507) );
  XNOR U42317 ( .A(n42014), .B(n42012), .Z(n42016) );
  AND U42318 ( .A(n42017), .B(n42018), .Z(n42012) );
  NANDN U42319 ( .A(n42019), .B(n42020), .Z(n42018) );
  NANDN U42320 ( .A(n42021), .B(n42022), .Z(n42020) );
  NANDN U42321 ( .A(n42022), .B(n42021), .Z(n42017) );
  ANDN U42322 ( .B(B[113]), .A(n54), .Z(n42014) );
  XNOR U42323 ( .A(n41809), .B(n42023), .Z(n42015) );
  XNOR U42324 ( .A(n41808), .B(n41806), .Z(n42023) );
  AND U42325 ( .A(n42024), .B(n42025), .Z(n41806) );
  NANDN U42326 ( .A(n42026), .B(n42027), .Z(n42025) );
  OR U42327 ( .A(n42028), .B(n42029), .Z(n42027) );
  NAND U42328 ( .A(n42029), .B(n42028), .Z(n42024) );
  ANDN U42329 ( .B(B[114]), .A(n55), .Z(n41808) );
  XNOR U42330 ( .A(n41816), .B(n42030), .Z(n41809) );
  XNOR U42331 ( .A(n41815), .B(n41813), .Z(n42030) );
  AND U42332 ( .A(n42031), .B(n42032), .Z(n41813) );
  NANDN U42333 ( .A(n42033), .B(n42034), .Z(n42032) );
  NANDN U42334 ( .A(n42035), .B(n42036), .Z(n42034) );
  NANDN U42335 ( .A(n42036), .B(n42035), .Z(n42031) );
  ANDN U42336 ( .B(B[115]), .A(n56), .Z(n41815) );
  XNOR U42337 ( .A(n41823), .B(n42037), .Z(n41816) );
  XNOR U42338 ( .A(n41822), .B(n41820), .Z(n42037) );
  AND U42339 ( .A(n42038), .B(n42039), .Z(n41820) );
  NANDN U42340 ( .A(n42040), .B(n42041), .Z(n42039) );
  OR U42341 ( .A(n42042), .B(n42043), .Z(n42041) );
  NAND U42342 ( .A(n42043), .B(n42042), .Z(n42038) );
  ANDN U42343 ( .B(B[116]), .A(n57), .Z(n41822) );
  XNOR U42344 ( .A(n41830), .B(n42044), .Z(n41823) );
  XNOR U42345 ( .A(n41829), .B(n41827), .Z(n42044) );
  AND U42346 ( .A(n42045), .B(n42046), .Z(n41827) );
  NANDN U42347 ( .A(n42047), .B(n42048), .Z(n42046) );
  NANDN U42348 ( .A(n42049), .B(n42050), .Z(n42048) );
  NANDN U42349 ( .A(n42050), .B(n42049), .Z(n42045) );
  ANDN U42350 ( .B(B[117]), .A(n58), .Z(n41829) );
  XNOR U42351 ( .A(n41837), .B(n42051), .Z(n41830) );
  XNOR U42352 ( .A(n41836), .B(n41834), .Z(n42051) );
  AND U42353 ( .A(n42052), .B(n42053), .Z(n41834) );
  NANDN U42354 ( .A(n42054), .B(n42055), .Z(n42053) );
  OR U42355 ( .A(n42056), .B(n42057), .Z(n42055) );
  NAND U42356 ( .A(n42057), .B(n42056), .Z(n42052) );
  ANDN U42357 ( .B(B[118]), .A(n59), .Z(n41836) );
  XNOR U42358 ( .A(n41844), .B(n42058), .Z(n41837) );
  XNOR U42359 ( .A(n41843), .B(n41841), .Z(n42058) );
  AND U42360 ( .A(n42059), .B(n42060), .Z(n41841) );
  NANDN U42361 ( .A(n42061), .B(n42062), .Z(n42060) );
  NANDN U42362 ( .A(n42063), .B(n42064), .Z(n42062) );
  NANDN U42363 ( .A(n42064), .B(n42063), .Z(n42059) );
  ANDN U42364 ( .B(B[119]), .A(n60), .Z(n41843) );
  XNOR U42365 ( .A(n41851), .B(n42065), .Z(n41844) );
  XNOR U42366 ( .A(n41850), .B(n41848), .Z(n42065) );
  AND U42367 ( .A(n42066), .B(n42067), .Z(n41848) );
  NANDN U42368 ( .A(n42068), .B(n42069), .Z(n42067) );
  OR U42369 ( .A(n42070), .B(n42071), .Z(n42069) );
  NAND U42370 ( .A(n42071), .B(n42070), .Z(n42066) );
  ANDN U42371 ( .B(B[120]), .A(n61), .Z(n41850) );
  XNOR U42372 ( .A(n41858), .B(n42072), .Z(n41851) );
  XNOR U42373 ( .A(n41857), .B(n41855), .Z(n42072) );
  AND U42374 ( .A(n42073), .B(n42074), .Z(n41855) );
  NANDN U42375 ( .A(n42075), .B(n42076), .Z(n42074) );
  NANDN U42376 ( .A(n42077), .B(n42078), .Z(n42076) );
  NANDN U42377 ( .A(n42078), .B(n42077), .Z(n42073) );
  ANDN U42378 ( .B(B[121]), .A(n62), .Z(n41857) );
  XNOR U42379 ( .A(n41865), .B(n42079), .Z(n41858) );
  XNOR U42380 ( .A(n41864), .B(n41862), .Z(n42079) );
  AND U42381 ( .A(n42080), .B(n42081), .Z(n41862) );
  NANDN U42382 ( .A(n42082), .B(n42083), .Z(n42081) );
  OR U42383 ( .A(n42084), .B(n42085), .Z(n42083) );
  NAND U42384 ( .A(n42085), .B(n42084), .Z(n42080) );
  ANDN U42385 ( .B(B[122]), .A(n63), .Z(n41864) );
  XNOR U42386 ( .A(n41872), .B(n42086), .Z(n41865) );
  XNOR U42387 ( .A(n41871), .B(n41869), .Z(n42086) );
  AND U42388 ( .A(n42087), .B(n42088), .Z(n41869) );
  NANDN U42389 ( .A(n42089), .B(n42090), .Z(n42088) );
  NANDN U42390 ( .A(n42091), .B(n42092), .Z(n42090) );
  NANDN U42391 ( .A(n42092), .B(n42091), .Z(n42087) );
  ANDN U42392 ( .B(B[123]), .A(n64), .Z(n41871) );
  XNOR U42393 ( .A(n41879), .B(n42093), .Z(n41872) );
  XNOR U42394 ( .A(n41878), .B(n41876), .Z(n42093) );
  AND U42395 ( .A(n42094), .B(n42095), .Z(n41876) );
  NANDN U42396 ( .A(n42096), .B(n42097), .Z(n42095) );
  OR U42397 ( .A(n42098), .B(n42099), .Z(n42097) );
  NAND U42398 ( .A(n42099), .B(n42098), .Z(n42094) );
  ANDN U42399 ( .B(B[124]), .A(n65), .Z(n41878) );
  XNOR U42400 ( .A(n41886), .B(n42100), .Z(n41879) );
  XNOR U42401 ( .A(n41885), .B(n41883), .Z(n42100) );
  AND U42402 ( .A(n42101), .B(n42102), .Z(n41883) );
  NANDN U42403 ( .A(n42103), .B(n42104), .Z(n42102) );
  NANDN U42404 ( .A(n42105), .B(n42106), .Z(n42104) );
  NANDN U42405 ( .A(n42106), .B(n42105), .Z(n42101) );
  ANDN U42406 ( .B(B[125]), .A(n66), .Z(n41885) );
  XNOR U42407 ( .A(n41893), .B(n42107), .Z(n41886) );
  XNOR U42408 ( .A(n41892), .B(n41890), .Z(n42107) );
  AND U42409 ( .A(n42108), .B(n42109), .Z(n41890) );
  NANDN U42410 ( .A(n42110), .B(n42111), .Z(n42109) );
  OR U42411 ( .A(n42112), .B(n42113), .Z(n42111) );
  NAND U42412 ( .A(n42113), .B(n42112), .Z(n42108) );
  ANDN U42413 ( .B(B[126]), .A(n67), .Z(n41892) );
  XNOR U42414 ( .A(n41900), .B(n42114), .Z(n41893) );
  XNOR U42415 ( .A(n41899), .B(n41897), .Z(n42114) );
  AND U42416 ( .A(n42115), .B(n42116), .Z(n41897) );
  NANDN U42417 ( .A(n42117), .B(n42118), .Z(n42116) );
  NANDN U42418 ( .A(n42119), .B(n42120), .Z(n42118) );
  NANDN U42419 ( .A(n42120), .B(n42119), .Z(n42115) );
  ANDN U42420 ( .B(B[127]), .A(n68), .Z(n41899) );
  XNOR U42421 ( .A(n41907), .B(n42121), .Z(n41900) );
  XNOR U42422 ( .A(n41906), .B(n41904), .Z(n42121) );
  AND U42423 ( .A(n42122), .B(n42123), .Z(n41904) );
  NANDN U42424 ( .A(n42124), .B(n42125), .Z(n42123) );
  OR U42425 ( .A(n42126), .B(n42127), .Z(n42125) );
  NAND U42426 ( .A(n42127), .B(n42126), .Z(n42122) );
  ANDN U42427 ( .B(B[128]), .A(n69), .Z(n41906) );
  XNOR U42428 ( .A(n41914), .B(n42128), .Z(n41907) );
  XNOR U42429 ( .A(n41913), .B(n41911), .Z(n42128) );
  AND U42430 ( .A(n42129), .B(n42130), .Z(n41911) );
  NANDN U42431 ( .A(n42131), .B(n42132), .Z(n42130) );
  NANDN U42432 ( .A(n42133), .B(n42134), .Z(n42132) );
  NANDN U42433 ( .A(n42134), .B(n42133), .Z(n42129) );
  ANDN U42434 ( .B(B[129]), .A(n70), .Z(n41913) );
  XNOR U42435 ( .A(n41921), .B(n42135), .Z(n41914) );
  XNOR U42436 ( .A(n41920), .B(n41918), .Z(n42135) );
  AND U42437 ( .A(n42136), .B(n42137), .Z(n41918) );
  NANDN U42438 ( .A(n42138), .B(n42139), .Z(n42137) );
  OR U42439 ( .A(n42140), .B(n42141), .Z(n42139) );
  NAND U42440 ( .A(n42141), .B(n42140), .Z(n42136) );
  ANDN U42441 ( .B(B[130]), .A(n71), .Z(n41920) );
  XNOR U42442 ( .A(n41928), .B(n42142), .Z(n41921) );
  XNOR U42443 ( .A(n41927), .B(n41925), .Z(n42142) );
  AND U42444 ( .A(n42143), .B(n42144), .Z(n41925) );
  NANDN U42445 ( .A(n42145), .B(n42146), .Z(n42144) );
  NANDN U42446 ( .A(n42147), .B(n42148), .Z(n42146) );
  NANDN U42447 ( .A(n42148), .B(n42147), .Z(n42143) );
  ANDN U42448 ( .B(B[131]), .A(n72), .Z(n41927) );
  XNOR U42449 ( .A(n41935), .B(n42149), .Z(n41928) );
  XNOR U42450 ( .A(n41934), .B(n41932), .Z(n42149) );
  AND U42451 ( .A(n42150), .B(n42151), .Z(n41932) );
  NANDN U42452 ( .A(n42152), .B(n42153), .Z(n42151) );
  OR U42453 ( .A(n42154), .B(n42155), .Z(n42153) );
  NAND U42454 ( .A(n42155), .B(n42154), .Z(n42150) );
  ANDN U42455 ( .B(B[132]), .A(n73), .Z(n41934) );
  XNOR U42456 ( .A(n41942), .B(n42156), .Z(n41935) );
  XNOR U42457 ( .A(n41941), .B(n41939), .Z(n42156) );
  AND U42458 ( .A(n42157), .B(n42158), .Z(n41939) );
  NANDN U42459 ( .A(n42159), .B(n42160), .Z(n42158) );
  NANDN U42460 ( .A(n42161), .B(n42162), .Z(n42160) );
  NANDN U42461 ( .A(n42162), .B(n42161), .Z(n42157) );
  ANDN U42462 ( .B(B[133]), .A(n74), .Z(n41941) );
  XNOR U42463 ( .A(n41949), .B(n42163), .Z(n41942) );
  XNOR U42464 ( .A(n41948), .B(n41946), .Z(n42163) );
  AND U42465 ( .A(n42164), .B(n42165), .Z(n41946) );
  NANDN U42466 ( .A(n42166), .B(n42167), .Z(n42165) );
  OR U42467 ( .A(n42168), .B(n42169), .Z(n42167) );
  NAND U42468 ( .A(n42169), .B(n42168), .Z(n42164) );
  ANDN U42469 ( .B(B[134]), .A(n75), .Z(n41948) );
  XNOR U42470 ( .A(n41956), .B(n42170), .Z(n41949) );
  XNOR U42471 ( .A(n41955), .B(n41953), .Z(n42170) );
  AND U42472 ( .A(n42171), .B(n42172), .Z(n41953) );
  NANDN U42473 ( .A(n42173), .B(n42174), .Z(n42172) );
  NANDN U42474 ( .A(n42175), .B(n42176), .Z(n42174) );
  NANDN U42475 ( .A(n42176), .B(n42175), .Z(n42171) );
  ANDN U42476 ( .B(B[135]), .A(n76), .Z(n41955) );
  XNOR U42477 ( .A(n41963), .B(n42177), .Z(n41956) );
  XNOR U42478 ( .A(n41962), .B(n41960), .Z(n42177) );
  AND U42479 ( .A(n42178), .B(n42179), .Z(n41960) );
  NANDN U42480 ( .A(n42180), .B(n42181), .Z(n42179) );
  OR U42481 ( .A(n42182), .B(n42183), .Z(n42181) );
  NAND U42482 ( .A(n42183), .B(n42182), .Z(n42178) );
  ANDN U42483 ( .B(B[136]), .A(n77), .Z(n41962) );
  XNOR U42484 ( .A(n41970), .B(n42184), .Z(n41963) );
  XNOR U42485 ( .A(n41969), .B(n41967), .Z(n42184) );
  AND U42486 ( .A(n42185), .B(n42186), .Z(n41967) );
  NANDN U42487 ( .A(n42187), .B(n42188), .Z(n42186) );
  NANDN U42488 ( .A(n42189), .B(n42190), .Z(n42188) );
  NANDN U42489 ( .A(n42190), .B(n42189), .Z(n42185) );
  ANDN U42490 ( .B(B[137]), .A(n78), .Z(n41969) );
  XNOR U42491 ( .A(n41977), .B(n42191), .Z(n41970) );
  XNOR U42492 ( .A(n41976), .B(n41974), .Z(n42191) );
  AND U42493 ( .A(n42192), .B(n42193), .Z(n41974) );
  NANDN U42494 ( .A(n42194), .B(n42195), .Z(n42193) );
  OR U42495 ( .A(n42196), .B(n42197), .Z(n42195) );
  NAND U42496 ( .A(n42197), .B(n42196), .Z(n42192) );
  ANDN U42497 ( .B(B[138]), .A(n79), .Z(n41976) );
  XNOR U42498 ( .A(n41984), .B(n42198), .Z(n41977) );
  XNOR U42499 ( .A(n41983), .B(n41981), .Z(n42198) );
  AND U42500 ( .A(n42199), .B(n42200), .Z(n41981) );
  NANDN U42501 ( .A(n42201), .B(n42202), .Z(n42200) );
  NANDN U42502 ( .A(n42203), .B(n42204), .Z(n42202) );
  NANDN U42503 ( .A(n42204), .B(n42203), .Z(n42199) );
  ANDN U42504 ( .B(B[139]), .A(n80), .Z(n41983) );
  XNOR U42505 ( .A(n41991), .B(n42205), .Z(n41984) );
  XNOR U42506 ( .A(n41990), .B(n41988), .Z(n42205) );
  AND U42507 ( .A(n42206), .B(n42207), .Z(n41988) );
  NANDN U42508 ( .A(n42208), .B(n42209), .Z(n42207) );
  OR U42509 ( .A(n42210), .B(n42211), .Z(n42209) );
  NAND U42510 ( .A(n42211), .B(n42210), .Z(n42206) );
  ANDN U42511 ( .B(B[140]), .A(n81), .Z(n41990) );
  XNOR U42512 ( .A(n41998), .B(n42212), .Z(n41991) );
  XNOR U42513 ( .A(n41997), .B(n41995), .Z(n42212) );
  AND U42514 ( .A(n42213), .B(n42214), .Z(n41995) );
  NANDN U42515 ( .A(n42215), .B(n42216), .Z(n42214) );
  NAND U42516 ( .A(n42217), .B(n42218), .Z(n42216) );
  ANDN U42517 ( .B(B[141]), .A(n82), .Z(n41997) );
  XOR U42518 ( .A(n42004), .B(n42219), .Z(n41998) );
  XNOR U42519 ( .A(n42002), .B(n42005), .Z(n42219) );
  NAND U42520 ( .A(A[2]), .B(B[142]), .Z(n42005) );
  NANDN U42521 ( .A(n42220), .B(n42221), .Z(n42002) );
  AND U42522 ( .A(A[0]), .B(B[143]), .Z(n42221) );
  XNOR U42523 ( .A(n42007), .B(n42222), .Z(n42004) );
  NAND U42524 ( .A(A[0]), .B(B[144]), .Z(n42222) );
  NAND U42525 ( .A(B[143]), .B(A[1]), .Z(n42007) );
  NAND U42526 ( .A(n42223), .B(n42224), .Z(n508) );
  NANDN U42527 ( .A(n42225), .B(n42226), .Z(n42224) );
  OR U42528 ( .A(n42227), .B(n42228), .Z(n42226) );
  NAND U42529 ( .A(n42228), .B(n42227), .Z(n42223) );
  XOR U42530 ( .A(n510), .B(n509), .Z(\A1[141] ) );
  XOR U42531 ( .A(n42228), .B(n42229), .Z(n509) );
  XNOR U42532 ( .A(n42227), .B(n42225), .Z(n42229) );
  AND U42533 ( .A(n42230), .B(n42231), .Z(n42225) );
  NANDN U42534 ( .A(n42232), .B(n42233), .Z(n42231) );
  NANDN U42535 ( .A(n42234), .B(n42235), .Z(n42233) );
  NANDN U42536 ( .A(n42235), .B(n42234), .Z(n42230) );
  ANDN U42537 ( .B(B[112]), .A(n54), .Z(n42227) );
  XNOR U42538 ( .A(n42022), .B(n42236), .Z(n42228) );
  XNOR U42539 ( .A(n42021), .B(n42019), .Z(n42236) );
  AND U42540 ( .A(n42237), .B(n42238), .Z(n42019) );
  NANDN U42541 ( .A(n42239), .B(n42240), .Z(n42238) );
  OR U42542 ( .A(n42241), .B(n42242), .Z(n42240) );
  NAND U42543 ( .A(n42242), .B(n42241), .Z(n42237) );
  ANDN U42544 ( .B(B[113]), .A(n55), .Z(n42021) );
  XNOR U42545 ( .A(n42029), .B(n42243), .Z(n42022) );
  XNOR U42546 ( .A(n42028), .B(n42026), .Z(n42243) );
  AND U42547 ( .A(n42244), .B(n42245), .Z(n42026) );
  NANDN U42548 ( .A(n42246), .B(n42247), .Z(n42245) );
  NANDN U42549 ( .A(n42248), .B(n42249), .Z(n42247) );
  NANDN U42550 ( .A(n42249), .B(n42248), .Z(n42244) );
  ANDN U42551 ( .B(B[114]), .A(n56), .Z(n42028) );
  XNOR U42552 ( .A(n42036), .B(n42250), .Z(n42029) );
  XNOR U42553 ( .A(n42035), .B(n42033), .Z(n42250) );
  AND U42554 ( .A(n42251), .B(n42252), .Z(n42033) );
  NANDN U42555 ( .A(n42253), .B(n42254), .Z(n42252) );
  OR U42556 ( .A(n42255), .B(n42256), .Z(n42254) );
  NAND U42557 ( .A(n42256), .B(n42255), .Z(n42251) );
  ANDN U42558 ( .B(B[115]), .A(n57), .Z(n42035) );
  XNOR U42559 ( .A(n42043), .B(n42257), .Z(n42036) );
  XNOR U42560 ( .A(n42042), .B(n42040), .Z(n42257) );
  AND U42561 ( .A(n42258), .B(n42259), .Z(n42040) );
  NANDN U42562 ( .A(n42260), .B(n42261), .Z(n42259) );
  NANDN U42563 ( .A(n42262), .B(n42263), .Z(n42261) );
  NANDN U42564 ( .A(n42263), .B(n42262), .Z(n42258) );
  ANDN U42565 ( .B(B[116]), .A(n58), .Z(n42042) );
  XNOR U42566 ( .A(n42050), .B(n42264), .Z(n42043) );
  XNOR U42567 ( .A(n42049), .B(n42047), .Z(n42264) );
  AND U42568 ( .A(n42265), .B(n42266), .Z(n42047) );
  NANDN U42569 ( .A(n42267), .B(n42268), .Z(n42266) );
  OR U42570 ( .A(n42269), .B(n42270), .Z(n42268) );
  NAND U42571 ( .A(n42270), .B(n42269), .Z(n42265) );
  ANDN U42572 ( .B(B[117]), .A(n59), .Z(n42049) );
  XNOR U42573 ( .A(n42057), .B(n42271), .Z(n42050) );
  XNOR U42574 ( .A(n42056), .B(n42054), .Z(n42271) );
  AND U42575 ( .A(n42272), .B(n42273), .Z(n42054) );
  NANDN U42576 ( .A(n42274), .B(n42275), .Z(n42273) );
  NANDN U42577 ( .A(n42276), .B(n42277), .Z(n42275) );
  NANDN U42578 ( .A(n42277), .B(n42276), .Z(n42272) );
  ANDN U42579 ( .B(B[118]), .A(n60), .Z(n42056) );
  XNOR U42580 ( .A(n42064), .B(n42278), .Z(n42057) );
  XNOR U42581 ( .A(n42063), .B(n42061), .Z(n42278) );
  AND U42582 ( .A(n42279), .B(n42280), .Z(n42061) );
  NANDN U42583 ( .A(n42281), .B(n42282), .Z(n42280) );
  OR U42584 ( .A(n42283), .B(n42284), .Z(n42282) );
  NAND U42585 ( .A(n42284), .B(n42283), .Z(n42279) );
  ANDN U42586 ( .B(B[119]), .A(n61), .Z(n42063) );
  XNOR U42587 ( .A(n42071), .B(n42285), .Z(n42064) );
  XNOR U42588 ( .A(n42070), .B(n42068), .Z(n42285) );
  AND U42589 ( .A(n42286), .B(n42287), .Z(n42068) );
  NANDN U42590 ( .A(n42288), .B(n42289), .Z(n42287) );
  NANDN U42591 ( .A(n42290), .B(n42291), .Z(n42289) );
  NANDN U42592 ( .A(n42291), .B(n42290), .Z(n42286) );
  ANDN U42593 ( .B(B[120]), .A(n62), .Z(n42070) );
  XNOR U42594 ( .A(n42078), .B(n42292), .Z(n42071) );
  XNOR U42595 ( .A(n42077), .B(n42075), .Z(n42292) );
  AND U42596 ( .A(n42293), .B(n42294), .Z(n42075) );
  NANDN U42597 ( .A(n42295), .B(n42296), .Z(n42294) );
  OR U42598 ( .A(n42297), .B(n42298), .Z(n42296) );
  NAND U42599 ( .A(n42298), .B(n42297), .Z(n42293) );
  ANDN U42600 ( .B(B[121]), .A(n63), .Z(n42077) );
  XNOR U42601 ( .A(n42085), .B(n42299), .Z(n42078) );
  XNOR U42602 ( .A(n42084), .B(n42082), .Z(n42299) );
  AND U42603 ( .A(n42300), .B(n42301), .Z(n42082) );
  NANDN U42604 ( .A(n42302), .B(n42303), .Z(n42301) );
  NANDN U42605 ( .A(n42304), .B(n42305), .Z(n42303) );
  NANDN U42606 ( .A(n42305), .B(n42304), .Z(n42300) );
  ANDN U42607 ( .B(B[122]), .A(n64), .Z(n42084) );
  XNOR U42608 ( .A(n42092), .B(n42306), .Z(n42085) );
  XNOR U42609 ( .A(n42091), .B(n42089), .Z(n42306) );
  AND U42610 ( .A(n42307), .B(n42308), .Z(n42089) );
  NANDN U42611 ( .A(n42309), .B(n42310), .Z(n42308) );
  OR U42612 ( .A(n42311), .B(n42312), .Z(n42310) );
  NAND U42613 ( .A(n42312), .B(n42311), .Z(n42307) );
  ANDN U42614 ( .B(B[123]), .A(n65), .Z(n42091) );
  XNOR U42615 ( .A(n42099), .B(n42313), .Z(n42092) );
  XNOR U42616 ( .A(n42098), .B(n42096), .Z(n42313) );
  AND U42617 ( .A(n42314), .B(n42315), .Z(n42096) );
  NANDN U42618 ( .A(n42316), .B(n42317), .Z(n42315) );
  NANDN U42619 ( .A(n42318), .B(n42319), .Z(n42317) );
  NANDN U42620 ( .A(n42319), .B(n42318), .Z(n42314) );
  ANDN U42621 ( .B(B[124]), .A(n66), .Z(n42098) );
  XNOR U42622 ( .A(n42106), .B(n42320), .Z(n42099) );
  XNOR U42623 ( .A(n42105), .B(n42103), .Z(n42320) );
  AND U42624 ( .A(n42321), .B(n42322), .Z(n42103) );
  NANDN U42625 ( .A(n42323), .B(n42324), .Z(n42322) );
  OR U42626 ( .A(n42325), .B(n42326), .Z(n42324) );
  NAND U42627 ( .A(n42326), .B(n42325), .Z(n42321) );
  ANDN U42628 ( .B(B[125]), .A(n67), .Z(n42105) );
  XNOR U42629 ( .A(n42113), .B(n42327), .Z(n42106) );
  XNOR U42630 ( .A(n42112), .B(n42110), .Z(n42327) );
  AND U42631 ( .A(n42328), .B(n42329), .Z(n42110) );
  NANDN U42632 ( .A(n42330), .B(n42331), .Z(n42329) );
  NANDN U42633 ( .A(n42332), .B(n42333), .Z(n42331) );
  NANDN U42634 ( .A(n42333), .B(n42332), .Z(n42328) );
  ANDN U42635 ( .B(B[126]), .A(n68), .Z(n42112) );
  XNOR U42636 ( .A(n42120), .B(n42334), .Z(n42113) );
  XNOR U42637 ( .A(n42119), .B(n42117), .Z(n42334) );
  AND U42638 ( .A(n42335), .B(n42336), .Z(n42117) );
  NANDN U42639 ( .A(n42337), .B(n42338), .Z(n42336) );
  OR U42640 ( .A(n42339), .B(n42340), .Z(n42338) );
  NAND U42641 ( .A(n42340), .B(n42339), .Z(n42335) );
  ANDN U42642 ( .B(B[127]), .A(n69), .Z(n42119) );
  XNOR U42643 ( .A(n42127), .B(n42341), .Z(n42120) );
  XNOR U42644 ( .A(n42126), .B(n42124), .Z(n42341) );
  AND U42645 ( .A(n42342), .B(n42343), .Z(n42124) );
  NANDN U42646 ( .A(n42344), .B(n42345), .Z(n42343) );
  NANDN U42647 ( .A(n42346), .B(n42347), .Z(n42345) );
  NANDN U42648 ( .A(n42347), .B(n42346), .Z(n42342) );
  ANDN U42649 ( .B(B[128]), .A(n70), .Z(n42126) );
  XNOR U42650 ( .A(n42134), .B(n42348), .Z(n42127) );
  XNOR U42651 ( .A(n42133), .B(n42131), .Z(n42348) );
  AND U42652 ( .A(n42349), .B(n42350), .Z(n42131) );
  NANDN U42653 ( .A(n42351), .B(n42352), .Z(n42350) );
  OR U42654 ( .A(n42353), .B(n42354), .Z(n42352) );
  NAND U42655 ( .A(n42354), .B(n42353), .Z(n42349) );
  ANDN U42656 ( .B(B[129]), .A(n71), .Z(n42133) );
  XNOR U42657 ( .A(n42141), .B(n42355), .Z(n42134) );
  XNOR U42658 ( .A(n42140), .B(n42138), .Z(n42355) );
  AND U42659 ( .A(n42356), .B(n42357), .Z(n42138) );
  NANDN U42660 ( .A(n42358), .B(n42359), .Z(n42357) );
  NANDN U42661 ( .A(n42360), .B(n42361), .Z(n42359) );
  NANDN U42662 ( .A(n42361), .B(n42360), .Z(n42356) );
  ANDN U42663 ( .B(B[130]), .A(n72), .Z(n42140) );
  XNOR U42664 ( .A(n42148), .B(n42362), .Z(n42141) );
  XNOR U42665 ( .A(n42147), .B(n42145), .Z(n42362) );
  AND U42666 ( .A(n42363), .B(n42364), .Z(n42145) );
  NANDN U42667 ( .A(n42365), .B(n42366), .Z(n42364) );
  OR U42668 ( .A(n42367), .B(n42368), .Z(n42366) );
  NAND U42669 ( .A(n42368), .B(n42367), .Z(n42363) );
  ANDN U42670 ( .B(B[131]), .A(n73), .Z(n42147) );
  XNOR U42671 ( .A(n42155), .B(n42369), .Z(n42148) );
  XNOR U42672 ( .A(n42154), .B(n42152), .Z(n42369) );
  AND U42673 ( .A(n42370), .B(n42371), .Z(n42152) );
  NANDN U42674 ( .A(n42372), .B(n42373), .Z(n42371) );
  NANDN U42675 ( .A(n42374), .B(n42375), .Z(n42373) );
  NANDN U42676 ( .A(n42375), .B(n42374), .Z(n42370) );
  ANDN U42677 ( .B(B[132]), .A(n74), .Z(n42154) );
  XNOR U42678 ( .A(n42162), .B(n42376), .Z(n42155) );
  XNOR U42679 ( .A(n42161), .B(n42159), .Z(n42376) );
  AND U42680 ( .A(n42377), .B(n42378), .Z(n42159) );
  NANDN U42681 ( .A(n42379), .B(n42380), .Z(n42378) );
  OR U42682 ( .A(n42381), .B(n42382), .Z(n42380) );
  NAND U42683 ( .A(n42382), .B(n42381), .Z(n42377) );
  ANDN U42684 ( .B(B[133]), .A(n75), .Z(n42161) );
  XNOR U42685 ( .A(n42169), .B(n42383), .Z(n42162) );
  XNOR U42686 ( .A(n42168), .B(n42166), .Z(n42383) );
  AND U42687 ( .A(n42384), .B(n42385), .Z(n42166) );
  NANDN U42688 ( .A(n42386), .B(n42387), .Z(n42385) );
  NANDN U42689 ( .A(n42388), .B(n42389), .Z(n42387) );
  NANDN U42690 ( .A(n42389), .B(n42388), .Z(n42384) );
  ANDN U42691 ( .B(B[134]), .A(n76), .Z(n42168) );
  XNOR U42692 ( .A(n42176), .B(n42390), .Z(n42169) );
  XNOR U42693 ( .A(n42175), .B(n42173), .Z(n42390) );
  AND U42694 ( .A(n42391), .B(n42392), .Z(n42173) );
  NANDN U42695 ( .A(n42393), .B(n42394), .Z(n42392) );
  OR U42696 ( .A(n42395), .B(n42396), .Z(n42394) );
  NAND U42697 ( .A(n42396), .B(n42395), .Z(n42391) );
  ANDN U42698 ( .B(B[135]), .A(n77), .Z(n42175) );
  XNOR U42699 ( .A(n42183), .B(n42397), .Z(n42176) );
  XNOR U42700 ( .A(n42182), .B(n42180), .Z(n42397) );
  AND U42701 ( .A(n42398), .B(n42399), .Z(n42180) );
  NANDN U42702 ( .A(n42400), .B(n42401), .Z(n42399) );
  NANDN U42703 ( .A(n42402), .B(n42403), .Z(n42401) );
  NANDN U42704 ( .A(n42403), .B(n42402), .Z(n42398) );
  ANDN U42705 ( .B(B[136]), .A(n78), .Z(n42182) );
  XNOR U42706 ( .A(n42190), .B(n42404), .Z(n42183) );
  XNOR U42707 ( .A(n42189), .B(n42187), .Z(n42404) );
  AND U42708 ( .A(n42405), .B(n42406), .Z(n42187) );
  NANDN U42709 ( .A(n42407), .B(n42408), .Z(n42406) );
  OR U42710 ( .A(n42409), .B(n42410), .Z(n42408) );
  NAND U42711 ( .A(n42410), .B(n42409), .Z(n42405) );
  ANDN U42712 ( .B(B[137]), .A(n79), .Z(n42189) );
  XNOR U42713 ( .A(n42197), .B(n42411), .Z(n42190) );
  XNOR U42714 ( .A(n42196), .B(n42194), .Z(n42411) );
  AND U42715 ( .A(n42412), .B(n42413), .Z(n42194) );
  NANDN U42716 ( .A(n42414), .B(n42415), .Z(n42413) );
  NANDN U42717 ( .A(n42416), .B(n42417), .Z(n42415) );
  NANDN U42718 ( .A(n42417), .B(n42416), .Z(n42412) );
  ANDN U42719 ( .B(B[138]), .A(n80), .Z(n42196) );
  XNOR U42720 ( .A(n42204), .B(n42418), .Z(n42197) );
  XNOR U42721 ( .A(n42203), .B(n42201), .Z(n42418) );
  AND U42722 ( .A(n42419), .B(n42420), .Z(n42201) );
  NANDN U42723 ( .A(n42421), .B(n42422), .Z(n42420) );
  OR U42724 ( .A(n42423), .B(n42424), .Z(n42422) );
  NAND U42725 ( .A(n42424), .B(n42423), .Z(n42419) );
  ANDN U42726 ( .B(B[139]), .A(n81), .Z(n42203) );
  XNOR U42727 ( .A(n42211), .B(n42425), .Z(n42204) );
  XNOR U42728 ( .A(n42210), .B(n42208), .Z(n42425) );
  AND U42729 ( .A(n42426), .B(n42427), .Z(n42208) );
  NANDN U42730 ( .A(n42428), .B(n42429), .Z(n42427) );
  NAND U42731 ( .A(n42430), .B(n42431), .Z(n42429) );
  ANDN U42732 ( .B(B[140]), .A(n82), .Z(n42210) );
  XOR U42733 ( .A(n42217), .B(n42432), .Z(n42211) );
  XNOR U42734 ( .A(n42215), .B(n42218), .Z(n42432) );
  NAND U42735 ( .A(A[2]), .B(B[141]), .Z(n42218) );
  NANDN U42736 ( .A(n42433), .B(n42434), .Z(n42215) );
  AND U42737 ( .A(A[0]), .B(B[142]), .Z(n42434) );
  XNOR U42738 ( .A(n42220), .B(n42435), .Z(n42217) );
  NAND U42739 ( .A(A[0]), .B(B[143]), .Z(n42435) );
  NAND U42740 ( .A(B[142]), .B(A[1]), .Z(n42220) );
  NAND U42741 ( .A(n42436), .B(n42437), .Z(n510) );
  NANDN U42742 ( .A(n42438), .B(n42439), .Z(n42437) );
  OR U42743 ( .A(n42440), .B(n42441), .Z(n42439) );
  NAND U42744 ( .A(n42441), .B(n42440), .Z(n42436) );
  XOR U42745 ( .A(n512), .B(n511), .Z(\A1[140] ) );
  XOR U42746 ( .A(n42441), .B(n42442), .Z(n511) );
  XNOR U42747 ( .A(n42440), .B(n42438), .Z(n42442) );
  AND U42748 ( .A(n42443), .B(n42444), .Z(n42438) );
  NANDN U42749 ( .A(n42445), .B(n42446), .Z(n42444) );
  NANDN U42750 ( .A(n42447), .B(n42448), .Z(n42446) );
  NANDN U42751 ( .A(n42448), .B(n42447), .Z(n42443) );
  ANDN U42752 ( .B(B[111]), .A(n54), .Z(n42440) );
  XNOR U42753 ( .A(n42235), .B(n42449), .Z(n42441) );
  XNOR U42754 ( .A(n42234), .B(n42232), .Z(n42449) );
  AND U42755 ( .A(n42450), .B(n42451), .Z(n42232) );
  NANDN U42756 ( .A(n42452), .B(n42453), .Z(n42451) );
  OR U42757 ( .A(n42454), .B(n42455), .Z(n42453) );
  NAND U42758 ( .A(n42455), .B(n42454), .Z(n42450) );
  ANDN U42759 ( .B(B[112]), .A(n55), .Z(n42234) );
  XNOR U42760 ( .A(n42242), .B(n42456), .Z(n42235) );
  XNOR U42761 ( .A(n42241), .B(n42239), .Z(n42456) );
  AND U42762 ( .A(n42457), .B(n42458), .Z(n42239) );
  NANDN U42763 ( .A(n42459), .B(n42460), .Z(n42458) );
  NANDN U42764 ( .A(n42461), .B(n42462), .Z(n42460) );
  NANDN U42765 ( .A(n42462), .B(n42461), .Z(n42457) );
  ANDN U42766 ( .B(B[113]), .A(n56), .Z(n42241) );
  XNOR U42767 ( .A(n42249), .B(n42463), .Z(n42242) );
  XNOR U42768 ( .A(n42248), .B(n42246), .Z(n42463) );
  AND U42769 ( .A(n42464), .B(n42465), .Z(n42246) );
  NANDN U42770 ( .A(n42466), .B(n42467), .Z(n42465) );
  OR U42771 ( .A(n42468), .B(n42469), .Z(n42467) );
  NAND U42772 ( .A(n42469), .B(n42468), .Z(n42464) );
  ANDN U42773 ( .B(B[114]), .A(n57), .Z(n42248) );
  XNOR U42774 ( .A(n42256), .B(n42470), .Z(n42249) );
  XNOR U42775 ( .A(n42255), .B(n42253), .Z(n42470) );
  AND U42776 ( .A(n42471), .B(n42472), .Z(n42253) );
  NANDN U42777 ( .A(n42473), .B(n42474), .Z(n42472) );
  NANDN U42778 ( .A(n42475), .B(n42476), .Z(n42474) );
  NANDN U42779 ( .A(n42476), .B(n42475), .Z(n42471) );
  ANDN U42780 ( .B(B[115]), .A(n58), .Z(n42255) );
  XNOR U42781 ( .A(n42263), .B(n42477), .Z(n42256) );
  XNOR U42782 ( .A(n42262), .B(n42260), .Z(n42477) );
  AND U42783 ( .A(n42478), .B(n42479), .Z(n42260) );
  NANDN U42784 ( .A(n42480), .B(n42481), .Z(n42479) );
  OR U42785 ( .A(n42482), .B(n42483), .Z(n42481) );
  NAND U42786 ( .A(n42483), .B(n42482), .Z(n42478) );
  ANDN U42787 ( .B(B[116]), .A(n59), .Z(n42262) );
  XNOR U42788 ( .A(n42270), .B(n42484), .Z(n42263) );
  XNOR U42789 ( .A(n42269), .B(n42267), .Z(n42484) );
  AND U42790 ( .A(n42485), .B(n42486), .Z(n42267) );
  NANDN U42791 ( .A(n42487), .B(n42488), .Z(n42486) );
  NANDN U42792 ( .A(n42489), .B(n42490), .Z(n42488) );
  NANDN U42793 ( .A(n42490), .B(n42489), .Z(n42485) );
  ANDN U42794 ( .B(B[117]), .A(n60), .Z(n42269) );
  XNOR U42795 ( .A(n42277), .B(n42491), .Z(n42270) );
  XNOR U42796 ( .A(n42276), .B(n42274), .Z(n42491) );
  AND U42797 ( .A(n42492), .B(n42493), .Z(n42274) );
  NANDN U42798 ( .A(n42494), .B(n42495), .Z(n42493) );
  OR U42799 ( .A(n42496), .B(n42497), .Z(n42495) );
  NAND U42800 ( .A(n42497), .B(n42496), .Z(n42492) );
  ANDN U42801 ( .B(B[118]), .A(n61), .Z(n42276) );
  XNOR U42802 ( .A(n42284), .B(n42498), .Z(n42277) );
  XNOR U42803 ( .A(n42283), .B(n42281), .Z(n42498) );
  AND U42804 ( .A(n42499), .B(n42500), .Z(n42281) );
  NANDN U42805 ( .A(n42501), .B(n42502), .Z(n42500) );
  NANDN U42806 ( .A(n42503), .B(n42504), .Z(n42502) );
  NANDN U42807 ( .A(n42504), .B(n42503), .Z(n42499) );
  ANDN U42808 ( .B(B[119]), .A(n62), .Z(n42283) );
  XNOR U42809 ( .A(n42291), .B(n42505), .Z(n42284) );
  XNOR U42810 ( .A(n42290), .B(n42288), .Z(n42505) );
  AND U42811 ( .A(n42506), .B(n42507), .Z(n42288) );
  NANDN U42812 ( .A(n42508), .B(n42509), .Z(n42507) );
  OR U42813 ( .A(n42510), .B(n42511), .Z(n42509) );
  NAND U42814 ( .A(n42511), .B(n42510), .Z(n42506) );
  ANDN U42815 ( .B(B[120]), .A(n63), .Z(n42290) );
  XNOR U42816 ( .A(n42298), .B(n42512), .Z(n42291) );
  XNOR U42817 ( .A(n42297), .B(n42295), .Z(n42512) );
  AND U42818 ( .A(n42513), .B(n42514), .Z(n42295) );
  NANDN U42819 ( .A(n42515), .B(n42516), .Z(n42514) );
  NANDN U42820 ( .A(n42517), .B(n42518), .Z(n42516) );
  NANDN U42821 ( .A(n42518), .B(n42517), .Z(n42513) );
  ANDN U42822 ( .B(B[121]), .A(n64), .Z(n42297) );
  XNOR U42823 ( .A(n42305), .B(n42519), .Z(n42298) );
  XNOR U42824 ( .A(n42304), .B(n42302), .Z(n42519) );
  AND U42825 ( .A(n42520), .B(n42521), .Z(n42302) );
  NANDN U42826 ( .A(n42522), .B(n42523), .Z(n42521) );
  OR U42827 ( .A(n42524), .B(n42525), .Z(n42523) );
  NAND U42828 ( .A(n42525), .B(n42524), .Z(n42520) );
  ANDN U42829 ( .B(B[122]), .A(n65), .Z(n42304) );
  XNOR U42830 ( .A(n42312), .B(n42526), .Z(n42305) );
  XNOR U42831 ( .A(n42311), .B(n42309), .Z(n42526) );
  AND U42832 ( .A(n42527), .B(n42528), .Z(n42309) );
  NANDN U42833 ( .A(n42529), .B(n42530), .Z(n42528) );
  NANDN U42834 ( .A(n42531), .B(n42532), .Z(n42530) );
  NANDN U42835 ( .A(n42532), .B(n42531), .Z(n42527) );
  ANDN U42836 ( .B(B[123]), .A(n66), .Z(n42311) );
  XNOR U42837 ( .A(n42319), .B(n42533), .Z(n42312) );
  XNOR U42838 ( .A(n42318), .B(n42316), .Z(n42533) );
  AND U42839 ( .A(n42534), .B(n42535), .Z(n42316) );
  NANDN U42840 ( .A(n42536), .B(n42537), .Z(n42535) );
  OR U42841 ( .A(n42538), .B(n42539), .Z(n42537) );
  NAND U42842 ( .A(n42539), .B(n42538), .Z(n42534) );
  ANDN U42843 ( .B(B[124]), .A(n67), .Z(n42318) );
  XNOR U42844 ( .A(n42326), .B(n42540), .Z(n42319) );
  XNOR U42845 ( .A(n42325), .B(n42323), .Z(n42540) );
  AND U42846 ( .A(n42541), .B(n42542), .Z(n42323) );
  NANDN U42847 ( .A(n42543), .B(n42544), .Z(n42542) );
  NANDN U42848 ( .A(n42545), .B(n42546), .Z(n42544) );
  NANDN U42849 ( .A(n42546), .B(n42545), .Z(n42541) );
  ANDN U42850 ( .B(B[125]), .A(n68), .Z(n42325) );
  XNOR U42851 ( .A(n42333), .B(n42547), .Z(n42326) );
  XNOR U42852 ( .A(n42332), .B(n42330), .Z(n42547) );
  AND U42853 ( .A(n42548), .B(n42549), .Z(n42330) );
  NANDN U42854 ( .A(n42550), .B(n42551), .Z(n42549) );
  OR U42855 ( .A(n42552), .B(n42553), .Z(n42551) );
  NAND U42856 ( .A(n42553), .B(n42552), .Z(n42548) );
  ANDN U42857 ( .B(B[126]), .A(n69), .Z(n42332) );
  XNOR U42858 ( .A(n42340), .B(n42554), .Z(n42333) );
  XNOR U42859 ( .A(n42339), .B(n42337), .Z(n42554) );
  AND U42860 ( .A(n42555), .B(n42556), .Z(n42337) );
  NANDN U42861 ( .A(n42557), .B(n42558), .Z(n42556) );
  NANDN U42862 ( .A(n42559), .B(n42560), .Z(n42558) );
  NANDN U42863 ( .A(n42560), .B(n42559), .Z(n42555) );
  ANDN U42864 ( .B(B[127]), .A(n70), .Z(n42339) );
  XNOR U42865 ( .A(n42347), .B(n42561), .Z(n42340) );
  XNOR U42866 ( .A(n42346), .B(n42344), .Z(n42561) );
  AND U42867 ( .A(n42562), .B(n42563), .Z(n42344) );
  NANDN U42868 ( .A(n42564), .B(n42565), .Z(n42563) );
  OR U42869 ( .A(n42566), .B(n42567), .Z(n42565) );
  NAND U42870 ( .A(n42567), .B(n42566), .Z(n42562) );
  ANDN U42871 ( .B(B[128]), .A(n71), .Z(n42346) );
  XNOR U42872 ( .A(n42354), .B(n42568), .Z(n42347) );
  XNOR U42873 ( .A(n42353), .B(n42351), .Z(n42568) );
  AND U42874 ( .A(n42569), .B(n42570), .Z(n42351) );
  NANDN U42875 ( .A(n42571), .B(n42572), .Z(n42570) );
  NANDN U42876 ( .A(n42573), .B(n42574), .Z(n42572) );
  NANDN U42877 ( .A(n42574), .B(n42573), .Z(n42569) );
  ANDN U42878 ( .B(B[129]), .A(n72), .Z(n42353) );
  XNOR U42879 ( .A(n42361), .B(n42575), .Z(n42354) );
  XNOR U42880 ( .A(n42360), .B(n42358), .Z(n42575) );
  AND U42881 ( .A(n42576), .B(n42577), .Z(n42358) );
  NANDN U42882 ( .A(n42578), .B(n42579), .Z(n42577) );
  OR U42883 ( .A(n42580), .B(n42581), .Z(n42579) );
  NAND U42884 ( .A(n42581), .B(n42580), .Z(n42576) );
  ANDN U42885 ( .B(B[130]), .A(n73), .Z(n42360) );
  XNOR U42886 ( .A(n42368), .B(n42582), .Z(n42361) );
  XNOR U42887 ( .A(n42367), .B(n42365), .Z(n42582) );
  AND U42888 ( .A(n42583), .B(n42584), .Z(n42365) );
  NANDN U42889 ( .A(n42585), .B(n42586), .Z(n42584) );
  NANDN U42890 ( .A(n42587), .B(n42588), .Z(n42586) );
  NANDN U42891 ( .A(n42588), .B(n42587), .Z(n42583) );
  ANDN U42892 ( .B(B[131]), .A(n74), .Z(n42367) );
  XNOR U42893 ( .A(n42375), .B(n42589), .Z(n42368) );
  XNOR U42894 ( .A(n42374), .B(n42372), .Z(n42589) );
  AND U42895 ( .A(n42590), .B(n42591), .Z(n42372) );
  NANDN U42896 ( .A(n42592), .B(n42593), .Z(n42591) );
  OR U42897 ( .A(n42594), .B(n42595), .Z(n42593) );
  NAND U42898 ( .A(n42595), .B(n42594), .Z(n42590) );
  ANDN U42899 ( .B(B[132]), .A(n75), .Z(n42374) );
  XNOR U42900 ( .A(n42382), .B(n42596), .Z(n42375) );
  XNOR U42901 ( .A(n42381), .B(n42379), .Z(n42596) );
  AND U42902 ( .A(n42597), .B(n42598), .Z(n42379) );
  NANDN U42903 ( .A(n42599), .B(n42600), .Z(n42598) );
  NANDN U42904 ( .A(n42601), .B(n42602), .Z(n42600) );
  NANDN U42905 ( .A(n42602), .B(n42601), .Z(n42597) );
  ANDN U42906 ( .B(B[133]), .A(n76), .Z(n42381) );
  XNOR U42907 ( .A(n42389), .B(n42603), .Z(n42382) );
  XNOR U42908 ( .A(n42388), .B(n42386), .Z(n42603) );
  AND U42909 ( .A(n42604), .B(n42605), .Z(n42386) );
  NANDN U42910 ( .A(n42606), .B(n42607), .Z(n42605) );
  OR U42911 ( .A(n42608), .B(n42609), .Z(n42607) );
  NAND U42912 ( .A(n42609), .B(n42608), .Z(n42604) );
  ANDN U42913 ( .B(B[134]), .A(n77), .Z(n42388) );
  XNOR U42914 ( .A(n42396), .B(n42610), .Z(n42389) );
  XNOR U42915 ( .A(n42395), .B(n42393), .Z(n42610) );
  AND U42916 ( .A(n42611), .B(n42612), .Z(n42393) );
  NANDN U42917 ( .A(n42613), .B(n42614), .Z(n42612) );
  NANDN U42918 ( .A(n42615), .B(n42616), .Z(n42614) );
  NANDN U42919 ( .A(n42616), .B(n42615), .Z(n42611) );
  ANDN U42920 ( .B(B[135]), .A(n78), .Z(n42395) );
  XNOR U42921 ( .A(n42403), .B(n42617), .Z(n42396) );
  XNOR U42922 ( .A(n42402), .B(n42400), .Z(n42617) );
  AND U42923 ( .A(n42618), .B(n42619), .Z(n42400) );
  NANDN U42924 ( .A(n42620), .B(n42621), .Z(n42619) );
  OR U42925 ( .A(n42622), .B(n42623), .Z(n42621) );
  NAND U42926 ( .A(n42623), .B(n42622), .Z(n42618) );
  ANDN U42927 ( .B(B[136]), .A(n79), .Z(n42402) );
  XNOR U42928 ( .A(n42410), .B(n42624), .Z(n42403) );
  XNOR U42929 ( .A(n42409), .B(n42407), .Z(n42624) );
  AND U42930 ( .A(n42625), .B(n42626), .Z(n42407) );
  NANDN U42931 ( .A(n42627), .B(n42628), .Z(n42626) );
  NANDN U42932 ( .A(n42629), .B(n42630), .Z(n42628) );
  NANDN U42933 ( .A(n42630), .B(n42629), .Z(n42625) );
  ANDN U42934 ( .B(B[137]), .A(n80), .Z(n42409) );
  XNOR U42935 ( .A(n42417), .B(n42631), .Z(n42410) );
  XNOR U42936 ( .A(n42416), .B(n42414), .Z(n42631) );
  AND U42937 ( .A(n42632), .B(n42633), .Z(n42414) );
  NANDN U42938 ( .A(n42634), .B(n42635), .Z(n42633) );
  OR U42939 ( .A(n42636), .B(n42637), .Z(n42635) );
  NAND U42940 ( .A(n42637), .B(n42636), .Z(n42632) );
  ANDN U42941 ( .B(B[138]), .A(n81), .Z(n42416) );
  XNOR U42942 ( .A(n42424), .B(n42638), .Z(n42417) );
  XNOR U42943 ( .A(n42423), .B(n42421), .Z(n42638) );
  AND U42944 ( .A(n42639), .B(n42640), .Z(n42421) );
  NANDN U42945 ( .A(n42641), .B(n42642), .Z(n42640) );
  NAND U42946 ( .A(n42643), .B(n42644), .Z(n42642) );
  ANDN U42947 ( .B(B[139]), .A(n82), .Z(n42423) );
  XOR U42948 ( .A(n42430), .B(n42645), .Z(n42424) );
  XNOR U42949 ( .A(n42428), .B(n42431), .Z(n42645) );
  NAND U42950 ( .A(A[2]), .B(B[140]), .Z(n42431) );
  NANDN U42951 ( .A(n42646), .B(n42647), .Z(n42428) );
  AND U42952 ( .A(A[0]), .B(B[141]), .Z(n42647) );
  XNOR U42953 ( .A(n42433), .B(n42648), .Z(n42430) );
  NAND U42954 ( .A(A[0]), .B(B[142]), .Z(n42648) );
  NAND U42955 ( .A(B[141]), .B(A[1]), .Z(n42433) );
  NAND U42956 ( .A(n42649), .B(n42650), .Z(n512) );
  NANDN U42957 ( .A(n42651), .B(n42652), .Z(n42650) );
  OR U42958 ( .A(n42653), .B(n42654), .Z(n42652) );
  NAND U42959 ( .A(n42654), .B(n42653), .Z(n42649) );
  XOR U42960 ( .A(n40429), .B(n42655), .Z(\A1[13] ) );
  XNOR U42961 ( .A(n40428), .B(n40426), .Z(n42655) );
  AND U42962 ( .A(n42656), .B(n42657), .Z(n40426) );
  NAND U42963 ( .A(n42658), .B(n42659), .Z(n42657) );
  NANDN U42964 ( .A(n42660), .B(n42661), .Z(n42658) );
  NANDN U42965 ( .A(n42661), .B(n42660), .Z(n42656) );
  ANDN U42966 ( .B(B[0]), .A(n70), .Z(n40428) );
  XNOR U42967 ( .A(n40436), .B(n42662), .Z(n40429) );
  XNOR U42968 ( .A(n40435), .B(n40433), .Z(n42662) );
  AND U42969 ( .A(n42663), .B(n42664), .Z(n40433) );
  NANDN U42970 ( .A(n42665), .B(n42666), .Z(n42664) );
  OR U42971 ( .A(n42667), .B(n42668), .Z(n42666) );
  NAND U42972 ( .A(n42668), .B(n42667), .Z(n42663) );
  ANDN U42973 ( .B(B[1]), .A(n71), .Z(n40435) );
  XNOR U42974 ( .A(n40443), .B(n42669), .Z(n40436) );
  XNOR U42975 ( .A(n40442), .B(n40440), .Z(n42669) );
  AND U42976 ( .A(n42670), .B(n42671), .Z(n40440) );
  NANDN U42977 ( .A(n42672), .B(n42673), .Z(n42671) );
  NANDN U42978 ( .A(n42674), .B(n42675), .Z(n42673) );
  NANDN U42979 ( .A(n42675), .B(n42674), .Z(n42670) );
  ANDN U42980 ( .B(B[2]), .A(n72), .Z(n40442) );
  XNOR U42981 ( .A(n40450), .B(n42676), .Z(n40443) );
  XNOR U42982 ( .A(n40449), .B(n40447), .Z(n42676) );
  AND U42983 ( .A(n42677), .B(n42678), .Z(n40447) );
  NANDN U42984 ( .A(n42679), .B(n42680), .Z(n42678) );
  OR U42985 ( .A(n42681), .B(n42682), .Z(n42680) );
  NAND U42986 ( .A(n42682), .B(n42681), .Z(n42677) );
  ANDN U42987 ( .B(B[3]), .A(n73), .Z(n40449) );
  XNOR U42988 ( .A(n40457), .B(n42683), .Z(n40450) );
  XNOR U42989 ( .A(n40456), .B(n40454), .Z(n42683) );
  AND U42990 ( .A(n42684), .B(n42685), .Z(n40454) );
  NANDN U42991 ( .A(n42686), .B(n42687), .Z(n42685) );
  NANDN U42992 ( .A(n42688), .B(n42689), .Z(n42687) );
  NANDN U42993 ( .A(n42689), .B(n42688), .Z(n42684) );
  ANDN U42994 ( .B(B[4]), .A(n74), .Z(n40456) );
  XNOR U42995 ( .A(n40464), .B(n42690), .Z(n40457) );
  XNOR U42996 ( .A(n40463), .B(n40461), .Z(n42690) );
  AND U42997 ( .A(n42691), .B(n42692), .Z(n40461) );
  NANDN U42998 ( .A(n42693), .B(n42694), .Z(n42692) );
  OR U42999 ( .A(n42695), .B(n42696), .Z(n42694) );
  NAND U43000 ( .A(n42696), .B(n42695), .Z(n42691) );
  ANDN U43001 ( .B(B[5]), .A(n75), .Z(n40463) );
  XNOR U43002 ( .A(n40471), .B(n42697), .Z(n40464) );
  XNOR U43003 ( .A(n40470), .B(n40468), .Z(n42697) );
  AND U43004 ( .A(n42698), .B(n42699), .Z(n40468) );
  NANDN U43005 ( .A(n42700), .B(n42701), .Z(n42699) );
  NANDN U43006 ( .A(n42702), .B(n42703), .Z(n42701) );
  NANDN U43007 ( .A(n42703), .B(n42702), .Z(n42698) );
  ANDN U43008 ( .B(B[6]), .A(n76), .Z(n40470) );
  XNOR U43009 ( .A(n40478), .B(n42704), .Z(n40471) );
  XNOR U43010 ( .A(n40477), .B(n40475), .Z(n42704) );
  AND U43011 ( .A(n42705), .B(n42706), .Z(n40475) );
  NANDN U43012 ( .A(n42707), .B(n42708), .Z(n42706) );
  OR U43013 ( .A(n42709), .B(n42710), .Z(n42708) );
  NAND U43014 ( .A(n42710), .B(n42709), .Z(n42705) );
  ANDN U43015 ( .B(B[7]), .A(n77), .Z(n40477) );
  XNOR U43016 ( .A(n40485), .B(n42711), .Z(n40478) );
  XNOR U43017 ( .A(n40484), .B(n40482), .Z(n42711) );
  AND U43018 ( .A(n42712), .B(n42713), .Z(n40482) );
  NANDN U43019 ( .A(n42714), .B(n42715), .Z(n42713) );
  NANDN U43020 ( .A(n42716), .B(n42717), .Z(n42715) );
  NANDN U43021 ( .A(n42717), .B(n42716), .Z(n42712) );
  ANDN U43022 ( .B(B[8]), .A(n78), .Z(n40484) );
  XNOR U43023 ( .A(n40492), .B(n42718), .Z(n40485) );
  XNOR U43024 ( .A(n40491), .B(n40489), .Z(n42718) );
  AND U43025 ( .A(n42719), .B(n42720), .Z(n40489) );
  NANDN U43026 ( .A(n42721), .B(n42722), .Z(n42720) );
  OR U43027 ( .A(n42723), .B(n42724), .Z(n42722) );
  NAND U43028 ( .A(n42724), .B(n42723), .Z(n42719) );
  ANDN U43029 ( .B(B[9]), .A(n79), .Z(n40491) );
  XNOR U43030 ( .A(n40499), .B(n42725), .Z(n40492) );
  XNOR U43031 ( .A(n40498), .B(n40496), .Z(n42725) );
  AND U43032 ( .A(n42726), .B(n42727), .Z(n40496) );
  NANDN U43033 ( .A(n42728), .B(n42729), .Z(n42727) );
  NANDN U43034 ( .A(n42730), .B(n42731), .Z(n42729) );
  NANDN U43035 ( .A(n42731), .B(n42730), .Z(n42726) );
  ANDN U43036 ( .B(B[10]), .A(n80), .Z(n40498) );
  XNOR U43037 ( .A(n40506), .B(n42732), .Z(n40499) );
  XNOR U43038 ( .A(n40505), .B(n40503), .Z(n42732) );
  AND U43039 ( .A(n42733), .B(n42734), .Z(n40503) );
  NANDN U43040 ( .A(n42735), .B(n42736), .Z(n42734) );
  OR U43041 ( .A(n42737), .B(n42738), .Z(n42736) );
  NAND U43042 ( .A(n42738), .B(n42737), .Z(n42733) );
  ANDN U43043 ( .B(B[11]), .A(n81), .Z(n40505) );
  XNOR U43044 ( .A(n40513), .B(n42739), .Z(n40506) );
  XNOR U43045 ( .A(n40512), .B(n40510), .Z(n42739) );
  AND U43046 ( .A(n42740), .B(n42741), .Z(n40510) );
  NANDN U43047 ( .A(n42742), .B(n42743), .Z(n42741) );
  NAND U43048 ( .A(n42744), .B(n42745), .Z(n42743) );
  ANDN U43049 ( .B(B[12]), .A(n82), .Z(n40512) );
  XOR U43050 ( .A(n40519), .B(n42746), .Z(n40513) );
  XNOR U43051 ( .A(n40517), .B(n40520), .Z(n42746) );
  NAND U43052 ( .A(A[2]), .B(B[13]), .Z(n40520) );
  NANDN U43053 ( .A(n42747), .B(n42748), .Z(n40517) );
  AND U43054 ( .A(A[0]), .B(B[14]), .Z(n42748) );
  XNOR U43055 ( .A(n40522), .B(n42749), .Z(n40519) );
  NAND U43056 ( .A(A[0]), .B(B[15]), .Z(n42749) );
  NAND U43057 ( .A(B[14]), .B(A[1]), .Z(n40522) );
  XOR U43058 ( .A(n514), .B(n513), .Z(\A1[139] ) );
  XOR U43059 ( .A(n42654), .B(n42750), .Z(n513) );
  XNOR U43060 ( .A(n42653), .B(n42651), .Z(n42750) );
  AND U43061 ( .A(n42751), .B(n42752), .Z(n42651) );
  NANDN U43062 ( .A(n42753), .B(n42754), .Z(n42752) );
  NANDN U43063 ( .A(n42755), .B(n42756), .Z(n42754) );
  NANDN U43064 ( .A(n42756), .B(n42755), .Z(n42751) );
  ANDN U43065 ( .B(B[110]), .A(n54), .Z(n42653) );
  XNOR U43066 ( .A(n42448), .B(n42757), .Z(n42654) );
  XNOR U43067 ( .A(n42447), .B(n42445), .Z(n42757) );
  AND U43068 ( .A(n42758), .B(n42759), .Z(n42445) );
  NANDN U43069 ( .A(n42760), .B(n42761), .Z(n42759) );
  OR U43070 ( .A(n42762), .B(n42763), .Z(n42761) );
  NAND U43071 ( .A(n42763), .B(n42762), .Z(n42758) );
  ANDN U43072 ( .B(B[111]), .A(n55), .Z(n42447) );
  XNOR U43073 ( .A(n42455), .B(n42764), .Z(n42448) );
  XNOR U43074 ( .A(n42454), .B(n42452), .Z(n42764) );
  AND U43075 ( .A(n42765), .B(n42766), .Z(n42452) );
  NANDN U43076 ( .A(n42767), .B(n42768), .Z(n42766) );
  NANDN U43077 ( .A(n42769), .B(n42770), .Z(n42768) );
  NANDN U43078 ( .A(n42770), .B(n42769), .Z(n42765) );
  ANDN U43079 ( .B(B[112]), .A(n56), .Z(n42454) );
  XNOR U43080 ( .A(n42462), .B(n42771), .Z(n42455) );
  XNOR U43081 ( .A(n42461), .B(n42459), .Z(n42771) );
  AND U43082 ( .A(n42772), .B(n42773), .Z(n42459) );
  NANDN U43083 ( .A(n42774), .B(n42775), .Z(n42773) );
  OR U43084 ( .A(n42776), .B(n42777), .Z(n42775) );
  NAND U43085 ( .A(n42777), .B(n42776), .Z(n42772) );
  ANDN U43086 ( .B(B[113]), .A(n57), .Z(n42461) );
  XNOR U43087 ( .A(n42469), .B(n42778), .Z(n42462) );
  XNOR U43088 ( .A(n42468), .B(n42466), .Z(n42778) );
  AND U43089 ( .A(n42779), .B(n42780), .Z(n42466) );
  NANDN U43090 ( .A(n42781), .B(n42782), .Z(n42780) );
  NANDN U43091 ( .A(n42783), .B(n42784), .Z(n42782) );
  NANDN U43092 ( .A(n42784), .B(n42783), .Z(n42779) );
  ANDN U43093 ( .B(B[114]), .A(n58), .Z(n42468) );
  XNOR U43094 ( .A(n42476), .B(n42785), .Z(n42469) );
  XNOR U43095 ( .A(n42475), .B(n42473), .Z(n42785) );
  AND U43096 ( .A(n42786), .B(n42787), .Z(n42473) );
  NANDN U43097 ( .A(n42788), .B(n42789), .Z(n42787) );
  OR U43098 ( .A(n42790), .B(n42791), .Z(n42789) );
  NAND U43099 ( .A(n42791), .B(n42790), .Z(n42786) );
  ANDN U43100 ( .B(B[115]), .A(n59), .Z(n42475) );
  XNOR U43101 ( .A(n42483), .B(n42792), .Z(n42476) );
  XNOR U43102 ( .A(n42482), .B(n42480), .Z(n42792) );
  AND U43103 ( .A(n42793), .B(n42794), .Z(n42480) );
  NANDN U43104 ( .A(n42795), .B(n42796), .Z(n42794) );
  NANDN U43105 ( .A(n42797), .B(n42798), .Z(n42796) );
  NANDN U43106 ( .A(n42798), .B(n42797), .Z(n42793) );
  ANDN U43107 ( .B(B[116]), .A(n60), .Z(n42482) );
  XNOR U43108 ( .A(n42490), .B(n42799), .Z(n42483) );
  XNOR U43109 ( .A(n42489), .B(n42487), .Z(n42799) );
  AND U43110 ( .A(n42800), .B(n42801), .Z(n42487) );
  NANDN U43111 ( .A(n42802), .B(n42803), .Z(n42801) );
  OR U43112 ( .A(n42804), .B(n42805), .Z(n42803) );
  NAND U43113 ( .A(n42805), .B(n42804), .Z(n42800) );
  ANDN U43114 ( .B(B[117]), .A(n61), .Z(n42489) );
  XNOR U43115 ( .A(n42497), .B(n42806), .Z(n42490) );
  XNOR U43116 ( .A(n42496), .B(n42494), .Z(n42806) );
  AND U43117 ( .A(n42807), .B(n42808), .Z(n42494) );
  NANDN U43118 ( .A(n42809), .B(n42810), .Z(n42808) );
  NANDN U43119 ( .A(n42811), .B(n42812), .Z(n42810) );
  NANDN U43120 ( .A(n42812), .B(n42811), .Z(n42807) );
  ANDN U43121 ( .B(B[118]), .A(n62), .Z(n42496) );
  XNOR U43122 ( .A(n42504), .B(n42813), .Z(n42497) );
  XNOR U43123 ( .A(n42503), .B(n42501), .Z(n42813) );
  AND U43124 ( .A(n42814), .B(n42815), .Z(n42501) );
  NANDN U43125 ( .A(n42816), .B(n42817), .Z(n42815) );
  OR U43126 ( .A(n42818), .B(n42819), .Z(n42817) );
  NAND U43127 ( .A(n42819), .B(n42818), .Z(n42814) );
  ANDN U43128 ( .B(B[119]), .A(n63), .Z(n42503) );
  XNOR U43129 ( .A(n42511), .B(n42820), .Z(n42504) );
  XNOR U43130 ( .A(n42510), .B(n42508), .Z(n42820) );
  AND U43131 ( .A(n42821), .B(n42822), .Z(n42508) );
  NANDN U43132 ( .A(n42823), .B(n42824), .Z(n42822) );
  NANDN U43133 ( .A(n42825), .B(n42826), .Z(n42824) );
  NANDN U43134 ( .A(n42826), .B(n42825), .Z(n42821) );
  ANDN U43135 ( .B(B[120]), .A(n64), .Z(n42510) );
  XNOR U43136 ( .A(n42518), .B(n42827), .Z(n42511) );
  XNOR U43137 ( .A(n42517), .B(n42515), .Z(n42827) );
  AND U43138 ( .A(n42828), .B(n42829), .Z(n42515) );
  NANDN U43139 ( .A(n42830), .B(n42831), .Z(n42829) );
  OR U43140 ( .A(n42832), .B(n42833), .Z(n42831) );
  NAND U43141 ( .A(n42833), .B(n42832), .Z(n42828) );
  ANDN U43142 ( .B(B[121]), .A(n65), .Z(n42517) );
  XNOR U43143 ( .A(n42525), .B(n42834), .Z(n42518) );
  XNOR U43144 ( .A(n42524), .B(n42522), .Z(n42834) );
  AND U43145 ( .A(n42835), .B(n42836), .Z(n42522) );
  NANDN U43146 ( .A(n42837), .B(n42838), .Z(n42836) );
  NANDN U43147 ( .A(n42839), .B(n42840), .Z(n42838) );
  NANDN U43148 ( .A(n42840), .B(n42839), .Z(n42835) );
  ANDN U43149 ( .B(B[122]), .A(n66), .Z(n42524) );
  XNOR U43150 ( .A(n42532), .B(n42841), .Z(n42525) );
  XNOR U43151 ( .A(n42531), .B(n42529), .Z(n42841) );
  AND U43152 ( .A(n42842), .B(n42843), .Z(n42529) );
  NANDN U43153 ( .A(n42844), .B(n42845), .Z(n42843) );
  OR U43154 ( .A(n42846), .B(n42847), .Z(n42845) );
  NAND U43155 ( .A(n42847), .B(n42846), .Z(n42842) );
  ANDN U43156 ( .B(B[123]), .A(n67), .Z(n42531) );
  XNOR U43157 ( .A(n42539), .B(n42848), .Z(n42532) );
  XNOR U43158 ( .A(n42538), .B(n42536), .Z(n42848) );
  AND U43159 ( .A(n42849), .B(n42850), .Z(n42536) );
  NANDN U43160 ( .A(n42851), .B(n42852), .Z(n42850) );
  NANDN U43161 ( .A(n42853), .B(n42854), .Z(n42852) );
  NANDN U43162 ( .A(n42854), .B(n42853), .Z(n42849) );
  ANDN U43163 ( .B(B[124]), .A(n68), .Z(n42538) );
  XNOR U43164 ( .A(n42546), .B(n42855), .Z(n42539) );
  XNOR U43165 ( .A(n42545), .B(n42543), .Z(n42855) );
  AND U43166 ( .A(n42856), .B(n42857), .Z(n42543) );
  NANDN U43167 ( .A(n42858), .B(n42859), .Z(n42857) );
  OR U43168 ( .A(n42860), .B(n42861), .Z(n42859) );
  NAND U43169 ( .A(n42861), .B(n42860), .Z(n42856) );
  ANDN U43170 ( .B(B[125]), .A(n69), .Z(n42545) );
  XNOR U43171 ( .A(n42553), .B(n42862), .Z(n42546) );
  XNOR U43172 ( .A(n42552), .B(n42550), .Z(n42862) );
  AND U43173 ( .A(n42863), .B(n42864), .Z(n42550) );
  NANDN U43174 ( .A(n42865), .B(n42866), .Z(n42864) );
  NANDN U43175 ( .A(n42867), .B(n42868), .Z(n42866) );
  NANDN U43176 ( .A(n42868), .B(n42867), .Z(n42863) );
  ANDN U43177 ( .B(B[126]), .A(n70), .Z(n42552) );
  XNOR U43178 ( .A(n42560), .B(n42869), .Z(n42553) );
  XNOR U43179 ( .A(n42559), .B(n42557), .Z(n42869) );
  AND U43180 ( .A(n42870), .B(n42871), .Z(n42557) );
  NANDN U43181 ( .A(n42872), .B(n42873), .Z(n42871) );
  OR U43182 ( .A(n42874), .B(n42875), .Z(n42873) );
  NAND U43183 ( .A(n42875), .B(n42874), .Z(n42870) );
  ANDN U43184 ( .B(B[127]), .A(n71), .Z(n42559) );
  XNOR U43185 ( .A(n42567), .B(n42876), .Z(n42560) );
  XNOR U43186 ( .A(n42566), .B(n42564), .Z(n42876) );
  AND U43187 ( .A(n42877), .B(n42878), .Z(n42564) );
  NANDN U43188 ( .A(n42879), .B(n42880), .Z(n42878) );
  NANDN U43189 ( .A(n42881), .B(n42882), .Z(n42880) );
  NANDN U43190 ( .A(n42882), .B(n42881), .Z(n42877) );
  ANDN U43191 ( .B(B[128]), .A(n72), .Z(n42566) );
  XNOR U43192 ( .A(n42574), .B(n42883), .Z(n42567) );
  XNOR U43193 ( .A(n42573), .B(n42571), .Z(n42883) );
  AND U43194 ( .A(n42884), .B(n42885), .Z(n42571) );
  NANDN U43195 ( .A(n42886), .B(n42887), .Z(n42885) );
  OR U43196 ( .A(n42888), .B(n42889), .Z(n42887) );
  NAND U43197 ( .A(n42889), .B(n42888), .Z(n42884) );
  ANDN U43198 ( .B(B[129]), .A(n73), .Z(n42573) );
  XNOR U43199 ( .A(n42581), .B(n42890), .Z(n42574) );
  XNOR U43200 ( .A(n42580), .B(n42578), .Z(n42890) );
  AND U43201 ( .A(n42891), .B(n42892), .Z(n42578) );
  NANDN U43202 ( .A(n42893), .B(n42894), .Z(n42892) );
  NANDN U43203 ( .A(n42895), .B(n42896), .Z(n42894) );
  NANDN U43204 ( .A(n42896), .B(n42895), .Z(n42891) );
  ANDN U43205 ( .B(B[130]), .A(n74), .Z(n42580) );
  XNOR U43206 ( .A(n42588), .B(n42897), .Z(n42581) );
  XNOR U43207 ( .A(n42587), .B(n42585), .Z(n42897) );
  AND U43208 ( .A(n42898), .B(n42899), .Z(n42585) );
  NANDN U43209 ( .A(n42900), .B(n42901), .Z(n42899) );
  OR U43210 ( .A(n42902), .B(n42903), .Z(n42901) );
  NAND U43211 ( .A(n42903), .B(n42902), .Z(n42898) );
  ANDN U43212 ( .B(B[131]), .A(n75), .Z(n42587) );
  XNOR U43213 ( .A(n42595), .B(n42904), .Z(n42588) );
  XNOR U43214 ( .A(n42594), .B(n42592), .Z(n42904) );
  AND U43215 ( .A(n42905), .B(n42906), .Z(n42592) );
  NANDN U43216 ( .A(n42907), .B(n42908), .Z(n42906) );
  NANDN U43217 ( .A(n42909), .B(n42910), .Z(n42908) );
  NANDN U43218 ( .A(n42910), .B(n42909), .Z(n42905) );
  ANDN U43219 ( .B(B[132]), .A(n76), .Z(n42594) );
  XNOR U43220 ( .A(n42602), .B(n42911), .Z(n42595) );
  XNOR U43221 ( .A(n42601), .B(n42599), .Z(n42911) );
  AND U43222 ( .A(n42912), .B(n42913), .Z(n42599) );
  NANDN U43223 ( .A(n42914), .B(n42915), .Z(n42913) );
  OR U43224 ( .A(n42916), .B(n42917), .Z(n42915) );
  NAND U43225 ( .A(n42917), .B(n42916), .Z(n42912) );
  ANDN U43226 ( .B(B[133]), .A(n77), .Z(n42601) );
  XNOR U43227 ( .A(n42609), .B(n42918), .Z(n42602) );
  XNOR U43228 ( .A(n42608), .B(n42606), .Z(n42918) );
  AND U43229 ( .A(n42919), .B(n42920), .Z(n42606) );
  NANDN U43230 ( .A(n42921), .B(n42922), .Z(n42920) );
  NANDN U43231 ( .A(n42923), .B(n42924), .Z(n42922) );
  NANDN U43232 ( .A(n42924), .B(n42923), .Z(n42919) );
  ANDN U43233 ( .B(B[134]), .A(n78), .Z(n42608) );
  XNOR U43234 ( .A(n42616), .B(n42925), .Z(n42609) );
  XNOR U43235 ( .A(n42615), .B(n42613), .Z(n42925) );
  AND U43236 ( .A(n42926), .B(n42927), .Z(n42613) );
  NANDN U43237 ( .A(n42928), .B(n42929), .Z(n42927) );
  OR U43238 ( .A(n42930), .B(n42931), .Z(n42929) );
  NAND U43239 ( .A(n42931), .B(n42930), .Z(n42926) );
  ANDN U43240 ( .B(B[135]), .A(n79), .Z(n42615) );
  XNOR U43241 ( .A(n42623), .B(n42932), .Z(n42616) );
  XNOR U43242 ( .A(n42622), .B(n42620), .Z(n42932) );
  AND U43243 ( .A(n42933), .B(n42934), .Z(n42620) );
  NANDN U43244 ( .A(n42935), .B(n42936), .Z(n42934) );
  NANDN U43245 ( .A(n42937), .B(n42938), .Z(n42936) );
  NANDN U43246 ( .A(n42938), .B(n42937), .Z(n42933) );
  ANDN U43247 ( .B(B[136]), .A(n80), .Z(n42622) );
  XNOR U43248 ( .A(n42630), .B(n42939), .Z(n42623) );
  XNOR U43249 ( .A(n42629), .B(n42627), .Z(n42939) );
  AND U43250 ( .A(n42940), .B(n42941), .Z(n42627) );
  NANDN U43251 ( .A(n42942), .B(n42943), .Z(n42941) );
  OR U43252 ( .A(n42944), .B(n42945), .Z(n42943) );
  NAND U43253 ( .A(n42945), .B(n42944), .Z(n42940) );
  ANDN U43254 ( .B(B[137]), .A(n81), .Z(n42629) );
  XNOR U43255 ( .A(n42637), .B(n42946), .Z(n42630) );
  XNOR U43256 ( .A(n42636), .B(n42634), .Z(n42946) );
  AND U43257 ( .A(n42947), .B(n42948), .Z(n42634) );
  NANDN U43258 ( .A(n42949), .B(n42950), .Z(n42948) );
  NAND U43259 ( .A(n42951), .B(n42952), .Z(n42950) );
  ANDN U43260 ( .B(B[138]), .A(n82), .Z(n42636) );
  XOR U43261 ( .A(n42643), .B(n42953), .Z(n42637) );
  XNOR U43262 ( .A(n42641), .B(n42644), .Z(n42953) );
  NAND U43263 ( .A(A[2]), .B(B[139]), .Z(n42644) );
  NANDN U43264 ( .A(n42954), .B(n42955), .Z(n42641) );
  AND U43265 ( .A(A[0]), .B(B[140]), .Z(n42955) );
  XNOR U43266 ( .A(n42646), .B(n42956), .Z(n42643) );
  NAND U43267 ( .A(A[0]), .B(B[141]), .Z(n42956) );
  NAND U43268 ( .A(B[140]), .B(A[1]), .Z(n42646) );
  NAND U43269 ( .A(n42957), .B(n42958), .Z(n514) );
  NANDN U43270 ( .A(n42959), .B(n42960), .Z(n42958) );
  OR U43271 ( .A(n42961), .B(n42962), .Z(n42960) );
  NAND U43272 ( .A(n42962), .B(n42961), .Z(n42957) );
  XOR U43273 ( .A(n516), .B(n515), .Z(\A1[138] ) );
  XOR U43274 ( .A(n42962), .B(n42963), .Z(n515) );
  XNOR U43275 ( .A(n42961), .B(n42959), .Z(n42963) );
  AND U43276 ( .A(n42964), .B(n42965), .Z(n42959) );
  NANDN U43277 ( .A(n42966), .B(n42967), .Z(n42965) );
  NANDN U43278 ( .A(n42968), .B(n42969), .Z(n42967) );
  NANDN U43279 ( .A(n42969), .B(n42968), .Z(n42964) );
  ANDN U43280 ( .B(B[109]), .A(n54), .Z(n42961) );
  XNOR U43281 ( .A(n42756), .B(n42970), .Z(n42962) );
  XNOR U43282 ( .A(n42755), .B(n42753), .Z(n42970) );
  AND U43283 ( .A(n42971), .B(n42972), .Z(n42753) );
  NANDN U43284 ( .A(n42973), .B(n42974), .Z(n42972) );
  OR U43285 ( .A(n42975), .B(n42976), .Z(n42974) );
  NAND U43286 ( .A(n42976), .B(n42975), .Z(n42971) );
  ANDN U43287 ( .B(B[110]), .A(n55), .Z(n42755) );
  XNOR U43288 ( .A(n42763), .B(n42977), .Z(n42756) );
  XNOR U43289 ( .A(n42762), .B(n42760), .Z(n42977) );
  AND U43290 ( .A(n42978), .B(n42979), .Z(n42760) );
  NANDN U43291 ( .A(n42980), .B(n42981), .Z(n42979) );
  NANDN U43292 ( .A(n42982), .B(n42983), .Z(n42981) );
  NANDN U43293 ( .A(n42983), .B(n42982), .Z(n42978) );
  ANDN U43294 ( .B(B[111]), .A(n56), .Z(n42762) );
  XNOR U43295 ( .A(n42770), .B(n42984), .Z(n42763) );
  XNOR U43296 ( .A(n42769), .B(n42767), .Z(n42984) );
  AND U43297 ( .A(n42985), .B(n42986), .Z(n42767) );
  NANDN U43298 ( .A(n42987), .B(n42988), .Z(n42986) );
  OR U43299 ( .A(n42989), .B(n42990), .Z(n42988) );
  NAND U43300 ( .A(n42990), .B(n42989), .Z(n42985) );
  ANDN U43301 ( .B(B[112]), .A(n57), .Z(n42769) );
  XNOR U43302 ( .A(n42777), .B(n42991), .Z(n42770) );
  XNOR U43303 ( .A(n42776), .B(n42774), .Z(n42991) );
  AND U43304 ( .A(n42992), .B(n42993), .Z(n42774) );
  NANDN U43305 ( .A(n42994), .B(n42995), .Z(n42993) );
  NANDN U43306 ( .A(n42996), .B(n42997), .Z(n42995) );
  NANDN U43307 ( .A(n42997), .B(n42996), .Z(n42992) );
  ANDN U43308 ( .B(B[113]), .A(n58), .Z(n42776) );
  XNOR U43309 ( .A(n42784), .B(n42998), .Z(n42777) );
  XNOR U43310 ( .A(n42783), .B(n42781), .Z(n42998) );
  AND U43311 ( .A(n42999), .B(n43000), .Z(n42781) );
  NANDN U43312 ( .A(n43001), .B(n43002), .Z(n43000) );
  OR U43313 ( .A(n43003), .B(n43004), .Z(n43002) );
  NAND U43314 ( .A(n43004), .B(n43003), .Z(n42999) );
  ANDN U43315 ( .B(B[114]), .A(n59), .Z(n42783) );
  XNOR U43316 ( .A(n42791), .B(n43005), .Z(n42784) );
  XNOR U43317 ( .A(n42790), .B(n42788), .Z(n43005) );
  AND U43318 ( .A(n43006), .B(n43007), .Z(n42788) );
  NANDN U43319 ( .A(n43008), .B(n43009), .Z(n43007) );
  NANDN U43320 ( .A(n43010), .B(n43011), .Z(n43009) );
  NANDN U43321 ( .A(n43011), .B(n43010), .Z(n43006) );
  ANDN U43322 ( .B(B[115]), .A(n60), .Z(n42790) );
  XNOR U43323 ( .A(n42798), .B(n43012), .Z(n42791) );
  XNOR U43324 ( .A(n42797), .B(n42795), .Z(n43012) );
  AND U43325 ( .A(n43013), .B(n43014), .Z(n42795) );
  NANDN U43326 ( .A(n43015), .B(n43016), .Z(n43014) );
  OR U43327 ( .A(n43017), .B(n43018), .Z(n43016) );
  NAND U43328 ( .A(n43018), .B(n43017), .Z(n43013) );
  ANDN U43329 ( .B(B[116]), .A(n61), .Z(n42797) );
  XNOR U43330 ( .A(n42805), .B(n43019), .Z(n42798) );
  XNOR U43331 ( .A(n42804), .B(n42802), .Z(n43019) );
  AND U43332 ( .A(n43020), .B(n43021), .Z(n42802) );
  NANDN U43333 ( .A(n43022), .B(n43023), .Z(n43021) );
  NANDN U43334 ( .A(n43024), .B(n43025), .Z(n43023) );
  NANDN U43335 ( .A(n43025), .B(n43024), .Z(n43020) );
  ANDN U43336 ( .B(B[117]), .A(n62), .Z(n42804) );
  XNOR U43337 ( .A(n42812), .B(n43026), .Z(n42805) );
  XNOR U43338 ( .A(n42811), .B(n42809), .Z(n43026) );
  AND U43339 ( .A(n43027), .B(n43028), .Z(n42809) );
  NANDN U43340 ( .A(n43029), .B(n43030), .Z(n43028) );
  OR U43341 ( .A(n43031), .B(n43032), .Z(n43030) );
  NAND U43342 ( .A(n43032), .B(n43031), .Z(n43027) );
  ANDN U43343 ( .B(B[118]), .A(n63), .Z(n42811) );
  XNOR U43344 ( .A(n42819), .B(n43033), .Z(n42812) );
  XNOR U43345 ( .A(n42818), .B(n42816), .Z(n43033) );
  AND U43346 ( .A(n43034), .B(n43035), .Z(n42816) );
  NANDN U43347 ( .A(n43036), .B(n43037), .Z(n43035) );
  NANDN U43348 ( .A(n43038), .B(n43039), .Z(n43037) );
  NANDN U43349 ( .A(n43039), .B(n43038), .Z(n43034) );
  ANDN U43350 ( .B(B[119]), .A(n64), .Z(n42818) );
  XNOR U43351 ( .A(n42826), .B(n43040), .Z(n42819) );
  XNOR U43352 ( .A(n42825), .B(n42823), .Z(n43040) );
  AND U43353 ( .A(n43041), .B(n43042), .Z(n42823) );
  NANDN U43354 ( .A(n43043), .B(n43044), .Z(n43042) );
  OR U43355 ( .A(n43045), .B(n43046), .Z(n43044) );
  NAND U43356 ( .A(n43046), .B(n43045), .Z(n43041) );
  ANDN U43357 ( .B(B[120]), .A(n65), .Z(n42825) );
  XNOR U43358 ( .A(n42833), .B(n43047), .Z(n42826) );
  XNOR U43359 ( .A(n42832), .B(n42830), .Z(n43047) );
  AND U43360 ( .A(n43048), .B(n43049), .Z(n42830) );
  NANDN U43361 ( .A(n43050), .B(n43051), .Z(n43049) );
  NANDN U43362 ( .A(n43052), .B(n43053), .Z(n43051) );
  NANDN U43363 ( .A(n43053), .B(n43052), .Z(n43048) );
  ANDN U43364 ( .B(B[121]), .A(n66), .Z(n42832) );
  XNOR U43365 ( .A(n42840), .B(n43054), .Z(n42833) );
  XNOR U43366 ( .A(n42839), .B(n42837), .Z(n43054) );
  AND U43367 ( .A(n43055), .B(n43056), .Z(n42837) );
  NANDN U43368 ( .A(n43057), .B(n43058), .Z(n43056) );
  OR U43369 ( .A(n43059), .B(n43060), .Z(n43058) );
  NAND U43370 ( .A(n43060), .B(n43059), .Z(n43055) );
  ANDN U43371 ( .B(B[122]), .A(n67), .Z(n42839) );
  XNOR U43372 ( .A(n42847), .B(n43061), .Z(n42840) );
  XNOR U43373 ( .A(n42846), .B(n42844), .Z(n43061) );
  AND U43374 ( .A(n43062), .B(n43063), .Z(n42844) );
  NANDN U43375 ( .A(n43064), .B(n43065), .Z(n43063) );
  NANDN U43376 ( .A(n43066), .B(n43067), .Z(n43065) );
  NANDN U43377 ( .A(n43067), .B(n43066), .Z(n43062) );
  ANDN U43378 ( .B(B[123]), .A(n68), .Z(n42846) );
  XNOR U43379 ( .A(n42854), .B(n43068), .Z(n42847) );
  XNOR U43380 ( .A(n42853), .B(n42851), .Z(n43068) );
  AND U43381 ( .A(n43069), .B(n43070), .Z(n42851) );
  NANDN U43382 ( .A(n43071), .B(n43072), .Z(n43070) );
  OR U43383 ( .A(n43073), .B(n43074), .Z(n43072) );
  NAND U43384 ( .A(n43074), .B(n43073), .Z(n43069) );
  ANDN U43385 ( .B(B[124]), .A(n69), .Z(n42853) );
  XNOR U43386 ( .A(n42861), .B(n43075), .Z(n42854) );
  XNOR U43387 ( .A(n42860), .B(n42858), .Z(n43075) );
  AND U43388 ( .A(n43076), .B(n43077), .Z(n42858) );
  NANDN U43389 ( .A(n43078), .B(n43079), .Z(n43077) );
  NANDN U43390 ( .A(n43080), .B(n43081), .Z(n43079) );
  NANDN U43391 ( .A(n43081), .B(n43080), .Z(n43076) );
  ANDN U43392 ( .B(B[125]), .A(n70), .Z(n42860) );
  XNOR U43393 ( .A(n42868), .B(n43082), .Z(n42861) );
  XNOR U43394 ( .A(n42867), .B(n42865), .Z(n43082) );
  AND U43395 ( .A(n43083), .B(n43084), .Z(n42865) );
  NANDN U43396 ( .A(n43085), .B(n43086), .Z(n43084) );
  OR U43397 ( .A(n43087), .B(n43088), .Z(n43086) );
  NAND U43398 ( .A(n43088), .B(n43087), .Z(n43083) );
  ANDN U43399 ( .B(B[126]), .A(n71), .Z(n42867) );
  XNOR U43400 ( .A(n42875), .B(n43089), .Z(n42868) );
  XNOR U43401 ( .A(n42874), .B(n42872), .Z(n43089) );
  AND U43402 ( .A(n43090), .B(n43091), .Z(n42872) );
  NANDN U43403 ( .A(n43092), .B(n43093), .Z(n43091) );
  NANDN U43404 ( .A(n43094), .B(n43095), .Z(n43093) );
  NANDN U43405 ( .A(n43095), .B(n43094), .Z(n43090) );
  ANDN U43406 ( .B(B[127]), .A(n72), .Z(n42874) );
  XNOR U43407 ( .A(n42882), .B(n43096), .Z(n42875) );
  XNOR U43408 ( .A(n42881), .B(n42879), .Z(n43096) );
  AND U43409 ( .A(n43097), .B(n43098), .Z(n42879) );
  NANDN U43410 ( .A(n43099), .B(n43100), .Z(n43098) );
  OR U43411 ( .A(n43101), .B(n43102), .Z(n43100) );
  NAND U43412 ( .A(n43102), .B(n43101), .Z(n43097) );
  ANDN U43413 ( .B(B[128]), .A(n73), .Z(n42881) );
  XNOR U43414 ( .A(n42889), .B(n43103), .Z(n42882) );
  XNOR U43415 ( .A(n42888), .B(n42886), .Z(n43103) );
  AND U43416 ( .A(n43104), .B(n43105), .Z(n42886) );
  NANDN U43417 ( .A(n43106), .B(n43107), .Z(n43105) );
  NANDN U43418 ( .A(n43108), .B(n43109), .Z(n43107) );
  NANDN U43419 ( .A(n43109), .B(n43108), .Z(n43104) );
  ANDN U43420 ( .B(B[129]), .A(n74), .Z(n42888) );
  XNOR U43421 ( .A(n42896), .B(n43110), .Z(n42889) );
  XNOR U43422 ( .A(n42895), .B(n42893), .Z(n43110) );
  AND U43423 ( .A(n43111), .B(n43112), .Z(n42893) );
  NANDN U43424 ( .A(n43113), .B(n43114), .Z(n43112) );
  OR U43425 ( .A(n43115), .B(n43116), .Z(n43114) );
  NAND U43426 ( .A(n43116), .B(n43115), .Z(n43111) );
  ANDN U43427 ( .B(B[130]), .A(n75), .Z(n42895) );
  XNOR U43428 ( .A(n42903), .B(n43117), .Z(n42896) );
  XNOR U43429 ( .A(n42902), .B(n42900), .Z(n43117) );
  AND U43430 ( .A(n43118), .B(n43119), .Z(n42900) );
  NANDN U43431 ( .A(n43120), .B(n43121), .Z(n43119) );
  NANDN U43432 ( .A(n43122), .B(n43123), .Z(n43121) );
  NANDN U43433 ( .A(n43123), .B(n43122), .Z(n43118) );
  ANDN U43434 ( .B(B[131]), .A(n76), .Z(n42902) );
  XNOR U43435 ( .A(n42910), .B(n43124), .Z(n42903) );
  XNOR U43436 ( .A(n42909), .B(n42907), .Z(n43124) );
  AND U43437 ( .A(n43125), .B(n43126), .Z(n42907) );
  NANDN U43438 ( .A(n43127), .B(n43128), .Z(n43126) );
  OR U43439 ( .A(n43129), .B(n43130), .Z(n43128) );
  NAND U43440 ( .A(n43130), .B(n43129), .Z(n43125) );
  ANDN U43441 ( .B(B[132]), .A(n77), .Z(n42909) );
  XNOR U43442 ( .A(n42917), .B(n43131), .Z(n42910) );
  XNOR U43443 ( .A(n42916), .B(n42914), .Z(n43131) );
  AND U43444 ( .A(n43132), .B(n43133), .Z(n42914) );
  NANDN U43445 ( .A(n43134), .B(n43135), .Z(n43133) );
  NANDN U43446 ( .A(n43136), .B(n43137), .Z(n43135) );
  NANDN U43447 ( .A(n43137), .B(n43136), .Z(n43132) );
  ANDN U43448 ( .B(B[133]), .A(n78), .Z(n42916) );
  XNOR U43449 ( .A(n42924), .B(n43138), .Z(n42917) );
  XNOR U43450 ( .A(n42923), .B(n42921), .Z(n43138) );
  AND U43451 ( .A(n43139), .B(n43140), .Z(n42921) );
  NANDN U43452 ( .A(n43141), .B(n43142), .Z(n43140) );
  OR U43453 ( .A(n43143), .B(n43144), .Z(n43142) );
  NAND U43454 ( .A(n43144), .B(n43143), .Z(n43139) );
  ANDN U43455 ( .B(B[134]), .A(n79), .Z(n42923) );
  XNOR U43456 ( .A(n42931), .B(n43145), .Z(n42924) );
  XNOR U43457 ( .A(n42930), .B(n42928), .Z(n43145) );
  AND U43458 ( .A(n43146), .B(n43147), .Z(n42928) );
  NANDN U43459 ( .A(n43148), .B(n43149), .Z(n43147) );
  NANDN U43460 ( .A(n43150), .B(n43151), .Z(n43149) );
  NANDN U43461 ( .A(n43151), .B(n43150), .Z(n43146) );
  ANDN U43462 ( .B(B[135]), .A(n80), .Z(n42930) );
  XNOR U43463 ( .A(n42938), .B(n43152), .Z(n42931) );
  XNOR U43464 ( .A(n42937), .B(n42935), .Z(n43152) );
  AND U43465 ( .A(n43153), .B(n43154), .Z(n42935) );
  NANDN U43466 ( .A(n43155), .B(n43156), .Z(n43154) );
  OR U43467 ( .A(n43157), .B(n43158), .Z(n43156) );
  NAND U43468 ( .A(n43158), .B(n43157), .Z(n43153) );
  ANDN U43469 ( .B(B[136]), .A(n81), .Z(n42937) );
  XNOR U43470 ( .A(n42945), .B(n43159), .Z(n42938) );
  XNOR U43471 ( .A(n42944), .B(n42942), .Z(n43159) );
  AND U43472 ( .A(n43160), .B(n43161), .Z(n42942) );
  NANDN U43473 ( .A(n43162), .B(n43163), .Z(n43161) );
  NAND U43474 ( .A(n43164), .B(n43165), .Z(n43163) );
  ANDN U43475 ( .B(B[137]), .A(n82), .Z(n42944) );
  XOR U43476 ( .A(n42951), .B(n43166), .Z(n42945) );
  XNOR U43477 ( .A(n42949), .B(n42952), .Z(n43166) );
  NAND U43478 ( .A(A[2]), .B(B[138]), .Z(n42952) );
  NANDN U43479 ( .A(n43167), .B(n43168), .Z(n42949) );
  AND U43480 ( .A(A[0]), .B(B[139]), .Z(n43168) );
  XNOR U43481 ( .A(n42954), .B(n43169), .Z(n42951) );
  NAND U43482 ( .A(A[0]), .B(B[140]), .Z(n43169) );
  NAND U43483 ( .A(B[139]), .B(A[1]), .Z(n42954) );
  NAND U43484 ( .A(n43170), .B(n43171), .Z(n516) );
  NANDN U43485 ( .A(n43172), .B(n43173), .Z(n43171) );
  OR U43486 ( .A(n43174), .B(n43175), .Z(n43173) );
  NAND U43487 ( .A(n43175), .B(n43174), .Z(n43170) );
  XOR U43488 ( .A(n518), .B(n517), .Z(\A1[137] ) );
  XOR U43489 ( .A(n43175), .B(n43176), .Z(n517) );
  XNOR U43490 ( .A(n43174), .B(n43172), .Z(n43176) );
  AND U43491 ( .A(n43177), .B(n43178), .Z(n43172) );
  NANDN U43492 ( .A(n43179), .B(n43180), .Z(n43178) );
  NANDN U43493 ( .A(n43181), .B(n43182), .Z(n43180) );
  NANDN U43494 ( .A(n43182), .B(n43181), .Z(n43177) );
  ANDN U43495 ( .B(B[108]), .A(n54), .Z(n43174) );
  XNOR U43496 ( .A(n42969), .B(n43183), .Z(n43175) );
  XNOR U43497 ( .A(n42968), .B(n42966), .Z(n43183) );
  AND U43498 ( .A(n43184), .B(n43185), .Z(n42966) );
  NANDN U43499 ( .A(n43186), .B(n43187), .Z(n43185) );
  OR U43500 ( .A(n43188), .B(n43189), .Z(n43187) );
  NAND U43501 ( .A(n43189), .B(n43188), .Z(n43184) );
  ANDN U43502 ( .B(B[109]), .A(n55), .Z(n42968) );
  XNOR U43503 ( .A(n42976), .B(n43190), .Z(n42969) );
  XNOR U43504 ( .A(n42975), .B(n42973), .Z(n43190) );
  AND U43505 ( .A(n43191), .B(n43192), .Z(n42973) );
  NANDN U43506 ( .A(n43193), .B(n43194), .Z(n43192) );
  NANDN U43507 ( .A(n43195), .B(n43196), .Z(n43194) );
  NANDN U43508 ( .A(n43196), .B(n43195), .Z(n43191) );
  ANDN U43509 ( .B(B[110]), .A(n56), .Z(n42975) );
  XNOR U43510 ( .A(n42983), .B(n43197), .Z(n42976) );
  XNOR U43511 ( .A(n42982), .B(n42980), .Z(n43197) );
  AND U43512 ( .A(n43198), .B(n43199), .Z(n42980) );
  NANDN U43513 ( .A(n43200), .B(n43201), .Z(n43199) );
  OR U43514 ( .A(n43202), .B(n43203), .Z(n43201) );
  NAND U43515 ( .A(n43203), .B(n43202), .Z(n43198) );
  ANDN U43516 ( .B(B[111]), .A(n57), .Z(n42982) );
  XNOR U43517 ( .A(n42990), .B(n43204), .Z(n42983) );
  XNOR U43518 ( .A(n42989), .B(n42987), .Z(n43204) );
  AND U43519 ( .A(n43205), .B(n43206), .Z(n42987) );
  NANDN U43520 ( .A(n43207), .B(n43208), .Z(n43206) );
  NANDN U43521 ( .A(n43209), .B(n43210), .Z(n43208) );
  NANDN U43522 ( .A(n43210), .B(n43209), .Z(n43205) );
  ANDN U43523 ( .B(B[112]), .A(n58), .Z(n42989) );
  XNOR U43524 ( .A(n42997), .B(n43211), .Z(n42990) );
  XNOR U43525 ( .A(n42996), .B(n42994), .Z(n43211) );
  AND U43526 ( .A(n43212), .B(n43213), .Z(n42994) );
  NANDN U43527 ( .A(n43214), .B(n43215), .Z(n43213) );
  OR U43528 ( .A(n43216), .B(n43217), .Z(n43215) );
  NAND U43529 ( .A(n43217), .B(n43216), .Z(n43212) );
  ANDN U43530 ( .B(B[113]), .A(n59), .Z(n42996) );
  XNOR U43531 ( .A(n43004), .B(n43218), .Z(n42997) );
  XNOR U43532 ( .A(n43003), .B(n43001), .Z(n43218) );
  AND U43533 ( .A(n43219), .B(n43220), .Z(n43001) );
  NANDN U43534 ( .A(n43221), .B(n43222), .Z(n43220) );
  NANDN U43535 ( .A(n43223), .B(n43224), .Z(n43222) );
  NANDN U43536 ( .A(n43224), .B(n43223), .Z(n43219) );
  ANDN U43537 ( .B(B[114]), .A(n60), .Z(n43003) );
  XNOR U43538 ( .A(n43011), .B(n43225), .Z(n43004) );
  XNOR U43539 ( .A(n43010), .B(n43008), .Z(n43225) );
  AND U43540 ( .A(n43226), .B(n43227), .Z(n43008) );
  NANDN U43541 ( .A(n43228), .B(n43229), .Z(n43227) );
  OR U43542 ( .A(n43230), .B(n43231), .Z(n43229) );
  NAND U43543 ( .A(n43231), .B(n43230), .Z(n43226) );
  ANDN U43544 ( .B(B[115]), .A(n61), .Z(n43010) );
  XNOR U43545 ( .A(n43018), .B(n43232), .Z(n43011) );
  XNOR U43546 ( .A(n43017), .B(n43015), .Z(n43232) );
  AND U43547 ( .A(n43233), .B(n43234), .Z(n43015) );
  NANDN U43548 ( .A(n43235), .B(n43236), .Z(n43234) );
  NANDN U43549 ( .A(n43237), .B(n43238), .Z(n43236) );
  NANDN U43550 ( .A(n43238), .B(n43237), .Z(n43233) );
  ANDN U43551 ( .B(B[116]), .A(n62), .Z(n43017) );
  XNOR U43552 ( .A(n43025), .B(n43239), .Z(n43018) );
  XNOR U43553 ( .A(n43024), .B(n43022), .Z(n43239) );
  AND U43554 ( .A(n43240), .B(n43241), .Z(n43022) );
  NANDN U43555 ( .A(n43242), .B(n43243), .Z(n43241) );
  OR U43556 ( .A(n43244), .B(n43245), .Z(n43243) );
  NAND U43557 ( .A(n43245), .B(n43244), .Z(n43240) );
  ANDN U43558 ( .B(B[117]), .A(n63), .Z(n43024) );
  XNOR U43559 ( .A(n43032), .B(n43246), .Z(n43025) );
  XNOR U43560 ( .A(n43031), .B(n43029), .Z(n43246) );
  AND U43561 ( .A(n43247), .B(n43248), .Z(n43029) );
  NANDN U43562 ( .A(n43249), .B(n43250), .Z(n43248) );
  NANDN U43563 ( .A(n43251), .B(n43252), .Z(n43250) );
  NANDN U43564 ( .A(n43252), .B(n43251), .Z(n43247) );
  ANDN U43565 ( .B(B[118]), .A(n64), .Z(n43031) );
  XNOR U43566 ( .A(n43039), .B(n43253), .Z(n43032) );
  XNOR U43567 ( .A(n43038), .B(n43036), .Z(n43253) );
  AND U43568 ( .A(n43254), .B(n43255), .Z(n43036) );
  NANDN U43569 ( .A(n43256), .B(n43257), .Z(n43255) );
  OR U43570 ( .A(n43258), .B(n43259), .Z(n43257) );
  NAND U43571 ( .A(n43259), .B(n43258), .Z(n43254) );
  ANDN U43572 ( .B(B[119]), .A(n65), .Z(n43038) );
  XNOR U43573 ( .A(n43046), .B(n43260), .Z(n43039) );
  XNOR U43574 ( .A(n43045), .B(n43043), .Z(n43260) );
  AND U43575 ( .A(n43261), .B(n43262), .Z(n43043) );
  NANDN U43576 ( .A(n43263), .B(n43264), .Z(n43262) );
  NANDN U43577 ( .A(n43265), .B(n43266), .Z(n43264) );
  NANDN U43578 ( .A(n43266), .B(n43265), .Z(n43261) );
  ANDN U43579 ( .B(B[120]), .A(n66), .Z(n43045) );
  XNOR U43580 ( .A(n43053), .B(n43267), .Z(n43046) );
  XNOR U43581 ( .A(n43052), .B(n43050), .Z(n43267) );
  AND U43582 ( .A(n43268), .B(n43269), .Z(n43050) );
  NANDN U43583 ( .A(n43270), .B(n43271), .Z(n43269) );
  OR U43584 ( .A(n43272), .B(n43273), .Z(n43271) );
  NAND U43585 ( .A(n43273), .B(n43272), .Z(n43268) );
  ANDN U43586 ( .B(B[121]), .A(n67), .Z(n43052) );
  XNOR U43587 ( .A(n43060), .B(n43274), .Z(n43053) );
  XNOR U43588 ( .A(n43059), .B(n43057), .Z(n43274) );
  AND U43589 ( .A(n43275), .B(n43276), .Z(n43057) );
  NANDN U43590 ( .A(n43277), .B(n43278), .Z(n43276) );
  NANDN U43591 ( .A(n43279), .B(n43280), .Z(n43278) );
  NANDN U43592 ( .A(n43280), .B(n43279), .Z(n43275) );
  ANDN U43593 ( .B(B[122]), .A(n68), .Z(n43059) );
  XNOR U43594 ( .A(n43067), .B(n43281), .Z(n43060) );
  XNOR U43595 ( .A(n43066), .B(n43064), .Z(n43281) );
  AND U43596 ( .A(n43282), .B(n43283), .Z(n43064) );
  NANDN U43597 ( .A(n43284), .B(n43285), .Z(n43283) );
  OR U43598 ( .A(n43286), .B(n43287), .Z(n43285) );
  NAND U43599 ( .A(n43287), .B(n43286), .Z(n43282) );
  ANDN U43600 ( .B(B[123]), .A(n69), .Z(n43066) );
  XNOR U43601 ( .A(n43074), .B(n43288), .Z(n43067) );
  XNOR U43602 ( .A(n43073), .B(n43071), .Z(n43288) );
  AND U43603 ( .A(n43289), .B(n43290), .Z(n43071) );
  NANDN U43604 ( .A(n43291), .B(n43292), .Z(n43290) );
  NANDN U43605 ( .A(n43293), .B(n43294), .Z(n43292) );
  NANDN U43606 ( .A(n43294), .B(n43293), .Z(n43289) );
  ANDN U43607 ( .B(B[124]), .A(n70), .Z(n43073) );
  XNOR U43608 ( .A(n43081), .B(n43295), .Z(n43074) );
  XNOR U43609 ( .A(n43080), .B(n43078), .Z(n43295) );
  AND U43610 ( .A(n43296), .B(n43297), .Z(n43078) );
  NANDN U43611 ( .A(n43298), .B(n43299), .Z(n43297) );
  OR U43612 ( .A(n43300), .B(n43301), .Z(n43299) );
  NAND U43613 ( .A(n43301), .B(n43300), .Z(n43296) );
  ANDN U43614 ( .B(B[125]), .A(n71), .Z(n43080) );
  XNOR U43615 ( .A(n43088), .B(n43302), .Z(n43081) );
  XNOR U43616 ( .A(n43087), .B(n43085), .Z(n43302) );
  AND U43617 ( .A(n43303), .B(n43304), .Z(n43085) );
  NANDN U43618 ( .A(n43305), .B(n43306), .Z(n43304) );
  NANDN U43619 ( .A(n43307), .B(n43308), .Z(n43306) );
  NANDN U43620 ( .A(n43308), .B(n43307), .Z(n43303) );
  ANDN U43621 ( .B(B[126]), .A(n72), .Z(n43087) );
  XNOR U43622 ( .A(n43095), .B(n43309), .Z(n43088) );
  XNOR U43623 ( .A(n43094), .B(n43092), .Z(n43309) );
  AND U43624 ( .A(n43310), .B(n43311), .Z(n43092) );
  NANDN U43625 ( .A(n43312), .B(n43313), .Z(n43311) );
  OR U43626 ( .A(n43314), .B(n43315), .Z(n43313) );
  NAND U43627 ( .A(n43315), .B(n43314), .Z(n43310) );
  ANDN U43628 ( .B(B[127]), .A(n73), .Z(n43094) );
  XNOR U43629 ( .A(n43102), .B(n43316), .Z(n43095) );
  XNOR U43630 ( .A(n43101), .B(n43099), .Z(n43316) );
  AND U43631 ( .A(n43317), .B(n43318), .Z(n43099) );
  NANDN U43632 ( .A(n43319), .B(n43320), .Z(n43318) );
  NANDN U43633 ( .A(n43321), .B(n43322), .Z(n43320) );
  NANDN U43634 ( .A(n43322), .B(n43321), .Z(n43317) );
  ANDN U43635 ( .B(B[128]), .A(n74), .Z(n43101) );
  XNOR U43636 ( .A(n43109), .B(n43323), .Z(n43102) );
  XNOR U43637 ( .A(n43108), .B(n43106), .Z(n43323) );
  AND U43638 ( .A(n43324), .B(n43325), .Z(n43106) );
  NANDN U43639 ( .A(n43326), .B(n43327), .Z(n43325) );
  OR U43640 ( .A(n43328), .B(n43329), .Z(n43327) );
  NAND U43641 ( .A(n43329), .B(n43328), .Z(n43324) );
  ANDN U43642 ( .B(B[129]), .A(n75), .Z(n43108) );
  XNOR U43643 ( .A(n43116), .B(n43330), .Z(n43109) );
  XNOR U43644 ( .A(n43115), .B(n43113), .Z(n43330) );
  AND U43645 ( .A(n43331), .B(n43332), .Z(n43113) );
  NANDN U43646 ( .A(n43333), .B(n43334), .Z(n43332) );
  NANDN U43647 ( .A(n43335), .B(n43336), .Z(n43334) );
  NANDN U43648 ( .A(n43336), .B(n43335), .Z(n43331) );
  ANDN U43649 ( .B(B[130]), .A(n76), .Z(n43115) );
  XNOR U43650 ( .A(n43123), .B(n43337), .Z(n43116) );
  XNOR U43651 ( .A(n43122), .B(n43120), .Z(n43337) );
  AND U43652 ( .A(n43338), .B(n43339), .Z(n43120) );
  NANDN U43653 ( .A(n43340), .B(n43341), .Z(n43339) );
  OR U43654 ( .A(n43342), .B(n43343), .Z(n43341) );
  NAND U43655 ( .A(n43343), .B(n43342), .Z(n43338) );
  ANDN U43656 ( .B(B[131]), .A(n77), .Z(n43122) );
  XNOR U43657 ( .A(n43130), .B(n43344), .Z(n43123) );
  XNOR U43658 ( .A(n43129), .B(n43127), .Z(n43344) );
  AND U43659 ( .A(n43345), .B(n43346), .Z(n43127) );
  NANDN U43660 ( .A(n43347), .B(n43348), .Z(n43346) );
  NANDN U43661 ( .A(n43349), .B(n43350), .Z(n43348) );
  NANDN U43662 ( .A(n43350), .B(n43349), .Z(n43345) );
  ANDN U43663 ( .B(B[132]), .A(n78), .Z(n43129) );
  XNOR U43664 ( .A(n43137), .B(n43351), .Z(n43130) );
  XNOR U43665 ( .A(n43136), .B(n43134), .Z(n43351) );
  AND U43666 ( .A(n43352), .B(n43353), .Z(n43134) );
  NANDN U43667 ( .A(n43354), .B(n43355), .Z(n43353) );
  OR U43668 ( .A(n43356), .B(n43357), .Z(n43355) );
  NAND U43669 ( .A(n43357), .B(n43356), .Z(n43352) );
  ANDN U43670 ( .B(B[133]), .A(n79), .Z(n43136) );
  XNOR U43671 ( .A(n43144), .B(n43358), .Z(n43137) );
  XNOR U43672 ( .A(n43143), .B(n43141), .Z(n43358) );
  AND U43673 ( .A(n43359), .B(n43360), .Z(n43141) );
  NANDN U43674 ( .A(n43361), .B(n43362), .Z(n43360) );
  NANDN U43675 ( .A(n43363), .B(n43364), .Z(n43362) );
  NANDN U43676 ( .A(n43364), .B(n43363), .Z(n43359) );
  ANDN U43677 ( .B(B[134]), .A(n80), .Z(n43143) );
  XNOR U43678 ( .A(n43151), .B(n43365), .Z(n43144) );
  XNOR U43679 ( .A(n43150), .B(n43148), .Z(n43365) );
  AND U43680 ( .A(n43366), .B(n43367), .Z(n43148) );
  NANDN U43681 ( .A(n43368), .B(n43369), .Z(n43367) );
  OR U43682 ( .A(n43370), .B(n43371), .Z(n43369) );
  NAND U43683 ( .A(n43371), .B(n43370), .Z(n43366) );
  ANDN U43684 ( .B(B[135]), .A(n81), .Z(n43150) );
  XNOR U43685 ( .A(n43158), .B(n43372), .Z(n43151) );
  XNOR U43686 ( .A(n43157), .B(n43155), .Z(n43372) );
  AND U43687 ( .A(n43373), .B(n43374), .Z(n43155) );
  NANDN U43688 ( .A(n43375), .B(n43376), .Z(n43374) );
  NAND U43689 ( .A(n43377), .B(n43378), .Z(n43376) );
  ANDN U43690 ( .B(B[136]), .A(n82), .Z(n43157) );
  XOR U43691 ( .A(n43164), .B(n43379), .Z(n43158) );
  XNOR U43692 ( .A(n43162), .B(n43165), .Z(n43379) );
  NAND U43693 ( .A(A[2]), .B(B[137]), .Z(n43165) );
  NANDN U43694 ( .A(n43380), .B(n43381), .Z(n43162) );
  AND U43695 ( .A(A[0]), .B(B[138]), .Z(n43381) );
  XNOR U43696 ( .A(n43167), .B(n43382), .Z(n43164) );
  NAND U43697 ( .A(A[0]), .B(B[139]), .Z(n43382) );
  NAND U43698 ( .A(B[138]), .B(A[1]), .Z(n43167) );
  NAND U43699 ( .A(n43383), .B(n43384), .Z(n518) );
  NANDN U43700 ( .A(n43385), .B(n43386), .Z(n43384) );
  OR U43701 ( .A(n43387), .B(n43388), .Z(n43386) );
  NAND U43702 ( .A(n43388), .B(n43387), .Z(n43383) );
  XOR U43703 ( .A(n520), .B(n519), .Z(\A1[136] ) );
  XOR U43704 ( .A(n43388), .B(n43389), .Z(n519) );
  XNOR U43705 ( .A(n43387), .B(n43385), .Z(n43389) );
  AND U43706 ( .A(n43390), .B(n43391), .Z(n43385) );
  NANDN U43707 ( .A(n43392), .B(n43393), .Z(n43391) );
  NANDN U43708 ( .A(n43394), .B(n43395), .Z(n43393) );
  NANDN U43709 ( .A(n43395), .B(n43394), .Z(n43390) );
  ANDN U43710 ( .B(B[107]), .A(n54), .Z(n43387) );
  XNOR U43711 ( .A(n43182), .B(n43396), .Z(n43388) );
  XNOR U43712 ( .A(n43181), .B(n43179), .Z(n43396) );
  AND U43713 ( .A(n43397), .B(n43398), .Z(n43179) );
  NANDN U43714 ( .A(n43399), .B(n43400), .Z(n43398) );
  OR U43715 ( .A(n43401), .B(n43402), .Z(n43400) );
  NAND U43716 ( .A(n43402), .B(n43401), .Z(n43397) );
  ANDN U43717 ( .B(B[108]), .A(n55), .Z(n43181) );
  XNOR U43718 ( .A(n43189), .B(n43403), .Z(n43182) );
  XNOR U43719 ( .A(n43188), .B(n43186), .Z(n43403) );
  AND U43720 ( .A(n43404), .B(n43405), .Z(n43186) );
  NANDN U43721 ( .A(n43406), .B(n43407), .Z(n43405) );
  NANDN U43722 ( .A(n43408), .B(n43409), .Z(n43407) );
  NANDN U43723 ( .A(n43409), .B(n43408), .Z(n43404) );
  ANDN U43724 ( .B(B[109]), .A(n56), .Z(n43188) );
  XNOR U43725 ( .A(n43196), .B(n43410), .Z(n43189) );
  XNOR U43726 ( .A(n43195), .B(n43193), .Z(n43410) );
  AND U43727 ( .A(n43411), .B(n43412), .Z(n43193) );
  NANDN U43728 ( .A(n43413), .B(n43414), .Z(n43412) );
  OR U43729 ( .A(n43415), .B(n43416), .Z(n43414) );
  NAND U43730 ( .A(n43416), .B(n43415), .Z(n43411) );
  ANDN U43731 ( .B(B[110]), .A(n57), .Z(n43195) );
  XNOR U43732 ( .A(n43203), .B(n43417), .Z(n43196) );
  XNOR U43733 ( .A(n43202), .B(n43200), .Z(n43417) );
  AND U43734 ( .A(n43418), .B(n43419), .Z(n43200) );
  NANDN U43735 ( .A(n43420), .B(n43421), .Z(n43419) );
  NANDN U43736 ( .A(n43422), .B(n43423), .Z(n43421) );
  NANDN U43737 ( .A(n43423), .B(n43422), .Z(n43418) );
  ANDN U43738 ( .B(B[111]), .A(n58), .Z(n43202) );
  XNOR U43739 ( .A(n43210), .B(n43424), .Z(n43203) );
  XNOR U43740 ( .A(n43209), .B(n43207), .Z(n43424) );
  AND U43741 ( .A(n43425), .B(n43426), .Z(n43207) );
  NANDN U43742 ( .A(n43427), .B(n43428), .Z(n43426) );
  OR U43743 ( .A(n43429), .B(n43430), .Z(n43428) );
  NAND U43744 ( .A(n43430), .B(n43429), .Z(n43425) );
  ANDN U43745 ( .B(B[112]), .A(n59), .Z(n43209) );
  XNOR U43746 ( .A(n43217), .B(n43431), .Z(n43210) );
  XNOR U43747 ( .A(n43216), .B(n43214), .Z(n43431) );
  AND U43748 ( .A(n43432), .B(n43433), .Z(n43214) );
  NANDN U43749 ( .A(n43434), .B(n43435), .Z(n43433) );
  NANDN U43750 ( .A(n43436), .B(n43437), .Z(n43435) );
  NANDN U43751 ( .A(n43437), .B(n43436), .Z(n43432) );
  ANDN U43752 ( .B(B[113]), .A(n60), .Z(n43216) );
  XNOR U43753 ( .A(n43224), .B(n43438), .Z(n43217) );
  XNOR U43754 ( .A(n43223), .B(n43221), .Z(n43438) );
  AND U43755 ( .A(n43439), .B(n43440), .Z(n43221) );
  NANDN U43756 ( .A(n43441), .B(n43442), .Z(n43440) );
  OR U43757 ( .A(n43443), .B(n43444), .Z(n43442) );
  NAND U43758 ( .A(n43444), .B(n43443), .Z(n43439) );
  ANDN U43759 ( .B(B[114]), .A(n61), .Z(n43223) );
  XNOR U43760 ( .A(n43231), .B(n43445), .Z(n43224) );
  XNOR U43761 ( .A(n43230), .B(n43228), .Z(n43445) );
  AND U43762 ( .A(n43446), .B(n43447), .Z(n43228) );
  NANDN U43763 ( .A(n43448), .B(n43449), .Z(n43447) );
  NANDN U43764 ( .A(n43450), .B(n43451), .Z(n43449) );
  NANDN U43765 ( .A(n43451), .B(n43450), .Z(n43446) );
  ANDN U43766 ( .B(B[115]), .A(n62), .Z(n43230) );
  XNOR U43767 ( .A(n43238), .B(n43452), .Z(n43231) );
  XNOR U43768 ( .A(n43237), .B(n43235), .Z(n43452) );
  AND U43769 ( .A(n43453), .B(n43454), .Z(n43235) );
  NANDN U43770 ( .A(n43455), .B(n43456), .Z(n43454) );
  OR U43771 ( .A(n43457), .B(n43458), .Z(n43456) );
  NAND U43772 ( .A(n43458), .B(n43457), .Z(n43453) );
  ANDN U43773 ( .B(B[116]), .A(n63), .Z(n43237) );
  XNOR U43774 ( .A(n43245), .B(n43459), .Z(n43238) );
  XNOR U43775 ( .A(n43244), .B(n43242), .Z(n43459) );
  AND U43776 ( .A(n43460), .B(n43461), .Z(n43242) );
  NANDN U43777 ( .A(n43462), .B(n43463), .Z(n43461) );
  NANDN U43778 ( .A(n43464), .B(n43465), .Z(n43463) );
  NANDN U43779 ( .A(n43465), .B(n43464), .Z(n43460) );
  ANDN U43780 ( .B(B[117]), .A(n64), .Z(n43244) );
  XNOR U43781 ( .A(n43252), .B(n43466), .Z(n43245) );
  XNOR U43782 ( .A(n43251), .B(n43249), .Z(n43466) );
  AND U43783 ( .A(n43467), .B(n43468), .Z(n43249) );
  NANDN U43784 ( .A(n43469), .B(n43470), .Z(n43468) );
  OR U43785 ( .A(n43471), .B(n43472), .Z(n43470) );
  NAND U43786 ( .A(n43472), .B(n43471), .Z(n43467) );
  ANDN U43787 ( .B(B[118]), .A(n65), .Z(n43251) );
  XNOR U43788 ( .A(n43259), .B(n43473), .Z(n43252) );
  XNOR U43789 ( .A(n43258), .B(n43256), .Z(n43473) );
  AND U43790 ( .A(n43474), .B(n43475), .Z(n43256) );
  NANDN U43791 ( .A(n43476), .B(n43477), .Z(n43475) );
  NANDN U43792 ( .A(n43478), .B(n43479), .Z(n43477) );
  NANDN U43793 ( .A(n43479), .B(n43478), .Z(n43474) );
  ANDN U43794 ( .B(B[119]), .A(n66), .Z(n43258) );
  XNOR U43795 ( .A(n43266), .B(n43480), .Z(n43259) );
  XNOR U43796 ( .A(n43265), .B(n43263), .Z(n43480) );
  AND U43797 ( .A(n43481), .B(n43482), .Z(n43263) );
  NANDN U43798 ( .A(n43483), .B(n43484), .Z(n43482) );
  OR U43799 ( .A(n43485), .B(n43486), .Z(n43484) );
  NAND U43800 ( .A(n43486), .B(n43485), .Z(n43481) );
  ANDN U43801 ( .B(B[120]), .A(n67), .Z(n43265) );
  XNOR U43802 ( .A(n43273), .B(n43487), .Z(n43266) );
  XNOR U43803 ( .A(n43272), .B(n43270), .Z(n43487) );
  AND U43804 ( .A(n43488), .B(n43489), .Z(n43270) );
  NANDN U43805 ( .A(n43490), .B(n43491), .Z(n43489) );
  NANDN U43806 ( .A(n43492), .B(n43493), .Z(n43491) );
  NANDN U43807 ( .A(n43493), .B(n43492), .Z(n43488) );
  ANDN U43808 ( .B(B[121]), .A(n68), .Z(n43272) );
  XNOR U43809 ( .A(n43280), .B(n43494), .Z(n43273) );
  XNOR U43810 ( .A(n43279), .B(n43277), .Z(n43494) );
  AND U43811 ( .A(n43495), .B(n43496), .Z(n43277) );
  NANDN U43812 ( .A(n43497), .B(n43498), .Z(n43496) );
  OR U43813 ( .A(n43499), .B(n43500), .Z(n43498) );
  NAND U43814 ( .A(n43500), .B(n43499), .Z(n43495) );
  ANDN U43815 ( .B(B[122]), .A(n69), .Z(n43279) );
  XNOR U43816 ( .A(n43287), .B(n43501), .Z(n43280) );
  XNOR U43817 ( .A(n43286), .B(n43284), .Z(n43501) );
  AND U43818 ( .A(n43502), .B(n43503), .Z(n43284) );
  NANDN U43819 ( .A(n43504), .B(n43505), .Z(n43503) );
  NANDN U43820 ( .A(n43506), .B(n43507), .Z(n43505) );
  NANDN U43821 ( .A(n43507), .B(n43506), .Z(n43502) );
  ANDN U43822 ( .B(B[123]), .A(n70), .Z(n43286) );
  XNOR U43823 ( .A(n43294), .B(n43508), .Z(n43287) );
  XNOR U43824 ( .A(n43293), .B(n43291), .Z(n43508) );
  AND U43825 ( .A(n43509), .B(n43510), .Z(n43291) );
  NANDN U43826 ( .A(n43511), .B(n43512), .Z(n43510) );
  OR U43827 ( .A(n43513), .B(n43514), .Z(n43512) );
  NAND U43828 ( .A(n43514), .B(n43513), .Z(n43509) );
  ANDN U43829 ( .B(B[124]), .A(n71), .Z(n43293) );
  XNOR U43830 ( .A(n43301), .B(n43515), .Z(n43294) );
  XNOR U43831 ( .A(n43300), .B(n43298), .Z(n43515) );
  AND U43832 ( .A(n43516), .B(n43517), .Z(n43298) );
  NANDN U43833 ( .A(n43518), .B(n43519), .Z(n43517) );
  NANDN U43834 ( .A(n43520), .B(n43521), .Z(n43519) );
  NANDN U43835 ( .A(n43521), .B(n43520), .Z(n43516) );
  ANDN U43836 ( .B(B[125]), .A(n72), .Z(n43300) );
  XNOR U43837 ( .A(n43308), .B(n43522), .Z(n43301) );
  XNOR U43838 ( .A(n43307), .B(n43305), .Z(n43522) );
  AND U43839 ( .A(n43523), .B(n43524), .Z(n43305) );
  NANDN U43840 ( .A(n43525), .B(n43526), .Z(n43524) );
  OR U43841 ( .A(n43527), .B(n43528), .Z(n43526) );
  NAND U43842 ( .A(n43528), .B(n43527), .Z(n43523) );
  ANDN U43843 ( .B(B[126]), .A(n73), .Z(n43307) );
  XNOR U43844 ( .A(n43315), .B(n43529), .Z(n43308) );
  XNOR U43845 ( .A(n43314), .B(n43312), .Z(n43529) );
  AND U43846 ( .A(n43530), .B(n43531), .Z(n43312) );
  NANDN U43847 ( .A(n43532), .B(n43533), .Z(n43531) );
  NANDN U43848 ( .A(n43534), .B(n43535), .Z(n43533) );
  NANDN U43849 ( .A(n43535), .B(n43534), .Z(n43530) );
  ANDN U43850 ( .B(B[127]), .A(n74), .Z(n43314) );
  XNOR U43851 ( .A(n43322), .B(n43536), .Z(n43315) );
  XNOR U43852 ( .A(n43321), .B(n43319), .Z(n43536) );
  AND U43853 ( .A(n43537), .B(n43538), .Z(n43319) );
  NANDN U43854 ( .A(n43539), .B(n43540), .Z(n43538) );
  OR U43855 ( .A(n43541), .B(n43542), .Z(n43540) );
  NAND U43856 ( .A(n43542), .B(n43541), .Z(n43537) );
  ANDN U43857 ( .B(B[128]), .A(n75), .Z(n43321) );
  XNOR U43858 ( .A(n43329), .B(n43543), .Z(n43322) );
  XNOR U43859 ( .A(n43328), .B(n43326), .Z(n43543) );
  AND U43860 ( .A(n43544), .B(n43545), .Z(n43326) );
  NANDN U43861 ( .A(n43546), .B(n43547), .Z(n43545) );
  NANDN U43862 ( .A(n43548), .B(n43549), .Z(n43547) );
  NANDN U43863 ( .A(n43549), .B(n43548), .Z(n43544) );
  ANDN U43864 ( .B(B[129]), .A(n76), .Z(n43328) );
  XNOR U43865 ( .A(n43336), .B(n43550), .Z(n43329) );
  XNOR U43866 ( .A(n43335), .B(n43333), .Z(n43550) );
  AND U43867 ( .A(n43551), .B(n43552), .Z(n43333) );
  NANDN U43868 ( .A(n43553), .B(n43554), .Z(n43552) );
  OR U43869 ( .A(n43555), .B(n43556), .Z(n43554) );
  NAND U43870 ( .A(n43556), .B(n43555), .Z(n43551) );
  ANDN U43871 ( .B(B[130]), .A(n77), .Z(n43335) );
  XNOR U43872 ( .A(n43343), .B(n43557), .Z(n43336) );
  XNOR U43873 ( .A(n43342), .B(n43340), .Z(n43557) );
  AND U43874 ( .A(n43558), .B(n43559), .Z(n43340) );
  NANDN U43875 ( .A(n43560), .B(n43561), .Z(n43559) );
  NANDN U43876 ( .A(n43562), .B(n43563), .Z(n43561) );
  NANDN U43877 ( .A(n43563), .B(n43562), .Z(n43558) );
  ANDN U43878 ( .B(B[131]), .A(n78), .Z(n43342) );
  XNOR U43879 ( .A(n43350), .B(n43564), .Z(n43343) );
  XNOR U43880 ( .A(n43349), .B(n43347), .Z(n43564) );
  AND U43881 ( .A(n43565), .B(n43566), .Z(n43347) );
  NANDN U43882 ( .A(n43567), .B(n43568), .Z(n43566) );
  OR U43883 ( .A(n43569), .B(n43570), .Z(n43568) );
  NAND U43884 ( .A(n43570), .B(n43569), .Z(n43565) );
  ANDN U43885 ( .B(B[132]), .A(n79), .Z(n43349) );
  XNOR U43886 ( .A(n43357), .B(n43571), .Z(n43350) );
  XNOR U43887 ( .A(n43356), .B(n43354), .Z(n43571) );
  AND U43888 ( .A(n43572), .B(n43573), .Z(n43354) );
  NANDN U43889 ( .A(n43574), .B(n43575), .Z(n43573) );
  NANDN U43890 ( .A(n43576), .B(n43577), .Z(n43575) );
  NANDN U43891 ( .A(n43577), .B(n43576), .Z(n43572) );
  ANDN U43892 ( .B(B[133]), .A(n80), .Z(n43356) );
  XNOR U43893 ( .A(n43364), .B(n43578), .Z(n43357) );
  XNOR U43894 ( .A(n43363), .B(n43361), .Z(n43578) );
  AND U43895 ( .A(n43579), .B(n43580), .Z(n43361) );
  NANDN U43896 ( .A(n43581), .B(n43582), .Z(n43580) );
  OR U43897 ( .A(n43583), .B(n43584), .Z(n43582) );
  NAND U43898 ( .A(n43584), .B(n43583), .Z(n43579) );
  ANDN U43899 ( .B(B[134]), .A(n81), .Z(n43363) );
  XNOR U43900 ( .A(n43371), .B(n43585), .Z(n43364) );
  XNOR U43901 ( .A(n43370), .B(n43368), .Z(n43585) );
  AND U43902 ( .A(n43586), .B(n43587), .Z(n43368) );
  NANDN U43903 ( .A(n43588), .B(n43589), .Z(n43587) );
  NAND U43904 ( .A(n43590), .B(n43591), .Z(n43589) );
  ANDN U43905 ( .B(B[135]), .A(n82), .Z(n43370) );
  XOR U43906 ( .A(n43377), .B(n43592), .Z(n43371) );
  XNOR U43907 ( .A(n43375), .B(n43378), .Z(n43592) );
  NAND U43908 ( .A(A[2]), .B(B[136]), .Z(n43378) );
  NANDN U43909 ( .A(n43593), .B(n43594), .Z(n43375) );
  AND U43910 ( .A(A[0]), .B(B[137]), .Z(n43594) );
  XNOR U43911 ( .A(n43380), .B(n43595), .Z(n43377) );
  NAND U43912 ( .A(A[0]), .B(B[138]), .Z(n43595) );
  NAND U43913 ( .A(B[137]), .B(A[1]), .Z(n43380) );
  NAND U43914 ( .A(n43596), .B(n43597), .Z(n520) );
  NANDN U43915 ( .A(n43598), .B(n43599), .Z(n43597) );
  OR U43916 ( .A(n43600), .B(n43601), .Z(n43599) );
  NAND U43917 ( .A(n43601), .B(n43600), .Z(n43596) );
  XOR U43918 ( .A(n522), .B(n521), .Z(\A1[135] ) );
  XOR U43919 ( .A(n43601), .B(n43602), .Z(n521) );
  XNOR U43920 ( .A(n43600), .B(n43598), .Z(n43602) );
  AND U43921 ( .A(n43603), .B(n43604), .Z(n43598) );
  NANDN U43922 ( .A(n43605), .B(n43606), .Z(n43604) );
  NANDN U43923 ( .A(n43607), .B(n43608), .Z(n43606) );
  NANDN U43924 ( .A(n43608), .B(n43607), .Z(n43603) );
  ANDN U43925 ( .B(B[106]), .A(n54), .Z(n43600) );
  XNOR U43926 ( .A(n43395), .B(n43609), .Z(n43601) );
  XNOR U43927 ( .A(n43394), .B(n43392), .Z(n43609) );
  AND U43928 ( .A(n43610), .B(n43611), .Z(n43392) );
  NANDN U43929 ( .A(n43612), .B(n43613), .Z(n43611) );
  OR U43930 ( .A(n43614), .B(n43615), .Z(n43613) );
  NAND U43931 ( .A(n43615), .B(n43614), .Z(n43610) );
  ANDN U43932 ( .B(B[107]), .A(n55), .Z(n43394) );
  XNOR U43933 ( .A(n43402), .B(n43616), .Z(n43395) );
  XNOR U43934 ( .A(n43401), .B(n43399), .Z(n43616) );
  AND U43935 ( .A(n43617), .B(n43618), .Z(n43399) );
  NANDN U43936 ( .A(n43619), .B(n43620), .Z(n43618) );
  NANDN U43937 ( .A(n43621), .B(n43622), .Z(n43620) );
  NANDN U43938 ( .A(n43622), .B(n43621), .Z(n43617) );
  ANDN U43939 ( .B(B[108]), .A(n56), .Z(n43401) );
  XNOR U43940 ( .A(n43409), .B(n43623), .Z(n43402) );
  XNOR U43941 ( .A(n43408), .B(n43406), .Z(n43623) );
  AND U43942 ( .A(n43624), .B(n43625), .Z(n43406) );
  NANDN U43943 ( .A(n43626), .B(n43627), .Z(n43625) );
  OR U43944 ( .A(n43628), .B(n43629), .Z(n43627) );
  NAND U43945 ( .A(n43629), .B(n43628), .Z(n43624) );
  ANDN U43946 ( .B(B[109]), .A(n57), .Z(n43408) );
  XNOR U43947 ( .A(n43416), .B(n43630), .Z(n43409) );
  XNOR U43948 ( .A(n43415), .B(n43413), .Z(n43630) );
  AND U43949 ( .A(n43631), .B(n43632), .Z(n43413) );
  NANDN U43950 ( .A(n43633), .B(n43634), .Z(n43632) );
  NANDN U43951 ( .A(n43635), .B(n43636), .Z(n43634) );
  NANDN U43952 ( .A(n43636), .B(n43635), .Z(n43631) );
  ANDN U43953 ( .B(B[110]), .A(n58), .Z(n43415) );
  XNOR U43954 ( .A(n43423), .B(n43637), .Z(n43416) );
  XNOR U43955 ( .A(n43422), .B(n43420), .Z(n43637) );
  AND U43956 ( .A(n43638), .B(n43639), .Z(n43420) );
  NANDN U43957 ( .A(n43640), .B(n43641), .Z(n43639) );
  OR U43958 ( .A(n43642), .B(n43643), .Z(n43641) );
  NAND U43959 ( .A(n43643), .B(n43642), .Z(n43638) );
  ANDN U43960 ( .B(B[111]), .A(n59), .Z(n43422) );
  XNOR U43961 ( .A(n43430), .B(n43644), .Z(n43423) );
  XNOR U43962 ( .A(n43429), .B(n43427), .Z(n43644) );
  AND U43963 ( .A(n43645), .B(n43646), .Z(n43427) );
  NANDN U43964 ( .A(n43647), .B(n43648), .Z(n43646) );
  NANDN U43965 ( .A(n43649), .B(n43650), .Z(n43648) );
  NANDN U43966 ( .A(n43650), .B(n43649), .Z(n43645) );
  ANDN U43967 ( .B(B[112]), .A(n60), .Z(n43429) );
  XNOR U43968 ( .A(n43437), .B(n43651), .Z(n43430) );
  XNOR U43969 ( .A(n43436), .B(n43434), .Z(n43651) );
  AND U43970 ( .A(n43652), .B(n43653), .Z(n43434) );
  NANDN U43971 ( .A(n43654), .B(n43655), .Z(n43653) );
  OR U43972 ( .A(n43656), .B(n43657), .Z(n43655) );
  NAND U43973 ( .A(n43657), .B(n43656), .Z(n43652) );
  ANDN U43974 ( .B(B[113]), .A(n61), .Z(n43436) );
  XNOR U43975 ( .A(n43444), .B(n43658), .Z(n43437) );
  XNOR U43976 ( .A(n43443), .B(n43441), .Z(n43658) );
  AND U43977 ( .A(n43659), .B(n43660), .Z(n43441) );
  NANDN U43978 ( .A(n43661), .B(n43662), .Z(n43660) );
  NANDN U43979 ( .A(n43663), .B(n43664), .Z(n43662) );
  NANDN U43980 ( .A(n43664), .B(n43663), .Z(n43659) );
  ANDN U43981 ( .B(B[114]), .A(n62), .Z(n43443) );
  XNOR U43982 ( .A(n43451), .B(n43665), .Z(n43444) );
  XNOR U43983 ( .A(n43450), .B(n43448), .Z(n43665) );
  AND U43984 ( .A(n43666), .B(n43667), .Z(n43448) );
  NANDN U43985 ( .A(n43668), .B(n43669), .Z(n43667) );
  OR U43986 ( .A(n43670), .B(n43671), .Z(n43669) );
  NAND U43987 ( .A(n43671), .B(n43670), .Z(n43666) );
  ANDN U43988 ( .B(B[115]), .A(n63), .Z(n43450) );
  XNOR U43989 ( .A(n43458), .B(n43672), .Z(n43451) );
  XNOR U43990 ( .A(n43457), .B(n43455), .Z(n43672) );
  AND U43991 ( .A(n43673), .B(n43674), .Z(n43455) );
  NANDN U43992 ( .A(n43675), .B(n43676), .Z(n43674) );
  NANDN U43993 ( .A(n43677), .B(n43678), .Z(n43676) );
  NANDN U43994 ( .A(n43678), .B(n43677), .Z(n43673) );
  ANDN U43995 ( .B(B[116]), .A(n64), .Z(n43457) );
  XNOR U43996 ( .A(n43465), .B(n43679), .Z(n43458) );
  XNOR U43997 ( .A(n43464), .B(n43462), .Z(n43679) );
  AND U43998 ( .A(n43680), .B(n43681), .Z(n43462) );
  NANDN U43999 ( .A(n43682), .B(n43683), .Z(n43681) );
  OR U44000 ( .A(n43684), .B(n43685), .Z(n43683) );
  NAND U44001 ( .A(n43685), .B(n43684), .Z(n43680) );
  ANDN U44002 ( .B(B[117]), .A(n65), .Z(n43464) );
  XNOR U44003 ( .A(n43472), .B(n43686), .Z(n43465) );
  XNOR U44004 ( .A(n43471), .B(n43469), .Z(n43686) );
  AND U44005 ( .A(n43687), .B(n43688), .Z(n43469) );
  NANDN U44006 ( .A(n43689), .B(n43690), .Z(n43688) );
  NANDN U44007 ( .A(n43691), .B(n43692), .Z(n43690) );
  NANDN U44008 ( .A(n43692), .B(n43691), .Z(n43687) );
  ANDN U44009 ( .B(B[118]), .A(n66), .Z(n43471) );
  XNOR U44010 ( .A(n43479), .B(n43693), .Z(n43472) );
  XNOR U44011 ( .A(n43478), .B(n43476), .Z(n43693) );
  AND U44012 ( .A(n43694), .B(n43695), .Z(n43476) );
  NANDN U44013 ( .A(n43696), .B(n43697), .Z(n43695) );
  OR U44014 ( .A(n43698), .B(n43699), .Z(n43697) );
  NAND U44015 ( .A(n43699), .B(n43698), .Z(n43694) );
  ANDN U44016 ( .B(B[119]), .A(n67), .Z(n43478) );
  XNOR U44017 ( .A(n43486), .B(n43700), .Z(n43479) );
  XNOR U44018 ( .A(n43485), .B(n43483), .Z(n43700) );
  AND U44019 ( .A(n43701), .B(n43702), .Z(n43483) );
  NANDN U44020 ( .A(n43703), .B(n43704), .Z(n43702) );
  NANDN U44021 ( .A(n43705), .B(n43706), .Z(n43704) );
  NANDN U44022 ( .A(n43706), .B(n43705), .Z(n43701) );
  ANDN U44023 ( .B(B[120]), .A(n68), .Z(n43485) );
  XNOR U44024 ( .A(n43493), .B(n43707), .Z(n43486) );
  XNOR U44025 ( .A(n43492), .B(n43490), .Z(n43707) );
  AND U44026 ( .A(n43708), .B(n43709), .Z(n43490) );
  NANDN U44027 ( .A(n43710), .B(n43711), .Z(n43709) );
  OR U44028 ( .A(n43712), .B(n43713), .Z(n43711) );
  NAND U44029 ( .A(n43713), .B(n43712), .Z(n43708) );
  ANDN U44030 ( .B(B[121]), .A(n69), .Z(n43492) );
  XNOR U44031 ( .A(n43500), .B(n43714), .Z(n43493) );
  XNOR U44032 ( .A(n43499), .B(n43497), .Z(n43714) );
  AND U44033 ( .A(n43715), .B(n43716), .Z(n43497) );
  NANDN U44034 ( .A(n43717), .B(n43718), .Z(n43716) );
  NANDN U44035 ( .A(n43719), .B(n43720), .Z(n43718) );
  NANDN U44036 ( .A(n43720), .B(n43719), .Z(n43715) );
  ANDN U44037 ( .B(B[122]), .A(n70), .Z(n43499) );
  XNOR U44038 ( .A(n43507), .B(n43721), .Z(n43500) );
  XNOR U44039 ( .A(n43506), .B(n43504), .Z(n43721) );
  AND U44040 ( .A(n43722), .B(n43723), .Z(n43504) );
  NANDN U44041 ( .A(n43724), .B(n43725), .Z(n43723) );
  OR U44042 ( .A(n43726), .B(n43727), .Z(n43725) );
  NAND U44043 ( .A(n43727), .B(n43726), .Z(n43722) );
  ANDN U44044 ( .B(B[123]), .A(n71), .Z(n43506) );
  XNOR U44045 ( .A(n43514), .B(n43728), .Z(n43507) );
  XNOR U44046 ( .A(n43513), .B(n43511), .Z(n43728) );
  AND U44047 ( .A(n43729), .B(n43730), .Z(n43511) );
  NANDN U44048 ( .A(n43731), .B(n43732), .Z(n43730) );
  NANDN U44049 ( .A(n43733), .B(n43734), .Z(n43732) );
  NANDN U44050 ( .A(n43734), .B(n43733), .Z(n43729) );
  ANDN U44051 ( .B(B[124]), .A(n72), .Z(n43513) );
  XNOR U44052 ( .A(n43521), .B(n43735), .Z(n43514) );
  XNOR U44053 ( .A(n43520), .B(n43518), .Z(n43735) );
  AND U44054 ( .A(n43736), .B(n43737), .Z(n43518) );
  NANDN U44055 ( .A(n43738), .B(n43739), .Z(n43737) );
  OR U44056 ( .A(n43740), .B(n43741), .Z(n43739) );
  NAND U44057 ( .A(n43741), .B(n43740), .Z(n43736) );
  ANDN U44058 ( .B(B[125]), .A(n73), .Z(n43520) );
  XNOR U44059 ( .A(n43528), .B(n43742), .Z(n43521) );
  XNOR U44060 ( .A(n43527), .B(n43525), .Z(n43742) );
  AND U44061 ( .A(n43743), .B(n43744), .Z(n43525) );
  NANDN U44062 ( .A(n43745), .B(n43746), .Z(n43744) );
  NANDN U44063 ( .A(n43747), .B(n43748), .Z(n43746) );
  NANDN U44064 ( .A(n43748), .B(n43747), .Z(n43743) );
  ANDN U44065 ( .B(B[126]), .A(n74), .Z(n43527) );
  XNOR U44066 ( .A(n43535), .B(n43749), .Z(n43528) );
  XNOR U44067 ( .A(n43534), .B(n43532), .Z(n43749) );
  AND U44068 ( .A(n43750), .B(n43751), .Z(n43532) );
  NANDN U44069 ( .A(n43752), .B(n43753), .Z(n43751) );
  OR U44070 ( .A(n43754), .B(n43755), .Z(n43753) );
  NAND U44071 ( .A(n43755), .B(n43754), .Z(n43750) );
  ANDN U44072 ( .B(B[127]), .A(n75), .Z(n43534) );
  XNOR U44073 ( .A(n43542), .B(n43756), .Z(n43535) );
  XNOR U44074 ( .A(n43541), .B(n43539), .Z(n43756) );
  AND U44075 ( .A(n43757), .B(n43758), .Z(n43539) );
  NANDN U44076 ( .A(n43759), .B(n43760), .Z(n43758) );
  NANDN U44077 ( .A(n43761), .B(n43762), .Z(n43760) );
  NANDN U44078 ( .A(n43762), .B(n43761), .Z(n43757) );
  ANDN U44079 ( .B(B[128]), .A(n76), .Z(n43541) );
  XNOR U44080 ( .A(n43549), .B(n43763), .Z(n43542) );
  XNOR U44081 ( .A(n43548), .B(n43546), .Z(n43763) );
  AND U44082 ( .A(n43764), .B(n43765), .Z(n43546) );
  NANDN U44083 ( .A(n43766), .B(n43767), .Z(n43765) );
  OR U44084 ( .A(n43768), .B(n43769), .Z(n43767) );
  NAND U44085 ( .A(n43769), .B(n43768), .Z(n43764) );
  ANDN U44086 ( .B(B[129]), .A(n77), .Z(n43548) );
  XNOR U44087 ( .A(n43556), .B(n43770), .Z(n43549) );
  XNOR U44088 ( .A(n43555), .B(n43553), .Z(n43770) );
  AND U44089 ( .A(n43771), .B(n43772), .Z(n43553) );
  NANDN U44090 ( .A(n43773), .B(n43774), .Z(n43772) );
  NANDN U44091 ( .A(n43775), .B(n43776), .Z(n43774) );
  NANDN U44092 ( .A(n43776), .B(n43775), .Z(n43771) );
  ANDN U44093 ( .B(B[130]), .A(n78), .Z(n43555) );
  XNOR U44094 ( .A(n43563), .B(n43777), .Z(n43556) );
  XNOR U44095 ( .A(n43562), .B(n43560), .Z(n43777) );
  AND U44096 ( .A(n43778), .B(n43779), .Z(n43560) );
  NANDN U44097 ( .A(n43780), .B(n43781), .Z(n43779) );
  OR U44098 ( .A(n43782), .B(n43783), .Z(n43781) );
  NAND U44099 ( .A(n43783), .B(n43782), .Z(n43778) );
  ANDN U44100 ( .B(B[131]), .A(n79), .Z(n43562) );
  XNOR U44101 ( .A(n43570), .B(n43784), .Z(n43563) );
  XNOR U44102 ( .A(n43569), .B(n43567), .Z(n43784) );
  AND U44103 ( .A(n43785), .B(n43786), .Z(n43567) );
  NANDN U44104 ( .A(n43787), .B(n43788), .Z(n43786) );
  NANDN U44105 ( .A(n43789), .B(n43790), .Z(n43788) );
  NANDN U44106 ( .A(n43790), .B(n43789), .Z(n43785) );
  ANDN U44107 ( .B(B[132]), .A(n80), .Z(n43569) );
  XNOR U44108 ( .A(n43577), .B(n43791), .Z(n43570) );
  XNOR U44109 ( .A(n43576), .B(n43574), .Z(n43791) );
  AND U44110 ( .A(n43792), .B(n43793), .Z(n43574) );
  NANDN U44111 ( .A(n43794), .B(n43795), .Z(n43793) );
  OR U44112 ( .A(n43796), .B(n43797), .Z(n43795) );
  NAND U44113 ( .A(n43797), .B(n43796), .Z(n43792) );
  ANDN U44114 ( .B(B[133]), .A(n81), .Z(n43576) );
  XNOR U44115 ( .A(n43584), .B(n43798), .Z(n43577) );
  XNOR U44116 ( .A(n43583), .B(n43581), .Z(n43798) );
  AND U44117 ( .A(n43799), .B(n43800), .Z(n43581) );
  NANDN U44118 ( .A(n43801), .B(n43802), .Z(n43800) );
  NAND U44119 ( .A(n43803), .B(n43804), .Z(n43802) );
  ANDN U44120 ( .B(B[134]), .A(n82), .Z(n43583) );
  XOR U44121 ( .A(n43590), .B(n43805), .Z(n43584) );
  XNOR U44122 ( .A(n43588), .B(n43591), .Z(n43805) );
  NAND U44123 ( .A(A[2]), .B(B[135]), .Z(n43591) );
  NANDN U44124 ( .A(n43806), .B(n43807), .Z(n43588) );
  AND U44125 ( .A(A[0]), .B(B[136]), .Z(n43807) );
  XNOR U44126 ( .A(n43593), .B(n43808), .Z(n43590) );
  NAND U44127 ( .A(A[0]), .B(B[137]), .Z(n43808) );
  NAND U44128 ( .A(B[136]), .B(A[1]), .Z(n43593) );
  NAND U44129 ( .A(n43809), .B(n43810), .Z(n522) );
  NANDN U44130 ( .A(n43811), .B(n43812), .Z(n43810) );
  OR U44131 ( .A(n43813), .B(n43814), .Z(n43812) );
  NAND U44132 ( .A(n43814), .B(n43813), .Z(n43809) );
  XOR U44133 ( .A(n524), .B(n523), .Z(\A1[134] ) );
  XOR U44134 ( .A(n43814), .B(n43815), .Z(n523) );
  XNOR U44135 ( .A(n43813), .B(n43811), .Z(n43815) );
  AND U44136 ( .A(n43816), .B(n43817), .Z(n43811) );
  NANDN U44137 ( .A(n43818), .B(n43819), .Z(n43817) );
  NANDN U44138 ( .A(n43820), .B(n43821), .Z(n43819) );
  NANDN U44139 ( .A(n43821), .B(n43820), .Z(n43816) );
  ANDN U44140 ( .B(B[105]), .A(n54), .Z(n43813) );
  XNOR U44141 ( .A(n43608), .B(n43822), .Z(n43814) );
  XNOR U44142 ( .A(n43607), .B(n43605), .Z(n43822) );
  AND U44143 ( .A(n43823), .B(n43824), .Z(n43605) );
  NANDN U44144 ( .A(n43825), .B(n43826), .Z(n43824) );
  OR U44145 ( .A(n43827), .B(n43828), .Z(n43826) );
  NAND U44146 ( .A(n43828), .B(n43827), .Z(n43823) );
  ANDN U44147 ( .B(B[106]), .A(n55), .Z(n43607) );
  XNOR U44148 ( .A(n43615), .B(n43829), .Z(n43608) );
  XNOR U44149 ( .A(n43614), .B(n43612), .Z(n43829) );
  AND U44150 ( .A(n43830), .B(n43831), .Z(n43612) );
  NANDN U44151 ( .A(n43832), .B(n43833), .Z(n43831) );
  NANDN U44152 ( .A(n43834), .B(n43835), .Z(n43833) );
  NANDN U44153 ( .A(n43835), .B(n43834), .Z(n43830) );
  ANDN U44154 ( .B(B[107]), .A(n56), .Z(n43614) );
  XNOR U44155 ( .A(n43622), .B(n43836), .Z(n43615) );
  XNOR U44156 ( .A(n43621), .B(n43619), .Z(n43836) );
  AND U44157 ( .A(n43837), .B(n43838), .Z(n43619) );
  NANDN U44158 ( .A(n43839), .B(n43840), .Z(n43838) );
  OR U44159 ( .A(n43841), .B(n43842), .Z(n43840) );
  NAND U44160 ( .A(n43842), .B(n43841), .Z(n43837) );
  ANDN U44161 ( .B(B[108]), .A(n57), .Z(n43621) );
  XNOR U44162 ( .A(n43629), .B(n43843), .Z(n43622) );
  XNOR U44163 ( .A(n43628), .B(n43626), .Z(n43843) );
  AND U44164 ( .A(n43844), .B(n43845), .Z(n43626) );
  NANDN U44165 ( .A(n43846), .B(n43847), .Z(n43845) );
  NANDN U44166 ( .A(n43848), .B(n43849), .Z(n43847) );
  NANDN U44167 ( .A(n43849), .B(n43848), .Z(n43844) );
  ANDN U44168 ( .B(B[109]), .A(n58), .Z(n43628) );
  XNOR U44169 ( .A(n43636), .B(n43850), .Z(n43629) );
  XNOR U44170 ( .A(n43635), .B(n43633), .Z(n43850) );
  AND U44171 ( .A(n43851), .B(n43852), .Z(n43633) );
  NANDN U44172 ( .A(n43853), .B(n43854), .Z(n43852) );
  OR U44173 ( .A(n43855), .B(n43856), .Z(n43854) );
  NAND U44174 ( .A(n43856), .B(n43855), .Z(n43851) );
  ANDN U44175 ( .B(B[110]), .A(n59), .Z(n43635) );
  XNOR U44176 ( .A(n43643), .B(n43857), .Z(n43636) );
  XNOR U44177 ( .A(n43642), .B(n43640), .Z(n43857) );
  AND U44178 ( .A(n43858), .B(n43859), .Z(n43640) );
  NANDN U44179 ( .A(n43860), .B(n43861), .Z(n43859) );
  NANDN U44180 ( .A(n43862), .B(n43863), .Z(n43861) );
  NANDN U44181 ( .A(n43863), .B(n43862), .Z(n43858) );
  ANDN U44182 ( .B(B[111]), .A(n60), .Z(n43642) );
  XNOR U44183 ( .A(n43650), .B(n43864), .Z(n43643) );
  XNOR U44184 ( .A(n43649), .B(n43647), .Z(n43864) );
  AND U44185 ( .A(n43865), .B(n43866), .Z(n43647) );
  NANDN U44186 ( .A(n43867), .B(n43868), .Z(n43866) );
  OR U44187 ( .A(n43869), .B(n43870), .Z(n43868) );
  NAND U44188 ( .A(n43870), .B(n43869), .Z(n43865) );
  ANDN U44189 ( .B(B[112]), .A(n61), .Z(n43649) );
  XNOR U44190 ( .A(n43657), .B(n43871), .Z(n43650) );
  XNOR U44191 ( .A(n43656), .B(n43654), .Z(n43871) );
  AND U44192 ( .A(n43872), .B(n43873), .Z(n43654) );
  NANDN U44193 ( .A(n43874), .B(n43875), .Z(n43873) );
  NANDN U44194 ( .A(n43876), .B(n43877), .Z(n43875) );
  NANDN U44195 ( .A(n43877), .B(n43876), .Z(n43872) );
  ANDN U44196 ( .B(B[113]), .A(n62), .Z(n43656) );
  XNOR U44197 ( .A(n43664), .B(n43878), .Z(n43657) );
  XNOR U44198 ( .A(n43663), .B(n43661), .Z(n43878) );
  AND U44199 ( .A(n43879), .B(n43880), .Z(n43661) );
  NANDN U44200 ( .A(n43881), .B(n43882), .Z(n43880) );
  OR U44201 ( .A(n43883), .B(n43884), .Z(n43882) );
  NAND U44202 ( .A(n43884), .B(n43883), .Z(n43879) );
  ANDN U44203 ( .B(B[114]), .A(n63), .Z(n43663) );
  XNOR U44204 ( .A(n43671), .B(n43885), .Z(n43664) );
  XNOR U44205 ( .A(n43670), .B(n43668), .Z(n43885) );
  AND U44206 ( .A(n43886), .B(n43887), .Z(n43668) );
  NANDN U44207 ( .A(n43888), .B(n43889), .Z(n43887) );
  NANDN U44208 ( .A(n43890), .B(n43891), .Z(n43889) );
  NANDN U44209 ( .A(n43891), .B(n43890), .Z(n43886) );
  ANDN U44210 ( .B(B[115]), .A(n64), .Z(n43670) );
  XNOR U44211 ( .A(n43678), .B(n43892), .Z(n43671) );
  XNOR U44212 ( .A(n43677), .B(n43675), .Z(n43892) );
  AND U44213 ( .A(n43893), .B(n43894), .Z(n43675) );
  NANDN U44214 ( .A(n43895), .B(n43896), .Z(n43894) );
  OR U44215 ( .A(n43897), .B(n43898), .Z(n43896) );
  NAND U44216 ( .A(n43898), .B(n43897), .Z(n43893) );
  ANDN U44217 ( .B(B[116]), .A(n65), .Z(n43677) );
  XNOR U44218 ( .A(n43685), .B(n43899), .Z(n43678) );
  XNOR U44219 ( .A(n43684), .B(n43682), .Z(n43899) );
  AND U44220 ( .A(n43900), .B(n43901), .Z(n43682) );
  NANDN U44221 ( .A(n43902), .B(n43903), .Z(n43901) );
  NANDN U44222 ( .A(n43904), .B(n43905), .Z(n43903) );
  NANDN U44223 ( .A(n43905), .B(n43904), .Z(n43900) );
  ANDN U44224 ( .B(B[117]), .A(n66), .Z(n43684) );
  XNOR U44225 ( .A(n43692), .B(n43906), .Z(n43685) );
  XNOR U44226 ( .A(n43691), .B(n43689), .Z(n43906) );
  AND U44227 ( .A(n43907), .B(n43908), .Z(n43689) );
  NANDN U44228 ( .A(n43909), .B(n43910), .Z(n43908) );
  OR U44229 ( .A(n43911), .B(n43912), .Z(n43910) );
  NAND U44230 ( .A(n43912), .B(n43911), .Z(n43907) );
  ANDN U44231 ( .B(B[118]), .A(n67), .Z(n43691) );
  XNOR U44232 ( .A(n43699), .B(n43913), .Z(n43692) );
  XNOR U44233 ( .A(n43698), .B(n43696), .Z(n43913) );
  AND U44234 ( .A(n43914), .B(n43915), .Z(n43696) );
  NANDN U44235 ( .A(n43916), .B(n43917), .Z(n43915) );
  NANDN U44236 ( .A(n43918), .B(n43919), .Z(n43917) );
  NANDN U44237 ( .A(n43919), .B(n43918), .Z(n43914) );
  ANDN U44238 ( .B(B[119]), .A(n68), .Z(n43698) );
  XNOR U44239 ( .A(n43706), .B(n43920), .Z(n43699) );
  XNOR U44240 ( .A(n43705), .B(n43703), .Z(n43920) );
  AND U44241 ( .A(n43921), .B(n43922), .Z(n43703) );
  NANDN U44242 ( .A(n43923), .B(n43924), .Z(n43922) );
  OR U44243 ( .A(n43925), .B(n43926), .Z(n43924) );
  NAND U44244 ( .A(n43926), .B(n43925), .Z(n43921) );
  ANDN U44245 ( .B(B[120]), .A(n69), .Z(n43705) );
  XNOR U44246 ( .A(n43713), .B(n43927), .Z(n43706) );
  XNOR U44247 ( .A(n43712), .B(n43710), .Z(n43927) );
  AND U44248 ( .A(n43928), .B(n43929), .Z(n43710) );
  NANDN U44249 ( .A(n43930), .B(n43931), .Z(n43929) );
  NANDN U44250 ( .A(n43932), .B(n43933), .Z(n43931) );
  NANDN U44251 ( .A(n43933), .B(n43932), .Z(n43928) );
  ANDN U44252 ( .B(B[121]), .A(n70), .Z(n43712) );
  XNOR U44253 ( .A(n43720), .B(n43934), .Z(n43713) );
  XNOR U44254 ( .A(n43719), .B(n43717), .Z(n43934) );
  AND U44255 ( .A(n43935), .B(n43936), .Z(n43717) );
  NANDN U44256 ( .A(n43937), .B(n43938), .Z(n43936) );
  OR U44257 ( .A(n43939), .B(n43940), .Z(n43938) );
  NAND U44258 ( .A(n43940), .B(n43939), .Z(n43935) );
  ANDN U44259 ( .B(B[122]), .A(n71), .Z(n43719) );
  XNOR U44260 ( .A(n43727), .B(n43941), .Z(n43720) );
  XNOR U44261 ( .A(n43726), .B(n43724), .Z(n43941) );
  AND U44262 ( .A(n43942), .B(n43943), .Z(n43724) );
  NANDN U44263 ( .A(n43944), .B(n43945), .Z(n43943) );
  NANDN U44264 ( .A(n43946), .B(n43947), .Z(n43945) );
  NANDN U44265 ( .A(n43947), .B(n43946), .Z(n43942) );
  ANDN U44266 ( .B(B[123]), .A(n72), .Z(n43726) );
  XNOR U44267 ( .A(n43734), .B(n43948), .Z(n43727) );
  XNOR U44268 ( .A(n43733), .B(n43731), .Z(n43948) );
  AND U44269 ( .A(n43949), .B(n43950), .Z(n43731) );
  NANDN U44270 ( .A(n43951), .B(n43952), .Z(n43950) );
  OR U44271 ( .A(n43953), .B(n43954), .Z(n43952) );
  NAND U44272 ( .A(n43954), .B(n43953), .Z(n43949) );
  ANDN U44273 ( .B(B[124]), .A(n73), .Z(n43733) );
  XNOR U44274 ( .A(n43741), .B(n43955), .Z(n43734) );
  XNOR U44275 ( .A(n43740), .B(n43738), .Z(n43955) );
  AND U44276 ( .A(n43956), .B(n43957), .Z(n43738) );
  NANDN U44277 ( .A(n43958), .B(n43959), .Z(n43957) );
  NANDN U44278 ( .A(n43960), .B(n43961), .Z(n43959) );
  NANDN U44279 ( .A(n43961), .B(n43960), .Z(n43956) );
  ANDN U44280 ( .B(B[125]), .A(n74), .Z(n43740) );
  XNOR U44281 ( .A(n43748), .B(n43962), .Z(n43741) );
  XNOR U44282 ( .A(n43747), .B(n43745), .Z(n43962) );
  AND U44283 ( .A(n43963), .B(n43964), .Z(n43745) );
  NANDN U44284 ( .A(n43965), .B(n43966), .Z(n43964) );
  OR U44285 ( .A(n43967), .B(n43968), .Z(n43966) );
  NAND U44286 ( .A(n43968), .B(n43967), .Z(n43963) );
  ANDN U44287 ( .B(B[126]), .A(n75), .Z(n43747) );
  XNOR U44288 ( .A(n43755), .B(n43969), .Z(n43748) );
  XNOR U44289 ( .A(n43754), .B(n43752), .Z(n43969) );
  AND U44290 ( .A(n43970), .B(n43971), .Z(n43752) );
  NANDN U44291 ( .A(n43972), .B(n43973), .Z(n43971) );
  NANDN U44292 ( .A(n43974), .B(n43975), .Z(n43973) );
  NANDN U44293 ( .A(n43975), .B(n43974), .Z(n43970) );
  ANDN U44294 ( .B(B[127]), .A(n76), .Z(n43754) );
  XNOR U44295 ( .A(n43762), .B(n43976), .Z(n43755) );
  XNOR U44296 ( .A(n43761), .B(n43759), .Z(n43976) );
  AND U44297 ( .A(n43977), .B(n43978), .Z(n43759) );
  NANDN U44298 ( .A(n43979), .B(n43980), .Z(n43978) );
  OR U44299 ( .A(n43981), .B(n43982), .Z(n43980) );
  NAND U44300 ( .A(n43982), .B(n43981), .Z(n43977) );
  ANDN U44301 ( .B(B[128]), .A(n77), .Z(n43761) );
  XNOR U44302 ( .A(n43769), .B(n43983), .Z(n43762) );
  XNOR U44303 ( .A(n43768), .B(n43766), .Z(n43983) );
  AND U44304 ( .A(n43984), .B(n43985), .Z(n43766) );
  NANDN U44305 ( .A(n43986), .B(n43987), .Z(n43985) );
  NANDN U44306 ( .A(n43988), .B(n43989), .Z(n43987) );
  NANDN U44307 ( .A(n43989), .B(n43988), .Z(n43984) );
  ANDN U44308 ( .B(B[129]), .A(n78), .Z(n43768) );
  XNOR U44309 ( .A(n43776), .B(n43990), .Z(n43769) );
  XNOR U44310 ( .A(n43775), .B(n43773), .Z(n43990) );
  AND U44311 ( .A(n43991), .B(n43992), .Z(n43773) );
  NANDN U44312 ( .A(n43993), .B(n43994), .Z(n43992) );
  OR U44313 ( .A(n43995), .B(n43996), .Z(n43994) );
  NAND U44314 ( .A(n43996), .B(n43995), .Z(n43991) );
  ANDN U44315 ( .B(B[130]), .A(n79), .Z(n43775) );
  XNOR U44316 ( .A(n43783), .B(n43997), .Z(n43776) );
  XNOR U44317 ( .A(n43782), .B(n43780), .Z(n43997) );
  AND U44318 ( .A(n43998), .B(n43999), .Z(n43780) );
  NANDN U44319 ( .A(n44000), .B(n44001), .Z(n43999) );
  NANDN U44320 ( .A(n44002), .B(n44003), .Z(n44001) );
  NANDN U44321 ( .A(n44003), .B(n44002), .Z(n43998) );
  ANDN U44322 ( .B(B[131]), .A(n80), .Z(n43782) );
  XNOR U44323 ( .A(n43790), .B(n44004), .Z(n43783) );
  XNOR U44324 ( .A(n43789), .B(n43787), .Z(n44004) );
  AND U44325 ( .A(n44005), .B(n44006), .Z(n43787) );
  NANDN U44326 ( .A(n44007), .B(n44008), .Z(n44006) );
  OR U44327 ( .A(n44009), .B(n44010), .Z(n44008) );
  NAND U44328 ( .A(n44010), .B(n44009), .Z(n44005) );
  ANDN U44329 ( .B(B[132]), .A(n81), .Z(n43789) );
  XNOR U44330 ( .A(n43797), .B(n44011), .Z(n43790) );
  XNOR U44331 ( .A(n43796), .B(n43794), .Z(n44011) );
  AND U44332 ( .A(n44012), .B(n44013), .Z(n43794) );
  NANDN U44333 ( .A(n44014), .B(n44015), .Z(n44013) );
  NAND U44334 ( .A(n44016), .B(n44017), .Z(n44015) );
  ANDN U44335 ( .B(B[133]), .A(n82), .Z(n43796) );
  XOR U44336 ( .A(n43803), .B(n44018), .Z(n43797) );
  XNOR U44337 ( .A(n43801), .B(n43804), .Z(n44018) );
  NAND U44338 ( .A(A[2]), .B(B[134]), .Z(n43804) );
  NANDN U44339 ( .A(n44019), .B(n44020), .Z(n43801) );
  AND U44340 ( .A(A[0]), .B(B[135]), .Z(n44020) );
  XNOR U44341 ( .A(n43806), .B(n44021), .Z(n43803) );
  NAND U44342 ( .A(A[0]), .B(B[136]), .Z(n44021) );
  NAND U44343 ( .A(B[135]), .B(A[1]), .Z(n43806) );
  NAND U44344 ( .A(n44022), .B(n44023), .Z(n524) );
  NANDN U44345 ( .A(n44024), .B(n44025), .Z(n44023) );
  OR U44346 ( .A(n44026), .B(n44027), .Z(n44025) );
  NAND U44347 ( .A(n44027), .B(n44026), .Z(n44022) );
  XOR U44348 ( .A(n526), .B(n525), .Z(\A1[133] ) );
  XOR U44349 ( .A(n44027), .B(n44028), .Z(n525) );
  XNOR U44350 ( .A(n44026), .B(n44024), .Z(n44028) );
  AND U44351 ( .A(n44029), .B(n44030), .Z(n44024) );
  NANDN U44352 ( .A(n44031), .B(n44032), .Z(n44030) );
  NANDN U44353 ( .A(n44033), .B(n44034), .Z(n44032) );
  NANDN U44354 ( .A(n44034), .B(n44033), .Z(n44029) );
  ANDN U44355 ( .B(B[104]), .A(n54), .Z(n44026) );
  XNOR U44356 ( .A(n43821), .B(n44035), .Z(n44027) );
  XNOR U44357 ( .A(n43820), .B(n43818), .Z(n44035) );
  AND U44358 ( .A(n44036), .B(n44037), .Z(n43818) );
  NANDN U44359 ( .A(n44038), .B(n44039), .Z(n44037) );
  OR U44360 ( .A(n44040), .B(n44041), .Z(n44039) );
  NAND U44361 ( .A(n44041), .B(n44040), .Z(n44036) );
  ANDN U44362 ( .B(B[105]), .A(n55), .Z(n43820) );
  XNOR U44363 ( .A(n43828), .B(n44042), .Z(n43821) );
  XNOR U44364 ( .A(n43827), .B(n43825), .Z(n44042) );
  AND U44365 ( .A(n44043), .B(n44044), .Z(n43825) );
  NANDN U44366 ( .A(n44045), .B(n44046), .Z(n44044) );
  NANDN U44367 ( .A(n44047), .B(n44048), .Z(n44046) );
  NANDN U44368 ( .A(n44048), .B(n44047), .Z(n44043) );
  ANDN U44369 ( .B(B[106]), .A(n56), .Z(n43827) );
  XNOR U44370 ( .A(n43835), .B(n44049), .Z(n43828) );
  XNOR U44371 ( .A(n43834), .B(n43832), .Z(n44049) );
  AND U44372 ( .A(n44050), .B(n44051), .Z(n43832) );
  NANDN U44373 ( .A(n44052), .B(n44053), .Z(n44051) );
  OR U44374 ( .A(n44054), .B(n44055), .Z(n44053) );
  NAND U44375 ( .A(n44055), .B(n44054), .Z(n44050) );
  ANDN U44376 ( .B(B[107]), .A(n57), .Z(n43834) );
  XNOR U44377 ( .A(n43842), .B(n44056), .Z(n43835) );
  XNOR U44378 ( .A(n43841), .B(n43839), .Z(n44056) );
  AND U44379 ( .A(n44057), .B(n44058), .Z(n43839) );
  NANDN U44380 ( .A(n44059), .B(n44060), .Z(n44058) );
  NANDN U44381 ( .A(n44061), .B(n44062), .Z(n44060) );
  NANDN U44382 ( .A(n44062), .B(n44061), .Z(n44057) );
  ANDN U44383 ( .B(B[108]), .A(n58), .Z(n43841) );
  XNOR U44384 ( .A(n43849), .B(n44063), .Z(n43842) );
  XNOR U44385 ( .A(n43848), .B(n43846), .Z(n44063) );
  AND U44386 ( .A(n44064), .B(n44065), .Z(n43846) );
  NANDN U44387 ( .A(n44066), .B(n44067), .Z(n44065) );
  OR U44388 ( .A(n44068), .B(n44069), .Z(n44067) );
  NAND U44389 ( .A(n44069), .B(n44068), .Z(n44064) );
  ANDN U44390 ( .B(B[109]), .A(n59), .Z(n43848) );
  XNOR U44391 ( .A(n43856), .B(n44070), .Z(n43849) );
  XNOR U44392 ( .A(n43855), .B(n43853), .Z(n44070) );
  AND U44393 ( .A(n44071), .B(n44072), .Z(n43853) );
  NANDN U44394 ( .A(n44073), .B(n44074), .Z(n44072) );
  NANDN U44395 ( .A(n44075), .B(n44076), .Z(n44074) );
  NANDN U44396 ( .A(n44076), .B(n44075), .Z(n44071) );
  ANDN U44397 ( .B(B[110]), .A(n60), .Z(n43855) );
  XNOR U44398 ( .A(n43863), .B(n44077), .Z(n43856) );
  XNOR U44399 ( .A(n43862), .B(n43860), .Z(n44077) );
  AND U44400 ( .A(n44078), .B(n44079), .Z(n43860) );
  NANDN U44401 ( .A(n44080), .B(n44081), .Z(n44079) );
  OR U44402 ( .A(n44082), .B(n44083), .Z(n44081) );
  NAND U44403 ( .A(n44083), .B(n44082), .Z(n44078) );
  ANDN U44404 ( .B(B[111]), .A(n61), .Z(n43862) );
  XNOR U44405 ( .A(n43870), .B(n44084), .Z(n43863) );
  XNOR U44406 ( .A(n43869), .B(n43867), .Z(n44084) );
  AND U44407 ( .A(n44085), .B(n44086), .Z(n43867) );
  NANDN U44408 ( .A(n44087), .B(n44088), .Z(n44086) );
  NANDN U44409 ( .A(n44089), .B(n44090), .Z(n44088) );
  NANDN U44410 ( .A(n44090), .B(n44089), .Z(n44085) );
  ANDN U44411 ( .B(B[112]), .A(n62), .Z(n43869) );
  XNOR U44412 ( .A(n43877), .B(n44091), .Z(n43870) );
  XNOR U44413 ( .A(n43876), .B(n43874), .Z(n44091) );
  AND U44414 ( .A(n44092), .B(n44093), .Z(n43874) );
  NANDN U44415 ( .A(n44094), .B(n44095), .Z(n44093) );
  OR U44416 ( .A(n44096), .B(n44097), .Z(n44095) );
  NAND U44417 ( .A(n44097), .B(n44096), .Z(n44092) );
  ANDN U44418 ( .B(B[113]), .A(n63), .Z(n43876) );
  XNOR U44419 ( .A(n43884), .B(n44098), .Z(n43877) );
  XNOR U44420 ( .A(n43883), .B(n43881), .Z(n44098) );
  AND U44421 ( .A(n44099), .B(n44100), .Z(n43881) );
  NANDN U44422 ( .A(n44101), .B(n44102), .Z(n44100) );
  NANDN U44423 ( .A(n44103), .B(n44104), .Z(n44102) );
  NANDN U44424 ( .A(n44104), .B(n44103), .Z(n44099) );
  ANDN U44425 ( .B(B[114]), .A(n64), .Z(n43883) );
  XNOR U44426 ( .A(n43891), .B(n44105), .Z(n43884) );
  XNOR U44427 ( .A(n43890), .B(n43888), .Z(n44105) );
  AND U44428 ( .A(n44106), .B(n44107), .Z(n43888) );
  NANDN U44429 ( .A(n44108), .B(n44109), .Z(n44107) );
  OR U44430 ( .A(n44110), .B(n44111), .Z(n44109) );
  NAND U44431 ( .A(n44111), .B(n44110), .Z(n44106) );
  ANDN U44432 ( .B(B[115]), .A(n65), .Z(n43890) );
  XNOR U44433 ( .A(n43898), .B(n44112), .Z(n43891) );
  XNOR U44434 ( .A(n43897), .B(n43895), .Z(n44112) );
  AND U44435 ( .A(n44113), .B(n44114), .Z(n43895) );
  NANDN U44436 ( .A(n44115), .B(n44116), .Z(n44114) );
  NANDN U44437 ( .A(n44117), .B(n44118), .Z(n44116) );
  NANDN U44438 ( .A(n44118), .B(n44117), .Z(n44113) );
  ANDN U44439 ( .B(B[116]), .A(n66), .Z(n43897) );
  XNOR U44440 ( .A(n43905), .B(n44119), .Z(n43898) );
  XNOR U44441 ( .A(n43904), .B(n43902), .Z(n44119) );
  AND U44442 ( .A(n44120), .B(n44121), .Z(n43902) );
  NANDN U44443 ( .A(n44122), .B(n44123), .Z(n44121) );
  OR U44444 ( .A(n44124), .B(n44125), .Z(n44123) );
  NAND U44445 ( .A(n44125), .B(n44124), .Z(n44120) );
  ANDN U44446 ( .B(B[117]), .A(n67), .Z(n43904) );
  XNOR U44447 ( .A(n43912), .B(n44126), .Z(n43905) );
  XNOR U44448 ( .A(n43911), .B(n43909), .Z(n44126) );
  AND U44449 ( .A(n44127), .B(n44128), .Z(n43909) );
  NANDN U44450 ( .A(n44129), .B(n44130), .Z(n44128) );
  NANDN U44451 ( .A(n44131), .B(n44132), .Z(n44130) );
  NANDN U44452 ( .A(n44132), .B(n44131), .Z(n44127) );
  ANDN U44453 ( .B(B[118]), .A(n68), .Z(n43911) );
  XNOR U44454 ( .A(n43919), .B(n44133), .Z(n43912) );
  XNOR U44455 ( .A(n43918), .B(n43916), .Z(n44133) );
  AND U44456 ( .A(n44134), .B(n44135), .Z(n43916) );
  NANDN U44457 ( .A(n44136), .B(n44137), .Z(n44135) );
  OR U44458 ( .A(n44138), .B(n44139), .Z(n44137) );
  NAND U44459 ( .A(n44139), .B(n44138), .Z(n44134) );
  ANDN U44460 ( .B(B[119]), .A(n69), .Z(n43918) );
  XNOR U44461 ( .A(n43926), .B(n44140), .Z(n43919) );
  XNOR U44462 ( .A(n43925), .B(n43923), .Z(n44140) );
  AND U44463 ( .A(n44141), .B(n44142), .Z(n43923) );
  NANDN U44464 ( .A(n44143), .B(n44144), .Z(n44142) );
  NANDN U44465 ( .A(n44145), .B(n44146), .Z(n44144) );
  NANDN U44466 ( .A(n44146), .B(n44145), .Z(n44141) );
  ANDN U44467 ( .B(B[120]), .A(n70), .Z(n43925) );
  XNOR U44468 ( .A(n43933), .B(n44147), .Z(n43926) );
  XNOR U44469 ( .A(n43932), .B(n43930), .Z(n44147) );
  AND U44470 ( .A(n44148), .B(n44149), .Z(n43930) );
  NANDN U44471 ( .A(n44150), .B(n44151), .Z(n44149) );
  OR U44472 ( .A(n44152), .B(n44153), .Z(n44151) );
  NAND U44473 ( .A(n44153), .B(n44152), .Z(n44148) );
  ANDN U44474 ( .B(B[121]), .A(n71), .Z(n43932) );
  XNOR U44475 ( .A(n43940), .B(n44154), .Z(n43933) );
  XNOR U44476 ( .A(n43939), .B(n43937), .Z(n44154) );
  AND U44477 ( .A(n44155), .B(n44156), .Z(n43937) );
  NANDN U44478 ( .A(n44157), .B(n44158), .Z(n44156) );
  NANDN U44479 ( .A(n44159), .B(n44160), .Z(n44158) );
  NANDN U44480 ( .A(n44160), .B(n44159), .Z(n44155) );
  ANDN U44481 ( .B(B[122]), .A(n72), .Z(n43939) );
  XNOR U44482 ( .A(n43947), .B(n44161), .Z(n43940) );
  XNOR U44483 ( .A(n43946), .B(n43944), .Z(n44161) );
  AND U44484 ( .A(n44162), .B(n44163), .Z(n43944) );
  NANDN U44485 ( .A(n44164), .B(n44165), .Z(n44163) );
  OR U44486 ( .A(n44166), .B(n44167), .Z(n44165) );
  NAND U44487 ( .A(n44167), .B(n44166), .Z(n44162) );
  ANDN U44488 ( .B(B[123]), .A(n73), .Z(n43946) );
  XNOR U44489 ( .A(n43954), .B(n44168), .Z(n43947) );
  XNOR U44490 ( .A(n43953), .B(n43951), .Z(n44168) );
  AND U44491 ( .A(n44169), .B(n44170), .Z(n43951) );
  NANDN U44492 ( .A(n44171), .B(n44172), .Z(n44170) );
  NANDN U44493 ( .A(n44173), .B(n44174), .Z(n44172) );
  NANDN U44494 ( .A(n44174), .B(n44173), .Z(n44169) );
  ANDN U44495 ( .B(B[124]), .A(n74), .Z(n43953) );
  XNOR U44496 ( .A(n43961), .B(n44175), .Z(n43954) );
  XNOR U44497 ( .A(n43960), .B(n43958), .Z(n44175) );
  AND U44498 ( .A(n44176), .B(n44177), .Z(n43958) );
  NANDN U44499 ( .A(n44178), .B(n44179), .Z(n44177) );
  OR U44500 ( .A(n44180), .B(n44181), .Z(n44179) );
  NAND U44501 ( .A(n44181), .B(n44180), .Z(n44176) );
  ANDN U44502 ( .B(B[125]), .A(n75), .Z(n43960) );
  XNOR U44503 ( .A(n43968), .B(n44182), .Z(n43961) );
  XNOR U44504 ( .A(n43967), .B(n43965), .Z(n44182) );
  AND U44505 ( .A(n44183), .B(n44184), .Z(n43965) );
  NANDN U44506 ( .A(n44185), .B(n44186), .Z(n44184) );
  NANDN U44507 ( .A(n44187), .B(n44188), .Z(n44186) );
  NANDN U44508 ( .A(n44188), .B(n44187), .Z(n44183) );
  ANDN U44509 ( .B(B[126]), .A(n76), .Z(n43967) );
  XNOR U44510 ( .A(n43975), .B(n44189), .Z(n43968) );
  XNOR U44511 ( .A(n43974), .B(n43972), .Z(n44189) );
  AND U44512 ( .A(n44190), .B(n44191), .Z(n43972) );
  NANDN U44513 ( .A(n44192), .B(n44193), .Z(n44191) );
  OR U44514 ( .A(n44194), .B(n44195), .Z(n44193) );
  NAND U44515 ( .A(n44195), .B(n44194), .Z(n44190) );
  ANDN U44516 ( .B(B[127]), .A(n77), .Z(n43974) );
  XNOR U44517 ( .A(n43982), .B(n44196), .Z(n43975) );
  XNOR U44518 ( .A(n43981), .B(n43979), .Z(n44196) );
  AND U44519 ( .A(n44197), .B(n44198), .Z(n43979) );
  NANDN U44520 ( .A(n44199), .B(n44200), .Z(n44198) );
  NANDN U44521 ( .A(n44201), .B(n44202), .Z(n44200) );
  NANDN U44522 ( .A(n44202), .B(n44201), .Z(n44197) );
  ANDN U44523 ( .B(B[128]), .A(n78), .Z(n43981) );
  XNOR U44524 ( .A(n43989), .B(n44203), .Z(n43982) );
  XNOR U44525 ( .A(n43988), .B(n43986), .Z(n44203) );
  AND U44526 ( .A(n44204), .B(n44205), .Z(n43986) );
  NANDN U44527 ( .A(n44206), .B(n44207), .Z(n44205) );
  OR U44528 ( .A(n44208), .B(n44209), .Z(n44207) );
  NAND U44529 ( .A(n44209), .B(n44208), .Z(n44204) );
  ANDN U44530 ( .B(B[129]), .A(n79), .Z(n43988) );
  XNOR U44531 ( .A(n43996), .B(n44210), .Z(n43989) );
  XNOR U44532 ( .A(n43995), .B(n43993), .Z(n44210) );
  AND U44533 ( .A(n44211), .B(n44212), .Z(n43993) );
  NANDN U44534 ( .A(n44213), .B(n44214), .Z(n44212) );
  NANDN U44535 ( .A(n44215), .B(n44216), .Z(n44214) );
  NANDN U44536 ( .A(n44216), .B(n44215), .Z(n44211) );
  ANDN U44537 ( .B(B[130]), .A(n80), .Z(n43995) );
  XNOR U44538 ( .A(n44003), .B(n44217), .Z(n43996) );
  XNOR U44539 ( .A(n44002), .B(n44000), .Z(n44217) );
  AND U44540 ( .A(n44218), .B(n44219), .Z(n44000) );
  NANDN U44541 ( .A(n44220), .B(n44221), .Z(n44219) );
  OR U44542 ( .A(n44222), .B(n44223), .Z(n44221) );
  NAND U44543 ( .A(n44223), .B(n44222), .Z(n44218) );
  ANDN U44544 ( .B(B[131]), .A(n81), .Z(n44002) );
  XNOR U44545 ( .A(n44010), .B(n44224), .Z(n44003) );
  XNOR U44546 ( .A(n44009), .B(n44007), .Z(n44224) );
  AND U44547 ( .A(n44225), .B(n44226), .Z(n44007) );
  NANDN U44548 ( .A(n44227), .B(n44228), .Z(n44226) );
  NAND U44549 ( .A(n44229), .B(n44230), .Z(n44228) );
  ANDN U44550 ( .B(B[132]), .A(n82), .Z(n44009) );
  XOR U44551 ( .A(n44016), .B(n44231), .Z(n44010) );
  XNOR U44552 ( .A(n44014), .B(n44017), .Z(n44231) );
  NAND U44553 ( .A(A[2]), .B(B[133]), .Z(n44017) );
  NANDN U44554 ( .A(n44232), .B(n44233), .Z(n44014) );
  AND U44555 ( .A(A[0]), .B(B[134]), .Z(n44233) );
  XNOR U44556 ( .A(n44019), .B(n44234), .Z(n44016) );
  NAND U44557 ( .A(A[0]), .B(B[135]), .Z(n44234) );
  NAND U44558 ( .A(B[134]), .B(A[1]), .Z(n44019) );
  NAND U44559 ( .A(n44235), .B(n44236), .Z(n526) );
  NANDN U44560 ( .A(n44237), .B(n44238), .Z(n44236) );
  OR U44561 ( .A(n44239), .B(n44240), .Z(n44238) );
  NAND U44562 ( .A(n44240), .B(n44239), .Z(n44235) );
  XOR U44563 ( .A(n528), .B(n527), .Z(\A1[132] ) );
  XOR U44564 ( .A(n44240), .B(n44241), .Z(n527) );
  XNOR U44565 ( .A(n44239), .B(n44237), .Z(n44241) );
  AND U44566 ( .A(n44242), .B(n44243), .Z(n44237) );
  NANDN U44567 ( .A(n44244), .B(n44245), .Z(n44243) );
  NANDN U44568 ( .A(n44246), .B(n44247), .Z(n44245) );
  NANDN U44569 ( .A(n44247), .B(n44246), .Z(n44242) );
  ANDN U44570 ( .B(B[103]), .A(n54), .Z(n44239) );
  XNOR U44571 ( .A(n44034), .B(n44248), .Z(n44240) );
  XNOR U44572 ( .A(n44033), .B(n44031), .Z(n44248) );
  AND U44573 ( .A(n44249), .B(n44250), .Z(n44031) );
  NANDN U44574 ( .A(n44251), .B(n44252), .Z(n44250) );
  OR U44575 ( .A(n44253), .B(n44254), .Z(n44252) );
  NAND U44576 ( .A(n44254), .B(n44253), .Z(n44249) );
  ANDN U44577 ( .B(B[104]), .A(n55), .Z(n44033) );
  XNOR U44578 ( .A(n44041), .B(n44255), .Z(n44034) );
  XNOR U44579 ( .A(n44040), .B(n44038), .Z(n44255) );
  AND U44580 ( .A(n44256), .B(n44257), .Z(n44038) );
  NANDN U44581 ( .A(n44258), .B(n44259), .Z(n44257) );
  NANDN U44582 ( .A(n44260), .B(n44261), .Z(n44259) );
  NANDN U44583 ( .A(n44261), .B(n44260), .Z(n44256) );
  ANDN U44584 ( .B(B[105]), .A(n56), .Z(n44040) );
  XNOR U44585 ( .A(n44048), .B(n44262), .Z(n44041) );
  XNOR U44586 ( .A(n44047), .B(n44045), .Z(n44262) );
  AND U44587 ( .A(n44263), .B(n44264), .Z(n44045) );
  NANDN U44588 ( .A(n44265), .B(n44266), .Z(n44264) );
  OR U44589 ( .A(n44267), .B(n44268), .Z(n44266) );
  NAND U44590 ( .A(n44268), .B(n44267), .Z(n44263) );
  ANDN U44591 ( .B(B[106]), .A(n57), .Z(n44047) );
  XNOR U44592 ( .A(n44055), .B(n44269), .Z(n44048) );
  XNOR U44593 ( .A(n44054), .B(n44052), .Z(n44269) );
  AND U44594 ( .A(n44270), .B(n44271), .Z(n44052) );
  NANDN U44595 ( .A(n44272), .B(n44273), .Z(n44271) );
  NANDN U44596 ( .A(n44274), .B(n44275), .Z(n44273) );
  NANDN U44597 ( .A(n44275), .B(n44274), .Z(n44270) );
  ANDN U44598 ( .B(B[107]), .A(n58), .Z(n44054) );
  XNOR U44599 ( .A(n44062), .B(n44276), .Z(n44055) );
  XNOR U44600 ( .A(n44061), .B(n44059), .Z(n44276) );
  AND U44601 ( .A(n44277), .B(n44278), .Z(n44059) );
  NANDN U44602 ( .A(n44279), .B(n44280), .Z(n44278) );
  OR U44603 ( .A(n44281), .B(n44282), .Z(n44280) );
  NAND U44604 ( .A(n44282), .B(n44281), .Z(n44277) );
  ANDN U44605 ( .B(B[108]), .A(n59), .Z(n44061) );
  XNOR U44606 ( .A(n44069), .B(n44283), .Z(n44062) );
  XNOR U44607 ( .A(n44068), .B(n44066), .Z(n44283) );
  AND U44608 ( .A(n44284), .B(n44285), .Z(n44066) );
  NANDN U44609 ( .A(n44286), .B(n44287), .Z(n44285) );
  NANDN U44610 ( .A(n44288), .B(n44289), .Z(n44287) );
  NANDN U44611 ( .A(n44289), .B(n44288), .Z(n44284) );
  ANDN U44612 ( .B(B[109]), .A(n60), .Z(n44068) );
  XNOR U44613 ( .A(n44076), .B(n44290), .Z(n44069) );
  XNOR U44614 ( .A(n44075), .B(n44073), .Z(n44290) );
  AND U44615 ( .A(n44291), .B(n44292), .Z(n44073) );
  NANDN U44616 ( .A(n44293), .B(n44294), .Z(n44292) );
  OR U44617 ( .A(n44295), .B(n44296), .Z(n44294) );
  NAND U44618 ( .A(n44296), .B(n44295), .Z(n44291) );
  ANDN U44619 ( .B(B[110]), .A(n61), .Z(n44075) );
  XNOR U44620 ( .A(n44083), .B(n44297), .Z(n44076) );
  XNOR U44621 ( .A(n44082), .B(n44080), .Z(n44297) );
  AND U44622 ( .A(n44298), .B(n44299), .Z(n44080) );
  NANDN U44623 ( .A(n44300), .B(n44301), .Z(n44299) );
  NANDN U44624 ( .A(n44302), .B(n44303), .Z(n44301) );
  NANDN U44625 ( .A(n44303), .B(n44302), .Z(n44298) );
  ANDN U44626 ( .B(B[111]), .A(n62), .Z(n44082) );
  XNOR U44627 ( .A(n44090), .B(n44304), .Z(n44083) );
  XNOR U44628 ( .A(n44089), .B(n44087), .Z(n44304) );
  AND U44629 ( .A(n44305), .B(n44306), .Z(n44087) );
  NANDN U44630 ( .A(n44307), .B(n44308), .Z(n44306) );
  OR U44631 ( .A(n44309), .B(n44310), .Z(n44308) );
  NAND U44632 ( .A(n44310), .B(n44309), .Z(n44305) );
  ANDN U44633 ( .B(B[112]), .A(n63), .Z(n44089) );
  XNOR U44634 ( .A(n44097), .B(n44311), .Z(n44090) );
  XNOR U44635 ( .A(n44096), .B(n44094), .Z(n44311) );
  AND U44636 ( .A(n44312), .B(n44313), .Z(n44094) );
  NANDN U44637 ( .A(n44314), .B(n44315), .Z(n44313) );
  NANDN U44638 ( .A(n44316), .B(n44317), .Z(n44315) );
  NANDN U44639 ( .A(n44317), .B(n44316), .Z(n44312) );
  ANDN U44640 ( .B(B[113]), .A(n64), .Z(n44096) );
  XNOR U44641 ( .A(n44104), .B(n44318), .Z(n44097) );
  XNOR U44642 ( .A(n44103), .B(n44101), .Z(n44318) );
  AND U44643 ( .A(n44319), .B(n44320), .Z(n44101) );
  NANDN U44644 ( .A(n44321), .B(n44322), .Z(n44320) );
  OR U44645 ( .A(n44323), .B(n44324), .Z(n44322) );
  NAND U44646 ( .A(n44324), .B(n44323), .Z(n44319) );
  ANDN U44647 ( .B(B[114]), .A(n65), .Z(n44103) );
  XNOR U44648 ( .A(n44111), .B(n44325), .Z(n44104) );
  XNOR U44649 ( .A(n44110), .B(n44108), .Z(n44325) );
  AND U44650 ( .A(n44326), .B(n44327), .Z(n44108) );
  NANDN U44651 ( .A(n44328), .B(n44329), .Z(n44327) );
  NANDN U44652 ( .A(n44330), .B(n44331), .Z(n44329) );
  NANDN U44653 ( .A(n44331), .B(n44330), .Z(n44326) );
  ANDN U44654 ( .B(B[115]), .A(n66), .Z(n44110) );
  XNOR U44655 ( .A(n44118), .B(n44332), .Z(n44111) );
  XNOR U44656 ( .A(n44117), .B(n44115), .Z(n44332) );
  AND U44657 ( .A(n44333), .B(n44334), .Z(n44115) );
  NANDN U44658 ( .A(n44335), .B(n44336), .Z(n44334) );
  OR U44659 ( .A(n44337), .B(n44338), .Z(n44336) );
  NAND U44660 ( .A(n44338), .B(n44337), .Z(n44333) );
  ANDN U44661 ( .B(B[116]), .A(n67), .Z(n44117) );
  XNOR U44662 ( .A(n44125), .B(n44339), .Z(n44118) );
  XNOR U44663 ( .A(n44124), .B(n44122), .Z(n44339) );
  AND U44664 ( .A(n44340), .B(n44341), .Z(n44122) );
  NANDN U44665 ( .A(n44342), .B(n44343), .Z(n44341) );
  NANDN U44666 ( .A(n44344), .B(n44345), .Z(n44343) );
  NANDN U44667 ( .A(n44345), .B(n44344), .Z(n44340) );
  ANDN U44668 ( .B(B[117]), .A(n68), .Z(n44124) );
  XNOR U44669 ( .A(n44132), .B(n44346), .Z(n44125) );
  XNOR U44670 ( .A(n44131), .B(n44129), .Z(n44346) );
  AND U44671 ( .A(n44347), .B(n44348), .Z(n44129) );
  NANDN U44672 ( .A(n44349), .B(n44350), .Z(n44348) );
  OR U44673 ( .A(n44351), .B(n44352), .Z(n44350) );
  NAND U44674 ( .A(n44352), .B(n44351), .Z(n44347) );
  ANDN U44675 ( .B(B[118]), .A(n69), .Z(n44131) );
  XNOR U44676 ( .A(n44139), .B(n44353), .Z(n44132) );
  XNOR U44677 ( .A(n44138), .B(n44136), .Z(n44353) );
  AND U44678 ( .A(n44354), .B(n44355), .Z(n44136) );
  NANDN U44679 ( .A(n44356), .B(n44357), .Z(n44355) );
  NANDN U44680 ( .A(n44358), .B(n44359), .Z(n44357) );
  NANDN U44681 ( .A(n44359), .B(n44358), .Z(n44354) );
  ANDN U44682 ( .B(B[119]), .A(n70), .Z(n44138) );
  XNOR U44683 ( .A(n44146), .B(n44360), .Z(n44139) );
  XNOR U44684 ( .A(n44145), .B(n44143), .Z(n44360) );
  AND U44685 ( .A(n44361), .B(n44362), .Z(n44143) );
  NANDN U44686 ( .A(n44363), .B(n44364), .Z(n44362) );
  OR U44687 ( .A(n44365), .B(n44366), .Z(n44364) );
  NAND U44688 ( .A(n44366), .B(n44365), .Z(n44361) );
  ANDN U44689 ( .B(B[120]), .A(n71), .Z(n44145) );
  XNOR U44690 ( .A(n44153), .B(n44367), .Z(n44146) );
  XNOR U44691 ( .A(n44152), .B(n44150), .Z(n44367) );
  AND U44692 ( .A(n44368), .B(n44369), .Z(n44150) );
  NANDN U44693 ( .A(n44370), .B(n44371), .Z(n44369) );
  NANDN U44694 ( .A(n44372), .B(n44373), .Z(n44371) );
  NANDN U44695 ( .A(n44373), .B(n44372), .Z(n44368) );
  ANDN U44696 ( .B(B[121]), .A(n72), .Z(n44152) );
  XNOR U44697 ( .A(n44160), .B(n44374), .Z(n44153) );
  XNOR U44698 ( .A(n44159), .B(n44157), .Z(n44374) );
  AND U44699 ( .A(n44375), .B(n44376), .Z(n44157) );
  NANDN U44700 ( .A(n44377), .B(n44378), .Z(n44376) );
  OR U44701 ( .A(n44379), .B(n44380), .Z(n44378) );
  NAND U44702 ( .A(n44380), .B(n44379), .Z(n44375) );
  ANDN U44703 ( .B(B[122]), .A(n73), .Z(n44159) );
  XNOR U44704 ( .A(n44167), .B(n44381), .Z(n44160) );
  XNOR U44705 ( .A(n44166), .B(n44164), .Z(n44381) );
  AND U44706 ( .A(n44382), .B(n44383), .Z(n44164) );
  NANDN U44707 ( .A(n44384), .B(n44385), .Z(n44383) );
  NANDN U44708 ( .A(n44386), .B(n44387), .Z(n44385) );
  NANDN U44709 ( .A(n44387), .B(n44386), .Z(n44382) );
  ANDN U44710 ( .B(B[123]), .A(n74), .Z(n44166) );
  XNOR U44711 ( .A(n44174), .B(n44388), .Z(n44167) );
  XNOR U44712 ( .A(n44173), .B(n44171), .Z(n44388) );
  AND U44713 ( .A(n44389), .B(n44390), .Z(n44171) );
  NANDN U44714 ( .A(n44391), .B(n44392), .Z(n44390) );
  OR U44715 ( .A(n44393), .B(n44394), .Z(n44392) );
  NAND U44716 ( .A(n44394), .B(n44393), .Z(n44389) );
  ANDN U44717 ( .B(B[124]), .A(n75), .Z(n44173) );
  XNOR U44718 ( .A(n44181), .B(n44395), .Z(n44174) );
  XNOR U44719 ( .A(n44180), .B(n44178), .Z(n44395) );
  AND U44720 ( .A(n44396), .B(n44397), .Z(n44178) );
  NANDN U44721 ( .A(n44398), .B(n44399), .Z(n44397) );
  NANDN U44722 ( .A(n44400), .B(n44401), .Z(n44399) );
  NANDN U44723 ( .A(n44401), .B(n44400), .Z(n44396) );
  ANDN U44724 ( .B(B[125]), .A(n76), .Z(n44180) );
  XNOR U44725 ( .A(n44188), .B(n44402), .Z(n44181) );
  XNOR U44726 ( .A(n44187), .B(n44185), .Z(n44402) );
  AND U44727 ( .A(n44403), .B(n44404), .Z(n44185) );
  NANDN U44728 ( .A(n44405), .B(n44406), .Z(n44404) );
  OR U44729 ( .A(n44407), .B(n44408), .Z(n44406) );
  NAND U44730 ( .A(n44408), .B(n44407), .Z(n44403) );
  ANDN U44731 ( .B(B[126]), .A(n77), .Z(n44187) );
  XNOR U44732 ( .A(n44195), .B(n44409), .Z(n44188) );
  XNOR U44733 ( .A(n44194), .B(n44192), .Z(n44409) );
  AND U44734 ( .A(n44410), .B(n44411), .Z(n44192) );
  NANDN U44735 ( .A(n44412), .B(n44413), .Z(n44411) );
  NANDN U44736 ( .A(n44414), .B(n44415), .Z(n44413) );
  NANDN U44737 ( .A(n44415), .B(n44414), .Z(n44410) );
  ANDN U44738 ( .B(B[127]), .A(n78), .Z(n44194) );
  XNOR U44739 ( .A(n44202), .B(n44416), .Z(n44195) );
  XNOR U44740 ( .A(n44201), .B(n44199), .Z(n44416) );
  AND U44741 ( .A(n44417), .B(n44418), .Z(n44199) );
  NANDN U44742 ( .A(n44419), .B(n44420), .Z(n44418) );
  OR U44743 ( .A(n44421), .B(n44422), .Z(n44420) );
  NAND U44744 ( .A(n44422), .B(n44421), .Z(n44417) );
  ANDN U44745 ( .B(B[128]), .A(n79), .Z(n44201) );
  XNOR U44746 ( .A(n44209), .B(n44423), .Z(n44202) );
  XNOR U44747 ( .A(n44208), .B(n44206), .Z(n44423) );
  AND U44748 ( .A(n44424), .B(n44425), .Z(n44206) );
  NANDN U44749 ( .A(n44426), .B(n44427), .Z(n44425) );
  NANDN U44750 ( .A(n44428), .B(n44429), .Z(n44427) );
  NANDN U44751 ( .A(n44429), .B(n44428), .Z(n44424) );
  ANDN U44752 ( .B(B[129]), .A(n80), .Z(n44208) );
  XNOR U44753 ( .A(n44216), .B(n44430), .Z(n44209) );
  XNOR U44754 ( .A(n44215), .B(n44213), .Z(n44430) );
  AND U44755 ( .A(n44431), .B(n44432), .Z(n44213) );
  NANDN U44756 ( .A(n44433), .B(n44434), .Z(n44432) );
  OR U44757 ( .A(n44435), .B(n44436), .Z(n44434) );
  NAND U44758 ( .A(n44436), .B(n44435), .Z(n44431) );
  ANDN U44759 ( .B(B[130]), .A(n81), .Z(n44215) );
  XNOR U44760 ( .A(n44223), .B(n44437), .Z(n44216) );
  XNOR U44761 ( .A(n44222), .B(n44220), .Z(n44437) );
  AND U44762 ( .A(n44438), .B(n44439), .Z(n44220) );
  NANDN U44763 ( .A(n44440), .B(n44441), .Z(n44439) );
  NAND U44764 ( .A(n44442), .B(n44443), .Z(n44441) );
  ANDN U44765 ( .B(B[131]), .A(n82), .Z(n44222) );
  XOR U44766 ( .A(n44229), .B(n44444), .Z(n44223) );
  XNOR U44767 ( .A(n44227), .B(n44230), .Z(n44444) );
  NAND U44768 ( .A(A[2]), .B(B[132]), .Z(n44230) );
  NANDN U44769 ( .A(n44445), .B(n44446), .Z(n44227) );
  AND U44770 ( .A(A[0]), .B(B[133]), .Z(n44446) );
  XNOR U44771 ( .A(n44232), .B(n44447), .Z(n44229) );
  NAND U44772 ( .A(A[0]), .B(B[134]), .Z(n44447) );
  NAND U44773 ( .A(B[133]), .B(A[1]), .Z(n44232) );
  NAND U44774 ( .A(n44448), .B(n44449), .Z(n528) );
  NANDN U44775 ( .A(n44450), .B(n44451), .Z(n44449) );
  OR U44776 ( .A(n44452), .B(n44453), .Z(n44451) );
  NAND U44777 ( .A(n44453), .B(n44452), .Z(n44448) );
  XOR U44778 ( .A(n530), .B(n529), .Z(\A1[131] ) );
  XOR U44779 ( .A(n44453), .B(n44454), .Z(n529) );
  XNOR U44780 ( .A(n44452), .B(n44450), .Z(n44454) );
  AND U44781 ( .A(n44455), .B(n44456), .Z(n44450) );
  NANDN U44782 ( .A(n44457), .B(n44458), .Z(n44456) );
  NANDN U44783 ( .A(n44459), .B(n44460), .Z(n44458) );
  NANDN U44784 ( .A(n44460), .B(n44459), .Z(n44455) );
  ANDN U44785 ( .B(B[102]), .A(n54), .Z(n44452) );
  XNOR U44786 ( .A(n44247), .B(n44461), .Z(n44453) );
  XNOR U44787 ( .A(n44246), .B(n44244), .Z(n44461) );
  AND U44788 ( .A(n44462), .B(n44463), .Z(n44244) );
  NANDN U44789 ( .A(n44464), .B(n44465), .Z(n44463) );
  OR U44790 ( .A(n44466), .B(n44467), .Z(n44465) );
  NAND U44791 ( .A(n44467), .B(n44466), .Z(n44462) );
  ANDN U44792 ( .B(B[103]), .A(n55), .Z(n44246) );
  XNOR U44793 ( .A(n44254), .B(n44468), .Z(n44247) );
  XNOR U44794 ( .A(n44253), .B(n44251), .Z(n44468) );
  AND U44795 ( .A(n44469), .B(n44470), .Z(n44251) );
  NANDN U44796 ( .A(n44471), .B(n44472), .Z(n44470) );
  NANDN U44797 ( .A(n44473), .B(n44474), .Z(n44472) );
  NANDN U44798 ( .A(n44474), .B(n44473), .Z(n44469) );
  ANDN U44799 ( .B(B[104]), .A(n56), .Z(n44253) );
  XNOR U44800 ( .A(n44261), .B(n44475), .Z(n44254) );
  XNOR U44801 ( .A(n44260), .B(n44258), .Z(n44475) );
  AND U44802 ( .A(n44476), .B(n44477), .Z(n44258) );
  NANDN U44803 ( .A(n44478), .B(n44479), .Z(n44477) );
  OR U44804 ( .A(n44480), .B(n44481), .Z(n44479) );
  NAND U44805 ( .A(n44481), .B(n44480), .Z(n44476) );
  ANDN U44806 ( .B(B[105]), .A(n57), .Z(n44260) );
  XNOR U44807 ( .A(n44268), .B(n44482), .Z(n44261) );
  XNOR U44808 ( .A(n44267), .B(n44265), .Z(n44482) );
  AND U44809 ( .A(n44483), .B(n44484), .Z(n44265) );
  NANDN U44810 ( .A(n44485), .B(n44486), .Z(n44484) );
  NANDN U44811 ( .A(n44487), .B(n44488), .Z(n44486) );
  NANDN U44812 ( .A(n44488), .B(n44487), .Z(n44483) );
  ANDN U44813 ( .B(B[106]), .A(n58), .Z(n44267) );
  XNOR U44814 ( .A(n44275), .B(n44489), .Z(n44268) );
  XNOR U44815 ( .A(n44274), .B(n44272), .Z(n44489) );
  AND U44816 ( .A(n44490), .B(n44491), .Z(n44272) );
  NANDN U44817 ( .A(n44492), .B(n44493), .Z(n44491) );
  OR U44818 ( .A(n44494), .B(n44495), .Z(n44493) );
  NAND U44819 ( .A(n44495), .B(n44494), .Z(n44490) );
  ANDN U44820 ( .B(B[107]), .A(n59), .Z(n44274) );
  XNOR U44821 ( .A(n44282), .B(n44496), .Z(n44275) );
  XNOR U44822 ( .A(n44281), .B(n44279), .Z(n44496) );
  AND U44823 ( .A(n44497), .B(n44498), .Z(n44279) );
  NANDN U44824 ( .A(n44499), .B(n44500), .Z(n44498) );
  NANDN U44825 ( .A(n44501), .B(n44502), .Z(n44500) );
  NANDN U44826 ( .A(n44502), .B(n44501), .Z(n44497) );
  ANDN U44827 ( .B(B[108]), .A(n60), .Z(n44281) );
  XNOR U44828 ( .A(n44289), .B(n44503), .Z(n44282) );
  XNOR U44829 ( .A(n44288), .B(n44286), .Z(n44503) );
  AND U44830 ( .A(n44504), .B(n44505), .Z(n44286) );
  NANDN U44831 ( .A(n44506), .B(n44507), .Z(n44505) );
  OR U44832 ( .A(n44508), .B(n44509), .Z(n44507) );
  NAND U44833 ( .A(n44509), .B(n44508), .Z(n44504) );
  ANDN U44834 ( .B(B[109]), .A(n61), .Z(n44288) );
  XNOR U44835 ( .A(n44296), .B(n44510), .Z(n44289) );
  XNOR U44836 ( .A(n44295), .B(n44293), .Z(n44510) );
  AND U44837 ( .A(n44511), .B(n44512), .Z(n44293) );
  NANDN U44838 ( .A(n44513), .B(n44514), .Z(n44512) );
  NANDN U44839 ( .A(n44515), .B(n44516), .Z(n44514) );
  NANDN U44840 ( .A(n44516), .B(n44515), .Z(n44511) );
  ANDN U44841 ( .B(B[110]), .A(n62), .Z(n44295) );
  XNOR U44842 ( .A(n44303), .B(n44517), .Z(n44296) );
  XNOR U44843 ( .A(n44302), .B(n44300), .Z(n44517) );
  AND U44844 ( .A(n44518), .B(n44519), .Z(n44300) );
  NANDN U44845 ( .A(n44520), .B(n44521), .Z(n44519) );
  OR U44846 ( .A(n44522), .B(n44523), .Z(n44521) );
  NAND U44847 ( .A(n44523), .B(n44522), .Z(n44518) );
  ANDN U44848 ( .B(B[111]), .A(n63), .Z(n44302) );
  XNOR U44849 ( .A(n44310), .B(n44524), .Z(n44303) );
  XNOR U44850 ( .A(n44309), .B(n44307), .Z(n44524) );
  AND U44851 ( .A(n44525), .B(n44526), .Z(n44307) );
  NANDN U44852 ( .A(n44527), .B(n44528), .Z(n44526) );
  NANDN U44853 ( .A(n44529), .B(n44530), .Z(n44528) );
  NANDN U44854 ( .A(n44530), .B(n44529), .Z(n44525) );
  ANDN U44855 ( .B(B[112]), .A(n64), .Z(n44309) );
  XNOR U44856 ( .A(n44317), .B(n44531), .Z(n44310) );
  XNOR U44857 ( .A(n44316), .B(n44314), .Z(n44531) );
  AND U44858 ( .A(n44532), .B(n44533), .Z(n44314) );
  NANDN U44859 ( .A(n44534), .B(n44535), .Z(n44533) );
  OR U44860 ( .A(n44536), .B(n44537), .Z(n44535) );
  NAND U44861 ( .A(n44537), .B(n44536), .Z(n44532) );
  ANDN U44862 ( .B(B[113]), .A(n65), .Z(n44316) );
  XNOR U44863 ( .A(n44324), .B(n44538), .Z(n44317) );
  XNOR U44864 ( .A(n44323), .B(n44321), .Z(n44538) );
  AND U44865 ( .A(n44539), .B(n44540), .Z(n44321) );
  NANDN U44866 ( .A(n44541), .B(n44542), .Z(n44540) );
  NANDN U44867 ( .A(n44543), .B(n44544), .Z(n44542) );
  NANDN U44868 ( .A(n44544), .B(n44543), .Z(n44539) );
  ANDN U44869 ( .B(B[114]), .A(n66), .Z(n44323) );
  XNOR U44870 ( .A(n44331), .B(n44545), .Z(n44324) );
  XNOR U44871 ( .A(n44330), .B(n44328), .Z(n44545) );
  AND U44872 ( .A(n44546), .B(n44547), .Z(n44328) );
  NANDN U44873 ( .A(n44548), .B(n44549), .Z(n44547) );
  OR U44874 ( .A(n44550), .B(n44551), .Z(n44549) );
  NAND U44875 ( .A(n44551), .B(n44550), .Z(n44546) );
  ANDN U44876 ( .B(B[115]), .A(n67), .Z(n44330) );
  XNOR U44877 ( .A(n44338), .B(n44552), .Z(n44331) );
  XNOR U44878 ( .A(n44337), .B(n44335), .Z(n44552) );
  AND U44879 ( .A(n44553), .B(n44554), .Z(n44335) );
  NANDN U44880 ( .A(n44555), .B(n44556), .Z(n44554) );
  NANDN U44881 ( .A(n44557), .B(n44558), .Z(n44556) );
  NANDN U44882 ( .A(n44558), .B(n44557), .Z(n44553) );
  ANDN U44883 ( .B(B[116]), .A(n68), .Z(n44337) );
  XNOR U44884 ( .A(n44345), .B(n44559), .Z(n44338) );
  XNOR U44885 ( .A(n44344), .B(n44342), .Z(n44559) );
  AND U44886 ( .A(n44560), .B(n44561), .Z(n44342) );
  NANDN U44887 ( .A(n44562), .B(n44563), .Z(n44561) );
  OR U44888 ( .A(n44564), .B(n44565), .Z(n44563) );
  NAND U44889 ( .A(n44565), .B(n44564), .Z(n44560) );
  ANDN U44890 ( .B(B[117]), .A(n69), .Z(n44344) );
  XNOR U44891 ( .A(n44352), .B(n44566), .Z(n44345) );
  XNOR U44892 ( .A(n44351), .B(n44349), .Z(n44566) );
  AND U44893 ( .A(n44567), .B(n44568), .Z(n44349) );
  NANDN U44894 ( .A(n44569), .B(n44570), .Z(n44568) );
  NANDN U44895 ( .A(n44571), .B(n44572), .Z(n44570) );
  NANDN U44896 ( .A(n44572), .B(n44571), .Z(n44567) );
  ANDN U44897 ( .B(B[118]), .A(n70), .Z(n44351) );
  XNOR U44898 ( .A(n44359), .B(n44573), .Z(n44352) );
  XNOR U44899 ( .A(n44358), .B(n44356), .Z(n44573) );
  AND U44900 ( .A(n44574), .B(n44575), .Z(n44356) );
  NANDN U44901 ( .A(n44576), .B(n44577), .Z(n44575) );
  OR U44902 ( .A(n44578), .B(n44579), .Z(n44577) );
  NAND U44903 ( .A(n44579), .B(n44578), .Z(n44574) );
  ANDN U44904 ( .B(B[119]), .A(n71), .Z(n44358) );
  XNOR U44905 ( .A(n44366), .B(n44580), .Z(n44359) );
  XNOR U44906 ( .A(n44365), .B(n44363), .Z(n44580) );
  AND U44907 ( .A(n44581), .B(n44582), .Z(n44363) );
  NANDN U44908 ( .A(n44583), .B(n44584), .Z(n44582) );
  NANDN U44909 ( .A(n44585), .B(n44586), .Z(n44584) );
  NANDN U44910 ( .A(n44586), .B(n44585), .Z(n44581) );
  ANDN U44911 ( .B(B[120]), .A(n72), .Z(n44365) );
  XNOR U44912 ( .A(n44373), .B(n44587), .Z(n44366) );
  XNOR U44913 ( .A(n44372), .B(n44370), .Z(n44587) );
  AND U44914 ( .A(n44588), .B(n44589), .Z(n44370) );
  NANDN U44915 ( .A(n44590), .B(n44591), .Z(n44589) );
  OR U44916 ( .A(n44592), .B(n44593), .Z(n44591) );
  NAND U44917 ( .A(n44593), .B(n44592), .Z(n44588) );
  ANDN U44918 ( .B(B[121]), .A(n73), .Z(n44372) );
  XNOR U44919 ( .A(n44380), .B(n44594), .Z(n44373) );
  XNOR U44920 ( .A(n44379), .B(n44377), .Z(n44594) );
  AND U44921 ( .A(n44595), .B(n44596), .Z(n44377) );
  NANDN U44922 ( .A(n44597), .B(n44598), .Z(n44596) );
  NANDN U44923 ( .A(n44599), .B(n44600), .Z(n44598) );
  NANDN U44924 ( .A(n44600), .B(n44599), .Z(n44595) );
  ANDN U44925 ( .B(B[122]), .A(n74), .Z(n44379) );
  XNOR U44926 ( .A(n44387), .B(n44601), .Z(n44380) );
  XNOR U44927 ( .A(n44386), .B(n44384), .Z(n44601) );
  AND U44928 ( .A(n44602), .B(n44603), .Z(n44384) );
  NANDN U44929 ( .A(n44604), .B(n44605), .Z(n44603) );
  OR U44930 ( .A(n44606), .B(n44607), .Z(n44605) );
  NAND U44931 ( .A(n44607), .B(n44606), .Z(n44602) );
  ANDN U44932 ( .B(B[123]), .A(n75), .Z(n44386) );
  XNOR U44933 ( .A(n44394), .B(n44608), .Z(n44387) );
  XNOR U44934 ( .A(n44393), .B(n44391), .Z(n44608) );
  AND U44935 ( .A(n44609), .B(n44610), .Z(n44391) );
  NANDN U44936 ( .A(n44611), .B(n44612), .Z(n44610) );
  NANDN U44937 ( .A(n44613), .B(n44614), .Z(n44612) );
  NANDN U44938 ( .A(n44614), .B(n44613), .Z(n44609) );
  ANDN U44939 ( .B(B[124]), .A(n76), .Z(n44393) );
  XNOR U44940 ( .A(n44401), .B(n44615), .Z(n44394) );
  XNOR U44941 ( .A(n44400), .B(n44398), .Z(n44615) );
  AND U44942 ( .A(n44616), .B(n44617), .Z(n44398) );
  NANDN U44943 ( .A(n44618), .B(n44619), .Z(n44617) );
  OR U44944 ( .A(n44620), .B(n44621), .Z(n44619) );
  NAND U44945 ( .A(n44621), .B(n44620), .Z(n44616) );
  ANDN U44946 ( .B(B[125]), .A(n77), .Z(n44400) );
  XNOR U44947 ( .A(n44408), .B(n44622), .Z(n44401) );
  XNOR U44948 ( .A(n44407), .B(n44405), .Z(n44622) );
  AND U44949 ( .A(n44623), .B(n44624), .Z(n44405) );
  NANDN U44950 ( .A(n44625), .B(n44626), .Z(n44624) );
  NANDN U44951 ( .A(n44627), .B(n44628), .Z(n44626) );
  NANDN U44952 ( .A(n44628), .B(n44627), .Z(n44623) );
  ANDN U44953 ( .B(B[126]), .A(n78), .Z(n44407) );
  XNOR U44954 ( .A(n44415), .B(n44629), .Z(n44408) );
  XNOR U44955 ( .A(n44414), .B(n44412), .Z(n44629) );
  AND U44956 ( .A(n44630), .B(n44631), .Z(n44412) );
  NANDN U44957 ( .A(n44632), .B(n44633), .Z(n44631) );
  OR U44958 ( .A(n44634), .B(n44635), .Z(n44633) );
  NAND U44959 ( .A(n44635), .B(n44634), .Z(n44630) );
  ANDN U44960 ( .B(B[127]), .A(n79), .Z(n44414) );
  XNOR U44961 ( .A(n44422), .B(n44636), .Z(n44415) );
  XNOR U44962 ( .A(n44421), .B(n44419), .Z(n44636) );
  AND U44963 ( .A(n44637), .B(n44638), .Z(n44419) );
  NANDN U44964 ( .A(n44639), .B(n44640), .Z(n44638) );
  NANDN U44965 ( .A(n44641), .B(n44642), .Z(n44640) );
  NANDN U44966 ( .A(n44642), .B(n44641), .Z(n44637) );
  ANDN U44967 ( .B(B[128]), .A(n80), .Z(n44421) );
  XNOR U44968 ( .A(n44429), .B(n44643), .Z(n44422) );
  XNOR U44969 ( .A(n44428), .B(n44426), .Z(n44643) );
  AND U44970 ( .A(n44644), .B(n44645), .Z(n44426) );
  NANDN U44971 ( .A(n44646), .B(n44647), .Z(n44645) );
  OR U44972 ( .A(n44648), .B(n44649), .Z(n44647) );
  NAND U44973 ( .A(n44649), .B(n44648), .Z(n44644) );
  ANDN U44974 ( .B(B[129]), .A(n81), .Z(n44428) );
  XNOR U44975 ( .A(n44436), .B(n44650), .Z(n44429) );
  XNOR U44976 ( .A(n44435), .B(n44433), .Z(n44650) );
  AND U44977 ( .A(n44651), .B(n44652), .Z(n44433) );
  NANDN U44978 ( .A(n44653), .B(n44654), .Z(n44652) );
  NAND U44979 ( .A(n44655), .B(n44656), .Z(n44654) );
  ANDN U44980 ( .B(B[130]), .A(n82), .Z(n44435) );
  XOR U44981 ( .A(n44442), .B(n44657), .Z(n44436) );
  XNOR U44982 ( .A(n44440), .B(n44443), .Z(n44657) );
  NAND U44983 ( .A(A[2]), .B(B[131]), .Z(n44443) );
  NANDN U44984 ( .A(n44658), .B(n44659), .Z(n44440) );
  AND U44985 ( .A(A[0]), .B(B[132]), .Z(n44659) );
  XNOR U44986 ( .A(n44445), .B(n44660), .Z(n44442) );
  NAND U44987 ( .A(A[0]), .B(B[133]), .Z(n44660) );
  NAND U44988 ( .A(B[132]), .B(A[1]), .Z(n44445) );
  NAND U44989 ( .A(n44661), .B(n44662), .Z(n530) );
  NANDN U44990 ( .A(n44663), .B(n44664), .Z(n44662) );
  OR U44991 ( .A(n44665), .B(n44666), .Z(n44664) );
  NAND U44992 ( .A(n44666), .B(n44665), .Z(n44661) );
  XOR U44993 ( .A(n532), .B(n531), .Z(\A1[130] ) );
  XOR U44994 ( .A(n44666), .B(n44667), .Z(n531) );
  XNOR U44995 ( .A(n44665), .B(n44663), .Z(n44667) );
  AND U44996 ( .A(n44668), .B(n44669), .Z(n44663) );
  NANDN U44997 ( .A(n44670), .B(n44671), .Z(n44669) );
  NANDN U44998 ( .A(n44672), .B(n44673), .Z(n44671) );
  NANDN U44999 ( .A(n44673), .B(n44672), .Z(n44668) );
  ANDN U45000 ( .B(B[101]), .A(n54), .Z(n44665) );
  XNOR U45001 ( .A(n44460), .B(n44674), .Z(n44666) );
  XNOR U45002 ( .A(n44459), .B(n44457), .Z(n44674) );
  AND U45003 ( .A(n44675), .B(n44676), .Z(n44457) );
  NANDN U45004 ( .A(n44677), .B(n44678), .Z(n44676) );
  OR U45005 ( .A(n44679), .B(n44680), .Z(n44678) );
  NAND U45006 ( .A(n44680), .B(n44679), .Z(n44675) );
  ANDN U45007 ( .B(B[102]), .A(n55), .Z(n44459) );
  XNOR U45008 ( .A(n44467), .B(n44681), .Z(n44460) );
  XNOR U45009 ( .A(n44466), .B(n44464), .Z(n44681) );
  AND U45010 ( .A(n44682), .B(n44683), .Z(n44464) );
  NANDN U45011 ( .A(n44684), .B(n44685), .Z(n44683) );
  NANDN U45012 ( .A(n44686), .B(n44687), .Z(n44685) );
  NANDN U45013 ( .A(n44687), .B(n44686), .Z(n44682) );
  ANDN U45014 ( .B(B[103]), .A(n56), .Z(n44466) );
  XNOR U45015 ( .A(n44474), .B(n44688), .Z(n44467) );
  XNOR U45016 ( .A(n44473), .B(n44471), .Z(n44688) );
  AND U45017 ( .A(n44689), .B(n44690), .Z(n44471) );
  NANDN U45018 ( .A(n44691), .B(n44692), .Z(n44690) );
  OR U45019 ( .A(n44693), .B(n44694), .Z(n44692) );
  NAND U45020 ( .A(n44694), .B(n44693), .Z(n44689) );
  ANDN U45021 ( .B(B[104]), .A(n57), .Z(n44473) );
  XNOR U45022 ( .A(n44481), .B(n44695), .Z(n44474) );
  XNOR U45023 ( .A(n44480), .B(n44478), .Z(n44695) );
  AND U45024 ( .A(n44696), .B(n44697), .Z(n44478) );
  NANDN U45025 ( .A(n44698), .B(n44699), .Z(n44697) );
  NANDN U45026 ( .A(n44700), .B(n44701), .Z(n44699) );
  NANDN U45027 ( .A(n44701), .B(n44700), .Z(n44696) );
  ANDN U45028 ( .B(B[105]), .A(n58), .Z(n44480) );
  XNOR U45029 ( .A(n44488), .B(n44702), .Z(n44481) );
  XNOR U45030 ( .A(n44487), .B(n44485), .Z(n44702) );
  AND U45031 ( .A(n44703), .B(n44704), .Z(n44485) );
  NANDN U45032 ( .A(n44705), .B(n44706), .Z(n44704) );
  OR U45033 ( .A(n44707), .B(n44708), .Z(n44706) );
  NAND U45034 ( .A(n44708), .B(n44707), .Z(n44703) );
  ANDN U45035 ( .B(B[106]), .A(n59), .Z(n44487) );
  XNOR U45036 ( .A(n44495), .B(n44709), .Z(n44488) );
  XNOR U45037 ( .A(n44494), .B(n44492), .Z(n44709) );
  AND U45038 ( .A(n44710), .B(n44711), .Z(n44492) );
  NANDN U45039 ( .A(n44712), .B(n44713), .Z(n44711) );
  NANDN U45040 ( .A(n44714), .B(n44715), .Z(n44713) );
  NANDN U45041 ( .A(n44715), .B(n44714), .Z(n44710) );
  ANDN U45042 ( .B(B[107]), .A(n60), .Z(n44494) );
  XNOR U45043 ( .A(n44502), .B(n44716), .Z(n44495) );
  XNOR U45044 ( .A(n44501), .B(n44499), .Z(n44716) );
  AND U45045 ( .A(n44717), .B(n44718), .Z(n44499) );
  NANDN U45046 ( .A(n44719), .B(n44720), .Z(n44718) );
  OR U45047 ( .A(n44721), .B(n44722), .Z(n44720) );
  NAND U45048 ( .A(n44722), .B(n44721), .Z(n44717) );
  ANDN U45049 ( .B(B[108]), .A(n61), .Z(n44501) );
  XNOR U45050 ( .A(n44509), .B(n44723), .Z(n44502) );
  XNOR U45051 ( .A(n44508), .B(n44506), .Z(n44723) );
  AND U45052 ( .A(n44724), .B(n44725), .Z(n44506) );
  NANDN U45053 ( .A(n44726), .B(n44727), .Z(n44725) );
  NANDN U45054 ( .A(n44728), .B(n44729), .Z(n44727) );
  NANDN U45055 ( .A(n44729), .B(n44728), .Z(n44724) );
  ANDN U45056 ( .B(B[109]), .A(n62), .Z(n44508) );
  XNOR U45057 ( .A(n44516), .B(n44730), .Z(n44509) );
  XNOR U45058 ( .A(n44515), .B(n44513), .Z(n44730) );
  AND U45059 ( .A(n44731), .B(n44732), .Z(n44513) );
  NANDN U45060 ( .A(n44733), .B(n44734), .Z(n44732) );
  OR U45061 ( .A(n44735), .B(n44736), .Z(n44734) );
  NAND U45062 ( .A(n44736), .B(n44735), .Z(n44731) );
  ANDN U45063 ( .B(B[110]), .A(n63), .Z(n44515) );
  XNOR U45064 ( .A(n44523), .B(n44737), .Z(n44516) );
  XNOR U45065 ( .A(n44522), .B(n44520), .Z(n44737) );
  AND U45066 ( .A(n44738), .B(n44739), .Z(n44520) );
  NANDN U45067 ( .A(n44740), .B(n44741), .Z(n44739) );
  NANDN U45068 ( .A(n44742), .B(n44743), .Z(n44741) );
  NANDN U45069 ( .A(n44743), .B(n44742), .Z(n44738) );
  ANDN U45070 ( .B(B[111]), .A(n64), .Z(n44522) );
  XNOR U45071 ( .A(n44530), .B(n44744), .Z(n44523) );
  XNOR U45072 ( .A(n44529), .B(n44527), .Z(n44744) );
  AND U45073 ( .A(n44745), .B(n44746), .Z(n44527) );
  NANDN U45074 ( .A(n44747), .B(n44748), .Z(n44746) );
  OR U45075 ( .A(n44749), .B(n44750), .Z(n44748) );
  NAND U45076 ( .A(n44750), .B(n44749), .Z(n44745) );
  ANDN U45077 ( .B(B[112]), .A(n65), .Z(n44529) );
  XNOR U45078 ( .A(n44537), .B(n44751), .Z(n44530) );
  XNOR U45079 ( .A(n44536), .B(n44534), .Z(n44751) );
  AND U45080 ( .A(n44752), .B(n44753), .Z(n44534) );
  NANDN U45081 ( .A(n44754), .B(n44755), .Z(n44753) );
  NANDN U45082 ( .A(n44756), .B(n44757), .Z(n44755) );
  NANDN U45083 ( .A(n44757), .B(n44756), .Z(n44752) );
  ANDN U45084 ( .B(B[113]), .A(n66), .Z(n44536) );
  XNOR U45085 ( .A(n44544), .B(n44758), .Z(n44537) );
  XNOR U45086 ( .A(n44543), .B(n44541), .Z(n44758) );
  AND U45087 ( .A(n44759), .B(n44760), .Z(n44541) );
  NANDN U45088 ( .A(n44761), .B(n44762), .Z(n44760) );
  OR U45089 ( .A(n44763), .B(n44764), .Z(n44762) );
  NAND U45090 ( .A(n44764), .B(n44763), .Z(n44759) );
  ANDN U45091 ( .B(B[114]), .A(n67), .Z(n44543) );
  XNOR U45092 ( .A(n44551), .B(n44765), .Z(n44544) );
  XNOR U45093 ( .A(n44550), .B(n44548), .Z(n44765) );
  AND U45094 ( .A(n44766), .B(n44767), .Z(n44548) );
  NANDN U45095 ( .A(n44768), .B(n44769), .Z(n44767) );
  NANDN U45096 ( .A(n44770), .B(n44771), .Z(n44769) );
  NANDN U45097 ( .A(n44771), .B(n44770), .Z(n44766) );
  ANDN U45098 ( .B(B[115]), .A(n68), .Z(n44550) );
  XNOR U45099 ( .A(n44558), .B(n44772), .Z(n44551) );
  XNOR U45100 ( .A(n44557), .B(n44555), .Z(n44772) );
  AND U45101 ( .A(n44773), .B(n44774), .Z(n44555) );
  NANDN U45102 ( .A(n44775), .B(n44776), .Z(n44774) );
  OR U45103 ( .A(n44777), .B(n44778), .Z(n44776) );
  NAND U45104 ( .A(n44778), .B(n44777), .Z(n44773) );
  ANDN U45105 ( .B(B[116]), .A(n69), .Z(n44557) );
  XNOR U45106 ( .A(n44565), .B(n44779), .Z(n44558) );
  XNOR U45107 ( .A(n44564), .B(n44562), .Z(n44779) );
  AND U45108 ( .A(n44780), .B(n44781), .Z(n44562) );
  NANDN U45109 ( .A(n44782), .B(n44783), .Z(n44781) );
  NANDN U45110 ( .A(n44784), .B(n44785), .Z(n44783) );
  NANDN U45111 ( .A(n44785), .B(n44784), .Z(n44780) );
  ANDN U45112 ( .B(B[117]), .A(n70), .Z(n44564) );
  XNOR U45113 ( .A(n44572), .B(n44786), .Z(n44565) );
  XNOR U45114 ( .A(n44571), .B(n44569), .Z(n44786) );
  AND U45115 ( .A(n44787), .B(n44788), .Z(n44569) );
  NANDN U45116 ( .A(n44789), .B(n44790), .Z(n44788) );
  OR U45117 ( .A(n44791), .B(n44792), .Z(n44790) );
  NAND U45118 ( .A(n44792), .B(n44791), .Z(n44787) );
  ANDN U45119 ( .B(B[118]), .A(n71), .Z(n44571) );
  XNOR U45120 ( .A(n44579), .B(n44793), .Z(n44572) );
  XNOR U45121 ( .A(n44578), .B(n44576), .Z(n44793) );
  AND U45122 ( .A(n44794), .B(n44795), .Z(n44576) );
  NANDN U45123 ( .A(n44796), .B(n44797), .Z(n44795) );
  NANDN U45124 ( .A(n44798), .B(n44799), .Z(n44797) );
  NANDN U45125 ( .A(n44799), .B(n44798), .Z(n44794) );
  ANDN U45126 ( .B(B[119]), .A(n72), .Z(n44578) );
  XNOR U45127 ( .A(n44586), .B(n44800), .Z(n44579) );
  XNOR U45128 ( .A(n44585), .B(n44583), .Z(n44800) );
  AND U45129 ( .A(n44801), .B(n44802), .Z(n44583) );
  NANDN U45130 ( .A(n44803), .B(n44804), .Z(n44802) );
  OR U45131 ( .A(n44805), .B(n44806), .Z(n44804) );
  NAND U45132 ( .A(n44806), .B(n44805), .Z(n44801) );
  ANDN U45133 ( .B(B[120]), .A(n73), .Z(n44585) );
  XNOR U45134 ( .A(n44593), .B(n44807), .Z(n44586) );
  XNOR U45135 ( .A(n44592), .B(n44590), .Z(n44807) );
  AND U45136 ( .A(n44808), .B(n44809), .Z(n44590) );
  NANDN U45137 ( .A(n44810), .B(n44811), .Z(n44809) );
  NANDN U45138 ( .A(n44812), .B(n44813), .Z(n44811) );
  NANDN U45139 ( .A(n44813), .B(n44812), .Z(n44808) );
  ANDN U45140 ( .B(B[121]), .A(n74), .Z(n44592) );
  XNOR U45141 ( .A(n44600), .B(n44814), .Z(n44593) );
  XNOR U45142 ( .A(n44599), .B(n44597), .Z(n44814) );
  AND U45143 ( .A(n44815), .B(n44816), .Z(n44597) );
  NANDN U45144 ( .A(n44817), .B(n44818), .Z(n44816) );
  OR U45145 ( .A(n44819), .B(n44820), .Z(n44818) );
  NAND U45146 ( .A(n44820), .B(n44819), .Z(n44815) );
  ANDN U45147 ( .B(B[122]), .A(n75), .Z(n44599) );
  XNOR U45148 ( .A(n44607), .B(n44821), .Z(n44600) );
  XNOR U45149 ( .A(n44606), .B(n44604), .Z(n44821) );
  AND U45150 ( .A(n44822), .B(n44823), .Z(n44604) );
  NANDN U45151 ( .A(n44824), .B(n44825), .Z(n44823) );
  NANDN U45152 ( .A(n44826), .B(n44827), .Z(n44825) );
  NANDN U45153 ( .A(n44827), .B(n44826), .Z(n44822) );
  ANDN U45154 ( .B(B[123]), .A(n76), .Z(n44606) );
  XNOR U45155 ( .A(n44614), .B(n44828), .Z(n44607) );
  XNOR U45156 ( .A(n44613), .B(n44611), .Z(n44828) );
  AND U45157 ( .A(n44829), .B(n44830), .Z(n44611) );
  NANDN U45158 ( .A(n44831), .B(n44832), .Z(n44830) );
  OR U45159 ( .A(n44833), .B(n44834), .Z(n44832) );
  NAND U45160 ( .A(n44834), .B(n44833), .Z(n44829) );
  ANDN U45161 ( .B(B[124]), .A(n77), .Z(n44613) );
  XNOR U45162 ( .A(n44621), .B(n44835), .Z(n44614) );
  XNOR U45163 ( .A(n44620), .B(n44618), .Z(n44835) );
  AND U45164 ( .A(n44836), .B(n44837), .Z(n44618) );
  NANDN U45165 ( .A(n44838), .B(n44839), .Z(n44837) );
  NANDN U45166 ( .A(n44840), .B(n44841), .Z(n44839) );
  NANDN U45167 ( .A(n44841), .B(n44840), .Z(n44836) );
  ANDN U45168 ( .B(B[125]), .A(n78), .Z(n44620) );
  XNOR U45169 ( .A(n44628), .B(n44842), .Z(n44621) );
  XNOR U45170 ( .A(n44627), .B(n44625), .Z(n44842) );
  AND U45171 ( .A(n44843), .B(n44844), .Z(n44625) );
  NANDN U45172 ( .A(n44845), .B(n44846), .Z(n44844) );
  OR U45173 ( .A(n44847), .B(n44848), .Z(n44846) );
  NAND U45174 ( .A(n44848), .B(n44847), .Z(n44843) );
  ANDN U45175 ( .B(B[126]), .A(n79), .Z(n44627) );
  XNOR U45176 ( .A(n44635), .B(n44849), .Z(n44628) );
  XNOR U45177 ( .A(n44634), .B(n44632), .Z(n44849) );
  AND U45178 ( .A(n44850), .B(n44851), .Z(n44632) );
  NANDN U45179 ( .A(n44852), .B(n44853), .Z(n44851) );
  NANDN U45180 ( .A(n44854), .B(n44855), .Z(n44853) );
  NANDN U45181 ( .A(n44855), .B(n44854), .Z(n44850) );
  ANDN U45182 ( .B(B[127]), .A(n80), .Z(n44634) );
  XNOR U45183 ( .A(n44642), .B(n44856), .Z(n44635) );
  XNOR U45184 ( .A(n44641), .B(n44639), .Z(n44856) );
  AND U45185 ( .A(n44857), .B(n44858), .Z(n44639) );
  NANDN U45186 ( .A(n44859), .B(n44860), .Z(n44858) );
  OR U45187 ( .A(n44861), .B(n44862), .Z(n44860) );
  NAND U45188 ( .A(n44862), .B(n44861), .Z(n44857) );
  ANDN U45189 ( .B(B[128]), .A(n81), .Z(n44641) );
  XNOR U45190 ( .A(n44649), .B(n44863), .Z(n44642) );
  XNOR U45191 ( .A(n44648), .B(n44646), .Z(n44863) );
  AND U45192 ( .A(n44864), .B(n44865), .Z(n44646) );
  NANDN U45193 ( .A(n44866), .B(n44867), .Z(n44865) );
  NAND U45194 ( .A(n44868), .B(n44869), .Z(n44867) );
  ANDN U45195 ( .B(B[129]), .A(n82), .Z(n44648) );
  XOR U45196 ( .A(n44655), .B(n44870), .Z(n44649) );
  XNOR U45197 ( .A(n44653), .B(n44656), .Z(n44870) );
  NAND U45198 ( .A(A[2]), .B(B[130]), .Z(n44656) );
  NANDN U45199 ( .A(n44871), .B(n44872), .Z(n44653) );
  AND U45200 ( .A(A[0]), .B(B[131]), .Z(n44872) );
  XNOR U45201 ( .A(n44658), .B(n44873), .Z(n44655) );
  NAND U45202 ( .A(A[0]), .B(B[132]), .Z(n44873) );
  NAND U45203 ( .A(B[131]), .B(A[1]), .Z(n44658) );
  NAND U45204 ( .A(n44874), .B(n44875), .Z(n532) );
  NANDN U45205 ( .A(n44876), .B(n44877), .Z(n44875) );
  OR U45206 ( .A(n44878), .B(n44879), .Z(n44877) );
  NAND U45207 ( .A(n44879), .B(n44878), .Z(n44874) );
  XOR U45208 ( .A(n42661), .B(n44880), .Z(\A1[12] ) );
  XNOR U45209 ( .A(n42660), .B(n42659), .Z(n44880) );
  NAND U45210 ( .A(n44881), .B(n44882), .Z(n42659) );
  NANDN U45211 ( .A(n44883), .B(n44884), .Z(n44882) );
  OR U45212 ( .A(n44885), .B(n44886), .Z(n44884) );
  NAND U45213 ( .A(n44886), .B(n44885), .Z(n44881) );
  ANDN U45214 ( .B(B[0]), .A(n71), .Z(n42660) );
  XNOR U45215 ( .A(n42668), .B(n44887), .Z(n42661) );
  XNOR U45216 ( .A(n42667), .B(n42665), .Z(n44887) );
  AND U45217 ( .A(n44888), .B(n44889), .Z(n42665) );
  NANDN U45218 ( .A(n44890), .B(n44891), .Z(n44889) );
  NANDN U45219 ( .A(n44892), .B(n44893), .Z(n44891) );
  NANDN U45220 ( .A(n44893), .B(n44892), .Z(n44888) );
  ANDN U45221 ( .B(B[1]), .A(n72), .Z(n42667) );
  XNOR U45222 ( .A(n42675), .B(n44894), .Z(n42668) );
  XNOR U45223 ( .A(n42674), .B(n42672), .Z(n44894) );
  AND U45224 ( .A(n44895), .B(n44896), .Z(n42672) );
  NANDN U45225 ( .A(n44897), .B(n44898), .Z(n44896) );
  OR U45226 ( .A(n44899), .B(n44900), .Z(n44898) );
  NAND U45227 ( .A(n44900), .B(n44899), .Z(n44895) );
  ANDN U45228 ( .B(B[2]), .A(n73), .Z(n42674) );
  XNOR U45229 ( .A(n42682), .B(n44901), .Z(n42675) );
  XNOR U45230 ( .A(n42681), .B(n42679), .Z(n44901) );
  AND U45231 ( .A(n44902), .B(n44903), .Z(n42679) );
  NANDN U45232 ( .A(n44904), .B(n44905), .Z(n44903) );
  NANDN U45233 ( .A(n44906), .B(n44907), .Z(n44905) );
  NANDN U45234 ( .A(n44907), .B(n44906), .Z(n44902) );
  ANDN U45235 ( .B(B[3]), .A(n74), .Z(n42681) );
  XNOR U45236 ( .A(n42689), .B(n44908), .Z(n42682) );
  XNOR U45237 ( .A(n42688), .B(n42686), .Z(n44908) );
  AND U45238 ( .A(n44909), .B(n44910), .Z(n42686) );
  NANDN U45239 ( .A(n44911), .B(n44912), .Z(n44910) );
  OR U45240 ( .A(n44913), .B(n44914), .Z(n44912) );
  NAND U45241 ( .A(n44914), .B(n44913), .Z(n44909) );
  ANDN U45242 ( .B(B[4]), .A(n75), .Z(n42688) );
  XNOR U45243 ( .A(n42696), .B(n44915), .Z(n42689) );
  XNOR U45244 ( .A(n42695), .B(n42693), .Z(n44915) );
  AND U45245 ( .A(n44916), .B(n44917), .Z(n42693) );
  NANDN U45246 ( .A(n44918), .B(n44919), .Z(n44917) );
  NANDN U45247 ( .A(n44920), .B(n44921), .Z(n44919) );
  NANDN U45248 ( .A(n44921), .B(n44920), .Z(n44916) );
  ANDN U45249 ( .B(B[5]), .A(n76), .Z(n42695) );
  XNOR U45250 ( .A(n42703), .B(n44922), .Z(n42696) );
  XNOR U45251 ( .A(n42702), .B(n42700), .Z(n44922) );
  AND U45252 ( .A(n44923), .B(n44924), .Z(n42700) );
  NANDN U45253 ( .A(n44925), .B(n44926), .Z(n44924) );
  OR U45254 ( .A(n44927), .B(n44928), .Z(n44926) );
  NAND U45255 ( .A(n44928), .B(n44927), .Z(n44923) );
  ANDN U45256 ( .B(B[6]), .A(n77), .Z(n42702) );
  XNOR U45257 ( .A(n42710), .B(n44929), .Z(n42703) );
  XNOR U45258 ( .A(n42709), .B(n42707), .Z(n44929) );
  AND U45259 ( .A(n44930), .B(n44931), .Z(n42707) );
  NANDN U45260 ( .A(n44932), .B(n44933), .Z(n44931) );
  NANDN U45261 ( .A(n44934), .B(n44935), .Z(n44933) );
  NANDN U45262 ( .A(n44935), .B(n44934), .Z(n44930) );
  ANDN U45263 ( .B(B[7]), .A(n78), .Z(n42709) );
  XNOR U45264 ( .A(n42717), .B(n44936), .Z(n42710) );
  XNOR U45265 ( .A(n42716), .B(n42714), .Z(n44936) );
  AND U45266 ( .A(n44937), .B(n44938), .Z(n42714) );
  NANDN U45267 ( .A(n44939), .B(n44940), .Z(n44938) );
  OR U45268 ( .A(n44941), .B(n44942), .Z(n44940) );
  NAND U45269 ( .A(n44942), .B(n44941), .Z(n44937) );
  ANDN U45270 ( .B(B[8]), .A(n79), .Z(n42716) );
  XNOR U45271 ( .A(n42724), .B(n44943), .Z(n42717) );
  XNOR U45272 ( .A(n42723), .B(n42721), .Z(n44943) );
  AND U45273 ( .A(n44944), .B(n44945), .Z(n42721) );
  NANDN U45274 ( .A(n44946), .B(n44947), .Z(n44945) );
  NANDN U45275 ( .A(n44948), .B(n44949), .Z(n44947) );
  NANDN U45276 ( .A(n44949), .B(n44948), .Z(n44944) );
  ANDN U45277 ( .B(B[9]), .A(n80), .Z(n42723) );
  XNOR U45278 ( .A(n42731), .B(n44950), .Z(n42724) );
  XNOR U45279 ( .A(n42730), .B(n42728), .Z(n44950) );
  AND U45280 ( .A(n44951), .B(n44952), .Z(n42728) );
  NANDN U45281 ( .A(n44953), .B(n44954), .Z(n44952) );
  OR U45282 ( .A(n44955), .B(n44956), .Z(n44954) );
  NAND U45283 ( .A(n44956), .B(n44955), .Z(n44951) );
  ANDN U45284 ( .B(B[10]), .A(n81), .Z(n42730) );
  XNOR U45285 ( .A(n42738), .B(n44957), .Z(n42731) );
  XNOR U45286 ( .A(n42737), .B(n42735), .Z(n44957) );
  AND U45287 ( .A(n44958), .B(n44959), .Z(n42735) );
  NANDN U45288 ( .A(n44960), .B(n44961), .Z(n44959) );
  NAND U45289 ( .A(n44962), .B(n44963), .Z(n44961) );
  ANDN U45290 ( .B(B[11]), .A(n82), .Z(n42737) );
  XOR U45291 ( .A(n42744), .B(n44964), .Z(n42738) );
  XNOR U45292 ( .A(n42742), .B(n42745), .Z(n44964) );
  NAND U45293 ( .A(A[2]), .B(B[12]), .Z(n42745) );
  NANDN U45294 ( .A(n44965), .B(n44966), .Z(n42742) );
  AND U45295 ( .A(A[0]), .B(B[13]), .Z(n44966) );
  XNOR U45296 ( .A(n42747), .B(n44967), .Z(n42744) );
  NAND U45297 ( .A(A[0]), .B(B[14]), .Z(n44967) );
  NAND U45298 ( .A(B[13]), .B(A[1]), .Z(n42747) );
  XOR U45299 ( .A(n534), .B(n533), .Z(\A1[129] ) );
  XOR U45300 ( .A(n44879), .B(n44968), .Z(n533) );
  XNOR U45301 ( .A(n44878), .B(n44876), .Z(n44968) );
  AND U45302 ( .A(n44969), .B(n44970), .Z(n44876) );
  NANDN U45303 ( .A(n44971), .B(n44972), .Z(n44970) );
  NANDN U45304 ( .A(n44973), .B(n44974), .Z(n44972) );
  NANDN U45305 ( .A(n44974), .B(n44973), .Z(n44969) );
  ANDN U45306 ( .B(A[31]), .A(n4), .Z(n44878) );
  XNOR U45307 ( .A(n44673), .B(n44975), .Z(n44879) );
  XNOR U45308 ( .A(n44672), .B(n44670), .Z(n44975) );
  AND U45309 ( .A(n44976), .B(n44977), .Z(n44670) );
  NANDN U45310 ( .A(n44978), .B(n44979), .Z(n44977) );
  OR U45311 ( .A(n44980), .B(n44981), .Z(n44979) );
  NAND U45312 ( .A(n44981), .B(n44980), .Z(n44976) );
  ANDN U45313 ( .B(B[101]), .A(n55), .Z(n44672) );
  XNOR U45314 ( .A(n44680), .B(n44982), .Z(n44673) );
  XNOR U45315 ( .A(n44679), .B(n44677), .Z(n44982) );
  AND U45316 ( .A(n44983), .B(n44984), .Z(n44677) );
  NANDN U45317 ( .A(n44985), .B(n44986), .Z(n44984) );
  NANDN U45318 ( .A(n44987), .B(n44988), .Z(n44986) );
  NANDN U45319 ( .A(n44988), .B(n44987), .Z(n44983) );
  ANDN U45320 ( .B(B[102]), .A(n56), .Z(n44679) );
  XNOR U45321 ( .A(n44687), .B(n44989), .Z(n44680) );
  XNOR U45322 ( .A(n44686), .B(n44684), .Z(n44989) );
  AND U45323 ( .A(n44990), .B(n44991), .Z(n44684) );
  NANDN U45324 ( .A(n44992), .B(n44993), .Z(n44991) );
  OR U45325 ( .A(n44994), .B(n44995), .Z(n44993) );
  NAND U45326 ( .A(n44995), .B(n44994), .Z(n44990) );
  ANDN U45327 ( .B(B[103]), .A(n57), .Z(n44686) );
  XNOR U45328 ( .A(n44694), .B(n44996), .Z(n44687) );
  XNOR U45329 ( .A(n44693), .B(n44691), .Z(n44996) );
  AND U45330 ( .A(n44997), .B(n44998), .Z(n44691) );
  NANDN U45331 ( .A(n44999), .B(n45000), .Z(n44998) );
  NANDN U45332 ( .A(n45001), .B(n45002), .Z(n45000) );
  NANDN U45333 ( .A(n45002), .B(n45001), .Z(n44997) );
  ANDN U45334 ( .B(B[104]), .A(n58), .Z(n44693) );
  XNOR U45335 ( .A(n44701), .B(n45003), .Z(n44694) );
  XNOR U45336 ( .A(n44700), .B(n44698), .Z(n45003) );
  AND U45337 ( .A(n45004), .B(n45005), .Z(n44698) );
  NANDN U45338 ( .A(n45006), .B(n45007), .Z(n45005) );
  OR U45339 ( .A(n45008), .B(n45009), .Z(n45007) );
  NAND U45340 ( .A(n45009), .B(n45008), .Z(n45004) );
  ANDN U45341 ( .B(B[105]), .A(n59), .Z(n44700) );
  XNOR U45342 ( .A(n44708), .B(n45010), .Z(n44701) );
  XNOR U45343 ( .A(n44707), .B(n44705), .Z(n45010) );
  AND U45344 ( .A(n45011), .B(n45012), .Z(n44705) );
  NANDN U45345 ( .A(n45013), .B(n45014), .Z(n45012) );
  NANDN U45346 ( .A(n45015), .B(n45016), .Z(n45014) );
  NANDN U45347 ( .A(n45016), .B(n45015), .Z(n45011) );
  ANDN U45348 ( .B(B[106]), .A(n60), .Z(n44707) );
  XNOR U45349 ( .A(n44715), .B(n45017), .Z(n44708) );
  XNOR U45350 ( .A(n44714), .B(n44712), .Z(n45017) );
  AND U45351 ( .A(n45018), .B(n45019), .Z(n44712) );
  NANDN U45352 ( .A(n45020), .B(n45021), .Z(n45019) );
  OR U45353 ( .A(n45022), .B(n45023), .Z(n45021) );
  NAND U45354 ( .A(n45023), .B(n45022), .Z(n45018) );
  ANDN U45355 ( .B(B[107]), .A(n61), .Z(n44714) );
  XNOR U45356 ( .A(n44722), .B(n45024), .Z(n44715) );
  XNOR U45357 ( .A(n44721), .B(n44719), .Z(n45024) );
  AND U45358 ( .A(n45025), .B(n45026), .Z(n44719) );
  NANDN U45359 ( .A(n45027), .B(n45028), .Z(n45026) );
  NANDN U45360 ( .A(n45029), .B(n45030), .Z(n45028) );
  NANDN U45361 ( .A(n45030), .B(n45029), .Z(n45025) );
  ANDN U45362 ( .B(B[108]), .A(n62), .Z(n44721) );
  XNOR U45363 ( .A(n44729), .B(n45031), .Z(n44722) );
  XNOR U45364 ( .A(n44728), .B(n44726), .Z(n45031) );
  AND U45365 ( .A(n45032), .B(n45033), .Z(n44726) );
  NANDN U45366 ( .A(n45034), .B(n45035), .Z(n45033) );
  OR U45367 ( .A(n45036), .B(n45037), .Z(n45035) );
  NAND U45368 ( .A(n45037), .B(n45036), .Z(n45032) );
  ANDN U45369 ( .B(B[109]), .A(n63), .Z(n44728) );
  XNOR U45370 ( .A(n44736), .B(n45038), .Z(n44729) );
  XNOR U45371 ( .A(n44735), .B(n44733), .Z(n45038) );
  AND U45372 ( .A(n45039), .B(n45040), .Z(n44733) );
  NANDN U45373 ( .A(n45041), .B(n45042), .Z(n45040) );
  NANDN U45374 ( .A(n45043), .B(n45044), .Z(n45042) );
  NANDN U45375 ( .A(n45044), .B(n45043), .Z(n45039) );
  ANDN U45376 ( .B(B[110]), .A(n64), .Z(n44735) );
  XNOR U45377 ( .A(n44743), .B(n45045), .Z(n44736) );
  XNOR U45378 ( .A(n44742), .B(n44740), .Z(n45045) );
  AND U45379 ( .A(n45046), .B(n45047), .Z(n44740) );
  NANDN U45380 ( .A(n45048), .B(n45049), .Z(n45047) );
  OR U45381 ( .A(n45050), .B(n45051), .Z(n45049) );
  NAND U45382 ( .A(n45051), .B(n45050), .Z(n45046) );
  ANDN U45383 ( .B(B[111]), .A(n65), .Z(n44742) );
  XNOR U45384 ( .A(n44750), .B(n45052), .Z(n44743) );
  XNOR U45385 ( .A(n44749), .B(n44747), .Z(n45052) );
  AND U45386 ( .A(n45053), .B(n45054), .Z(n44747) );
  NANDN U45387 ( .A(n45055), .B(n45056), .Z(n45054) );
  NANDN U45388 ( .A(n45057), .B(n45058), .Z(n45056) );
  NANDN U45389 ( .A(n45058), .B(n45057), .Z(n45053) );
  ANDN U45390 ( .B(B[112]), .A(n66), .Z(n44749) );
  XNOR U45391 ( .A(n44757), .B(n45059), .Z(n44750) );
  XNOR U45392 ( .A(n44756), .B(n44754), .Z(n45059) );
  AND U45393 ( .A(n45060), .B(n45061), .Z(n44754) );
  NANDN U45394 ( .A(n45062), .B(n45063), .Z(n45061) );
  OR U45395 ( .A(n45064), .B(n45065), .Z(n45063) );
  NAND U45396 ( .A(n45065), .B(n45064), .Z(n45060) );
  ANDN U45397 ( .B(B[113]), .A(n67), .Z(n44756) );
  XNOR U45398 ( .A(n44764), .B(n45066), .Z(n44757) );
  XNOR U45399 ( .A(n44763), .B(n44761), .Z(n45066) );
  AND U45400 ( .A(n45067), .B(n45068), .Z(n44761) );
  NANDN U45401 ( .A(n45069), .B(n45070), .Z(n45068) );
  NANDN U45402 ( .A(n45071), .B(n45072), .Z(n45070) );
  NANDN U45403 ( .A(n45072), .B(n45071), .Z(n45067) );
  ANDN U45404 ( .B(B[114]), .A(n68), .Z(n44763) );
  XNOR U45405 ( .A(n44771), .B(n45073), .Z(n44764) );
  XNOR U45406 ( .A(n44770), .B(n44768), .Z(n45073) );
  AND U45407 ( .A(n45074), .B(n45075), .Z(n44768) );
  NANDN U45408 ( .A(n45076), .B(n45077), .Z(n45075) );
  OR U45409 ( .A(n45078), .B(n45079), .Z(n45077) );
  NAND U45410 ( .A(n45079), .B(n45078), .Z(n45074) );
  ANDN U45411 ( .B(B[115]), .A(n69), .Z(n44770) );
  XNOR U45412 ( .A(n44778), .B(n45080), .Z(n44771) );
  XNOR U45413 ( .A(n44777), .B(n44775), .Z(n45080) );
  AND U45414 ( .A(n45081), .B(n45082), .Z(n44775) );
  NANDN U45415 ( .A(n45083), .B(n45084), .Z(n45082) );
  NANDN U45416 ( .A(n45085), .B(n45086), .Z(n45084) );
  NANDN U45417 ( .A(n45086), .B(n45085), .Z(n45081) );
  ANDN U45418 ( .B(B[116]), .A(n70), .Z(n44777) );
  XNOR U45419 ( .A(n44785), .B(n45087), .Z(n44778) );
  XNOR U45420 ( .A(n44784), .B(n44782), .Z(n45087) );
  AND U45421 ( .A(n45088), .B(n45089), .Z(n44782) );
  NANDN U45422 ( .A(n45090), .B(n45091), .Z(n45089) );
  OR U45423 ( .A(n45092), .B(n45093), .Z(n45091) );
  NAND U45424 ( .A(n45093), .B(n45092), .Z(n45088) );
  ANDN U45425 ( .B(B[117]), .A(n71), .Z(n44784) );
  XNOR U45426 ( .A(n44792), .B(n45094), .Z(n44785) );
  XNOR U45427 ( .A(n44791), .B(n44789), .Z(n45094) );
  AND U45428 ( .A(n45095), .B(n45096), .Z(n44789) );
  NANDN U45429 ( .A(n45097), .B(n45098), .Z(n45096) );
  NANDN U45430 ( .A(n45099), .B(n45100), .Z(n45098) );
  NANDN U45431 ( .A(n45100), .B(n45099), .Z(n45095) );
  ANDN U45432 ( .B(B[118]), .A(n72), .Z(n44791) );
  XNOR U45433 ( .A(n44799), .B(n45101), .Z(n44792) );
  XNOR U45434 ( .A(n44798), .B(n44796), .Z(n45101) );
  AND U45435 ( .A(n45102), .B(n45103), .Z(n44796) );
  NANDN U45436 ( .A(n45104), .B(n45105), .Z(n45103) );
  OR U45437 ( .A(n45106), .B(n45107), .Z(n45105) );
  NAND U45438 ( .A(n45107), .B(n45106), .Z(n45102) );
  ANDN U45439 ( .B(B[119]), .A(n73), .Z(n44798) );
  XNOR U45440 ( .A(n44806), .B(n45108), .Z(n44799) );
  XNOR U45441 ( .A(n44805), .B(n44803), .Z(n45108) );
  AND U45442 ( .A(n45109), .B(n45110), .Z(n44803) );
  NANDN U45443 ( .A(n45111), .B(n45112), .Z(n45110) );
  NANDN U45444 ( .A(n45113), .B(n45114), .Z(n45112) );
  NANDN U45445 ( .A(n45114), .B(n45113), .Z(n45109) );
  ANDN U45446 ( .B(B[120]), .A(n74), .Z(n44805) );
  XNOR U45447 ( .A(n44813), .B(n45115), .Z(n44806) );
  XNOR U45448 ( .A(n44812), .B(n44810), .Z(n45115) );
  AND U45449 ( .A(n45116), .B(n45117), .Z(n44810) );
  NANDN U45450 ( .A(n45118), .B(n45119), .Z(n45117) );
  OR U45451 ( .A(n45120), .B(n45121), .Z(n45119) );
  NAND U45452 ( .A(n45121), .B(n45120), .Z(n45116) );
  ANDN U45453 ( .B(B[121]), .A(n75), .Z(n44812) );
  XNOR U45454 ( .A(n44820), .B(n45122), .Z(n44813) );
  XNOR U45455 ( .A(n44819), .B(n44817), .Z(n45122) );
  AND U45456 ( .A(n45123), .B(n45124), .Z(n44817) );
  NANDN U45457 ( .A(n45125), .B(n45126), .Z(n45124) );
  NANDN U45458 ( .A(n45127), .B(n45128), .Z(n45126) );
  NANDN U45459 ( .A(n45128), .B(n45127), .Z(n45123) );
  ANDN U45460 ( .B(B[122]), .A(n76), .Z(n44819) );
  XNOR U45461 ( .A(n44827), .B(n45129), .Z(n44820) );
  XNOR U45462 ( .A(n44826), .B(n44824), .Z(n45129) );
  AND U45463 ( .A(n45130), .B(n45131), .Z(n44824) );
  NANDN U45464 ( .A(n45132), .B(n45133), .Z(n45131) );
  OR U45465 ( .A(n45134), .B(n45135), .Z(n45133) );
  NAND U45466 ( .A(n45135), .B(n45134), .Z(n45130) );
  ANDN U45467 ( .B(B[123]), .A(n77), .Z(n44826) );
  XNOR U45468 ( .A(n44834), .B(n45136), .Z(n44827) );
  XNOR U45469 ( .A(n44833), .B(n44831), .Z(n45136) );
  AND U45470 ( .A(n45137), .B(n45138), .Z(n44831) );
  NANDN U45471 ( .A(n45139), .B(n45140), .Z(n45138) );
  NANDN U45472 ( .A(n45141), .B(n45142), .Z(n45140) );
  NANDN U45473 ( .A(n45142), .B(n45141), .Z(n45137) );
  ANDN U45474 ( .B(B[124]), .A(n78), .Z(n44833) );
  XNOR U45475 ( .A(n44841), .B(n45143), .Z(n44834) );
  XNOR U45476 ( .A(n44840), .B(n44838), .Z(n45143) );
  AND U45477 ( .A(n45144), .B(n45145), .Z(n44838) );
  NANDN U45478 ( .A(n45146), .B(n45147), .Z(n45145) );
  OR U45479 ( .A(n45148), .B(n45149), .Z(n45147) );
  NAND U45480 ( .A(n45149), .B(n45148), .Z(n45144) );
  ANDN U45481 ( .B(B[125]), .A(n79), .Z(n44840) );
  XNOR U45482 ( .A(n44848), .B(n45150), .Z(n44841) );
  XNOR U45483 ( .A(n44847), .B(n44845), .Z(n45150) );
  AND U45484 ( .A(n45151), .B(n45152), .Z(n44845) );
  NANDN U45485 ( .A(n45153), .B(n45154), .Z(n45152) );
  NANDN U45486 ( .A(n45155), .B(n45156), .Z(n45154) );
  NANDN U45487 ( .A(n45156), .B(n45155), .Z(n45151) );
  ANDN U45488 ( .B(B[126]), .A(n80), .Z(n44847) );
  XNOR U45489 ( .A(n44855), .B(n45157), .Z(n44848) );
  XNOR U45490 ( .A(n44854), .B(n44852), .Z(n45157) );
  AND U45491 ( .A(n45158), .B(n45159), .Z(n44852) );
  NANDN U45492 ( .A(n45160), .B(n45161), .Z(n45159) );
  OR U45493 ( .A(n45162), .B(n45163), .Z(n45161) );
  NAND U45494 ( .A(n45163), .B(n45162), .Z(n45158) );
  ANDN U45495 ( .B(B[127]), .A(n81), .Z(n44854) );
  XNOR U45496 ( .A(n44862), .B(n45164), .Z(n44855) );
  XNOR U45497 ( .A(n44861), .B(n44859), .Z(n45164) );
  AND U45498 ( .A(n45165), .B(n45166), .Z(n44859) );
  NANDN U45499 ( .A(n45167), .B(n45168), .Z(n45166) );
  NAND U45500 ( .A(n45169), .B(n45170), .Z(n45168) );
  ANDN U45501 ( .B(B[128]), .A(n82), .Z(n44861) );
  XOR U45502 ( .A(n44868), .B(n45171), .Z(n44862) );
  XNOR U45503 ( .A(n44866), .B(n44869), .Z(n45171) );
  NAND U45504 ( .A(A[2]), .B(B[129]), .Z(n44869) );
  NANDN U45505 ( .A(n45172), .B(n45173), .Z(n44866) );
  AND U45506 ( .A(A[0]), .B(B[130]), .Z(n45173) );
  XNOR U45507 ( .A(n44871), .B(n45174), .Z(n44868) );
  NAND U45508 ( .A(A[0]), .B(B[131]), .Z(n45174) );
  NAND U45509 ( .A(B[130]), .B(A[1]), .Z(n44871) );
  NAND U45510 ( .A(n45175), .B(n45176), .Z(n534) );
  NANDN U45511 ( .A(n45177), .B(n45178), .Z(n45176) );
  OR U45512 ( .A(n45179), .B(n45180), .Z(n45178) );
  NAND U45513 ( .A(n45180), .B(n45179), .Z(n45175) );
  XOR U45514 ( .A(n536), .B(n535), .Z(\A1[128] ) );
  XOR U45515 ( .A(n45180), .B(n45181), .Z(n535) );
  XNOR U45516 ( .A(n45179), .B(n45177), .Z(n45181) );
  AND U45517 ( .A(n45182), .B(n45183), .Z(n45177) );
  NANDN U45518 ( .A(n45184), .B(n45185), .Z(n45183) );
  NANDN U45519 ( .A(n45186), .B(n45187), .Z(n45185) );
  NANDN U45520 ( .A(n45187), .B(n45186), .Z(n45182) );
  ANDN U45521 ( .B(A[31]), .A(n6), .Z(n45179) );
  XNOR U45522 ( .A(n44974), .B(n45188), .Z(n45180) );
  XNOR U45523 ( .A(n44973), .B(n44971), .Z(n45188) );
  AND U45524 ( .A(n45189), .B(n45190), .Z(n44971) );
  NANDN U45525 ( .A(n45191), .B(n45192), .Z(n45190) );
  OR U45526 ( .A(n45193), .B(n45194), .Z(n45192) );
  NAND U45527 ( .A(n45194), .B(n45193), .Z(n45189) );
  ANDN U45528 ( .B(A[30]), .A(n4), .Z(n44973) );
  XNOR U45529 ( .A(n44981), .B(n45195), .Z(n44974) );
  XNOR U45530 ( .A(n44980), .B(n44978), .Z(n45195) );
  AND U45531 ( .A(n45196), .B(n45197), .Z(n44978) );
  NANDN U45532 ( .A(n45198), .B(n45199), .Z(n45197) );
  NANDN U45533 ( .A(n45200), .B(n45201), .Z(n45199) );
  NANDN U45534 ( .A(n45201), .B(n45200), .Z(n45196) );
  ANDN U45535 ( .B(B[101]), .A(n56), .Z(n44980) );
  XNOR U45536 ( .A(n44988), .B(n45202), .Z(n44981) );
  XNOR U45537 ( .A(n44987), .B(n44985), .Z(n45202) );
  AND U45538 ( .A(n45203), .B(n45204), .Z(n44985) );
  NANDN U45539 ( .A(n45205), .B(n45206), .Z(n45204) );
  OR U45540 ( .A(n45207), .B(n45208), .Z(n45206) );
  NAND U45541 ( .A(n45208), .B(n45207), .Z(n45203) );
  ANDN U45542 ( .B(B[102]), .A(n57), .Z(n44987) );
  XNOR U45543 ( .A(n44995), .B(n45209), .Z(n44988) );
  XNOR U45544 ( .A(n44994), .B(n44992), .Z(n45209) );
  AND U45545 ( .A(n45210), .B(n45211), .Z(n44992) );
  NANDN U45546 ( .A(n45212), .B(n45213), .Z(n45211) );
  NANDN U45547 ( .A(n45214), .B(n45215), .Z(n45213) );
  NANDN U45548 ( .A(n45215), .B(n45214), .Z(n45210) );
  ANDN U45549 ( .B(B[103]), .A(n58), .Z(n44994) );
  XNOR U45550 ( .A(n45002), .B(n45216), .Z(n44995) );
  XNOR U45551 ( .A(n45001), .B(n44999), .Z(n45216) );
  AND U45552 ( .A(n45217), .B(n45218), .Z(n44999) );
  NANDN U45553 ( .A(n45219), .B(n45220), .Z(n45218) );
  OR U45554 ( .A(n45221), .B(n45222), .Z(n45220) );
  NAND U45555 ( .A(n45222), .B(n45221), .Z(n45217) );
  ANDN U45556 ( .B(B[104]), .A(n59), .Z(n45001) );
  XNOR U45557 ( .A(n45009), .B(n45223), .Z(n45002) );
  XNOR U45558 ( .A(n45008), .B(n45006), .Z(n45223) );
  AND U45559 ( .A(n45224), .B(n45225), .Z(n45006) );
  NANDN U45560 ( .A(n45226), .B(n45227), .Z(n45225) );
  NANDN U45561 ( .A(n45228), .B(n45229), .Z(n45227) );
  NANDN U45562 ( .A(n45229), .B(n45228), .Z(n45224) );
  ANDN U45563 ( .B(B[105]), .A(n60), .Z(n45008) );
  XNOR U45564 ( .A(n45016), .B(n45230), .Z(n45009) );
  XNOR U45565 ( .A(n45015), .B(n45013), .Z(n45230) );
  AND U45566 ( .A(n45231), .B(n45232), .Z(n45013) );
  NANDN U45567 ( .A(n45233), .B(n45234), .Z(n45232) );
  OR U45568 ( .A(n45235), .B(n45236), .Z(n45234) );
  NAND U45569 ( .A(n45236), .B(n45235), .Z(n45231) );
  ANDN U45570 ( .B(B[106]), .A(n61), .Z(n45015) );
  XNOR U45571 ( .A(n45023), .B(n45237), .Z(n45016) );
  XNOR U45572 ( .A(n45022), .B(n45020), .Z(n45237) );
  AND U45573 ( .A(n45238), .B(n45239), .Z(n45020) );
  NANDN U45574 ( .A(n45240), .B(n45241), .Z(n45239) );
  NANDN U45575 ( .A(n45242), .B(n45243), .Z(n45241) );
  NANDN U45576 ( .A(n45243), .B(n45242), .Z(n45238) );
  ANDN U45577 ( .B(B[107]), .A(n62), .Z(n45022) );
  XNOR U45578 ( .A(n45030), .B(n45244), .Z(n45023) );
  XNOR U45579 ( .A(n45029), .B(n45027), .Z(n45244) );
  AND U45580 ( .A(n45245), .B(n45246), .Z(n45027) );
  NANDN U45581 ( .A(n45247), .B(n45248), .Z(n45246) );
  OR U45582 ( .A(n45249), .B(n45250), .Z(n45248) );
  NAND U45583 ( .A(n45250), .B(n45249), .Z(n45245) );
  ANDN U45584 ( .B(B[108]), .A(n63), .Z(n45029) );
  XNOR U45585 ( .A(n45037), .B(n45251), .Z(n45030) );
  XNOR U45586 ( .A(n45036), .B(n45034), .Z(n45251) );
  AND U45587 ( .A(n45252), .B(n45253), .Z(n45034) );
  NANDN U45588 ( .A(n45254), .B(n45255), .Z(n45253) );
  NANDN U45589 ( .A(n45256), .B(n45257), .Z(n45255) );
  NANDN U45590 ( .A(n45257), .B(n45256), .Z(n45252) );
  ANDN U45591 ( .B(B[109]), .A(n64), .Z(n45036) );
  XNOR U45592 ( .A(n45044), .B(n45258), .Z(n45037) );
  XNOR U45593 ( .A(n45043), .B(n45041), .Z(n45258) );
  AND U45594 ( .A(n45259), .B(n45260), .Z(n45041) );
  NANDN U45595 ( .A(n45261), .B(n45262), .Z(n45260) );
  OR U45596 ( .A(n45263), .B(n45264), .Z(n45262) );
  NAND U45597 ( .A(n45264), .B(n45263), .Z(n45259) );
  ANDN U45598 ( .B(B[110]), .A(n65), .Z(n45043) );
  XNOR U45599 ( .A(n45051), .B(n45265), .Z(n45044) );
  XNOR U45600 ( .A(n45050), .B(n45048), .Z(n45265) );
  AND U45601 ( .A(n45266), .B(n45267), .Z(n45048) );
  NANDN U45602 ( .A(n45268), .B(n45269), .Z(n45267) );
  NANDN U45603 ( .A(n45270), .B(n45271), .Z(n45269) );
  NANDN U45604 ( .A(n45271), .B(n45270), .Z(n45266) );
  ANDN U45605 ( .B(B[111]), .A(n66), .Z(n45050) );
  XNOR U45606 ( .A(n45058), .B(n45272), .Z(n45051) );
  XNOR U45607 ( .A(n45057), .B(n45055), .Z(n45272) );
  AND U45608 ( .A(n45273), .B(n45274), .Z(n45055) );
  NANDN U45609 ( .A(n45275), .B(n45276), .Z(n45274) );
  OR U45610 ( .A(n45277), .B(n45278), .Z(n45276) );
  NAND U45611 ( .A(n45278), .B(n45277), .Z(n45273) );
  ANDN U45612 ( .B(B[112]), .A(n67), .Z(n45057) );
  XNOR U45613 ( .A(n45065), .B(n45279), .Z(n45058) );
  XNOR U45614 ( .A(n45064), .B(n45062), .Z(n45279) );
  AND U45615 ( .A(n45280), .B(n45281), .Z(n45062) );
  NANDN U45616 ( .A(n45282), .B(n45283), .Z(n45281) );
  NANDN U45617 ( .A(n45284), .B(n45285), .Z(n45283) );
  NANDN U45618 ( .A(n45285), .B(n45284), .Z(n45280) );
  ANDN U45619 ( .B(B[113]), .A(n68), .Z(n45064) );
  XNOR U45620 ( .A(n45072), .B(n45286), .Z(n45065) );
  XNOR U45621 ( .A(n45071), .B(n45069), .Z(n45286) );
  AND U45622 ( .A(n45287), .B(n45288), .Z(n45069) );
  NANDN U45623 ( .A(n45289), .B(n45290), .Z(n45288) );
  OR U45624 ( .A(n45291), .B(n45292), .Z(n45290) );
  NAND U45625 ( .A(n45292), .B(n45291), .Z(n45287) );
  ANDN U45626 ( .B(B[114]), .A(n69), .Z(n45071) );
  XNOR U45627 ( .A(n45079), .B(n45293), .Z(n45072) );
  XNOR U45628 ( .A(n45078), .B(n45076), .Z(n45293) );
  AND U45629 ( .A(n45294), .B(n45295), .Z(n45076) );
  NANDN U45630 ( .A(n45296), .B(n45297), .Z(n45295) );
  NANDN U45631 ( .A(n45298), .B(n45299), .Z(n45297) );
  NANDN U45632 ( .A(n45299), .B(n45298), .Z(n45294) );
  ANDN U45633 ( .B(B[115]), .A(n70), .Z(n45078) );
  XNOR U45634 ( .A(n45086), .B(n45300), .Z(n45079) );
  XNOR U45635 ( .A(n45085), .B(n45083), .Z(n45300) );
  AND U45636 ( .A(n45301), .B(n45302), .Z(n45083) );
  NANDN U45637 ( .A(n45303), .B(n45304), .Z(n45302) );
  OR U45638 ( .A(n45305), .B(n45306), .Z(n45304) );
  NAND U45639 ( .A(n45306), .B(n45305), .Z(n45301) );
  ANDN U45640 ( .B(B[116]), .A(n71), .Z(n45085) );
  XNOR U45641 ( .A(n45093), .B(n45307), .Z(n45086) );
  XNOR U45642 ( .A(n45092), .B(n45090), .Z(n45307) );
  AND U45643 ( .A(n45308), .B(n45309), .Z(n45090) );
  NANDN U45644 ( .A(n45310), .B(n45311), .Z(n45309) );
  NANDN U45645 ( .A(n45312), .B(n45313), .Z(n45311) );
  NANDN U45646 ( .A(n45313), .B(n45312), .Z(n45308) );
  ANDN U45647 ( .B(B[117]), .A(n72), .Z(n45092) );
  XNOR U45648 ( .A(n45100), .B(n45314), .Z(n45093) );
  XNOR U45649 ( .A(n45099), .B(n45097), .Z(n45314) );
  AND U45650 ( .A(n45315), .B(n45316), .Z(n45097) );
  NANDN U45651 ( .A(n45317), .B(n45318), .Z(n45316) );
  OR U45652 ( .A(n45319), .B(n45320), .Z(n45318) );
  NAND U45653 ( .A(n45320), .B(n45319), .Z(n45315) );
  ANDN U45654 ( .B(B[118]), .A(n73), .Z(n45099) );
  XNOR U45655 ( .A(n45107), .B(n45321), .Z(n45100) );
  XNOR U45656 ( .A(n45106), .B(n45104), .Z(n45321) );
  AND U45657 ( .A(n45322), .B(n45323), .Z(n45104) );
  NANDN U45658 ( .A(n45324), .B(n45325), .Z(n45323) );
  NANDN U45659 ( .A(n45326), .B(n45327), .Z(n45325) );
  NANDN U45660 ( .A(n45327), .B(n45326), .Z(n45322) );
  ANDN U45661 ( .B(B[119]), .A(n74), .Z(n45106) );
  XNOR U45662 ( .A(n45114), .B(n45328), .Z(n45107) );
  XNOR U45663 ( .A(n45113), .B(n45111), .Z(n45328) );
  AND U45664 ( .A(n45329), .B(n45330), .Z(n45111) );
  NANDN U45665 ( .A(n45331), .B(n45332), .Z(n45330) );
  OR U45666 ( .A(n45333), .B(n45334), .Z(n45332) );
  NAND U45667 ( .A(n45334), .B(n45333), .Z(n45329) );
  ANDN U45668 ( .B(B[120]), .A(n75), .Z(n45113) );
  XNOR U45669 ( .A(n45121), .B(n45335), .Z(n45114) );
  XNOR U45670 ( .A(n45120), .B(n45118), .Z(n45335) );
  AND U45671 ( .A(n45336), .B(n45337), .Z(n45118) );
  NANDN U45672 ( .A(n45338), .B(n45339), .Z(n45337) );
  NANDN U45673 ( .A(n45340), .B(n45341), .Z(n45339) );
  NANDN U45674 ( .A(n45341), .B(n45340), .Z(n45336) );
  ANDN U45675 ( .B(B[121]), .A(n76), .Z(n45120) );
  XNOR U45676 ( .A(n45128), .B(n45342), .Z(n45121) );
  XNOR U45677 ( .A(n45127), .B(n45125), .Z(n45342) );
  AND U45678 ( .A(n45343), .B(n45344), .Z(n45125) );
  NANDN U45679 ( .A(n45345), .B(n45346), .Z(n45344) );
  OR U45680 ( .A(n45347), .B(n45348), .Z(n45346) );
  NAND U45681 ( .A(n45348), .B(n45347), .Z(n45343) );
  ANDN U45682 ( .B(B[122]), .A(n77), .Z(n45127) );
  XNOR U45683 ( .A(n45135), .B(n45349), .Z(n45128) );
  XNOR U45684 ( .A(n45134), .B(n45132), .Z(n45349) );
  AND U45685 ( .A(n45350), .B(n45351), .Z(n45132) );
  NANDN U45686 ( .A(n45352), .B(n45353), .Z(n45351) );
  NANDN U45687 ( .A(n45354), .B(n45355), .Z(n45353) );
  NANDN U45688 ( .A(n45355), .B(n45354), .Z(n45350) );
  ANDN U45689 ( .B(B[123]), .A(n78), .Z(n45134) );
  XNOR U45690 ( .A(n45142), .B(n45356), .Z(n45135) );
  XNOR U45691 ( .A(n45141), .B(n45139), .Z(n45356) );
  AND U45692 ( .A(n45357), .B(n45358), .Z(n45139) );
  NANDN U45693 ( .A(n45359), .B(n45360), .Z(n45358) );
  OR U45694 ( .A(n45361), .B(n45362), .Z(n45360) );
  NAND U45695 ( .A(n45362), .B(n45361), .Z(n45357) );
  ANDN U45696 ( .B(B[124]), .A(n79), .Z(n45141) );
  XNOR U45697 ( .A(n45149), .B(n45363), .Z(n45142) );
  XNOR U45698 ( .A(n45148), .B(n45146), .Z(n45363) );
  AND U45699 ( .A(n45364), .B(n45365), .Z(n45146) );
  NANDN U45700 ( .A(n45366), .B(n45367), .Z(n45365) );
  NANDN U45701 ( .A(n45368), .B(n45369), .Z(n45367) );
  NANDN U45702 ( .A(n45369), .B(n45368), .Z(n45364) );
  ANDN U45703 ( .B(B[125]), .A(n80), .Z(n45148) );
  XNOR U45704 ( .A(n45156), .B(n45370), .Z(n45149) );
  XNOR U45705 ( .A(n45155), .B(n45153), .Z(n45370) );
  AND U45706 ( .A(n45371), .B(n45372), .Z(n45153) );
  NANDN U45707 ( .A(n45373), .B(n45374), .Z(n45372) );
  OR U45708 ( .A(n45375), .B(n45376), .Z(n45374) );
  NAND U45709 ( .A(n45376), .B(n45375), .Z(n45371) );
  ANDN U45710 ( .B(B[126]), .A(n81), .Z(n45155) );
  XNOR U45711 ( .A(n45163), .B(n45377), .Z(n45156) );
  XNOR U45712 ( .A(n45162), .B(n45160), .Z(n45377) );
  AND U45713 ( .A(n45378), .B(n45379), .Z(n45160) );
  NANDN U45714 ( .A(n45380), .B(n45381), .Z(n45379) );
  NAND U45715 ( .A(n45382), .B(n45383), .Z(n45381) );
  ANDN U45716 ( .B(B[127]), .A(n82), .Z(n45162) );
  XOR U45717 ( .A(n45169), .B(n45384), .Z(n45163) );
  XNOR U45718 ( .A(n45167), .B(n45170), .Z(n45384) );
  NAND U45719 ( .A(A[2]), .B(B[128]), .Z(n45170) );
  NANDN U45720 ( .A(n45385), .B(n45386), .Z(n45167) );
  AND U45721 ( .A(A[0]), .B(B[129]), .Z(n45386) );
  XNOR U45722 ( .A(n45172), .B(n45387), .Z(n45169) );
  NAND U45723 ( .A(A[0]), .B(B[130]), .Z(n45387) );
  NAND U45724 ( .A(B[129]), .B(A[1]), .Z(n45172) );
  NAND U45725 ( .A(n45388), .B(n45389), .Z(n536) );
  NANDN U45726 ( .A(n45390), .B(n45391), .Z(n45389) );
  OR U45727 ( .A(n45392), .B(n45393), .Z(n45391) );
  NAND U45728 ( .A(n45393), .B(n45392), .Z(n45388) );
  XOR U45729 ( .A(n538), .B(n537), .Z(\A1[127] ) );
  XOR U45730 ( .A(n45393), .B(n45394), .Z(n537) );
  XNOR U45731 ( .A(n45392), .B(n45390), .Z(n45394) );
  AND U45732 ( .A(n45395), .B(n45396), .Z(n45390) );
  NANDN U45733 ( .A(n45397), .B(n45398), .Z(n45396) );
  NANDN U45734 ( .A(n45399), .B(n45400), .Z(n45398) );
  NANDN U45735 ( .A(n45400), .B(n45399), .Z(n45395) );
  ANDN U45736 ( .B(B[98]), .A(n54), .Z(n45392) );
  XNOR U45737 ( .A(n45187), .B(n45401), .Z(n45393) );
  XNOR U45738 ( .A(n45186), .B(n45184), .Z(n45401) );
  AND U45739 ( .A(n45402), .B(n45403), .Z(n45184) );
  NANDN U45740 ( .A(n45404), .B(n45405), .Z(n45403) );
  OR U45741 ( .A(n45406), .B(n45407), .Z(n45405) );
  NAND U45742 ( .A(n45407), .B(n45406), .Z(n45402) );
  ANDN U45743 ( .B(A[30]), .A(n6), .Z(n45186) );
  XNOR U45744 ( .A(n45194), .B(n45408), .Z(n45187) );
  XNOR U45745 ( .A(n45193), .B(n45191), .Z(n45408) );
  AND U45746 ( .A(n45409), .B(n45410), .Z(n45191) );
  NANDN U45747 ( .A(n45411), .B(n45412), .Z(n45410) );
  NANDN U45748 ( .A(n45413), .B(n45414), .Z(n45412) );
  NANDN U45749 ( .A(n45414), .B(n45413), .Z(n45409) );
  ANDN U45750 ( .B(A[29]), .A(n4), .Z(n45193) );
  XNOR U45751 ( .A(n45201), .B(n45415), .Z(n45194) );
  XNOR U45752 ( .A(n45200), .B(n45198), .Z(n45415) );
  AND U45753 ( .A(n45416), .B(n45417), .Z(n45198) );
  NANDN U45754 ( .A(n45418), .B(n45419), .Z(n45417) );
  OR U45755 ( .A(n45420), .B(n45421), .Z(n45419) );
  NAND U45756 ( .A(n45421), .B(n45420), .Z(n45416) );
  ANDN U45757 ( .B(B[101]), .A(n57), .Z(n45200) );
  XNOR U45758 ( .A(n45208), .B(n45422), .Z(n45201) );
  XNOR U45759 ( .A(n45207), .B(n45205), .Z(n45422) );
  AND U45760 ( .A(n45423), .B(n45424), .Z(n45205) );
  NANDN U45761 ( .A(n45425), .B(n45426), .Z(n45424) );
  NANDN U45762 ( .A(n45427), .B(n45428), .Z(n45426) );
  NANDN U45763 ( .A(n45428), .B(n45427), .Z(n45423) );
  ANDN U45764 ( .B(B[102]), .A(n58), .Z(n45207) );
  XNOR U45765 ( .A(n45215), .B(n45429), .Z(n45208) );
  XNOR U45766 ( .A(n45214), .B(n45212), .Z(n45429) );
  AND U45767 ( .A(n45430), .B(n45431), .Z(n45212) );
  NANDN U45768 ( .A(n45432), .B(n45433), .Z(n45431) );
  OR U45769 ( .A(n45434), .B(n45435), .Z(n45433) );
  NAND U45770 ( .A(n45435), .B(n45434), .Z(n45430) );
  ANDN U45771 ( .B(B[103]), .A(n59), .Z(n45214) );
  XNOR U45772 ( .A(n45222), .B(n45436), .Z(n45215) );
  XNOR U45773 ( .A(n45221), .B(n45219), .Z(n45436) );
  AND U45774 ( .A(n45437), .B(n45438), .Z(n45219) );
  NANDN U45775 ( .A(n45439), .B(n45440), .Z(n45438) );
  NANDN U45776 ( .A(n45441), .B(n45442), .Z(n45440) );
  NANDN U45777 ( .A(n45442), .B(n45441), .Z(n45437) );
  ANDN U45778 ( .B(B[104]), .A(n60), .Z(n45221) );
  XNOR U45779 ( .A(n45229), .B(n45443), .Z(n45222) );
  XNOR U45780 ( .A(n45228), .B(n45226), .Z(n45443) );
  AND U45781 ( .A(n45444), .B(n45445), .Z(n45226) );
  NANDN U45782 ( .A(n45446), .B(n45447), .Z(n45445) );
  OR U45783 ( .A(n45448), .B(n45449), .Z(n45447) );
  NAND U45784 ( .A(n45449), .B(n45448), .Z(n45444) );
  ANDN U45785 ( .B(B[105]), .A(n61), .Z(n45228) );
  XNOR U45786 ( .A(n45236), .B(n45450), .Z(n45229) );
  XNOR U45787 ( .A(n45235), .B(n45233), .Z(n45450) );
  AND U45788 ( .A(n45451), .B(n45452), .Z(n45233) );
  NANDN U45789 ( .A(n45453), .B(n45454), .Z(n45452) );
  NANDN U45790 ( .A(n45455), .B(n45456), .Z(n45454) );
  NANDN U45791 ( .A(n45456), .B(n45455), .Z(n45451) );
  ANDN U45792 ( .B(B[106]), .A(n62), .Z(n45235) );
  XNOR U45793 ( .A(n45243), .B(n45457), .Z(n45236) );
  XNOR U45794 ( .A(n45242), .B(n45240), .Z(n45457) );
  AND U45795 ( .A(n45458), .B(n45459), .Z(n45240) );
  NANDN U45796 ( .A(n45460), .B(n45461), .Z(n45459) );
  OR U45797 ( .A(n45462), .B(n45463), .Z(n45461) );
  NAND U45798 ( .A(n45463), .B(n45462), .Z(n45458) );
  ANDN U45799 ( .B(B[107]), .A(n63), .Z(n45242) );
  XNOR U45800 ( .A(n45250), .B(n45464), .Z(n45243) );
  XNOR U45801 ( .A(n45249), .B(n45247), .Z(n45464) );
  AND U45802 ( .A(n45465), .B(n45466), .Z(n45247) );
  NANDN U45803 ( .A(n45467), .B(n45468), .Z(n45466) );
  NANDN U45804 ( .A(n45469), .B(n45470), .Z(n45468) );
  NANDN U45805 ( .A(n45470), .B(n45469), .Z(n45465) );
  ANDN U45806 ( .B(B[108]), .A(n64), .Z(n45249) );
  XNOR U45807 ( .A(n45257), .B(n45471), .Z(n45250) );
  XNOR U45808 ( .A(n45256), .B(n45254), .Z(n45471) );
  AND U45809 ( .A(n45472), .B(n45473), .Z(n45254) );
  NANDN U45810 ( .A(n45474), .B(n45475), .Z(n45473) );
  OR U45811 ( .A(n45476), .B(n45477), .Z(n45475) );
  NAND U45812 ( .A(n45477), .B(n45476), .Z(n45472) );
  ANDN U45813 ( .B(B[109]), .A(n65), .Z(n45256) );
  XNOR U45814 ( .A(n45264), .B(n45478), .Z(n45257) );
  XNOR U45815 ( .A(n45263), .B(n45261), .Z(n45478) );
  AND U45816 ( .A(n45479), .B(n45480), .Z(n45261) );
  NANDN U45817 ( .A(n45481), .B(n45482), .Z(n45480) );
  NANDN U45818 ( .A(n45483), .B(n45484), .Z(n45482) );
  NANDN U45819 ( .A(n45484), .B(n45483), .Z(n45479) );
  ANDN U45820 ( .B(B[110]), .A(n66), .Z(n45263) );
  XNOR U45821 ( .A(n45271), .B(n45485), .Z(n45264) );
  XNOR U45822 ( .A(n45270), .B(n45268), .Z(n45485) );
  AND U45823 ( .A(n45486), .B(n45487), .Z(n45268) );
  NANDN U45824 ( .A(n45488), .B(n45489), .Z(n45487) );
  OR U45825 ( .A(n45490), .B(n45491), .Z(n45489) );
  NAND U45826 ( .A(n45491), .B(n45490), .Z(n45486) );
  ANDN U45827 ( .B(B[111]), .A(n67), .Z(n45270) );
  XNOR U45828 ( .A(n45278), .B(n45492), .Z(n45271) );
  XNOR U45829 ( .A(n45277), .B(n45275), .Z(n45492) );
  AND U45830 ( .A(n45493), .B(n45494), .Z(n45275) );
  NANDN U45831 ( .A(n45495), .B(n45496), .Z(n45494) );
  NANDN U45832 ( .A(n45497), .B(n45498), .Z(n45496) );
  NANDN U45833 ( .A(n45498), .B(n45497), .Z(n45493) );
  ANDN U45834 ( .B(B[112]), .A(n68), .Z(n45277) );
  XNOR U45835 ( .A(n45285), .B(n45499), .Z(n45278) );
  XNOR U45836 ( .A(n45284), .B(n45282), .Z(n45499) );
  AND U45837 ( .A(n45500), .B(n45501), .Z(n45282) );
  NANDN U45838 ( .A(n45502), .B(n45503), .Z(n45501) );
  OR U45839 ( .A(n45504), .B(n45505), .Z(n45503) );
  NAND U45840 ( .A(n45505), .B(n45504), .Z(n45500) );
  ANDN U45841 ( .B(B[113]), .A(n69), .Z(n45284) );
  XNOR U45842 ( .A(n45292), .B(n45506), .Z(n45285) );
  XNOR U45843 ( .A(n45291), .B(n45289), .Z(n45506) );
  AND U45844 ( .A(n45507), .B(n45508), .Z(n45289) );
  NANDN U45845 ( .A(n45509), .B(n45510), .Z(n45508) );
  NANDN U45846 ( .A(n45511), .B(n45512), .Z(n45510) );
  NANDN U45847 ( .A(n45512), .B(n45511), .Z(n45507) );
  ANDN U45848 ( .B(B[114]), .A(n70), .Z(n45291) );
  XNOR U45849 ( .A(n45299), .B(n45513), .Z(n45292) );
  XNOR U45850 ( .A(n45298), .B(n45296), .Z(n45513) );
  AND U45851 ( .A(n45514), .B(n45515), .Z(n45296) );
  NANDN U45852 ( .A(n45516), .B(n45517), .Z(n45515) );
  OR U45853 ( .A(n45518), .B(n45519), .Z(n45517) );
  NAND U45854 ( .A(n45519), .B(n45518), .Z(n45514) );
  ANDN U45855 ( .B(B[115]), .A(n71), .Z(n45298) );
  XNOR U45856 ( .A(n45306), .B(n45520), .Z(n45299) );
  XNOR U45857 ( .A(n45305), .B(n45303), .Z(n45520) );
  AND U45858 ( .A(n45521), .B(n45522), .Z(n45303) );
  NANDN U45859 ( .A(n45523), .B(n45524), .Z(n45522) );
  NANDN U45860 ( .A(n45525), .B(n45526), .Z(n45524) );
  NANDN U45861 ( .A(n45526), .B(n45525), .Z(n45521) );
  ANDN U45862 ( .B(B[116]), .A(n72), .Z(n45305) );
  XNOR U45863 ( .A(n45313), .B(n45527), .Z(n45306) );
  XNOR U45864 ( .A(n45312), .B(n45310), .Z(n45527) );
  AND U45865 ( .A(n45528), .B(n45529), .Z(n45310) );
  NANDN U45866 ( .A(n45530), .B(n45531), .Z(n45529) );
  OR U45867 ( .A(n45532), .B(n45533), .Z(n45531) );
  NAND U45868 ( .A(n45533), .B(n45532), .Z(n45528) );
  ANDN U45869 ( .B(B[117]), .A(n73), .Z(n45312) );
  XNOR U45870 ( .A(n45320), .B(n45534), .Z(n45313) );
  XNOR U45871 ( .A(n45319), .B(n45317), .Z(n45534) );
  AND U45872 ( .A(n45535), .B(n45536), .Z(n45317) );
  NANDN U45873 ( .A(n45537), .B(n45538), .Z(n45536) );
  NANDN U45874 ( .A(n45539), .B(n45540), .Z(n45538) );
  NANDN U45875 ( .A(n45540), .B(n45539), .Z(n45535) );
  ANDN U45876 ( .B(B[118]), .A(n74), .Z(n45319) );
  XNOR U45877 ( .A(n45327), .B(n45541), .Z(n45320) );
  XNOR U45878 ( .A(n45326), .B(n45324), .Z(n45541) );
  AND U45879 ( .A(n45542), .B(n45543), .Z(n45324) );
  NANDN U45880 ( .A(n45544), .B(n45545), .Z(n45543) );
  OR U45881 ( .A(n45546), .B(n45547), .Z(n45545) );
  NAND U45882 ( .A(n45547), .B(n45546), .Z(n45542) );
  ANDN U45883 ( .B(B[119]), .A(n75), .Z(n45326) );
  XNOR U45884 ( .A(n45334), .B(n45548), .Z(n45327) );
  XNOR U45885 ( .A(n45333), .B(n45331), .Z(n45548) );
  AND U45886 ( .A(n45549), .B(n45550), .Z(n45331) );
  NANDN U45887 ( .A(n45551), .B(n45552), .Z(n45550) );
  NANDN U45888 ( .A(n45553), .B(n45554), .Z(n45552) );
  NANDN U45889 ( .A(n45554), .B(n45553), .Z(n45549) );
  ANDN U45890 ( .B(B[120]), .A(n76), .Z(n45333) );
  XNOR U45891 ( .A(n45341), .B(n45555), .Z(n45334) );
  XNOR U45892 ( .A(n45340), .B(n45338), .Z(n45555) );
  AND U45893 ( .A(n45556), .B(n45557), .Z(n45338) );
  NANDN U45894 ( .A(n45558), .B(n45559), .Z(n45557) );
  OR U45895 ( .A(n45560), .B(n45561), .Z(n45559) );
  NAND U45896 ( .A(n45561), .B(n45560), .Z(n45556) );
  ANDN U45897 ( .B(B[121]), .A(n77), .Z(n45340) );
  XNOR U45898 ( .A(n45348), .B(n45562), .Z(n45341) );
  XNOR U45899 ( .A(n45347), .B(n45345), .Z(n45562) );
  AND U45900 ( .A(n45563), .B(n45564), .Z(n45345) );
  NANDN U45901 ( .A(n45565), .B(n45566), .Z(n45564) );
  NANDN U45902 ( .A(n45567), .B(n45568), .Z(n45566) );
  NANDN U45903 ( .A(n45568), .B(n45567), .Z(n45563) );
  ANDN U45904 ( .B(B[122]), .A(n78), .Z(n45347) );
  XNOR U45905 ( .A(n45355), .B(n45569), .Z(n45348) );
  XNOR U45906 ( .A(n45354), .B(n45352), .Z(n45569) );
  AND U45907 ( .A(n45570), .B(n45571), .Z(n45352) );
  NANDN U45908 ( .A(n45572), .B(n45573), .Z(n45571) );
  OR U45909 ( .A(n45574), .B(n45575), .Z(n45573) );
  NAND U45910 ( .A(n45575), .B(n45574), .Z(n45570) );
  ANDN U45911 ( .B(B[123]), .A(n79), .Z(n45354) );
  XNOR U45912 ( .A(n45362), .B(n45576), .Z(n45355) );
  XNOR U45913 ( .A(n45361), .B(n45359), .Z(n45576) );
  AND U45914 ( .A(n45577), .B(n45578), .Z(n45359) );
  NANDN U45915 ( .A(n45579), .B(n45580), .Z(n45578) );
  NANDN U45916 ( .A(n45581), .B(n45582), .Z(n45580) );
  NANDN U45917 ( .A(n45582), .B(n45581), .Z(n45577) );
  ANDN U45918 ( .B(B[124]), .A(n80), .Z(n45361) );
  XNOR U45919 ( .A(n45369), .B(n45583), .Z(n45362) );
  XNOR U45920 ( .A(n45368), .B(n45366), .Z(n45583) );
  AND U45921 ( .A(n45584), .B(n45585), .Z(n45366) );
  NANDN U45922 ( .A(n45586), .B(n45587), .Z(n45585) );
  OR U45923 ( .A(n45588), .B(n45589), .Z(n45587) );
  NAND U45924 ( .A(n45589), .B(n45588), .Z(n45584) );
  ANDN U45925 ( .B(B[125]), .A(n81), .Z(n45368) );
  XNOR U45926 ( .A(n45376), .B(n45590), .Z(n45369) );
  XNOR U45927 ( .A(n45375), .B(n45373), .Z(n45590) );
  AND U45928 ( .A(n45591), .B(n45592), .Z(n45373) );
  NANDN U45929 ( .A(n45593), .B(n45594), .Z(n45592) );
  NAND U45930 ( .A(n45595), .B(n45596), .Z(n45594) );
  ANDN U45931 ( .B(B[126]), .A(n82), .Z(n45375) );
  XOR U45932 ( .A(n45382), .B(n45597), .Z(n45376) );
  XNOR U45933 ( .A(n45380), .B(n45383), .Z(n45597) );
  NAND U45934 ( .A(A[2]), .B(B[127]), .Z(n45383) );
  NANDN U45935 ( .A(n45598), .B(n45599), .Z(n45380) );
  AND U45936 ( .A(A[0]), .B(B[128]), .Z(n45599) );
  XNOR U45937 ( .A(n45385), .B(n45600), .Z(n45382) );
  NAND U45938 ( .A(A[0]), .B(B[129]), .Z(n45600) );
  NAND U45939 ( .A(B[128]), .B(A[1]), .Z(n45385) );
  NAND U45940 ( .A(n45601), .B(n45602), .Z(n538) );
  NANDN U45941 ( .A(n45603), .B(n45604), .Z(n45602) );
  OR U45942 ( .A(n45605), .B(n45606), .Z(n45604) );
  NAND U45943 ( .A(n45606), .B(n45605), .Z(n45601) );
  XOR U45944 ( .A(n540), .B(n539), .Z(\A1[126] ) );
  XOR U45945 ( .A(n45606), .B(n45607), .Z(n539) );
  XNOR U45946 ( .A(n45605), .B(n45603), .Z(n45607) );
  AND U45947 ( .A(n45608), .B(n45609), .Z(n45603) );
  NANDN U45948 ( .A(n45610), .B(n45611), .Z(n45609) );
  NANDN U45949 ( .A(n45612), .B(n45613), .Z(n45611) );
  NANDN U45950 ( .A(n45613), .B(n45612), .Z(n45608) );
  ANDN U45951 ( .B(B[97]), .A(n54), .Z(n45605) );
  XNOR U45952 ( .A(n45400), .B(n45614), .Z(n45606) );
  XNOR U45953 ( .A(n45399), .B(n45397), .Z(n45614) );
  AND U45954 ( .A(n45615), .B(n45616), .Z(n45397) );
  NANDN U45955 ( .A(n45617), .B(n45618), .Z(n45616) );
  OR U45956 ( .A(n45619), .B(n45620), .Z(n45618) );
  NAND U45957 ( .A(n45620), .B(n45619), .Z(n45615) );
  ANDN U45958 ( .B(B[98]), .A(n55), .Z(n45399) );
  XNOR U45959 ( .A(n45407), .B(n45621), .Z(n45400) );
  XNOR U45960 ( .A(n45406), .B(n45404), .Z(n45621) );
  AND U45961 ( .A(n45622), .B(n45623), .Z(n45404) );
  NANDN U45962 ( .A(n45624), .B(n45625), .Z(n45623) );
  NANDN U45963 ( .A(n45626), .B(n45627), .Z(n45625) );
  NANDN U45964 ( .A(n45627), .B(n45626), .Z(n45622) );
  ANDN U45965 ( .B(A[29]), .A(n6), .Z(n45406) );
  XNOR U45966 ( .A(n45414), .B(n45628), .Z(n45407) );
  XNOR U45967 ( .A(n45413), .B(n45411), .Z(n45628) );
  AND U45968 ( .A(n45629), .B(n45630), .Z(n45411) );
  NANDN U45969 ( .A(n45631), .B(n45632), .Z(n45630) );
  OR U45970 ( .A(n45633), .B(n45634), .Z(n45632) );
  NAND U45971 ( .A(n45634), .B(n45633), .Z(n45629) );
  ANDN U45972 ( .B(A[28]), .A(n4), .Z(n45413) );
  XNOR U45973 ( .A(n45421), .B(n45635), .Z(n45414) );
  XNOR U45974 ( .A(n45420), .B(n45418), .Z(n45635) );
  AND U45975 ( .A(n45636), .B(n45637), .Z(n45418) );
  NANDN U45976 ( .A(n45638), .B(n45639), .Z(n45637) );
  NANDN U45977 ( .A(n45640), .B(n45641), .Z(n45639) );
  NANDN U45978 ( .A(n45641), .B(n45640), .Z(n45636) );
  ANDN U45979 ( .B(B[101]), .A(n58), .Z(n45420) );
  XNOR U45980 ( .A(n45428), .B(n45642), .Z(n45421) );
  XNOR U45981 ( .A(n45427), .B(n45425), .Z(n45642) );
  AND U45982 ( .A(n45643), .B(n45644), .Z(n45425) );
  NANDN U45983 ( .A(n45645), .B(n45646), .Z(n45644) );
  OR U45984 ( .A(n45647), .B(n45648), .Z(n45646) );
  NAND U45985 ( .A(n45648), .B(n45647), .Z(n45643) );
  ANDN U45986 ( .B(B[102]), .A(n59), .Z(n45427) );
  XNOR U45987 ( .A(n45435), .B(n45649), .Z(n45428) );
  XNOR U45988 ( .A(n45434), .B(n45432), .Z(n45649) );
  AND U45989 ( .A(n45650), .B(n45651), .Z(n45432) );
  NANDN U45990 ( .A(n45652), .B(n45653), .Z(n45651) );
  NANDN U45991 ( .A(n45654), .B(n45655), .Z(n45653) );
  NANDN U45992 ( .A(n45655), .B(n45654), .Z(n45650) );
  ANDN U45993 ( .B(B[103]), .A(n60), .Z(n45434) );
  XNOR U45994 ( .A(n45442), .B(n45656), .Z(n45435) );
  XNOR U45995 ( .A(n45441), .B(n45439), .Z(n45656) );
  AND U45996 ( .A(n45657), .B(n45658), .Z(n45439) );
  NANDN U45997 ( .A(n45659), .B(n45660), .Z(n45658) );
  OR U45998 ( .A(n45661), .B(n45662), .Z(n45660) );
  NAND U45999 ( .A(n45662), .B(n45661), .Z(n45657) );
  ANDN U46000 ( .B(B[104]), .A(n61), .Z(n45441) );
  XNOR U46001 ( .A(n45449), .B(n45663), .Z(n45442) );
  XNOR U46002 ( .A(n45448), .B(n45446), .Z(n45663) );
  AND U46003 ( .A(n45664), .B(n45665), .Z(n45446) );
  NANDN U46004 ( .A(n45666), .B(n45667), .Z(n45665) );
  NANDN U46005 ( .A(n45668), .B(n45669), .Z(n45667) );
  NANDN U46006 ( .A(n45669), .B(n45668), .Z(n45664) );
  ANDN U46007 ( .B(B[105]), .A(n62), .Z(n45448) );
  XNOR U46008 ( .A(n45456), .B(n45670), .Z(n45449) );
  XNOR U46009 ( .A(n45455), .B(n45453), .Z(n45670) );
  AND U46010 ( .A(n45671), .B(n45672), .Z(n45453) );
  NANDN U46011 ( .A(n45673), .B(n45674), .Z(n45672) );
  OR U46012 ( .A(n45675), .B(n45676), .Z(n45674) );
  NAND U46013 ( .A(n45676), .B(n45675), .Z(n45671) );
  ANDN U46014 ( .B(B[106]), .A(n63), .Z(n45455) );
  XNOR U46015 ( .A(n45463), .B(n45677), .Z(n45456) );
  XNOR U46016 ( .A(n45462), .B(n45460), .Z(n45677) );
  AND U46017 ( .A(n45678), .B(n45679), .Z(n45460) );
  NANDN U46018 ( .A(n45680), .B(n45681), .Z(n45679) );
  NANDN U46019 ( .A(n45682), .B(n45683), .Z(n45681) );
  NANDN U46020 ( .A(n45683), .B(n45682), .Z(n45678) );
  ANDN U46021 ( .B(B[107]), .A(n64), .Z(n45462) );
  XNOR U46022 ( .A(n45470), .B(n45684), .Z(n45463) );
  XNOR U46023 ( .A(n45469), .B(n45467), .Z(n45684) );
  AND U46024 ( .A(n45685), .B(n45686), .Z(n45467) );
  NANDN U46025 ( .A(n45687), .B(n45688), .Z(n45686) );
  OR U46026 ( .A(n45689), .B(n45690), .Z(n45688) );
  NAND U46027 ( .A(n45690), .B(n45689), .Z(n45685) );
  ANDN U46028 ( .B(B[108]), .A(n65), .Z(n45469) );
  XNOR U46029 ( .A(n45477), .B(n45691), .Z(n45470) );
  XNOR U46030 ( .A(n45476), .B(n45474), .Z(n45691) );
  AND U46031 ( .A(n45692), .B(n45693), .Z(n45474) );
  NANDN U46032 ( .A(n45694), .B(n45695), .Z(n45693) );
  NANDN U46033 ( .A(n45696), .B(n45697), .Z(n45695) );
  NANDN U46034 ( .A(n45697), .B(n45696), .Z(n45692) );
  ANDN U46035 ( .B(B[109]), .A(n66), .Z(n45476) );
  XNOR U46036 ( .A(n45484), .B(n45698), .Z(n45477) );
  XNOR U46037 ( .A(n45483), .B(n45481), .Z(n45698) );
  AND U46038 ( .A(n45699), .B(n45700), .Z(n45481) );
  NANDN U46039 ( .A(n45701), .B(n45702), .Z(n45700) );
  OR U46040 ( .A(n45703), .B(n45704), .Z(n45702) );
  NAND U46041 ( .A(n45704), .B(n45703), .Z(n45699) );
  ANDN U46042 ( .B(B[110]), .A(n67), .Z(n45483) );
  XNOR U46043 ( .A(n45491), .B(n45705), .Z(n45484) );
  XNOR U46044 ( .A(n45490), .B(n45488), .Z(n45705) );
  AND U46045 ( .A(n45706), .B(n45707), .Z(n45488) );
  NANDN U46046 ( .A(n45708), .B(n45709), .Z(n45707) );
  NANDN U46047 ( .A(n45710), .B(n45711), .Z(n45709) );
  NANDN U46048 ( .A(n45711), .B(n45710), .Z(n45706) );
  ANDN U46049 ( .B(B[111]), .A(n68), .Z(n45490) );
  XNOR U46050 ( .A(n45498), .B(n45712), .Z(n45491) );
  XNOR U46051 ( .A(n45497), .B(n45495), .Z(n45712) );
  AND U46052 ( .A(n45713), .B(n45714), .Z(n45495) );
  NANDN U46053 ( .A(n45715), .B(n45716), .Z(n45714) );
  OR U46054 ( .A(n45717), .B(n45718), .Z(n45716) );
  NAND U46055 ( .A(n45718), .B(n45717), .Z(n45713) );
  ANDN U46056 ( .B(B[112]), .A(n69), .Z(n45497) );
  XNOR U46057 ( .A(n45505), .B(n45719), .Z(n45498) );
  XNOR U46058 ( .A(n45504), .B(n45502), .Z(n45719) );
  AND U46059 ( .A(n45720), .B(n45721), .Z(n45502) );
  NANDN U46060 ( .A(n45722), .B(n45723), .Z(n45721) );
  NANDN U46061 ( .A(n45724), .B(n45725), .Z(n45723) );
  NANDN U46062 ( .A(n45725), .B(n45724), .Z(n45720) );
  ANDN U46063 ( .B(B[113]), .A(n70), .Z(n45504) );
  XNOR U46064 ( .A(n45512), .B(n45726), .Z(n45505) );
  XNOR U46065 ( .A(n45511), .B(n45509), .Z(n45726) );
  AND U46066 ( .A(n45727), .B(n45728), .Z(n45509) );
  NANDN U46067 ( .A(n45729), .B(n45730), .Z(n45728) );
  OR U46068 ( .A(n45731), .B(n45732), .Z(n45730) );
  NAND U46069 ( .A(n45732), .B(n45731), .Z(n45727) );
  ANDN U46070 ( .B(B[114]), .A(n71), .Z(n45511) );
  XNOR U46071 ( .A(n45519), .B(n45733), .Z(n45512) );
  XNOR U46072 ( .A(n45518), .B(n45516), .Z(n45733) );
  AND U46073 ( .A(n45734), .B(n45735), .Z(n45516) );
  NANDN U46074 ( .A(n45736), .B(n45737), .Z(n45735) );
  NANDN U46075 ( .A(n45738), .B(n45739), .Z(n45737) );
  NANDN U46076 ( .A(n45739), .B(n45738), .Z(n45734) );
  ANDN U46077 ( .B(B[115]), .A(n72), .Z(n45518) );
  XNOR U46078 ( .A(n45526), .B(n45740), .Z(n45519) );
  XNOR U46079 ( .A(n45525), .B(n45523), .Z(n45740) );
  AND U46080 ( .A(n45741), .B(n45742), .Z(n45523) );
  NANDN U46081 ( .A(n45743), .B(n45744), .Z(n45742) );
  OR U46082 ( .A(n45745), .B(n45746), .Z(n45744) );
  NAND U46083 ( .A(n45746), .B(n45745), .Z(n45741) );
  ANDN U46084 ( .B(B[116]), .A(n73), .Z(n45525) );
  XNOR U46085 ( .A(n45533), .B(n45747), .Z(n45526) );
  XNOR U46086 ( .A(n45532), .B(n45530), .Z(n45747) );
  AND U46087 ( .A(n45748), .B(n45749), .Z(n45530) );
  NANDN U46088 ( .A(n45750), .B(n45751), .Z(n45749) );
  NANDN U46089 ( .A(n45752), .B(n45753), .Z(n45751) );
  NANDN U46090 ( .A(n45753), .B(n45752), .Z(n45748) );
  ANDN U46091 ( .B(B[117]), .A(n74), .Z(n45532) );
  XNOR U46092 ( .A(n45540), .B(n45754), .Z(n45533) );
  XNOR U46093 ( .A(n45539), .B(n45537), .Z(n45754) );
  AND U46094 ( .A(n45755), .B(n45756), .Z(n45537) );
  NANDN U46095 ( .A(n45757), .B(n45758), .Z(n45756) );
  OR U46096 ( .A(n45759), .B(n45760), .Z(n45758) );
  NAND U46097 ( .A(n45760), .B(n45759), .Z(n45755) );
  ANDN U46098 ( .B(B[118]), .A(n75), .Z(n45539) );
  XNOR U46099 ( .A(n45547), .B(n45761), .Z(n45540) );
  XNOR U46100 ( .A(n45546), .B(n45544), .Z(n45761) );
  AND U46101 ( .A(n45762), .B(n45763), .Z(n45544) );
  NANDN U46102 ( .A(n45764), .B(n45765), .Z(n45763) );
  NANDN U46103 ( .A(n45766), .B(n45767), .Z(n45765) );
  NANDN U46104 ( .A(n45767), .B(n45766), .Z(n45762) );
  ANDN U46105 ( .B(B[119]), .A(n76), .Z(n45546) );
  XNOR U46106 ( .A(n45554), .B(n45768), .Z(n45547) );
  XNOR U46107 ( .A(n45553), .B(n45551), .Z(n45768) );
  AND U46108 ( .A(n45769), .B(n45770), .Z(n45551) );
  NANDN U46109 ( .A(n45771), .B(n45772), .Z(n45770) );
  OR U46110 ( .A(n45773), .B(n45774), .Z(n45772) );
  NAND U46111 ( .A(n45774), .B(n45773), .Z(n45769) );
  ANDN U46112 ( .B(B[120]), .A(n77), .Z(n45553) );
  XNOR U46113 ( .A(n45561), .B(n45775), .Z(n45554) );
  XNOR U46114 ( .A(n45560), .B(n45558), .Z(n45775) );
  AND U46115 ( .A(n45776), .B(n45777), .Z(n45558) );
  NANDN U46116 ( .A(n45778), .B(n45779), .Z(n45777) );
  NANDN U46117 ( .A(n45780), .B(n45781), .Z(n45779) );
  NANDN U46118 ( .A(n45781), .B(n45780), .Z(n45776) );
  ANDN U46119 ( .B(B[121]), .A(n78), .Z(n45560) );
  XNOR U46120 ( .A(n45568), .B(n45782), .Z(n45561) );
  XNOR U46121 ( .A(n45567), .B(n45565), .Z(n45782) );
  AND U46122 ( .A(n45783), .B(n45784), .Z(n45565) );
  NANDN U46123 ( .A(n45785), .B(n45786), .Z(n45784) );
  OR U46124 ( .A(n45787), .B(n45788), .Z(n45786) );
  NAND U46125 ( .A(n45788), .B(n45787), .Z(n45783) );
  ANDN U46126 ( .B(B[122]), .A(n79), .Z(n45567) );
  XNOR U46127 ( .A(n45575), .B(n45789), .Z(n45568) );
  XNOR U46128 ( .A(n45574), .B(n45572), .Z(n45789) );
  AND U46129 ( .A(n45790), .B(n45791), .Z(n45572) );
  NANDN U46130 ( .A(n45792), .B(n45793), .Z(n45791) );
  NANDN U46131 ( .A(n45794), .B(n45795), .Z(n45793) );
  NANDN U46132 ( .A(n45795), .B(n45794), .Z(n45790) );
  ANDN U46133 ( .B(B[123]), .A(n80), .Z(n45574) );
  XNOR U46134 ( .A(n45582), .B(n45796), .Z(n45575) );
  XNOR U46135 ( .A(n45581), .B(n45579), .Z(n45796) );
  AND U46136 ( .A(n45797), .B(n45798), .Z(n45579) );
  NANDN U46137 ( .A(n45799), .B(n45800), .Z(n45798) );
  OR U46138 ( .A(n45801), .B(n45802), .Z(n45800) );
  NAND U46139 ( .A(n45802), .B(n45801), .Z(n45797) );
  ANDN U46140 ( .B(B[124]), .A(n81), .Z(n45581) );
  XNOR U46141 ( .A(n45589), .B(n45803), .Z(n45582) );
  XNOR U46142 ( .A(n45588), .B(n45586), .Z(n45803) );
  AND U46143 ( .A(n45804), .B(n45805), .Z(n45586) );
  NANDN U46144 ( .A(n45806), .B(n45807), .Z(n45805) );
  NAND U46145 ( .A(n45808), .B(n45809), .Z(n45807) );
  ANDN U46146 ( .B(B[125]), .A(n82), .Z(n45588) );
  XOR U46147 ( .A(n45595), .B(n45810), .Z(n45589) );
  XNOR U46148 ( .A(n45593), .B(n45596), .Z(n45810) );
  NAND U46149 ( .A(A[2]), .B(B[126]), .Z(n45596) );
  NANDN U46150 ( .A(n45811), .B(n45812), .Z(n45593) );
  AND U46151 ( .A(A[0]), .B(B[127]), .Z(n45812) );
  XNOR U46152 ( .A(n45598), .B(n45813), .Z(n45595) );
  NAND U46153 ( .A(A[0]), .B(B[128]), .Z(n45813) );
  NAND U46154 ( .A(B[127]), .B(A[1]), .Z(n45598) );
  NAND U46155 ( .A(n45814), .B(n45815), .Z(n540) );
  NANDN U46156 ( .A(n45816), .B(n45817), .Z(n45815) );
  OR U46157 ( .A(n45818), .B(n45819), .Z(n45817) );
  NAND U46158 ( .A(n45819), .B(n45818), .Z(n45814) );
  XOR U46159 ( .A(n542), .B(n541), .Z(\A1[125] ) );
  XOR U46160 ( .A(n45819), .B(n45820), .Z(n541) );
  XNOR U46161 ( .A(n45818), .B(n45816), .Z(n45820) );
  AND U46162 ( .A(n45821), .B(n45822), .Z(n45816) );
  NANDN U46163 ( .A(n45823), .B(n45824), .Z(n45822) );
  NANDN U46164 ( .A(n45825), .B(n45826), .Z(n45824) );
  NANDN U46165 ( .A(n45826), .B(n45825), .Z(n45821) );
  ANDN U46166 ( .B(B[96]), .A(n54), .Z(n45818) );
  XNOR U46167 ( .A(n45613), .B(n45827), .Z(n45819) );
  XNOR U46168 ( .A(n45612), .B(n45610), .Z(n45827) );
  AND U46169 ( .A(n45828), .B(n45829), .Z(n45610) );
  NANDN U46170 ( .A(n45830), .B(n45831), .Z(n45829) );
  OR U46171 ( .A(n45832), .B(n45833), .Z(n45831) );
  NAND U46172 ( .A(n45833), .B(n45832), .Z(n45828) );
  ANDN U46173 ( .B(B[97]), .A(n55), .Z(n45612) );
  XNOR U46174 ( .A(n45620), .B(n45834), .Z(n45613) );
  XNOR U46175 ( .A(n45619), .B(n45617), .Z(n45834) );
  AND U46176 ( .A(n45835), .B(n45836), .Z(n45617) );
  NANDN U46177 ( .A(n45837), .B(n45838), .Z(n45836) );
  NANDN U46178 ( .A(n45839), .B(n45840), .Z(n45838) );
  NANDN U46179 ( .A(n45840), .B(n45839), .Z(n45835) );
  ANDN U46180 ( .B(B[98]), .A(n56), .Z(n45619) );
  XNOR U46181 ( .A(n45627), .B(n45841), .Z(n45620) );
  XNOR U46182 ( .A(n45626), .B(n45624), .Z(n45841) );
  AND U46183 ( .A(n45842), .B(n45843), .Z(n45624) );
  NANDN U46184 ( .A(n45844), .B(n45845), .Z(n45843) );
  OR U46185 ( .A(n45846), .B(n45847), .Z(n45845) );
  NAND U46186 ( .A(n45847), .B(n45846), .Z(n45842) );
  ANDN U46187 ( .B(A[28]), .A(n6), .Z(n45626) );
  XNOR U46188 ( .A(n45634), .B(n45848), .Z(n45627) );
  XNOR U46189 ( .A(n45633), .B(n45631), .Z(n45848) );
  AND U46190 ( .A(n45849), .B(n45850), .Z(n45631) );
  NANDN U46191 ( .A(n45851), .B(n45852), .Z(n45850) );
  NANDN U46192 ( .A(n45853), .B(n45854), .Z(n45852) );
  NANDN U46193 ( .A(n45854), .B(n45853), .Z(n45849) );
  ANDN U46194 ( .B(A[27]), .A(n4), .Z(n45633) );
  XNOR U46195 ( .A(n45641), .B(n45855), .Z(n45634) );
  XNOR U46196 ( .A(n45640), .B(n45638), .Z(n45855) );
  AND U46197 ( .A(n45856), .B(n45857), .Z(n45638) );
  NANDN U46198 ( .A(n45858), .B(n45859), .Z(n45857) );
  OR U46199 ( .A(n45860), .B(n45861), .Z(n45859) );
  NAND U46200 ( .A(n45861), .B(n45860), .Z(n45856) );
  ANDN U46201 ( .B(B[101]), .A(n59), .Z(n45640) );
  XNOR U46202 ( .A(n45648), .B(n45862), .Z(n45641) );
  XNOR U46203 ( .A(n45647), .B(n45645), .Z(n45862) );
  AND U46204 ( .A(n45863), .B(n45864), .Z(n45645) );
  NANDN U46205 ( .A(n45865), .B(n45866), .Z(n45864) );
  NANDN U46206 ( .A(n45867), .B(n45868), .Z(n45866) );
  NANDN U46207 ( .A(n45868), .B(n45867), .Z(n45863) );
  ANDN U46208 ( .B(B[102]), .A(n60), .Z(n45647) );
  XNOR U46209 ( .A(n45655), .B(n45869), .Z(n45648) );
  XNOR U46210 ( .A(n45654), .B(n45652), .Z(n45869) );
  AND U46211 ( .A(n45870), .B(n45871), .Z(n45652) );
  NANDN U46212 ( .A(n45872), .B(n45873), .Z(n45871) );
  OR U46213 ( .A(n45874), .B(n45875), .Z(n45873) );
  NAND U46214 ( .A(n45875), .B(n45874), .Z(n45870) );
  ANDN U46215 ( .B(B[103]), .A(n61), .Z(n45654) );
  XNOR U46216 ( .A(n45662), .B(n45876), .Z(n45655) );
  XNOR U46217 ( .A(n45661), .B(n45659), .Z(n45876) );
  AND U46218 ( .A(n45877), .B(n45878), .Z(n45659) );
  NANDN U46219 ( .A(n45879), .B(n45880), .Z(n45878) );
  NANDN U46220 ( .A(n45881), .B(n45882), .Z(n45880) );
  NANDN U46221 ( .A(n45882), .B(n45881), .Z(n45877) );
  ANDN U46222 ( .B(B[104]), .A(n62), .Z(n45661) );
  XNOR U46223 ( .A(n45669), .B(n45883), .Z(n45662) );
  XNOR U46224 ( .A(n45668), .B(n45666), .Z(n45883) );
  AND U46225 ( .A(n45884), .B(n45885), .Z(n45666) );
  NANDN U46226 ( .A(n45886), .B(n45887), .Z(n45885) );
  OR U46227 ( .A(n45888), .B(n45889), .Z(n45887) );
  NAND U46228 ( .A(n45889), .B(n45888), .Z(n45884) );
  ANDN U46229 ( .B(B[105]), .A(n63), .Z(n45668) );
  XNOR U46230 ( .A(n45676), .B(n45890), .Z(n45669) );
  XNOR U46231 ( .A(n45675), .B(n45673), .Z(n45890) );
  AND U46232 ( .A(n45891), .B(n45892), .Z(n45673) );
  NANDN U46233 ( .A(n45893), .B(n45894), .Z(n45892) );
  NANDN U46234 ( .A(n45895), .B(n45896), .Z(n45894) );
  NANDN U46235 ( .A(n45896), .B(n45895), .Z(n45891) );
  ANDN U46236 ( .B(B[106]), .A(n64), .Z(n45675) );
  XNOR U46237 ( .A(n45683), .B(n45897), .Z(n45676) );
  XNOR U46238 ( .A(n45682), .B(n45680), .Z(n45897) );
  AND U46239 ( .A(n45898), .B(n45899), .Z(n45680) );
  NANDN U46240 ( .A(n45900), .B(n45901), .Z(n45899) );
  OR U46241 ( .A(n45902), .B(n45903), .Z(n45901) );
  NAND U46242 ( .A(n45903), .B(n45902), .Z(n45898) );
  ANDN U46243 ( .B(B[107]), .A(n65), .Z(n45682) );
  XNOR U46244 ( .A(n45690), .B(n45904), .Z(n45683) );
  XNOR U46245 ( .A(n45689), .B(n45687), .Z(n45904) );
  AND U46246 ( .A(n45905), .B(n45906), .Z(n45687) );
  NANDN U46247 ( .A(n45907), .B(n45908), .Z(n45906) );
  NANDN U46248 ( .A(n45909), .B(n45910), .Z(n45908) );
  NANDN U46249 ( .A(n45910), .B(n45909), .Z(n45905) );
  ANDN U46250 ( .B(B[108]), .A(n66), .Z(n45689) );
  XNOR U46251 ( .A(n45697), .B(n45911), .Z(n45690) );
  XNOR U46252 ( .A(n45696), .B(n45694), .Z(n45911) );
  AND U46253 ( .A(n45912), .B(n45913), .Z(n45694) );
  NANDN U46254 ( .A(n45914), .B(n45915), .Z(n45913) );
  OR U46255 ( .A(n45916), .B(n45917), .Z(n45915) );
  NAND U46256 ( .A(n45917), .B(n45916), .Z(n45912) );
  ANDN U46257 ( .B(B[109]), .A(n67), .Z(n45696) );
  XNOR U46258 ( .A(n45704), .B(n45918), .Z(n45697) );
  XNOR U46259 ( .A(n45703), .B(n45701), .Z(n45918) );
  AND U46260 ( .A(n45919), .B(n45920), .Z(n45701) );
  NANDN U46261 ( .A(n45921), .B(n45922), .Z(n45920) );
  NANDN U46262 ( .A(n45923), .B(n45924), .Z(n45922) );
  NANDN U46263 ( .A(n45924), .B(n45923), .Z(n45919) );
  ANDN U46264 ( .B(B[110]), .A(n68), .Z(n45703) );
  XNOR U46265 ( .A(n45711), .B(n45925), .Z(n45704) );
  XNOR U46266 ( .A(n45710), .B(n45708), .Z(n45925) );
  AND U46267 ( .A(n45926), .B(n45927), .Z(n45708) );
  NANDN U46268 ( .A(n45928), .B(n45929), .Z(n45927) );
  OR U46269 ( .A(n45930), .B(n45931), .Z(n45929) );
  NAND U46270 ( .A(n45931), .B(n45930), .Z(n45926) );
  ANDN U46271 ( .B(B[111]), .A(n69), .Z(n45710) );
  XNOR U46272 ( .A(n45718), .B(n45932), .Z(n45711) );
  XNOR U46273 ( .A(n45717), .B(n45715), .Z(n45932) );
  AND U46274 ( .A(n45933), .B(n45934), .Z(n45715) );
  NANDN U46275 ( .A(n45935), .B(n45936), .Z(n45934) );
  NANDN U46276 ( .A(n45937), .B(n45938), .Z(n45936) );
  NANDN U46277 ( .A(n45938), .B(n45937), .Z(n45933) );
  ANDN U46278 ( .B(B[112]), .A(n70), .Z(n45717) );
  XNOR U46279 ( .A(n45725), .B(n45939), .Z(n45718) );
  XNOR U46280 ( .A(n45724), .B(n45722), .Z(n45939) );
  AND U46281 ( .A(n45940), .B(n45941), .Z(n45722) );
  NANDN U46282 ( .A(n45942), .B(n45943), .Z(n45941) );
  OR U46283 ( .A(n45944), .B(n45945), .Z(n45943) );
  NAND U46284 ( .A(n45945), .B(n45944), .Z(n45940) );
  ANDN U46285 ( .B(B[113]), .A(n71), .Z(n45724) );
  XNOR U46286 ( .A(n45732), .B(n45946), .Z(n45725) );
  XNOR U46287 ( .A(n45731), .B(n45729), .Z(n45946) );
  AND U46288 ( .A(n45947), .B(n45948), .Z(n45729) );
  NANDN U46289 ( .A(n45949), .B(n45950), .Z(n45948) );
  NANDN U46290 ( .A(n45951), .B(n45952), .Z(n45950) );
  NANDN U46291 ( .A(n45952), .B(n45951), .Z(n45947) );
  ANDN U46292 ( .B(B[114]), .A(n72), .Z(n45731) );
  XNOR U46293 ( .A(n45739), .B(n45953), .Z(n45732) );
  XNOR U46294 ( .A(n45738), .B(n45736), .Z(n45953) );
  AND U46295 ( .A(n45954), .B(n45955), .Z(n45736) );
  NANDN U46296 ( .A(n45956), .B(n45957), .Z(n45955) );
  OR U46297 ( .A(n45958), .B(n45959), .Z(n45957) );
  NAND U46298 ( .A(n45959), .B(n45958), .Z(n45954) );
  ANDN U46299 ( .B(B[115]), .A(n73), .Z(n45738) );
  XNOR U46300 ( .A(n45746), .B(n45960), .Z(n45739) );
  XNOR U46301 ( .A(n45745), .B(n45743), .Z(n45960) );
  AND U46302 ( .A(n45961), .B(n45962), .Z(n45743) );
  NANDN U46303 ( .A(n45963), .B(n45964), .Z(n45962) );
  NANDN U46304 ( .A(n45965), .B(n45966), .Z(n45964) );
  NANDN U46305 ( .A(n45966), .B(n45965), .Z(n45961) );
  ANDN U46306 ( .B(B[116]), .A(n74), .Z(n45745) );
  XNOR U46307 ( .A(n45753), .B(n45967), .Z(n45746) );
  XNOR U46308 ( .A(n45752), .B(n45750), .Z(n45967) );
  AND U46309 ( .A(n45968), .B(n45969), .Z(n45750) );
  NANDN U46310 ( .A(n45970), .B(n45971), .Z(n45969) );
  OR U46311 ( .A(n45972), .B(n45973), .Z(n45971) );
  NAND U46312 ( .A(n45973), .B(n45972), .Z(n45968) );
  ANDN U46313 ( .B(B[117]), .A(n75), .Z(n45752) );
  XNOR U46314 ( .A(n45760), .B(n45974), .Z(n45753) );
  XNOR U46315 ( .A(n45759), .B(n45757), .Z(n45974) );
  AND U46316 ( .A(n45975), .B(n45976), .Z(n45757) );
  NANDN U46317 ( .A(n45977), .B(n45978), .Z(n45976) );
  NANDN U46318 ( .A(n45979), .B(n45980), .Z(n45978) );
  NANDN U46319 ( .A(n45980), .B(n45979), .Z(n45975) );
  ANDN U46320 ( .B(B[118]), .A(n76), .Z(n45759) );
  XNOR U46321 ( .A(n45767), .B(n45981), .Z(n45760) );
  XNOR U46322 ( .A(n45766), .B(n45764), .Z(n45981) );
  AND U46323 ( .A(n45982), .B(n45983), .Z(n45764) );
  NANDN U46324 ( .A(n45984), .B(n45985), .Z(n45983) );
  OR U46325 ( .A(n45986), .B(n45987), .Z(n45985) );
  NAND U46326 ( .A(n45987), .B(n45986), .Z(n45982) );
  ANDN U46327 ( .B(B[119]), .A(n77), .Z(n45766) );
  XNOR U46328 ( .A(n45774), .B(n45988), .Z(n45767) );
  XNOR U46329 ( .A(n45773), .B(n45771), .Z(n45988) );
  AND U46330 ( .A(n45989), .B(n45990), .Z(n45771) );
  NANDN U46331 ( .A(n45991), .B(n45992), .Z(n45990) );
  NANDN U46332 ( .A(n45993), .B(n45994), .Z(n45992) );
  NANDN U46333 ( .A(n45994), .B(n45993), .Z(n45989) );
  ANDN U46334 ( .B(B[120]), .A(n78), .Z(n45773) );
  XNOR U46335 ( .A(n45781), .B(n45995), .Z(n45774) );
  XNOR U46336 ( .A(n45780), .B(n45778), .Z(n45995) );
  AND U46337 ( .A(n45996), .B(n45997), .Z(n45778) );
  NANDN U46338 ( .A(n45998), .B(n45999), .Z(n45997) );
  OR U46339 ( .A(n46000), .B(n46001), .Z(n45999) );
  NAND U46340 ( .A(n46001), .B(n46000), .Z(n45996) );
  ANDN U46341 ( .B(B[121]), .A(n79), .Z(n45780) );
  XNOR U46342 ( .A(n45788), .B(n46002), .Z(n45781) );
  XNOR U46343 ( .A(n45787), .B(n45785), .Z(n46002) );
  AND U46344 ( .A(n46003), .B(n46004), .Z(n45785) );
  NANDN U46345 ( .A(n46005), .B(n46006), .Z(n46004) );
  NANDN U46346 ( .A(n46007), .B(n46008), .Z(n46006) );
  NANDN U46347 ( .A(n46008), .B(n46007), .Z(n46003) );
  ANDN U46348 ( .B(B[122]), .A(n80), .Z(n45787) );
  XNOR U46349 ( .A(n45795), .B(n46009), .Z(n45788) );
  XNOR U46350 ( .A(n45794), .B(n45792), .Z(n46009) );
  AND U46351 ( .A(n46010), .B(n46011), .Z(n45792) );
  NANDN U46352 ( .A(n46012), .B(n46013), .Z(n46011) );
  OR U46353 ( .A(n46014), .B(n46015), .Z(n46013) );
  NAND U46354 ( .A(n46015), .B(n46014), .Z(n46010) );
  ANDN U46355 ( .B(B[123]), .A(n81), .Z(n45794) );
  XNOR U46356 ( .A(n45802), .B(n46016), .Z(n45795) );
  XNOR U46357 ( .A(n45801), .B(n45799), .Z(n46016) );
  AND U46358 ( .A(n46017), .B(n46018), .Z(n45799) );
  NANDN U46359 ( .A(n46019), .B(n46020), .Z(n46018) );
  NAND U46360 ( .A(n46021), .B(n46022), .Z(n46020) );
  ANDN U46361 ( .B(B[124]), .A(n82), .Z(n45801) );
  XOR U46362 ( .A(n45808), .B(n46023), .Z(n45802) );
  XNOR U46363 ( .A(n45806), .B(n45809), .Z(n46023) );
  NAND U46364 ( .A(A[2]), .B(B[125]), .Z(n45809) );
  NANDN U46365 ( .A(n46024), .B(n46025), .Z(n45806) );
  AND U46366 ( .A(A[0]), .B(B[126]), .Z(n46025) );
  XNOR U46367 ( .A(n45811), .B(n46026), .Z(n45808) );
  NAND U46368 ( .A(A[0]), .B(B[127]), .Z(n46026) );
  NAND U46369 ( .A(B[126]), .B(A[1]), .Z(n45811) );
  NAND U46370 ( .A(n46027), .B(n46028), .Z(n542) );
  NANDN U46371 ( .A(n46029), .B(n46030), .Z(n46028) );
  OR U46372 ( .A(n46031), .B(n46032), .Z(n46030) );
  NAND U46373 ( .A(n46032), .B(n46031), .Z(n46027) );
  XOR U46374 ( .A(n544), .B(n543), .Z(\A1[124] ) );
  XOR U46375 ( .A(n46032), .B(n46033), .Z(n543) );
  XNOR U46376 ( .A(n46031), .B(n46029), .Z(n46033) );
  AND U46377 ( .A(n46034), .B(n46035), .Z(n46029) );
  NANDN U46378 ( .A(n46036), .B(n46037), .Z(n46035) );
  NANDN U46379 ( .A(n46038), .B(n46039), .Z(n46037) );
  NANDN U46380 ( .A(n46039), .B(n46038), .Z(n46034) );
  ANDN U46381 ( .B(B[95]), .A(n54), .Z(n46031) );
  XNOR U46382 ( .A(n45826), .B(n46040), .Z(n46032) );
  XNOR U46383 ( .A(n45825), .B(n45823), .Z(n46040) );
  AND U46384 ( .A(n46041), .B(n46042), .Z(n45823) );
  NANDN U46385 ( .A(n46043), .B(n46044), .Z(n46042) );
  OR U46386 ( .A(n46045), .B(n46046), .Z(n46044) );
  NAND U46387 ( .A(n46046), .B(n46045), .Z(n46041) );
  ANDN U46388 ( .B(B[96]), .A(n55), .Z(n45825) );
  XNOR U46389 ( .A(n45833), .B(n46047), .Z(n45826) );
  XNOR U46390 ( .A(n45832), .B(n45830), .Z(n46047) );
  AND U46391 ( .A(n46048), .B(n46049), .Z(n45830) );
  NANDN U46392 ( .A(n46050), .B(n46051), .Z(n46049) );
  NANDN U46393 ( .A(n46052), .B(n46053), .Z(n46051) );
  NANDN U46394 ( .A(n46053), .B(n46052), .Z(n46048) );
  ANDN U46395 ( .B(A[29]), .A(n9), .Z(n45832) );
  XNOR U46396 ( .A(n45840), .B(n46054), .Z(n45833) );
  XNOR U46397 ( .A(n45839), .B(n45837), .Z(n46054) );
  AND U46398 ( .A(n46055), .B(n46056), .Z(n45837) );
  NANDN U46399 ( .A(n46057), .B(n46058), .Z(n46056) );
  OR U46400 ( .A(n46059), .B(n46060), .Z(n46058) );
  NAND U46401 ( .A(n46060), .B(n46059), .Z(n46055) );
  ANDN U46402 ( .B(B[98]), .A(n57), .Z(n45839) );
  XNOR U46403 ( .A(n45847), .B(n46061), .Z(n45840) );
  XNOR U46404 ( .A(n45846), .B(n45844), .Z(n46061) );
  AND U46405 ( .A(n46062), .B(n46063), .Z(n45844) );
  NANDN U46406 ( .A(n46064), .B(n46065), .Z(n46063) );
  NANDN U46407 ( .A(n46066), .B(n46067), .Z(n46065) );
  NANDN U46408 ( .A(n46067), .B(n46066), .Z(n46062) );
  ANDN U46409 ( .B(A[27]), .A(n6), .Z(n45846) );
  XNOR U46410 ( .A(n45854), .B(n46068), .Z(n45847) );
  XNOR U46411 ( .A(n45853), .B(n45851), .Z(n46068) );
  AND U46412 ( .A(n46069), .B(n46070), .Z(n45851) );
  NANDN U46413 ( .A(n46071), .B(n46072), .Z(n46070) );
  OR U46414 ( .A(n46073), .B(n46074), .Z(n46072) );
  NAND U46415 ( .A(n46074), .B(n46073), .Z(n46069) );
  ANDN U46416 ( .B(A[26]), .A(n4), .Z(n45853) );
  XNOR U46417 ( .A(n45861), .B(n46075), .Z(n45854) );
  XNOR U46418 ( .A(n45860), .B(n45858), .Z(n46075) );
  AND U46419 ( .A(n46076), .B(n46077), .Z(n45858) );
  NANDN U46420 ( .A(n46078), .B(n46079), .Z(n46077) );
  NANDN U46421 ( .A(n46080), .B(n46081), .Z(n46079) );
  NANDN U46422 ( .A(n46081), .B(n46080), .Z(n46076) );
  ANDN U46423 ( .B(B[101]), .A(n60), .Z(n45860) );
  XNOR U46424 ( .A(n45868), .B(n46082), .Z(n45861) );
  XNOR U46425 ( .A(n45867), .B(n45865), .Z(n46082) );
  AND U46426 ( .A(n46083), .B(n46084), .Z(n45865) );
  NANDN U46427 ( .A(n46085), .B(n46086), .Z(n46084) );
  OR U46428 ( .A(n46087), .B(n46088), .Z(n46086) );
  NAND U46429 ( .A(n46088), .B(n46087), .Z(n46083) );
  ANDN U46430 ( .B(B[102]), .A(n61), .Z(n45867) );
  XNOR U46431 ( .A(n45875), .B(n46089), .Z(n45868) );
  XNOR U46432 ( .A(n45874), .B(n45872), .Z(n46089) );
  AND U46433 ( .A(n46090), .B(n46091), .Z(n45872) );
  NANDN U46434 ( .A(n46092), .B(n46093), .Z(n46091) );
  NANDN U46435 ( .A(n46094), .B(n46095), .Z(n46093) );
  NANDN U46436 ( .A(n46095), .B(n46094), .Z(n46090) );
  ANDN U46437 ( .B(B[103]), .A(n62), .Z(n45874) );
  XNOR U46438 ( .A(n45882), .B(n46096), .Z(n45875) );
  XNOR U46439 ( .A(n45881), .B(n45879), .Z(n46096) );
  AND U46440 ( .A(n46097), .B(n46098), .Z(n45879) );
  NANDN U46441 ( .A(n46099), .B(n46100), .Z(n46098) );
  OR U46442 ( .A(n46101), .B(n46102), .Z(n46100) );
  NAND U46443 ( .A(n46102), .B(n46101), .Z(n46097) );
  ANDN U46444 ( .B(B[104]), .A(n63), .Z(n45881) );
  XNOR U46445 ( .A(n45889), .B(n46103), .Z(n45882) );
  XNOR U46446 ( .A(n45888), .B(n45886), .Z(n46103) );
  AND U46447 ( .A(n46104), .B(n46105), .Z(n45886) );
  NANDN U46448 ( .A(n46106), .B(n46107), .Z(n46105) );
  NANDN U46449 ( .A(n46108), .B(n46109), .Z(n46107) );
  NANDN U46450 ( .A(n46109), .B(n46108), .Z(n46104) );
  ANDN U46451 ( .B(B[105]), .A(n64), .Z(n45888) );
  XNOR U46452 ( .A(n45896), .B(n46110), .Z(n45889) );
  XNOR U46453 ( .A(n45895), .B(n45893), .Z(n46110) );
  AND U46454 ( .A(n46111), .B(n46112), .Z(n45893) );
  NANDN U46455 ( .A(n46113), .B(n46114), .Z(n46112) );
  OR U46456 ( .A(n46115), .B(n46116), .Z(n46114) );
  NAND U46457 ( .A(n46116), .B(n46115), .Z(n46111) );
  ANDN U46458 ( .B(B[106]), .A(n65), .Z(n45895) );
  XNOR U46459 ( .A(n45903), .B(n46117), .Z(n45896) );
  XNOR U46460 ( .A(n45902), .B(n45900), .Z(n46117) );
  AND U46461 ( .A(n46118), .B(n46119), .Z(n45900) );
  NANDN U46462 ( .A(n46120), .B(n46121), .Z(n46119) );
  NANDN U46463 ( .A(n46122), .B(n46123), .Z(n46121) );
  NANDN U46464 ( .A(n46123), .B(n46122), .Z(n46118) );
  ANDN U46465 ( .B(B[107]), .A(n66), .Z(n45902) );
  XNOR U46466 ( .A(n45910), .B(n46124), .Z(n45903) );
  XNOR U46467 ( .A(n45909), .B(n45907), .Z(n46124) );
  AND U46468 ( .A(n46125), .B(n46126), .Z(n45907) );
  NANDN U46469 ( .A(n46127), .B(n46128), .Z(n46126) );
  OR U46470 ( .A(n46129), .B(n46130), .Z(n46128) );
  NAND U46471 ( .A(n46130), .B(n46129), .Z(n46125) );
  ANDN U46472 ( .B(B[108]), .A(n67), .Z(n45909) );
  XNOR U46473 ( .A(n45917), .B(n46131), .Z(n45910) );
  XNOR U46474 ( .A(n45916), .B(n45914), .Z(n46131) );
  AND U46475 ( .A(n46132), .B(n46133), .Z(n45914) );
  NANDN U46476 ( .A(n46134), .B(n46135), .Z(n46133) );
  NANDN U46477 ( .A(n46136), .B(n46137), .Z(n46135) );
  NANDN U46478 ( .A(n46137), .B(n46136), .Z(n46132) );
  ANDN U46479 ( .B(B[109]), .A(n68), .Z(n45916) );
  XNOR U46480 ( .A(n45924), .B(n46138), .Z(n45917) );
  XNOR U46481 ( .A(n45923), .B(n45921), .Z(n46138) );
  AND U46482 ( .A(n46139), .B(n46140), .Z(n45921) );
  NANDN U46483 ( .A(n46141), .B(n46142), .Z(n46140) );
  OR U46484 ( .A(n46143), .B(n46144), .Z(n46142) );
  NAND U46485 ( .A(n46144), .B(n46143), .Z(n46139) );
  ANDN U46486 ( .B(B[110]), .A(n69), .Z(n45923) );
  XNOR U46487 ( .A(n45931), .B(n46145), .Z(n45924) );
  XNOR U46488 ( .A(n45930), .B(n45928), .Z(n46145) );
  AND U46489 ( .A(n46146), .B(n46147), .Z(n45928) );
  NANDN U46490 ( .A(n46148), .B(n46149), .Z(n46147) );
  NANDN U46491 ( .A(n46150), .B(n46151), .Z(n46149) );
  NANDN U46492 ( .A(n46151), .B(n46150), .Z(n46146) );
  ANDN U46493 ( .B(B[111]), .A(n70), .Z(n45930) );
  XNOR U46494 ( .A(n45938), .B(n46152), .Z(n45931) );
  XNOR U46495 ( .A(n45937), .B(n45935), .Z(n46152) );
  AND U46496 ( .A(n46153), .B(n46154), .Z(n45935) );
  NANDN U46497 ( .A(n46155), .B(n46156), .Z(n46154) );
  OR U46498 ( .A(n46157), .B(n46158), .Z(n46156) );
  NAND U46499 ( .A(n46158), .B(n46157), .Z(n46153) );
  ANDN U46500 ( .B(B[112]), .A(n71), .Z(n45937) );
  XNOR U46501 ( .A(n45945), .B(n46159), .Z(n45938) );
  XNOR U46502 ( .A(n45944), .B(n45942), .Z(n46159) );
  AND U46503 ( .A(n46160), .B(n46161), .Z(n45942) );
  NANDN U46504 ( .A(n46162), .B(n46163), .Z(n46161) );
  NANDN U46505 ( .A(n46164), .B(n46165), .Z(n46163) );
  NANDN U46506 ( .A(n46165), .B(n46164), .Z(n46160) );
  ANDN U46507 ( .B(B[113]), .A(n72), .Z(n45944) );
  XNOR U46508 ( .A(n45952), .B(n46166), .Z(n45945) );
  XNOR U46509 ( .A(n45951), .B(n45949), .Z(n46166) );
  AND U46510 ( .A(n46167), .B(n46168), .Z(n45949) );
  NANDN U46511 ( .A(n46169), .B(n46170), .Z(n46168) );
  OR U46512 ( .A(n46171), .B(n46172), .Z(n46170) );
  NAND U46513 ( .A(n46172), .B(n46171), .Z(n46167) );
  ANDN U46514 ( .B(B[114]), .A(n73), .Z(n45951) );
  XNOR U46515 ( .A(n45959), .B(n46173), .Z(n45952) );
  XNOR U46516 ( .A(n45958), .B(n45956), .Z(n46173) );
  AND U46517 ( .A(n46174), .B(n46175), .Z(n45956) );
  NANDN U46518 ( .A(n46176), .B(n46177), .Z(n46175) );
  NANDN U46519 ( .A(n46178), .B(n46179), .Z(n46177) );
  NANDN U46520 ( .A(n46179), .B(n46178), .Z(n46174) );
  ANDN U46521 ( .B(B[115]), .A(n74), .Z(n45958) );
  XNOR U46522 ( .A(n45966), .B(n46180), .Z(n45959) );
  XNOR U46523 ( .A(n45965), .B(n45963), .Z(n46180) );
  AND U46524 ( .A(n46181), .B(n46182), .Z(n45963) );
  NANDN U46525 ( .A(n46183), .B(n46184), .Z(n46182) );
  OR U46526 ( .A(n46185), .B(n46186), .Z(n46184) );
  NAND U46527 ( .A(n46186), .B(n46185), .Z(n46181) );
  ANDN U46528 ( .B(B[116]), .A(n75), .Z(n45965) );
  XNOR U46529 ( .A(n45973), .B(n46187), .Z(n45966) );
  XNOR U46530 ( .A(n45972), .B(n45970), .Z(n46187) );
  AND U46531 ( .A(n46188), .B(n46189), .Z(n45970) );
  NANDN U46532 ( .A(n46190), .B(n46191), .Z(n46189) );
  NANDN U46533 ( .A(n46192), .B(n46193), .Z(n46191) );
  NANDN U46534 ( .A(n46193), .B(n46192), .Z(n46188) );
  ANDN U46535 ( .B(B[117]), .A(n76), .Z(n45972) );
  XNOR U46536 ( .A(n45980), .B(n46194), .Z(n45973) );
  XNOR U46537 ( .A(n45979), .B(n45977), .Z(n46194) );
  AND U46538 ( .A(n46195), .B(n46196), .Z(n45977) );
  NANDN U46539 ( .A(n46197), .B(n46198), .Z(n46196) );
  OR U46540 ( .A(n46199), .B(n46200), .Z(n46198) );
  NAND U46541 ( .A(n46200), .B(n46199), .Z(n46195) );
  ANDN U46542 ( .B(B[118]), .A(n77), .Z(n45979) );
  XNOR U46543 ( .A(n45987), .B(n46201), .Z(n45980) );
  XNOR U46544 ( .A(n45986), .B(n45984), .Z(n46201) );
  AND U46545 ( .A(n46202), .B(n46203), .Z(n45984) );
  NANDN U46546 ( .A(n46204), .B(n46205), .Z(n46203) );
  NANDN U46547 ( .A(n46206), .B(n46207), .Z(n46205) );
  NANDN U46548 ( .A(n46207), .B(n46206), .Z(n46202) );
  ANDN U46549 ( .B(B[119]), .A(n78), .Z(n45986) );
  XNOR U46550 ( .A(n45994), .B(n46208), .Z(n45987) );
  XNOR U46551 ( .A(n45993), .B(n45991), .Z(n46208) );
  AND U46552 ( .A(n46209), .B(n46210), .Z(n45991) );
  NANDN U46553 ( .A(n46211), .B(n46212), .Z(n46210) );
  OR U46554 ( .A(n46213), .B(n46214), .Z(n46212) );
  NAND U46555 ( .A(n46214), .B(n46213), .Z(n46209) );
  ANDN U46556 ( .B(B[120]), .A(n79), .Z(n45993) );
  XNOR U46557 ( .A(n46001), .B(n46215), .Z(n45994) );
  XNOR U46558 ( .A(n46000), .B(n45998), .Z(n46215) );
  AND U46559 ( .A(n46216), .B(n46217), .Z(n45998) );
  NANDN U46560 ( .A(n46218), .B(n46219), .Z(n46217) );
  NANDN U46561 ( .A(n46220), .B(n46221), .Z(n46219) );
  NANDN U46562 ( .A(n46221), .B(n46220), .Z(n46216) );
  ANDN U46563 ( .B(B[121]), .A(n80), .Z(n46000) );
  XNOR U46564 ( .A(n46008), .B(n46222), .Z(n46001) );
  XNOR U46565 ( .A(n46007), .B(n46005), .Z(n46222) );
  AND U46566 ( .A(n46223), .B(n46224), .Z(n46005) );
  NANDN U46567 ( .A(n46225), .B(n46226), .Z(n46224) );
  OR U46568 ( .A(n46227), .B(n46228), .Z(n46226) );
  NAND U46569 ( .A(n46228), .B(n46227), .Z(n46223) );
  ANDN U46570 ( .B(B[122]), .A(n81), .Z(n46007) );
  XNOR U46571 ( .A(n46015), .B(n46229), .Z(n46008) );
  XNOR U46572 ( .A(n46014), .B(n46012), .Z(n46229) );
  AND U46573 ( .A(n46230), .B(n46231), .Z(n46012) );
  NANDN U46574 ( .A(n46232), .B(n46233), .Z(n46231) );
  NAND U46575 ( .A(n46234), .B(n46235), .Z(n46233) );
  ANDN U46576 ( .B(B[123]), .A(n82), .Z(n46014) );
  XOR U46577 ( .A(n46021), .B(n46236), .Z(n46015) );
  XNOR U46578 ( .A(n46019), .B(n46022), .Z(n46236) );
  NAND U46579 ( .A(A[2]), .B(B[124]), .Z(n46022) );
  NANDN U46580 ( .A(n46237), .B(n46238), .Z(n46019) );
  AND U46581 ( .A(A[0]), .B(B[125]), .Z(n46238) );
  XNOR U46582 ( .A(n46024), .B(n46239), .Z(n46021) );
  NAND U46583 ( .A(A[0]), .B(B[126]), .Z(n46239) );
  NAND U46584 ( .A(B[125]), .B(A[1]), .Z(n46024) );
  NAND U46585 ( .A(n46240), .B(n46241), .Z(n544) );
  NANDN U46586 ( .A(n46242), .B(n46243), .Z(n46241) );
  OR U46587 ( .A(n46244), .B(n46245), .Z(n46243) );
  NAND U46588 ( .A(n46245), .B(n46244), .Z(n46240) );
  XOR U46589 ( .A(n546), .B(n545), .Z(\A1[123] ) );
  XOR U46590 ( .A(n46245), .B(n46246), .Z(n545) );
  XNOR U46591 ( .A(n46244), .B(n46242), .Z(n46246) );
  AND U46592 ( .A(n46247), .B(n46248), .Z(n46242) );
  NANDN U46593 ( .A(n46249), .B(n46250), .Z(n46248) );
  NANDN U46594 ( .A(n46251), .B(n46252), .Z(n46250) );
  NANDN U46595 ( .A(n46252), .B(n46251), .Z(n46247) );
  ANDN U46596 ( .B(B[94]), .A(n54), .Z(n46244) );
  XNOR U46597 ( .A(n46039), .B(n46253), .Z(n46245) );
  XNOR U46598 ( .A(n46038), .B(n46036), .Z(n46253) );
  AND U46599 ( .A(n46254), .B(n46255), .Z(n46036) );
  NANDN U46600 ( .A(n46256), .B(n46257), .Z(n46255) );
  OR U46601 ( .A(n46258), .B(n46259), .Z(n46257) );
  NAND U46602 ( .A(n46259), .B(n46258), .Z(n46254) );
  ANDN U46603 ( .B(B[95]), .A(n55), .Z(n46038) );
  XNOR U46604 ( .A(n46046), .B(n46260), .Z(n46039) );
  XNOR U46605 ( .A(n46045), .B(n46043), .Z(n46260) );
  AND U46606 ( .A(n46261), .B(n46262), .Z(n46043) );
  NANDN U46607 ( .A(n46263), .B(n46264), .Z(n46262) );
  NANDN U46608 ( .A(n46265), .B(n46266), .Z(n46264) );
  NANDN U46609 ( .A(n46266), .B(n46265), .Z(n46261) );
  ANDN U46610 ( .B(B[96]), .A(n56), .Z(n46045) );
  XNOR U46611 ( .A(n46053), .B(n46267), .Z(n46046) );
  XNOR U46612 ( .A(n46052), .B(n46050), .Z(n46267) );
  AND U46613 ( .A(n46268), .B(n46269), .Z(n46050) );
  NANDN U46614 ( .A(n46270), .B(n46271), .Z(n46269) );
  OR U46615 ( .A(n46272), .B(n46273), .Z(n46271) );
  NAND U46616 ( .A(n46273), .B(n46272), .Z(n46268) );
  ANDN U46617 ( .B(A[28]), .A(n9), .Z(n46052) );
  XNOR U46618 ( .A(n46060), .B(n46274), .Z(n46053) );
  XNOR U46619 ( .A(n46059), .B(n46057), .Z(n46274) );
  AND U46620 ( .A(n46275), .B(n46276), .Z(n46057) );
  NANDN U46621 ( .A(n46277), .B(n46278), .Z(n46276) );
  NANDN U46622 ( .A(n46279), .B(n46280), .Z(n46278) );
  NANDN U46623 ( .A(n46280), .B(n46279), .Z(n46275) );
  ANDN U46624 ( .B(B[98]), .A(n58), .Z(n46059) );
  XNOR U46625 ( .A(n46067), .B(n46281), .Z(n46060) );
  XNOR U46626 ( .A(n46066), .B(n46064), .Z(n46281) );
  AND U46627 ( .A(n46282), .B(n46283), .Z(n46064) );
  NANDN U46628 ( .A(n46284), .B(n46285), .Z(n46283) );
  OR U46629 ( .A(n46286), .B(n46287), .Z(n46285) );
  NAND U46630 ( .A(n46287), .B(n46286), .Z(n46282) );
  ANDN U46631 ( .B(A[26]), .A(n6), .Z(n46066) );
  XNOR U46632 ( .A(n46074), .B(n46288), .Z(n46067) );
  XNOR U46633 ( .A(n46073), .B(n46071), .Z(n46288) );
  AND U46634 ( .A(n46289), .B(n46290), .Z(n46071) );
  NANDN U46635 ( .A(n46291), .B(n46292), .Z(n46290) );
  NANDN U46636 ( .A(n46293), .B(n46294), .Z(n46292) );
  NANDN U46637 ( .A(n46294), .B(n46293), .Z(n46289) );
  ANDN U46638 ( .B(A[25]), .A(n4), .Z(n46073) );
  XNOR U46639 ( .A(n46081), .B(n46295), .Z(n46074) );
  XNOR U46640 ( .A(n46080), .B(n46078), .Z(n46295) );
  AND U46641 ( .A(n46296), .B(n46297), .Z(n46078) );
  NANDN U46642 ( .A(n46298), .B(n46299), .Z(n46297) );
  OR U46643 ( .A(n46300), .B(n46301), .Z(n46299) );
  NAND U46644 ( .A(n46301), .B(n46300), .Z(n46296) );
  ANDN U46645 ( .B(B[101]), .A(n61), .Z(n46080) );
  XNOR U46646 ( .A(n46088), .B(n46302), .Z(n46081) );
  XNOR U46647 ( .A(n46087), .B(n46085), .Z(n46302) );
  AND U46648 ( .A(n46303), .B(n46304), .Z(n46085) );
  NANDN U46649 ( .A(n46305), .B(n46306), .Z(n46304) );
  NANDN U46650 ( .A(n46307), .B(n46308), .Z(n46306) );
  NANDN U46651 ( .A(n46308), .B(n46307), .Z(n46303) );
  ANDN U46652 ( .B(B[102]), .A(n62), .Z(n46087) );
  XNOR U46653 ( .A(n46095), .B(n46309), .Z(n46088) );
  XNOR U46654 ( .A(n46094), .B(n46092), .Z(n46309) );
  AND U46655 ( .A(n46310), .B(n46311), .Z(n46092) );
  NANDN U46656 ( .A(n46312), .B(n46313), .Z(n46311) );
  OR U46657 ( .A(n46314), .B(n46315), .Z(n46313) );
  NAND U46658 ( .A(n46315), .B(n46314), .Z(n46310) );
  ANDN U46659 ( .B(B[103]), .A(n63), .Z(n46094) );
  XNOR U46660 ( .A(n46102), .B(n46316), .Z(n46095) );
  XNOR U46661 ( .A(n46101), .B(n46099), .Z(n46316) );
  AND U46662 ( .A(n46317), .B(n46318), .Z(n46099) );
  NANDN U46663 ( .A(n46319), .B(n46320), .Z(n46318) );
  NANDN U46664 ( .A(n46321), .B(n46322), .Z(n46320) );
  NANDN U46665 ( .A(n46322), .B(n46321), .Z(n46317) );
  ANDN U46666 ( .B(B[104]), .A(n64), .Z(n46101) );
  XNOR U46667 ( .A(n46109), .B(n46323), .Z(n46102) );
  XNOR U46668 ( .A(n46108), .B(n46106), .Z(n46323) );
  AND U46669 ( .A(n46324), .B(n46325), .Z(n46106) );
  NANDN U46670 ( .A(n46326), .B(n46327), .Z(n46325) );
  OR U46671 ( .A(n46328), .B(n46329), .Z(n46327) );
  NAND U46672 ( .A(n46329), .B(n46328), .Z(n46324) );
  ANDN U46673 ( .B(B[105]), .A(n65), .Z(n46108) );
  XNOR U46674 ( .A(n46116), .B(n46330), .Z(n46109) );
  XNOR U46675 ( .A(n46115), .B(n46113), .Z(n46330) );
  AND U46676 ( .A(n46331), .B(n46332), .Z(n46113) );
  NANDN U46677 ( .A(n46333), .B(n46334), .Z(n46332) );
  NANDN U46678 ( .A(n46335), .B(n46336), .Z(n46334) );
  NANDN U46679 ( .A(n46336), .B(n46335), .Z(n46331) );
  ANDN U46680 ( .B(B[106]), .A(n66), .Z(n46115) );
  XNOR U46681 ( .A(n46123), .B(n46337), .Z(n46116) );
  XNOR U46682 ( .A(n46122), .B(n46120), .Z(n46337) );
  AND U46683 ( .A(n46338), .B(n46339), .Z(n46120) );
  NANDN U46684 ( .A(n46340), .B(n46341), .Z(n46339) );
  OR U46685 ( .A(n46342), .B(n46343), .Z(n46341) );
  NAND U46686 ( .A(n46343), .B(n46342), .Z(n46338) );
  ANDN U46687 ( .B(B[107]), .A(n67), .Z(n46122) );
  XNOR U46688 ( .A(n46130), .B(n46344), .Z(n46123) );
  XNOR U46689 ( .A(n46129), .B(n46127), .Z(n46344) );
  AND U46690 ( .A(n46345), .B(n46346), .Z(n46127) );
  NANDN U46691 ( .A(n46347), .B(n46348), .Z(n46346) );
  NANDN U46692 ( .A(n46349), .B(n46350), .Z(n46348) );
  NANDN U46693 ( .A(n46350), .B(n46349), .Z(n46345) );
  ANDN U46694 ( .B(B[108]), .A(n68), .Z(n46129) );
  XNOR U46695 ( .A(n46137), .B(n46351), .Z(n46130) );
  XNOR U46696 ( .A(n46136), .B(n46134), .Z(n46351) );
  AND U46697 ( .A(n46352), .B(n46353), .Z(n46134) );
  NANDN U46698 ( .A(n46354), .B(n46355), .Z(n46353) );
  OR U46699 ( .A(n46356), .B(n46357), .Z(n46355) );
  NAND U46700 ( .A(n46357), .B(n46356), .Z(n46352) );
  ANDN U46701 ( .B(B[109]), .A(n69), .Z(n46136) );
  XNOR U46702 ( .A(n46144), .B(n46358), .Z(n46137) );
  XNOR U46703 ( .A(n46143), .B(n46141), .Z(n46358) );
  AND U46704 ( .A(n46359), .B(n46360), .Z(n46141) );
  NANDN U46705 ( .A(n46361), .B(n46362), .Z(n46360) );
  NANDN U46706 ( .A(n46363), .B(n46364), .Z(n46362) );
  NANDN U46707 ( .A(n46364), .B(n46363), .Z(n46359) );
  ANDN U46708 ( .B(B[110]), .A(n70), .Z(n46143) );
  XNOR U46709 ( .A(n46151), .B(n46365), .Z(n46144) );
  XNOR U46710 ( .A(n46150), .B(n46148), .Z(n46365) );
  AND U46711 ( .A(n46366), .B(n46367), .Z(n46148) );
  NANDN U46712 ( .A(n46368), .B(n46369), .Z(n46367) );
  OR U46713 ( .A(n46370), .B(n46371), .Z(n46369) );
  NAND U46714 ( .A(n46371), .B(n46370), .Z(n46366) );
  ANDN U46715 ( .B(B[111]), .A(n71), .Z(n46150) );
  XNOR U46716 ( .A(n46158), .B(n46372), .Z(n46151) );
  XNOR U46717 ( .A(n46157), .B(n46155), .Z(n46372) );
  AND U46718 ( .A(n46373), .B(n46374), .Z(n46155) );
  NANDN U46719 ( .A(n46375), .B(n46376), .Z(n46374) );
  NANDN U46720 ( .A(n46377), .B(n46378), .Z(n46376) );
  NANDN U46721 ( .A(n46378), .B(n46377), .Z(n46373) );
  ANDN U46722 ( .B(B[112]), .A(n72), .Z(n46157) );
  XNOR U46723 ( .A(n46165), .B(n46379), .Z(n46158) );
  XNOR U46724 ( .A(n46164), .B(n46162), .Z(n46379) );
  AND U46725 ( .A(n46380), .B(n46381), .Z(n46162) );
  NANDN U46726 ( .A(n46382), .B(n46383), .Z(n46381) );
  OR U46727 ( .A(n46384), .B(n46385), .Z(n46383) );
  NAND U46728 ( .A(n46385), .B(n46384), .Z(n46380) );
  ANDN U46729 ( .B(B[113]), .A(n73), .Z(n46164) );
  XNOR U46730 ( .A(n46172), .B(n46386), .Z(n46165) );
  XNOR U46731 ( .A(n46171), .B(n46169), .Z(n46386) );
  AND U46732 ( .A(n46387), .B(n46388), .Z(n46169) );
  NANDN U46733 ( .A(n46389), .B(n46390), .Z(n46388) );
  NANDN U46734 ( .A(n46391), .B(n46392), .Z(n46390) );
  NANDN U46735 ( .A(n46392), .B(n46391), .Z(n46387) );
  ANDN U46736 ( .B(B[114]), .A(n74), .Z(n46171) );
  XNOR U46737 ( .A(n46179), .B(n46393), .Z(n46172) );
  XNOR U46738 ( .A(n46178), .B(n46176), .Z(n46393) );
  AND U46739 ( .A(n46394), .B(n46395), .Z(n46176) );
  NANDN U46740 ( .A(n46396), .B(n46397), .Z(n46395) );
  OR U46741 ( .A(n46398), .B(n46399), .Z(n46397) );
  NAND U46742 ( .A(n46399), .B(n46398), .Z(n46394) );
  ANDN U46743 ( .B(B[115]), .A(n75), .Z(n46178) );
  XNOR U46744 ( .A(n46186), .B(n46400), .Z(n46179) );
  XNOR U46745 ( .A(n46185), .B(n46183), .Z(n46400) );
  AND U46746 ( .A(n46401), .B(n46402), .Z(n46183) );
  NANDN U46747 ( .A(n46403), .B(n46404), .Z(n46402) );
  NANDN U46748 ( .A(n46405), .B(n46406), .Z(n46404) );
  NANDN U46749 ( .A(n46406), .B(n46405), .Z(n46401) );
  ANDN U46750 ( .B(B[116]), .A(n76), .Z(n46185) );
  XNOR U46751 ( .A(n46193), .B(n46407), .Z(n46186) );
  XNOR U46752 ( .A(n46192), .B(n46190), .Z(n46407) );
  AND U46753 ( .A(n46408), .B(n46409), .Z(n46190) );
  NANDN U46754 ( .A(n46410), .B(n46411), .Z(n46409) );
  OR U46755 ( .A(n46412), .B(n46413), .Z(n46411) );
  NAND U46756 ( .A(n46413), .B(n46412), .Z(n46408) );
  ANDN U46757 ( .B(B[117]), .A(n77), .Z(n46192) );
  XNOR U46758 ( .A(n46200), .B(n46414), .Z(n46193) );
  XNOR U46759 ( .A(n46199), .B(n46197), .Z(n46414) );
  AND U46760 ( .A(n46415), .B(n46416), .Z(n46197) );
  NANDN U46761 ( .A(n46417), .B(n46418), .Z(n46416) );
  NANDN U46762 ( .A(n46419), .B(n46420), .Z(n46418) );
  NANDN U46763 ( .A(n46420), .B(n46419), .Z(n46415) );
  ANDN U46764 ( .B(B[118]), .A(n78), .Z(n46199) );
  XNOR U46765 ( .A(n46207), .B(n46421), .Z(n46200) );
  XNOR U46766 ( .A(n46206), .B(n46204), .Z(n46421) );
  AND U46767 ( .A(n46422), .B(n46423), .Z(n46204) );
  NANDN U46768 ( .A(n46424), .B(n46425), .Z(n46423) );
  OR U46769 ( .A(n46426), .B(n46427), .Z(n46425) );
  NAND U46770 ( .A(n46427), .B(n46426), .Z(n46422) );
  ANDN U46771 ( .B(B[119]), .A(n79), .Z(n46206) );
  XNOR U46772 ( .A(n46214), .B(n46428), .Z(n46207) );
  XNOR U46773 ( .A(n46213), .B(n46211), .Z(n46428) );
  AND U46774 ( .A(n46429), .B(n46430), .Z(n46211) );
  NANDN U46775 ( .A(n46431), .B(n46432), .Z(n46430) );
  NANDN U46776 ( .A(n46433), .B(n46434), .Z(n46432) );
  NANDN U46777 ( .A(n46434), .B(n46433), .Z(n46429) );
  ANDN U46778 ( .B(B[120]), .A(n80), .Z(n46213) );
  XNOR U46779 ( .A(n46221), .B(n46435), .Z(n46214) );
  XNOR U46780 ( .A(n46220), .B(n46218), .Z(n46435) );
  AND U46781 ( .A(n46436), .B(n46437), .Z(n46218) );
  NANDN U46782 ( .A(n46438), .B(n46439), .Z(n46437) );
  OR U46783 ( .A(n46440), .B(n46441), .Z(n46439) );
  NAND U46784 ( .A(n46441), .B(n46440), .Z(n46436) );
  ANDN U46785 ( .B(B[121]), .A(n81), .Z(n46220) );
  XNOR U46786 ( .A(n46228), .B(n46442), .Z(n46221) );
  XNOR U46787 ( .A(n46227), .B(n46225), .Z(n46442) );
  AND U46788 ( .A(n46443), .B(n46444), .Z(n46225) );
  NANDN U46789 ( .A(n46445), .B(n46446), .Z(n46444) );
  NAND U46790 ( .A(n46447), .B(n46448), .Z(n46446) );
  ANDN U46791 ( .B(B[122]), .A(n82), .Z(n46227) );
  XOR U46792 ( .A(n46234), .B(n46449), .Z(n46228) );
  XNOR U46793 ( .A(n46232), .B(n46235), .Z(n46449) );
  NAND U46794 ( .A(A[2]), .B(B[123]), .Z(n46235) );
  NANDN U46795 ( .A(n46450), .B(n46451), .Z(n46232) );
  AND U46796 ( .A(A[0]), .B(B[124]), .Z(n46451) );
  XNOR U46797 ( .A(n46237), .B(n46452), .Z(n46234) );
  NAND U46798 ( .A(A[0]), .B(B[125]), .Z(n46452) );
  NAND U46799 ( .A(B[124]), .B(A[1]), .Z(n46237) );
  NAND U46800 ( .A(n46453), .B(n46454), .Z(n546) );
  NANDN U46801 ( .A(n46455), .B(n46456), .Z(n46454) );
  OR U46802 ( .A(n46457), .B(n46458), .Z(n46456) );
  NAND U46803 ( .A(n46458), .B(n46457), .Z(n46453) );
  XOR U46804 ( .A(n548), .B(n547), .Z(\A1[122] ) );
  XOR U46805 ( .A(n46458), .B(n46459), .Z(n547) );
  XNOR U46806 ( .A(n46457), .B(n46455), .Z(n46459) );
  AND U46807 ( .A(n46460), .B(n46461), .Z(n46455) );
  NANDN U46808 ( .A(n46462), .B(n46463), .Z(n46461) );
  NANDN U46809 ( .A(n46464), .B(n46465), .Z(n46463) );
  NANDN U46810 ( .A(n46465), .B(n46464), .Z(n46460) );
  ANDN U46811 ( .B(B[93]), .A(n54), .Z(n46457) );
  XNOR U46812 ( .A(n46252), .B(n46466), .Z(n46458) );
  XNOR U46813 ( .A(n46251), .B(n46249), .Z(n46466) );
  AND U46814 ( .A(n46467), .B(n46468), .Z(n46249) );
  NANDN U46815 ( .A(n46469), .B(n46470), .Z(n46468) );
  OR U46816 ( .A(n46471), .B(n46472), .Z(n46470) );
  NAND U46817 ( .A(n46472), .B(n46471), .Z(n46467) );
  ANDN U46818 ( .B(B[94]), .A(n55), .Z(n46251) );
  XNOR U46819 ( .A(n46259), .B(n46473), .Z(n46252) );
  XNOR U46820 ( .A(n46258), .B(n46256), .Z(n46473) );
  AND U46821 ( .A(n46474), .B(n46475), .Z(n46256) );
  NANDN U46822 ( .A(n46476), .B(n46477), .Z(n46475) );
  NANDN U46823 ( .A(n46478), .B(n46479), .Z(n46477) );
  NANDN U46824 ( .A(n46479), .B(n46478), .Z(n46474) );
  ANDN U46825 ( .B(B[95]), .A(n56), .Z(n46258) );
  XNOR U46826 ( .A(n46266), .B(n46480), .Z(n46259) );
  XNOR U46827 ( .A(n46265), .B(n46263), .Z(n46480) );
  AND U46828 ( .A(n46481), .B(n46482), .Z(n46263) );
  NANDN U46829 ( .A(n46483), .B(n46484), .Z(n46482) );
  OR U46830 ( .A(n46485), .B(n46486), .Z(n46484) );
  NAND U46831 ( .A(n46486), .B(n46485), .Z(n46481) );
  ANDN U46832 ( .B(A[28]), .A(n11), .Z(n46265) );
  XNOR U46833 ( .A(n46273), .B(n46487), .Z(n46266) );
  XNOR U46834 ( .A(n46272), .B(n46270), .Z(n46487) );
  AND U46835 ( .A(n46488), .B(n46489), .Z(n46270) );
  NANDN U46836 ( .A(n46490), .B(n46491), .Z(n46489) );
  NANDN U46837 ( .A(n46492), .B(n46493), .Z(n46491) );
  NANDN U46838 ( .A(n46493), .B(n46492), .Z(n46488) );
  ANDN U46839 ( .B(A[27]), .A(n9), .Z(n46272) );
  XNOR U46840 ( .A(n46280), .B(n46494), .Z(n46273) );
  XNOR U46841 ( .A(n46279), .B(n46277), .Z(n46494) );
  AND U46842 ( .A(n46495), .B(n46496), .Z(n46277) );
  NANDN U46843 ( .A(n46497), .B(n46498), .Z(n46496) );
  OR U46844 ( .A(n46499), .B(n46500), .Z(n46498) );
  NAND U46845 ( .A(n46500), .B(n46499), .Z(n46495) );
  ANDN U46846 ( .B(B[98]), .A(n59), .Z(n46279) );
  XNOR U46847 ( .A(n46287), .B(n46501), .Z(n46280) );
  XNOR U46848 ( .A(n46286), .B(n46284), .Z(n46501) );
  AND U46849 ( .A(n46502), .B(n46503), .Z(n46284) );
  NANDN U46850 ( .A(n46504), .B(n46505), .Z(n46503) );
  NANDN U46851 ( .A(n46506), .B(n46507), .Z(n46505) );
  NANDN U46852 ( .A(n46507), .B(n46506), .Z(n46502) );
  ANDN U46853 ( .B(A[25]), .A(n6), .Z(n46286) );
  XNOR U46854 ( .A(n46294), .B(n46508), .Z(n46287) );
  XNOR U46855 ( .A(n46293), .B(n46291), .Z(n46508) );
  AND U46856 ( .A(n46509), .B(n46510), .Z(n46291) );
  NANDN U46857 ( .A(n46511), .B(n46512), .Z(n46510) );
  OR U46858 ( .A(n46513), .B(n46514), .Z(n46512) );
  NAND U46859 ( .A(n46514), .B(n46513), .Z(n46509) );
  ANDN U46860 ( .B(A[24]), .A(n4), .Z(n46293) );
  XNOR U46861 ( .A(n46301), .B(n46515), .Z(n46294) );
  XNOR U46862 ( .A(n46300), .B(n46298), .Z(n46515) );
  AND U46863 ( .A(n46516), .B(n46517), .Z(n46298) );
  NANDN U46864 ( .A(n46518), .B(n46519), .Z(n46517) );
  NANDN U46865 ( .A(n46520), .B(n46521), .Z(n46519) );
  NANDN U46866 ( .A(n46521), .B(n46520), .Z(n46516) );
  ANDN U46867 ( .B(B[101]), .A(n62), .Z(n46300) );
  XNOR U46868 ( .A(n46308), .B(n46522), .Z(n46301) );
  XNOR U46869 ( .A(n46307), .B(n46305), .Z(n46522) );
  AND U46870 ( .A(n46523), .B(n46524), .Z(n46305) );
  NANDN U46871 ( .A(n46525), .B(n46526), .Z(n46524) );
  OR U46872 ( .A(n46527), .B(n46528), .Z(n46526) );
  NAND U46873 ( .A(n46528), .B(n46527), .Z(n46523) );
  ANDN U46874 ( .B(B[102]), .A(n63), .Z(n46307) );
  XNOR U46875 ( .A(n46315), .B(n46529), .Z(n46308) );
  XNOR U46876 ( .A(n46314), .B(n46312), .Z(n46529) );
  AND U46877 ( .A(n46530), .B(n46531), .Z(n46312) );
  NANDN U46878 ( .A(n46532), .B(n46533), .Z(n46531) );
  NANDN U46879 ( .A(n46534), .B(n46535), .Z(n46533) );
  NANDN U46880 ( .A(n46535), .B(n46534), .Z(n46530) );
  ANDN U46881 ( .B(B[103]), .A(n64), .Z(n46314) );
  XNOR U46882 ( .A(n46322), .B(n46536), .Z(n46315) );
  XNOR U46883 ( .A(n46321), .B(n46319), .Z(n46536) );
  AND U46884 ( .A(n46537), .B(n46538), .Z(n46319) );
  NANDN U46885 ( .A(n46539), .B(n46540), .Z(n46538) );
  OR U46886 ( .A(n46541), .B(n46542), .Z(n46540) );
  NAND U46887 ( .A(n46542), .B(n46541), .Z(n46537) );
  ANDN U46888 ( .B(B[104]), .A(n65), .Z(n46321) );
  XNOR U46889 ( .A(n46329), .B(n46543), .Z(n46322) );
  XNOR U46890 ( .A(n46328), .B(n46326), .Z(n46543) );
  AND U46891 ( .A(n46544), .B(n46545), .Z(n46326) );
  NANDN U46892 ( .A(n46546), .B(n46547), .Z(n46545) );
  NANDN U46893 ( .A(n46548), .B(n46549), .Z(n46547) );
  NANDN U46894 ( .A(n46549), .B(n46548), .Z(n46544) );
  ANDN U46895 ( .B(B[105]), .A(n66), .Z(n46328) );
  XNOR U46896 ( .A(n46336), .B(n46550), .Z(n46329) );
  XNOR U46897 ( .A(n46335), .B(n46333), .Z(n46550) );
  AND U46898 ( .A(n46551), .B(n46552), .Z(n46333) );
  NANDN U46899 ( .A(n46553), .B(n46554), .Z(n46552) );
  OR U46900 ( .A(n46555), .B(n46556), .Z(n46554) );
  NAND U46901 ( .A(n46556), .B(n46555), .Z(n46551) );
  ANDN U46902 ( .B(B[106]), .A(n67), .Z(n46335) );
  XNOR U46903 ( .A(n46343), .B(n46557), .Z(n46336) );
  XNOR U46904 ( .A(n46342), .B(n46340), .Z(n46557) );
  AND U46905 ( .A(n46558), .B(n46559), .Z(n46340) );
  NANDN U46906 ( .A(n46560), .B(n46561), .Z(n46559) );
  NANDN U46907 ( .A(n46562), .B(n46563), .Z(n46561) );
  NANDN U46908 ( .A(n46563), .B(n46562), .Z(n46558) );
  ANDN U46909 ( .B(B[107]), .A(n68), .Z(n46342) );
  XNOR U46910 ( .A(n46350), .B(n46564), .Z(n46343) );
  XNOR U46911 ( .A(n46349), .B(n46347), .Z(n46564) );
  AND U46912 ( .A(n46565), .B(n46566), .Z(n46347) );
  NANDN U46913 ( .A(n46567), .B(n46568), .Z(n46566) );
  OR U46914 ( .A(n46569), .B(n46570), .Z(n46568) );
  NAND U46915 ( .A(n46570), .B(n46569), .Z(n46565) );
  ANDN U46916 ( .B(B[108]), .A(n69), .Z(n46349) );
  XNOR U46917 ( .A(n46357), .B(n46571), .Z(n46350) );
  XNOR U46918 ( .A(n46356), .B(n46354), .Z(n46571) );
  AND U46919 ( .A(n46572), .B(n46573), .Z(n46354) );
  NANDN U46920 ( .A(n46574), .B(n46575), .Z(n46573) );
  NANDN U46921 ( .A(n46576), .B(n46577), .Z(n46575) );
  NANDN U46922 ( .A(n46577), .B(n46576), .Z(n46572) );
  ANDN U46923 ( .B(B[109]), .A(n70), .Z(n46356) );
  XNOR U46924 ( .A(n46364), .B(n46578), .Z(n46357) );
  XNOR U46925 ( .A(n46363), .B(n46361), .Z(n46578) );
  AND U46926 ( .A(n46579), .B(n46580), .Z(n46361) );
  NANDN U46927 ( .A(n46581), .B(n46582), .Z(n46580) );
  OR U46928 ( .A(n46583), .B(n46584), .Z(n46582) );
  NAND U46929 ( .A(n46584), .B(n46583), .Z(n46579) );
  ANDN U46930 ( .B(B[110]), .A(n71), .Z(n46363) );
  XNOR U46931 ( .A(n46371), .B(n46585), .Z(n46364) );
  XNOR U46932 ( .A(n46370), .B(n46368), .Z(n46585) );
  AND U46933 ( .A(n46586), .B(n46587), .Z(n46368) );
  NANDN U46934 ( .A(n46588), .B(n46589), .Z(n46587) );
  NANDN U46935 ( .A(n46590), .B(n46591), .Z(n46589) );
  NANDN U46936 ( .A(n46591), .B(n46590), .Z(n46586) );
  ANDN U46937 ( .B(B[111]), .A(n72), .Z(n46370) );
  XNOR U46938 ( .A(n46378), .B(n46592), .Z(n46371) );
  XNOR U46939 ( .A(n46377), .B(n46375), .Z(n46592) );
  AND U46940 ( .A(n46593), .B(n46594), .Z(n46375) );
  NANDN U46941 ( .A(n46595), .B(n46596), .Z(n46594) );
  OR U46942 ( .A(n46597), .B(n46598), .Z(n46596) );
  NAND U46943 ( .A(n46598), .B(n46597), .Z(n46593) );
  ANDN U46944 ( .B(B[112]), .A(n73), .Z(n46377) );
  XNOR U46945 ( .A(n46385), .B(n46599), .Z(n46378) );
  XNOR U46946 ( .A(n46384), .B(n46382), .Z(n46599) );
  AND U46947 ( .A(n46600), .B(n46601), .Z(n46382) );
  NANDN U46948 ( .A(n46602), .B(n46603), .Z(n46601) );
  NANDN U46949 ( .A(n46604), .B(n46605), .Z(n46603) );
  NANDN U46950 ( .A(n46605), .B(n46604), .Z(n46600) );
  ANDN U46951 ( .B(B[113]), .A(n74), .Z(n46384) );
  XNOR U46952 ( .A(n46392), .B(n46606), .Z(n46385) );
  XNOR U46953 ( .A(n46391), .B(n46389), .Z(n46606) );
  AND U46954 ( .A(n46607), .B(n46608), .Z(n46389) );
  NANDN U46955 ( .A(n46609), .B(n46610), .Z(n46608) );
  OR U46956 ( .A(n46611), .B(n46612), .Z(n46610) );
  NAND U46957 ( .A(n46612), .B(n46611), .Z(n46607) );
  ANDN U46958 ( .B(B[114]), .A(n75), .Z(n46391) );
  XNOR U46959 ( .A(n46399), .B(n46613), .Z(n46392) );
  XNOR U46960 ( .A(n46398), .B(n46396), .Z(n46613) );
  AND U46961 ( .A(n46614), .B(n46615), .Z(n46396) );
  NANDN U46962 ( .A(n46616), .B(n46617), .Z(n46615) );
  NANDN U46963 ( .A(n46618), .B(n46619), .Z(n46617) );
  NANDN U46964 ( .A(n46619), .B(n46618), .Z(n46614) );
  ANDN U46965 ( .B(B[115]), .A(n76), .Z(n46398) );
  XNOR U46966 ( .A(n46406), .B(n46620), .Z(n46399) );
  XNOR U46967 ( .A(n46405), .B(n46403), .Z(n46620) );
  AND U46968 ( .A(n46621), .B(n46622), .Z(n46403) );
  NANDN U46969 ( .A(n46623), .B(n46624), .Z(n46622) );
  OR U46970 ( .A(n46625), .B(n46626), .Z(n46624) );
  NAND U46971 ( .A(n46626), .B(n46625), .Z(n46621) );
  ANDN U46972 ( .B(B[116]), .A(n77), .Z(n46405) );
  XNOR U46973 ( .A(n46413), .B(n46627), .Z(n46406) );
  XNOR U46974 ( .A(n46412), .B(n46410), .Z(n46627) );
  AND U46975 ( .A(n46628), .B(n46629), .Z(n46410) );
  NANDN U46976 ( .A(n46630), .B(n46631), .Z(n46629) );
  NANDN U46977 ( .A(n46632), .B(n46633), .Z(n46631) );
  NANDN U46978 ( .A(n46633), .B(n46632), .Z(n46628) );
  ANDN U46979 ( .B(B[117]), .A(n78), .Z(n46412) );
  XNOR U46980 ( .A(n46420), .B(n46634), .Z(n46413) );
  XNOR U46981 ( .A(n46419), .B(n46417), .Z(n46634) );
  AND U46982 ( .A(n46635), .B(n46636), .Z(n46417) );
  NANDN U46983 ( .A(n46637), .B(n46638), .Z(n46636) );
  OR U46984 ( .A(n46639), .B(n46640), .Z(n46638) );
  NAND U46985 ( .A(n46640), .B(n46639), .Z(n46635) );
  ANDN U46986 ( .B(B[118]), .A(n79), .Z(n46419) );
  XNOR U46987 ( .A(n46427), .B(n46641), .Z(n46420) );
  XNOR U46988 ( .A(n46426), .B(n46424), .Z(n46641) );
  AND U46989 ( .A(n46642), .B(n46643), .Z(n46424) );
  NANDN U46990 ( .A(n46644), .B(n46645), .Z(n46643) );
  NANDN U46991 ( .A(n46646), .B(n46647), .Z(n46645) );
  NANDN U46992 ( .A(n46647), .B(n46646), .Z(n46642) );
  ANDN U46993 ( .B(B[119]), .A(n80), .Z(n46426) );
  XNOR U46994 ( .A(n46434), .B(n46648), .Z(n46427) );
  XNOR U46995 ( .A(n46433), .B(n46431), .Z(n46648) );
  AND U46996 ( .A(n46649), .B(n46650), .Z(n46431) );
  NANDN U46997 ( .A(n46651), .B(n46652), .Z(n46650) );
  OR U46998 ( .A(n46653), .B(n46654), .Z(n46652) );
  NAND U46999 ( .A(n46654), .B(n46653), .Z(n46649) );
  ANDN U47000 ( .B(B[120]), .A(n81), .Z(n46433) );
  XNOR U47001 ( .A(n46441), .B(n46655), .Z(n46434) );
  XNOR U47002 ( .A(n46440), .B(n46438), .Z(n46655) );
  AND U47003 ( .A(n46656), .B(n46657), .Z(n46438) );
  NANDN U47004 ( .A(n46658), .B(n46659), .Z(n46657) );
  NAND U47005 ( .A(n46660), .B(n46661), .Z(n46659) );
  ANDN U47006 ( .B(B[121]), .A(n82), .Z(n46440) );
  XOR U47007 ( .A(n46447), .B(n46662), .Z(n46441) );
  XNOR U47008 ( .A(n46445), .B(n46448), .Z(n46662) );
  NAND U47009 ( .A(A[2]), .B(B[122]), .Z(n46448) );
  NANDN U47010 ( .A(n46663), .B(n46664), .Z(n46445) );
  AND U47011 ( .A(A[0]), .B(B[123]), .Z(n46664) );
  XNOR U47012 ( .A(n46450), .B(n46665), .Z(n46447) );
  NAND U47013 ( .A(A[0]), .B(B[124]), .Z(n46665) );
  NAND U47014 ( .A(B[123]), .B(A[1]), .Z(n46450) );
  NAND U47015 ( .A(n46666), .B(n46667), .Z(n548) );
  NANDN U47016 ( .A(n46668), .B(n46669), .Z(n46667) );
  OR U47017 ( .A(n46670), .B(n46671), .Z(n46669) );
  NAND U47018 ( .A(n46671), .B(n46670), .Z(n46666) );
  XOR U47019 ( .A(n550), .B(n549), .Z(\A1[121] ) );
  XOR U47020 ( .A(n46671), .B(n46672), .Z(n549) );
  XNOR U47021 ( .A(n46670), .B(n46668), .Z(n46672) );
  AND U47022 ( .A(n46673), .B(n46674), .Z(n46668) );
  NANDN U47023 ( .A(n46675), .B(n46676), .Z(n46674) );
  NANDN U47024 ( .A(n46677), .B(n46678), .Z(n46676) );
  NANDN U47025 ( .A(n46678), .B(n46677), .Z(n46673) );
  ANDN U47026 ( .B(B[92]), .A(n54), .Z(n46670) );
  XNOR U47027 ( .A(n46465), .B(n46679), .Z(n46671) );
  XNOR U47028 ( .A(n46464), .B(n46462), .Z(n46679) );
  AND U47029 ( .A(n46680), .B(n46681), .Z(n46462) );
  NANDN U47030 ( .A(n46682), .B(n46683), .Z(n46681) );
  OR U47031 ( .A(n46684), .B(n46685), .Z(n46683) );
  NAND U47032 ( .A(n46685), .B(n46684), .Z(n46680) );
  ANDN U47033 ( .B(B[93]), .A(n55), .Z(n46464) );
  XNOR U47034 ( .A(n46472), .B(n46686), .Z(n46465) );
  XNOR U47035 ( .A(n46471), .B(n46469), .Z(n46686) );
  AND U47036 ( .A(n46687), .B(n46688), .Z(n46469) );
  NANDN U47037 ( .A(n46689), .B(n46690), .Z(n46688) );
  NANDN U47038 ( .A(n46691), .B(n46692), .Z(n46690) );
  NANDN U47039 ( .A(n46692), .B(n46691), .Z(n46687) );
  ANDN U47040 ( .B(B[94]), .A(n56), .Z(n46471) );
  XNOR U47041 ( .A(n46479), .B(n46693), .Z(n46472) );
  XNOR U47042 ( .A(n46478), .B(n46476), .Z(n46693) );
  AND U47043 ( .A(n46694), .B(n46695), .Z(n46476) );
  NANDN U47044 ( .A(n46696), .B(n46697), .Z(n46695) );
  OR U47045 ( .A(n46698), .B(n46699), .Z(n46697) );
  NAND U47046 ( .A(n46699), .B(n46698), .Z(n46694) );
  ANDN U47047 ( .B(B[95]), .A(n57), .Z(n46478) );
  XNOR U47048 ( .A(n46486), .B(n46700), .Z(n46479) );
  XNOR U47049 ( .A(n46485), .B(n46483), .Z(n46700) );
  AND U47050 ( .A(n46701), .B(n46702), .Z(n46483) );
  NANDN U47051 ( .A(n46703), .B(n46704), .Z(n46702) );
  NANDN U47052 ( .A(n46705), .B(n46706), .Z(n46704) );
  NANDN U47053 ( .A(n46706), .B(n46705), .Z(n46701) );
  ANDN U47054 ( .B(A[27]), .A(n11), .Z(n46485) );
  XNOR U47055 ( .A(n46493), .B(n46707), .Z(n46486) );
  XNOR U47056 ( .A(n46492), .B(n46490), .Z(n46707) );
  AND U47057 ( .A(n46708), .B(n46709), .Z(n46490) );
  NANDN U47058 ( .A(n46710), .B(n46711), .Z(n46709) );
  OR U47059 ( .A(n46712), .B(n46713), .Z(n46711) );
  NAND U47060 ( .A(n46713), .B(n46712), .Z(n46708) );
  ANDN U47061 ( .B(A[26]), .A(n9), .Z(n46492) );
  XNOR U47062 ( .A(n46500), .B(n46714), .Z(n46493) );
  XNOR U47063 ( .A(n46499), .B(n46497), .Z(n46714) );
  AND U47064 ( .A(n46715), .B(n46716), .Z(n46497) );
  NANDN U47065 ( .A(n46717), .B(n46718), .Z(n46716) );
  NANDN U47066 ( .A(n46719), .B(n46720), .Z(n46718) );
  NANDN U47067 ( .A(n46720), .B(n46719), .Z(n46715) );
  ANDN U47068 ( .B(B[98]), .A(n60), .Z(n46499) );
  XNOR U47069 ( .A(n46507), .B(n46721), .Z(n46500) );
  XNOR U47070 ( .A(n46506), .B(n46504), .Z(n46721) );
  AND U47071 ( .A(n46722), .B(n46723), .Z(n46504) );
  NANDN U47072 ( .A(n46724), .B(n46725), .Z(n46723) );
  OR U47073 ( .A(n46726), .B(n46727), .Z(n46725) );
  NAND U47074 ( .A(n46727), .B(n46726), .Z(n46722) );
  ANDN U47075 ( .B(A[24]), .A(n6), .Z(n46506) );
  XNOR U47076 ( .A(n46514), .B(n46728), .Z(n46507) );
  XNOR U47077 ( .A(n46513), .B(n46511), .Z(n46728) );
  AND U47078 ( .A(n46729), .B(n46730), .Z(n46511) );
  NANDN U47079 ( .A(n46731), .B(n46732), .Z(n46730) );
  NANDN U47080 ( .A(n46733), .B(n46734), .Z(n46732) );
  NANDN U47081 ( .A(n46734), .B(n46733), .Z(n46729) );
  ANDN U47082 ( .B(A[23]), .A(n4), .Z(n46513) );
  XNOR U47083 ( .A(n46521), .B(n46735), .Z(n46514) );
  XNOR U47084 ( .A(n46520), .B(n46518), .Z(n46735) );
  AND U47085 ( .A(n46736), .B(n46737), .Z(n46518) );
  NANDN U47086 ( .A(n46738), .B(n46739), .Z(n46737) );
  OR U47087 ( .A(n46740), .B(n46741), .Z(n46739) );
  NAND U47088 ( .A(n46741), .B(n46740), .Z(n46736) );
  ANDN U47089 ( .B(B[101]), .A(n63), .Z(n46520) );
  XNOR U47090 ( .A(n46528), .B(n46742), .Z(n46521) );
  XNOR U47091 ( .A(n46527), .B(n46525), .Z(n46742) );
  AND U47092 ( .A(n46743), .B(n46744), .Z(n46525) );
  NANDN U47093 ( .A(n46745), .B(n46746), .Z(n46744) );
  NANDN U47094 ( .A(n46747), .B(n46748), .Z(n46746) );
  NANDN U47095 ( .A(n46748), .B(n46747), .Z(n46743) );
  ANDN U47096 ( .B(B[102]), .A(n64), .Z(n46527) );
  XNOR U47097 ( .A(n46535), .B(n46749), .Z(n46528) );
  XNOR U47098 ( .A(n46534), .B(n46532), .Z(n46749) );
  AND U47099 ( .A(n46750), .B(n46751), .Z(n46532) );
  NANDN U47100 ( .A(n46752), .B(n46753), .Z(n46751) );
  OR U47101 ( .A(n46754), .B(n46755), .Z(n46753) );
  NAND U47102 ( .A(n46755), .B(n46754), .Z(n46750) );
  ANDN U47103 ( .B(B[103]), .A(n65), .Z(n46534) );
  XNOR U47104 ( .A(n46542), .B(n46756), .Z(n46535) );
  XNOR U47105 ( .A(n46541), .B(n46539), .Z(n46756) );
  AND U47106 ( .A(n46757), .B(n46758), .Z(n46539) );
  NANDN U47107 ( .A(n46759), .B(n46760), .Z(n46758) );
  NANDN U47108 ( .A(n46761), .B(n46762), .Z(n46760) );
  NANDN U47109 ( .A(n46762), .B(n46761), .Z(n46757) );
  ANDN U47110 ( .B(B[104]), .A(n66), .Z(n46541) );
  XNOR U47111 ( .A(n46549), .B(n46763), .Z(n46542) );
  XNOR U47112 ( .A(n46548), .B(n46546), .Z(n46763) );
  AND U47113 ( .A(n46764), .B(n46765), .Z(n46546) );
  NANDN U47114 ( .A(n46766), .B(n46767), .Z(n46765) );
  OR U47115 ( .A(n46768), .B(n46769), .Z(n46767) );
  NAND U47116 ( .A(n46769), .B(n46768), .Z(n46764) );
  ANDN U47117 ( .B(B[105]), .A(n67), .Z(n46548) );
  XNOR U47118 ( .A(n46556), .B(n46770), .Z(n46549) );
  XNOR U47119 ( .A(n46555), .B(n46553), .Z(n46770) );
  AND U47120 ( .A(n46771), .B(n46772), .Z(n46553) );
  NANDN U47121 ( .A(n46773), .B(n46774), .Z(n46772) );
  NANDN U47122 ( .A(n46775), .B(n46776), .Z(n46774) );
  NANDN U47123 ( .A(n46776), .B(n46775), .Z(n46771) );
  ANDN U47124 ( .B(B[106]), .A(n68), .Z(n46555) );
  XNOR U47125 ( .A(n46563), .B(n46777), .Z(n46556) );
  XNOR U47126 ( .A(n46562), .B(n46560), .Z(n46777) );
  AND U47127 ( .A(n46778), .B(n46779), .Z(n46560) );
  NANDN U47128 ( .A(n46780), .B(n46781), .Z(n46779) );
  OR U47129 ( .A(n46782), .B(n46783), .Z(n46781) );
  NAND U47130 ( .A(n46783), .B(n46782), .Z(n46778) );
  ANDN U47131 ( .B(B[107]), .A(n69), .Z(n46562) );
  XNOR U47132 ( .A(n46570), .B(n46784), .Z(n46563) );
  XNOR U47133 ( .A(n46569), .B(n46567), .Z(n46784) );
  AND U47134 ( .A(n46785), .B(n46786), .Z(n46567) );
  NANDN U47135 ( .A(n46787), .B(n46788), .Z(n46786) );
  NANDN U47136 ( .A(n46789), .B(n46790), .Z(n46788) );
  NANDN U47137 ( .A(n46790), .B(n46789), .Z(n46785) );
  ANDN U47138 ( .B(B[108]), .A(n70), .Z(n46569) );
  XNOR U47139 ( .A(n46577), .B(n46791), .Z(n46570) );
  XNOR U47140 ( .A(n46576), .B(n46574), .Z(n46791) );
  AND U47141 ( .A(n46792), .B(n46793), .Z(n46574) );
  NANDN U47142 ( .A(n46794), .B(n46795), .Z(n46793) );
  OR U47143 ( .A(n46796), .B(n46797), .Z(n46795) );
  NAND U47144 ( .A(n46797), .B(n46796), .Z(n46792) );
  ANDN U47145 ( .B(B[109]), .A(n71), .Z(n46576) );
  XNOR U47146 ( .A(n46584), .B(n46798), .Z(n46577) );
  XNOR U47147 ( .A(n46583), .B(n46581), .Z(n46798) );
  AND U47148 ( .A(n46799), .B(n46800), .Z(n46581) );
  NANDN U47149 ( .A(n46801), .B(n46802), .Z(n46800) );
  NANDN U47150 ( .A(n46803), .B(n46804), .Z(n46802) );
  NANDN U47151 ( .A(n46804), .B(n46803), .Z(n46799) );
  ANDN U47152 ( .B(B[110]), .A(n72), .Z(n46583) );
  XNOR U47153 ( .A(n46591), .B(n46805), .Z(n46584) );
  XNOR U47154 ( .A(n46590), .B(n46588), .Z(n46805) );
  AND U47155 ( .A(n46806), .B(n46807), .Z(n46588) );
  NANDN U47156 ( .A(n46808), .B(n46809), .Z(n46807) );
  OR U47157 ( .A(n46810), .B(n46811), .Z(n46809) );
  NAND U47158 ( .A(n46811), .B(n46810), .Z(n46806) );
  ANDN U47159 ( .B(B[111]), .A(n73), .Z(n46590) );
  XNOR U47160 ( .A(n46598), .B(n46812), .Z(n46591) );
  XNOR U47161 ( .A(n46597), .B(n46595), .Z(n46812) );
  AND U47162 ( .A(n46813), .B(n46814), .Z(n46595) );
  NANDN U47163 ( .A(n46815), .B(n46816), .Z(n46814) );
  NANDN U47164 ( .A(n46817), .B(n46818), .Z(n46816) );
  NANDN U47165 ( .A(n46818), .B(n46817), .Z(n46813) );
  ANDN U47166 ( .B(B[112]), .A(n74), .Z(n46597) );
  XNOR U47167 ( .A(n46605), .B(n46819), .Z(n46598) );
  XNOR U47168 ( .A(n46604), .B(n46602), .Z(n46819) );
  AND U47169 ( .A(n46820), .B(n46821), .Z(n46602) );
  NANDN U47170 ( .A(n46822), .B(n46823), .Z(n46821) );
  OR U47171 ( .A(n46824), .B(n46825), .Z(n46823) );
  NAND U47172 ( .A(n46825), .B(n46824), .Z(n46820) );
  ANDN U47173 ( .B(B[113]), .A(n75), .Z(n46604) );
  XNOR U47174 ( .A(n46612), .B(n46826), .Z(n46605) );
  XNOR U47175 ( .A(n46611), .B(n46609), .Z(n46826) );
  AND U47176 ( .A(n46827), .B(n46828), .Z(n46609) );
  NANDN U47177 ( .A(n46829), .B(n46830), .Z(n46828) );
  NANDN U47178 ( .A(n46831), .B(n46832), .Z(n46830) );
  NANDN U47179 ( .A(n46832), .B(n46831), .Z(n46827) );
  ANDN U47180 ( .B(B[114]), .A(n76), .Z(n46611) );
  XNOR U47181 ( .A(n46619), .B(n46833), .Z(n46612) );
  XNOR U47182 ( .A(n46618), .B(n46616), .Z(n46833) );
  AND U47183 ( .A(n46834), .B(n46835), .Z(n46616) );
  NANDN U47184 ( .A(n46836), .B(n46837), .Z(n46835) );
  OR U47185 ( .A(n46838), .B(n46839), .Z(n46837) );
  NAND U47186 ( .A(n46839), .B(n46838), .Z(n46834) );
  ANDN U47187 ( .B(B[115]), .A(n77), .Z(n46618) );
  XNOR U47188 ( .A(n46626), .B(n46840), .Z(n46619) );
  XNOR U47189 ( .A(n46625), .B(n46623), .Z(n46840) );
  AND U47190 ( .A(n46841), .B(n46842), .Z(n46623) );
  NANDN U47191 ( .A(n46843), .B(n46844), .Z(n46842) );
  NANDN U47192 ( .A(n46845), .B(n46846), .Z(n46844) );
  NANDN U47193 ( .A(n46846), .B(n46845), .Z(n46841) );
  ANDN U47194 ( .B(B[116]), .A(n78), .Z(n46625) );
  XNOR U47195 ( .A(n46633), .B(n46847), .Z(n46626) );
  XNOR U47196 ( .A(n46632), .B(n46630), .Z(n46847) );
  AND U47197 ( .A(n46848), .B(n46849), .Z(n46630) );
  NANDN U47198 ( .A(n46850), .B(n46851), .Z(n46849) );
  OR U47199 ( .A(n46852), .B(n46853), .Z(n46851) );
  NAND U47200 ( .A(n46853), .B(n46852), .Z(n46848) );
  ANDN U47201 ( .B(B[117]), .A(n79), .Z(n46632) );
  XNOR U47202 ( .A(n46640), .B(n46854), .Z(n46633) );
  XNOR U47203 ( .A(n46639), .B(n46637), .Z(n46854) );
  AND U47204 ( .A(n46855), .B(n46856), .Z(n46637) );
  NANDN U47205 ( .A(n46857), .B(n46858), .Z(n46856) );
  NANDN U47206 ( .A(n46859), .B(n46860), .Z(n46858) );
  NANDN U47207 ( .A(n46860), .B(n46859), .Z(n46855) );
  ANDN U47208 ( .B(B[118]), .A(n80), .Z(n46639) );
  XNOR U47209 ( .A(n46647), .B(n46861), .Z(n46640) );
  XNOR U47210 ( .A(n46646), .B(n46644), .Z(n46861) );
  AND U47211 ( .A(n46862), .B(n46863), .Z(n46644) );
  NANDN U47212 ( .A(n46864), .B(n46865), .Z(n46863) );
  OR U47213 ( .A(n46866), .B(n46867), .Z(n46865) );
  NAND U47214 ( .A(n46867), .B(n46866), .Z(n46862) );
  ANDN U47215 ( .B(B[119]), .A(n81), .Z(n46646) );
  XNOR U47216 ( .A(n46654), .B(n46868), .Z(n46647) );
  XNOR U47217 ( .A(n46653), .B(n46651), .Z(n46868) );
  AND U47218 ( .A(n46869), .B(n46870), .Z(n46651) );
  NANDN U47219 ( .A(n46871), .B(n46872), .Z(n46870) );
  NAND U47220 ( .A(n46873), .B(n46874), .Z(n46872) );
  ANDN U47221 ( .B(B[120]), .A(n82), .Z(n46653) );
  XOR U47222 ( .A(n46660), .B(n46875), .Z(n46654) );
  XNOR U47223 ( .A(n46658), .B(n46661), .Z(n46875) );
  NAND U47224 ( .A(A[2]), .B(B[121]), .Z(n46661) );
  NANDN U47225 ( .A(n46876), .B(n46877), .Z(n46658) );
  AND U47226 ( .A(A[0]), .B(B[122]), .Z(n46877) );
  XNOR U47227 ( .A(n46663), .B(n46878), .Z(n46660) );
  NAND U47228 ( .A(A[0]), .B(B[123]), .Z(n46878) );
  NAND U47229 ( .A(B[122]), .B(A[1]), .Z(n46663) );
  NAND U47230 ( .A(n46879), .B(n46880), .Z(n550) );
  NANDN U47231 ( .A(n46881), .B(n46882), .Z(n46880) );
  OR U47232 ( .A(n46883), .B(n46884), .Z(n46882) );
  NAND U47233 ( .A(n46884), .B(n46883), .Z(n46879) );
  XOR U47234 ( .A(n552), .B(n551), .Z(\A1[120] ) );
  XOR U47235 ( .A(n46884), .B(n46885), .Z(n551) );
  XNOR U47236 ( .A(n46883), .B(n46881), .Z(n46885) );
  AND U47237 ( .A(n46886), .B(n46887), .Z(n46881) );
  NANDN U47238 ( .A(n46888), .B(n46889), .Z(n46887) );
  NANDN U47239 ( .A(n46890), .B(n46891), .Z(n46889) );
  NANDN U47240 ( .A(n46891), .B(n46890), .Z(n46886) );
  ANDN U47241 ( .B(B[91]), .A(n54), .Z(n46883) );
  XNOR U47242 ( .A(n46678), .B(n46892), .Z(n46884) );
  XNOR U47243 ( .A(n46677), .B(n46675), .Z(n46892) );
  AND U47244 ( .A(n46893), .B(n46894), .Z(n46675) );
  NANDN U47245 ( .A(n46895), .B(n46896), .Z(n46894) );
  OR U47246 ( .A(n46897), .B(n46898), .Z(n46896) );
  NAND U47247 ( .A(n46898), .B(n46897), .Z(n46893) );
  ANDN U47248 ( .B(B[92]), .A(n55), .Z(n46677) );
  XNOR U47249 ( .A(n46685), .B(n46899), .Z(n46678) );
  XNOR U47250 ( .A(n46684), .B(n46682), .Z(n46899) );
  AND U47251 ( .A(n46900), .B(n46901), .Z(n46682) );
  NANDN U47252 ( .A(n46902), .B(n46903), .Z(n46901) );
  NANDN U47253 ( .A(n46904), .B(n46905), .Z(n46903) );
  NANDN U47254 ( .A(n46905), .B(n46904), .Z(n46900) );
  ANDN U47255 ( .B(B[93]), .A(n56), .Z(n46684) );
  XNOR U47256 ( .A(n46692), .B(n46906), .Z(n46685) );
  XNOR U47257 ( .A(n46691), .B(n46689), .Z(n46906) );
  AND U47258 ( .A(n46907), .B(n46908), .Z(n46689) );
  NANDN U47259 ( .A(n46909), .B(n46910), .Z(n46908) );
  OR U47260 ( .A(n46911), .B(n46912), .Z(n46910) );
  NAND U47261 ( .A(n46912), .B(n46911), .Z(n46907) );
  ANDN U47262 ( .B(B[94]), .A(n57), .Z(n46691) );
  XNOR U47263 ( .A(n46699), .B(n46913), .Z(n46692) );
  XNOR U47264 ( .A(n46698), .B(n46696), .Z(n46913) );
  AND U47265 ( .A(n46914), .B(n46915), .Z(n46696) );
  NANDN U47266 ( .A(n46916), .B(n46917), .Z(n46915) );
  NANDN U47267 ( .A(n46918), .B(n46919), .Z(n46917) );
  NANDN U47268 ( .A(n46919), .B(n46918), .Z(n46914) );
  ANDN U47269 ( .B(A[27]), .A(n13), .Z(n46698) );
  XNOR U47270 ( .A(n46706), .B(n46920), .Z(n46699) );
  XNOR U47271 ( .A(n46705), .B(n46703), .Z(n46920) );
  AND U47272 ( .A(n46921), .B(n46922), .Z(n46703) );
  NANDN U47273 ( .A(n46923), .B(n46924), .Z(n46922) );
  OR U47274 ( .A(n46925), .B(n46926), .Z(n46924) );
  NAND U47275 ( .A(n46926), .B(n46925), .Z(n46921) );
  ANDN U47276 ( .B(A[26]), .A(n11), .Z(n46705) );
  XNOR U47277 ( .A(n46713), .B(n46927), .Z(n46706) );
  XNOR U47278 ( .A(n46712), .B(n46710), .Z(n46927) );
  AND U47279 ( .A(n46928), .B(n46929), .Z(n46710) );
  NANDN U47280 ( .A(n46930), .B(n46931), .Z(n46929) );
  NANDN U47281 ( .A(n46932), .B(n46933), .Z(n46931) );
  NANDN U47282 ( .A(n46933), .B(n46932), .Z(n46928) );
  ANDN U47283 ( .B(A[25]), .A(n9), .Z(n46712) );
  XNOR U47284 ( .A(n46720), .B(n46934), .Z(n46713) );
  XNOR U47285 ( .A(n46719), .B(n46717), .Z(n46934) );
  AND U47286 ( .A(n46935), .B(n46936), .Z(n46717) );
  NANDN U47287 ( .A(n46937), .B(n46938), .Z(n46936) );
  OR U47288 ( .A(n46939), .B(n46940), .Z(n46938) );
  NAND U47289 ( .A(n46940), .B(n46939), .Z(n46935) );
  ANDN U47290 ( .B(B[98]), .A(n61), .Z(n46719) );
  XNOR U47291 ( .A(n46727), .B(n46941), .Z(n46720) );
  XNOR U47292 ( .A(n46726), .B(n46724), .Z(n46941) );
  AND U47293 ( .A(n46942), .B(n46943), .Z(n46724) );
  NANDN U47294 ( .A(n46944), .B(n46945), .Z(n46943) );
  NANDN U47295 ( .A(n46946), .B(n46947), .Z(n46945) );
  NANDN U47296 ( .A(n46947), .B(n46946), .Z(n46942) );
  ANDN U47297 ( .B(A[23]), .A(n6), .Z(n46726) );
  XNOR U47298 ( .A(n46734), .B(n46948), .Z(n46727) );
  XNOR U47299 ( .A(n46733), .B(n46731), .Z(n46948) );
  AND U47300 ( .A(n46949), .B(n46950), .Z(n46731) );
  NANDN U47301 ( .A(n46951), .B(n46952), .Z(n46950) );
  OR U47302 ( .A(n46953), .B(n46954), .Z(n46952) );
  NAND U47303 ( .A(n46954), .B(n46953), .Z(n46949) );
  ANDN U47304 ( .B(A[22]), .A(n4), .Z(n46733) );
  XNOR U47305 ( .A(n46741), .B(n46955), .Z(n46734) );
  XNOR U47306 ( .A(n46740), .B(n46738), .Z(n46955) );
  AND U47307 ( .A(n46956), .B(n46957), .Z(n46738) );
  NANDN U47308 ( .A(n46958), .B(n46959), .Z(n46957) );
  NANDN U47309 ( .A(n46960), .B(n46961), .Z(n46959) );
  NANDN U47310 ( .A(n46961), .B(n46960), .Z(n46956) );
  ANDN U47311 ( .B(B[101]), .A(n64), .Z(n46740) );
  XNOR U47312 ( .A(n46748), .B(n46962), .Z(n46741) );
  XNOR U47313 ( .A(n46747), .B(n46745), .Z(n46962) );
  AND U47314 ( .A(n46963), .B(n46964), .Z(n46745) );
  NANDN U47315 ( .A(n46965), .B(n46966), .Z(n46964) );
  OR U47316 ( .A(n46967), .B(n46968), .Z(n46966) );
  NAND U47317 ( .A(n46968), .B(n46967), .Z(n46963) );
  ANDN U47318 ( .B(B[102]), .A(n65), .Z(n46747) );
  XNOR U47319 ( .A(n46755), .B(n46969), .Z(n46748) );
  XNOR U47320 ( .A(n46754), .B(n46752), .Z(n46969) );
  AND U47321 ( .A(n46970), .B(n46971), .Z(n46752) );
  NANDN U47322 ( .A(n46972), .B(n46973), .Z(n46971) );
  NANDN U47323 ( .A(n46974), .B(n46975), .Z(n46973) );
  NANDN U47324 ( .A(n46975), .B(n46974), .Z(n46970) );
  ANDN U47325 ( .B(B[103]), .A(n66), .Z(n46754) );
  XNOR U47326 ( .A(n46762), .B(n46976), .Z(n46755) );
  XNOR U47327 ( .A(n46761), .B(n46759), .Z(n46976) );
  AND U47328 ( .A(n46977), .B(n46978), .Z(n46759) );
  NANDN U47329 ( .A(n46979), .B(n46980), .Z(n46978) );
  OR U47330 ( .A(n46981), .B(n46982), .Z(n46980) );
  NAND U47331 ( .A(n46982), .B(n46981), .Z(n46977) );
  ANDN U47332 ( .B(B[104]), .A(n67), .Z(n46761) );
  XNOR U47333 ( .A(n46769), .B(n46983), .Z(n46762) );
  XNOR U47334 ( .A(n46768), .B(n46766), .Z(n46983) );
  AND U47335 ( .A(n46984), .B(n46985), .Z(n46766) );
  NANDN U47336 ( .A(n46986), .B(n46987), .Z(n46985) );
  NANDN U47337 ( .A(n46988), .B(n46989), .Z(n46987) );
  NANDN U47338 ( .A(n46989), .B(n46988), .Z(n46984) );
  ANDN U47339 ( .B(B[105]), .A(n68), .Z(n46768) );
  XNOR U47340 ( .A(n46776), .B(n46990), .Z(n46769) );
  XNOR U47341 ( .A(n46775), .B(n46773), .Z(n46990) );
  AND U47342 ( .A(n46991), .B(n46992), .Z(n46773) );
  NANDN U47343 ( .A(n46993), .B(n46994), .Z(n46992) );
  OR U47344 ( .A(n46995), .B(n46996), .Z(n46994) );
  NAND U47345 ( .A(n46996), .B(n46995), .Z(n46991) );
  ANDN U47346 ( .B(B[106]), .A(n69), .Z(n46775) );
  XNOR U47347 ( .A(n46783), .B(n46997), .Z(n46776) );
  XNOR U47348 ( .A(n46782), .B(n46780), .Z(n46997) );
  AND U47349 ( .A(n46998), .B(n46999), .Z(n46780) );
  NANDN U47350 ( .A(n47000), .B(n47001), .Z(n46999) );
  NANDN U47351 ( .A(n47002), .B(n47003), .Z(n47001) );
  NANDN U47352 ( .A(n47003), .B(n47002), .Z(n46998) );
  ANDN U47353 ( .B(B[107]), .A(n70), .Z(n46782) );
  XNOR U47354 ( .A(n46790), .B(n47004), .Z(n46783) );
  XNOR U47355 ( .A(n46789), .B(n46787), .Z(n47004) );
  AND U47356 ( .A(n47005), .B(n47006), .Z(n46787) );
  NANDN U47357 ( .A(n47007), .B(n47008), .Z(n47006) );
  OR U47358 ( .A(n47009), .B(n47010), .Z(n47008) );
  NAND U47359 ( .A(n47010), .B(n47009), .Z(n47005) );
  ANDN U47360 ( .B(B[108]), .A(n71), .Z(n46789) );
  XNOR U47361 ( .A(n46797), .B(n47011), .Z(n46790) );
  XNOR U47362 ( .A(n46796), .B(n46794), .Z(n47011) );
  AND U47363 ( .A(n47012), .B(n47013), .Z(n46794) );
  NANDN U47364 ( .A(n47014), .B(n47015), .Z(n47013) );
  NANDN U47365 ( .A(n47016), .B(n47017), .Z(n47015) );
  NANDN U47366 ( .A(n47017), .B(n47016), .Z(n47012) );
  ANDN U47367 ( .B(B[109]), .A(n72), .Z(n46796) );
  XNOR U47368 ( .A(n46804), .B(n47018), .Z(n46797) );
  XNOR U47369 ( .A(n46803), .B(n46801), .Z(n47018) );
  AND U47370 ( .A(n47019), .B(n47020), .Z(n46801) );
  NANDN U47371 ( .A(n47021), .B(n47022), .Z(n47020) );
  OR U47372 ( .A(n47023), .B(n47024), .Z(n47022) );
  NAND U47373 ( .A(n47024), .B(n47023), .Z(n47019) );
  ANDN U47374 ( .B(B[110]), .A(n73), .Z(n46803) );
  XNOR U47375 ( .A(n46811), .B(n47025), .Z(n46804) );
  XNOR U47376 ( .A(n46810), .B(n46808), .Z(n47025) );
  AND U47377 ( .A(n47026), .B(n47027), .Z(n46808) );
  NANDN U47378 ( .A(n47028), .B(n47029), .Z(n47027) );
  NANDN U47379 ( .A(n47030), .B(n47031), .Z(n47029) );
  NANDN U47380 ( .A(n47031), .B(n47030), .Z(n47026) );
  ANDN U47381 ( .B(B[111]), .A(n74), .Z(n46810) );
  XNOR U47382 ( .A(n46818), .B(n47032), .Z(n46811) );
  XNOR U47383 ( .A(n46817), .B(n46815), .Z(n47032) );
  AND U47384 ( .A(n47033), .B(n47034), .Z(n46815) );
  NANDN U47385 ( .A(n47035), .B(n47036), .Z(n47034) );
  OR U47386 ( .A(n47037), .B(n47038), .Z(n47036) );
  NAND U47387 ( .A(n47038), .B(n47037), .Z(n47033) );
  ANDN U47388 ( .B(B[112]), .A(n75), .Z(n46817) );
  XNOR U47389 ( .A(n46825), .B(n47039), .Z(n46818) );
  XNOR U47390 ( .A(n46824), .B(n46822), .Z(n47039) );
  AND U47391 ( .A(n47040), .B(n47041), .Z(n46822) );
  NANDN U47392 ( .A(n47042), .B(n47043), .Z(n47041) );
  NANDN U47393 ( .A(n47044), .B(n47045), .Z(n47043) );
  NANDN U47394 ( .A(n47045), .B(n47044), .Z(n47040) );
  ANDN U47395 ( .B(B[113]), .A(n76), .Z(n46824) );
  XNOR U47396 ( .A(n46832), .B(n47046), .Z(n46825) );
  XNOR U47397 ( .A(n46831), .B(n46829), .Z(n47046) );
  AND U47398 ( .A(n47047), .B(n47048), .Z(n46829) );
  NANDN U47399 ( .A(n47049), .B(n47050), .Z(n47048) );
  OR U47400 ( .A(n47051), .B(n47052), .Z(n47050) );
  NAND U47401 ( .A(n47052), .B(n47051), .Z(n47047) );
  ANDN U47402 ( .B(B[114]), .A(n77), .Z(n46831) );
  XNOR U47403 ( .A(n46839), .B(n47053), .Z(n46832) );
  XNOR U47404 ( .A(n46838), .B(n46836), .Z(n47053) );
  AND U47405 ( .A(n47054), .B(n47055), .Z(n46836) );
  NANDN U47406 ( .A(n47056), .B(n47057), .Z(n47055) );
  NANDN U47407 ( .A(n47058), .B(n47059), .Z(n47057) );
  NANDN U47408 ( .A(n47059), .B(n47058), .Z(n47054) );
  ANDN U47409 ( .B(B[115]), .A(n78), .Z(n46838) );
  XNOR U47410 ( .A(n46846), .B(n47060), .Z(n46839) );
  XNOR U47411 ( .A(n46845), .B(n46843), .Z(n47060) );
  AND U47412 ( .A(n47061), .B(n47062), .Z(n46843) );
  NANDN U47413 ( .A(n47063), .B(n47064), .Z(n47062) );
  OR U47414 ( .A(n47065), .B(n47066), .Z(n47064) );
  NAND U47415 ( .A(n47066), .B(n47065), .Z(n47061) );
  ANDN U47416 ( .B(B[116]), .A(n79), .Z(n46845) );
  XNOR U47417 ( .A(n46853), .B(n47067), .Z(n46846) );
  XNOR U47418 ( .A(n46852), .B(n46850), .Z(n47067) );
  AND U47419 ( .A(n47068), .B(n47069), .Z(n46850) );
  NANDN U47420 ( .A(n47070), .B(n47071), .Z(n47069) );
  NANDN U47421 ( .A(n47072), .B(n47073), .Z(n47071) );
  NANDN U47422 ( .A(n47073), .B(n47072), .Z(n47068) );
  ANDN U47423 ( .B(B[117]), .A(n80), .Z(n46852) );
  XNOR U47424 ( .A(n46860), .B(n47074), .Z(n46853) );
  XNOR U47425 ( .A(n46859), .B(n46857), .Z(n47074) );
  AND U47426 ( .A(n47075), .B(n47076), .Z(n46857) );
  NANDN U47427 ( .A(n47077), .B(n47078), .Z(n47076) );
  OR U47428 ( .A(n47079), .B(n47080), .Z(n47078) );
  NAND U47429 ( .A(n47080), .B(n47079), .Z(n47075) );
  ANDN U47430 ( .B(B[118]), .A(n81), .Z(n46859) );
  XNOR U47431 ( .A(n46867), .B(n47081), .Z(n46860) );
  XNOR U47432 ( .A(n46866), .B(n46864), .Z(n47081) );
  AND U47433 ( .A(n47082), .B(n47083), .Z(n46864) );
  NANDN U47434 ( .A(n47084), .B(n47085), .Z(n47083) );
  NAND U47435 ( .A(n47086), .B(n47087), .Z(n47085) );
  ANDN U47436 ( .B(B[119]), .A(n82), .Z(n46866) );
  XOR U47437 ( .A(n46873), .B(n47088), .Z(n46867) );
  XNOR U47438 ( .A(n46871), .B(n46874), .Z(n47088) );
  NAND U47439 ( .A(A[2]), .B(B[120]), .Z(n46874) );
  NANDN U47440 ( .A(n47089), .B(n47090), .Z(n46871) );
  AND U47441 ( .A(A[0]), .B(B[121]), .Z(n47090) );
  XNOR U47442 ( .A(n46876), .B(n47091), .Z(n46873) );
  NAND U47443 ( .A(A[0]), .B(B[122]), .Z(n47091) );
  NAND U47444 ( .A(B[121]), .B(A[1]), .Z(n46876) );
  NAND U47445 ( .A(n47092), .B(n47093), .Z(n552) );
  NANDN U47446 ( .A(n47094), .B(n47095), .Z(n47093) );
  OR U47447 ( .A(n47096), .B(n47097), .Z(n47095) );
  NAND U47448 ( .A(n47097), .B(n47096), .Z(n47092) );
  XOR U47449 ( .A(n44886), .B(n47098), .Z(\A1[11] ) );
  XNOR U47450 ( .A(n44885), .B(n44883), .Z(n47098) );
  AND U47451 ( .A(n47099), .B(n47100), .Z(n44883) );
  NANDN U47452 ( .A(n47101), .B(n47102), .Z(n47100) );
  NANDN U47453 ( .A(n47103), .B(n47104), .Z(n47102) );
  NANDN U47454 ( .A(n47104), .B(n47103), .Z(n47099) );
  ANDN U47455 ( .B(B[0]), .A(n72), .Z(n44885) );
  XNOR U47456 ( .A(n44893), .B(n47105), .Z(n44886) );
  XNOR U47457 ( .A(n44892), .B(n44890), .Z(n47105) );
  AND U47458 ( .A(n47106), .B(n47107), .Z(n44890) );
  NANDN U47459 ( .A(n47108), .B(n47109), .Z(n47107) );
  OR U47460 ( .A(n47110), .B(n47111), .Z(n47109) );
  NAND U47461 ( .A(n47111), .B(n47110), .Z(n47106) );
  ANDN U47462 ( .B(B[1]), .A(n73), .Z(n44892) );
  XNOR U47463 ( .A(n44900), .B(n47112), .Z(n44893) );
  XNOR U47464 ( .A(n44899), .B(n44897), .Z(n47112) );
  AND U47465 ( .A(n47113), .B(n47114), .Z(n44897) );
  NANDN U47466 ( .A(n47115), .B(n47116), .Z(n47114) );
  NANDN U47467 ( .A(n47117), .B(n47118), .Z(n47116) );
  NANDN U47468 ( .A(n47118), .B(n47117), .Z(n47113) );
  ANDN U47469 ( .B(B[2]), .A(n74), .Z(n44899) );
  XNOR U47470 ( .A(n44907), .B(n47119), .Z(n44900) );
  XNOR U47471 ( .A(n44906), .B(n44904), .Z(n47119) );
  AND U47472 ( .A(n47120), .B(n47121), .Z(n44904) );
  NANDN U47473 ( .A(n47122), .B(n47123), .Z(n47121) );
  OR U47474 ( .A(n47124), .B(n47125), .Z(n47123) );
  NAND U47475 ( .A(n47125), .B(n47124), .Z(n47120) );
  ANDN U47476 ( .B(B[3]), .A(n75), .Z(n44906) );
  XNOR U47477 ( .A(n44914), .B(n47126), .Z(n44907) );
  XNOR U47478 ( .A(n44913), .B(n44911), .Z(n47126) );
  AND U47479 ( .A(n47127), .B(n47128), .Z(n44911) );
  NANDN U47480 ( .A(n47129), .B(n47130), .Z(n47128) );
  NANDN U47481 ( .A(n47131), .B(n47132), .Z(n47130) );
  NANDN U47482 ( .A(n47132), .B(n47131), .Z(n47127) );
  ANDN U47483 ( .B(B[4]), .A(n76), .Z(n44913) );
  XNOR U47484 ( .A(n44921), .B(n47133), .Z(n44914) );
  XNOR U47485 ( .A(n44920), .B(n44918), .Z(n47133) );
  AND U47486 ( .A(n47134), .B(n47135), .Z(n44918) );
  NANDN U47487 ( .A(n47136), .B(n47137), .Z(n47135) );
  OR U47488 ( .A(n47138), .B(n47139), .Z(n47137) );
  NAND U47489 ( .A(n47139), .B(n47138), .Z(n47134) );
  ANDN U47490 ( .B(B[5]), .A(n77), .Z(n44920) );
  XNOR U47491 ( .A(n44928), .B(n47140), .Z(n44921) );
  XNOR U47492 ( .A(n44927), .B(n44925), .Z(n47140) );
  AND U47493 ( .A(n47141), .B(n47142), .Z(n44925) );
  NANDN U47494 ( .A(n47143), .B(n47144), .Z(n47142) );
  NANDN U47495 ( .A(n47145), .B(n47146), .Z(n47144) );
  NANDN U47496 ( .A(n47146), .B(n47145), .Z(n47141) );
  ANDN U47497 ( .B(B[6]), .A(n78), .Z(n44927) );
  XNOR U47498 ( .A(n44935), .B(n47147), .Z(n44928) );
  XNOR U47499 ( .A(n44934), .B(n44932), .Z(n47147) );
  AND U47500 ( .A(n47148), .B(n47149), .Z(n44932) );
  NANDN U47501 ( .A(n47150), .B(n47151), .Z(n47149) );
  OR U47502 ( .A(n47152), .B(n47153), .Z(n47151) );
  NAND U47503 ( .A(n47153), .B(n47152), .Z(n47148) );
  ANDN U47504 ( .B(B[7]), .A(n79), .Z(n44934) );
  XNOR U47505 ( .A(n44942), .B(n47154), .Z(n44935) );
  XNOR U47506 ( .A(n44941), .B(n44939), .Z(n47154) );
  AND U47507 ( .A(n47155), .B(n47156), .Z(n44939) );
  NANDN U47508 ( .A(n47157), .B(n47158), .Z(n47156) );
  NANDN U47509 ( .A(n47159), .B(n47160), .Z(n47158) );
  NANDN U47510 ( .A(n47160), .B(n47159), .Z(n47155) );
  ANDN U47511 ( .B(B[8]), .A(n80), .Z(n44941) );
  XNOR U47512 ( .A(n44949), .B(n47161), .Z(n44942) );
  XNOR U47513 ( .A(n44948), .B(n44946), .Z(n47161) );
  AND U47514 ( .A(n47162), .B(n47163), .Z(n44946) );
  NANDN U47515 ( .A(n47164), .B(n47165), .Z(n47163) );
  OR U47516 ( .A(n47166), .B(n47167), .Z(n47165) );
  NAND U47517 ( .A(n47167), .B(n47166), .Z(n47162) );
  ANDN U47518 ( .B(B[9]), .A(n81), .Z(n44948) );
  XNOR U47519 ( .A(n44956), .B(n47168), .Z(n44949) );
  XNOR U47520 ( .A(n44955), .B(n44953), .Z(n47168) );
  AND U47521 ( .A(n47169), .B(n47170), .Z(n44953) );
  NANDN U47522 ( .A(n47171), .B(n47172), .Z(n47170) );
  NAND U47523 ( .A(n47173), .B(n47174), .Z(n47172) );
  ANDN U47524 ( .B(B[10]), .A(n82), .Z(n44955) );
  XOR U47525 ( .A(n44962), .B(n47175), .Z(n44956) );
  XNOR U47526 ( .A(n44960), .B(n44963), .Z(n47175) );
  NAND U47527 ( .A(A[2]), .B(B[11]), .Z(n44963) );
  NANDN U47528 ( .A(n47176), .B(n47177), .Z(n44960) );
  AND U47529 ( .A(A[0]), .B(B[12]), .Z(n47177) );
  XNOR U47530 ( .A(n44965), .B(n47178), .Z(n44962) );
  NAND U47531 ( .A(A[0]), .B(B[13]), .Z(n47178) );
  NAND U47532 ( .A(B[12]), .B(A[1]), .Z(n44965) );
  XOR U47533 ( .A(n554), .B(n553), .Z(\A1[119] ) );
  XOR U47534 ( .A(n47097), .B(n47179), .Z(n553) );
  XNOR U47535 ( .A(n47096), .B(n47094), .Z(n47179) );
  AND U47536 ( .A(n47180), .B(n47181), .Z(n47094) );
  NANDN U47537 ( .A(n47182), .B(n47183), .Z(n47181) );
  NANDN U47538 ( .A(n47184), .B(n47185), .Z(n47183) );
  NANDN U47539 ( .A(n47185), .B(n47184), .Z(n47180) );
  ANDN U47540 ( .B(B[90]), .A(n54), .Z(n47096) );
  XNOR U47541 ( .A(n46891), .B(n47186), .Z(n47097) );
  XNOR U47542 ( .A(n46890), .B(n46888), .Z(n47186) );
  AND U47543 ( .A(n47187), .B(n47188), .Z(n46888) );
  NANDN U47544 ( .A(n47189), .B(n47190), .Z(n47188) );
  OR U47545 ( .A(n47191), .B(n47192), .Z(n47190) );
  NAND U47546 ( .A(n47192), .B(n47191), .Z(n47187) );
  ANDN U47547 ( .B(B[91]), .A(n55), .Z(n46890) );
  XNOR U47548 ( .A(n46898), .B(n47193), .Z(n46891) );
  XNOR U47549 ( .A(n46897), .B(n46895), .Z(n47193) );
  AND U47550 ( .A(n47194), .B(n47195), .Z(n46895) );
  NANDN U47551 ( .A(n47196), .B(n47197), .Z(n47195) );
  NANDN U47552 ( .A(n47198), .B(n47199), .Z(n47197) );
  NANDN U47553 ( .A(n47199), .B(n47198), .Z(n47194) );
  ANDN U47554 ( .B(B[92]), .A(n56), .Z(n46897) );
  XNOR U47555 ( .A(n46905), .B(n47200), .Z(n46898) );
  XNOR U47556 ( .A(n46904), .B(n46902), .Z(n47200) );
  AND U47557 ( .A(n47201), .B(n47202), .Z(n46902) );
  NANDN U47558 ( .A(n47203), .B(n47204), .Z(n47202) );
  OR U47559 ( .A(n47205), .B(n47206), .Z(n47204) );
  NAND U47560 ( .A(n47206), .B(n47205), .Z(n47201) );
  ANDN U47561 ( .B(B[93]), .A(n57), .Z(n46904) );
  XNOR U47562 ( .A(n46912), .B(n47207), .Z(n46905) );
  XNOR U47563 ( .A(n46911), .B(n46909), .Z(n47207) );
  AND U47564 ( .A(n47208), .B(n47209), .Z(n46909) );
  NANDN U47565 ( .A(n47210), .B(n47211), .Z(n47209) );
  NANDN U47566 ( .A(n47212), .B(n47213), .Z(n47211) );
  NANDN U47567 ( .A(n47213), .B(n47212), .Z(n47208) );
  ANDN U47568 ( .B(B[94]), .A(n58), .Z(n46911) );
  XNOR U47569 ( .A(n46919), .B(n47214), .Z(n46912) );
  XNOR U47570 ( .A(n46918), .B(n46916), .Z(n47214) );
  AND U47571 ( .A(n47215), .B(n47216), .Z(n46916) );
  NANDN U47572 ( .A(n47217), .B(n47218), .Z(n47216) );
  OR U47573 ( .A(n47219), .B(n47220), .Z(n47218) );
  NAND U47574 ( .A(n47220), .B(n47219), .Z(n47215) );
  ANDN U47575 ( .B(A[26]), .A(n13), .Z(n46918) );
  XNOR U47576 ( .A(n46926), .B(n47221), .Z(n46919) );
  XNOR U47577 ( .A(n46925), .B(n46923), .Z(n47221) );
  AND U47578 ( .A(n47222), .B(n47223), .Z(n46923) );
  NANDN U47579 ( .A(n47224), .B(n47225), .Z(n47223) );
  NANDN U47580 ( .A(n47226), .B(n47227), .Z(n47225) );
  NANDN U47581 ( .A(n47227), .B(n47226), .Z(n47222) );
  ANDN U47582 ( .B(A[25]), .A(n11), .Z(n46925) );
  XNOR U47583 ( .A(n46933), .B(n47228), .Z(n46926) );
  XNOR U47584 ( .A(n46932), .B(n46930), .Z(n47228) );
  AND U47585 ( .A(n47229), .B(n47230), .Z(n46930) );
  NANDN U47586 ( .A(n47231), .B(n47232), .Z(n47230) );
  OR U47587 ( .A(n47233), .B(n47234), .Z(n47232) );
  NAND U47588 ( .A(n47234), .B(n47233), .Z(n47229) );
  ANDN U47589 ( .B(A[24]), .A(n9), .Z(n46932) );
  XNOR U47590 ( .A(n46940), .B(n47235), .Z(n46933) );
  XNOR U47591 ( .A(n46939), .B(n46937), .Z(n47235) );
  AND U47592 ( .A(n47236), .B(n47237), .Z(n46937) );
  NANDN U47593 ( .A(n47238), .B(n47239), .Z(n47237) );
  NANDN U47594 ( .A(n47240), .B(n47241), .Z(n47239) );
  NANDN U47595 ( .A(n47241), .B(n47240), .Z(n47236) );
  ANDN U47596 ( .B(B[98]), .A(n62), .Z(n46939) );
  XNOR U47597 ( .A(n46947), .B(n47242), .Z(n46940) );
  XNOR U47598 ( .A(n46946), .B(n46944), .Z(n47242) );
  AND U47599 ( .A(n47243), .B(n47244), .Z(n46944) );
  NANDN U47600 ( .A(n47245), .B(n47246), .Z(n47244) );
  OR U47601 ( .A(n47247), .B(n47248), .Z(n47246) );
  NAND U47602 ( .A(n47248), .B(n47247), .Z(n47243) );
  ANDN U47603 ( .B(A[22]), .A(n6), .Z(n46946) );
  XNOR U47604 ( .A(n46954), .B(n47249), .Z(n46947) );
  XNOR U47605 ( .A(n46953), .B(n46951), .Z(n47249) );
  AND U47606 ( .A(n47250), .B(n47251), .Z(n46951) );
  NANDN U47607 ( .A(n47252), .B(n47253), .Z(n47251) );
  NANDN U47608 ( .A(n47254), .B(n47255), .Z(n47253) );
  NANDN U47609 ( .A(n47255), .B(n47254), .Z(n47250) );
  ANDN U47610 ( .B(A[21]), .A(n4), .Z(n46953) );
  XNOR U47611 ( .A(n46961), .B(n47256), .Z(n46954) );
  XNOR U47612 ( .A(n46960), .B(n46958), .Z(n47256) );
  AND U47613 ( .A(n47257), .B(n47258), .Z(n46958) );
  NANDN U47614 ( .A(n47259), .B(n47260), .Z(n47258) );
  OR U47615 ( .A(n47261), .B(n47262), .Z(n47260) );
  NAND U47616 ( .A(n47262), .B(n47261), .Z(n47257) );
  ANDN U47617 ( .B(B[101]), .A(n65), .Z(n46960) );
  XNOR U47618 ( .A(n46968), .B(n47263), .Z(n46961) );
  XNOR U47619 ( .A(n46967), .B(n46965), .Z(n47263) );
  AND U47620 ( .A(n47264), .B(n47265), .Z(n46965) );
  NANDN U47621 ( .A(n47266), .B(n47267), .Z(n47265) );
  NANDN U47622 ( .A(n47268), .B(n47269), .Z(n47267) );
  NANDN U47623 ( .A(n47269), .B(n47268), .Z(n47264) );
  ANDN U47624 ( .B(B[102]), .A(n66), .Z(n46967) );
  XNOR U47625 ( .A(n46975), .B(n47270), .Z(n46968) );
  XNOR U47626 ( .A(n46974), .B(n46972), .Z(n47270) );
  AND U47627 ( .A(n47271), .B(n47272), .Z(n46972) );
  NANDN U47628 ( .A(n47273), .B(n47274), .Z(n47272) );
  OR U47629 ( .A(n47275), .B(n47276), .Z(n47274) );
  NAND U47630 ( .A(n47276), .B(n47275), .Z(n47271) );
  ANDN U47631 ( .B(B[103]), .A(n67), .Z(n46974) );
  XNOR U47632 ( .A(n46982), .B(n47277), .Z(n46975) );
  XNOR U47633 ( .A(n46981), .B(n46979), .Z(n47277) );
  AND U47634 ( .A(n47278), .B(n47279), .Z(n46979) );
  NANDN U47635 ( .A(n47280), .B(n47281), .Z(n47279) );
  NANDN U47636 ( .A(n47282), .B(n47283), .Z(n47281) );
  NANDN U47637 ( .A(n47283), .B(n47282), .Z(n47278) );
  ANDN U47638 ( .B(B[104]), .A(n68), .Z(n46981) );
  XNOR U47639 ( .A(n46989), .B(n47284), .Z(n46982) );
  XNOR U47640 ( .A(n46988), .B(n46986), .Z(n47284) );
  AND U47641 ( .A(n47285), .B(n47286), .Z(n46986) );
  NANDN U47642 ( .A(n47287), .B(n47288), .Z(n47286) );
  OR U47643 ( .A(n47289), .B(n47290), .Z(n47288) );
  NAND U47644 ( .A(n47290), .B(n47289), .Z(n47285) );
  ANDN U47645 ( .B(B[105]), .A(n69), .Z(n46988) );
  XNOR U47646 ( .A(n46996), .B(n47291), .Z(n46989) );
  XNOR U47647 ( .A(n46995), .B(n46993), .Z(n47291) );
  AND U47648 ( .A(n47292), .B(n47293), .Z(n46993) );
  NANDN U47649 ( .A(n47294), .B(n47295), .Z(n47293) );
  NANDN U47650 ( .A(n47296), .B(n47297), .Z(n47295) );
  NANDN U47651 ( .A(n47297), .B(n47296), .Z(n47292) );
  ANDN U47652 ( .B(B[106]), .A(n70), .Z(n46995) );
  XNOR U47653 ( .A(n47003), .B(n47298), .Z(n46996) );
  XNOR U47654 ( .A(n47002), .B(n47000), .Z(n47298) );
  AND U47655 ( .A(n47299), .B(n47300), .Z(n47000) );
  NANDN U47656 ( .A(n47301), .B(n47302), .Z(n47300) );
  OR U47657 ( .A(n47303), .B(n47304), .Z(n47302) );
  NAND U47658 ( .A(n47304), .B(n47303), .Z(n47299) );
  ANDN U47659 ( .B(B[107]), .A(n71), .Z(n47002) );
  XNOR U47660 ( .A(n47010), .B(n47305), .Z(n47003) );
  XNOR U47661 ( .A(n47009), .B(n47007), .Z(n47305) );
  AND U47662 ( .A(n47306), .B(n47307), .Z(n47007) );
  NANDN U47663 ( .A(n47308), .B(n47309), .Z(n47307) );
  NANDN U47664 ( .A(n47310), .B(n47311), .Z(n47309) );
  NANDN U47665 ( .A(n47311), .B(n47310), .Z(n47306) );
  ANDN U47666 ( .B(B[108]), .A(n72), .Z(n47009) );
  XNOR U47667 ( .A(n47017), .B(n47312), .Z(n47010) );
  XNOR U47668 ( .A(n47016), .B(n47014), .Z(n47312) );
  AND U47669 ( .A(n47313), .B(n47314), .Z(n47014) );
  NANDN U47670 ( .A(n47315), .B(n47316), .Z(n47314) );
  OR U47671 ( .A(n47317), .B(n47318), .Z(n47316) );
  NAND U47672 ( .A(n47318), .B(n47317), .Z(n47313) );
  ANDN U47673 ( .B(B[109]), .A(n73), .Z(n47016) );
  XNOR U47674 ( .A(n47024), .B(n47319), .Z(n47017) );
  XNOR U47675 ( .A(n47023), .B(n47021), .Z(n47319) );
  AND U47676 ( .A(n47320), .B(n47321), .Z(n47021) );
  NANDN U47677 ( .A(n47322), .B(n47323), .Z(n47321) );
  NANDN U47678 ( .A(n47324), .B(n47325), .Z(n47323) );
  NANDN U47679 ( .A(n47325), .B(n47324), .Z(n47320) );
  ANDN U47680 ( .B(B[110]), .A(n74), .Z(n47023) );
  XNOR U47681 ( .A(n47031), .B(n47326), .Z(n47024) );
  XNOR U47682 ( .A(n47030), .B(n47028), .Z(n47326) );
  AND U47683 ( .A(n47327), .B(n47328), .Z(n47028) );
  NANDN U47684 ( .A(n47329), .B(n47330), .Z(n47328) );
  OR U47685 ( .A(n47331), .B(n47332), .Z(n47330) );
  NAND U47686 ( .A(n47332), .B(n47331), .Z(n47327) );
  ANDN U47687 ( .B(B[111]), .A(n75), .Z(n47030) );
  XNOR U47688 ( .A(n47038), .B(n47333), .Z(n47031) );
  XNOR U47689 ( .A(n47037), .B(n47035), .Z(n47333) );
  AND U47690 ( .A(n47334), .B(n47335), .Z(n47035) );
  NANDN U47691 ( .A(n47336), .B(n47337), .Z(n47335) );
  NANDN U47692 ( .A(n47338), .B(n47339), .Z(n47337) );
  NANDN U47693 ( .A(n47339), .B(n47338), .Z(n47334) );
  ANDN U47694 ( .B(B[112]), .A(n76), .Z(n47037) );
  XNOR U47695 ( .A(n47045), .B(n47340), .Z(n47038) );
  XNOR U47696 ( .A(n47044), .B(n47042), .Z(n47340) );
  AND U47697 ( .A(n47341), .B(n47342), .Z(n47042) );
  NANDN U47698 ( .A(n47343), .B(n47344), .Z(n47342) );
  OR U47699 ( .A(n47345), .B(n47346), .Z(n47344) );
  NAND U47700 ( .A(n47346), .B(n47345), .Z(n47341) );
  ANDN U47701 ( .B(B[113]), .A(n77), .Z(n47044) );
  XNOR U47702 ( .A(n47052), .B(n47347), .Z(n47045) );
  XNOR U47703 ( .A(n47051), .B(n47049), .Z(n47347) );
  AND U47704 ( .A(n47348), .B(n47349), .Z(n47049) );
  NANDN U47705 ( .A(n47350), .B(n47351), .Z(n47349) );
  NANDN U47706 ( .A(n47352), .B(n47353), .Z(n47351) );
  NANDN U47707 ( .A(n47353), .B(n47352), .Z(n47348) );
  ANDN U47708 ( .B(B[114]), .A(n78), .Z(n47051) );
  XNOR U47709 ( .A(n47059), .B(n47354), .Z(n47052) );
  XNOR U47710 ( .A(n47058), .B(n47056), .Z(n47354) );
  AND U47711 ( .A(n47355), .B(n47356), .Z(n47056) );
  NANDN U47712 ( .A(n47357), .B(n47358), .Z(n47356) );
  OR U47713 ( .A(n47359), .B(n47360), .Z(n47358) );
  NAND U47714 ( .A(n47360), .B(n47359), .Z(n47355) );
  ANDN U47715 ( .B(B[115]), .A(n79), .Z(n47058) );
  XNOR U47716 ( .A(n47066), .B(n47361), .Z(n47059) );
  XNOR U47717 ( .A(n47065), .B(n47063), .Z(n47361) );
  AND U47718 ( .A(n47362), .B(n47363), .Z(n47063) );
  NANDN U47719 ( .A(n47364), .B(n47365), .Z(n47363) );
  NANDN U47720 ( .A(n47366), .B(n47367), .Z(n47365) );
  NANDN U47721 ( .A(n47367), .B(n47366), .Z(n47362) );
  ANDN U47722 ( .B(B[116]), .A(n80), .Z(n47065) );
  XNOR U47723 ( .A(n47073), .B(n47368), .Z(n47066) );
  XNOR U47724 ( .A(n47072), .B(n47070), .Z(n47368) );
  AND U47725 ( .A(n47369), .B(n47370), .Z(n47070) );
  NANDN U47726 ( .A(n47371), .B(n47372), .Z(n47370) );
  OR U47727 ( .A(n47373), .B(n47374), .Z(n47372) );
  NAND U47728 ( .A(n47374), .B(n47373), .Z(n47369) );
  ANDN U47729 ( .B(B[117]), .A(n81), .Z(n47072) );
  XNOR U47730 ( .A(n47080), .B(n47375), .Z(n47073) );
  XNOR U47731 ( .A(n47079), .B(n47077), .Z(n47375) );
  AND U47732 ( .A(n47376), .B(n47377), .Z(n47077) );
  NANDN U47733 ( .A(n47378), .B(n47379), .Z(n47377) );
  NAND U47734 ( .A(n47380), .B(n47381), .Z(n47379) );
  ANDN U47735 ( .B(B[118]), .A(n82), .Z(n47079) );
  XOR U47736 ( .A(n47086), .B(n47382), .Z(n47080) );
  XNOR U47737 ( .A(n47084), .B(n47087), .Z(n47382) );
  NAND U47738 ( .A(A[2]), .B(B[119]), .Z(n47087) );
  NANDN U47739 ( .A(n47383), .B(n47384), .Z(n47084) );
  AND U47740 ( .A(A[0]), .B(B[120]), .Z(n47384) );
  XNOR U47741 ( .A(n47089), .B(n47385), .Z(n47086) );
  NAND U47742 ( .A(A[0]), .B(B[121]), .Z(n47385) );
  NAND U47743 ( .A(B[120]), .B(A[1]), .Z(n47089) );
  NAND U47744 ( .A(n47386), .B(n47387), .Z(n554) );
  NANDN U47745 ( .A(n47388), .B(n47389), .Z(n47387) );
  OR U47746 ( .A(n47390), .B(n47391), .Z(n47389) );
  NAND U47747 ( .A(n47391), .B(n47390), .Z(n47386) );
  XOR U47748 ( .A(n556), .B(n555), .Z(\A1[118] ) );
  XOR U47749 ( .A(n47391), .B(n47392), .Z(n555) );
  XNOR U47750 ( .A(n47390), .B(n47388), .Z(n47392) );
  AND U47751 ( .A(n47393), .B(n47394), .Z(n47388) );
  NANDN U47752 ( .A(n47395), .B(n47396), .Z(n47394) );
  NANDN U47753 ( .A(n47397), .B(n47398), .Z(n47396) );
  NANDN U47754 ( .A(n47398), .B(n47397), .Z(n47393) );
  ANDN U47755 ( .B(B[89]), .A(n54), .Z(n47390) );
  XNOR U47756 ( .A(n47185), .B(n47399), .Z(n47391) );
  XNOR U47757 ( .A(n47184), .B(n47182), .Z(n47399) );
  AND U47758 ( .A(n47400), .B(n47401), .Z(n47182) );
  NANDN U47759 ( .A(n47402), .B(n47403), .Z(n47401) );
  OR U47760 ( .A(n47404), .B(n47405), .Z(n47403) );
  NAND U47761 ( .A(n47405), .B(n47404), .Z(n47400) );
  ANDN U47762 ( .B(B[90]), .A(n55), .Z(n47184) );
  XNOR U47763 ( .A(n47192), .B(n47406), .Z(n47185) );
  XNOR U47764 ( .A(n47191), .B(n47189), .Z(n47406) );
  AND U47765 ( .A(n47407), .B(n47408), .Z(n47189) );
  NANDN U47766 ( .A(n47409), .B(n47410), .Z(n47408) );
  NANDN U47767 ( .A(n47411), .B(n47412), .Z(n47410) );
  NANDN U47768 ( .A(n47412), .B(n47411), .Z(n47407) );
  ANDN U47769 ( .B(B[91]), .A(n56), .Z(n47191) );
  XNOR U47770 ( .A(n47199), .B(n47413), .Z(n47192) );
  XNOR U47771 ( .A(n47198), .B(n47196), .Z(n47413) );
  AND U47772 ( .A(n47414), .B(n47415), .Z(n47196) );
  NANDN U47773 ( .A(n47416), .B(n47417), .Z(n47415) );
  OR U47774 ( .A(n47418), .B(n47419), .Z(n47417) );
  NAND U47775 ( .A(n47419), .B(n47418), .Z(n47414) );
  ANDN U47776 ( .B(B[92]), .A(n57), .Z(n47198) );
  XNOR U47777 ( .A(n47206), .B(n47420), .Z(n47199) );
  XNOR U47778 ( .A(n47205), .B(n47203), .Z(n47420) );
  AND U47779 ( .A(n47421), .B(n47422), .Z(n47203) );
  NANDN U47780 ( .A(n47423), .B(n47424), .Z(n47422) );
  NANDN U47781 ( .A(n47425), .B(n47426), .Z(n47424) );
  NANDN U47782 ( .A(n47426), .B(n47425), .Z(n47421) );
  ANDN U47783 ( .B(B[93]), .A(n58), .Z(n47205) );
  XNOR U47784 ( .A(n47213), .B(n47427), .Z(n47206) );
  XNOR U47785 ( .A(n47212), .B(n47210), .Z(n47427) );
  AND U47786 ( .A(n47428), .B(n47429), .Z(n47210) );
  NANDN U47787 ( .A(n47430), .B(n47431), .Z(n47429) );
  OR U47788 ( .A(n47432), .B(n47433), .Z(n47431) );
  NAND U47789 ( .A(n47433), .B(n47432), .Z(n47428) );
  ANDN U47790 ( .B(A[26]), .A(n15), .Z(n47212) );
  XNOR U47791 ( .A(n47220), .B(n47434), .Z(n47213) );
  XNOR U47792 ( .A(n47219), .B(n47217), .Z(n47434) );
  AND U47793 ( .A(n47435), .B(n47436), .Z(n47217) );
  NANDN U47794 ( .A(n47437), .B(n47438), .Z(n47436) );
  NANDN U47795 ( .A(n47439), .B(n47440), .Z(n47438) );
  NANDN U47796 ( .A(n47440), .B(n47439), .Z(n47435) );
  ANDN U47797 ( .B(A[25]), .A(n13), .Z(n47219) );
  XNOR U47798 ( .A(n47227), .B(n47441), .Z(n47220) );
  XNOR U47799 ( .A(n47226), .B(n47224), .Z(n47441) );
  AND U47800 ( .A(n47442), .B(n47443), .Z(n47224) );
  NANDN U47801 ( .A(n47444), .B(n47445), .Z(n47443) );
  OR U47802 ( .A(n47446), .B(n47447), .Z(n47445) );
  NAND U47803 ( .A(n47447), .B(n47446), .Z(n47442) );
  ANDN U47804 ( .B(A[24]), .A(n11), .Z(n47226) );
  XNOR U47805 ( .A(n47234), .B(n47448), .Z(n47227) );
  XNOR U47806 ( .A(n47233), .B(n47231), .Z(n47448) );
  AND U47807 ( .A(n47449), .B(n47450), .Z(n47231) );
  NANDN U47808 ( .A(n47451), .B(n47452), .Z(n47450) );
  NANDN U47809 ( .A(n47453), .B(n47454), .Z(n47452) );
  NANDN U47810 ( .A(n47454), .B(n47453), .Z(n47449) );
  ANDN U47811 ( .B(A[23]), .A(n9), .Z(n47233) );
  XNOR U47812 ( .A(n47241), .B(n47455), .Z(n47234) );
  XNOR U47813 ( .A(n47240), .B(n47238), .Z(n47455) );
  AND U47814 ( .A(n47456), .B(n47457), .Z(n47238) );
  NANDN U47815 ( .A(n47458), .B(n47459), .Z(n47457) );
  OR U47816 ( .A(n47460), .B(n47461), .Z(n47459) );
  NAND U47817 ( .A(n47461), .B(n47460), .Z(n47456) );
  ANDN U47818 ( .B(B[98]), .A(n63), .Z(n47240) );
  XNOR U47819 ( .A(n47248), .B(n47462), .Z(n47241) );
  XNOR U47820 ( .A(n47247), .B(n47245), .Z(n47462) );
  AND U47821 ( .A(n47463), .B(n47464), .Z(n47245) );
  NANDN U47822 ( .A(n47465), .B(n47466), .Z(n47464) );
  NANDN U47823 ( .A(n47467), .B(n47468), .Z(n47466) );
  NANDN U47824 ( .A(n47468), .B(n47467), .Z(n47463) );
  ANDN U47825 ( .B(A[21]), .A(n6), .Z(n47247) );
  XNOR U47826 ( .A(n47255), .B(n47469), .Z(n47248) );
  XNOR U47827 ( .A(n47254), .B(n47252), .Z(n47469) );
  AND U47828 ( .A(n47470), .B(n47471), .Z(n47252) );
  NANDN U47829 ( .A(n47472), .B(n47473), .Z(n47471) );
  OR U47830 ( .A(n47474), .B(n47475), .Z(n47473) );
  NAND U47831 ( .A(n47475), .B(n47474), .Z(n47470) );
  ANDN U47832 ( .B(A[20]), .A(n4), .Z(n47254) );
  XNOR U47833 ( .A(n47262), .B(n47476), .Z(n47255) );
  XNOR U47834 ( .A(n47261), .B(n47259), .Z(n47476) );
  AND U47835 ( .A(n47477), .B(n47478), .Z(n47259) );
  NANDN U47836 ( .A(n47479), .B(n47480), .Z(n47478) );
  NANDN U47837 ( .A(n47481), .B(n47482), .Z(n47480) );
  NANDN U47838 ( .A(n47482), .B(n47481), .Z(n47477) );
  ANDN U47839 ( .B(B[101]), .A(n66), .Z(n47261) );
  XNOR U47840 ( .A(n47269), .B(n47483), .Z(n47262) );
  XNOR U47841 ( .A(n47268), .B(n47266), .Z(n47483) );
  AND U47842 ( .A(n47484), .B(n47485), .Z(n47266) );
  NANDN U47843 ( .A(n47486), .B(n47487), .Z(n47485) );
  OR U47844 ( .A(n47488), .B(n47489), .Z(n47487) );
  NAND U47845 ( .A(n47489), .B(n47488), .Z(n47484) );
  ANDN U47846 ( .B(B[102]), .A(n67), .Z(n47268) );
  XNOR U47847 ( .A(n47276), .B(n47490), .Z(n47269) );
  XNOR U47848 ( .A(n47275), .B(n47273), .Z(n47490) );
  AND U47849 ( .A(n47491), .B(n47492), .Z(n47273) );
  NANDN U47850 ( .A(n47493), .B(n47494), .Z(n47492) );
  NANDN U47851 ( .A(n47495), .B(n47496), .Z(n47494) );
  NANDN U47852 ( .A(n47496), .B(n47495), .Z(n47491) );
  ANDN U47853 ( .B(B[103]), .A(n68), .Z(n47275) );
  XNOR U47854 ( .A(n47283), .B(n47497), .Z(n47276) );
  XNOR U47855 ( .A(n47282), .B(n47280), .Z(n47497) );
  AND U47856 ( .A(n47498), .B(n47499), .Z(n47280) );
  NANDN U47857 ( .A(n47500), .B(n47501), .Z(n47499) );
  OR U47858 ( .A(n47502), .B(n47503), .Z(n47501) );
  NAND U47859 ( .A(n47503), .B(n47502), .Z(n47498) );
  ANDN U47860 ( .B(B[104]), .A(n69), .Z(n47282) );
  XNOR U47861 ( .A(n47290), .B(n47504), .Z(n47283) );
  XNOR U47862 ( .A(n47289), .B(n47287), .Z(n47504) );
  AND U47863 ( .A(n47505), .B(n47506), .Z(n47287) );
  NANDN U47864 ( .A(n47507), .B(n47508), .Z(n47506) );
  NANDN U47865 ( .A(n47509), .B(n47510), .Z(n47508) );
  NANDN U47866 ( .A(n47510), .B(n47509), .Z(n47505) );
  ANDN U47867 ( .B(B[105]), .A(n70), .Z(n47289) );
  XNOR U47868 ( .A(n47297), .B(n47511), .Z(n47290) );
  XNOR U47869 ( .A(n47296), .B(n47294), .Z(n47511) );
  AND U47870 ( .A(n47512), .B(n47513), .Z(n47294) );
  NANDN U47871 ( .A(n47514), .B(n47515), .Z(n47513) );
  OR U47872 ( .A(n47516), .B(n47517), .Z(n47515) );
  NAND U47873 ( .A(n47517), .B(n47516), .Z(n47512) );
  ANDN U47874 ( .B(B[106]), .A(n71), .Z(n47296) );
  XNOR U47875 ( .A(n47304), .B(n47518), .Z(n47297) );
  XNOR U47876 ( .A(n47303), .B(n47301), .Z(n47518) );
  AND U47877 ( .A(n47519), .B(n47520), .Z(n47301) );
  NANDN U47878 ( .A(n47521), .B(n47522), .Z(n47520) );
  NANDN U47879 ( .A(n47523), .B(n47524), .Z(n47522) );
  NANDN U47880 ( .A(n47524), .B(n47523), .Z(n47519) );
  ANDN U47881 ( .B(B[107]), .A(n72), .Z(n47303) );
  XNOR U47882 ( .A(n47311), .B(n47525), .Z(n47304) );
  XNOR U47883 ( .A(n47310), .B(n47308), .Z(n47525) );
  AND U47884 ( .A(n47526), .B(n47527), .Z(n47308) );
  NANDN U47885 ( .A(n47528), .B(n47529), .Z(n47527) );
  OR U47886 ( .A(n47530), .B(n47531), .Z(n47529) );
  NAND U47887 ( .A(n47531), .B(n47530), .Z(n47526) );
  ANDN U47888 ( .B(B[108]), .A(n73), .Z(n47310) );
  XNOR U47889 ( .A(n47318), .B(n47532), .Z(n47311) );
  XNOR U47890 ( .A(n47317), .B(n47315), .Z(n47532) );
  AND U47891 ( .A(n47533), .B(n47534), .Z(n47315) );
  NANDN U47892 ( .A(n47535), .B(n47536), .Z(n47534) );
  NANDN U47893 ( .A(n47537), .B(n47538), .Z(n47536) );
  NANDN U47894 ( .A(n47538), .B(n47537), .Z(n47533) );
  ANDN U47895 ( .B(B[109]), .A(n74), .Z(n47317) );
  XNOR U47896 ( .A(n47325), .B(n47539), .Z(n47318) );
  XNOR U47897 ( .A(n47324), .B(n47322), .Z(n47539) );
  AND U47898 ( .A(n47540), .B(n47541), .Z(n47322) );
  NANDN U47899 ( .A(n47542), .B(n47543), .Z(n47541) );
  OR U47900 ( .A(n47544), .B(n47545), .Z(n47543) );
  NAND U47901 ( .A(n47545), .B(n47544), .Z(n47540) );
  ANDN U47902 ( .B(B[110]), .A(n75), .Z(n47324) );
  XNOR U47903 ( .A(n47332), .B(n47546), .Z(n47325) );
  XNOR U47904 ( .A(n47331), .B(n47329), .Z(n47546) );
  AND U47905 ( .A(n47547), .B(n47548), .Z(n47329) );
  NANDN U47906 ( .A(n47549), .B(n47550), .Z(n47548) );
  NANDN U47907 ( .A(n47551), .B(n47552), .Z(n47550) );
  NANDN U47908 ( .A(n47552), .B(n47551), .Z(n47547) );
  ANDN U47909 ( .B(B[111]), .A(n76), .Z(n47331) );
  XNOR U47910 ( .A(n47339), .B(n47553), .Z(n47332) );
  XNOR U47911 ( .A(n47338), .B(n47336), .Z(n47553) );
  AND U47912 ( .A(n47554), .B(n47555), .Z(n47336) );
  NANDN U47913 ( .A(n47556), .B(n47557), .Z(n47555) );
  OR U47914 ( .A(n47558), .B(n47559), .Z(n47557) );
  NAND U47915 ( .A(n47559), .B(n47558), .Z(n47554) );
  ANDN U47916 ( .B(B[112]), .A(n77), .Z(n47338) );
  XNOR U47917 ( .A(n47346), .B(n47560), .Z(n47339) );
  XNOR U47918 ( .A(n47345), .B(n47343), .Z(n47560) );
  AND U47919 ( .A(n47561), .B(n47562), .Z(n47343) );
  NANDN U47920 ( .A(n47563), .B(n47564), .Z(n47562) );
  NANDN U47921 ( .A(n47565), .B(n47566), .Z(n47564) );
  NANDN U47922 ( .A(n47566), .B(n47565), .Z(n47561) );
  ANDN U47923 ( .B(B[113]), .A(n78), .Z(n47345) );
  XNOR U47924 ( .A(n47353), .B(n47567), .Z(n47346) );
  XNOR U47925 ( .A(n47352), .B(n47350), .Z(n47567) );
  AND U47926 ( .A(n47568), .B(n47569), .Z(n47350) );
  NANDN U47927 ( .A(n47570), .B(n47571), .Z(n47569) );
  OR U47928 ( .A(n47572), .B(n47573), .Z(n47571) );
  NAND U47929 ( .A(n47573), .B(n47572), .Z(n47568) );
  ANDN U47930 ( .B(B[114]), .A(n79), .Z(n47352) );
  XNOR U47931 ( .A(n47360), .B(n47574), .Z(n47353) );
  XNOR U47932 ( .A(n47359), .B(n47357), .Z(n47574) );
  AND U47933 ( .A(n47575), .B(n47576), .Z(n47357) );
  NANDN U47934 ( .A(n47577), .B(n47578), .Z(n47576) );
  NANDN U47935 ( .A(n47579), .B(n47580), .Z(n47578) );
  NANDN U47936 ( .A(n47580), .B(n47579), .Z(n47575) );
  ANDN U47937 ( .B(B[115]), .A(n80), .Z(n47359) );
  XNOR U47938 ( .A(n47367), .B(n47581), .Z(n47360) );
  XNOR U47939 ( .A(n47366), .B(n47364), .Z(n47581) );
  AND U47940 ( .A(n47582), .B(n47583), .Z(n47364) );
  NANDN U47941 ( .A(n47584), .B(n47585), .Z(n47583) );
  OR U47942 ( .A(n47586), .B(n47587), .Z(n47585) );
  NAND U47943 ( .A(n47587), .B(n47586), .Z(n47582) );
  ANDN U47944 ( .B(B[116]), .A(n81), .Z(n47366) );
  XNOR U47945 ( .A(n47374), .B(n47588), .Z(n47367) );
  XNOR U47946 ( .A(n47373), .B(n47371), .Z(n47588) );
  AND U47947 ( .A(n47589), .B(n47590), .Z(n47371) );
  NANDN U47948 ( .A(n47591), .B(n47592), .Z(n47590) );
  NAND U47949 ( .A(n47593), .B(n47594), .Z(n47592) );
  ANDN U47950 ( .B(B[117]), .A(n82), .Z(n47373) );
  XOR U47951 ( .A(n47380), .B(n47595), .Z(n47374) );
  XNOR U47952 ( .A(n47378), .B(n47381), .Z(n47595) );
  NAND U47953 ( .A(A[2]), .B(B[118]), .Z(n47381) );
  NANDN U47954 ( .A(n47596), .B(n47597), .Z(n47378) );
  AND U47955 ( .A(A[0]), .B(B[119]), .Z(n47597) );
  XNOR U47956 ( .A(n47383), .B(n47598), .Z(n47380) );
  NAND U47957 ( .A(A[0]), .B(B[120]), .Z(n47598) );
  NAND U47958 ( .A(B[119]), .B(A[1]), .Z(n47383) );
  NAND U47959 ( .A(n47599), .B(n47600), .Z(n556) );
  NANDN U47960 ( .A(n47601), .B(n47602), .Z(n47600) );
  OR U47961 ( .A(n47603), .B(n47604), .Z(n47602) );
  NAND U47962 ( .A(n47604), .B(n47603), .Z(n47599) );
  XOR U47963 ( .A(n558), .B(n557), .Z(\A1[117] ) );
  XOR U47964 ( .A(n47604), .B(n47605), .Z(n557) );
  XNOR U47965 ( .A(n47603), .B(n47601), .Z(n47605) );
  AND U47966 ( .A(n47606), .B(n47607), .Z(n47601) );
  NANDN U47967 ( .A(n47608), .B(n47609), .Z(n47607) );
  NANDN U47968 ( .A(n47610), .B(n47611), .Z(n47609) );
  NANDN U47969 ( .A(n47611), .B(n47610), .Z(n47606) );
  ANDN U47970 ( .B(B[88]), .A(n54), .Z(n47603) );
  XNOR U47971 ( .A(n47398), .B(n47612), .Z(n47604) );
  XNOR U47972 ( .A(n47397), .B(n47395), .Z(n47612) );
  AND U47973 ( .A(n47613), .B(n47614), .Z(n47395) );
  NANDN U47974 ( .A(n47615), .B(n47616), .Z(n47614) );
  OR U47975 ( .A(n47617), .B(n47618), .Z(n47616) );
  NAND U47976 ( .A(n47618), .B(n47617), .Z(n47613) );
  ANDN U47977 ( .B(B[89]), .A(n55), .Z(n47397) );
  XNOR U47978 ( .A(n47405), .B(n47619), .Z(n47398) );
  XNOR U47979 ( .A(n47404), .B(n47402), .Z(n47619) );
  AND U47980 ( .A(n47620), .B(n47621), .Z(n47402) );
  NANDN U47981 ( .A(n47622), .B(n47623), .Z(n47621) );
  NANDN U47982 ( .A(n47624), .B(n47625), .Z(n47623) );
  NANDN U47983 ( .A(n47625), .B(n47624), .Z(n47620) );
  ANDN U47984 ( .B(B[90]), .A(n56), .Z(n47404) );
  XNOR U47985 ( .A(n47412), .B(n47626), .Z(n47405) );
  XNOR U47986 ( .A(n47411), .B(n47409), .Z(n47626) );
  AND U47987 ( .A(n47627), .B(n47628), .Z(n47409) );
  NANDN U47988 ( .A(n47629), .B(n47630), .Z(n47628) );
  OR U47989 ( .A(n47631), .B(n47632), .Z(n47630) );
  NAND U47990 ( .A(n47632), .B(n47631), .Z(n47627) );
  ANDN U47991 ( .B(B[91]), .A(n57), .Z(n47411) );
  XNOR U47992 ( .A(n47419), .B(n47633), .Z(n47412) );
  XNOR U47993 ( .A(n47418), .B(n47416), .Z(n47633) );
  AND U47994 ( .A(n47634), .B(n47635), .Z(n47416) );
  NANDN U47995 ( .A(n47636), .B(n47637), .Z(n47635) );
  NANDN U47996 ( .A(n47638), .B(n47639), .Z(n47637) );
  NANDN U47997 ( .A(n47639), .B(n47638), .Z(n47634) );
  ANDN U47998 ( .B(B[92]), .A(n58), .Z(n47418) );
  XNOR U47999 ( .A(n47426), .B(n47640), .Z(n47419) );
  XNOR U48000 ( .A(n47425), .B(n47423), .Z(n47640) );
  AND U48001 ( .A(n47641), .B(n47642), .Z(n47423) );
  NANDN U48002 ( .A(n47643), .B(n47644), .Z(n47642) );
  OR U48003 ( .A(n47645), .B(n47646), .Z(n47644) );
  NAND U48004 ( .A(n47646), .B(n47645), .Z(n47641) );
  ANDN U48005 ( .B(B[93]), .A(n59), .Z(n47425) );
  XNOR U48006 ( .A(n47433), .B(n47647), .Z(n47426) );
  XNOR U48007 ( .A(n47432), .B(n47430), .Z(n47647) );
  AND U48008 ( .A(n47648), .B(n47649), .Z(n47430) );
  NANDN U48009 ( .A(n47650), .B(n47651), .Z(n47649) );
  NANDN U48010 ( .A(n47652), .B(n47653), .Z(n47651) );
  NANDN U48011 ( .A(n47653), .B(n47652), .Z(n47648) );
  ANDN U48012 ( .B(A[25]), .A(n15), .Z(n47432) );
  XNOR U48013 ( .A(n47440), .B(n47654), .Z(n47433) );
  XNOR U48014 ( .A(n47439), .B(n47437), .Z(n47654) );
  AND U48015 ( .A(n47655), .B(n47656), .Z(n47437) );
  NANDN U48016 ( .A(n47657), .B(n47658), .Z(n47656) );
  OR U48017 ( .A(n47659), .B(n47660), .Z(n47658) );
  NAND U48018 ( .A(n47660), .B(n47659), .Z(n47655) );
  ANDN U48019 ( .B(A[24]), .A(n13), .Z(n47439) );
  XNOR U48020 ( .A(n47447), .B(n47661), .Z(n47440) );
  XNOR U48021 ( .A(n47446), .B(n47444), .Z(n47661) );
  AND U48022 ( .A(n47662), .B(n47663), .Z(n47444) );
  NANDN U48023 ( .A(n47664), .B(n47665), .Z(n47663) );
  NANDN U48024 ( .A(n47666), .B(n47667), .Z(n47665) );
  NANDN U48025 ( .A(n47667), .B(n47666), .Z(n47662) );
  ANDN U48026 ( .B(A[23]), .A(n11), .Z(n47446) );
  XNOR U48027 ( .A(n47454), .B(n47668), .Z(n47447) );
  XNOR U48028 ( .A(n47453), .B(n47451), .Z(n47668) );
  AND U48029 ( .A(n47669), .B(n47670), .Z(n47451) );
  NANDN U48030 ( .A(n47671), .B(n47672), .Z(n47670) );
  OR U48031 ( .A(n47673), .B(n47674), .Z(n47672) );
  NAND U48032 ( .A(n47674), .B(n47673), .Z(n47669) );
  ANDN U48033 ( .B(A[22]), .A(n9), .Z(n47453) );
  XNOR U48034 ( .A(n47461), .B(n47675), .Z(n47454) );
  XNOR U48035 ( .A(n47460), .B(n47458), .Z(n47675) );
  AND U48036 ( .A(n47676), .B(n47677), .Z(n47458) );
  NANDN U48037 ( .A(n47678), .B(n47679), .Z(n47677) );
  NANDN U48038 ( .A(n47680), .B(n47681), .Z(n47679) );
  NANDN U48039 ( .A(n47681), .B(n47680), .Z(n47676) );
  ANDN U48040 ( .B(B[98]), .A(n64), .Z(n47460) );
  XNOR U48041 ( .A(n47468), .B(n47682), .Z(n47461) );
  XNOR U48042 ( .A(n47467), .B(n47465), .Z(n47682) );
  AND U48043 ( .A(n47683), .B(n47684), .Z(n47465) );
  NANDN U48044 ( .A(n47685), .B(n47686), .Z(n47684) );
  OR U48045 ( .A(n47687), .B(n47688), .Z(n47686) );
  NAND U48046 ( .A(n47688), .B(n47687), .Z(n47683) );
  ANDN U48047 ( .B(A[20]), .A(n6), .Z(n47467) );
  XNOR U48048 ( .A(n47475), .B(n47689), .Z(n47468) );
  XNOR U48049 ( .A(n47474), .B(n47472), .Z(n47689) );
  AND U48050 ( .A(n47690), .B(n47691), .Z(n47472) );
  NANDN U48051 ( .A(n47692), .B(n47693), .Z(n47691) );
  NANDN U48052 ( .A(n47694), .B(n47695), .Z(n47693) );
  NANDN U48053 ( .A(n47695), .B(n47694), .Z(n47690) );
  ANDN U48054 ( .B(A[19]), .A(n4), .Z(n47474) );
  XNOR U48055 ( .A(n47482), .B(n47696), .Z(n47475) );
  XNOR U48056 ( .A(n47481), .B(n47479), .Z(n47696) );
  AND U48057 ( .A(n47697), .B(n47698), .Z(n47479) );
  NANDN U48058 ( .A(n47699), .B(n47700), .Z(n47698) );
  OR U48059 ( .A(n47701), .B(n47702), .Z(n47700) );
  NAND U48060 ( .A(n47702), .B(n47701), .Z(n47697) );
  ANDN U48061 ( .B(B[101]), .A(n67), .Z(n47481) );
  XNOR U48062 ( .A(n47489), .B(n47703), .Z(n47482) );
  XNOR U48063 ( .A(n47488), .B(n47486), .Z(n47703) );
  AND U48064 ( .A(n47704), .B(n47705), .Z(n47486) );
  NANDN U48065 ( .A(n47706), .B(n47707), .Z(n47705) );
  NANDN U48066 ( .A(n47708), .B(n47709), .Z(n47707) );
  NANDN U48067 ( .A(n47709), .B(n47708), .Z(n47704) );
  ANDN U48068 ( .B(B[102]), .A(n68), .Z(n47488) );
  XNOR U48069 ( .A(n47496), .B(n47710), .Z(n47489) );
  XNOR U48070 ( .A(n47495), .B(n47493), .Z(n47710) );
  AND U48071 ( .A(n47711), .B(n47712), .Z(n47493) );
  NANDN U48072 ( .A(n47713), .B(n47714), .Z(n47712) );
  OR U48073 ( .A(n47715), .B(n47716), .Z(n47714) );
  NAND U48074 ( .A(n47716), .B(n47715), .Z(n47711) );
  ANDN U48075 ( .B(B[103]), .A(n69), .Z(n47495) );
  XNOR U48076 ( .A(n47503), .B(n47717), .Z(n47496) );
  XNOR U48077 ( .A(n47502), .B(n47500), .Z(n47717) );
  AND U48078 ( .A(n47718), .B(n47719), .Z(n47500) );
  NANDN U48079 ( .A(n47720), .B(n47721), .Z(n47719) );
  NANDN U48080 ( .A(n47722), .B(n47723), .Z(n47721) );
  NANDN U48081 ( .A(n47723), .B(n47722), .Z(n47718) );
  ANDN U48082 ( .B(B[104]), .A(n70), .Z(n47502) );
  XNOR U48083 ( .A(n47510), .B(n47724), .Z(n47503) );
  XNOR U48084 ( .A(n47509), .B(n47507), .Z(n47724) );
  AND U48085 ( .A(n47725), .B(n47726), .Z(n47507) );
  NANDN U48086 ( .A(n47727), .B(n47728), .Z(n47726) );
  OR U48087 ( .A(n47729), .B(n47730), .Z(n47728) );
  NAND U48088 ( .A(n47730), .B(n47729), .Z(n47725) );
  ANDN U48089 ( .B(B[105]), .A(n71), .Z(n47509) );
  XNOR U48090 ( .A(n47517), .B(n47731), .Z(n47510) );
  XNOR U48091 ( .A(n47516), .B(n47514), .Z(n47731) );
  AND U48092 ( .A(n47732), .B(n47733), .Z(n47514) );
  NANDN U48093 ( .A(n47734), .B(n47735), .Z(n47733) );
  NANDN U48094 ( .A(n47736), .B(n47737), .Z(n47735) );
  NANDN U48095 ( .A(n47737), .B(n47736), .Z(n47732) );
  ANDN U48096 ( .B(B[106]), .A(n72), .Z(n47516) );
  XNOR U48097 ( .A(n47524), .B(n47738), .Z(n47517) );
  XNOR U48098 ( .A(n47523), .B(n47521), .Z(n47738) );
  AND U48099 ( .A(n47739), .B(n47740), .Z(n47521) );
  NANDN U48100 ( .A(n47741), .B(n47742), .Z(n47740) );
  OR U48101 ( .A(n47743), .B(n47744), .Z(n47742) );
  NAND U48102 ( .A(n47744), .B(n47743), .Z(n47739) );
  ANDN U48103 ( .B(B[107]), .A(n73), .Z(n47523) );
  XNOR U48104 ( .A(n47531), .B(n47745), .Z(n47524) );
  XNOR U48105 ( .A(n47530), .B(n47528), .Z(n47745) );
  AND U48106 ( .A(n47746), .B(n47747), .Z(n47528) );
  NANDN U48107 ( .A(n47748), .B(n47749), .Z(n47747) );
  NANDN U48108 ( .A(n47750), .B(n47751), .Z(n47749) );
  NANDN U48109 ( .A(n47751), .B(n47750), .Z(n47746) );
  ANDN U48110 ( .B(B[108]), .A(n74), .Z(n47530) );
  XNOR U48111 ( .A(n47538), .B(n47752), .Z(n47531) );
  XNOR U48112 ( .A(n47537), .B(n47535), .Z(n47752) );
  AND U48113 ( .A(n47753), .B(n47754), .Z(n47535) );
  NANDN U48114 ( .A(n47755), .B(n47756), .Z(n47754) );
  OR U48115 ( .A(n47757), .B(n47758), .Z(n47756) );
  NAND U48116 ( .A(n47758), .B(n47757), .Z(n47753) );
  ANDN U48117 ( .B(B[109]), .A(n75), .Z(n47537) );
  XNOR U48118 ( .A(n47545), .B(n47759), .Z(n47538) );
  XNOR U48119 ( .A(n47544), .B(n47542), .Z(n47759) );
  AND U48120 ( .A(n47760), .B(n47761), .Z(n47542) );
  NANDN U48121 ( .A(n47762), .B(n47763), .Z(n47761) );
  NANDN U48122 ( .A(n47764), .B(n47765), .Z(n47763) );
  NANDN U48123 ( .A(n47765), .B(n47764), .Z(n47760) );
  ANDN U48124 ( .B(B[110]), .A(n76), .Z(n47544) );
  XNOR U48125 ( .A(n47552), .B(n47766), .Z(n47545) );
  XNOR U48126 ( .A(n47551), .B(n47549), .Z(n47766) );
  AND U48127 ( .A(n47767), .B(n47768), .Z(n47549) );
  NANDN U48128 ( .A(n47769), .B(n47770), .Z(n47768) );
  OR U48129 ( .A(n47771), .B(n47772), .Z(n47770) );
  NAND U48130 ( .A(n47772), .B(n47771), .Z(n47767) );
  ANDN U48131 ( .B(B[111]), .A(n77), .Z(n47551) );
  XNOR U48132 ( .A(n47559), .B(n47773), .Z(n47552) );
  XNOR U48133 ( .A(n47558), .B(n47556), .Z(n47773) );
  AND U48134 ( .A(n47774), .B(n47775), .Z(n47556) );
  NANDN U48135 ( .A(n47776), .B(n47777), .Z(n47775) );
  NANDN U48136 ( .A(n47778), .B(n47779), .Z(n47777) );
  NANDN U48137 ( .A(n47779), .B(n47778), .Z(n47774) );
  ANDN U48138 ( .B(B[112]), .A(n78), .Z(n47558) );
  XNOR U48139 ( .A(n47566), .B(n47780), .Z(n47559) );
  XNOR U48140 ( .A(n47565), .B(n47563), .Z(n47780) );
  AND U48141 ( .A(n47781), .B(n47782), .Z(n47563) );
  NANDN U48142 ( .A(n47783), .B(n47784), .Z(n47782) );
  OR U48143 ( .A(n47785), .B(n47786), .Z(n47784) );
  NAND U48144 ( .A(n47786), .B(n47785), .Z(n47781) );
  ANDN U48145 ( .B(B[113]), .A(n79), .Z(n47565) );
  XNOR U48146 ( .A(n47573), .B(n47787), .Z(n47566) );
  XNOR U48147 ( .A(n47572), .B(n47570), .Z(n47787) );
  AND U48148 ( .A(n47788), .B(n47789), .Z(n47570) );
  NANDN U48149 ( .A(n47790), .B(n47791), .Z(n47789) );
  NANDN U48150 ( .A(n47792), .B(n47793), .Z(n47791) );
  NANDN U48151 ( .A(n47793), .B(n47792), .Z(n47788) );
  ANDN U48152 ( .B(B[114]), .A(n80), .Z(n47572) );
  XNOR U48153 ( .A(n47580), .B(n47794), .Z(n47573) );
  XNOR U48154 ( .A(n47579), .B(n47577), .Z(n47794) );
  AND U48155 ( .A(n47795), .B(n47796), .Z(n47577) );
  NANDN U48156 ( .A(n47797), .B(n47798), .Z(n47796) );
  OR U48157 ( .A(n47799), .B(n47800), .Z(n47798) );
  NAND U48158 ( .A(n47800), .B(n47799), .Z(n47795) );
  ANDN U48159 ( .B(B[115]), .A(n81), .Z(n47579) );
  XNOR U48160 ( .A(n47587), .B(n47801), .Z(n47580) );
  XNOR U48161 ( .A(n47586), .B(n47584), .Z(n47801) );
  AND U48162 ( .A(n47802), .B(n47803), .Z(n47584) );
  NANDN U48163 ( .A(n47804), .B(n47805), .Z(n47803) );
  NAND U48164 ( .A(n47806), .B(n47807), .Z(n47805) );
  ANDN U48165 ( .B(B[116]), .A(n82), .Z(n47586) );
  XOR U48166 ( .A(n47593), .B(n47808), .Z(n47587) );
  XNOR U48167 ( .A(n47591), .B(n47594), .Z(n47808) );
  NAND U48168 ( .A(A[2]), .B(B[117]), .Z(n47594) );
  NANDN U48169 ( .A(n47809), .B(n47810), .Z(n47591) );
  AND U48170 ( .A(A[0]), .B(B[118]), .Z(n47810) );
  XNOR U48171 ( .A(n47596), .B(n47811), .Z(n47593) );
  NAND U48172 ( .A(A[0]), .B(B[119]), .Z(n47811) );
  NAND U48173 ( .A(B[118]), .B(A[1]), .Z(n47596) );
  NAND U48174 ( .A(n47812), .B(n47813), .Z(n558) );
  NANDN U48175 ( .A(n47814), .B(n47815), .Z(n47813) );
  OR U48176 ( .A(n47816), .B(n47817), .Z(n47815) );
  NAND U48177 ( .A(n47817), .B(n47816), .Z(n47812) );
  XOR U48178 ( .A(n560), .B(n559), .Z(\A1[116] ) );
  XOR U48179 ( .A(n47817), .B(n47818), .Z(n559) );
  XNOR U48180 ( .A(n47816), .B(n47814), .Z(n47818) );
  AND U48181 ( .A(n47819), .B(n47820), .Z(n47814) );
  NANDN U48182 ( .A(n47821), .B(n47822), .Z(n47820) );
  NANDN U48183 ( .A(n47823), .B(n47824), .Z(n47822) );
  NANDN U48184 ( .A(n47824), .B(n47823), .Z(n47819) );
  ANDN U48185 ( .B(B[87]), .A(n54), .Z(n47816) );
  XNOR U48186 ( .A(n47611), .B(n47825), .Z(n47817) );
  XNOR U48187 ( .A(n47610), .B(n47608), .Z(n47825) );
  AND U48188 ( .A(n47826), .B(n47827), .Z(n47608) );
  NANDN U48189 ( .A(n47828), .B(n47829), .Z(n47827) );
  OR U48190 ( .A(n47830), .B(n47831), .Z(n47829) );
  NAND U48191 ( .A(n47831), .B(n47830), .Z(n47826) );
  ANDN U48192 ( .B(B[88]), .A(n55), .Z(n47610) );
  XNOR U48193 ( .A(n47618), .B(n47832), .Z(n47611) );
  XNOR U48194 ( .A(n47617), .B(n47615), .Z(n47832) );
  AND U48195 ( .A(n47833), .B(n47834), .Z(n47615) );
  NANDN U48196 ( .A(n47835), .B(n47836), .Z(n47834) );
  NANDN U48197 ( .A(n47837), .B(n47838), .Z(n47836) );
  NANDN U48198 ( .A(n47838), .B(n47837), .Z(n47833) );
  ANDN U48199 ( .B(B[89]), .A(n56), .Z(n47617) );
  XNOR U48200 ( .A(n47625), .B(n47839), .Z(n47618) );
  XNOR U48201 ( .A(n47624), .B(n47622), .Z(n47839) );
  AND U48202 ( .A(n47840), .B(n47841), .Z(n47622) );
  NANDN U48203 ( .A(n47842), .B(n47843), .Z(n47841) );
  OR U48204 ( .A(n47844), .B(n47845), .Z(n47843) );
  NAND U48205 ( .A(n47845), .B(n47844), .Z(n47840) );
  ANDN U48206 ( .B(B[90]), .A(n57), .Z(n47624) );
  XNOR U48207 ( .A(n47632), .B(n47846), .Z(n47625) );
  XNOR U48208 ( .A(n47631), .B(n47629), .Z(n47846) );
  AND U48209 ( .A(n47847), .B(n47848), .Z(n47629) );
  NANDN U48210 ( .A(n47849), .B(n47850), .Z(n47848) );
  NANDN U48211 ( .A(n47851), .B(n47852), .Z(n47850) );
  NANDN U48212 ( .A(n47852), .B(n47851), .Z(n47847) );
  ANDN U48213 ( .B(B[91]), .A(n58), .Z(n47631) );
  XNOR U48214 ( .A(n47639), .B(n47853), .Z(n47632) );
  XNOR U48215 ( .A(n47638), .B(n47636), .Z(n47853) );
  AND U48216 ( .A(n47854), .B(n47855), .Z(n47636) );
  NANDN U48217 ( .A(n47856), .B(n47857), .Z(n47855) );
  OR U48218 ( .A(n47858), .B(n47859), .Z(n47857) );
  NAND U48219 ( .A(n47859), .B(n47858), .Z(n47854) );
  ANDN U48220 ( .B(B[92]), .A(n59), .Z(n47638) );
  XNOR U48221 ( .A(n47646), .B(n47860), .Z(n47639) );
  XNOR U48222 ( .A(n47645), .B(n47643), .Z(n47860) );
  AND U48223 ( .A(n47861), .B(n47862), .Z(n47643) );
  NANDN U48224 ( .A(n47863), .B(n47864), .Z(n47862) );
  NANDN U48225 ( .A(n47865), .B(n47866), .Z(n47864) );
  NANDN U48226 ( .A(n47866), .B(n47865), .Z(n47861) );
  ANDN U48227 ( .B(A[25]), .A(n17), .Z(n47645) );
  XNOR U48228 ( .A(n47653), .B(n47867), .Z(n47646) );
  XNOR U48229 ( .A(n47652), .B(n47650), .Z(n47867) );
  AND U48230 ( .A(n47868), .B(n47869), .Z(n47650) );
  NANDN U48231 ( .A(n47870), .B(n47871), .Z(n47869) );
  OR U48232 ( .A(n47872), .B(n47873), .Z(n47871) );
  NAND U48233 ( .A(n47873), .B(n47872), .Z(n47868) );
  ANDN U48234 ( .B(A[24]), .A(n15), .Z(n47652) );
  XNOR U48235 ( .A(n47660), .B(n47874), .Z(n47653) );
  XNOR U48236 ( .A(n47659), .B(n47657), .Z(n47874) );
  AND U48237 ( .A(n47875), .B(n47876), .Z(n47657) );
  NANDN U48238 ( .A(n47877), .B(n47878), .Z(n47876) );
  NANDN U48239 ( .A(n47879), .B(n47880), .Z(n47878) );
  NANDN U48240 ( .A(n47880), .B(n47879), .Z(n47875) );
  ANDN U48241 ( .B(A[23]), .A(n13), .Z(n47659) );
  XNOR U48242 ( .A(n47667), .B(n47881), .Z(n47660) );
  XNOR U48243 ( .A(n47666), .B(n47664), .Z(n47881) );
  AND U48244 ( .A(n47882), .B(n47883), .Z(n47664) );
  NANDN U48245 ( .A(n47884), .B(n47885), .Z(n47883) );
  OR U48246 ( .A(n47886), .B(n47887), .Z(n47885) );
  NAND U48247 ( .A(n47887), .B(n47886), .Z(n47882) );
  ANDN U48248 ( .B(A[22]), .A(n11), .Z(n47666) );
  XNOR U48249 ( .A(n47674), .B(n47888), .Z(n47667) );
  XNOR U48250 ( .A(n47673), .B(n47671), .Z(n47888) );
  AND U48251 ( .A(n47889), .B(n47890), .Z(n47671) );
  NANDN U48252 ( .A(n47891), .B(n47892), .Z(n47890) );
  NANDN U48253 ( .A(n47893), .B(n47894), .Z(n47892) );
  NANDN U48254 ( .A(n47894), .B(n47893), .Z(n47889) );
  ANDN U48255 ( .B(A[21]), .A(n9), .Z(n47673) );
  XNOR U48256 ( .A(n47681), .B(n47895), .Z(n47674) );
  XNOR U48257 ( .A(n47680), .B(n47678), .Z(n47895) );
  AND U48258 ( .A(n47896), .B(n47897), .Z(n47678) );
  NANDN U48259 ( .A(n47898), .B(n47899), .Z(n47897) );
  OR U48260 ( .A(n47900), .B(n47901), .Z(n47899) );
  NAND U48261 ( .A(n47901), .B(n47900), .Z(n47896) );
  ANDN U48262 ( .B(B[98]), .A(n65), .Z(n47680) );
  XNOR U48263 ( .A(n47688), .B(n47902), .Z(n47681) );
  XNOR U48264 ( .A(n47687), .B(n47685), .Z(n47902) );
  AND U48265 ( .A(n47903), .B(n47904), .Z(n47685) );
  NANDN U48266 ( .A(n47905), .B(n47906), .Z(n47904) );
  NANDN U48267 ( .A(n47907), .B(n47908), .Z(n47906) );
  NANDN U48268 ( .A(n47908), .B(n47907), .Z(n47903) );
  ANDN U48269 ( .B(A[19]), .A(n6), .Z(n47687) );
  XNOR U48270 ( .A(n47695), .B(n47909), .Z(n47688) );
  XNOR U48271 ( .A(n47694), .B(n47692), .Z(n47909) );
  AND U48272 ( .A(n47910), .B(n47911), .Z(n47692) );
  NANDN U48273 ( .A(n47912), .B(n47913), .Z(n47911) );
  OR U48274 ( .A(n47914), .B(n47915), .Z(n47913) );
  NAND U48275 ( .A(n47915), .B(n47914), .Z(n47910) );
  ANDN U48276 ( .B(A[18]), .A(n4), .Z(n47694) );
  XNOR U48277 ( .A(n47702), .B(n47916), .Z(n47695) );
  XNOR U48278 ( .A(n47701), .B(n47699), .Z(n47916) );
  AND U48279 ( .A(n47917), .B(n47918), .Z(n47699) );
  NANDN U48280 ( .A(n47919), .B(n47920), .Z(n47918) );
  NANDN U48281 ( .A(n47921), .B(n47922), .Z(n47920) );
  NANDN U48282 ( .A(n47922), .B(n47921), .Z(n47917) );
  ANDN U48283 ( .B(B[101]), .A(n68), .Z(n47701) );
  XNOR U48284 ( .A(n47709), .B(n47923), .Z(n47702) );
  XNOR U48285 ( .A(n47708), .B(n47706), .Z(n47923) );
  AND U48286 ( .A(n47924), .B(n47925), .Z(n47706) );
  NANDN U48287 ( .A(n47926), .B(n47927), .Z(n47925) );
  OR U48288 ( .A(n47928), .B(n47929), .Z(n47927) );
  NAND U48289 ( .A(n47929), .B(n47928), .Z(n47924) );
  ANDN U48290 ( .B(B[102]), .A(n69), .Z(n47708) );
  XNOR U48291 ( .A(n47716), .B(n47930), .Z(n47709) );
  XNOR U48292 ( .A(n47715), .B(n47713), .Z(n47930) );
  AND U48293 ( .A(n47931), .B(n47932), .Z(n47713) );
  NANDN U48294 ( .A(n47933), .B(n47934), .Z(n47932) );
  NANDN U48295 ( .A(n47935), .B(n47936), .Z(n47934) );
  NANDN U48296 ( .A(n47936), .B(n47935), .Z(n47931) );
  ANDN U48297 ( .B(B[103]), .A(n70), .Z(n47715) );
  XNOR U48298 ( .A(n47723), .B(n47937), .Z(n47716) );
  XNOR U48299 ( .A(n47722), .B(n47720), .Z(n47937) );
  AND U48300 ( .A(n47938), .B(n47939), .Z(n47720) );
  NANDN U48301 ( .A(n47940), .B(n47941), .Z(n47939) );
  OR U48302 ( .A(n47942), .B(n47943), .Z(n47941) );
  NAND U48303 ( .A(n47943), .B(n47942), .Z(n47938) );
  ANDN U48304 ( .B(B[104]), .A(n71), .Z(n47722) );
  XNOR U48305 ( .A(n47730), .B(n47944), .Z(n47723) );
  XNOR U48306 ( .A(n47729), .B(n47727), .Z(n47944) );
  AND U48307 ( .A(n47945), .B(n47946), .Z(n47727) );
  NANDN U48308 ( .A(n47947), .B(n47948), .Z(n47946) );
  NANDN U48309 ( .A(n47949), .B(n47950), .Z(n47948) );
  NANDN U48310 ( .A(n47950), .B(n47949), .Z(n47945) );
  ANDN U48311 ( .B(B[105]), .A(n72), .Z(n47729) );
  XNOR U48312 ( .A(n47737), .B(n47951), .Z(n47730) );
  XNOR U48313 ( .A(n47736), .B(n47734), .Z(n47951) );
  AND U48314 ( .A(n47952), .B(n47953), .Z(n47734) );
  NANDN U48315 ( .A(n47954), .B(n47955), .Z(n47953) );
  OR U48316 ( .A(n47956), .B(n47957), .Z(n47955) );
  NAND U48317 ( .A(n47957), .B(n47956), .Z(n47952) );
  ANDN U48318 ( .B(B[106]), .A(n73), .Z(n47736) );
  XNOR U48319 ( .A(n47744), .B(n47958), .Z(n47737) );
  XNOR U48320 ( .A(n47743), .B(n47741), .Z(n47958) );
  AND U48321 ( .A(n47959), .B(n47960), .Z(n47741) );
  NANDN U48322 ( .A(n47961), .B(n47962), .Z(n47960) );
  NANDN U48323 ( .A(n47963), .B(n47964), .Z(n47962) );
  NANDN U48324 ( .A(n47964), .B(n47963), .Z(n47959) );
  ANDN U48325 ( .B(B[107]), .A(n74), .Z(n47743) );
  XNOR U48326 ( .A(n47751), .B(n47965), .Z(n47744) );
  XNOR U48327 ( .A(n47750), .B(n47748), .Z(n47965) );
  AND U48328 ( .A(n47966), .B(n47967), .Z(n47748) );
  NANDN U48329 ( .A(n47968), .B(n47969), .Z(n47967) );
  OR U48330 ( .A(n47970), .B(n47971), .Z(n47969) );
  NAND U48331 ( .A(n47971), .B(n47970), .Z(n47966) );
  ANDN U48332 ( .B(B[108]), .A(n75), .Z(n47750) );
  XNOR U48333 ( .A(n47758), .B(n47972), .Z(n47751) );
  XNOR U48334 ( .A(n47757), .B(n47755), .Z(n47972) );
  AND U48335 ( .A(n47973), .B(n47974), .Z(n47755) );
  NANDN U48336 ( .A(n47975), .B(n47976), .Z(n47974) );
  NANDN U48337 ( .A(n47977), .B(n47978), .Z(n47976) );
  NANDN U48338 ( .A(n47978), .B(n47977), .Z(n47973) );
  ANDN U48339 ( .B(B[109]), .A(n76), .Z(n47757) );
  XNOR U48340 ( .A(n47765), .B(n47979), .Z(n47758) );
  XNOR U48341 ( .A(n47764), .B(n47762), .Z(n47979) );
  AND U48342 ( .A(n47980), .B(n47981), .Z(n47762) );
  NANDN U48343 ( .A(n47982), .B(n47983), .Z(n47981) );
  OR U48344 ( .A(n47984), .B(n47985), .Z(n47983) );
  NAND U48345 ( .A(n47985), .B(n47984), .Z(n47980) );
  ANDN U48346 ( .B(B[110]), .A(n77), .Z(n47764) );
  XNOR U48347 ( .A(n47772), .B(n47986), .Z(n47765) );
  XNOR U48348 ( .A(n47771), .B(n47769), .Z(n47986) );
  AND U48349 ( .A(n47987), .B(n47988), .Z(n47769) );
  NANDN U48350 ( .A(n47989), .B(n47990), .Z(n47988) );
  NANDN U48351 ( .A(n47991), .B(n47992), .Z(n47990) );
  NANDN U48352 ( .A(n47992), .B(n47991), .Z(n47987) );
  ANDN U48353 ( .B(B[111]), .A(n78), .Z(n47771) );
  XNOR U48354 ( .A(n47779), .B(n47993), .Z(n47772) );
  XNOR U48355 ( .A(n47778), .B(n47776), .Z(n47993) );
  AND U48356 ( .A(n47994), .B(n47995), .Z(n47776) );
  NANDN U48357 ( .A(n47996), .B(n47997), .Z(n47995) );
  OR U48358 ( .A(n47998), .B(n47999), .Z(n47997) );
  NAND U48359 ( .A(n47999), .B(n47998), .Z(n47994) );
  ANDN U48360 ( .B(B[112]), .A(n79), .Z(n47778) );
  XNOR U48361 ( .A(n47786), .B(n48000), .Z(n47779) );
  XNOR U48362 ( .A(n47785), .B(n47783), .Z(n48000) );
  AND U48363 ( .A(n48001), .B(n48002), .Z(n47783) );
  NANDN U48364 ( .A(n48003), .B(n48004), .Z(n48002) );
  NANDN U48365 ( .A(n48005), .B(n48006), .Z(n48004) );
  NANDN U48366 ( .A(n48006), .B(n48005), .Z(n48001) );
  ANDN U48367 ( .B(B[113]), .A(n80), .Z(n47785) );
  XNOR U48368 ( .A(n47793), .B(n48007), .Z(n47786) );
  XNOR U48369 ( .A(n47792), .B(n47790), .Z(n48007) );
  AND U48370 ( .A(n48008), .B(n48009), .Z(n47790) );
  NANDN U48371 ( .A(n48010), .B(n48011), .Z(n48009) );
  OR U48372 ( .A(n48012), .B(n48013), .Z(n48011) );
  NAND U48373 ( .A(n48013), .B(n48012), .Z(n48008) );
  ANDN U48374 ( .B(B[114]), .A(n81), .Z(n47792) );
  XNOR U48375 ( .A(n47800), .B(n48014), .Z(n47793) );
  XNOR U48376 ( .A(n47799), .B(n47797), .Z(n48014) );
  AND U48377 ( .A(n48015), .B(n48016), .Z(n47797) );
  NANDN U48378 ( .A(n48017), .B(n48018), .Z(n48016) );
  NAND U48379 ( .A(n48019), .B(n48020), .Z(n48018) );
  ANDN U48380 ( .B(B[115]), .A(n82), .Z(n47799) );
  XOR U48381 ( .A(n47806), .B(n48021), .Z(n47800) );
  XNOR U48382 ( .A(n47804), .B(n47807), .Z(n48021) );
  NAND U48383 ( .A(A[2]), .B(B[116]), .Z(n47807) );
  NANDN U48384 ( .A(n48022), .B(n48023), .Z(n47804) );
  AND U48385 ( .A(A[0]), .B(B[117]), .Z(n48023) );
  XNOR U48386 ( .A(n47809), .B(n48024), .Z(n47806) );
  NAND U48387 ( .A(A[0]), .B(B[118]), .Z(n48024) );
  NAND U48388 ( .A(B[117]), .B(A[1]), .Z(n47809) );
  NAND U48389 ( .A(n48025), .B(n48026), .Z(n560) );
  NANDN U48390 ( .A(n48027), .B(n48028), .Z(n48026) );
  OR U48391 ( .A(n48029), .B(n48030), .Z(n48028) );
  NAND U48392 ( .A(n48030), .B(n48029), .Z(n48025) );
  XOR U48393 ( .A(n562), .B(n561), .Z(\A1[115] ) );
  XOR U48394 ( .A(n48030), .B(n48031), .Z(n561) );
  XNOR U48395 ( .A(n48029), .B(n48027), .Z(n48031) );
  AND U48396 ( .A(n48032), .B(n48033), .Z(n48027) );
  NANDN U48397 ( .A(n48034), .B(n48035), .Z(n48033) );
  NANDN U48398 ( .A(n48036), .B(n48037), .Z(n48035) );
  NANDN U48399 ( .A(n48037), .B(n48036), .Z(n48032) );
  ANDN U48400 ( .B(B[86]), .A(n54), .Z(n48029) );
  XNOR U48401 ( .A(n47824), .B(n48038), .Z(n48030) );
  XNOR U48402 ( .A(n47823), .B(n47821), .Z(n48038) );
  AND U48403 ( .A(n48039), .B(n48040), .Z(n47821) );
  NANDN U48404 ( .A(n48041), .B(n48042), .Z(n48040) );
  OR U48405 ( .A(n48043), .B(n48044), .Z(n48042) );
  NAND U48406 ( .A(n48044), .B(n48043), .Z(n48039) );
  ANDN U48407 ( .B(B[87]), .A(n55), .Z(n47823) );
  XNOR U48408 ( .A(n47831), .B(n48045), .Z(n47824) );
  XNOR U48409 ( .A(n47830), .B(n47828), .Z(n48045) );
  AND U48410 ( .A(n48046), .B(n48047), .Z(n47828) );
  NANDN U48411 ( .A(n48048), .B(n48049), .Z(n48047) );
  NANDN U48412 ( .A(n48050), .B(n48051), .Z(n48049) );
  NANDN U48413 ( .A(n48051), .B(n48050), .Z(n48046) );
  ANDN U48414 ( .B(B[88]), .A(n56), .Z(n47830) );
  XNOR U48415 ( .A(n47838), .B(n48052), .Z(n47831) );
  XNOR U48416 ( .A(n47837), .B(n47835), .Z(n48052) );
  AND U48417 ( .A(n48053), .B(n48054), .Z(n47835) );
  NANDN U48418 ( .A(n48055), .B(n48056), .Z(n48054) );
  OR U48419 ( .A(n48057), .B(n48058), .Z(n48056) );
  NAND U48420 ( .A(n48058), .B(n48057), .Z(n48053) );
  ANDN U48421 ( .B(B[89]), .A(n57), .Z(n47837) );
  XNOR U48422 ( .A(n47845), .B(n48059), .Z(n47838) );
  XNOR U48423 ( .A(n47844), .B(n47842), .Z(n48059) );
  AND U48424 ( .A(n48060), .B(n48061), .Z(n47842) );
  NANDN U48425 ( .A(n48062), .B(n48063), .Z(n48061) );
  NANDN U48426 ( .A(n48064), .B(n48065), .Z(n48063) );
  NANDN U48427 ( .A(n48065), .B(n48064), .Z(n48060) );
  ANDN U48428 ( .B(B[90]), .A(n58), .Z(n47844) );
  XNOR U48429 ( .A(n47852), .B(n48066), .Z(n47845) );
  XNOR U48430 ( .A(n47851), .B(n47849), .Z(n48066) );
  AND U48431 ( .A(n48067), .B(n48068), .Z(n47849) );
  NANDN U48432 ( .A(n48069), .B(n48070), .Z(n48068) );
  OR U48433 ( .A(n48071), .B(n48072), .Z(n48070) );
  NAND U48434 ( .A(n48072), .B(n48071), .Z(n48067) );
  ANDN U48435 ( .B(B[91]), .A(n59), .Z(n47851) );
  XNOR U48436 ( .A(n47859), .B(n48073), .Z(n47852) );
  XNOR U48437 ( .A(n47858), .B(n47856), .Z(n48073) );
  AND U48438 ( .A(n48074), .B(n48075), .Z(n47856) );
  NANDN U48439 ( .A(n48076), .B(n48077), .Z(n48075) );
  NANDN U48440 ( .A(n48078), .B(n48079), .Z(n48077) );
  NANDN U48441 ( .A(n48079), .B(n48078), .Z(n48074) );
  ANDN U48442 ( .B(B[92]), .A(n60), .Z(n47858) );
  XNOR U48443 ( .A(n47866), .B(n48080), .Z(n47859) );
  XNOR U48444 ( .A(n47865), .B(n47863), .Z(n48080) );
  AND U48445 ( .A(n48081), .B(n48082), .Z(n47863) );
  NANDN U48446 ( .A(n48083), .B(n48084), .Z(n48082) );
  OR U48447 ( .A(n48085), .B(n48086), .Z(n48084) );
  NAND U48448 ( .A(n48086), .B(n48085), .Z(n48081) );
  ANDN U48449 ( .B(A[24]), .A(n17), .Z(n47865) );
  XNOR U48450 ( .A(n47873), .B(n48087), .Z(n47866) );
  XNOR U48451 ( .A(n47872), .B(n47870), .Z(n48087) );
  AND U48452 ( .A(n48088), .B(n48089), .Z(n47870) );
  NANDN U48453 ( .A(n48090), .B(n48091), .Z(n48089) );
  NANDN U48454 ( .A(n48092), .B(n48093), .Z(n48091) );
  NANDN U48455 ( .A(n48093), .B(n48092), .Z(n48088) );
  ANDN U48456 ( .B(A[23]), .A(n15), .Z(n47872) );
  XNOR U48457 ( .A(n47880), .B(n48094), .Z(n47873) );
  XNOR U48458 ( .A(n47879), .B(n47877), .Z(n48094) );
  AND U48459 ( .A(n48095), .B(n48096), .Z(n47877) );
  NANDN U48460 ( .A(n48097), .B(n48098), .Z(n48096) );
  OR U48461 ( .A(n48099), .B(n48100), .Z(n48098) );
  NAND U48462 ( .A(n48100), .B(n48099), .Z(n48095) );
  ANDN U48463 ( .B(A[22]), .A(n13), .Z(n47879) );
  XNOR U48464 ( .A(n47887), .B(n48101), .Z(n47880) );
  XNOR U48465 ( .A(n47886), .B(n47884), .Z(n48101) );
  AND U48466 ( .A(n48102), .B(n48103), .Z(n47884) );
  NANDN U48467 ( .A(n48104), .B(n48105), .Z(n48103) );
  NANDN U48468 ( .A(n48106), .B(n48107), .Z(n48105) );
  NANDN U48469 ( .A(n48107), .B(n48106), .Z(n48102) );
  ANDN U48470 ( .B(A[21]), .A(n11), .Z(n47886) );
  XNOR U48471 ( .A(n47894), .B(n48108), .Z(n47887) );
  XNOR U48472 ( .A(n47893), .B(n47891), .Z(n48108) );
  AND U48473 ( .A(n48109), .B(n48110), .Z(n47891) );
  NANDN U48474 ( .A(n48111), .B(n48112), .Z(n48110) );
  OR U48475 ( .A(n48113), .B(n48114), .Z(n48112) );
  NAND U48476 ( .A(n48114), .B(n48113), .Z(n48109) );
  ANDN U48477 ( .B(A[20]), .A(n9), .Z(n47893) );
  XNOR U48478 ( .A(n47901), .B(n48115), .Z(n47894) );
  XNOR U48479 ( .A(n47900), .B(n47898), .Z(n48115) );
  AND U48480 ( .A(n48116), .B(n48117), .Z(n47898) );
  NANDN U48481 ( .A(n48118), .B(n48119), .Z(n48117) );
  NANDN U48482 ( .A(n48120), .B(n48121), .Z(n48119) );
  NANDN U48483 ( .A(n48121), .B(n48120), .Z(n48116) );
  ANDN U48484 ( .B(B[98]), .A(n66), .Z(n47900) );
  XNOR U48485 ( .A(n47908), .B(n48122), .Z(n47901) );
  XNOR U48486 ( .A(n47907), .B(n47905), .Z(n48122) );
  AND U48487 ( .A(n48123), .B(n48124), .Z(n47905) );
  NANDN U48488 ( .A(n48125), .B(n48126), .Z(n48124) );
  OR U48489 ( .A(n48127), .B(n48128), .Z(n48126) );
  NAND U48490 ( .A(n48128), .B(n48127), .Z(n48123) );
  ANDN U48491 ( .B(A[18]), .A(n6), .Z(n47907) );
  XNOR U48492 ( .A(n47915), .B(n48129), .Z(n47908) );
  XNOR U48493 ( .A(n47914), .B(n47912), .Z(n48129) );
  AND U48494 ( .A(n48130), .B(n48131), .Z(n47912) );
  NANDN U48495 ( .A(n48132), .B(n48133), .Z(n48131) );
  NANDN U48496 ( .A(n48134), .B(n48135), .Z(n48133) );
  NANDN U48497 ( .A(n48135), .B(n48134), .Z(n48130) );
  ANDN U48498 ( .B(A[17]), .A(n4), .Z(n47914) );
  XNOR U48499 ( .A(n47922), .B(n48136), .Z(n47915) );
  XNOR U48500 ( .A(n47921), .B(n47919), .Z(n48136) );
  AND U48501 ( .A(n48137), .B(n48138), .Z(n47919) );
  NANDN U48502 ( .A(n48139), .B(n48140), .Z(n48138) );
  OR U48503 ( .A(n48141), .B(n48142), .Z(n48140) );
  NAND U48504 ( .A(n48142), .B(n48141), .Z(n48137) );
  ANDN U48505 ( .B(B[101]), .A(n69), .Z(n47921) );
  XNOR U48506 ( .A(n47929), .B(n48143), .Z(n47922) );
  XNOR U48507 ( .A(n47928), .B(n47926), .Z(n48143) );
  AND U48508 ( .A(n48144), .B(n48145), .Z(n47926) );
  NANDN U48509 ( .A(n48146), .B(n48147), .Z(n48145) );
  NANDN U48510 ( .A(n48148), .B(n48149), .Z(n48147) );
  NANDN U48511 ( .A(n48149), .B(n48148), .Z(n48144) );
  ANDN U48512 ( .B(B[102]), .A(n70), .Z(n47928) );
  XNOR U48513 ( .A(n47936), .B(n48150), .Z(n47929) );
  XNOR U48514 ( .A(n47935), .B(n47933), .Z(n48150) );
  AND U48515 ( .A(n48151), .B(n48152), .Z(n47933) );
  NANDN U48516 ( .A(n48153), .B(n48154), .Z(n48152) );
  OR U48517 ( .A(n48155), .B(n48156), .Z(n48154) );
  NAND U48518 ( .A(n48156), .B(n48155), .Z(n48151) );
  ANDN U48519 ( .B(B[103]), .A(n71), .Z(n47935) );
  XNOR U48520 ( .A(n47943), .B(n48157), .Z(n47936) );
  XNOR U48521 ( .A(n47942), .B(n47940), .Z(n48157) );
  AND U48522 ( .A(n48158), .B(n48159), .Z(n47940) );
  NANDN U48523 ( .A(n48160), .B(n48161), .Z(n48159) );
  NANDN U48524 ( .A(n48162), .B(n48163), .Z(n48161) );
  NANDN U48525 ( .A(n48163), .B(n48162), .Z(n48158) );
  ANDN U48526 ( .B(B[104]), .A(n72), .Z(n47942) );
  XNOR U48527 ( .A(n47950), .B(n48164), .Z(n47943) );
  XNOR U48528 ( .A(n47949), .B(n47947), .Z(n48164) );
  AND U48529 ( .A(n48165), .B(n48166), .Z(n47947) );
  NANDN U48530 ( .A(n48167), .B(n48168), .Z(n48166) );
  OR U48531 ( .A(n48169), .B(n48170), .Z(n48168) );
  NAND U48532 ( .A(n48170), .B(n48169), .Z(n48165) );
  ANDN U48533 ( .B(B[105]), .A(n73), .Z(n47949) );
  XNOR U48534 ( .A(n47957), .B(n48171), .Z(n47950) );
  XNOR U48535 ( .A(n47956), .B(n47954), .Z(n48171) );
  AND U48536 ( .A(n48172), .B(n48173), .Z(n47954) );
  NANDN U48537 ( .A(n48174), .B(n48175), .Z(n48173) );
  NANDN U48538 ( .A(n48176), .B(n48177), .Z(n48175) );
  NANDN U48539 ( .A(n48177), .B(n48176), .Z(n48172) );
  ANDN U48540 ( .B(B[106]), .A(n74), .Z(n47956) );
  XNOR U48541 ( .A(n47964), .B(n48178), .Z(n47957) );
  XNOR U48542 ( .A(n47963), .B(n47961), .Z(n48178) );
  AND U48543 ( .A(n48179), .B(n48180), .Z(n47961) );
  NANDN U48544 ( .A(n48181), .B(n48182), .Z(n48180) );
  OR U48545 ( .A(n48183), .B(n48184), .Z(n48182) );
  NAND U48546 ( .A(n48184), .B(n48183), .Z(n48179) );
  ANDN U48547 ( .B(B[107]), .A(n75), .Z(n47963) );
  XNOR U48548 ( .A(n47971), .B(n48185), .Z(n47964) );
  XNOR U48549 ( .A(n47970), .B(n47968), .Z(n48185) );
  AND U48550 ( .A(n48186), .B(n48187), .Z(n47968) );
  NANDN U48551 ( .A(n48188), .B(n48189), .Z(n48187) );
  NANDN U48552 ( .A(n48190), .B(n48191), .Z(n48189) );
  NANDN U48553 ( .A(n48191), .B(n48190), .Z(n48186) );
  ANDN U48554 ( .B(B[108]), .A(n76), .Z(n47970) );
  XNOR U48555 ( .A(n47978), .B(n48192), .Z(n47971) );
  XNOR U48556 ( .A(n47977), .B(n47975), .Z(n48192) );
  AND U48557 ( .A(n48193), .B(n48194), .Z(n47975) );
  NANDN U48558 ( .A(n48195), .B(n48196), .Z(n48194) );
  OR U48559 ( .A(n48197), .B(n48198), .Z(n48196) );
  NAND U48560 ( .A(n48198), .B(n48197), .Z(n48193) );
  ANDN U48561 ( .B(B[109]), .A(n77), .Z(n47977) );
  XNOR U48562 ( .A(n47985), .B(n48199), .Z(n47978) );
  XNOR U48563 ( .A(n47984), .B(n47982), .Z(n48199) );
  AND U48564 ( .A(n48200), .B(n48201), .Z(n47982) );
  NANDN U48565 ( .A(n48202), .B(n48203), .Z(n48201) );
  NANDN U48566 ( .A(n48204), .B(n48205), .Z(n48203) );
  NANDN U48567 ( .A(n48205), .B(n48204), .Z(n48200) );
  ANDN U48568 ( .B(B[110]), .A(n78), .Z(n47984) );
  XNOR U48569 ( .A(n47992), .B(n48206), .Z(n47985) );
  XNOR U48570 ( .A(n47991), .B(n47989), .Z(n48206) );
  AND U48571 ( .A(n48207), .B(n48208), .Z(n47989) );
  NANDN U48572 ( .A(n48209), .B(n48210), .Z(n48208) );
  OR U48573 ( .A(n48211), .B(n48212), .Z(n48210) );
  NAND U48574 ( .A(n48212), .B(n48211), .Z(n48207) );
  ANDN U48575 ( .B(B[111]), .A(n79), .Z(n47991) );
  XNOR U48576 ( .A(n47999), .B(n48213), .Z(n47992) );
  XNOR U48577 ( .A(n47998), .B(n47996), .Z(n48213) );
  AND U48578 ( .A(n48214), .B(n48215), .Z(n47996) );
  NANDN U48579 ( .A(n48216), .B(n48217), .Z(n48215) );
  NANDN U48580 ( .A(n48218), .B(n48219), .Z(n48217) );
  NANDN U48581 ( .A(n48219), .B(n48218), .Z(n48214) );
  ANDN U48582 ( .B(B[112]), .A(n80), .Z(n47998) );
  XNOR U48583 ( .A(n48006), .B(n48220), .Z(n47999) );
  XNOR U48584 ( .A(n48005), .B(n48003), .Z(n48220) );
  AND U48585 ( .A(n48221), .B(n48222), .Z(n48003) );
  NANDN U48586 ( .A(n48223), .B(n48224), .Z(n48222) );
  OR U48587 ( .A(n48225), .B(n48226), .Z(n48224) );
  NAND U48588 ( .A(n48226), .B(n48225), .Z(n48221) );
  ANDN U48589 ( .B(B[113]), .A(n81), .Z(n48005) );
  XNOR U48590 ( .A(n48013), .B(n48227), .Z(n48006) );
  XNOR U48591 ( .A(n48012), .B(n48010), .Z(n48227) );
  AND U48592 ( .A(n48228), .B(n48229), .Z(n48010) );
  NANDN U48593 ( .A(n48230), .B(n48231), .Z(n48229) );
  NAND U48594 ( .A(n48232), .B(n48233), .Z(n48231) );
  ANDN U48595 ( .B(B[114]), .A(n82), .Z(n48012) );
  XOR U48596 ( .A(n48019), .B(n48234), .Z(n48013) );
  XNOR U48597 ( .A(n48017), .B(n48020), .Z(n48234) );
  NAND U48598 ( .A(A[2]), .B(B[115]), .Z(n48020) );
  NANDN U48599 ( .A(n48235), .B(n48236), .Z(n48017) );
  AND U48600 ( .A(A[0]), .B(B[116]), .Z(n48236) );
  XNOR U48601 ( .A(n48022), .B(n48237), .Z(n48019) );
  NAND U48602 ( .A(A[0]), .B(B[117]), .Z(n48237) );
  NAND U48603 ( .A(B[116]), .B(A[1]), .Z(n48022) );
  NAND U48604 ( .A(n48238), .B(n48239), .Z(n562) );
  NANDN U48605 ( .A(n48240), .B(n48241), .Z(n48239) );
  OR U48606 ( .A(n48242), .B(n48243), .Z(n48241) );
  NAND U48607 ( .A(n48243), .B(n48242), .Z(n48238) );
  XOR U48608 ( .A(n564), .B(n563), .Z(\A1[114] ) );
  XOR U48609 ( .A(n48243), .B(n48244), .Z(n563) );
  XNOR U48610 ( .A(n48242), .B(n48240), .Z(n48244) );
  AND U48611 ( .A(n48245), .B(n48246), .Z(n48240) );
  NANDN U48612 ( .A(n48247), .B(n48248), .Z(n48246) );
  NANDN U48613 ( .A(n48249), .B(n48250), .Z(n48248) );
  NANDN U48614 ( .A(n48250), .B(n48249), .Z(n48245) );
  ANDN U48615 ( .B(B[85]), .A(n54), .Z(n48242) );
  XNOR U48616 ( .A(n48037), .B(n48251), .Z(n48243) );
  XNOR U48617 ( .A(n48036), .B(n48034), .Z(n48251) );
  AND U48618 ( .A(n48252), .B(n48253), .Z(n48034) );
  NANDN U48619 ( .A(n48254), .B(n48255), .Z(n48253) );
  OR U48620 ( .A(n48256), .B(n48257), .Z(n48255) );
  NAND U48621 ( .A(n48257), .B(n48256), .Z(n48252) );
  ANDN U48622 ( .B(B[86]), .A(n55), .Z(n48036) );
  XNOR U48623 ( .A(n48044), .B(n48258), .Z(n48037) );
  XNOR U48624 ( .A(n48043), .B(n48041), .Z(n48258) );
  AND U48625 ( .A(n48259), .B(n48260), .Z(n48041) );
  NANDN U48626 ( .A(n48261), .B(n48262), .Z(n48260) );
  NANDN U48627 ( .A(n48263), .B(n48264), .Z(n48262) );
  NANDN U48628 ( .A(n48264), .B(n48263), .Z(n48259) );
  ANDN U48629 ( .B(B[87]), .A(n56), .Z(n48043) );
  XNOR U48630 ( .A(n48051), .B(n48265), .Z(n48044) );
  XNOR U48631 ( .A(n48050), .B(n48048), .Z(n48265) );
  AND U48632 ( .A(n48266), .B(n48267), .Z(n48048) );
  NANDN U48633 ( .A(n48268), .B(n48269), .Z(n48267) );
  OR U48634 ( .A(n48270), .B(n48271), .Z(n48269) );
  NAND U48635 ( .A(n48271), .B(n48270), .Z(n48266) );
  ANDN U48636 ( .B(B[88]), .A(n57), .Z(n48050) );
  XNOR U48637 ( .A(n48058), .B(n48272), .Z(n48051) );
  XNOR U48638 ( .A(n48057), .B(n48055), .Z(n48272) );
  AND U48639 ( .A(n48273), .B(n48274), .Z(n48055) );
  NANDN U48640 ( .A(n48275), .B(n48276), .Z(n48274) );
  NANDN U48641 ( .A(n48277), .B(n48278), .Z(n48276) );
  NANDN U48642 ( .A(n48278), .B(n48277), .Z(n48273) );
  ANDN U48643 ( .B(B[89]), .A(n58), .Z(n48057) );
  XNOR U48644 ( .A(n48065), .B(n48279), .Z(n48058) );
  XNOR U48645 ( .A(n48064), .B(n48062), .Z(n48279) );
  AND U48646 ( .A(n48280), .B(n48281), .Z(n48062) );
  NANDN U48647 ( .A(n48282), .B(n48283), .Z(n48281) );
  OR U48648 ( .A(n48284), .B(n48285), .Z(n48283) );
  NAND U48649 ( .A(n48285), .B(n48284), .Z(n48280) );
  ANDN U48650 ( .B(B[90]), .A(n59), .Z(n48064) );
  XNOR U48651 ( .A(n48072), .B(n48286), .Z(n48065) );
  XNOR U48652 ( .A(n48071), .B(n48069), .Z(n48286) );
  AND U48653 ( .A(n48287), .B(n48288), .Z(n48069) );
  NANDN U48654 ( .A(n48289), .B(n48290), .Z(n48288) );
  NANDN U48655 ( .A(n48291), .B(n48292), .Z(n48290) );
  NANDN U48656 ( .A(n48292), .B(n48291), .Z(n48287) );
  ANDN U48657 ( .B(B[91]), .A(n60), .Z(n48071) );
  XNOR U48658 ( .A(n48079), .B(n48293), .Z(n48072) );
  XNOR U48659 ( .A(n48078), .B(n48076), .Z(n48293) );
  AND U48660 ( .A(n48294), .B(n48295), .Z(n48076) );
  NANDN U48661 ( .A(n48296), .B(n48297), .Z(n48295) );
  OR U48662 ( .A(n48298), .B(n48299), .Z(n48297) );
  NAND U48663 ( .A(n48299), .B(n48298), .Z(n48294) );
  ANDN U48664 ( .B(A[24]), .A(n19), .Z(n48078) );
  XNOR U48665 ( .A(n48086), .B(n48300), .Z(n48079) );
  XNOR U48666 ( .A(n48085), .B(n48083), .Z(n48300) );
  AND U48667 ( .A(n48301), .B(n48302), .Z(n48083) );
  NANDN U48668 ( .A(n48303), .B(n48304), .Z(n48302) );
  NANDN U48669 ( .A(n48305), .B(n48306), .Z(n48304) );
  NANDN U48670 ( .A(n48306), .B(n48305), .Z(n48301) );
  ANDN U48671 ( .B(A[23]), .A(n17), .Z(n48085) );
  XNOR U48672 ( .A(n48093), .B(n48307), .Z(n48086) );
  XNOR U48673 ( .A(n48092), .B(n48090), .Z(n48307) );
  AND U48674 ( .A(n48308), .B(n48309), .Z(n48090) );
  NANDN U48675 ( .A(n48310), .B(n48311), .Z(n48309) );
  OR U48676 ( .A(n48312), .B(n48313), .Z(n48311) );
  NAND U48677 ( .A(n48313), .B(n48312), .Z(n48308) );
  ANDN U48678 ( .B(A[22]), .A(n15), .Z(n48092) );
  XNOR U48679 ( .A(n48100), .B(n48314), .Z(n48093) );
  XNOR U48680 ( .A(n48099), .B(n48097), .Z(n48314) );
  AND U48681 ( .A(n48315), .B(n48316), .Z(n48097) );
  NANDN U48682 ( .A(n48317), .B(n48318), .Z(n48316) );
  NANDN U48683 ( .A(n48319), .B(n48320), .Z(n48318) );
  NANDN U48684 ( .A(n48320), .B(n48319), .Z(n48315) );
  ANDN U48685 ( .B(A[21]), .A(n13), .Z(n48099) );
  XNOR U48686 ( .A(n48107), .B(n48321), .Z(n48100) );
  XNOR U48687 ( .A(n48106), .B(n48104), .Z(n48321) );
  AND U48688 ( .A(n48322), .B(n48323), .Z(n48104) );
  NANDN U48689 ( .A(n48324), .B(n48325), .Z(n48323) );
  OR U48690 ( .A(n48326), .B(n48327), .Z(n48325) );
  NAND U48691 ( .A(n48327), .B(n48326), .Z(n48322) );
  ANDN U48692 ( .B(A[20]), .A(n11), .Z(n48106) );
  XNOR U48693 ( .A(n48114), .B(n48328), .Z(n48107) );
  XNOR U48694 ( .A(n48113), .B(n48111), .Z(n48328) );
  AND U48695 ( .A(n48329), .B(n48330), .Z(n48111) );
  NANDN U48696 ( .A(n48331), .B(n48332), .Z(n48330) );
  NANDN U48697 ( .A(n48333), .B(n48334), .Z(n48332) );
  NANDN U48698 ( .A(n48334), .B(n48333), .Z(n48329) );
  ANDN U48699 ( .B(A[19]), .A(n9), .Z(n48113) );
  XNOR U48700 ( .A(n48121), .B(n48335), .Z(n48114) );
  XNOR U48701 ( .A(n48120), .B(n48118), .Z(n48335) );
  AND U48702 ( .A(n48336), .B(n48337), .Z(n48118) );
  NANDN U48703 ( .A(n48338), .B(n48339), .Z(n48337) );
  OR U48704 ( .A(n48340), .B(n48341), .Z(n48339) );
  NAND U48705 ( .A(n48341), .B(n48340), .Z(n48336) );
  ANDN U48706 ( .B(B[98]), .A(n67), .Z(n48120) );
  XNOR U48707 ( .A(n48128), .B(n48342), .Z(n48121) );
  XNOR U48708 ( .A(n48127), .B(n48125), .Z(n48342) );
  AND U48709 ( .A(n48343), .B(n48344), .Z(n48125) );
  NANDN U48710 ( .A(n48345), .B(n48346), .Z(n48344) );
  NANDN U48711 ( .A(n48347), .B(n48348), .Z(n48346) );
  NANDN U48712 ( .A(n48348), .B(n48347), .Z(n48343) );
  ANDN U48713 ( .B(A[17]), .A(n6), .Z(n48127) );
  XNOR U48714 ( .A(n48135), .B(n48349), .Z(n48128) );
  XNOR U48715 ( .A(n48134), .B(n48132), .Z(n48349) );
  AND U48716 ( .A(n48350), .B(n48351), .Z(n48132) );
  NANDN U48717 ( .A(n48352), .B(n48353), .Z(n48351) );
  OR U48718 ( .A(n48354), .B(n48355), .Z(n48353) );
  NAND U48719 ( .A(n48355), .B(n48354), .Z(n48350) );
  ANDN U48720 ( .B(A[16]), .A(n4), .Z(n48134) );
  XNOR U48721 ( .A(n48142), .B(n48356), .Z(n48135) );
  XNOR U48722 ( .A(n48141), .B(n48139), .Z(n48356) );
  AND U48723 ( .A(n48357), .B(n48358), .Z(n48139) );
  NANDN U48724 ( .A(n48359), .B(n48360), .Z(n48358) );
  NANDN U48725 ( .A(n48361), .B(n48362), .Z(n48360) );
  NANDN U48726 ( .A(n48362), .B(n48361), .Z(n48357) );
  ANDN U48727 ( .B(B[101]), .A(n70), .Z(n48141) );
  XNOR U48728 ( .A(n48149), .B(n48363), .Z(n48142) );
  XNOR U48729 ( .A(n48148), .B(n48146), .Z(n48363) );
  AND U48730 ( .A(n48364), .B(n48365), .Z(n48146) );
  NANDN U48731 ( .A(n48366), .B(n48367), .Z(n48365) );
  OR U48732 ( .A(n48368), .B(n48369), .Z(n48367) );
  NAND U48733 ( .A(n48369), .B(n48368), .Z(n48364) );
  ANDN U48734 ( .B(B[102]), .A(n71), .Z(n48148) );
  XNOR U48735 ( .A(n48156), .B(n48370), .Z(n48149) );
  XNOR U48736 ( .A(n48155), .B(n48153), .Z(n48370) );
  AND U48737 ( .A(n48371), .B(n48372), .Z(n48153) );
  NANDN U48738 ( .A(n48373), .B(n48374), .Z(n48372) );
  NANDN U48739 ( .A(n48375), .B(n48376), .Z(n48374) );
  NANDN U48740 ( .A(n48376), .B(n48375), .Z(n48371) );
  ANDN U48741 ( .B(B[103]), .A(n72), .Z(n48155) );
  XNOR U48742 ( .A(n48163), .B(n48377), .Z(n48156) );
  XNOR U48743 ( .A(n48162), .B(n48160), .Z(n48377) );
  AND U48744 ( .A(n48378), .B(n48379), .Z(n48160) );
  NANDN U48745 ( .A(n48380), .B(n48381), .Z(n48379) );
  OR U48746 ( .A(n48382), .B(n48383), .Z(n48381) );
  NAND U48747 ( .A(n48383), .B(n48382), .Z(n48378) );
  ANDN U48748 ( .B(B[104]), .A(n73), .Z(n48162) );
  XNOR U48749 ( .A(n48170), .B(n48384), .Z(n48163) );
  XNOR U48750 ( .A(n48169), .B(n48167), .Z(n48384) );
  AND U48751 ( .A(n48385), .B(n48386), .Z(n48167) );
  NANDN U48752 ( .A(n48387), .B(n48388), .Z(n48386) );
  NANDN U48753 ( .A(n48389), .B(n48390), .Z(n48388) );
  NANDN U48754 ( .A(n48390), .B(n48389), .Z(n48385) );
  ANDN U48755 ( .B(B[105]), .A(n74), .Z(n48169) );
  XNOR U48756 ( .A(n48177), .B(n48391), .Z(n48170) );
  XNOR U48757 ( .A(n48176), .B(n48174), .Z(n48391) );
  AND U48758 ( .A(n48392), .B(n48393), .Z(n48174) );
  NANDN U48759 ( .A(n48394), .B(n48395), .Z(n48393) );
  OR U48760 ( .A(n48396), .B(n48397), .Z(n48395) );
  NAND U48761 ( .A(n48397), .B(n48396), .Z(n48392) );
  ANDN U48762 ( .B(B[106]), .A(n75), .Z(n48176) );
  XNOR U48763 ( .A(n48184), .B(n48398), .Z(n48177) );
  XNOR U48764 ( .A(n48183), .B(n48181), .Z(n48398) );
  AND U48765 ( .A(n48399), .B(n48400), .Z(n48181) );
  NANDN U48766 ( .A(n48401), .B(n48402), .Z(n48400) );
  NANDN U48767 ( .A(n48403), .B(n48404), .Z(n48402) );
  NANDN U48768 ( .A(n48404), .B(n48403), .Z(n48399) );
  ANDN U48769 ( .B(B[107]), .A(n76), .Z(n48183) );
  XNOR U48770 ( .A(n48191), .B(n48405), .Z(n48184) );
  XNOR U48771 ( .A(n48190), .B(n48188), .Z(n48405) );
  AND U48772 ( .A(n48406), .B(n48407), .Z(n48188) );
  NANDN U48773 ( .A(n48408), .B(n48409), .Z(n48407) );
  OR U48774 ( .A(n48410), .B(n48411), .Z(n48409) );
  NAND U48775 ( .A(n48411), .B(n48410), .Z(n48406) );
  ANDN U48776 ( .B(B[108]), .A(n77), .Z(n48190) );
  XNOR U48777 ( .A(n48198), .B(n48412), .Z(n48191) );
  XNOR U48778 ( .A(n48197), .B(n48195), .Z(n48412) );
  AND U48779 ( .A(n48413), .B(n48414), .Z(n48195) );
  NANDN U48780 ( .A(n48415), .B(n48416), .Z(n48414) );
  NANDN U48781 ( .A(n48417), .B(n48418), .Z(n48416) );
  NANDN U48782 ( .A(n48418), .B(n48417), .Z(n48413) );
  ANDN U48783 ( .B(B[109]), .A(n78), .Z(n48197) );
  XNOR U48784 ( .A(n48205), .B(n48419), .Z(n48198) );
  XNOR U48785 ( .A(n48204), .B(n48202), .Z(n48419) );
  AND U48786 ( .A(n48420), .B(n48421), .Z(n48202) );
  NANDN U48787 ( .A(n48422), .B(n48423), .Z(n48421) );
  OR U48788 ( .A(n48424), .B(n48425), .Z(n48423) );
  NAND U48789 ( .A(n48425), .B(n48424), .Z(n48420) );
  ANDN U48790 ( .B(B[110]), .A(n79), .Z(n48204) );
  XNOR U48791 ( .A(n48212), .B(n48426), .Z(n48205) );
  XNOR U48792 ( .A(n48211), .B(n48209), .Z(n48426) );
  AND U48793 ( .A(n48427), .B(n48428), .Z(n48209) );
  NANDN U48794 ( .A(n48429), .B(n48430), .Z(n48428) );
  NANDN U48795 ( .A(n48431), .B(n48432), .Z(n48430) );
  NANDN U48796 ( .A(n48432), .B(n48431), .Z(n48427) );
  ANDN U48797 ( .B(B[111]), .A(n80), .Z(n48211) );
  XNOR U48798 ( .A(n48219), .B(n48433), .Z(n48212) );
  XNOR U48799 ( .A(n48218), .B(n48216), .Z(n48433) );
  AND U48800 ( .A(n48434), .B(n48435), .Z(n48216) );
  NANDN U48801 ( .A(n48436), .B(n48437), .Z(n48435) );
  OR U48802 ( .A(n48438), .B(n48439), .Z(n48437) );
  NAND U48803 ( .A(n48439), .B(n48438), .Z(n48434) );
  ANDN U48804 ( .B(B[112]), .A(n81), .Z(n48218) );
  XNOR U48805 ( .A(n48226), .B(n48440), .Z(n48219) );
  XNOR U48806 ( .A(n48225), .B(n48223), .Z(n48440) );
  AND U48807 ( .A(n48441), .B(n48442), .Z(n48223) );
  NANDN U48808 ( .A(n48443), .B(n48444), .Z(n48442) );
  NAND U48809 ( .A(n48445), .B(n48446), .Z(n48444) );
  ANDN U48810 ( .B(B[113]), .A(n82), .Z(n48225) );
  XOR U48811 ( .A(n48232), .B(n48447), .Z(n48226) );
  XNOR U48812 ( .A(n48230), .B(n48233), .Z(n48447) );
  NAND U48813 ( .A(A[2]), .B(B[114]), .Z(n48233) );
  NANDN U48814 ( .A(n48448), .B(n48449), .Z(n48230) );
  AND U48815 ( .A(A[0]), .B(B[115]), .Z(n48449) );
  XNOR U48816 ( .A(n48235), .B(n48450), .Z(n48232) );
  NAND U48817 ( .A(A[0]), .B(B[116]), .Z(n48450) );
  NAND U48818 ( .A(B[115]), .B(A[1]), .Z(n48235) );
  NAND U48819 ( .A(n48451), .B(n48452), .Z(n564) );
  NANDN U48820 ( .A(n48453), .B(n48454), .Z(n48452) );
  OR U48821 ( .A(n48455), .B(n48456), .Z(n48454) );
  NAND U48822 ( .A(n48456), .B(n48455), .Z(n48451) );
  XOR U48823 ( .A(n566), .B(n565), .Z(\A1[113] ) );
  XOR U48824 ( .A(n48456), .B(n48457), .Z(n565) );
  XNOR U48825 ( .A(n48455), .B(n48453), .Z(n48457) );
  AND U48826 ( .A(n48458), .B(n48459), .Z(n48453) );
  NANDN U48827 ( .A(n48460), .B(n48461), .Z(n48459) );
  NANDN U48828 ( .A(n48462), .B(n48463), .Z(n48461) );
  NANDN U48829 ( .A(n48463), .B(n48462), .Z(n48458) );
  ANDN U48830 ( .B(B[84]), .A(n54), .Z(n48455) );
  XNOR U48831 ( .A(n48250), .B(n48464), .Z(n48456) );
  XNOR U48832 ( .A(n48249), .B(n48247), .Z(n48464) );
  AND U48833 ( .A(n48465), .B(n48466), .Z(n48247) );
  NANDN U48834 ( .A(n48467), .B(n48468), .Z(n48466) );
  OR U48835 ( .A(n48469), .B(n48470), .Z(n48468) );
  NAND U48836 ( .A(n48470), .B(n48469), .Z(n48465) );
  ANDN U48837 ( .B(B[85]), .A(n55), .Z(n48249) );
  XNOR U48838 ( .A(n48257), .B(n48471), .Z(n48250) );
  XNOR U48839 ( .A(n48256), .B(n48254), .Z(n48471) );
  AND U48840 ( .A(n48472), .B(n48473), .Z(n48254) );
  NANDN U48841 ( .A(n48474), .B(n48475), .Z(n48473) );
  NANDN U48842 ( .A(n48476), .B(n48477), .Z(n48475) );
  NANDN U48843 ( .A(n48477), .B(n48476), .Z(n48472) );
  ANDN U48844 ( .B(B[86]), .A(n56), .Z(n48256) );
  XNOR U48845 ( .A(n48264), .B(n48478), .Z(n48257) );
  XNOR U48846 ( .A(n48263), .B(n48261), .Z(n48478) );
  AND U48847 ( .A(n48479), .B(n48480), .Z(n48261) );
  NANDN U48848 ( .A(n48481), .B(n48482), .Z(n48480) );
  OR U48849 ( .A(n48483), .B(n48484), .Z(n48482) );
  NAND U48850 ( .A(n48484), .B(n48483), .Z(n48479) );
  ANDN U48851 ( .B(B[87]), .A(n57), .Z(n48263) );
  XNOR U48852 ( .A(n48271), .B(n48485), .Z(n48264) );
  XNOR U48853 ( .A(n48270), .B(n48268), .Z(n48485) );
  AND U48854 ( .A(n48486), .B(n48487), .Z(n48268) );
  NANDN U48855 ( .A(n48488), .B(n48489), .Z(n48487) );
  NANDN U48856 ( .A(n48490), .B(n48491), .Z(n48489) );
  NANDN U48857 ( .A(n48491), .B(n48490), .Z(n48486) );
  ANDN U48858 ( .B(B[88]), .A(n58), .Z(n48270) );
  XNOR U48859 ( .A(n48278), .B(n48492), .Z(n48271) );
  XNOR U48860 ( .A(n48277), .B(n48275), .Z(n48492) );
  AND U48861 ( .A(n48493), .B(n48494), .Z(n48275) );
  NANDN U48862 ( .A(n48495), .B(n48496), .Z(n48494) );
  OR U48863 ( .A(n48497), .B(n48498), .Z(n48496) );
  NAND U48864 ( .A(n48498), .B(n48497), .Z(n48493) );
  ANDN U48865 ( .B(B[89]), .A(n59), .Z(n48277) );
  XNOR U48866 ( .A(n48285), .B(n48499), .Z(n48278) );
  XNOR U48867 ( .A(n48284), .B(n48282), .Z(n48499) );
  AND U48868 ( .A(n48500), .B(n48501), .Z(n48282) );
  NANDN U48869 ( .A(n48502), .B(n48503), .Z(n48501) );
  NANDN U48870 ( .A(n48504), .B(n48505), .Z(n48503) );
  NANDN U48871 ( .A(n48505), .B(n48504), .Z(n48500) );
  ANDN U48872 ( .B(B[90]), .A(n60), .Z(n48284) );
  XNOR U48873 ( .A(n48292), .B(n48506), .Z(n48285) );
  XNOR U48874 ( .A(n48291), .B(n48289), .Z(n48506) );
  AND U48875 ( .A(n48507), .B(n48508), .Z(n48289) );
  NANDN U48876 ( .A(n48509), .B(n48510), .Z(n48508) );
  OR U48877 ( .A(n48511), .B(n48512), .Z(n48510) );
  NAND U48878 ( .A(n48512), .B(n48511), .Z(n48507) );
  ANDN U48879 ( .B(B[91]), .A(n61), .Z(n48291) );
  XNOR U48880 ( .A(n48299), .B(n48513), .Z(n48292) );
  XNOR U48881 ( .A(n48298), .B(n48296), .Z(n48513) );
  AND U48882 ( .A(n48514), .B(n48515), .Z(n48296) );
  NANDN U48883 ( .A(n48516), .B(n48517), .Z(n48515) );
  NANDN U48884 ( .A(n48518), .B(n48519), .Z(n48517) );
  NANDN U48885 ( .A(n48519), .B(n48518), .Z(n48514) );
  ANDN U48886 ( .B(A[23]), .A(n19), .Z(n48298) );
  XNOR U48887 ( .A(n48306), .B(n48520), .Z(n48299) );
  XNOR U48888 ( .A(n48305), .B(n48303), .Z(n48520) );
  AND U48889 ( .A(n48521), .B(n48522), .Z(n48303) );
  NANDN U48890 ( .A(n48523), .B(n48524), .Z(n48522) );
  OR U48891 ( .A(n48525), .B(n48526), .Z(n48524) );
  NAND U48892 ( .A(n48526), .B(n48525), .Z(n48521) );
  ANDN U48893 ( .B(A[22]), .A(n17), .Z(n48305) );
  XNOR U48894 ( .A(n48313), .B(n48527), .Z(n48306) );
  XNOR U48895 ( .A(n48312), .B(n48310), .Z(n48527) );
  AND U48896 ( .A(n48528), .B(n48529), .Z(n48310) );
  NANDN U48897 ( .A(n48530), .B(n48531), .Z(n48529) );
  NANDN U48898 ( .A(n48532), .B(n48533), .Z(n48531) );
  NANDN U48899 ( .A(n48533), .B(n48532), .Z(n48528) );
  ANDN U48900 ( .B(A[21]), .A(n15), .Z(n48312) );
  XNOR U48901 ( .A(n48320), .B(n48534), .Z(n48313) );
  XNOR U48902 ( .A(n48319), .B(n48317), .Z(n48534) );
  AND U48903 ( .A(n48535), .B(n48536), .Z(n48317) );
  NANDN U48904 ( .A(n48537), .B(n48538), .Z(n48536) );
  OR U48905 ( .A(n48539), .B(n48540), .Z(n48538) );
  NAND U48906 ( .A(n48540), .B(n48539), .Z(n48535) );
  ANDN U48907 ( .B(A[20]), .A(n13), .Z(n48319) );
  XNOR U48908 ( .A(n48327), .B(n48541), .Z(n48320) );
  XNOR U48909 ( .A(n48326), .B(n48324), .Z(n48541) );
  AND U48910 ( .A(n48542), .B(n48543), .Z(n48324) );
  NANDN U48911 ( .A(n48544), .B(n48545), .Z(n48543) );
  NANDN U48912 ( .A(n48546), .B(n48547), .Z(n48545) );
  NANDN U48913 ( .A(n48547), .B(n48546), .Z(n48542) );
  ANDN U48914 ( .B(A[19]), .A(n11), .Z(n48326) );
  XNOR U48915 ( .A(n48334), .B(n48548), .Z(n48327) );
  XNOR U48916 ( .A(n48333), .B(n48331), .Z(n48548) );
  AND U48917 ( .A(n48549), .B(n48550), .Z(n48331) );
  NANDN U48918 ( .A(n48551), .B(n48552), .Z(n48550) );
  OR U48919 ( .A(n48553), .B(n48554), .Z(n48552) );
  NAND U48920 ( .A(n48554), .B(n48553), .Z(n48549) );
  ANDN U48921 ( .B(A[18]), .A(n9), .Z(n48333) );
  XNOR U48922 ( .A(n48341), .B(n48555), .Z(n48334) );
  XNOR U48923 ( .A(n48340), .B(n48338), .Z(n48555) );
  AND U48924 ( .A(n48556), .B(n48557), .Z(n48338) );
  NANDN U48925 ( .A(n48558), .B(n48559), .Z(n48557) );
  NANDN U48926 ( .A(n48560), .B(n48561), .Z(n48559) );
  NANDN U48927 ( .A(n48561), .B(n48560), .Z(n48556) );
  ANDN U48928 ( .B(B[98]), .A(n68), .Z(n48340) );
  XNOR U48929 ( .A(n48348), .B(n48562), .Z(n48341) );
  XNOR U48930 ( .A(n48347), .B(n48345), .Z(n48562) );
  AND U48931 ( .A(n48563), .B(n48564), .Z(n48345) );
  NANDN U48932 ( .A(n48565), .B(n48566), .Z(n48564) );
  OR U48933 ( .A(n48567), .B(n48568), .Z(n48566) );
  NAND U48934 ( .A(n48568), .B(n48567), .Z(n48563) );
  ANDN U48935 ( .B(A[16]), .A(n6), .Z(n48347) );
  XNOR U48936 ( .A(n48355), .B(n48569), .Z(n48348) );
  XNOR U48937 ( .A(n48354), .B(n48352), .Z(n48569) );
  AND U48938 ( .A(n48570), .B(n48571), .Z(n48352) );
  NANDN U48939 ( .A(n48572), .B(n48573), .Z(n48571) );
  NANDN U48940 ( .A(n48574), .B(n48575), .Z(n48573) );
  NANDN U48941 ( .A(n48575), .B(n48574), .Z(n48570) );
  ANDN U48942 ( .B(A[15]), .A(n4), .Z(n48354) );
  XNOR U48943 ( .A(n48362), .B(n48576), .Z(n48355) );
  XNOR U48944 ( .A(n48361), .B(n48359), .Z(n48576) );
  AND U48945 ( .A(n48577), .B(n48578), .Z(n48359) );
  NANDN U48946 ( .A(n48579), .B(n48580), .Z(n48578) );
  OR U48947 ( .A(n48581), .B(n48582), .Z(n48580) );
  NAND U48948 ( .A(n48582), .B(n48581), .Z(n48577) );
  ANDN U48949 ( .B(B[101]), .A(n71), .Z(n48361) );
  XNOR U48950 ( .A(n48369), .B(n48583), .Z(n48362) );
  XNOR U48951 ( .A(n48368), .B(n48366), .Z(n48583) );
  AND U48952 ( .A(n48584), .B(n48585), .Z(n48366) );
  NANDN U48953 ( .A(n48586), .B(n48587), .Z(n48585) );
  NANDN U48954 ( .A(n48588), .B(n48589), .Z(n48587) );
  NANDN U48955 ( .A(n48589), .B(n48588), .Z(n48584) );
  ANDN U48956 ( .B(B[102]), .A(n72), .Z(n48368) );
  XNOR U48957 ( .A(n48376), .B(n48590), .Z(n48369) );
  XNOR U48958 ( .A(n48375), .B(n48373), .Z(n48590) );
  AND U48959 ( .A(n48591), .B(n48592), .Z(n48373) );
  NANDN U48960 ( .A(n48593), .B(n48594), .Z(n48592) );
  OR U48961 ( .A(n48595), .B(n48596), .Z(n48594) );
  NAND U48962 ( .A(n48596), .B(n48595), .Z(n48591) );
  ANDN U48963 ( .B(B[103]), .A(n73), .Z(n48375) );
  XNOR U48964 ( .A(n48383), .B(n48597), .Z(n48376) );
  XNOR U48965 ( .A(n48382), .B(n48380), .Z(n48597) );
  AND U48966 ( .A(n48598), .B(n48599), .Z(n48380) );
  NANDN U48967 ( .A(n48600), .B(n48601), .Z(n48599) );
  NANDN U48968 ( .A(n48602), .B(n48603), .Z(n48601) );
  NANDN U48969 ( .A(n48603), .B(n48602), .Z(n48598) );
  ANDN U48970 ( .B(B[104]), .A(n74), .Z(n48382) );
  XNOR U48971 ( .A(n48390), .B(n48604), .Z(n48383) );
  XNOR U48972 ( .A(n48389), .B(n48387), .Z(n48604) );
  AND U48973 ( .A(n48605), .B(n48606), .Z(n48387) );
  NANDN U48974 ( .A(n48607), .B(n48608), .Z(n48606) );
  OR U48975 ( .A(n48609), .B(n48610), .Z(n48608) );
  NAND U48976 ( .A(n48610), .B(n48609), .Z(n48605) );
  ANDN U48977 ( .B(B[105]), .A(n75), .Z(n48389) );
  XNOR U48978 ( .A(n48397), .B(n48611), .Z(n48390) );
  XNOR U48979 ( .A(n48396), .B(n48394), .Z(n48611) );
  AND U48980 ( .A(n48612), .B(n48613), .Z(n48394) );
  NANDN U48981 ( .A(n48614), .B(n48615), .Z(n48613) );
  NANDN U48982 ( .A(n48616), .B(n48617), .Z(n48615) );
  NANDN U48983 ( .A(n48617), .B(n48616), .Z(n48612) );
  ANDN U48984 ( .B(B[106]), .A(n76), .Z(n48396) );
  XNOR U48985 ( .A(n48404), .B(n48618), .Z(n48397) );
  XNOR U48986 ( .A(n48403), .B(n48401), .Z(n48618) );
  AND U48987 ( .A(n48619), .B(n48620), .Z(n48401) );
  NANDN U48988 ( .A(n48621), .B(n48622), .Z(n48620) );
  OR U48989 ( .A(n48623), .B(n48624), .Z(n48622) );
  NAND U48990 ( .A(n48624), .B(n48623), .Z(n48619) );
  ANDN U48991 ( .B(B[107]), .A(n77), .Z(n48403) );
  XNOR U48992 ( .A(n48411), .B(n48625), .Z(n48404) );
  XNOR U48993 ( .A(n48410), .B(n48408), .Z(n48625) );
  AND U48994 ( .A(n48626), .B(n48627), .Z(n48408) );
  NANDN U48995 ( .A(n48628), .B(n48629), .Z(n48627) );
  NANDN U48996 ( .A(n48630), .B(n48631), .Z(n48629) );
  NANDN U48997 ( .A(n48631), .B(n48630), .Z(n48626) );
  ANDN U48998 ( .B(B[108]), .A(n78), .Z(n48410) );
  XNOR U48999 ( .A(n48418), .B(n48632), .Z(n48411) );
  XNOR U49000 ( .A(n48417), .B(n48415), .Z(n48632) );
  AND U49001 ( .A(n48633), .B(n48634), .Z(n48415) );
  NANDN U49002 ( .A(n48635), .B(n48636), .Z(n48634) );
  OR U49003 ( .A(n48637), .B(n48638), .Z(n48636) );
  NAND U49004 ( .A(n48638), .B(n48637), .Z(n48633) );
  ANDN U49005 ( .B(B[109]), .A(n79), .Z(n48417) );
  XNOR U49006 ( .A(n48425), .B(n48639), .Z(n48418) );
  XNOR U49007 ( .A(n48424), .B(n48422), .Z(n48639) );
  AND U49008 ( .A(n48640), .B(n48641), .Z(n48422) );
  NANDN U49009 ( .A(n48642), .B(n48643), .Z(n48641) );
  NANDN U49010 ( .A(n48644), .B(n48645), .Z(n48643) );
  NANDN U49011 ( .A(n48645), .B(n48644), .Z(n48640) );
  ANDN U49012 ( .B(B[110]), .A(n80), .Z(n48424) );
  XNOR U49013 ( .A(n48432), .B(n48646), .Z(n48425) );
  XNOR U49014 ( .A(n48431), .B(n48429), .Z(n48646) );
  AND U49015 ( .A(n48647), .B(n48648), .Z(n48429) );
  NANDN U49016 ( .A(n48649), .B(n48650), .Z(n48648) );
  OR U49017 ( .A(n48651), .B(n48652), .Z(n48650) );
  NAND U49018 ( .A(n48652), .B(n48651), .Z(n48647) );
  ANDN U49019 ( .B(B[111]), .A(n81), .Z(n48431) );
  XNOR U49020 ( .A(n48439), .B(n48653), .Z(n48432) );
  XNOR U49021 ( .A(n48438), .B(n48436), .Z(n48653) );
  AND U49022 ( .A(n48654), .B(n48655), .Z(n48436) );
  NANDN U49023 ( .A(n48656), .B(n48657), .Z(n48655) );
  NAND U49024 ( .A(n48658), .B(n48659), .Z(n48657) );
  ANDN U49025 ( .B(B[112]), .A(n82), .Z(n48438) );
  XOR U49026 ( .A(n48445), .B(n48660), .Z(n48439) );
  XNOR U49027 ( .A(n48443), .B(n48446), .Z(n48660) );
  NAND U49028 ( .A(A[2]), .B(B[113]), .Z(n48446) );
  NANDN U49029 ( .A(n48661), .B(n48662), .Z(n48443) );
  AND U49030 ( .A(A[0]), .B(B[114]), .Z(n48662) );
  XNOR U49031 ( .A(n48448), .B(n48663), .Z(n48445) );
  NAND U49032 ( .A(A[0]), .B(B[115]), .Z(n48663) );
  NAND U49033 ( .A(B[114]), .B(A[1]), .Z(n48448) );
  NAND U49034 ( .A(n48664), .B(n48665), .Z(n566) );
  NANDN U49035 ( .A(n48666), .B(n48667), .Z(n48665) );
  OR U49036 ( .A(n48668), .B(n48669), .Z(n48667) );
  NAND U49037 ( .A(n48669), .B(n48668), .Z(n48664) );
  XOR U49038 ( .A(n568), .B(n567), .Z(\A1[112] ) );
  XOR U49039 ( .A(n48669), .B(n48670), .Z(n567) );
  XNOR U49040 ( .A(n48668), .B(n48666), .Z(n48670) );
  AND U49041 ( .A(n48671), .B(n48672), .Z(n48666) );
  NANDN U49042 ( .A(n48673), .B(n48674), .Z(n48672) );
  NANDN U49043 ( .A(n48675), .B(n48676), .Z(n48674) );
  NANDN U49044 ( .A(n48676), .B(n48675), .Z(n48671) );
  ANDN U49045 ( .B(B[83]), .A(n54), .Z(n48668) );
  XNOR U49046 ( .A(n48463), .B(n48677), .Z(n48669) );
  XNOR U49047 ( .A(n48462), .B(n48460), .Z(n48677) );
  AND U49048 ( .A(n48678), .B(n48679), .Z(n48460) );
  NANDN U49049 ( .A(n48680), .B(n48681), .Z(n48679) );
  OR U49050 ( .A(n48682), .B(n48683), .Z(n48681) );
  NAND U49051 ( .A(n48683), .B(n48682), .Z(n48678) );
  ANDN U49052 ( .B(B[84]), .A(n55), .Z(n48462) );
  XNOR U49053 ( .A(n48470), .B(n48684), .Z(n48463) );
  XNOR U49054 ( .A(n48469), .B(n48467), .Z(n48684) );
  AND U49055 ( .A(n48685), .B(n48686), .Z(n48467) );
  NANDN U49056 ( .A(n48687), .B(n48688), .Z(n48686) );
  NANDN U49057 ( .A(n48689), .B(n48690), .Z(n48688) );
  NANDN U49058 ( .A(n48690), .B(n48689), .Z(n48685) );
  ANDN U49059 ( .B(B[85]), .A(n56), .Z(n48469) );
  XNOR U49060 ( .A(n48477), .B(n48691), .Z(n48470) );
  XNOR U49061 ( .A(n48476), .B(n48474), .Z(n48691) );
  AND U49062 ( .A(n48692), .B(n48693), .Z(n48474) );
  NANDN U49063 ( .A(n48694), .B(n48695), .Z(n48693) );
  OR U49064 ( .A(n48696), .B(n48697), .Z(n48695) );
  NAND U49065 ( .A(n48697), .B(n48696), .Z(n48692) );
  ANDN U49066 ( .B(B[86]), .A(n57), .Z(n48476) );
  XNOR U49067 ( .A(n48484), .B(n48698), .Z(n48477) );
  XNOR U49068 ( .A(n48483), .B(n48481), .Z(n48698) );
  AND U49069 ( .A(n48699), .B(n48700), .Z(n48481) );
  NANDN U49070 ( .A(n48701), .B(n48702), .Z(n48700) );
  NANDN U49071 ( .A(n48703), .B(n48704), .Z(n48702) );
  NANDN U49072 ( .A(n48704), .B(n48703), .Z(n48699) );
  ANDN U49073 ( .B(B[87]), .A(n58), .Z(n48483) );
  XNOR U49074 ( .A(n48491), .B(n48705), .Z(n48484) );
  XNOR U49075 ( .A(n48490), .B(n48488), .Z(n48705) );
  AND U49076 ( .A(n48706), .B(n48707), .Z(n48488) );
  NANDN U49077 ( .A(n48708), .B(n48709), .Z(n48707) );
  OR U49078 ( .A(n48710), .B(n48711), .Z(n48709) );
  NAND U49079 ( .A(n48711), .B(n48710), .Z(n48706) );
  ANDN U49080 ( .B(B[88]), .A(n59), .Z(n48490) );
  XNOR U49081 ( .A(n48498), .B(n48712), .Z(n48491) );
  XNOR U49082 ( .A(n48497), .B(n48495), .Z(n48712) );
  AND U49083 ( .A(n48713), .B(n48714), .Z(n48495) );
  NANDN U49084 ( .A(n48715), .B(n48716), .Z(n48714) );
  NANDN U49085 ( .A(n48717), .B(n48718), .Z(n48716) );
  NANDN U49086 ( .A(n48718), .B(n48717), .Z(n48713) );
  ANDN U49087 ( .B(B[89]), .A(n60), .Z(n48497) );
  XNOR U49088 ( .A(n48505), .B(n48719), .Z(n48498) );
  XNOR U49089 ( .A(n48504), .B(n48502), .Z(n48719) );
  AND U49090 ( .A(n48720), .B(n48721), .Z(n48502) );
  NANDN U49091 ( .A(n48722), .B(n48723), .Z(n48721) );
  OR U49092 ( .A(n48724), .B(n48725), .Z(n48723) );
  NAND U49093 ( .A(n48725), .B(n48724), .Z(n48720) );
  ANDN U49094 ( .B(B[90]), .A(n61), .Z(n48504) );
  XNOR U49095 ( .A(n48512), .B(n48726), .Z(n48505) );
  XNOR U49096 ( .A(n48511), .B(n48509), .Z(n48726) );
  AND U49097 ( .A(n48727), .B(n48728), .Z(n48509) );
  NANDN U49098 ( .A(n48729), .B(n48730), .Z(n48728) );
  NANDN U49099 ( .A(n48731), .B(n48732), .Z(n48730) );
  NANDN U49100 ( .A(n48732), .B(n48731), .Z(n48727) );
  ANDN U49101 ( .B(A[23]), .A(n21), .Z(n48511) );
  XNOR U49102 ( .A(n48519), .B(n48733), .Z(n48512) );
  XNOR U49103 ( .A(n48518), .B(n48516), .Z(n48733) );
  AND U49104 ( .A(n48734), .B(n48735), .Z(n48516) );
  NANDN U49105 ( .A(n48736), .B(n48737), .Z(n48735) );
  OR U49106 ( .A(n48738), .B(n48739), .Z(n48737) );
  NAND U49107 ( .A(n48739), .B(n48738), .Z(n48734) );
  ANDN U49108 ( .B(A[22]), .A(n19), .Z(n48518) );
  XNOR U49109 ( .A(n48526), .B(n48740), .Z(n48519) );
  XNOR U49110 ( .A(n48525), .B(n48523), .Z(n48740) );
  AND U49111 ( .A(n48741), .B(n48742), .Z(n48523) );
  NANDN U49112 ( .A(n48743), .B(n48744), .Z(n48742) );
  NANDN U49113 ( .A(n48745), .B(n48746), .Z(n48744) );
  NANDN U49114 ( .A(n48746), .B(n48745), .Z(n48741) );
  ANDN U49115 ( .B(A[21]), .A(n17), .Z(n48525) );
  XNOR U49116 ( .A(n48533), .B(n48747), .Z(n48526) );
  XNOR U49117 ( .A(n48532), .B(n48530), .Z(n48747) );
  AND U49118 ( .A(n48748), .B(n48749), .Z(n48530) );
  NANDN U49119 ( .A(n48750), .B(n48751), .Z(n48749) );
  OR U49120 ( .A(n48752), .B(n48753), .Z(n48751) );
  NAND U49121 ( .A(n48753), .B(n48752), .Z(n48748) );
  ANDN U49122 ( .B(A[20]), .A(n15), .Z(n48532) );
  XNOR U49123 ( .A(n48540), .B(n48754), .Z(n48533) );
  XNOR U49124 ( .A(n48539), .B(n48537), .Z(n48754) );
  AND U49125 ( .A(n48755), .B(n48756), .Z(n48537) );
  NANDN U49126 ( .A(n48757), .B(n48758), .Z(n48756) );
  NANDN U49127 ( .A(n48759), .B(n48760), .Z(n48758) );
  NANDN U49128 ( .A(n48760), .B(n48759), .Z(n48755) );
  ANDN U49129 ( .B(A[19]), .A(n13), .Z(n48539) );
  XNOR U49130 ( .A(n48547), .B(n48761), .Z(n48540) );
  XNOR U49131 ( .A(n48546), .B(n48544), .Z(n48761) );
  AND U49132 ( .A(n48762), .B(n48763), .Z(n48544) );
  NANDN U49133 ( .A(n48764), .B(n48765), .Z(n48763) );
  OR U49134 ( .A(n48766), .B(n48767), .Z(n48765) );
  NAND U49135 ( .A(n48767), .B(n48766), .Z(n48762) );
  ANDN U49136 ( .B(A[18]), .A(n11), .Z(n48546) );
  XNOR U49137 ( .A(n48554), .B(n48768), .Z(n48547) );
  XNOR U49138 ( .A(n48553), .B(n48551), .Z(n48768) );
  AND U49139 ( .A(n48769), .B(n48770), .Z(n48551) );
  NANDN U49140 ( .A(n48771), .B(n48772), .Z(n48770) );
  NANDN U49141 ( .A(n48773), .B(n48774), .Z(n48772) );
  NANDN U49142 ( .A(n48774), .B(n48773), .Z(n48769) );
  ANDN U49143 ( .B(A[17]), .A(n9), .Z(n48553) );
  XNOR U49144 ( .A(n48561), .B(n48775), .Z(n48554) );
  XNOR U49145 ( .A(n48560), .B(n48558), .Z(n48775) );
  AND U49146 ( .A(n48776), .B(n48777), .Z(n48558) );
  NANDN U49147 ( .A(n48778), .B(n48779), .Z(n48777) );
  OR U49148 ( .A(n48780), .B(n48781), .Z(n48779) );
  NAND U49149 ( .A(n48781), .B(n48780), .Z(n48776) );
  ANDN U49150 ( .B(B[98]), .A(n69), .Z(n48560) );
  XNOR U49151 ( .A(n48568), .B(n48782), .Z(n48561) );
  XNOR U49152 ( .A(n48567), .B(n48565), .Z(n48782) );
  AND U49153 ( .A(n48783), .B(n48784), .Z(n48565) );
  NANDN U49154 ( .A(n48785), .B(n48786), .Z(n48784) );
  NANDN U49155 ( .A(n48787), .B(n48788), .Z(n48786) );
  NANDN U49156 ( .A(n48788), .B(n48787), .Z(n48783) );
  ANDN U49157 ( .B(A[15]), .A(n6), .Z(n48567) );
  XNOR U49158 ( .A(n48575), .B(n48789), .Z(n48568) );
  XNOR U49159 ( .A(n48574), .B(n48572), .Z(n48789) );
  AND U49160 ( .A(n48790), .B(n48791), .Z(n48572) );
  NANDN U49161 ( .A(n48792), .B(n48793), .Z(n48791) );
  OR U49162 ( .A(n48794), .B(n48795), .Z(n48793) );
  NAND U49163 ( .A(n48795), .B(n48794), .Z(n48790) );
  ANDN U49164 ( .B(A[14]), .A(n4), .Z(n48574) );
  XNOR U49165 ( .A(n48582), .B(n48796), .Z(n48575) );
  XNOR U49166 ( .A(n48581), .B(n48579), .Z(n48796) );
  AND U49167 ( .A(n48797), .B(n48798), .Z(n48579) );
  NANDN U49168 ( .A(n48799), .B(n48800), .Z(n48798) );
  NANDN U49169 ( .A(n48801), .B(n48802), .Z(n48800) );
  NANDN U49170 ( .A(n48802), .B(n48801), .Z(n48797) );
  ANDN U49171 ( .B(B[101]), .A(n72), .Z(n48581) );
  XNOR U49172 ( .A(n48589), .B(n48803), .Z(n48582) );
  XNOR U49173 ( .A(n48588), .B(n48586), .Z(n48803) );
  AND U49174 ( .A(n48804), .B(n48805), .Z(n48586) );
  NANDN U49175 ( .A(n48806), .B(n48807), .Z(n48805) );
  OR U49176 ( .A(n48808), .B(n48809), .Z(n48807) );
  NAND U49177 ( .A(n48809), .B(n48808), .Z(n48804) );
  ANDN U49178 ( .B(B[102]), .A(n73), .Z(n48588) );
  XNOR U49179 ( .A(n48596), .B(n48810), .Z(n48589) );
  XNOR U49180 ( .A(n48595), .B(n48593), .Z(n48810) );
  AND U49181 ( .A(n48811), .B(n48812), .Z(n48593) );
  NANDN U49182 ( .A(n48813), .B(n48814), .Z(n48812) );
  NANDN U49183 ( .A(n48815), .B(n48816), .Z(n48814) );
  NANDN U49184 ( .A(n48816), .B(n48815), .Z(n48811) );
  ANDN U49185 ( .B(B[103]), .A(n74), .Z(n48595) );
  XNOR U49186 ( .A(n48603), .B(n48817), .Z(n48596) );
  XNOR U49187 ( .A(n48602), .B(n48600), .Z(n48817) );
  AND U49188 ( .A(n48818), .B(n48819), .Z(n48600) );
  NANDN U49189 ( .A(n48820), .B(n48821), .Z(n48819) );
  OR U49190 ( .A(n48822), .B(n48823), .Z(n48821) );
  NAND U49191 ( .A(n48823), .B(n48822), .Z(n48818) );
  ANDN U49192 ( .B(B[104]), .A(n75), .Z(n48602) );
  XNOR U49193 ( .A(n48610), .B(n48824), .Z(n48603) );
  XNOR U49194 ( .A(n48609), .B(n48607), .Z(n48824) );
  AND U49195 ( .A(n48825), .B(n48826), .Z(n48607) );
  NANDN U49196 ( .A(n48827), .B(n48828), .Z(n48826) );
  NANDN U49197 ( .A(n48829), .B(n48830), .Z(n48828) );
  NANDN U49198 ( .A(n48830), .B(n48829), .Z(n48825) );
  ANDN U49199 ( .B(B[105]), .A(n76), .Z(n48609) );
  XNOR U49200 ( .A(n48617), .B(n48831), .Z(n48610) );
  XNOR U49201 ( .A(n48616), .B(n48614), .Z(n48831) );
  AND U49202 ( .A(n48832), .B(n48833), .Z(n48614) );
  NANDN U49203 ( .A(n48834), .B(n48835), .Z(n48833) );
  OR U49204 ( .A(n48836), .B(n48837), .Z(n48835) );
  NAND U49205 ( .A(n48837), .B(n48836), .Z(n48832) );
  ANDN U49206 ( .B(B[106]), .A(n77), .Z(n48616) );
  XNOR U49207 ( .A(n48624), .B(n48838), .Z(n48617) );
  XNOR U49208 ( .A(n48623), .B(n48621), .Z(n48838) );
  AND U49209 ( .A(n48839), .B(n48840), .Z(n48621) );
  NANDN U49210 ( .A(n48841), .B(n48842), .Z(n48840) );
  NANDN U49211 ( .A(n48843), .B(n48844), .Z(n48842) );
  NANDN U49212 ( .A(n48844), .B(n48843), .Z(n48839) );
  ANDN U49213 ( .B(B[107]), .A(n78), .Z(n48623) );
  XNOR U49214 ( .A(n48631), .B(n48845), .Z(n48624) );
  XNOR U49215 ( .A(n48630), .B(n48628), .Z(n48845) );
  AND U49216 ( .A(n48846), .B(n48847), .Z(n48628) );
  NANDN U49217 ( .A(n48848), .B(n48849), .Z(n48847) );
  OR U49218 ( .A(n48850), .B(n48851), .Z(n48849) );
  NAND U49219 ( .A(n48851), .B(n48850), .Z(n48846) );
  ANDN U49220 ( .B(B[108]), .A(n79), .Z(n48630) );
  XNOR U49221 ( .A(n48638), .B(n48852), .Z(n48631) );
  XNOR U49222 ( .A(n48637), .B(n48635), .Z(n48852) );
  AND U49223 ( .A(n48853), .B(n48854), .Z(n48635) );
  NANDN U49224 ( .A(n48855), .B(n48856), .Z(n48854) );
  NANDN U49225 ( .A(n48857), .B(n48858), .Z(n48856) );
  NANDN U49226 ( .A(n48858), .B(n48857), .Z(n48853) );
  ANDN U49227 ( .B(B[109]), .A(n80), .Z(n48637) );
  XNOR U49228 ( .A(n48645), .B(n48859), .Z(n48638) );
  XNOR U49229 ( .A(n48644), .B(n48642), .Z(n48859) );
  AND U49230 ( .A(n48860), .B(n48861), .Z(n48642) );
  NANDN U49231 ( .A(n48862), .B(n48863), .Z(n48861) );
  OR U49232 ( .A(n48864), .B(n48865), .Z(n48863) );
  NAND U49233 ( .A(n48865), .B(n48864), .Z(n48860) );
  ANDN U49234 ( .B(B[110]), .A(n81), .Z(n48644) );
  XNOR U49235 ( .A(n48652), .B(n48866), .Z(n48645) );
  XNOR U49236 ( .A(n48651), .B(n48649), .Z(n48866) );
  AND U49237 ( .A(n48867), .B(n48868), .Z(n48649) );
  NANDN U49238 ( .A(n48869), .B(n48870), .Z(n48868) );
  NAND U49239 ( .A(n48871), .B(n48872), .Z(n48870) );
  ANDN U49240 ( .B(B[111]), .A(n82), .Z(n48651) );
  XOR U49241 ( .A(n48658), .B(n48873), .Z(n48652) );
  XNOR U49242 ( .A(n48656), .B(n48659), .Z(n48873) );
  NAND U49243 ( .A(A[2]), .B(B[112]), .Z(n48659) );
  NANDN U49244 ( .A(n48874), .B(n48875), .Z(n48656) );
  AND U49245 ( .A(A[0]), .B(B[113]), .Z(n48875) );
  XNOR U49246 ( .A(n48661), .B(n48876), .Z(n48658) );
  NAND U49247 ( .A(A[0]), .B(B[114]), .Z(n48876) );
  NAND U49248 ( .A(B[113]), .B(A[1]), .Z(n48661) );
  NAND U49249 ( .A(n48877), .B(n48878), .Z(n568) );
  NANDN U49250 ( .A(n48879), .B(n48880), .Z(n48878) );
  OR U49251 ( .A(n48881), .B(n48882), .Z(n48880) );
  NAND U49252 ( .A(n48882), .B(n48881), .Z(n48877) );
  XOR U49253 ( .A(n570), .B(n569), .Z(\A1[111] ) );
  XOR U49254 ( .A(n48882), .B(n48883), .Z(n569) );
  XNOR U49255 ( .A(n48881), .B(n48879), .Z(n48883) );
  AND U49256 ( .A(n48884), .B(n48885), .Z(n48879) );
  NANDN U49257 ( .A(n48886), .B(n48887), .Z(n48885) );
  NANDN U49258 ( .A(n48888), .B(n48889), .Z(n48887) );
  NANDN U49259 ( .A(n48889), .B(n48888), .Z(n48884) );
  ANDN U49260 ( .B(B[82]), .A(n54), .Z(n48881) );
  XNOR U49261 ( .A(n48676), .B(n48890), .Z(n48882) );
  XNOR U49262 ( .A(n48675), .B(n48673), .Z(n48890) );
  AND U49263 ( .A(n48891), .B(n48892), .Z(n48673) );
  NANDN U49264 ( .A(n48893), .B(n48894), .Z(n48892) );
  OR U49265 ( .A(n48895), .B(n48896), .Z(n48894) );
  NAND U49266 ( .A(n48896), .B(n48895), .Z(n48891) );
  ANDN U49267 ( .B(B[83]), .A(n55), .Z(n48675) );
  XNOR U49268 ( .A(n48683), .B(n48897), .Z(n48676) );
  XNOR U49269 ( .A(n48682), .B(n48680), .Z(n48897) );
  AND U49270 ( .A(n48898), .B(n48899), .Z(n48680) );
  NANDN U49271 ( .A(n48900), .B(n48901), .Z(n48899) );
  NANDN U49272 ( .A(n48902), .B(n48903), .Z(n48901) );
  NANDN U49273 ( .A(n48903), .B(n48902), .Z(n48898) );
  ANDN U49274 ( .B(B[84]), .A(n56), .Z(n48682) );
  XNOR U49275 ( .A(n48690), .B(n48904), .Z(n48683) );
  XNOR U49276 ( .A(n48689), .B(n48687), .Z(n48904) );
  AND U49277 ( .A(n48905), .B(n48906), .Z(n48687) );
  NANDN U49278 ( .A(n48907), .B(n48908), .Z(n48906) );
  OR U49279 ( .A(n48909), .B(n48910), .Z(n48908) );
  NAND U49280 ( .A(n48910), .B(n48909), .Z(n48905) );
  ANDN U49281 ( .B(B[85]), .A(n57), .Z(n48689) );
  XNOR U49282 ( .A(n48697), .B(n48911), .Z(n48690) );
  XNOR U49283 ( .A(n48696), .B(n48694), .Z(n48911) );
  AND U49284 ( .A(n48912), .B(n48913), .Z(n48694) );
  NANDN U49285 ( .A(n48914), .B(n48915), .Z(n48913) );
  NANDN U49286 ( .A(n48916), .B(n48917), .Z(n48915) );
  NANDN U49287 ( .A(n48917), .B(n48916), .Z(n48912) );
  ANDN U49288 ( .B(B[86]), .A(n58), .Z(n48696) );
  XNOR U49289 ( .A(n48704), .B(n48918), .Z(n48697) );
  XNOR U49290 ( .A(n48703), .B(n48701), .Z(n48918) );
  AND U49291 ( .A(n48919), .B(n48920), .Z(n48701) );
  NANDN U49292 ( .A(n48921), .B(n48922), .Z(n48920) );
  OR U49293 ( .A(n48923), .B(n48924), .Z(n48922) );
  NAND U49294 ( .A(n48924), .B(n48923), .Z(n48919) );
  ANDN U49295 ( .B(B[87]), .A(n59), .Z(n48703) );
  XNOR U49296 ( .A(n48711), .B(n48925), .Z(n48704) );
  XNOR U49297 ( .A(n48710), .B(n48708), .Z(n48925) );
  AND U49298 ( .A(n48926), .B(n48927), .Z(n48708) );
  NANDN U49299 ( .A(n48928), .B(n48929), .Z(n48927) );
  NANDN U49300 ( .A(n48930), .B(n48931), .Z(n48929) );
  NANDN U49301 ( .A(n48931), .B(n48930), .Z(n48926) );
  ANDN U49302 ( .B(B[88]), .A(n60), .Z(n48710) );
  XNOR U49303 ( .A(n48718), .B(n48932), .Z(n48711) );
  XNOR U49304 ( .A(n48717), .B(n48715), .Z(n48932) );
  AND U49305 ( .A(n48933), .B(n48934), .Z(n48715) );
  NANDN U49306 ( .A(n48935), .B(n48936), .Z(n48934) );
  OR U49307 ( .A(n48937), .B(n48938), .Z(n48936) );
  NAND U49308 ( .A(n48938), .B(n48937), .Z(n48933) );
  ANDN U49309 ( .B(B[89]), .A(n61), .Z(n48717) );
  XNOR U49310 ( .A(n48725), .B(n48939), .Z(n48718) );
  XNOR U49311 ( .A(n48724), .B(n48722), .Z(n48939) );
  AND U49312 ( .A(n48940), .B(n48941), .Z(n48722) );
  NANDN U49313 ( .A(n48942), .B(n48943), .Z(n48941) );
  NANDN U49314 ( .A(n48944), .B(n48945), .Z(n48943) );
  NANDN U49315 ( .A(n48945), .B(n48944), .Z(n48940) );
  ANDN U49316 ( .B(B[90]), .A(n62), .Z(n48724) );
  XNOR U49317 ( .A(n48732), .B(n48946), .Z(n48725) );
  XNOR U49318 ( .A(n48731), .B(n48729), .Z(n48946) );
  AND U49319 ( .A(n48947), .B(n48948), .Z(n48729) );
  NANDN U49320 ( .A(n48949), .B(n48950), .Z(n48948) );
  OR U49321 ( .A(n48951), .B(n48952), .Z(n48950) );
  NAND U49322 ( .A(n48952), .B(n48951), .Z(n48947) );
  ANDN U49323 ( .B(A[22]), .A(n21), .Z(n48731) );
  XNOR U49324 ( .A(n48739), .B(n48953), .Z(n48732) );
  XNOR U49325 ( .A(n48738), .B(n48736), .Z(n48953) );
  AND U49326 ( .A(n48954), .B(n48955), .Z(n48736) );
  NANDN U49327 ( .A(n48956), .B(n48957), .Z(n48955) );
  NANDN U49328 ( .A(n48958), .B(n48959), .Z(n48957) );
  NANDN U49329 ( .A(n48959), .B(n48958), .Z(n48954) );
  ANDN U49330 ( .B(A[21]), .A(n19), .Z(n48738) );
  XNOR U49331 ( .A(n48746), .B(n48960), .Z(n48739) );
  XNOR U49332 ( .A(n48745), .B(n48743), .Z(n48960) );
  AND U49333 ( .A(n48961), .B(n48962), .Z(n48743) );
  NANDN U49334 ( .A(n48963), .B(n48964), .Z(n48962) );
  OR U49335 ( .A(n48965), .B(n48966), .Z(n48964) );
  NAND U49336 ( .A(n48966), .B(n48965), .Z(n48961) );
  ANDN U49337 ( .B(A[20]), .A(n17), .Z(n48745) );
  XNOR U49338 ( .A(n48753), .B(n48967), .Z(n48746) );
  XNOR U49339 ( .A(n48752), .B(n48750), .Z(n48967) );
  AND U49340 ( .A(n48968), .B(n48969), .Z(n48750) );
  NANDN U49341 ( .A(n48970), .B(n48971), .Z(n48969) );
  NANDN U49342 ( .A(n48972), .B(n48973), .Z(n48971) );
  NANDN U49343 ( .A(n48973), .B(n48972), .Z(n48968) );
  ANDN U49344 ( .B(A[19]), .A(n15), .Z(n48752) );
  XNOR U49345 ( .A(n48760), .B(n48974), .Z(n48753) );
  XNOR U49346 ( .A(n48759), .B(n48757), .Z(n48974) );
  AND U49347 ( .A(n48975), .B(n48976), .Z(n48757) );
  NANDN U49348 ( .A(n48977), .B(n48978), .Z(n48976) );
  OR U49349 ( .A(n48979), .B(n48980), .Z(n48978) );
  NAND U49350 ( .A(n48980), .B(n48979), .Z(n48975) );
  ANDN U49351 ( .B(A[18]), .A(n13), .Z(n48759) );
  XNOR U49352 ( .A(n48767), .B(n48981), .Z(n48760) );
  XNOR U49353 ( .A(n48766), .B(n48764), .Z(n48981) );
  AND U49354 ( .A(n48982), .B(n48983), .Z(n48764) );
  NANDN U49355 ( .A(n48984), .B(n48985), .Z(n48983) );
  NANDN U49356 ( .A(n48986), .B(n48987), .Z(n48985) );
  NANDN U49357 ( .A(n48987), .B(n48986), .Z(n48982) );
  ANDN U49358 ( .B(A[17]), .A(n11), .Z(n48766) );
  XNOR U49359 ( .A(n48774), .B(n48988), .Z(n48767) );
  XNOR U49360 ( .A(n48773), .B(n48771), .Z(n48988) );
  AND U49361 ( .A(n48989), .B(n48990), .Z(n48771) );
  NANDN U49362 ( .A(n48991), .B(n48992), .Z(n48990) );
  OR U49363 ( .A(n48993), .B(n48994), .Z(n48992) );
  NAND U49364 ( .A(n48994), .B(n48993), .Z(n48989) );
  ANDN U49365 ( .B(A[16]), .A(n9), .Z(n48773) );
  XNOR U49366 ( .A(n48781), .B(n48995), .Z(n48774) );
  XNOR U49367 ( .A(n48780), .B(n48778), .Z(n48995) );
  AND U49368 ( .A(n48996), .B(n48997), .Z(n48778) );
  NANDN U49369 ( .A(n48998), .B(n48999), .Z(n48997) );
  NANDN U49370 ( .A(n49000), .B(n49001), .Z(n48999) );
  NANDN U49371 ( .A(n49001), .B(n49000), .Z(n48996) );
  ANDN U49372 ( .B(B[98]), .A(n70), .Z(n48780) );
  XNOR U49373 ( .A(n48788), .B(n49002), .Z(n48781) );
  XNOR U49374 ( .A(n48787), .B(n48785), .Z(n49002) );
  AND U49375 ( .A(n49003), .B(n49004), .Z(n48785) );
  NANDN U49376 ( .A(n49005), .B(n49006), .Z(n49004) );
  OR U49377 ( .A(n49007), .B(n49008), .Z(n49006) );
  NAND U49378 ( .A(n49008), .B(n49007), .Z(n49003) );
  ANDN U49379 ( .B(A[14]), .A(n6), .Z(n48787) );
  XNOR U49380 ( .A(n48795), .B(n49009), .Z(n48788) );
  XNOR U49381 ( .A(n48794), .B(n48792), .Z(n49009) );
  AND U49382 ( .A(n49010), .B(n49011), .Z(n48792) );
  NANDN U49383 ( .A(n49012), .B(n49013), .Z(n49011) );
  NANDN U49384 ( .A(n49014), .B(n49015), .Z(n49013) );
  NANDN U49385 ( .A(n49015), .B(n49014), .Z(n49010) );
  ANDN U49386 ( .B(A[13]), .A(n4), .Z(n48794) );
  XNOR U49387 ( .A(n48802), .B(n49016), .Z(n48795) );
  XNOR U49388 ( .A(n48801), .B(n48799), .Z(n49016) );
  AND U49389 ( .A(n49017), .B(n49018), .Z(n48799) );
  NANDN U49390 ( .A(n49019), .B(n49020), .Z(n49018) );
  OR U49391 ( .A(n49021), .B(n49022), .Z(n49020) );
  NAND U49392 ( .A(n49022), .B(n49021), .Z(n49017) );
  ANDN U49393 ( .B(B[101]), .A(n73), .Z(n48801) );
  XNOR U49394 ( .A(n48809), .B(n49023), .Z(n48802) );
  XNOR U49395 ( .A(n48808), .B(n48806), .Z(n49023) );
  AND U49396 ( .A(n49024), .B(n49025), .Z(n48806) );
  NANDN U49397 ( .A(n49026), .B(n49027), .Z(n49025) );
  NANDN U49398 ( .A(n49028), .B(n49029), .Z(n49027) );
  NANDN U49399 ( .A(n49029), .B(n49028), .Z(n49024) );
  ANDN U49400 ( .B(B[102]), .A(n74), .Z(n48808) );
  XNOR U49401 ( .A(n48816), .B(n49030), .Z(n48809) );
  XNOR U49402 ( .A(n48815), .B(n48813), .Z(n49030) );
  AND U49403 ( .A(n49031), .B(n49032), .Z(n48813) );
  NANDN U49404 ( .A(n49033), .B(n49034), .Z(n49032) );
  OR U49405 ( .A(n49035), .B(n49036), .Z(n49034) );
  NAND U49406 ( .A(n49036), .B(n49035), .Z(n49031) );
  ANDN U49407 ( .B(B[103]), .A(n75), .Z(n48815) );
  XNOR U49408 ( .A(n48823), .B(n49037), .Z(n48816) );
  XNOR U49409 ( .A(n48822), .B(n48820), .Z(n49037) );
  AND U49410 ( .A(n49038), .B(n49039), .Z(n48820) );
  NANDN U49411 ( .A(n49040), .B(n49041), .Z(n49039) );
  NANDN U49412 ( .A(n49042), .B(n49043), .Z(n49041) );
  NANDN U49413 ( .A(n49043), .B(n49042), .Z(n49038) );
  ANDN U49414 ( .B(B[104]), .A(n76), .Z(n48822) );
  XNOR U49415 ( .A(n48830), .B(n49044), .Z(n48823) );
  XNOR U49416 ( .A(n48829), .B(n48827), .Z(n49044) );
  AND U49417 ( .A(n49045), .B(n49046), .Z(n48827) );
  NANDN U49418 ( .A(n49047), .B(n49048), .Z(n49046) );
  OR U49419 ( .A(n49049), .B(n49050), .Z(n49048) );
  NAND U49420 ( .A(n49050), .B(n49049), .Z(n49045) );
  ANDN U49421 ( .B(B[105]), .A(n77), .Z(n48829) );
  XNOR U49422 ( .A(n48837), .B(n49051), .Z(n48830) );
  XNOR U49423 ( .A(n48836), .B(n48834), .Z(n49051) );
  AND U49424 ( .A(n49052), .B(n49053), .Z(n48834) );
  NANDN U49425 ( .A(n49054), .B(n49055), .Z(n49053) );
  NANDN U49426 ( .A(n49056), .B(n49057), .Z(n49055) );
  NANDN U49427 ( .A(n49057), .B(n49056), .Z(n49052) );
  ANDN U49428 ( .B(B[106]), .A(n78), .Z(n48836) );
  XNOR U49429 ( .A(n48844), .B(n49058), .Z(n48837) );
  XNOR U49430 ( .A(n48843), .B(n48841), .Z(n49058) );
  AND U49431 ( .A(n49059), .B(n49060), .Z(n48841) );
  NANDN U49432 ( .A(n49061), .B(n49062), .Z(n49060) );
  OR U49433 ( .A(n49063), .B(n49064), .Z(n49062) );
  NAND U49434 ( .A(n49064), .B(n49063), .Z(n49059) );
  ANDN U49435 ( .B(B[107]), .A(n79), .Z(n48843) );
  XNOR U49436 ( .A(n48851), .B(n49065), .Z(n48844) );
  XNOR U49437 ( .A(n48850), .B(n48848), .Z(n49065) );
  AND U49438 ( .A(n49066), .B(n49067), .Z(n48848) );
  NANDN U49439 ( .A(n49068), .B(n49069), .Z(n49067) );
  NANDN U49440 ( .A(n49070), .B(n49071), .Z(n49069) );
  NANDN U49441 ( .A(n49071), .B(n49070), .Z(n49066) );
  ANDN U49442 ( .B(B[108]), .A(n80), .Z(n48850) );
  XNOR U49443 ( .A(n48858), .B(n49072), .Z(n48851) );
  XNOR U49444 ( .A(n48857), .B(n48855), .Z(n49072) );
  AND U49445 ( .A(n49073), .B(n49074), .Z(n48855) );
  NANDN U49446 ( .A(n49075), .B(n49076), .Z(n49074) );
  OR U49447 ( .A(n49077), .B(n49078), .Z(n49076) );
  NAND U49448 ( .A(n49078), .B(n49077), .Z(n49073) );
  ANDN U49449 ( .B(B[109]), .A(n81), .Z(n48857) );
  XNOR U49450 ( .A(n48865), .B(n49079), .Z(n48858) );
  XNOR U49451 ( .A(n48864), .B(n48862), .Z(n49079) );
  AND U49452 ( .A(n49080), .B(n49081), .Z(n48862) );
  NANDN U49453 ( .A(n49082), .B(n49083), .Z(n49081) );
  NAND U49454 ( .A(n49084), .B(n49085), .Z(n49083) );
  ANDN U49455 ( .B(B[110]), .A(n82), .Z(n48864) );
  XOR U49456 ( .A(n48871), .B(n49086), .Z(n48865) );
  XNOR U49457 ( .A(n48869), .B(n48872), .Z(n49086) );
  NAND U49458 ( .A(A[2]), .B(B[111]), .Z(n48872) );
  NANDN U49459 ( .A(n49087), .B(n49088), .Z(n48869) );
  AND U49460 ( .A(A[0]), .B(B[112]), .Z(n49088) );
  XNOR U49461 ( .A(n48874), .B(n49089), .Z(n48871) );
  NAND U49462 ( .A(A[0]), .B(B[113]), .Z(n49089) );
  NAND U49463 ( .A(B[112]), .B(A[1]), .Z(n48874) );
  NAND U49464 ( .A(n49090), .B(n49091), .Z(n570) );
  NANDN U49465 ( .A(n49092), .B(n49093), .Z(n49091) );
  OR U49466 ( .A(n49094), .B(n49095), .Z(n49093) );
  NAND U49467 ( .A(n49095), .B(n49094), .Z(n49090) );
  XOR U49468 ( .A(n572), .B(n571), .Z(\A1[110] ) );
  XOR U49469 ( .A(n49095), .B(n49096), .Z(n571) );
  XNOR U49470 ( .A(n49094), .B(n49092), .Z(n49096) );
  AND U49471 ( .A(n49097), .B(n49098), .Z(n49092) );
  NANDN U49472 ( .A(n49099), .B(n49100), .Z(n49098) );
  NANDN U49473 ( .A(n49101), .B(n49102), .Z(n49100) );
  NANDN U49474 ( .A(n49102), .B(n49101), .Z(n49097) );
  ANDN U49475 ( .B(B[81]), .A(n54), .Z(n49094) );
  XNOR U49476 ( .A(n48889), .B(n49103), .Z(n49095) );
  XNOR U49477 ( .A(n48888), .B(n48886), .Z(n49103) );
  AND U49478 ( .A(n49104), .B(n49105), .Z(n48886) );
  NANDN U49479 ( .A(n49106), .B(n49107), .Z(n49105) );
  OR U49480 ( .A(n49108), .B(n49109), .Z(n49107) );
  NAND U49481 ( .A(n49109), .B(n49108), .Z(n49104) );
  ANDN U49482 ( .B(B[82]), .A(n55), .Z(n48888) );
  XNOR U49483 ( .A(n48896), .B(n49110), .Z(n48889) );
  XNOR U49484 ( .A(n48895), .B(n48893), .Z(n49110) );
  AND U49485 ( .A(n49111), .B(n49112), .Z(n48893) );
  NANDN U49486 ( .A(n49113), .B(n49114), .Z(n49112) );
  NANDN U49487 ( .A(n49115), .B(n49116), .Z(n49114) );
  NANDN U49488 ( .A(n49116), .B(n49115), .Z(n49111) );
  ANDN U49489 ( .B(B[83]), .A(n56), .Z(n48895) );
  XNOR U49490 ( .A(n48903), .B(n49117), .Z(n48896) );
  XNOR U49491 ( .A(n48902), .B(n48900), .Z(n49117) );
  AND U49492 ( .A(n49118), .B(n49119), .Z(n48900) );
  NANDN U49493 ( .A(n49120), .B(n49121), .Z(n49119) );
  OR U49494 ( .A(n49122), .B(n49123), .Z(n49121) );
  NAND U49495 ( .A(n49123), .B(n49122), .Z(n49118) );
  ANDN U49496 ( .B(B[84]), .A(n57), .Z(n48902) );
  XNOR U49497 ( .A(n48910), .B(n49124), .Z(n48903) );
  XNOR U49498 ( .A(n48909), .B(n48907), .Z(n49124) );
  AND U49499 ( .A(n49125), .B(n49126), .Z(n48907) );
  NANDN U49500 ( .A(n49127), .B(n49128), .Z(n49126) );
  NANDN U49501 ( .A(n49129), .B(n49130), .Z(n49128) );
  NANDN U49502 ( .A(n49130), .B(n49129), .Z(n49125) );
  ANDN U49503 ( .B(B[85]), .A(n58), .Z(n48909) );
  XNOR U49504 ( .A(n48917), .B(n49131), .Z(n48910) );
  XNOR U49505 ( .A(n48916), .B(n48914), .Z(n49131) );
  AND U49506 ( .A(n49132), .B(n49133), .Z(n48914) );
  NANDN U49507 ( .A(n49134), .B(n49135), .Z(n49133) );
  OR U49508 ( .A(n49136), .B(n49137), .Z(n49135) );
  NAND U49509 ( .A(n49137), .B(n49136), .Z(n49132) );
  ANDN U49510 ( .B(B[86]), .A(n59), .Z(n48916) );
  XNOR U49511 ( .A(n48924), .B(n49138), .Z(n48917) );
  XNOR U49512 ( .A(n48923), .B(n48921), .Z(n49138) );
  AND U49513 ( .A(n49139), .B(n49140), .Z(n48921) );
  NANDN U49514 ( .A(n49141), .B(n49142), .Z(n49140) );
  NANDN U49515 ( .A(n49143), .B(n49144), .Z(n49142) );
  NANDN U49516 ( .A(n49144), .B(n49143), .Z(n49139) );
  ANDN U49517 ( .B(B[87]), .A(n60), .Z(n48923) );
  XNOR U49518 ( .A(n48931), .B(n49145), .Z(n48924) );
  XNOR U49519 ( .A(n48930), .B(n48928), .Z(n49145) );
  AND U49520 ( .A(n49146), .B(n49147), .Z(n48928) );
  NANDN U49521 ( .A(n49148), .B(n49149), .Z(n49147) );
  OR U49522 ( .A(n49150), .B(n49151), .Z(n49149) );
  NAND U49523 ( .A(n49151), .B(n49150), .Z(n49146) );
  ANDN U49524 ( .B(B[88]), .A(n61), .Z(n48930) );
  XNOR U49525 ( .A(n48938), .B(n49152), .Z(n48931) );
  XNOR U49526 ( .A(n48937), .B(n48935), .Z(n49152) );
  AND U49527 ( .A(n49153), .B(n49154), .Z(n48935) );
  NANDN U49528 ( .A(n49155), .B(n49156), .Z(n49154) );
  NANDN U49529 ( .A(n49157), .B(n49158), .Z(n49156) );
  NANDN U49530 ( .A(n49158), .B(n49157), .Z(n49153) );
  ANDN U49531 ( .B(B[89]), .A(n62), .Z(n48937) );
  XNOR U49532 ( .A(n48945), .B(n49159), .Z(n48938) );
  XNOR U49533 ( .A(n48944), .B(n48942), .Z(n49159) );
  AND U49534 ( .A(n49160), .B(n49161), .Z(n48942) );
  NANDN U49535 ( .A(n49162), .B(n49163), .Z(n49161) );
  OR U49536 ( .A(n49164), .B(n49165), .Z(n49163) );
  NAND U49537 ( .A(n49165), .B(n49164), .Z(n49160) );
  ANDN U49538 ( .B(A[22]), .A(n23), .Z(n48944) );
  XNOR U49539 ( .A(n48952), .B(n49166), .Z(n48945) );
  XNOR U49540 ( .A(n48951), .B(n48949), .Z(n49166) );
  AND U49541 ( .A(n49167), .B(n49168), .Z(n48949) );
  NANDN U49542 ( .A(n49169), .B(n49170), .Z(n49168) );
  NANDN U49543 ( .A(n49171), .B(n49172), .Z(n49170) );
  NANDN U49544 ( .A(n49172), .B(n49171), .Z(n49167) );
  ANDN U49545 ( .B(A[21]), .A(n21), .Z(n48951) );
  XNOR U49546 ( .A(n48959), .B(n49173), .Z(n48952) );
  XNOR U49547 ( .A(n48958), .B(n48956), .Z(n49173) );
  AND U49548 ( .A(n49174), .B(n49175), .Z(n48956) );
  NANDN U49549 ( .A(n49176), .B(n49177), .Z(n49175) );
  OR U49550 ( .A(n49178), .B(n49179), .Z(n49177) );
  NAND U49551 ( .A(n49179), .B(n49178), .Z(n49174) );
  ANDN U49552 ( .B(A[20]), .A(n19), .Z(n48958) );
  XNOR U49553 ( .A(n48966), .B(n49180), .Z(n48959) );
  XNOR U49554 ( .A(n48965), .B(n48963), .Z(n49180) );
  AND U49555 ( .A(n49181), .B(n49182), .Z(n48963) );
  NANDN U49556 ( .A(n49183), .B(n49184), .Z(n49182) );
  NANDN U49557 ( .A(n49185), .B(n49186), .Z(n49184) );
  NANDN U49558 ( .A(n49186), .B(n49185), .Z(n49181) );
  ANDN U49559 ( .B(A[19]), .A(n17), .Z(n48965) );
  XNOR U49560 ( .A(n48973), .B(n49187), .Z(n48966) );
  XNOR U49561 ( .A(n48972), .B(n48970), .Z(n49187) );
  AND U49562 ( .A(n49188), .B(n49189), .Z(n48970) );
  NANDN U49563 ( .A(n49190), .B(n49191), .Z(n49189) );
  OR U49564 ( .A(n49192), .B(n49193), .Z(n49191) );
  NAND U49565 ( .A(n49193), .B(n49192), .Z(n49188) );
  ANDN U49566 ( .B(A[18]), .A(n15), .Z(n48972) );
  XNOR U49567 ( .A(n48980), .B(n49194), .Z(n48973) );
  XNOR U49568 ( .A(n48979), .B(n48977), .Z(n49194) );
  AND U49569 ( .A(n49195), .B(n49196), .Z(n48977) );
  NANDN U49570 ( .A(n49197), .B(n49198), .Z(n49196) );
  NANDN U49571 ( .A(n49199), .B(n49200), .Z(n49198) );
  NANDN U49572 ( .A(n49200), .B(n49199), .Z(n49195) );
  ANDN U49573 ( .B(A[17]), .A(n13), .Z(n48979) );
  XNOR U49574 ( .A(n48987), .B(n49201), .Z(n48980) );
  XNOR U49575 ( .A(n48986), .B(n48984), .Z(n49201) );
  AND U49576 ( .A(n49202), .B(n49203), .Z(n48984) );
  NANDN U49577 ( .A(n49204), .B(n49205), .Z(n49203) );
  OR U49578 ( .A(n49206), .B(n49207), .Z(n49205) );
  NAND U49579 ( .A(n49207), .B(n49206), .Z(n49202) );
  ANDN U49580 ( .B(A[16]), .A(n11), .Z(n48986) );
  XNOR U49581 ( .A(n48994), .B(n49208), .Z(n48987) );
  XNOR U49582 ( .A(n48993), .B(n48991), .Z(n49208) );
  AND U49583 ( .A(n49209), .B(n49210), .Z(n48991) );
  NANDN U49584 ( .A(n49211), .B(n49212), .Z(n49210) );
  NANDN U49585 ( .A(n49213), .B(n49214), .Z(n49212) );
  NANDN U49586 ( .A(n49214), .B(n49213), .Z(n49209) );
  ANDN U49587 ( .B(A[15]), .A(n9), .Z(n48993) );
  XNOR U49588 ( .A(n49001), .B(n49215), .Z(n48994) );
  XNOR U49589 ( .A(n49000), .B(n48998), .Z(n49215) );
  AND U49590 ( .A(n49216), .B(n49217), .Z(n48998) );
  NANDN U49591 ( .A(n49218), .B(n49219), .Z(n49217) );
  OR U49592 ( .A(n49220), .B(n49221), .Z(n49219) );
  NAND U49593 ( .A(n49221), .B(n49220), .Z(n49216) );
  ANDN U49594 ( .B(B[98]), .A(n71), .Z(n49000) );
  XNOR U49595 ( .A(n49008), .B(n49222), .Z(n49001) );
  XNOR U49596 ( .A(n49007), .B(n49005), .Z(n49222) );
  AND U49597 ( .A(n49223), .B(n49224), .Z(n49005) );
  NANDN U49598 ( .A(n49225), .B(n49226), .Z(n49224) );
  NANDN U49599 ( .A(n49227), .B(n49228), .Z(n49226) );
  NANDN U49600 ( .A(n49228), .B(n49227), .Z(n49223) );
  ANDN U49601 ( .B(A[13]), .A(n6), .Z(n49007) );
  XNOR U49602 ( .A(n49015), .B(n49229), .Z(n49008) );
  XNOR U49603 ( .A(n49014), .B(n49012), .Z(n49229) );
  AND U49604 ( .A(n49230), .B(n49231), .Z(n49012) );
  NANDN U49605 ( .A(n49232), .B(n49233), .Z(n49231) );
  OR U49606 ( .A(n49234), .B(n49235), .Z(n49233) );
  NAND U49607 ( .A(n49235), .B(n49234), .Z(n49230) );
  ANDN U49608 ( .B(A[12]), .A(n4), .Z(n49014) );
  XNOR U49609 ( .A(n49022), .B(n49236), .Z(n49015) );
  XNOR U49610 ( .A(n49021), .B(n49019), .Z(n49236) );
  AND U49611 ( .A(n49237), .B(n49238), .Z(n49019) );
  NANDN U49612 ( .A(n49239), .B(n49240), .Z(n49238) );
  NANDN U49613 ( .A(n49241), .B(n49242), .Z(n49240) );
  NANDN U49614 ( .A(n49242), .B(n49241), .Z(n49237) );
  ANDN U49615 ( .B(B[101]), .A(n74), .Z(n49021) );
  XNOR U49616 ( .A(n49029), .B(n49243), .Z(n49022) );
  XNOR U49617 ( .A(n49028), .B(n49026), .Z(n49243) );
  AND U49618 ( .A(n49244), .B(n49245), .Z(n49026) );
  NANDN U49619 ( .A(n49246), .B(n49247), .Z(n49245) );
  OR U49620 ( .A(n49248), .B(n49249), .Z(n49247) );
  NAND U49621 ( .A(n49249), .B(n49248), .Z(n49244) );
  ANDN U49622 ( .B(B[102]), .A(n75), .Z(n49028) );
  XNOR U49623 ( .A(n49036), .B(n49250), .Z(n49029) );
  XNOR U49624 ( .A(n49035), .B(n49033), .Z(n49250) );
  AND U49625 ( .A(n49251), .B(n49252), .Z(n49033) );
  NANDN U49626 ( .A(n49253), .B(n49254), .Z(n49252) );
  NANDN U49627 ( .A(n49255), .B(n49256), .Z(n49254) );
  NANDN U49628 ( .A(n49256), .B(n49255), .Z(n49251) );
  ANDN U49629 ( .B(B[103]), .A(n76), .Z(n49035) );
  XNOR U49630 ( .A(n49043), .B(n49257), .Z(n49036) );
  XNOR U49631 ( .A(n49042), .B(n49040), .Z(n49257) );
  AND U49632 ( .A(n49258), .B(n49259), .Z(n49040) );
  NANDN U49633 ( .A(n49260), .B(n49261), .Z(n49259) );
  OR U49634 ( .A(n49262), .B(n49263), .Z(n49261) );
  NAND U49635 ( .A(n49263), .B(n49262), .Z(n49258) );
  ANDN U49636 ( .B(B[104]), .A(n77), .Z(n49042) );
  XNOR U49637 ( .A(n49050), .B(n49264), .Z(n49043) );
  XNOR U49638 ( .A(n49049), .B(n49047), .Z(n49264) );
  AND U49639 ( .A(n49265), .B(n49266), .Z(n49047) );
  NANDN U49640 ( .A(n49267), .B(n49268), .Z(n49266) );
  NANDN U49641 ( .A(n49269), .B(n49270), .Z(n49268) );
  NANDN U49642 ( .A(n49270), .B(n49269), .Z(n49265) );
  ANDN U49643 ( .B(B[105]), .A(n78), .Z(n49049) );
  XNOR U49644 ( .A(n49057), .B(n49271), .Z(n49050) );
  XNOR U49645 ( .A(n49056), .B(n49054), .Z(n49271) );
  AND U49646 ( .A(n49272), .B(n49273), .Z(n49054) );
  NANDN U49647 ( .A(n49274), .B(n49275), .Z(n49273) );
  OR U49648 ( .A(n49276), .B(n49277), .Z(n49275) );
  NAND U49649 ( .A(n49277), .B(n49276), .Z(n49272) );
  ANDN U49650 ( .B(B[106]), .A(n79), .Z(n49056) );
  XNOR U49651 ( .A(n49064), .B(n49278), .Z(n49057) );
  XNOR U49652 ( .A(n49063), .B(n49061), .Z(n49278) );
  AND U49653 ( .A(n49279), .B(n49280), .Z(n49061) );
  NANDN U49654 ( .A(n49281), .B(n49282), .Z(n49280) );
  NANDN U49655 ( .A(n49283), .B(n49284), .Z(n49282) );
  NANDN U49656 ( .A(n49284), .B(n49283), .Z(n49279) );
  ANDN U49657 ( .B(B[107]), .A(n80), .Z(n49063) );
  XNOR U49658 ( .A(n49071), .B(n49285), .Z(n49064) );
  XNOR U49659 ( .A(n49070), .B(n49068), .Z(n49285) );
  AND U49660 ( .A(n49286), .B(n49287), .Z(n49068) );
  NANDN U49661 ( .A(n49288), .B(n49289), .Z(n49287) );
  OR U49662 ( .A(n49290), .B(n49291), .Z(n49289) );
  NAND U49663 ( .A(n49291), .B(n49290), .Z(n49286) );
  ANDN U49664 ( .B(B[108]), .A(n81), .Z(n49070) );
  XNOR U49665 ( .A(n49078), .B(n49292), .Z(n49071) );
  XNOR U49666 ( .A(n49077), .B(n49075), .Z(n49292) );
  AND U49667 ( .A(n49293), .B(n49294), .Z(n49075) );
  NANDN U49668 ( .A(n49295), .B(n49296), .Z(n49294) );
  NAND U49669 ( .A(n49297), .B(n49298), .Z(n49296) );
  ANDN U49670 ( .B(B[109]), .A(n82), .Z(n49077) );
  XOR U49671 ( .A(n49084), .B(n49299), .Z(n49078) );
  XNOR U49672 ( .A(n49082), .B(n49085), .Z(n49299) );
  NAND U49673 ( .A(A[2]), .B(B[110]), .Z(n49085) );
  NANDN U49674 ( .A(n49300), .B(n49301), .Z(n49082) );
  AND U49675 ( .A(A[0]), .B(B[111]), .Z(n49301) );
  XNOR U49676 ( .A(n49087), .B(n49302), .Z(n49084) );
  NAND U49677 ( .A(A[0]), .B(B[112]), .Z(n49302) );
  NAND U49678 ( .A(B[111]), .B(A[1]), .Z(n49087) );
  NAND U49679 ( .A(n49303), .B(n49304), .Z(n572) );
  NANDN U49680 ( .A(n49305), .B(n49306), .Z(n49304) );
  OR U49681 ( .A(n49307), .B(n49308), .Z(n49306) );
  NAND U49682 ( .A(n49308), .B(n49307), .Z(n49303) );
  XNOR U49683 ( .A(n47103), .B(n49309), .Z(\A1[10] ) );
  XNOR U49684 ( .A(n47101), .B(n47104), .Z(n49309) );
  AND U49685 ( .A(n49310), .B(n49311), .Z(n47104) );
  NANDN U49686 ( .A(n597), .B(n49312), .Z(n49311) );
  NANDN U49687 ( .A(n595), .B(n49313), .Z(n49312) );
  NAND U49688 ( .A(A[11]), .B(B[0]), .Z(n597) );
  NAND U49689 ( .A(n49), .B(n595), .Z(n49310) );
  XOR U49690 ( .A(n49314), .B(n49315), .Z(n595) );
  XNOR U49691 ( .A(n49316), .B(n49317), .Z(n49315) );
  AND U49692 ( .A(n49318), .B(n49319), .Z(n49313) );
  NANDN U49693 ( .A(n1006), .B(n49320), .Z(n49319) );
  NANDN U49694 ( .A(n1004), .B(n1007), .Z(n49320) );
  NAND U49695 ( .A(A[10]), .B(B[0]), .Z(n1006) );
  NANDN U49696 ( .A(n1007), .B(n1004), .Z(n49318) );
  XOR U49697 ( .A(n49321), .B(n49322), .Z(n1004) );
  XNOR U49698 ( .A(n49323), .B(n49324), .Z(n49322) );
  AND U49699 ( .A(n49325), .B(n49326), .Z(n1007) );
  NANDN U49700 ( .A(n2115), .B(n49327), .Z(n49326) );
  NANDN U49701 ( .A(n2113), .B(n49328), .Z(n49327) );
  NAND U49702 ( .A(A[9]), .B(B[0]), .Z(n2115) );
  NAND U49703 ( .A(n50), .B(n2113), .Z(n49325) );
  XOR U49704 ( .A(n49329), .B(n49330), .Z(n2113) );
  XNOR U49705 ( .A(n49331), .B(n49332), .Z(n49330) );
  AND U49706 ( .A(n49333), .B(n49334), .Z(n49328) );
  NANDN U49707 ( .A(n3924), .B(n49335), .Z(n49334) );
  NANDN U49708 ( .A(n3922), .B(n3925), .Z(n49335) );
  NAND U49709 ( .A(A[8]), .B(B[0]), .Z(n3924) );
  NANDN U49710 ( .A(n3925), .B(n3922), .Z(n49333) );
  XOR U49711 ( .A(n49336), .B(n49337), .Z(n3922) );
  XNOR U49712 ( .A(n49338), .B(n49339), .Z(n49337) );
  AND U49713 ( .A(n49340), .B(n49341), .Z(n3925) );
  NANDN U49714 ( .A(n6059), .B(n49342), .Z(n49341) );
  NANDN U49715 ( .A(n6057), .B(n49343), .Z(n49342) );
  NAND U49716 ( .A(A[7]), .B(B[0]), .Z(n6059) );
  NAND U49717 ( .A(n51), .B(n6057), .Z(n49340) );
  XOR U49718 ( .A(n49344), .B(n49345), .Z(n6057) );
  XNOR U49719 ( .A(n49346), .B(n49347), .Z(n49345) );
  AND U49720 ( .A(n49348), .B(n49349), .Z(n49343) );
  NANDN U49721 ( .A(n8192), .B(n49350), .Z(n49349) );
  NANDN U49722 ( .A(n8190), .B(n8193), .Z(n49350) );
  NAND U49723 ( .A(A[6]), .B(B[0]), .Z(n8192) );
  NANDN U49724 ( .A(n8193), .B(n8190), .Z(n49348) );
  XOR U49725 ( .A(n49351), .B(n49352), .Z(n8190) );
  XNOR U49726 ( .A(n49353), .B(n49354), .Z(n49352) );
  AND U49727 ( .A(n49355), .B(n49356), .Z(n8193) );
  NANDN U49728 ( .A(n10326), .B(n49357), .Z(n49356) );
  NANDN U49729 ( .A(n10324), .B(n49358), .Z(n49357) );
  NAND U49730 ( .A(A[5]), .B(B[0]), .Z(n10326) );
  NAND U49731 ( .A(n52), .B(n10324), .Z(n49355) );
  XOR U49732 ( .A(n49359), .B(n49360), .Z(n10324) );
  XNOR U49733 ( .A(n49361), .B(n49362), .Z(n49360) );
  AND U49734 ( .A(n49363), .B(n49364), .Z(n49358) );
  NANDN U49735 ( .A(n12459), .B(n49365), .Z(n49364) );
  NANDN U49736 ( .A(n12457), .B(n12460), .Z(n49365) );
  NAND U49737 ( .A(A[4]), .B(B[0]), .Z(n12459) );
  NANDN U49738 ( .A(n12460), .B(n12457), .Z(n49363) );
  XOR U49739 ( .A(n49366), .B(n49367), .Z(n12457) );
  XNOR U49740 ( .A(n49368), .B(n49369), .Z(n49367) );
  AND U49741 ( .A(n49370), .B(n49371), .Z(n12460) );
  NANDN U49742 ( .A(n29157), .B(n49372), .Z(n49371) );
  OR U49743 ( .A(n29156), .B(n29154), .Z(n49372) );
  AND U49744 ( .A(n49373), .B(n49374), .Z(n29157) );
  NANDN U49745 ( .A(n49375), .B(n49376), .Z(n49374) );
  OR U49746 ( .A(n49377), .B(n53), .Z(n49376) );
  NAND U49747 ( .A(n53), .B(n49377), .Z(n49373) );
  NAND U49748 ( .A(n29154), .B(n29156), .Z(n49370) );
  ANDN U49749 ( .B(B[0]), .A(n82), .Z(n29156) );
  XOR U49750 ( .A(n49379), .B(n49380), .Z(n29154) );
  XNOR U49751 ( .A(n49381), .B(n49382), .Z(n49380) );
  NAND U49752 ( .A(A[12]), .B(B[0]), .Z(n47101) );
  XOR U49753 ( .A(n47111), .B(n49383), .Z(n47103) );
  XNOR U49754 ( .A(n47110), .B(n47108), .Z(n49383) );
  AND U49755 ( .A(n49384), .B(n49385), .Z(n47108) );
  NANDN U49756 ( .A(n49317), .B(n49386), .Z(n49385) );
  AND U49757 ( .A(n49387), .B(n49388), .Z(n49317) );
  NANDN U49758 ( .A(n49324), .B(n49389), .Z(n49388) );
  OR U49759 ( .A(n49323), .B(n49321), .Z(n49389) );
  AND U49760 ( .A(n49390), .B(n49391), .Z(n49324) );
  NANDN U49761 ( .A(n49332), .B(n49392), .Z(n49391) );
  AND U49762 ( .A(n49393), .B(n49394), .Z(n49332) );
  NANDN U49763 ( .A(n49339), .B(n49395), .Z(n49394) );
  OR U49764 ( .A(n49338), .B(n49336), .Z(n49395) );
  AND U49765 ( .A(n49396), .B(n49397), .Z(n49339) );
  NANDN U49766 ( .A(n49347), .B(n49398), .Z(n49397) );
  AND U49767 ( .A(n49399), .B(n49400), .Z(n49347) );
  NANDN U49768 ( .A(n49354), .B(n49401), .Z(n49400) );
  OR U49769 ( .A(n49353), .B(n49351), .Z(n49401) );
  AND U49770 ( .A(n49402), .B(n49403), .Z(n49354) );
  NANDN U49771 ( .A(n49362), .B(n49404), .Z(n49403) );
  AND U49772 ( .A(n49405), .B(n49406), .Z(n49362) );
  NANDN U49773 ( .A(n49369), .B(n49407), .Z(n49406) );
  OR U49774 ( .A(n49368), .B(n49366), .Z(n49407) );
  AND U49775 ( .A(n49408), .B(n49409), .Z(n49369) );
  NANDN U49776 ( .A(n49381), .B(n49410), .Z(n49409) );
  NAND U49777 ( .A(n49379), .B(n49382), .Z(n49410) );
  NANDN U49778 ( .A(n49411), .B(n49412), .Z(n49381) );
  AND U49779 ( .A(A[0]), .B(B[2]), .Z(n49412) );
  XNOR U49780 ( .A(n49413), .B(n49414), .Z(n49379) );
  NAND U49781 ( .A(A[0]), .B(B[3]), .Z(n49414) );
  NAND U49782 ( .A(B[1]), .B(A[2]), .Z(n49382) );
  NAND U49783 ( .A(n49366), .B(n49368), .Z(n49405) );
  ANDN U49784 ( .B(B[1]), .A(n82), .Z(n49368) );
  XOR U49785 ( .A(n49415), .B(n49416), .Z(n49366) );
  XNOR U49786 ( .A(n49417), .B(n49418), .Z(n49416) );
  NAND U49787 ( .A(n49359), .B(n49361), .Z(n49402) );
  ANDN U49788 ( .B(B[1]), .A(n81), .Z(n49361) );
  XOR U49789 ( .A(n49419), .B(n49420), .Z(n49359) );
  XNOR U49790 ( .A(n49421), .B(n49422), .Z(n49420) );
  NAND U49791 ( .A(n49351), .B(n49353), .Z(n49399) );
  ANDN U49792 ( .B(B[1]), .A(n80), .Z(n49353) );
  XNOR U49793 ( .A(n49423), .B(n49424), .Z(n49351) );
  XNOR U49794 ( .A(n49425), .B(n49426), .Z(n49424) );
  NAND U49795 ( .A(n49344), .B(n49346), .Z(n49396) );
  ANDN U49796 ( .B(B[1]), .A(n79), .Z(n49346) );
  XOR U49797 ( .A(n49427), .B(n49428), .Z(n49344) );
  XNOR U49798 ( .A(n49429), .B(n49430), .Z(n49428) );
  NAND U49799 ( .A(n49336), .B(n49338), .Z(n49393) );
  ANDN U49800 ( .B(B[1]), .A(n78), .Z(n49338) );
  XNOR U49801 ( .A(n49431), .B(n49432), .Z(n49336) );
  XNOR U49802 ( .A(n49433), .B(n49434), .Z(n49432) );
  NAND U49803 ( .A(n49329), .B(n49331), .Z(n49390) );
  ANDN U49804 ( .B(B[1]), .A(n77), .Z(n49331) );
  XOR U49805 ( .A(n49435), .B(n49436), .Z(n49329) );
  XNOR U49806 ( .A(n49437), .B(n49438), .Z(n49436) );
  NAND U49807 ( .A(n49321), .B(n49323), .Z(n49387) );
  ANDN U49808 ( .B(B[1]), .A(n76), .Z(n49323) );
  XNOR U49809 ( .A(n49439), .B(n49440), .Z(n49321) );
  XNOR U49810 ( .A(n49441), .B(n49442), .Z(n49440) );
  NAND U49811 ( .A(n49314), .B(n49316), .Z(n49384) );
  ANDN U49812 ( .B(B[1]), .A(n75), .Z(n49316) );
  XOR U49813 ( .A(n49443), .B(n49444), .Z(n49314) );
  XNOR U49814 ( .A(n49445), .B(n49446), .Z(n49444) );
  ANDN U49815 ( .B(B[1]), .A(n74), .Z(n47110) );
  XNOR U49816 ( .A(n47118), .B(n49447), .Z(n47111) );
  XNOR U49817 ( .A(n47117), .B(n47115), .Z(n49447) );
  AND U49818 ( .A(n49448), .B(n49449), .Z(n47115) );
  NANDN U49819 ( .A(n49446), .B(n49450), .Z(n49449) );
  OR U49820 ( .A(n49445), .B(n49443), .Z(n49450) );
  AND U49821 ( .A(n49451), .B(n49452), .Z(n49446) );
  NANDN U49822 ( .A(n49442), .B(n49453), .Z(n49452) );
  NANDN U49823 ( .A(n49441), .B(n49439), .Z(n49453) );
  AND U49824 ( .A(n49454), .B(n49455), .Z(n49442) );
  NANDN U49825 ( .A(n49438), .B(n49456), .Z(n49455) );
  OR U49826 ( .A(n49437), .B(n49435), .Z(n49456) );
  AND U49827 ( .A(n49457), .B(n49458), .Z(n49438) );
  NANDN U49828 ( .A(n49434), .B(n49459), .Z(n49458) );
  NANDN U49829 ( .A(n49433), .B(n49431), .Z(n49459) );
  AND U49830 ( .A(n49460), .B(n49461), .Z(n49434) );
  NANDN U49831 ( .A(n49430), .B(n49462), .Z(n49461) );
  OR U49832 ( .A(n49429), .B(n49427), .Z(n49462) );
  AND U49833 ( .A(n49463), .B(n49464), .Z(n49430) );
  NANDN U49834 ( .A(n49426), .B(n49465), .Z(n49464) );
  NANDN U49835 ( .A(n49425), .B(n49423), .Z(n49465) );
  AND U49836 ( .A(n49466), .B(n49467), .Z(n49426) );
  NANDN U49837 ( .A(n49422), .B(n49468), .Z(n49467) );
  OR U49838 ( .A(n49421), .B(n49419), .Z(n49468) );
  AND U49839 ( .A(n49469), .B(n49470), .Z(n49422) );
  NANDN U49840 ( .A(n49417), .B(n49471), .Z(n49470) );
  NAND U49841 ( .A(n49415), .B(n49418), .Z(n49471) );
  NANDN U49842 ( .A(n49413), .B(n49472), .Z(n49417) );
  AND U49843 ( .A(A[0]), .B(B[3]), .Z(n49472) );
  NAND U49844 ( .A(B[2]), .B(A[1]), .Z(n49413) );
  XNOR U49845 ( .A(n49473), .B(n49474), .Z(n49415) );
  NAND U49846 ( .A(A[0]), .B(B[4]), .Z(n49474) );
  NAND U49847 ( .A(A[2]), .B(B[2]), .Z(n49418) );
  NAND U49848 ( .A(n49419), .B(n49421), .Z(n49466) );
  ANDN U49849 ( .B(B[2]), .A(n82), .Z(n49421) );
  XOR U49850 ( .A(n49475), .B(n49476), .Z(n49419) );
  XNOR U49851 ( .A(n49477), .B(n49478), .Z(n49476) );
  NANDN U49852 ( .A(n49423), .B(n49425), .Z(n49463) );
  ANDN U49853 ( .B(B[2]), .A(n81), .Z(n49425) );
  XNOR U49854 ( .A(n49479), .B(n49480), .Z(n49423) );
  XNOR U49855 ( .A(n49481), .B(n49482), .Z(n49480) );
  NAND U49856 ( .A(n49427), .B(n49429), .Z(n49460) );
  ANDN U49857 ( .B(B[2]), .A(n80), .Z(n49429) );
  XNOR U49858 ( .A(n49483), .B(n49484), .Z(n49427) );
  XNOR U49859 ( .A(n49485), .B(n49486), .Z(n49484) );
  NANDN U49860 ( .A(n49431), .B(n49433), .Z(n49457) );
  ANDN U49861 ( .B(B[2]), .A(n79), .Z(n49433) );
  XNOR U49862 ( .A(n49487), .B(n49488), .Z(n49431) );
  XNOR U49863 ( .A(n49489), .B(n49490), .Z(n49488) );
  NAND U49864 ( .A(n49435), .B(n49437), .Z(n49454) );
  ANDN U49865 ( .B(B[2]), .A(n78), .Z(n49437) );
  XNOR U49866 ( .A(n49491), .B(n49492), .Z(n49435) );
  XNOR U49867 ( .A(n49493), .B(n49494), .Z(n49492) );
  NANDN U49868 ( .A(n49439), .B(n49441), .Z(n49451) );
  ANDN U49869 ( .B(B[2]), .A(n77), .Z(n49441) );
  XNOR U49870 ( .A(n49495), .B(n49496), .Z(n49439) );
  XNOR U49871 ( .A(n49497), .B(n49498), .Z(n49496) );
  NAND U49872 ( .A(n49443), .B(n49445), .Z(n49448) );
  ANDN U49873 ( .B(B[2]), .A(n76), .Z(n49445) );
  XNOR U49874 ( .A(n49499), .B(n49500), .Z(n49443) );
  XNOR U49875 ( .A(n49501), .B(n49502), .Z(n49500) );
  ANDN U49876 ( .B(B[2]), .A(n75), .Z(n47117) );
  XNOR U49877 ( .A(n47125), .B(n49503), .Z(n47118) );
  XNOR U49878 ( .A(n47124), .B(n47122), .Z(n49503) );
  AND U49879 ( .A(n49504), .B(n49505), .Z(n47122) );
  NANDN U49880 ( .A(n49502), .B(n49506), .Z(n49505) );
  NANDN U49881 ( .A(n49501), .B(n49499), .Z(n49506) );
  AND U49882 ( .A(n49507), .B(n49508), .Z(n49502) );
  NANDN U49883 ( .A(n49498), .B(n49509), .Z(n49508) );
  OR U49884 ( .A(n49497), .B(n49495), .Z(n49509) );
  AND U49885 ( .A(n49510), .B(n49511), .Z(n49498) );
  NANDN U49886 ( .A(n49494), .B(n49512), .Z(n49511) );
  NANDN U49887 ( .A(n49493), .B(n49491), .Z(n49512) );
  AND U49888 ( .A(n49513), .B(n49514), .Z(n49494) );
  NANDN U49889 ( .A(n49490), .B(n49515), .Z(n49514) );
  OR U49890 ( .A(n49489), .B(n49487), .Z(n49515) );
  AND U49891 ( .A(n49516), .B(n49517), .Z(n49490) );
  NANDN U49892 ( .A(n49486), .B(n49518), .Z(n49517) );
  NANDN U49893 ( .A(n49485), .B(n49483), .Z(n49518) );
  AND U49894 ( .A(n49519), .B(n49520), .Z(n49486) );
  NANDN U49895 ( .A(n49482), .B(n49521), .Z(n49520) );
  OR U49896 ( .A(n49481), .B(n49479), .Z(n49521) );
  AND U49897 ( .A(n49522), .B(n49523), .Z(n49482) );
  NANDN U49898 ( .A(n49477), .B(n49524), .Z(n49523) );
  NAND U49899 ( .A(n49475), .B(n49478), .Z(n49524) );
  NANDN U49900 ( .A(n49473), .B(n49525), .Z(n49477) );
  AND U49901 ( .A(A[0]), .B(B[4]), .Z(n49525) );
  NAND U49902 ( .A(B[3]), .B(A[1]), .Z(n49473) );
  XNOR U49903 ( .A(n49526), .B(n49527), .Z(n49475) );
  NAND U49904 ( .A(A[0]), .B(B[5]), .Z(n49527) );
  NAND U49905 ( .A(A[2]), .B(B[3]), .Z(n49478) );
  NAND U49906 ( .A(n49479), .B(n49481), .Z(n49519) );
  ANDN U49907 ( .B(B[3]), .A(n82), .Z(n49481) );
  XOR U49908 ( .A(n49528), .B(n49529), .Z(n49479) );
  XNOR U49909 ( .A(n49530), .B(n49531), .Z(n49529) );
  NANDN U49910 ( .A(n49483), .B(n49485), .Z(n49516) );
  ANDN U49911 ( .B(B[3]), .A(n81), .Z(n49485) );
  XNOR U49912 ( .A(n49532), .B(n49533), .Z(n49483) );
  XNOR U49913 ( .A(n49534), .B(n49535), .Z(n49533) );
  NAND U49914 ( .A(n49487), .B(n49489), .Z(n49513) );
  ANDN U49915 ( .B(B[3]), .A(n80), .Z(n49489) );
  XNOR U49916 ( .A(n49536), .B(n49537), .Z(n49487) );
  XNOR U49917 ( .A(n49538), .B(n49539), .Z(n49537) );
  NANDN U49918 ( .A(n49491), .B(n49493), .Z(n49510) );
  ANDN U49919 ( .B(B[3]), .A(n79), .Z(n49493) );
  XNOR U49920 ( .A(n49540), .B(n49541), .Z(n49491) );
  XNOR U49921 ( .A(n49542), .B(n49543), .Z(n49541) );
  NAND U49922 ( .A(n49495), .B(n49497), .Z(n49507) );
  ANDN U49923 ( .B(B[3]), .A(n78), .Z(n49497) );
  XNOR U49924 ( .A(n49544), .B(n49545), .Z(n49495) );
  XNOR U49925 ( .A(n49546), .B(n49547), .Z(n49545) );
  NANDN U49926 ( .A(n49499), .B(n49501), .Z(n49504) );
  ANDN U49927 ( .B(B[3]), .A(n77), .Z(n49501) );
  XNOR U49928 ( .A(n49548), .B(n49549), .Z(n49499) );
  XNOR U49929 ( .A(n49550), .B(n49551), .Z(n49549) );
  ANDN U49930 ( .B(B[3]), .A(n76), .Z(n47124) );
  XNOR U49931 ( .A(n47132), .B(n49552), .Z(n47125) );
  XNOR U49932 ( .A(n47131), .B(n47129), .Z(n49552) );
  AND U49933 ( .A(n49553), .B(n49554), .Z(n47129) );
  NANDN U49934 ( .A(n49551), .B(n49555), .Z(n49554) );
  OR U49935 ( .A(n49550), .B(n49548), .Z(n49555) );
  AND U49936 ( .A(n49556), .B(n49557), .Z(n49551) );
  NANDN U49937 ( .A(n49547), .B(n49558), .Z(n49557) );
  NANDN U49938 ( .A(n49546), .B(n49544), .Z(n49558) );
  AND U49939 ( .A(n49559), .B(n49560), .Z(n49547) );
  NANDN U49940 ( .A(n49543), .B(n49561), .Z(n49560) );
  OR U49941 ( .A(n49542), .B(n49540), .Z(n49561) );
  AND U49942 ( .A(n49562), .B(n49563), .Z(n49543) );
  NANDN U49943 ( .A(n49539), .B(n49564), .Z(n49563) );
  NANDN U49944 ( .A(n49538), .B(n49536), .Z(n49564) );
  AND U49945 ( .A(n49565), .B(n49566), .Z(n49539) );
  NANDN U49946 ( .A(n49535), .B(n49567), .Z(n49566) );
  OR U49947 ( .A(n49534), .B(n49532), .Z(n49567) );
  AND U49948 ( .A(n49568), .B(n49569), .Z(n49535) );
  NANDN U49949 ( .A(n49530), .B(n49570), .Z(n49569) );
  NAND U49950 ( .A(n49528), .B(n49531), .Z(n49570) );
  NANDN U49951 ( .A(n49526), .B(n49571), .Z(n49530) );
  AND U49952 ( .A(A[0]), .B(B[5]), .Z(n49571) );
  NAND U49953 ( .A(B[4]), .B(A[1]), .Z(n49526) );
  XNOR U49954 ( .A(n49572), .B(n49573), .Z(n49528) );
  NAND U49955 ( .A(A[0]), .B(B[6]), .Z(n49573) );
  NAND U49956 ( .A(A[2]), .B(B[4]), .Z(n49531) );
  NAND U49957 ( .A(n49532), .B(n49534), .Z(n49565) );
  ANDN U49958 ( .B(B[4]), .A(n82), .Z(n49534) );
  XOR U49959 ( .A(n49574), .B(n49575), .Z(n49532) );
  XNOR U49960 ( .A(n49576), .B(n49577), .Z(n49575) );
  NANDN U49961 ( .A(n49536), .B(n49538), .Z(n49562) );
  ANDN U49962 ( .B(B[4]), .A(n81), .Z(n49538) );
  XNOR U49963 ( .A(n49578), .B(n49579), .Z(n49536) );
  XNOR U49964 ( .A(n49580), .B(n49581), .Z(n49579) );
  NAND U49965 ( .A(n49540), .B(n49542), .Z(n49559) );
  ANDN U49966 ( .B(B[4]), .A(n80), .Z(n49542) );
  XNOR U49967 ( .A(n49582), .B(n49583), .Z(n49540) );
  XNOR U49968 ( .A(n49584), .B(n49585), .Z(n49583) );
  NANDN U49969 ( .A(n49544), .B(n49546), .Z(n49556) );
  ANDN U49970 ( .B(B[4]), .A(n79), .Z(n49546) );
  XNOR U49971 ( .A(n49586), .B(n49587), .Z(n49544) );
  XNOR U49972 ( .A(n49588), .B(n49589), .Z(n49587) );
  NAND U49973 ( .A(n49548), .B(n49550), .Z(n49553) );
  ANDN U49974 ( .B(B[4]), .A(n78), .Z(n49550) );
  XNOR U49975 ( .A(n49590), .B(n49591), .Z(n49548) );
  XNOR U49976 ( .A(n49592), .B(n49593), .Z(n49591) );
  ANDN U49977 ( .B(B[4]), .A(n77), .Z(n47131) );
  XNOR U49978 ( .A(n47139), .B(n49594), .Z(n47132) );
  XNOR U49979 ( .A(n47138), .B(n47136), .Z(n49594) );
  AND U49980 ( .A(n49595), .B(n49596), .Z(n47136) );
  NANDN U49981 ( .A(n49593), .B(n49597), .Z(n49596) );
  NANDN U49982 ( .A(n49592), .B(n49590), .Z(n49597) );
  AND U49983 ( .A(n49598), .B(n49599), .Z(n49593) );
  NANDN U49984 ( .A(n49589), .B(n49600), .Z(n49599) );
  OR U49985 ( .A(n49588), .B(n49586), .Z(n49600) );
  AND U49986 ( .A(n49601), .B(n49602), .Z(n49589) );
  NANDN U49987 ( .A(n49585), .B(n49603), .Z(n49602) );
  NANDN U49988 ( .A(n49584), .B(n49582), .Z(n49603) );
  AND U49989 ( .A(n49604), .B(n49605), .Z(n49585) );
  NANDN U49990 ( .A(n49581), .B(n49606), .Z(n49605) );
  OR U49991 ( .A(n49580), .B(n49578), .Z(n49606) );
  AND U49992 ( .A(n49607), .B(n49608), .Z(n49581) );
  NANDN U49993 ( .A(n49576), .B(n49609), .Z(n49608) );
  NAND U49994 ( .A(n49574), .B(n49577), .Z(n49609) );
  NANDN U49995 ( .A(n49572), .B(n49610), .Z(n49576) );
  AND U49996 ( .A(A[0]), .B(B[6]), .Z(n49610) );
  NAND U49997 ( .A(B[5]), .B(A[1]), .Z(n49572) );
  XNOR U49998 ( .A(n49611), .B(n49612), .Z(n49574) );
  NAND U49999 ( .A(A[0]), .B(B[7]), .Z(n49612) );
  NAND U50000 ( .A(A[2]), .B(B[5]), .Z(n49577) );
  NAND U50001 ( .A(n49578), .B(n49580), .Z(n49604) );
  ANDN U50002 ( .B(B[5]), .A(n82), .Z(n49580) );
  XOR U50003 ( .A(n49613), .B(n49614), .Z(n49578) );
  XNOR U50004 ( .A(n49615), .B(n49616), .Z(n49614) );
  NANDN U50005 ( .A(n49582), .B(n49584), .Z(n49601) );
  ANDN U50006 ( .B(B[5]), .A(n81), .Z(n49584) );
  XNOR U50007 ( .A(n49617), .B(n49618), .Z(n49582) );
  XNOR U50008 ( .A(n49619), .B(n49620), .Z(n49618) );
  NAND U50009 ( .A(n49586), .B(n49588), .Z(n49598) );
  ANDN U50010 ( .B(B[5]), .A(n80), .Z(n49588) );
  XNOR U50011 ( .A(n49621), .B(n49622), .Z(n49586) );
  XNOR U50012 ( .A(n49623), .B(n49624), .Z(n49622) );
  NANDN U50013 ( .A(n49590), .B(n49592), .Z(n49595) );
  ANDN U50014 ( .B(B[5]), .A(n79), .Z(n49592) );
  XNOR U50015 ( .A(n49625), .B(n49626), .Z(n49590) );
  XNOR U50016 ( .A(n49627), .B(n49628), .Z(n49626) );
  ANDN U50017 ( .B(B[5]), .A(n78), .Z(n47138) );
  XNOR U50018 ( .A(n47146), .B(n49629), .Z(n47139) );
  XNOR U50019 ( .A(n47145), .B(n47143), .Z(n49629) );
  AND U50020 ( .A(n49630), .B(n49631), .Z(n47143) );
  NANDN U50021 ( .A(n49628), .B(n49632), .Z(n49631) );
  OR U50022 ( .A(n49627), .B(n49625), .Z(n49632) );
  AND U50023 ( .A(n49633), .B(n49634), .Z(n49628) );
  NANDN U50024 ( .A(n49624), .B(n49635), .Z(n49634) );
  NANDN U50025 ( .A(n49623), .B(n49621), .Z(n49635) );
  AND U50026 ( .A(n49636), .B(n49637), .Z(n49624) );
  NANDN U50027 ( .A(n49620), .B(n49638), .Z(n49637) );
  OR U50028 ( .A(n49619), .B(n49617), .Z(n49638) );
  AND U50029 ( .A(n49639), .B(n49640), .Z(n49620) );
  NANDN U50030 ( .A(n49615), .B(n49641), .Z(n49640) );
  NAND U50031 ( .A(n49613), .B(n49616), .Z(n49641) );
  NANDN U50032 ( .A(n49611), .B(n49642), .Z(n49615) );
  AND U50033 ( .A(A[0]), .B(B[7]), .Z(n49642) );
  NAND U50034 ( .A(B[6]), .B(A[1]), .Z(n49611) );
  XNOR U50035 ( .A(n49643), .B(n49644), .Z(n49613) );
  NAND U50036 ( .A(A[0]), .B(B[8]), .Z(n49644) );
  NAND U50037 ( .A(A[2]), .B(B[6]), .Z(n49616) );
  NAND U50038 ( .A(n49617), .B(n49619), .Z(n49636) );
  ANDN U50039 ( .B(B[6]), .A(n82), .Z(n49619) );
  XOR U50040 ( .A(n49645), .B(n49646), .Z(n49617) );
  XNOR U50041 ( .A(n49647), .B(n49648), .Z(n49646) );
  NANDN U50042 ( .A(n49621), .B(n49623), .Z(n49633) );
  ANDN U50043 ( .B(B[6]), .A(n81), .Z(n49623) );
  XNOR U50044 ( .A(n49649), .B(n49650), .Z(n49621) );
  XNOR U50045 ( .A(n49651), .B(n49652), .Z(n49650) );
  NAND U50046 ( .A(n49625), .B(n49627), .Z(n49630) );
  ANDN U50047 ( .B(B[6]), .A(n80), .Z(n49627) );
  XNOR U50048 ( .A(n49653), .B(n49654), .Z(n49625) );
  XNOR U50049 ( .A(n49655), .B(n49656), .Z(n49654) );
  ANDN U50050 ( .B(B[6]), .A(n79), .Z(n47145) );
  XNOR U50051 ( .A(n47153), .B(n49657), .Z(n47146) );
  XNOR U50052 ( .A(n47152), .B(n47150), .Z(n49657) );
  AND U50053 ( .A(n49658), .B(n49659), .Z(n47150) );
  NANDN U50054 ( .A(n49656), .B(n49660), .Z(n49659) );
  NANDN U50055 ( .A(n49655), .B(n49653), .Z(n49660) );
  AND U50056 ( .A(n49661), .B(n49662), .Z(n49656) );
  NANDN U50057 ( .A(n49652), .B(n49663), .Z(n49662) );
  OR U50058 ( .A(n49651), .B(n49649), .Z(n49663) );
  AND U50059 ( .A(n49664), .B(n49665), .Z(n49652) );
  NANDN U50060 ( .A(n49647), .B(n49666), .Z(n49665) );
  NAND U50061 ( .A(n49645), .B(n49648), .Z(n49666) );
  NANDN U50062 ( .A(n49643), .B(n49667), .Z(n49647) );
  AND U50063 ( .A(A[0]), .B(B[8]), .Z(n49667) );
  NAND U50064 ( .A(B[7]), .B(A[1]), .Z(n49643) );
  XNOR U50065 ( .A(n49668), .B(n49669), .Z(n49645) );
  NAND U50066 ( .A(A[0]), .B(B[9]), .Z(n49669) );
  NAND U50067 ( .A(A[2]), .B(B[7]), .Z(n49648) );
  NAND U50068 ( .A(n49649), .B(n49651), .Z(n49661) );
  ANDN U50069 ( .B(B[7]), .A(n82), .Z(n49651) );
  XOR U50070 ( .A(n49670), .B(n49671), .Z(n49649) );
  XNOR U50071 ( .A(n49672), .B(n49673), .Z(n49671) );
  NANDN U50072 ( .A(n49653), .B(n49655), .Z(n49658) );
  ANDN U50073 ( .B(B[7]), .A(n81), .Z(n49655) );
  XNOR U50074 ( .A(n49674), .B(n49675), .Z(n49653) );
  XNOR U50075 ( .A(n49676), .B(n49677), .Z(n49675) );
  ANDN U50076 ( .B(B[7]), .A(n80), .Z(n47152) );
  XNOR U50077 ( .A(n47160), .B(n49678), .Z(n47153) );
  XNOR U50078 ( .A(n47159), .B(n47157), .Z(n49678) );
  AND U50079 ( .A(n49679), .B(n49680), .Z(n47157) );
  NANDN U50080 ( .A(n49677), .B(n49681), .Z(n49680) );
  OR U50081 ( .A(n49676), .B(n49674), .Z(n49681) );
  AND U50082 ( .A(n49682), .B(n49683), .Z(n49677) );
  NANDN U50083 ( .A(n49672), .B(n49684), .Z(n49683) );
  NAND U50084 ( .A(n49670), .B(n49673), .Z(n49684) );
  NANDN U50085 ( .A(n49668), .B(n49685), .Z(n49672) );
  AND U50086 ( .A(A[0]), .B(B[9]), .Z(n49685) );
  NAND U50087 ( .A(B[8]), .B(A[1]), .Z(n49668) );
  XNOR U50088 ( .A(n49686), .B(n49687), .Z(n49670) );
  NAND U50089 ( .A(A[0]), .B(B[10]), .Z(n49687) );
  NAND U50090 ( .A(A[2]), .B(B[8]), .Z(n49673) );
  NAND U50091 ( .A(n49674), .B(n49676), .Z(n49679) );
  ANDN U50092 ( .B(B[8]), .A(n82), .Z(n49676) );
  XOR U50093 ( .A(n49688), .B(n49689), .Z(n49674) );
  XNOR U50094 ( .A(n49690), .B(n49691), .Z(n49689) );
  ANDN U50095 ( .B(B[8]), .A(n81), .Z(n47159) );
  XNOR U50096 ( .A(n47167), .B(n49692), .Z(n47160) );
  XNOR U50097 ( .A(n47166), .B(n47164), .Z(n49692) );
  AND U50098 ( .A(n49693), .B(n49694), .Z(n47164) );
  NANDN U50099 ( .A(n49690), .B(n49695), .Z(n49694) );
  NAND U50100 ( .A(n49688), .B(n49691), .Z(n49695) );
  NANDN U50101 ( .A(n49686), .B(n49696), .Z(n49690) );
  AND U50102 ( .A(A[0]), .B(B[10]), .Z(n49696) );
  NAND U50103 ( .A(B[9]), .B(A[1]), .Z(n49686) );
  XNOR U50104 ( .A(n49697), .B(n49698), .Z(n49688) );
  NAND U50105 ( .A(A[0]), .B(B[11]), .Z(n49698) );
  NAND U50106 ( .A(A[2]), .B(B[9]), .Z(n49691) );
  ANDN U50107 ( .B(B[9]), .A(n82), .Z(n47166) );
  XOR U50108 ( .A(n47173), .B(n49699), .Z(n47167) );
  XNOR U50109 ( .A(n47171), .B(n47174), .Z(n49699) );
  NAND U50110 ( .A(A[2]), .B(B[10]), .Z(n47174) );
  NANDN U50111 ( .A(n49697), .B(n49700), .Z(n47171) );
  AND U50112 ( .A(A[0]), .B(B[11]), .Z(n49700) );
  NAND U50113 ( .A(B[10]), .B(A[1]), .Z(n49697) );
  XNOR U50114 ( .A(n47176), .B(n49701), .Z(n47173) );
  NAND U50115 ( .A(A[0]), .B(B[12]), .Z(n49701) );
  NAND U50116 ( .A(B[11]), .B(A[1]), .Z(n47176) );
  XOR U50117 ( .A(n574), .B(n573), .Z(\A1[109] ) );
  XOR U50118 ( .A(n49308), .B(n49702), .Z(n573) );
  XNOR U50119 ( .A(n49307), .B(n49305), .Z(n49702) );
  AND U50120 ( .A(n49703), .B(n49704), .Z(n49305) );
  NANDN U50121 ( .A(n49705), .B(n49706), .Z(n49704) );
  NANDN U50122 ( .A(n49707), .B(n49708), .Z(n49706) );
  NANDN U50123 ( .A(n49708), .B(n49707), .Z(n49703) );
  ANDN U50124 ( .B(B[80]), .A(n54), .Z(n49307) );
  XNOR U50125 ( .A(n49102), .B(n49709), .Z(n49308) );
  XNOR U50126 ( .A(n49101), .B(n49099), .Z(n49709) );
  AND U50127 ( .A(n49710), .B(n49711), .Z(n49099) );
  NANDN U50128 ( .A(n49712), .B(n49713), .Z(n49711) );
  OR U50129 ( .A(n49714), .B(n49715), .Z(n49713) );
  NAND U50130 ( .A(n49715), .B(n49714), .Z(n49710) );
  ANDN U50131 ( .B(B[81]), .A(n55), .Z(n49101) );
  XNOR U50132 ( .A(n49109), .B(n49716), .Z(n49102) );
  XNOR U50133 ( .A(n49108), .B(n49106), .Z(n49716) );
  AND U50134 ( .A(n49717), .B(n49718), .Z(n49106) );
  NANDN U50135 ( .A(n49719), .B(n49720), .Z(n49718) );
  NANDN U50136 ( .A(n49721), .B(n49722), .Z(n49720) );
  NANDN U50137 ( .A(n49722), .B(n49721), .Z(n49717) );
  ANDN U50138 ( .B(B[82]), .A(n56), .Z(n49108) );
  XNOR U50139 ( .A(n49116), .B(n49723), .Z(n49109) );
  XNOR U50140 ( .A(n49115), .B(n49113), .Z(n49723) );
  AND U50141 ( .A(n49724), .B(n49725), .Z(n49113) );
  NANDN U50142 ( .A(n49726), .B(n49727), .Z(n49725) );
  OR U50143 ( .A(n49728), .B(n49729), .Z(n49727) );
  NAND U50144 ( .A(n49729), .B(n49728), .Z(n49724) );
  ANDN U50145 ( .B(B[83]), .A(n57), .Z(n49115) );
  XNOR U50146 ( .A(n49123), .B(n49730), .Z(n49116) );
  XNOR U50147 ( .A(n49122), .B(n49120), .Z(n49730) );
  AND U50148 ( .A(n49731), .B(n49732), .Z(n49120) );
  NANDN U50149 ( .A(n49733), .B(n49734), .Z(n49732) );
  NANDN U50150 ( .A(n49735), .B(n49736), .Z(n49734) );
  NANDN U50151 ( .A(n49736), .B(n49735), .Z(n49731) );
  ANDN U50152 ( .B(B[84]), .A(n58), .Z(n49122) );
  XNOR U50153 ( .A(n49130), .B(n49737), .Z(n49123) );
  XNOR U50154 ( .A(n49129), .B(n49127), .Z(n49737) );
  AND U50155 ( .A(n49738), .B(n49739), .Z(n49127) );
  NANDN U50156 ( .A(n49740), .B(n49741), .Z(n49739) );
  OR U50157 ( .A(n49742), .B(n49743), .Z(n49741) );
  NAND U50158 ( .A(n49743), .B(n49742), .Z(n49738) );
  ANDN U50159 ( .B(B[85]), .A(n59), .Z(n49129) );
  XNOR U50160 ( .A(n49137), .B(n49744), .Z(n49130) );
  XNOR U50161 ( .A(n49136), .B(n49134), .Z(n49744) );
  AND U50162 ( .A(n49745), .B(n49746), .Z(n49134) );
  NANDN U50163 ( .A(n49747), .B(n49748), .Z(n49746) );
  NANDN U50164 ( .A(n49749), .B(n49750), .Z(n49748) );
  NANDN U50165 ( .A(n49750), .B(n49749), .Z(n49745) );
  ANDN U50166 ( .B(B[86]), .A(n60), .Z(n49136) );
  XNOR U50167 ( .A(n49144), .B(n49751), .Z(n49137) );
  XNOR U50168 ( .A(n49143), .B(n49141), .Z(n49751) );
  AND U50169 ( .A(n49752), .B(n49753), .Z(n49141) );
  NANDN U50170 ( .A(n49754), .B(n49755), .Z(n49753) );
  OR U50171 ( .A(n49756), .B(n49757), .Z(n49755) );
  NAND U50172 ( .A(n49757), .B(n49756), .Z(n49752) );
  ANDN U50173 ( .B(B[87]), .A(n61), .Z(n49143) );
  XNOR U50174 ( .A(n49151), .B(n49758), .Z(n49144) );
  XNOR U50175 ( .A(n49150), .B(n49148), .Z(n49758) );
  AND U50176 ( .A(n49759), .B(n49760), .Z(n49148) );
  NANDN U50177 ( .A(n49761), .B(n49762), .Z(n49760) );
  NANDN U50178 ( .A(n49763), .B(n49764), .Z(n49762) );
  NANDN U50179 ( .A(n49764), .B(n49763), .Z(n49759) );
  ANDN U50180 ( .B(B[88]), .A(n62), .Z(n49150) );
  XNOR U50181 ( .A(n49158), .B(n49765), .Z(n49151) );
  XNOR U50182 ( .A(n49157), .B(n49155), .Z(n49765) );
  AND U50183 ( .A(n49766), .B(n49767), .Z(n49155) );
  NANDN U50184 ( .A(n49768), .B(n49769), .Z(n49767) );
  OR U50185 ( .A(n49770), .B(n49771), .Z(n49769) );
  NAND U50186 ( .A(n49771), .B(n49770), .Z(n49766) );
  ANDN U50187 ( .B(B[89]), .A(n63), .Z(n49157) );
  XNOR U50188 ( .A(n49165), .B(n49772), .Z(n49158) );
  XNOR U50189 ( .A(n49164), .B(n49162), .Z(n49772) );
  AND U50190 ( .A(n49773), .B(n49774), .Z(n49162) );
  NANDN U50191 ( .A(n49775), .B(n49776), .Z(n49774) );
  NANDN U50192 ( .A(n49777), .B(n49778), .Z(n49776) );
  NANDN U50193 ( .A(n49778), .B(n49777), .Z(n49773) );
  ANDN U50194 ( .B(A[21]), .A(n23), .Z(n49164) );
  XNOR U50195 ( .A(n49172), .B(n49779), .Z(n49165) );
  XNOR U50196 ( .A(n49171), .B(n49169), .Z(n49779) );
  AND U50197 ( .A(n49780), .B(n49781), .Z(n49169) );
  NANDN U50198 ( .A(n49782), .B(n49783), .Z(n49781) );
  OR U50199 ( .A(n49784), .B(n49785), .Z(n49783) );
  NAND U50200 ( .A(n49785), .B(n49784), .Z(n49780) );
  ANDN U50201 ( .B(A[20]), .A(n21), .Z(n49171) );
  XNOR U50202 ( .A(n49179), .B(n49786), .Z(n49172) );
  XNOR U50203 ( .A(n49178), .B(n49176), .Z(n49786) );
  AND U50204 ( .A(n49787), .B(n49788), .Z(n49176) );
  NANDN U50205 ( .A(n49789), .B(n49790), .Z(n49788) );
  NANDN U50206 ( .A(n49791), .B(n49792), .Z(n49790) );
  NANDN U50207 ( .A(n49792), .B(n49791), .Z(n49787) );
  ANDN U50208 ( .B(A[19]), .A(n19), .Z(n49178) );
  XNOR U50209 ( .A(n49186), .B(n49793), .Z(n49179) );
  XNOR U50210 ( .A(n49185), .B(n49183), .Z(n49793) );
  AND U50211 ( .A(n49794), .B(n49795), .Z(n49183) );
  NANDN U50212 ( .A(n49796), .B(n49797), .Z(n49795) );
  OR U50213 ( .A(n49798), .B(n49799), .Z(n49797) );
  NAND U50214 ( .A(n49799), .B(n49798), .Z(n49794) );
  ANDN U50215 ( .B(A[18]), .A(n17), .Z(n49185) );
  XNOR U50216 ( .A(n49193), .B(n49800), .Z(n49186) );
  XNOR U50217 ( .A(n49192), .B(n49190), .Z(n49800) );
  AND U50218 ( .A(n49801), .B(n49802), .Z(n49190) );
  NANDN U50219 ( .A(n49803), .B(n49804), .Z(n49802) );
  NANDN U50220 ( .A(n49805), .B(n49806), .Z(n49804) );
  NANDN U50221 ( .A(n49806), .B(n49805), .Z(n49801) );
  ANDN U50222 ( .B(A[17]), .A(n15), .Z(n49192) );
  XNOR U50223 ( .A(n49200), .B(n49807), .Z(n49193) );
  XNOR U50224 ( .A(n49199), .B(n49197), .Z(n49807) );
  AND U50225 ( .A(n49808), .B(n49809), .Z(n49197) );
  NANDN U50226 ( .A(n49810), .B(n49811), .Z(n49809) );
  OR U50227 ( .A(n49812), .B(n49813), .Z(n49811) );
  NAND U50228 ( .A(n49813), .B(n49812), .Z(n49808) );
  ANDN U50229 ( .B(A[16]), .A(n13), .Z(n49199) );
  XNOR U50230 ( .A(n49207), .B(n49814), .Z(n49200) );
  XNOR U50231 ( .A(n49206), .B(n49204), .Z(n49814) );
  AND U50232 ( .A(n49815), .B(n49816), .Z(n49204) );
  NANDN U50233 ( .A(n49817), .B(n49818), .Z(n49816) );
  NANDN U50234 ( .A(n49819), .B(n49820), .Z(n49818) );
  NANDN U50235 ( .A(n49820), .B(n49819), .Z(n49815) );
  ANDN U50236 ( .B(A[15]), .A(n11), .Z(n49206) );
  XNOR U50237 ( .A(n49214), .B(n49821), .Z(n49207) );
  XNOR U50238 ( .A(n49213), .B(n49211), .Z(n49821) );
  AND U50239 ( .A(n49822), .B(n49823), .Z(n49211) );
  NANDN U50240 ( .A(n49824), .B(n49825), .Z(n49823) );
  OR U50241 ( .A(n49826), .B(n49827), .Z(n49825) );
  NAND U50242 ( .A(n49827), .B(n49826), .Z(n49822) );
  ANDN U50243 ( .B(A[14]), .A(n9), .Z(n49213) );
  XNOR U50244 ( .A(n49221), .B(n49828), .Z(n49214) );
  XNOR U50245 ( .A(n49220), .B(n49218), .Z(n49828) );
  AND U50246 ( .A(n49829), .B(n49830), .Z(n49218) );
  NANDN U50247 ( .A(n49831), .B(n49832), .Z(n49830) );
  NANDN U50248 ( .A(n49833), .B(n49834), .Z(n49832) );
  NANDN U50249 ( .A(n49834), .B(n49833), .Z(n49829) );
  ANDN U50250 ( .B(B[98]), .A(n72), .Z(n49220) );
  XNOR U50251 ( .A(n49228), .B(n49835), .Z(n49221) );
  XNOR U50252 ( .A(n49227), .B(n49225), .Z(n49835) );
  AND U50253 ( .A(n49836), .B(n49837), .Z(n49225) );
  NANDN U50254 ( .A(n49838), .B(n49839), .Z(n49837) );
  OR U50255 ( .A(n49840), .B(n49841), .Z(n49839) );
  NAND U50256 ( .A(n49841), .B(n49840), .Z(n49836) );
  ANDN U50257 ( .B(A[12]), .A(n6), .Z(n49227) );
  XNOR U50258 ( .A(n49235), .B(n49842), .Z(n49228) );
  XNOR U50259 ( .A(n49234), .B(n49232), .Z(n49842) );
  AND U50260 ( .A(n49843), .B(n49844), .Z(n49232) );
  NANDN U50261 ( .A(n49845), .B(n49846), .Z(n49844) );
  NANDN U50262 ( .A(n49847), .B(n49848), .Z(n49846) );
  NANDN U50263 ( .A(n49848), .B(n49847), .Z(n49843) );
  ANDN U50264 ( .B(A[11]), .A(n4), .Z(n49234) );
  XNOR U50265 ( .A(n49242), .B(n49849), .Z(n49235) );
  XNOR U50266 ( .A(n49241), .B(n49239), .Z(n49849) );
  AND U50267 ( .A(n49850), .B(n49851), .Z(n49239) );
  NANDN U50268 ( .A(n49852), .B(n49853), .Z(n49851) );
  OR U50269 ( .A(n49854), .B(n49855), .Z(n49853) );
  NAND U50270 ( .A(n49855), .B(n49854), .Z(n49850) );
  ANDN U50271 ( .B(B[101]), .A(n75), .Z(n49241) );
  XNOR U50272 ( .A(n49249), .B(n49856), .Z(n49242) );
  XNOR U50273 ( .A(n49248), .B(n49246), .Z(n49856) );
  AND U50274 ( .A(n49857), .B(n49858), .Z(n49246) );
  NANDN U50275 ( .A(n49859), .B(n49860), .Z(n49858) );
  NANDN U50276 ( .A(n49861), .B(n49862), .Z(n49860) );
  NANDN U50277 ( .A(n49862), .B(n49861), .Z(n49857) );
  ANDN U50278 ( .B(B[102]), .A(n76), .Z(n49248) );
  XNOR U50279 ( .A(n49256), .B(n49863), .Z(n49249) );
  XNOR U50280 ( .A(n49255), .B(n49253), .Z(n49863) );
  AND U50281 ( .A(n49864), .B(n49865), .Z(n49253) );
  NANDN U50282 ( .A(n49866), .B(n49867), .Z(n49865) );
  OR U50283 ( .A(n49868), .B(n49869), .Z(n49867) );
  NAND U50284 ( .A(n49869), .B(n49868), .Z(n49864) );
  ANDN U50285 ( .B(B[103]), .A(n77), .Z(n49255) );
  XNOR U50286 ( .A(n49263), .B(n49870), .Z(n49256) );
  XNOR U50287 ( .A(n49262), .B(n49260), .Z(n49870) );
  AND U50288 ( .A(n49871), .B(n49872), .Z(n49260) );
  NANDN U50289 ( .A(n49873), .B(n49874), .Z(n49872) );
  NANDN U50290 ( .A(n49875), .B(n49876), .Z(n49874) );
  NANDN U50291 ( .A(n49876), .B(n49875), .Z(n49871) );
  ANDN U50292 ( .B(B[104]), .A(n78), .Z(n49262) );
  XNOR U50293 ( .A(n49270), .B(n49877), .Z(n49263) );
  XNOR U50294 ( .A(n49269), .B(n49267), .Z(n49877) );
  AND U50295 ( .A(n49878), .B(n49879), .Z(n49267) );
  NANDN U50296 ( .A(n49880), .B(n49881), .Z(n49879) );
  OR U50297 ( .A(n49882), .B(n49883), .Z(n49881) );
  NAND U50298 ( .A(n49883), .B(n49882), .Z(n49878) );
  ANDN U50299 ( .B(B[105]), .A(n79), .Z(n49269) );
  XNOR U50300 ( .A(n49277), .B(n49884), .Z(n49270) );
  XNOR U50301 ( .A(n49276), .B(n49274), .Z(n49884) );
  AND U50302 ( .A(n49885), .B(n49886), .Z(n49274) );
  NANDN U50303 ( .A(n49887), .B(n49888), .Z(n49886) );
  NANDN U50304 ( .A(n49889), .B(n49890), .Z(n49888) );
  NANDN U50305 ( .A(n49890), .B(n49889), .Z(n49885) );
  ANDN U50306 ( .B(B[106]), .A(n80), .Z(n49276) );
  XNOR U50307 ( .A(n49284), .B(n49891), .Z(n49277) );
  XNOR U50308 ( .A(n49283), .B(n49281), .Z(n49891) );
  AND U50309 ( .A(n49892), .B(n49893), .Z(n49281) );
  NANDN U50310 ( .A(n49894), .B(n49895), .Z(n49893) );
  OR U50311 ( .A(n49896), .B(n49897), .Z(n49895) );
  NAND U50312 ( .A(n49897), .B(n49896), .Z(n49892) );
  ANDN U50313 ( .B(B[107]), .A(n81), .Z(n49283) );
  XNOR U50314 ( .A(n49291), .B(n49898), .Z(n49284) );
  XNOR U50315 ( .A(n49290), .B(n49288), .Z(n49898) );
  AND U50316 ( .A(n49899), .B(n49900), .Z(n49288) );
  NANDN U50317 ( .A(n49901), .B(n49902), .Z(n49900) );
  NAND U50318 ( .A(n49903), .B(n49904), .Z(n49902) );
  ANDN U50319 ( .B(B[108]), .A(n82), .Z(n49290) );
  XOR U50320 ( .A(n49297), .B(n49905), .Z(n49291) );
  XNOR U50321 ( .A(n49295), .B(n49298), .Z(n49905) );
  NAND U50322 ( .A(A[2]), .B(B[109]), .Z(n49298) );
  NANDN U50323 ( .A(n49906), .B(n49907), .Z(n49295) );
  AND U50324 ( .A(A[0]), .B(B[110]), .Z(n49907) );
  XNOR U50325 ( .A(n49300), .B(n49908), .Z(n49297) );
  NAND U50326 ( .A(A[0]), .B(B[111]), .Z(n49908) );
  NAND U50327 ( .A(B[110]), .B(A[1]), .Z(n49300) );
  NAND U50328 ( .A(n49909), .B(n49910), .Z(n574) );
  NANDN U50329 ( .A(n49911), .B(n49912), .Z(n49910) );
  OR U50330 ( .A(n49913), .B(n49914), .Z(n49912) );
  NAND U50331 ( .A(n49914), .B(n49913), .Z(n49909) );
  XOR U50332 ( .A(n576), .B(n575), .Z(\A1[108] ) );
  XOR U50333 ( .A(n49914), .B(n49915), .Z(n575) );
  XNOR U50334 ( .A(n49913), .B(n49911), .Z(n49915) );
  AND U50335 ( .A(n49916), .B(n49917), .Z(n49911) );
  NANDN U50336 ( .A(n49918), .B(n49919), .Z(n49917) );
  NANDN U50337 ( .A(n49920), .B(n49921), .Z(n49919) );
  NANDN U50338 ( .A(n49921), .B(n49920), .Z(n49916) );
  ANDN U50339 ( .B(B[79]), .A(n54), .Z(n49913) );
  XNOR U50340 ( .A(n49708), .B(n49922), .Z(n49914) );
  XNOR U50341 ( .A(n49707), .B(n49705), .Z(n49922) );
  AND U50342 ( .A(n49923), .B(n49924), .Z(n49705) );
  NANDN U50343 ( .A(n49925), .B(n49926), .Z(n49924) );
  OR U50344 ( .A(n49927), .B(n49928), .Z(n49926) );
  NAND U50345 ( .A(n49928), .B(n49927), .Z(n49923) );
  ANDN U50346 ( .B(B[80]), .A(n55), .Z(n49707) );
  XNOR U50347 ( .A(n49715), .B(n49929), .Z(n49708) );
  XNOR U50348 ( .A(n49714), .B(n49712), .Z(n49929) );
  AND U50349 ( .A(n49930), .B(n49931), .Z(n49712) );
  NANDN U50350 ( .A(n49932), .B(n49933), .Z(n49931) );
  NANDN U50351 ( .A(n49934), .B(n49935), .Z(n49933) );
  NANDN U50352 ( .A(n49935), .B(n49934), .Z(n49930) );
  ANDN U50353 ( .B(B[81]), .A(n56), .Z(n49714) );
  XNOR U50354 ( .A(n49722), .B(n49936), .Z(n49715) );
  XNOR U50355 ( .A(n49721), .B(n49719), .Z(n49936) );
  AND U50356 ( .A(n49937), .B(n49938), .Z(n49719) );
  NANDN U50357 ( .A(n49939), .B(n49940), .Z(n49938) );
  OR U50358 ( .A(n49941), .B(n49942), .Z(n49940) );
  NAND U50359 ( .A(n49942), .B(n49941), .Z(n49937) );
  ANDN U50360 ( .B(B[82]), .A(n57), .Z(n49721) );
  XNOR U50361 ( .A(n49729), .B(n49943), .Z(n49722) );
  XNOR U50362 ( .A(n49728), .B(n49726), .Z(n49943) );
  AND U50363 ( .A(n49944), .B(n49945), .Z(n49726) );
  NANDN U50364 ( .A(n49946), .B(n49947), .Z(n49945) );
  NANDN U50365 ( .A(n49948), .B(n49949), .Z(n49947) );
  NANDN U50366 ( .A(n49949), .B(n49948), .Z(n49944) );
  ANDN U50367 ( .B(B[83]), .A(n58), .Z(n49728) );
  XNOR U50368 ( .A(n49736), .B(n49950), .Z(n49729) );
  XNOR U50369 ( .A(n49735), .B(n49733), .Z(n49950) );
  AND U50370 ( .A(n49951), .B(n49952), .Z(n49733) );
  NANDN U50371 ( .A(n49953), .B(n49954), .Z(n49952) );
  OR U50372 ( .A(n49955), .B(n49956), .Z(n49954) );
  NAND U50373 ( .A(n49956), .B(n49955), .Z(n49951) );
  ANDN U50374 ( .B(B[84]), .A(n59), .Z(n49735) );
  XNOR U50375 ( .A(n49743), .B(n49957), .Z(n49736) );
  XNOR U50376 ( .A(n49742), .B(n49740), .Z(n49957) );
  AND U50377 ( .A(n49958), .B(n49959), .Z(n49740) );
  NANDN U50378 ( .A(n49960), .B(n49961), .Z(n49959) );
  NANDN U50379 ( .A(n49962), .B(n49963), .Z(n49961) );
  NANDN U50380 ( .A(n49963), .B(n49962), .Z(n49958) );
  ANDN U50381 ( .B(B[85]), .A(n60), .Z(n49742) );
  XNOR U50382 ( .A(n49750), .B(n49964), .Z(n49743) );
  XNOR U50383 ( .A(n49749), .B(n49747), .Z(n49964) );
  AND U50384 ( .A(n49965), .B(n49966), .Z(n49747) );
  NANDN U50385 ( .A(n49967), .B(n49968), .Z(n49966) );
  OR U50386 ( .A(n49969), .B(n49970), .Z(n49968) );
  NAND U50387 ( .A(n49970), .B(n49969), .Z(n49965) );
  ANDN U50388 ( .B(B[86]), .A(n61), .Z(n49749) );
  XNOR U50389 ( .A(n49757), .B(n49971), .Z(n49750) );
  XNOR U50390 ( .A(n49756), .B(n49754), .Z(n49971) );
  AND U50391 ( .A(n49972), .B(n49973), .Z(n49754) );
  NANDN U50392 ( .A(n49974), .B(n49975), .Z(n49973) );
  NANDN U50393 ( .A(n49976), .B(n49977), .Z(n49975) );
  NANDN U50394 ( .A(n49977), .B(n49976), .Z(n49972) );
  ANDN U50395 ( .B(B[87]), .A(n62), .Z(n49756) );
  XNOR U50396 ( .A(n49764), .B(n49978), .Z(n49757) );
  XNOR U50397 ( .A(n49763), .B(n49761), .Z(n49978) );
  AND U50398 ( .A(n49979), .B(n49980), .Z(n49761) );
  NANDN U50399 ( .A(n49981), .B(n49982), .Z(n49980) );
  OR U50400 ( .A(n49983), .B(n49984), .Z(n49982) );
  NAND U50401 ( .A(n49984), .B(n49983), .Z(n49979) );
  ANDN U50402 ( .B(B[88]), .A(n63), .Z(n49763) );
  XNOR U50403 ( .A(n49771), .B(n49985), .Z(n49764) );
  XNOR U50404 ( .A(n49770), .B(n49768), .Z(n49985) );
  AND U50405 ( .A(n49986), .B(n49987), .Z(n49768) );
  NANDN U50406 ( .A(n49988), .B(n49989), .Z(n49987) );
  NANDN U50407 ( .A(n49990), .B(n49991), .Z(n49989) );
  NANDN U50408 ( .A(n49991), .B(n49990), .Z(n49986) );
  ANDN U50409 ( .B(A[21]), .A(n25), .Z(n49770) );
  XNOR U50410 ( .A(n49778), .B(n49992), .Z(n49771) );
  XNOR U50411 ( .A(n49777), .B(n49775), .Z(n49992) );
  AND U50412 ( .A(n49993), .B(n49994), .Z(n49775) );
  NANDN U50413 ( .A(n49995), .B(n49996), .Z(n49994) );
  OR U50414 ( .A(n49997), .B(n49998), .Z(n49996) );
  NAND U50415 ( .A(n49998), .B(n49997), .Z(n49993) );
  ANDN U50416 ( .B(A[20]), .A(n23), .Z(n49777) );
  XNOR U50417 ( .A(n49785), .B(n49999), .Z(n49778) );
  XNOR U50418 ( .A(n49784), .B(n49782), .Z(n49999) );
  AND U50419 ( .A(n50000), .B(n50001), .Z(n49782) );
  NANDN U50420 ( .A(n50002), .B(n50003), .Z(n50001) );
  NANDN U50421 ( .A(n50004), .B(n50005), .Z(n50003) );
  NANDN U50422 ( .A(n50005), .B(n50004), .Z(n50000) );
  ANDN U50423 ( .B(A[19]), .A(n21), .Z(n49784) );
  XNOR U50424 ( .A(n49792), .B(n50006), .Z(n49785) );
  XNOR U50425 ( .A(n49791), .B(n49789), .Z(n50006) );
  AND U50426 ( .A(n50007), .B(n50008), .Z(n49789) );
  NANDN U50427 ( .A(n50009), .B(n50010), .Z(n50008) );
  OR U50428 ( .A(n50011), .B(n50012), .Z(n50010) );
  NAND U50429 ( .A(n50012), .B(n50011), .Z(n50007) );
  ANDN U50430 ( .B(A[18]), .A(n19), .Z(n49791) );
  XNOR U50431 ( .A(n49799), .B(n50013), .Z(n49792) );
  XNOR U50432 ( .A(n49798), .B(n49796), .Z(n50013) );
  AND U50433 ( .A(n50014), .B(n50015), .Z(n49796) );
  NANDN U50434 ( .A(n50016), .B(n50017), .Z(n50015) );
  NANDN U50435 ( .A(n50018), .B(n50019), .Z(n50017) );
  NANDN U50436 ( .A(n50019), .B(n50018), .Z(n50014) );
  ANDN U50437 ( .B(A[17]), .A(n17), .Z(n49798) );
  XNOR U50438 ( .A(n49806), .B(n50020), .Z(n49799) );
  XNOR U50439 ( .A(n49805), .B(n49803), .Z(n50020) );
  AND U50440 ( .A(n50021), .B(n50022), .Z(n49803) );
  NANDN U50441 ( .A(n50023), .B(n50024), .Z(n50022) );
  OR U50442 ( .A(n50025), .B(n50026), .Z(n50024) );
  NAND U50443 ( .A(n50026), .B(n50025), .Z(n50021) );
  ANDN U50444 ( .B(A[16]), .A(n15), .Z(n49805) );
  XNOR U50445 ( .A(n49813), .B(n50027), .Z(n49806) );
  XNOR U50446 ( .A(n49812), .B(n49810), .Z(n50027) );
  AND U50447 ( .A(n50028), .B(n50029), .Z(n49810) );
  NANDN U50448 ( .A(n50030), .B(n50031), .Z(n50029) );
  NANDN U50449 ( .A(n50032), .B(n50033), .Z(n50031) );
  NANDN U50450 ( .A(n50033), .B(n50032), .Z(n50028) );
  ANDN U50451 ( .B(A[15]), .A(n13), .Z(n49812) );
  XNOR U50452 ( .A(n49820), .B(n50034), .Z(n49813) );
  XNOR U50453 ( .A(n49819), .B(n49817), .Z(n50034) );
  AND U50454 ( .A(n50035), .B(n50036), .Z(n49817) );
  NANDN U50455 ( .A(n50037), .B(n50038), .Z(n50036) );
  OR U50456 ( .A(n50039), .B(n50040), .Z(n50038) );
  NAND U50457 ( .A(n50040), .B(n50039), .Z(n50035) );
  ANDN U50458 ( .B(A[14]), .A(n11), .Z(n49819) );
  XNOR U50459 ( .A(n49827), .B(n50041), .Z(n49820) );
  XNOR U50460 ( .A(n49826), .B(n49824), .Z(n50041) );
  AND U50461 ( .A(n50042), .B(n50043), .Z(n49824) );
  NANDN U50462 ( .A(n50044), .B(n50045), .Z(n50043) );
  NANDN U50463 ( .A(n50046), .B(n50047), .Z(n50045) );
  NANDN U50464 ( .A(n50047), .B(n50046), .Z(n50042) );
  ANDN U50465 ( .B(A[13]), .A(n9), .Z(n49826) );
  XNOR U50466 ( .A(n49834), .B(n50048), .Z(n49827) );
  XNOR U50467 ( .A(n49833), .B(n49831), .Z(n50048) );
  AND U50468 ( .A(n50049), .B(n50050), .Z(n49831) );
  NANDN U50469 ( .A(n50051), .B(n50052), .Z(n50050) );
  OR U50470 ( .A(n50053), .B(n50054), .Z(n50052) );
  NAND U50471 ( .A(n50054), .B(n50053), .Z(n50049) );
  ANDN U50472 ( .B(B[98]), .A(n73), .Z(n49833) );
  XNOR U50473 ( .A(n49841), .B(n50055), .Z(n49834) );
  XNOR U50474 ( .A(n49840), .B(n49838), .Z(n50055) );
  AND U50475 ( .A(n50056), .B(n50057), .Z(n49838) );
  NANDN U50476 ( .A(n50058), .B(n50059), .Z(n50057) );
  NANDN U50477 ( .A(n50060), .B(n50061), .Z(n50059) );
  NANDN U50478 ( .A(n50061), .B(n50060), .Z(n50056) );
  ANDN U50479 ( .B(A[11]), .A(n6), .Z(n49840) );
  XNOR U50480 ( .A(n49848), .B(n50062), .Z(n49841) );
  XNOR U50481 ( .A(n49847), .B(n49845), .Z(n50062) );
  AND U50482 ( .A(n50063), .B(n50064), .Z(n49845) );
  NANDN U50483 ( .A(n50065), .B(n50066), .Z(n50064) );
  OR U50484 ( .A(n50067), .B(n50068), .Z(n50066) );
  NAND U50485 ( .A(n50068), .B(n50067), .Z(n50063) );
  ANDN U50486 ( .B(A[10]), .A(n4), .Z(n49847) );
  XNOR U50487 ( .A(n49855), .B(n50069), .Z(n49848) );
  XNOR U50488 ( .A(n49854), .B(n49852), .Z(n50069) );
  AND U50489 ( .A(n50070), .B(n50071), .Z(n49852) );
  NANDN U50490 ( .A(n50072), .B(n50073), .Z(n50071) );
  NANDN U50491 ( .A(n50074), .B(n50075), .Z(n50073) );
  NANDN U50492 ( .A(n50075), .B(n50074), .Z(n50070) );
  ANDN U50493 ( .B(B[101]), .A(n76), .Z(n49854) );
  XNOR U50494 ( .A(n49862), .B(n50076), .Z(n49855) );
  XNOR U50495 ( .A(n49861), .B(n49859), .Z(n50076) );
  AND U50496 ( .A(n50077), .B(n50078), .Z(n49859) );
  NANDN U50497 ( .A(n50079), .B(n50080), .Z(n50078) );
  OR U50498 ( .A(n50081), .B(n50082), .Z(n50080) );
  NAND U50499 ( .A(n50082), .B(n50081), .Z(n50077) );
  ANDN U50500 ( .B(B[102]), .A(n77), .Z(n49861) );
  XNOR U50501 ( .A(n49869), .B(n50083), .Z(n49862) );
  XNOR U50502 ( .A(n49868), .B(n49866), .Z(n50083) );
  AND U50503 ( .A(n50084), .B(n50085), .Z(n49866) );
  NANDN U50504 ( .A(n50086), .B(n50087), .Z(n50085) );
  NANDN U50505 ( .A(n50088), .B(n50089), .Z(n50087) );
  NANDN U50506 ( .A(n50089), .B(n50088), .Z(n50084) );
  ANDN U50507 ( .B(B[103]), .A(n78), .Z(n49868) );
  XNOR U50508 ( .A(n49876), .B(n50090), .Z(n49869) );
  XNOR U50509 ( .A(n49875), .B(n49873), .Z(n50090) );
  AND U50510 ( .A(n50091), .B(n50092), .Z(n49873) );
  NANDN U50511 ( .A(n50093), .B(n50094), .Z(n50092) );
  OR U50512 ( .A(n50095), .B(n50096), .Z(n50094) );
  NAND U50513 ( .A(n50096), .B(n50095), .Z(n50091) );
  ANDN U50514 ( .B(B[104]), .A(n79), .Z(n49875) );
  XNOR U50515 ( .A(n49883), .B(n50097), .Z(n49876) );
  XNOR U50516 ( .A(n49882), .B(n49880), .Z(n50097) );
  AND U50517 ( .A(n50098), .B(n50099), .Z(n49880) );
  NANDN U50518 ( .A(n50100), .B(n50101), .Z(n50099) );
  NANDN U50519 ( .A(n50102), .B(n50103), .Z(n50101) );
  NANDN U50520 ( .A(n50103), .B(n50102), .Z(n50098) );
  ANDN U50521 ( .B(B[105]), .A(n80), .Z(n49882) );
  XNOR U50522 ( .A(n49890), .B(n50104), .Z(n49883) );
  XNOR U50523 ( .A(n49889), .B(n49887), .Z(n50104) );
  AND U50524 ( .A(n50105), .B(n50106), .Z(n49887) );
  NANDN U50525 ( .A(n50107), .B(n50108), .Z(n50106) );
  OR U50526 ( .A(n50109), .B(n50110), .Z(n50108) );
  NAND U50527 ( .A(n50110), .B(n50109), .Z(n50105) );
  ANDN U50528 ( .B(B[106]), .A(n81), .Z(n49889) );
  XNOR U50529 ( .A(n49897), .B(n50111), .Z(n49890) );
  XNOR U50530 ( .A(n49896), .B(n49894), .Z(n50111) );
  AND U50531 ( .A(n50112), .B(n50113), .Z(n49894) );
  NANDN U50532 ( .A(n50114), .B(n50115), .Z(n50113) );
  NAND U50533 ( .A(n50116), .B(n50117), .Z(n50115) );
  ANDN U50534 ( .B(B[107]), .A(n82), .Z(n49896) );
  XOR U50535 ( .A(n49903), .B(n50118), .Z(n49897) );
  XNOR U50536 ( .A(n49901), .B(n49904), .Z(n50118) );
  NAND U50537 ( .A(A[2]), .B(B[108]), .Z(n49904) );
  NANDN U50538 ( .A(n50119), .B(n50120), .Z(n49901) );
  AND U50539 ( .A(A[0]), .B(B[109]), .Z(n50120) );
  XNOR U50540 ( .A(n49906), .B(n50121), .Z(n49903) );
  NAND U50541 ( .A(A[0]), .B(B[110]), .Z(n50121) );
  NAND U50542 ( .A(B[109]), .B(A[1]), .Z(n49906) );
  NAND U50543 ( .A(n50122), .B(n50123), .Z(n576) );
  NANDN U50544 ( .A(n50124), .B(n50125), .Z(n50123) );
  OR U50545 ( .A(n50126), .B(n50127), .Z(n50125) );
  NAND U50546 ( .A(n50127), .B(n50126), .Z(n50122) );
  XOR U50547 ( .A(n578), .B(n577), .Z(\A1[107] ) );
  XOR U50548 ( .A(n50127), .B(n50128), .Z(n577) );
  XNOR U50549 ( .A(n50126), .B(n50124), .Z(n50128) );
  AND U50550 ( .A(n50129), .B(n50130), .Z(n50124) );
  NANDN U50551 ( .A(n50131), .B(n50132), .Z(n50130) );
  NANDN U50552 ( .A(n50133), .B(n50134), .Z(n50132) );
  NANDN U50553 ( .A(n50134), .B(n50133), .Z(n50129) );
  ANDN U50554 ( .B(B[78]), .A(n54), .Z(n50126) );
  XNOR U50555 ( .A(n49921), .B(n50135), .Z(n50127) );
  XNOR U50556 ( .A(n49920), .B(n49918), .Z(n50135) );
  AND U50557 ( .A(n50136), .B(n50137), .Z(n49918) );
  NANDN U50558 ( .A(n50138), .B(n50139), .Z(n50137) );
  OR U50559 ( .A(n50140), .B(n50141), .Z(n50139) );
  NAND U50560 ( .A(n50141), .B(n50140), .Z(n50136) );
  ANDN U50561 ( .B(B[79]), .A(n55), .Z(n49920) );
  XNOR U50562 ( .A(n49928), .B(n50142), .Z(n49921) );
  XNOR U50563 ( .A(n49927), .B(n49925), .Z(n50142) );
  AND U50564 ( .A(n50143), .B(n50144), .Z(n49925) );
  NANDN U50565 ( .A(n50145), .B(n50146), .Z(n50144) );
  NANDN U50566 ( .A(n50147), .B(n50148), .Z(n50146) );
  NANDN U50567 ( .A(n50148), .B(n50147), .Z(n50143) );
  ANDN U50568 ( .B(B[80]), .A(n56), .Z(n49927) );
  XNOR U50569 ( .A(n49935), .B(n50149), .Z(n49928) );
  XNOR U50570 ( .A(n49934), .B(n49932), .Z(n50149) );
  AND U50571 ( .A(n50150), .B(n50151), .Z(n49932) );
  NANDN U50572 ( .A(n50152), .B(n50153), .Z(n50151) );
  OR U50573 ( .A(n50154), .B(n50155), .Z(n50153) );
  NAND U50574 ( .A(n50155), .B(n50154), .Z(n50150) );
  ANDN U50575 ( .B(B[81]), .A(n57), .Z(n49934) );
  XNOR U50576 ( .A(n49942), .B(n50156), .Z(n49935) );
  XNOR U50577 ( .A(n49941), .B(n49939), .Z(n50156) );
  AND U50578 ( .A(n50157), .B(n50158), .Z(n49939) );
  NANDN U50579 ( .A(n50159), .B(n50160), .Z(n50158) );
  NANDN U50580 ( .A(n50161), .B(n50162), .Z(n50160) );
  NANDN U50581 ( .A(n50162), .B(n50161), .Z(n50157) );
  ANDN U50582 ( .B(B[82]), .A(n58), .Z(n49941) );
  XNOR U50583 ( .A(n49949), .B(n50163), .Z(n49942) );
  XNOR U50584 ( .A(n49948), .B(n49946), .Z(n50163) );
  AND U50585 ( .A(n50164), .B(n50165), .Z(n49946) );
  NANDN U50586 ( .A(n50166), .B(n50167), .Z(n50165) );
  OR U50587 ( .A(n50168), .B(n50169), .Z(n50167) );
  NAND U50588 ( .A(n50169), .B(n50168), .Z(n50164) );
  ANDN U50589 ( .B(B[83]), .A(n59), .Z(n49948) );
  XNOR U50590 ( .A(n49956), .B(n50170), .Z(n49949) );
  XNOR U50591 ( .A(n49955), .B(n49953), .Z(n50170) );
  AND U50592 ( .A(n50171), .B(n50172), .Z(n49953) );
  NANDN U50593 ( .A(n50173), .B(n50174), .Z(n50172) );
  NANDN U50594 ( .A(n50175), .B(n50176), .Z(n50174) );
  NANDN U50595 ( .A(n50176), .B(n50175), .Z(n50171) );
  ANDN U50596 ( .B(B[84]), .A(n60), .Z(n49955) );
  XNOR U50597 ( .A(n49963), .B(n50177), .Z(n49956) );
  XNOR U50598 ( .A(n49962), .B(n49960), .Z(n50177) );
  AND U50599 ( .A(n50178), .B(n50179), .Z(n49960) );
  NANDN U50600 ( .A(n50180), .B(n50181), .Z(n50179) );
  OR U50601 ( .A(n50182), .B(n50183), .Z(n50181) );
  NAND U50602 ( .A(n50183), .B(n50182), .Z(n50178) );
  ANDN U50603 ( .B(B[85]), .A(n61), .Z(n49962) );
  XNOR U50604 ( .A(n49970), .B(n50184), .Z(n49963) );
  XNOR U50605 ( .A(n49969), .B(n49967), .Z(n50184) );
  AND U50606 ( .A(n50185), .B(n50186), .Z(n49967) );
  NANDN U50607 ( .A(n50187), .B(n50188), .Z(n50186) );
  NANDN U50608 ( .A(n50189), .B(n50190), .Z(n50188) );
  NANDN U50609 ( .A(n50190), .B(n50189), .Z(n50185) );
  ANDN U50610 ( .B(B[86]), .A(n62), .Z(n49969) );
  XNOR U50611 ( .A(n49977), .B(n50191), .Z(n49970) );
  XNOR U50612 ( .A(n49976), .B(n49974), .Z(n50191) );
  AND U50613 ( .A(n50192), .B(n50193), .Z(n49974) );
  NANDN U50614 ( .A(n50194), .B(n50195), .Z(n50193) );
  OR U50615 ( .A(n50196), .B(n50197), .Z(n50195) );
  NAND U50616 ( .A(n50197), .B(n50196), .Z(n50192) );
  ANDN U50617 ( .B(B[87]), .A(n63), .Z(n49976) );
  XNOR U50618 ( .A(n49984), .B(n50198), .Z(n49977) );
  XNOR U50619 ( .A(n49983), .B(n49981), .Z(n50198) );
  AND U50620 ( .A(n50199), .B(n50200), .Z(n49981) );
  NANDN U50621 ( .A(n50201), .B(n50202), .Z(n50200) );
  NANDN U50622 ( .A(n50203), .B(n50204), .Z(n50202) );
  NANDN U50623 ( .A(n50204), .B(n50203), .Z(n50199) );
  ANDN U50624 ( .B(B[88]), .A(n64), .Z(n49983) );
  XNOR U50625 ( .A(n49991), .B(n50205), .Z(n49984) );
  XNOR U50626 ( .A(n49990), .B(n49988), .Z(n50205) );
  AND U50627 ( .A(n50206), .B(n50207), .Z(n49988) );
  NANDN U50628 ( .A(n50208), .B(n50209), .Z(n50207) );
  OR U50629 ( .A(n50210), .B(n50211), .Z(n50209) );
  NAND U50630 ( .A(n50211), .B(n50210), .Z(n50206) );
  ANDN U50631 ( .B(A[20]), .A(n25), .Z(n49990) );
  XNOR U50632 ( .A(n49998), .B(n50212), .Z(n49991) );
  XNOR U50633 ( .A(n49997), .B(n49995), .Z(n50212) );
  AND U50634 ( .A(n50213), .B(n50214), .Z(n49995) );
  NANDN U50635 ( .A(n50215), .B(n50216), .Z(n50214) );
  NANDN U50636 ( .A(n50217), .B(n50218), .Z(n50216) );
  NANDN U50637 ( .A(n50218), .B(n50217), .Z(n50213) );
  ANDN U50638 ( .B(A[19]), .A(n23), .Z(n49997) );
  XNOR U50639 ( .A(n50005), .B(n50219), .Z(n49998) );
  XNOR U50640 ( .A(n50004), .B(n50002), .Z(n50219) );
  AND U50641 ( .A(n50220), .B(n50221), .Z(n50002) );
  NANDN U50642 ( .A(n50222), .B(n50223), .Z(n50221) );
  OR U50643 ( .A(n50224), .B(n50225), .Z(n50223) );
  NAND U50644 ( .A(n50225), .B(n50224), .Z(n50220) );
  ANDN U50645 ( .B(A[18]), .A(n21), .Z(n50004) );
  XNOR U50646 ( .A(n50012), .B(n50226), .Z(n50005) );
  XNOR U50647 ( .A(n50011), .B(n50009), .Z(n50226) );
  AND U50648 ( .A(n50227), .B(n50228), .Z(n50009) );
  NANDN U50649 ( .A(n50229), .B(n50230), .Z(n50228) );
  NANDN U50650 ( .A(n50231), .B(n50232), .Z(n50230) );
  NANDN U50651 ( .A(n50232), .B(n50231), .Z(n50227) );
  ANDN U50652 ( .B(A[17]), .A(n19), .Z(n50011) );
  XNOR U50653 ( .A(n50019), .B(n50233), .Z(n50012) );
  XNOR U50654 ( .A(n50018), .B(n50016), .Z(n50233) );
  AND U50655 ( .A(n50234), .B(n50235), .Z(n50016) );
  NANDN U50656 ( .A(n50236), .B(n50237), .Z(n50235) );
  OR U50657 ( .A(n50238), .B(n50239), .Z(n50237) );
  NAND U50658 ( .A(n50239), .B(n50238), .Z(n50234) );
  ANDN U50659 ( .B(A[16]), .A(n17), .Z(n50018) );
  XNOR U50660 ( .A(n50026), .B(n50240), .Z(n50019) );
  XNOR U50661 ( .A(n50025), .B(n50023), .Z(n50240) );
  AND U50662 ( .A(n50241), .B(n50242), .Z(n50023) );
  NANDN U50663 ( .A(n50243), .B(n50244), .Z(n50242) );
  NANDN U50664 ( .A(n50245), .B(n50246), .Z(n50244) );
  NANDN U50665 ( .A(n50246), .B(n50245), .Z(n50241) );
  ANDN U50666 ( .B(A[15]), .A(n15), .Z(n50025) );
  XNOR U50667 ( .A(n50033), .B(n50247), .Z(n50026) );
  XNOR U50668 ( .A(n50032), .B(n50030), .Z(n50247) );
  AND U50669 ( .A(n50248), .B(n50249), .Z(n50030) );
  NANDN U50670 ( .A(n50250), .B(n50251), .Z(n50249) );
  OR U50671 ( .A(n50252), .B(n50253), .Z(n50251) );
  NAND U50672 ( .A(n50253), .B(n50252), .Z(n50248) );
  ANDN U50673 ( .B(A[14]), .A(n13), .Z(n50032) );
  XNOR U50674 ( .A(n50040), .B(n50254), .Z(n50033) );
  XNOR U50675 ( .A(n50039), .B(n50037), .Z(n50254) );
  AND U50676 ( .A(n50255), .B(n50256), .Z(n50037) );
  NANDN U50677 ( .A(n50257), .B(n50258), .Z(n50256) );
  NANDN U50678 ( .A(n50259), .B(n50260), .Z(n50258) );
  NANDN U50679 ( .A(n50260), .B(n50259), .Z(n50255) );
  ANDN U50680 ( .B(A[13]), .A(n11), .Z(n50039) );
  XNOR U50681 ( .A(n50047), .B(n50261), .Z(n50040) );
  XNOR U50682 ( .A(n50046), .B(n50044), .Z(n50261) );
  AND U50683 ( .A(n50262), .B(n50263), .Z(n50044) );
  NANDN U50684 ( .A(n50264), .B(n50265), .Z(n50263) );
  OR U50685 ( .A(n50266), .B(n50267), .Z(n50265) );
  NAND U50686 ( .A(n50267), .B(n50266), .Z(n50262) );
  ANDN U50687 ( .B(A[12]), .A(n9), .Z(n50046) );
  XNOR U50688 ( .A(n50054), .B(n50268), .Z(n50047) );
  XNOR U50689 ( .A(n50053), .B(n50051), .Z(n50268) );
  AND U50690 ( .A(n50269), .B(n50270), .Z(n50051) );
  NANDN U50691 ( .A(n50271), .B(n50272), .Z(n50270) );
  NANDN U50692 ( .A(n50273), .B(n50274), .Z(n50272) );
  NANDN U50693 ( .A(n50274), .B(n50273), .Z(n50269) );
  ANDN U50694 ( .B(B[98]), .A(n74), .Z(n50053) );
  XNOR U50695 ( .A(n50061), .B(n50275), .Z(n50054) );
  XNOR U50696 ( .A(n50060), .B(n50058), .Z(n50275) );
  AND U50697 ( .A(n50276), .B(n50277), .Z(n50058) );
  NANDN U50698 ( .A(n50278), .B(n50279), .Z(n50277) );
  OR U50699 ( .A(n50280), .B(n50281), .Z(n50279) );
  NAND U50700 ( .A(n50281), .B(n50280), .Z(n50276) );
  ANDN U50701 ( .B(A[10]), .A(n6), .Z(n50060) );
  XNOR U50702 ( .A(n50068), .B(n50282), .Z(n50061) );
  XNOR U50703 ( .A(n50067), .B(n50065), .Z(n50282) );
  AND U50704 ( .A(n50283), .B(n50284), .Z(n50065) );
  NANDN U50705 ( .A(n50285), .B(n50286), .Z(n50284) );
  NANDN U50706 ( .A(n50287), .B(n50288), .Z(n50286) );
  NANDN U50707 ( .A(n50288), .B(n50287), .Z(n50283) );
  ANDN U50708 ( .B(A[9]), .A(n4), .Z(n50067) );
  XNOR U50709 ( .A(n50075), .B(n50289), .Z(n50068) );
  XNOR U50710 ( .A(n50074), .B(n50072), .Z(n50289) );
  AND U50711 ( .A(n50290), .B(n50291), .Z(n50072) );
  NANDN U50712 ( .A(n50292), .B(n50293), .Z(n50291) );
  OR U50713 ( .A(n50294), .B(n50295), .Z(n50293) );
  NAND U50714 ( .A(n50295), .B(n50294), .Z(n50290) );
  ANDN U50715 ( .B(B[101]), .A(n77), .Z(n50074) );
  XNOR U50716 ( .A(n50082), .B(n50296), .Z(n50075) );
  XNOR U50717 ( .A(n50081), .B(n50079), .Z(n50296) );
  AND U50718 ( .A(n50297), .B(n50298), .Z(n50079) );
  NANDN U50719 ( .A(n50299), .B(n50300), .Z(n50298) );
  NANDN U50720 ( .A(n50301), .B(n50302), .Z(n50300) );
  NANDN U50721 ( .A(n50302), .B(n50301), .Z(n50297) );
  ANDN U50722 ( .B(B[102]), .A(n78), .Z(n50081) );
  XNOR U50723 ( .A(n50089), .B(n50303), .Z(n50082) );
  XNOR U50724 ( .A(n50088), .B(n50086), .Z(n50303) );
  AND U50725 ( .A(n50304), .B(n50305), .Z(n50086) );
  NANDN U50726 ( .A(n50306), .B(n50307), .Z(n50305) );
  OR U50727 ( .A(n50308), .B(n50309), .Z(n50307) );
  NAND U50728 ( .A(n50309), .B(n50308), .Z(n50304) );
  ANDN U50729 ( .B(B[103]), .A(n79), .Z(n50088) );
  XNOR U50730 ( .A(n50096), .B(n50310), .Z(n50089) );
  XNOR U50731 ( .A(n50095), .B(n50093), .Z(n50310) );
  AND U50732 ( .A(n50311), .B(n50312), .Z(n50093) );
  NANDN U50733 ( .A(n50313), .B(n50314), .Z(n50312) );
  NANDN U50734 ( .A(n50315), .B(n50316), .Z(n50314) );
  NANDN U50735 ( .A(n50316), .B(n50315), .Z(n50311) );
  ANDN U50736 ( .B(B[104]), .A(n80), .Z(n50095) );
  XNOR U50737 ( .A(n50103), .B(n50317), .Z(n50096) );
  XNOR U50738 ( .A(n50102), .B(n50100), .Z(n50317) );
  AND U50739 ( .A(n50318), .B(n50319), .Z(n50100) );
  NANDN U50740 ( .A(n50320), .B(n50321), .Z(n50319) );
  OR U50741 ( .A(n50322), .B(n50323), .Z(n50321) );
  NAND U50742 ( .A(n50323), .B(n50322), .Z(n50318) );
  ANDN U50743 ( .B(B[105]), .A(n81), .Z(n50102) );
  XNOR U50744 ( .A(n50110), .B(n50324), .Z(n50103) );
  XNOR U50745 ( .A(n50109), .B(n50107), .Z(n50324) );
  AND U50746 ( .A(n50325), .B(n50326), .Z(n50107) );
  NANDN U50747 ( .A(n50327), .B(n50328), .Z(n50326) );
  NAND U50748 ( .A(n50329), .B(n50330), .Z(n50328) );
  ANDN U50749 ( .B(B[106]), .A(n82), .Z(n50109) );
  XOR U50750 ( .A(n50116), .B(n50331), .Z(n50110) );
  XNOR U50751 ( .A(n50114), .B(n50117), .Z(n50331) );
  NAND U50752 ( .A(A[2]), .B(B[107]), .Z(n50117) );
  NANDN U50753 ( .A(n50332), .B(n50333), .Z(n50114) );
  AND U50754 ( .A(A[0]), .B(B[108]), .Z(n50333) );
  XNOR U50755 ( .A(n50119), .B(n50334), .Z(n50116) );
  NAND U50756 ( .A(A[0]), .B(B[109]), .Z(n50334) );
  NAND U50757 ( .A(B[108]), .B(A[1]), .Z(n50119) );
  NAND U50758 ( .A(n50335), .B(n50336), .Z(n578) );
  NANDN U50759 ( .A(n50337), .B(n50338), .Z(n50336) );
  OR U50760 ( .A(n50339), .B(n50340), .Z(n50338) );
  NAND U50761 ( .A(n50340), .B(n50339), .Z(n50335) );
  XOR U50762 ( .A(n580), .B(n579), .Z(\A1[106] ) );
  XOR U50763 ( .A(n50340), .B(n50341), .Z(n579) );
  XNOR U50764 ( .A(n50339), .B(n50337), .Z(n50341) );
  AND U50765 ( .A(n50342), .B(n50343), .Z(n50337) );
  NANDN U50766 ( .A(n50344), .B(n50345), .Z(n50343) );
  NANDN U50767 ( .A(n50346), .B(n50347), .Z(n50345) );
  NANDN U50768 ( .A(n50347), .B(n50346), .Z(n50342) );
  ANDN U50769 ( .B(B[77]), .A(n54), .Z(n50339) );
  XNOR U50770 ( .A(n50134), .B(n50348), .Z(n50340) );
  XNOR U50771 ( .A(n50133), .B(n50131), .Z(n50348) );
  AND U50772 ( .A(n50349), .B(n50350), .Z(n50131) );
  NANDN U50773 ( .A(n50351), .B(n50352), .Z(n50350) );
  OR U50774 ( .A(n50353), .B(n50354), .Z(n50352) );
  NAND U50775 ( .A(n50354), .B(n50353), .Z(n50349) );
  ANDN U50776 ( .B(B[78]), .A(n55), .Z(n50133) );
  XNOR U50777 ( .A(n50141), .B(n50355), .Z(n50134) );
  XNOR U50778 ( .A(n50140), .B(n50138), .Z(n50355) );
  AND U50779 ( .A(n50356), .B(n50357), .Z(n50138) );
  NANDN U50780 ( .A(n50358), .B(n50359), .Z(n50357) );
  NANDN U50781 ( .A(n50360), .B(n50361), .Z(n50359) );
  NANDN U50782 ( .A(n50361), .B(n50360), .Z(n50356) );
  ANDN U50783 ( .B(B[79]), .A(n56), .Z(n50140) );
  XNOR U50784 ( .A(n50148), .B(n50362), .Z(n50141) );
  XNOR U50785 ( .A(n50147), .B(n50145), .Z(n50362) );
  AND U50786 ( .A(n50363), .B(n50364), .Z(n50145) );
  NANDN U50787 ( .A(n50365), .B(n50366), .Z(n50364) );
  OR U50788 ( .A(n50367), .B(n50368), .Z(n50366) );
  NAND U50789 ( .A(n50368), .B(n50367), .Z(n50363) );
  ANDN U50790 ( .B(B[80]), .A(n57), .Z(n50147) );
  XNOR U50791 ( .A(n50155), .B(n50369), .Z(n50148) );
  XNOR U50792 ( .A(n50154), .B(n50152), .Z(n50369) );
  AND U50793 ( .A(n50370), .B(n50371), .Z(n50152) );
  NANDN U50794 ( .A(n50372), .B(n50373), .Z(n50371) );
  NANDN U50795 ( .A(n50374), .B(n50375), .Z(n50373) );
  NANDN U50796 ( .A(n50375), .B(n50374), .Z(n50370) );
  ANDN U50797 ( .B(B[81]), .A(n58), .Z(n50154) );
  XNOR U50798 ( .A(n50162), .B(n50376), .Z(n50155) );
  XNOR U50799 ( .A(n50161), .B(n50159), .Z(n50376) );
  AND U50800 ( .A(n50377), .B(n50378), .Z(n50159) );
  NANDN U50801 ( .A(n50379), .B(n50380), .Z(n50378) );
  OR U50802 ( .A(n50381), .B(n50382), .Z(n50380) );
  NAND U50803 ( .A(n50382), .B(n50381), .Z(n50377) );
  ANDN U50804 ( .B(B[82]), .A(n59), .Z(n50161) );
  XNOR U50805 ( .A(n50169), .B(n50383), .Z(n50162) );
  XNOR U50806 ( .A(n50168), .B(n50166), .Z(n50383) );
  AND U50807 ( .A(n50384), .B(n50385), .Z(n50166) );
  NANDN U50808 ( .A(n50386), .B(n50387), .Z(n50385) );
  NANDN U50809 ( .A(n50388), .B(n50389), .Z(n50387) );
  NANDN U50810 ( .A(n50389), .B(n50388), .Z(n50384) );
  ANDN U50811 ( .B(B[83]), .A(n60), .Z(n50168) );
  XNOR U50812 ( .A(n50176), .B(n50390), .Z(n50169) );
  XNOR U50813 ( .A(n50175), .B(n50173), .Z(n50390) );
  AND U50814 ( .A(n50391), .B(n50392), .Z(n50173) );
  NANDN U50815 ( .A(n50393), .B(n50394), .Z(n50392) );
  OR U50816 ( .A(n50395), .B(n50396), .Z(n50394) );
  NAND U50817 ( .A(n50396), .B(n50395), .Z(n50391) );
  ANDN U50818 ( .B(B[84]), .A(n61), .Z(n50175) );
  XNOR U50819 ( .A(n50183), .B(n50397), .Z(n50176) );
  XNOR U50820 ( .A(n50182), .B(n50180), .Z(n50397) );
  AND U50821 ( .A(n50398), .B(n50399), .Z(n50180) );
  NANDN U50822 ( .A(n50400), .B(n50401), .Z(n50399) );
  NANDN U50823 ( .A(n50402), .B(n50403), .Z(n50401) );
  NANDN U50824 ( .A(n50403), .B(n50402), .Z(n50398) );
  ANDN U50825 ( .B(B[85]), .A(n62), .Z(n50182) );
  XNOR U50826 ( .A(n50190), .B(n50404), .Z(n50183) );
  XNOR U50827 ( .A(n50189), .B(n50187), .Z(n50404) );
  AND U50828 ( .A(n50405), .B(n50406), .Z(n50187) );
  NANDN U50829 ( .A(n50407), .B(n50408), .Z(n50406) );
  OR U50830 ( .A(n50409), .B(n50410), .Z(n50408) );
  NAND U50831 ( .A(n50410), .B(n50409), .Z(n50405) );
  ANDN U50832 ( .B(B[86]), .A(n63), .Z(n50189) );
  XNOR U50833 ( .A(n50197), .B(n50411), .Z(n50190) );
  XNOR U50834 ( .A(n50196), .B(n50194), .Z(n50411) );
  AND U50835 ( .A(n50412), .B(n50413), .Z(n50194) );
  NANDN U50836 ( .A(n50414), .B(n50415), .Z(n50413) );
  NANDN U50837 ( .A(n50416), .B(n50417), .Z(n50415) );
  NANDN U50838 ( .A(n50417), .B(n50416), .Z(n50412) );
  ANDN U50839 ( .B(B[87]), .A(n64), .Z(n50196) );
  XNOR U50840 ( .A(n50204), .B(n50418), .Z(n50197) );
  XNOR U50841 ( .A(n50203), .B(n50201), .Z(n50418) );
  AND U50842 ( .A(n50419), .B(n50420), .Z(n50201) );
  NANDN U50843 ( .A(n50421), .B(n50422), .Z(n50420) );
  OR U50844 ( .A(n50423), .B(n50424), .Z(n50422) );
  NAND U50845 ( .A(n50424), .B(n50423), .Z(n50419) );
  ANDN U50846 ( .B(A[20]), .A(n27), .Z(n50203) );
  XNOR U50847 ( .A(n50211), .B(n50425), .Z(n50204) );
  XNOR U50848 ( .A(n50210), .B(n50208), .Z(n50425) );
  AND U50849 ( .A(n50426), .B(n50427), .Z(n50208) );
  NANDN U50850 ( .A(n50428), .B(n50429), .Z(n50427) );
  NANDN U50851 ( .A(n50430), .B(n50431), .Z(n50429) );
  NANDN U50852 ( .A(n50431), .B(n50430), .Z(n50426) );
  ANDN U50853 ( .B(A[19]), .A(n25), .Z(n50210) );
  XNOR U50854 ( .A(n50218), .B(n50432), .Z(n50211) );
  XNOR U50855 ( .A(n50217), .B(n50215), .Z(n50432) );
  AND U50856 ( .A(n50433), .B(n50434), .Z(n50215) );
  NANDN U50857 ( .A(n50435), .B(n50436), .Z(n50434) );
  OR U50858 ( .A(n50437), .B(n50438), .Z(n50436) );
  NAND U50859 ( .A(n50438), .B(n50437), .Z(n50433) );
  ANDN U50860 ( .B(A[18]), .A(n23), .Z(n50217) );
  XNOR U50861 ( .A(n50225), .B(n50439), .Z(n50218) );
  XNOR U50862 ( .A(n50224), .B(n50222), .Z(n50439) );
  AND U50863 ( .A(n50440), .B(n50441), .Z(n50222) );
  NANDN U50864 ( .A(n50442), .B(n50443), .Z(n50441) );
  NANDN U50865 ( .A(n50444), .B(n50445), .Z(n50443) );
  NANDN U50866 ( .A(n50445), .B(n50444), .Z(n50440) );
  ANDN U50867 ( .B(A[17]), .A(n21), .Z(n50224) );
  XNOR U50868 ( .A(n50232), .B(n50446), .Z(n50225) );
  XNOR U50869 ( .A(n50231), .B(n50229), .Z(n50446) );
  AND U50870 ( .A(n50447), .B(n50448), .Z(n50229) );
  NANDN U50871 ( .A(n50449), .B(n50450), .Z(n50448) );
  OR U50872 ( .A(n50451), .B(n50452), .Z(n50450) );
  NAND U50873 ( .A(n50452), .B(n50451), .Z(n50447) );
  ANDN U50874 ( .B(A[16]), .A(n19), .Z(n50231) );
  XNOR U50875 ( .A(n50239), .B(n50453), .Z(n50232) );
  XNOR U50876 ( .A(n50238), .B(n50236), .Z(n50453) );
  AND U50877 ( .A(n50454), .B(n50455), .Z(n50236) );
  NANDN U50878 ( .A(n50456), .B(n50457), .Z(n50455) );
  NANDN U50879 ( .A(n50458), .B(n50459), .Z(n50457) );
  NANDN U50880 ( .A(n50459), .B(n50458), .Z(n50454) );
  ANDN U50881 ( .B(A[15]), .A(n17), .Z(n50238) );
  XNOR U50882 ( .A(n50246), .B(n50460), .Z(n50239) );
  XNOR U50883 ( .A(n50245), .B(n50243), .Z(n50460) );
  AND U50884 ( .A(n50461), .B(n50462), .Z(n50243) );
  NANDN U50885 ( .A(n50463), .B(n50464), .Z(n50462) );
  OR U50886 ( .A(n50465), .B(n50466), .Z(n50464) );
  NAND U50887 ( .A(n50466), .B(n50465), .Z(n50461) );
  ANDN U50888 ( .B(A[14]), .A(n15), .Z(n50245) );
  XNOR U50889 ( .A(n50253), .B(n50467), .Z(n50246) );
  XNOR U50890 ( .A(n50252), .B(n50250), .Z(n50467) );
  AND U50891 ( .A(n50468), .B(n50469), .Z(n50250) );
  NANDN U50892 ( .A(n50470), .B(n50471), .Z(n50469) );
  NANDN U50893 ( .A(n50472), .B(n50473), .Z(n50471) );
  NANDN U50894 ( .A(n50473), .B(n50472), .Z(n50468) );
  ANDN U50895 ( .B(A[13]), .A(n13), .Z(n50252) );
  XNOR U50896 ( .A(n50260), .B(n50474), .Z(n50253) );
  XNOR U50897 ( .A(n50259), .B(n50257), .Z(n50474) );
  AND U50898 ( .A(n50475), .B(n50476), .Z(n50257) );
  NANDN U50899 ( .A(n50477), .B(n50478), .Z(n50476) );
  OR U50900 ( .A(n50479), .B(n50480), .Z(n50478) );
  NAND U50901 ( .A(n50480), .B(n50479), .Z(n50475) );
  ANDN U50902 ( .B(A[12]), .A(n11), .Z(n50259) );
  XNOR U50903 ( .A(n50267), .B(n50481), .Z(n50260) );
  XNOR U50904 ( .A(n50266), .B(n50264), .Z(n50481) );
  AND U50905 ( .A(n50482), .B(n50483), .Z(n50264) );
  NANDN U50906 ( .A(n50484), .B(n50485), .Z(n50483) );
  NANDN U50907 ( .A(n50486), .B(n50487), .Z(n50485) );
  NANDN U50908 ( .A(n50487), .B(n50486), .Z(n50482) );
  ANDN U50909 ( .B(A[11]), .A(n9), .Z(n50266) );
  XNOR U50910 ( .A(n50274), .B(n50488), .Z(n50267) );
  XNOR U50911 ( .A(n50273), .B(n50271), .Z(n50488) );
  AND U50912 ( .A(n50489), .B(n50490), .Z(n50271) );
  NANDN U50913 ( .A(n50491), .B(n50492), .Z(n50490) );
  OR U50914 ( .A(n50493), .B(n50494), .Z(n50492) );
  NAND U50915 ( .A(n50494), .B(n50493), .Z(n50489) );
  ANDN U50916 ( .B(B[98]), .A(n75), .Z(n50273) );
  XNOR U50917 ( .A(n50281), .B(n50495), .Z(n50274) );
  XNOR U50918 ( .A(n50280), .B(n50278), .Z(n50495) );
  AND U50919 ( .A(n50496), .B(n50497), .Z(n50278) );
  NANDN U50920 ( .A(n50498), .B(n50499), .Z(n50497) );
  NANDN U50921 ( .A(n50500), .B(n50501), .Z(n50499) );
  NANDN U50922 ( .A(n50501), .B(n50500), .Z(n50496) );
  ANDN U50923 ( .B(A[9]), .A(n6), .Z(n50280) );
  XNOR U50924 ( .A(n50288), .B(n50502), .Z(n50281) );
  XNOR U50925 ( .A(n50287), .B(n50285), .Z(n50502) );
  AND U50926 ( .A(n50503), .B(n50504), .Z(n50285) );
  NANDN U50927 ( .A(n50505), .B(n50506), .Z(n50504) );
  OR U50928 ( .A(n50507), .B(n50508), .Z(n50506) );
  NAND U50929 ( .A(n50508), .B(n50507), .Z(n50503) );
  ANDN U50930 ( .B(A[8]), .A(n4), .Z(n50287) );
  XNOR U50931 ( .A(n50295), .B(n50509), .Z(n50288) );
  XNOR U50932 ( .A(n50294), .B(n50292), .Z(n50509) );
  AND U50933 ( .A(n50510), .B(n50511), .Z(n50292) );
  NANDN U50934 ( .A(n50512), .B(n50513), .Z(n50511) );
  NANDN U50935 ( .A(n50514), .B(n50515), .Z(n50513) );
  NANDN U50936 ( .A(n50515), .B(n50514), .Z(n50510) );
  ANDN U50937 ( .B(B[101]), .A(n78), .Z(n50294) );
  XNOR U50938 ( .A(n50302), .B(n50516), .Z(n50295) );
  XNOR U50939 ( .A(n50301), .B(n50299), .Z(n50516) );
  AND U50940 ( .A(n50517), .B(n50518), .Z(n50299) );
  NANDN U50941 ( .A(n50519), .B(n50520), .Z(n50518) );
  OR U50942 ( .A(n50521), .B(n50522), .Z(n50520) );
  NAND U50943 ( .A(n50522), .B(n50521), .Z(n50517) );
  ANDN U50944 ( .B(B[102]), .A(n79), .Z(n50301) );
  XNOR U50945 ( .A(n50309), .B(n50523), .Z(n50302) );
  XNOR U50946 ( .A(n50308), .B(n50306), .Z(n50523) );
  AND U50947 ( .A(n50524), .B(n50525), .Z(n50306) );
  NANDN U50948 ( .A(n50526), .B(n50527), .Z(n50525) );
  NANDN U50949 ( .A(n50528), .B(n50529), .Z(n50527) );
  NANDN U50950 ( .A(n50529), .B(n50528), .Z(n50524) );
  ANDN U50951 ( .B(B[103]), .A(n80), .Z(n50308) );
  XNOR U50952 ( .A(n50316), .B(n50530), .Z(n50309) );
  XNOR U50953 ( .A(n50315), .B(n50313), .Z(n50530) );
  AND U50954 ( .A(n50531), .B(n50532), .Z(n50313) );
  NANDN U50955 ( .A(n50533), .B(n50534), .Z(n50532) );
  OR U50956 ( .A(n50535), .B(n50536), .Z(n50534) );
  NAND U50957 ( .A(n50536), .B(n50535), .Z(n50531) );
  ANDN U50958 ( .B(B[104]), .A(n81), .Z(n50315) );
  XNOR U50959 ( .A(n50323), .B(n50537), .Z(n50316) );
  XNOR U50960 ( .A(n50322), .B(n50320), .Z(n50537) );
  AND U50961 ( .A(n50538), .B(n50539), .Z(n50320) );
  NANDN U50962 ( .A(n50540), .B(n50541), .Z(n50539) );
  NAND U50963 ( .A(n50542), .B(n50543), .Z(n50541) );
  ANDN U50964 ( .B(B[105]), .A(n82), .Z(n50322) );
  XOR U50965 ( .A(n50329), .B(n50544), .Z(n50323) );
  XNOR U50966 ( .A(n50327), .B(n50330), .Z(n50544) );
  NAND U50967 ( .A(A[2]), .B(B[106]), .Z(n50330) );
  NANDN U50968 ( .A(n50545), .B(n50546), .Z(n50327) );
  AND U50969 ( .A(A[0]), .B(B[107]), .Z(n50546) );
  XNOR U50970 ( .A(n50332), .B(n50547), .Z(n50329) );
  NAND U50971 ( .A(A[0]), .B(B[108]), .Z(n50547) );
  NAND U50972 ( .A(B[107]), .B(A[1]), .Z(n50332) );
  NAND U50973 ( .A(n50548), .B(n50549), .Z(n580) );
  NANDN U50974 ( .A(n50550), .B(n50551), .Z(n50549) );
  OR U50975 ( .A(n50552), .B(n50553), .Z(n50551) );
  NAND U50976 ( .A(n50553), .B(n50552), .Z(n50548) );
  XOR U50977 ( .A(n582), .B(n581), .Z(\A1[105] ) );
  XOR U50978 ( .A(n50553), .B(n50554), .Z(n581) );
  XNOR U50979 ( .A(n50552), .B(n50550), .Z(n50554) );
  AND U50980 ( .A(n50555), .B(n50556), .Z(n50550) );
  NANDN U50981 ( .A(n50557), .B(n50558), .Z(n50556) );
  NANDN U50982 ( .A(n50559), .B(n50560), .Z(n50558) );
  NANDN U50983 ( .A(n50560), .B(n50559), .Z(n50555) );
  ANDN U50984 ( .B(B[76]), .A(n54), .Z(n50552) );
  XNOR U50985 ( .A(n50347), .B(n50561), .Z(n50553) );
  XNOR U50986 ( .A(n50346), .B(n50344), .Z(n50561) );
  AND U50987 ( .A(n50562), .B(n50563), .Z(n50344) );
  NANDN U50988 ( .A(n50564), .B(n50565), .Z(n50563) );
  OR U50989 ( .A(n50566), .B(n50567), .Z(n50565) );
  NAND U50990 ( .A(n50567), .B(n50566), .Z(n50562) );
  ANDN U50991 ( .B(B[77]), .A(n55), .Z(n50346) );
  XNOR U50992 ( .A(n50354), .B(n50568), .Z(n50347) );
  XNOR U50993 ( .A(n50353), .B(n50351), .Z(n50568) );
  AND U50994 ( .A(n50569), .B(n50570), .Z(n50351) );
  NANDN U50995 ( .A(n50571), .B(n50572), .Z(n50570) );
  NANDN U50996 ( .A(n50573), .B(n50574), .Z(n50572) );
  NANDN U50997 ( .A(n50574), .B(n50573), .Z(n50569) );
  ANDN U50998 ( .B(B[78]), .A(n56), .Z(n50353) );
  XNOR U50999 ( .A(n50361), .B(n50575), .Z(n50354) );
  XNOR U51000 ( .A(n50360), .B(n50358), .Z(n50575) );
  AND U51001 ( .A(n50576), .B(n50577), .Z(n50358) );
  NANDN U51002 ( .A(n50578), .B(n50579), .Z(n50577) );
  OR U51003 ( .A(n50580), .B(n50581), .Z(n50579) );
  NAND U51004 ( .A(n50581), .B(n50580), .Z(n50576) );
  ANDN U51005 ( .B(B[79]), .A(n57), .Z(n50360) );
  XNOR U51006 ( .A(n50368), .B(n50582), .Z(n50361) );
  XNOR U51007 ( .A(n50367), .B(n50365), .Z(n50582) );
  AND U51008 ( .A(n50583), .B(n50584), .Z(n50365) );
  NANDN U51009 ( .A(n50585), .B(n50586), .Z(n50584) );
  NANDN U51010 ( .A(n50587), .B(n50588), .Z(n50586) );
  NANDN U51011 ( .A(n50588), .B(n50587), .Z(n50583) );
  ANDN U51012 ( .B(B[80]), .A(n58), .Z(n50367) );
  XNOR U51013 ( .A(n50375), .B(n50589), .Z(n50368) );
  XNOR U51014 ( .A(n50374), .B(n50372), .Z(n50589) );
  AND U51015 ( .A(n50590), .B(n50591), .Z(n50372) );
  NANDN U51016 ( .A(n50592), .B(n50593), .Z(n50591) );
  OR U51017 ( .A(n50594), .B(n50595), .Z(n50593) );
  NAND U51018 ( .A(n50595), .B(n50594), .Z(n50590) );
  ANDN U51019 ( .B(B[81]), .A(n59), .Z(n50374) );
  XNOR U51020 ( .A(n50382), .B(n50596), .Z(n50375) );
  XNOR U51021 ( .A(n50381), .B(n50379), .Z(n50596) );
  AND U51022 ( .A(n50597), .B(n50598), .Z(n50379) );
  NANDN U51023 ( .A(n50599), .B(n50600), .Z(n50598) );
  NANDN U51024 ( .A(n50601), .B(n50602), .Z(n50600) );
  NANDN U51025 ( .A(n50602), .B(n50601), .Z(n50597) );
  ANDN U51026 ( .B(B[82]), .A(n60), .Z(n50381) );
  XNOR U51027 ( .A(n50389), .B(n50603), .Z(n50382) );
  XNOR U51028 ( .A(n50388), .B(n50386), .Z(n50603) );
  AND U51029 ( .A(n50604), .B(n50605), .Z(n50386) );
  NANDN U51030 ( .A(n50606), .B(n50607), .Z(n50605) );
  OR U51031 ( .A(n50608), .B(n50609), .Z(n50607) );
  NAND U51032 ( .A(n50609), .B(n50608), .Z(n50604) );
  ANDN U51033 ( .B(B[83]), .A(n61), .Z(n50388) );
  XNOR U51034 ( .A(n50396), .B(n50610), .Z(n50389) );
  XNOR U51035 ( .A(n50395), .B(n50393), .Z(n50610) );
  AND U51036 ( .A(n50611), .B(n50612), .Z(n50393) );
  NANDN U51037 ( .A(n50613), .B(n50614), .Z(n50612) );
  NANDN U51038 ( .A(n50615), .B(n50616), .Z(n50614) );
  NANDN U51039 ( .A(n50616), .B(n50615), .Z(n50611) );
  ANDN U51040 ( .B(B[84]), .A(n62), .Z(n50395) );
  XNOR U51041 ( .A(n50403), .B(n50617), .Z(n50396) );
  XNOR U51042 ( .A(n50402), .B(n50400), .Z(n50617) );
  AND U51043 ( .A(n50618), .B(n50619), .Z(n50400) );
  NANDN U51044 ( .A(n50620), .B(n50621), .Z(n50619) );
  OR U51045 ( .A(n50622), .B(n50623), .Z(n50621) );
  NAND U51046 ( .A(n50623), .B(n50622), .Z(n50618) );
  ANDN U51047 ( .B(B[85]), .A(n63), .Z(n50402) );
  XNOR U51048 ( .A(n50410), .B(n50624), .Z(n50403) );
  XNOR U51049 ( .A(n50409), .B(n50407), .Z(n50624) );
  AND U51050 ( .A(n50625), .B(n50626), .Z(n50407) );
  NANDN U51051 ( .A(n50627), .B(n50628), .Z(n50626) );
  NANDN U51052 ( .A(n50629), .B(n50630), .Z(n50628) );
  NANDN U51053 ( .A(n50630), .B(n50629), .Z(n50625) );
  ANDN U51054 ( .B(B[86]), .A(n64), .Z(n50409) );
  XNOR U51055 ( .A(n50417), .B(n50631), .Z(n50410) );
  XNOR U51056 ( .A(n50416), .B(n50414), .Z(n50631) );
  AND U51057 ( .A(n50632), .B(n50633), .Z(n50414) );
  NANDN U51058 ( .A(n50634), .B(n50635), .Z(n50633) );
  OR U51059 ( .A(n50636), .B(n50637), .Z(n50635) );
  NAND U51060 ( .A(n50637), .B(n50636), .Z(n50632) );
  ANDN U51061 ( .B(B[87]), .A(n65), .Z(n50416) );
  XNOR U51062 ( .A(n50424), .B(n50638), .Z(n50417) );
  XNOR U51063 ( .A(n50423), .B(n50421), .Z(n50638) );
  AND U51064 ( .A(n50639), .B(n50640), .Z(n50421) );
  NANDN U51065 ( .A(n50641), .B(n50642), .Z(n50640) );
  NANDN U51066 ( .A(n50643), .B(n50644), .Z(n50642) );
  NANDN U51067 ( .A(n50644), .B(n50643), .Z(n50639) );
  ANDN U51068 ( .B(A[19]), .A(n27), .Z(n50423) );
  XNOR U51069 ( .A(n50431), .B(n50645), .Z(n50424) );
  XNOR U51070 ( .A(n50430), .B(n50428), .Z(n50645) );
  AND U51071 ( .A(n50646), .B(n50647), .Z(n50428) );
  NANDN U51072 ( .A(n50648), .B(n50649), .Z(n50647) );
  OR U51073 ( .A(n50650), .B(n50651), .Z(n50649) );
  NAND U51074 ( .A(n50651), .B(n50650), .Z(n50646) );
  ANDN U51075 ( .B(A[18]), .A(n25), .Z(n50430) );
  XNOR U51076 ( .A(n50438), .B(n50652), .Z(n50431) );
  XNOR U51077 ( .A(n50437), .B(n50435), .Z(n50652) );
  AND U51078 ( .A(n50653), .B(n50654), .Z(n50435) );
  NANDN U51079 ( .A(n50655), .B(n50656), .Z(n50654) );
  NANDN U51080 ( .A(n50657), .B(n50658), .Z(n50656) );
  NANDN U51081 ( .A(n50658), .B(n50657), .Z(n50653) );
  ANDN U51082 ( .B(A[17]), .A(n23), .Z(n50437) );
  XNOR U51083 ( .A(n50445), .B(n50659), .Z(n50438) );
  XNOR U51084 ( .A(n50444), .B(n50442), .Z(n50659) );
  AND U51085 ( .A(n50660), .B(n50661), .Z(n50442) );
  NANDN U51086 ( .A(n50662), .B(n50663), .Z(n50661) );
  OR U51087 ( .A(n50664), .B(n50665), .Z(n50663) );
  NAND U51088 ( .A(n50665), .B(n50664), .Z(n50660) );
  ANDN U51089 ( .B(A[16]), .A(n21), .Z(n50444) );
  XNOR U51090 ( .A(n50452), .B(n50666), .Z(n50445) );
  XNOR U51091 ( .A(n50451), .B(n50449), .Z(n50666) );
  AND U51092 ( .A(n50667), .B(n50668), .Z(n50449) );
  NANDN U51093 ( .A(n50669), .B(n50670), .Z(n50668) );
  NANDN U51094 ( .A(n50671), .B(n50672), .Z(n50670) );
  NANDN U51095 ( .A(n50672), .B(n50671), .Z(n50667) );
  ANDN U51096 ( .B(A[15]), .A(n19), .Z(n50451) );
  XNOR U51097 ( .A(n50459), .B(n50673), .Z(n50452) );
  XNOR U51098 ( .A(n50458), .B(n50456), .Z(n50673) );
  AND U51099 ( .A(n50674), .B(n50675), .Z(n50456) );
  NANDN U51100 ( .A(n50676), .B(n50677), .Z(n50675) );
  OR U51101 ( .A(n50678), .B(n50679), .Z(n50677) );
  NAND U51102 ( .A(n50679), .B(n50678), .Z(n50674) );
  ANDN U51103 ( .B(A[14]), .A(n17), .Z(n50458) );
  XNOR U51104 ( .A(n50466), .B(n50680), .Z(n50459) );
  XNOR U51105 ( .A(n50465), .B(n50463), .Z(n50680) );
  AND U51106 ( .A(n50681), .B(n50682), .Z(n50463) );
  NANDN U51107 ( .A(n50683), .B(n50684), .Z(n50682) );
  NANDN U51108 ( .A(n50685), .B(n50686), .Z(n50684) );
  NANDN U51109 ( .A(n50686), .B(n50685), .Z(n50681) );
  ANDN U51110 ( .B(A[13]), .A(n15), .Z(n50465) );
  XNOR U51111 ( .A(n50473), .B(n50687), .Z(n50466) );
  XNOR U51112 ( .A(n50472), .B(n50470), .Z(n50687) );
  AND U51113 ( .A(n50688), .B(n50689), .Z(n50470) );
  NANDN U51114 ( .A(n50690), .B(n50691), .Z(n50689) );
  OR U51115 ( .A(n50692), .B(n50693), .Z(n50691) );
  NAND U51116 ( .A(n50693), .B(n50692), .Z(n50688) );
  ANDN U51117 ( .B(A[12]), .A(n13), .Z(n50472) );
  XNOR U51118 ( .A(n50480), .B(n50694), .Z(n50473) );
  XNOR U51119 ( .A(n50479), .B(n50477), .Z(n50694) );
  AND U51120 ( .A(n50695), .B(n50696), .Z(n50477) );
  NANDN U51121 ( .A(n50697), .B(n50698), .Z(n50696) );
  NANDN U51122 ( .A(n50699), .B(n50700), .Z(n50698) );
  NANDN U51123 ( .A(n50700), .B(n50699), .Z(n50695) );
  ANDN U51124 ( .B(A[11]), .A(n11), .Z(n50479) );
  XNOR U51125 ( .A(n50487), .B(n50701), .Z(n50480) );
  XNOR U51126 ( .A(n50486), .B(n50484), .Z(n50701) );
  AND U51127 ( .A(n50702), .B(n50703), .Z(n50484) );
  NANDN U51128 ( .A(n50704), .B(n50705), .Z(n50703) );
  OR U51129 ( .A(n50706), .B(n50707), .Z(n50705) );
  NAND U51130 ( .A(n50707), .B(n50706), .Z(n50702) );
  ANDN U51131 ( .B(A[10]), .A(n9), .Z(n50486) );
  XNOR U51132 ( .A(n50494), .B(n50708), .Z(n50487) );
  XNOR U51133 ( .A(n50493), .B(n50491), .Z(n50708) );
  AND U51134 ( .A(n50709), .B(n50710), .Z(n50491) );
  NANDN U51135 ( .A(n50711), .B(n50712), .Z(n50710) );
  NANDN U51136 ( .A(n50713), .B(n50714), .Z(n50712) );
  NANDN U51137 ( .A(n50714), .B(n50713), .Z(n50709) );
  ANDN U51138 ( .B(B[98]), .A(n76), .Z(n50493) );
  XNOR U51139 ( .A(n50501), .B(n50715), .Z(n50494) );
  XNOR U51140 ( .A(n50500), .B(n50498), .Z(n50715) );
  AND U51141 ( .A(n50716), .B(n50717), .Z(n50498) );
  NANDN U51142 ( .A(n50718), .B(n50719), .Z(n50717) );
  OR U51143 ( .A(n50720), .B(n50721), .Z(n50719) );
  NAND U51144 ( .A(n50721), .B(n50720), .Z(n50716) );
  ANDN U51145 ( .B(A[8]), .A(n6), .Z(n50500) );
  XNOR U51146 ( .A(n50508), .B(n50722), .Z(n50501) );
  XNOR U51147 ( .A(n50507), .B(n50505), .Z(n50722) );
  AND U51148 ( .A(n50723), .B(n50724), .Z(n50505) );
  NANDN U51149 ( .A(n50725), .B(n50726), .Z(n50724) );
  NANDN U51150 ( .A(n50727), .B(n50728), .Z(n50726) );
  NANDN U51151 ( .A(n50728), .B(n50727), .Z(n50723) );
  ANDN U51152 ( .B(A[7]), .A(n4), .Z(n50507) );
  XNOR U51153 ( .A(n50515), .B(n50729), .Z(n50508) );
  XNOR U51154 ( .A(n50514), .B(n50512), .Z(n50729) );
  AND U51155 ( .A(n50730), .B(n50731), .Z(n50512) );
  NANDN U51156 ( .A(n50732), .B(n50733), .Z(n50731) );
  OR U51157 ( .A(n50734), .B(n50735), .Z(n50733) );
  NAND U51158 ( .A(n50735), .B(n50734), .Z(n50730) );
  ANDN U51159 ( .B(B[101]), .A(n79), .Z(n50514) );
  XNOR U51160 ( .A(n50522), .B(n50736), .Z(n50515) );
  XNOR U51161 ( .A(n50521), .B(n50519), .Z(n50736) );
  AND U51162 ( .A(n50737), .B(n50738), .Z(n50519) );
  NANDN U51163 ( .A(n50739), .B(n50740), .Z(n50738) );
  NANDN U51164 ( .A(n50741), .B(n50742), .Z(n50740) );
  NANDN U51165 ( .A(n50742), .B(n50741), .Z(n50737) );
  ANDN U51166 ( .B(B[102]), .A(n80), .Z(n50521) );
  XNOR U51167 ( .A(n50529), .B(n50743), .Z(n50522) );
  XNOR U51168 ( .A(n50528), .B(n50526), .Z(n50743) );
  AND U51169 ( .A(n50744), .B(n50745), .Z(n50526) );
  NANDN U51170 ( .A(n50746), .B(n50747), .Z(n50745) );
  OR U51171 ( .A(n50748), .B(n50749), .Z(n50747) );
  NAND U51172 ( .A(n50749), .B(n50748), .Z(n50744) );
  ANDN U51173 ( .B(B[103]), .A(n81), .Z(n50528) );
  XNOR U51174 ( .A(n50536), .B(n50750), .Z(n50529) );
  XNOR U51175 ( .A(n50535), .B(n50533), .Z(n50750) );
  AND U51176 ( .A(n50751), .B(n50752), .Z(n50533) );
  NANDN U51177 ( .A(n50753), .B(n50754), .Z(n50752) );
  NAND U51178 ( .A(n50755), .B(n50756), .Z(n50754) );
  ANDN U51179 ( .B(B[104]), .A(n82), .Z(n50535) );
  XOR U51180 ( .A(n50542), .B(n50757), .Z(n50536) );
  XNOR U51181 ( .A(n50540), .B(n50543), .Z(n50757) );
  NAND U51182 ( .A(A[2]), .B(B[105]), .Z(n50543) );
  NANDN U51183 ( .A(n50758), .B(n50759), .Z(n50540) );
  AND U51184 ( .A(A[0]), .B(B[106]), .Z(n50759) );
  XNOR U51185 ( .A(n50545), .B(n50760), .Z(n50542) );
  NAND U51186 ( .A(A[0]), .B(B[107]), .Z(n50760) );
  NAND U51187 ( .A(B[106]), .B(A[1]), .Z(n50545) );
  NAND U51188 ( .A(n50761), .B(n50762), .Z(n582) );
  NANDN U51189 ( .A(n50763), .B(n50764), .Z(n50762) );
  OR U51190 ( .A(n50765), .B(n50766), .Z(n50764) );
  NAND U51191 ( .A(n50766), .B(n50765), .Z(n50761) );
  XOR U51192 ( .A(n584), .B(n583), .Z(\A1[104] ) );
  XOR U51193 ( .A(n50766), .B(n50767), .Z(n583) );
  XNOR U51194 ( .A(n50765), .B(n50763), .Z(n50767) );
  AND U51195 ( .A(n50768), .B(n50769), .Z(n50763) );
  NANDN U51196 ( .A(n50770), .B(n50771), .Z(n50769) );
  NANDN U51197 ( .A(n50772), .B(n50773), .Z(n50771) );
  NANDN U51198 ( .A(n50773), .B(n50772), .Z(n50768) );
  ANDN U51199 ( .B(B[75]), .A(n54), .Z(n50765) );
  XNOR U51200 ( .A(n50560), .B(n50774), .Z(n50766) );
  XNOR U51201 ( .A(n50559), .B(n50557), .Z(n50774) );
  AND U51202 ( .A(n50775), .B(n50776), .Z(n50557) );
  NANDN U51203 ( .A(n50777), .B(n50778), .Z(n50776) );
  OR U51204 ( .A(n50779), .B(n50780), .Z(n50778) );
  NAND U51205 ( .A(n50780), .B(n50779), .Z(n50775) );
  ANDN U51206 ( .B(B[76]), .A(n55), .Z(n50559) );
  XNOR U51207 ( .A(n50567), .B(n50781), .Z(n50560) );
  XNOR U51208 ( .A(n50566), .B(n50564), .Z(n50781) );
  AND U51209 ( .A(n50782), .B(n50783), .Z(n50564) );
  NANDN U51210 ( .A(n50784), .B(n50785), .Z(n50783) );
  NANDN U51211 ( .A(n50786), .B(n50787), .Z(n50785) );
  NANDN U51212 ( .A(n50787), .B(n50786), .Z(n50782) );
  ANDN U51213 ( .B(B[77]), .A(n56), .Z(n50566) );
  XNOR U51214 ( .A(n50574), .B(n50788), .Z(n50567) );
  XNOR U51215 ( .A(n50573), .B(n50571), .Z(n50788) );
  AND U51216 ( .A(n50789), .B(n50790), .Z(n50571) );
  NANDN U51217 ( .A(n50791), .B(n50792), .Z(n50790) );
  OR U51218 ( .A(n50793), .B(n50794), .Z(n50792) );
  NAND U51219 ( .A(n50794), .B(n50793), .Z(n50789) );
  ANDN U51220 ( .B(B[78]), .A(n57), .Z(n50573) );
  XNOR U51221 ( .A(n50581), .B(n50795), .Z(n50574) );
  XNOR U51222 ( .A(n50580), .B(n50578), .Z(n50795) );
  AND U51223 ( .A(n50796), .B(n50797), .Z(n50578) );
  NANDN U51224 ( .A(n50798), .B(n50799), .Z(n50797) );
  NANDN U51225 ( .A(n50800), .B(n50801), .Z(n50799) );
  NANDN U51226 ( .A(n50801), .B(n50800), .Z(n50796) );
  ANDN U51227 ( .B(B[79]), .A(n58), .Z(n50580) );
  XNOR U51228 ( .A(n50588), .B(n50802), .Z(n50581) );
  XNOR U51229 ( .A(n50587), .B(n50585), .Z(n50802) );
  AND U51230 ( .A(n50803), .B(n50804), .Z(n50585) );
  NANDN U51231 ( .A(n50805), .B(n50806), .Z(n50804) );
  OR U51232 ( .A(n50807), .B(n50808), .Z(n50806) );
  NAND U51233 ( .A(n50808), .B(n50807), .Z(n50803) );
  ANDN U51234 ( .B(B[80]), .A(n59), .Z(n50587) );
  XNOR U51235 ( .A(n50595), .B(n50809), .Z(n50588) );
  XNOR U51236 ( .A(n50594), .B(n50592), .Z(n50809) );
  AND U51237 ( .A(n50810), .B(n50811), .Z(n50592) );
  NANDN U51238 ( .A(n50812), .B(n50813), .Z(n50811) );
  NANDN U51239 ( .A(n50814), .B(n50815), .Z(n50813) );
  NANDN U51240 ( .A(n50815), .B(n50814), .Z(n50810) );
  ANDN U51241 ( .B(B[81]), .A(n60), .Z(n50594) );
  XNOR U51242 ( .A(n50602), .B(n50816), .Z(n50595) );
  XNOR U51243 ( .A(n50601), .B(n50599), .Z(n50816) );
  AND U51244 ( .A(n50817), .B(n50818), .Z(n50599) );
  NANDN U51245 ( .A(n50819), .B(n50820), .Z(n50818) );
  OR U51246 ( .A(n50821), .B(n50822), .Z(n50820) );
  NAND U51247 ( .A(n50822), .B(n50821), .Z(n50817) );
  ANDN U51248 ( .B(B[82]), .A(n61), .Z(n50601) );
  XNOR U51249 ( .A(n50609), .B(n50823), .Z(n50602) );
  XNOR U51250 ( .A(n50608), .B(n50606), .Z(n50823) );
  AND U51251 ( .A(n50824), .B(n50825), .Z(n50606) );
  NANDN U51252 ( .A(n50826), .B(n50827), .Z(n50825) );
  NANDN U51253 ( .A(n50828), .B(n50829), .Z(n50827) );
  NANDN U51254 ( .A(n50829), .B(n50828), .Z(n50824) );
  ANDN U51255 ( .B(B[83]), .A(n62), .Z(n50608) );
  XNOR U51256 ( .A(n50616), .B(n50830), .Z(n50609) );
  XNOR U51257 ( .A(n50615), .B(n50613), .Z(n50830) );
  AND U51258 ( .A(n50831), .B(n50832), .Z(n50613) );
  NANDN U51259 ( .A(n50833), .B(n50834), .Z(n50832) );
  OR U51260 ( .A(n50835), .B(n50836), .Z(n50834) );
  NAND U51261 ( .A(n50836), .B(n50835), .Z(n50831) );
  ANDN U51262 ( .B(B[84]), .A(n63), .Z(n50615) );
  XNOR U51263 ( .A(n50623), .B(n50837), .Z(n50616) );
  XNOR U51264 ( .A(n50622), .B(n50620), .Z(n50837) );
  AND U51265 ( .A(n50838), .B(n50839), .Z(n50620) );
  NANDN U51266 ( .A(n50840), .B(n50841), .Z(n50839) );
  NANDN U51267 ( .A(n50842), .B(n50843), .Z(n50841) );
  NANDN U51268 ( .A(n50843), .B(n50842), .Z(n50838) );
  ANDN U51269 ( .B(B[85]), .A(n64), .Z(n50622) );
  XNOR U51270 ( .A(n50630), .B(n50844), .Z(n50623) );
  XNOR U51271 ( .A(n50629), .B(n50627), .Z(n50844) );
  AND U51272 ( .A(n50845), .B(n50846), .Z(n50627) );
  NANDN U51273 ( .A(n50847), .B(n50848), .Z(n50846) );
  OR U51274 ( .A(n50849), .B(n50850), .Z(n50848) );
  NAND U51275 ( .A(n50850), .B(n50849), .Z(n50845) );
  ANDN U51276 ( .B(B[86]), .A(n65), .Z(n50629) );
  XNOR U51277 ( .A(n50637), .B(n50851), .Z(n50630) );
  XNOR U51278 ( .A(n50636), .B(n50634), .Z(n50851) );
  AND U51279 ( .A(n50852), .B(n50853), .Z(n50634) );
  NANDN U51280 ( .A(n50854), .B(n50855), .Z(n50853) );
  NANDN U51281 ( .A(n50856), .B(n50857), .Z(n50855) );
  NANDN U51282 ( .A(n50857), .B(n50856), .Z(n50852) );
  ANDN U51283 ( .B(A[19]), .A(n29), .Z(n50636) );
  XNOR U51284 ( .A(n50644), .B(n50858), .Z(n50637) );
  XNOR U51285 ( .A(n50643), .B(n50641), .Z(n50858) );
  AND U51286 ( .A(n50859), .B(n50860), .Z(n50641) );
  NANDN U51287 ( .A(n50861), .B(n50862), .Z(n50860) );
  OR U51288 ( .A(n50863), .B(n50864), .Z(n50862) );
  NAND U51289 ( .A(n50864), .B(n50863), .Z(n50859) );
  ANDN U51290 ( .B(A[18]), .A(n27), .Z(n50643) );
  XNOR U51291 ( .A(n50651), .B(n50865), .Z(n50644) );
  XNOR U51292 ( .A(n50650), .B(n50648), .Z(n50865) );
  AND U51293 ( .A(n50866), .B(n50867), .Z(n50648) );
  NANDN U51294 ( .A(n50868), .B(n50869), .Z(n50867) );
  NANDN U51295 ( .A(n50870), .B(n50871), .Z(n50869) );
  NANDN U51296 ( .A(n50871), .B(n50870), .Z(n50866) );
  ANDN U51297 ( .B(A[17]), .A(n25), .Z(n50650) );
  XNOR U51298 ( .A(n50658), .B(n50872), .Z(n50651) );
  XNOR U51299 ( .A(n50657), .B(n50655), .Z(n50872) );
  AND U51300 ( .A(n50873), .B(n50874), .Z(n50655) );
  NANDN U51301 ( .A(n50875), .B(n50876), .Z(n50874) );
  OR U51302 ( .A(n50877), .B(n50878), .Z(n50876) );
  NAND U51303 ( .A(n50878), .B(n50877), .Z(n50873) );
  ANDN U51304 ( .B(A[16]), .A(n23), .Z(n50657) );
  XNOR U51305 ( .A(n50665), .B(n50879), .Z(n50658) );
  XNOR U51306 ( .A(n50664), .B(n50662), .Z(n50879) );
  AND U51307 ( .A(n50880), .B(n50881), .Z(n50662) );
  NANDN U51308 ( .A(n50882), .B(n50883), .Z(n50881) );
  NANDN U51309 ( .A(n50884), .B(n50885), .Z(n50883) );
  NANDN U51310 ( .A(n50885), .B(n50884), .Z(n50880) );
  ANDN U51311 ( .B(A[15]), .A(n21), .Z(n50664) );
  XNOR U51312 ( .A(n50672), .B(n50886), .Z(n50665) );
  XNOR U51313 ( .A(n50671), .B(n50669), .Z(n50886) );
  AND U51314 ( .A(n50887), .B(n50888), .Z(n50669) );
  NANDN U51315 ( .A(n50889), .B(n50890), .Z(n50888) );
  OR U51316 ( .A(n50891), .B(n50892), .Z(n50890) );
  NAND U51317 ( .A(n50892), .B(n50891), .Z(n50887) );
  ANDN U51318 ( .B(A[14]), .A(n19), .Z(n50671) );
  XNOR U51319 ( .A(n50679), .B(n50893), .Z(n50672) );
  XNOR U51320 ( .A(n50678), .B(n50676), .Z(n50893) );
  AND U51321 ( .A(n50894), .B(n50895), .Z(n50676) );
  NANDN U51322 ( .A(n50896), .B(n50897), .Z(n50895) );
  NANDN U51323 ( .A(n50898), .B(n50899), .Z(n50897) );
  NANDN U51324 ( .A(n50899), .B(n50898), .Z(n50894) );
  ANDN U51325 ( .B(A[13]), .A(n17), .Z(n50678) );
  XNOR U51326 ( .A(n50686), .B(n50900), .Z(n50679) );
  XNOR U51327 ( .A(n50685), .B(n50683), .Z(n50900) );
  AND U51328 ( .A(n50901), .B(n50902), .Z(n50683) );
  NANDN U51329 ( .A(n50903), .B(n50904), .Z(n50902) );
  OR U51330 ( .A(n50905), .B(n50906), .Z(n50904) );
  NAND U51331 ( .A(n50906), .B(n50905), .Z(n50901) );
  ANDN U51332 ( .B(A[12]), .A(n15), .Z(n50685) );
  XNOR U51333 ( .A(n50693), .B(n50907), .Z(n50686) );
  XNOR U51334 ( .A(n50692), .B(n50690), .Z(n50907) );
  AND U51335 ( .A(n50908), .B(n50909), .Z(n50690) );
  NANDN U51336 ( .A(n50910), .B(n50911), .Z(n50909) );
  NANDN U51337 ( .A(n50912), .B(n50913), .Z(n50911) );
  NANDN U51338 ( .A(n50913), .B(n50912), .Z(n50908) );
  ANDN U51339 ( .B(A[11]), .A(n13), .Z(n50692) );
  XNOR U51340 ( .A(n50700), .B(n50914), .Z(n50693) );
  XNOR U51341 ( .A(n50699), .B(n50697), .Z(n50914) );
  AND U51342 ( .A(n50915), .B(n50916), .Z(n50697) );
  NANDN U51343 ( .A(n50917), .B(n50918), .Z(n50916) );
  OR U51344 ( .A(n50919), .B(n50920), .Z(n50918) );
  NAND U51345 ( .A(n50920), .B(n50919), .Z(n50915) );
  ANDN U51346 ( .B(A[10]), .A(n11), .Z(n50699) );
  XNOR U51347 ( .A(n50707), .B(n50921), .Z(n50700) );
  XNOR U51348 ( .A(n50706), .B(n50704), .Z(n50921) );
  AND U51349 ( .A(n50922), .B(n50923), .Z(n50704) );
  NANDN U51350 ( .A(n50924), .B(n50925), .Z(n50923) );
  NANDN U51351 ( .A(n50926), .B(n50927), .Z(n50925) );
  NANDN U51352 ( .A(n50927), .B(n50926), .Z(n50922) );
  ANDN U51353 ( .B(A[9]), .A(n9), .Z(n50706) );
  XNOR U51354 ( .A(n50714), .B(n50928), .Z(n50707) );
  XNOR U51355 ( .A(n50713), .B(n50711), .Z(n50928) );
  AND U51356 ( .A(n50929), .B(n50930), .Z(n50711) );
  NANDN U51357 ( .A(n50931), .B(n50932), .Z(n50930) );
  OR U51358 ( .A(n50933), .B(n50934), .Z(n50932) );
  NAND U51359 ( .A(n50934), .B(n50933), .Z(n50929) );
  ANDN U51360 ( .B(B[98]), .A(n77), .Z(n50713) );
  XNOR U51361 ( .A(n50721), .B(n50935), .Z(n50714) );
  XNOR U51362 ( .A(n50720), .B(n50718), .Z(n50935) );
  AND U51363 ( .A(n50936), .B(n50937), .Z(n50718) );
  NANDN U51364 ( .A(n50938), .B(n50939), .Z(n50937) );
  NANDN U51365 ( .A(n50940), .B(n50941), .Z(n50939) );
  NANDN U51366 ( .A(n50941), .B(n50940), .Z(n50936) );
  ANDN U51367 ( .B(A[7]), .A(n6), .Z(n50720) );
  XNOR U51368 ( .A(n50728), .B(n50942), .Z(n50721) );
  XNOR U51369 ( .A(n50727), .B(n50725), .Z(n50942) );
  AND U51370 ( .A(n50943), .B(n50944), .Z(n50725) );
  NANDN U51371 ( .A(n50945), .B(n50946), .Z(n50944) );
  OR U51372 ( .A(n50947), .B(n50948), .Z(n50946) );
  NAND U51373 ( .A(n50948), .B(n50947), .Z(n50943) );
  ANDN U51374 ( .B(A[6]), .A(n4), .Z(n50727) );
  XNOR U51375 ( .A(n50735), .B(n50949), .Z(n50728) );
  XNOR U51376 ( .A(n50734), .B(n50732), .Z(n50949) );
  AND U51377 ( .A(n50950), .B(n50951), .Z(n50732) );
  NANDN U51378 ( .A(n50952), .B(n50953), .Z(n50951) );
  NANDN U51379 ( .A(n50954), .B(n50955), .Z(n50953) );
  NANDN U51380 ( .A(n50955), .B(n50954), .Z(n50950) );
  ANDN U51381 ( .B(B[101]), .A(n80), .Z(n50734) );
  XNOR U51382 ( .A(n50742), .B(n50956), .Z(n50735) );
  XNOR U51383 ( .A(n50741), .B(n50739), .Z(n50956) );
  AND U51384 ( .A(n50957), .B(n50958), .Z(n50739) );
  NANDN U51385 ( .A(n50959), .B(n50960), .Z(n50958) );
  OR U51386 ( .A(n50961), .B(n50962), .Z(n50960) );
  NAND U51387 ( .A(n50962), .B(n50961), .Z(n50957) );
  ANDN U51388 ( .B(B[102]), .A(n81), .Z(n50741) );
  XNOR U51389 ( .A(n50749), .B(n50963), .Z(n50742) );
  XNOR U51390 ( .A(n50748), .B(n50746), .Z(n50963) );
  AND U51391 ( .A(n50964), .B(n50965), .Z(n50746) );
  NANDN U51392 ( .A(n50966), .B(n50967), .Z(n50965) );
  NAND U51393 ( .A(n50968), .B(n50969), .Z(n50967) );
  ANDN U51394 ( .B(B[103]), .A(n82), .Z(n50748) );
  XOR U51395 ( .A(n50755), .B(n50970), .Z(n50749) );
  XNOR U51396 ( .A(n50753), .B(n50756), .Z(n50970) );
  NAND U51397 ( .A(A[2]), .B(B[104]), .Z(n50756) );
  NANDN U51398 ( .A(n50971), .B(n50972), .Z(n50753) );
  AND U51399 ( .A(A[0]), .B(B[105]), .Z(n50972) );
  XNOR U51400 ( .A(n50758), .B(n50973), .Z(n50755) );
  NAND U51401 ( .A(A[0]), .B(B[106]), .Z(n50973) );
  NAND U51402 ( .A(B[105]), .B(A[1]), .Z(n50758) );
  NAND U51403 ( .A(n50974), .B(n50975), .Z(n584) );
  NANDN U51404 ( .A(n50976), .B(n50977), .Z(n50975) );
  OR U51405 ( .A(n50978), .B(n50979), .Z(n50977) );
  NAND U51406 ( .A(n50979), .B(n50978), .Z(n50974) );
  XOR U51407 ( .A(n586), .B(n585), .Z(\A1[103] ) );
  XOR U51408 ( .A(n50979), .B(n50980), .Z(n585) );
  XNOR U51409 ( .A(n50978), .B(n50976), .Z(n50980) );
  AND U51410 ( .A(n50981), .B(n50982), .Z(n50976) );
  NANDN U51411 ( .A(n50983), .B(n50984), .Z(n50982) );
  NANDN U51412 ( .A(n50985), .B(n50986), .Z(n50984) );
  NANDN U51413 ( .A(n50986), .B(n50985), .Z(n50981) );
  ANDN U51414 ( .B(B[74]), .A(n54), .Z(n50978) );
  XNOR U51415 ( .A(n50773), .B(n50987), .Z(n50979) );
  XNOR U51416 ( .A(n50772), .B(n50770), .Z(n50987) );
  AND U51417 ( .A(n50988), .B(n50989), .Z(n50770) );
  NANDN U51418 ( .A(n50990), .B(n50991), .Z(n50989) );
  OR U51419 ( .A(n50992), .B(n50993), .Z(n50991) );
  NAND U51420 ( .A(n50993), .B(n50992), .Z(n50988) );
  ANDN U51421 ( .B(B[75]), .A(n55), .Z(n50772) );
  XNOR U51422 ( .A(n50780), .B(n50994), .Z(n50773) );
  XNOR U51423 ( .A(n50779), .B(n50777), .Z(n50994) );
  AND U51424 ( .A(n50995), .B(n50996), .Z(n50777) );
  NANDN U51425 ( .A(n50997), .B(n50998), .Z(n50996) );
  NANDN U51426 ( .A(n50999), .B(n51000), .Z(n50998) );
  NANDN U51427 ( .A(n51000), .B(n50999), .Z(n50995) );
  ANDN U51428 ( .B(B[76]), .A(n56), .Z(n50779) );
  XNOR U51429 ( .A(n50787), .B(n51001), .Z(n50780) );
  XNOR U51430 ( .A(n50786), .B(n50784), .Z(n51001) );
  AND U51431 ( .A(n51002), .B(n51003), .Z(n50784) );
  NANDN U51432 ( .A(n51004), .B(n51005), .Z(n51003) );
  OR U51433 ( .A(n51006), .B(n51007), .Z(n51005) );
  NAND U51434 ( .A(n51007), .B(n51006), .Z(n51002) );
  ANDN U51435 ( .B(B[77]), .A(n57), .Z(n50786) );
  XNOR U51436 ( .A(n50794), .B(n51008), .Z(n50787) );
  XNOR U51437 ( .A(n50793), .B(n50791), .Z(n51008) );
  AND U51438 ( .A(n51009), .B(n51010), .Z(n50791) );
  NANDN U51439 ( .A(n51011), .B(n51012), .Z(n51010) );
  NANDN U51440 ( .A(n51013), .B(n51014), .Z(n51012) );
  NANDN U51441 ( .A(n51014), .B(n51013), .Z(n51009) );
  ANDN U51442 ( .B(B[78]), .A(n58), .Z(n50793) );
  XNOR U51443 ( .A(n50801), .B(n51015), .Z(n50794) );
  XNOR U51444 ( .A(n50800), .B(n50798), .Z(n51015) );
  AND U51445 ( .A(n51016), .B(n51017), .Z(n50798) );
  NANDN U51446 ( .A(n51018), .B(n51019), .Z(n51017) );
  OR U51447 ( .A(n51020), .B(n51021), .Z(n51019) );
  NAND U51448 ( .A(n51021), .B(n51020), .Z(n51016) );
  ANDN U51449 ( .B(B[79]), .A(n59), .Z(n50800) );
  XNOR U51450 ( .A(n50808), .B(n51022), .Z(n50801) );
  XNOR U51451 ( .A(n50807), .B(n50805), .Z(n51022) );
  AND U51452 ( .A(n51023), .B(n51024), .Z(n50805) );
  NANDN U51453 ( .A(n51025), .B(n51026), .Z(n51024) );
  NANDN U51454 ( .A(n51027), .B(n51028), .Z(n51026) );
  NANDN U51455 ( .A(n51028), .B(n51027), .Z(n51023) );
  ANDN U51456 ( .B(B[80]), .A(n60), .Z(n50807) );
  XNOR U51457 ( .A(n50815), .B(n51029), .Z(n50808) );
  XNOR U51458 ( .A(n50814), .B(n50812), .Z(n51029) );
  AND U51459 ( .A(n51030), .B(n51031), .Z(n50812) );
  NANDN U51460 ( .A(n51032), .B(n51033), .Z(n51031) );
  OR U51461 ( .A(n51034), .B(n51035), .Z(n51033) );
  NAND U51462 ( .A(n51035), .B(n51034), .Z(n51030) );
  ANDN U51463 ( .B(B[81]), .A(n61), .Z(n50814) );
  XNOR U51464 ( .A(n50822), .B(n51036), .Z(n50815) );
  XNOR U51465 ( .A(n50821), .B(n50819), .Z(n51036) );
  AND U51466 ( .A(n51037), .B(n51038), .Z(n50819) );
  NANDN U51467 ( .A(n51039), .B(n51040), .Z(n51038) );
  NANDN U51468 ( .A(n51041), .B(n51042), .Z(n51040) );
  NANDN U51469 ( .A(n51042), .B(n51041), .Z(n51037) );
  ANDN U51470 ( .B(B[82]), .A(n62), .Z(n50821) );
  XNOR U51471 ( .A(n50829), .B(n51043), .Z(n50822) );
  XNOR U51472 ( .A(n50828), .B(n50826), .Z(n51043) );
  AND U51473 ( .A(n51044), .B(n51045), .Z(n50826) );
  NANDN U51474 ( .A(n51046), .B(n51047), .Z(n51045) );
  OR U51475 ( .A(n51048), .B(n51049), .Z(n51047) );
  NAND U51476 ( .A(n51049), .B(n51048), .Z(n51044) );
  ANDN U51477 ( .B(B[83]), .A(n63), .Z(n50828) );
  XNOR U51478 ( .A(n50836), .B(n51050), .Z(n50829) );
  XNOR U51479 ( .A(n50835), .B(n50833), .Z(n51050) );
  AND U51480 ( .A(n51051), .B(n51052), .Z(n50833) );
  NANDN U51481 ( .A(n51053), .B(n51054), .Z(n51052) );
  NANDN U51482 ( .A(n51055), .B(n51056), .Z(n51054) );
  NANDN U51483 ( .A(n51056), .B(n51055), .Z(n51051) );
  ANDN U51484 ( .B(B[84]), .A(n64), .Z(n50835) );
  XNOR U51485 ( .A(n50843), .B(n51057), .Z(n50836) );
  XNOR U51486 ( .A(n50842), .B(n50840), .Z(n51057) );
  AND U51487 ( .A(n51058), .B(n51059), .Z(n50840) );
  NANDN U51488 ( .A(n51060), .B(n51061), .Z(n51059) );
  OR U51489 ( .A(n51062), .B(n51063), .Z(n51061) );
  NAND U51490 ( .A(n51063), .B(n51062), .Z(n51058) );
  ANDN U51491 ( .B(B[85]), .A(n65), .Z(n50842) );
  XNOR U51492 ( .A(n50850), .B(n51064), .Z(n50843) );
  XNOR U51493 ( .A(n50849), .B(n50847), .Z(n51064) );
  AND U51494 ( .A(n51065), .B(n51066), .Z(n50847) );
  NANDN U51495 ( .A(n51067), .B(n51068), .Z(n51066) );
  NANDN U51496 ( .A(n51069), .B(n51070), .Z(n51068) );
  NANDN U51497 ( .A(n51070), .B(n51069), .Z(n51065) );
  ANDN U51498 ( .B(B[86]), .A(n66), .Z(n50849) );
  XNOR U51499 ( .A(n50857), .B(n51071), .Z(n50850) );
  XNOR U51500 ( .A(n50856), .B(n50854), .Z(n51071) );
  AND U51501 ( .A(n51072), .B(n51073), .Z(n50854) );
  NANDN U51502 ( .A(n51074), .B(n51075), .Z(n51073) );
  OR U51503 ( .A(n51076), .B(n51077), .Z(n51075) );
  NAND U51504 ( .A(n51077), .B(n51076), .Z(n51072) );
  ANDN U51505 ( .B(A[18]), .A(n29), .Z(n50856) );
  XNOR U51506 ( .A(n50864), .B(n51078), .Z(n50857) );
  XNOR U51507 ( .A(n50863), .B(n50861), .Z(n51078) );
  AND U51508 ( .A(n51079), .B(n51080), .Z(n50861) );
  NANDN U51509 ( .A(n51081), .B(n51082), .Z(n51080) );
  NANDN U51510 ( .A(n51083), .B(n51084), .Z(n51082) );
  NANDN U51511 ( .A(n51084), .B(n51083), .Z(n51079) );
  ANDN U51512 ( .B(A[17]), .A(n27), .Z(n50863) );
  XNOR U51513 ( .A(n50871), .B(n51085), .Z(n50864) );
  XNOR U51514 ( .A(n50870), .B(n50868), .Z(n51085) );
  AND U51515 ( .A(n51086), .B(n51087), .Z(n50868) );
  NANDN U51516 ( .A(n51088), .B(n51089), .Z(n51087) );
  OR U51517 ( .A(n51090), .B(n51091), .Z(n51089) );
  NAND U51518 ( .A(n51091), .B(n51090), .Z(n51086) );
  ANDN U51519 ( .B(A[16]), .A(n25), .Z(n50870) );
  XNOR U51520 ( .A(n50878), .B(n51092), .Z(n50871) );
  XNOR U51521 ( .A(n50877), .B(n50875), .Z(n51092) );
  AND U51522 ( .A(n51093), .B(n51094), .Z(n50875) );
  NANDN U51523 ( .A(n51095), .B(n51096), .Z(n51094) );
  NANDN U51524 ( .A(n51097), .B(n51098), .Z(n51096) );
  NANDN U51525 ( .A(n51098), .B(n51097), .Z(n51093) );
  ANDN U51526 ( .B(A[15]), .A(n23), .Z(n50877) );
  XNOR U51527 ( .A(n50885), .B(n51099), .Z(n50878) );
  XNOR U51528 ( .A(n50884), .B(n50882), .Z(n51099) );
  AND U51529 ( .A(n51100), .B(n51101), .Z(n50882) );
  NANDN U51530 ( .A(n51102), .B(n51103), .Z(n51101) );
  OR U51531 ( .A(n51104), .B(n51105), .Z(n51103) );
  NAND U51532 ( .A(n51105), .B(n51104), .Z(n51100) );
  ANDN U51533 ( .B(A[14]), .A(n21), .Z(n50884) );
  XNOR U51534 ( .A(n50892), .B(n51106), .Z(n50885) );
  XNOR U51535 ( .A(n50891), .B(n50889), .Z(n51106) );
  AND U51536 ( .A(n51107), .B(n51108), .Z(n50889) );
  NANDN U51537 ( .A(n51109), .B(n51110), .Z(n51108) );
  NANDN U51538 ( .A(n51111), .B(n51112), .Z(n51110) );
  NANDN U51539 ( .A(n51112), .B(n51111), .Z(n51107) );
  ANDN U51540 ( .B(A[13]), .A(n19), .Z(n50891) );
  XNOR U51541 ( .A(n50899), .B(n51113), .Z(n50892) );
  XNOR U51542 ( .A(n50898), .B(n50896), .Z(n51113) );
  AND U51543 ( .A(n51114), .B(n51115), .Z(n50896) );
  NANDN U51544 ( .A(n51116), .B(n51117), .Z(n51115) );
  OR U51545 ( .A(n51118), .B(n51119), .Z(n51117) );
  NAND U51546 ( .A(n51119), .B(n51118), .Z(n51114) );
  ANDN U51547 ( .B(A[12]), .A(n17), .Z(n50898) );
  XNOR U51548 ( .A(n50906), .B(n51120), .Z(n50899) );
  XNOR U51549 ( .A(n50905), .B(n50903), .Z(n51120) );
  AND U51550 ( .A(n51121), .B(n51122), .Z(n50903) );
  NANDN U51551 ( .A(n51123), .B(n51124), .Z(n51122) );
  NANDN U51552 ( .A(n51125), .B(n51126), .Z(n51124) );
  NANDN U51553 ( .A(n51126), .B(n51125), .Z(n51121) );
  ANDN U51554 ( .B(A[11]), .A(n15), .Z(n50905) );
  XNOR U51555 ( .A(n50913), .B(n51127), .Z(n50906) );
  XNOR U51556 ( .A(n50912), .B(n50910), .Z(n51127) );
  AND U51557 ( .A(n51128), .B(n51129), .Z(n50910) );
  NANDN U51558 ( .A(n51130), .B(n51131), .Z(n51129) );
  OR U51559 ( .A(n51132), .B(n51133), .Z(n51131) );
  NAND U51560 ( .A(n51133), .B(n51132), .Z(n51128) );
  ANDN U51561 ( .B(A[10]), .A(n13), .Z(n50912) );
  XNOR U51562 ( .A(n50920), .B(n51134), .Z(n50913) );
  XNOR U51563 ( .A(n50919), .B(n50917), .Z(n51134) );
  AND U51564 ( .A(n51135), .B(n51136), .Z(n50917) );
  NANDN U51565 ( .A(n51137), .B(n51138), .Z(n51136) );
  NANDN U51566 ( .A(n51139), .B(n51140), .Z(n51138) );
  NANDN U51567 ( .A(n51140), .B(n51139), .Z(n51135) );
  ANDN U51568 ( .B(A[9]), .A(n11), .Z(n50919) );
  XNOR U51569 ( .A(n50927), .B(n51141), .Z(n50920) );
  XNOR U51570 ( .A(n50926), .B(n50924), .Z(n51141) );
  AND U51571 ( .A(n51142), .B(n51143), .Z(n50924) );
  NANDN U51572 ( .A(n51144), .B(n51145), .Z(n51143) );
  OR U51573 ( .A(n51146), .B(n51147), .Z(n51145) );
  NAND U51574 ( .A(n51147), .B(n51146), .Z(n51142) );
  ANDN U51575 ( .B(A[8]), .A(n9), .Z(n50926) );
  XNOR U51576 ( .A(n50934), .B(n51148), .Z(n50927) );
  XNOR U51577 ( .A(n50933), .B(n50931), .Z(n51148) );
  AND U51578 ( .A(n51149), .B(n51150), .Z(n50931) );
  NANDN U51579 ( .A(n51151), .B(n51152), .Z(n51150) );
  NANDN U51580 ( .A(n51153), .B(n51154), .Z(n51152) );
  NANDN U51581 ( .A(n51154), .B(n51153), .Z(n51149) );
  ANDN U51582 ( .B(B[98]), .A(n78), .Z(n50933) );
  XNOR U51583 ( .A(n50941), .B(n51155), .Z(n50934) );
  XNOR U51584 ( .A(n50940), .B(n50938), .Z(n51155) );
  AND U51585 ( .A(n51156), .B(n51157), .Z(n50938) );
  NANDN U51586 ( .A(n51158), .B(n51159), .Z(n51157) );
  OR U51587 ( .A(n51160), .B(n51161), .Z(n51159) );
  NAND U51588 ( .A(n51161), .B(n51160), .Z(n51156) );
  ANDN U51589 ( .B(A[6]), .A(n6), .Z(n50940) );
  XNOR U51590 ( .A(n50948), .B(n51162), .Z(n50941) );
  XNOR U51591 ( .A(n50947), .B(n50945), .Z(n51162) );
  AND U51592 ( .A(n51163), .B(n51164), .Z(n50945) );
  NANDN U51593 ( .A(n51165), .B(n51166), .Z(n51164) );
  NANDN U51594 ( .A(n51167), .B(n51168), .Z(n51166) );
  NANDN U51595 ( .A(n51168), .B(n51167), .Z(n51163) );
  ANDN U51596 ( .B(A[5]), .A(n4), .Z(n50947) );
  XNOR U51597 ( .A(n50955), .B(n51169), .Z(n50948) );
  XNOR U51598 ( .A(n50954), .B(n50952), .Z(n51169) );
  AND U51599 ( .A(n51170), .B(n51171), .Z(n50952) );
  NANDN U51600 ( .A(n51172), .B(n51173), .Z(n51171) );
  OR U51601 ( .A(n51174), .B(n51175), .Z(n51173) );
  NAND U51602 ( .A(n51175), .B(n51174), .Z(n51170) );
  ANDN U51603 ( .B(B[101]), .A(n81), .Z(n50954) );
  XNOR U51604 ( .A(n50962), .B(n51176), .Z(n50955) );
  XNOR U51605 ( .A(n50961), .B(n50959), .Z(n51176) );
  AND U51606 ( .A(n51177), .B(n51178), .Z(n50959) );
  NANDN U51607 ( .A(n51179), .B(n51180), .Z(n51178) );
  NAND U51608 ( .A(n51181), .B(n51182), .Z(n51180) );
  ANDN U51609 ( .B(B[102]), .A(n82), .Z(n50961) );
  XOR U51610 ( .A(n50968), .B(n51183), .Z(n50962) );
  XNOR U51611 ( .A(n50966), .B(n50969), .Z(n51183) );
  NAND U51612 ( .A(A[2]), .B(B[103]), .Z(n50969) );
  NANDN U51613 ( .A(n51184), .B(n51185), .Z(n50966) );
  AND U51614 ( .A(A[0]), .B(B[104]), .Z(n51185) );
  XNOR U51615 ( .A(n50971), .B(n51186), .Z(n50968) );
  NAND U51616 ( .A(A[0]), .B(B[105]), .Z(n51186) );
  NAND U51617 ( .A(B[104]), .B(A[1]), .Z(n50971) );
  NAND U51618 ( .A(n51187), .B(n51188), .Z(n586) );
  NANDN U51619 ( .A(n51189), .B(n51190), .Z(n51188) );
  OR U51620 ( .A(n51191), .B(n51192), .Z(n51190) );
  NAND U51621 ( .A(n51192), .B(n51191), .Z(n51187) );
  XOR U51622 ( .A(n588), .B(n587), .Z(\A1[102] ) );
  XOR U51623 ( .A(n51192), .B(n51193), .Z(n587) );
  XNOR U51624 ( .A(n51191), .B(n51189), .Z(n51193) );
  AND U51625 ( .A(n51194), .B(n51195), .Z(n51189) );
  NANDN U51626 ( .A(n51196), .B(n51197), .Z(n51195) );
  NANDN U51627 ( .A(n51198), .B(n51199), .Z(n51197) );
  NANDN U51628 ( .A(n51199), .B(n51198), .Z(n51194) );
  ANDN U51629 ( .B(B[73]), .A(n54), .Z(n51191) );
  XNOR U51630 ( .A(n50986), .B(n51200), .Z(n51192) );
  XNOR U51631 ( .A(n50985), .B(n50983), .Z(n51200) );
  AND U51632 ( .A(n51201), .B(n51202), .Z(n50983) );
  NANDN U51633 ( .A(n51203), .B(n51204), .Z(n51202) );
  OR U51634 ( .A(n51205), .B(n51206), .Z(n51204) );
  NAND U51635 ( .A(n51206), .B(n51205), .Z(n51201) );
  ANDN U51636 ( .B(B[74]), .A(n55), .Z(n50985) );
  XNOR U51637 ( .A(n50993), .B(n51207), .Z(n50986) );
  XNOR U51638 ( .A(n50992), .B(n50990), .Z(n51207) );
  AND U51639 ( .A(n51208), .B(n51209), .Z(n50990) );
  NANDN U51640 ( .A(n51210), .B(n51211), .Z(n51209) );
  NANDN U51641 ( .A(n51212), .B(n51213), .Z(n51211) );
  NANDN U51642 ( .A(n51213), .B(n51212), .Z(n51208) );
  ANDN U51643 ( .B(B[75]), .A(n56), .Z(n50992) );
  XNOR U51644 ( .A(n51000), .B(n51214), .Z(n50993) );
  XNOR U51645 ( .A(n50999), .B(n50997), .Z(n51214) );
  AND U51646 ( .A(n51215), .B(n51216), .Z(n50997) );
  NANDN U51647 ( .A(n51217), .B(n51218), .Z(n51216) );
  OR U51648 ( .A(n51219), .B(n51220), .Z(n51218) );
  NAND U51649 ( .A(n51220), .B(n51219), .Z(n51215) );
  ANDN U51650 ( .B(B[76]), .A(n57), .Z(n50999) );
  XNOR U51651 ( .A(n51007), .B(n51221), .Z(n51000) );
  XNOR U51652 ( .A(n51006), .B(n51004), .Z(n51221) );
  AND U51653 ( .A(n51222), .B(n51223), .Z(n51004) );
  NANDN U51654 ( .A(n51224), .B(n51225), .Z(n51223) );
  NANDN U51655 ( .A(n51226), .B(n51227), .Z(n51225) );
  NANDN U51656 ( .A(n51227), .B(n51226), .Z(n51222) );
  ANDN U51657 ( .B(B[77]), .A(n58), .Z(n51006) );
  XNOR U51658 ( .A(n51014), .B(n51228), .Z(n51007) );
  XNOR U51659 ( .A(n51013), .B(n51011), .Z(n51228) );
  AND U51660 ( .A(n51229), .B(n51230), .Z(n51011) );
  NANDN U51661 ( .A(n51231), .B(n51232), .Z(n51230) );
  OR U51662 ( .A(n51233), .B(n51234), .Z(n51232) );
  NAND U51663 ( .A(n51234), .B(n51233), .Z(n51229) );
  ANDN U51664 ( .B(B[78]), .A(n59), .Z(n51013) );
  XNOR U51665 ( .A(n51021), .B(n51235), .Z(n51014) );
  XNOR U51666 ( .A(n51020), .B(n51018), .Z(n51235) );
  AND U51667 ( .A(n51236), .B(n51237), .Z(n51018) );
  NANDN U51668 ( .A(n51238), .B(n51239), .Z(n51237) );
  NANDN U51669 ( .A(n51240), .B(n51241), .Z(n51239) );
  NANDN U51670 ( .A(n51241), .B(n51240), .Z(n51236) );
  ANDN U51671 ( .B(B[79]), .A(n60), .Z(n51020) );
  XNOR U51672 ( .A(n51028), .B(n51242), .Z(n51021) );
  XNOR U51673 ( .A(n51027), .B(n51025), .Z(n51242) );
  AND U51674 ( .A(n51243), .B(n51244), .Z(n51025) );
  NANDN U51675 ( .A(n51245), .B(n51246), .Z(n51244) );
  OR U51676 ( .A(n51247), .B(n51248), .Z(n51246) );
  NAND U51677 ( .A(n51248), .B(n51247), .Z(n51243) );
  ANDN U51678 ( .B(B[80]), .A(n61), .Z(n51027) );
  XNOR U51679 ( .A(n51035), .B(n51249), .Z(n51028) );
  XNOR U51680 ( .A(n51034), .B(n51032), .Z(n51249) );
  AND U51681 ( .A(n51250), .B(n51251), .Z(n51032) );
  NANDN U51682 ( .A(n51252), .B(n51253), .Z(n51251) );
  NANDN U51683 ( .A(n51254), .B(n51255), .Z(n51253) );
  NANDN U51684 ( .A(n51255), .B(n51254), .Z(n51250) );
  ANDN U51685 ( .B(B[81]), .A(n62), .Z(n51034) );
  XNOR U51686 ( .A(n51042), .B(n51256), .Z(n51035) );
  XNOR U51687 ( .A(n51041), .B(n51039), .Z(n51256) );
  AND U51688 ( .A(n51257), .B(n51258), .Z(n51039) );
  NANDN U51689 ( .A(n51259), .B(n51260), .Z(n51258) );
  OR U51690 ( .A(n51261), .B(n51262), .Z(n51260) );
  NAND U51691 ( .A(n51262), .B(n51261), .Z(n51257) );
  ANDN U51692 ( .B(B[82]), .A(n63), .Z(n51041) );
  XNOR U51693 ( .A(n51049), .B(n51263), .Z(n51042) );
  XNOR U51694 ( .A(n51048), .B(n51046), .Z(n51263) );
  AND U51695 ( .A(n51264), .B(n51265), .Z(n51046) );
  NANDN U51696 ( .A(n51266), .B(n51267), .Z(n51265) );
  NANDN U51697 ( .A(n51268), .B(n51269), .Z(n51267) );
  NANDN U51698 ( .A(n51269), .B(n51268), .Z(n51264) );
  ANDN U51699 ( .B(B[83]), .A(n64), .Z(n51048) );
  XNOR U51700 ( .A(n51056), .B(n51270), .Z(n51049) );
  XNOR U51701 ( .A(n51055), .B(n51053), .Z(n51270) );
  AND U51702 ( .A(n51271), .B(n51272), .Z(n51053) );
  NANDN U51703 ( .A(n51273), .B(n51274), .Z(n51272) );
  OR U51704 ( .A(n51275), .B(n51276), .Z(n51274) );
  NAND U51705 ( .A(n51276), .B(n51275), .Z(n51271) );
  ANDN U51706 ( .B(B[84]), .A(n65), .Z(n51055) );
  XNOR U51707 ( .A(n51063), .B(n51277), .Z(n51056) );
  XNOR U51708 ( .A(n51062), .B(n51060), .Z(n51277) );
  AND U51709 ( .A(n51278), .B(n51279), .Z(n51060) );
  NANDN U51710 ( .A(n51280), .B(n51281), .Z(n51279) );
  NANDN U51711 ( .A(n51282), .B(n51283), .Z(n51281) );
  NANDN U51712 ( .A(n51283), .B(n51282), .Z(n51278) );
  ANDN U51713 ( .B(B[85]), .A(n66), .Z(n51062) );
  XNOR U51714 ( .A(n51070), .B(n51284), .Z(n51063) );
  XNOR U51715 ( .A(n51069), .B(n51067), .Z(n51284) );
  AND U51716 ( .A(n51285), .B(n51286), .Z(n51067) );
  NANDN U51717 ( .A(n51287), .B(n51288), .Z(n51286) );
  OR U51718 ( .A(n51289), .B(n51290), .Z(n51288) );
  NAND U51719 ( .A(n51290), .B(n51289), .Z(n51285) );
  ANDN U51720 ( .B(A[18]), .A(n31), .Z(n51069) );
  XNOR U51721 ( .A(n51077), .B(n51291), .Z(n51070) );
  XNOR U51722 ( .A(n51076), .B(n51074), .Z(n51291) );
  AND U51723 ( .A(n51292), .B(n51293), .Z(n51074) );
  NANDN U51724 ( .A(n51294), .B(n51295), .Z(n51293) );
  NANDN U51725 ( .A(n51296), .B(n51297), .Z(n51295) );
  NANDN U51726 ( .A(n51297), .B(n51296), .Z(n51292) );
  ANDN U51727 ( .B(A[17]), .A(n29), .Z(n51076) );
  XNOR U51728 ( .A(n51084), .B(n51298), .Z(n51077) );
  XNOR U51729 ( .A(n51083), .B(n51081), .Z(n51298) );
  AND U51730 ( .A(n51299), .B(n51300), .Z(n51081) );
  NANDN U51731 ( .A(n51301), .B(n51302), .Z(n51300) );
  OR U51732 ( .A(n51303), .B(n51304), .Z(n51302) );
  NAND U51733 ( .A(n51304), .B(n51303), .Z(n51299) );
  ANDN U51734 ( .B(A[16]), .A(n27), .Z(n51083) );
  XNOR U51735 ( .A(n51091), .B(n51305), .Z(n51084) );
  XNOR U51736 ( .A(n51090), .B(n51088), .Z(n51305) );
  AND U51737 ( .A(n51306), .B(n51307), .Z(n51088) );
  NANDN U51738 ( .A(n51308), .B(n51309), .Z(n51307) );
  NANDN U51739 ( .A(n51310), .B(n51311), .Z(n51309) );
  NANDN U51740 ( .A(n51311), .B(n51310), .Z(n51306) );
  ANDN U51741 ( .B(A[15]), .A(n25), .Z(n51090) );
  XNOR U51742 ( .A(n51098), .B(n51312), .Z(n51091) );
  XNOR U51743 ( .A(n51097), .B(n51095), .Z(n51312) );
  AND U51744 ( .A(n51313), .B(n51314), .Z(n51095) );
  NANDN U51745 ( .A(n51315), .B(n51316), .Z(n51314) );
  OR U51746 ( .A(n51317), .B(n51318), .Z(n51316) );
  NAND U51747 ( .A(n51318), .B(n51317), .Z(n51313) );
  ANDN U51748 ( .B(A[14]), .A(n23), .Z(n51097) );
  XNOR U51749 ( .A(n51105), .B(n51319), .Z(n51098) );
  XNOR U51750 ( .A(n51104), .B(n51102), .Z(n51319) );
  AND U51751 ( .A(n51320), .B(n51321), .Z(n51102) );
  NANDN U51752 ( .A(n51322), .B(n51323), .Z(n51321) );
  NANDN U51753 ( .A(n51324), .B(n51325), .Z(n51323) );
  NANDN U51754 ( .A(n51325), .B(n51324), .Z(n51320) );
  ANDN U51755 ( .B(A[13]), .A(n21), .Z(n51104) );
  XNOR U51756 ( .A(n51112), .B(n51326), .Z(n51105) );
  XNOR U51757 ( .A(n51111), .B(n51109), .Z(n51326) );
  AND U51758 ( .A(n51327), .B(n51328), .Z(n51109) );
  NANDN U51759 ( .A(n51329), .B(n51330), .Z(n51328) );
  OR U51760 ( .A(n51331), .B(n51332), .Z(n51330) );
  NAND U51761 ( .A(n51332), .B(n51331), .Z(n51327) );
  ANDN U51762 ( .B(A[12]), .A(n19), .Z(n51111) );
  XNOR U51763 ( .A(n51119), .B(n51333), .Z(n51112) );
  XNOR U51764 ( .A(n51118), .B(n51116), .Z(n51333) );
  AND U51765 ( .A(n51334), .B(n51335), .Z(n51116) );
  NANDN U51766 ( .A(n51336), .B(n51337), .Z(n51335) );
  NANDN U51767 ( .A(n51338), .B(n51339), .Z(n51337) );
  NANDN U51768 ( .A(n51339), .B(n51338), .Z(n51334) );
  ANDN U51769 ( .B(A[11]), .A(n17), .Z(n51118) );
  XNOR U51770 ( .A(n51126), .B(n51340), .Z(n51119) );
  XNOR U51771 ( .A(n51125), .B(n51123), .Z(n51340) );
  AND U51772 ( .A(n51341), .B(n51342), .Z(n51123) );
  NANDN U51773 ( .A(n51343), .B(n51344), .Z(n51342) );
  OR U51774 ( .A(n51345), .B(n51346), .Z(n51344) );
  NAND U51775 ( .A(n51346), .B(n51345), .Z(n51341) );
  ANDN U51776 ( .B(A[10]), .A(n15), .Z(n51125) );
  XNOR U51777 ( .A(n51133), .B(n51347), .Z(n51126) );
  XNOR U51778 ( .A(n51132), .B(n51130), .Z(n51347) );
  AND U51779 ( .A(n51348), .B(n51349), .Z(n51130) );
  NANDN U51780 ( .A(n51350), .B(n51351), .Z(n51349) );
  NANDN U51781 ( .A(n51352), .B(n51353), .Z(n51351) );
  NANDN U51782 ( .A(n51353), .B(n51352), .Z(n51348) );
  ANDN U51783 ( .B(A[9]), .A(n13), .Z(n51132) );
  XNOR U51784 ( .A(n51140), .B(n51354), .Z(n51133) );
  XNOR U51785 ( .A(n51139), .B(n51137), .Z(n51354) );
  AND U51786 ( .A(n51355), .B(n51356), .Z(n51137) );
  NANDN U51787 ( .A(n51357), .B(n51358), .Z(n51356) );
  OR U51788 ( .A(n51359), .B(n51360), .Z(n51358) );
  NAND U51789 ( .A(n51360), .B(n51359), .Z(n51355) );
  ANDN U51790 ( .B(A[8]), .A(n11), .Z(n51139) );
  XNOR U51791 ( .A(n51147), .B(n51361), .Z(n51140) );
  XNOR U51792 ( .A(n51146), .B(n51144), .Z(n51361) );
  AND U51793 ( .A(n51362), .B(n51363), .Z(n51144) );
  NANDN U51794 ( .A(n51364), .B(n51365), .Z(n51363) );
  NANDN U51795 ( .A(n51366), .B(n51367), .Z(n51365) );
  NANDN U51796 ( .A(n51367), .B(n51366), .Z(n51362) );
  ANDN U51797 ( .B(A[7]), .A(n9), .Z(n51146) );
  XNOR U51798 ( .A(n51154), .B(n51368), .Z(n51147) );
  XNOR U51799 ( .A(n51153), .B(n51151), .Z(n51368) );
  AND U51800 ( .A(n51369), .B(n51370), .Z(n51151) );
  NANDN U51801 ( .A(n51371), .B(n51372), .Z(n51370) );
  OR U51802 ( .A(n51373), .B(n51374), .Z(n51372) );
  NAND U51803 ( .A(n51374), .B(n51373), .Z(n51369) );
  ANDN U51804 ( .B(B[98]), .A(n79), .Z(n51153) );
  XNOR U51805 ( .A(n51161), .B(n51375), .Z(n51154) );
  XNOR U51806 ( .A(n51160), .B(n51158), .Z(n51375) );
  AND U51807 ( .A(n51376), .B(n51377), .Z(n51158) );
  NANDN U51808 ( .A(n51378), .B(n51379), .Z(n51377) );
  NANDN U51809 ( .A(n51380), .B(n51381), .Z(n51379) );
  NANDN U51810 ( .A(n51381), .B(n51380), .Z(n51376) );
  ANDN U51811 ( .B(A[5]), .A(n6), .Z(n51160) );
  XNOR U51812 ( .A(n51168), .B(n51382), .Z(n51161) );
  XNOR U51813 ( .A(n51167), .B(n51165), .Z(n51382) );
  AND U51814 ( .A(n51383), .B(n51384), .Z(n51165) );
  NANDN U51815 ( .A(n51385), .B(n51386), .Z(n51384) );
  OR U51816 ( .A(n51387), .B(n51388), .Z(n51386) );
  NAND U51817 ( .A(n51388), .B(n51387), .Z(n51383) );
  ANDN U51818 ( .B(A[4]), .A(n4), .Z(n51167) );
  XNOR U51819 ( .A(n51175), .B(n51389), .Z(n51168) );
  XNOR U51820 ( .A(n51174), .B(n51172), .Z(n51389) );
  AND U51821 ( .A(n51390), .B(n51391), .Z(n51172) );
  NANDN U51822 ( .A(n51392), .B(n51393), .Z(n51391) );
  NAND U51823 ( .A(n51394), .B(n51395), .Z(n51393) );
  ANDN U51824 ( .B(B[101]), .A(n82), .Z(n51174) );
  XOR U51825 ( .A(n51181), .B(n51396), .Z(n51175) );
  XNOR U51826 ( .A(n51179), .B(n51182), .Z(n51396) );
  NAND U51827 ( .A(A[2]), .B(B[102]), .Z(n51182) );
  NANDN U51828 ( .A(n51397), .B(n51398), .Z(n51179) );
  AND U51829 ( .A(A[0]), .B(B[103]), .Z(n51398) );
  XNOR U51830 ( .A(n51184), .B(n51399), .Z(n51181) );
  NAND U51831 ( .A(A[0]), .B(B[104]), .Z(n51399) );
  NAND U51832 ( .A(B[103]), .B(A[1]), .Z(n51184) );
  NAND U51833 ( .A(n51400), .B(n51401), .Z(n588) );
  NANDN U51834 ( .A(n51402), .B(n51403), .Z(n51401) );
  OR U51835 ( .A(n51404), .B(n51405), .Z(n51403) );
  NAND U51836 ( .A(n51405), .B(n51404), .Z(n51400) );
  XOR U51837 ( .A(n590), .B(n589), .Z(\A1[101] ) );
  XOR U51838 ( .A(n51405), .B(n51406), .Z(n589) );
  XNOR U51839 ( .A(n51404), .B(n51402), .Z(n51406) );
  AND U51840 ( .A(n51407), .B(n51408), .Z(n51402) );
  NANDN U51841 ( .A(n51409), .B(n51410), .Z(n51408) );
  NANDN U51842 ( .A(n51411), .B(n51412), .Z(n51410) );
  NANDN U51843 ( .A(n51412), .B(n51411), .Z(n51407) );
  ANDN U51844 ( .B(B[72]), .A(n54), .Z(n51404) );
  XNOR U51845 ( .A(n51199), .B(n51413), .Z(n51405) );
  XNOR U51846 ( .A(n51198), .B(n51196), .Z(n51413) );
  AND U51847 ( .A(n51414), .B(n51415), .Z(n51196) );
  NANDN U51848 ( .A(n51416), .B(n51417), .Z(n51415) );
  OR U51849 ( .A(n51418), .B(n51419), .Z(n51417) );
  NAND U51850 ( .A(n51419), .B(n51418), .Z(n51414) );
  ANDN U51851 ( .B(B[73]), .A(n55), .Z(n51198) );
  XNOR U51852 ( .A(n51206), .B(n51420), .Z(n51199) );
  XNOR U51853 ( .A(n51205), .B(n51203), .Z(n51420) );
  AND U51854 ( .A(n51421), .B(n51422), .Z(n51203) );
  NANDN U51855 ( .A(n51423), .B(n51424), .Z(n51422) );
  NANDN U51856 ( .A(n51425), .B(n51426), .Z(n51424) );
  NANDN U51857 ( .A(n51426), .B(n51425), .Z(n51421) );
  ANDN U51858 ( .B(B[74]), .A(n56), .Z(n51205) );
  XNOR U51859 ( .A(n51213), .B(n51427), .Z(n51206) );
  XNOR U51860 ( .A(n51212), .B(n51210), .Z(n51427) );
  AND U51861 ( .A(n51428), .B(n51429), .Z(n51210) );
  NANDN U51862 ( .A(n51430), .B(n51431), .Z(n51429) );
  OR U51863 ( .A(n51432), .B(n51433), .Z(n51431) );
  NAND U51864 ( .A(n51433), .B(n51432), .Z(n51428) );
  ANDN U51865 ( .B(B[75]), .A(n57), .Z(n51212) );
  XNOR U51866 ( .A(n51220), .B(n51434), .Z(n51213) );
  XNOR U51867 ( .A(n51219), .B(n51217), .Z(n51434) );
  AND U51868 ( .A(n51435), .B(n51436), .Z(n51217) );
  NANDN U51869 ( .A(n51437), .B(n51438), .Z(n51436) );
  NANDN U51870 ( .A(n51439), .B(n51440), .Z(n51438) );
  NANDN U51871 ( .A(n51440), .B(n51439), .Z(n51435) );
  ANDN U51872 ( .B(B[76]), .A(n58), .Z(n51219) );
  XNOR U51873 ( .A(n51227), .B(n51441), .Z(n51220) );
  XNOR U51874 ( .A(n51226), .B(n51224), .Z(n51441) );
  AND U51875 ( .A(n51442), .B(n51443), .Z(n51224) );
  NANDN U51876 ( .A(n51444), .B(n51445), .Z(n51443) );
  OR U51877 ( .A(n51446), .B(n51447), .Z(n51445) );
  NAND U51878 ( .A(n51447), .B(n51446), .Z(n51442) );
  ANDN U51879 ( .B(B[77]), .A(n59), .Z(n51226) );
  XNOR U51880 ( .A(n51234), .B(n51448), .Z(n51227) );
  XNOR U51881 ( .A(n51233), .B(n51231), .Z(n51448) );
  AND U51882 ( .A(n51449), .B(n51450), .Z(n51231) );
  NANDN U51883 ( .A(n51451), .B(n51452), .Z(n51450) );
  NANDN U51884 ( .A(n51453), .B(n51454), .Z(n51452) );
  NANDN U51885 ( .A(n51454), .B(n51453), .Z(n51449) );
  ANDN U51886 ( .B(B[78]), .A(n60), .Z(n51233) );
  XNOR U51887 ( .A(n51241), .B(n51455), .Z(n51234) );
  XNOR U51888 ( .A(n51240), .B(n51238), .Z(n51455) );
  AND U51889 ( .A(n51456), .B(n51457), .Z(n51238) );
  NANDN U51890 ( .A(n51458), .B(n51459), .Z(n51457) );
  OR U51891 ( .A(n51460), .B(n51461), .Z(n51459) );
  NAND U51892 ( .A(n51461), .B(n51460), .Z(n51456) );
  ANDN U51893 ( .B(B[79]), .A(n61), .Z(n51240) );
  XNOR U51894 ( .A(n51248), .B(n51462), .Z(n51241) );
  XNOR U51895 ( .A(n51247), .B(n51245), .Z(n51462) );
  AND U51896 ( .A(n51463), .B(n51464), .Z(n51245) );
  NANDN U51897 ( .A(n51465), .B(n51466), .Z(n51464) );
  NANDN U51898 ( .A(n51467), .B(n51468), .Z(n51466) );
  NANDN U51899 ( .A(n51468), .B(n51467), .Z(n51463) );
  ANDN U51900 ( .B(B[80]), .A(n62), .Z(n51247) );
  XNOR U51901 ( .A(n51255), .B(n51469), .Z(n51248) );
  XNOR U51902 ( .A(n51254), .B(n51252), .Z(n51469) );
  AND U51903 ( .A(n51470), .B(n51471), .Z(n51252) );
  NANDN U51904 ( .A(n51472), .B(n51473), .Z(n51471) );
  OR U51905 ( .A(n51474), .B(n51475), .Z(n51473) );
  NAND U51906 ( .A(n51475), .B(n51474), .Z(n51470) );
  ANDN U51907 ( .B(B[81]), .A(n63), .Z(n51254) );
  XNOR U51908 ( .A(n51262), .B(n51476), .Z(n51255) );
  XNOR U51909 ( .A(n51261), .B(n51259), .Z(n51476) );
  AND U51910 ( .A(n51477), .B(n51478), .Z(n51259) );
  NANDN U51911 ( .A(n51479), .B(n51480), .Z(n51478) );
  NANDN U51912 ( .A(n51481), .B(n51482), .Z(n51480) );
  NANDN U51913 ( .A(n51482), .B(n51481), .Z(n51477) );
  ANDN U51914 ( .B(B[82]), .A(n64), .Z(n51261) );
  XNOR U51915 ( .A(n51269), .B(n51483), .Z(n51262) );
  XNOR U51916 ( .A(n51268), .B(n51266), .Z(n51483) );
  AND U51917 ( .A(n51484), .B(n51485), .Z(n51266) );
  NANDN U51918 ( .A(n51486), .B(n51487), .Z(n51485) );
  OR U51919 ( .A(n51488), .B(n51489), .Z(n51487) );
  NAND U51920 ( .A(n51489), .B(n51488), .Z(n51484) );
  ANDN U51921 ( .B(B[83]), .A(n65), .Z(n51268) );
  XNOR U51922 ( .A(n51276), .B(n51490), .Z(n51269) );
  XNOR U51923 ( .A(n51275), .B(n51273), .Z(n51490) );
  AND U51924 ( .A(n51491), .B(n51492), .Z(n51273) );
  NANDN U51925 ( .A(n51493), .B(n51494), .Z(n51492) );
  NANDN U51926 ( .A(n51495), .B(n51496), .Z(n51494) );
  NANDN U51927 ( .A(n51496), .B(n51495), .Z(n51491) );
  ANDN U51928 ( .B(B[84]), .A(n66), .Z(n51275) );
  XNOR U51929 ( .A(n51283), .B(n51497), .Z(n51276) );
  XNOR U51930 ( .A(n51282), .B(n51280), .Z(n51497) );
  AND U51931 ( .A(n51498), .B(n51499), .Z(n51280) );
  NANDN U51932 ( .A(n51500), .B(n51501), .Z(n51499) );
  OR U51933 ( .A(n51502), .B(n51503), .Z(n51501) );
  NAND U51934 ( .A(n51503), .B(n51502), .Z(n51498) );
  ANDN U51935 ( .B(B[85]), .A(n67), .Z(n51282) );
  XNOR U51936 ( .A(n51290), .B(n51504), .Z(n51283) );
  XNOR U51937 ( .A(n51289), .B(n51287), .Z(n51504) );
  AND U51938 ( .A(n51505), .B(n51506), .Z(n51287) );
  NANDN U51939 ( .A(n51507), .B(n51508), .Z(n51506) );
  NANDN U51940 ( .A(n51509), .B(n51510), .Z(n51508) );
  NANDN U51941 ( .A(n51510), .B(n51509), .Z(n51505) );
  ANDN U51942 ( .B(A[17]), .A(n31), .Z(n51289) );
  XNOR U51943 ( .A(n51297), .B(n51511), .Z(n51290) );
  XNOR U51944 ( .A(n51296), .B(n51294), .Z(n51511) );
  AND U51945 ( .A(n51512), .B(n51513), .Z(n51294) );
  NANDN U51946 ( .A(n51514), .B(n51515), .Z(n51513) );
  OR U51947 ( .A(n51516), .B(n51517), .Z(n51515) );
  NAND U51948 ( .A(n51517), .B(n51516), .Z(n51512) );
  ANDN U51949 ( .B(A[16]), .A(n29), .Z(n51296) );
  XNOR U51950 ( .A(n51304), .B(n51518), .Z(n51297) );
  XNOR U51951 ( .A(n51303), .B(n51301), .Z(n51518) );
  AND U51952 ( .A(n51519), .B(n51520), .Z(n51301) );
  NANDN U51953 ( .A(n51521), .B(n51522), .Z(n51520) );
  NANDN U51954 ( .A(n51523), .B(n51524), .Z(n51522) );
  NANDN U51955 ( .A(n51524), .B(n51523), .Z(n51519) );
  ANDN U51956 ( .B(A[15]), .A(n27), .Z(n51303) );
  XNOR U51957 ( .A(n51311), .B(n51525), .Z(n51304) );
  XNOR U51958 ( .A(n51310), .B(n51308), .Z(n51525) );
  AND U51959 ( .A(n51526), .B(n51527), .Z(n51308) );
  NANDN U51960 ( .A(n51528), .B(n51529), .Z(n51527) );
  OR U51961 ( .A(n51530), .B(n51531), .Z(n51529) );
  NAND U51962 ( .A(n51531), .B(n51530), .Z(n51526) );
  ANDN U51963 ( .B(A[14]), .A(n25), .Z(n51310) );
  XNOR U51964 ( .A(n51318), .B(n51532), .Z(n51311) );
  XNOR U51965 ( .A(n51317), .B(n51315), .Z(n51532) );
  AND U51966 ( .A(n51533), .B(n51534), .Z(n51315) );
  NANDN U51967 ( .A(n51535), .B(n51536), .Z(n51534) );
  NANDN U51968 ( .A(n51537), .B(n51538), .Z(n51536) );
  NANDN U51969 ( .A(n51538), .B(n51537), .Z(n51533) );
  ANDN U51970 ( .B(A[13]), .A(n23), .Z(n51317) );
  XNOR U51971 ( .A(n51325), .B(n51539), .Z(n51318) );
  XNOR U51972 ( .A(n51324), .B(n51322), .Z(n51539) );
  AND U51973 ( .A(n51540), .B(n51541), .Z(n51322) );
  NANDN U51974 ( .A(n51542), .B(n51543), .Z(n51541) );
  OR U51975 ( .A(n51544), .B(n51545), .Z(n51543) );
  NAND U51976 ( .A(n51545), .B(n51544), .Z(n51540) );
  ANDN U51977 ( .B(A[12]), .A(n21), .Z(n51324) );
  XNOR U51978 ( .A(n51332), .B(n51546), .Z(n51325) );
  XNOR U51979 ( .A(n51331), .B(n51329), .Z(n51546) );
  AND U51980 ( .A(n51547), .B(n51548), .Z(n51329) );
  NANDN U51981 ( .A(n51549), .B(n51550), .Z(n51548) );
  NANDN U51982 ( .A(n51551), .B(n51552), .Z(n51550) );
  NANDN U51983 ( .A(n51552), .B(n51551), .Z(n51547) );
  ANDN U51984 ( .B(A[11]), .A(n19), .Z(n51331) );
  XNOR U51985 ( .A(n51339), .B(n51553), .Z(n51332) );
  XNOR U51986 ( .A(n51338), .B(n51336), .Z(n51553) );
  AND U51987 ( .A(n51554), .B(n51555), .Z(n51336) );
  NANDN U51988 ( .A(n51556), .B(n51557), .Z(n51555) );
  OR U51989 ( .A(n51558), .B(n51559), .Z(n51557) );
  NAND U51990 ( .A(n51559), .B(n51558), .Z(n51554) );
  ANDN U51991 ( .B(A[10]), .A(n17), .Z(n51338) );
  XNOR U51992 ( .A(n51346), .B(n51560), .Z(n51339) );
  XNOR U51993 ( .A(n51345), .B(n51343), .Z(n51560) );
  AND U51994 ( .A(n51561), .B(n51562), .Z(n51343) );
  NANDN U51995 ( .A(n51563), .B(n51564), .Z(n51562) );
  NANDN U51996 ( .A(n51565), .B(n51566), .Z(n51564) );
  NANDN U51997 ( .A(n51566), .B(n51565), .Z(n51561) );
  ANDN U51998 ( .B(A[9]), .A(n15), .Z(n51345) );
  XNOR U51999 ( .A(n51353), .B(n51567), .Z(n51346) );
  XNOR U52000 ( .A(n51352), .B(n51350), .Z(n51567) );
  AND U52001 ( .A(n51568), .B(n51569), .Z(n51350) );
  NANDN U52002 ( .A(n51570), .B(n51571), .Z(n51569) );
  OR U52003 ( .A(n51572), .B(n51573), .Z(n51571) );
  NAND U52004 ( .A(n51573), .B(n51572), .Z(n51568) );
  ANDN U52005 ( .B(A[8]), .A(n13), .Z(n51352) );
  XNOR U52006 ( .A(n51360), .B(n51574), .Z(n51353) );
  XNOR U52007 ( .A(n51359), .B(n51357), .Z(n51574) );
  AND U52008 ( .A(n51575), .B(n51576), .Z(n51357) );
  NANDN U52009 ( .A(n51577), .B(n51578), .Z(n51576) );
  NANDN U52010 ( .A(n51579), .B(n51580), .Z(n51578) );
  NANDN U52011 ( .A(n51580), .B(n51579), .Z(n51575) );
  ANDN U52012 ( .B(A[7]), .A(n11), .Z(n51359) );
  XNOR U52013 ( .A(n51367), .B(n51581), .Z(n51360) );
  XNOR U52014 ( .A(n51366), .B(n51364), .Z(n51581) );
  AND U52015 ( .A(n51582), .B(n51583), .Z(n51364) );
  NANDN U52016 ( .A(n51584), .B(n51585), .Z(n51583) );
  OR U52017 ( .A(n51586), .B(n51587), .Z(n51585) );
  NAND U52018 ( .A(n51587), .B(n51586), .Z(n51582) );
  ANDN U52019 ( .B(A[6]), .A(n9), .Z(n51366) );
  XNOR U52020 ( .A(n51374), .B(n51588), .Z(n51367) );
  XNOR U52021 ( .A(n51373), .B(n51371), .Z(n51588) );
  AND U52022 ( .A(n51589), .B(n51590), .Z(n51371) );
  NANDN U52023 ( .A(n51591), .B(n51592), .Z(n51590) );
  NANDN U52024 ( .A(n51593), .B(n51594), .Z(n51592) );
  NANDN U52025 ( .A(n51594), .B(n51593), .Z(n51589) );
  ANDN U52026 ( .B(B[98]), .A(n80), .Z(n51373) );
  XNOR U52027 ( .A(n51381), .B(n51595), .Z(n51374) );
  XNOR U52028 ( .A(n51380), .B(n51378), .Z(n51595) );
  AND U52029 ( .A(n51596), .B(n51597), .Z(n51378) );
  NANDN U52030 ( .A(n51598), .B(n51599), .Z(n51597) );
  OR U52031 ( .A(n51600), .B(n51601), .Z(n51599) );
  NAND U52032 ( .A(n51601), .B(n51600), .Z(n51596) );
  ANDN U52033 ( .B(A[4]), .A(n6), .Z(n51380) );
  XNOR U52034 ( .A(n51388), .B(n51602), .Z(n51381) );
  XNOR U52035 ( .A(n51387), .B(n51385), .Z(n51602) );
  AND U52036 ( .A(n51603), .B(n51604), .Z(n51385) );
  NANDN U52037 ( .A(n51605), .B(n51606), .Z(n51604) );
  NAND U52038 ( .A(n51607), .B(n51608), .Z(n51606) );
  ANDN U52039 ( .B(A[3]), .A(n4), .Z(n51387) );
  XOR U52040 ( .A(n51394), .B(n51609), .Z(n51388) );
  XNOR U52041 ( .A(n51392), .B(n51395), .Z(n51609) );
  NAND U52042 ( .A(A[2]), .B(B[101]), .Z(n51395) );
  NANDN U52043 ( .A(n51610), .B(n51611), .Z(n51392) );
  AND U52044 ( .A(A[0]), .B(B[102]), .Z(n51611) );
  XNOR U52045 ( .A(n51397), .B(n51612), .Z(n51394) );
  NAND U52046 ( .A(A[0]), .B(B[103]), .Z(n51612) );
  NAND U52047 ( .A(B[102]), .B(A[1]), .Z(n51397) );
  NAND U52048 ( .A(n51613), .B(n51614), .Z(n590) );
  NANDN U52049 ( .A(n51615), .B(n51616), .Z(n51614) );
  OR U52050 ( .A(n51617), .B(n51618), .Z(n51616) );
  NAND U52051 ( .A(n51618), .B(n51617), .Z(n51613) );
  XOR U52052 ( .A(n592), .B(n591), .Z(\A1[100] ) );
  XOR U52053 ( .A(n51618), .B(n51619), .Z(n591) );
  XNOR U52054 ( .A(n51617), .B(n51615), .Z(n51619) );
  AND U52055 ( .A(n51620), .B(n51621), .Z(n51615) );
  NANDN U52056 ( .A(n51622), .B(n51623), .Z(n51621) );
  NAND U52057 ( .A(n51625), .B(n51624), .Z(n51620) );
  ANDN U52058 ( .B(B[71]), .A(n54), .Z(n51617) );
  XNOR U52059 ( .A(n51412), .B(n51626), .Z(n51618) );
  XNOR U52060 ( .A(n51411), .B(n51409), .Z(n51626) );
  AND U52061 ( .A(n51627), .B(n51628), .Z(n51409) );
  NANDN U52062 ( .A(n51629), .B(n51630), .Z(n51628) );
  OR U52063 ( .A(n51631), .B(n51632), .Z(n51630) );
  NAND U52064 ( .A(n51632), .B(n51631), .Z(n51627) );
  ANDN U52065 ( .B(B[72]), .A(n55), .Z(n51411) );
  XNOR U52066 ( .A(n51419), .B(n51633), .Z(n51412) );
  XNOR U52067 ( .A(n51418), .B(n51416), .Z(n51633) );
  AND U52068 ( .A(n51634), .B(n51635), .Z(n51416) );
  NANDN U52069 ( .A(n51636), .B(n51637), .Z(n51635) );
  NANDN U52070 ( .A(n51638), .B(n51639), .Z(n51637) );
  NANDN U52071 ( .A(n51639), .B(n51638), .Z(n51634) );
  ANDN U52072 ( .B(B[73]), .A(n56), .Z(n51418) );
  XNOR U52073 ( .A(n51426), .B(n51640), .Z(n51419) );
  XNOR U52074 ( .A(n51425), .B(n51423), .Z(n51640) );
  AND U52075 ( .A(n51641), .B(n51642), .Z(n51423) );
  NANDN U52076 ( .A(n51643), .B(n51644), .Z(n51642) );
  OR U52077 ( .A(n51645), .B(n51646), .Z(n51644) );
  NAND U52078 ( .A(n51646), .B(n51645), .Z(n51641) );
  ANDN U52079 ( .B(B[74]), .A(n57), .Z(n51425) );
  XNOR U52080 ( .A(n51433), .B(n51647), .Z(n51426) );
  XNOR U52081 ( .A(n51432), .B(n51430), .Z(n51647) );
  AND U52082 ( .A(n51648), .B(n51649), .Z(n51430) );
  NANDN U52083 ( .A(n51650), .B(n51651), .Z(n51649) );
  NANDN U52084 ( .A(n51652), .B(n51653), .Z(n51651) );
  NANDN U52085 ( .A(n51653), .B(n51652), .Z(n51648) );
  ANDN U52086 ( .B(B[75]), .A(n58), .Z(n51432) );
  XNOR U52087 ( .A(n51440), .B(n51654), .Z(n51433) );
  XNOR U52088 ( .A(n51439), .B(n51437), .Z(n51654) );
  AND U52089 ( .A(n51655), .B(n51656), .Z(n51437) );
  NANDN U52090 ( .A(n51657), .B(n51658), .Z(n51656) );
  OR U52091 ( .A(n51659), .B(n51660), .Z(n51658) );
  NAND U52092 ( .A(n51660), .B(n51659), .Z(n51655) );
  ANDN U52093 ( .B(B[76]), .A(n59), .Z(n51439) );
  XNOR U52094 ( .A(n51447), .B(n51661), .Z(n51440) );
  XNOR U52095 ( .A(n51446), .B(n51444), .Z(n51661) );
  AND U52096 ( .A(n51662), .B(n51663), .Z(n51444) );
  NANDN U52097 ( .A(n51664), .B(n51665), .Z(n51663) );
  NANDN U52098 ( .A(n51666), .B(n51667), .Z(n51665) );
  NANDN U52099 ( .A(n51667), .B(n51666), .Z(n51662) );
  ANDN U52100 ( .B(B[77]), .A(n60), .Z(n51446) );
  XNOR U52101 ( .A(n51454), .B(n51668), .Z(n51447) );
  XNOR U52102 ( .A(n51453), .B(n51451), .Z(n51668) );
  AND U52103 ( .A(n51669), .B(n51670), .Z(n51451) );
  NANDN U52104 ( .A(n51671), .B(n51672), .Z(n51670) );
  OR U52105 ( .A(n51673), .B(n51674), .Z(n51672) );
  NAND U52106 ( .A(n51674), .B(n51673), .Z(n51669) );
  ANDN U52107 ( .B(B[78]), .A(n61), .Z(n51453) );
  XNOR U52108 ( .A(n51461), .B(n51675), .Z(n51454) );
  XNOR U52109 ( .A(n51460), .B(n51458), .Z(n51675) );
  AND U52110 ( .A(n51676), .B(n51677), .Z(n51458) );
  NANDN U52111 ( .A(n51678), .B(n51679), .Z(n51677) );
  NANDN U52112 ( .A(n51680), .B(n51681), .Z(n51679) );
  NANDN U52113 ( .A(n51681), .B(n51680), .Z(n51676) );
  ANDN U52114 ( .B(B[79]), .A(n62), .Z(n51460) );
  XNOR U52115 ( .A(n51468), .B(n51682), .Z(n51461) );
  XNOR U52116 ( .A(n51467), .B(n51465), .Z(n51682) );
  AND U52117 ( .A(n51683), .B(n51684), .Z(n51465) );
  NANDN U52118 ( .A(n51685), .B(n51686), .Z(n51684) );
  OR U52119 ( .A(n51687), .B(n51688), .Z(n51686) );
  NAND U52120 ( .A(n51688), .B(n51687), .Z(n51683) );
  ANDN U52121 ( .B(B[80]), .A(n63), .Z(n51467) );
  XNOR U52122 ( .A(n51475), .B(n51689), .Z(n51468) );
  XNOR U52123 ( .A(n51474), .B(n51472), .Z(n51689) );
  AND U52124 ( .A(n51690), .B(n51691), .Z(n51472) );
  NANDN U52125 ( .A(n51692), .B(n51693), .Z(n51691) );
  NANDN U52126 ( .A(n51694), .B(n51695), .Z(n51693) );
  NANDN U52127 ( .A(n51695), .B(n51694), .Z(n51690) );
  ANDN U52128 ( .B(B[81]), .A(n64), .Z(n51474) );
  XNOR U52129 ( .A(n51482), .B(n51696), .Z(n51475) );
  XNOR U52130 ( .A(n51481), .B(n51479), .Z(n51696) );
  AND U52131 ( .A(n51697), .B(n51698), .Z(n51479) );
  NANDN U52132 ( .A(n51699), .B(n51700), .Z(n51698) );
  OR U52133 ( .A(n51701), .B(n51702), .Z(n51700) );
  NAND U52134 ( .A(n51702), .B(n51701), .Z(n51697) );
  ANDN U52135 ( .B(B[82]), .A(n65), .Z(n51481) );
  XNOR U52136 ( .A(n51489), .B(n51703), .Z(n51482) );
  XNOR U52137 ( .A(n51488), .B(n51486), .Z(n51703) );
  AND U52138 ( .A(n51704), .B(n51705), .Z(n51486) );
  NANDN U52139 ( .A(n51706), .B(n51707), .Z(n51705) );
  NANDN U52140 ( .A(n51708), .B(n51709), .Z(n51707) );
  NANDN U52141 ( .A(n51709), .B(n51708), .Z(n51704) );
  ANDN U52142 ( .B(B[83]), .A(n66), .Z(n51488) );
  XNOR U52143 ( .A(n51496), .B(n51710), .Z(n51489) );
  XNOR U52144 ( .A(n51495), .B(n51493), .Z(n51710) );
  AND U52145 ( .A(n51711), .B(n51712), .Z(n51493) );
  NANDN U52146 ( .A(n51713), .B(n51714), .Z(n51712) );
  OR U52147 ( .A(n51715), .B(n51716), .Z(n51714) );
  NAND U52148 ( .A(n51716), .B(n51715), .Z(n51711) );
  ANDN U52149 ( .B(B[84]), .A(n67), .Z(n51495) );
  XNOR U52150 ( .A(n51503), .B(n51717), .Z(n51496) );
  XNOR U52151 ( .A(n51502), .B(n51500), .Z(n51717) );
  AND U52152 ( .A(n51718), .B(n51719), .Z(n51500) );
  NANDN U52153 ( .A(n51720), .B(n51721), .Z(n51719) );
  NANDN U52154 ( .A(n51722), .B(n51723), .Z(n51721) );
  NANDN U52155 ( .A(n51723), .B(n51722), .Z(n51718) );
  ANDN U52156 ( .B(A[17]), .A(n33), .Z(n51502) );
  XNOR U52157 ( .A(n51510), .B(n51724), .Z(n51503) );
  XNOR U52158 ( .A(n51509), .B(n51507), .Z(n51724) );
  AND U52159 ( .A(n51725), .B(n51726), .Z(n51507) );
  NANDN U52160 ( .A(n51727), .B(n51728), .Z(n51726) );
  OR U52161 ( .A(n51729), .B(n51730), .Z(n51728) );
  NAND U52162 ( .A(n51730), .B(n51729), .Z(n51725) );
  ANDN U52163 ( .B(A[16]), .A(n31), .Z(n51509) );
  XNOR U52164 ( .A(n51517), .B(n51731), .Z(n51510) );
  XNOR U52165 ( .A(n51516), .B(n51514), .Z(n51731) );
  AND U52166 ( .A(n51732), .B(n51733), .Z(n51514) );
  NANDN U52167 ( .A(n51734), .B(n51735), .Z(n51733) );
  NANDN U52168 ( .A(n51736), .B(n51737), .Z(n51735) );
  NANDN U52169 ( .A(n51737), .B(n51736), .Z(n51732) );
  ANDN U52170 ( .B(A[15]), .A(n29), .Z(n51516) );
  XNOR U52171 ( .A(n51524), .B(n51738), .Z(n51517) );
  XNOR U52172 ( .A(n51523), .B(n51521), .Z(n51738) );
  AND U52173 ( .A(n51739), .B(n51740), .Z(n51521) );
  NANDN U52174 ( .A(n51741), .B(n51742), .Z(n51740) );
  OR U52175 ( .A(n51743), .B(n51744), .Z(n51742) );
  NAND U52176 ( .A(n51744), .B(n51743), .Z(n51739) );
  ANDN U52177 ( .B(A[14]), .A(n27), .Z(n51523) );
  XNOR U52178 ( .A(n51531), .B(n51745), .Z(n51524) );
  XNOR U52179 ( .A(n51530), .B(n51528), .Z(n51745) );
  AND U52180 ( .A(n51746), .B(n51747), .Z(n51528) );
  NANDN U52181 ( .A(n51748), .B(n51749), .Z(n51747) );
  NANDN U52182 ( .A(n51750), .B(n51751), .Z(n51749) );
  NANDN U52183 ( .A(n51751), .B(n51750), .Z(n51746) );
  ANDN U52184 ( .B(A[13]), .A(n25), .Z(n51530) );
  XNOR U52185 ( .A(n51538), .B(n51752), .Z(n51531) );
  XNOR U52186 ( .A(n51537), .B(n51535), .Z(n51752) );
  AND U52187 ( .A(n51753), .B(n51754), .Z(n51535) );
  NANDN U52188 ( .A(n51755), .B(n51756), .Z(n51754) );
  OR U52189 ( .A(n51757), .B(n51758), .Z(n51756) );
  NAND U52190 ( .A(n51758), .B(n51757), .Z(n51753) );
  ANDN U52191 ( .B(A[12]), .A(n23), .Z(n51537) );
  XNOR U52192 ( .A(n51545), .B(n51759), .Z(n51538) );
  XNOR U52193 ( .A(n51544), .B(n51542), .Z(n51759) );
  AND U52194 ( .A(n51760), .B(n51761), .Z(n51542) );
  NANDN U52195 ( .A(n51762), .B(n51763), .Z(n51761) );
  NANDN U52196 ( .A(n51764), .B(n51765), .Z(n51763) );
  NANDN U52197 ( .A(n51765), .B(n51764), .Z(n51760) );
  ANDN U52198 ( .B(A[11]), .A(n21), .Z(n51544) );
  XNOR U52199 ( .A(n51552), .B(n51766), .Z(n51545) );
  XNOR U52200 ( .A(n51551), .B(n51549), .Z(n51766) );
  AND U52201 ( .A(n51767), .B(n51768), .Z(n51549) );
  NANDN U52202 ( .A(n51769), .B(n51770), .Z(n51768) );
  OR U52203 ( .A(n51771), .B(n51772), .Z(n51770) );
  NAND U52204 ( .A(n51772), .B(n51771), .Z(n51767) );
  ANDN U52205 ( .B(A[10]), .A(n19), .Z(n51551) );
  XNOR U52206 ( .A(n51559), .B(n51773), .Z(n51552) );
  XNOR U52207 ( .A(n51558), .B(n51556), .Z(n51773) );
  AND U52208 ( .A(n51774), .B(n51775), .Z(n51556) );
  NANDN U52209 ( .A(n51776), .B(n51777), .Z(n51775) );
  NANDN U52210 ( .A(n51778), .B(n51779), .Z(n51777) );
  NANDN U52211 ( .A(n51779), .B(n51778), .Z(n51774) );
  ANDN U52212 ( .B(A[9]), .A(n17), .Z(n51558) );
  XNOR U52213 ( .A(n51566), .B(n51780), .Z(n51559) );
  XNOR U52214 ( .A(n51565), .B(n51563), .Z(n51780) );
  AND U52215 ( .A(n51781), .B(n51782), .Z(n51563) );
  NANDN U52216 ( .A(n51783), .B(n51784), .Z(n51782) );
  OR U52217 ( .A(n51785), .B(n51786), .Z(n51784) );
  NAND U52218 ( .A(n51786), .B(n51785), .Z(n51781) );
  ANDN U52219 ( .B(A[8]), .A(n15), .Z(n51565) );
  XNOR U52220 ( .A(n51573), .B(n51787), .Z(n51566) );
  XNOR U52221 ( .A(n51572), .B(n51570), .Z(n51787) );
  AND U52222 ( .A(n51788), .B(n51789), .Z(n51570) );
  NANDN U52223 ( .A(n51790), .B(n51791), .Z(n51789) );
  NANDN U52224 ( .A(n51792), .B(n51793), .Z(n51791) );
  NANDN U52225 ( .A(n51793), .B(n51792), .Z(n51788) );
  ANDN U52226 ( .B(A[7]), .A(n13), .Z(n51572) );
  XNOR U52227 ( .A(n51580), .B(n51794), .Z(n51573) );
  XNOR U52228 ( .A(n51579), .B(n51577), .Z(n51794) );
  AND U52229 ( .A(n51795), .B(n51796), .Z(n51577) );
  NANDN U52230 ( .A(n51797), .B(n51798), .Z(n51796) );
  OR U52231 ( .A(n51799), .B(n51800), .Z(n51798) );
  NAND U52232 ( .A(n51800), .B(n51799), .Z(n51795) );
  ANDN U52233 ( .B(A[6]), .A(n11), .Z(n51579) );
  XNOR U52234 ( .A(n51587), .B(n51801), .Z(n51580) );
  XNOR U52235 ( .A(n51586), .B(n51584), .Z(n51801) );
  AND U52236 ( .A(n51802), .B(n51803), .Z(n51584) );
  NANDN U52237 ( .A(n51804), .B(n51805), .Z(n51803) );
  NANDN U52238 ( .A(n51806), .B(n51807), .Z(n51805) );
  NANDN U52239 ( .A(n51807), .B(n51806), .Z(n51802) );
  ANDN U52240 ( .B(A[5]), .A(n9), .Z(n51586) );
  XNOR U52241 ( .A(n51594), .B(n51808), .Z(n51587) );
  XNOR U52242 ( .A(n51593), .B(n51591), .Z(n51808) );
  AND U52243 ( .A(n51809), .B(n51810), .Z(n51591) );
  NANDN U52244 ( .A(n51811), .B(n51812), .Z(n51810) );
  OR U52245 ( .A(n51813), .B(n51814), .Z(n51812) );
  NAND U52246 ( .A(n51814), .B(n51813), .Z(n51809) );
  ANDN U52247 ( .B(B[98]), .A(n81), .Z(n51593) );
  XNOR U52248 ( .A(n51601), .B(n51815), .Z(n51594) );
  XNOR U52249 ( .A(n51600), .B(n51598), .Z(n51815) );
  AND U52250 ( .A(n51816), .B(n51817), .Z(n51598) );
  NANDN U52251 ( .A(n51818), .B(n51819), .Z(n51817) );
  NAND U52252 ( .A(n51820), .B(n51821), .Z(n51819) );
  ANDN U52253 ( .B(A[3]), .A(n6), .Z(n51600) );
  XOR U52254 ( .A(n51607), .B(n51822), .Z(n51601) );
  XNOR U52255 ( .A(n51605), .B(n51608), .Z(n51822) );
  NAND U52256 ( .A(B[100]), .B(A[2]), .Z(n51608) );
  NANDN U52257 ( .A(n51823), .B(n51824), .Z(n51605) );
  AND U52258 ( .A(A[0]), .B(B[101]), .Z(n51824) );
  XNOR U52259 ( .A(n51610), .B(n51825), .Z(n51607) );
  NAND U52260 ( .A(A[0]), .B(B[102]), .Z(n51825) );
  NAND U52261 ( .A(B[101]), .B(A[1]), .Z(n51610) );
  NAND U52262 ( .A(n51826), .B(n51827), .Z(n592) );
  NANDN U52263 ( .A(n600), .B(n51828), .Z(n51827) );
  NANDN U52264 ( .A(n598), .B(n51829), .Z(n51828) );
  NAND U52265 ( .A(A[31]), .B(B[70]), .Z(n600) );
  NAND U52266 ( .A(n5), .B(n598), .Z(n51826) );
  XOR U52267 ( .A(n51625), .B(n51830), .Z(n598) );
  XNOR U52268 ( .A(n51624), .B(n51622), .Z(n51830) );
  AND U52269 ( .A(n51831), .B(n51832), .Z(n51622) );
  NANDN U52270 ( .A(n51833), .B(n51834), .Z(n51832) );
  OR U52271 ( .A(n51835), .B(n51836), .Z(n51834) );
  NAND U52272 ( .A(n51836), .B(n51835), .Z(n51831) );
  ANDN U52273 ( .B(B[71]), .A(n55), .Z(n51624) );
  XOR U52274 ( .A(n51632), .B(n51837), .Z(n51625) );
  XNOR U52275 ( .A(n51631), .B(n51629), .Z(n51837) );
  AND U52276 ( .A(n51838), .B(n51839), .Z(n51629) );
  NANDN U52277 ( .A(n51840), .B(n51841), .Z(n51839) );
  NANDN U52278 ( .A(n51842), .B(n51843), .Z(n51841) );
  ANDN U52279 ( .B(B[72]), .A(n56), .Z(n51631) );
  XNOR U52280 ( .A(n51639), .B(n51844), .Z(n51632) );
  XNOR U52281 ( .A(n51638), .B(n51636), .Z(n51844) );
  AND U52282 ( .A(n51845), .B(n51846), .Z(n51636) );
  NANDN U52283 ( .A(n51847), .B(n51848), .Z(n51846) );
  OR U52284 ( .A(n51849), .B(n51850), .Z(n51848) );
  NAND U52285 ( .A(n51850), .B(n51849), .Z(n51845) );
  ANDN U52286 ( .B(B[73]), .A(n57), .Z(n51638) );
  XNOR U52287 ( .A(n51646), .B(n51851), .Z(n51639) );
  XNOR U52288 ( .A(n51645), .B(n51643), .Z(n51851) );
  AND U52289 ( .A(n51852), .B(n51853), .Z(n51643) );
  NANDN U52290 ( .A(n51854), .B(n51855), .Z(n51853) );
  NANDN U52291 ( .A(n51856), .B(n51857), .Z(n51855) );
  ANDN U52292 ( .B(B[74]), .A(n58), .Z(n51645) );
  XNOR U52293 ( .A(n51653), .B(n51858), .Z(n51646) );
  XNOR U52294 ( .A(n51652), .B(n51650), .Z(n51858) );
  AND U52295 ( .A(n51859), .B(n51860), .Z(n51650) );
  NANDN U52296 ( .A(n51861), .B(n51862), .Z(n51860) );
  OR U52297 ( .A(n51863), .B(n51864), .Z(n51862) );
  NAND U52298 ( .A(n51864), .B(n51863), .Z(n51859) );
  ANDN U52299 ( .B(B[75]), .A(n59), .Z(n51652) );
  XNOR U52300 ( .A(n51660), .B(n51865), .Z(n51653) );
  XNOR U52301 ( .A(n51659), .B(n51657), .Z(n51865) );
  AND U52302 ( .A(n51866), .B(n51867), .Z(n51657) );
  NANDN U52303 ( .A(n51868), .B(n51869), .Z(n51867) );
  NANDN U52304 ( .A(n51870), .B(n51871), .Z(n51869) );
  ANDN U52305 ( .B(B[76]), .A(n60), .Z(n51659) );
  XNOR U52306 ( .A(n51667), .B(n51872), .Z(n51660) );
  XNOR U52307 ( .A(n51666), .B(n51664), .Z(n51872) );
  AND U52308 ( .A(n51873), .B(n51874), .Z(n51664) );
  NANDN U52309 ( .A(n51875), .B(n51876), .Z(n51874) );
  OR U52310 ( .A(n51877), .B(n51878), .Z(n51876) );
  NAND U52311 ( .A(n51878), .B(n51877), .Z(n51873) );
  ANDN U52312 ( .B(B[77]), .A(n61), .Z(n51666) );
  XNOR U52313 ( .A(n51674), .B(n51879), .Z(n51667) );
  XNOR U52314 ( .A(n51673), .B(n51671), .Z(n51879) );
  AND U52315 ( .A(n51880), .B(n51881), .Z(n51671) );
  NANDN U52316 ( .A(n51882), .B(n51883), .Z(n51881) );
  NANDN U52317 ( .A(n51884), .B(n51885), .Z(n51883) );
  ANDN U52318 ( .B(B[78]), .A(n62), .Z(n51673) );
  XNOR U52319 ( .A(n51681), .B(n51886), .Z(n51674) );
  XNOR U52320 ( .A(n51680), .B(n51678), .Z(n51886) );
  AND U52321 ( .A(n51887), .B(n51888), .Z(n51678) );
  NANDN U52322 ( .A(n51889), .B(n51890), .Z(n51888) );
  OR U52323 ( .A(n51891), .B(n51892), .Z(n51890) );
  NAND U52324 ( .A(n51892), .B(n51891), .Z(n51887) );
  ANDN U52325 ( .B(B[79]), .A(n63), .Z(n51680) );
  XNOR U52326 ( .A(n51688), .B(n51893), .Z(n51681) );
  XNOR U52327 ( .A(n51687), .B(n51685), .Z(n51893) );
  AND U52328 ( .A(n51894), .B(n51895), .Z(n51685) );
  NANDN U52329 ( .A(n51896), .B(n51897), .Z(n51895) );
  NANDN U52330 ( .A(n51898), .B(n51899), .Z(n51897) );
  ANDN U52331 ( .B(B[80]), .A(n64), .Z(n51687) );
  XNOR U52332 ( .A(n51695), .B(n51900), .Z(n51688) );
  XNOR U52333 ( .A(n51694), .B(n51692), .Z(n51900) );
  AND U52334 ( .A(n51901), .B(n51902), .Z(n51692) );
  NANDN U52335 ( .A(n51903), .B(n51904), .Z(n51902) );
  OR U52336 ( .A(n51905), .B(n51906), .Z(n51904) );
  NAND U52337 ( .A(n51906), .B(n51905), .Z(n51901) );
  ANDN U52338 ( .B(B[81]), .A(n65), .Z(n51694) );
  XNOR U52339 ( .A(n51702), .B(n51907), .Z(n51695) );
  XNOR U52340 ( .A(n51701), .B(n51699), .Z(n51907) );
  AND U52341 ( .A(n51908), .B(n51909), .Z(n51699) );
  NANDN U52342 ( .A(n51910), .B(n51911), .Z(n51909) );
  NANDN U52343 ( .A(n51912), .B(n51913), .Z(n51911) );
  ANDN U52344 ( .B(B[82]), .A(n66), .Z(n51701) );
  XNOR U52345 ( .A(n51709), .B(n51914), .Z(n51702) );
  XNOR U52346 ( .A(n51708), .B(n51706), .Z(n51914) );
  AND U52347 ( .A(n51915), .B(n51916), .Z(n51706) );
  NANDN U52348 ( .A(n51917), .B(n51918), .Z(n51916) );
  OR U52349 ( .A(n51919), .B(n51920), .Z(n51918) );
  NAND U52350 ( .A(n51920), .B(n51919), .Z(n51915) );
  ANDN U52351 ( .B(B[83]), .A(n67), .Z(n51708) );
  XNOR U52352 ( .A(n51716), .B(n51921), .Z(n51709) );
  XNOR U52353 ( .A(n51715), .B(n51713), .Z(n51921) );
  AND U52354 ( .A(n51922), .B(n51923), .Z(n51713) );
  NANDN U52355 ( .A(n51924), .B(n51925), .Z(n51923) );
  NANDN U52356 ( .A(n51926), .B(n51927), .Z(n51925) );
  ANDN U52357 ( .B(B[84]), .A(n68), .Z(n51715) );
  XNOR U52358 ( .A(n51723), .B(n51928), .Z(n51716) );
  XNOR U52359 ( .A(n51722), .B(n51720), .Z(n51928) );
  AND U52360 ( .A(n51929), .B(n51930), .Z(n51720) );
  NANDN U52361 ( .A(n51931), .B(n51932), .Z(n51930) );
  OR U52362 ( .A(n51933), .B(n51934), .Z(n51932) );
  NAND U52363 ( .A(n51934), .B(n51933), .Z(n51929) );
  ANDN U52364 ( .B(A[16]), .A(n33), .Z(n51722) );
  XNOR U52365 ( .A(n51730), .B(n51935), .Z(n51723) );
  XNOR U52366 ( .A(n51729), .B(n51727), .Z(n51935) );
  AND U52367 ( .A(n51936), .B(n51937), .Z(n51727) );
  NANDN U52368 ( .A(n51938), .B(n51939), .Z(n51937) );
  NANDN U52369 ( .A(n51940), .B(n51941), .Z(n51939) );
  ANDN U52370 ( .B(A[15]), .A(n31), .Z(n51729) );
  XNOR U52371 ( .A(n51737), .B(n51942), .Z(n51730) );
  XNOR U52372 ( .A(n51736), .B(n51734), .Z(n51942) );
  AND U52373 ( .A(n51943), .B(n51944), .Z(n51734) );
  NANDN U52374 ( .A(n51945), .B(n51946), .Z(n51944) );
  OR U52375 ( .A(n51947), .B(n51948), .Z(n51946) );
  NAND U52376 ( .A(n51948), .B(n51947), .Z(n51943) );
  ANDN U52377 ( .B(A[14]), .A(n29), .Z(n51736) );
  XNOR U52378 ( .A(n51744), .B(n51949), .Z(n51737) );
  XNOR U52379 ( .A(n51743), .B(n51741), .Z(n51949) );
  AND U52380 ( .A(n51950), .B(n51951), .Z(n51741) );
  NANDN U52381 ( .A(n51952), .B(n51953), .Z(n51951) );
  NANDN U52382 ( .A(n51954), .B(n51955), .Z(n51953) );
  ANDN U52383 ( .B(A[13]), .A(n27), .Z(n51743) );
  XNOR U52384 ( .A(n51751), .B(n51956), .Z(n51744) );
  XNOR U52385 ( .A(n51750), .B(n51748), .Z(n51956) );
  AND U52386 ( .A(n51957), .B(n51958), .Z(n51748) );
  NANDN U52387 ( .A(n51959), .B(n51960), .Z(n51958) );
  OR U52388 ( .A(n51961), .B(n51962), .Z(n51960) );
  NAND U52389 ( .A(n51962), .B(n51961), .Z(n51957) );
  ANDN U52390 ( .B(A[12]), .A(n25), .Z(n51750) );
  XNOR U52391 ( .A(n51758), .B(n51963), .Z(n51751) );
  XNOR U52392 ( .A(n51757), .B(n51755), .Z(n51963) );
  AND U52393 ( .A(n51964), .B(n51965), .Z(n51755) );
  NANDN U52394 ( .A(n51966), .B(n51967), .Z(n51965) );
  NANDN U52395 ( .A(n51968), .B(n51969), .Z(n51967) );
  ANDN U52396 ( .B(A[11]), .A(n23), .Z(n51757) );
  XNOR U52397 ( .A(n51765), .B(n51970), .Z(n51758) );
  XNOR U52398 ( .A(n51764), .B(n51762), .Z(n51970) );
  AND U52399 ( .A(n51971), .B(n51972), .Z(n51762) );
  NANDN U52400 ( .A(n51973), .B(n51974), .Z(n51972) );
  OR U52401 ( .A(n51975), .B(n51976), .Z(n51974) );
  NAND U52402 ( .A(n51976), .B(n51975), .Z(n51971) );
  ANDN U52403 ( .B(A[10]), .A(n21), .Z(n51764) );
  XNOR U52404 ( .A(n51772), .B(n51977), .Z(n51765) );
  XNOR U52405 ( .A(n51771), .B(n51769), .Z(n51977) );
  AND U52406 ( .A(n51978), .B(n51979), .Z(n51769) );
  NANDN U52407 ( .A(n51980), .B(n51981), .Z(n51979) );
  NANDN U52408 ( .A(n51982), .B(n51983), .Z(n51981) );
  ANDN U52409 ( .B(A[9]), .A(n19), .Z(n51771) );
  XNOR U52410 ( .A(n51779), .B(n51984), .Z(n51772) );
  XNOR U52411 ( .A(n51778), .B(n51776), .Z(n51984) );
  AND U52412 ( .A(n51985), .B(n51986), .Z(n51776) );
  NANDN U52413 ( .A(n51987), .B(n51988), .Z(n51986) );
  OR U52414 ( .A(n51989), .B(n51990), .Z(n51988) );
  NAND U52415 ( .A(n51990), .B(n51989), .Z(n51985) );
  ANDN U52416 ( .B(A[8]), .A(n17), .Z(n51778) );
  XNOR U52417 ( .A(n51786), .B(n51991), .Z(n51779) );
  XNOR U52418 ( .A(n51785), .B(n51783), .Z(n51991) );
  AND U52419 ( .A(n51992), .B(n51993), .Z(n51783) );
  NANDN U52420 ( .A(n51994), .B(n51995), .Z(n51993) );
  NANDN U52421 ( .A(n51996), .B(n51997), .Z(n51995) );
  ANDN U52422 ( .B(A[7]), .A(n15), .Z(n51785) );
  XNOR U52423 ( .A(n51793), .B(n51998), .Z(n51786) );
  XNOR U52424 ( .A(n51792), .B(n51790), .Z(n51998) );
  AND U52425 ( .A(n51999), .B(n52000), .Z(n51790) );
  NANDN U52426 ( .A(n52001), .B(n52002), .Z(n52000) );
  OR U52427 ( .A(n52003), .B(n52004), .Z(n52002) );
  NAND U52428 ( .A(n52004), .B(n52003), .Z(n51999) );
  ANDN U52429 ( .B(A[6]), .A(n13), .Z(n51792) );
  XNOR U52430 ( .A(n51800), .B(n52005), .Z(n51793) );
  XNOR U52431 ( .A(n51799), .B(n51797), .Z(n52005) );
  AND U52432 ( .A(n52006), .B(n52007), .Z(n51797) );
  NANDN U52433 ( .A(n52008), .B(n52009), .Z(n52007) );
  NANDN U52434 ( .A(n52010), .B(n52011), .Z(n52009) );
  ANDN U52435 ( .B(A[5]), .A(n11), .Z(n51799) );
  XNOR U52436 ( .A(n51807), .B(n52012), .Z(n51800) );
  XNOR U52437 ( .A(n51806), .B(n51804), .Z(n52012) );
  AND U52438 ( .A(n52013), .B(n52014), .Z(n51804) );
  NANDN U52439 ( .A(n52015), .B(n52016), .Z(n52014) );
  OR U52440 ( .A(n52017), .B(n52018), .Z(n52016) );
  NAND U52441 ( .A(n52018), .B(n52017), .Z(n52013) );
  ANDN U52442 ( .B(A[4]), .A(n9), .Z(n51806) );
  XNOR U52443 ( .A(n51814), .B(n52019), .Z(n51807) );
  XNOR U52444 ( .A(n51813), .B(n51811), .Z(n52019) );
  AND U52445 ( .A(n52020), .B(n52021), .Z(n51811) );
  NANDN U52446 ( .A(n52022), .B(n52023), .Z(n52021) );
  NANDN U52447 ( .A(n52024), .B(n52025), .Z(n52023) );
  NANDN U52448 ( .A(n52025), .B(n52024), .Z(n52020) );
  ANDN U52449 ( .B(B[98]), .A(n82), .Z(n51813) );
  XOR U52450 ( .A(n51820), .B(n52026), .Z(n51814) );
  XNOR U52451 ( .A(n51818), .B(n51821), .Z(n52026) );
  NAND U52452 ( .A(B[99]), .B(A[2]), .Z(n51821) );
  NANDN U52453 ( .A(n52027), .B(n52028), .Z(n51818) );
  AND U52454 ( .A(A[0]), .B(B[100]), .Z(n52028) );
  XNOR U52455 ( .A(n51823), .B(n52029), .Z(n51820) );
  NAND U52456 ( .A(A[0]), .B(B[101]), .Z(n52029) );
  NAND U52457 ( .A(B[100]), .B(A[1]), .Z(n51823) );
  AND U52458 ( .A(n52030), .B(n52031), .Z(n51829) );
  NANDN U52459 ( .A(n616), .B(n52032), .Z(n52031) );
  NAND U52460 ( .A(n617), .B(n614), .Z(n52032) );
  NAND U52461 ( .A(A[30]), .B(B[70]), .Z(n616) );
  AND U52462 ( .A(n52033), .B(n52034), .Z(n617) );
  NANDN U52463 ( .A(n640), .B(n52035), .Z(n52034) );
  NANDN U52464 ( .A(n638), .B(n52036), .Z(n52035) );
  NAND U52465 ( .A(A[29]), .B(B[70]), .Z(n640) );
  NAND U52466 ( .A(n7), .B(n638), .Z(n52033) );
  XOR U52467 ( .A(n52037), .B(n52038), .Z(n638) );
  XNOR U52468 ( .A(n52039), .B(n52040), .Z(n52038) );
  AND U52469 ( .A(n52041), .B(n52042), .Z(n52036) );
  NANDN U52470 ( .A(n670), .B(n52043), .Z(n52042) );
  NANDN U52471 ( .A(n668), .B(n52044), .Z(n52043) );
  NAND U52472 ( .A(A[28]), .B(B[70]), .Z(n670) );
  NAND U52473 ( .A(n8), .B(n668), .Z(n52041) );
  XOR U52474 ( .A(n52045), .B(n52046), .Z(n668) );
  XNOR U52475 ( .A(n52047), .B(n52048), .Z(n52046) );
  AND U52476 ( .A(n52049), .B(n52050), .Z(n52044) );
  NANDN U52477 ( .A(n707), .B(n52051), .Z(n52050) );
  NANDN U52478 ( .A(n705), .B(n52052), .Z(n52051) );
  NAND U52479 ( .A(A[27]), .B(B[70]), .Z(n707) );
  NAND U52480 ( .A(n10), .B(n705), .Z(n52049) );
  XOR U52481 ( .A(n52053), .B(n52054), .Z(n705) );
  XNOR U52482 ( .A(n52055), .B(n52056), .Z(n52054) );
  AND U52483 ( .A(n52057), .B(n52058), .Z(n52052) );
  NANDN U52484 ( .A(n751), .B(n52059), .Z(n52058) );
  NANDN U52485 ( .A(n749), .B(n52060), .Z(n52059) );
  NAND U52486 ( .A(A[26]), .B(B[70]), .Z(n751) );
  NAND U52487 ( .A(n12), .B(n749), .Z(n52057) );
  XOR U52488 ( .A(n52061), .B(n52062), .Z(n749) );
  XNOR U52489 ( .A(n52063), .B(n52064), .Z(n52062) );
  AND U52490 ( .A(n52065), .B(n52066), .Z(n52060) );
  NANDN U52491 ( .A(n802), .B(n52067), .Z(n52066) );
  NANDN U52492 ( .A(n800), .B(n52068), .Z(n52067) );
  NAND U52493 ( .A(A[25]), .B(B[70]), .Z(n802) );
  NAND U52494 ( .A(n14), .B(n800), .Z(n52065) );
  XOR U52495 ( .A(n52069), .B(n52070), .Z(n800) );
  XNOR U52496 ( .A(n52071), .B(n52072), .Z(n52070) );
  AND U52497 ( .A(n52073), .B(n52074), .Z(n52068) );
  NANDN U52498 ( .A(n860), .B(n52075), .Z(n52074) );
  NANDN U52499 ( .A(n858), .B(n52076), .Z(n52075) );
  NAND U52500 ( .A(A[24]), .B(B[70]), .Z(n860) );
  NAND U52501 ( .A(n16), .B(n858), .Z(n52073) );
  XOR U52502 ( .A(n52077), .B(n52078), .Z(n858) );
  XNOR U52503 ( .A(n52079), .B(n52080), .Z(n52078) );
  AND U52504 ( .A(n52081), .B(n52082), .Z(n52076) );
  NANDN U52505 ( .A(n925), .B(n52083), .Z(n52082) );
  NANDN U52506 ( .A(n923), .B(n52084), .Z(n52083) );
  NAND U52507 ( .A(A[23]), .B(B[70]), .Z(n925) );
  NAND U52508 ( .A(n18), .B(n923), .Z(n52081) );
  XOR U52509 ( .A(n52085), .B(n52086), .Z(n923) );
  XNOR U52510 ( .A(n52087), .B(n52088), .Z(n52086) );
  AND U52511 ( .A(n52089), .B(n52090), .Z(n52084) );
  NANDN U52512 ( .A(n997), .B(n52091), .Z(n52090) );
  NANDN U52513 ( .A(n995), .B(n52092), .Z(n52091) );
  NAND U52514 ( .A(A[22]), .B(B[70]), .Z(n997) );
  NAND U52515 ( .A(n20), .B(n995), .Z(n52089) );
  XOR U52516 ( .A(n52093), .B(n52094), .Z(n995) );
  XNOR U52517 ( .A(n52095), .B(n52096), .Z(n52094) );
  AND U52518 ( .A(n52097), .B(n52098), .Z(n52092) );
  NANDN U52519 ( .A(n1080), .B(n52099), .Z(n52098) );
  NANDN U52520 ( .A(n1078), .B(n52100), .Z(n52099) );
  NAND U52521 ( .A(A[21]), .B(B[70]), .Z(n1080) );
  NAND U52522 ( .A(n22), .B(n1078), .Z(n52097) );
  XOR U52523 ( .A(n52101), .B(n52102), .Z(n1078) );
  XNOR U52524 ( .A(n52103), .B(n52104), .Z(n52102) );
  AND U52525 ( .A(n52105), .B(n52106), .Z(n52100) );
  NANDN U52526 ( .A(n1166), .B(n52107), .Z(n52106) );
  NANDN U52527 ( .A(n1164), .B(n52108), .Z(n52107) );
  NAND U52528 ( .A(A[20]), .B(B[70]), .Z(n1166) );
  NAND U52529 ( .A(n24), .B(n1164), .Z(n52105) );
  XOR U52530 ( .A(n52109), .B(n52110), .Z(n1164) );
  XNOR U52531 ( .A(n52111), .B(n52112), .Z(n52110) );
  AND U52532 ( .A(n52113), .B(n52114), .Z(n52108) );
  NANDN U52533 ( .A(n1259), .B(n52115), .Z(n52114) );
  NANDN U52534 ( .A(n1257), .B(n52116), .Z(n52115) );
  NAND U52535 ( .A(A[19]), .B(B[70]), .Z(n1259) );
  NAND U52536 ( .A(n26), .B(n1257), .Z(n52113) );
  XOR U52537 ( .A(n52117), .B(n52118), .Z(n1257) );
  XNOR U52538 ( .A(n52119), .B(n52120), .Z(n52118) );
  AND U52539 ( .A(n52121), .B(n52122), .Z(n52116) );
  NANDN U52540 ( .A(n1359), .B(n52123), .Z(n52122) );
  NANDN U52541 ( .A(n1357), .B(n52124), .Z(n52123) );
  NAND U52542 ( .A(A[18]), .B(B[70]), .Z(n1359) );
  NAND U52543 ( .A(n28), .B(n1357), .Z(n52121) );
  XOR U52544 ( .A(n52125), .B(n52126), .Z(n1357) );
  XNOR U52545 ( .A(n52127), .B(n52128), .Z(n52126) );
  AND U52546 ( .A(n52129), .B(n52130), .Z(n52124) );
  NANDN U52547 ( .A(n1466), .B(n52131), .Z(n52130) );
  NANDN U52548 ( .A(n1464), .B(n52132), .Z(n52131) );
  NAND U52549 ( .A(A[17]), .B(B[70]), .Z(n1466) );
  NAND U52550 ( .A(n30), .B(n1464), .Z(n52129) );
  XOR U52551 ( .A(n52133), .B(n52134), .Z(n1464) );
  XNOR U52552 ( .A(n52135), .B(n52136), .Z(n52134) );
  AND U52553 ( .A(n52137), .B(n52138), .Z(n52132) );
  NANDN U52554 ( .A(n1580), .B(n52139), .Z(n52138) );
  NANDN U52555 ( .A(n1578), .B(n52140), .Z(n52139) );
  NAND U52556 ( .A(A[16]), .B(B[70]), .Z(n1580) );
  NAND U52557 ( .A(n32), .B(n1578), .Z(n52137) );
  XOR U52558 ( .A(n52141), .B(n52142), .Z(n1578) );
  XNOR U52559 ( .A(n52143), .B(n52144), .Z(n52142) );
  AND U52560 ( .A(n52145), .B(n52146), .Z(n52140) );
  NANDN U52561 ( .A(n1701), .B(n52147), .Z(n52146) );
  NANDN U52562 ( .A(n1699), .B(n52148), .Z(n52147) );
  NAND U52563 ( .A(A[15]), .B(B[70]), .Z(n1701) );
  NAND U52564 ( .A(n34), .B(n1699), .Z(n52145) );
  XOR U52565 ( .A(n52149), .B(n52150), .Z(n1699) );
  XNOR U52566 ( .A(n52151), .B(n52152), .Z(n52150) );
  AND U52567 ( .A(n52153), .B(n52154), .Z(n52148) );
  NANDN U52568 ( .A(n1829), .B(n52155), .Z(n52154) );
  NANDN U52569 ( .A(n1827), .B(n52156), .Z(n52155) );
  NAND U52570 ( .A(A[14]), .B(B[70]), .Z(n1829) );
  NAND U52571 ( .A(n35), .B(n1827), .Z(n52153) );
  XOR U52572 ( .A(n52157), .B(n52158), .Z(n1827) );
  XNOR U52573 ( .A(n52159), .B(n52160), .Z(n52158) );
  AND U52574 ( .A(n52161), .B(n52162), .Z(n52156) );
  NANDN U52575 ( .A(n1964), .B(n52163), .Z(n52162) );
  NANDN U52576 ( .A(n1962), .B(n52164), .Z(n52163) );
  NAND U52577 ( .A(A[13]), .B(B[70]), .Z(n1964) );
  NAND U52578 ( .A(n36), .B(n1962), .Z(n52161) );
  XOR U52579 ( .A(n52165), .B(n52166), .Z(n1962) );
  XNOR U52580 ( .A(n52167), .B(n52168), .Z(n52166) );
  AND U52581 ( .A(n52169), .B(n52170), .Z(n52164) );
  NANDN U52582 ( .A(n2106), .B(n52171), .Z(n52170) );
  NANDN U52583 ( .A(n2104), .B(n52172), .Z(n52171) );
  NAND U52584 ( .A(A[12]), .B(B[70]), .Z(n2106) );
  NAND U52585 ( .A(n37), .B(n2104), .Z(n52169) );
  XOR U52586 ( .A(n52173), .B(n52174), .Z(n2104) );
  XNOR U52587 ( .A(n52175), .B(n52176), .Z(n52174) );
  AND U52588 ( .A(n52177), .B(n52178), .Z(n52172) );
  NANDN U52589 ( .A(n2258), .B(n52179), .Z(n52178) );
  NANDN U52590 ( .A(n2256), .B(n52180), .Z(n52179) );
  NAND U52591 ( .A(A[11]), .B(B[70]), .Z(n2258) );
  NAND U52592 ( .A(n38), .B(n2256), .Z(n52177) );
  XOR U52593 ( .A(n52181), .B(n52182), .Z(n2256) );
  XNOR U52594 ( .A(n52183), .B(n52184), .Z(n52182) );
  AND U52595 ( .A(n52185), .B(n52186), .Z(n52180) );
  NANDN U52596 ( .A(n2414), .B(n52187), .Z(n52186) );
  NANDN U52597 ( .A(n2412), .B(n52188), .Z(n52187) );
  NAND U52598 ( .A(A[10]), .B(B[70]), .Z(n2414) );
  NAND U52599 ( .A(n39), .B(n2412), .Z(n52185) );
  XOR U52600 ( .A(n52189), .B(n52190), .Z(n2412) );
  XNOR U52601 ( .A(n52191), .B(n52192), .Z(n52190) );
  AND U52602 ( .A(n52193), .B(n52194), .Z(n52188) );
  NANDN U52603 ( .A(n2577), .B(n52195), .Z(n52194) );
  NANDN U52604 ( .A(n2575), .B(n52196), .Z(n52195) );
  NAND U52605 ( .A(A[9]), .B(B[70]), .Z(n2577) );
  NAND U52606 ( .A(n40), .B(n2575), .Z(n52193) );
  XOR U52607 ( .A(n52197), .B(n52198), .Z(n2575) );
  XNOR U52608 ( .A(n52199), .B(n52200), .Z(n52198) );
  AND U52609 ( .A(n52201), .B(n52202), .Z(n52196) );
  NANDN U52610 ( .A(n2747), .B(n52203), .Z(n52202) );
  NANDN U52611 ( .A(n2745), .B(n52204), .Z(n52203) );
  NAND U52612 ( .A(A[8]), .B(B[70]), .Z(n2747) );
  NAND U52613 ( .A(n41), .B(n2745), .Z(n52201) );
  XOR U52614 ( .A(n52205), .B(n52206), .Z(n2745) );
  XNOR U52615 ( .A(n52207), .B(n52208), .Z(n52206) );
  AND U52616 ( .A(n52209), .B(n52210), .Z(n52204) );
  NANDN U52617 ( .A(n2924), .B(n52211), .Z(n52210) );
  NANDN U52618 ( .A(n2922), .B(n52212), .Z(n52211) );
  NAND U52619 ( .A(A[7]), .B(B[70]), .Z(n2924) );
  NAND U52620 ( .A(n42), .B(n2922), .Z(n52209) );
  XOR U52621 ( .A(n52213), .B(n52214), .Z(n2922) );
  XNOR U52622 ( .A(n52215), .B(n52216), .Z(n52214) );
  AND U52623 ( .A(n52217), .B(n52218), .Z(n52212) );
  NANDN U52624 ( .A(n3108), .B(n52219), .Z(n52218) );
  NANDN U52625 ( .A(n3106), .B(n52220), .Z(n52219) );
  NAND U52626 ( .A(A[6]), .B(B[70]), .Z(n3108) );
  NAND U52627 ( .A(n43), .B(n3106), .Z(n52217) );
  XOR U52628 ( .A(n52221), .B(n52222), .Z(n3106) );
  XNOR U52629 ( .A(n52223), .B(n52224), .Z(n52222) );
  AND U52630 ( .A(n52225), .B(n52226), .Z(n52220) );
  NANDN U52631 ( .A(n3299), .B(n52227), .Z(n52226) );
  NANDN U52632 ( .A(n3297), .B(n52228), .Z(n52227) );
  NAND U52633 ( .A(A[5]), .B(B[70]), .Z(n3299) );
  NAND U52634 ( .A(n44), .B(n3297), .Z(n52225) );
  XOR U52635 ( .A(n52229), .B(n52230), .Z(n3297) );
  XNOR U52636 ( .A(n52231), .B(n52232), .Z(n52230) );
  AND U52637 ( .A(n52233), .B(n52234), .Z(n52228) );
  NANDN U52638 ( .A(n3497), .B(n52235), .Z(n52234) );
  NANDN U52639 ( .A(n3495), .B(n52236), .Z(n52235) );
  NAND U52640 ( .A(A[4]), .B(B[70]), .Z(n3497) );
  NAND U52641 ( .A(n45), .B(n3495), .Z(n52233) );
  XOR U52642 ( .A(n52237), .B(n52238), .Z(n3495) );
  XNOR U52643 ( .A(n52239), .B(n52240), .Z(n52238) );
  AND U52644 ( .A(n52241), .B(n52242), .Z(n52236) );
  NANDN U52645 ( .A(n3702), .B(n52243), .Z(n52242) );
  NAND U52646 ( .A(n52244), .B(n3700), .Z(n52243) );
  NAND U52647 ( .A(A[3]), .B(B[70]), .Z(n3702) );
  NANDN U52648 ( .A(n3700), .B(n47), .Z(n52241) );
  AND U52649 ( .A(n52245), .B(n52246), .Z(n52244) );
  NANDN U52650 ( .A(n3914), .B(n52247), .Z(n52246) );
  NANDN U52651 ( .A(n3915), .B(n3912), .Z(n52247) );
  NAND U52652 ( .A(B[70]), .B(A[2]), .Z(n3914) );
  ANDN U52653 ( .B(n52248), .A(n4132), .Z(n3915) );
  NAND U52654 ( .A(B[70]), .B(A[1]), .Z(n4132) );
  AND U52655 ( .A(A[0]), .B(B[71]), .Z(n52248) );
  XNOR U52656 ( .A(n52249), .B(n52250), .Z(n3912) );
  NAND U52657 ( .A(B[72]), .B(A[0]), .Z(n52250) );
  XOR U52658 ( .A(n46), .B(n52251), .Z(n3700) );
  XNOR U52659 ( .A(n52252), .B(n52253), .Z(n52251) );
  XNOR U52660 ( .A(n51836), .B(n52254), .Z(n614) );
  XNOR U52661 ( .A(n51835), .B(n51833), .Z(n52254) );
  AND U52662 ( .A(n52255), .B(n52256), .Z(n51833) );
  NANDN U52663 ( .A(n52040), .B(n52257), .Z(n52256) );
  AND U52664 ( .A(n52258), .B(n52259), .Z(n52040) );
  NANDN U52665 ( .A(n52048), .B(n52260), .Z(n52259) );
  OR U52666 ( .A(n52047), .B(n52045), .Z(n52260) );
  AND U52667 ( .A(n52261), .B(n52262), .Z(n52048) );
  NANDN U52668 ( .A(n52056), .B(n52263), .Z(n52262) );
  AND U52669 ( .A(n52264), .B(n52265), .Z(n52056) );
  NANDN U52670 ( .A(n52064), .B(n52266), .Z(n52265) );
  OR U52671 ( .A(n52063), .B(n52061), .Z(n52266) );
  AND U52672 ( .A(n52267), .B(n52268), .Z(n52064) );
  NANDN U52673 ( .A(n52072), .B(n52269), .Z(n52268) );
  AND U52674 ( .A(n52270), .B(n52271), .Z(n52072) );
  NANDN U52675 ( .A(n52080), .B(n52272), .Z(n52271) );
  OR U52676 ( .A(n52079), .B(n52077), .Z(n52272) );
  AND U52677 ( .A(n52273), .B(n52274), .Z(n52080) );
  NANDN U52678 ( .A(n52088), .B(n52275), .Z(n52274) );
  AND U52679 ( .A(n52276), .B(n52277), .Z(n52088) );
  NANDN U52680 ( .A(n52096), .B(n52278), .Z(n52277) );
  OR U52681 ( .A(n52095), .B(n52093), .Z(n52278) );
  AND U52682 ( .A(n52279), .B(n52280), .Z(n52096) );
  NANDN U52683 ( .A(n52104), .B(n52281), .Z(n52280) );
  AND U52684 ( .A(n52282), .B(n52283), .Z(n52104) );
  NANDN U52685 ( .A(n52112), .B(n52284), .Z(n52283) );
  OR U52686 ( .A(n52111), .B(n52109), .Z(n52284) );
  AND U52687 ( .A(n52285), .B(n52286), .Z(n52112) );
  NANDN U52688 ( .A(n52120), .B(n52287), .Z(n52286) );
  AND U52689 ( .A(n52288), .B(n52289), .Z(n52120) );
  NANDN U52690 ( .A(n52128), .B(n52290), .Z(n52289) );
  OR U52691 ( .A(n52127), .B(n52125), .Z(n52290) );
  AND U52692 ( .A(n52291), .B(n52292), .Z(n52128) );
  NANDN U52693 ( .A(n52136), .B(n52293), .Z(n52292) );
  AND U52694 ( .A(n52294), .B(n52295), .Z(n52136) );
  NANDN U52695 ( .A(n52144), .B(n52296), .Z(n52295) );
  OR U52696 ( .A(n52143), .B(n52141), .Z(n52296) );
  AND U52697 ( .A(n52297), .B(n52298), .Z(n52144) );
  NANDN U52698 ( .A(n52152), .B(n52299), .Z(n52298) );
  AND U52699 ( .A(n52300), .B(n52301), .Z(n52152) );
  NANDN U52700 ( .A(n52160), .B(n52302), .Z(n52301) );
  OR U52701 ( .A(n52159), .B(n52157), .Z(n52302) );
  AND U52702 ( .A(n52303), .B(n52304), .Z(n52160) );
  NANDN U52703 ( .A(n52168), .B(n52305), .Z(n52304) );
  AND U52704 ( .A(n52306), .B(n52307), .Z(n52168) );
  NANDN U52705 ( .A(n52176), .B(n52308), .Z(n52307) );
  OR U52706 ( .A(n52175), .B(n52173), .Z(n52308) );
  AND U52707 ( .A(n52309), .B(n52310), .Z(n52176) );
  NANDN U52708 ( .A(n52184), .B(n52311), .Z(n52310) );
  AND U52709 ( .A(n52312), .B(n52313), .Z(n52184) );
  NANDN U52710 ( .A(n52192), .B(n52314), .Z(n52313) );
  OR U52711 ( .A(n52191), .B(n52189), .Z(n52314) );
  AND U52712 ( .A(n52315), .B(n52316), .Z(n52192) );
  NANDN U52713 ( .A(n52200), .B(n52317), .Z(n52316) );
  AND U52714 ( .A(n52318), .B(n52319), .Z(n52200) );
  NANDN U52715 ( .A(n52208), .B(n52320), .Z(n52319) );
  OR U52716 ( .A(n52207), .B(n52205), .Z(n52320) );
  AND U52717 ( .A(n52321), .B(n52322), .Z(n52208) );
  NANDN U52718 ( .A(n52216), .B(n52323), .Z(n52322) );
  AND U52719 ( .A(n52324), .B(n52325), .Z(n52216) );
  NANDN U52720 ( .A(n52224), .B(n52326), .Z(n52325) );
  OR U52721 ( .A(n52223), .B(n52221), .Z(n52326) );
  AND U52722 ( .A(n52327), .B(n52328), .Z(n52224) );
  NANDN U52723 ( .A(n52232), .B(n52329), .Z(n52328) );
  AND U52724 ( .A(n52330), .B(n52331), .Z(n52232) );
  NANDN U52725 ( .A(n52240), .B(n52332), .Z(n52331) );
  OR U52726 ( .A(n52239), .B(n52237), .Z(n52332) );
  AND U52727 ( .A(n52333), .B(n52334), .Z(n52240) );
  NANDN U52728 ( .A(n52252), .B(n52335), .Z(n52334) );
  NAND U52729 ( .A(n52336), .B(n52253), .Z(n52335) );
  NANDN U52730 ( .A(n52249), .B(n52337), .Z(n52252) );
  AND U52731 ( .A(A[0]), .B(B[72]), .Z(n52337) );
  NAND U52732 ( .A(B[71]), .B(A[1]), .Z(n52249) );
  NANDN U52733 ( .A(n52253), .B(n46), .Z(n52333) );
  XNOR U52734 ( .A(n52338), .B(n52339), .Z(n52336) );
  NAND U52735 ( .A(B[73]), .B(A[0]), .Z(n52339) );
  NAND U52736 ( .A(B[71]), .B(A[2]), .Z(n52253) );
  NAND U52737 ( .A(n52237), .B(n52239), .Z(n52330) );
  ANDN U52738 ( .B(B[71]), .A(n82), .Z(n52239) );
  XOR U52739 ( .A(n52340), .B(n52341), .Z(n52237) );
  XNOR U52740 ( .A(n52342), .B(n52343), .Z(n52341) );
  NAND U52741 ( .A(n52229), .B(n52231), .Z(n52327) );
  ANDN U52742 ( .B(B[71]), .A(n81), .Z(n52231) );
  XOR U52743 ( .A(n52344), .B(n52345), .Z(n52229) );
  XNOR U52744 ( .A(n52346), .B(n52347), .Z(n52345) );
  NAND U52745 ( .A(n52221), .B(n52223), .Z(n52324) );
  ANDN U52746 ( .B(B[71]), .A(n80), .Z(n52223) );
  XNOR U52747 ( .A(n52348), .B(n52349), .Z(n52221) );
  XNOR U52748 ( .A(n52350), .B(n52351), .Z(n52349) );
  NAND U52749 ( .A(n52213), .B(n52215), .Z(n52321) );
  ANDN U52750 ( .B(B[71]), .A(n79), .Z(n52215) );
  XOR U52751 ( .A(n52352), .B(n52353), .Z(n52213) );
  XNOR U52752 ( .A(n52354), .B(n52355), .Z(n52353) );
  NAND U52753 ( .A(n52205), .B(n52207), .Z(n52318) );
  ANDN U52754 ( .B(B[71]), .A(n78), .Z(n52207) );
  XNOR U52755 ( .A(n52356), .B(n52357), .Z(n52205) );
  XNOR U52756 ( .A(n52358), .B(n52359), .Z(n52357) );
  NAND U52757 ( .A(n52197), .B(n52199), .Z(n52315) );
  ANDN U52758 ( .B(B[71]), .A(n77), .Z(n52199) );
  XOR U52759 ( .A(n52360), .B(n52361), .Z(n52197) );
  XNOR U52760 ( .A(n52362), .B(n52363), .Z(n52361) );
  NAND U52761 ( .A(n52189), .B(n52191), .Z(n52312) );
  ANDN U52762 ( .B(B[71]), .A(n76), .Z(n52191) );
  XNOR U52763 ( .A(n52364), .B(n52365), .Z(n52189) );
  XNOR U52764 ( .A(n52366), .B(n52367), .Z(n52365) );
  NAND U52765 ( .A(n52181), .B(n52183), .Z(n52309) );
  ANDN U52766 ( .B(B[71]), .A(n75), .Z(n52183) );
  XOR U52767 ( .A(n52368), .B(n52369), .Z(n52181) );
  XNOR U52768 ( .A(n52370), .B(n52371), .Z(n52369) );
  NAND U52769 ( .A(n52173), .B(n52175), .Z(n52306) );
  ANDN U52770 ( .B(B[71]), .A(n74), .Z(n52175) );
  XNOR U52771 ( .A(n52372), .B(n52373), .Z(n52173) );
  XNOR U52772 ( .A(n52374), .B(n52375), .Z(n52373) );
  NAND U52773 ( .A(n52165), .B(n52167), .Z(n52303) );
  ANDN U52774 ( .B(B[71]), .A(n73), .Z(n52167) );
  XOR U52775 ( .A(n52376), .B(n52377), .Z(n52165) );
  XNOR U52776 ( .A(n52378), .B(n52379), .Z(n52377) );
  NAND U52777 ( .A(n52157), .B(n52159), .Z(n52300) );
  ANDN U52778 ( .B(B[71]), .A(n72), .Z(n52159) );
  XNOR U52779 ( .A(n52380), .B(n52381), .Z(n52157) );
  XNOR U52780 ( .A(n52382), .B(n52383), .Z(n52381) );
  NAND U52781 ( .A(n52149), .B(n52151), .Z(n52297) );
  ANDN U52782 ( .B(B[71]), .A(n71), .Z(n52151) );
  XOR U52783 ( .A(n52384), .B(n52385), .Z(n52149) );
  XNOR U52784 ( .A(n52386), .B(n52387), .Z(n52385) );
  NAND U52785 ( .A(n52141), .B(n52143), .Z(n52294) );
  ANDN U52786 ( .B(B[71]), .A(n70), .Z(n52143) );
  XNOR U52787 ( .A(n52388), .B(n52389), .Z(n52141) );
  XNOR U52788 ( .A(n52390), .B(n52391), .Z(n52389) );
  NAND U52789 ( .A(n52133), .B(n52135), .Z(n52291) );
  ANDN U52790 ( .B(B[71]), .A(n69), .Z(n52135) );
  XOR U52791 ( .A(n52392), .B(n52393), .Z(n52133) );
  XNOR U52792 ( .A(n52394), .B(n52395), .Z(n52393) );
  NAND U52793 ( .A(n52125), .B(n52127), .Z(n52288) );
  ANDN U52794 ( .B(B[71]), .A(n68), .Z(n52127) );
  XNOR U52795 ( .A(n52396), .B(n52397), .Z(n52125) );
  XNOR U52796 ( .A(n52398), .B(n52399), .Z(n52397) );
  NAND U52797 ( .A(n52117), .B(n52119), .Z(n52285) );
  ANDN U52798 ( .B(B[71]), .A(n67), .Z(n52119) );
  XOR U52799 ( .A(n52400), .B(n52401), .Z(n52117) );
  XNOR U52800 ( .A(n52402), .B(n52403), .Z(n52401) );
  NAND U52801 ( .A(n52109), .B(n52111), .Z(n52282) );
  ANDN U52802 ( .B(B[71]), .A(n66), .Z(n52111) );
  XNOR U52803 ( .A(n52404), .B(n52405), .Z(n52109) );
  XNOR U52804 ( .A(n52406), .B(n52407), .Z(n52405) );
  NAND U52805 ( .A(n52101), .B(n52103), .Z(n52279) );
  ANDN U52806 ( .B(B[71]), .A(n65), .Z(n52103) );
  XOR U52807 ( .A(n52408), .B(n52409), .Z(n52101) );
  XNOR U52808 ( .A(n52410), .B(n52411), .Z(n52409) );
  NAND U52809 ( .A(n52093), .B(n52095), .Z(n52276) );
  ANDN U52810 ( .B(B[71]), .A(n64), .Z(n52095) );
  XNOR U52811 ( .A(n52412), .B(n52413), .Z(n52093) );
  XNOR U52812 ( .A(n52414), .B(n52415), .Z(n52413) );
  NAND U52813 ( .A(n52085), .B(n52087), .Z(n52273) );
  ANDN U52814 ( .B(B[71]), .A(n63), .Z(n52087) );
  XOR U52815 ( .A(n52416), .B(n52417), .Z(n52085) );
  XNOR U52816 ( .A(n52418), .B(n52419), .Z(n52417) );
  NAND U52817 ( .A(n52077), .B(n52079), .Z(n52270) );
  ANDN U52818 ( .B(B[71]), .A(n62), .Z(n52079) );
  XNOR U52819 ( .A(n52420), .B(n52421), .Z(n52077) );
  XNOR U52820 ( .A(n52422), .B(n52423), .Z(n52421) );
  NAND U52821 ( .A(n52069), .B(n52071), .Z(n52267) );
  ANDN U52822 ( .B(B[71]), .A(n61), .Z(n52071) );
  XOR U52823 ( .A(n52424), .B(n52425), .Z(n52069) );
  XNOR U52824 ( .A(n52426), .B(n52427), .Z(n52425) );
  NAND U52825 ( .A(n52061), .B(n52063), .Z(n52264) );
  ANDN U52826 ( .B(B[71]), .A(n60), .Z(n52063) );
  XNOR U52827 ( .A(n52428), .B(n52429), .Z(n52061) );
  XNOR U52828 ( .A(n52430), .B(n52431), .Z(n52429) );
  NAND U52829 ( .A(n52053), .B(n52055), .Z(n52261) );
  ANDN U52830 ( .B(B[71]), .A(n59), .Z(n52055) );
  XOR U52831 ( .A(n52432), .B(n52433), .Z(n52053) );
  XNOR U52832 ( .A(n52434), .B(n52435), .Z(n52433) );
  NAND U52833 ( .A(n52045), .B(n52047), .Z(n52258) );
  ANDN U52834 ( .B(B[71]), .A(n58), .Z(n52047) );
  XNOR U52835 ( .A(n52436), .B(n52437), .Z(n52045) );
  XNOR U52836 ( .A(n52438), .B(n52439), .Z(n52437) );
  NAND U52837 ( .A(n52037), .B(n52039), .Z(n52255) );
  ANDN U52838 ( .B(B[71]), .A(n57), .Z(n52039) );
  XOR U52839 ( .A(n52440), .B(n52441), .Z(n52037) );
  XNOR U52840 ( .A(n52442), .B(n52443), .Z(n52441) );
  ANDN U52841 ( .B(B[71]), .A(n56), .Z(n51835) );
  XNOR U52842 ( .A(n51843), .B(n52444), .Z(n51836) );
  XNOR U52843 ( .A(n51842), .B(n51840), .Z(n52444) );
  AND U52844 ( .A(n52445), .B(n52446), .Z(n51840) );
  NANDN U52845 ( .A(n52443), .B(n52447), .Z(n52446) );
  OR U52846 ( .A(n52442), .B(n52440), .Z(n52447) );
  AND U52847 ( .A(n52448), .B(n52449), .Z(n52443) );
  NANDN U52848 ( .A(n52439), .B(n52450), .Z(n52449) );
  NANDN U52849 ( .A(n52438), .B(n52436), .Z(n52450) );
  AND U52850 ( .A(n52451), .B(n52452), .Z(n52439) );
  NANDN U52851 ( .A(n52435), .B(n52453), .Z(n52452) );
  OR U52852 ( .A(n52434), .B(n52432), .Z(n52453) );
  AND U52853 ( .A(n52454), .B(n52455), .Z(n52435) );
  NANDN U52854 ( .A(n52431), .B(n52456), .Z(n52455) );
  NANDN U52855 ( .A(n52430), .B(n52428), .Z(n52456) );
  AND U52856 ( .A(n52457), .B(n52458), .Z(n52431) );
  NANDN U52857 ( .A(n52427), .B(n52459), .Z(n52458) );
  OR U52858 ( .A(n52426), .B(n52424), .Z(n52459) );
  AND U52859 ( .A(n52460), .B(n52461), .Z(n52427) );
  NANDN U52860 ( .A(n52423), .B(n52462), .Z(n52461) );
  NANDN U52861 ( .A(n52422), .B(n52420), .Z(n52462) );
  AND U52862 ( .A(n52463), .B(n52464), .Z(n52423) );
  NANDN U52863 ( .A(n52419), .B(n52465), .Z(n52464) );
  OR U52864 ( .A(n52418), .B(n52416), .Z(n52465) );
  AND U52865 ( .A(n52466), .B(n52467), .Z(n52419) );
  NANDN U52866 ( .A(n52415), .B(n52468), .Z(n52467) );
  NANDN U52867 ( .A(n52414), .B(n52412), .Z(n52468) );
  AND U52868 ( .A(n52469), .B(n52470), .Z(n52415) );
  NANDN U52869 ( .A(n52411), .B(n52471), .Z(n52470) );
  OR U52870 ( .A(n52410), .B(n52408), .Z(n52471) );
  AND U52871 ( .A(n52472), .B(n52473), .Z(n52411) );
  NANDN U52872 ( .A(n52407), .B(n52474), .Z(n52473) );
  NANDN U52873 ( .A(n52406), .B(n52404), .Z(n52474) );
  AND U52874 ( .A(n52475), .B(n52476), .Z(n52407) );
  NANDN U52875 ( .A(n52403), .B(n52477), .Z(n52476) );
  OR U52876 ( .A(n52402), .B(n52400), .Z(n52477) );
  AND U52877 ( .A(n52478), .B(n52479), .Z(n52403) );
  NANDN U52878 ( .A(n52399), .B(n52480), .Z(n52479) );
  NANDN U52879 ( .A(n52398), .B(n52396), .Z(n52480) );
  AND U52880 ( .A(n52481), .B(n52482), .Z(n52399) );
  NANDN U52881 ( .A(n52395), .B(n52483), .Z(n52482) );
  OR U52882 ( .A(n52394), .B(n52392), .Z(n52483) );
  AND U52883 ( .A(n52484), .B(n52485), .Z(n52395) );
  NANDN U52884 ( .A(n52391), .B(n52486), .Z(n52485) );
  NANDN U52885 ( .A(n52390), .B(n52388), .Z(n52486) );
  AND U52886 ( .A(n52487), .B(n52488), .Z(n52391) );
  NANDN U52887 ( .A(n52387), .B(n52489), .Z(n52488) );
  OR U52888 ( .A(n52386), .B(n52384), .Z(n52489) );
  AND U52889 ( .A(n52490), .B(n52491), .Z(n52387) );
  NANDN U52890 ( .A(n52383), .B(n52492), .Z(n52491) );
  NANDN U52891 ( .A(n52382), .B(n52380), .Z(n52492) );
  AND U52892 ( .A(n52493), .B(n52494), .Z(n52383) );
  NANDN U52893 ( .A(n52379), .B(n52495), .Z(n52494) );
  OR U52894 ( .A(n52378), .B(n52376), .Z(n52495) );
  AND U52895 ( .A(n52496), .B(n52497), .Z(n52379) );
  NANDN U52896 ( .A(n52375), .B(n52498), .Z(n52497) );
  NANDN U52897 ( .A(n52374), .B(n52372), .Z(n52498) );
  AND U52898 ( .A(n52499), .B(n52500), .Z(n52375) );
  NANDN U52899 ( .A(n52371), .B(n52501), .Z(n52500) );
  OR U52900 ( .A(n52370), .B(n52368), .Z(n52501) );
  AND U52901 ( .A(n52502), .B(n52503), .Z(n52371) );
  NANDN U52902 ( .A(n52367), .B(n52504), .Z(n52503) );
  NANDN U52903 ( .A(n52366), .B(n52364), .Z(n52504) );
  AND U52904 ( .A(n52505), .B(n52506), .Z(n52367) );
  NANDN U52905 ( .A(n52363), .B(n52507), .Z(n52506) );
  OR U52906 ( .A(n52362), .B(n52360), .Z(n52507) );
  AND U52907 ( .A(n52508), .B(n52509), .Z(n52363) );
  NANDN U52908 ( .A(n52359), .B(n52510), .Z(n52509) );
  NANDN U52909 ( .A(n52358), .B(n52356), .Z(n52510) );
  AND U52910 ( .A(n52511), .B(n52512), .Z(n52359) );
  NANDN U52911 ( .A(n52355), .B(n52513), .Z(n52512) );
  OR U52912 ( .A(n52354), .B(n52352), .Z(n52513) );
  AND U52913 ( .A(n52514), .B(n52515), .Z(n52355) );
  NANDN U52914 ( .A(n52351), .B(n52516), .Z(n52515) );
  NANDN U52915 ( .A(n52350), .B(n52348), .Z(n52516) );
  AND U52916 ( .A(n52517), .B(n52518), .Z(n52351) );
  NANDN U52917 ( .A(n52347), .B(n52519), .Z(n52518) );
  OR U52918 ( .A(n52346), .B(n52344), .Z(n52519) );
  AND U52919 ( .A(n52520), .B(n52521), .Z(n52347) );
  NANDN U52920 ( .A(n52342), .B(n52522), .Z(n52521) );
  NAND U52921 ( .A(n52340), .B(n52343), .Z(n52522) );
  NANDN U52922 ( .A(n52338), .B(n52523), .Z(n52342) );
  AND U52923 ( .A(A[0]), .B(B[73]), .Z(n52523) );
  NAND U52924 ( .A(B[72]), .B(A[1]), .Z(n52338) );
  XNOR U52925 ( .A(n52524), .B(n52525), .Z(n52340) );
  NAND U52926 ( .A(B[74]), .B(A[0]), .Z(n52525) );
  NAND U52927 ( .A(B[72]), .B(A[2]), .Z(n52343) );
  NAND U52928 ( .A(n52344), .B(n52346), .Z(n52517) );
  ANDN U52929 ( .B(B[72]), .A(n82), .Z(n52346) );
  XOR U52930 ( .A(n52526), .B(n52527), .Z(n52344) );
  XNOR U52931 ( .A(n52528), .B(n52529), .Z(n52527) );
  NANDN U52932 ( .A(n52348), .B(n52350), .Z(n52514) );
  ANDN U52933 ( .B(B[72]), .A(n81), .Z(n52350) );
  XNOR U52934 ( .A(n52530), .B(n52531), .Z(n52348) );
  XNOR U52935 ( .A(n52532), .B(n52533), .Z(n52531) );
  NAND U52936 ( .A(n52352), .B(n52354), .Z(n52511) );
  ANDN U52937 ( .B(B[72]), .A(n80), .Z(n52354) );
  XNOR U52938 ( .A(n52534), .B(n52535), .Z(n52352) );
  XNOR U52939 ( .A(n52536), .B(n52537), .Z(n52535) );
  NANDN U52940 ( .A(n52356), .B(n52358), .Z(n52508) );
  ANDN U52941 ( .B(B[72]), .A(n79), .Z(n52358) );
  XNOR U52942 ( .A(n52538), .B(n52539), .Z(n52356) );
  XNOR U52943 ( .A(n52540), .B(n52541), .Z(n52539) );
  NAND U52944 ( .A(n52360), .B(n52362), .Z(n52505) );
  ANDN U52945 ( .B(B[72]), .A(n78), .Z(n52362) );
  XNOR U52946 ( .A(n52542), .B(n52543), .Z(n52360) );
  XNOR U52947 ( .A(n52544), .B(n52545), .Z(n52543) );
  NANDN U52948 ( .A(n52364), .B(n52366), .Z(n52502) );
  ANDN U52949 ( .B(B[72]), .A(n77), .Z(n52366) );
  XNOR U52950 ( .A(n52546), .B(n52547), .Z(n52364) );
  XNOR U52951 ( .A(n52548), .B(n52549), .Z(n52547) );
  NAND U52952 ( .A(n52368), .B(n52370), .Z(n52499) );
  ANDN U52953 ( .B(B[72]), .A(n76), .Z(n52370) );
  XNOR U52954 ( .A(n52550), .B(n52551), .Z(n52368) );
  XNOR U52955 ( .A(n52552), .B(n52553), .Z(n52551) );
  NANDN U52956 ( .A(n52372), .B(n52374), .Z(n52496) );
  ANDN U52957 ( .B(B[72]), .A(n75), .Z(n52374) );
  XNOR U52958 ( .A(n52554), .B(n52555), .Z(n52372) );
  XNOR U52959 ( .A(n52556), .B(n52557), .Z(n52555) );
  NAND U52960 ( .A(n52376), .B(n52378), .Z(n52493) );
  ANDN U52961 ( .B(B[72]), .A(n74), .Z(n52378) );
  XNOR U52962 ( .A(n52558), .B(n52559), .Z(n52376) );
  XNOR U52963 ( .A(n52560), .B(n52561), .Z(n52559) );
  NANDN U52964 ( .A(n52380), .B(n52382), .Z(n52490) );
  ANDN U52965 ( .B(B[72]), .A(n73), .Z(n52382) );
  XNOR U52966 ( .A(n52562), .B(n52563), .Z(n52380) );
  XNOR U52967 ( .A(n52564), .B(n52565), .Z(n52563) );
  NAND U52968 ( .A(n52384), .B(n52386), .Z(n52487) );
  ANDN U52969 ( .B(B[72]), .A(n72), .Z(n52386) );
  XNOR U52970 ( .A(n52566), .B(n52567), .Z(n52384) );
  XNOR U52971 ( .A(n52568), .B(n52569), .Z(n52567) );
  NANDN U52972 ( .A(n52388), .B(n52390), .Z(n52484) );
  ANDN U52973 ( .B(B[72]), .A(n71), .Z(n52390) );
  XNOR U52974 ( .A(n52570), .B(n52571), .Z(n52388) );
  XNOR U52975 ( .A(n52572), .B(n52573), .Z(n52571) );
  NAND U52976 ( .A(n52392), .B(n52394), .Z(n52481) );
  ANDN U52977 ( .B(B[72]), .A(n70), .Z(n52394) );
  XNOR U52978 ( .A(n52574), .B(n52575), .Z(n52392) );
  XNOR U52979 ( .A(n52576), .B(n52577), .Z(n52575) );
  NANDN U52980 ( .A(n52396), .B(n52398), .Z(n52478) );
  ANDN U52981 ( .B(B[72]), .A(n69), .Z(n52398) );
  XNOR U52982 ( .A(n52578), .B(n52579), .Z(n52396) );
  XNOR U52983 ( .A(n52580), .B(n52581), .Z(n52579) );
  NAND U52984 ( .A(n52400), .B(n52402), .Z(n52475) );
  ANDN U52985 ( .B(B[72]), .A(n68), .Z(n52402) );
  XNOR U52986 ( .A(n52582), .B(n52583), .Z(n52400) );
  XNOR U52987 ( .A(n52584), .B(n52585), .Z(n52583) );
  NANDN U52988 ( .A(n52404), .B(n52406), .Z(n52472) );
  ANDN U52989 ( .B(B[72]), .A(n67), .Z(n52406) );
  XNOR U52990 ( .A(n52586), .B(n52587), .Z(n52404) );
  XNOR U52991 ( .A(n52588), .B(n52589), .Z(n52587) );
  NAND U52992 ( .A(n52408), .B(n52410), .Z(n52469) );
  ANDN U52993 ( .B(B[72]), .A(n66), .Z(n52410) );
  XNOR U52994 ( .A(n52590), .B(n52591), .Z(n52408) );
  XNOR U52995 ( .A(n52592), .B(n52593), .Z(n52591) );
  NANDN U52996 ( .A(n52412), .B(n52414), .Z(n52466) );
  ANDN U52997 ( .B(B[72]), .A(n65), .Z(n52414) );
  XNOR U52998 ( .A(n52594), .B(n52595), .Z(n52412) );
  XNOR U52999 ( .A(n52596), .B(n52597), .Z(n52595) );
  NAND U53000 ( .A(n52416), .B(n52418), .Z(n52463) );
  ANDN U53001 ( .B(B[72]), .A(n64), .Z(n52418) );
  XNOR U53002 ( .A(n52598), .B(n52599), .Z(n52416) );
  XNOR U53003 ( .A(n52600), .B(n52601), .Z(n52599) );
  NANDN U53004 ( .A(n52420), .B(n52422), .Z(n52460) );
  ANDN U53005 ( .B(B[72]), .A(n63), .Z(n52422) );
  XNOR U53006 ( .A(n52602), .B(n52603), .Z(n52420) );
  XNOR U53007 ( .A(n52604), .B(n52605), .Z(n52603) );
  NAND U53008 ( .A(n52424), .B(n52426), .Z(n52457) );
  ANDN U53009 ( .B(B[72]), .A(n62), .Z(n52426) );
  XNOR U53010 ( .A(n52606), .B(n52607), .Z(n52424) );
  XNOR U53011 ( .A(n52608), .B(n52609), .Z(n52607) );
  NANDN U53012 ( .A(n52428), .B(n52430), .Z(n52454) );
  ANDN U53013 ( .B(B[72]), .A(n61), .Z(n52430) );
  XNOR U53014 ( .A(n52610), .B(n52611), .Z(n52428) );
  XNOR U53015 ( .A(n52612), .B(n52613), .Z(n52611) );
  NAND U53016 ( .A(n52432), .B(n52434), .Z(n52451) );
  ANDN U53017 ( .B(B[72]), .A(n60), .Z(n52434) );
  XNOR U53018 ( .A(n52614), .B(n52615), .Z(n52432) );
  XNOR U53019 ( .A(n52616), .B(n52617), .Z(n52615) );
  NANDN U53020 ( .A(n52436), .B(n52438), .Z(n52448) );
  ANDN U53021 ( .B(B[72]), .A(n59), .Z(n52438) );
  XNOR U53022 ( .A(n52618), .B(n52619), .Z(n52436) );
  XNOR U53023 ( .A(n52620), .B(n52621), .Z(n52619) );
  NAND U53024 ( .A(n52440), .B(n52442), .Z(n52445) );
  ANDN U53025 ( .B(B[72]), .A(n58), .Z(n52442) );
  XNOR U53026 ( .A(n52622), .B(n52623), .Z(n52440) );
  XNOR U53027 ( .A(n52624), .B(n52625), .Z(n52623) );
  ANDN U53028 ( .B(B[72]), .A(n57), .Z(n51842) );
  XNOR U53029 ( .A(n51850), .B(n52626), .Z(n51843) );
  XNOR U53030 ( .A(n51849), .B(n51847), .Z(n52626) );
  AND U53031 ( .A(n52627), .B(n52628), .Z(n51847) );
  NANDN U53032 ( .A(n52625), .B(n52629), .Z(n52628) );
  NANDN U53033 ( .A(n52624), .B(n52622), .Z(n52629) );
  AND U53034 ( .A(n52630), .B(n52631), .Z(n52625) );
  NANDN U53035 ( .A(n52621), .B(n52632), .Z(n52631) );
  OR U53036 ( .A(n52620), .B(n52618), .Z(n52632) );
  AND U53037 ( .A(n52633), .B(n52634), .Z(n52621) );
  NANDN U53038 ( .A(n52617), .B(n52635), .Z(n52634) );
  NANDN U53039 ( .A(n52616), .B(n52614), .Z(n52635) );
  AND U53040 ( .A(n52636), .B(n52637), .Z(n52617) );
  NANDN U53041 ( .A(n52613), .B(n52638), .Z(n52637) );
  OR U53042 ( .A(n52612), .B(n52610), .Z(n52638) );
  AND U53043 ( .A(n52639), .B(n52640), .Z(n52613) );
  NANDN U53044 ( .A(n52609), .B(n52641), .Z(n52640) );
  NANDN U53045 ( .A(n52608), .B(n52606), .Z(n52641) );
  AND U53046 ( .A(n52642), .B(n52643), .Z(n52609) );
  NANDN U53047 ( .A(n52605), .B(n52644), .Z(n52643) );
  OR U53048 ( .A(n52604), .B(n52602), .Z(n52644) );
  AND U53049 ( .A(n52645), .B(n52646), .Z(n52605) );
  NANDN U53050 ( .A(n52601), .B(n52647), .Z(n52646) );
  NANDN U53051 ( .A(n52600), .B(n52598), .Z(n52647) );
  AND U53052 ( .A(n52648), .B(n52649), .Z(n52601) );
  NANDN U53053 ( .A(n52597), .B(n52650), .Z(n52649) );
  OR U53054 ( .A(n52596), .B(n52594), .Z(n52650) );
  AND U53055 ( .A(n52651), .B(n52652), .Z(n52597) );
  NANDN U53056 ( .A(n52593), .B(n52653), .Z(n52652) );
  NANDN U53057 ( .A(n52592), .B(n52590), .Z(n52653) );
  AND U53058 ( .A(n52654), .B(n52655), .Z(n52593) );
  NANDN U53059 ( .A(n52589), .B(n52656), .Z(n52655) );
  OR U53060 ( .A(n52588), .B(n52586), .Z(n52656) );
  AND U53061 ( .A(n52657), .B(n52658), .Z(n52589) );
  NANDN U53062 ( .A(n52585), .B(n52659), .Z(n52658) );
  NANDN U53063 ( .A(n52584), .B(n52582), .Z(n52659) );
  AND U53064 ( .A(n52660), .B(n52661), .Z(n52585) );
  NANDN U53065 ( .A(n52581), .B(n52662), .Z(n52661) );
  OR U53066 ( .A(n52580), .B(n52578), .Z(n52662) );
  AND U53067 ( .A(n52663), .B(n52664), .Z(n52581) );
  NANDN U53068 ( .A(n52577), .B(n52665), .Z(n52664) );
  NANDN U53069 ( .A(n52576), .B(n52574), .Z(n52665) );
  AND U53070 ( .A(n52666), .B(n52667), .Z(n52577) );
  NANDN U53071 ( .A(n52573), .B(n52668), .Z(n52667) );
  OR U53072 ( .A(n52572), .B(n52570), .Z(n52668) );
  AND U53073 ( .A(n52669), .B(n52670), .Z(n52573) );
  NANDN U53074 ( .A(n52569), .B(n52671), .Z(n52670) );
  NANDN U53075 ( .A(n52568), .B(n52566), .Z(n52671) );
  AND U53076 ( .A(n52672), .B(n52673), .Z(n52569) );
  NANDN U53077 ( .A(n52565), .B(n52674), .Z(n52673) );
  OR U53078 ( .A(n52564), .B(n52562), .Z(n52674) );
  AND U53079 ( .A(n52675), .B(n52676), .Z(n52565) );
  NANDN U53080 ( .A(n52561), .B(n52677), .Z(n52676) );
  NANDN U53081 ( .A(n52560), .B(n52558), .Z(n52677) );
  AND U53082 ( .A(n52678), .B(n52679), .Z(n52561) );
  NANDN U53083 ( .A(n52557), .B(n52680), .Z(n52679) );
  OR U53084 ( .A(n52556), .B(n52554), .Z(n52680) );
  AND U53085 ( .A(n52681), .B(n52682), .Z(n52557) );
  NANDN U53086 ( .A(n52553), .B(n52683), .Z(n52682) );
  NANDN U53087 ( .A(n52552), .B(n52550), .Z(n52683) );
  AND U53088 ( .A(n52684), .B(n52685), .Z(n52553) );
  NANDN U53089 ( .A(n52549), .B(n52686), .Z(n52685) );
  OR U53090 ( .A(n52548), .B(n52546), .Z(n52686) );
  AND U53091 ( .A(n52687), .B(n52688), .Z(n52549) );
  NANDN U53092 ( .A(n52545), .B(n52689), .Z(n52688) );
  NANDN U53093 ( .A(n52544), .B(n52542), .Z(n52689) );
  AND U53094 ( .A(n52690), .B(n52691), .Z(n52545) );
  NANDN U53095 ( .A(n52541), .B(n52692), .Z(n52691) );
  OR U53096 ( .A(n52540), .B(n52538), .Z(n52692) );
  AND U53097 ( .A(n52693), .B(n52694), .Z(n52541) );
  NANDN U53098 ( .A(n52537), .B(n52695), .Z(n52694) );
  NANDN U53099 ( .A(n52536), .B(n52534), .Z(n52695) );
  AND U53100 ( .A(n52696), .B(n52697), .Z(n52537) );
  NANDN U53101 ( .A(n52533), .B(n52698), .Z(n52697) );
  OR U53102 ( .A(n52532), .B(n52530), .Z(n52698) );
  AND U53103 ( .A(n52699), .B(n52700), .Z(n52533) );
  NANDN U53104 ( .A(n52528), .B(n52701), .Z(n52700) );
  NAND U53105 ( .A(n52526), .B(n52529), .Z(n52701) );
  NANDN U53106 ( .A(n52524), .B(n52702), .Z(n52528) );
  AND U53107 ( .A(A[0]), .B(B[74]), .Z(n52702) );
  NAND U53108 ( .A(B[73]), .B(A[1]), .Z(n52524) );
  XNOR U53109 ( .A(n52703), .B(n52704), .Z(n52526) );
  NAND U53110 ( .A(B[75]), .B(A[0]), .Z(n52704) );
  NAND U53111 ( .A(B[73]), .B(A[2]), .Z(n52529) );
  NAND U53112 ( .A(n52530), .B(n52532), .Z(n52696) );
  ANDN U53113 ( .B(B[73]), .A(n82), .Z(n52532) );
  XOR U53114 ( .A(n52705), .B(n52706), .Z(n52530) );
  XNOR U53115 ( .A(n52707), .B(n52708), .Z(n52706) );
  NANDN U53116 ( .A(n52534), .B(n52536), .Z(n52693) );
  ANDN U53117 ( .B(B[73]), .A(n81), .Z(n52536) );
  XNOR U53118 ( .A(n52709), .B(n52710), .Z(n52534) );
  XNOR U53119 ( .A(n52711), .B(n52712), .Z(n52710) );
  NAND U53120 ( .A(n52538), .B(n52540), .Z(n52690) );
  ANDN U53121 ( .B(B[73]), .A(n80), .Z(n52540) );
  XNOR U53122 ( .A(n52713), .B(n52714), .Z(n52538) );
  XNOR U53123 ( .A(n52715), .B(n52716), .Z(n52714) );
  NANDN U53124 ( .A(n52542), .B(n52544), .Z(n52687) );
  ANDN U53125 ( .B(B[73]), .A(n79), .Z(n52544) );
  XNOR U53126 ( .A(n52717), .B(n52718), .Z(n52542) );
  XNOR U53127 ( .A(n52719), .B(n52720), .Z(n52718) );
  NAND U53128 ( .A(n52546), .B(n52548), .Z(n52684) );
  ANDN U53129 ( .B(B[73]), .A(n78), .Z(n52548) );
  XNOR U53130 ( .A(n52721), .B(n52722), .Z(n52546) );
  XNOR U53131 ( .A(n52723), .B(n52724), .Z(n52722) );
  NANDN U53132 ( .A(n52550), .B(n52552), .Z(n52681) );
  ANDN U53133 ( .B(B[73]), .A(n77), .Z(n52552) );
  XNOR U53134 ( .A(n52725), .B(n52726), .Z(n52550) );
  XNOR U53135 ( .A(n52727), .B(n52728), .Z(n52726) );
  NAND U53136 ( .A(n52554), .B(n52556), .Z(n52678) );
  ANDN U53137 ( .B(B[73]), .A(n76), .Z(n52556) );
  XNOR U53138 ( .A(n52729), .B(n52730), .Z(n52554) );
  XNOR U53139 ( .A(n52731), .B(n52732), .Z(n52730) );
  NANDN U53140 ( .A(n52558), .B(n52560), .Z(n52675) );
  ANDN U53141 ( .B(B[73]), .A(n75), .Z(n52560) );
  XNOR U53142 ( .A(n52733), .B(n52734), .Z(n52558) );
  XNOR U53143 ( .A(n52735), .B(n52736), .Z(n52734) );
  NAND U53144 ( .A(n52562), .B(n52564), .Z(n52672) );
  ANDN U53145 ( .B(B[73]), .A(n74), .Z(n52564) );
  XNOR U53146 ( .A(n52737), .B(n52738), .Z(n52562) );
  XNOR U53147 ( .A(n52739), .B(n52740), .Z(n52738) );
  NANDN U53148 ( .A(n52566), .B(n52568), .Z(n52669) );
  ANDN U53149 ( .B(B[73]), .A(n73), .Z(n52568) );
  XNOR U53150 ( .A(n52741), .B(n52742), .Z(n52566) );
  XNOR U53151 ( .A(n52743), .B(n52744), .Z(n52742) );
  NAND U53152 ( .A(n52570), .B(n52572), .Z(n52666) );
  ANDN U53153 ( .B(B[73]), .A(n72), .Z(n52572) );
  XNOR U53154 ( .A(n52745), .B(n52746), .Z(n52570) );
  XNOR U53155 ( .A(n52747), .B(n52748), .Z(n52746) );
  NANDN U53156 ( .A(n52574), .B(n52576), .Z(n52663) );
  ANDN U53157 ( .B(B[73]), .A(n71), .Z(n52576) );
  XNOR U53158 ( .A(n52749), .B(n52750), .Z(n52574) );
  XNOR U53159 ( .A(n52751), .B(n52752), .Z(n52750) );
  NAND U53160 ( .A(n52578), .B(n52580), .Z(n52660) );
  ANDN U53161 ( .B(B[73]), .A(n70), .Z(n52580) );
  XNOR U53162 ( .A(n52753), .B(n52754), .Z(n52578) );
  XNOR U53163 ( .A(n52755), .B(n52756), .Z(n52754) );
  NANDN U53164 ( .A(n52582), .B(n52584), .Z(n52657) );
  ANDN U53165 ( .B(B[73]), .A(n69), .Z(n52584) );
  XNOR U53166 ( .A(n52757), .B(n52758), .Z(n52582) );
  XNOR U53167 ( .A(n52759), .B(n52760), .Z(n52758) );
  NAND U53168 ( .A(n52586), .B(n52588), .Z(n52654) );
  ANDN U53169 ( .B(B[73]), .A(n68), .Z(n52588) );
  XNOR U53170 ( .A(n52761), .B(n52762), .Z(n52586) );
  XNOR U53171 ( .A(n52763), .B(n52764), .Z(n52762) );
  NANDN U53172 ( .A(n52590), .B(n52592), .Z(n52651) );
  ANDN U53173 ( .B(B[73]), .A(n67), .Z(n52592) );
  XNOR U53174 ( .A(n52765), .B(n52766), .Z(n52590) );
  XNOR U53175 ( .A(n52767), .B(n52768), .Z(n52766) );
  NAND U53176 ( .A(n52594), .B(n52596), .Z(n52648) );
  ANDN U53177 ( .B(B[73]), .A(n66), .Z(n52596) );
  XNOR U53178 ( .A(n52769), .B(n52770), .Z(n52594) );
  XNOR U53179 ( .A(n52771), .B(n52772), .Z(n52770) );
  NANDN U53180 ( .A(n52598), .B(n52600), .Z(n52645) );
  ANDN U53181 ( .B(B[73]), .A(n65), .Z(n52600) );
  XNOR U53182 ( .A(n52773), .B(n52774), .Z(n52598) );
  XNOR U53183 ( .A(n52775), .B(n52776), .Z(n52774) );
  NAND U53184 ( .A(n52602), .B(n52604), .Z(n52642) );
  ANDN U53185 ( .B(B[73]), .A(n64), .Z(n52604) );
  XNOR U53186 ( .A(n52777), .B(n52778), .Z(n52602) );
  XNOR U53187 ( .A(n52779), .B(n52780), .Z(n52778) );
  NANDN U53188 ( .A(n52606), .B(n52608), .Z(n52639) );
  ANDN U53189 ( .B(B[73]), .A(n63), .Z(n52608) );
  XNOR U53190 ( .A(n52781), .B(n52782), .Z(n52606) );
  XNOR U53191 ( .A(n52783), .B(n52784), .Z(n52782) );
  NAND U53192 ( .A(n52610), .B(n52612), .Z(n52636) );
  ANDN U53193 ( .B(B[73]), .A(n62), .Z(n52612) );
  XNOR U53194 ( .A(n52785), .B(n52786), .Z(n52610) );
  XNOR U53195 ( .A(n52787), .B(n52788), .Z(n52786) );
  NANDN U53196 ( .A(n52614), .B(n52616), .Z(n52633) );
  ANDN U53197 ( .B(B[73]), .A(n61), .Z(n52616) );
  XNOR U53198 ( .A(n52789), .B(n52790), .Z(n52614) );
  XNOR U53199 ( .A(n52791), .B(n52792), .Z(n52790) );
  NAND U53200 ( .A(n52618), .B(n52620), .Z(n52630) );
  ANDN U53201 ( .B(B[73]), .A(n60), .Z(n52620) );
  XNOR U53202 ( .A(n52793), .B(n52794), .Z(n52618) );
  XNOR U53203 ( .A(n52795), .B(n52796), .Z(n52794) );
  NANDN U53204 ( .A(n52622), .B(n52624), .Z(n52627) );
  ANDN U53205 ( .B(B[73]), .A(n59), .Z(n52624) );
  XNOR U53206 ( .A(n52797), .B(n52798), .Z(n52622) );
  XNOR U53207 ( .A(n52799), .B(n52800), .Z(n52798) );
  ANDN U53208 ( .B(B[73]), .A(n58), .Z(n51849) );
  XNOR U53209 ( .A(n51857), .B(n52801), .Z(n51850) );
  XNOR U53210 ( .A(n51856), .B(n51854), .Z(n52801) );
  AND U53211 ( .A(n52802), .B(n52803), .Z(n51854) );
  NANDN U53212 ( .A(n52800), .B(n52804), .Z(n52803) );
  OR U53213 ( .A(n52799), .B(n52797), .Z(n52804) );
  AND U53214 ( .A(n52805), .B(n52806), .Z(n52800) );
  NANDN U53215 ( .A(n52796), .B(n52807), .Z(n52806) );
  NANDN U53216 ( .A(n52795), .B(n52793), .Z(n52807) );
  AND U53217 ( .A(n52808), .B(n52809), .Z(n52796) );
  NANDN U53218 ( .A(n52792), .B(n52810), .Z(n52809) );
  OR U53219 ( .A(n52791), .B(n52789), .Z(n52810) );
  AND U53220 ( .A(n52811), .B(n52812), .Z(n52792) );
  NANDN U53221 ( .A(n52788), .B(n52813), .Z(n52812) );
  NANDN U53222 ( .A(n52787), .B(n52785), .Z(n52813) );
  AND U53223 ( .A(n52814), .B(n52815), .Z(n52788) );
  NANDN U53224 ( .A(n52784), .B(n52816), .Z(n52815) );
  OR U53225 ( .A(n52783), .B(n52781), .Z(n52816) );
  AND U53226 ( .A(n52817), .B(n52818), .Z(n52784) );
  NANDN U53227 ( .A(n52780), .B(n52819), .Z(n52818) );
  NANDN U53228 ( .A(n52779), .B(n52777), .Z(n52819) );
  AND U53229 ( .A(n52820), .B(n52821), .Z(n52780) );
  NANDN U53230 ( .A(n52776), .B(n52822), .Z(n52821) );
  OR U53231 ( .A(n52775), .B(n52773), .Z(n52822) );
  AND U53232 ( .A(n52823), .B(n52824), .Z(n52776) );
  NANDN U53233 ( .A(n52772), .B(n52825), .Z(n52824) );
  NANDN U53234 ( .A(n52771), .B(n52769), .Z(n52825) );
  AND U53235 ( .A(n52826), .B(n52827), .Z(n52772) );
  NANDN U53236 ( .A(n52768), .B(n52828), .Z(n52827) );
  OR U53237 ( .A(n52767), .B(n52765), .Z(n52828) );
  AND U53238 ( .A(n52829), .B(n52830), .Z(n52768) );
  NANDN U53239 ( .A(n52764), .B(n52831), .Z(n52830) );
  NANDN U53240 ( .A(n52763), .B(n52761), .Z(n52831) );
  AND U53241 ( .A(n52832), .B(n52833), .Z(n52764) );
  NANDN U53242 ( .A(n52760), .B(n52834), .Z(n52833) );
  OR U53243 ( .A(n52759), .B(n52757), .Z(n52834) );
  AND U53244 ( .A(n52835), .B(n52836), .Z(n52760) );
  NANDN U53245 ( .A(n52756), .B(n52837), .Z(n52836) );
  NANDN U53246 ( .A(n52755), .B(n52753), .Z(n52837) );
  AND U53247 ( .A(n52838), .B(n52839), .Z(n52756) );
  NANDN U53248 ( .A(n52752), .B(n52840), .Z(n52839) );
  OR U53249 ( .A(n52751), .B(n52749), .Z(n52840) );
  AND U53250 ( .A(n52841), .B(n52842), .Z(n52752) );
  NANDN U53251 ( .A(n52748), .B(n52843), .Z(n52842) );
  NANDN U53252 ( .A(n52747), .B(n52745), .Z(n52843) );
  AND U53253 ( .A(n52844), .B(n52845), .Z(n52748) );
  NANDN U53254 ( .A(n52744), .B(n52846), .Z(n52845) );
  OR U53255 ( .A(n52743), .B(n52741), .Z(n52846) );
  AND U53256 ( .A(n52847), .B(n52848), .Z(n52744) );
  NANDN U53257 ( .A(n52740), .B(n52849), .Z(n52848) );
  NANDN U53258 ( .A(n52739), .B(n52737), .Z(n52849) );
  AND U53259 ( .A(n52850), .B(n52851), .Z(n52740) );
  NANDN U53260 ( .A(n52736), .B(n52852), .Z(n52851) );
  OR U53261 ( .A(n52735), .B(n52733), .Z(n52852) );
  AND U53262 ( .A(n52853), .B(n52854), .Z(n52736) );
  NANDN U53263 ( .A(n52732), .B(n52855), .Z(n52854) );
  NANDN U53264 ( .A(n52731), .B(n52729), .Z(n52855) );
  AND U53265 ( .A(n52856), .B(n52857), .Z(n52732) );
  NANDN U53266 ( .A(n52728), .B(n52858), .Z(n52857) );
  OR U53267 ( .A(n52727), .B(n52725), .Z(n52858) );
  AND U53268 ( .A(n52859), .B(n52860), .Z(n52728) );
  NANDN U53269 ( .A(n52724), .B(n52861), .Z(n52860) );
  NANDN U53270 ( .A(n52723), .B(n52721), .Z(n52861) );
  AND U53271 ( .A(n52862), .B(n52863), .Z(n52724) );
  NANDN U53272 ( .A(n52720), .B(n52864), .Z(n52863) );
  OR U53273 ( .A(n52719), .B(n52717), .Z(n52864) );
  AND U53274 ( .A(n52865), .B(n52866), .Z(n52720) );
  NANDN U53275 ( .A(n52716), .B(n52867), .Z(n52866) );
  NANDN U53276 ( .A(n52715), .B(n52713), .Z(n52867) );
  AND U53277 ( .A(n52868), .B(n52869), .Z(n52716) );
  NANDN U53278 ( .A(n52712), .B(n52870), .Z(n52869) );
  OR U53279 ( .A(n52711), .B(n52709), .Z(n52870) );
  AND U53280 ( .A(n52871), .B(n52872), .Z(n52712) );
  NANDN U53281 ( .A(n52707), .B(n52873), .Z(n52872) );
  NAND U53282 ( .A(n52705), .B(n52708), .Z(n52873) );
  NANDN U53283 ( .A(n52703), .B(n52874), .Z(n52707) );
  AND U53284 ( .A(A[0]), .B(B[75]), .Z(n52874) );
  NAND U53285 ( .A(B[74]), .B(A[1]), .Z(n52703) );
  XNOR U53286 ( .A(n52875), .B(n52876), .Z(n52705) );
  NAND U53287 ( .A(B[76]), .B(A[0]), .Z(n52876) );
  NAND U53288 ( .A(B[74]), .B(A[2]), .Z(n52708) );
  NAND U53289 ( .A(n52709), .B(n52711), .Z(n52868) );
  ANDN U53290 ( .B(B[74]), .A(n82), .Z(n52711) );
  XOR U53291 ( .A(n52877), .B(n52878), .Z(n52709) );
  XNOR U53292 ( .A(n52879), .B(n52880), .Z(n52878) );
  NANDN U53293 ( .A(n52713), .B(n52715), .Z(n52865) );
  ANDN U53294 ( .B(B[74]), .A(n81), .Z(n52715) );
  XNOR U53295 ( .A(n52881), .B(n52882), .Z(n52713) );
  XNOR U53296 ( .A(n52883), .B(n52884), .Z(n52882) );
  NAND U53297 ( .A(n52717), .B(n52719), .Z(n52862) );
  ANDN U53298 ( .B(B[74]), .A(n80), .Z(n52719) );
  XNOR U53299 ( .A(n52885), .B(n52886), .Z(n52717) );
  XNOR U53300 ( .A(n52887), .B(n52888), .Z(n52886) );
  NANDN U53301 ( .A(n52721), .B(n52723), .Z(n52859) );
  ANDN U53302 ( .B(B[74]), .A(n79), .Z(n52723) );
  XNOR U53303 ( .A(n52889), .B(n52890), .Z(n52721) );
  XNOR U53304 ( .A(n52891), .B(n52892), .Z(n52890) );
  NAND U53305 ( .A(n52725), .B(n52727), .Z(n52856) );
  ANDN U53306 ( .B(B[74]), .A(n78), .Z(n52727) );
  XNOR U53307 ( .A(n52893), .B(n52894), .Z(n52725) );
  XNOR U53308 ( .A(n52895), .B(n52896), .Z(n52894) );
  NANDN U53309 ( .A(n52729), .B(n52731), .Z(n52853) );
  ANDN U53310 ( .B(B[74]), .A(n77), .Z(n52731) );
  XNOR U53311 ( .A(n52897), .B(n52898), .Z(n52729) );
  XNOR U53312 ( .A(n52899), .B(n52900), .Z(n52898) );
  NAND U53313 ( .A(n52733), .B(n52735), .Z(n52850) );
  ANDN U53314 ( .B(B[74]), .A(n76), .Z(n52735) );
  XNOR U53315 ( .A(n52901), .B(n52902), .Z(n52733) );
  XNOR U53316 ( .A(n52903), .B(n52904), .Z(n52902) );
  NANDN U53317 ( .A(n52737), .B(n52739), .Z(n52847) );
  ANDN U53318 ( .B(B[74]), .A(n75), .Z(n52739) );
  XNOR U53319 ( .A(n52905), .B(n52906), .Z(n52737) );
  XNOR U53320 ( .A(n52907), .B(n52908), .Z(n52906) );
  NAND U53321 ( .A(n52741), .B(n52743), .Z(n52844) );
  ANDN U53322 ( .B(B[74]), .A(n74), .Z(n52743) );
  XNOR U53323 ( .A(n52909), .B(n52910), .Z(n52741) );
  XNOR U53324 ( .A(n52911), .B(n52912), .Z(n52910) );
  NANDN U53325 ( .A(n52745), .B(n52747), .Z(n52841) );
  ANDN U53326 ( .B(B[74]), .A(n73), .Z(n52747) );
  XNOR U53327 ( .A(n52913), .B(n52914), .Z(n52745) );
  XNOR U53328 ( .A(n52915), .B(n52916), .Z(n52914) );
  NAND U53329 ( .A(n52749), .B(n52751), .Z(n52838) );
  ANDN U53330 ( .B(B[74]), .A(n72), .Z(n52751) );
  XNOR U53331 ( .A(n52917), .B(n52918), .Z(n52749) );
  XNOR U53332 ( .A(n52919), .B(n52920), .Z(n52918) );
  NANDN U53333 ( .A(n52753), .B(n52755), .Z(n52835) );
  ANDN U53334 ( .B(B[74]), .A(n71), .Z(n52755) );
  XNOR U53335 ( .A(n52921), .B(n52922), .Z(n52753) );
  XNOR U53336 ( .A(n52923), .B(n52924), .Z(n52922) );
  NAND U53337 ( .A(n52757), .B(n52759), .Z(n52832) );
  ANDN U53338 ( .B(B[74]), .A(n70), .Z(n52759) );
  XNOR U53339 ( .A(n52925), .B(n52926), .Z(n52757) );
  XNOR U53340 ( .A(n52927), .B(n52928), .Z(n52926) );
  NANDN U53341 ( .A(n52761), .B(n52763), .Z(n52829) );
  ANDN U53342 ( .B(B[74]), .A(n69), .Z(n52763) );
  XNOR U53343 ( .A(n52929), .B(n52930), .Z(n52761) );
  XNOR U53344 ( .A(n52931), .B(n52932), .Z(n52930) );
  NAND U53345 ( .A(n52765), .B(n52767), .Z(n52826) );
  ANDN U53346 ( .B(B[74]), .A(n68), .Z(n52767) );
  XNOR U53347 ( .A(n52933), .B(n52934), .Z(n52765) );
  XNOR U53348 ( .A(n52935), .B(n52936), .Z(n52934) );
  NANDN U53349 ( .A(n52769), .B(n52771), .Z(n52823) );
  ANDN U53350 ( .B(B[74]), .A(n67), .Z(n52771) );
  XNOR U53351 ( .A(n52937), .B(n52938), .Z(n52769) );
  XNOR U53352 ( .A(n52939), .B(n52940), .Z(n52938) );
  NAND U53353 ( .A(n52773), .B(n52775), .Z(n52820) );
  ANDN U53354 ( .B(B[74]), .A(n66), .Z(n52775) );
  XNOR U53355 ( .A(n52941), .B(n52942), .Z(n52773) );
  XNOR U53356 ( .A(n52943), .B(n52944), .Z(n52942) );
  NANDN U53357 ( .A(n52777), .B(n52779), .Z(n52817) );
  ANDN U53358 ( .B(B[74]), .A(n65), .Z(n52779) );
  XNOR U53359 ( .A(n52945), .B(n52946), .Z(n52777) );
  XNOR U53360 ( .A(n52947), .B(n52948), .Z(n52946) );
  NAND U53361 ( .A(n52781), .B(n52783), .Z(n52814) );
  ANDN U53362 ( .B(B[74]), .A(n64), .Z(n52783) );
  XNOR U53363 ( .A(n52949), .B(n52950), .Z(n52781) );
  XNOR U53364 ( .A(n52951), .B(n52952), .Z(n52950) );
  NANDN U53365 ( .A(n52785), .B(n52787), .Z(n52811) );
  ANDN U53366 ( .B(B[74]), .A(n63), .Z(n52787) );
  XNOR U53367 ( .A(n52953), .B(n52954), .Z(n52785) );
  XNOR U53368 ( .A(n52955), .B(n52956), .Z(n52954) );
  NAND U53369 ( .A(n52789), .B(n52791), .Z(n52808) );
  ANDN U53370 ( .B(B[74]), .A(n62), .Z(n52791) );
  XNOR U53371 ( .A(n52957), .B(n52958), .Z(n52789) );
  XNOR U53372 ( .A(n52959), .B(n52960), .Z(n52958) );
  NANDN U53373 ( .A(n52793), .B(n52795), .Z(n52805) );
  ANDN U53374 ( .B(B[74]), .A(n61), .Z(n52795) );
  XNOR U53375 ( .A(n52961), .B(n52962), .Z(n52793) );
  XNOR U53376 ( .A(n52963), .B(n52964), .Z(n52962) );
  NAND U53377 ( .A(n52797), .B(n52799), .Z(n52802) );
  ANDN U53378 ( .B(B[74]), .A(n60), .Z(n52799) );
  XNOR U53379 ( .A(n52965), .B(n52966), .Z(n52797) );
  XNOR U53380 ( .A(n52967), .B(n52968), .Z(n52966) );
  ANDN U53381 ( .B(B[74]), .A(n59), .Z(n51856) );
  XNOR U53382 ( .A(n51864), .B(n52969), .Z(n51857) );
  XNOR U53383 ( .A(n51863), .B(n51861), .Z(n52969) );
  AND U53384 ( .A(n52970), .B(n52971), .Z(n51861) );
  NANDN U53385 ( .A(n52968), .B(n52972), .Z(n52971) );
  NANDN U53386 ( .A(n52967), .B(n52965), .Z(n52972) );
  AND U53387 ( .A(n52973), .B(n52974), .Z(n52968) );
  NANDN U53388 ( .A(n52964), .B(n52975), .Z(n52974) );
  OR U53389 ( .A(n52963), .B(n52961), .Z(n52975) );
  AND U53390 ( .A(n52976), .B(n52977), .Z(n52964) );
  NANDN U53391 ( .A(n52960), .B(n52978), .Z(n52977) );
  NANDN U53392 ( .A(n52959), .B(n52957), .Z(n52978) );
  AND U53393 ( .A(n52979), .B(n52980), .Z(n52960) );
  NANDN U53394 ( .A(n52956), .B(n52981), .Z(n52980) );
  OR U53395 ( .A(n52955), .B(n52953), .Z(n52981) );
  AND U53396 ( .A(n52982), .B(n52983), .Z(n52956) );
  NANDN U53397 ( .A(n52952), .B(n52984), .Z(n52983) );
  NANDN U53398 ( .A(n52951), .B(n52949), .Z(n52984) );
  AND U53399 ( .A(n52985), .B(n52986), .Z(n52952) );
  NANDN U53400 ( .A(n52948), .B(n52987), .Z(n52986) );
  OR U53401 ( .A(n52947), .B(n52945), .Z(n52987) );
  AND U53402 ( .A(n52988), .B(n52989), .Z(n52948) );
  NANDN U53403 ( .A(n52944), .B(n52990), .Z(n52989) );
  NANDN U53404 ( .A(n52943), .B(n52941), .Z(n52990) );
  AND U53405 ( .A(n52991), .B(n52992), .Z(n52944) );
  NANDN U53406 ( .A(n52940), .B(n52993), .Z(n52992) );
  OR U53407 ( .A(n52939), .B(n52937), .Z(n52993) );
  AND U53408 ( .A(n52994), .B(n52995), .Z(n52940) );
  NANDN U53409 ( .A(n52936), .B(n52996), .Z(n52995) );
  NANDN U53410 ( .A(n52935), .B(n52933), .Z(n52996) );
  AND U53411 ( .A(n52997), .B(n52998), .Z(n52936) );
  NANDN U53412 ( .A(n52932), .B(n52999), .Z(n52998) );
  OR U53413 ( .A(n52931), .B(n52929), .Z(n52999) );
  AND U53414 ( .A(n53000), .B(n53001), .Z(n52932) );
  NANDN U53415 ( .A(n52928), .B(n53002), .Z(n53001) );
  NANDN U53416 ( .A(n52927), .B(n52925), .Z(n53002) );
  AND U53417 ( .A(n53003), .B(n53004), .Z(n52928) );
  NANDN U53418 ( .A(n52924), .B(n53005), .Z(n53004) );
  OR U53419 ( .A(n52923), .B(n52921), .Z(n53005) );
  AND U53420 ( .A(n53006), .B(n53007), .Z(n52924) );
  NANDN U53421 ( .A(n52920), .B(n53008), .Z(n53007) );
  NANDN U53422 ( .A(n52919), .B(n52917), .Z(n53008) );
  AND U53423 ( .A(n53009), .B(n53010), .Z(n52920) );
  NANDN U53424 ( .A(n52916), .B(n53011), .Z(n53010) );
  OR U53425 ( .A(n52915), .B(n52913), .Z(n53011) );
  AND U53426 ( .A(n53012), .B(n53013), .Z(n52916) );
  NANDN U53427 ( .A(n52912), .B(n53014), .Z(n53013) );
  NANDN U53428 ( .A(n52911), .B(n52909), .Z(n53014) );
  AND U53429 ( .A(n53015), .B(n53016), .Z(n52912) );
  NANDN U53430 ( .A(n52908), .B(n53017), .Z(n53016) );
  OR U53431 ( .A(n52907), .B(n52905), .Z(n53017) );
  AND U53432 ( .A(n53018), .B(n53019), .Z(n52908) );
  NANDN U53433 ( .A(n52904), .B(n53020), .Z(n53019) );
  NANDN U53434 ( .A(n52903), .B(n52901), .Z(n53020) );
  AND U53435 ( .A(n53021), .B(n53022), .Z(n52904) );
  NANDN U53436 ( .A(n52900), .B(n53023), .Z(n53022) );
  OR U53437 ( .A(n52899), .B(n52897), .Z(n53023) );
  AND U53438 ( .A(n53024), .B(n53025), .Z(n52900) );
  NANDN U53439 ( .A(n52896), .B(n53026), .Z(n53025) );
  NANDN U53440 ( .A(n52895), .B(n52893), .Z(n53026) );
  AND U53441 ( .A(n53027), .B(n53028), .Z(n52896) );
  NANDN U53442 ( .A(n52892), .B(n53029), .Z(n53028) );
  OR U53443 ( .A(n52891), .B(n52889), .Z(n53029) );
  AND U53444 ( .A(n53030), .B(n53031), .Z(n52892) );
  NANDN U53445 ( .A(n52888), .B(n53032), .Z(n53031) );
  NANDN U53446 ( .A(n52887), .B(n52885), .Z(n53032) );
  AND U53447 ( .A(n53033), .B(n53034), .Z(n52888) );
  NANDN U53448 ( .A(n52884), .B(n53035), .Z(n53034) );
  OR U53449 ( .A(n52883), .B(n52881), .Z(n53035) );
  AND U53450 ( .A(n53036), .B(n53037), .Z(n52884) );
  NANDN U53451 ( .A(n52879), .B(n53038), .Z(n53037) );
  NAND U53452 ( .A(n52877), .B(n52880), .Z(n53038) );
  NANDN U53453 ( .A(n52875), .B(n53039), .Z(n52879) );
  AND U53454 ( .A(A[0]), .B(B[76]), .Z(n53039) );
  NAND U53455 ( .A(B[75]), .B(A[1]), .Z(n52875) );
  XNOR U53456 ( .A(n53040), .B(n53041), .Z(n52877) );
  NAND U53457 ( .A(B[77]), .B(A[0]), .Z(n53041) );
  NAND U53458 ( .A(B[75]), .B(A[2]), .Z(n52880) );
  NAND U53459 ( .A(n52881), .B(n52883), .Z(n53033) );
  ANDN U53460 ( .B(B[75]), .A(n82), .Z(n52883) );
  XOR U53461 ( .A(n53042), .B(n53043), .Z(n52881) );
  XNOR U53462 ( .A(n53044), .B(n53045), .Z(n53043) );
  NANDN U53463 ( .A(n52885), .B(n52887), .Z(n53030) );
  ANDN U53464 ( .B(B[75]), .A(n81), .Z(n52887) );
  XNOR U53465 ( .A(n53046), .B(n53047), .Z(n52885) );
  XNOR U53466 ( .A(n53048), .B(n53049), .Z(n53047) );
  NAND U53467 ( .A(n52889), .B(n52891), .Z(n53027) );
  ANDN U53468 ( .B(B[75]), .A(n80), .Z(n52891) );
  XNOR U53469 ( .A(n53050), .B(n53051), .Z(n52889) );
  XNOR U53470 ( .A(n53052), .B(n53053), .Z(n53051) );
  NANDN U53471 ( .A(n52893), .B(n52895), .Z(n53024) );
  ANDN U53472 ( .B(B[75]), .A(n79), .Z(n52895) );
  XNOR U53473 ( .A(n53054), .B(n53055), .Z(n52893) );
  XNOR U53474 ( .A(n53056), .B(n53057), .Z(n53055) );
  NAND U53475 ( .A(n52897), .B(n52899), .Z(n53021) );
  ANDN U53476 ( .B(B[75]), .A(n78), .Z(n52899) );
  XNOR U53477 ( .A(n53058), .B(n53059), .Z(n52897) );
  XNOR U53478 ( .A(n53060), .B(n53061), .Z(n53059) );
  NANDN U53479 ( .A(n52901), .B(n52903), .Z(n53018) );
  ANDN U53480 ( .B(B[75]), .A(n77), .Z(n52903) );
  XNOR U53481 ( .A(n53062), .B(n53063), .Z(n52901) );
  XNOR U53482 ( .A(n53064), .B(n53065), .Z(n53063) );
  NAND U53483 ( .A(n52905), .B(n52907), .Z(n53015) );
  ANDN U53484 ( .B(B[75]), .A(n76), .Z(n52907) );
  XNOR U53485 ( .A(n53066), .B(n53067), .Z(n52905) );
  XNOR U53486 ( .A(n53068), .B(n53069), .Z(n53067) );
  NANDN U53487 ( .A(n52909), .B(n52911), .Z(n53012) );
  ANDN U53488 ( .B(B[75]), .A(n75), .Z(n52911) );
  XNOR U53489 ( .A(n53070), .B(n53071), .Z(n52909) );
  XNOR U53490 ( .A(n53072), .B(n53073), .Z(n53071) );
  NAND U53491 ( .A(n52913), .B(n52915), .Z(n53009) );
  ANDN U53492 ( .B(B[75]), .A(n74), .Z(n52915) );
  XNOR U53493 ( .A(n53074), .B(n53075), .Z(n52913) );
  XNOR U53494 ( .A(n53076), .B(n53077), .Z(n53075) );
  NANDN U53495 ( .A(n52917), .B(n52919), .Z(n53006) );
  ANDN U53496 ( .B(B[75]), .A(n73), .Z(n52919) );
  XNOR U53497 ( .A(n53078), .B(n53079), .Z(n52917) );
  XNOR U53498 ( .A(n53080), .B(n53081), .Z(n53079) );
  NAND U53499 ( .A(n52921), .B(n52923), .Z(n53003) );
  ANDN U53500 ( .B(B[75]), .A(n72), .Z(n52923) );
  XNOR U53501 ( .A(n53082), .B(n53083), .Z(n52921) );
  XNOR U53502 ( .A(n53084), .B(n53085), .Z(n53083) );
  NANDN U53503 ( .A(n52925), .B(n52927), .Z(n53000) );
  ANDN U53504 ( .B(B[75]), .A(n71), .Z(n52927) );
  XNOR U53505 ( .A(n53086), .B(n53087), .Z(n52925) );
  XNOR U53506 ( .A(n53088), .B(n53089), .Z(n53087) );
  NAND U53507 ( .A(n52929), .B(n52931), .Z(n52997) );
  ANDN U53508 ( .B(B[75]), .A(n70), .Z(n52931) );
  XNOR U53509 ( .A(n53090), .B(n53091), .Z(n52929) );
  XNOR U53510 ( .A(n53092), .B(n53093), .Z(n53091) );
  NANDN U53511 ( .A(n52933), .B(n52935), .Z(n52994) );
  ANDN U53512 ( .B(B[75]), .A(n69), .Z(n52935) );
  XNOR U53513 ( .A(n53094), .B(n53095), .Z(n52933) );
  XNOR U53514 ( .A(n53096), .B(n53097), .Z(n53095) );
  NAND U53515 ( .A(n52937), .B(n52939), .Z(n52991) );
  ANDN U53516 ( .B(B[75]), .A(n68), .Z(n52939) );
  XNOR U53517 ( .A(n53098), .B(n53099), .Z(n52937) );
  XNOR U53518 ( .A(n53100), .B(n53101), .Z(n53099) );
  NANDN U53519 ( .A(n52941), .B(n52943), .Z(n52988) );
  ANDN U53520 ( .B(B[75]), .A(n67), .Z(n52943) );
  XNOR U53521 ( .A(n53102), .B(n53103), .Z(n52941) );
  XNOR U53522 ( .A(n53104), .B(n53105), .Z(n53103) );
  NAND U53523 ( .A(n52945), .B(n52947), .Z(n52985) );
  ANDN U53524 ( .B(B[75]), .A(n66), .Z(n52947) );
  XNOR U53525 ( .A(n53106), .B(n53107), .Z(n52945) );
  XNOR U53526 ( .A(n53108), .B(n53109), .Z(n53107) );
  NANDN U53527 ( .A(n52949), .B(n52951), .Z(n52982) );
  ANDN U53528 ( .B(B[75]), .A(n65), .Z(n52951) );
  XNOR U53529 ( .A(n53110), .B(n53111), .Z(n52949) );
  XNOR U53530 ( .A(n53112), .B(n53113), .Z(n53111) );
  NAND U53531 ( .A(n52953), .B(n52955), .Z(n52979) );
  ANDN U53532 ( .B(B[75]), .A(n64), .Z(n52955) );
  XNOR U53533 ( .A(n53114), .B(n53115), .Z(n52953) );
  XNOR U53534 ( .A(n53116), .B(n53117), .Z(n53115) );
  NANDN U53535 ( .A(n52957), .B(n52959), .Z(n52976) );
  ANDN U53536 ( .B(B[75]), .A(n63), .Z(n52959) );
  XNOR U53537 ( .A(n53118), .B(n53119), .Z(n52957) );
  XNOR U53538 ( .A(n53120), .B(n53121), .Z(n53119) );
  NAND U53539 ( .A(n52961), .B(n52963), .Z(n52973) );
  ANDN U53540 ( .B(B[75]), .A(n62), .Z(n52963) );
  XNOR U53541 ( .A(n53122), .B(n53123), .Z(n52961) );
  XNOR U53542 ( .A(n53124), .B(n53125), .Z(n53123) );
  NANDN U53543 ( .A(n52965), .B(n52967), .Z(n52970) );
  ANDN U53544 ( .B(B[75]), .A(n61), .Z(n52967) );
  XNOR U53545 ( .A(n53126), .B(n53127), .Z(n52965) );
  XNOR U53546 ( .A(n53128), .B(n53129), .Z(n53127) );
  ANDN U53547 ( .B(B[75]), .A(n60), .Z(n51863) );
  XNOR U53548 ( .A(n51871), .B(n53130), .Z(n51864) );
  XNOR U53549 ( .A(n51870), .B(n51868), .Z(n53130) );
  AND U53550 ( .A(n53131), .B(n53132), .Z(n51868) );
  NANDN U53551 ( .A(n53129), .B(n53133), .Z(n53132) );
  OR U53552 ( .A(n53128), .B(n53126), .Z(n53133) );
  AND U53553 ( .A(n53134), .B(n53135), .Z(n53129) );
  NANDN U53554 ( .A(n53125), .B(n53136), .Z(n53135) );
  NANDN U53555 ( .A(n53124), .B(n53122), .Z(n53136) );
  AND U53556 ( .A(n53137), .B(n53138), .Z(n53125) );
  NANDN U53557 ( .A(n53121), .B(n53139), .Z(n53138) );
  OR U53558 ( .A(n53120), .B(n53118), .Z(n53139) );
  AND U53559 ( .A(n53140), .B(n53141), .Z(n53121) );
  NANDN U53560 ( .A(n53117), .B(n53142), .Z(n53141) );
  NANDN U53561 ( .A(n53116), .B(n53114), .Z(n53142) );
  AND U53562 ( .A(n53143), .B(n53144), .Z(n53117) );
  NANDN U53563 ( .A(n53113), .B(n53145), .Z(n53144) );
  OR U53564 ( .A(n53112), .B(n53110), .Z(n53145) );
  AND U53565 ( .A(n53146), .B(n53147), .Z(n53113) );
  NANDN U53566 ( .A(n53109), .B(n53148), .Z(n53147) );
  NANDN U53567 ( .A(n53108), .B(n53106), .Z(n53148) );
  AND U53568 ( .A(n53149), .B(n53150), .Z(n53109) );
  NANDN U53569 ( .A(n53105), .B(n53151), .Z(n53150) );
  OR U53570 ( .A(n53104), .B(n53102), .Z(n53151) );
  AND U53571 ( .A(n53152), .B(n53153), .Z(n53105) );
  NANDN U53572 ( .A(n53101), .B(n53154), .Z(n53153) );
  NANDN U53573 ( .A(n53100), .B(n53098), .Z(n53154) );
  AND U53574 ( .A(n53155), .B(n53156), .Z(n53101) );
  NANDN U53575 ( .A(n53097), .B(n53157), .Z(n53156) );
  OR U53576 ( .A(n53096), .B(n53094), .Z(n53157) );
  AND U53577 ( .A(n53158), .B(n53159), .Z(n53097) );
  NANDN U53578 ( .A(n53093), .B(n53160), .Z(n53159) );
  NANDN U53579 ( .A(n53092), .B(n53090), .Z(n53160) );
  AND U53580 ( .A(n53161), .B(n53162), .Z(n53093) );
  NANDN U53581 ( .A(n53089), .B(n53163), .Z(n53162) );
  OR U53582 ( .A(n53088), .B(n53086), .Z(n53163) );
  AND U53583 ( .A(n53164), .B(n53165), .Z(n53089) );
  NANDN U53584 ( .A(n53085), .B(n53166), .Z(n53165) );
  NANDN U53585 ( .A(n53084), .B(n53082), .Z(n53166) );
  AND U53586 ( .A(n53167), .B(n53168), .Z(n53085) );
  NANDN U53587 ( .A(n53081), .B(n53169), .Z(n53168) );
  OR U53588 ( .A(n53080), .B(n53078), .Z(n53169) );
  AND U53589 ( .A(n53170), .B(n53171), .Z(n53081) );
  NANDN U53590 ( .A(n53077), .B(n53172), .Z(n53171) );
  NANDN U53591 ( .A(n53076), .B(n53074), .Z(n53172) );
  AND U53592 ( .A(n53173), .B(n53174), .Z(n53077) );
  NANDN U53593 ( .A(n53073), .B(n53175), .Z(n53174) );
  OR U53594 ( .A(n53072), .B(n53070), .Z(n53175) );
  AND U53595 ( .A(n53176), .B(n53177), .Z(n53073) );
  NANDN U53596 ( .A(n53069), .B(n53178), .Z(n53177) );
  NANDN U53597 ( .A(n53068), .B(n53066), .Z(n53178) );
  AND U53598 ( .A(n53179), .B(n53180), .Z(n53069) );
  NANDN U53599 ( .A(n53065), .B(n53181), .Z(n53180) );
  OR U53600 ( .A(n53064), .B(n53062), .Z(n53181) );
  AND U53601 ( .A(n53182), .B(n53183), .Z(n53065) );
  NANDN U53602 ( .A(n53061), .B(n53184), .Z(n53183) );
  NANDN U53603 ( .A(n53060), .B(n53058), .Z(n53184) );
  AND U53604 ( .A(n53185), .B(n53186), .Z(n53061) );
  NANDN U53605 ( .A(n53057), .B(n53187), .Z(n53186) );
  OR U53606 ( .A(n53056), .B(n53054), .Z(n53187) );
  AND U53607 ( .A(n53188), .B(n53189), .Z(n53057) );
  NANDN U53608 ( .A(n53053), .B(n53190), .Z(n53189) );
  NANDN U53609 ( .A(n53052), .B(n53050), .Z(n53190) );
  AND U53610 ( .A(n53191), .B(n53192), .Z(n53053) );
  NANDN U53611 ( .A(n53049), .B(n53193), .Z(n53192) );
  OR U53612 ( .A(n53048), .B(n53046), .Z(n53193) );
  AND U53613 ( .A(n53194), .B(n53195), .Z(n53049) );
  NANDN U53614 ( .A(n53044), .B(n53196), .Z(n53195) );
  NAND U53615 ( .A(n53042), .B(n53045), .Z(n53196) );
  NANDN U53616 ( .A(n53040), .B(n53197), .Z(n53044) );
  AND U53617 ( .A(A[0]), .B(B[77]), .Z(n53197) );
  NAND U53618 ( .A(B[76]), .B(A[1]), .Z(n53040) );
  XNOR U53619 ( .A(n53198), .B(n53199), .Z(n53042) );
  NAND U53620 ( .A(B[78]), .B(A[0]), .Z(n53199) );
  NAND U53621 ( .A(B[76]), .B(A[2]), .Z(n53045) );
  NAND U53622 ( .A(n53046), .B(n53048), .Z(n53191) );
  ANDN U53623 ( .B(B[76]), .A(n82), .Z(n53048) );
  XOR U53624 ( .A(n53200), .B(n53201), .Z(n53046) );
  XNOR U53625 ( .A(n53202), .B(n53203), .Z(n53201) );
  NANDN U53626 ( .A(n53050), .B(n53052), .Z(n53188) );
  ANDN U53627 ( .B(B[76]), .A(n81), .Z(n53052) );
  XNOR U53628 ( .A(n53204), .B(n53205), .Z(n53050) );
  XNOR U53629 ( .A(n53206), .B(n53207), .Z(n53205) );
  NAND U53630 ( .A(n53054), .B(n53056), .Z(n53185) );
  ANDN U53631 ( .B(B[76]), .A(n80), .Z(n53056) );
  XNOR U53632 ( .A(n53208), .B(n53209), .Z(n53054) );
  XNOR U53633 ( .A(n53210), .B(n53211), .Z(n53209) );
  NANDN U53634 ( .A(n53058), .B(n53060), .Z(n53182) );
  ANDN U53635 ( .B(B[76]), .A(n79), .Z(n53060) );
  XNOR U53636 ( .A(n53212), .B(n53213), .Z(n53058) );
  XNOR U53637 ( .A(n53214), .B(n53215), .Z(n53213) );
  NAND U53638 ( .A(n53062), .B(n53064), .Z(n53179) );
  ANDN U53639 ( .B(B[76]), .A(n78), .Z(n53064) );
  XNOR U53640 ( .A(n53216), .B(n53217), .Z(n53062) );
  XNOR U53641 ( .A(n53218), .B(n53219), .Z(n53217) );
  NANDN U53642 ( .A(n53066), .B(n53068), .Z(n53176) );
  ANDN U53643 ( .B(B[76]), .A(n77), .Z(n53068) );
  XNOR U53644 ( .A(n53220), .B(n53221), .Z(n53066) );
  XNOR U53645 ( .A(n53222), .B(n53223), .Z(n53221) );
  NAND U53646 ( .A(n53070), .B(n53072), .Z(n53173) );
  ANDN U53647 ( .B(B[76]), .A(n76), .Z(n53072) );
  XNOR U53648 ( .A(n53224), .B(n53225), .Z(n53070) );
  XNOR U53649 ( .A(n53226), .B(n53227), .Z(n53225) );
  NANDN U53650 ( .A(n53074), .B(n53076), .Z(n53170) );
  ANDN U53651 ( .B(B[76]), .A(n75), .Z(n53076) );
  XNOR U53652 ( .A(n53228), .B(n53229), .Z(n53074) );
  XNOR U53653 ( .A(n53230), .B(n53231), .Z(n53229) );
  NAND U53654 ( .A(n53078), .B(n53080), .Z(n53167) );
  ANDN U53655 ( .B(B[76]), .A(n74), .Z(n53080) );
  XNOR U53656 ( .A(n53232), .B(n53233), .Z(n53078) );
  XNOR U53657 ( .A(n53234), .B(n53235), .Z(n53233) );
  NANDN U53658 ( .A(n53082), .B(n53084), .Z(n53164) );
  ANDN U53659 ( .B(B[76]), .A(n73), .Z(n53084) );
  XNOR U53660 ( .A(n53236), .B(n53237), .Z(n53082) );
  XNOR U53661 ( .A(n53238), .B(n53239), .Z(n53237) );
  NAND U53662 ( .A(n53086), .B(n53088), .Z(n53161) );
  ANDN U53663 ( .B(B[76]), .A(n72), .Z(n53088) );
  XNOR U53664 ( .A(n53240), .B(n53241), .Z(n53086) );
  XNOR U53665 ( .A(n53242), .B(n53243), .Z(n53241) );
  NANDN U53666 ( .A(n53090), .B(n53092), .Z(n53158) );
  ANDN U53667 ( .B(B[76]), .A(n71), .Z(n53092) );
  XNOR U53668 ( .A(n53244), .B(n53245), .Z(n53090) );
  XNOR U53669 ( .A(n53246), .B(n53247), .Z(n53245) );
  NAND U53670 ( .A(n53094), .B(n53096), .Z(n53155) );
  ANDN U53671 ( .B(B[76]), .A(n70), .Z(n53096) );
  XNOR U53672 ( .A(n53248), .B(n53249), .Z(n53094) );
  XNOR U53673 ( .A(n53250), .B(n53251), .Z(n53249) );
  NANDN U53674 ( .A(n53098), .B(n53100), .Z(n53152) );
  ANDN U53675 ( .B(B[76]), .A(n69), .Z(n53100) );
  XNOR U53676 ( .A(n53252), .B(n53253), .Z(n53098) );
  XNOR U53677 ( .A(n53254), .B(n53255), .Z(n53253) );
  NAND U53678 ( .A(n53102), .B(n53104), .Z(n53149) );
  ANDN U53679 ( .B(B[76]), .A(n68), .Z(n53104) );
  XNOR U53680 ( .A(n53256), .B(n53257), .Z(n53102) );
  XNOR U53681 ( .A(n53258), .B(n53259), .Z(n53257) );
  NANDN U53682 ( .A(n53106), .B(n53108), .Z(n53146) );
  ANDN U53683 ( .B(B[76]), .A(n67), .Z(n53108) );
  XNOR U53684 ( .A(n53260), .B(n53261), .Z(n53106) );
  XNOR U53685 ( .A(n53262), .B(n53263), .Z(n53261) );
  NAND U53686 ( .A(n53110), .B(n53112), .Z(n53143) );
  ANDN U53687 ( .B(B[76]), .A(n66), .Z(n53112) );
  XNOR U53688 ( .A(n53264), .B(n53265), .Z(n53110) );
  XNOR U53689 ( .A(n53266), .B(n53267), .Z(n53265) );
  NANDN U53690 ( .A(n53114), .B(n53116), .Z(n53140) );
  ANDN U53691 ( .B(B[76]), .A(n65), .Z(n53116) );
  XNOR U53692 ( .A(n53268), .B(n53269), .Z(n53114) );
  XNOR U53693 ( .A(n53270), .B(n53271), .Z(n53269) );
  NAND U53694 ( .A(n53118), .B(n53120), .Z(n53137) );
  ANDN U53695 ( .B(B[76]), .A(n64), .Z(n53120) );
  XNOR U53696 ( .A(n53272), .B(n53273), .Z(n53118) );
  XNOR U53697 ( .A(n53274), .B(n53275), .Z(n53273) );
  NANDN U53698 ( .A(n53122), .B(n53124), .Z(n53134) );
  ANDN U53699 ( .B(B[76]), .A(n63), .Z(n53124) );
  XNOR U53700 ( .A(n53276), .B(n53277), .Z(n53122) );
  XNOR U53701 ( .A(n53278), .B(n53279), .Z(n53277) );
  NAND U53702 ( .A(n53126), .B(n53128), .Z(n53131) );
  ANDN U53703 ( .B(B[76]), .A(n62), .Z(n53128) );
  XNOR U53704 ( .A(n53280), .B(n53281), .Z(n53126) );
  XNOR U53705 ( .A(n53282), .B(n53283), .Z(n53281) );
  ANDN U53706 ( .B(B[76]), .A(n61), .Z(n51870) );
  XNOR U53707 ( .A(n51878), .B(n53284), .Z(n51871) );
  XNOR U53708 ( .A(n51877), .B(n51875), .Z(n53284) );
  AND U53709 ( .A(n53285), .B(n53286), .Z(n51875) );
  NANDN U53710 ( .A(n53283), .B(n53287), .Z(n53286) );
  NANDN U53711 ( .A(n53282), .B(n53280), .Z(n53287) );
  AND U53712 ( .A(n53288), .B(n53289), .Z(n53283) );
  NANDN U53713 ( .A(n53279), .B(n53290), .Z(n53289) );
  OR U53714 ( .A(n53278), .B(n53276), .Z(n53290) );
  AND U53715 ( .A(n53291), .B(n53292), .Z(n53279) );
  NANDN U53716 ( .A(n53275), .B(n53293), .Z(n53292) );
  NANDN U53717 ( .A(n53274), .B(n53272), .Z(n53293) );
  AND U53718 ( .A(n53294), .B(n53295), .Z(n53275) );
  NANDN U53719 ( .A(n53271), .B(n53296), .Z(n53295) );
  OR U53720 ( .A(n53270), .B(n53268), .Z(n53296) );
  AND U53721 ( .A(n53297), .B(n53298), .Z(n53271) );
  NANDN U53722 ( .A(n53267), .B(n53299), .Z(n53298) );
  NANDN U53723 ( .A(n53266), .B(n53264), .Z(n53299) );
  AND U53724 ( .A(n53300), .B(n53301), .Z(n53267) );
  NANDN U53725 ( .A(n53263), .B(n53302), .Z(n53301) );
  OR U53726 ( .A(n53262), .B(n53260), .Z(n53302) );
  AND U53727 ( .A(n53303), .B(n53304), .Z(n53263) );
  NANDN U53728 ( .A(n53259), .B(n53305), .Z(n53304) );
  NANDN U53729 ( .A(n53258), .B(n53256), .Z(n53305) );
  AND U53730 ( .A(n53306), .B(n53307), .Z(n53259) );
  NANDN U53731 ( .A(n53255), .B(n53308), .Z(n53307) );
  OR U53732 ( .A(n53254), .B(n53252), .Z(n53308) );
  AND U53733 ( .A(n53309), .B(n53310), .Z(n53255) );
  NANDN U53734 ( .A(n53251), .B(n53311), .Z(n53310) );
  NANDN U53735 ( .A(n53250), .B(n53248), .Z(n53311) );
  AND U53736 ( .A(n53312), .B(n53313), .Z(n53251) );
  NANDN U53737 ( .A(n53247), .B(n53314), .Z(n53313) );
  OR U53738 ( .A(n53246), .B(n53244), .Z(n53314) );
  AND U53739 ( .A(n53315), .B(n53316), .Z(n53247) );
  NANDN U53740 ( .A(n53243), .B(n53317), .Z(n53316) );
  NANDN U53741 ( .A(n53242), .B(n53240), .Z(n53317) );
  AND U53742 ( .A(n53318), .B(n53319), .Z(n53243) );
  NANDN U53743 ( .A(n53239), .B(n53320), .Z(n53319) );
  OR U53744 ( .A(n53238), .B(n53236), .Z(n53320) );
  AND U53745 ( .A(n53321), .B(n53322), .Z(n53239) );
  NANDN U53746 ( .A(n53235), .B(n53323), .Z(n53322) );
  NANDN U53747 ( .A(n53234), .B(n53232), .Z(n53323) );
  AND U53748 ( .A(n53324), .B(n53325), .Z(n53235) );
  NANDN U53749 ( .A(n53231), .B(n53326), .Z(n53325) );
  OR U53750 ( .A(n53230), .B(n53228), .Z(n53326) );
  AND U53751 ( .A(n53327), .B(n53328), .Z(n53231) );
  NANDN U53752 ( .A(n53227), .B(n53329), .Z(n53328) );
  NANDN U53753 ( .A(n53226), .B(n53224), .Z(n53329) );
  AND U53754 ( .A(n53330), .B(n53331), .Z(n53227) );
  NANDN U53755 ( .A(n53223), .B(n53332), .Z(n53331) );
  OR U53756 ( .A(n53222), .B(n53220), .Z(n53332) );
  AND U53757 ( .A(n53333), .B(n53334), .Z(n53223) );
  NANDN U53758 ( .A(n53219), .B(n53335), .Z(n53334) );
  NANDN U53759 ( .A(n53218), .B(n53216), .Z(n53335) );
  AND U53760 ( .A(n53336), .B(n53337), .Z(n53219) );
  NANDN U53761 ( .A(n53215), .B(n53338), .Z(n53337) );
  OR U53762 ( .A(n53214), .B(n53212), .Z(n53338) );
  AND U53763 ( .A(n53339), .B(n53340), .Z(n53215) );
  NANDN U53764 ( .A(n53211), .B(n53341), .Z(n53340) );
  NANDN U53765 ( .A(n53210), .B(n53208), .Z(n53341) );
  AND U53766 ( .A(n53342), .B(n53343), .Z(n53211) );
  NANDN U53767 ( .A(n53207), .B(n53344), .Z(n53343) );
  OR U53768 ( .A(n53206), .B(n53204), .Z(n53344) );
  AND U53769 ( .A(n53345), .B(n53346), .Z(n53207) );
  NANDN U53770 ( .A(n53202), .B(n53347), .Z(n53346) );
  NAND U53771 ( .A(n53200), .B(n53203), .Z(n53347) );
  NANDN U53772 ( .A(n53198), .B(n53348), .Z(n53202) );
  AND U53773 ( .A(A[0]), .B(B[78]), .Z(n53348) );
  NAND U53774 ( .A(B[77]), .B(A[1]), .Z(n53198) );
  XNOR U53775 ( .A(n53349), .B(n53350), .Z(n53200) );
  NAND U53776 ( .A(B[79]), .B(A[0]), .Z(n53350) );
  NAND U53777 ( .A(B[77]), .B(A[2]), .Z(n53203) );
  NAND U53778 ( .A(n53204), .B(n53206), .Z(n53342) );
  ANDN U53779 ( .B(B[77]), .A(n82), .Z(n53206) );
  XOR U53780 ( .A(n53351), .B(n53352), .Z(n53204) );
  XNOR U53781 ( .A(n53353), .B(n53354), .Z(n53352) );
  NANDN U53782 ( .A(n53208), .B(n53210), .Z(n53339) );
  ANDN U53783 ( .B(B[77]), .A(n81), .Z(n53210) );
  XNOR U53784 ( .A(n53355), .B(n53356), .Z(n53208) );
  XNOR U53785 ( .A(n53357), .B(n53358), .Z(n53356) );
  NAND U53786 ( .A(n53212), .B(n53214), .Z(n53336) );
  ANDN U53787 ( .B(B[77]), .A(n80), .Z(n53214) );
  XNOR U53788 ( .A(n53359), .B(n53360), .Z(n53212) );
  XNOR U53789 ( .A(n53361), .B(n53362), .Z(n53360) );
  NANDN U53790 ( .A(n53216), .B(n53218), .Z(n53333) );
  ANDN U53791 ( .B(B[77]), .A(n79), .Z(n53218) );
  XNOR U53792 ( .A(n53363), .B(n53364), .Z(n53216) );
  XNOR U53793 ( .A(n53365), .B(n53366), .Z(n53364) );
  NAND U53794 ( .A(n53220), .B(n53222), .Z(n53330) );
  ANDN U53795 ( .B(B[77]), .A(n78), .Z(n53222) );
  XNOR U53796 ( .A(n53367), .B(n53368), .Z(n53220) );
  XNOR U53797 ( .A(n53369), .B(n53370), .Z(n53368) );
  NANDN U53798 ( .A(n53224), .B(n53226), .Z(n53327) );
  ANDN U53799 ( .B(B[77]), .A(n77), .Z(n53226) );
  XNOR U53800 ( .A(n53371), .B(n53372), .Z(n53224) );
  XNOR U53801 ( .A(n53373), .B(n53374), .Z(n53372) );
  NAND U53802 ( .A(n53228), .B(n53230), .Z(n53324) );
  ANDN U53803 ( .B(B[77]), .A(n76), .Z(n53230) );
  XNOR U53804 ( .A(n53375), .B(n53376), .Z(n53228) );
  XNOR U53805 ( .A(n53377), .B(n53378), .Z(n53376) );
  NANDN U53806 ( .A(n53232), .B(n53234), .Z(n53321) );
  ANDN U53807 ( .B(B[77]), .A(n75), .Z(n53234) );
  XNOR U53808 ( .A(n53379), .B(n53380), .Z(n53232) );
  XNOR U53809 ( .A(n53381), .B(n53382), .Z(n53380) );
  NAND U53810 ( .A(n53236), .B(n53238), .Z(n53318) );
  ANDN U53811 ( .B(B[77]), .A(n74), .Z(n53238) );
  XNOR U53812 ( .A(n53383), .B(n53384), .Z(n53236) );
  XNOR U53813 ( .A(n53385), .B(n53386), .Z(n53384) );
  NANDN U53814 ( .A(n53240), .B(n53242), .Z(n53315) );
  ANDN U53815 ( .B(B[77]), .A(n73), .Z(n53242) );
  XNOR U53816 ( .A(n53387), .B(n53388), .Z(n53240) );
  XNOR U53817 ( .A(n53389), .B(n53390), .Z(n53388) );
  NAND U53818 ( .A(n53244), .B(n53246), .Z(n53312) );
  ANDN U53819 ( .B(B[77]), .A(n72), .Z(n53246) );
  XNOR U53820 ( .A(n53391), .B(n53392), .Z(n53244) );
  XNOR U53821 ( .A(n53393), .B(n53394), .Z(n53392) );
  NANDN U53822 ( .A(n53248), .B(n53250), .Z(n53309) );
  ANDN U53823 ( .B(B[77]), .A(n71), .Z(n53250) );
  XNOR U53824 ( .A(n53395), .B(n53396), .Z(n53248) );
  XNOR U53825 ( .A(n53397), .B(n53398), .Z(n53396) );
  NAND U53826 ( .A(n53252), .B(n53254), .Z(n53306) );
  ANDN U53827 ( .B(B[77]), .A(n70), .Z(n53254) );
  XNOR U53828 ( .A(n53399), .B(n53400), .Z(n53252) );
  XNOR U53829 ( .A(n53401), .B(n53402), .Z(n53400) );
  NANDN U53830 ( .A(n53256), .B(n53258), .Z(n53303) );
  ANDN U53831 ( .B(B[77]), .A(n69), .Z(n53258) );
  XNOR U53832 ( .A(n53403), .B(n53404), .Z(n53256) );
  XNOR U53833 ( .A(n53405), .B(n53406), .Z(n53404) );
  NAND U53834 ( .A(n53260), .B(n53262), .Z(n53300) );
  ANDN U53835 ( .B(B[77]), .A(n68), .Z(n53262) );
  XNOR U53836 ( .A(n53407), .B(n53408), .Z(n53260) );
  XNOR U53837 ( .A(n53409), .B(n53410), .Z(n53408) );
  NANDN U53838 ( .A(n53264), .B(n53266), .Z(n53297) );
  ANDN U53839 ( .B(B[77]), .A(n67), .Z(n53266) );
  XNOR U53840 ( .A(n53411), .B(n53412), .Z(n53264) );
  XNOR U53841 ( .A(n53413), .B(n53414), .Z(n53412) );
  NAND U53842 ( .A(n53268), .B(n53270), .Z(n53294) );
  ANDN U53843 ( .B(B[77]), .A(n66), .Z(n53270) );
  XNOR U53844 ( .A(n53415), .B(n53416), .Z(n53268) );
  XNOR U53845 ( .A(n53417), .B(n53418), .Z(n53416) );
  NANDN U53846 ( .A(n53272), .B(n53274), .Z(n53291) );
  ANDN U53847 ( .B(B[77]), .A(n65), .Z(n53274) );
  XNOR U53848 ( .A(n53419), .B(n53420), .Z(n53272) );
  XNOR U53849 ( .A(n53421), .B(n53422), .Z(n53420) );
  NAND U53850 ( .A(n53276), .B(n53278), .Z(n53288) );
  ANDN U53851 ( .B(B[77]), .A(n64), .Z(n53278) );
  XNOR U53852 ( .A(n53423), .B(n53424), .Z(n53276) );
  XNOR U53853 ( .A(n53425), .B(n53426), .Z(n53424) );
  NANDN U53854 ( .A(n53280), .B(n53282), .Z(n53285) );
  ANDN U53855 ( .B(B[77]), .A(n63), .Z(n53282) );
  XNOR U53856 ( .A(n53427), .B(n53428), .Z(n53280) );
  XNOR U53857 ( .A(n53429), .B(n53430), .Z(n53428) );
  ANDN U53858 ( .B(B[77]), .A(n62), .Z(n51877) );
  XNOR U53859 ( .A(n51885), .B(n53431), .Z(n51878) );
  XNOR U53860 ( .A(n51884), .B(n51882), .Z(n53431) );
  AND U53861 ( .A(n53432), .B(n53433), .Z(n51882) );
  NANDN U53862 ( .A(n53430), .B(n53434), .Z(n53433) );
  OR U53863 ( .A(n53429), .B(n53427), .Z(n53434) );
  AND U53864 ( .A(n53435), .B(n53436), .Z(n53430) );
  NANDN U53865 ( .A(n53426), .B(n53437), .Z(n53436) );
  NANDN U53866 ( .A(n53425), .B(n53423), .Z(n53437) );
  AND U53867 ( .A(n53438), .B(n53439), .Z(n53426) );
  NANDN U53868 ( .A(n53422), .B(n53440), .Z(n53439) );
  OR U53869 ( .A(n53421), .B(n53419), .Z(n53440) );
  AND U53870 ( .A(n53441), .B(n53442), .Z(n53422) );
  NANDN U53871 ( .A(n53418), .B(n53443), .Z(n53442) );
  NANDN U53872 ( .A(n53417), .B(n53415), .Z(n53443) );
  AND U53873 ( .A(n53444), .B(n53445), .Z(n53418) );
  NANDN U53874 ( .A(n53414), .B(n53446), .Z(n53445) );
  OR U53875 ( .A(n53413), .B(n53411), .Z(n53446) );
  AND U53876 ( .A(n53447), .B(n53448), .Z(n53414) );
  NANDN U53877 ( .A(n53410), .B(n53449), .Z(n53448) );
  NANDN U53878 ( .A(n53409), .B(n53407), .Z(n53449) );
  AND U53879 ( .A(n53450), .B(n53451), .Z(n53410) );
  NANDN U53880 ( .A(n53406), .B(n53452), .Z(n53451) );
  OR U53881 ( .A(n53405), .B(n53403), .Z(n53452) );
  AND U53882 ( .A(n53453), .B(n53454), .Z(n53406) );
  NANDN U53883 ( .A(n53402), .B(n53455), .Z(n53454) );
  NANDN U53884 ( .A(n53401), .B(n53399), .Z(n53455) );
  AND U53885 ( .A(n53456), .B(n53457), .Z(n53402) );
  NANDN U53886 ( .A(n53398), .B(n53458), .Z(n53457) );
  OR U53887 ( .A(n53397), .B(n53395), .Z(n53458) );
  AND U53888 ( .A(n53459), .B(n53460), .Z(n53398) );
  NANDN U53889 ( .A(n53394), .B(n53461), .Z(n53460) );
  NANDN U53890 ( .A(n53393), .B(n53391), .Z(n53461) );
  AND U53891 ( .A(n53462), .B(n53463), .Z(n53394) );
  NANDN U53892 ( .A(n53390), .B(n53464), .Z(n53463) );
  OR U53893 ( .A(n53389), .B(n53387), .Z(n53464) );
  AND U53894 ( .A(n53465), .B(n53466), .Z(n53390) );
  NANDN U53895 ( .A(n53386), .B(n53467), .Z(n53466) );
  NANDN U53896 ( .A(n53385), .B(n53383), .Z(n53467) );
  AND U53897 ( .A(n53468), .B(n53469), .Z(n53386) );
  NANDN U53898 ( .A(n53382), .B(n53470), .Z(n53469) );
  OR U53899 ( .A(n53381), .B(n53379), .Z(n53470) );
  AND U53900 ( .A(n53471), .B(n53472), .Z(n53382) );
  NANDN U53901 ( .A(n53378), .B(n53473), .Z(n53472) );
  NANDN U53902 ( .A(n53377), .B(n53375), .Z(n53473) );
  AND U53903 ( .A(n53474), .B(n53475), .Z(n53378) );
  NANDN U53904 ( .A(n53374), .B(n53476), .Z(n53475) );
  OR U53905 ( .A(n53373), .B(n53371), .Z(n53476) );
  AND U53906 ( .A(n53477), .B(n53478), .Z(n53374) );
  NANDN U53907 ( .A(n53370), .B(n53479), .Z(n53478) );
  NANDN U53908 ( .A(n53369), .B(n53367), .Z(n53479) );
  AND U53909 ( .A(n53480), .B(n53481), .Z(n53370) );
  NANDN U53910 ( .A(n53366), .B(n53482), .Z(n53481) );
  OR U53911 ( .A(n53365), .B(n53363), .Z(n53482) );
  AND U53912 ( .A(n53483), .B(n53484), .Z(n53366) );
  NANDN U53913 ( .A(n53362), .B(n53485), .Z(n53484) );
  NANDN U53914 ( .A(n53361), .B(n53359), .Z(n53485) );
  AND U53915 ( .A(n53486), .B(n53487), .Z(n53362) );
  NANDN U53916 ( .A(n53358), .B(n53488), .Z(n53487) );
  OR U53917 ( .A(n53357), .B(n53355), .Z(n53488) );
  AND U53918 ( .A(n53489), .B(n53490), .Z(n53358) );
  NANDN U53919 ( .A(n53353), .B(n53491), .Z(n53490) );
  NAND U53920 ( .A(n53351), .B(n53354), .Z(n53491) );
  NANDN U53921 ( .A(n53349), .B(n53492), .Z(n53353) );
  AND U53922 ( .A(A[0]), .B(B[79]), .Z(n53492) );
  NAND U53923 ( .A(B[78]), .B(A[1]), .Z(n53349) );
  XNOR U53924 ( .A(n53493), .B(n53494), .Z(n53351) );
  NAND U53925 ( .A(B[80]), .B(A[0]), .Z(n53494) );
  NAND U53926 ( .A(B[78]), .B(A[2]), .Z(n53354) );
  NAND U53927 ( .A(n53355), .B(n53357), .Z(n53486) );
  ANDN U53928 ( .B(B[78]), .A(n82), .Z(n53357) );
  XOR U53929 ( .A(n53495), .B(n53496), .Z(n53355) );
  XNOR U53930 ( .A(n53497), .B(n53498), .Z(n53496) );
  NANDN U53931 ( .A(n53359), .B(n53361), .Z(n53483) );
  ANDN U53932 ( .B(B[78]), .A(n81), .Z(n53361) );
  XNOR U53933 ( .A(n53499), .B(n53500), .Z(n53359) );
  XNOR U53934 ( .A(n53501), .B(n53502), .Z(n53500) );
  NAND U53935 ( .A(n53363), .B(n53365), .Z(n53480) );
  ANDN U53936 ( .B(B[78]), .A(n80), .Z(n53365) );
  XNOR U53937 ( .A(n53503), .B(n53504), .Z(n53363) );
  XNOR U53938 ( .A(n53505), .B(n53506), .Z(n53504) );
  NANDN U53939 ( .A(n53367), .B(n53369), .Z(n53477) );
  ANDN U53940 ( .B(B[78]), .A(n79), .Z(n53369) );
  XNOR U53941 ( .A(n53507), .B(n53508), .Z(n53367) );
  XNOR U53942 ( .A(n53509), .B(n53510), .Z(n53508) );
  NAND U53943 ( .A(n53371), .B(n53373), .Z(n53474) );
  ANDN U53944 ( .B(B[78]), .A(n78), .Z(n53373) );
  XNOR U53945 ( .A(n53511), .B(n53512), .Z(n53371) );
  XNOR U53946 ( .A(n53513), .B(n53514), .Z(n53512) );
  NANDN U53947 ( .A(n53375), .B(n53377), .Z(n53471) );
  ANDN U53948 ( .B(B[78]), .A(n77), .Z(n53377) );
  XNOR U53949 ( .A(n53515), .B(n53516), .Z(n53375) );
  XNOR U53950 ( .A(n53517), .B(n53518), .Z(n53516) );
  NAND U53951 ( .A(n53379), .B(n53381), .Z(n53468) );
  ANDN U53952 ( .B(B[78]), .A(n76), .Z(n53381) );
  XNOR U53953 ( .A(n53519), .B(n53520), .Z(n53379) );
  XNOR U53954 ( .A(n53521), .B(n53522), .Z(n53520) );
  NANDN U53955 ( .A(n53383), .B(n53385), .Z(n53465) );
  ANDN U53956 ( .B(B[78]), .A(n75), .Z(n53385) );
  XNOR U53957 ( .A(n53523), .B(n53524), .Z(n53383) );
  XNOR U53958 ( .A(n53525), .B(n53526), .Z(n53524) );
  NAND U53959 ( .A(n53387), .B(n53389), .Z(n53462) );
  ANDN U53960 ( .B(B[78]), .A(n74), .Z(n53389) );
  XNOR U53961 ( .A(n53527), .B(n53528), .Z(n53387) );
  XNOR U53962 ( .A(n53529), .B(n53530), .Z(n53528) );
  NANDN U53963 ( .A(n53391), .B(n53393), .Z(n53459) );
  ANDN U53964 ( .B(B[78]), .A(n73), .Z(n53393) );
  XNOR U53965 ( .A(n53531), .B(n53532), .Z(n53391) );
  XNOR U53966 ( .A(n53533), .B(n53534), .Z(n53532) );
  NAND U53967 ( .A(n53395), .B(n53397), .Z(n53456) );
  ANDN U53968 ( .B(B[78]), .A(n72), .Z(n53397) );
  XNOR U53969 ( .A(n53535), .B(n53536), .Z(n53395) );
  XNOR U53970 ( .A(n53537), .B(n53538), .Z(n53536) );
  NANDN U53971 ( .A(n53399), .B(n53401), .Z(n53453) );
  ANDN U53972 ( .B(B[78]), .A(n71), .Z(n53401) );
  XNOR U53973 ( .A(n53539), .B(n53540), .Z(n53399) );
  XNOR U53974 ( .A(n53541), .B(n53542), .Z(n53540) );
  NAND U53975 ( .A(n53403), .B(n53405), .Z(n53450) );
  ANDN U53976 ( .B(B[78]), .A(n70), .Z(n53405) );
  XNOR U53977 ( .A(n53543), .B(n53544), .Z(n53403) );
  XNOR U53978 ( .A(n53545), .B(n53546), .Z(n53544) );
  NANDN U53979 ( .A(n53407), .B(n53409), .Z(n53447) );
  ANDN U53980 ( .B(B[78]), .A(n69), .Z(n53409) );
  XNOR U53981 ( .A(n53547), .B(n53548), .Z(n53407) );
  XNOR U53982 ( .A(n53549), .B(n53550), .Z(n53548) );
  NAND U53983 ( .A(n53411), .B(n53413), .Z(n53444) );
  ANDN U53984 ( .B(B[78]), .A(n68), .Z(n53413) );
  XNOR U53985 ( .A(n53551), .B(n53552), .Z(n53411) );
  XNOR U53986 ( .A(n53553), .B(n53554), .Z(n53552) );
  NANDN U53987 ( .A(n53415), .B(n53417), .Z(n53441) );
  ANDN U53988 ( .B(B[78]), .A(n67), .Z(n53417) );
  XNOR U53989 ( .A(n53555), .B(n53556), .Z(n53415) );
  XNOR U53990 ( .A(n53557), .B(n53558), .Z(n53556) );
  NAND U53991 ( .A(n53419), .B(n53421), .Z(n53438) );
  ANDN U53992 ( .B(B[78]), .A(n66), .Z(n53421) );
  XNOR U53993 ( .A(n53559), .B(n53560), .Z(n53419) );
  XNOR U53994 ( .A(n53561), .B(n53562), .Z(n53560) );
  NANDN U53995 ( .A(n53423), .B(n53425), .Z(n53435) );
  ANDN U53996 ( .B(B[78]), .A(n65), .Z(n53425) );
  XNOR U53997 ( .A(n53563), .B(n53564), .Z(n53423) );
  XNOR U53998 ( .A(n53565), .B(n53566), .Z(n53564) );
  NAND U53999 ( .A(n53427), .B(n53429), .Z(n53432) );
  ANDN U54000 ( .B(B[78]), .A(n64), .Z(n53429) );
  XNOR U54001 ( .A(n53567), .B(n53568), .Z(n53427) );
  XNOR U54002 ( .A(n53569), .B(n53570), .Z(n53568) );
  ANDN U54003 ( .B(B[78]), .A(n63), .Z(n51884) );
  XNOR U54004 ( .A(n51892), .B(n53571), .Z(n51885) );
  XNOR U54005 ( .A(n51891), .B(n51889), .Z(n53571) );
  AND U54006 ( .A(n53572), .B(n53573), .Z(n51889) );
  NANDN U54007 ( .A(n53570), .B(n53574), .Z(n53573) );
  NANDN U54008 ( .A(n53569), .B(n53567), .Z(n53574) );
  AND U54009 ( .A(n53575), .B(n53576), .Z(n53570) );
  NANDN U54010 ( .A(n53566), .B(n53577), .Z(n53576) );
  OR U54011 ( .A(n53565), .B(n53563), .Z(n53577) );
  AND U54012 ( .A(n53578), .B(n53579), .Z(n53566) );
  NANDN U54013 ( .A(n53562), .B(n53580), .Z(n53579) );
  NANDN U54014 ( .A(n53561), .B(n53559), .Z(n53580) );
  AND U54015 ( .A(n53581), .B(n53582), .Z(n53562) );
  NANDN U54016 ( .A(n53558), .B(n53583), .Z(n53582) );
  OR U54017 ( .A(n53557), .B(n53555), .Z(n53583) );
  AND U54018 ( .A(n53584), .B(n53585), .Z(n53558) );
  NANDN U54019 ( .A(n53554), .B(n53586), .Z(n53585) );
  NANDN U54020 ( .A(n53553), .B(n53551), .Z(n53586) );
  AND U54021 ( .A(n53587), .B(n53588), .Z(n53554) );
  NANDN U54022 ( .A(n53550), .B(n53589), .Z(n53588) );
  OR U54023 ( .A(n53549), .B(n53547), .Z(n53589) );
  AND U54024 ( .A(n53590), .B(n53591), .Z(n53550) );
  NANDN U54025 ( .A(n53546), .B(n53592), .Z(n53591) );
  NANDN U54026 ( .A(n53545), .B(n53543), .Z(n53592) );
  AND U54027 ( .A(n53593), .B(n53594), .Z(n53546) );
  NANDN U54028 ( .A(n53542), .B(n53595), .Z(n53594) );
  OR U54029 ( .A(n53541), .B(n53539), .Z(n53595) );
  AND U54030 ( .A(n53596), .B(n53597), .Z(n53542) );
  NANDN U54031 ( .A(n53538), .B(n53598), .Z(n53597) );
  NANDN U54032 ( .A(n53537), .B(n53535), .Z(n53598) );
  AND U54033 ( .A(n53599), .B(n53600), .Z(n53538) );
  NANDN U54034 ( .A(n53534), .B(n53601), .Z(n53600) );
  OR U54035 ( .A(n53533), .B(n53531), .Z(n53601) );
  AND U54036 ( .A(n53602), .B(n53603), .Z(n53534) );
  NANDN U54037 ( .A(n53530), .B(n53604), .Z(n53603) );
  NANDN U54038 ( .A(n53529), .B(n53527), .Z(n53604) );
  AND U54039 ( .A(n53605), .B(n53606), .Z(n53530) );
  NANDN U54040 ( .A(n53526), .B(n53607), .Z(n53606) );
  OR U54041 ( .A(n53525), .B(n53523), .Z(n53607) );
  AND U54042 ( .A(n53608), .B(n53609), .Z(n53526) );
  NANDN U54043 ( .A(n53522), .B(n53610), .Z(n53609) );
  NANDN U54044 ( .A(n53521), .B(n53519), .Z(n53610) );
  AND U54045 ( .A(n53611), .B(n53612), .Z(n53522) );
  NANDN U54046 ( .A(n53518), .B(n53613), .Z(n53612) );
  OR U54047 ( .A(n53517), .B(n53515), .Z(n53613) );
  AND U54048 ( .A(n53614), .B(n53615), .Z(n53518) );
  NANDN U54049 ( .A(n53514), .B(n53616), .Z(n53615) );
  NANDN U54050 ( .A(n53513), .B(n53511), .Z(n53616) );
  AND U54051 ( .A(n53617), .B(n53618), .Z(n53514) );
  NANDN U54052 ( .A(n53510), .B(n53619), .Z(n53618) );
  OR U54053 ( .A(n53509), .B(n53507), .Z(n53619) );
  AND U54054 ( .A(n53620), .B(n53621), .Z(n53510) );
  NANDN U54055 ( .A(n53506), .B(n53622), .Z(n53621) );
  NANDN U54056 ( .A(n53505), .B(n53503), .Z(n53622) );
  AND U54057 ( .A(n53623), .B(n53624), .Z(n53506) );
  NANDN U54058 ( .A(n53502), .B(n53625), .Z(n53624) );
  OR U54059 ( .A(n53501), .B(n53499), .Z(n53625) );
  AND U54060 ( .A(n53626), .B(n53627), .Z(n53502) );
  NANDN U54061 ( .A(n53497), .B(n53628), .Z(n53627) );
  NAND U54062 ( .A(n53495), .B(n53498), .Z(n53628) );
  NANDN U54063 ( .A(n53493), .B(n53629), .Z(n53497) );
  AND U54064 ( .A(A[0]), .B(B[80]), .Z(n53629) );
  NAND U54065 ( .A(B[79]), .B(A[1]), .Z(n53493) );
  XNOR U54066 ( .A(n53630), .B(n53631), .Z(n53495) );
  NAND U54067 ( .A(B[81]), .B(A[0]), .Z(n53631) );
  NAND U54068 ( .A(B[79]), .B(A[2]), .Z(n53498) );
  NAND U54069 ( .A(n53499), .B(n53501), .Z(n53623) );
  ANDN U54070 ( .B(B[79]), .A(n82), .Z(n53501) );
  XOR U54071 ( .A(n53632), .B(n53633), .Z(n53499) );
  XNOR U54072 ( .A(n53634), .B(n53635), .Z(n53633) );
  NANDN U54073 ( .A(n53503), .B(n53505), .Z(n53620) );
  ANDN U54074 ( .B(B[79]), .A(n81), .Z(n53505) );
  XNOR U54075 ( .A(n53636), .B(n53637), .Z(n53503) );
  XNOR U54076 ( .A(n53638), .B(n53639), .Z(n53637) );
  NAND U54077 ( .A(n53507), .B(n53509), .Z(n53617) );
  ANDN U54078 ( .B(B[79]), .A(n80), .Z(n53509) );
  XNOR U54079 ( .A(n53640), .B(n53641), .Z(n53507) );
  XNOR U54080 ( .A(n53642), .B(n53643), .Z(n53641) );
  NANDN U54081 ( .A(n53511), .B(n53513), .Z(n53614) );
  ANDN U54082 ( .B(B[79]), .A(n79), .Z(n53513) );
  XNOR U54083 ( .A(n53644), .B(n53645), .Z(n53511) );
  XNOR U54084 ( .A(n53646), .B(n53647), .Z(n53645) );
  NAND U54085 ( .A(n53515), .B(n53517), .Z(n53611) );
  ANDN U54086 ( .B(B[79]), .A(n78), .Z(n53517) );
  XNOR U54087 ( .A(n53648), .B(n53649), .Z(n53515) );
  XNOR U54088 ( .A(n53650), .B(n53651), .Z(n53649) );
  NANDN U54089 ( .A(n53519), .B(n53521), .Z(n53608) );
  ANDN U54090 ( .B(B[79]), .A(n77), .Z(n53521) );
  XNOR U54091 ( .A(n53652), .B(n53653), .Z(n53519) );
  XNOR U54092 ( .A(n53654), .B(n53655), .Z(n53653) );
  NAND U54093 ( .A(n53523), .B(n53525), .Z(n53605) );
  ANDN U54094 ( .B(B[79]), .A(n76), .Z(n53525) );
  XNOR U54095 ( .A(n53656), .B(n53657), .Z(n53523) );
  XNOR U54096 ( .A(n53658), .B(n53659), .Z(n53657) );
  NANDN U54097 ( .A(n53527), .B(n53529), .Z(n53602) );
  ANDN U54098 ( .B(B[79]), .A(n75), .Z(n53529) );
  XNOR U54099 ( .A(n53660), .B(n53661), .Z(n53527) );
  XNOR U54100 ( .A(n53662), .B(n53663), .Z(n53661) );
  NAND U54101 ( .A(n53531), .B(n53533), .Z(n53599) );
  ANDN U54102 ( .B(B[79]), .A(n74), .Z(n53533) );
  XNOR U54103 ( .A(n53664), .B(n53665), .Z(n53531) );
  XNOR U54104 ( .A(n53666), .B(n53667), .Z(n53665) );
  NANDN U54105 ( .A(n53535), .B(n53537), .Z(n53596) );
  ANDN U54106 ( .B(B[79]), .A(n73), .Z(n53537) );
  XNOR U54107 ( .A(n53668), .B(n53669), .Z(n53535) );
  XNOR U54108 ( .A(n53670), .B(n53671), .Z(n53669) );
  NAND U54109 ( .A(n53539), .B(n53541), .Z(n53593) );
  ANDN U54110 ( .B(B[79]), .A(n72), .Z(n53541) );
  XNOR U54111 ( .A(n53672), .B(n53673), .Z(n53539) );
  XNOR U54112 ( .A(n53674), .B(n53675), .Z(n53673) );
  NANDN U54113 ( .A(n53543), .B(n53545), .Z(n53590) );
  ANDN U54114 ( .B(B[79]), .A(n71), .Z(n53545) );
  XNOR U54115 ( .A(n53676), .B(n53677), .Z(n53543) );
  XNOR U54116 ( .A(n53678), .B(n53679), .Z(n53677) );
  NAND U54117 ( .A(n53547), .B(n53549), .Z(n53587) );
  ANDN U54118 ( .B(B[79]), .A(n70), .Z(n53549) );
  XNOR U54119 ( .A(n53680), .B(n53681), .Z(n53547) );
  XNOR U54120 ( .A(n53682), .B(n53683), .Z(n53681) );
  NANDN U54121 ( .A(n53551), .B(n53553), .Z(n53584) );
  ANDN U54122 ( .B(B[79]), .A(n69), .Z(n53553) );
  XNOR U54123 ( .A(n53684), .B(n53685), .Z(n53551) );
  XNOR U54124 ( .A(n53686), .B(n53687), .Z(n53685) );
  NAND U54125 ( .A(n53555), .B(n53557), .Z(n53581) );
  ANDN U54126 ( .B(B[79]), .A(n68), .Z(n53557) );
  XNOR U54127 ( .A(n53688), .B(n53689), .Z(n53555) );
  XNOR U54128 ( .A(n53690), .B(n53691), .Z(n53689) );
  NANDN U54129 ( .A(n53559), .B(n53561), .Z(n53578) );
  ANDN U54130 ( .B(B[79]), .A(n67), .Z(n53561) );
  XNOR U54131 ( .A(n53692), .B(n53693), .Z(n53559) );
  XNOR U54132 ( .A(n53694), .B(n53695), .Z(n53693) );
  NAND U54133 ( .A(n53563), .B(n53565), .Z(n53575) );
  ANDN U54134 ( .B(B[79]), .A(n66), .Z(n53565) );
  XNOR U54135 ( .A(n53696), .B(n53697), .Z(n53563) );
  XNOR U54136 ( .A(n53698), .B(n53699), .Z(n53697) );
  NANDN U54137 ( .A(n53567), .B(n53569), .Z(n53572) );
  ANDN U54138 ( .B(B[79]), .A(n65), .Z(n53569) );
  XNOR U54139 ( .A(n53700), .B(n53701), .Z(n53567) );
  XNOR U54140 ( .A(n53702), .B(n53703), .Z(n53701) );
  ANDN U54141 ( .B(B[79]), .A(n64), .Z(n51891) );
  XNOR U54142 ( .A(n51899), .B(n53704), .Z(n51892) );
  XNOR U54143 ( .A(n51898), .B(n51896), .Z(n53704) );
  AND U54144 ( .A(n53705), .B(n53706), .Z(n51896) );
  NANDN U54145 ( .A(n53703), .B(n53707), .Z(n53706) );
  OR U54146 ( .A(n53702), .B(n53700), .Z(n53707) );
  AND U54147 ( .A(n53708), .B(n53709), .Z(n53703) );
  NANDN U54148 ( .A(n53699), .B(n53710), .Z(n53709) );
  NANDN U54149 ( .A(n53698), .B(n53696), .Z(n53710) );
  AND U54150 ( .A(n53711), .B(n53712), .Z(n53699) );
  NANDN U54151 ( .A(n53695), .B(n53713), .Z(n53712) );
  OR U54152 ( .A(n53694), .B(n53692), .Z(n53713) );
  AND U54153 ( .A(n53714), .B(n53715), .Z(n53695) );
  NANDN U54154 ( .A(n53691), .B(n53716), .Z(n53715) );
  NANDN U54155 ( .A(n53690), .B(n53688), .Z(n53716) );
  AND U54156 ( .A(n53717), .B(n53718), .Z(n53691) );
  NANDN U54157 ( .A(n53687), .B(n53719), .Z(n53718) );
  OR U54158 ( .A(n53686), .B(n53684), .Z(n53719) );
  AND U54159 ( .A(n53720), .B(n53721), .Z(n53687) );
  NANDN U54160 ( .A(n53683), .B(n53722), .Z(n53721) );
  NANDN U54161 ( .A(n53682), .B(n53680), .Z(n53722) );
  AND U54162 ( .A(n53723), .B(n53724), .Z(n53683) );
  NANDN U54163 ( .A(n53679), .B(n53725), .Z(n53724) );
  OR U54164 ( .A(n53678), .B(n53676), .Z(n53725) );
  AND U54165 ( .A(n53726), .B(n53727), .Z(n53679) );
  NANDN U54166 ( .A(n53675), .B(n53728), .Z(n53727) );
  NANDN U54167 ( .A(n53674), .B(n53672), .Z(n53728) );
  AND U54168 ( .A(n53729), .B(n53730), .Z(n53675) );
  NANDN U54169 ( .A(n53671), .B(n53731), .Z(n53730) );
  OR U54170 ( .A(n53670), .B(n53668), .Z(n53731) );
  AND U54171 ( .A(n53732), .B(n53733), .Z(n53671) );
  NANDN U54172 ( .A(n53667), .B(n53734), .Z(n53733) );
  NANDN U54173 ( .A(n53666), .B(n53664), .Z(n53734) );
  AND U54174 ( .A(n53735), .B(n53736), .Z(n53667) );
  NANDN U54175 ( .A(n53663), .B(n53737), .Z(n53736) );
  OR U54176 ( .A(n53662), .B(n53660), .Z(n53737) );
  AND U54177 ( .A(n53738), .B(n53739), .Z(n53663) );
  NANDN U54178 ( .A(n53659), .B(n53740), .Z(n53739) );
  NANDN U54179 ( .A(n53658), .B(n53656), .Z(n53740) );
  AND U54180 ( .A(n53741), .B(n53742), .Z(n53659) );
  NANDN U54181 ( .A(n53655), .B(n53743), .Z(n53742) );
  OR U54182 ( .A(n53654), .B(n53652), .Z(n53743) );
  AND U54183 ( .A(n53744), .B(n53745), .Z(n53655) );
  NANDN U54184 ( .A(n53651), .B(n53746), .Z(n53745) );
  NANDN U54185 ( .A(n53650), .B(n53648), .Z(n53746) );
  AND U54186 ( .A(n53747), .B(n53748), .Z(n53651) );
  NANDN U54187 ( .A(n53647), .B(n53749), .Z(n53748) );
  OR U54188 ( .A(n53646), .B(n53644), .Z(n53749) );
  AND U54189 ( .A(n53750), .B(n53751), .Z(n53647) );
  NANDN U54190 ( .A(n53643), .B(n53752), .Z(n53751) );
  NANDN U54191 ( .A(n53642), .B(n53640), .Z(n53752) );
  AND U54192 ( .A(n53753), .B(n53754), .Z(n53643) );
  NANDN U54193 ( .A(n53639), .B(n53755), .Z(n53754) );
  OR U54194 ( .A(n53638), .B(n53636), .Z(n53755) );
  AND U54195 ( .A(n53756), .B(n53757), .Z(n53639) );
  NANDN U54196 ( .A(n53634), .B(n53758), .Z(n53757) );
  NAND U54197 ( .A(n53632), .B(n53635), .Z(n53758) );
  NANDN U54198 ( .A(n53630), .B(n53759), .Z(n53634) );
  AND U54199 ( .A(A[0]), .B(B[81]), .Z(n53759) );
  NAND U54200 ( .A(B[80]), .B(A[1]), .Z(n53630) );
  XNOR U54201 ( .A(n53760), .B(n53761), .Z(n53632) );
  NAND U54202 ( .A(B[82]), .B(A[0]), .Z(n53761) );
  NAND U54203 ( .A(B[80]), .B(A[2]), .Z(n53635) );
  NAND U54204 ( .A(n53636), .B(n53638), .Z(n53753) );
  ANDN U54205 ( .B(B[80]), .A(n82), .Z(n53638) );
  XOR U54206 ( .A(n53762), .B(n53763), .Z(n53636) );
  XNOR U54207 ( .A(n53764), .B(n53765), .Z(n53763) );
  NANDN U54208 ( .A(n53640), .B(n53642), .Z(n53750) );
  ANDN U54209 ( .B(B[80]), .A(n81), .Z(n53642) );
  XNOR U54210 ( .A(n53766), .B(n53767), .Z(n53640) );
  XNOR U54211 ( .A(n53768), .B(n53769), .Z(n53767) );
  NAND U54212 ( .A(n53644), .B(n53646), .Z(n53747) );
  ANDN U54213 ( .B(B[80]), .A(n80), .Z(n53646) );
  XNOR U54214 ( .A(n53770), .B(n53771), .Z(n53644) );
  XNOR U54215 ( .A(n53772), .B(n53773), .Z(n53771) );
  NANDN U54216 ( .A(n53648), .B(n53650), .Z(n53744) );
  ANDN U54217 ( .B(B[80]), .A(n79), .Z(n53650) );
  XNOR U54218 ( .A(n53774), .B(n53775), .Z(n53648) );
  XNOR U54219 ( .A(n53776), .B(n53777), .Z(n53775) );
  NAND U54220 ( .A(n53652), .B(n53654), .Z(n53741) );
  ANDN U54221 ( .B(B[80]), .A(n78), .Z(n53654) );
  XNOR U54222 ( .A(n53778), .B(n53779), .Z(n53652) );
  XNOR U54223 ( .A(n53780), .B(n53781), .Z(n53779) );
  NANDN U54224 ( .A(n53656), .B(n53658), .Z(n53738) );
  ANDN U54225 ( .B(B[80]), .A(n77), .Z(n53658) );
  XNOR U54226 ( .A(n53782), .B(n53783), .Z(n53656) );
  XNOR U54227 ( .A(n53784), .B(n53785), .Z(n53783) );
  NAND U54228 ( .A(n53660), .B(n53662), .Z(n53735) );
  ANDN U54229 ( .B(B[80]), .A(n76), .Z(n53662) );
  XNOR U54230 ( .A(n53786), .B(n53787), .Z(n53660) );
  XNOR U54231 ( .A(n53788), .B(n53789), .Z(n53787) );
  NANDN U54232 ( .A(n53664), .B(n53666), .Z(n53732) );
  ANDN U54233 ( .B(B[80]), .A(n75), .Z(n53666) );
  XNOR U54234 ( .A(n53790), .B(n53791), .Z(n53664) );
  XNOR U54235 ( .A(n53792), .B(n53793), .Z(n53791) );
  NAND U54236 ( .A(n53668), .B(n53670), .Z(n53729) );
  ANDN U54237 ( .B(B[80]), .A(n74), .Z(n53670) );
  XNOR U54238 ( .A(n53794), .B(n53795), .Z(n53668) );
  XNOR U54239 ( .A(n53796), .B(n53797), .Z(n53795) );
  NANDN U54240 ( .A(n53672), .B(n53674), .Z(n53726) );
  ANDN U54241 ( .B(B[80]), .A(n73), .Z(n53674) );
  XNOR U54242 ( .A(n53798), .B(n53799), .Z(n53672) );
  XNOR U54243 ( .A(n53800), .B(n53801), .Z(n53799) );
  NAND U54244 ( .A(n53676), .B(n53678), .Z(n53723) );
  ANDN U54245 ( .B(B[80]), .A(n72), .Z(n53678) );
  XNOR U54246 ( .A(n53802), .B(n53803), .Z(n53676) );
  XNOR U54247 ( .A(n53804), .B(n53805), .Z(n53803) );
  NANDN U54248 ( .A(n53680), .B(n53682), .Z(n53720) );
  ANDN U54249 ( .B(B[80]), .A(n71), .Z(n53682) );
  XNOR U54250 ( .A(n53806), .B(n53807), .Z(n53680) );
  XNOR U54251 ( .A(n53808), .B(n53809), .Z(n53807) );
  NAND U54252 ( .A(n53684), .B(n53686), .Z(n53717) );
  ANDN U54253 ( .B(B[80]), .A(n70), .Z(n53686) );
  XNOR U54254 ( .A(n53810), .B(n53811), .Z(n53684) );
  XNOR U54255 ( .A(n53812), .B(n53813), .Z(n53811) );
  NANDN U54256 ( .A(n53688), .B(n53690), .Z(n53714) );
  ANDN U54257 ( .B(B[80]), .A(n69), .Z(n53690) );
  XNOR U54258 ( .A(n53814), .B(n53815), .Z(n53688) );
  XNOR U54259 ( .A(n53816), .B(n53817), .Z(n53815) );
  NAND U54260 ( .A(n53692), .B(n53694), .Z(n53711) );
  ANDN U54261 ( .B(B[80]), .A(n68), .Z(n53694) );
  XNOR U54262 ( .A(n53818), .B(n53819), .Z(n53692) );
  XNOR U54263 ( .A(n53820), .B(n53821), .Z(n53819) );
  NANDN U54264 ( .A(n53696), .B(n53698), .Z(n53708) );
  ANDN U54265 ( .B(B[80]), .A(n67), .Z(n53698) );
  XNOR U54266 ( .A(n53822), .B(n53823), .Z(n53696) );
  XNOR U54267 ( .A(n53824), .B(n53825), .Z(n53823) );
  NAND U54268 ( .A(n53700), .B(n53702), .Z(n53705) );
  ANDN U54269 ( .B(B[80]), .A(n66), .Z(n53702) );
  XNOR U54270 ( .A(n53826), .B(n53827), .Z(n53700) );
  XNOR U54271 ( .A(n53828), .B(n53829), .Z(n53827) );
  ANDN U54272 ( .B(B[80]), .A(n65), .Z(n51898) );
  XNOR U54273 ( .A(n51906), .B(n53830), .Z(n51899) );
  XNOR U54274 ( .A(n51905), .B(n51903), .Z(n53830) );
  AND U54275 ( .A(n53831), .B(n53832), .Z(n51903) );
  NANDN U54276 ( .A(n53829), .B(n53833), .Z(n53832) );
  NANDN U54277 ( .A(n53828), .B(n53826), .Z(n53833) );
  AND U54278 ( .A(n53834), .B(n53835), .Z(n53829) );
  NANDN U54279 ( .A(n53825), .B(n53836), .Z(n53835) );
  OR U54280 ( .A(n53824), .B(n53822), .Z(n53836) );
  AND U54281 ( .A(n53837), .B(n53838), .Z(n53825) );
  NANDN U54282 ( .A(n53821), .B(n53839), .Z(n53838) );
  NANDN U54283 ( .A(n53820), .B(n53818), .Z(n53839) );
  AND U54284 ( .A(n53840), .B(n53841), .Z(n53821) );
  NANDN U54285 ( .A(n53817), .B(n53842), .Z(n53841) );
  OR U54286 ( .A(n53816), .B(n53814), .Z(n53842) );
  AND U54287 ( .A(n53843), .B(n53844), .Z(n53817) );
  NANDN U54288 ( .A(n53813), .B(n53845), .Z(n53844) );
  NANDN U54289 ( .A(n53812), .B(n53810), .Z(n53845) );
  AND U54290 ( .A(n53846), .B(n53847), .Z(n53813) );
  NANDN U54291 ( .A(n53809), .B(n53848), .Z(n53847) );
  OR U54292 ( .A(n53808), .B(n53806), .Z(n53848) );
  AND U54293 ( .A(n53849), .B(n53850), .Z(n53809) );
  NANDN U54294 ( .A(n53805), .B(n53851), .Z(n53850) );
  NANDN U54295 ( .A(n53804), .B(n53802), .Z(n53851) );
  AND U54296 ( .A(n53852), .B(n53853), .Z(n53805) );
  NANDN U54297 ( .A(n53801), .B(n53854), .Z(n53853) );
  OR U54298 ( .A(n53800), .B(n53798), .Z(n53854) );
  AND U54299 ( .A(n53855), .B(n53856), .Z(n53801) );
  NANDN U54300 ( .A(n53797), .B(n53857), .Z(n53856) );
  NANDN U54301 ( .A(n53796), .B(n53794), .Z(n53857) );
  AND U54302 ( .A(n53858), .B(n53859), .Z(n53797) );
  NANDN U54303 ( .A(n53793), .B(n53860), .Z(n53859) );
  OR U54304 ( .A(n53792), .B(n53790), .Z(n53860) );
  AND U54305 ( .A(n53861), .B(n53862), .Z(n53793) );
  NANDN U54306 ( .A(n53789), .B(n53863), .Z(n53862) );
  NANDN U54307 ( .A(n53788), .B(n53786), .Z(n53863) );
  AND U54308 ( .A(n53864), .B(n53865), .Z(n53789) );
  NANDN U54309 ( .A(n53785), .B(n53866), .Z(n53865) );
  OR U54310 ( .A(n53784), .B(n53782), .Z(n53866) );
  AND U54311 ( .A(n53867), .B(n53868), .Z(n53785) );
  NANDN U54312 ( .A(n53781), .B(n53869), .Z(n53868) );
  NANDN U54313 ( .A(n53780), .B(n53778), .Z(n53869) );
  AND U54314 ( .A(n53870), .B(n53871), .Z(n53781) );
  NANDN U54315 ( .A(n53777), .B(n53872), .Z(n53871) );
  OR U54316 ( .A(n53776), .B(n53774), .Z(n53872) );
  AND U54317 ( .A(n53873), .B(n53874), .Z(n53777) );
  NANDN U54318 ( .A(n53773), .B(n53875), .Z(n53874) );
  NANDN U54319 ( .A(n53772), .B(n53770), .Z(n53875) );
  AND U54320 ( .A(n53876), .B(n53877), .Z(n53773) );
  NANDN U54321 ( .A(n53769), .B(n53878), .Z(n53877) );
  OR U54322 ( .A(n53768), .B(n53766), .Z(n53878) );
  AND U54323 ( .A(n53879), .B(n53880), .Z(n53769) );
  NANDN U54324 ( .A(n53764), .B(n53881), .Z(n53880) );
  NAND U54325 ( .A(n53762), .B(n53765), .Z(n53881) );
  NANDN U54326 ( .A(n53760), .B(n53882), .Z(n53764) );
  AND U54327 ( .A(A[0]), .B(B[82]), .Z(n53882) );
  NAND U54328 ( .A(B[81]), .B(A[1]), .Z(n53760) );
  XNOR U54329 ( .A(n53883), .B(n53884), .Z(n53762) );
  NAND U54330 ( .A(B[83]), .B(A[0]), .Z(n53884) );
  NAND U54331 ( .A(B[81]), .B(A[2]), .Z(n53765) );
  NAND U54332 ( .A(n53766), .B(n53768), .Z(n53876) );
  ANDN U54333 ( .B(B[81]), .A(n82), .Z(n53768) );
  XOR U54334 ( .A(n53885), .B(n53886), .Z(n53766) );
  XNOR U54335 ( .A(n53887), .B(n53888), .Z(n53886) );
  NANDN U54336 ( .A(n53770), .B(n53772), .Z(n53873) );
  ANDN U54337 ( .B(B[81]), .A(n81), .Z(n53772) );
  XNOR U54338 ( .A(n53889), .B(n53890), .Z(n53770) );
  XNOR U54339 ( .A(n53891), .B(n53892), .Z(n53890) );
  NAND U54340 ( .A(n53774), .B(n53776), .Z(n53870) );
  ANDN U54341 ( .B(B[81]), .A(n80), .Z(n53776) );
  XNOR U54342 ( .A(n53893), .B(n53894), .Z(n53774) );
  XNOR U54343 ( .A(n53895), .B(n53896), .Z(n53894) );
  NANDN U54344 ( .A(n53778), .B(n53780), .Z(n53867) );
  ANDN U54345 ( .B(B[81]), .A(n79), .Z(n53780) );
  XNOR U54346 ( .A(n53897), .B(n53898), .Z(n53778) );
  XNOR U54347 ( .A(n53899), .B(n53900), .Z(n53898) );
  NAND U54348 ( .A(n53782), .B(n53784), .Z(n53864) );
  ANDN U54349 ( .B(B[81]), .A(n78), .Z(n53784) );
  XNOR U54350 ( .A(n53901), .B(n53902), .Z(n53782) );
  XNOR U54351 ( .A(n53903), .B(n53904), .Z(n53902) );
  NANDN U54352 ( .A(n53786), .B(n53788), .Z(n53861) );
  ANDN U54353 ( .B(B[81]), .A(n77), .Z(n53788) );
  XNOR U54354 ( .A(n53905), .B(n53906), .Z(n53786) );
  XNOR U54355 ( .A(n53907), .B(n53908), .Z(n53906) );
  NAND U54356 ( .A(n53790), .B(n53792), .Z(n53858) );
  ANDN U54357 ( .B(B[81]), .A(n76), .Z(n53792) );
  XNOR U54358 ( .A(n53909), .B(n53910), .Z(n53790) );
  XNOR U54359 ( .A(n53911), .B(n53912), .Z(n53910) );
  NANDN U54360 ( .A(n53794), .B(n53796), .Z(n53855) );
  ANDN U54361 ( .B(B[81]), .A(n75), .Z(n53796) );
  XNOR U54362 ( .A(n53913), .B(n53914), .Z(n53794) );
  XNOR U54363 ( .A(n53915), .B(n53916), .Z(n53914) );
  NAND U54364 ( .A(n53798), .B(n53800), .Z(n53852) );
  ANDN U54365 ( .B(B[81]), .A(n74), .Z(n53800) );
  XNOR U54366 ( .A(n53917), .B(n53918), .Z(n53798) );
  XNOR U54367 ( .A(n53919), .B(n53920), .Z(n53918) );
  NANDN U54368 ( .A(n53802), .B(n53804), .Z(n53849) );
  ANDN U54369 ( .B(B[81]), .A(n73), .Z(n53804) );
  XNOR U54370 ( .A(n53921), .B(n53922), .Z(n53802) );
  XNOR U54371 ( .A(n53923), .B(n53924), .Z(n53922) );
  NAND U54372 ( .A(n53806), .B(n53808), .Z(n53846) );
  ANDN U54373 ( .B(B[81]), .A(n72), .Z(n53808) );
  XNOR U54374 ( .A(n53925), .B(n53926), .Z(n53806) );
  XNOR U54375 ( .A(n53927), .B(n53928), .Z(n53926) );
  NANDN U54376 ( .A(n53810), .B(n53812), .Z(n53843) );
  ANDN U54377 ( .B(B[81]), .A(n71), .Z(n53812) );
  XNOR U54378 ( .A(n53929), .B(n53930), .Z(n53810) );
  XNOR U54379 ( .A(n53931), .B(n53932), .Z(n53930) );
  NAND U54380 ( .A(n53814), .B(n53816), .Z(n53840) );
  ANDN U54381 ( .B(B[81]), .A(n70), .Z(n53816) );
  XNOR U54382 ( .A(n53933), .B(n53934), .Z(n53814) );
  XNOR U54383 ( .A(n53935), .B(n53936), .Z(n53934) );
  NANDN U54384 ( .A(n53818), .B(n53820), .Z(n53837) );
  ANDN U54385 ( .B(B[81]), .A(n69), .Z(n53820) );
  XNOR U54386 ( .A(n53937), .B(n53938), .Z(n53818) );
  XNOR U54387 ( .A(n53939), .B(n53940), .Z(n53938) );
  NAND U54388 ( .A(n53822), .B(n53824), .Z(n53834) );
  ANDN U54389 ( .B(B[81]), .A(n68), .Z(n53824) );
  XNOR U54390 ( .A(n53941), .B(n53942), .Z(n53822) );
  XNOR U54391 ( .A(n53943), .B(n53944), .Z(n53942) );
  NANDN U54392 ( .A(n53826), .B(n53828), .Z(n53831) );
  ANDN U54393 ( .B(B[81]), .A(n67), .Z(n53828) );
  XNOR U54394 ( .A(n53945), .B(n53946), .Z(n53826) );
  XNOR U54395 ( .A(n53947), .B(n53948), .Z(n53946) );
  ANDN U54396 ( .B(B[81]), .A(n66), .Z(n51905) );
  XNOR U54397 ( .A(n51913), .B(n53949), .Z(n51906) );
  XNOR U54398 ( .A(n51912), .B(n51910), .Z(n53949) );
  AND U54399 ( .A(n53950), .B(n53951), .Z(n51910) );
  NANDN U54400 ( .A(n53948), .B(n53952), .Z(n53951) );
  OR U54401 ( .A(n53947), .B(n53945), .Z(n53952) );
  AND U54402 ( .A(n53953), .B(n53954), .Z(n53948) );
  NANDN U54403 ( .A(n53944), .B(n53955), .Z(n53954) );
  NANDN U54404 ( .A(n53943), .B(n53941), .Z(n53955) );
  AND U54405 ( .A(n53956), .B(n53957), .Z(n53944) );
  NANDN U54406 ( .A(n53940), .B(n53958), .Z(n53957) );
  OR U54407 ( .A(n53939), .B(n53937), .Z(n53958) );
  AND U54408 ( .A(n53959), .B(n53960), .Z(n53940) );
  NANDN U54409 ( .A(n53936), .B(n53961), .Z(n53960) );
  NANDN U54410 ( .A(n53935), .B(n53933), .Z(n53961) );
  AND U54411 ( .A(n53962), .B(n53963), .Z(n53936) );
  NANDN U54412 ( .A(n53932), .B(n53964), .Z(n53963) );
  OR U54413 ( .A(n53931), .B(n53929), .Z(n53964) );
  AND U54414 ( .A(n53965), .B(n53966), .Z(n53932) );
  NANDN U54415 ( .A(n53928), .B(n53967), .Z(n53966) );
  NANDN U54416 ( .A(n53927), .B(n53925), .Z(n53967) );
  AND U54417 ( .A(n53968), .B(n53969), .Z(n53928) );
  NANDN U54418 ( .A(n53924), .B(n53970), .Z(n53969) );
  OR U54419 ( .A(n53923), .B(n53921), .Z(n53970) );
  AND U54420 ( .A(n53971), .B(n53972), .Z(n53924) );
  NANDN U54421 ( .A(n53920), .B(n53973), .Z(n53972) );
  NANDN U54422 ( .A(n53919), .B(n53917), .Z(n53973) );
  AND U54423 ( .A(n53974), .B(n53975), .Z(n53920) );
  NANDN U54424 ( .A(n53916), .B(n53976), .Z(n53975) );
  OR U54425 ( .A(n53915), .B(n53913), .Z(n53976) );
  AND U54426 ( .A(n53977), .B(n53978), .Z(n53916) );
  NANDN U54427 ( .A(n53912), .B(n53979), .Z(n53978) );
  NANDN U54428 ( .A(n53911), .B(n53909), .Z(n53979) );
  AND U54429 ( .A(n53980), .B(n53981), .Z(n53912) );
  NANDN U54430 ( .A(n53908), .B(n53982), .Z(n53981) );
  OR U54431 ( .A(n53907), .B(n53905), .Z(n53982) );
  AND U54432 ( .A(n53983), .B(n53984), .Z(n53908) );
  NANDN U54433 ( .A(n53904), .B(n53985), .Z(n53984) );
  NANDN U54434 ( .A(n53903), .B(n53901), .Z(n53985) );
  AND U54435 ( .A(n53986), .B(n53987), .Z(n53904) );
  NANDN U54436 ( .A(n53900), .B(n53988), .Z(n53987) );
  OR U54437 ( .A(n53899), .B(n53897), .Z(n53988) );
  AND U54438 ( .A(n53989), .B(n53990), .Z(n53900) );
  NANDN U54439 ( .A(n53896), .B(n53991), .Z(n53990) );
  NANDN U54440 ( .A(n53895), .B(n53893), .Z(n53991) );
  AND U54441 ( .A(n53992), .B(n53993), .Z(n53896) );
  NANDN U54442 ( .A(n53892), .B(n53994), .Z(n53993) );
  OR U54443 ( .A(n53891), .B(n53889), .Z(n53994) );
  AND U54444 ( .A(n53995), .B(n53996), .Z(n53892) );
  NANDN U54445 ( .A(n53887), .B(n53997), .Z(n53996) );
  NAND U54446 ( .A(n53885), .B(n53888), .Z(n53997) );
  NANDN U54447 ( .A(n53883), .B(n53998), .Z(n53887) );
  AND U54448 ( .A(A[0]), .B(B[83]), .Z(n53998) );
  NAND U54449 ( .A(B[82]), .B(A[1]), .Z(n53883) );
  XNOR U54450 ( .A(n53999), .B(n54000), .Z(n53885) );
  NAND U54451 ( .A(B[84]), .B(A[0]), .Z(n54000) );
  NAND U54452 ( .A(B[82]), .B(A[2]), .Z(n53888) );
  NAND U54453 ( .A(n53889), .B(n53891), .Z(n53992) );
  ANDN U54454 ( .B(B[82]), .A(n82), .Z(n53891) );
  XOR U54455 ( .A(n54001), .B(n54002), .Z(n53889) );
  XNOR U54456 ( .A(n54003), .B(n54004), .Z(n54002) );
  NANDN U54457 ( .A(n53893), .B(n53895), .Z(n53989) );
  ANDN U54458 ( .B(B[82]), .A(n81), .Z(n53895) );
  XNOR U54459 ( .A(n54005), .B(n54006), .Z(n53893) );
  XNOR U54460 ( .A(n54007), .B(n54008), .Z(n54006) );
  NAND U54461 ( .A(n53897), .B(n53899), .Z(n53986) );
  ANDN U54462 ( .B(B[82]), .A(n80), .Z(n53899) );
  XNOR U54463 ( .A(n54009), .B(n54010), .Z(n53897) );
  XNOR U54464 ( .A(n54011), .B(n54012), .Z(n54010) );
  NANDN U54465 ( .A(n53901), .B(n53903), .Z(n53983) );
  ANDN U54466 ( .B(B[82]), .A(n79), .Z(n53903) );
  XNOR U54467 ( .A(n54013), .B(n54014), .Z(n53901) );
  XNOR U54468 ( .A(n54015), .B(n54016), .Z(n54014) );
  NAND U54469 ( .A(n53905), .B(n53907), .Z(n53980) );
  ANDN U54470 ( .B(B[82]), .A(n78), .Z(n53907) );
  XNOR U54471 ( .A(n54017), .B(n54018), .Z(n53905) );
  XNOR U54472 ( .A(n54019), .B(n54020), .Z(n54018) );
  NANDN U54473 ( .A(n53909), .B(n53911), .Z(n53977) );
  ANDN U54474 ( .B(B[82]), .A(n77), .Z(n53911) );
  XNOR U54475 ( .A(n54021), .B(n54022), .Z(n53909) );
  XNOR U54476 ( .A(n54023), .B(n54024), .Z(n54022) );
  NAND U54477 ( .A(n53913), .B(n53915), .Z(n53974) );
  ANDN U54478 ( .B(B[82]), .A(n76), .Z(n53915) );
  XNOR U54479 ( .A(n54025), .B(n54026), .Z(n53913) );
  XNOR U54480 ( .A(n54027), .B(n54028), .Z(n54026) );
  NANDN U54481 ( .A(n53917), .B(n53919), .Z(n53971) );
  ANDN U54482 ( .B(B[82]), .A(n75), .Z(n53919) );
  XNOR U54483 ( .A(n54029), .B(n54030), .Z(n53917) );
  XNOR U54484 ( .A(n54031), .B(n54032), .Z(n54030) );
  NAND U54485 ( .A(n53921), .B(n53923), .Z(n53968) );
  ANDN U54486 ( .B(B[82]), .A(n74), .Z(n53923) );
  XNOR U54487 ( .A(n54033), .B(n54034), .Z(n53921) );
  XNOR U54488 ( .A(n54035), .B(n54036), .Z(n54034) );
  NANDN U54489 ( .A(n53925), .B(n53927), .Z(n53965) );
  ANDN U54490 ( .B(B[82]), .A(n73), .Z(n53927) );
  XNOR U54491 ( .A(n54037), .B(n54038), .Z(n53925) );
  XNOR U54492 ( .A(n54039), .B(n54040), .Z(n54038) );
  NAND U54493 ( .A(n53929), .B(n53931), .Z(n53962) );
  ANDN U54494 ( .B(B[82]), .A(n72), .Z(n53931) );
  XNOR U54495 ( .A(n54041), .B(n54042), .Z(n53929) );
  XNOR U54496 ( .A(n54043), .B(n54044), .Z(n54042) );
  NANDN U54497 ( .A(n53933), .B(n53935), .Z(n53959) );
  ANDN U54498 ( .B(B[82]), .A(n71), .Z(n53935) );
  XNOR U54499 ( .A(n54045), .B(n54046), .Z(n53933) );
  XNOR U54500 ( .A(n54047), .B(n54048), .Z(n54046) );
  NAND U54501 ( .A(n53937), .B(n53939), .Z(n53956) );
  ANDN U54502 ( .B(B[82]), .A(n70), .Z(n53939) );
  XNOR U54503 ( .A(n54049), .B(n54050), .Z(n53937) );
  XNOR U54504 ( .A(n54051), .B(n54052), .Z(n54050) );
  NANDN U54505 ( .A(n53941), .B(n53943), .Z(n53953) );
  ANDN U54506 ( .B(B[82]), .A(n69), .Z(n53943) );
  XNOR U54507 ( .A(n54053), .B(n54054), .Z(n53941) );
  XNOR U54508 ( .A(n54055), .B(n54056), .Z(n54054) );
  NAND U54509 ( .A(n53945), .B(n53947), .Z(n53950) );
  ANDN U54510 ( .B(B[82]), .A(n68), .Z(n53947) );
  XNOR U54511 ( .A(n54057), .B(n54058), .Z(n53945) );
  XNOR U54512 ( .A(n54059), .B(n54060), .Z(n54058) );
  ANDN U54513 ( .B(B[82]), .A(n67), .Z(n51912) );
  XNOR U54514 ( .A(n51920), .B(n54061), .Z(n51913) );
  XNOR U54515 ( .A(n51919), .B(n51917), .Z(n54061) );
  AND U54516 ( .A(n54062), .B(n54063), .Z(n51917) );
  NANDN U54517 ( .A(n54060), .B(n54064), .Z(n54063) );
  NANDN U54518 ( .A(n54059), .B(n54057), .Z(n54064) );
  AND U54519 ( .A(n54065), .B(n54066), .Z(n54060) );
  NANDN U54520 ( .A(n54056), .B(n54067), .Z(n54066) );
  OR U54521 ( .A(n54055), .B(n54053), .Z(n54067) );
  AND U54522 ( .A(n54068), .B(n54069), .Z(n54056) );
  NANDN U54523 ( .A(n54052), .B(n54070), .Z(n54069) );
  NANDN U54524 ( .A(n54051), .B(n54049), .Z(n54070) );
  AND U54525 ( .A(n54071), .B(n54072), .Z(n54052) );
  NANDN U54526 ( .A(n54048), .B(n54073), .Z(n54072) );
  OR U54527 ( .A(n54047), .B(n54045), .Z(n54073) );
  AND U54528 ( .A(n54074), .B(n54075), .Z(n54048) );
  NANDN U54529 ( .A(n54044), .B(n54076), .Z(n54075) );
  NANDN U54530 ( .A(n54043), .B(n54041), .Z(n54076) );
  AND U54531 ( .A(n54077), .B(n54078), .Z(n54044) );
  NANDN U54532 ( .A(n54040), .B(n54079), .Z(n54078) );
  OR U54533 ( .A(n54039), .B(n54037), .Z(n54079) );
  AND U54534 ( .A(n54080), .B(n54081), .Z(n54040) );
  NANDN U54535 ( .A(n54036), .B(n54082), .Z(n54081) );
  NANDN U54536 ( .A(n54035), .B(n54033), .Z(n54082) );
  AND U54537 ( .A(n54083), .B(n54084), .Z(n54036) );
  NANDN U54538 ( .A(n54032), .B(n54085), .Z(n54084) );
  OR U54539 ( .A(n54031), .B(n54029), .Z(n54085) );
  AND U54540 ( .A(n54086), .B(n54087), .Z(n54032) );
  NANDN U54541 ( .A(n54028), .B(n54088), .Z(n54087) );
  NANDN U54542 ( .A(n54027), .B(n54025), .Z(n54088) );
  AND U54543 ( .A(n54089), .B(n54090), .Z(n54028) );
  NANDN U54544 ( .A(n54024), .B(n54091), .Z(n54090) );
  OR U54545 ( .A(n54023), .B(n54021), .Z(n54091) );
  AND U54546 ( .A(n54092), .B(n54093), .Z(n54024) );
  NANDN U54547 ( .A(n54020), .B(n54094), .Z(n54093) );
  NANDN U54548 ( .A(n54019), .B(n54017), .Z(n54094) );
  AND U54549 ( .A(n54095), .B(n54096), .Z(n54020) );
  NANDN U54550 ( .A(n54016), .B(n54097), .Z(n54096) );
  OR U54551 ( .A(n54015), .B(n54013), .Z(n54097) );
  AND U54552 ( .A(n54098), .B(n54099), .Z(n54016) );
  NANDN U54553 ( .A(n54012), .B(n54100), .Z(n54099) );
  NANDN U54554 ( .A(n54011), .B(n54009), .Z(n54100) );
  AND U54555 ( .A(n54101), .B(n54102), .Z(n54012) );
  NANDN U54556 ( .A(n54008), .B(n54103), .Z(n54102) );
  OR U54557 ( .A(n54007), .B(n54005), .Z(n54103) );
  AND U54558 ( .A(n54104), .B(n54105), .Z(n54008) );
  NANDN U54559 ( .A(n54003), .B(n54106), .Z(n54105) );
  NAND U54560 ( .A(n54001), .B(n54004), .Z(n54106) );
  NANDN U54561 ( .A(n53999), .B(n54107), .Z(n54003) );
  AND U54562 ( .A(A[0]), .B(B[84]), .Z(n54107) );
  NAND U54563 ( .A(B[83]), .B(A[1]), .Z(n53999) );
  XNOR U54564 ( .A(n54108), .B(n54109), .Z(n54001) );
  NAND U54565 ( .A(B[85]), .B(A[0]), .Z(n54109) );
  NAND U54566 ( .A(B[83]), .B(A[2]), .Z(n54004) );
  NAND U54567 ( .A(n54005), .B(n54007), .Z(n54101) );
  ANDN U54568 ( .B(B[83]), .A(n82), .Z(n54007) );
  XOR U54569 ( .A(n54110), .B(n54111), .Z(n54005) );
  XNOR U54570 ( .A(n54112), .B(n54113), .Z(n54111) );
  NANDN U54571 ( .A(n54009), .B(n54011), .Z(n54098) );
  ANDN U54572 ( .B(B[83]), .A(n81), .Z(n54011) );
  XNOR U54573 ( .A(n54114), .B(n54115), .Z(n54009) );
  XNOR U54574 ( .A(n54116), .B(n54117), .Z(n54115) );
  NAND U54575 ( .A(n54013), .B(n54015), .Z(n54095) );
  ANDN U54576 ( .B(B[83]), .A(n80), .Z(n54015) );
  XNOR U54577 ( .A(n54118), .B(n54119), .Z(n54013) );
  XNOR U54578 ( .A(n54120), .B(n54121), .Z(n54119) );
  NANDN U54579 ( .A(n54017), .B(n54019), .Z(n54092) );
  ANDN U54580 ( .B(B[83]), .A(n79), .Z(n54019) );
  XNOR U54581 ( .A(n54122), .B(n54123), .Z(n54017) );
  XNOR U54582 ( .A(n54124), .B(n54125), .Z(n54123) );
  NAND U54583 ( .A(n54021), .B(n54023), .Z(n54089) );
  ANDN U54584 ( .B(B[83]), .A(n78), .Z(n54023) );
  XNOR U54585 ( .A(n54126), .B(n54127), .Z(n54021) );
  XNOR U54586 ( .A(n54128), .B(n54129), .Z(n54127) );
  NANDN U54587 ( .A(n54025), .B(n54027), .Z(n54086) );
  ANDN U54588 ( .B(B[83]), .A(n77), .Z(n54027) );
  XNOR U54589 ( .A(n54130), .B(n54131), .Z(n54025) );
  XNOR U54590 ( .A(n54132), .B(n54133), .Z(n54131) );
  NAND U54591 ( .A(n54029), .B(n54031), .Z(n54083) );
  ANDN U54592 ( .B(B[83]), .A(n76), .Z(n54031) );
  XNOR U54593 ( .A(n54134), .B(n54135), .Z(n54029) );
  XNOR U54594 ( .A(n54136), .B(n54137), .Z(n54135) );
  NANDN U54595 ( .A(n54033), .B(n54035), .Z(n54080) );
  ANDN U54596 ( .B(B[83]), .A(n75), .Z(n54035) );
  XNOR U54597 ( .A(n54138), .B(n54139), .Z(n54033) );
  XNOR U54598 ( .A(n54140), .B(n54141), .Z(n54139) );
  NAND U54599 ( .A(n54037), .B(n54039), .Z(n54077) );
  ANDN U54600 ( .B(B[83]), .A(n74), .Z(n54039) );
  XNOR U54601 ( .A(n54142), .B(n54143), .Z(n54037) );
  XNOR U54602 ( .A(n54144), .B(n54145), .Z(n54143) );
  NANDN U54603 ( .A(n54041), .B(n54043), .Z(n54074) );
  ANDN U54604 ( .B(B[83]), .A(n73), .Z(n54043) );
  XNOR U54605 ( .A(n54146), .B(n54147), .Z(n54041) );
  XNOR U54606 ( .A(n54148), .B(n54149), .Z(n54147) );
  NAND U54607 ( .A(n54045), .B(n54047), .Z(n54071) );
  ANDN U54608 ( .B(B[83]), .A(n72), .Z(n54047) );
  XNOR U54609 ( .A(n54150), .B(n54151), .Z(n54045) );
  XNOR U54610 ( .A(n54152), .B(n54153), .Z(n54151) );
  NANDN U54611 ( .A(n54049), .B(n54051), .Z(n54068) );
  ANDN U54612 ( .B(B[83]), .A(n71), .Z(n54051) );
  XNOR U54613 ( .A(n54154), .B(n54155), .Z(n54049) );
  XNOR U54614 ( .A(n54156), .B(n54157), .Z(n54155) );
  NAND U54615 ( .A(n54053), .B(n54055), .Z(n54065) );
  ANDN U54616 ( .B(B[83]), .A(n70), .Z(n54055) );
  XNOR U54617 ( .A(n54158), .B(n54159), .Z(n54053) );
  XNOR U54618 ( .A(n54160), .B(n54161), .Z(n54159) );
  NANDN U54619 ( .A(n54057), .B(n54059), .Z(n54062) );
  ANDN U54620 ( .B(B[83]), .A(n69), .Z(n54059) );
  XNOR U54621 ( .A(n54162), .B(n54163), .Z(n54057) );
  XNOR U54622 ( .A(n54164), .B(n54165), .Z(n54163) );
  ANDN U54623 ( .B(B[83]), .A(n68), .Z(n51919) );
  XNOR U54624 ( .A(n51927), .B(n54166), .Z(n51920) );
  XNOR U54625 ( .A(n51926), .B(n51924), .Z(n54166) );
  AND U54626 ( .A(n54167), .B(n54168), .Z(n51924) );
  NANDN U54627 ( .A(n54165), .B(n54169), .Z(n54168) );
  OR U54628 ( .A(n54164), .B(n54162), .Z(n54169) );
  AND U54629 ( .A(n54170), .B(n54171), .Z(n54165) );
  NANDN U54630 ( .A(n54161), .B(n54172), .Z(n54171) );
  NANDN U54631 ( .A(n54160), .B(n54158), .Z(n54172) );
  AND U54632 ( .A(n54173), .B(n54174), .Z(n54161) );
  NANDN U54633 ( .A(n54157), .B(n54175), .Z(n54174) );
  OR U54634 ( .A(n54156), .B(n54154), .Z(n54175) );
  AND U54635 ( .A(n54176), .B(n54177), .Z(n54157) );
  NANDN U54636 ( .A(n54153), .B(n54178), .Z(n54177) );
  NANDN U54637 ( .A(n54152), .B(n54150), .Z(n54178) );
  AND U54638 ( .A(n54179), .B(n54180), .Z(n54153) );
  NANDN U54639 ( .A(n54149), .B(n54181), .Z(n54180) );
  OR U54640 ( .A(n54148), .B(n54146), .Z(n54181) );
  AND U54641 ( .A(n54182), .B(n54183), .Z(n54149) );
  NANDN U54642 ( .A(n54145), .B(n54184), .Z(n54183) );
  NANDN U54643 ( .A(n54144), .B(n54142), .Z(n54184) );
  AND U54644 ( .A(n54185), .B(n54186), .Z(n54145) );
  NANDN U54645 ( .A(n54141), .B(n54187), .Z(n54186) );
  OR U54646 ( .A(n54140), .B(n54138), .Z(n54187) );
  AND U54647 ( .A(n54188), .B(n54189), .Z(n54141) );
  NANDN U54648 ( .A(n54137), .B(n54190), .Z(n54189) );
  NANDN U54649 ( .A(n54136), .B(n54134), .Z(n54190) );
  AND U54650 ( .A(n54191), .B(n54192), .Z(n54137) );
  NANDN U54651 ( .A(n54133), .B(n54193), .Z(n54192) );
  OR U54652 ( .A(n54132), .B(n54130), .Z(n54193) );
  AND U54653 ( .A(n54194), .B(n54195), .Z(n54133) );
  NANDN U54654 ( .A(n54129), .B(n54196), .Z(n54195) );
  NANDN U54655 ( .A(n54128), .B(n54126), .Z(n54196) );
  AND U54656 ( .A(n54197), .B(n54198), .Z(n54129) );
  NANDN U54657 ( .A(n54125), .B(n54199), .Z(n54198) );
  OR U54658 ( .A(n54124), .B(n54122), .Z(n54199) );
  AND U54659 ( .A(n54200), .B(n54201), .Z(n54125) );
  NANDN U54660 ( .A(n54121), .B(n54202), .Z(n54201) );
  NANDN U54661 ( .A(n54120), .B(n54118), .Z(n54202) );
  AND U54662 ( .A(n54203), .B(n54204), .Z(n54121) );
  NANDN U54663 ( .A(n54117), .B(n54205), .Z(n54204) );
  OR U54664 ( .A(n54116), .B(n54114), .Z(n54205) );
  AND U54665 ( .A(n54206), .B(n54207), .Z(n54117) );
  NANDN U54666 ( .A(n54112), .B(n54208), .Z(n54207) );
  NAND U54667 ( .A(n54110), .B(n54113), .Z(n54208) );
  NANDN U54668 ( .A(n54108), .B(n54209), .Z(n54112) );
  AND U54669 ( .A(A[0]), .B(B[85]), .Z(n54209) );
  NAND U54670 ( .A(B[84]), .B(A[1]), .Z(n54108) );
  XNOR U54671 ( .A(n54210), .B(n54211), .Z(n54110) );
  NAND U54672 ( .A(B[86]), .B(A[0]), .Z(n54211) );
  NAND U54673 ( .A(B[84]), .B(A[2]), .Z(n54113) );
  NAND U54674 ( .A(n54114), .B(n54116), .Z(n54203) );
  ANDN U54675 ( .B(B[84]), .A(n82), .Z(n54116) );
  XOR U54676 ( .A(n54212), .B(n54213), .Z(n54114) );
  XNOR U54677 ( .A(n54214), .B(n54215), .Z(n54213) );
  NANDN U54678 ( .A(n54118), .B(n54120), .Z(n54200) );
  ANDN U54679 ( .B(B[84]), .A(n81), .Z(n54120) );
  XNOR U54680 ( .A(n54216), .B(n54217), .Z(n54118) );
  XNOR U54681 ( .A(n54218), .B(n54219), .Z(n54217) );
  NAND U54682 ( .A(n54122), .B(n54124), .Z(n54197) );
  ANDN U54683 ( .B(B[84]), .A(n80), .Z(n54124) );
  XNOR U54684 ( .A(n54220), .B(n54221), .Z(n54122) );
  XNOR U54685 ( .A(n54222), .B(n54223), .Z(n54221) );
  NANDN U54686 ( .A(n54126), .B(n54128), .Z(n54194) );
  ANDN U54687 ( .B(B[84]), .A(n79), .Z(n54128) );
  XNOR U54688 ( .A(n54224), .B(n54225), .Z(n54126) );
  XNOR U54689 ( .A(n54226), .B(n54227), .Z(n54225) );
  NAND U54690 ( .A(n54130), .B(n54132), .Z(n54191) );
  ANDN U54691 ( .B(B[84]), .A(n78), .Z(n54132) );
  XNOR U54692 ( .A(n54228), .B(n54229), .Z(n54130) );
  XNOR U54693 ( .A(n54230), .B(n54231), .Z(n54229) );
  NANDN U54694 ( .A(n54134), .B(n54136), .Z(n54188) );
  ANDN U54695 ( .B(B[84]), .A(n77), .Z(n54136) );
  XNOR U54696 ( .A(n54232), .B(n54233), .Z(n54134) );
  XNOR U54697 ( .A(n54234), .B(n54235), .Z(n54233) );
  NAND U54698 ( .A(n54138), .B(n54140), .Z(n54185) );
  ANDN U54699 ( .B(B[84]), .A(n76), .Z(n54140) );
  XNOR U54700 ( .A(n54236), .B(n54237), .Z(n54138) );
  XNOR U54701 ( .A(n54238), .B(n54239), .Z(n54237) );
  NANDN U54702 ( .A(n54142), .B(n54144), .Z(n54182) );
  ANDN U54703 ( .B(B[84]), .A(n75), .Z(n54144) );
  XNOR U54704 ( .A(n54240), .B(n54241), .Z(n54142) );
  XNOR U54705 ( .A(n54242), .B(n54243), .Z(n54241) );
  NAND U54706 ( .A(n54146), .B(n54148), .Z(n54179) );
  ANDN U54707 ( .B(B[84]), .A(n74), .Z(n54148) );
  XNOR U54708 ( .A(n54244), .B(n54245), .Z(n54146) );
  XNOR U54709 ( .A(n54246), .B(n54247), .Z(n54245) );
  NANDN U54710 ( .A(n54150), .B(n54152), .Z(n54176) );
  ANDN U54711 ( .B(B[84]), .A(n73), .Z(n54152) );
  XNOR U54712 ( .A(n54248), .B(n54249), .Z(n54150) );
  XNOR U54713 ( .A(n54250), .B(n54251), .Z(n54249) );
  NAND U54714 ( .A(n54154), .B(n54156), .Z(n54173) );
  ANDN U54715 ( .B(B[84]), .A(n72), .Z(n54156) );
  XNOR U54716 ( .A(n54252), .B(n54253), .Z(n54154) );
  XNOR U54717 ( .A(n54254), .B(n54255), .Z(n54253) );
  NANDN U54718 ( .A(n54158), .B(n54160), .Z(n54170) );
  ANDN U54719 ( .B(B[84]), .A(n71), .Z(n54160) );
  XNOR U54720 ( .A(n54256), .B(n54257), .Z(n54158) );
  XNOR U54721 ( .A(n54258), .B(n54259), .Z(n54257) );
  NAND U54722 ( .A(n54162), .B(n54164), .Z(n54167) );
  ANDN U54723 ( .B(B[84]), .A(n70), .Z(n54164) );
  XNOR U54724 ( .A(n54260), .B(n54261), .Z(n54162) );
  XNOR U54725 ( .A(n54262), .B(n54263), .Z(n54261) );
  ANDN U54726 ( .B(B[84]), .A(n69), .Z(n51926) );
  XNOR U54727 ( .A(n51934), .B(n54264), .Z(n51927) );
  XNOR U54728 ( .A(n51933), .B(n51931), .Z(n54264) );
  AND U54729 ( .A(n54265), .B(n54266), .Z(n51931) );
  NANDN U54730 ( .A(n54263), .B(n54267), .Z(n54266) );
  NANDN U54731 ( .A(n54262), .B(n54260), .Z(n54267) );
  AND U54732 ( .A(n54268), .B(n54269), .Z(n54263) );
  NANDN U54733 ( .A(n54259), .B(n54270), .Z(n54269) );
  OR U54734 ( .A(n54258), .B(n54256), .Z(n54270) );
  AND U54735 ( .A(n54271), .B(n54272), .Z(n54259) );
  NANDN U54736 ( .A(n54255), .B(n54273), .Z(n54272) );
  NANDN U54737 ( .A(n54254), .B(n54252), .Z(n54273) );
  AND U54738 ( .A(n54274), .B(n54275), .Z(n54255) );
  NANDN U54739 ( .A(n54251), .B(n54276), .Z(n54275) );
  OR U54740 ( .A(n54250), .B(n54248), .Z(n54276) );
  AND U54741 ( .A(n54277), .B(n54278), .Z(n54251) );
  NANDN U54742 ( .A(n54247), .B(n54279), .Z(n54278) );
  NANDN U54743 ( .A(n54246), .B(n54244), .Z(n54279) );
  AND U54744 ( .A(n54280), .B(n54281), .Z(n54247) );
  NANDN U54745 ( .A(n54243), .B(n54282), .Z(n54281) );
  OR U54746 ( .A(n54242), .B(n54240), .Z(n54282) );
  AND U54747 ( .A(n54283), .B(n54284), .Z(n54243) );
  NANDN U54748 ( .A(n54239), .B(n54285), .Z(n54284) );
  NANDN U54749 ( .A(n54238), .B(n54236), .Z(n54285) );
  AND U54750 ( .A(n54286), .B(n54287), .Z(n54239) );
  NANDN U54751 ( .A(n54235), .B(n54288), .Z(n54287) );
  OR U54752 ( .A(n54234), .B(n54232), .Z(n54288) );
  AND U54753 ( .A(n54289), .B(n54290), .Z(n54235) );
  NANDN U54754 ( .A(n54231), .B(n54291), .Z(n54290) );
  NANDN U54755 ( .A(n54230), .B(n54228), .Z(n54291) );
  AND U54756 ( .A(n54292), .B(n54293), .Z(n54231) );
  NANDN U54757 ( .A(n54227), .B(n54294), .Z(n54293) );
  OR U54758 ( .A(n54226), .B(n54224), .Z(n54294) );
  AND U54759 ( .A(n54295), .B(n54296), .Z(n54227) );
  NANDN U54760 ( .A(n54223), .B(n54297), .Z(n54296) );
  NANDN U54761 ( .A(n54222), .B(n54220), .Z(n54297) );
  AND U54762 ( .A(n54298), .B(n54299), .Z(n54223) );
  NANDN U54763 ( .A(n54219), .B(n54300), .Z(n54299) );
  OR U54764 ( .A(n54218), .B(n54216), .Z(n54300) );
  AND U54765 ( .A(n54301), .B(n54302), .Z(n54219) );
  NANDN U54766 ( .A(n54214), .B(n54303), .Z(n54302) );
  NAND U54767 ( .A(n54212), .B(n54215), .Z(n54303) );
  NANDN U54768 ( .A(n54210), .B(n54304), .Z(n54214) );
  AND U54769 ( .A(A[0]), .B(B[86]), .Z(n54304) );
  NAND U54770 ( .A(B[85]), .B(A[1]), .Z(n54210) );
  XNOR U54771 ( .A(n54305), .B(n54306), .Z(n54212) );
  NAND U54772 ( .A(B[87]), .B(A[0]), .Z(n54306) );
  NAND U54773 ( .A(B[85]), .B(A[2]), .Z(n54215) );
  NAND U54774 ( .A(n54216), .B(n54218), .Z(n54298) );
  ANDN U54775 ( .B(A[3]), .A(n33), .Z(n54218) );
  XOR U54776 ( .A(n54307), .B(n54308), .Z(n54216) );
  XNOR U54777 ( .A(n54309), .B(n54310), .Z(n54308) );
  NANDN U54778 ( .A(n54220), .B(n54222), .Z(n54295) );
  ANDN U54779 ( .B(A[4]), .A(n33), .Z(n54222) );
  XNOR U54780 ( .A(n54311), .B(n54312), .Z(n54220) );
  XNOR U54781 ( .A(n54313), .B(n54314), .Z(n54312) );
  NAND U54782 ( .A(n54224), .B(n54226), .Z(n54292) );
  ANDN U54783 ( .B(A[5]), .A(n33), .Z(n54226) );
  XNOR U54784 ( .A(n54315), .B(n54316), .Z(n54224) );
  XNOR U54785 ( .A(n54317), .B(n54318), .Z(n54316) );
  NANDN U54786 ( .A(n54228), .B(n54230), .Z(n54289) );
  ANDN U54787 ( .B(A[6]), .A(n33), .Z(n54230) );
  XNOR U54788 ( .A(n54319), .B(n54320), .Z(n54228) );
  XNOR U54789 ( .A(n54321), .B(n54322), .Z(n54320) );
  NAND U54790 ( .A(n54232), .B(n54234), .Z(n54286) );
  ANDN U54791 ( .B(A[7]), .A(n33), .Z(n54234) );
  XNOR U54792 ( .A(n54323), .B(n54324), .Z(n54232) );
  XNOR U54793 ( .A(n54325), .B(n54326), .Z(n54324) );
  NANDN U54794 ( .A(n54236), .B(n54238), .Z(n54283) );
  ANDN U54795 ( .B(A[8]), .A(n33), .Z(n54238) );
  XNOR U54796 ( .A(n54327), .B(n54328), .Z(n54236) );
  XNOR U54797 ( .A(n54329), .B(n54330), .Z(n54328) );
  NAND U54798 ( .A(n54240), .B(n54242), .Z(n54280) );
  ANDN U54799 ( .B(A[9]), .A(n33), .Z(n54242) );
  XNOR U54800 ( .A(n54331), .B(n54332), .Z(n54240) );
  XNOR U54801 ( .A(n54333), .B(n54334), .Z(n54332) );
  NANDN U54802 ( .A(n54244), .B(n54246), .Z(n54277) );
  ANDN U54803 ( .B(A[10]), .A(n33), .Z(n54246) );
  XNOR U54804 ( .A(n54335), .B(n54336), .Z(n54244) );
  XNOR U54805 ( .A(n54337), .B(n54338), .Z(n54336) );
  NAND U54806 ( .A(n54248), .B(n54250), .Z(n54274) );
  ANDN U54807 ( .B(A[11]), .A(n33), .Z(n54250) );
  XNOR U54808 ( .A(n54339), .B(n54340), .Z(n54248) );
  XNOR U54809 ( .A(n54341), .B(n54342), .Z(n54340) );
  NANDN U54810 ( .A(n54252), .B(n54254), .Z(n54271) );
  ANDN U54811 ( .B(A[12]), .A(n33), .Z(n54254) );
  XNOR U54812 ( .A(n54343), .B(n54344), .Z(n54252) );
  XNOR U54813 ( .A(n54345), .B(n54346), .Z(n54344) );
  NAND U54814 ( .A(n54256), .B(n54258), .Z(n54268) );
  ANDN U54815 ( .B(A[13]), .A(n33), .Z(n54258) );
  XNOR U54816 ( .A(n54347), .B(n54348), .Z(n54256) );
  XNOR U54817 ( .A(n54349), .B(n54350), .Z(n54348) );
  NANDN U54818 ( .A(n54260), .B(n54262), .Z(n54265) );
  ANDN U54819 ( .B(A[14]), .A(n33), .Z(n54262) );
  XNOR U54820 ( .A(n54351), .B(n54352), .Z(n54260) );
  XNOR U54821 ( .A(n54353), .B(n54354), .Z(n54352) );
  ANDN U54822 ( .B(A[15]), .A(n33), .Z(n51933) );
  XNOR U54823 ( .A(n51941), .B(n54355), .Z(n51934) );
  XNOR U54824 ( .A(n51940), .B(n51938), .Z(n54355) );
  AND U54825 ( .A(n54356), .B(n54357), .Z(n51938) );
  NANDN U54826 ( .A(n54354), .B(n54358), .Z(n54357) );
  OR U54827 ( .A(n54353), .B(n54351), .Z(n54358) );
  AND U54828 ( .A(n54359), .B(n54360), .Z(n54354) );
  NANDN U54829 ( .A(n54350), .B(n54361), .Z(n54360) );
  NANDN U54830 ( .A(n54349), .B(n54347), .Z(n54361) );
  AND U54831 ( .A(n54362), .B(n54363), .Z(n54350) );
  NANDN U54832 ( .A(n54346), .B(n54364), .Z(n54363) );
  OR U54833 ( .A(n54345), .B(n54343), .Z(n54364) );
  AND U54834 ( .A(n54365), .B(n54366), .Z(n54346) );
  NANDN U54835 ( .A(n54342), .B(n54367), .Z(n54366) );
  NANDN U54836 ( .A(n54341), .B(n54339), .Z(n54367) );
  AND U54837 ( .A(n54368), .B(n54369), .Z(n54342) );
  NANDN U54838 ( .A(n54338), .B(n54370), .Z(n54369) );
  OR U54839 ( .A(n54337), .B(n54335), .Z(n54370) );
  AND U54840 ( .A(n54371), .B(n54372), .Z(n54338) );
  NANDN U54841 ( .A(n54334), .B(n54373), .Z(n54372) );
  NANDN U54842 ( .A(n54333), .B(n54331), .Z(n54373) );
  AND U54843 ( .A(n54374), .B(n54375), .Z(n54334) );
  NANDN U54844 ( .A(n54330), .B(n54376), .Z(n54375) );
  OR U54845 ( .A(n54329), .B(n54327), .Z(n54376) );
  AND U54846 ( .A(n54377), .B(n54378), .Z(n54330) );
  NANDN U54847 ( .A(n54326), .B(n54379), .Z(n54378) );
  NANDN U54848 ( .A(n54325), .B(n54323), .Z(n54379) );
  AND U54849 ( .A(n54380), .B(n54381), .Z(n54326) );
  NANDN U54850 ( .A(n54322), .B(n54382), .Z(n54381) );
  OR U54851 ( .A(n54321), .B(n54319), .Z(n54382) );
  AND U54852 ( .A(n54383), .B(n54384), .Z(n54322) );
  NANDN U54853 ( .A(n54318), .B(n54385), .Z(n54384) );
  NANDN U54854 ( .A(n54317), .B(n54315), .Z(n54385) );
  AND U54855 ( .A(n54386), .B(n54387), .Z(n54318) );
  NANDN U54856 ( .A(n54314), .B(n54388), .Z(n54387) );
  OR U54857 ( .A(n54313), .B(n54311), .Z(n54388) );
  AND U54858 ( .A(n54389), .B(n54390), .Z(n54314) );
  NANDN U54859 ( .A(n54309), .B(n54391), .Z(n54390) );
  NAND U54860 ( .A(n54307), .B(n54310), .Z(n54391) );
  NANDN U54861 ( .A(n54305), .B(n54392), .Z(n54309) );
  AND U54862 ( .A(A[0]), .B(B[87]), .Z(n54392) );
  NAND U54863 ( .A(B[86]), .B(A[1]), .Z(n54305) );
  XNOR U54864 ( .A(n54393), .B(n54394), .Z(n54307) );
  NAND U54865 ( .A(B[88]), .B(A[0]), .Z(n54394) );
  NAND U54866 ( .A(B[86]), .B(A[2]), .Z(n54310) );
  NAND U54867 ( .A(n54311), .B(n54313), .Z(n54386) );
  ANDN U54868 ( .B(A[3]), .A(n31), .Z(n54313) );
  XOR U54869 ( .A(n54395), .B(n54396), .Z(n54311) );
  XNOR U54870 ( .A(n54397), .B(n54398), .Z(n54396) );
  NANDN U54871 ( .A(n54315), .B(n54317), .Z(n54383) );
  ANDN U54872 ( .B(A[4]), .A(n31), .Z(n54317) );
  XNOR U54873 ( .A(n54399), .B(n54400), .Z(n54315) );
  XNOR U54874 ( .A(n54401), .B(n54402), .Z(n54400) );
  NAND U54875 ( .A(n54319), .B(n54321), .Z(n54380) );
  ANDN U54876 ( .B(A[5]), .A(n31), .Z(n54321) );
  XNOR U54877 ( .A(n54403), .B(n54404), .Z(n54319) );
  XNOR U54878 ( .A(n54405), .B(n54406), .Z(n54404) );
  NANDN U54879 ( .A(n54323), .B(n54325), .Z(n54377) );
  ANDN U54880 ( .B(A[6]), .A(n31), .Z(n54325) );
  XNOR U54881 ( .A(n54407), .B(n54408), .Z(n54323) );
  XNOR U54882 ( .A(n54409), .B(n54410), .Z(n54408) );
  NAND U54883 ( .A(n54327), .B(n54329), .Z(n54374) );
  ANDN U54884 ( .B(A[7]), .A(n31), .Z(n54329) );
  XNOR U54885 ( .A(n54411), .B(n54412), .Z(n54327) );
  XNOR U54886 ( .A(n54413), .B(n54414), .Z(n54412) );
  NANDN U54887 ( .A(n54331), .B(n54333), .Z(n54371) );
  ANDN U54888 ( .B(A[8]), .A(n31), .Z(n54333) );
  XNOR U54889 ( .A(n54415), .B(n54416), .Z(n54331) );
  XNOR U54890 ( .A(n54417), .B(n54418), .Z(n54416) );
  NAND U54891 ( .A(n54335), .B(n54337), .Z(n54368) );
  ANDN U54892 ( .B(A[9]), .A(n31), .Z(n54337) );
  XNOR U54893 ( .A(n54419), .B(n54420), .Z(n54335) );
  XNOR U54894 ( .A(n54421), .B(n54422), .Z(n54420) );
  NANDN U54895 ( .A(n54339), .B(n54341), .Z(n54365) );
  ANDN U54896 ( .B(A[10]), .A(n31), .Z(n54341) );
  XNOR U54897 ( .A(n54423), .B(n54424), .Z(n54339) );
  XNOR U54898 ( .A(n54425), .B(n54426), .Z(n54424) );
  NAND U54899 ( .A(n54343), .B(n54345), .Z(n54362) );
  ANDN U54900 ( .B(A[11]), .A(n31), .Z(n54345) );
  XNOR U54901 ( .A(n54427), .B(n54428), .Z(n54343) );
  XNOR U54902 ( .A(n54429), .B(n54430), .Z(n54428) );
  NANDN U54903 ( .A(n54347), .B(n54349), .Z(n54359) );
  ANDN U54904 ( .B(A[12]), .A(n31), .Z(n54349) );
  XNOR U54905 ( .A(n54431), .B(n54432), .Z(n54347) );
  XNOR U54906 ( .A(n54433), .B(n54434), .Z(n54432) );
  NAND U54907 ( .A(n54351), .B(n54353), .Z(n54356) );
  ANDN U54908 ( .B(A[13]), .A(n31), .Z(n54353) );
  XNOR U54909 ( .A(n54435), .B(n54436), .Z(n54351) );
  XNOR U54910 ( .A(n54437), .B(n54438), .Z(n54436) );
  ANDN U54911 ( .B(A[14]), .A(n31), .Z(n51940) );
  XNOR U54912 ( .A(n51948), .B(n54439), .Z(n51941) );
  XNOR U54913 ( .A(n51947), .B(n51945), .Z(n54439) );
  AND U54914 ( .A(n54440), .B(n54441), .Z(n51945) );
  NANDN U54915 ( .A(n54438), .B(n54442), .Z(n54441) );
  NANDN U54916 ( .A(n54437), .B(n54435), .Z(n54442) );
  AND U54917 ( .A(n54443), .B(n54444), .Z(n54438) );
  NANDN U54918 ( .A(n54434), .B(n54445), .Z(n54444) );
  OR U54919 ( .A(n54433), .B(n54431), .Z(n54445) );
  AND U54920 ( .A(n54446), .B(n54447), .Z(n54434) );
  NANDN U54921 ( .A(n54430), .B(n54448), .Z(n54447) );
  NANDN U54922 ( .A(n54429), .B(n54427), .Z(n54448) );
  AND U54923 ( .A(n54449), .B(n54450), .Z(n54430) );
  NANDN U54924 ( .A(n54426), .B(n54451), .Z(n54450) );
  OR U54925 ( .A(n54425), .B(n54423), .Z(n54451) );
  AND U54926 ( .A(n54452), .B(n54453), .Z(n54426) );
  NANDN U54927 ( .A(n54422), .B(n54454), .Z(n54453) );
  NANDN U54928 ( .A(n54421), .B(n54419), .Z(n54454) );
  AND U54929 ( .A(n54455), .B(n54456), .Z(n54422) );
  NANDN U54930 ( .A(n54418), .B(n54457), .Z(n54456) );
  OR U54931 ( .A(n54417), .B(n54415), .Z(n54457) );
  AND U54932 ( .A(n54458), .B(n54459), .Z(n54418) );
  NANDN U54933 ( .A(n54414), .B(n54460), .Z(n54459) );
  NANDN U54934 ( .A(n54413), .B(n54411), .Z(n54460) );
  AND U54935 ( .A(n54461), .B(n54462), .Z(n54414) );
  NANDN U54936 ( .A(n54410), .B(n54463), .Z(n54462) );
  OR U54937 ( .A(n54409), .B(n54407), .Z(n54463) );
  AND U54938 ( .A(n54464), .B(n54465), .Z(n54410) );
  NANDN U54939 ( .A(n54406), .B(n54466), .Z(n54465) );
  NANDN U54940 ( .A(n54405), .B(n54403), .Z(n54466) );
  AND U54941 ( .A(n54467), .B(n54468), .Z(n54406) );
  NANDN U54942 ( .A(n54402), .B(n54469), .Z(n54468) );
  OR U54943 ( .A(n54401), .B(n54399), .Z(n54469) );
  AND U54944 ( .A(n54470), .B(n54471), .Z(n54402) );
  NANDN U54945 ( .A(n54397), .B(n54472), .Z(n54471) );
  NAND U54946 ( .A(n54395), .B(n54398), .Z(n54472) );
  NANDN U54947 ( .A(n54393), .B(n54473), .Z(n54397) );
  AND U54948 ( .A(A[0]), .B(B[88]), .Z(n54473) );
  NAND U54949 ( .A(B[87]), .B(A[1]), .Z(n54393) );
  XNOR U54950 ( .A(n54474), .B(n54475), .Z(n54395) );
  NAND U54951 ( .A(B[89]), .B(A[0]), .Z(n54475) );
  NAND U54952 ( .A(B[87]), .B(A[2]), .Z(n54398) );
  NAND U54953 ( .A(n54399), .B(n54401), .Z(n54467) );
  ANDN U54954 ( .B(A[3]), .A(n29), .Z(n54401) );
  XOR U54955 ( .A(n54476), .B(n54477), .Z(n54399) );
  XNOR U54956 ( .A(n54478), .B(n54479), .Z(n54477) );
  NANDN U54957 ( .A(n54403), .B(n54405), .Z(n54464) );
  ANDN U54958 ( .B(A[4]), .A(n29), .Z(n54405) );
  XNOR U54959 ( .A(n54480), .B(n54481), .Z(n54403) );
  XNOR U54960 ( .A(n54482), .B(n54483), .Z(n54481) );
  NAND U54961 ( .A(n54407), .B(n54409), .Z(n54461) );
  ANDN U54962 ( .B(A[5]), .A(n29), .Z(n54409) );
  XNOR U54963 ( .A(n54484), .B(n54485), .Z(n54407) );
  XNOR U54964 ( .A(n54486), .B(n54487), .Z(n54485) );
  NANDN U54965 ( .A(n54411), .B(n54413), .Z(n54458) );
  ANDN U54966 ( .B(A[6]), .A(n29), .Z(n54413) );
  XNOR U54967 ( .A(n54488), .B(n54489), .Z(n54411) );
  XNOR U54968 ( .A(n54490), .B(n54491), .Z(n54489) );
  NAND U54969 ( .A(n54415), .B(n54417), .Z(n54455) );
  ANDN U54970 ( .B(A[7]), .A(n29), .Z(n54417) );
  XNOR U54971 ( .A(n54492), .B(n54493), .Z(n54415) );
  XNOR U54972 ( .A(n54494), .B(n54495), .Z(n54493) );
  NANDN U54973 ( .A(n54419), .B(n54421), .Z(n54452) );
  ANDN U54974 ( .B(A[8]), .A(n29), .Z(n54421) );
  XNOR U54975 ( .A(n54496), .B(n54497), .Z(n54419) );
  XNOR U54976 ( .A(n54498), .B(n54499), .Z(n54497) );
  NAND U54977 ( .A(n54423), .B(n54425), .Z(n54449) );
  ANDN U54978 ( .B(A[9]), .A(n29), .Z(n54425) );
  XNOR U54979 ( .A(n54500), .B(n54501), .Z(n54423) );
  XNOR U54980 ( .A(n54502), .B(n54503), .Z(n54501) );
  NANDN U54981 ( .A(n54427), .B(n54429), .Z(n54446) );
  ANDN U54982 ( .B(A[10]), .A(n29), .Z(n54429) );
  XNOR U54983 ( .A(n54504), .B(n54505), .Z(n54427) );
  XNOR U54984 ( .A(n54506), .B(n54507), .Z(n54505) );
  NAND U54985 ( .A(n54431), .B(n54433), .Z(n54443) );
  ANDN U54986 ( .B(A[11]), .A(n29), .Z(n54433) );
  XNOR U54987 ( .A(n54508), .B(n54509), .Z(n54431) );
  XNOR U54988 ( .A(n54510), .B(n54511), .Z(n54509) );
  NANDN U54989 ( .A(n54435), .B(n54437), .Z(n54440) );
  ANDN U54990 ( .B(A[12]), .A(n29), .Z(n54437) );
  XNOR U54991 ( .A(n54512), .B(n54513), .Z(n54435) );
  XNOR U54992 ( .A(n54514), .B(n54515), .Z(n54513) );
  ANDN U54993 ( .B(A[13]), .A(n29), .Z(n51947) );
  XNOR U54994 ( .A(n51955), .B(n54516), .Z(n51948) );
  XNOR U54995 ( .A(n51954), .B(n51952), .Z(n54516) );
  AND U54996 ( .A(n54517), .B(n54518), .Z(n51952) );
  NANDN U54997 ( .A(n54515), .B(n54519), .Z(n54518) );
  OR U54998 ( .A(n54514), .B(n54512), .Z(n54519) );
  AND U54999 ( .A(n54520), .B(n54521), .Z(n54515) );
  NANDN U55000 ( .A(n54511), .B(n54522), .Z(n54521) );
  NANDN U55001 ( .A(n54510), .B(n54508), .Z(n54522) );
  AND U55002 ( .A(n54523), .B(n54524), .Z(n54511) );
  NANDN U55003 ( .A(n54507), .B(n54525), .Z(n54524) );
  OR U55004 ( .A(n54506), .B(n54504), .Z(n54525) );
  AND U55005 ( .A(n54526), .B(n54527), .Z(n54507) );
  NANDN U55006 ( .A(n54503), .B(n54528), .Z(n54527) );
  NANDN U55007 ( .A(n54502), .B(n54500), .Z(n54528) );
  AND U55008 ( .A(n54529), .B(n54530), .Z(n54503) );
  NANDN U55009 ( .A(n54499), .B(n54531), .Z(n54530) );
  OR U55010 ( .A(n54498), .B(n54496), .Z(n54531) );
  AND U55011 ( .A(n54532), .B(n54533), .Z(n54499) );
  NANDN U55012 ( .A(n54495), .B(n54534), .Z(n54533) );
  NANDN U55013 ( .A(n54494), .B(n54492), .Z(n54534) );
  AND U55014 ( .A(n54535), .B(n54536), .Z(n54495) );
  NANDN U55015 ( .A(n54491), .B(n54537), .Z(n54536) );
  OR U55016 ( .A(n54490), .B(n54488), .Z(n54537) );
  AND U55017 ( .A(n54538), .B(n54539), .Z(n54491) );
  NANDN U55018 ( .A(n54487), .B(n54540), .Z(n54539) );
  NANDN U55019 ( .A(n54486), .B(n54484), .Z(n54540) );
  AND U55020 ( .A(n54541), .B(n54542), .Z(n54487) );
  NANDN U55021 ( .A(n54483), .B(n54543), .Z(n54542) );
  OR U55022 ( .A(n54482), .B(n54480), .Z(n54543) );
  AND U55023 ( .A(n54544), .B(n54545), .Z(n54483) );
  NANDN U55024 ( .A(n54478), .B(n54546), .Z(n54545) );
  NAND U55025 ( .A(n54476), .B(n54479), .Z(n54546) );
  NANDN U55026 ( .A(n54474), .B(n54547), .Z(n54478) );
  AND U55027 ( .A(A[0]), .B(B[89]), .Z(n54547) );
  NAND U55028 ( .A(B[88]), .B(A[1]), .Z(n54474) );
  XNOR U55029 ( .A(n54548), .B(n54549), .Z(n54476) );
  NAND U55030 ( .A(B[90]), .B(A[0]), .Z(n54549) );
  NAND U55031 ( .A(B[88]), .B(A[2]), .Z(n54479) );
  NAND U55032 ( .A(n54480), .B(n54482), .Z(n54541) );
  ANDN U55033 ( .B(A[3]), .A(n27), .Z(n54482) );
  XOR U55034 ( .A(n54550), .B(n54551), .Z(n54480) );
  XNOR U55035 ( .A(n54552), .B(n54553), .Z(n54551) );
  NANDN U55036 ( .A(n54484), .B(n54486), .Z(n54538) );
  ANDN U55037 ( .B(A[4]), .A(n27), .Z(n54486) );
  XNOR U55038 ( .A(n54554), .B(n54555), .Z(n54484) );
  XNOR U55039 ( .A(n54556), .B(n54557), .Z(n54555) );
  NAND U55040 ( .A(n54488), .B(n54490), .Z(n54535) );
  ANDN U55041 ( .B(A[5]), .A(n27), .Z(n54490) );
  XNOR U55042 ( .A(n54558), .B(n54559), .Z(n54488) );
  XNOR U55043 ( .A(n54560), .B(n54561), .Z(n54559) );
  NANDN U55044 ( .A(n54492), .B(n54494), .Z(n54532) );
  ANDN U55045 ( .B(A[6]), .A(n27), .Z(n54494) );
  XNOR U55046 ( .A(n54562), .B(n54563), .Z(n54492) );
  XNOR U55047 ( .A(n54564), .B(n54565), .Z(n54563) );
  NAND U55048 ( .A(n54496), .B(n54498), .Z(n54529) );
  ANDN U55049 ( .B(A[7]), .A(n27), .Z(n54498) );
  XNOR U55050 ( .A(n54566), .B(n54567), .Z(n54496) );
  XNOR U55051 ( .A(n54568), .B(n54569), .Z(n54567) );
  NANDN U55052 ( .A(n54500), .B(n54502), .Z(n54526) );
  ANDN U55053 ( .B(A[8]), .A(n27), .Z(n54502) );
  XNOR U55054 ( .A(n54570), .B(n54571), .Z(n54500) );
  XNOR U55055 ( .A(n54572), .B(n54573), .Z(n54571) );
  NAND U55056 ( .A(n54504), .B(n54506), .Z(n54523) );
  ANDN U55057 ( .B(A[9]), .A(n27), .Z(n54506) );
  XNOR U55058 ( .A(n54574), .B(n54575), .Z(n54504) );
  XNOR U55059 ( .A(n54576), .B(n54577), .Z(n54575) );
  NANDN U55060 ( .A(n54508), .B(n54510), .Z(n54520) );
  ANDN U55061 ( .B(A[10]), .A(n27), .Z(n54510) );
  XNOR U55062 ( .A(n54578), .B(n54579), .Z(n54508) );
  XNOR U55063 ( .A(n54580), .B(n54581), .Z(n54579) );
  NAND U55064 ( .A(n54512), .B(n54514), .Z(n54517) );
  ANDN U55065 ( .B(A[11]), .A(n27), .Z(n54514) );
  XNOR U55066 ( .A(n54582), .B(n54583), .Z(n54512) );
  XNOR U55067 ( .A(n54584), .B(n54585), .Z(n54583) );
  ANDN U55068 ( .B(A[12]), .A(n27), .Z(n51954) );
  XNOR U55069 ( .A(n51962), .B(n54586), .Z(n51955) );
  XNOR U55070 ( .A(n51961), .B(n51959), .Z(n54586) );
  AND U55071 ( .A(n54587), .B(n54588), .Z(n51959) );
  NANDN U55072 ( .A(n54585), .B(n54589), .Z(n54588) );
  NANDN U55073 ( .A(n54584), .B(n54582), .Z(n54589) );
  AND U55074 ( .A(n54590), .B(n54591), .Z(n54585) );
  NANDN U55075 ( .A(n54581), .B(n54592), .Z(n54591) );
  OR U55076 ( .A(n54580), .B(n54578), .Z(n54592) );
  AND U55077 ( .A(n54593), .B(n54594), .Z(n54581) );
  NANDN U55078 ( .A(n54577), .B(n54595), .Z(n54594) );
  NANDN U55079 ( .A(n54576), .B(n54574), .Z(n54595) );
  AND U55080 ( .A(n54596), .B(n54597), .Z(n54577) );
  NANDN U55081 ( .A(n54573), .B(n54598), .Z(n54597) );
  OR U55082 ( .A(n54572), .B(n54570), .Z(n54598) );
  AND U55083 ( .A(n54599), .B(n54600), .Z(n54573) );
  NANDN U55084 ( .A(n54569), .B(n54601), .Z(n54600) );
  NANDN U55085 ( .A(n54568), .B(n54566), .Z(n54601) );
  AND U55086 ( .A(n54602), .B(n54603), .Z(n54569) );
  NANDN U55087 ( .A(n54565), .B(n54604), .Z(n54603) );
  OR U55088 ( .A(n54564), .B(n54562), .Z(n54604) );
  AND U55089 ( .A(n54605), .B(n54606), .Z(n54565) );
  NANDN U55090 ( .A(n54561), .B(n54607), .Z(n54606) );
  NANDN U55091 ( .A(n54560), .B(n54558), .Z(n54607) );
  AND U55092 ( .A(n54608), .B(n54609), .Z(n54561) );
  NANDN U55093 ( .A(n54557), .B(n54610), .Z(n54609) );
  OR U55094 ( .A(n54556), .B(n54554), .Z(n54610) );
  AND U55095 ( .A(n54611), .B(n54612), .Z(n54557) );
  NANDN U55096 ( .A(n54552), .B(n54613), .Z(n54612) );
  NAND U55097 ( .A(n54550), .B(n54553), .Z(n54613) );
  NANDN U55098 ( .A(n54548), .B(n54614), .Z(n54552) );
  AND U55099 ( .A(A[0]), .B(B[90]), .Z(n54614) );
  NAND U55100 ( .A(B[89]), .B(A[1]), .Z(n54548) );
  XNOR U55101 ( .A(n54615), .B(n54616), .Z(n54550) );
  NAND U55102 ( .A(B[91]), .B(A[0]), .Z(n54616) );
  NAND U55103 ( .A(B[89]), .B(A[2]), .Z(n54553) );
  NAND U55104 ( .A(n54554), .B(n54556), .Z(n54608) );
  ANDN U55105 ( .B(A[3]), .A(n25), .Z(n54556) );
  XOR U55106 ( .A(n54617), .B(n54618), .Z(n54554) );
  XNOR U55107 ( .A(n54619), .B(n54620), .Z(n54618) );
  NANDN U55108 ( .A(n54558), .B(n54560), .Z(n54605) );
  ANDN U55109 ( .B(A[4]), .A(n25), .Z(n54560) );
  XNOR U55110 ( .A(n54621), .B(n54622), .Z(n54558) );
  XNOR U55111 ( .A(n54623), .B(n54624), .Z(n54622) );
  NAND U55112 ( .A(n54562), .B(n54564), .Z(n54602) );
  ANDN U55113 ( .B(A[5]), .A(n25), .Z(n54564) );
  XNOR U55114 ( .A(n54625), .B(n54626), .Z(n54562) );
  XNOR U55115 ( .A(n54627), .B(n54628), .Z(n54626) );
  NANDN U55116 ( .A(n54566), .B(n54568), .Z(n54599) );
  ANDN U55117 ( .B(A[6]), .A(n25), .Z(n54568) );
  XNOR U55118 ( .A(n54629), .B(n54630), .Z(n54566) );
  XNOR U55119 ( .A(n54631), .B(n54632), .Z(n54630) );
  NAND U55120 ( .A(n54570), .B(n54572), .Z(n54596) );
  ANDN U55121 ( .B(A[7]), .A(n25), .Z(n54572) );
  XNOR U55122 ( .A(n54633), .B(n54634), .Z(n54570) );
  XNOR U55123 ( .A(n54635), .B(n54636), .Z(n54634) );
  NANDN U55124 ( .A(n54574), .B(n54576), .Z(n54593) );
  ANDN U55125 ( .B(A[8]), .A(n25), .Z(n54576) );
  XNOR U55126 ( .A(n54637), .B(n54638), .Z(n54574) );
  XNOR U55127 ( .A(n54639), .B(n54640), .Z(n54638) );
  NAND U55128 ( .A(n54578), .B(n54580), .Z(n54590) );
  ANDN U55129 ( .B(A[9]), .A(n25), .Z(n54580) );
  XNOR U55130 ( .A(n54641), .B(n54642), .Z(n54578) );
  XNOR U55131 ( .A(n54643), .B(n54644), .Z(n54642) );
  NANDN U55132 ( .A(n54582), .B(n54584), .Z(n54587) );
  ANDN U55133 ( .B(A[10]), .A(n25), .Z(n54584) );
  XNOR U55134 ( .A(n54645), .B(n54646), .Z(n54582) );
  XNOR U55135 ( .A(n54647), .B(n54648), .Z(n54646) );
  ANDN U55136 ( .B(A[11]), .A(n25), .Z(n51961) );
  XNOR U55137 ( .A(n51969), .B(n54649), .Z(n51962) );
  XNOR U55138 ( .A(n51968), .B(n51966), .Z(n54649) );
  AND U55139 ( .A(n54650), .B(n54651), .Z(n51966) );
  NANDN U55140 ( .A(n54648), .B(n54652), .Z(n54651) );
  OR U55141 ( .A(n54647), .B(n54645), .Z(n54652) );
  AND U55142 ( .A(n54653), .B(n54654), .Z(n54648) );
  NANDN U55143 ( .A(n54644), .B(n54655), .Z(n54654) );
  NANDN U55144 ( .A(n54643), .B(n54641), .Z(n54655) );
  AND U55145 ( .A(n54656), .B(n54657), .Z(n54644) );
  NANDN U55146 ( .A(n54640), .B(n54658), .Z(n54657) );
  OR U55147 ( .A(n54639), .B(n54637), .Z(n54658) );
  AND U55148 ( .A(n54659), .B(n54660), .Z(n54640) );
  NANDN U55149 ( .A(n54636), .B(n54661), .Z(n54660) );
  NANDN U55150 ( .A(n54635), .B(n54633), .Z(n54661) );
  AND U55151 ( .A(n54662), .B(n54663), .Z(n54636) );
  NANDN U55152 ( .A(n54632), .B(n54664), .Z(n54663) );
  OR U55153 ( .A(n54631), .B(n54629), .Z(n54664) );
  AND U55154 ( .A(n54665), .B(n54666), .Z(n54632) );
  NANDN U55155 ( .A(n54628), .B(n54667), .Z(n54666) );
  NANDN U55156 ( .A(n54627), .B(n54625), .Z(n54667) );
  AND U55157 ( .A(n54668), .B(n54669), .Z(n54628) );
  NANDN U55158 ( .A(n54624), .B(n54670), .Z(n54669) );
  OR U55159 ( .A(n54623), .B(n54621), .Z(n54670) );
  AND U55160 ( .A(n54671), .B(n54672), .Z(n54624) );
  NANDN U55161 ( .A(n54619), .B(n54673), .Z(n54672) );
  NAND U55162 ( .A(n54617), .B(n54620), .Z(n54673) );
  NANDN U55163 ( .A(n54615), .B(n54674), .Z(n54619) );
  AND U55164 ( .A(A[0]), .B(B[91]), .Z(n54674) );
  NAND U55165 ( .A(B[90]), .B(A[1]), .Z(n54615) );
  XNOR U55166 ( .A(n54675), .B(n54676), .Z(n54617) );
  NAND U55167 ( .A(B[92]), .B(A[0]), .Z(n54676) );
  NAND U55168 ( .A(B[90]), .B(A[2]), .Z(n54620) );
  NAND U55169 ( .A(n54621), .B(n54623), .Z(n54668) );
  ANDN U55170 ( .B(A[3]), .A(n23), .Z(n54623) );
  XOR U55171 ( .A(n54677), .B(n54678), .Z(n54621) );
  XNOR U55172 ( .A(n54679), .B(n54680), .Z(n54678) );
  NANDN U55173 ( .A(n54625), .B(n54627), .Z(n54665) );
  ANDN U55174 ( .B(A[4]), .A(n23), .Z(n54627) );
  XNOR U55175 ( .A(n54681), .B(n54682), .Z(n54625) );
  XNOR U55176 ( .A(n54683), .B(n54684), .Z(n54682) );
  NAND U55177 ( .A(n54629), .B(n54631), .Z(n54662) );
  ANDN U55178 ( .B(A[5]), .A(n23), .Z(n54631) );
  XNOR U55179 ( .A(n54685), .B(n54686), .Z(n54629) );
  XNOR U55180 ( .A(n54687), .B(n54688), .Z(n54686) );
  NANDN U55181 ( .A(n54633), .B(n54635), .Z(n54659) );
  ANDN U55182 ( .B(A[6]), .A(n23), .Z(n54635) );
  XNOR U55183 ( .A(n54689), .B(n54690), .Z(n54633) );
  XNOR U55184 ( .A(n54691), .B(n54692), .Z(n54690) );
  NAND U55185 ( .A(n54637), .B(n54639), .Z(n54656) );
  ANDN U55186 ( .B(A[7]), .A(n23), .Z(n54639) );
  XNOR U55187 ( .A(n54693), .B(n54694), .Z(n54637) );
  XNOR U55188 ( .A(n54695), .B(n54696), .Z(n54694) );
  NANDN U55189 ( .A(n54641), .B(n54643), .Z(n54653) );
  ANDN U55190 ( .B(A[8]), .A(n23), .Z(n54643) );
  XNOR U55191 ( .A(n54697), .B(n54698), .Z(n54641) );
  XNOR U55192 ( .A(n54699), .B(n54700), .Z(n54698) );
  NAND U55193 ( .A(n54645), .B(n54647), .Z(n54650) );
  ANDN U55194 ( .B(A[9]), .A(n23), .Z(n54647) );
  XNOR U55195 ( .A(n54701), .B(n54702), .Z(n54645) );
  XNOR U55196 ( .A(n54703), .B(n54704), .Z(n54702) );
  ANDN U55197 ( .B(A[10]), .A(n23), .Z(n51968) );
  XNOR U55198 ( .A(n51976), .B(n54705), .Z(n51969) );
  XNOR U55199 ( .A(n51975), .B(n51973), .Z(n54705) );
  AND U55200 ( .A(n54706), .B(n54707), .Z(n51973) );
  NANDN U55201 ( .A(n54704), .B(n54708), .Z(n54707) );
  NANDN U55202 ( .A(n54703), .B(n54701), .Z(n54708) );
  AND U55203 ( .A(n54709), .B(n54710), .Z(n54704) );
  NANDN U55204 ( .A(n54700), .B(n54711), .Z(n54710) );
  OR U55205 ( .A(n54699), .B(n54697), .Z(n54711) );
  AND U55206 ( .A(n54712), .B(n54713), .Z(n54700) );
  NANDN U55207 ( .A(n54696), .B(n54714), .Z(n54713) );
  NANDN U55208 ( .A(n54695), .B(n54693), .Z(n54714) );
  AND U55209 ( .A(n54715), .B(n54716), .Z(n54696) );
  NANDN U55210 ( .A(n54692), .B(n54717), .Z(n54716) );
  OR U55211 ( .A(n54691), .B(n54689), .Z(n54717) );
  AND U55212 ( .A(n54718), .B(n54719), .Z(n54692) );
  NANDN U55213 ( .A(n54688), .B(n54720), .Z(n54719) );
  NANDN U55214 ( .A(n54687), .B(n54685), .Z(n54720) );
  AND U55215 ( .A(n54721), .B(n54722), .Z(n54688) );
  NANDN U55216 ( .A(n54684), .B(n54723), .Z(n54722) );
  OR U55217 ( .A(n54683), .B(n54681), .Z(n54723) );
  AND U55218 ( .A(n54724), .B(n54725), .Z(n54684) );
  NANDN U55219 ( .A(n54679), .B(n54726), .Z(n54725) );
  NAND U55220 ( .A(n54677), .B(n54680), .Z(n54726) );
  NANDN U55221 ( .A(n54675), .B(n54727), .Z(n54679) );
  AND U55222 ( .A(A[0]), .B(B[92]), .Z(n54727) );
  NAND U55223 ( .A(B[91]), .B(A[1]), .Z(n54675) );
  XNOR U55224 ( .A(n54728), .B(n54729), .Z(n54677) );
  NAND U55225 ( .A(B[93]), .B(A[0]), .Z(n54729) );
  NAND U55226 ( .A(B[91]), .B(A[2]), .Z(n54680) );
  NAND U55227 ( .A(n54681), .B(n54683), .Z(n54721) );
  ANDN U55228 ( .B(A[3]), .A(n21), .Z(n54683) );
  XOR U55229 ( .A(n54730), .B(n54731), .Z(n54681) );
  XNOR U55230 ( .A(n54732), .B(n54733), .Z(n54731) );
  NANDN U55231 ( .A(n54685), .B(n54687), .Z(n54718) );
  ANDN U55232 ( .B(A[4]), .A(n21), .Z(n54687) );
  XNOR U55233 ( .A(n54734), .B(n54735), .Z(n54685) );
  XNOR U55234 ( .A(n54736), .B(n54737), .Z(n54735) );
  NAND U55235 ( .A(n54689), .B(n54691), .Z(n54715) );
  ANDN U55236 ( .B(A[5]), .A(n21), .Z(n54691) );
  XNOR U55237 ( .A(n54738), .B(n54739), .Z(n54689) );
  XNOR U55238 ( .A(n54740), .B(n54741), .Z(n54739) );
  NANDN U55239 ( .A(n54693), .B(n54695), .Z(n54712) );
  ANDN U55240 ( .B(A[6]), .A(n21), .Z(n54695) );
  XNOR U55241 ( .A(n54742), .B(n54743), .Z(n54693) );
  XNOR U55242 ( .A(n54744), .B(n54745), .Z(n54743) );
  NAND U55243 ( .A(n54697), .B(n54699), .Z(n54709) );
  ANDN U55244 ( .B(A[7]), .A(n21), .Z(n54699) );
  XNOR U55245 ( .A(n54746), .B(n54747), .Z(n54697) );
  XNOR U55246 ( .A(n54748), .B(n54749), .Z(n54747) );
  NANDN U55247 ( .A(n54701), .B(n54703), .Z(n54706) );
  ANDN U55248 ( .B(A[8]), .A(n21), .Z(n54703) );
  XNOR U55249 ( .A(n54750), .B(n54751), .Z(n54701) );
  XNOR U55250 ( .A(n54752), .B(n54753), .Z(n54751) );
  ANDN U55251 ( .B(A[9]), .A(n21), .Z(n51975) );
  XNOR U55252 ( .A(n51983), .B(n54754), .Z(n51976) );
  XNOR U55253 ( .A(n51982), .B(n51980), .Z(n54754) );
  AND U55254 ( .A(n54755), .B(n54756), .Z(n51980) );
  NANDN U55255 ( .A(n54753), .B(n54757), .Z(n54756) );
  OR U55256 ( .A(n54752), .B(n54750), .Z(n54757) );
  AND U55257 ( .A(n54758), .B(n54759), .Z(n54753) );
  NANDN U55258 ( .A(n54749), .B(n54760), .Z(n54759) );
  NANDN U55259 ( .A(n54748), .B(n54746), .Z(n54760) );
  AND U55260 ( .A(n54761), .B(n54762), .Z(n54749) );
  NANDN U55261 ( .A(n54745), .B(n54763), .Z(n54762) );
  OR U55262 ( .A(n54744), .B(n54742), .Z(n54763) );
  AND U55263 ( .A(n54764), .B(n54765), .Z(n54745) );
  NANDN U55264 ( .A(n54741), .B(n54766), .Z(n54765) );
  NANDN U55265 ( .A(n54740), .B(n54738), .Z(n54766) );
  AND U55266 ( .A(n54767), .B(n54768), .Z(n54741) );
  NANDN U55267 ( .A(n54737), .B(n54769), .Z(n54768) );
  OR U55268 ( .A(n54736), .B(n54734), .Z(n54769) );
  AND U55269 ( .A(n54770), .B(n54771), .Z(n54737) );
  NANDN U55270 ( .A(n54732), .B(n54772), .Z(n54771) );
  NAND U55271 ( .A(n54730), .B(n54733), .Z(n54772) );
  NANDN U55272 ( .A(n54728), .B(n54773), .Z(n54732) );
  AND U55273 ( .A(A[0]), .B(B[93]), .Z(n54773) );
  NAND U55274 ( .A(B[92]), .B(A[1]), .Z(n54728) );
  XNOR U55275 ( .A(n54774), .B(n54775), .Z(n54730) );
  NAND U55276 ( .A(B[94]), .B(A[0]), .Z(n54775) );
  NAND U55277 ( .A(B[92]), .B(A[2]), .Z(n54733) );
  NAND U55278 ( .A(n54734), .B(n54736), .Z(n54767) );
  ANDN U55279 ( .B(A[3]), .A(n19), .Z(n54736) );
  XOR U55280 ( .A(n54776), .B(n54777), .Z(n54734) );
  XNOR U55281 ( .A(n54778), .B(n54779), .Z(n54777) );
  NANDN U55282 ( .A(n54738), .B(n54740), .Z(n54764) );
  ANDN U55283 ( .B(A[4]), .A(n19), .Z(n54740) );
  XNOR U55284 ( .A(n54780), .B(n54781), .Z(n54738) );
  XNOR U55285 ( .A(n54782), .B(n54783), .Z(n54781) );
  NAND U55286 ( .A(n54742), .B(n54744), .Z(n54761) );
  ANDN U55287 ( .B(A[5]), .A(n19), .Z(n54744) );
  XNOR U55288 ( .A(n54784), .B(n54785), .Z(n54742) );
  XNOR U55289 ( .A(n54786), .B(n54787), .Z(n54785) );
  NANDN U55290 ( .A(n54746), .B(n54748), .Z(n54758) );
  ANDN U55291 ( .B(A[6]), .A(n19), .Z(n54748) );
  XNOR U55292 ( .A(n54788), .B(n54789), .Z(n54746) );
  XNOR U55293 ( .A(n54790), .B(n54791), .Z(n54789) );
  NAND U55294 ( .A(n54750), .B(n54752), .Z(n54755) );
  ANDN U55295 ( .B(A[7]), .A(n19), .Z(n54752) );
  XNOR U55296 ( .A(n54792), .B(n54793), .Z(n54750) );
  XNOR U55297 ( .A(n54794), .B(n54795), .Z(n54793) );
  ANDN U55298 ( .B(A[8]), .A(n19), .Z(n51982) );
  XNOR U55299 ( .A(n51990), .B(n54796), .Z(n51983) );
  XNOR U55300 ( .A(n51989), .B(n51987), .Z(n54796) );
  AND U55301 ( .A(n54797), .B(n54798), .Z(n51987) );
  NANDN U55302 ( .A(n54795), .B(n54799), .Z(n54798) );
  NANDN U55303 ( .A(n54794), .B(n54792), .Z(n54799) );
  AND U55304 ( .A(n54800), .B(n54801), .Z(n54795) );
  NANDN U55305 ( .A(n54791), .B(n54802), .Z(n54801) );
  OR U55306 ( .A(n54790), .B(n54788), .Z(n54802) );
  AND U55307 ( .A(n54803), .B(n54804), .Z(n54791) );
  NANDN U55308 ( .A(n54787), .B(n54805), .Z(n54804) );
  NANDN U55309 ( .A(n54786), .B(n54784), .Z(n54805) );
  AND U55310 ( .A(n54806), .B(n54807), .Z(n54787) );
  NANDN U55311 ( .A(n54783), .B(n54808), .Z(n54807) );
  OR U55312 ( .A(n54782), .B(n54780), .Z(n54808) );
  AND U55313 ( .A(n54809), .B(n54810), .Z(n54783) );
  NANDN U55314 ( .A(n54778), .B(n54811), .Z(n54810) );
  NAND U55315 ( .A(n54776), .B(n54779), .Z(n54811) );
  NANDN U55316 ( .A(n54774), .B(n54812), .Z(n54778) );
  AND U55317 ( .A(A[0]), .B(B[94]), .Z(n54812) );
  NAND U55318 ( .A(B[93]), .B(A[1]), .Z(n54774) );
  XNOR U55319 ( .A(n54813), .B(n54814), .Z(n54776) );
  NAND U55320 ( .A(B[95]), .B(A[0]), .Z(n54814) );
  NAND U55321 ( .A(B[93]), .B(A[2]), .Z(n54779) );
  NAND U55322 ( .A(n54780), .B(n54782), .Z(n54806) );
  ANDN U55323 ( .B(A[3]), .A(n17), .Z(n54782) );
  XOR U55324 ( .A(n54815), .B(n54816), .Z(n54780) );
  XNOR U55325 ( .A(n54817), .B(n54818), .Z(n54816) );
  NANDN U55326 ( .A(n54784), .B(n54786), .Z(n54803) );
  ANDN U55327 ( .B(A[4]), .A(n17), .Z(n54786) );
  XNOR U55328 ( .A(n54819), .B(n54820), .Z(n54784) );
  XNOR U55329 ( .A(n54821), .B(n54822), .Z(n54820) );
  NAND U55330 ( .A(n54788), .B(n54790), .Z(n54800) );
  ANDN U55331 ( .B(A[5]), .A(n17), .Z(n54790) );
  XNOR U55332 ( .A(n54823), .B(n54824), .Z(n54788) );
  XNOR U55333 ( .A(n54825), .B(n54826), .Z(n54824) );
  NANDN U55334 ( .A(n54792), .B(n54794), .Z(n54797) );
  ANDN U55335 ( .B(A[6]), .A(n17), .Z(n54794) );
  XNOR U55336 ( .A(n54827), .B(n54828), .Z(n54792) );
  XNOR U55337 ( .A(n54829), .B(n54830), .Z(n54828) );
  ANDN U55338 ( .B(A[7]), .A(n17), .Z(n51989) );
  XNOR U55339 ( .A(n51997), .B(n54831), .Z(n51990) );
  XNOR U55340 ( .A(n51996), .B(n51994), .Z(n54831) );
  AND U55341 ( .A(n54832), .B(n54833), .Z(n51994) );
  NANDN U55342 ( .A(n54830), .B(n54834), .Z(n54833) );
  OR U55343 ( .A(n54829), .B(n54827), .Z(n54834) );
  AND U55344 ( .A(n54835), .B(n54836), .Z(n54830) );
  NANDN U55345 ( .A(n54826), .B(n54837), .Z(n54836) );
  NANDN U55346 ( .A(n54825), .B(n54823), .Z(n54837) );
  AND U55347 ( .A(n54838), .B(n54839), .Z(n54826) );
  NANDN U55348 ( .A(n54822), .B(n54840), .Z(n54839) );
  OR U55349 ( .A(n54821), .B(n54819), .Z(n54840) );
  AND U55350 ( .A(n54841), .B(n54842), .Z(n54822) );
  NANDN U55351 ( .A(n54817), .B(n54843), .Z(n54842) );
  NAND U55352 ( .A(n54815), .B(n54818), .Z(n54843) );
  NANDN U55353 ( .A(n54813), .B(n54844), .Z(n54817) );
  AND U55354 ( .A(A[0]), .B(B[95]), .Z(n54844) );
  NAND U55355 ( .A(B[94]), .B(A[1]), .Z(n54813) );
  XNOR U55356 ( .A(n54845), .B(n54846), .Z(n54815) );
  NAND U55357 ( .A(B[96]), .B(A[0]), .Z(n54846) );
  NAND U55358 ( .A(B[94]), .B(A[2]), .Z(n54818) );
  NAND U55359 ( .A(n54819), .B(n54821), .Z(n54838) );
  ANDN U55360 ( .B(A[3]), .A(n15), .Z(n54821) );
  XOR U55361 ( .A(n54847), .B(n54848), .Z(n54819) );
  XNOR U55362 ( .A(n54849), .B(n54850), .Z(n54848) );
  NANDN U55363 ( .A(n54823), .B(n54825), .Z(n54835) );
  ANDN U55364 ( .B(A[4]), .A(n15), .Z(n54825) );
  XNOR U55365 ( .A(n54851), .B(n54852), .Z(n54823) );
  XNOR U55366 ( .A(n54853), .B(n54854), .Z(n54852) );
  NAND U55367 ( .A(n54827), .B(n54829), .Z(n54832) );
  ANDN U55368 ( .B(A[5]), .A(n15), .Z(n54829) );
  XNOR U55369 ( .A(n54855), .B(n54856), .Z(n54827) );
  XNOR U55370 ( .A(n54857), .B(n54858), .Z(n54856) );
  ANDN U55371 ( .B(A[6]), .A(n15), .Z(n51996) );
  XNOR U55372 ( .A(n52004), .B(n54859), .Z(n51997) );
  XNOR U55373 ( .A(n52003), .B(n52001), .Z(n54859) );
  AND U55374 ( .A(n54860), .B(n54861), .Z(n52001) );
  NANDN U55375 ( .A(n54858), .B(n54862), .Z(n54861) );
  NANDN U55376 ( .A(n54857), .B(n54855), .Z(n54862) );
  AND U55377 ( .A(n54863), .B(n54864), .Z(n54858) );
  NANDN U55378 ( .A(n54854), .B(n54865), .Z(n54864) );
  OR U55379 ( .A(n54853), .B(n54851), .Z(n54865) );
  AND U55380 ( .A(n54866), .B(n54867), .Z(n54854) );
  NANDN U55381 ( .A(n54849), .B(n54868), .Z(n54867) );
  NAND U55382 ( .A(n54847), .B(n54850), .Z(n54868) );
  NANDN U55383 ( .A(n54845), .B(n54869), .Z(n54849) );
  AND U55384 ( .A(A[0]), .B(B[96]), .Z(n54869) );
  NAND U55385 ( .A(B[95]), .B(A[1]), .Z(n54845) );
  XNOR U55386 ( .A(n54870), .B(n54871), .Z(n54847) );
  NAND U55387 ( .A(B[97]), .B(A[0]), .Z(n54871) );
  NAND U55388 ( .A(B[95]), .B(A[2]), .Z(n54850) );
  NAND U55389 ( .A(n54851), .B(n54853), .Z(n54863) );
  ANDN U55390 ( .B(A[3]), .A(n13), .Z(n54853) );
  XOR U55391 ( .A(n54872), .B(n54873), .Z(n54851) );
  XNOR U55392 ( .A(n54874), .B(n54875), .Z(n54873) );
  NANDN U55393 ( .A(n54855), .B(n54857), .Z(n54860) );
  ANDN U55394 ( .B(A[4]), .A(n13), .Z(n54857) );
  XNOR U55395 ( .A(n54876), .B(n54877), .Z(n54855) );
  XNOR U55396 ( .A(n54878), .B(n54879), .Z(n54877) );
  ANDN U55397 ( .B(A[5]), .A(n13), .Z(n52003) );
  XNOR U55398 ( .A(n52011), .B(n54880), .Z(n52004) );
  XNOR U55399 ( .A(n52010), .B(n52008), .Z(n54880) );
  AND U55400 ( .A(n54881), .B(n54882), .Z(n52008) );
  NANDN U55401 ( .A(n54879), .B(n54883), .Z(n54882) );
  OR U55402 ( .A(n54878), .B(n54876), .Z(n54883) );
  AND U55403 ( .A(n54884), .B(n54885), .Z(n54879) );
  NANDN U55404 ( .A(n54874), .B(n54886), .Z(n54885) );
  NAND U55405 ( .A(n54872), .B(n54875), .Z(n54886) );
  NANDN U55406 ( .A(n54870), .B(n54887), .Z(n54874) );
  AND U55407 ( .A(A[0]), .B(B[97]), .Z(n54887) );
  NAND U55408 ( .A(B[96]), .B(A[1]), .Z(n54870) );
  XNOR U55409 ( .A(n54888), .B(n54889), .Z(n54872) );
  NAND U55410 ( .A(B[98]), .B(A[0]), .Z(n54889) );
  NAND U55411 ( .A(B[96]), .B(A[2]), .Z(n54875) );
  NAND U55412 ( .A(n54876), .B(n54878), .Z(n54881) );
  ANDN U55413 ( .B(A[3]), .A(n11), .Z(n54878) );
  XOR U55414 ( .A(n54890), .B(n54891), .Z(n54876) );
  XNOR U55415 ( .A(n54892), .B(n54893), .Z(n54891) );
  ANDN U55416 ( .B(A[4]), .A(n11), .Z(n52010) );
  XNOR U55417 ( .A(n52018), .B(n54894), .Z(n52011) );
  XNOR U55418 ( .A(n52017), .B(n52015), .Z(n54894) );
  AND U55419 ( .A(n54895), .B(n54896), .Z(n52015) );
  NANDN U55420 ( .A(n54892), .B(n54897), .Z(n54896) );
  NAND U55421 ( .A(n54890), .B(n54893), .Z(n54897) );
  NANDN U55422 ( .A(n54888), .B(n54898), .Z(n54892) );
  AND U55423 ( .A(A[0]), .B(B[98]), .Z(n54898) );
  NAND U55424 ( .A(B[97]), .B(A[1]), .Z(n54888) );
  XNOR U55425 ( .A(n54899), .B(n54900), .Z(n54890) );
  NAND U55426 ( .A(B[99]), .B(A[0]), .Z(n54900) );
  NAND U55427 ( .A(B[97]), .B(A[2]), .Z(n54893) );
  ANDN U55428 ( .B(A[3]), .A(n9), .Z(n52017) );
  XNOR U55429 ( .A(n52024), .B(n54901), .Z(n52018) );
  XNOR U55430 ( .A(n52022), .B(n52025), .Z(n54901) );
  NAND U55431 ( .A(B[98]), .B(A[2]), .Z(n52025) );
  NANDN U55432 ( .A(n54899), .B(n54902), .Z(n52022) );
  AND U55433 ( .A(A[0]), .B(B[99]), .Z(n54902) );
  NAND U55434 ( .A(B[98]), .B(A[1]), .Z(n54899) );
  XOR U55435 ( .A(n52027), .B(n54903), .Z(n52024) );
  NAND U55436 ( .A(B[100]), .B(A[0]), .Z(n54903) );
  NAND U55437 ( .A(B[99]), .B(A[1]), .Z(n52027) );
  XNOR U55438 ( .A(n49378), .B(n54904), .Z(\A1[0] ) );
  XNOR U55439 ( .A(n49375), .B(n49377), .Z(n54904) );
  ANDN U55440 ( .B(n85), .A(n84), .Z(n49377) );
  NAND U55441 ( .A(B[0]), .B(A[1]), .Z(n84) );
  AND U55442 ( .A(A[0]), .B(B[1]), .Z(n85) );
  NAND U55443 ( .A(B[0]), .B(A[2]), .Z(n49375) );
  XNOR U55444 ( .A(n49411), .B(n54905), .Z(n49378) );
  NAND U55445 ( .A(A[0]), .B(B[2]), .Z(n54905) );
  NAND U55446 ( .A(B[1]), .B(A[1]), .Z(n49411) );
endmodule


module mult_N256_CC8 ( clk, rst, a, b, c );
  input [255:0] a;
  input [31:0] b;
  output [255:0] c;
  input clk, rst;

  wire   [255:32] swire;
  wire   [511:256] sreg;
  wire   [255:0] clocal;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31;

  DFF \sreg_reg[256]  ( .D(swire[32]), .CLK(clk), .RST(rst), .Q(sreg[256]) );
  DFF \sreg_reg[257]  ( .D(swire[33]), .CLK(clk), .RST(rst), .Q(sreg[257]) );
  DFF \sreg_reg[258]  ( .D(swire[34]), .CLK(clk), .RST(rst), .Q(sreg[258]) );
  DFF \sreg_reg[259]  ( .D(swire[35]), .CLK(clk), .RST(rst), .Q(sreg[259]) );
  DFF \sreg_reg[260]  ( .D(swire[36]), .CLK(clk), .RST(rst), .Q(sreg[260]) );
  DFF \sreg_reg[261]  ( .D(swire[37]), .CLK(clk), .RST(rst), .Q(sreg[261]) );
  DFF \sreg_reg[262]  ( .D(swire[38]), .CLK(clk), .RST(rst), .Q(sreg[262]) );
  DFF \sreg_reg[263]  ( .D(swire[39]), .CLK(clk), .RST(rst), .Q(sreg[263]) );
  DFF \sreg_reg[264]  ( .D(swire[40]), .CLK(clk), .RST(rst), .Q(sreg[264]) );
  DFF \sreg_reg[265]  ( .D(swire[41]), .CLK(clk), .RST(rst), .Q(sreg[265]) );
  DFF \sreg_reg[266]  ( .D(swire[42]), .CLK(clk), .RST(rst), .Q(sreg[266]) );
  DFF \sreg_reg[267]  ( .D(swire[43]), .CLK(clk), .RST(rst), .Q(sreg[267]) );
  DFF \sreg_reg[268]  ( .D(swire[44]), .CLK(clk), .RST(rst), .Q(sreg[268]) );
  DFF \sreg_reg[269]  ( .D(swire[45]), .CLK(clk), .RST(rst), .Q(sreg[269]) );
  DFF \sreg_reg[270]  ( .D(swire[46]), .CLK(clk), .RST(rst), .Q(sreg[270]) );
  DFF \sreg_reg[271]  ( .D(swire[47]), .CLK(clk), .RST(rst), .Q(sreg[271]) );
  DFF \sreg_reg[272]  ( .D(swire[48]), .CLK(clk), .RST(rst), .Q(sreg[272]) );
  DFF \sreg_reg[273]  ( .D(swire[49]), .CLK(clk), .RST(rst), .Q(sreg[273]) );
  DFF \sreg_reg[274]  ( .D(swire[50]), .CLK(clk), .RST(rst), .Q(sreg[274]) );
  DFF \sreg_reg[275]  ( .D(swire[51]), .CLK(clk), .RST(rst), .Q(sreg[275]) );
  DFF \sreg_reg[276]  ( .D(swire[52]), .CLK(clk), .RST(rst), .Q(sreg[276]) );
  DFF \sreg_reg[277]  ( .D(swire[53]), .CLK(clk), .RST(rst), .Q(sreg[277]) );
  DFF \sreg_reg[278]  ( .D(swire[54]), .CLK(clk), .RST(rst), .Q(sreg[278]) );
  DFF \sreg_reg[279]  ( .D(swire[55]), .CLK(clk), .RST(rst), .Q(sreg[279]) );
  DFF \sreg_reg[280]  ( .D(swire[56]), .CLK(clk), .RST(rst), .Q(sreg[280]) );
  DFF \sreg_reg[281]  ( .D(swire[57]), .CLK(clk), .RST(rst), .Q(sreg[281]) );
  DFF \sreg_reg[282]  ( .D(swire[58]), .CLK(clk), .RST(rst), .Q(sreg[282]) );
  DFF \sreg_reg[283]  ( .D(swire[59]), .CLK(clk), .RST(rst), .Q(sreg[283]) );
  DFF \sreg_reg[284]  ( .D(swire[60]), .CLK(clk), .RST(rst), .Q(sreg[284]) );
  DFF \sreg_reg[285]  ( .D(swire[61]), .CLK(clk), .RST(rst), .Q(sreg[285]) );
  DFF \sreg_reg[286]  ( .D(swire[62]), .CLK(clk), .RST(rst), .Q(sreg[286]) );
  DFF \sreg_reg[287]  ( .D(swire[63]), .CLK(clk), .RST(rst), .Q(sreg[287]) );
  DFF \sreg_reg[288]  ( .D(swire[64]), .CLK(clk), .RST(rst), .Q(sreg[288]) );
  DFF \sreg_reg[289]  ( .D(swire[65]), .CLK(clk), .RST(rst), .Q(sreg[289]) );
  DFF \sreg_reg[290]  ( .D(swire[66]), .CLK(clk), .RST(rst), .Q(sreg[290]) );
  DFF \sreg_reg[291]  ( .D(swire[67]), .CLK(clk), .RST(rst), .Q(sreg[291]) );
  DFF \sreg_reg[292]  ( .D(swire[68]), .CLK(clk), .RST(rst), .Q(sreg[292]) );
  DFF \sreg_reg[293]  ( .D(swire[69]), .CLK(clk), .RST(rst), .Q(sreg[293]) );
  DFF \sreg_reg[294]  ( .D(swire[70]), .CLK(clk), .RST(rst), .Q(sreg[294]) );
  DFF \sreg_reg[295]  ( .D(swire[71]), .CLK(clk), .RST(rst), .Q(sreg[295]) );
  DFF \sreg_reg[296]  ( .D(swire[72]), .CLK(clk), .RST(rst), .Q(sreg[296]) );
  DFF \sreg_reg[297]  ( .D(swire[73]), .CLK(clk), .RST(rst), .Q(sreg[297]) );
  DFF \sreg_reg[298]  ( .D(swire[74]), .CLK(clk), .RST(rst), .Q(sreg[298]) );
  DFF \sreg_reg[299]  ( .D(swire[75]), .CLK(clk), .RST(rst), .Q(sreg[299]) );
  DFF \sreg_reg[300]  ( .D(swire[76]), .CLK(clk), .RST(rst), .Q(sreg[300]) );
  DFF \sreg_reg[301]  ( .D(swire[77]), .CLK(clk), .RST(rst), .Q(sreg[301]) );
  DFF \sreg_reg[302]  ( .D(swire[78]), .CLK(clk), .RST(rst), .Q(sreg[302]) );
  DFF \sreg_reg[303]  ( .D(swire[79]), .CLK(clk), .RST(rst), .Q(sreg[303]) );
  DFF \sreg_reg[304]  ( .D(swire[80]), .CLK(clk), .RST(rst), .Q(sreg[304]) );
  DFF \sreg_reg[305]  ( .D(swire[81]), .CLK(clk), .RST(rst), .Q(sreg[305]) );
  DFF \sreg_reg[306]  ( .D(swire[82]), .CLK(clk), .RST(rst), .Q(sreg[306]) );
  DFF \sreg_reg[307]  ( .D(swire[83]), .CLK(clk), .RST(rst), .Q(sreg[307]) );
  DFF \sreg_reg[308]  ( .D(swire[84]), .CLK(clk), .RST(rst), .Q(sreg[308]) );
  DFF \sreg_reg[309]  ( .D(swire[85]), .CLK(clk), .RST(rst), .Q(sreg[309]) );
  DFF \sreg_reg[310]  ( .D(swire[86]), .CLK(clk), .RST(rst), .Q(sreg[310]) );
  DFF \sreg_reg[311]  ( .D(swire[87]), .CLK(clk), .RST(rst), .Q(sreg[311]) );
  DFF \sreg_reg[312]  ( .D(swire[88]), .CLK(clk), .RST(rst), .Q(sreg[312]) );
  DFF \sreg_reg[313]  ( .D(swire[89]), .CLK(clk), .RST(rst), .Q(sreg[313]) );
  DFF \sreg_reg[314]  ( .D(swire[90]), .CLK(clk), .RST(rst), .Q(sreg[314]) );
  DFF \sreg_reg[315]  ( .D(swire[91]), .CLK(clk), .RST(rst), .Q(sreg[315]) );
  DFF \sreg_reg[316]  ( .D(swire[92]), .CLK(clk), .RST(rst), .Q(sreg[316]) );
  DFF \sreg_reg[317]  ( .D(swire[93]), .CLK(clk), .RST(rst), .Q(sreg[317]) );
  DFF \sreg_reg[318]  ( .D(swire[94]), .CLK(clk), .RST(rst), .Q(sreg[318]) );
  DFF \sreg_reg[319]  ( .D(swire[95]), .CLK(clk), .RST(rst), .Q(sreg[319]) );
  DFF \sreg_reg[320]  ( .D(swire[96]), .CLK(clk), .RST(rst), .Q(sreg[320]) );
  DFF \sreg_reg[321]  ( .D(swire[97]), .CLK(clk), .RST(rst), .Q(sreg[321]) );
  DFF \sreg_reg[322]  ( .D(swire[98]), .CLK(clk), .RST(rst), .Q(sreg[322]) );
  DFF \sreg_reg[323]  ( .D(swire[99]), .CLK(clk), .RST(rst), .Q(sreg[323]) );
  DFF \sreg_reg[324]  ( .D(swire[100]), .CLK(clk), .RST(rst), .Q(sreg[324]) );
  DFF \sreg_reg[325]  ( .D(swire[101]), .CLK(clk), .RST(rst), .Q(sreg[325]) );
  DFF \sreg_reg[326]  ( .D(swire[102]), .CLK(clk), .RST(rst), .Q(sreg[326]) );
  DFF \sreg_reg[327]  ( .D(swire[103]), .CLK(clk), .RST(rst), .Q(sreg[327]) );
  DFF \sreg_reg[328]  ( .D(swire[104]), .CLK(clk), .RST(rst), .Q(sreg[328]) );
  DFF \sreg_reg[329]  ( .D(swire[105]), .CLK(clk), .RST(rst), .Q(sreg[329]) );
  DFF \sreg_reg[330]  ( .D(swire[106]), .CLK(clk), .RST(rst), .Q(sreg[330]) );
  DFF \sreg_reg[331]  ( .D(swire[107]), .CLK(clk), .RST(rst), .Q(sreg[331]) );
  DFF \sreg_reg[332]  ( .D(swire[108]), .CLK(clk), .RST(rst), .Q(sreg[332]) );
  DFF \sreg_reg[333]  ( .D(swire[109]), .CLK(clk), .RST(rst), .Q(sreg[333]) );
  DFF \sreg_reg[334]  ( .D(swire[110]), .CLK(clk), .RST(rst), .Q(sreg[334]) );
  DFF \sreg_reg[335]  ( .D(swire[111]), .CLK(clk), .RST(rst), .Q(sreg[335]) );
  DFF \sreg_reg[336]  ( .D(swire[112]), .CLK(clk), .RST(rst), .Q(sreg[336]) );
  DFF \sreg_reg[337]  ( .D(swire[113]), .CLK(clk), .RST(rst), .Q(sreg[337]) );
  DFF \sreg_reg[338]  ( .D(swire[114]), .CLK(clk), .RST(rst), .Q(sreg[338]) );
  DFF \sreg_reg[339]  ( .D(swire[115]), .CLK(clk), .RST(rst), .Q(sreg[339]) );
  DFF \sreg_reg[340]  ( .D(swire[116]), .CLK(clk), .RST(rst), .Q(sreg[340]) );
  DFF \sreg_reg[341]  ( .D(swire[117]), .CLK(clk), .RST(rst), .Q(sreg[341]) );
  DFF \sreg_reg[342]  ( .D(swire[118]), .CLK(clk), .RST(rst), .Q(sreg[342]) );
  DFF \sreg_reg[343]  ( .D(swire[119]), .CLK(clk), .RST(rst), .Q(sreg[343]) );
  DFF \sreg_reg[344]  ( .D(swire[120]), .CLK(clk), .RST(rst), .Q(sreg[344]) );
  DFF \sreg_reg[345]  ( .D(swire[121]), .CLK(clk), .RST(rst), .Q(sreg[345]) );
  DFF \sreg_reg[346]  ( .D(swire[122]), .CLK(clk), .RST(rst), .Q(sreg[346]) );
  DFF \sreg_reg[347]  ( .D(swire[123]), .CLK(clk), .RST(rst), .Q(sreg[347]) );
  DFF \sreg_reg[348]  ( .D(swire[124]), .CLK(clk), .RST(rst), .Q(sreg[348]) );
  DFF \sreg_reg[349]  ( .D(swire[125]), .CLK(clk), .RST(rst), .Q(sreg[349]) );
  DFF \sreg_reg[350]  ( .D(swire[126]), .CLK(clk), .RST(rst), .Q(sreg[350]) );
  DFF \sreg_reg[351]  ( .D(swire[127]), .CLK(clk), .RST(rst), .Q(sreg[351]) );
  DFF \sreg_reg[352]  ( .D(swire[128]), .CLK(clk), .RST(rst), .Q(sreg[352]) );
  DFF \sreg_reg[353]  ( .D(swire[129]), .CLK(clk), .RST(rst), .Q(sreg[353]) );
  DFF \sreg_reg[354]  ( .D(swire[130]), .CLK(clk), .RST(rst), .Q(sreg[354]) );
  DFF \sreg_reg[355]  ( .D(swire[131]), .CLK(clk), .RST(rst), .Q(sreg[355]) );
  DFF \sreg_reg[356]  ( .D(swire[132]), .CLK(clk), .RST(rst), .Q(sreg[356]) );
  DFF \sreg_reg[357]  ( .D(swire[133]), .CLK(clk), .RST(rst), .Q(sreg[357]) );
  DFF \sreg_reg[358]  ( .D(swire[134]), .CLK(clk), .RST(rst), .Q(sreg[358]) );
  DFF \sreg_reg[359]  ( .D(swire[135]), .CLK(clk), .RST(rst), .Q(sreg[359]) );
  DFF \sreg_reg[360]  ( .D(swire[136]), .CLK(clk), .RST(rst), .Q(sreg[360]) );
  DFF \sreg_reg[361]  ( .D(swire[137]), .CLK(clk), .RST(rst), .Q(sreg[361]) );
  DFF \sreg_reg[362]  ( .D(swire[138]), .CLK(clk), .RST(rst), .Q(sreg[362]) );
  DFF \sreg_reg[363]  ( .D(swire[139]), .CLK(clk), .RST(rst), .Q(sreg[363]) );
  DFF \sreg_reg[364]  ( .D(swire[140]), .CLK(clk), .RST(rst), .Q(sreg[364]) );
  DFF \sreg_reg[365]  ( .D(swire[141]), .CLK(clk), .RST(rst), .Q(sreg[365]) );
  DFF \sreg_reg[366]  ( .D(swire[142]), .CLK(clk), .RST(rst), .Q(sreg[366]) );
  DFF \sreg_reg[367]  ( .D(swire[143]), .CLK(clk), .RST(rst), .Q(sreg[367]) );
  DFF \sreg_reg[368]  ( .D(swire[144]), .CLK(clk), .RST(rst), .Q(sreg[368]) );
  DFF \sreg_reg[369]  ( .D(swire[145]), .CLK(clk), .RST(rst), .Q(sreg[369]) );
  DFF \sreg_reg[370]  ( .D(swire[146]), .CLK(clk), .RST(rst), .Q(sreg[370]) );
  DFF \sreg_reg[371]  ( .D(swire[147]), .CLK(clk), .RST(rst), .Q(sreg[371]) );
  DFF \sreg_reg[372]  ( .D(swire[148]), .CLK(clk), .RST(rst), .Q(sreg[372]) );
  DFF \sreg_reg[373]  ( .D(swire[149]), .CLK(clk), .RST(rst), .Q(sreg[373]) );
  DFF \sreg_reg[374]  ( .D(swire[150]), .CLK(clk), .RST(rst), .Q(sreg[374]) );
  DFF \sreg_reg[375]  ( .D(swire[151]), .CLK(clk), .RST(rst), .Q(sreg[375]) );
  DFF \sreg_reg[376]  ( .D(swire[152]), .CLK(clk), .RST(rst), .Q(sreg[376]) );
  DFF \sreg_reg[377]  ( .D(swire[153]), .CLK(clk), .RST(rst), .Q(sreg[377]) );
  DFF \sreg_reg[378]  ( .D(swire[154]), .CLK(clk), .RST(rst), .Q(sreg[378]) );
  DFF \sreg_reg[379]  ( .D(swire[155]), .CLK(clk), .RST(rst), .Q(sreg[379]) );
  DFF \sreg_reg[380]  ( .D(swire[156]), .CLK(clk), .RST(rst), .Q(sreg[380]) );
  DFF \sreg_reg[381]  ( .D(swire[157]), .CLK(clk), .RST(rst), .Q(sreg[381]) );
  DFF \sreg_reg[382]  ( .D(swire[158]), .CLK(clk), .RST(rst), .Q(sreg[382]) );
  DFF \sreg_reg[383]  ( .D(swire[159]), .CLK(clk), .RST(rst), .Q(sreg[383]) );
  DFF \sreg_reg[384]  ( .D(swire[160]), .CLK(clk), .RST(rst), .Q(sreg[384]) );
  DFF \sreg_reg[385]  ( .D(swire[161]), .CLK(clk), .RST(rst), .Q(sreg[385]) );
  DFF \sreg_reg[386]  ( .D(swire[162]), .CLK(clk), .RST(rst), .Q(sreg[386]) );
  DFF \sreg_reg[387]  ( .D(swire[163]), .CLK(clk), .RST(rst), .Q(sreg[387]) );
  DFF \sreg_reg[388]  ( .D(swire[164]), .CLK(clk), .RST(rst), .Q(sreg[388]) );
  DFF \sreg_reg[389]  ( .D(swire[165]), .CLK(clk), .RST(rst), .Q(sreg[389]) );
  DFF \sreg_reg[390]  ( .D(swire[166]), .CLK(clk), .RST(rst), .Q(sreg[390]) );
  DFF \sreg_reg[391]  ( .D(swire[167]), .CLK(clk), .RST(rst), .Q(sreg[391]) );
  DFF \sreg_reg[392]  ( .D(swire[168]), .CLK(clk), .RST(rst), .Q(sreg[392]) );
  DFF \sreg_reg[393]  ( .D(swire[169]), .CLK(clk), .RST(rst), .Q(sreg[393]) );
  DFF \sreg_reg[394]  ( .D(swire[170]), .CLK(clk), .RST(rst), .Q(sreg[394]) );
  DFF \sreg_reg[395]  ( .D(swire[171]), .CLK(clk), .RST(rst), .Q(sreg[395]) );
  DFF \sreg_reg[396]  ( .D(swire[172]), .CLK(clk), .RST(rst), .Q(sreg[396]) );
  DFF \sreg_reg[397]  ( .D(swire[173]), .CLK(clk), .RST(rst), .Q(sreg[397]) );
  DFF \sreg_reg[398]  ( .D(swire[174]), .CLK(clk), .RST(rst), .Q(sreg[398]) );
  DFF \sreg_reg[399]  ( .D(swire[175]), .CLK(clk), .RST(rst), .Q(sreg[399]) );
  DFF \sreg_reg[400]  ( .D(swire[176]), .CLK(clk), .RST(rst), .Q(sreg[400]) );
  DFF \sreg_reg[401]  ( .D(swire[177]), .CLK(clk), .RST(rst), .Q(sreg[401]) );
  DFF \sreg_reg[402]  ( .D(swire[178]), .CLK(clk), .RST(rst), .Q(sreg[402]) );
  DFF \sreg_reg[403]  ( .D(swire[179]), .CLK(clk), .RST(rst), .Q(sreg[403]) );
  DFF \sreg_reg[404]  ( .D(swire[180]), .CLK(clk), .RST(rst), .Q(sreg[404]) );
  DFF \sreg_reg[405]  ( .D(swire[181]), .CLK(clk), .RST(rst), .Q(sreg[405]) );
  DFF \sreg_reg[406]  ( .D(swire[182]), .CLK(clk), .RST(rst), .Q(sreg[406]) );
  DFF \sreg_reg[407]  ( .D(swire[183]), .CLK(clk), .RST(rst), .Q(sreg[407]) );
  DFF \sreg_reg[408]  ( .D(swire[184]), .CLK(clk), .RST(rst), .Q(sreg[408]) );
  DFF \sreg_reg[409]  ( .D(swire[185]), .CLK(clk), .RST(rst), .Q(sreg[409]) );
  DFF \sreg_reg[410]  ( .D(swire[186]), .CLK(clk), .RST(rst), .Q(sreg[410]) );
  DFF \sreg_reg[411]  ( .D(swire[187]), .CLK(clk), .RST(rst), .Q(sreg[411]) );
  DFF \sreg_reg[412]  ( .D(swire[188]), .CLK(clk), .RST(rst), .Q(sreg[412]) );
  DFF \sreg_reg[413]  ( .D(swire[189]), .CLK(clk), .RST(rst), .Q(sreg[413]) );
  DFF \sreg_reg[414]  ( .D(swire[190]), .CLK(clk), .RST(rst), .Q(sreg[414]) );
  DFF \sreg_reg[415]  ( .D(swire[191]), .CLK(clk), .RST(rst), .Q(sreg[415]) );
  DFF \sreg_reg[416]  ( .D(swire[192]), .CLK(clk), .RST(rst), .Q(sreg[416]) );
  DFF \sreg_reg[417]  ( .D(swire[193]), .CLK(clk), .RST(rst), .Q(sreg[417]) );
  DFF \sreg_reg[418]  ( .D(swire[194]), .CLK(clk), .RST(rst), .Q(sreg[418]) );
  DFF \sreg_reg[419]  ( .D(swire[195]), .CLK(clk), .RST(rst), .Q(sreg[419]) );
  DFF \sreg_reg[420]  ( .D(swire[196]), .CLK(clk), .RST(rst), .Q(sreg[420]) );
  DFF \sreg_reg[421]  ( .D(swire[197]), .CLK(clk), .RST(rst), .Q(sreg[421]) );
  DFF \sreg_reg[422]  ( .D(swire[198]), .CLK(clk), .RST(rst), .Q(sreg[422]) );
  DFF \sreg_reg[423]  ( .D(swire[199]), .CLK(clk), .RST(rst), .Q(sreg[423]) );
  DFF \sreg_reg[424]  ( .D(swire[200]), .CLK(clk), .RST(rst), .Q(sreg[424]) );
  DFF \sreg_reg[425]  ( .D(swire[201]), .CLK(clk), .RST(rst), .Q(sreg[425]) );
  DFF \sreg_reg[426]  ( .D(swire[202]), .CLK(clk), .RST(rst), .Q(sreg[426]) );
  DFF \sreg_reg[427]  ( .D(swire[203]), .CLK(clk), .RST(rst), .Q(sreg[427]) );
  DFF \sreg_reg[428]  ( .D(swire[204]), .CLK(clk), .RST(rst), .Q(sreg[428]) );
  DFF \sreg_reg[429]  ( .D(swire[205]), .CLK(clk), .RST(rst), .Q(sreg[429]) );
  DFF \sreg_reg[430]  ( .D(swire[206]), .CLK(clk), .RST(rst), .Q(sreg[430]) );
  DFF \sreg_reg[431]  ( .D(swire[207]), .CLK(clk), .RST(rst), .Q(sreg[431]) );
  DFF \sreg_reg[432]  ( .D(swire[208]), .CLK(clk), .RST(rst), .Q(sreg[432]) );
  DFF \sreg_reg[433]  ( .D(swire[209]), .CLK(clk), .RST(rst), .Q(sreg[433]) );
  DFF \sreg_reg[434]  ( .D(swire[210]), .CLK(clk), .RST(rst), .Q(sreg[434]) );
  DFF \sreg_reg[435]  ( .D(swire[211]), .CLK(clk), .RST(rst), .Q(sreg[435]) );
  DFF \sreg_reg[436]  ( .D(swire[212]), .CLK(clk), .RST(rst), .Q(sreg[436]) );
  DFF \sreg_reg[437]  ( .D(swire[213]), .CLK(clk), .RST(rst), .Q(sreg[437]) );
  DFF \sreg_reg[438]  ( .D(swire[214]), .CLK(clk), .RST(rst), .Q(sreg[438]) );
  DFF \sreg_reg[439]  ( .D(swire[215]), .CLK(clk), .RST(rst), .Q(sreg[439]) );
  DFF \sreg_reg[440]  ( .D(swire[216]), .CLK(clk), .RST(rst), .Q(sreg[440]) );
  DFF \sreg_reg[441]  ( .D(swire[217]), .CLK(clk), .RST(rst), .Q(sreg[441]) );
  DFF \sreg_reg[442]  ( .D(swire[218]), .CLK(clk), .RST(rst), .Q(sreg[442]) );
  DFF \sreg_reg[443]  ( .D(swire[219]), .CLK(clk), .RST(rst), .Q(sreg[443]) );
  DFF \sreg_reg[444]  ( .D(swire[220]), .CLK(clk), .RST(rst), .Q(sreg[444]) );
  DFF \sreg_reg[445]  ( .D(swire[221]), .CLK(clk), .RST(rst), .Q(sreg[445]) );
  DFF \sreg_reg[446]  ( .D(swire[222]), .CLK(clk), .RST(rst), .Q(sreg[446]) );
  DFF \sreg_reg[447]  ( .D(swire[223]), .CLK(clk), .RST(rst), .Q(sreg[447]) );
  DFF \sreg_reg[448]  ( .D(swire[224]), .CLK(clk), .RST(rst), .Q(sreg[448]) );
  DFF \sreg_reg[449]  ( .D(swire[225]), .CLK(clk), .RST(rst), .Q(sreg[449]) );
  DFF \sreg_reg[450]  ( .D(swire[226]), .CLK(clk), .RST(rst), .Q(sreg[450]) );
  DFF \sreg_reg[451]  ( .D(swire[227]), .CLK(clk), .RST(rst), .Q(sreg[451]) );
  DFF \sreg_reg[452]  ( .D(swire[228]), .CLK(clk), .RST(rst), .Q(sreg[452]) );
  DFF \sreg_reg[453]  ( .D(swire[229]), .CLK(clk), .RST(rst), .Q(sreg[453]) );
  DFF \sreg_reg[454]  ( .D(swire[230]), .CLK(clk), .RST(rst), .Q(sreg[454]) );
  DFF \sreg_reg[455]  ( .D(swire[231]), .CLK(clk), .RST(rst), .Q(sreg[455]) );
  DFF \sreg_reg[456]  ( .D(swire[232]), .CLK(clk), .RST(rst), .Q(sreg[456]) );
  DFF \sreg_reg[457]  ( .D(swire[233]), .CLK(clk), .RST(rst), .Q(sreg[457]) );
  DFF \sreg_reg[458]  ( .D(swire[234]), .CLK(clk), .RST(rst), .Q(sreg[458]) );
  DFF \sreg_reg[459]  ( .D(swire[235]), .CLK(clk), .RST(rst), .Q(sreg[459]) );
  DFF \sreg_reg[460]  ( .D(swire[236]), .CLK(clk), .RST(rst), .Q(sreg[460]) );
  DFF \sreg_reg[461]  ( .D(swire[237]), .CLK(clk), .RST(rst), .Q(sreg[461]) );
  DFF \sreg_reg[462]  ( .D(swire[238]), .CLK(clk), .RST(rst), .Q(sreg[462]) );
  DFF \sreg_reg[463]  ( .D(swire[239]), .CLK(clk), .RST(rst), .Q(sreg[463]) );
  DFF \sreg_reg[464]  ( .D(swire[240]), .CLK(clk), .RST(rst), .Q(sreg[464]) );
  DFF \sreg_reg[465]  ( .D(swire[241]), .CLK(clk), .RST(rst), .Q(sreg[465]) );
  DFF \sreg_reg[466]  ( .D(swire[242]), .CLK(clk), .RST(rst), .Q(sreg[466]) );
  DFF \sreg_reg[467]  ( .D(swire[243]), .CLK(clk), .RST(rst), .Q(sreg[467]) );
  DFF \sreg_reg[468]  ( .D(swire[244]), .CLK(clk), .RST(rst), .Q(sreg[468]) );
  DFF \sreg_reg[469]  ( .D(swire[245]), .CLK(clk), .RST(rst), .Q(sreg[469]) );
  DFF \sreg_reg[470]  ( .D(swire[246]), .CLK(clk), .RST(rst), .Q(sreg[470]) );
  DFF \sreg_reg[471]  ( .D(swire[247]), .CLK(clk), .RST(rst), .Q(sreg[471]) );
  DFF \sreg_reg[472]  ( .D(swire[248]), .CLK(clk), .RST(rst), .Q(sreg[472]) );
  DFF \sreg_reg[473]  ( .D(swire[249]), .CLK(clk), .RST(rst), .Q(sreg[473]) );
  DFF \sreg_reg[474]  ( .D(swire[250]), .CLK(clk), .RST(rst), .Q(sreg[474]) );
  DFF \sreg_reg[475]  ( .D(swire[251]), .CLK(clk), .RST(rst), .Q(sreg[475]) );
  DFF \sreg_reg[476]  ( .D(swire[252]), .CLK(clk), .RST(rst), .Q(sreg[476]) );
  DFF \sreg_reg[477]  ( .D(swire[253]), .CLK(clk), .RST(rst), .Q(sreg[477]) );
  DFF \sreg_reg[478]  ( .D(swire[254]), .CLK(clk), .RST(rst), .Q(sreg[478]) );
  DFF \sreg_reg[479]  ( .D(swire[255]), .CLK(clk), .RST(rst), .Q(sreg[479]) );
  DFF \sreg_reg[255]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(c[223]) );
  DFF \sreg_reg[254]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(c[222]) );
  DFF \sreg_reg[253]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(c[221]) );
  DFF \sreg_reg[252]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(c[220]) );
  DFF \sreg_reg[251]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(c[219]) );
  DFF \sreg_reg[250]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(c[218]) );
  DFF \sreg_reg[249]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(c[217]) );
  DFF \sreg_reg[248]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(c[216]) );
  DFF \sreg_reg[247]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(c[215]) );
  DFF \sreg_reg[246]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(c[214]) );
  DFF \sreg_reg[245]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(c[213]) );
  DFF \sreg_reg[244]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(c[212]) );
  DFF \sreg_reg[243]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(c[211]) );
  DFF \sreg_reg[242]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(c[210]) );
  DFF \sreg_reg[241]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(c[209]) );
  DFF \sreg_reg[240]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(c[208]) );
  DFF \sreg_reg[239]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(c[207]) );
  DFF \sreg_reg[238]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(c[206]) );
  DFF \sreg_reg[237]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(c[205]) );
  DFF \sreg_reg[236]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(c[204]) );
  DFF \sreg_reg[235]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(c[203]) );
  DFF \sreg_reg[234]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(c[202]) );
  DFF \sreg_reg[233]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(c[201]) );
  DFF \sreg_reg[232]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(c[200]) );
  DFF \sreg_reg[231]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(c[199]) );
  DFF \sreg_reg[230]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(c[198]) );
  DFF \sreg_reg[229]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(c[197]) );
  DFF \sreg_reg[228]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(c[196]) );
  DFF \sreg_reg[227]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(c[195]) );
  DFF \sreg_reg[226]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(c[194]) );
  DFF \sreg_reg[225]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(c[193]) );
  DFF \sreg_reg[224]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(c[192]) );
  DFF \sreg_reg[223]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(c[191]) );
  DFF \sreg_reg[222]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(c[190]) );
  DFF \sreg_reg[221]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(c[189]) );
  DFF \sreg_reg[220]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(c[188]) );
  DFF \sreg_reg[219]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(c[187]) );
  DFF \sreg_reg[218]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(c[186]) );
  DFF \sreg_reg[217]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(c[185]) );
  DFF \sreg_reg[216]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(c[184]) );
  DFF \sreg_reg[215]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(c[183]) );
  DFF \sreg_reg[214]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(c[182]) );
  DFF \sreg_reg[213]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(c[181]) );
  DFF \sreg_reg[212]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(c[180]) );
  DFF \sreg_reg[211]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(c[179]) );
  DFF \sreg_reg[210]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(c[178]) );
  DFF \sreg_reg[209]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(c[177]) );
  DFF \sreg_reg[208]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(c[176]) );
  DFF \sreg_reg[207]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(c[175]) );
  DFF \sreg_reg[206]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(c[174]) );
  DFF \sreg_reg[205]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(c[173]) );
  DFF \sreg_reg[204]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(c[172]) );
  DFF \sreg_reg[203]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(c[171]) );
  DFF \sreg_reg[202]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(c[170]) );
  DFF \sreg_reg[201]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(c[169]) );
  DFF \sreg_reg[200]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(c[168]) );
  DFF \sreg_reg[199]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(c[167]) );
  DFF \sreg_reg[198]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(c[166]) );
  DFF \sreg_reg[197]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(c[165]) );
  DFF \sreg_reg[196]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(c[164]) );
  DFF \sreg_reg[195]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(c[163]) );
  DFF \sreg_reg[194]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(c[162]) );
  DFF \sreg_reg[193]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(c[161]) );
  DFF \sreg_reg[192]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(c[160]) );
  DFF \sreg_reg[191]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(c[159]) );
  DFF \sreg_reg[190]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(c[158]) );
  DFF \sreg_reg[189]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(c[157]) );
  DFF \sreg_reg[188]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(c[156]) );
  DFF \sreg_reg[187]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(c[155]) );
  DFF \sreg_reg[186]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(c[154]) );
  DFF \sreg_reg[185]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(c[153]) );
  DFF \sreg_reg[184]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(c[152]) );
  DFF \sreg_reg[183]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(c[151]) );
  DFF \sreg_reg[182]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(c[150]) );
  DFF \sreg_reg[181]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(c[149]) );
  DFF \sreg_reg[180]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(c[148]) );
  DFF \sreg_reg[179]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(c[147]) );
  DFF \sreg_reg[178]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(c[146]) );
  DFF \sreg_reg[177]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(c[145]) );
  DFF \sreg_reg[176]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(c[144]) );
  DFF \sreg_reg[175]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(c[143]) );
  DFF \sreg_reg[174]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(c[142]) );
  DFF \sreg_reg[173]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(c[141]) );
  DFF \sreg_reg[172]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(c[140]) );
  DFF \sreg_reg[171]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(c[139]) );
  DFF \sreg_reg[170]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(c[138]) );
  DFF \sreg_reg[169]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(c[137]) );
  DFF \sreg_reg[168]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(c[136]) );
  DFF \sreg_reg[167]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(c[135]) );
  DFF \sreg_reg[166]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(c[134]) );
  DFF \sreg_reg[165]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(c[133]) );
  DFF \sreg_reg[164]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(c[132]) );
  DFF \sreg_reg[163]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(c[131]) );
  DFF \sreg_reg[162]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(c[130]) );
  DFF \sreg_reg[161]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(c[129]) );
  DFF \sreg_reg[160]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(c[128]) );
  DFF \sreg_reg[159]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(c[127]) );
  DFF \sreg_reg[158]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(c[126]) );
  DFF \sreg_reg[157]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(c[125]) );
  DFF \sreg_reg[156]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(c[124]) );
  DFF \sreg_reg[155]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[154]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[153]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[152]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[151]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[150]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[149]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[148]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[147]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[146]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[145]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[144]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[143]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[142]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[141]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[140]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[139]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[138]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[137]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[136]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[135]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[134]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[133]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[132]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[131]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[130]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[129]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[128]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[127]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[126]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[125]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[124]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[123]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[122]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[121]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[120]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[119]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[118]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[117]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[116]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[115]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[114]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[113]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[112]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[111]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[110]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[109]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[108]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[107]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[106]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[105]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[104]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[103]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[102]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[101]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[100]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[99]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[98]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[97]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[96]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[95]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[94]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[93]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[92]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[91]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[90]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[89]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[88]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[87]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[86]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[85]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[84]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[83]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[82]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[81]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[80]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[79]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[78]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[77]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[76]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[75]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[74]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[73]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[72]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[71]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[70]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[69]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[68]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[67]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[66]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[65]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[64]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[0]) );
  ADD_N256_1 ADD_ ( .A({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        sreg[479:256]}), .B(clocal), .CI(1'b0), .S({swire, c[255:224]}) );
  mult_N256_CC8_DW02_mult_0 mult_44 ( .A(b), .B(a), .TC(1'b0), .PRODUCT({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, SYNOPSYS_UNCONNECTED__31, clocal}) );
endmodule

