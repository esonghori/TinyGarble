
module k_nns_seq_W15_K8 ( clk, rst, q, DB, min_val_out );
  input [14:0] q;
  input [14:0] DB;
  output [119:0] min_val_out;
  input clk, rst;
  wire   \min_dist_reg[7][3] , \min_dist_reg[7][2] , \min_dist_reg[7][1] ,
         \min_dist_reg[7][0] , \min_dist_reg[6][3] , \min_dist_reg[6][2] ,
         \min_dist_reg[6][1] , \min_dist_reg[6][0] , \min_dist_reg[5][3] ,
         \min_dist_reg[5][2] , \min_dist_reg[5][1] , \min_dist_reg[5][0] ,
         \min_dist_reg[4][3] , \min_dist_reg[4][2] , \min_dist_reg[4][1] ,
         \min_dist_reg[4][0] , \min_dist_reg[3][3] , \min_dist_reg[3][2] ,
         \min_dist_reg[3][1] , \min_dist_reg[3][0] , \min_dist_reg[2][3] ,
         \min_dist_reg[2][2] , \min_dist_reg[2][1] , \min_dist_reg[2][0] ,
         \min_dist_reg[1][3] , \min_dist_reg[1][2] , \min_dist_reg[1][1] ,
         \min_dist_reg[1][0] , \min_dist_reg[0][3] , \min_dist_reg[0][2] ,
         \min_dist_reg[0][1] , \min_dist_reg[0][0] , \local_min_dist[0][3] ,
         \local_min_dist[0][2] , \local_min_dist[0][1] ,
         \local_min_dist[0][0] , \min_dist[7][3] , \min_dist[7][2] ,
         \min_dist[7][1] , \min_dist[7][0] , \min_dist[6][3] ,
         \min_dist[6][2] , \min_dist[6][1] , \min_dist[6][0] ,
         \min_dist[5][3] , \min_dist[5][2] , \min_dist[5][1] ,
         \min_dist[5][0] , \min_dist[4][3] , \min_dist[4][2] ,
         \min_dist[4][1] , \min_dist[4][0] , \min_dist[3][3] ,
         \min_dist[3][2] , \min_dist[3][1] , \min_dist[3][0] ,
         \min_dist[2][3] , \min_dist[2][2] , \min_dist[2][1] ,
         \min_dist[2][0] , \min_dist[1][3] , \min_dist[1][2] ,
         \min_dist[1][1] , \min_dist[1][0] , \min_val_reg[7][14] ,
         \min_val_reg[7][13] , \min_val_reg[7][12] , \min_val_reg[7][11] ,
         \min_val_reg[7][10] , \min_val_reg[7][9] , \min_val_reg[7][8] ,
         \min_val_reg[7][7] , \min_val_reg[7][6] , \min_val_reg[7][5] ,
         \min_val_reg[7][4] , \min_val_reg[7][3] , \min_val_reg[7][2] ,
         \min_val_reg[7][1] , \min_val_reg[7][0] , \min_val_reg[6][14] ,
         \min_val_reg[6][13] , \min_val_reg[6][12] , \min_val_reg[6][11] ,
         \min_val_reg[6][10] , \min_val_reg[6][9] , \min_val_reg[6][8] ,
         \min_val_reg[6][7] , \min_val_reg[6][6] , \min_val_reg[6][5] ,
         \min_val_reg[6][4] , \min_val_reg[6][3] , \min_val_reg[6][2] ,
         \min_val_reg[6][1] , \min_val_reg[6][0] , \min_val_reg[5][14] ,
         \min_val_reg[5][13] , \min_val_reg[5][12] , \min_val_reg[5][11] ,
         \min_val_reg[5][10] , \min_val_reg[5][9] , \min_val_reg[5][8] ,
         \min_val_reg[5][7] , \min_val_reg[5][6] , \min_val_reg[5][5] ,
         \min_val_reg[5][4] , \min_val_reg[5][3] , \min_val_reg[5][2] ,
         \min_val_reg[5][1] , \min_val_reg[5][0] , \min_val_reg[4][14] ,
         \min_val_reg[4][13] , \min_val_reg[4][12] , \min_val_reg[4][11] ,
         \min_val_reg[4][10] , \min_val_reg[4][9] , \min_val_reg[4][8] ,
         \min_val_reg[4][7] , \min_val_reg[4][6] , \min_val_reg[4][5] ,
         \min_val_reg[4][4] , \min_val_reg[4][3] , \min_val_reg[4][2] ,
         \min_val_reg[4][1] , \min_val_reg[4][0] , \min_val_reg[3][14] ,
         \min_val_reg[3][13] , \min_val_reg[3][12] , \min_val_reg[3][11] ,
         \min_val_reg[3][10] , \min_val_reg[3][9] , \min_val_reg[3][8] ,
         \min_val_reg[3][7] , \min_val_reg[3][6] , \min_val_reg[3][5] ,
         \min_val_reg[3][4] , \min_val_reg[3][3] , \min_val_reg[3][2] ,
         \min_val_reg[3][1] , \min_val_reg[3][0] , \min_val_reg[2][14] ,
         \min_val_reg[2][13] , \min_val_reg[2][12] , \min_val_reg[2][11] ,
         \min_val_reg[2][10] , \min_val_reg[2][9] , \min_val_reg[2][8] ,
         \min_val_reg[2][7] , \min_val_reg[2][6] , \min_val_reg[2][5] ,
         \min_val_reg[2][4] , \min_val_reg[2][3] , \min_val_reg[2][2] ,
         \min_val_reg[2][1] , \min_val_reg[2][0] , \min_val_reg[1][14] ,
         \min_val_reg[1][13] , \min_val_reg[1][12] , \min_val_reg[1][11] ,
         \min_val_reg[1][10] , \min_val_reg[1][9] , \min_val_reg[1][8] ,
         \min_val_reg[1][7] , \min_val_reg[1][6] , \min_val_reg[1][5] ,
         \min_val_reg[1][4] , \min_val_reg[1][3] , \min_val_reg[1][2] ,
         \min_val_reg[1][1] , \min_val_reg[1][0] , \min_val_reg[0][14] ,
         \min_val_reg[0][13] , \min_val_reg[0][12] , \min_val_reg[0][11] ,
         \min_val_reg[0][10] , \min_val_reg[0][9] , \min_val_reg[0][8] ,
         \min_val_reg[0][7] , \min_val_reg[0][6] , \min_val_reg[0][5] ,
         \min_val_reg[0][4] , \min_val_reg[0][3] , \min_val_reg[0][2] ,
         \min_val_reg[0][1] , \min_val_reg[0][0] , n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963;

  DFF \min_dist_reg_reg[0][0]  ( .D(\local_min_dist[0][0] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][0] ) );
  DFF \min_dist_reg_reg[0][1]  ( .D(\local_min_dist[0][1] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][1] ) );
  DFF \min_dist_reg_reg[0][2]  ( .D(\local_min_dist[0][2] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][2] ) );
  DFF \min_dist_reg_reg[0][3]  ( .D(\local_min_dist[0][3] ), .CLK(clk), .RST(
        rst), .I(1'b1), .Q(\min_dist_reg[0][3] ) );
  DFF \min_dist_reg_reg[1][0]  ( .D(\min_dist[1][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][0] ) );
  DFF \min_dist_reg_reg[1][1]  ( .D(\min_dist[1][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][1] ) );
  DFF \min_dist_reg_reg[1][2]  ( .D(\min_dist[1][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][2] ) );
  DFF \min_dist_reg_reg[1][3]  ( .D(\min_dist[1][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[1][3] ) );
  DFF \min_dist_reg_reg[2][0]  ( .D(\min_dist[2][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][0] ) );
  DFF \min_dist_reg_reg[2][1]  ( .D(\min_dist[2][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][1] ) );
  DFF \min_dist_reg_reg[2][2]  ( .D(\min_dist[2][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][2] ) );
  DFF \min_dist_reg_reg[2][3]  ( .D(\min_dist[2][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[2][3] ) );
  DFF \min_dist_reg_reg[3][0]  ( .D(\min_dist[3][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][0] ) );
  DFF \min_dist_reg_reg[3][1]  ( .D(\min_dist[3][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][1] ) );
  DFF \min_dist_reg_reg[3][2]  ( .D(\min_dist[3][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][2] ) );
  DFF \min_dist_reg_reg[3][3]  ( .D(\min_dist[3][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[3][3] ) );
  DFF \min_dist_reg_reg[4][0]  ( .D(\min_dist[4][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[4][0] ) );
  DFF \min_dist_reg_reg[4][1]  ( .D(\min_dist[4][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[4][1] ) );
  DFF \min_dist_reg_reg[4][2]  ( .D(\min_dist[4][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[4][2] ) );
  DFF \min_dist_reg_reg[4][3]  ( .D(\min_dist[4][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[4][3] ) );
  DFF \min_dist_reg_reg[5][0]  ( .D(\min_dist[5][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[5][0] ) );
  DFF \min_dist_reg_reg[5][1]  ( .D(\min_dist[5][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[5][1] ) );
  DFF \min_dist_reg_reg[5][2]  ( .D(\min_dist[5][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[5][2] ) );
  DFF \min_dist_reg_reg[5][3]  ( .D(\min_dist[5][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[5][3] ) );
  DFF \min_dist_reg_reg[6][0]  ( .D(\min_dist[6][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[6][0] ) );
  DFF \min_dist_reg_reg[6][1]  ( .D(\min_dist[6][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[6][1] ) );
  DFF \min_dist_reg_reg[6][2]  ( .D(\min_dist[6][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[6][2] ) );
  DFF \min_dist_reg_reg[6][3]  ( .D(\min_dist[6][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[6][3] ) );
  DFF \min_dist_reg_reg[7][0]  ( .D(\min_dist[7][0] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[7][0] ) );
  DFF \min_dist_reg_reg[7][1]  ( .D(\min_dist[7][1] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[7][1] ) );
  DFF \min_dist_reg_reg[7][2]  ( .D(\min_dist[7][2] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[7][2] ) );
  DFF \min_dist_reg_reg[7][3]  ( .D(\min_dist[7][3] ), .CLK(clk), .RST(rst), 
        .I(1'b1), .Q(\min_dist_reg[7][3] ) );
  DFF \min_val_reg_reg[0][0]  ( .D(min_val_out[0]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][0] ) );
  DFF \min_val_reg_reg[0][1]  ( .D(min_val_out[1]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][1] ) );
  DFF \min_val_reg_reg[0][2]  ( .D(min_val_out[2]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][2] ) );
  DFF \min_val_reg_reg[0][3]  ( .D(min_val_out[3]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][3] ) );
  DFF \min_val_reg_reg[0][4]  ( .D(min_val_out[4]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][4] ) );
  DFF \min_val_reg_reg[0][5]  ( .D(min_val_out[5]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][5] ) );
  DFF \min_val_reg_reg[0][6]  ( .D(min_val_out[6]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][6] ) );
  DFF \min_val_reg_reg[0][7]  ( .D(min_val_out[7]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][7] ) );
  DFF \min_val_reg_reg[0][8]  ( .D(min_val_out[8]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][8] ) );
  DFF \min_val_reg_reg[0][9]  ( .D(min_val_out[9]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[0][9] ) );
  DFF \min_val_reg_reg[0][10]  ( .D(min_val_out[10]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][10] ) );
  DFF \min_val_reg_reg[0][11]  ( .D(min_val_out[11]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][11] ) );
  DFF \min_val_reg_reg[0][12]  ( .D(min_val_out[12]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][12] ) );
  DFF \min_val_reg_reg[0][13]  ( .D(min_val_out[13]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][13] ) );
  DFF \min_val_reg_reg[0][14]  ( .D(min_val_out[14]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[0][14] ) );
  DFF \min_val_reg_reg[1][0]  ( .D(min_val_out[15]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][0] ) );
  DFF \min_val_reg_reg[1][1]  ( .D(min_val_out[16]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][1] ) );
  DFF \min_val_reg_reg[1][2]  ( .D(min_val_out[17]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][2] ) );
  DFF \min_val_reg_reg[1][3]  ( .D(min_val_out[18]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][3] ) );
  DFF \min_val_reg_reg[1][4]  ( .D(min_val_out[19]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][4] ) );
  DFF \min_val_reg_reg[1][5]  ( .D(min_val_out[20]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][5] ) );
  DFF \min_val_reg_reg[1][6]  ( .D(min_val_out[21]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][6] ) );
  DFF \min_val_reg_reg[1][7]  ( .D(min_val_out[22]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][7] ) );
  DFF \min_val_reg_reg[1][8]  ( .D(min_val_out[23]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][8] ) );
  DFF \min_val_reg_reg[1][9]  ( .D(min_val_out[24]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[1][9] ) );
  DFF \min_val_reg_reg[1][10]  ( .D(min_val_out[25]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][10] ) );
  DFF \min_val_reg_reg[1][11]  ( .D(min_val_out[26]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][11] ) );
  DFF \min_val_reg_reg[1][12]  ( .D(min_val_out[27]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][12] ) );
  DFF \min_val_reg_reg[1][13]  ( .D(min_val_out[28]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][13] ) );
  DFF \min_val_reg_reg[1][14]  ( .D(min_val_out[29]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[1][14] ) );
  DFF \min_val_reg_reg[2][0]  ( .D(min_val_out[30]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][0] ) );
  DFF \min_val_reg_reg[2][1]  ( .D(min_val_out[31]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][1] ) );
  DFF \min_val_reg_reg[2][2]  ( .D(min_val_out[32]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][2] ) );
  DFF \min_val_reg_reg[2][3]  ( .D(min_val_out[33]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][3] ) );
  DFF \min_val_reg_reg[2][4]  ( .D(min_val_out[34]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][4] ) );
  DFF \min_val_reg_reg[2][5]  ( .D(min_val_out[35]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][5] ) );
  DFF \min_val_reg_reg[2][6]  ( .D(min_val_out[36]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][6] ) );
  DFF \min_val_reg_reg[2][7]  ( .D(min_val_out[37]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][7] ) );
  DFF \min_val_reg_reg[2][8]  ( .D(min_val_out[38]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][8] ) );
  DFF \min_val_reg_reg[2][9]  ( .D(min_val_out[39]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[2][9] ) );
  DFF \min_val_reg_reg[2][10]  ( .D(min_val_out[40]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][10] ) );
  DFF \min_val_reg_reg[2][11]  ( .D(min_val_out[41]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][11] ) );
  DFF \min_val_reg_reg[2][12]  ( .D(min_val_out[42]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][12] ) );
  DFF \min_val_reg_reg[2][13]  ( .D(min_val_out[43]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][13] ) );
  DFF \min_val_reg_reg[2][14]  ( .D(min_val_out[44]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[2][14] ) );
  DFF \min_val_reg_reg[3][0]  ( .D(min_val_out[45]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][0] ) );
  DFF \min_val_reg_reg[3][1]  ( .D(min_val_out[46]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][1] ) );
  DFF \min_val_reg_reg[3][2]  ( .D(min_val_out[47]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][2] ) );
  DFF \min_val_reg_reg[3][3]  ( .D(min_val_out[48]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][3] ) );
  DFF \min_val_reg_reg[3][4]  ( .D(min_val_out[49]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][4] ) );
  DFF \min_val_reg_reg[3][5]  ( .D(min_val_out[50]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][5] ) );
  DFF \min_val_reg_reg[3][6]  ( .D(min_val_out[51]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][6] ) );
  DFF \min_val_reg_reg[3][7]  ( .D(min_val_out[52]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][7] ) );
  DFF \min_val_reg_reg[3][8]  ( .D(min_val_out[53]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][8] ) );
  DFF \min_val_reg_reg[3][9]  ( .D(min_val_out[54]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[3][9] ) );
  DFF \min_val_reg_reg[3][10]  ( .D(min_val_out[55]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][10] ) );
  DFF \min_val_reg_reg[3][11]  ( .D(min_val_out[56]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][11] ) );
  DFF \min_val_reg_reg[3][12]  ( .D(min_val_out[57]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][12] ) );
  DFF \min_val_reg_reg[3][13]  ( .D(min_val_out[58]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][13] ) );
  DFF \min_val_reg_reg[3][14]  ( .D(min_val_out[59]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[3][14] ) );
  DFF \min_val_reg_reg[4][0]  ( .D(min_val_out[60]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[4][0] ) );
  DFF \min_val_reg_reg[4][1]  ( .D(min_val_out[61]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[4][1] ) );
  DFF \min_val_reg_reg[4][2]  ( .D(min_val_out[62]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[4][2] ) );
  DFF \min_val_reg_reg[4][3]  ( .D(min_val_out[63]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[4][3] ) );
  DFF \min_val_reg_reg[4][4]  ( .D(min_val_out[64]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[4][4] ) );
  DFF \min_val_reg_reg[4][5]  ( .D(min_val_out[65]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[4][5] ) );
  DFF \min_val_reg_reg[4][6]  ( .D(min_val_out[66]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[4][6] ) );
  DFF \min_val_reg_reg[4][7]  ( .D(min_val_out[67]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[4][7] ) );
  DFF \min_val_reg_reg[4][8]  ( .D(min_val_out[68]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[4][8] ) );
  DFF \min_val_reg_reg[4][9]  ( .D(min_val_out[69]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[4][9] ) );
  DFF \min_val_reg_reg[4][10]  ( .D(min_val_out[70]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][10] ) );
  DFF \min_val_reg_reg[4][11]  ( .D(min_val_out[71]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][11] ) );
  DFF \min_val_reg_reg[4][12]  ( .D(min_val_out[72]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][12] ) );
  DFF \min_val_reg_reg[4][13]  ( .D(min_val_out[73]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][13] ) );
  DFF \min_val_reg_reg[4][14]  ( .D(min_val_out[74]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[4][14] ) );
  DFF \min_val_reg_reg[5][0]  ( .D(min_val_out[75]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[5][0] ) );
  DFF \min_val_reg_reg[5][1]  ( .D(min_val_out[76]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[5][1] ) );
  DFF \min_val_reg_reg[5][2]  ( .D(min_val_out[77]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[5][2] ) );
  DFF \min_val_reg_reg[5][3]  ( .D(min_val_out[78]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[5][3] ) );
  DFF \min_val_reg_reg[5][4]  ( .D(min_val_out[79]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[5][4] ) );
  DFF \min_val_reg_reg[5][5]  ( .D(min_val_out[80]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[5][5] ) );
  DFF \min_val_reg_reg[5][6]  ( .D(min_val_out[81]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[5][6] ) );
  DFF \min_val_reg_reg[5][7]  ( .D(min_val_out[82]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[5][7] ) );
  DFF \min_val_reg_reg[5][8]  ( .D(min_val_out[83]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[5][8] ) );
  DFF \min_val_reg_reg[5][9]  ( .D(min_val_out[84]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[5][9] ) );
  DFF \min_val_reg_reg[5][10]  ( .D(min_val_out[85]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][10] ) );
  DFF \min_val_reg_reg[5][11]  ( .D(min_val_out[86]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][11] ) );
  DFF \min_val_reg_reg[5][12]  ( .D(min_val_out[87]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][12] ) );
  DFF \min_val_reg_reg[5][13]  ( .D(min_val_out[88]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][13] ) );
  DFF \min_val_reg_reg[5][14]  ( .D(min_val_out[89]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[5][14] ) );
  DFF \min_val_reg_reg[6][0]  ( .D(min_val_out[90]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[6][0] ) );
  DFF \min_val_reg_reg[6][1]  ( .D(min_val_out[91]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[6][1] ) );
  DFF \min_val_reg_reg[6][2]  ( .D(min_val_out[92]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[6][2] ) );
  DFF \min_val_reg_reg[6][3]  ( .D(min_val_out[93]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[6][3] ) );
  DFF \min_val_reg_reg[6][4]  ( .D(min_val_out[94]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[6][4] ) );
  DFF \min_val_reg_reg[6][5]  ( .D(min_val_out[95]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[6][5] ) );
  DFF \min_val_reg_reg[6][6]  ( .D(min_val_out[96]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[6][6] ) );
  DFF \min_val_reg_reg[6][7]  ( .D(min_val_out[97]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[6][7] ) );
  DFF \min_val_reg_reg[6][8]  ( .D(min_val_out[98]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[6][8] ) );
  DFF \min_val_reg_reg[6][9]  ( .D(min_val_out[99]), .CLK(clk), .RST(rst), .I(
        1'b0), .Q(\min_val_reg[6][9] ) );
  DFF \min_val_reg_reg[6][10]  ( .D(min_val_out[100]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][10] ) );
  DFF \min_val_reg_reg[6][11]  ( .D(min_val_out[101]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][11] ) );
  DFF \min_val_reg_reg[6][12]  ( .D(min_val_out[102]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][12] ) );
  DFF \min_val_reg_reg[6][13]  ( .D(min_val_out[103]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][13] ) );
  DFF \min_val_reg_reg[6][14]  ( .D(min_val_out[104]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[6][14] ) );
  DFF \min_val_reg_reg[7][0]  ( .D(min_val_out[105]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][0] ) );
  DFF \min_val_reg_reg[7][1]  ( .D(min_val_out[106]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][1] ) );
  DFF \min_val_reg_reg[7][2]  ( .D(min_val_out[107]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][2] ) );
  DFF \min_val_reg_reg[7][3]  ( .D(min_val_out[108]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][3] ) );
  DFF \min_val_reg_reg[7][4]  ( .D(min_val_out[109]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][4] ) );
  DFF \min_val_reg_reg[7][5]  ( .D(min_val_out[110]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][5] ) );
  DFF \min_val_reg_reg[7][6]  ( .D(min_val_out[111]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][6] ) );
  DFF \min_val_reg_reg[7][7]  ( .D(min_val_out[112]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][7] ) );
  DFF \min_val_reg_reg[7][8]  ( .D(min_val_out[113]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][8] ) );
  DFF \min_val_reg_reg[7][9]  ( .D(min_val_out[114]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][9] ) );
  DFF \min_val_reg_reg[7][10]  ( .D(min_val_out[115]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][10] ) );
  DFF \min_val_reg_reg[7][11]  ( .D(min_val_out[116]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][11] ) );
  DFF \min_val_reg_reg[7][12]  ( .D(min_val_out[117]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][12] ) );
  DFF \min_val_reg_reg[7][13]  ( .D(min_val_out[118]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][13] ) );
  DFF \min_val_reg_reg[7][14]  ( .D(min_val_out[119]), .CLK(clk), .RST(rst), 
        .I(1'b0), .Q(\min_val_reg[7][14] ) );
  XOR U170 ( .A(\min_val_reg[0][9] ), .B(n153), .Z(min_val_out[9]) );
  AND U171 ( .A(n154), .B(n155), .Z(n153) );
  XOR U172 ( .A(n156), .B(n157), .Z(min_val_out[99]) );
  AND U173 ( .A(n158), .B(n159), .Z(n156) );
  XOR U174 ( .A(n160), .B(n161), .Z(min_val_out[98]) );
  AND U175 ( .A(n158), .B(n162), .Z(n160) );
  XOR U176 ( .A(n163), .B(n164), .Z(min_val_out[97]) );
  AND U177 ( .A(n158), .B(n165), .Z(n163) );
  XOR U178 ( .A(n166), .B(n167), .Z(min_val_out[96]) );
  AND U179 ( .A(n158), .B(n168), .Z(n166) );
  XOR U180 ( .A(n169), .B(n170), .Z(min_val_out[95]) );
  AND U181 ( .A(n158), .B(n171), .Z(n169) );
  XOR U182 ( .A(n172), .B(n173), .Z(min_val_out[94]) );
  AND U183 ( .A(n158), .B(n174), .Z(n172) );
  XOR U184 ( .A(n175), .B(n176), .Z(min_val_out[93]) );
  AND U185 ( .A(n158), .B(n177), .Z(n175) );
  XOR U186 ( .A(n178), .B(n179), .Z(min_val_out[92]) );
  AND U187 ( .A(n158), .B(n180), .Z(n178) );
  XOR U188 ( .A(n181), .B(n182), .Z(min_val_out[91]) );
  AND U189 ( .A(n158), .B(n183), .Z(n181) );
  XOR U190 ( .A(n184), .B(n185), .Z(min_val_out[90]) );
  AND U191 ( .A(n158), .B(n186), .Z(n184) );
  XOR U192 ( .A(\min_val_reg[0][8] ), .B(n187), .Z(min_val_out[8]) );
  AND U193 ( .A(n154), .B(n188), .Z(n187) );
  XOR U194 ( .A(n189), .B(n190), .Z(min_val_out[89]) );
  AND U195 ( .A(n191), .B(n192), .Z(n189) );
  XOR U196 ( .A(n193), .B(n194), .Z(min_val_out[88]) );
  AND U197 ( .A(n191), .B(n195), .Z(n193) );
  XOR U198 ( .A(n196), .B(n197), .Z(min_val_out[87]) );
  AND U199 ( .A(n191), .B(n198), .Z(n196) );
  XOR U200 ( .A(n199), .B(n200), .Z(min_val_out[86]) );
  AND U201 ( .A(n191), .B(n201), .Z(n199) );
  XOR U202 ( .A(n202), .B(n203), .Z(min_val_out[85]) );
  AND U203 ( .A(n191), .B(n204), .Z(n202) );
  XOR U204 ( .A(n205), .B(n206), .Z(min_val_out[84]) );
  AND U205 ( .A(n191), .B(n207), .Z(n205) );
  XNOR U206 ( .A(n208), .B(n209), .Z(min_val_out[83]) );
  AND U207 ( .A(n191), .B(n210), .Z(n208) );
  XNOR U208 ( .A(n211), .B(n212), .Z(min_val_out[82]) );
  AND U209 ( .A(n191), .B(n213), .Z(n211) );
  XNOR U210 ( .A(n214), .B(n215), .Z(min_val_out[81]) );
  AND U211 ( .A(n191), .B(n216), .Z(n214) );
  XNOR U212 ( .A(n217), .B(n218), .Z(min_val_out[80]) );
  AND U213 ( .A(n191), .B(n219), .Z(n217) );
  XOR U214 ( .A(\min_val_reg[0][7] ), .B(n220), .Z(min_val_out[7]) );
  AND U215 ( .A(n154), .B(n221), .Z(n220) );
  XNOR U216 ( .A(n222), .B(n223), .Z(min_val_out[79]) );
  AND U217 ( .A(n191), .B(n224), .Z(n222) );
  XNOR U218 ( .A(n225), .B(n226), .Z(min_val_out[78]) );
  AND U219 ( .A(n191), .B(n227), .Z(n225) );
  XNOR U220 ( .A(n228), .B(n229), .Z(min_val_out[77]) );
  AND U221 ( .A(n191), .B(n230), .Z(n228) );
  XNOR U222 ( .A(n231), .B(n232), .Z(min_val_out[76]) );
  AND U223 ( .A(n191), .B(n233), .Z(n231) );
  XNOR U224 ( .A(n234), .B(n235), .Z(min_val_out[75]) );
  AND U225 ( .A(n191), .B(n236), .Z(n234) );
  XNOR U226 ( .A(n237), .B(n238), .Z(min_val_out[74]) );
  AND U227 ( .A(n239), .B(n240), .Z(n237) );
  XNOR U228 ( .A(n241), .B(n242), .Z(min_val_out[73]) );
  AND U229 ( .A(n239), .B(n243), .Z(n241) );
  XNOR U230 ( .A(n244), .B(n245), .Z(min_val_out[72]) );
  AND U231 ( .A(n239), .B(n246), .Z(n244) );
  XNOR U232 ( .A(n247), .B(n248), .Z(min_val_out[71]) );
  AND U233 ( .A(n239), .B(n249), .Z(n247) );
  XNOR U234 ( .A(n250), .B(n251), .Z(min_val_out[70]) );
  AND U235 ( .A(n239), .B(n252), .Z(n250) );
  XOR U236 ( .A(\min_val_reg[0][6] ), .B(n253), .Z(min_val_out[6]) );
  AND U237 ( .A(n154), .B(n254), .Z(n253) );
  XOR U238 ( .A(n255), .B(n256), .Z(min_val_out[69]) );
  AND U239 ( .A(n239), .B(n257), .Z(n255) );
  XOR U240 ( .A(n258), .B(n259), .Z(min_val_out[68]) );
  AND U241 ( .A(n239), .B(n260), .Z(n258) );
  XNOR U242 ( .A(n261), .B(n262), .Z(min_val_out[67]) );
  AND U243 ( .A(n239), .B(n263), .Z(n261) );
  XNOR U244 ( .A(n264), .B(n265), .Z(min_val_out[66]) );
  AND U245 ( .A(n239), .B(n266), .Z(n264) );
  XNOR U246 ( .A(n267), .B(n268), .Z(min_val_out[65]) );
  AND U247 ( .A(n239), .B(n269), .Z(n267) );
  XNOR U248 ( .A(n270), .B(n271), .Z(min_val_out[64]) );
  AND U249 ( .A(n239), .B(n272), .Z(n270) );
  XNOR U250 ( .A(n273), .B(n274), .Z(min_val_out[63]) );
  AND U251 ( .A(n239), .B(n275), .Z(n273) );
  XNOR U252 ( .A(n276), .B(n277), .Z(min_val_out[62]) );
  AND U253 ( .A(n239), .B(n278), .Z(n276) );
  XNOR U254 ( .A(n279), .B(n280), .Z(min_val_out[61]) );
  AND U255 ( .A(n239), .B(n281), .Z(n279) );
  XNOR U256 ( .A(n282), .B(n283), .Z(min_val_out[60]) );
  AND U257 ( .A(n239), .B(n284), .Z(n282) );
  XOR U258 ( .A(\min_val_reg[0][5] ), .B(n285), .Z(min_val_out[5]) );
  AND U259 ( .A(n154), .B(n286), .Z(n285) );
  XNOR U260 ( .A(n287), .B(n288), .Z(min_val_out[59]) );
  AND U261 ( .A(n289), .B(n290), .Z(n287) );
  XNOR U262 ( .A(n291), .B(n292), .Z(min_val_out[58]) );
  AND U263 ( .A(n289), .B(n293), .Z(n291) );
  XNOR U264 ( .A(n294), .B(n295), .Z(min_val_out[57]) );
  AND U265 ( .A(n289), .B(n296), .Z(n294) );
  XNOR U266 ( .A(n297), .B(n298), .Z(min_val_out[56]) );
  AND U267 ( .A(n289), .B(n299), .Z(n297) );
  XNOR U268 ( .A(n300), .B(n301), .Z(min_val_out[55]) );
  AND U269 ( .A(n289), .B(n302), .Z(n300) );
  XOR U270 ( .A(n303), .B(n304), .Z(min_val_out[54]) );
  AND U271 ( .A(n289), .B(n305), .Z(n303) );
  XOR U272 ( .A(n306), .B(n307), .Z(min_val_out[53]) );
  AND U273 ( .A(n289), .B(n308), .Z(n306) );
  XOR U274 ( .A(n309), .B(n310), .Z(min_val_out[52]) );
  AND U275 ( .A(n289), .B(n311), .Z(n309) );
  XOR U276 ( .A(n312), .B(n313), .Z(min_val_out[51]) );
  AND U277 ( .A(n289), .B(n314), .Z(n312) );
  XNOR U278 ( .A(n315), .B(n316), .Z(min_val_out[50]) );
  AND U279 ( .A(n289), .B(n317), .Z(n315) );
  XOR U280 ( .A(\min_val_reg[0][4] ), .B(n318), .Z(min_val_out[4]) );
  AND U281 ( .A(n154), .B(n319), .Z(n318) );
  XNOR U282 ( .A(n320), .B(n321), .Z(min_val_out[49]) );
  AND U283 ( .A(n289), .B(n322), .Z(n320) );
  XNOR U284 ( .A(n323), .B(n324), .Z(min_val_out[48]) );
  AND U285 ( .A(n289), .B(n325), .Z(n323) );
  XNOR U286 ( .A(n326), .B(n327), .Z(min_val_out[47]) );
  AND U287 ( .A(n289), .B(n328), .Z(n326) );
  XNOR U288 ( .A(n329), .B(n330), .Z(min_val_out[46]) );
  AND U289 ( .A(n289), .B(n331), .Z(n329) );
  XNOR U290 ( .A(n332), .B(n333), .Z(min_val_out[45]) );
  AND U291 ( .A(n289), .B(n334), .Z(n332) );
  XNOR U292 ( .A(n335), .B(n336), .Z(min_val_out[44]) );
  AND U293 ( .A(n337), .B(n338), .Z(n335) );
  XNOR U294 ( .A(n339), .B(n340), .Z(min_val_out[43]) );
  AND U295 ( .A(n337), .B(n341), .Z(n339) );
  XNOR U296 ( .A(n342), .B(n343), .Z(min_val_out[42]) );
  AND U297 ( .A(n337), .B(n344), .Z(n342) );
  XNOR U298 ( .A(n345), .B(n346), .Z(min_val_out[41]) );
  AND U299 ( .A(n337), .B(n347), .Z(n345) );
  XNOR U300 ( .A(n348), .B(n349), .Z(min_val_out[40]) );
  AND U301 ( .A(n337), .B(n350), .Z(n348) );
  XOR U302 ( .A(\min_val_reg[0][3] ), .B(n351), .Z(min_val_out[3]) );
  AND U303 ( .A(n154), .B(n352), .Z(n351) );
  XOR U304 ( .A(n353), .B(n354), .Z(min_val_out[39]) );
  AND U305 ( .A(n337), .B(n355), .Z(n353) );
  XOR U306 ( .A(n356), .B(n357), .Z(min_val_out[38]) );
  AND U307 ( .A(n337), .B(n358), .Z(n356) );
  XOR U308 ( .A(n359), .B(n360), .Z(min_val_out[37]) );
  AND U309 ( .A(n337), .B(n361), .Z(n359) );
  XOR U310 ( .A(n362), .B(n363), .Z(min_val_out[36]) );
  AND U311 ( .A(n337), .B(n364), .Z(n362) );
  XOR U312 ( .A(n365), .B(n366), .Z(min_val_out[35]) );
  AND U313 ( .A(n337), .B(n367), .Z(n365) );
  XOR U314 ( .A(n368), .B(n369), .Z(min_val_out[34]) );
  AND U315 ( .A(n337), .B(n370), .Z(n368) );
  XNOR U316 ( .A(n371), .B(n372), .Z(min_val_out[33]) );
  AND U317 ( .A(n337), .B(n373), .Z(n371) );
  XNOR U318 ( .A(n374), .B(n375), .Z(min_val_out[32]) );
  AND U319 ( .A(n337), .B(n376), .Z(n374) );
  XNOR U320 ( .A(n377), .B(n378), .Z(min_val_out[31]) );
  AND U321 ( .A(n337), .B(n379), .Z(n377) );
  XNOR U322 ( .A(n380), .B(n381), .Z(min_val_out[30]) );
  AND U323 ( .A(n337), .B(n382), .Z(n380) );
  XOR U324 ( .A(\min_val_reg[0][2] ), .B(n383), .Z(min_val_out[2]) );
  AND U325 ( .A(n154), .B(n384), .Z(n383) );
  XNOR U326 ( .A(n385), .B(n386), .Z(min_val_out[29]) );
  AND U327 ( .A(n387), .B(n388), .Z(n385) );
  XNOR U328 ( .A(n389), .B(n390), .Z(min_val_out[28]) );
  AND U329 ( .A(n387), .B(n391), .Z(n389) );
  XNOR U330 ( .A(n392), .B(n393), .Z(min_val_out[27]) );
  AND U331 ( .A(n387), .B(n394), .Z(n392) );
  XNOR U332 ( .A(n395), .B(n396), .Z(min_val_out[26]) );
  AND U333 ( .A(n387), .B(n397), .Z(n395) );
  XNOR U334 ( .A(n398), .B(n399), .Z(min_val_out[25]) );
  AND U335 ( .A(n387), .B(n400), .Z(n398) );
  XOR U336 ( .A(n401), .B(n402), .Z(min_val_out[24]) );
  AND U337 ( .A(n387), .B(n155), .Z(n401) );
  XOR U338 ( .A(\min_val_reg[0][9] ), .B(n402), .Z(n155) );
  XNOR U339 ( .A(\min_val_reg[1][9] ), .B(n403), .Z(n402) );
  NAND U340 ( .A(n355), .B(n337), .Z(n403) );
  XOR U341 ( .A(\min_val_reg[1][9] ), .B(n354), .Z(n355) );
  XNOR U342 ( .A(\min_val_reg[2][9] ), .B(n404), .Z(n354) );
  NAND U343 ( .A(n305), .B(n289), .Z(n404) );
  XOR U344 ( .A(\min_val_reg[2][9] ), .B(n304), .Z(n305) );
  XNOR U345 ( .A(\min_val_reg[3][9] ), .B(n405), .Z(n304) );
  NAND U346 ( .A(n257), .B(n239), .Z(n405) );
  XOR U347 ( .A(\min_val_reg[3][9] ), .B(n256), .Z(n257) );
  XNOR U348 ( .A(\min_val_reg[4][9] ), .B(n406), .Z(n256) );
  NAND U349 ( .A(n207), .B(n191), .Z(n406) );
  XOR U350 ( .A(\min_val_reg[4][9] ), .B(n206), .Z(n207) );
  XNOR U351 ( .A(\min_val_reg[5][9] ), .B(n407), .Z(n206) );
  NAND U352 ( .A(n159), .B(n158), .Z(n407) );
  XOR U353 ( .A(\min_val_reg[5][9] ), .B(n157), .Z(n159) );
  XNOR U354 ( .A(\min_val_reg[6][9] ), .B(n408), .Z(n157) );
  NAND U355 ( .A(n409), .B(n410), .Z(n408) );
  XOR U356 ( .A(n411), .B(n412), .Z(min_val_out[23]) );
  AND U357 ( .A(n387), .B(n188), .Z(n411) );
  XOR U358 ( .A(\min_val_reg[0][8] ), .B(n412), .Z(n188) );
  XNOR U359 ( .A(\min_val_reg[1][8] ), .B(n413), .Z(n412) );
  NAND U360 ( .A(n358), .B(n337), .Z(n413) );
  XOR U361 ( .A(\min_val_reg[1][8] ), .B(n357), .Z(n358) );
  XNOR U362 ( .A(\min_val_reg[2][8] ), .B(n414), .Z(n357) );
  NAND U363 ( .A(n308), .B(n289), .Z(n414) );
  XOR U364 ( .A(\min_val_reg[2][8] ), .B(n307), .Z(n308) );
  XNOR U365 ( .A(\min_val_reg[3][8] ), .B(n415), .Z(n307) );
  NAND U366 ( .A(n260), .B(n239), .Z(n415) );
  XOR U367 ( .A(\min_val_reg[3][8] ), .B(n259), .Z(n260) );
  XNOR U368 ( .A(\min_val_reg[4][8] ), .B(n416), .Z(n259) );
  NAND U369 ( .A(n210), .B(n191), .Z(n416) );
  XNOR U370 ( .A(\min_val_reg[4][8] ), .B(n209), .Z(n210) );
  XOR U371 ( .A(\min_val_reg[5][8] ), .B(n417), .Z(n209) );
  NAND U372 ( .A(n162), .B(n158), .Z(n417) );
  XOR U373 ( .A(\min_val_reg[5][8] ), .B(n161), .Z(n162) );
  XNOR U374 ( .A(\min_val_reg[6][8] ), .B(n418), .Z(n161) );
  NAND U375 ( .A(n419), .B(n410), .Z(n418) );
  XOR U376 ( .A(n420), .B(n421), .Z(min_val_out[22]) );
  AND U377 ( .A(n387), .B(n221), .Z(n420) );
  XOR U378 ( .A(\min_val_reg[0][7] ), .B(n421), .Z(n221) );
  XNOR U379 ( .A(\min_val_reg[1][7] ), .B(n422), .Z(n421) );
  NAND U380 ( .A(n361), .B(n337), .Z(n422) );
  XOR U381 ( .A(\min_val_reg[1][7] ), .B(n360), .Z(n361) );
  XNOR U382 ( .A(\min_val_reg[2][7] ), .B(n423), .Z(n360) );
  NAND U383 ( .A(n311), .B(n289), .Z(n423) );
  XOR U384 ( .A(\min_val_reg[2][7] ), .B(n310), .Z(n311) );
  XNOR U385 ( .A(\min_val_reg[3][7] ), .B(n424), .Z(n310) );
  NAND U386 ( .A(n263), .B(n239), .Z(n424) );
  XNOR U387 ( .A(\min_val_reg[3][7] ), .B(n262), .Z(n263) );
  XOR U388 ( .A(\min_val_reg[4][7] ), .B(n425), .Z(n262) );
  NAND U389 ( .A(n213), .B(n191), .Z(n425) );
  XNOR U390 ( .A(\min_val_reg[4][7] ), .B(n212), .Z(n213) );
  XOR U391 ( .A(\min_val_reg[5][7] ), .B(n426), .Z(n212) );
  NAND U392 ( .A(n165), .B(n158), .Z(n426) );
  XOR U393 ( .A(\min_val_reg[5][7] ), .B(n164), .Z(n165) );
  XNOR U394 ( .A(\min_val_reg[6][7] ), .B(n427), .Z(n164) );
  NAND U395 ( .A(n428), .B(n410), .Z(n427) );
  XOR U396 ( .A(n429), .B(n430), .Z(min_val_out[21]) );
  AND U397 ( .A(n387), .B(n254), .Z(n429) );
  XOR U398 ( .A(\min_val_reg[0][6] ), .B(n430), .Z(n254) );
  XNOR U399 ( .A(\min_val_reg[1][6] ), .B(n431), .Z(n430) );
  NAND U400 ( .A(n364), .B(n337), .Z(n431) );
  XOR U401 ( .A(\min_val_reg[1][6] ), .B(n363), .Z(n364) );
  XNOR U402 ( .A(\min_val_reg[2][6] ), .B(n432), .Z(n363) );
  NAND U403 ( .A(n314), .B(n289), .Z(n432) );
  XOR U404 ( .A(\min_val_reg[2][6] ), .B(n313), .Z(n314) );
  XNOR U405 ( .A(\min_val_reg[3][6] ), .B(n433), .Z(n313) );
  NAND U406 ( .A(n266), .B(n239), .Z(n433) );
  XNOR U407 ( .A(\min_val_reg[3][6] ), .B(n265), .Z(n266) );
  XOR U408 ( .A(\min_val_reg[4][6] ), .B(n434), .Z(n265) );
  NAND U409 ( .A(n216), .B(n191), .Z(n434) );
  XNOR U410 ( .A(\min_val_reg[4][6] ), .B(n215), .Z(n216) );
  XOR U411 ( .A(\min_val_reg[5][6] ), .B(n435), .Z(n215) );
  NAND U412 ( .A(n168), .B(n158), .Z(n435) );
  XOR U413 ( .A(\min_val_reg[5][6] ), .B(n167), .Z(n168) );
  XNOR U414 ( .A(\min_val_reg[6][6] ), .B(n436), .Z(n167) );
  NAND U415 ( .A(n437), .B(n410), .Z(n436) );
  XOR U416 ( .A(n438), .B(n439), .Z(min_val_out[20]) );
  AND U417 ( .A(n387), .B(n286), .Z(n438) );
  XOR U418 ( .A(\min_val_reg[0][5] ), .B(n439), .Z(n286) );
  XNOR U419 ( .A(\min_val_reg[1][5] ), .B(n440), .Z(n439) );
  NAND U420 ( .A(n367), .B(n337), .Z(n440) );
  XOR U421 ( .A(\min_val_reg[1][5] ), .B(n366), .Z(n367) );
  XNOR U422 ( .A(\min_val_reg[2][5] ), .B(n441), .Z(n366) );
  NAND U423 ( .A(n317), .B(n289), .Z(n441) );
  XNOR U424 ( .A(\min_val_reg[2][5] ), .B(n316), .Z(n317) );
  XOR U425 ( .A(\min_val_reg[3][5] ), .B(n442), .Z(n316) );
  NAND U426 ( .A(n269), .B(n239), .Z(n442) );
  XNOR U427 ( .A(\min_val_reg[3][5] ), .B(n268), .Z(n269) );
  XOR U428 ( .A(\min_val_reg[4][5] ), .B(n443), .Z(n268) );
  NAND U429 ( .A(n219), .B(n191), .Z(n443) );
  XNOR U430 ( .A(\min_val_reg[4][5] ), .B(n218), .Z(n219) );
  XOR U431 ( .A(\min_val_reg[5][5] ), .B(n444), .Z(n218) );
  NAND U432 ( .A(n171), .B(n158), .Z(n444) );
  XOR U433 ( .A(\min_val_reg[5][5] ), .B(n170), .Z(n171) );
  XNOR U434 ( .A(\min_val_reg[6][5] ), .B(n445), .Z(n170) );
  NAND U435 ( .A(n446), .B(n410), .Z(n445) );
  XOR U436 ( .A(\min_val_reg[0][1] ), .B(n447), .Z(min_val_out[1]) );
  AND U437 ( .A(n154), .B(n448), .Z(n447) );
  XOR U438 ( .A(n449), .B(n450), .Z(min_val_out[19]) );
  AND U439 ( .A(n387), .B(n319), .Z(n449) );
  XOR U440 ( .A(\min_val_reg[0][4] ), .B(n450), .Z(n319) );
  XNOR U441 ( .A(\min_val_reg[1][4] ), .B(n451), .Z(n450) );
  NAND U442 ( .A(n370), .B(n337), .Z(n451) );
  XOR U443 ( .A(\min_val_reg[1][4] ), .B(n369), .Z(n370) );
  XNOR U444 ( .A(\min_val_reg[2][4] ), .B(n452), .Z(n369) );
  NAND U445 ( .A(n322), .B(n289), .Z(n452) );
  XNOR U446 ( .A(\min_val_reg[2][4] ), .B(n321), .Z(n322) );
  XOR U447 ( .A(\min_val_reg[3][4] ), .B(n453), .Z(n321) );
  NAND U448 ( .A(n272), .B(n239), .Z(n453) );
  XNOR U449 ( .A(\min_val_reg[3][4] ), .B(n271), .Z(n272) );
  XOR U450 ( .A(\min_val_reg[4][4] ), .B(n454), .Z(n271) );
  NAND U451 ( .A(n224), .B(n191), .Z(n454) );
  XNOR U452 ( .A(\min_val_reg[4][4] ), .B(n223), .Z(n224) );
  XOR U453 ( .A(\min_val_reg[5][4] ), .B(n455), .Z(n223) );
  NAND U454 ( .A(n174), .B(n158), .Z(n455) );
  XOR U455 ( .A(\min_val_reg[5][4] ), .B(n173), .Z(n174) );
  XNOR U456 ( .A(\min_val_reg[6][4] ), .B(n456), .Z(n173) );
  NAND U457 ( .A(n457), .B(n410), .Z(n456) );
  XOR U458 ( .A(n458), .B(n459), .Z(min_val_out[18]) );
  AND U459 ( .A(n387), .B(n352), .Z(n458) );
  XOR U460 ( .A(\min_val_reg[0][3] ), .B(n459), .Z(n352) );
  XNOR U461 ( .A(\min_val_reg[1][3] ), .B(n460), .Z(n459) );
  NAND U462 ( .A(n373), .B(n337), .Z(n460) );
  XNOR U463 ( .A(\min_val_reg[1][3] ), .B(n372), .Z(n373) );
  XOR U464 ( .A(\min_val_reg[2][3] ), .B(n461), .Z(n372) );
  NAND U465 ( .A(n325), .B(n289), .Z(n461) );
  XNOR U466 ( .A(\min_val_reg[2][3] ), .B(n324), .Z(n325) );
  XOR U467 ( .A(\min_val_reg[3][3] ), .B(n462), .Z(n324) );
  NAND U468 ( .A(n275), .B(n239), .Z(n462) );
  XNOR U469 ( .A(\min_val_reg[3][3] ), .B(n274), .Z(n275) );
  XOR U470 ( .A(\min_val_reg[4][3] ), .B(n463), .Z(n274) );
  NAND U471 ( .A(n227), .B(n191), .Z(n463) );
  XNOR U472 ( .A(\min_val_reg[4][3] ), .B(n226), .Z(n227) );
  XOR U473 ( .A(\min_val_reg[5][3] ), .B(n464), .Z(n226) );
  NAND U474 ( .A(n177), .B(n158), .Z(n464) );
  XOR U475 ( .A(\min_val_reg[5][3] ), .B(n176), .Z(n177) );
  XNOR U476 ( .A(\min_val_reg[6][3] ), .B(n465), .Z(n176) );
  NAND U477 ( .A(n466), .B(n410), .Z(n465) );
  XNOR U478 ( .A(n467), .B(n468), .Z(min_val_out[17]) );
  AND U479 ( .A(n387), .B(n384), .Z(n467) );
  XNOR U480 ( .A(\min_val_reg[0][2] ), .B(n468), .Z(n384) );
  XOR U481 ( .A(\min_val_reg[1][2] ), .B(n469), .Z(n468) );
  NAND U482 ( .A(n376), .B(n337), .Z(n469) );
  XNOR U483 ( .A(\min_val_reg[1][2] ), .B(n375), .Z(n376) );
  XOR U484 ( .A(\min_val_reg[2][2] ), .B(n470), .Z(n375) );
  NAND U485 ( .A(n328), .B(n289), .Z(n470) );
  XNOR U486 ( .A(\min_val_reg[2][2] ), .B(n327), .Z(n328) );
  XOR U487 ( .A(\min_val_reg[3][2] ), .B(n471), .Z(n327) );
  NAND U488 ( .A(n278), .B(n239), .Z(n471) );
  XNOR U489 ( .A(\min_val_reg[3][2] ), .B(n277), .Z(n278) );
  XOR U490 ( .A(\min_val_reg[4][2] ), .B(n472), .Z(n277) );
  NAND U491 ( .A(n230), .B(n191), .Z(n472) );
  XNOR U492 ( .A(\min_val_reg[4][2] ), .B(n229), .Z(n230) );
  XOR U493 ( .A(\min_val_reg[5][2] ), .B(n473), .Z(n229) );
  NAND U494 ( .A(n180), .B(n158), .Z(n473) );
  XOR U495 ( .A(\min_val_reg[5][2] ), .B(n179), .Z(n180) );
  XNOR U496 ( .A(\min_val_reg[6][2] ), .B(n474), .Z(n179) );
  NAND U497 ( .A(n475), .B(n410), .Z(n474) );
  XNOR U498 ( .A(n476), .B(n477), .Z(min_val_out[16]) );
  AND U499 ( .A(n387), .B(n448), .Z(n476) );
  XNOR U500 ( .A(\min_val_reg[0][1] ), .B(n477), .Z(n448) );
  XOR U501 ( .A(\min_val_reg[1][1] ), .B(n478), .Z(n477) );
  NAND U502 ( .A(n379), .B(n337), .Z(n478) );
  XNOR U503 ( .A(\min_val_reg[1][1] ), .B(n378), .Z(n379) );
  XOR U504 ( .A(\min_val_reg[2][1] ), .B(n479), .Z(n378) );
  NAND U505 ( .A(n331), .B(n289), .Z(n479) );
  XNOR U506 ( .A(\min_val_reg[2][1] ), .B(n330), .Z(n331) );
  XOR U507 ( .A(\min_val_reg[3][1] ), .B(n480), .Z(n330) );
  NAND U508 ( .A(n281), .B(n239), .Z(n480) );
  XNOR U509 ( .A(\min_val_reg[3][1] ), .B(n280), .Z(n281) );
  XOR U510 ( .A(\min_val_reg[4][1] ), .B(n481), .Z(n280) );
  NAND U511 ( .A(n233), .B(n191), .Z(n481) );
  XNOR U512 ( .A(\min_val_reg[4][1] ), .B(n232), .Z(n233) );
  XOR U513 ( .A(\min_val_reg[5][1] ), .B(n482), .Z(n232) );
  NAND U514 ( .A(n183), .B(n158), .Z(n482) );
  XOR U515 ( .A(\min_val_reg[5][1] ), .B(n182), .Z(n183) );
  XNOR U516 ( .A(\min_val_reg[6][1] ), .B(n483), .Z(n182) );
  NAND U517 ( .A(n484), .B(n410), .Z(n483) );
  XNOR U518 ( .A(n485), .B(n486), .Z(min_val_out[15]) );
  AND U519 ( .A(n387), .B(n487), .Z(n485) );
  XOR U520 ( .A(\min_val_reg[0][14] ), .B(n488), .Z(min_val_out[14]) );
  AND U521 ( .A(n154), .B(n388), .Z(n488) );
  XNOR U522 ( .A(\min_val_reg[0][14] ), .B(n386), .Z(n388) );
  XOR U523 ( .A(\min_val_reg[1][14] ), .B(n489), .Z(n386) );
  NAND U524 ( .A(n338), .B(n337), .Z(n489) );
  XNOR U525 ( .A(\min_val_reg[1][14] ), .B(n336), .Z(n338) );
  XOR U526 ( .A(\min_val_reg[2][14] ), .B(n490), .Z(n336) );
  NAND U527 ( .A(n290), .B(n289), .Z(n490) );
  XNOR U528 ( .A(\min_val_reg[2][14] ), .B(n288), .Z(n290) );
  XOR U529 ( .A(\min_val_reg[3][14] ), .B(n491), .Z(n288) );
  NAND U530 ( .A(n240), .B(n239), .Z(n491) );
  XNOR U531 ( .A(\min_val_reg[3][14] ), .B(n238), .Z(n240) );
  XOR U532 ( .A(\min_val_reg[4][14] ), .B(n492), .Z(n238) );
  NAND U533 ( .A(n192), .B(n191), .Z(n492) );
  XOR U534 ( .A(\min_val_reg[4][14] ), .B(n190), .Z(n192) );
  XNOR U535 ( .A(\min_val_reg[5][14] ), .B(n493), .Z(n190) );
  NAND U536 ( .A(n494), .B(n158), .Z(n493) );
  XOR U537 ( .A(\min_val_reg[0][13] ), .B(n495), .Z(min_val_out[13]) );
  AND U538 ( .A(n154), .B(n391), .Z(n495) );
  XNOR U539 ( .A(\min_val_reg[0][13] ), .B(n390), .Z(n391) );
  XOR U540 ( .A(\min_val_reg[1][13] ), .B(n496), .Z(n390) );
  NAND U541 ( .A(n341), .B(n337), .Z(n496) );
  XNOR U542 ( .A(\min_val_reg[1][13] ), .B(n340), .Z(n341) );
  XOR U543 ( .A(\min_val_reg[2][13] ), .B(n497), .Z(n340) );
  NAND U544 ( .A(n293), .B(n289), .Z(n497) );
  XNOR U545 ( .A(\min_val_reg[2][13] ), .B(n292), .Z(n293) );
  XOR U546 ( .A(\min_val_reg[3][13] ), .B(n498), .Z(n292) );
  NAND U547 ( .A(n243), .B(n239), .Z(n498) );
  XNOR U548 ( .A(\min_val_reg[3][13] ), .B(n242), .Z(n243) );
  XOR U549 ( .A(\min_val_reg[4][13] ), .B(n499), .Z(n242) );
  NAND U550 ( .A(n195), .B(n191), .Z(n499) );
  XOR U551 ( .A(\min_val_reg[4][13] ), .B(n194), .Z(n195) );
  XNOR U552 ( .A(\min_val_reg[5][13] ), .B(n500), .Z(n194) );
  NAND U553 ( .A(n501), .B(n158), .Z(n500) );
  XOR U554 ( .A(\min_val_reg[0][12] ), .B(n502), .Z(min_val_out[12]) );
  AND U555 ( .A(n154), .B(n394), .Z(n502) );
  XNOR U556 ( .A(\min_val_reg[0][12] ), .B(n393), .Z(n394) );
  XOR U557 ( .A(\min_val_reg[1][12] ), .B(n503), .Z(n393) );
  NAND U558 ( .A(n344), .B(n337), .Z(n503) );
  XNOR U559 ( .A(\min_val_reg[1][12] ), .B(n343), .Z(n344) );
  XOR U560 ( .A(\min_val_reg[2][12] ), .B(n504), .Z(n343) );
  NAND U561 ( .A(n296), .B(n289), .Z(n504) );
  XNOR U562 ( .A(\min_val_reg[2][12] ), .B(n295), .Z(n296) );
  XOR U563 ( .A(\min_val_reg[3][12] ), .B(n505), .Z(n295) );
  NAND U564 ( .A(n246), .B(n239), .Z(n505) );
  XNOR U565 ( .A(\min_val_reg[3][12] ), .B(n245), .Z(n246) );
  XOR U566 ( .A(\min_val_reg[4][12] ), .B(n506), .Z(n245) );
  NAND U567 ( .A(n198), .B(n191), .Z(n506) );
  XOR U568 ( .A(\min_val_reg[4][12] ), .B(n197), .Z(n198) );
  XNOR U569 ( .A(\min_val_reg[5][12] ), .B(n507), .Z(n197) );
  NAND U570 ( .A(n508), .B(n158), .Z(n507) );
  XOR U571 ( .A(\min_val_reg[0][11] ), .B(n509), .Z(min_val_out[11]) );
  AND U572 ( .A(n154), .B(n397), .Z(n509) );
  XNOR U573 ( .A(\min_val_reg[0][11] ), .B(n396), .Z(n397) );
  XOR U574 ( .A(\min_val_reg[1][11] ), .B(n510), .Z(n396) );
  NAND U575 ( .A(n347), .B(n337), .Z(n510) );
  XNOR U576 ( .A(\min_val_reg[1][11] ), .B(n346), .Z(n347) );
  XOR U577 ( .A(\min_val_reg[2][11] ), .B(n511), .Z(n346) );
  NAND U578 ( .A(n299), .B(n289), .Z(n511) );
  XNOR U579 ( .A(\min_val_reg[2][11] ), .B(n298), .Z(n299) );
  XOR U580 ( .A(\min_val_reg[3][11] ), .B(n512), .Z(n298) );
  NAND U581 ( .A(n249), .B(n239), .Z(n512) );
  XNOR U582 ( .A(\min_val_reg[3][11] ), .B(n248), .Z(n249) );
  XOR U583 ( .A(\min_val_reg[4][11] ), .B(n513), .Z(n248) );
  NAND U584 ( .A(n201), .B(n191), .Z(n513) );
  XOR U585 ( .A(\min_val_reg[4][11] ), .B(n200), .Z(n201) );
  XNOR U586 ( .A(\min_val_reg[5][11] ), .B(n514), .Z(n200) );
  NAND U587 ( .A(n515), .B(n158), .Z(n514) );
  XNOR U588 ( .A(n516), .B(n517), .Z(min_val_out[119]) );
  AND U589 ( .A(n410), .B(n518), .Z(n516) );
  XNOR U590 ( .A(n519), .B(n520), .Z(min_val_out[118]) );
  AND U591 ( .A(n410), .B(n521), .Z(n519) );
  XNOR U592 ( .A(n522), .B(n523), .Z(min_val_out[117]) );
  AND U593 ( .A(n410), .B(n524), .Z(n522) );
  XNOR U594 ( .A(n525), .B(n526), .Z(min_val_out[116]) );
  AND U595 ( .A(n410), .B(n527), .Z(n525) );
  XNOR U596 ( .A(n528), .B(n529), .Z(min_val_out[115]) );
  AND U597 ( .A(n410), .B(n530), .Z(n528) );
  XNOR U598 ( .A(n531), .B(n532), .Z(min_val_out[114]) );
  AND U599 ( .A(n410), .B(n409), .Z(n531) );
  XNOR U600 ( .A(\min_val_reg[6][9] ), .B(n532), .Z(n409) );
  XOR U601 ( .A(\min_val_reg[7][9] ), .B(n533), .Z(n532) );
  NAND U602 ( .A(n534), .B(n535), .Z(n533) );
  XOR U603 ( .A(\min_val_reg[7][9] ), .B(DB[9]), .Z(n534) );
  XNOR U604 ( .A(n536), .B(n537), .Z(min_val_out[113]) );
  AND U605 ( .A(n410), .B(n419), .Z(n536) );
  XNOR U606 ( .A(\min_val_reg[6][8] ), .B(n537), .Z(n419) );
  XOR U607 ( .A(\min_val_reg[7][8] ), .B(n538), .Z(n537) );
  NAND U608 ( .A(n539), .B(n535), .Z(n538) );
  XOR U609 ( .A(\min_val_reg[7][8] ), .B(DB[8]), .Z(n539) );
  XNOR U610 ( .A(n540), .B(n541), .Z(min_val_out[112]) );
  AND U611 ( .A(n410), .B(n428), .Z(n540) );
  XNOR U612 ( .A(\min_val_reg[6][7] ), .B(n541), .Z(n428) );
  XOR U613 ( .A(\min_val_reg[7][7] ), .B(n542), .Z(n541) );
  NAND U614 ( .A(n543), .B(n535), .Z(n542) );
  XOR U615 ( .A(\min_val_reg[7][7] ), .B(DB[7]), .Z(n543) );
  XNOR U616 ( .A(n544), .B(n545), .Z(min_val_out[111]) );
  AND U617 ( .A(n410), .B(n437), .Z(n544) );
  XNOR U618 ( .A(\min_val_reg[6][6] ), .B(n545), .Z(n437) );
  XOR U619 ( .A(\min_val_reg[7][6] ), .B(n546), .Z(n545) );
  NAND U620 ( .A(n547), .B(n535), .Z(n546) );
  XOR U621 ( .A(\min_val_reg[7][6] ), .B(DB[6]), .Z(n547) );
  XNOR U622 ( .A(n548), .B(n549), .Z(min_val_out[110]) );
  AND U623 ( .A(n410), .B(n446), .Z(n548) );
  XNOR U624 ( .A(\min_val_reg[6][5] ), .B(n549), .Z(n446) );
  XOR U625 ( .A(\min_val_reg[7][5] ), .B(n550), .Z(n549) );
  NAND U626 ( .A(n551), .B(n535), .Z(n550) );
  XOR U627 ( .A(\min_val_reg[7][5] ), .B(DB[5]), .Z(n551) );
  XOR U628 ( .A(\min_val_reg[0][10] ), .B(n552), .Z(min_val_out[10]) );
  AND U629 ( .A(n154), .B(n400), .Z(n552) );
  XNOR U630 ( .A(\min_val_reg[0][10] ), .B(n399), .Z(n400) );
  XOR U631 ( .A(\min_val_reg[1][10] ), .B(n553), .Z(n399) );
  NAND U632 ( .A(n350), .B(n337), .Z(n553) );
  XNOR U633 ( .A(\min_val_reg[1][10] ), .B(n349), .Z(n350) );
  XOR U634 ( .A(\min_val_reg[2][10] ), .B(n554), .Z(n349) );
  NAND U635 ( .A(n302), .B(n289), .Z(n554) );
  XNOR U636 ( .A(\min_val_reg[2][10] ), .B(n301), .Z(n302) );
  XOR U637 ( .A(\min_val_reg[3][10] ), .B(n555), .Z(n301) );
  NAND U638 ( .A(n252), .B(n239), .Z(n555) );
  XNOR U639 ( .A(\min_val_reg[3][10] ), .B(n251), .Z(n252) );
  XOR U640 ( .A(\min_val_reg[4][10] ), .B(n556), .Z(n251) );
  NAND U641 ( .A(n204), .B(n191), .Z(n556) );
  XOR U642 ( .A(\min_val_reg[4][10] ), .B(n203), .Z(n204) );
  XNOR U643 ( .A(\min_val_reg[5][10] ), .B(n557), .Z(n203) );
  NAND U644 ( .A(n558), .B(n158), .Z(n557) );
  XNOR U645 ( .A(n559), .B(n560), .Z(min_val_out[109]) );
  AND U646 ( .A(n410), .B(n457), .Z(n559) );
  XNOR U647 ( .A(\min_val_reg[6][4] ), .B(n560), .Z(n457) );
  XOR U648 ( .A(\min_val_reg[7][4] ), .B(n561), .Z(n560) );
  NAND U649 ( .A(n562), .B(n535), .Z(n561) );
  XOR U650 ( .A(\min_val_reg[7][4] ), .B(DB[4]), .Z(n562) );
  XNOR U651 ( .A(n563), .B(n564), .Z(min_val_out[108]) );
  AND U652 ( .A(n410), .B(n466), .Z(n563) );
  XNOR U653 ( .A(\min_val_reg[6][3] ), .B(n564), .Z(n466) );
  XOR U654 ( .A(\min_val_reg[7][3] ), .B(n565), .Z(n564) );
  NAND U655 ( .A(n566), .B(n535), .Z(n565) );
  XOR U656 ( .A(\min_val_reg[7][3] ), .B(DB[3]), .Z(n566) );
  XNOR U657 ( .A(n567), .B(n568), .Z(min_val_out[107]) );
  AND U658 ( .A(n410), .B(n475), .Z(n567) );
  XNOR U659 ( .A(\min_val_reg[6][2] ), .B(n568), .Z(n475) );
  XOR U660 ( .A(\min_val_reg[7][2] ), .B(n569), .Z(n568) );
  NAND U661 ( .A(n570), .B(n535), .Z(n569) );
  XOR U662 ( .A(\min_val_reg[7][2] ), .B(DB[2]), .Z(n570) );
  XNOR U663 ( .A(n571), .B(n572), .Z(min_val_out[106]) );
  AND U664 ( .A(n410), .B(n484), .Z(n571) );
  XNOR U665 ( .A(\min_val_reg[6][1] ), .B(n572), .Z(n484) );
  XOR U666 ( .A(\min_val_reg[7][1] ), .B(n573), .Z(n572) );
  NAND U667 ( .A(n574), .B(n535), .Z(n573) );
  XOR U668 ( .A(\min_val_reg[7][1] ), .B(DB[1]), .Z(n574) );
  XNOR U669 ( .A(n575), .B(n576), .Z(min_val_out[105]) );
  AND U670 ( .A(n410), .B(n577), .Z(n575) );
  XOR U671 ( .A(n578), .B(n579), .Z(min_val_out[104]) );
  AND U672 ( .A(n158), .B(n494), .Z(n578) );
  XOR U673 ( .A(\min_val_reg[5][14] ), .B(n579), .Z(n494) );
  XNOR U674 ( .A(\min_val_reg[6][14] ), .B(n580), .Z(n579) );
  NAND U675 ( .A(n518), .B(n410), .Z(n580) );
  XNOR U676 ( .A(\min_val_reg[6][14] ), .B(n517), .Z(n518) );
  XOR U677 ( .A(\min_val_reg[7][14] ), .B(n581), .Z(n517) );
  NAND U678 ( .A(n582), .B(n535), .Z(n581) );
  XOR U679 ( .A(\min_val_reg[7][14] ), .B(DB[14]), .Z(n582) );
  XOR U680 ( .A(n583), .B(n584), .Z(min_val_out[103]) );
  AND U681 ( .A(n158), .B(n501), .Z(n583) );
  XOR U682 ( .A(\min_val_reg[5][13] ), .B(n584), .Z(n501) );
  XNOR U683 ( .A(\min_val_reg[6][13] ), .B(n585), .Z(n584) );
  NAND U684 ( .A(n521), .B(n410), .Z(n585) );
  XNOR U685 ( .A(\min_val_reg[6][13] ), .B(n520), .Z(n521) );
  XOR U686 ( .A(\min_val_reg[7][13] ), .B(n586), .Z(n520) );
  NAND U687 ( .A(n587), .B(n535), .Z(n586) );
  XOR U688 ( .A(\min_val_reg[7][13] ), .B(DB[13]), .Z(n587) );
  XOR U689 ( .A(n588), .B(n589), .Z(min_val_out[102]) );
  AND U690 ( .A(n158), .B(n508), .Z(n588) );
  XOR U691 ( .A(\min_val_reg[5][12] ), .B(n589), .Z(n508) );
  XNOR U692 ( .A(\min_val_reg[6][12] ), .B(n590), .Z(n589) );
  NAND U693 ( .A(n524), .B(n410), .Z(n590) );
  XNOR U694 ( .A(\min_val_reg[6][12] ), .B(n523), .Z(n524) );
  XOR U695 ( .A(\min_val_reg[7][12] ), .B(n591), .Z(n523) );
  NAND U696 ( .A(n592), .B(n535), .Z(n591) );
  XOR U697 ( .A(\min_val_reg[7][12] ), .B(DB[12]), .Z(n592) );
  XOR U698 ( .A(n593), .B(n594), .Z(min_val_out[101]) );
  AND U699 ( .A(n158), .B(n515), .Z(n593) );
  XOR U700 ( .A(\min_val_reg[5][11] ), .B(n594), .Z(n515) );
  XNOR U701 ( .A(\min_val_reg[6][11] ), .B(n595), .Z(n594) );
  NAND U702 ( .A(n527), .B(n410), .Z(n595) );
  XNOR U703 ( .A(\min_val_reg[6][11] ), .B(n526), .Z(n527) );
  XOR U704 ( .A(\min_val_reg[7][11] ), .B(n596), .Z(n526) );
  NAND U705 ( .A(n597), .B(n535), .Z(n596) );
  XOR U706 ( .A(\min_val_reg[7][11] ), .B(DB[11]), .Z(n597) );
  XOR U707 ( .A(n598), .B(n599), .Z(min_val_out[100]) );
  AND U708 ( .A(n158), .B(n558), .Z(n598) );
  XOR U709 ( .A(\min_val_reg[5][10] ), .B(n599), .Z(n558) );
  XNOR U710 ( .A(\min_val_reg[6][10] ), .B(n600), .Z(n599) );
  NAND U711 ( .A(n530), .B(n410), .Z(n600) );
  XNOR U712 ( .A(\min_val_reg[6][10] ), .B(n529), .Z(n530) );
  XOR U713 ( .A(\min_val_reg[7][10] ), .B(n601), .Z(n529) );
  NAND U714 ( .A(n602), .B(n535), .Z(n601) );
  XOR U715 ( .A(\min_val_reg[7][10] ), .B(DB[10]), .Z(n602) );
  XOR U716 ( .A(\min_val_reg[0][0] ), .B(n603), .Z(min_val_out[0]) );
  AND U717 ( .A(n154), .B(n487), .Z(n603) );
  XNOR U718 ( .A(\min_val_reg[0][0] ), .B(n486), .Z(n487) );
  XOR U719 ( .A(\min_val_reg[1][0] ), .B(n604), .Z(n486) );
  NAND U720 ( .A(n382), .B(n337), .Z(n604) );
  XNOR U721 ( .A(\min_val_reg[1][0] ), .B(n381), .Z(n382) );
  XOR U722 ( .A(\min_val_reg[2][0] ), .B(n605), .Z(n381) );
  NAND U723 ( .A(n334), .B(n289), .Z(n605) );
  XNOR U724 ( .A(\min_val_reg[2][0] ), .B(n333), .Z(n334) );
  XOR U725 ( .A(\min_val_reg[3][0] ), .B(n606), .Z(n333) );
  NAND U726 ( .A(n284), .B(n239), .Z(n606) );
  XNOR U727 ( .A(\min_val_reg[3][0] ), .B(n283), .Z(n284) );
  XOR U728 ( .A(\min_val_reg[4][0] ), .B(n607), .Z(n283) );
  NAND U729 ( .A(n236), .B(n191), .Z(n607) );
  XNOR U730 ( .A(\min_val_reg[4][0] ), .B(n235), .Z(n236) );
  XOR U731 ( .A(\min_val_reg[5][0] ), .B(n608), .Z(n235) );
  NAND U732 ( .A(n186), .B(n158), .Z(n608) );
  XOR U733 ( .A(\min_val_reg[5][0] ), .B(n185), .Z(n186) );
  XNOR U734 ( .A(\min_val_reg[6][0] ), .B(n609), .Z(n185) );
  NAND U735 ( .A(n577), .B(n410), .Z(n609) );
  XNOR U736 ( .A(\min_val_reg[6][0] ), .B(n576), .Z(n577) );
  XOR U737 ( .A(\min_val_reg[7][0] ), .B(n610), .Z(n576) );
  NAND U738 ( .A(n611), .B(n535), .Z(n610) );
  XOR U739 ( .A(\min_val_reg[7][0] ), .B(DB[0]), .Z(n611) );
  XOR U740 ( .A(n612), .B(n613), .Z(\min_dist[7][3] ) );
  AND U741 ( .A(n410), .B(n614), .Z(n612) );
  XOR U742 ( .A(\min_dist_reg[6][3] ), .B(n613), .Z(n614) );
  XOR U743 ( .A(n615), .B(n616), .Z(\min_dist[7][2] ) );
  AND U744 ( .A(n410), .B(n617), .Z(n615) );
  XNOR U745 ( .A(\min_dist_reg[6][2] ), .B(n618), .Z(n617) );
  XOR U746 ( .A(n619), .B(n620), .Z(\min_dist[7][1] ) );
  AND U747 ( .A(n410), .B(n621), .Z(n619) );
  XNOR U748 ( .A(\min_dist_reg[6][1] ), .B(n622), .Z(n621) );
  XOR U749 ( .A(n623), .B(n624), .Z(\min_dist[7][0] ) );
  AND U750 ( .A(n410), .B(n625), .Z(n623) );
  XOR U751 ( .A(n626), .B(n627), .Z(\min_dist[6][3] ) );
  AND U752 ( .A(n158), .B(n628), .Z(n626) );
  XOR U753 ( .A(\min_dist_reg[5][3] ), .B(n627), .Z(n628) );
  XOR U754 ( .A(n629), .B(n630), .Z(\min_dist[6][2] ) );
  AND U755 ( .A(n158), .B(n631), .Z(n629) );
  XOR U756 ( .A(\min_dist_reg[5][2] ), .B(n630), .Z(n631) );
  XOR U757 ( .A(n632), .B(n633), .Z(\min_dist[6][1] ) );
  AND U758 ( .A(n158), .B(n634), .Z(n632) );
  XOR U759 ( .A(\min_dist_reg[5][1] ), .B(n633), .Z(n634) );
  XOR U760 ( .A(n635), .B(n636), .Z(\min_dist[6][0] ) );
  AND U761 ( .A(n158), .B(n637), .Z(n635) );
  XOR U762 ( .A(n638), .B(n639), .Z(\min_dist[5][3] ) );
  AND U763 ( .A(n191), .B(n640), .Z(n638) );
  XOR U764 ( .A(\min_dist_reg[4][3] ), .B(n639), .Z(n640) );
  XOR U765 ( .A(n641), .B(n642), .Z(\min_dist[5][2] ) );
  AND U766 ( .A(n191), .B(n643), .Z(n641) );
  XOR U767 ( .A(\min_dist_reg[4][2] ), .B(n642), .Z(n643) );
  XOR U768 ( .A(n644), .B(n645), .Z(\min_dist[5][1] ) );
  AND U769 ( .A(n191), .B(n646), .Z(n644) );
  XOR U770 ( .A(\min_dist_reg[4][1] ), .B(n645), .Z(n646) );
  XOR U771 ( .A(n647), .B(n648), .Z(\min_dist[5][0] ) );
  AND U772 ( .A(n191), .B(n649), .Z(n647) );
  XOR U773 ( .A(n650), .B(n651), .Z(\min_dist[4][3] ) );
  AND U774 ( .A(n239), .B(n652), .Z(n650) );
  XOR U775 ( .A(\min_dist_reg[3][3] ), .B(n651), .Z(n652) );
  XOR U776 ( .A(n653), .B(n654), .Z(\min_dist[4][2] ) );
  AND U777 ( .A(n239), .B(n655), .Z(n653) );
  XOR U778 ( .A(\min_dist_reg[3][2] ), .B(n654), .Z(n655) );
  XOR U779 ( .A(n656), .B(n657), .Z(\min_dist[4][1] ) );
  AND U780 ( .A(n239), .B(n658), .Z(n656) );
  XOR U781 ( .A(\min_dist_reg[3][1] ), .B(n657), .Z(n658) );
  XOR U782 ( .A(n659), .B(n660), .Z(\min_dist[4][0] ) );
  AND U783 ( .A(n239), .B(n661), .Z(n659) );
  XOR U784 ( .A(n662), .B(n663), .Z(\min_dist[3][3] ) );
  AND U785 ( .A(n289), .B(n664), .Z(n662) );
  XOR U786 ( .A(\min_dist_reg[2][3] ), .B(n663), .Z(n664) );
  XOR U787 ( .A(n665), .B(n666), .Z(\min_dist[3][2] ) );
  AND U788 ( .A(n289), .B(n667), .Z(n665) );
  XOR U789 ( .A(\min_dist_reg[2][2] ), .B(n666), .Z(n667) );
  XOR U790 ( .A(n668), .B(n669), .Z(\min_dist[3][1] ) );
  AND U791 ( .A(n289), .B(n670), .Z(n668) );
  XOR U792 ( .A(\min_dist_reg[2][1] ), .B(n669), .Z(n670) );
  XOR U793 ( .A(n671), .B(n672), .Z(\min_dist[3][0] ) );
  AND U794 ( .A(n289), .B(n673), .Z(n671) );
  XOR U795 ( .A(n674), .B(n675), .Z(\min_dist[2][3] ) );
  AND U796 ( .A(n337), .B(n676), .Z(n674) );
  XOR U797 ( .A(\min_dist_reg[1][3] ), .B(n675), .Z(n676) );
  XOR U798 ( .A(n677), .B(n678), .Z(\min_dist[2][2] ) );
  AND U799 ( .A(n337), .B(n679), .Z(n677) );
  XOR U800 ( .A(\min_dist_reg[1][2] ), .B(n678), .Z(n679) );
  XOR U801 ( .A(n680), .B(n681), .Z(\min_dist[2][1] ) );
  AND U802 ( .A(n337), .B(n682), .Z(n680) );
  XOR U803 ( .A(\min_dist_reg[1][1] ), .B(n681), .Z(n682) );
  XOR U804 ( .A(n683), .B(n684), .Z(\min_dist[2][0] ) );
  AND U805 ( .A(n337), .B(n685), .Z(n683) );
  XOR U806 ( .A(n686), .B(n687), .Z(\min_dist[1][3] ) );
  AND U807 ( .A(n387), .B(n688), .Z(n686) );
  XOR U808 ( .A(\min_dist_reg[0][3] ), .B(n687), .Z(n688) );
  XOR U809 ( .A(n689), .B(n690), .Z(\min_dist[1][2] ) );
  AND U810 ( .A(n387), .B(n691), .Z(n689) );
  XOR U811 ( .A(n692), .B(n693), .Z(\min_dist[1][1] ) );
  AND U812 ( .A(n387), .B(n694), .Z(n692) );
  XNOR U813 ( .A(n695), .B(n696), .Z(\min_dist[1][0] ) );
  AND U814 ( .A(n387), .B(n697), .Z(n695) );
  XNOR U815 ( .A(\min_dist_reg[0][0] ), .B(n696), .Z(n697) );
  XNOR U816 ( .A(n698), .B(n699), .Z(n387) );
  AND U817 ( .A(n700), .B(n701), .Z(n698) );
  XOR U818 ( .A(n687), .B(n699), .Z(n701) );
  XNOR U819 ( .A(\min_dist_reg[0][3] ), .B(n699), .Z(n700) );
  XNOR U820 ( .A(n702), .B(n703), .Z(n699) );
  AND U821 ( .A(n704), .B(n705), .Z(n702) );
  XNOR U822 ( .A(n690), .B(n703), .Z(n705) );
  XOR U823 ( .A(\min_dist_reg[0][2] ), .B(n703), .Z(n704) );
  XOR U824 ( .A(n706), .B(n707), .Z(n703) );
  NAND U825 ( .A(n708), .B(n709), .Z(n707) );
  XOR U826 ( .A(n706), .B(n693), .Z(n709) );
  XNOR U827 ( .A(\min_dist_reg[0][1] ), .B(n706), .Z(n708) );
  NOR U828 ( .A(n696), .B(\min_dist_reg[0][0] ), .Z(n706) );
  AND U829 ( .A(\min_dist_reg[0][3] ), .B(n710), .Z(\local_min_dist[0][3] ) );
  NANDN U830 ( .A(n687), .B(n154), .Z(n710) );
  XOR U831 ( .A(\min_dist_reg[0][2] ), .B(n711), .Z(\local_min_dist[0][2] ) );
  AND U832 ( .A(n154), .B(n691), .Z(n711) );
  XOR U833 ( .A(\min_dist_reg[0][2] ), .B(n690), .Z(n691) );
  XOR U834 ( .A(\min_dist_reg[0][1] ), .B(n712), .Z(\local_min_dist[0][1] ) );
  AND U835 ( .A(n154), .B(n694), .Z(n712) );
  XOR U836 ( .A(\min_dist_reg[0][1] ), .B(n693), .Z(n694) );
  XOR U837 ( .A(\min_dist_reg[0][0] ), .B(n713), .Z(\local_min_dist[0][0] ) );
  AND U838 ( .A(n154), .B(n714), .Z(n713) );
  XOR U839 ( .A(\min_dist_reg[0][0] ), .B(n715), .Z(n714) );
  XNOR U840 ( .A(n716), .B(n717), .Z(n154) );
  AND U841 ( .A(n718), .B(n719), .Z(n716) );
  XOR U842 ( .A(n687), .B(n717), .Z(n719) );
  AND U843 ( .A(n720), .B(\min_dist_reg[1][3] ), .Z(n687) );
  NANDN U844 ( .A(n675), .B(n337), .Z(n720) );
  XNOR U845 ( .A(\min_dist_reg[0][3] ), .B(n717), .Z(n718) );
  XNOR U846 ( .A(n721), .B(n722), .Z(n717) );
  AND U847 ( .A(n723), .B(n724), .Z(n721) );
  XNOR U848 ( .A(n722), .B(n690), .Z(n724) );
  XNOR U849 ( .A(\min_dist_reg[1][2] ), .B(n725), .Z(n690) );
  NAND U850 ( .A(n726), .B(n337), .Z(n725) );
  XNOR U851 ( .A(n727), .B(n678), .Z(n726) );
  XOR U852 ( .A(\min_dist_reg[0][2] ), .B(n722), .Z(n723) );
  XOR U853 ( .A(n728), .B(n729), .Z(n722) );
  NAND U854 ( .A(n730), .B(n731), .Z(n729) );
  XOR U855 ( .A(n728), .B(n693), .Z(n731) );
  XNOR U856 ( .A(\min_dist_reg[1][1] ), .B(n732), .Z(n693) );
  NAND U857 ( .A(n733), .B(n337), .Z(n732) );
  XNOR U858 ( .A(n734), .B(n681), .Z(n733) );
  XNOR U859 ( .A(\min_dist_reg[0][1] ), .B(n728), .Z(n730) );
  ANDN U860 ( .B(n715), .A(\min_dist_reg[0][0] ), .Z(n728) );
  IV U861 ( .A(n696), .Z(n715) );
  XOR U862 ( .A(\min_dist_reg[1][0] ), .B(n735), .Z(n696) );
  NAND U863 ( .A(n685), .B(n337), .Z(n735) );
  XOR U864 ( .A(n736), .B(n737), .Z(n337) );
  AND U865 ( .A(n738), .B(n739), .Z(n736) );
  XNOR U866 ( .A(n675), .B(n737), .Z(n739) );
  AND U867 ( .A(n740), .B(\min_dist_reg[2][3] ), .Z(n675) );
  NANDN U868 ( .A(n663), .B(n289), .Z(n740) );
  XNOR U869 ( .A(n741), .B(n737), .Z(n738) );
  XOR U870 ( .A(n742), .B(n743), .Z(n737) );
  AND U871 ( .A(n744), .B(n745), .Z(n742) );
  XNOR U872 ( .A(n678), .B(n743), .Z(n745) );
  XNOR U873 ( .A(\min_dist_reg[2][2] ), .B(n746), .Z(n678) );
  NAND U874 ( .A(n747), .B(n289), .Z(n746) );
  XNOR U875 ( .A(n748), .B(n666), .Z(n747) );
  XNOR U876 ( .A(n727), .B(n743), .Z(n744) );
  XOR U877 ( .A(n749), .B(n750), .Z(n743) );
  NAND U878 ( .A(n751), .B(n752), .Z(n750) );
  XOR U879 ( .A(n749), .B(n681), .Z(n752) );
  XNOR U880 ( .A(\min_dist_reg[2][1] ), .B(n753), .Z(n681) );
  NAND U881 ( .A(n754), .B(n289), .Z(n753) );
  XNOR U882 ( .A(n755), .B(n669), .Z(n754) );
  XOR U883 ( .A(n734), .B(n749), .Z(n751) );
  IV U884 ( .A(\min_dist_reg[1][1] ), .Z(n734) );
  AND U885 ( .A(n684), .B(n756), .Z(n749) );
  IV U886 ( .A(\min_dist_reg[1][2] ), .Z(n727) );
  IV U887 ( .A(\min_dist_reg[1][3] ), .Z(n741) );
  XNOR U888 ( .A(n756), .B(n684), .Z(n685) );
  XNOR U889 ( .A(\min_dist_reg[2][0] ), .B(n757), .Z(n684) );
  NAND U890 ( .A(n673), .B(n289), .Z(n757) );
  XOR U891 ( .A(n758), .B(n759), .Z(n289) );
  AND U892 ( .A(n760), .B(n761), .Z(n758) );
  XNOR U893 ( .A(n663), .B(n759), .Z(n761) );
  AND U894 ( .A(n762), .B(\min_dist_reg[3][3] ), .Z(n663) );
  NANDN U895 ( .A(n651), .B(n239), .Z(n762) );
  XNOR U896 ( .A(n763), .B(n759), .Z(n760) );
  XOR U897 ( .A(n764), .B(n765), .Z(n759) );
  AND U898 ( .A(n766), .B(n767), .Z(n764) );
  XNOR U899 ( .A(n666), .B(n765), .Z(n767) );
  XNOR U900 ( .A(\min_dist_reg[3][2] ), .B(n768), .Z(n666) );
  NAND U901 ( .A(n769), .B(n239), .Z(n768) );
  XNOR U902 ( .A(n770), .B(n654), .Z(n769) );
  XNOR U903 ( .A(n748), .B(n765), .Z(n766) );
  XOR U904 ( .A(n771), .B(n772), .Z(n765) );
  NAND U905 ( .A(n773), .B(n774), .Z(n772) );
  XOR U906 ( .A(n771), .B(n669), .Z(n774) );
  XNOR U907 ( .A(\min_dist_reg[3][1] ), .B(n775), .Z(n669) );
  NAND U908 ( .A(n776), .B(n239), .Z(n775) );
  XNOR U909 ( .A(n777), .B(n657), .Z(n776) );
  XOR U910 ( .A(n755), .B(n771), .Z(n773) );
  IV U911 ( .A(\min_dist_reg[2][1] ), .Z(n755) );
  ANDN U912 ( .B(n672), .A(\min_dist_reg[2][0] ), .Z(n771) );
  IV U913 ( .A(\min_dist_reg[2][2] ), .Z(n748) );
  IV U914 ( .A(\min_dist_reg[2][3] ), .Z(n763) );
  XOR U915 ( .A(\min_dist_reg[2][0] ), .B(n672), .Z(n673) );
  XNOR U916 ( .A(\min_dist_reg[3][0] ), .B(n778), .Z(n672) );
  NAND U917 ( .A(n661), .B(n239), .Z(n778) );
  XOR U918 ( .A(n779), .B(n780), .Z(n239) );
  AND U919 ( .A(n781), .B(n782), .Z(n779) );
  XNOR U920 ( .A(n651), .B(n780), .Z(n782) );
  AND U921 ( .A(n783), .B(\min_dist_reg[4][3] ), .Z(n651) );
  NANDN U922 ( .A(n639), .B(n191), .Z(n783) );
  XNOR U923 ( .A(n784), .B(n780), .Z(n781) );
  XOR U924 ( .A(n785), .B(n786), .Z(n780) );
  AND U925 ( .A(n787), .B(n788), .Z(n785) );
  XNOR U926 ( .A(n654), .B(n786), .Z(n788) );
  XNOR U927 ( .A(\min_dist_reg[4][2] ), .B(n789), .Z(n654) );
  NAND U928 ( .A(n790), .B(n191), .Z(n789) );
  XNOR U929 ( .A(n791), .B(n642), .Z(n790) );
  XNOR U930 ( .A(n770), .B(n786), .Z(n787) );
  XOR U931 ( .A(n792), .B(n793), .Z(n786) );
  NAND U932 ( .A(n794), .B(n795), .Z(n793) );
  XOR U933 ( .A(n792), .B(n657), .Z(n795) );
  XNOR U934 ( .A(\min_dist_reg[4][1] ), .B(n796), .Z(n657) );
  NAND U935 ( .A(n797), .B(n191), .Z(n796) );
  XNOR U936 ( .A(n798), .B(n645), .Z(n797) );
  XOR U937 ( .A(n777), .B(n792), .Z(n794) );
  IV U938 ( .A(\min_dist_reg[3][1] ), .Z(n777) );
  ANDN U939 ( .B(n660), .A(\min_dist_reg[3][0] ), .Z(n792) );
  IV U940 ( .A(\min_dist_reg[3][2] ), .Z(n770) );
  IV U941 ( .A(\min_dist_reg[3][3] ), .Z(n784) );
  XOR U942 ( .A(\min_dist_reg[3][0] ), .B(n660), .Z(n661) );
  XNOR U943 ( .A(\min_dist_reg[4][0] ), .B(n799), .Z(n660) );
  NAND U944 ( .A(n649), .B(n191), .Z(n799) );
  XOR U945 ( .A(n800), .B(n801), .Z(n191) );
  AND U946 ( .A(n802), .B(n803), .Z(n800) );
  XNOR U947 ( .A(n639), .B(n801), .Z(n803) );
  AND U948 ( .A(n804), .B(\min_dist_reg[5][3] ), .Z(n639) );
  NANDN U949 ( .A(n627), .B(n158), .Z(n804) );
  XNOR U950 ( .A(n805), .B(n801), .Z(n802) );
  XOR U951 ( .A(n806), .B(n807), .Z(n801) );
  AND U952 ( .A(n808), .B(n809), .Z(n806) );
  XNOR U953 ( .A(n642), .B(n807), .Z(n809) );
  XNOR U954 ( .A(\min_dist_reg[5][2] ), .B(n810), .Z(n642) );
  NAND U955 ( .A(n811), .B(n158), .Z(n810) );
  XNOR U956 ( .A(n812), .B(n630), .Z(n811) );
  XNOR U957 ( .A(n791), .B(n807), .Z(n808) );
  XOR U958 ( .A(n813), .B(n814), .Z(n807) );
  NAND U959 ( .A(n815), .B(n816), .Z(n814) );
  XOR U960 ( .A(n813), .B(n645), .Z(n816) );
  XNOR U961 ( .A(\min_dist_reg[5][1] ), .B(n817), .Z(n645) );
  NAND U962 ( .A(n818), .B(n158), .Z(n817) );
  XNOR U963 ( .A(n819), .B(n633), .Z(n818) );
  XOR U964 ( .A(n798), .B(n813), .Z(n815) );
  IV U965 ( .A(\min_dist_reg[4][1] ), .Z(n798) );
  ANDN U966 ( .B(n648), .A(\min_dist_reg[4][0] ), .Z(n813) );
  IV U967 ( .A(\min_dist_reg[4][2] ), .Z(n791) );
  IV U968 ( .A(\min_dist_reg[4][3] ), .Z(n805) );
  XOR U969 ( .A(\min_dist_reg[4][0] ), .B(n648), .Z(n649) );
  XNOR U970 ( .A(\min_dist_reg[5][0] ), .B(n820), .Z(n648) );
  NAND U971 ( .A(n637), .B(n158), .Z(n820) );
  XOR U972 ( .A(n821), .B(n822), .Z(n158) );
  AND U973 ( .A(n823), .B(n824), .Z(n821) );
  XNOR U974 ( .A(n627), .B(n822), .Z(n824) );
  AND U975 ( .A(n825), .B(\min_dist_reg[6][3] ), .Z(n627) );
  NANDN U976 ( .A(n613), .B(n410), .Z(n825) );
  XNOR U977 ( .A(n826), .B(n822), .Z(n823) );
  XOR U978 ( .A(n827), .B(n828), .Z(n822) );
  AND U979 ( .A(n829), .B(n830), .Z(n827) );
  XNOR U980 ( .A(n630), .B(n828), .Z(n830) );
  XNOR U981 ( .A(\min_dist_reg[6][2] ), .B(n831), .Z(n630) );
  NAND U982 ( .A(n832), .B(n410), .Z(n831) );
  XNOR U983 ( .A(n833), .B(n616), .Z(n832) );
  XNOR U984 ( .A(n812), .B(n828), .Z(n829) );
  XOR U985 ( .A(n834), .B(n835), .Z(n828) );
  NAND U986 ( .A(n836), .B(n837), .Z(n835) );
  XOR U987 ( .A(n834), .B(n633), .Z(n837) );
  XNOR U988 ( .A(\min_dist_reg[6][1] ), .B(n838), .Z(n633) );
  NAND U989 ( .A(n839), .B(n410), .Z(n838) );
  XNOR U990 ( .A(n840), .B(n620), .Z(n839) );
  XOR U991 ( .A(n819), .B(n834), .Z(n836) );
  IV U992 ( .A(\min_dist_reg[5][1] ), .Z(n819) );
  ANDN U993 ( .B(n636), .A(\min_dist_reg[5][0] ), .Z(n834) );
  IV U994 ( .A(\min_dist_reg[5][2] ), .Z(n812) );
  IV U995 ( .A(\min_dist_reg[5][3] ), .Z(n826) );
  XOR U996 ( .A(\min_dist_reg[5][0] ), .B(n636), .Z(n637) );
  XNOR U997 ( .A(\min_dist_reg[6][0] ), .B(n841), .Z(n636) );
  NAND U998 ( .A(n625), .B(n410), .Z(n841) );
  XOR U999 ( .A(n842), .B(n843), .Z(n410) );
  AND U1000 ( .A(n844), .B(n845), .Z(n842) );
  XNOR U1001 ( .A(n613), .B(n843), .Z(n845) );
  XNOR U1002 ( .A(\min_dist_reg[7][3] ), .B(n846), .Z(n613) );
  NAND U1003 ( .A(n847), .B(n535), .Z(n846) );
  XOR U1004 ( .A(\min_dist_reg[7][3] ), .B(n848), .Z(n847) );
  XNOR U1005 ( .A(n849), .B(n843), .Z(n844) );
  XOR U1006 ( .A(n850), .B(n851), .Z(n843) );
  AND U1007 ( .A(n852), .B(n853), .Z(n850) );
  XOR U1008 ( .A(n618), .B(n851), .Z(n853) );
  IV U1009 ( .A(n616), .Z(n618) );
  XNOR U1010 ( .A(\min_dist_reg[7][2] ), .B(n854), .Z(n616) );
  NAND U1011 ( .A(n855), .B(n535), .Z(n854) );
  XNOR U1012 ( .A(\min_dist_reg[7][2] ), .B(n856), .Z(n855) );
  XNOR U1013 ( .A(n833), .B(n851), .Z(n852) );
  XOR U1014 ( .A(n857), .B(n858), .Z(n851) );
  NAND U1015 ( .A(n859), .B(n860), .Z(n858) );
  XNOR U1016 ( .A(n857), .B(n622), .Z(n860) );
  IV U1017 ( .A(n620), .Z(n622) );
  XNOR U1018 ( .A(\min_dist_reg[7][1] ), .B(n861), .Z(n620) );
  NAND U1019 ( .A(n862), .B(n535), .Z(n861) );
  XNOR U1020 ( .A(\min_dist_reg[7][1] ), .B(n863), .Z(n862) );
  XOR U1021 ( .A(n840), .B(n857), .Z(n859) );
  IV U1022 ( .A(\min_dist_reg[6][1] ), .Z(n840) );
  ANDN U1023 ( .B(n624), .A(\min_dist_reg[6][0] ), .Z(n857) );
  IV U1024 ( .A(\min_dist_reg[6][2] ), .Z(n833) );
  IV U1025 ( .A(\min_dist_reg[6][3] ), .Z(n849) );
  XOR U1026 ( .A(\min_dist_reg[6][0] ), .B(n624), .Z(n625) );
  XOR U1027 ( .A(n864), .B(n865), .Z(n624) );
  NAND U1028 ( .A(n866), .B(n535), .Z(n865) );
  XNOR U1029 ( .A(n867), .B(n868), .Z(n535) );
  AND U1030 ( .A(n869), .B(n870), .Z(n867) );
  XNOR U1031 ( .A(n871), .B(n848), .Z(n870) );
  XNOR U1032 ( .A(n872), .B(n873), .Z(n848) );
  ANDN U1033 ( .B(n874), .A(n875), .Z(n872) );
  XOR U1034 ( .A(n873), .B(n876), .Z(n874) );
  XNOR U1035 ( .A(\min_dist_reg[7][3] ), .B(n868), .Z(n869) );
  IV U1036 ( .A(n871), .Z(n868) );
  XOR U1037 ( .A(n877), .B(n878), .Z(n871) );
  AND U1038 ( .A(n879), .B(n880), .Z(n877) );
  XOR U1039 ( .A(n878), .B(n856), .Z(n880) );
  XOR U1040 ( .A(n881), .B(n876), .Z(n856) );
  XNOR U1041 ( .A(n882), .B(n883), .Z(n876) );
  ANDN U1042 ( .B(n884), .A(n885), .Z(n882) );
  XOR U1043 ( .A(n886), .B(n887), .Z(n884) );
  IV U1044 ( .A(n875), .Z(n881) );
  XOR U1045 ( .A(n888), .B(n889), .Z(n875) );
  XNOR U1046 ( .A(n890), .B(n891), .Z(n889) );
  ANDN U1047 ( .B(n892), .A(n893), .Z(n890) );
  XNOR U1048 ( .A(n894), .B(n895), .Z(n892) );
  IV U1049 ( .A(n873), .Z(n888) );
  XOR U1050 ( .A(n896), .B(n897), .Z(n873) );
  ANDN U1051 ( .B(n898), .A(n899), .Z(n896) );
  XOR U1052 ( .A(n897), .B(n900), .Z(n898) );
  XOR U1053 ( .A(\min_dist_reg[7][2] ), .B(n878), .Z(n879) );
  XOR U1054 ( .A(n901), .B(n902), .Z(n878) );
  NAND U1055 ( .A(n903), .B(n904), .Z(n902) );
  XNOR U1056 ( .A(n901), .B(n863), .Z(n904) );
  XOR U1057 ( .A(n905), .B(n900), .Z(n863) );
  XOR U1058 ( .A(n906), .B(n887), .Z(n900) );
  XNOR U1059 ( .A(n907), .B(n908), .Z(n887) );
  ANDN U1060 ( .B(n909), .A(n910), .Z(n907) );
  XNOR U1061 ( .A(n908), .B(n911), .Z(n909) );
  IV U1062 ( .A(n885), .Z(n906) );
  XOR U1063 ( .A(n883), .B(n912), .Z(n885) );
  XNOR U1064 ( .A(n913), .B(n914), .Z(n912) );
  ANDN U1065 ( .B(n915), .A(n916), .Z(n913) );
  XNOR U1066 ( .A(n917), .B(n918), .Z(n915) );
  IV U1067 ( .A(n914), .Z(n918) );
  IV U1068 ( .A(n886), .Z(n883) );
  XNOR U1069 ( .A(n919), .B(n920), .Z(n886) );
  ANDN U1070 ( .B(n921), .A(n922), .Z(n919) );
  XNOR U1071 ( .A(n920), .B(n923), .Z(n921) );
  IV U1072 ( .A(n899), .Z(n905) );
  XOR U1073 ( .A(n924), .B(n925), .Z(n899) );
  XNOR U1074 ( .A(n894), .B(n926), .Z(n925) );
  IV U1075 ( .A(n897), .Z(n926) );
  XNOR U1076 ( .A(n927), .B(n928), .Z(n897) );
  ANDN U1077 ( .B(n929), .A(n930), .Z(n927) );
  XNOR U1078 ( .A(n928), .B(n931), .Z(n929) );
  XOR U1079 ( .A(n932), .B(n933), .Z(n894) );
  ANDN U1080 ( .B(n934), .A(n935), .Z(n932) );
  XNOR U1081 ( .A(n933), .B(n936), .Z(n934) );
  IV U1082 ( .A(n893), .Z(n924) );
  XOR U1083 ( .A(n891), .B(n937), .Z(n893) );
  XNOR U1084 ( .A(n938), .B(n939), .Z(n937) );
  ANDN U1085 ( .B(n940), .A(n941), .Z(n938) );
  XNOR U1086 ( .A(n942), .B(n943), .Z(n940) );
  IV U1087 ( .A(n939), .Z(n943) );
  IV U1088 ( .A(n895), .Z(n891) );
  XNOR U1089 ( .A(n944), .B(n945), .Z(n895) );
  ANDN U1090 ( .B(n946), .A(n947), .Z(n944) );
  XNOR U1091 ( .A(n948), .B(n945), .Z(n946) );
  XNOR U1092 ( .A(\min_dist_reg[7][1] ), .B(n901), .Z(n903) );
  NOR U1093 ( .A(\min_dist_reg[7][0] ), .B(n949), .Z(n901) );
  XOR U1094 ( .A(n864), .B(n949), .Z(n866) );
  XOR U1095 ( .A(n950), .B(n931), .Z(n949) );
  XOR U1096 ( .A(n951), .B(n923), .Z(n931) );
  XOR U1097 ( .A(n952), .B(n911), .Z(n923) );
  XNOR U1098 ( .A(q[14]), .B(DB[14]), .Z(n911) );
  IV U1099 ( .A(n910), .Z(n952) );
  XOR U1100 ( .A(n908), .B(n953), .Z(n910) );
  XNOR U1101 ( .A(q[13]), .B(DB[13]), .Z(n953) );
  XOR U1102 ( .A(q[12]), .B(DB[12]), .Z(n908) );
  IV U1103 ( .A(n922), .Z(n951) );
  XOR U1104 ( .A(n954), .B(n955), .Z(n922) );
  XNOR U1105 ( .A(n917), .B(n920), .Z(n955) );
  XOR U1106 ( .A(q[8]), .B(DB[8]), .Z(n920) );
  XOR U1107 ( .A(q[11]), .B(DB[11]), .Z(n917) );
  IV U1108 ( .A(n916), .Z(n954) );
  XOR U1109 ( .A(n914), .B(n956), .Z(n916) );
  XNOR U1110 ( .A(q[10]), .B(DB[10]), .Z(n956) );
  XOR U1111 ( .A(q[9]), .B(DB[9]), .Z(n914) );
  IV U1112 ( .A(n930), .Z(n950) );
  XOR U1113 ( .A(n957), .B(n958), .Z(n930) );
  XOR U1114 ( .A(n948), .B(n928), .Z(n958) );
  XOR U1115 ( .A(q[0]), .B(DB[0]), .Z(n928) );
  XOR U1116 ( .A(n959), .B(n936), .Z(n948) );
  XNOR U1117 ( .A(q[7]), .B(DB[7]), .Z(n936) );
  IV U1118 ( .A(n935), .Z(n959) );
  XOR U1119 ( .A(n933), .B(n960), .Z(n935) );
  XNOR U1120 ( .A(q[6]), .B(DB[6]), .Z(n960) );
  XOR U1121 ( .A(q[5]), .B(DB[5]), .Z(n933) );
  IV U1122 ( .A(n947), .Z(n957) );
  XOR U1123 ( .A(n961), .B(n962), .Z(n947) );
  XNOR U1124 ( .A(n942), .B(n945), .Z(n962) );
  XOR U1125 ( .A(q[1]), .B(DB[1]), .Z(n945) );
  XOR U1126 ( .A(q[4]), .B(DB[4]), .Z(n942) );
  IV U1127 ( .A(n941), .Z(n961) );
  XOR U1128 ( .A(n939), .B(n963), .Z(n941) );
  XNOR U1129 ( .A(q[3]), .B(DB[3]), .Z(n963) );
  XOR U1130 ( .A(q[2]), .B(DB[2]), .Z(n939) );
  IV U1131 ( .A(\min_dist_reg[7][0] ), .Z(n864) );
  IV U1132 ( .A(\min_dist_reg[1][0] ), .Z(n756) );
endmodule

