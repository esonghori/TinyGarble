
module mult_N128_CC32 ( clk, rst, a, b, c );
  input [127:0] a;
  input [3:0] b;
  output [255:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014;
  wire   [255:0] sreg;

  DFF \sreg_reg[251]  ( .D(c[255]), .CLK(clk), .RST(rst), .Q(sreg[251]) );
  DFF \sreg_reg[250]  ( .D(c[254]), .CLK(clk), .RST(rst), .Q(sreg[250]) );
  DFF \sreg_reg[249]  ( .D(c[253]), .CLK(clk), .RST(rst), .Q(sreg[249]) );
  DFF \sreg_reg[248]  ( .D(c[252]), .CLK(clk), .RST(rst), .Q(sreg[248]) );
  DFF \sreg_reg[247]  ( .D(c[251]), .CLK(clk), .RST(rst), .Q(sreg[247]) );
  DFF \sreg_reg[246]  ( .D(c[250]), .CLK(clk), .RST(rst), .Q(sreg[246]) );
  DFF \sreg_reg[245]  ( .D(c[249]), .CLK(clk), .RST(rst), .Q(sreg[245]) );
  DFF \sreg_reg[244]  ( .D(c[248]), .CLK(clk), .RST(rst), .Q(sreg[244]) );
  DFF \sreg_reg[243]  ( .D(c[247]), .CLK(clk), .RST(rst), .Q(sreg[243]) );
  DFF \sreg_reg[242]  ( .D(c[246]), .CLK(clk), .RST(rst), .Q(sreg[242]) );
  DFF \sreg_reg[241]  ( .D(c[245]), .CLK(clk), .RST(rst), .Q(sreg[241]) );
  DFF \sreg_reg[240]  ( .D(c[244]), .CLK(clk), .RST(rst), .Q(sreg[240]) );
  DFF \sreg_reg[239]  ( .D(c[243]), .CLK(clk), .RST(rst), .Q(sreg[239]) );
  DFF \sreg_reg[238]  ( .D(c[242]), .CLK(clk), .RST(rst), .Q(sreg[238]) );
  DFF \sreg_reg[237]  ( .D(c[241]), .CLK(clk), .RST(rst), .Q(sreg[237]) );
  DFF \sreg_reg[236]  ( .D(c[240]), .CLK(clk), .RST(rst), .Q(sreg[236]) );
  DFF \sreg_reg[235]  ( .D(c[239]), .CLK(clk), .RST(rst), .Q(sreg[235]) );
  DFF \sreg_reg[234]  ( .D(c[238]), .CLK(clk), .RST(rst), .Q(sreg[234]) );
  DFF \sreg_reg[233]  ( .D(c[237]), .CLK(clk), .RST(rst), .Q(sreg[233]) );
  DFF \sreg_reg[232]  ( .D(c[236]), .CLK(clk), .RST(rst), .Q(sreg[232]) );
  DFF \sreg_reg[231]  ( .D(c[235]), .CLK(clk), .RST(rst), .Q(sreg[231]) );
  DFF \sreg_reg[230]  ( .D(c[234]), .CLK(clk), .RST(rst), .Q(sreg[230]) );
  DFF \sreg_reg[229]  ( .D(c[233]), .CLK(clk), .RST(rst), .Q(sreg[229]) );
  DFF \sreg_reg[228]  ( .D(c[232]), .CLK(clk), .RST(rst), .Q(sreg[228]) );
  DFF \sreg_reg[227]  ( .D(c[231]), .CLK(clk), .RST(rst), .Q(sreg[227]) );
  DFF \sreg_reg[226]  ( .D(c[230]), .CLK(clk), .RST(rst), .Q(sreg[226]) );
  DFF \sreg_reg[225]  ( .D(c[229]), .CLK(clk), .RST(rst), .Q(sreg[225]) );
  DFF \sreg_reg[224]  ( .D(c[228]), .CLK(clk), .RST(rst), .Q(sreg[224]) );
  DFF \sreg_reg[223]  ( .D(c[227]), .CLK(clk), .RST(rst), .Q(sreg[223]) );
  DFF \sreg_reg[222]  ( .D(c[226]), .CLK(clk), .RST(rst), .Q(sreg[222]) );
  DFF \sreg_reg[221]  ( .D(c[225]), .CLK(clk), .RST(rst), .Q(sreg[221]) );
  DFF \sreg_reg[220]  ( .D(c[224]), .CLK(clk), .RST(rst), .Q(sreg[220]) );
  DFF \sreg_reg[219]  ( .D(c[223]), .CLK(clk), .RST(rst), .Q(sreg[219]) );
  DFF \sreg_reg[218]  ( .D(c[222]), .CLK(clk), .RST(rst), .Q(sreg[218]) );
  DFF \sreg_reg[217]  ( .D(c[221]), .CLK(clk), .RST(rst), .Q(sreg[217]) );
  DFF \sreg_reg[216]  ( .D(c[220]), .CLK(clk), .RST(rst), .Q(sreg[216]) );
  DFF \sreg_reg[215]  ( .D(c[219]), .CLK(clk), .RST(rst), .Q(sreg[215]) );
  DFF \sreg_reg[214]  ( .D(c[218]), .CLK(clk), .RST(rst), .Q(sreg[214]) );
  DFF \sreg_reg[213]  ( .D(c[217]), .CLK(clk), .RST(rst), .Q(sreg[213]) );
  DFF \sreg_reg[212]  ( .D(c[216]), .CLK(clk), .RST(rst), .Q(sreg[212]) );
  DFF \sreg_reg[211]  ( .D(c[215]), .CLK(clk), .RST(rst), .Q(sreg[211]) );
  DFF \sreg_reg[210]  ( .D(c[214]), .CLK(clk), .RST(rst), .Q(sreg[210]) );
  DFF \sreg_reg[209]  ( .D(c[213]), .CLK(clk), .RST(rst), .Q(sreg[209]) );
  DFF \sreg_reg[208]  ( .D(c[212]), .CLK(clk), .RST(rst), .Q(sreg[208]) );
  DFF \sreg_reg[207]  ( .D(c[211]), .CLK(clk), .RST(rst), .Q(sreg[207]) );
  DFF \sreg_reg[206]  ( .D(c[210]), .CLK(clk), .RST(rst), .Q(sreg[206]) );
  DFF \sreg_reg[205]  ( .D(c[209]), .CLK(clk), .RST(rst), .Q(sreg[205]) );
  DFF \sreg_reg[204]  ( .D(c[208]), .CLK(clk), .RST(rst), .Q(sreg[204]) );
  DFF \sreg_reg[203]  ( .D(c[207]), .CLK(clk), .RST(rst), .Q(sreg[203]) );
  DFF \sreg_reg[202]  ( .D(c[206]), .CLK(clk), .RST(rst), .Q(sreg[202]) );
  DFF \sreg_reg[201]  ( .D(c[205]), .CLK(clk), .RST(rst), .Q(sreg[201]) );
  DFF \sreg_reg[200]  ( .D(c[204]), .CLK(clk), .RST(rst), .Q(sreg[200]) );
  DFF \sreg_reg[199]  ( .D(c[203]), .CLK(clk), .RST(rst), .Q(sreg[199]) );
  DFF \sreg_reg[198]  ( .D(c[202]), .CLK(clk), .RST(rst), .Q(sreg[198]) );
  DFF \sreg_reg[197]  ( .D(c[201]), .CLK(clk), .RST(rst), .Q(sreg[197]) );
  DFF \sreg_reg[196]  ( .D(c[200]), .CLK(clk), .RST(rst), .Q(sreg[196]) );
  DFF \sreg_reg[195]  ( .D(c[199]), .CLK(clk), .RST(rst), .Q(sreg[195]) );
  DFF \sreg_reg[194]  ( .D(c[198]), .CLK(clk), .RST(rst), .Q(sreg[194]) );
  DFF \sreg_reg[193]  ( .D(c[197]), .CLK(clk), .RST(rst), .Q(sreg[193]) );
  DFF \sreg_reg[192]  ( .D(c[196]), .CLK(clk), .RST(rst), .Q(sreg[192]) );
  DFF \sreg_reg[191]  ( .D(c[195]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[190]  ( .D(c[194]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[189]  ( .D(c[193]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[188]  ( .D(c[192]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[187]  ( .D(c[191]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[186]  ( .D(c[190]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[185]  ( .D(c[189]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[184]  ( .D(c[188]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[183]  ( .D(c[187]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[182]  ( .D(c[186]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[181]  ( .D(c[185]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[180]  ( .D(c[184]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[179]  ( .D(c[183]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[178]  ( .D(c[182]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[177]  ( .D(c[181]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[176]  ( .D(c[180]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[175]  ( .D(c[179]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[174]  ( .D(c[178]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[173]  ( .D(c[177]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[172]  ( .D(c[176]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[171]  ( .D(c[175]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[170]  ( .D(c[174]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[169]  ( .D(c[173]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[168]  ( .D(c[172]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[167]  ( .D(c[171]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[166]  ( .D(c[170]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[165]  ( .D(c[169]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[164]  ( .D(c[168]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[163]  ( .D(c[167]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[162]  ( .D(c[166]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[161]  ( .D(c[165]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[160]  ( .D(c[164]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[159]  ( .D(c[163]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[158]  ( .D(c[162]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[157]  ( .D(c[161]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[156]  ( .D(c[160]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[155]  ( .D(c[159]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[154]  ( .D(c[158]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[153]  ( .D(c[157]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[152]  ( .D(c[156]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[151]  ( .D(c[155]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[150]  ( .D(c[154]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[149]  ( .D(c[153]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[148]  ( .D(c[152]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[147]  ( .D(c[151]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[146]  ( .D(c[150]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[145]  ( .D(c[149]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[144]  ( .D(c[148]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[143]  ( .D(c[147]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[142]  ( .D(c[146]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[141]  ( .D(c[145]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[140]  ( .D(c[144]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[139]  ( .D(c[143]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[138]  ( .D(c[142]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[137]  ( .D(c[141]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[136]  ( .D(c[140]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[135]  ( .D(c[139]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[134]  ( .D(c[138]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[133]  ( .D(c[137]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[132]  ( .D(c[136]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[131]  ( .D(c[135]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[130]  ( .D(c[134]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[129]  ( .D(c[133]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[128]  ( .D(c[132]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[127]  ( .D(c[131]), .CLK(clk), .RST(rst), .Q(sreg[127]) );
  DFF \sreg_reg[126]  ( .D(c[130]), .CLK(clk), .RST(rst), .Q(sreg[126]) );
  DFF \sreg_reg[125]  ( .D(c[129]), .CLK(clk), .RST(rst), .Q(sreg[125]) );
  DFF \sreg_reg[124]  ( .D(c[128]), .CLK(clk), .RST(rst), .Q(sreg[124]) );
  DFF \sreg_reg[123]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[122]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[121]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[120]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[119]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[118]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[117]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[116]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[115]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[114]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[113]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[112]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[111]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[110]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[109]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[108]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[107]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[106]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[105]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[104]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[103]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[102]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[101]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[100]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[99]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[98]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[97]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[96]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[95]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[94]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[93]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[92]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[91]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[90]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[89]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[88]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[87]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[86]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[85]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[84]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[83]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[82]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[81]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[80]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[79]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[78]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[77]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[76]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[75]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[74]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[73]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[72]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[71]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[70]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[69]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[68]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[67]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[66]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[65]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[64]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[63]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[62]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[61]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[60]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[59]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[58]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[57]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[56]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[55]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[54]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[53]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[52]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[51]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[50]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[49]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[48]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[47]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[46]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[45]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[44]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[43]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[42]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[41]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[40]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[39]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[38]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[37]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[36]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[35]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[34]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[33]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[32]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[31]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[30]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[29]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[28]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[27]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[26]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[25]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[24]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[23]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[22]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[21]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[20]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[19]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[18]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[17]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[16]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[15]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[14]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[13]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[12]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[11]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[10]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[9]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[8]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[7]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[6]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[5]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[4]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[3]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[2]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[1]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[0]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[0]) );
  NAND U7 ( .A(n2340), .B(n2338), .Z(n1) );
  XOR U8 ( .A(n2338), .B(n2340), .Z(n2) );
  NANDN U9 ( .A(n2339), .B(n2), .Z(n3) );
  NAND U10 ( .A(n1), .B(n3), .Z(n2359) );
  NAND U11 ( .A(n382), .B(n381), .Z(n4) );
  XOR U12 ( .A(n381), .B(n382), .Z(n5) );
  NAND U13 ( .A(n5), .B(sreg[132]), .Z(n6) );
  NAND U14 ( .A(n4), .B(n6), .Z(n402) );
  XOR U15 ( .A(n686), .B(n685), .Z(n7) );
  NANDN U16 ( .A(sreg[146]), .B(n7), .Z(n8) );
  NAND U17 ( .A(n686), .B(n685), .Z(n9) );
  AND U18 ( .A(n8), .B(n9), .Z(n706) );
  XOR U19 ( .A(n1237), .B(sreg[171]), .Z(n10) );
  NANDN U20 ( .A(n1236), .B(n10), .Z(n11) );
  NAND U21 ( .A(n1237), .B(sreg[171]), .Z(n12) );
  AND U22 ( .A(n11), .B(n12), .Z(n1257) );
  NAND U23 ( .A(sreg[221]), .B(n2335), .Z(n13) );
  XOR U24 ( .A(n2335), .B(sreg[221]), .Z(n14) );
  NANDN U25 ( .A(n2336), .B(n14), .Z(n15) );
  NAND U26 ( .A(n13), .B(n15), .Z(n2353) );
  NAND U27 ( .A(sreg[239]), .B(n2718), .Z(n16) );
  XOR U28 ( .A(n2718), .B(sreg[239]), .Z(n17) );
  NANDN U29 ( .A(n2719), .B(n17), .Z(n18) );
  NAND U30 ( .A(n16), .B(n18), .Z(n2739) );
  NAND U31 ( .A(b[1]), .B(a[125]), .Z(n2946) );
  OR U32 ( .A(n2966), .B(n2926), .Z(n19) );
  NANDN U33 ( .A(n2928), .B(n2927), .Z(n20) );
  AND U34 ( .A(n19), .B(n20), .Z(n2954) );
  NANDN U35 ( .A(n1683), .B(n1682), .Z(n21) );
  NANDN U36 ( .A(n1684), .B(n1685), .Z(n22) );
  NAND U37 ( .A(n21), .B(n22), .Z(n1692) );
  NAND U38 ( .A(n2391), .B(n2390), .Z(n23) );
  XOR U39 ( .A(n2390), .B(n2391), .Z(n24) );
  NANDN U40 ( .A(n2392), .B(n24), .Z(n25) );
  NAND U41 ( .A(n23), .B(n25), .Z(n2396) );
  NANDN U42 ( .A(n2404), .B(n2403), .Z(n26) );
  NANDN U43 ( .A(n2405), .B(n2406), .Z(n27) );
  NAND U44 ( .A(n26), .B(n27), .Z(n2418) );
  XOR U45 ( .A(n1613), .B(n1612), .Z(n28) );
  NANDN U46 ( .A(n1611), .B(n28), .Z(n29) );
  NAND U47 ( .A(n1613), .B(n1612), .Z(n30) );
  AND U48 ( .A(n29), .B(n30), .Z(n1634) );
  NAND U49 ( .A(n361), .B(n360), .Z(n31) );
  XOR U50 ( .A(n360), .B(n361), .Z(n32) );
  NAND U51 ( .A(n32), .B(sreg[131]), .Z(n33) );
  NAND U52 ( .A(n31), .B(n33), .Z(n381) );
  NAND U53 ( .A(n427), .B(n426), .Z(n34) );
  XOR U54 ( .A(n426), .B(n427), .Z(n35) );
  NAND U55 ( .A(n35), .B(sreg[135]), .Z(n36) );
  NAND U56 ( .A(n34), .B(n36), .Z(n465) );
  NAND U57 ( .A(sreg[144]), .B(n643), .Z(n37) );
  XOR U58 ( .A(n643), .B(sreg[144]), .Z(n38) );
  NANDN U59 ( .A(n644), .B(n38), .Z(n39) );
  NAND U60 ( .A(n37), .B(n39), .Z(n664) );
  NAND U61 ( .A(sreg[148]), .B(n727), .Z(n40) );
  XOR U62 ( .A(n727), .B(sreg[148]), .Z(n41) );
  NANDN U63 ( .A(n728), .B(n41), .Z(n42) );
  NAND U64 ( .A(n40), .B(n42), .Z(n730) );
  XOR U65 ( .A(n925), .B(sreg[157]), .Z(n43) );
  NANDN U66 ( .A(n924), .B(n43), .Z(n44) );
  NAND U67 ( .A(n925), .B(sreg[157]), .Z(n45) );
  AND U68 ( .A(n44), .B(n45), .Z(n927) );
  XOR U69 ( .A(n1258), .B(n1257), .Z(n46) );
  NANDN U70 ( .A(sreg[172]), .B(n46), .Z(n47) );
  NAND U71 ( .A(n1258), .B(n1257), .Z(n48) );
  AND U72 ( .A(n47), .B(n48), .Z(n1278) );
  NAND U73 ( .A(n1388), .B(n1387), .Z(n49) );
  XOR U74 ( .A(n1387), .B(n1388), .Z(n50) );
  NAND U75 ( .A(n50), .B(sreg[178]), .Z(n51) );
  NAND U76 ( .A(n49), .B(n51), .Z(n1390) );
  NAND U77 ( .A(sreg[188]), .B(n1608), .Z(n52) );
  XOR U78 ( .A(n1608), .B(sreg[188]), .Z(n53) );
  NANDN U79 ( .A(n1609), .B(n53), .Z(n54) );
  NAND U80 ( .A(n52), .B(n54), .Z(n1626) );
  XOR U81 ( .A(n2072), .B(sreg[210]), .Z(n55) );
  NAND U82 ( .A(n55), .B(n2071), .Z(n56) );
  NAND U83 ( .A(n2072), .B(sreg[210]), .Z(n57) );
  AND U84 ( .A(n56), .B(n57), .Z(n2111) );
  NAND U85 ( .A(n2354), .B(sreg[222]), .Z(n58) );
  XOR U86 ( .A(sreg[222]), .B(n2354), .Z(n59) );
  NAND U87 ( .A(n59), .B(n2353), .Z(n60) );
  NAND U88 ( .A(n58), .B(n60), .Z(n2375) );
  XOR U89 ( .A(sreg[230]), .B(n2501), .Z(n61) );
  NANDN U90 ( .A(n2502), .B(n61), .Z(n62) );
  NAND U91 ( .A(sreg[230]), .B(n2501), .Z(n63) );
  AND U92 ( .A(n62), .B(n63), .Z(n2541) );
  XOR U93 ( .A(n2760), .B(sreg[241]), .Z(n64) );
  NANDN U94 ( .A(n2761), .B(n64), .Z(n65) );
  NAND U95 ( .A(n2760), .B(sreg[241]), .Z(n66) );
  AND U96 ( .A(n65), .B(n66), .Z(n2763) );
  AND U97 ( .A(b[0]), .B(a[1]), .Z(n282) );
  NAND U98 ( .A(n1674), .B(n1673), .Z(n67) );
  XOR U99 ( .A(n1673), .B(n1674), .Z(n68) );
  NANDN U100 ( .A(n1675), .B(n68), .Z(n69) );
  NAND U101 ( .A(n67), .B(n69), .Z(n1693) );
  NANDN U102 ( .A(n2382), .B(n2383), .Z(n70) );
  NANDN U103 ( .A(n2381), .B(n2380), .Z(n71) );
  AND U104 ( .A(n70), .B(n71), .Z(n2394) );
  OR U105 ( .A(n2951), .B(n2952), .Z(n72) );
  NAND U106 ( .A(n2953), .B(n2954), .Z(n73) );
  AND U107 ( .A(n72), .B(n73), .Z(n2960) );
  XOR U108 ( .A(sreg[217]), .B(n2242), .Z(n74) );
  NANDN U109 ( .A(n2243), .B(n74), .Z(n75) );
  NAND U110 ( .A(sreg[217]), .B(n2242), .Z(n76) );
  AND U111 ( .A(n75), .B(n76), .Z(n2264) );
  XOR U112 ( .A(n340), .B(n339), .Z(n77) );
  NANDN U113 ( .A(sreg[130]), .B(n77), .Z(n78) );
  NAND U114 ( .A(n340), .B(n339), .Z(n79) );
  AND U115 ( .A(n78), .B(n79), .Z(n360) );
  NAND U116 ( .A(n424), .B(n423), .Z(n80) );
  XOR U117 ( .A(n423), .B(n424), .Z(n81) );
  NAND U118 ( .A(n81), .B(sreg[134]), .Z(n82) );
  NAND U119 ( .A(n80), .B(n82), .Z(n426) );
  NAND U120 ( .A(n492), .B(n491), .Z(n83) );
  XOR U121 ( .A(n491), .B(n492), .Z(n84) );
  NANDN U122 ( .A(sreg[138]), .B(n84), .Z(n85) );
  NAND U123 ( .A(n83), .B(n85), .Z(n513) );
  NAND U124 ( .A(sreg[143]), .B(n622), .Z(n86) );
  XOR U125 ( .A(n622), .B(sreg[143]), .Z(n87) );
  NANDN U126 ( .A(n623), .B(n87), .Z(n88) );
  NAND U127 ( .A(n86), .B(n88), .Z(n643) );
  NAND U128 ( .A(sreg[147]), .B(n706), .Z(n89) );
  XOR U129 ( .A(n706), .B(sreg[147]), .Z(n90) );
  NANDN U130 ( .A(n707), .B(n90), .Z(n91) );
  NAND U131 ( .A(n89), .B(n91), .Z(n727) );
  NAND U132 ( .A(n775), .B(sreg[151]), .Z(n92) );
  XOR U133 ( .A(sreg[151]), .B(n775), .Z(n93) );
  NANDN U134 ( .A(n774), .B(n93), .Z(n94) );
  NAND U135 ( .A(n92), .B(n94), .Z(n796) );
  XOR U136 ( .A(sreg[155]), .B(n862), .Z(n95) );
  NANDN U137 ( .A(n863), .B(n95), .Z(n96) );
  NAND U138 ( .A(sreg[155]), .B(n862), .Z(n97) );
  AND U139 ( .A(n96), .B(n97), .Z(n902) );
  XOR U140 ( .A(sreg[160]), .B(n971), .Z(n98) );
  NANDN U141 ( .A(n972), .B(n98), .Z(n99) );
  NAND U142 ( .A(sreg[160]), .B(n971), .Z(n100) );
  AND U143 ( .A(n99), .B(n100), .Z(n1011) );
  XOR U144 ( .A(sreg[174]), .B(n1281), .Z(n101) );
  NANDN U145 ( .A(n1282), .B(n101), .Z(n102) );
  NAND U146 ( .A(sreg[174]), .B(n1281), .Z(n103) );
  AND U147 ( .A(n102), .B(n103), .Z(n1321) );
  NAND U148 ( .A(n1391), .B(n1390), .Z(n104) );
  XOR U149 ( .A(n1390), .B(n1391), .Z(n105) );
  NAND U150 ( .A(n105), .B(sreg[179]), .Z(n106) );
  NAND U151 ( .A(n104), .B(n106), .Z(n1430) );
  XOR U152 ( .A(sreg[183]), .B(n1478), .Z(n107) );
  NANDN U153 ( .A(n1479), .B(n107), .Z(n108) );
  NAND U154 ( .A(sreg[183]), .B(n1478), .Z(n109) );
  AND U155 ( .A(n108), .B(n109), .Z(n1518) );
  XOR U156 ( .A(n1627), .B(n1626), .Z(n110) );
  NAND U157 ( .A(n110), .B(sreg[189]), .Z(n111) );
  NAND U158 ( .A(n1627), .B(n1626), .Z(n112) );
  AND U159 ( .A(n111), .B(n112), .Z(n1629) );
  XOR U160 ( .A(sreg[196]), .B(n1759), .Z(n113) );
  NANDN U161 ( .A(n1760), .B(n113), .Z(n114) );
  NAND U162 ( .A(sreg[196]), .B(n1759), .Z(n115) );
  AND U163 ( .A(n114), .B(n115), .Z(n1799) );
  XOR U164 ( .A(sreg[200]), .B(n1847), .Z(n116) );
  NANDN U165 ( .A(n1848), .B(n116), .Z(n117) );
  NAND U166 ( .A(sreg[200]), .B(n1847), .Z(n118) );
  AND U167 ( .A(n117), .B(n118), .Z(n1887) );
  NAND U168 ( .A(n2137), .B(n2136), .Z(n119) );
  XOR U169 ( .A(n2136), .B(n2137), .Z(n120) );
  NAND U170 ( .A(n120), .B(sreg[213]), .Z(n121) );
  NAND U171 ( .A(n119), .B(n121), .Z(n2175) );
  NAND U172 ( .A(n2376), .B(sreg[223]), .Z(n122) );
  XOR U173 ( .A(sreg[223]), .B(n2376), .Z(n123) );
  NAND U174 ( .A(n123), .B(n2375), .Z(n124) );
  NAND U175 ( .A(n122), .B(n124), .Z(n2378) );
  NAND U176 ( .A(n2455), .B(n2454), .Z(n125) );
  XOR U177 ( .A(n2454), .B(n2455), .Z(n126) );
  NAND U178 ( .A(n126), .B(sreg[227]), .Z(n127) );
  NAND U179 ( .A(n125), .B(n127), .Z(n2457) );
  NAND U180 ( .A(n2567), .B(n2566), .Z(n128) );
  XOR U181 ( .A(n2566), .B(n2567), .Z(n129) );
  NAND U182 ( .A(n129), .B(sreg[233]), .Z(n130) );
  NAND U183 ( .A(n128), .B(n130), .Z(n2605) );
  XOR U184 ( .A(n2764), .B(sreg[242]), .Z(n131) );
  NANDN U185 ( .A(n2763), .B(n131), .Z(n132) );
  NAND U186 ( .A(n2764), .B(sreg[242]), .Z(n133) );
  AND U187 ( .A(n132), .B(n133), .Z(n2803) );
  XOR U188 ( .A(sreg[247]), .B(n2874), .Z(n134) );
  NANDN U189 ( .A(n2875), .B(n134), .Z(n135) );
  NAND U190 ( .A(sreg[247]), .B(n2874), .Z(n136) );
  AND U191 ( .A(n135), .B(n136), .Z(n2914) );
  NAND U192 ( .A(b[2]), .B(a[2]), .Z(n285) );
  XOR U193 ( .A(n306), .B(n307), .Z(n308) );
  NAND U194 ( .A(n2396), .B(n2394), .Z(n137) );
  XOR U195 ( .A(n2394), .B(n2396), .Z(n138) );
  NAND U196 ( .A(n138), .B(n2395), .Z(n139) );
  NAND U197 ( .A(n137), .B(n139), .Z(n2419) );
  NANDN U198 ( .A(n2973), .B(n2974), .Z(n140) );
  NANDN U199 ( .A(n2972), .B(n2971), .Z(n141) );
  AND U200 ( .A(n140), .B(n141), .Z(n2977) );
  OR U201 ( .A(n247), .B(n248), .Z(n142) );
  NAND U202 ( .A(n245), .B(n246), .Z(n143) );
  AND U203 ( .A(n142), .B(n143), .Z(n257) );
  NANDN U204 ( .A(n2942), .B(n2943), .Z(n144) );
  NANDN U205 ( .A(n2940), .B(n2941), .Z(n145) );
  NAND U206 ( .A(n144), .B(n145), .Z(n2962) );
  NANDN U207 ( .A(n2984), .B(n2983), .Z(n146) );
  NANDN U208 ( .A(n2985), .B(n2986), .Z(n147) );
  NAND U209 ( .A(n146), .B(n147), .Z(n2989) );
  XOR U210 ( .A(n319), .B(sreg[129]), .Z(n148) );
  NANDN U211 ( .A(n318), .B(n148), .Z(n149) );
  NAND U212 ( .A(n319), .B(sreg[129]), .Z(n150) );
  AND U213 ( .A(n149), .B(n150), .Z(n339) );
  NAND U214 ( .A(n403), .B(n402), .Z(n151) );
  XOR U215 ( .A(n402), .B(n403), .Z(n152) );
  NAND U216 ( .A(n152), .B(sreg[133]), .Z(n153) );
  NAND U217 ( .A(n151), .B(n153), .Z(n423) );
  XOR U218 ( .A(n489), .B(sreg[137]), .Z(n154) );
  NANDN U219 ( .A(n488), .B(n154), .Z(n155) );
  NAND U220 ( .A(n489), .B(sreg[137]), .Z(n156) );
  AND U221 ( .A(n155), .B(n156), .Z(n491) );
  XOR U222 ( .A(sreg[141]), .B(n560), .Z(n157) );
  NANDN U223 ( .A(n561), .B(n157), .Z(n158) );
  NAND U224 ( .A(sreg[141]), .B(n560), .Z(n159) );
  AND U225 ( .A(n158), .B(n159), .Z(n600) );
  XOR U226 ( .A(n665), .B(n664), .Z(n160) );
  NAND U227 ( .A(n160), .B(sreg[145]), .Z(n161) );
  NAND U228 ( .A(n665), .B(n664), .Z(n162) );
  AND U229 ( .A(n161), .B(n162), .Z(n685) );
  XOR U230 ( .A(sreg[149]), .B(n730), .Z(n163) );
  NANDN U231 ( .A(n731), .B(n163), .Z(n164) );
  NAND U232 ( .A(sreg[149]), .B(n730), .Z(n165) );
  AND U233 ( .A(n164), .B(n165), .Z(n770) );
  NAND U234 ( .A(sreg[154]), .B(n859), .Z(n166) );
  XOR U235 ( .A(n859), .B(sreg[154]), .Z(n167) );
  NANDN U236 ( .A(n860), .B(n167), .Z(n168) );
  NAND U237 ( .A(n166), .B(n168), .Z(n862) );
  NAND U238 ( .A(n928), .B(n927), .Z(n169) );
  XOR U239 ( .A(n927), .B(n928), .Z(n170) );
  NANDN U240 ( .A(sreg[158]), .B(n170), .Z(n171) );
  NAND U241 ( .A(n169), .B(n171), .Z(n967) );
  XOR U242 ( .A(sreg[162]), .B(n1015), .Z(n172) );
  NANDN U243 ( .A(n1016), .B(n172), .Z(n173) );
  NAND U244 ( .A(sreg[162]), .B(n1015), .Z(n174) );
  AND U245 ( .A(n173), .B(n174), .Z(n1055) );
  XOR U246 ( .A(sreg[169]), .B(n1174), .Z(n175) );
  NANDN U247 ( .A(n1175), .B(n175), .Z(n176) );
  NAND U248 ( .A(sreg[169]), .B(n1174), .Z(n177) );
  AND U249 ( .A(n176), .B(n177), .Z(n1214) );
  NAND U250 ( .A(sreg[173]), .B(n1278), .Z(n178) );
  XOR U251 ( .A(n1278), .B(sreg[173]), .Z(n179) );
  NANDN U252 ( .A(n1279), .B(n179), .Z(n180) );
  NAND U253 ( .A(n178), .B(n180), .Z(n1281) );
  NAND U254 ( .A(n1367), .B(n1366), .Z(n181) );
  XOR U255 ( .A(n1366), .B(n1367), .Z(n182) );
  NAND U256 ( .A(n182), .B(sreg[177]), .Z(n183) );
  NAND U257 ( .A(n181), .B(n183), .Z(n1387) );
  XOR U258 ( .A(sreg[181]), .B(n1434), .Z(n184) );
  NANDN U259 ( .A(n1435), .B(n184), .Z(n185) );
  NAND U260 ( .A(sreg[181]), .B(n1434), .Z(n186) );
  AND U261 ( .A(n185), .B(n186), .Z(n1474) );
  NAND U262 ( .A(n1523), .B(sreg[185]), .Z(n187) );
  XOR U263 ( .A(sreg[185]), .B(n1523), .Z(n188) );
  NANDN U264 ( .A(n1522), .B(n188), .Z(n189) );
  NAND U265 ( .A(n187), .B(n189), .Z(n1561) );
  XOR U266 ( .A(n1630), .B(sreg[190]), .Z(n190) );
  NANDN U267 ( .A(n1629), .B(n190), .Z(n191) );
  NAND U268 ( .A(n1630), .B(sreg[190]), .Z(n192) );
  AND U269 ( .A(n191), .B(n192), .Z(n1670) );
  NAND U270 ( .A(n1716), .B(sreg[194]), .Z(n193) );
  XOR U271 ( .A(sreg[194]), .B(n1716), .Z(n194) );
  NANDN U272 ( .A(n1715), .B(n194), .Z(n195) );
  NAND U273 ( .A(n193), .B(n195), .Z(n1754) );
  NAND U274 ( .A(sreg[199]), .B(n1844), .Z(n196) );
  XOR U275 ( .A(n1844), .B(sreg[199]), .Z(n197) );
  NANDN U276 ( .A(n1845), .B(n197), .Z(n198) );
  NAND U277 ( .A(n196), .B(n198), .Z(n1847) );
  NAND U278 ( .A(n1915), .B(sreg[203]), .Z(n199) );
  XOR U279 ( .A(sreg[203]), .B(n1915), .Z(n200) );
  NANDN U280 ( .A(n1914), .B(n200), .Z(n201) );
  NAND U281 ( .A(n199), .B(n201), .Z(n1953) );
  XOR U282 ( .A(sreg[207]), .B(n2004), .Z(n202) );
  NANDN U283 ( .A(n2005), .B(n202), .Z(n203) );
  NAND U284 ( .A(sreg[207]), .B(n2004), .Z(n204) );
  AND U285 ( .A(n203), .B(n204), .Z(n2044) );
  XOR U286 ( .A(n2134), .B(n2133), .Z(n205) );
  NANDN U287 ( .A(sreg[212]), .B(n205), .Z(n206) );
  NAND U288 ( .A(n2134), .B(n2133), .Z(n207) );
  AND U289 ( .A(n206), .B(n207), .Z(n2136) );
  NAND U290 ( .A(n2222), .B(sreg[216]), .Z(n208) );
  XOR U291 ( .A(sreg[216]), .B(n2222), .Z(n209) );
  NAND U292 ( .A(n209), .B(n2221), .Z(n210) );
  NAND U293 ( .A(n208), .B(n210), .Z(n2242) );
  XOR U294 ( .A(sreg[224]), .B(n2378), .Z(n211) );
  NANDN U295 ( .A(n2379), .B(n211), .Z(n212) );
  NAND U296 ( .A(sreg[224]), .B(n2378), .Z(n213) );
  AND U297 ( .A(n212), .B(n213), .Z(n2409) );
  NAND U298 ( .A(n2458), .B(n2457), .Z(n214) );
  XOR U299 ( .A(n2457), .B(n2458), .Z(n215) );
  NAND U300 ( .A(n215), .B(sreg[228]), .Z(n216) );
  NAND U301 ( .A(n214), .B(n216), .Z(n2478) );
  NAND U302 ( .A(sreg[232]), .B(n2563), .Z(n217) );
  XOR U303 ( .A(n2563), .B(sreg[232]), .Z(n218) );
  NANDN U304 ( .A(n2564), .B(n218), .Z(n219) );
  NAND U305 ( .A(n217), .B(n219), .Z(n2566) );
  XOR U306 ( .A(sreg[236]), .B(n2633), .Z(n220) );
  NANDN U307 ( .A(n2634), .B(n220), .Z(n221) );
  NAND U308 ( .A(sreg[236]), .B(n2633), .Z(n222) );
  AND U309 ( .A(n221), .B(n222), .Z(n2673) );
  NAND U310 ( .A(n2740), .B(n2739), .Z(n223) );
  XOR U311 ( .A(n2739), .B(n2740), .Z(n224) );
  NAND U312 ( .A(n224), .B(sreg[240]), .Z(n225) );
  NAND U313 ( .A(n223), .B(n225), .Z(n2760) );
  XOR U314 ( .A(n2808), .B(n2807), .Z(n226) );
  NANDN U315 ( .A(sreg[244]), .B(n226), .Z(n227) );
  NAND U316 ( .A(n2808), .B(n2807), .Z(n228) );
  AND U317 ( .A(n227), .B(n228), .Z(n2846) );
  XOR U318 ( .A(n2919), .B(sreg[249]), .Z(n229) );
  NAND U319 ( .A(n229), .B(n2918), .Z(n230) );
  NAND U320 ( .A(n2919), .B(sreg[249]), .Z(n231) );
  AND U321 ( .A(n230), .B(n231), .Z(n2937) );
  IV U322 ( .A(b[1]), .Z(n232) );
  IV U323 ( .A(b[3]), .Z(n233) );
  NAND U324 ( .A(b[0]), .B(a[0]), .Z(n241) );
  XNOR U325 ( .A(n241), .B(sreg[124]), .Z(c[124]) );
  AND U326 ( .A(a[1]), .B(b[0]), .Z(n235) );
  NAND U327 ( .A(b[1]), .B(a[0]), .Z(n234) );
  XNOR U328 ( .A(n235), .B(n234), .Z(n236) );
  XNOR U329 ( .A(sreg[125]), .B(n236), .Z(n238) );
  NANDN U330 ( .A(n241), .B(sreg[124]), .Z(n237) );
  XOR U331 ( .A(n238), .B(n237), .Z(c[125]) );
  NAND U332 ( .A(n236), .B(sreg[125]), .Z(n240) );
  OR U333 ( .A(n238), .B(n237), .Z(n239) );
  NAND U334 ( .A(n240), .B(n239), .Z(n251) );
  ANDN U335 ( .B(a[1]), .A(n232), .Z(n265) );
  ANDN U336 ( .B(n265), .A(n241), .Z(n247) );
  NAND U337 ( .A(a[0]), .B(b[2]), .Z(n246) );
  NAND U338 ( .A(b[0]), .B(a[2]), .Z(n266) );
  XOR U339 ( .A(n266), .B(n265), .Z(n245) );
  XNOR U340 ( .A(n246), .B(n245), .Z(n248) );
  XOR U341 ( .A(n247), .B(n248), .Z(n250) );
  IV U342 ( .A(n250), .Z(n249) );
  XOR U343 ( .A(n249), .B(sreg[126]), .Z(n242) );
  XOR U344 ( .A(n251), .B(n242), .Z(c[126]) );
  ANDN U345 ( .B(a[2]), .A(n282), .Z(n243) );
  NAND U346 ( .A(b[1]), .B(n243), .Z(n268) );
  NAND U347 ( .A(b[3]), .B(a[0]), .Z(n267) );
  XOR U348 ( .A(n268), .B(n267), .Z(n255) );
  AND U349 ( .A(a[3]), .B(b[0]), .Z(n289) );
  NAND U350 ( .A(b[2]), .B(a[1]), .Z(n244) );
  XNOR U351 ( .A(n289), .B(n244), .Z(n256) );
  XNOR U352 ( .A(n255), .B(n256), .Z(n258) );
  XNOR U353 ( .A(n258), .B(n257), .Z(n272) );
  NAND U354 ( .A(n249), .B(sreg[126]), .Z(n254) );
  ANDN U355 ( .B(n250), .A(sreg[126]), .Z(n252) );
  NANDN U356 ( .A(n252), .B(n251), .Z(n253) );
  NAND U357 ( .A(n254), .B(n253), .Z(n271) );
  XNOR U358 ( .A(n271), .B(sreg[127]), .Z(n273) );
  XNOR U359 ( .A(n272), .B(n273), .Z(c[127]) );
  NAND U360 ( .A(n256), .B(n255), .Z(n260) );
  NANDN U361 ( .A(n258), .B(n257), .Z(n259) );
  NAND U362 ( .A(n260), .B(n259), .Z(n279) );
  AND U363 ( .A(b[2]), .B(a[3]), .Z(n309) );
  NAND U364 ( .A(b[0]), .B(n309), .Z(n261) );
  XNOR U365 ( .A(b[3]), .B(n261), .Z(n262) );
  NAND U366 ( .A(a[1]), .B(n262), .Z(n286) );
  XNOR U367 ( .A(n285), .B(n286), .Z(n291) );
  AND U368 ( .A(a[4]), .B(b[0]), .Z(n264) );
  NAND U369 ( .A(b[1]), .B(a[3]), .Z(n263) );
  XNOR U370 ( .A(n264), .B(n263), .Z(n290) );
  XNOR U371 ( .A(n291), .B(n290), .Z(n276) );
  NANDN U372 ( .A(n266), .B(n265), .Z(n270) );
  OR U373 ( .A(n268), .B(n267), .Z(n269) );
  NAND U374 ( .A(n270), .B(n269), .Z(n277) );
  XOR U375 ( .A(n276), .B(n277), .Z(n278) );
  XOR U376 ( .A(n279), .B(n278), .Z(n294) );
  XNOR U377 ( .A(n294), .B(sreg[128]), .Z(n296) );
  NAND U378 ( .A(sreg[127]), .B(n271), .Z(n275) );
  NANDN U379 ( .A(n273), .B(n272), .Z(n274) );
  AND U380 ( .A(n275), .B(n274), .Z(n295) );
  XOR U381 ( .A(n296), .B(n295), .Z(c[128]) );
  OR U382 ( .A(n277), .B(n276), .Z(n281) );
  NANDN U383 ( .A(n279), .B(n278), .Z(n280) );
  NAND U384 ( .A(n281), .B(n280), .Z(n303) );
  ANDN U385 ( .B(a[4]), .A(n232), .Z(n306) );
  AND U386 ( .A(b[3]), .B(a[2]), .Z(n307) );
  XNOR U387 ( .A(n309), .B(n308), .Z(n312) );
  NAND U388 ( .A(b[0]), .B(a[5]), .Z(n313) );
  XOR U389 ( .A(n312), .B(n313), .Z(n314) );
  NAND U390 ( .A(n309), .B(n282), .Z(n284) );
  NAND U391 ( .A(b[3]), .B(a[1]), .Z(n283) );
  AND U392 ( .A(n284), .B(n283), .Z(n288) );
  NANDN U393 ( .A(n286), .B(n285), .Z(n287) );
  NANDN U394 ( .A(n288), .B(n287), .Z(n315) );
  XOR U395 ( .A(n314), .B(n315), .Z(n300) );
  NAND U396 ( .A(n306), .B(n289), .Z(n293) );
  NANDN U397 ( .A(n291), .B(n290), .Z(n292) );
  NAND U398 ( .A(n293), .B(n292), .Z(n301) );
  XNOR U399 ( .A(n300), .B(n301), .Z(n302) );
  XNOR U400 ( .A(n303), .B(n302), .Z(n319) );
  NAND U401 ( .A(n294), .B(sreg[128]), .Z(n298) );
  OR U402 ( .A(n296), .B(n295), .Z(n297) );
  AND U403 ( .A(n298), .B(n297), .Z(n318) );
  XNOR U404 ( .A(n318), .B(sreg[129]), .Z(n299) );
  XOR U405 ( .A(n319), .B(n299), .Z(c[129]) );
  NANDN U406 ( .A(n301), .B(n300), .Z(n305) );
  NAND U407 ( .A(n303), .B(n302), .Z(n304) );
  NAND U408 ( .A(n305), .B(n304), .Z(n324) );
  AND U409 ( .A(b[2]), .B(a[4]), .Z(n330) );
  AND U410 ( .A(a[5]), .B(b[1]), .Z(n328) );
  AND U411 ( .A(a[3]), .B(b[3]), .Z(n327) );
  XOR U412 ( .A(n328), .B(n327), .Z(n329) );
  XOR U413 ( .A(n330), .B(n329), .Z(n333) );
  NAND U414 ( .A(b[0]), .B(a[6]), .Z(n334) );
  XOR U415 ( .A(n333), .B(n334), .Z(n336) );
  OR U416 ( .A(n307), .B(n306), .Z(n311) );
  NANDN U417 ( .A(n309), .B(n308), .Z(n310) );
  NAND U418 ( .A(n311), .B(n310), .Z(n335) );
  XNOR U419 ( .A(n336), .B(n335), .Z(n321) );
  OR U420 ( .A(n313), .B(n312), .Z(n317) );
  NANDN U421 ( .A(n315), .B(n314), .Z(n316) );
  NAND U422 ( .A(n317), .B(n316), .Z(n322) );
  XNOR U423 ( .A(n321), .B(n322), .Z(n323) );
  XOR U424 ( .A(n324), .B(n323), .Z(n340) );
  XOR U425 ( .A(sreg[130]), .B(n339), .Z(n320) );
  XOR U426 ( .A(n340), .B(n320), .Z(c[130]) );
  NANDN U427 ( .A(n322), .B(n321), .Z(n326) );
  NAND U428 ( .A(n324), .B(n323), .Z(n325) );
  NAND U429 ( .A(n326), .B(n325), .Z(n345) );
  AND U430 ( .A(b[2]), .B(a[5]), .Z(n351) );
  AND U431 ( .A(a[6]), .B(b[1]), .Z(n349) );
  AND U432 ( .A(a[4]), .B(b[3]), .Z(n348) );
  XOR U433 ( .A(n349), .B(n348), .Z(n350) );
  XOR U434 ( .A(n351), .B(n350), .Z(n354) );
  NAND U435 ( .A(b[0]), .B(a[7]), .Z(n355) );
  XOR U436 ( .A(n354), .B(n355), .Z(n357) );
  OR U437 ( .A(n328), .B(n327), .Z(n332) );
  NANDN U438 ( .A(n330), .B(n329), .Z(n331) );
  NAND U439 ( .A(n332), .B(n331), .Z(n356) );
  XNOR U440 ( .A(n357), .B(n356), .Z(n342) );
  NANDN U441 ( .A(n334), .B(n333), .Z(n338) );
  OR U442 ( .A(n336), .B(n335), .Z(n337) );
  NAND U443 ( .A(n338), .B(n337), .Z(n343) );
  XNOR U444 ( .A(n342), .B(n343), .Z(n344) );
  XNOR U445 ( .A(n345), .B(n344), .Z(n361) );
  XOR U446 ( .A(n360), .B(sreg[131]), .Z(n341) );
  XOR U447 ( .A(n361), .B(n341), .Z(c[131]) );
  NANDN U448 ( .A(n343), .B(n342), .Z(n347) );
  NAND U449 ( .A(n345), .B(n344), .Z(n346) );
  NAND U450 ( .A(n347), .B(n346), .Z(n366) );
  AND U451 ( .A(b[2]), .B(a[6]), .Z(n372) );
  AND U452 ( .A(a[7]), .B(b[1]), .Z(n370) );
  AND U453 ( .A(a[5]), .B(b[3]), .Z(n369) );
  XOR U454 ( .A(n370), .B(n369), .Z(n371) );
  XOR U455 ( .A(n372), .B(n371), .Z(n375) );
  NAND U456 ( .A(b[0]), .B(a[8]), .Z(n376) );
  XOR U457 ( .A(n375), .B(n376), .Z(n378) );
  OR U458 ( .A(n349), .B(n348), .Z(n353) );
  NANDN U459 ( .A(n351), .B(n350), .Z(n352) );
  NAND U460 ( .A(n353), .B(n352), .Z(n377) );
  XNOR U461 ( .A(n378), .B(n377), .Z(n363) );
  NANDN U462 ( .A(n355), .B(n354), .Z(n359) );
  OR U463 ( .A(n357), .B(n356), .Z(n358) );
  NAND U464 ( .A(n359), .B(n358), .Z(n364) );
  XNOR U465 ( .A(n363), .B(n364), .Z(n365) );
  XNOR U466 ( .A(n366), .B(n365), .Z(n382) );
  XOR U467 ( .A(n381), .B(sreg[132]), .Z(n362) );
  XOR U468 ( .A(n382), .B(n362), .Z(c[132]) );
  NANDN U469 ( .A(n364), .B(n363), .Z(n368) );
  NAND U470 ( .A(n366), .B(n365), .Z(n367) );
  NAND U471 ( .A(n368), .B(n367), .Z(n387) );
  AND U472 ( .A(b[2]), .B(a[7]), .Z(n393) );
  AND U473 ( .A(a[8]), .B(b[1]), .Z(n391) );
  AND U474 ( .A(a[6]), .B(b[3]), .Z(n390) );
  XOR U475 ( .A(n391), .B(n390), .Z(n392) );
  XOR U476 ( .A(n393), .B(n392), .Z(n396) );
  NAND U477 ( .A(b[0]), .B(a[9]), .Z(n397) );
  XOR U478 ( .A(n396), .B(n397), .Z(n399) );
  OR U479 ( .A(n370), .B(n369), .Z(n374) );
  NANDN U480 ( .A(n372), .B(n371), .Z(n373) );
  NAND U481 ( .A(n374), .B(n373), .Z(n398) );
  XNOR U482 ( .A(n399), .B(n398), .Z(n384) );
  NANDN U483 ( .A(n376), .B(n375), .Z(n380) );
  OR U484 ( .A(n378), .B(n377), .Z(n379) );
  NAND U485 ( .A(n380), .B(n379), .Z(n385) );
  XNOR U486 ( .A(n384), .B(n385), .Z(n386) );
  XNOR U487 ( .A(n387), .B(n386), .Z(n403) );
  XOR U488 ( .A(n402), .B(sreg[133]), .Z(n383) );
  XOR U489 ( .A(n403), .B(n383), .Z(c[133]) );
  NANDN U490 ( .A(n385), .B(n384), .Z(n389) );
  NAND U491 ( .A(n387), .B(n386), .Z(n388) );
  NAND U492 ( .A(n389), .B(n388), .Z(n408) );
  AND U493 ( .A(b[2]), .B(a[8]), .Z(n414) );
  AND U494 ( .A(a[9]), .B(b[1]), .Z(n412) );
  AND U495 ( .A(a[7]), .B(b[3]), .Z(n411) );
  XOR U496 ( .A(n412), .B(n411), .Z(n413) );
  XOR U497 ( .A(n414), .B(n413), .Z(n417) );
  NAND U498 ( .A(b[0]), .B(a[10]), .Z(n418) );
  XOR U499 ( .A(n417), .B(n418), .Z(n420) );
  OR U500 ( .A(n391), .B(n390), .Z(n395) );
  NANDN U501 ( .A(n393), .B(n392), .Z(n394) );
  NAND U502 ( .A(n395), .B(n394), .Z(n419) );
  XNOR U503 ( .A(n420), .B(n419), .Z(n405) );
  NANDN U504 ( .A(n397), .B(n396), .Z(n401) );
  OR U505 ( .A(n399), .B(n398), .Z(n400) );
  NAND U506 ( .A(n401), .B(n400), .Z(n406) );
  XNOR U507 ( .A(n405), .B(n406), .Z(n407) );
  XNOR U508 ( .A(n408), .B(n407), .Z(n424) );
  XOR U509 ( .A(n423), .B(sreg[134]), .Z(n404) );
  XOR U510 ( .A(n424), .B(n404), .Z(c[134]) );
  NANDN U511 ( .A(n406), .B(n405), .Z(n410) );
  NAND U512 ( .A(n408), .B(n407), .Z(n409) );
  NAND U513 ( .A(n410), .B(n409), .Z(n431) );
  AND U514 ( .A(b[2]), .B(a[9]), .Z(n437) );
  AND U515 ( .A(a[10]), .B(b[1]), .Z(n435) );
  AND U516 ( .A(a[8]), .B(b[3]), .Z(n434) );
  XOR U517 ( .A(n435), .B(n434), .Z(n436) );
  XOR U518 ( .A(n437), .B(n436), .Z(n440) );
  NAND U519 ( .A(b[0]), .B(a[11]), .Z(n441) );
  XOR U520 ( .A(n440), .B(n441), .Z(n443) );
  OR U521 ( .A(n412), .B(n411), .Z(n416) );
  NANDN U522 ( .A(n414), .B(n413), .Z(n415) );
  NAND U523 ( .A(n416), .B(n415), .Z(n442) );
  XNOR U524 ( .A(n443), .B(n442), .Z(n428) );
  NANDN U525 ( .A(n418), .B(n417), .Z(n422) );
  OR U526 ( .A(n420), .B(n419), .Z(n421) );
  NAND U527 ( .A(n422), .B(n421), .Z(n429) );
  XNOR U528 ( .A(n428), .B(n429), .Z(n430) );
  XNOR U529 ( .A(n431), .B(n430), .Z(n427) );
  XOR U530 ( .A(n426), .B(sreg[135]), .Z(n425) );
  XOR U531 ( .A(n427), .B(n425), .Z(c[135]) );
  NANDN U532 ( .A(n429), .B(n428), .Z(n433) );
  NAND U533 ( .A(n431), .B(n430), .Z(n432) );
  NAND U534 ( .A(n433), .B(n432), .Z(n449) );
  AND U535 ( .A(b[2]), .B(a[10]), .Z(n455) );
  AND U536 ( .A(a[11]), .B(b[1]), .Z(n453) );
  AND U537 ( .A(a[9]), .B(b[3]), .Z(n452) );
  XOR U538 ( .A(n453), .B(n452), .Z(n454) );
  XOR U539 ( .A(n455), .B(n454), .Z(n458) );
  NAND U540 ( .A(b[0]), .B(a[12]), .Z(n459) );
  XOR U541 ( .A(n458), .B(n459), .Z(n461) );
  OR U542 ( .A(n435), .B(n434), .Z(n439) );
  NANDN U543 ( .A(n437), .B(n436), .Z(n438) );
  NAND U544 ( .A(n439), .B(n438), .Z(n460) );
  XNOR U545 ( .A(n461), .B(n460), .Z(n446) );
  NANDN U546 ( .A(n441), .B(n440), .Z(n445) );
  OR U547 ( .A(n443), .B(n442), .Z(n444) );
  NAND U548 ( .A(n445), .B(n444), .Z(n447) );
  XNOR U549 ( .A(n446), .B(n447), .Z(n448) );
  XNOR U550 ( .A(n449), .B(n448), .Z(n464) );
  XNOR U551 ( .A(n464), .B(sreg[136]), .Z(n466) );
  XNOR U552 ( .A(n465), .B(n466), .Z(c[136]) );
  NANDN U553 ( .A(n447), .B(n446), .Z(n451) );
  NAND U554 ( .A(n449), .B(n448), .Z(n450) );
  NAND U555 ( .A(n451), .B(n450), .Z(n473) );
  AND U556 ( .A(b[2]), .B(a[11]), .Z(n479) );
  AND U557 ( .A(a[12]), .B(b[1]), .Z(n477) );
  AND U558 ( .A(a[10]), .B(b[3]), .Z(n476) );
  XOR U559 ( .A(n477), .B(n476), .Z(n478) );
  XOR U560 ( .A(n479), .B(n478), .Z(n482) );
  NAND U561 ( .A(b[0]), .B(a[13]), .Z(n483) );
  XOR U562 ( .A(n482), .B(n483), .Z(n485) );
  OR U563 ( .A(n453), .B(n452), .Z(n457) );
  NANDN U564 ( .A(n455), .B(n454), .Z(n456) );
  NAND U565 ( .A(n457), .B(n456), .Z(n484) );
  XNOR U566 ( .A(n485), .B(n484), .Z(n470) );
  NANDN U567 ( .A(n459), .B(n458), .Z(n463) );
  OR U568 ( .A(n461), .B(n460), .Z(n462) );
  NAND U569 ( .A(n463), .B(n462), .Z(n471) );
  XNOR U570 ( .A(n470), .B(n471), .Z(n472) );
  XNOR U571 ( .A(n473), .B(n472), .Z(n489) );
  NAND U572 ( .A(n464), .B(sreg[136]), .Z(n468) );
  NANDN U573 ( .A(n466), .B(n465), .Z(n467) );
  AND U574 ( .A(n468), .B(n467), .Z(n488) );
  XNOR U575 ( .A(n488), .B(sreg[137]), .Z(n469) );
  XOR U576 ( .A(n489), .B(n469), .Z(c[137]) );
  NANDN U577 ( .A(n471), .B(n470), .Z(n475) );
  NAND U578 ( .A(n473), .B(n472), .Z(n474) );
  NAND U579 ( .A(n475), .B(n474), .Z(n508) );
  AND U580 ( .A(b[2]), .B(a[12]), .Z(n502) );
  AND U581 ( .A(a[13]), .B(b[1]), .Z(n500) );
  AND U582 ( .A(a[11]), .B(b[3]), .Z(n499) );
  XOR U583 ( .A(n500), .B(n499), .Z(n501) );
  XOR U584 ( .A(n502), .B(n501), .Z(n493) );
  NAND U585 ( .A(b[0]), .B(a[14]), .Z(n494) );
  XOR U586 ( .A(n493), .B(n494), .Z(n496) );
  OR U587 ( .A(n477), .B(n476), .Z(n481) );
  NANDN U588 ( .A(n479), .B(n478), .Z(n480) );
  NAND U589 ( .A(n481), .B(n480), .Z(n495) );
  XNOR U590 ( .A(n496), .B(n495), .Z(n505) );
  NANDN U591 ( .A(n483), .B(n482), .Z(n487) );
  OR U592 ( .A(n485), .B(n484), .Z(n486) );
  NAND U593 ( .A(n487), .B(n486), .Z(n506) );
  XNOR U594 ( .A(n505), .B(n506), .Z(n507) );
  XOR U595 ( .A(n508), .B(n507), .Z(n492) );
  XOR U596 ( .A(sreg[138]), .B(n491), .Z(n490) );
  XOR U597 ( .A(n492), .B(n490), .Z(c[138]) );
  NANDN U598 ( .A(n494), .B(n493), .Z(n498) );
  OR U599 ( .A(n496), .B(n495), .Z(n497) );
  NAND U600 ( .A(n498), .B(n497), .Z(n516) );
  AND U601 ( .A(b[2]), .B(a[13]), .Z(n525) );
  AND U602 ( .A(a[14]), .B(b[1]), .Z(n523) );
  AND U603 ( .A(a[12]), .B(b[3]), .Z(n522) );
  XOR U604 ( .A(n523), .B(n522), .Z(n524) );
  XOR U605 ( .A(n525), .B(n524), .Z(n528) );
  NAND U606 ( .A(b[0]), .B(a[15]), .Z(n529) );
  XNOR U607 ( .A(n528), .B(n529), .Z(n530) );
  OR U608 ( .A(n500), .B(n499), .Z(n504) );
  NANDN U609 ( .A(n502), .B(n501), .Z(n503) );
  AND U610 ( .A(n504), .B(n503), .Z(n531) );
  XNOR U611 ( .A(n530), .B(n531), .Z(n517) );
  XNOR U612 ( .A(n516), .B(n517), .Z(n518) );
  NANDN U613 ( .A(n506), .B(n505), .Z(n510) );
  NAND U614 ( .A(n508), .B(n507), .Z(n509) );
  AND U615 ( .A(n510), .B(n509), .Z(n519) );
  XOR U616 ( .A(n518), .B(n519), .Z(n511) );
  XNOR U617 ( .A(sreg[139]), .B(n511), .Z(n512) );
  XOR U618 ( .A(n513), .B(n512), .Z(c[139]) );
  NAND U619 ( .A(sreg[139]), .B(n511), .Z(n515) );
  OR U620 ( .A(n513), .B(n512), .Z(n514) );
  AND U621 ( .A(n515), .B(n514), .Z(n555) );
  IV U622 ( .A(sreg[140]), .Z(n553) );
  NANDN U623 ( .A(n517), .B(n516), .Z(n521) );
  NAND U624 ( .A(n519), .B(n518), .Z(n520) );
  NAND U625 ( .A(n521), .B(n520), .Z(n538) );
  AND U626 ( .A(b[2]), .B(a[14]), .Z(n544) );
  AND U627 ( .A(a[15]), .B(b[1]), .Z(n542) );
  AND U628 ( .A(a[13]), .B(b[3]), .Z(n541) );
  XOR U629 ( .A(n542), .B(n541), .Z(n543) );
  XOR U630 ( .A(n544), .B(n543), .Z(n547) );
  NAND U631 ( .A(b[0]), .B(a[16]), .Z(n548) );
  XOR U632 ( .A(n547), .B(n548), .Z(n550) );
  OR U633 ( .A(n523), .B(n522), .Z(n527) );
  NANDN U634 ( .A(n525), .B(n524), .Z(n526) );
  NAND U635 ( .A(n527), .B(n526), .Z(n549) );
  XNOR U636 ( .A(n550), .B(n549), .Z(n535) );
  NANDN U637 ( .A(n529), .B(n528), .Z(n533) );
  NAND U638 ( .A(n531), .B(n530), .Z(n532) );
  NAND U639 ( .A(n533), .B(n532), .Z(n536) );
  XNOR U640 ( .A(n535), .B(n536), .Z(n537) );
  XOR U641 ( .A(n538), .B(n537), .Z(n554) );
  XOR U642 ( .A(n553), .B(n554), .Z(n534) );
  XOR U643 ( .A(n555), .B(n534), .Z(c[140]) );
  NANDN U644 ( .A(n536), .B(n535), .Z(n540) );
  NANDN U645 ( .A(n538), .B(n537), .Z(n539) );
  NAND U646 ( .A(n540), .B(n539), .Z(n565) );
  AND U647 ( .A(b[2]), .B(a[15]), .Z(n571) );
  AND U648 ( .A(a[16]), .B(b[1]), .Z(n569) );
  AND U649 ( .A(a[14]), .B(b[3]), .Z(n568) );
  XOR U650 ( .A(n569), .B(n568), .Z(n570) );
  XOR U651 ( .A(n571), .B(n570), .Z(n574) );
  NAND U652 ( .A(b[0]), .B(a[17]), .Z(n575) );
  XOR U653 ( .A(n574), .B(n575), .Z(n577) );
  OR U654 ( .A(n542), .B(n541), .Z(n546) );
  NANDN U655 ( .A(n544), .B(n543), .Z(n545) );
  NAND U656 ( .A(n546), .B(n545), .Z(n576) );
  XNOR U657 ( .A(n577), .B(n576), .Z(n562) );
  NANDN U658 ( .A(n548), .B(n547), .Z(n552) );
  OR U659 ( .A(n550), .B(n549), .Z(n551) );
  NAND U660 ( .A(n552), .B(n551), .Z(n563) );
  XNOR U661 ( .A(n562), .B(n563), .Z(n564) );
  XOR U662 ( .A(n565), .B(n564), .Z(n561) );
  NANDN U663 ( .A(n554), .B(n553), .Z(n558) );
  AND U664 ( .A(n554), .B(sreg[140]), .Z(n556) );
  NANDN U665 ( .A(n556), .B(n555), .Z(n557) );
  AND U666 ( .A(n558), .B(n557), .Z(n560) );
  XNOR U667 ( .A(sreg[141]), .B(n560), .Z(n559) );
  XOR U668 ( .A(n561), .B(n559), .Z(c[141]) );
  NANDN U669 ( .A(n563), .B(n562), .Z(n567) );
  NAND U670 ( .A(n565), .B(n564), .Z(n566) );
  NAND U671 ( .A(n567), .B(n566), .Z(n583) );
  AND U672 ( .A(b[2]), .B(a[16]), .Z(n589) );
  AND U673 ( .A(a[17]), .B(b[1]), .Z(n587) );
  AND U674 ( .A(a[15]), .B(b[3]), .Z(n586) );
  XOR U675 ( .A(n587), .B(n586), .Z(n588) );
  XOR U676 ( .A(n589), .B(n588), .Z(n592) );
  NAND U677 ( .A(b[0]), .B(a[18]), .Z(n593) );
  XOR U678 ( .A(n592), .B(n593), .Z(n595) );
  OR U679 ( .A(n569), .B(n568), .Z(n573) );
  NANDN U680 ( .A(n571), .B(n570), .Z(n572) );
  NAND U681 ( .A(n573), .B(n572), .Z(n594) );
  XNOR U682 ( .A(n595), .B(n594), .Z(n580) );
  NANDN U683 ( .A(n575), .B(n574), .Z(n579) );
  OR U684 ( .A(n577), .B(n576), .Z(n578) );
  NAND U685 ( .A(n579), .B(n578), .Z(n581) );
  XNOR U686 ( .A(n580), .B(n581), .Z(n582) );
  XNOR U687 ( .A(n583), .B(n582), .Z(n598) );
  XNOR U688 ( .A(n598), .B(sreg[142]), .Z(n599) );
  XOR U689 ( .A(n600), .B(n599), .Z(c[142]) );
  NANDN U690 ( .A(n581), .B(n580), .Z(n585) );
  NAND U691 ( .A(n583), .B(n582), .Z(n584) );
  NAND U692 ( .A(n585), .B(n584), .Z(n607) );
  AND U693 ( .A(b[2]), .B(a[17]), .Z(n613) );
  AND U694 ( .A(a[18]), .B(b[1]), .Z(n611) );
  AND U695 ( .A(a[16]), .B(b[3]), .Z(n610) );
  XOR U696 ( .A(n611), .B(n610), .Z(n612) );
  XOR U697 ( .A(n613), .B(n612), .Z(n616) );
  NAND U698 ( .A(b[0]), .B(a[19]), .Z(n617) );
  XOR U699 ( .A(n616), .B(n617), .Z(n619) );
  OR U700 ( .A(n587), .B(n586), .Z(n591) );
  NANDN U701 ( .A(n589), .B(n588), .Z(n590) );
  NAND U702 ( .A(n591), .B(n590), .Z(n618) );
  XNOR U703 ( .A(n619), .B(n618), .Z(n604) );
  NANDN U704 ( .A(n593), .B(n592), .Z(n597) );
  OR U705 ( .A(n595), .B(n594), .Z(n596) );
  NAND U706 ( .A(n597), .B(n596), .Z(n605) );
  XNOR U707 ( .A(n604), .B(n605), .Z(n606) );
  XOR U708 ( .A(n607), .B(n606), .Z(n623) );
  NAND U709 ( .A(n598), .B(sreg[142]), .Z(n602) );
  OR U710 ( .A(n600), .B(n599), .Z(n601) );
  NAND U711 ( .A(n602), .B(n601), .Z(n622) );
  XNOR U712 ( .A(sreg[143]), .B(n622), .Z(n603) );
  XOR U713 ( .A(n623), .B(n603), .Z(c[143]) );
  NANDN U714 ( .A(n605), .B(n604), .Z(n609) );
  NAND U715 ( .A(n607), .B(n606), .Z(n608) );
  NAND U716 ( .A(n609), .B(n608), .Z(n628) );
  AND U717 ( .A(b[2]), .B(a[18]), .Z(n634) );
  AND U718 ( .A(a[19]), .B(b[1]), .Z(n632) );
  AND U719 ( .A(a[17]), .B(b[3]), .Z(n631) );
  XOR U720 ( .A(n632), .B(n631), .Z(n633) );
  XOR U721 ( .A(n634), .B(n633), .Z(n637) );
  NAND U722 ( .A(b[0]), .B(a[20]), .Z(n638) );
  XOR U723 ( .A(n637), .B(n638), .Z(n640) );
  OR U724 ( .A(n611), .B(n610), .Z(n615) );
  NANDN U725 ( .A(n613), .B(n612), .Z(n614) );
  NAND U726 ( .A(n615), .B(n614), .Z(n639) );
  XNOR U727 ( .A(n640), .B(n639), .Z(n625) );
  NANDN U728 ( .A(n617), .B(n616), .Z(n621) );
  OR U729 ( .A(n619), .B(n618), .Z(n620) );
  NAND U730 ( .A(n621), .B(n620), .Z(n626) );
  XNOR U731 ( .A(n625), .B(n626), .Z(n627) );
  XOR U732 ( .A(n628), .B(n627), .Z(n644) );
  XNOR U733 ( .A(sreg[144]), .B(n643), .Z(n624) );
  XOR U734 ( .A(n644), .B(n624), .Z(c[144]) );
  NANDN U735 ( .A(n626), .B(n625), .Z(n630) );
  NAND U736 ( .A(n628), .B(n627), .Z(n629) );
  NAND U737 ( .A(n630), .B(n629), .Z(n649) );
  AND U738 ( .A(b[2]), .B(a[19]), .Z(n655) );
  AND U739 ( .A(a[20]), .B(b[1]), .Z(n653) );
  AND U740 ( .A(a[18]), .B(b[3]), .Z(n652) );
  XOR U741 ( .A(n653), .B(n652), .Z(n654) );
  XOR U742 ( .A(n655), .B(n654), .Z(n658) );
  NAND U743 ( .A(b[0]), .B(a[21]), .Z(n659) );
  XOR U744 ( .A(n658), .B(n659), .Z(n661) );
  OR U745 ( .A(n632), .B(n631), .Z(n636) );
  NANDN U746 ( .A(n634), .B(n633), .Z(n635) );
  NAND U747 ( .A(n636), .B(n635), .Z(n660) );
  XNOR U748 ( .A(n661), .B(n660), .Z(n646) );
  NANDN U749 ( .A(n638), .B(n637), .Z(n642) );
  OR U750 ( .A(n640), .B(n639), .Z(n641) );
  NAND U751 ( .A(n642), .B(n641), .Z(n647) );
  XNOR U752 ( .A(n646), .B(n647), .Z(n648) );
  XNOR U753 ( .A(n649), .B(n648), .Z(n665) );
  XOR U754 ( .A(n664), .B(sreg[145]), .Z(n645) );
  XOR U755 ( .A(n665), .B(n645), .Z(c[145]) );
  NANDN U756 ( .A(n647), .B(n646), .Z(n651) );
  NAND U757 ( .A(n649), .B(n648), .Z(n650) );
  NAND U758 ( .A(n651), .B(n650), .Z(n670) );
  AND U759 ( .A(b[2]), .B(a[20]), .Z(n676) );
  AND U760 ( .A(a[21]), .B(b[1]), .Z(n674) );
  AND U761 ( .A(a[19]), .B(b[3]), .Z(n673) );
  XOR U762 ( .A(n674), .B(n673), .Z(n675) );
  XOR U763 ( .A(n676), .B(n675), .Z(n679) );
  NAND U764 ( .A(b[0]), .B(a[22]), .Z(n680) );
  XOR U765 ( .A(n679), .B(n680), .Z(n682) );
  OR U766 ( .A(n653), .B(n652), .Z(n657) );
  NANDN U767 ( .A(n655), .B(n654), .Z(n656) );
  NAND U768 ( .A(n657), .B(n656), .Z(n681) );
  XNOR U769 ( .A(n682), .B(n681), .Z(n667) );
  NANDN U770 ( .A(n659), .B(n658), .Z(n663) );
  OR U771 ( .A(n661), .B(n660), .Z(n662) );
  NAND U772 ( .A(n663), .B(n662), .Z(n668) );
  XNOR U773 ( .A(n667), .B(n668), .Z(n669) );
  XOR U774 ( .A(n670), .B(n669), .Z(n686) );
  XOR U775 ( .A(sreg[146]), .B(n685), .Z(n666) );
  XOR U776 ( .A(n686), .B(n666), .Z(c[146]) );
  NANDN U777 ( .A(n668), .B(n667), .Z(n672) );
  NAND U778 ( .A(n670), .B(n669), .Z(n671) );
  NAND U779 ( .A(n672), .B(n671), .Z(n691) );
  AND U780 ( .A(b[2]), .B(a[21]), .Z(n697) );
  AND U781 ( .A(a[22]), .B(b[1]), .Z(n695) );
  AND U782 ( .A(a[20]), .B(b[3]), .Z(n694) );
  XOR U783 ( .A(n695), .B(n694), .Z(n696) );
  XOR U784 ( .A(n697), .B(n696), .Z(n700) );
  NAND U785 ( .A(b[0]), .B(a[23]), .Z(n701) );
  XOR U786 ( .A(n700), .B(n701), .Z(n703) );
  OR U787 ( .A(n674), .B(n673), .Z(n678) );
  NANDN U788 ( .A(n676), .B(n675), .Z(n677) );
  NAND U789 ( .A(n678), .B(n677), .Z(n702) );
  XNOR U790 ( .A(n703), .B(n702), .Z(n688) );
  NANDN U791 ( .A(n680), .B(n679), .Z(n684) );
  OR U792 ( .A(n682), .B(n681), .Z(n683) );
  NAND U793 ( .A(n684), .B(n683), .Z(n689) );
  XNOR U794 ( .A(n688), .B(n689), .Z(n690) );
  XOR U795 ( .A(n691), .B(n690), .Z(n707) );
  XNOR U796 ( .A(sreg[147]), .B(n706), .Z(n687) );
  XOR U797 ( .A(n707), .B(n687), .Z(c[147]) );
  NANDN U798 ( .A(n689), .B(n688), .Z(n693) );
  NAND U799 ( .A(n691), .B(n690), .Z(n692) );
  NAND U800 ( .A(n693), .B(n692), .Z(n712) );
  AND U801 ( .A(b[2]), .B(a[22]), .Z(n718) );
  AND U802 ( .A(a[23]), .B(b[1]), .Z(n716) );
  AND U803 ( .A(a[21]), .B(b[3]), .Z(n715) );
  XOR U804 ( .A(n716), .B(n715), .Z(n717) );
  XOR U805 ( .A(n718), .B(n717), .Z(n721) );
  NAND U806 ( .A(b[0]), .B(a[24]), .Z(n722) );
  XOR U807 ( .A(n721), .B(n722), .Z(n724) );
  OR U808 ( .A(n695), .B(n694), .Z(n699) );
  NANDN U809 ( .A(n697), .B(n696), .Z(n698) );
  NAND U810 ( .A(n699), .B(n698), .Z(n723) );
  XNOR U811 ( .A(n724), .B(n723), .Z(n709) );
  NANDN U812 ( .A(n701), .B(n700), .Z(n705) );
  OR U813 ( .A(n703), .B(n702), .Z(n704) );
  NAND U814 ( .A(n705), .B(n704), .Z(n710) );
  XNOR U815 ( .A(n709), .B(n710), .Z(n711) );
  XOR U816 ( .A(n712), .B(n711), .Z(n728) );
  XNOR U817 ( .A(sreg[148]), .B(n727), .Z(n708) );
  XOR U818 ( .A(n728), .B(n708), .Z(c[148]) );
  NANDN U819 ( .A(n710), .B(n709), .Z(n714) );
  NAND U820 ( .A(n712), .B(n711), .Z(n713) );
  NAND U821 ( .A(n714), .B(n713), .Z(n735) );
  AND U822 ( .A(b[2]), .B(a[23]), .Z(n741) );
  AND U823 ( .A(a[24]), .B(b[1]), .Z(n739) );
  AND U824 ( .A(a[22]), .B(b[3]), .Z(n738) );
  XOR U825 ( .A(n739), .B(n738), .Z(n740) );
  XOR U826 ( .A(n741), .B(n740), .Z(n744) );
  NAND U827 ( .A(b[0]), .B(a[25]), .Z(n745) );
  XOR U828 ( .A(n744), .B(n745), .Z(n747) );
  OR U829 ( .A(n716), .B(n715), .Z(n720) );
  NANDN U830 ( .A(n718), .B(n717), .Z(n719) );
  NAND U831 ( .A(n720), .B(n719), .Z(n746) );
  XNOR U832 ( .A(n747), .B(n746), .Z(n732) );
  NANDN U833 ( .A(n722), .B(n721), .Z(n726) );
  OR U834 ( .A(n724), .B(n723), .Z(n725) );
  NAND U835 ( .A(n726), .B(n725), .Z(n733) );
  XNOR U836 ( .A(n732), .B(n733), .Z(n734) );
  XOR U837 ( .A(n735), .B(n734), .Z(n731) );
  XNOR U838 ( .A(sreg[149]), .B(n730), .Z(n729) );
  XOR U839 ( .A(n731), .B(n729), .Z(c[149]) );
  NANDN U840 ( .A(n733), .B(n732), .Z(n737) );
  NAND U841 ( .A(n735), .B(n734), .Z(n736) );
  NAND U842 ( .A(n737), .B(n736), .Z(n753) );
  AND U843 ( .A(b[2]), .B(a[24]), .Z(n759) );
  AND U844 ( .A(a[25]), .B(b[1]), .Z(n757) );
  AND U845 ( .A(a[23]), .B(b[3]), .Z(n756) );
  XOR U846 ( .A(n757), .B(n756), .Z(n758) );
  XOR U847 ( .A(n759), .B(n758), .Z(n762) );
  NAND U848 ( .A(b[0]), .B(a[26]), .Z(n763) );
  XOR U849 ( .A(n762), .B(n763), .Z(n765) );
  OR U850 ( .A(n739), .B(n738), .Z(n743) );
  NANDN U851 ( .A(n741), .B(n740), .Z(n742) );
  NAND U852 ( .A(n743), .B(n742), .Z(n764) );
  XNOR U853 ( .A(n765), .B(n764), .Z(n750) );
  NANDN U854 ( .A(n745), .B(n744), .Z(n749) );
  OR U855 ( .A(n747), .B(n746), .Z(n748) );
  NAND U856 ( .A(n749), .B(n748), .Z(n751) );
  XNOR U857 ( .A(n750), .B(n751), .Z(n752) );
  XNOR U858 ( .A(n753), .B(n752), .Z(n768) );
  XNOR U859 ( .A(n768), .B(sreg[150]), .Z(n769) );
  XOR U860 ( .A(n770), .B(n769), .Z(c[150]) );
  NANDN U861 ( .A(n751), .B(n750), .Z(n755) );
  NAND U862 ( .A(n753), .B(n752), .Z(n754) );
  NAND U863 ( .A(n755), .B(n754), .Z(n779) );
  AND U864 ( .A(b[2]), .B(a[25]), .Z(n785) );
  AND U865 ( .A(a[26]), .B(b[1]), .Z(n783) );
  AND U866 ( .A(a[24]), .B(b[3]), .Z(n782) );
  XOR U867 ( .A(n783), .B(n782), .Z(n784) );
  XOR U868 ( .A(n785), .B(n784), .Z(n788) );
  NAND U869 ( .A(b[0]), .B(a[27]), .Z(n789) );
  XOR U870 ( .A(n788), .B(n789), .Z(n791) );
  OR U871 ( .A(n757), .B(n756), .Z(n761) );
  NANDN U872 ( .A(n759), .B(n758), .Z(n760) );
  NAND U873 ( .A(n761), .B(n760), .Z(n790) );
  XNOR U874 ( .A(n791), .B(n790), .Z(n776) );
  NANDN U875 ( .A(n763), .B(n762), .Z(n767) );
  OR U876 ( .A(n765), .B(n764), .Z(n766) );
  NAND U877 ( .A(n767), .B(n766), .Z(n777) );
  XNOR U878 ( .A(n776), .B(n777), .Z(n778) );
  XNOR U879 ( .A(n779), .B(n778), .Z(n775) );
  NAND U880 ( .A(n768), .B(sreg[150]), .Z(n772) );
  OR U881 ( .A(n770), .B(n769), .Z(n771) );
  AND U882 ( .A(n772), .B(n771), .Z(n774) );
  XNOR U883 ( .A(n774), .B(sreg[151]), .Z(n773) );
  XOR U884 ( .A(n775), .B(n773), .Z(c[151]) );
  NANDN U885 ( .A(n777), .B(n776), .Z(n781) );
  NAND U886 ( .A(n779), .B(n778), .Z(n780) );
  NAND U887 ( .A(n781), .B(n780), .Z(n802) );
  AND U888 ( .A(b[2]), .B(a[26]), .Z(n808) );
  AND U889 ( .A(a[27]), .B(b[1]), .Z(n806) );
  AND U890 ( .A(a[25]), .B(b[3]), .Z(n805) );
  XOR U891 ( .A(n806), .B(n805), .Z(n807) );
  XOR U892 ( .A(n808), .B(n807), .Z(n811) );
  NAND U893 ( .A(b[0]), .B(a[28]), .Z(n812) );
  XOR U894 ( .A(n811), .B(n812), .Z(n814) );
  OR U895 ( .A(n783), .B(n782), .Z(n787) );
  NANDN U896 ( .A(n785), .B(n784), .Z(n786) );
  NAND U897 ( .A(n787), .B(n786), .Z(n813) );
  XNOR U898 ( .A(n814), .B(n813), .Z(n799) );
  NANDN U899 ( .A(n789), .B(n788), .Z(n793) );
  OR U900 ( .A(n791), .B(n790), .Z(n792) );
  NAND U901 ( .A(n793), .B(n792), .Z(n800) );
  XNOR U902 ( .A(n799), .B(n800), .Z(n801) );
  XNOR U903 ( .A(n802), .B(n801), .Z(n794) );
  XOR U904 ( .A(sreg[152]), .B(n794), .Z(n795) );
  XOR U905 ( .A(n796), .B(n795), .Z(c[152]) );
  OR U906 ( .A(n794), .B(sreg[152]), .Z(n798) );
  NANDN U907 ( .A(n796), .B(n795), .Z(n797) );
  NAND U908 ( .A(n798), .B(n797), .Z(n837) );
  NANDN U909 ( .A(n800), .B(n799), .Z(n804) );
  NAND U910 ( .A(n802), .B(n801), .Z(n803) );
  NAND U911 ( .A(n804), .B(n803), .Z(n820) );
  AND U912 ( .A(b[2]), .B(a[27]), .Z(n826) );
  AND U913 ( .A(a[28]), .B(b[1]), .Z(n824) );
  AND U914 ( .A(a[26]), .B(b[3]), .Z(n823) );
  XOR U915 ( .A(n824), .B(n823), .Z(n825) );
  XOR U916 ( .A(n826), .B(n825), .Z(n829) );
  NAND U917 ( .A(b[0]), .B(a[29]), .Z(n830) );
  XOR U918 ( .A(n829), .B(n830), .Z(n832) );
  OR U919 ( .A(n806), .B(n805), .Z(n810) );
  NANDN U920 ( .A(n808), .B(n807), .Z(n809) );
  NAND U921 ( .A(n810), .B(n809), .Z(n831) );
  XNOR U922 ( .A(n832), .B(n831), .Z(n817) );
  NANDN U923 ( .A(n812), .B(n811), .Z(n816) );
  OR U924 ( .A(n814), .B(n813), .Z(n815) );
  NAND U925 ( .A(n816), .B(n815), .Z(n818) );
  XNOR U926 ( .A(n817), .B(n818), .Z(n819) );
  XNOR U927 ( .A(n820), .B(n819), .Z(n835) );
  XNOR U928 ( .A(n835), .B(sreg[153]), .Z(n836) );
  XOR U929 ( .A(n837), .B(n836), .Z(c[153]) );
  NANDN U930 ( .A(n818), .B(n817), .Z(n822) );
  NAND U931 ( .A(n820), .B(n819), .Z(n821) );
  NAND U932 ( .A(n822), .B(n821), .Z(n844) );
  AND U933 ( .A(b[2]), .B(a[28]), .Z(n850) );
  AND U934 ( .A(a[29]), .B(b[1]), .Z(n848) );
  AND U935 ( .A(a[27]), .B(b[3]), .Z(n847) );
  XOR U936 ( .A(n848), .B(n847), .Z(n849) );
  XOR U937 ( .A(n850), .B(n849), .Z(n853) );
  NAND U938 ( .A(b[0]), .B(a[30]), .Z(n854) );
  XOR U939 ( .A(n853), .B(n854), .Z(n856) );
  OR U940 ( .A(n824), .B(n823), .Z(n828) );
  NANDN U941 ( .A(n826), .B(n825), .Z(n827) );
  NAND U942 ( .A(n828), .B(n827), .Z(n855) );
  XNOR U943 ( .A(n856), .B(n855), .Z(n841) );
  NANDN U944 ( .A(n830), .B(n829), .Z(n834) );
  OR U945 ( .A(n832), .B(n831), .Z(n833) );
  NAND U946 ( .A(n834), .B(n833), .Z(n842) );
  XNOR U947 ( .A(n841), .B(n842), .Z(n843) );
  XOR U948 ( .A(n844), .B(n843), .Z(n860) );
  NAND U949 ( .A(n835), .B(sreg[153]), .Z(n839) );
  OR U950 ( .A(n837), .B(n836), .Z(n838) );
  NAND U951 ( .A(n839), .B(n838), .Z(n859) );
  XNOR U952 ( .A(sreg[154]), .B(n859), .Z(n840) );
  XOR U953 ( .A(n860), .B(n840), .Z(c[154]) );
  NANDN U954 ( .A(n842), .B(n841), .Z(n846) );
  NAND U955 ( .A(n844), .B(n843), .Z(n845) );
  NAND U956 ( .A(n846), .B(n845), .Z(n867) );
  AND U957 ( .A(b[2]), .B(a[29]), .Z(n873) );
  AND U958 ( .A(a[30]), .B(b[1]), .Z(n871) );
  AND U959 ( .A(a[28]), .B(b[3]), .Z(n870) );
  XOR U960 ( .A(n871), .B(n870), .Z(n872) );
  XOR U961 ( .A(n873), .B(n872), .Z(n876) );
  NAND U962 ( .A(b[0]), .B(a[31]), .Z(n877) );
  XOR U963 ( .A(n876), .B(n877), .Z(n879) );
  OR U964 ( .A(n848), .B(n847), .Z(n852) );
  NANDN U965 ( .A(n850), .B(n849), .Z(n851) );
  NAND U966 ( .A(n852), .B(n851), .Z(n878) );
  XNOR U967 ( .A(n879), .B(n878), .Z(n864) );
  NANDN U968 ( .A(n854), .B(n853), .Z(n858) );
  OR U969 ( .A(n856), .B(n855), .Z(n857) );
  NAND U970 ( .A(n858), .B(n857), .Z(n865) );
  XNOR U971 ( .A(n864), .B(n865), .Z(n866) );
  XOR U972 ( .A(n867), .B(n866), .Z(n863) );
  XNOR U973 ( .A(sreg[155]), .B(n862), .Z(n861) );
  XOR U974 ( .A(n863), .B(n861), .Z(c[155]) );
  NANDN U975 ( .A(n865), .B(n864), .Z(n869) );
  NAND U976 ( .A(n867), .B(n866), .Z(n868) );
  NAND U977 ( .A(n869), .B(n868), .Z(n885) );
  AND U978 ( .A(b[2]), .B(a[30]), .Z(n891) );
  AND U979 ( .A(a[31]), .B(b[1]), .Z(n889) );
  AND U980 ( .A(a[29]), .B(b[3]), .Z(n888) );
  XOR U981 ( .A(n889), .B(n888), .Z(n890) );
  XOR U982 ( .A(n891), .B(n890), .Z(n894) );
  NAND U983 ( .A(b[0]), .B(a[32]), .Z(n895) );
  XOR U984 ( .A(n894), .B(n895), .Z(n897) );
  OR U985 ( .A(n871), .B(n870), .Z(n875) );
  NANDN U986 ( .A(n873), .B(n872), .Z(n874) );
  NAND U987 ( .A(n875), .B(n874), .Z(n896) );
  XNOR U988 ( .A(n897), .B(n896), .Z(n882) );
  NANDN U989 ( .A(n877), .B(n876), .Z(n881) );
  OR U990 ( .A(n879), .B(n878), .Z(n880) );
  NAND U991 ( .A(n881), .B(n880), .Z(n883) );
  XNOR U992 ( .A(n882), .B(n883), .Z(n884) );
  XNOR U993 ( .A(n885), .B(n884), .Z(n900) );
  XNOR U994 ( .A(n900), .B(sreg[156]), .Z(n901) );
  XOR U995 ( .A(n902), .B(n901), .Z(c[156]) );
  NANDN U996 ( .A(n883), .B(n882), .Z(n887) );
  NAND U997 ( .A(n885), .B(n884), .Z(n886) );
  NAND U998 ( .A(n887), .B(n886), .Z(n909) );
  AND U999 ( .A(b[2]), .B(a[31]), .Z(n915) );
  AND U1000 ( .A(a[32]), .B(b[1]), .Z(n913) );
  AND U1001 ( .A(a[30]), .B(b[3]), .Z(n912) );
  XOR U1002 ( .A(n913), .B(n912), .Z(n914) );
  XOR U1003 ( .A(n915), .B(n914), .Z(n918) );
  NAND U1004 ( .A(b[0]), .B(a[33]), .Z(n919) );
  XOR U1005 ( .A(n918), .B(n919), .Z(n921) );
  OR U1006 ( .A(n889), .B(n888), .Z(n893) );
  NANDN U1007 ( .A(n891), .B(n890), .Z(n892) );
  NAND U1008 ( .A(n893), .B(n892), .Z(n920) );
  XNOR U1009 ( .A(n921), .B(n920), .Z(n906) );
  NANDN U1010 ( .A(n895), .B(n894), .Z(n899) );
  OR U1011 ( .A(n897), .B(n896), .Z(n898) );
  NAND U1012 ( .A(n899), .B(n898), .Z(n907) );
  XNOR U1013 ( .A(n906), .B(n907), .Z(n908) );
  XNOR U1014 ( .A(n909), .B(n908), .Z(n925) );
  NAND U1015 ( .A(n900), .B(sreg[156]), .Z(n904) );
  OR U1016 ( .A(n902), .B(n901), .Z(n903) );
  AND U1017 ( .A(n904), .B(n903), .Z(n924) );
  XNOR U1018 ( .A(n924), .B(sreg[157]), .Z(n905) );
  XOR U1019 ( .A(n925), .B(n905), .Z(c[157]) );
  NANDN U1020 ( .A(n907), .B(n906), .Z(n911) );
  NAND U1021 ( .A(n909), .B(n908), .Z(n910) );
  NAND U1022 ( .A(n911), .B(n910), .Z(n932) );
  AND U1023 ( .A(b[2]), .B(a[32]), .Z(n938) );
  AND U1024 ( .A(a[33]), .B(b[1]), .Z(n936) );
  AND U1025 ( .A(a[31]), .B(b[3]), .Z(n935) );
  XOR U1026 ( .A(n936), .B(n935), .Z(n937) );
  XOR U1027 ( .A(n938), .B(n937), .Z(n941) );
  NAND U1028 ( .A(b[0]), .B(a[34]), .Z(n942) );
  XOR U1029 ( .A(n941), .B(n942), .Z(n944) );
  OR U1030 ( .A(n913), .B(n912), .Z(n917) );
  NANDN U1031 ( .A(n915), .B(n914), .Z(n916) );
  NAND U1032 ( .A(n917), .B(n916), .Z(n943) );
  XNOR U1033 ( .A(n944), .B(n943), .Z(n929) );
  NANDN U1034 ( .A(n919), .B(n918), .Z(n923) );
  OR U1035 ( .A(n921), .B(n920), .Z(n922) );
  NAND U1036 ( .A(n923), .B(n922), .Z(n930) );
  XNOR U1037 ( .A(n929), .B(n930), .Z(n931) );
  XOR U1038 ( .A(n932), .B(n931), .Z(n928) );
  XOR U1039 ( .A(sreg[158]), .B(n927), .Z(n926) );
  XOR U1040 ( .A(n928), .B(n926), .Z(c[158]) );
  NANDN U1041 ( .A(n930), .B(n929), .Z(n934) );
  NAND U1042 ( .A(n932), .B(n931), .Z(n933) );
  NAND U1043 ( .A(n934), .B(n933), .Z(n950) );
  AND U1044 ( .A(b[2]), .B(a[33]), .Z(n956) );
  AND U1045 ( .A(a[34]), .B(b[1]), .Z(n954) );
  AND U1046 ( .A(a[32]), .B(b[3]), .Z(n953) );
  XOR U1047 ( .A(n954), .B(n953), .Z(n955) );
  XOR U1048 ( .A(n956), .B(n955), .Z(n959) );
  NAND U1049 ( .A(b[0]), .B(a[35]), .Z(n960) );
  XOR U1050 ( .A(n959), .B(n960), .Z(n962) );
  OR U1051 ( .A(n936), .B(n935), .Z(n940) );
  NANDN U1052 ( .A(n938), .B(n937), .Z(n939) );
  NAND U1053 ( .A(n940), .B(n939), .Z(n961) );
  XNOR U1054 ( .A(n962), .B(n961), .Z(n947) );
  NANDN U1055 ( .A(n942), .B(n941), .Z(n946) );
  OR U1056 ( .A(n944), .B(n943), .Z(n945) );
  NAND U1057 ( .A(n946), .B(n945), .Z(n948) );
  XNOR U1058 ( .A(n947), .B(n948), .Z(n949) );
  XNOR U1059 ( .A(n950), .B(n949), .Z(n965) );
  XNOR U1060 ( .A(n965), .B(sreg[159]), .Z(n966) );
  XOR U1061 ( .A(n967), .B(n966), .Z(c[159]) );
  NANDN U1062 ( .A(n948), .B(n947), .Z(n952) );
  NAND U1063 ( .A(n950), .B(n949), .Z(n951) );
  NAND U1064 ( .A(n952), .B(n951), .Z(n976) );
  AND U1065 ( .A(b[2]), .B(a[34]), .Z(n982) );
  AND U1066 ( .A(a[35]), .B(b[1]), .Z(n980) );
  AND U1067 ( .A(a[33]), .B(b[3]), .Z(n979) );
  XOR U1068 ( .A(n980), .B(n979), .Z(n981) );
  XOR U1069 ( .A(n982), .B(n981), .Z(n985) );
  NAND U1070 ( .A(b[0]), .B(a[36]), .Z(n986) );
  XOR U1071 ( .A(n985), .B(n986), .Z(n988) );
  OR U1072 ( .A(n954), .B(n953), .Z(n958) );
  NANDN U1073 ( .A(n956), .B(n955), .Z(n957) );
  NAND U1074 ( .A(n958), .B(n957), .Z(n987) );
  XNOR U1075 ( .A(n988), .B(n987), .Z(n973) );
  NANDN U1076 ( .A(n960), .B(n959), .Z(n964) );
  OR U1077 ( .A(n962), .B(n961), .Z(n963) );
  NAND U1078 ( .A(n964), .B(n963), .Z(n974) );
  XNOR U1079 ( .A(n973), .B(n974), .Z(n975) );
  XOR U1080 ( .A(n976), .B(n975), .Z(n972) );
  NAND U1081 ( .A(n965), .B(sreg[159]), .Z(n969) );
  OR U1082 ( .A(n967), .B(n966), .Z(n968) );
  NAND U1083 ( .A(n969), .B(n968), .Z(n971) );
  XNOR U1084 ( .A(sreg[160]), .B(n971), .Z(n970) );
  XOR U1085 ( .A(n972), .B(n970), .Z(c[160]) );
  NANDN U1086 ( .A(n974), .B(n973), .Z(n978) );
  NAND U1087 ( .A(n976), .B(n975), .Z(n977) );
  NAND U1088 ( .A(n978), .B(n977), .Z(n994) );
  AND U1089 ( .A(b[2]), .B(a[35]), .Z(n1000) );
  AND U1090 ( .A(a[36]), .B(b[1]), .Z(n998) );
  AND U1091 ( .A(a[34]), .B(b[3]), .Z(n997) );
  XOR U1092 ( .A(n998), .B(n997), .Z(n999) );
  XOR U1093 ( .A(n1000), .B(n999), .Z(n1003) );
  NAND U1094 ( .A(b[0]), .B(a[37]), .Z(n1004) );
  XOR U1095 ( .A(n1003), .B(n1004), .Z(n1006) );
  OR U1096 ( .A(n980), .B(n979), .Z(n984) );
  NANDN U1097 ( .A(n982), .B(n981), .Z(n983) );
  NAND U1098 ( .A(n984), .B(n983), .Z(n1005) );
  XNOR U1099 ( .A(n1006), .B(n1005), .Z(n991) );
  NANDN U1100 ( .A(n986), .B(n985), .Z(n990) );
  OR U1101 ( .A(n988), .B(n987), .Z(n989) );
  NAND U1102 ( .A(n990), .B(n989), .Z(n992) );
  XNOR U1103 ( .A(n991), .B(n992), .Z(n993) );
  XNOR U1104 ( .A(n994), .B(n993), .Z(n1009) );
  XNOR U1105 ( .A(n1009), .B(sreg[161]), .Z(n1010) );
  XOR U1106 ( .A(n1011), .B(n1010), .Z(c[161]) );
  NANDN U1107 ( .A(n992), .B(n991), .Z(n996) );
  NAND U1108 ( .A(n994), .B(n993), .Z(n995) );
  NAND U1109 ( .A(n996), .B(n995), .Z(n1020) );
  AND U1110 ( .A(b[2]), .B(a[36]), .Z(n1026) );
  AND U1111 ( .A(a[37]), .B(b[1]), .Z(n1024) );
  AND U1112 ( .A(a[35]), .B(b[3]), .Z(n1023) );
  XOR U1113 ( .A(n1024), .B(n1023), .Z(n1025) );
  XOR U1114 ( .A(n1026), .B(n1025), .Z(n1029) );
  NAND U1115 ( .A(b[0]), .B(a[38]), .Z(n1030) );
  XOR U1116 ( .A(n1029), .B(n1030), .Z(n1032) );
  OR U1117 ( .A(n998), .B(n997), .Z(n1002) );
  NANDN U1118 ( .A(n1000), .B(n999), .Z(n1001) );
  NAND U1119 ( .A(n1002), .B(n1001), .Z(n1031) );
  XNOR U1120 ( .A(n1032), .B(n1031), .Z(n1017) );
  NANDN U1121 ( .A(n1004), .B(n1003), .Z(n1008) );
  OR U1122 ( .A(n1006), .B(n1005), .Z(n1007) );
  NAND U1123 ( .A(n1008), .B(n1007), .Z(n1018) );
  XNOR U1124 ( .A(n1017), .B(n1018), .Z(n1019) );
  XOR U1125 ( .A(n1020), .B(n1019), .Z(n1016) );
  NAND U1126 ( .A(n1009), .B(sreg[161]), .Z(n1013) );
  OR U1127 ( .A(n1011), .B(n1010), .Z(n1012) );
  NAND U1128 ( .A(n1013), .B(n1012), .Z(n1015) );
  XNOR U1129 ( .A(sreg[162]), .B(n1015), .Z(n1014) );
  XOR U1130 ( .A(n1016), .B(n1014), .Z(c[162]) );
  NANDN U1131 ( .A(n1018), .B(n1017), .Z(n1022) );
  NAND U1132 ( .A(n1020), .B(n1019), .Z(n1021) );
  NAND U1133 ( .A(n1022), .B(n1021), .Z(n1038) );
  AND U1134 ( .A(b[2]), .B(a[37]), .Z(n1044) );
  AND U1135 ( .A(a[38]), .B(b[1]), .Z(n1042) );
  AND U1136 ( .A(a[36]), .B(b[3]), .Z(n1041) );
  XOR U1137 ( .A(n1042), .B(n1041), .Z(n1043) );
  XOR U1138 ( .A(n1044), .B(n1043), .Z(n1047) );
  NAND U1139 ( .A(b[0]), .B(a[39]), .Z(n1048) );
  XOR U1140 ( .A(n1047), .B(n1048), .Z(n1050) );
  OR U1141 ( .A(n1024), .B(n1023), .Z(n1028) );
  NANDN U1142 ( .A(n1026), .B(n1025), .Z(n1027) );
  NAND U1143 ( .A(n1028), .B(n1027), .Z(n1049) );
  XNOR U1144 ( .A(n1050), .B(n1049), .Z(n1035) );
  NANDN U1145 ( .A(n1030), .B(n1029), .Z(n1034) );
  OR U1146 ( .A(n1032), .B(n1031), .Z(n1033) );
  NAND U1147 ( .A(n1034), .B(n1033), .Z(n1036) );
  XNOR U1148 ( .A(n1035), .B(n1036), .Z(n1037) );
  XNOR U1149 ( .A(n1038), .B(n1037), .Z(n1053) );
  XNOR U1150 ( .A(n1053), .B(sreg[163]), .Z(n1054) );
  XOR U1151 ( .A(n1055), .B(n1054), .Z(c[163]) );
  NANDN U1152 ( .A(n1036), .B(n1035), .Z(n1040) );
  NAND U1153 ( .A(n1038), .B(n1037), .Z(n1039) );
  NAND U1154 ( .A(n1040), .B(n1039), .Z(n1061) );
  AND U1155 ( .A(b[2]), .B(a[38]), .Z(n1067) );
  AND U1156 ( .A(a[39]), .B(b[1]), .Z(n1065) );
  AND U1157 ( .A(a[37]), .B(b[3]), .Z(n1064) );
  XOR U1158 ( .A(n1065), .B(n1064), .Z(n1066) );
  XOR U1159 ( .A(n1067), .B(n1066), .Z(n1070) );
  NAND U1160 ( .A(b[0]), .B(a[40]), .Z(n1071) );
  XOR U1161 ( .A(n1070), .B(n1071), .Z(n1073) );
  OR U1162 ( .A(n1042), .B(n1041), .Z(n1046) );
  NANDN U1163 ( .A(n1044), .B(n1043), .Z(n1045) );
  NAND U1164 ( .A(n1046), .B(n1045), .Z(n1072) );
  XNOR U1165 ( .A(n1073), .B(n1072), .Z(n1058) );
  NANDN U1166 ( .A(n1048), .B(n1047), .Z(n1052) );
  OR U1167 ( .A(n1050), .B(n1049), .Z(n1051) );
  NAND U1168 ( .A(n1052), .B(n1051), .Z(n1059) );
  XNOR U1169 ( .A(n1058), .B(n1059), .Z(n1060) );
  XNOR U1170 ( .A(n1061), .B(n1060), .Z(n1076) );
  XNOR U1171 ( .A(n1076), .B(sreg[164]), .Z(n1078) );
  NAND U1172 ( .A(n1053), .B(sreg[163]), .Z(n1057) );
  OR U1173 ( .A(n1055), .B(n1054), .Z(n1056) );
  AND U1174 ( .A(n1057), .B(n1056), .Z(n1077) );
  XOR U1175 ( .A(n1078), .B(n1077), .Z(c[164]) );
  NANDN U1176 ( .A(n1059), .B(n1058), .Z(n1063) );
  NAND U1177 ( .A(n1061), .B(n1060), .Z(n1062) );
  NAND U1178 ( .A(n1063), .B(n1062), .Z(n1084) );
  AND U1179 ( .A(b[2]), .B(a[39]), .Z(n1090) );
  AND U1180 ( .A(a[40]), .B(b[1]), .Z(n1088) );
  AND U1181 ( .A(a[38]), .B(b[3]), .Z(n1087) );
  XOR U1182 ( .A(n1088), .B(n1087), .Z(n1089) );
  XOR U1183 ( .A(n1090), .B(n1089), .Z(n1093) );
  NAND U1184 ( .A(b[0]), .B(a[41]), .Z(n1094) );
  XOR U1185 ( .A(n1093), .B(n1094), .Z(n1096) );
  OR U1186 ( .A(n1065), .B(n1064), .Z(n1069) );
  NANDN U1187 ( .A(n1067), .B(n1066), .Z(n1068) );
  NAND U1188 ( .A(n1069), .B(n1068), .Z(n1095) );
  XNOR U1189 ( .A(n1096), .B(n1095), .Z(n1081) );
  NANDN U1190 ( .A(n1071), .B(n1070), .Z(n1075) );
  OR U1191 ( .A(n1073), .B(n1072), .Z(n1074) );
  NAND U1192 ( .A(n1075), .B(n1074), .Z(n1082) );
  XNOR U1193 ( .A(n1081), .B(n1082), .Z(n1083) );
  XNOR U1194 ( .A(n1084), .B(n1083), .Z(n1099) );
  XNOR U1195 ( .A(n1099), .B(sreg[165]), .Z(n1101) );
  NAND U1196 ( .A(n1076), .B(sreg[164]), .Z(n1080) );
  OR U1197 ( .A(n1078), .B(n1077), .Z(n1079) );
  AND U1198 ( .A(n1080), .B(n1079), .Z(n1100) );
  XOR U1199 ( .A(n1101), .B(n1100), .Z(c[165]) );
  NANDN U1200 ( .A(n1082), .B(n1081), .Z(n1086) );
  NAND U1201 ( .A(n1084), .B(n1083), .Z(n1085) );
  NAND U1202 ( .A(n1086), .B(n1085), .Z(n1107) );
  AND U1203 ( .A(b[2]), .B(a[40]), .Z(n1113) );
  AND U1204 ( .A(a[41]), .B(b[1]), .Z(n1111) );
  AND U1205 ( .A(a[39]), .B(b[3]), .Z(n1110) );
  XOR U1206 ( .A(n1111), .B(n1110), .Z(n1112) );
  XOR U1207 ( .A(n1113), .B(n1112), .Z(n1116) );
  NAND U1208 ( .A(b[0]), .B(a[42]), .Z(n1117) );
  XOR U1209 ( .A(n1116), .B(n1117), .Z(n1119) );
  OR U1210 ( .A(n1088), .B(n1087), .Z(n1092) );
  NANDN U1211 ( .A(n1090), .B(n1089), .Z(n1091) );
  NAND U1212 ( .A(n1092), .B(n1091), .Z(n1118) );
  XNOR U1213 ( .A(n1119), .B(n1118), .Z(n1104) );
  NANDN U1214 ( .A(n1094), .B(n1093), .Z(n1098) );
  OR U1215 ( .A(n1096), .B(n1095), .Z(n1097) );
  NAND U1216 ( .A(n1098), .B(n1097), .Z(n1105) );
  XNOR U1217 ( .A(n1104), .B(n1105), .Z(n1106) );
  XNOR U1218 ( .A(n1107), .B(n1106), .Z(n1122) );
  XNOR U1219 ( .A(n1122), .B(sreg[166]), .Z(n1124) );
  NAND U1220 ( .A(n1099), .B(sreg[165]), .Z(n1103) );
  OR U1221 ( .A(n1101), .B(n1100), .Z(n1102) );
  AND U1222 ( .A(n1103), .B(n1102), .Z(n1123) );
  XOR U1223 ( .A(n1124), .B(n1123), .Z(c[166]) );
  NANDN U1224 ( .A(n1105), .B(n1104), .Z(n1109) );
  NAND U1225 ( .A(n1107), .B(n1106), .Z(n1108) );
  NAND U1226 ( .A(n1109), .B(n1108), .Z(n1130) );
  AND U1227 ( .A(b[2]), .B(a[41]), .Z(n1136) );
  AND U1228 ( .A(a[42]), .B(b[1]), .Z(n1134) );
  AND U1229 ( .A(a[40]), .B(b[3]), .Z(n1133) );
  XOR U1230 ( .A(n1134), .B(n1133), .Z(n1135) );
  XOR U1231 ( .A(n1136), .B(n1135), .Z(n1139) );
  NAND U1232 ( .A(b[0]), .B(a[43]), .Z(n1140) );
  XOR U1233 ( .A(n1139), .B(n1140), .Z(n1142) );
  OR U1234 ( .A(n1111), .B(n1110), .Z(n1115) );
  NANDN U1235 ( .A(n1113), .B(n1112), .Z(n1114) );
  NAND U1236 ( .A(n1115), .B(n1114), .Z(n1141) );
  XNOR U1237 ( .A(n1142), .B(n1141), .Z(n1127) );
  NANDN U1238 ( .A(n1117), .B(n1116), .Z(n1121) );
  OR U1239 ( .A(n1119), .B(n1118), .Z(n1120) );
  NAND U1240 ( .A(n1121), .B(n1120), .Z(n1128) );
  XNOR U1241 ( .A(n1127), .B(n1128), .Z(n1129) );
  XNOR U1242 ( .A(n1130), .B(n1129), .Z(n1145) );
  XNOR U1243 ( .A(n1145), .B(sreg[167]), .Z(n1147) );
  NAND U1244 ( .A(n1122), .B(sreg[166]), .Z(n1126) );
  OR U1245 ( .A(n1124), .B(n1123), .Z(n1125) );
  AND U1246 ( .A(n1126), .B(n1125), .Z(n1146) );
  XOR U1247 ( .A(n1147), .B(n1146), .Z(c[167]) );
  NANDN U1248 ( .A(n1128), .B(n1127), .Z(n1132) );
  NAND U1249 ( .A(n1130), .B(n1129), .Z(n1131) );
  NAND U1250 ( .A(n1132), .B(n1131), .Z(n1153) );
  AND U1251 ( .A(b[2]), .B(a[42]), .Z(n1159) );
  AND U1252 ( .A(a[43]), .B(b[1]), .Z(n1157) );
  AND U1253 ( .A(a[41]), .B(b[3]), .Z(n1156) );
  XOR U1254 ( .A(n1157), .B(n1156), .Z(n1158) );
  XOR U1255 ( .A(n1159), .B(n1158), .Z(n1162) );
  NAND U1256 ( .A(b[0]), .B(a[44]), .Z(n1163) );
  XOR U1257 ( .A(n1162), .B(n1163), .Z(n1165) );
  OR U1258 ( .A(n1134), .B(n1133), .Z(n1138) );
  NANDN U1259 ( .A(n1136), .B(n1135), .Z(n1137) );
  NAND U1260 ( .A(n1138), .B(n1137), .Z(n1164) );
  XNOR U1261 ( .A(n1165), .B(n1164), .Z(n1150) );
  NANDN U1262 ( .A(n1140), .B(n1139), .Z(n1144) );
  OR U1263 ( .A(n1142), .B(n1141), .Z(n1143) );
  NAND U1264 ( .A(n1144), .B(n1143), .Z(n1151) );
  XNOR U1265 ( .A(n1150), .B(n1151), .Z(n1152) );
  XNOR U1266 ( .A(n1153), .B(n1152), .Z(n1168) );
  XNOR U1267 ( .A(n1168), .B(sreg[168]), .Z(n1170) );
  NAND U1268 ( .A(n1145), .B(sreg[167]), .Z(n1149) );
  OR U1269 ( .A(n1147), .B(n1146), .Z(n1148) );
  AND U1270 ( .A(n1149), .B(n1148), .Z(n1169) );
  XOR U1271 ( .A(n1170), .B(n1169), .Z(c[168]) );
  NANDN U1272 ( .A(n1151), .B(n1150), .Z(n1155) );
  NAND U1273 ( .A(n1153), .B(n1152), .Z(n1154) );
  NAND U1274 ( .A(n1155), .B(n1154), .Z(n1179) );
  AND U1275 ( .A(b[2]), .B(a[43]), .Z(n1185) );
  AND U1276 ( .A(a[44]), .B(b[1]), .Z(n1183) );
  AND U1277 ( .A(a[42]), .B(b[3]), .Z(n1182) );
  XOR U1278 ( .A(n1183), .B(n1182), .Z(n1184) );
  XOR U1279 ( .A(n1185), .B(n1184), .Z(n1188) );
  NAND U1280 ( .A(b[0]), .B(a[45]), .Z(n1189) );
  XOR U1281 ( .A(n1188), .B(n1189), .Z(n1191) );
  OR U1282 ( .A(n1157), .B(n1156), .Z(n1161) );
  NANDN U1283 ( .A(n1159), .B(n1158), .Z(n1160) );
  NAND U1284 ( .A(n1161), .B(n1160), .Z(n1190) );
  XNOR U1285 ( .A(n1191), .B(n1190), .Z(n1176) );
  NANDN U1286 ( .A(n1163), .B(n1162), .Z(n1167) );
  OR U1287 ( .A(n1165), .B(n1164), .Z(n1166) );
  NAND U1288 ( .A(n1167), .B(n1166), .Z(n1177) );
  XNOR U1289 ( .A(n1176), .B(n1177), .Z(n1178) );
  XOR U1290 ( .A(n1179), .B(n1178), .Z(n1175) );
  NAND U1291 ( .A(n1168), .B(sreg[168]), .Z(n1172) );
  OR U1292 ( .A(n1170), .B(n1169), .Z(n1171) );
  NAND U1293 ( .A(n1172), .B(n1171), .Z(n1174) );
  XNOR U1294 ( .A(sreg[169]), .B(n1174), .Z(n1173) );
  XOR U1295 ( .A(n1175), .B(n1173), .Z(c[169]) );
  NANDN U1296 ( .A(n1177), .B(n1176), .Z(n1181) );
  NAND U1297 ( .A(n1179), .B(n1178), .Z(n1180) );
  NAND U1298 ( .A(n1181), .B(n1180), .Z(n1197) );
  AND U1299 ( .A(b[2]), .B(a[44]), .Z(n1203) );
  AND U1300 ( .A(a[45]), .B(b[1]), .Z(n1201) );
  AND U1301 ( .A(a[43]), .B(b[3]), .Z(n1200) );
  XOR U1302 ( .A(n1201), .B(n1200), .Z(n1202) );
  XOR U1303 ( .A(n1203), .B(n1202), .Z(n1206) );
  NAND U1304 ( .A(b[0]), .B(a[46]), .Z(n1207) );
  XOR U1305 ( .A(n1206), .B(n1207), .Z(n1209) );
  OR U1306 ( .A(n1183), .B(n1182), .Z(n1187) );
  NANDN U1307 ( .A(n1185), .B(n1184), .Z(n1186) );
  NAND U1308 ( .A(n1187), .B(n1186), .Z(n1208) );
  XNOR U1309 ( .A(n1209), .B(n1208), .Z(n1194) );
  NANDN U1310 ( .A(n1189), .B(n1188), .Z(n1193) );
  OR U1311 ( .A(n1191), .B(n1190), .Z(n1192) );
  NAND U1312 ( .A(n1193), .B(n1192), .Z(n1195) );
  XNOR U1313 ( .A(n1194), .B(n1195), .Z(n1196) );
  XNOR U1314 ( .A(n1197), .B(n1196), .Z(n1212) );
  XNOR U1315 ( .A(n1212), .B(sreg[170]), .Z(n1213) );
  XOR U1316 ( .A(n1214), .B(n1213), .Z(c[170]) );
  NANDN U1317 ( .A(n1195), .B(n1194), .Z(n1199) );
  NAND U1318 ( .A(n1197), .B(n1196), .Z(n1198) );
  NAND U1319 ( .A(n1199), .B(n1198), .Z(n1221) );
  AND U1320 ( .A(b[2]), .B(a[45]), .Z(n1227) );
  AND U1321 ( .A(a[46]), .B(b[1]), .Z(n1225) );
  AND U1322 ( .A(a[44]), .B(b[3]), .Z(n1224) );
  XOR U1323 ( .A(n1225), .B(n1224), .Z(n1226) );
  XOR U1324 ( .A(n1227), .B(n1226), .Z(n1230) );
  NAND U1325 ( .A(b[0]), .B(a[47]), .Z(n1231) );
  XOR U1326 ( .A(n1230), .B(n1231), .Z(n1233) );
  OR U1327 ( .A(n1201), .B(n1200), .Z(n1205) );
  NANDN U1328 ( .A(n1203), .B(n1202), .Z(n1204) );
  NAND U1329 ( .A(n1205), .B(n1204), .Z(n1232) );
  XNOR U1330 ( .A(n1233), .B(n1232), .Z(n1218) );
  NANDN U1331 ( .A(n1207), .B(n1206), .Z(n1211) );
  OR U1332 ( .A(n1209), .B(n1208), .Z(n1210) );
  NAND U1333 ( .A(n1211), .B(n1210), .Z(n1219) );
  XNOR U1334 ( .A(n1218), .B(n1219), .Z(n1220) );
  XNOR U1335 ( .A(n1221), .B(n1220), .Z(n1237) );
  NAND U1336 ( .A(n1212), .B(sreg[170]), .Z(n1216) );
  OR U1337 ( .A(n1214), .B(n1213), .Z(n1215) );
  AND U1338 ( .A(n1216), .B(n1215), .Z(n1236) );
  XNOR U1339 ( .A(n1236), .B(sreg[171]), .Z(n1217) );
  XOR U1340 ( .A(n1237), .B(n1217), .Z(c[171]) );
  NANDN U1341 ( .A(n1219), .B(n1218), .Z(n1223) );
  NAND U1342 ( .A(n1221), .B(n1220), .Z(n1222) );
  NAND U1343 ( .A(n1223), .B(n1222), .Z(n1242) );
  AND U1344 ( .A(b[2]), .B(a[46]), .Z(n1248) );
  AND U1345 ( .A(a[47]), .B(b[1]), .Z(n1246) );
  AND U1346 ( .A(a[45]), .B(b[3]), .Z(n1245) );
  XOR U1347 ( .A(n1246), .B(n1245), .Z(n1247) );
  XOR U1348 ( .A(n1248), .B(n1247), .Z(n1251) );
  NAND U1349 ( .A(b[0]), .B(a[48]), .Z(n1252) );
  XOR U1350 ( .A(n1251), .B(n1252), .Z(n1254) );
  OR U1351 ( .A(n1225), .B(n1224), .Z(n1229) );
  NANDN U1352 ( .A(n1227), .B(n1226), .Z(n1228) );
  NAND U1353 ( .A(n1229), .B(n1228), .Z(n1253) );
  XNOR U1354 ( .A(n1254), .B(n1253), .Z(n1239) );
  NANDN U1355 ( .A(n1231), .B(n1230), .Z(n1235) );
  OR U1356 ( .A(n1233), .B(n1232), .Z(n1234) );
  NAND U1357 ( .A(n1235), .B(n1234), .Z(n1240) );
  XNOR U1358 ( .A(n1239), .B(n1240), .Z(n1241) );
  XOR U1359 ( .A(n1242), .B(n1241), .Z(n1258) );
  XOR U1360 ( .A(sreg[172]), .B(n1257), .Z(n1238) );
  XOR U1361 ( .A(n1258), .B(n1238), .Z(c[172]) );
  NANDN U1362 ( .A(n1240), .B(n1239), .Z(n1244) );
  NAND U1363 ( .A(n1242), .B(n1241), .Z(n1243) );
  NAND U1364 ( .A(n1244), .B(n1243), .Z(n1263) );
  AND U1365 ( .A(b[2]), .B(a[47]), .Z(n1269) );
  AND U1366 ( .A(a[48]), .B(b[1]), .Z(n1267) );
  AND U1367 ( .A(a[46]), .B(b[3]), .Z(n1266) );
  XOR U1368 ( .A(n1267), .B(n1266), .Z(n1268) );
  XOR U1369 ( .A(n1269), .B(n1268), .Z(n1272) );
  NAND U1370 ( .A(b[0]), .B(a[49]), .Z(n1273) );
  XOR U1371 ( .A(n1272), .B(n1273), .Z(n1275) );
  OR U1372 ( .A(n1246), .B(n1245), .Z(n1250) );
  NANDN U1373 ( .A(n1248), .B(n1247), .Z(n1249) );
  NAND U1374 ( .A(n1250), .B(n1249), .Z(n1274) );
  XNOR U1375 ( .A(n1275), .B(n1274), .Z(n1260) );
  NANDN U1376 ( .A(n1252), .B(n1251), .Z(n1256) );
  OR U1377 ( .A(n1254), .B(n1253), .Z(n1255) );
  NAND U1378 ( .A(n1256), .B(n1255), .Z(n1261) );
  XNOR U1379 ( .A(n1260), .B(n1261), .Z(n1262) );
  XOR U1380 ( .A(n1263), .B(n1262), .Z(n1279) );
  XNOR U1381 ( .A(sreg[173]), .B(n1278), .Z(n1259) );
  XOR U1382 ( .A(n1279), .B(n1259), .Z(c[173]) );
  NANDN U1383 ( .A(n1261), .B(n1260), .Z(n1265) );
  NAND U1384 ( .A(n1263), .B(n1262), .Z(n1264) );
  NAND U1385 ( .A(n1265), .B(n1264), .Z(n1286) );
  AND U1386 ( .A(b[2]), .B(a[48]), .Z(n1292) );
  AND U1387 ( .A(a[49]), .B(b[1]), .Z(n1290) );
  AND U1388 ( .A(a[47]), .B(b[3]), .Z(n1289) );
  XOR U1389 ( .A(n1290), .B(n1289), .Z(n1291) );
  XOR U1390 ( .A(n1292), .B(n1291), .Z(n1295) );
  NAND U1391 ( .A(b[0]), .B(a[50]), .Z(n1296) );
  XOR U1392 ( .A(n1295), .B(n1296), .Z(n1298) );
  OR U1393 ( .A(n1267), .B(n1266), .Z(n1271) );
  NANDN U1394 ( .A(n1269), .B(n1268), .Z(n1270) );
  NAND U1395 ( .A(n1271), .B(n1270), .Z(n1297) );
  XNOR U1396 ( .A(n1298), .B(n1297), .Z(n1283) );
  NANDN U1397 ( .A(n1273), .B(n1272), .Z(n1277) );
  OR U1398 ( .A(n1275), .B(n1274), .Z(n1276) );
  NAND U1399 ( .A(n1277), .B(n1276), .Z(n1284) );
  XNOR U1400 ( .A(n1283), .B(n1284), .Z(n1285) );
  XOR U1401 ( .A(n1286), .B(n1285), .Z(n1282) );
  XNOR U1402 ( .A(sreg[174]), .B(n1281), .Z(n1280) );
  XOR U1403 ( .A(n1282), .B(n1280), .Z(c[174]) );
  NANDN U1404 ( .A(n1284), .B(n1283), .Z(n1288) );
  NAND U1405 ( .A(n1286), .B(n1285), .Z(n1287) );
  NAND U1406 ( .A(n1288), .B(n1287), .Z(n1304) );
  AND U1407 ( .A(b[2]), .B(a[49]), .Z(n1310) );
  AND U1408 ( .A(a[50]), .B(b[1]), .Z(n1308) );
  AND U1409 ( .A(a[48]), .B(b[3]), .Z(n1307) );
  XOR U1410 ( .A(n1308), .B(n1307), .Z(n1309) );
  XOR U1411 ( .A(n1310), .B(n1309), .Z(n1313) );
  NAND U1412 ( .A(b[0]), .B(a[51]), .Z(n1314) );
  XOR U1413 ( .A(n1313), .B(n1314), .Z(n1316) );
  OR U1414 ( .A(n1290), .B(n1289), .Z(n1294) );
  NANDN U1415 ( .A(n1292), .B(n1291), .Z(n1293) );
  NAND U1416 ( .A(n1294), .B(n1293), .Z(n1315) );
  XNOR U1417 ( .A(n1316), .B(n1315), .Z(n1301) );
  NANDN U1418 ( .A(n1296), .B(n1295), .Z(n1300) );
  OR U1419 ( .A(n1298), .B(n1297), .Z(n1299) );
  NAND U1420 ( .A(n1300), .B(n1299), .Z(n1302) );
  XNOR U1421 ( .A(n1301), .B(n1302), .Z(n1303) );
  XNOR U1422 ( .A(n1304), .B(n1303), .Z(n1319) );
  XNOR U1423 ( .A(n1319), .B(sreg[175]), .Z(n1320) );
  XOR U1424 ( .A(n1321), .B(n1320), .Z(c[175]) );
  NANDN U1425 ( .A(n1302), .B(n1301), .Z(n1306) );
  NAND U1426 ( .A(n1304), .B(n1303), .Z(n1305) );
  NAND U1427 ( .A(n1306), .B(n1305), .Z(n1332) );
  AND U1428 ( .A(b[2]), .B(a[50]), .Z(n1338) );
  AND U1429 ( .A(a[51]), .B(b[1]), .Z(n1336) );
  AND U1430 ( .A(a[49]), .B(b[3]), .Z(n1335) );
  XOR U1431 ( .A(n1336), .B(n1335), .Z(n1337) );
  XOR U1432 ( .A(n1338), .B(n1337), .Z(n1341) );
  NAND U1433 ( .A(b[0]), .B(a[52]), .Z(n1342) );
  XOR U1434 ( .A(n1341), .B(n1342), .Z(n1344) );
  OR U1435 ( .A(n1308), .B(n1307), .Z(n1312) );
  NANDN U1436 ( .A(n1310), .B(n1309), .Z(n1311) );
  NAND U1437 ( .A(n1312), .B(n1311), .Z(n1343) );
  XNOR U1438 ( .A(n1344), .B(n1343), .Z(n1329) );
  NANDN U1439 ( .A(n1314), .B(n1313), .Z(n1318) );
  OR U1440 ( .A(n1316), .B(n1315), .Z(n1317) );
  NAND U1441 ( .A(n1318), .B(n1317), .Z(n1330) );
  XNOR U1442 ( .A(n1329), .B(n1330), .Z(n1331) );
  XNOR U1443 ( .A(n1332), .B(n1331), .Z(n1324) );
  XOR U1444 ( .A(sreg[176]), .B(n1324), .Z(n1325) );
  NAND U1445 ( .A(n1319), .B(sreg[175]), .Z(n1323) );
  OR U1446 ( .A(n1321), .B(n1320), .Z(n1322) );
  NAND U1447 ( .A(n1323), .B(n1322), .Z(n1326) );
  XOR U1448 ( .A(n1325), .B(n1326), .Z(c[176]) );
  OR U1449 ( .A(n1324), .B(sreg[176]), .Z(n1328) );
  NANDN U1450 ( .A(n1326), .B(n1325), .Z(n1327) );
  AND U1451 ( .A(n1328), .B(n1327), .Z(n1366) );
  NANDN U1452 ( .A(n1330), .B(n1329), .Z(n1334) );
  NAND U1453 ( .A(n1332), .B(n1331), .Z(n1333) );
  NAND U1454 ( .A(n1334), .B(n1333), .Z(n1351) );
  AND U1455 ( .A(b[2]), .B(a[51]), .Z(n1357) );
  AND U1456 ( .A(a[52]), .B(b[1]), .Z(n1355) );
  AND U1457 ( .A(a[50]), .B(b[3]), .Z(n1354) );
  XOR U1458 ( .A(n1355), .B(n1354), .Z(n1356) );
  XOR U1459 ( .A(n1357), .B(n1356), .Z(n1360) );
  NAND U1460 ( .A(b[0]), .B(a[53]), .Z(n1361) );
  XOR U1461 ( .A(n1360), .B(n1361), .Z(n1363) );
  OR U1462 ( .A(n1336), .B(n1335), .Z(n1340) );
  NANDN U1463 ( .A(n1338), .B(n1337), .Z(n1339) );
  NAND U1464 ( .A(n1340), .B(n1339), .Z(n1362) );
  XNOR U1465 ( .A(n1363), .B(n1362), .Z(n1348) );
  NANDN U1466 ( .A(n1342), .B(n1341), .Z(n1346) );
  OR U1467 ( .A(n1344), .B(n1343), .Z(n1345) );
  NAND U1468 ( .A(n1346), .B(n1345), .Z(n1349) );
  XNOR U1469 ( .A(n1348), .B(n1349), .Z(n1350) );
  XNOR U1470 ( .A(n1351), .B(n1350), .Z(n1367) );
  XOR U1471 ( .A(sreg[177]), .B(n1367), .Z(n1347) );
  XOR U1472 ( .A(n1366), .B(n1347), .Z(c[177]) );
  NANDN U1473 ( .A(n1349), .B(n1348), .Z(n1353) );
  NAND U1474 ( .A(n1351), .B(n1350), .Z(n1352) );
  NAND U1475 ( .A(n1353), .B(n1352), .Z(n1372) );
  AND U1476 ( .A(b[2]), .B(a[52]), .Z(n1378) );
  AND U1477 ( .A(a[53]), .B(b[1]), .Z(n1376) );
  AND U1478 ( .A(a[51]), .B(b[3]), .Z(n1375) );
  XOR U1479 ( .A(n1376), .B(n1375), .Z(n1377) );
  XOR U1480 ( .A(n1378), .B(n1377), .Z(n1381) );
  NAND U1481 ( .A(b[0]), .B(a[54]), .Z(n1382) );
  XOR U1482 ( .A(n1381), .B(n1382), .Z(n1384) );
  OR U1483 ( .A(n1355), .B(n1354), .Z(n1359) );
  NANDN U1484 ( .A(n1357), .B(n1356), .Z(n1358) );
  NAND U1485 ( .A(n1359), .B(n1358), .Z(n1383) );
  XNOR U1486 ( .A(n1384), .B(n1383), .Z(n1369) );
  NANDN U1487 ( .A(n1361), .B(n1360), .Z(n1365) );
  OR U1488 ( .A(n1363), .B(n1362), .Z(n1364) );
  NAND U1489 ( .A(n1365), .B(n1364), .Z(n1370) );
  XNOR U1490 ( .A(n1369), .B(n1370), .Z(n1371) );
  XNOR U1491 ( .A(n1372), .B(n1371), .Z(n1388) );
  XOR U1492 ( .A(n1387), .B(sreg[178]), .Z(n1368) );
  XOR U1493 ( .A(n1388), .B(n1368), .Z(c[178]) );
  NANDN U1494 ( .A(n1370), .B(n1369), .Z(n1374) );
  NAND U1495 ( .A(n1372), .B(n1371), .Z(n1373) );
  NAND U1496 ( .A(n1374), .B(n1373), .Z(n1395) );
  AND U1497 ( .A(b[2]), .B(a[53]), .Z(n1401) );
  AND U1498 ( .A(a[54]), .B(b[1]), .Z(n1399) );
  AND U1499 ( .A(a[52]), .B(b[3]), .Z(n1398) );
  XOR U1500 ( .A(n1399), .B(n1398), .Z(n1400) );
  XOR U1501 ( .A(n1401), .B(n1400), .Z(n1404) );
  NAND U1502 ( .A(b[0]), .B(a[55]), .Z(n1405) );
  XOR U1503 ( .A(n1404), .B(n1405), .Z(n1407) );
  OR U1504 ( .A(n1376), .B(n1375), .Z(n1380) );
  NANDN U1505 ( .A(n1378), .B(n1377), .Z(n1379) );
  NAND U1506 ( .A(n1380), .B(n1379), .Z(n1406) );
  XNOR U1507 ( .A(n1407), .B(n1406), .Z(n1392) );
  NANDN U1508 ( .A(n1382), .B(n1381), .Z(n1386) );
  OR U1509 ( .A(n1384), .B(n1383), .Z(n1385) );
  NAND U1510 ( .A(n1386), .B(n1385), .Z(n1393) );
  XNOR U1511 ( .A(n1392), .B(n1393), .Z(n1394) );
  XNOR U1512 ( .A(n1395), .B(n1394), .Z(n1391) );
  XOR U1513 ( .A(n1390), .B(sreg[179]), .Z(n1389) );
  XOR U1514 ( .A(n1391), .B(n1389), .Z(c[179]) );
  NANDN U1515 ( .A(n1393), .B(n1392), .Z(n1397) );
  NAND U1516 ( .A(n1395), .B(n1394), .Z(n1396) );
  NAND U1517 ( .A(n1397), .B(n1396), .Z(n1413) );
  AND U1518 ( .A(b[2]), .B(a[54]), .Z(n1419) );
  AND U1519 ( .A(a[55]), .B(b[1]), .Z(n1417) );
  AND U1520 ( .A(a[53]), .B(b[3]), .Z(n1416) );
  XOR U1521 ( .A(n1417), .B(n1416), .Z(n1418) );
  XOR U1522 ( .A(n1419), .B(n1418), .Z(n1422) );
  NAND U1523 ( .A(b[0]), .B(a[56]), .Z(n1423) );
  XOR U1524 ( .A(n1422), .B(n1423), .Z(n1425) );
  OR U1525 ( .A(n1399), .B(n1398), .Z(n1403) );
  NANDN U1526 ( .A(n1401), .B(n1400), .Z(n1402) );
  NAND U1527 ( .A(n1403), .B(n1402), .Z(n1424) );
  XNOR U1528 ( .A(n1425), .B(n1424), .Z(n1410) );
  NANDN U1529 ( .A(n1405), .B(n1404), .Z(n1409) );
  OR U1530 ( .A(n1407), .B(n1406), .Z(n1408) );
  NAND U1531 ( .A(n1409), .B(n1408), .Z(n1411) );
  XNOR U1532 ( .A(n1410), .B(n1411), .Z(n1412) );
  XNOR U1533 ( .A(n1413), .B(n1412), .Z(n1428) );
  XOR U1534 ( .A(sreg[180]), .B(n1428), .Z(n1429) );
  XOR U1535 ( .A(n1430), .B(n1429), .Z(c[180]) );
  NANDN U1536 ( .A(n1411), .B(n1410), .Z(n1415) );
  NAND U1537 ( .A(n1413), .B(n1412), .Z(n1414) );
  NAND U1538 ( .A(n1415), .B(n1414), .Z(n1439) );
  AND U1539 ( .A(b[2]), .B(a[55]), .Z(n1445) );
  AND U1540 ( .A(a[56]), .B(b[1]), .Z(n1443) );
  AND U1541 ( .A(a[54]), .B(b[3]), .Z(n1442) );
  XOR U1542 ( .A(n1443), .B(n1442), .Z(n1444) );
  XOR U1543 ( .A(n1445), .B(n1444), .Z(n1448) );
  NAND U1544 ( .A(b[0]), .B(a[57]), .Z(n1449) );
  XOR U1545 ( .A(n1448), .B(n1449), .Z(n1451) );
  OR U1546 ( .A(n1417), .B(n1416), .Z(n1421) );
  NANDN U1547 ( .A(n1419), .B(n1418), .Z(n1420) );
  NAND U1548 ( .A(n1421), .B(n1420), .Z(n1450) );
  XNOR U1549 ( .A(n1451), .B(n1450), .Z(n1436) );
  NANDN U1550 ( .A(n1423), .B(n1422), .Z(n1427) );
  OR U1551 ( .A(n1425), .B(n1424), .Z(n1426) );
  NAND U1552 ( .A(n1427), .B(n1426), .Z(n1437) );
  XNOR U1553 ( .A(n1436), .B(n1437), .Z(n1438) );
  XOR U1554 ( .A(n1439), .B(n1438), .Z(n1435) );
  OR U1555 ( .A(n1428), .B(sreg[180]), .Z(n1432) );
  NANDN U1556 ( .A(n1430), .B(n1429), .Z(n1431) );
  AND U1557 ( .A(n1432), .B(n1431), .Z(n1434) );
  XNOR U1558 ( .A(sreg[181]), .B(n1434), .Z(n1433) );
  XOR U1559 ( .A(n1435), .B(n1433), .Z(c[181]) );
  NANDN U1560 ( .A(n1437), .B(n1436), .Z(n1441) );
  NAND U1561 ( .A(n1439), .B(n1438), .Z(n1440) );
  NAND U1562 ( .A(n1441), .B(n1440), .Z(n1457) );
  AND U1563 ( .A(b[2]), .B(a[56]), .Z(n1463) );
  AND U1564 ( .A(a[57]), .B(b[1]), .Z(n1461) );
  AND U1565 ( .A(a[55]), .B(b[3]), .Z(n1460) );
  XOR U1566 ( .A(n1461), .B(n1460), .Z(n1462) );
  XOR U1567 ( .A(n1463), .B(n1462), .Z(n1466) );
  NAND U1568 ( .A(b[0]), .B(a[58]), .Z(n1467) );
  XOR U1569 ( .A(n1466), .B(n1467), .Z(n1469) );
  OR U1570 ( .A(n1443), .B(n1442), .Z(n1447) );
  NANDN U1571 ( .A(n1445), .B(n1444), .Z(n1446) );
  NAND U1572 ( .A(n1447), .B(n1446), .Z(n1468) );
  XNOR U1573 ( .A(n1469), .B(n1468), .Z(n1454) );
  NANDN U1574 ( .A(n1449), .B(n1448), .Z(n1453) );
  OR U1575 ( .A(n1451), .B(n1450), .Z(n1452) );
  NAND U1576 ( .A(n1453), .B(n1452), .Z(n1455) );
  XNOR U1577 ( .A(n1454), .B(n1455), .Z(n1456) );
  XNOR U1578 ( .A(n1457), .B(n1456), .Z(n1472) );
  XNOR U1579 ( .A(n1472), .B(sreg[182]), .Z(n1473) );
  XOR U1580 ( .A(n1474), .B(n1473), .Z(c[182]) );
  NANDN U1581 ( .A(n1455), .B(n1454), .Z(n1459) );
  NAND U1582 ( .A(n1457), .B(n1456), .Z(n1458) );
  NAND U1583 ( .A(n1459), .B(n1458), .Z(n1483) );
  AND U1584 ( .A(b[2]), .B(a[57]), .Z(n1489) );
  AND U1585 ( .A(a[58]), .B(b[1]), .Z(n1487) );
  AND U1586 ( .A(a[56]), .B(b[3]), .Z(n1486) );
  XOR U1587 ( .A(n1487), .B(n1486), .Z(n1488) );
  XOR U1588 ( .A(n1489), .B(n1488), .Z(n1492) );
  NAND U1589 ( .A(b[0]), .B(a[59]), .Z(n1493) );
  XOR U1590 ( .A(n1492), .B(n1493), .Z(n1495) );
  OR U1591 ( .A(n1461), .B(n1460), .Z(n1465) );
  NANDN U1592 ( .A(n1463), .B(n1462), .Z(n1464) );
  NAND U1593 ( .A(n1465), .B(n1464), .Z(n1494) );
  XNOR U1594 ( .A(n1495), .B(n1494), .Z(n1480) );
  NANDN U1595 ( .A(n1467), .B(n1466), .Z(n1471) );
  OR U1596 ( .A(n1469), .B(n1468), .Z(n1470) );
  NAND U1597 ( .A(n1471), .B(n1470), .Z(n1481) );
  XNOR U1598 ( .A(n1480), .B(n1481), .Z(n1482) );
  XOR U1599 ( .A(n1483), .B(n1482), .Z(n1479) );
  NAND U1600 ( .A(n1472), .B(sreg[182]), .Z(n1476) );
  OR U1601 ( .A(n1474), .B(n1473), .Z(n1475) );
  NAND U1602 ( .A(n1476), .B(n1475), .Z(n1478) );
  XNOR U1603 ( .A(sreg[183]), .B(n1478), .Z(n1477) );
  XOR U1604 ( .A(n1479), .B(n1477), .Z(c[183]) );
  NANDN U1605 ( .A(n1481), .B(n1480), .Z(n1485) );
  NAND U1606 ( .A(n1483), .B(n1482), .Z(n1484) );
  NAND U1607 ( .A(n1485), .B(n1484), .Z(n1501) );
  AND U1608 ( .A(b[2]), .B(a[58]), .Z(n1507) );
  AND U1609 ( .A(a[59]), .B(b[1]), .Z(n1505) );
  AND U1610 ( .A(a[57]), .B(b[3]), .Z(n1504) );
  XOR U1611 ( .A(n1505), .B(n1504), .Z(n1506) );
  XOR U1612 ( .A(n1507), .B(n1506), .Z(n1510) );
  NAND U1613 ( .A(b[0]), .B(a[60]), .Z(n1511) );
  XOR U1614 ( .A(n1510), .B(n1511), .Z(n1513) );
  OR U1615 ( .A(n1487), .B(n1486), .Z(n1491) );
  NANDN U1616 ( .A(n1489), .B(n1488), .Z(n1490) );
  NAND U1617 ( .A(n1491), .B(n1490), .Z(n1512) );
  XNOR U1618 ( .A(n1513), .B(n1512), .Z(n1498) );
  NANDN U1619 ( .A(n1493), .B(n1492), .Z(n1497) );
  OR U1620 ( .A(n1495), .B(n1494), .Z(n1496) );
  NAND U1621 ( .A(n1497), .B(n1496), .Z(n1499) );
  XNOR U1622 ( .A(n1498), .B(n1499), .Z(n1500) );
  XNOR U1623 ( .A(n1501), .B(n1500), .Z(n1516) );
  XNOR U1624 ( .A(n1516), .B(sreg[184]), .Z(n1517) );
  XOR U1625 ( .A(n1518), .B(n1517), .Z(c[184]) );
  NANDN U1626 ( .A(n1499), .B(n1498), .Z(n1503) );
  NAND U1627 ( .A(n1501), .B(n1500), .Z(n1502) );
  NAND U1628 ( .A(n1503), .B(n1502), .Z(n1527) );
  AND U1629 ( .A(b[2]), .B(a[59]), .Z(n1533) );
  AND U1630 ( .A(a[60]), .B(b[1]), .Z(n1531) );
  AND U1631 ( .A(a[58]), .B(b[3]), .Z(n1530) );
  XOR U1632 ( .A(n1531), .B(n1530), .Z(n1532) );
  XOR U1633 ( .A(n1533), .B(n1532), .Z(n1536) );
  NAND U1634 ( .A(b[0]), .B(a[61]), .Z(n1537) );
  XOR U1635 ( .A(n1536), .B(n1537), .Z(n1539) );
  OR U1636 ( .A(n1505), .B(n1504), .Z(n1509) );
  NANDN U1637 ( .A(n1507), .B(n1506), .Z(n1508) );
  NAND U1638 ( .A(n1509), .B(n1508), .Z(n1538) );
  XNOR U1639 ( .A(n1539), .B(n1538), .Z(n1524) );
  NANDN U1640 ( .A(n1511), .B(n1510), .Z(n1515) );
  OR U1641 ( .A(n1513), .B(n1512), .Z(n1514) );
  NAND U1642 ( .A(n1515), .B(n1514), .Z(n1525) );
  XNOR U1643 ( .A(n1524), .B(n1525), .Z(n1526) );
  XNOR U1644 ( .A(n1527), .B(n1526), .Z(n1523) );
  NAND U1645 ( .A(n1516), .B(sreg[184]), .Z(n1520) );
  OR U1646 ( .A(n1518), .B(n1517), .Z(n1519) );
  AND U1647 ( .A(n1520), .B(n1519), .Z(n1522) );
  XNOR U1648 ( .A(n1522), .B(sreg[185]), .Z(n1521) );
  XOR U1649 ( .A(n1523), .B(n1521), .Z(c[185]) );
  NANDN U1650 ( .A(n1525), .B(n1524), .Z(n1529) );
  NAND U1651 ( .A(n1527), .B(n1526), .Z(n1528) );
  NAND U1652 ( .A(n1529), .B(n1528), .Z(n1545) );
  AND U1653 ( .A(b[2]), .B(a[60]), .Z(n1551) );
  AND U1654 ( .A(a[61]), .B(b[1]), .Z(n1549) );
  AND U1655 ( .A(a[59]), .B(b[3]), .Z(n1548) );
  XOR U1656 ( .A(n1549), .B(n1548), .Z(n1550) );
  XOR U1657 ( .A(n1551), .B(n1550), .Z(n1554) );
  NAND U1658 ( .A(b[0]), .B(a[62]), .Z(n1555) );
  XOR U1659 ( .A(n1554), .B(n1555), .Z(n1557) );
  OR U1660 ( .A(n1531), .B(n1530), .Z(n1535) );
  NANDN U1661 ( .A(n1533), .B(n1532), .Z(n1534) );
  NAND U1662 ( .A(n1535), .B(n1534), .Z(n1556) );
  XNOR U1663 ( .A(n1557), .B(n1556), .Z(n1542) );
  NANDN U1664 ( .A(n1537), .B(n1536), .Z(n1541) );
  OR U1665 ( .A(n1539), .B(n1538), .Z(n1540) );
  NAND U1666 ( .A(n1541), .B(n1540), .Z(n1543) );
  XNOR U1667 ( .A(n1542), .B(n1543), .Z(n1544) );
  XNOR U1668 ( .A(n1545), .B(n1544), .Z(n1560) );
  XNOR U1669 ( .A(n1560), .B(sreg[186]), .Z(n1562) );
  XNOR U1670 ( .A(n1561), .B(n1562), .Z(c[186]) );
  NANDN U1671 ( .A(n1543), .B(n1542), .Z(n1547) );
  NAND U1672 ( .A(n1545), .B(n1544), .Z(n1546) );
  NAND U1673 ( .A(n1547), .B(n1546), .Z(n1573) );
  AND U1674 ( .A(b[2]), .B(a[61]), .Z(n1579) );
  AND U1675 ( .A(a[62]), .B(b[1]), .Z(n1577) );
  AND U1676 ( .A(a[60]), .B(b[3]), .Z(n1576) );
  XOR U1677 ( .A(n1577), .B(n1576), .Z(n1578) );
  XOR U1678 ( .A(n1579), .B(n1578), .Z(n1582) );
  NAND U1679 ( .A(b[0]), .B(a[63]), .Z(n1583) );
  XOR U1680 ( .A(n1582), .B(n1583), .Z(n1585) );
  OR U1681 ( .A(n1549), .B(n1548), .Z(n1553) );
  NANDN U1682 ( .A(n1551), .B(n1550), .Z(n1552) );
  NAND U1683 ( .A(n1553), .B(n1552), .Z(n1584) );
  XNOR U1684 ( .A(n1585), .B(n1584), .Z(n1570) );
  NANDN U1685 ( .A(n1555), .B(n1554), .Z(n1559) );
  OR U1686 ( .A(n1557), .B(n1556), .Z(n1558) );
  NAND U1687 ( .A(n1559), .B(n1558), .Z(n1571) );
  XNOR U1688 ( .A(n1570), .B(n1571), .Z(n1572) );
  XNOR U1689 ( .A(n1573), .B(n1572), .Z(n1565) );
  XNOR U1690 ( .A(n1565), .B(sreg[187]), .Z(n1567) );
  NAND U1691 ( .A(n1560), .B(sreg[186]), .Z(n1564) );
  NANDN U1692 ( .A(n1562), .B(n1561), .Z(n1563) );
  AND U1693 ( .A(n1564), .B(n1563), .Z(n1566) );
  XOR U1694 ( .A(n1567), .B(n1566), .Z(c[187]) );
  NAND U1695 ( .A(n1565), .B(sreg[187]), .Z(n1569) );
  OR U1696 ( .A(n1567), .B(n1566), .Z(n1568) );
  AND U1697 ( .A(n1569), .B(n1568), .Z(n1609) );
  NANDN U1698 ( .A(n1571), .B(n1570), .Z(n1575) );
  NAND U1699 ( .A(n1573), .B(n1572), .Z(n1574) );
  NAND U1700 ( .A(n1575), .B(n1574), .Z(n1592) );
  AND U1701 ( .A(b[2]), .B(a[62]), .Z(n1604) );
  AND U1702 ( .A(a[63]), .B(b[1]), .Z(n1602) );
  AND U1703 ( .A(a[61]), .B(b[3]), .Z(n1601) );
  XOR U1704 ( .A(n1602), .B(n1601), .Z(n1603) );
  XOR U1705 ( .A(n1604), .B(n1603), .Z(n1595) );
  NAND U1706 ( .A(b[0]), .B(a[64]), .Z(n1596) );
  XOR U1707 ( .A(n1595), .B(n1596), .Z(n1598) );
  OR U1708 ( .A(n1577), .B(n1576), .Z(n1581) );
  NANDN U1709 ( .A(n1579), .B(n1578), .Z(n1580) );
  NAND U1710 ( .A(n1581), .B(n1580), .Z(n1597) );
  XNOR U1711 ( .A(n1598), .B(n1597), .Z(n1589) );
  NANDN U1712 ( .A(n1583), .B(n1582), .Z(n1587) );
  OR U1713 ( .A(n1585), .B(n1584), .Z(n1586) );
  NAND U1714 ( .A(n1587), .B(n1586), .Z(n1590) );
  XNOR U1715 ( .A(n1589), .B(n1590), .Z(n1591) );
  XNOR U1716 ( .A(n1592), .B(n1591), .Z(n1608) );
  XNOR U1717 ( .A(sreg[188]), .B(n1608), .Z(n1588) );
  XOR U1718 ( .A(n1609), .B(n1588), .Z(c[188]) );
  NANDN U1719 ( .A(n1590), .B(n1589), .Z(n1594) );
  NAND U1720 ( .A(n1592), .B(n1591), .Z(n1593) );
  NAND U1721 ( .A(n1594), .B(n1593), .Z(n1613) );
  NANDN U1722 ( .A(n1596), .B(n1595), .Z(n1600) );
  OR U1723 ( .A(n1598), .B(n1597), .Z(n1599) );
  AND U1724 ( .A(n1600), .B(n1599), .Z(n1612) );
  AND U1725 ( .A(b[2]), .B(a[63]), .Z(n1617) );
  AND U1726 ( .A(a[64]), .B(b[1]), .Z(n1615) );
  AND U1727 ( .A(a[62]), .B(b[3]), .Z(n1614) );
  XOR U1728 ( .A(n1615), .B(n1614), .Z(n1616) );
  XOR U1729 ( .A(n1617), .B(n1616), .Z(n1620) );
  NAND U1730 ( .A(b[0]), .B(a[65]), .Z(n1621) );
  XOR U1731 ( .A(n1620), .B(n1621), .Z(n1623) );
  OR U1732 ( .A(n1602), .B(n1601), .Z(n1606) );
  NANDN U1733 ( .A(n1604), .B(n1603), .Z(n1605) );
  NAND U1734 ( .A(n1606), .B(n1605), .Z(n1622) );
  XOR U1735 ( .A(n1623), .B(n1622), .Z(n1611) );
  XNOR U1736 ( .A(n1612), .B(n1611), .Z(n1607) );
  XNOR U1737 ( .A(n1613), .B(n1607), .Z(n1627) );
  XOR U1738 ( .A(n1626), .B(sreg[189]), .Z(n1610) );
  XOR U1739 ( .A(n1627), .B(n1610), .Z(c[189]) );
  AND U1740 ( .A(b[2]), .B(a[64]), .Z(n1640) );
  AND U1741 ( .A(a[65]), .B(b[1]), .Z(n1638) );
  AND U1742 ( .A(a[63]), .B(b[3]), .Z(n1637) );
  XOR U1743 ( .A(n1638), .B(n1637), .Z(n1639) );
  XOR U1744 ( .A(n1640), .B(n1639), .Z(n1643) );
  NAND U1745 ( .A(b[0]), .B(a[66]), .Z(n1644) );
  XOR U1746 ( .A(n1643), .B(n1644), .Z(n1646) );
  OR U1747 ( .A(n1615), .B(n1614), .Z(n1619) );
  NANDN U1748 ( .A(n1617), .B(n1616), .Z(n1618) );
  NAND U1749 ( .A(n1619), .B(n1618), .Z(n1645) );
  XNOR U1750 ( .A(n1646), .B(n1645), .Z(n1631) );
  NANDN U1751 ( .A(n1621), .B(n1620), .Z(n1625) );
  OR U1752 ( .A(n1623), .B(n1622), .Z(n1624) );
  NAND U1753 ( .A(n1625), .B(n1624), .Z(n1632) );
  XNOR U1754 ( .A(n1631), .B(n1632), .Z(n1633) );
  XOR U1755 ( .A(n1634), .B(n1633), .Z(n1630) );
  XOR U1756 ( .A(sreg[190]), .B(n1629), .Z(n1628) );
  XNOR U1757 ( .A(n1630), .B(n1628), .Z(c[190]) );
  NANDN U1758 ( .A(n1632), .B(n1631), .Z(n1636) );
  NANDN U1759 ( .A(n1634), .B(n1633), .Z(n1635) );
  NAND U1760 ( .A(n1636), .B(n1635), .Z(n1652) );
  AND U1761 ( .A(b[2]), .B(a[65]), .Z(n1658) );
  AND U1762 ( .A(a[66]), .B(b[1]), .Z(n1656) );
  AND U1763 ( .A(a[64]), .B(b[3]), .Z(n1655) );
  XOR U1764 ( .A(n1656), .B(n1655), .Z(n1657) );
  XOR U1765 ( .A(n1658), .B(n1657), .Z(n1661) );
  NAND U1766 ( .A(b[0]), .B(a[67]), .Z(n1662) );
  XOR U1767 ( .A(n1661), .B(n1662), .Z(n1664) );
  OR U1768 ( .A(n1638), .B(n1637), .Z(n1642) );
  NANDN U1769 ( .A(n1640), .B(n1639), .Z(n1641) );
  NAND U1770 ( .A(n1642), .B(n1641), .Z(n1663) );
  XNOR U1771 ( .A(n1664), .B(n1663), .Z(n1649) );
  NANDN U1772 ( .A(n1644), .B(n1643), .Z(n1648) );
  OR U1773 ( .A(n1646), .B(n1645), .Z(n1647) );
  NAND U1774 ( .A(n1648), .B(n1647), .Z(n1650) );
  XNOR U1775 ( .A(n1649), .B(n1650), .Z(n1651) );
  XNOR U1776 ( .A(n1652), .B(n1651), .Z(n1668) );
  XNOR U1777 ( .A(n1668), .B(sreg[191]), .Z(n1669) );
  XOR U1778 ( .A(n1670), .B(n1669), .Z(c[191]) );
  NANDN U1779 ( .A(n1650), .B(n1649), .Z(n1654) );
  NAND U1780 ( .A(n1652), .B(n1651), .Z(n1653) );
  AND U1781 ( .A(n1654), .B(n1653), .Z(n1675) );
  AND U1782 ( .A(b[2]), .B(a[66]), .Z(n1679) );
  AND U1783 ( .A(a[67]), .B(b[1]), .Z(n1677) );
  AND U1784 ( .A(a[65]), .B(b[3]), .Z(n1676) );
  XOR U1785 ( .A(n1677), .B(n1676), .Z(n1678) );
  XOR U1786 ( .A(n1679), .B(n1678), .Z(n1682) );
  NAND U1787 ( .A(b[0]), .B(a[68]), .Z(n1683) );
  XOR U1788 ( .A(n1682), .B(n1683), .Z(n1684) );
  OR U1789 ( .A(n1656), .B(n1655), .Z(n1660) );
  NANDN U1790 ( .A(n1658), .B(n1657), .Z(n1659) );
  AND U1791 ( .A(n1660), .B(n1659), .Z(n1685) );
  XOR U1792 ( .A(n1684), .B(n1685), .Z(n1673) );
  NANDN U1793 ( .A(n1662), .B(n1661), .Z(n1666) );
  OR U1794 ( .A(n1664), .B(n1663), .Z(n1665) );
  AND U1795 ( .A(n1666), .B(n1665), .Z(n1674) );
  XOR U1796 ( .A(n1673), .B(n1674), .Z(n1667) );
  XOR U1797 ( .A(n1675), .B(n1667), .Z(n1686) );
  XNOR U1798 ( .A(sreg[192]), .B(n1686), .Z(n1688) );
  NAND U1799 ( .A(n1668), .B(sreg[191]), .Z(n1672) );
  OR U1800 ( .A(n1670), .B(n1669), .Z(n1671) );
  AND U1801 ( .A(n1672), .B(n1671), .Z(n1687) );
  XOR U1802 ( .A(n1688), .B(n1687), .Z(c[192]) );
  AND U1803 ( .A(b[2]), .B(a[67]), .Z(n1700) );
  AND U1804 ( .A(a[68]), .B(b[1]), .Z(n1698) );
  AND U1805 ( .A(a[66]), .B(b[3]), .Z(n1697) );
  XOR U1806 ( .A(n1698), .B(n1697), .Z(n1699) );
  XOR U1807 ( .A(n1700), .B(n1699), .Z(n1703) );
  NAND U1808 ( .A(b[0]), .B(a[69]), .Z(n1704) );
  XOR U1809 ( .A(n1703), .B(n1704), .Z(n1706) );
  OR U1810 ( .A(n1677), .B(n1676), .Z(n1681) );
  NANDN U1811 ( .A(n1679), .B(n1678), .Z(n1680) );
  NAND U1812 ( .A(n1681), .B(n1680), .Z(n1705) );
  XNOR U1813 ( .A(n1706), .B(n1705), .Z(n1691) );
  XNOR U1814 ( .A(n1691), .B(n1692), .Z(n1694) );
  XOR U1815 ( .A(n1693), .B(n1694), .Z(n1709) );
  XOR U1816 ( .A(n1709), .B(sreg[193]), .Z(n1711) );
  NAND U1817 ( .A(sreg[192]), .B(n1686), .Z(n1690) );
  OR U1818 ( .A(n1688), .B(n1687), .Z(n1689) );
  AND U1819 ( .A(n1690), .B(n1689), .Z(n1710) );
  XOR U1820 ( .A(n1711), .B(n1710), .Z(c[193]) );
  NANDN U1821 ( .A(n1692), .B(n1691), .Z(n1696) );
  NAND U1822 ( .A(n1694), .B(n1693), .Z(n1695) );
  NAND U1823 ( .A(n1696), .B(n1695), .Z(n1720) );
  AND U1824 ( .A(b[2]), .B(a[68]), .Z(n1726) );
  AND U1825 ( .A(a[69]), .B(b[1]), .Z(n1724) );
  AND U1826 ( .A(a[67]), .B(b[3]), .Z(n1723) );
  XOR U1827 ( .A(n1724), .B(n1723), .Z(n1725) );
  XOR U1828 ( .A(n1726), .B(n1725), .Z(n1729) );
  NAND U1829 ( .A(b[0]), .B(a[70]), .Z(n1730) );
  XOR U1830 ( .A(n1729), .B(n1730), .Z(n1732) );
  OR U1831 ( .A(n1698), .B(n1697), .Z(n1702) );
  NANDN U1832 ( .A(n1700), .B(n1699), .Z(n1701) );
  NAND U1833 ( .A(n1702), .B(n1701), .Z(n1731) );
  XNOR U1834 ( .A(n1732), .B(n1731), .Z(n1717) );
  NANDN U1835 ( .A(n1704), .B(n1703), .Z(n1708) );
  OR U1836 ( .A(n1706), .B(n1705), .Z(n1707) );
  NAND U1837 ( .A(n1708), .B(n1707), .Z(n1718) );
  XNOR U1838 ( .A(n1717), .B(n1718), .Z(n1719) );
  XNOR U1839 ( .A(n1720), .B(n1719), .Z(n1716) );
  NANDN U1840 ( .A(n1709), .B(sreg[193]), .Z(n1713) );
  OR U1841 ( .A(n1711), .B(n1710), .Z(n1712) );
  AND U1842 ( .A(n1713), .B(n1712), .Z(n1715) );
  XNOR U1843 ( .A(n1715), .B(sreg[194]), .Z(n1714) );
  XOR U1844 ( .A(n1716), .B(n1714), .Z(c[194]) );
  NANDN U1845 ( .A(n1718), .B(n1717), .Z(n1722) );
  NAND U1846 ( .A(n1720), .B(n1719), .Z(n1721) );
  NAND U1847 ( .A(n1722), .B(n1721), .Z(n1738) );
  AND U1848 ( .A(b[2]), .B(a[69]), .Z(n1744) );
  AND U1849 ( .A(a[70]), .B(b[1]), .Z(n1742) );
  AND U1850 ( .A(a[68]), .B(b[3]), .Z(n1741) );
  XOR U1851 ( .A(n1742), .B(n1741), .Z(n1743) );
  XOR U1852 ( .A(n1744), .B(n1743), .Z(n1747) );
  NAND U1853 ( .A(b[0]), .B(a[71]), .Z(n1748) );
  XOR U1854 ( .A(n1747), .B(n1748), .Z(n1750) );
  OR U1855 ( .A(n1724), .B(n1723), .Z(n1728) );
  NANDN U1856 ( .A(n1726), .B(n1725), .Z(n1727) );
  NAND U1857 ( .A(n1728), .B(n1727), .Z(n1749) );
  XNOR U1858 ( .A(n1750), .B(n1749), .Z(n1735) );
  NANDN U1859 ( .A(n1730), .B(n1729), .Z(n1734) );
  OR U1860 ( .A(n1732), .B(n1731), .Z(n1733) );
  NAND U1861 ( .A(n1734), .B(n1733), .Z(n1736) );
  XNOR U1862 ( .A(n1735), .B(n1736), .Z(n1737) );
  XNOR U1863 ( .A(n1738), .B(n1737), .Z(n1753) );
  XNOR U1864 ( .A(n1753), .B(sreg[195]), .Z(n1755) );
  XNOR U1865 ( .A(n1754), .B(n1755), .Z(c[195]) );
  NANDN U1866 ( .A(n1736), .B(n1735), .Z(n1740) );
  NAND U1867 ( .A(n1738), .B(n1737), .Z(n1739) );
  NAND U1868 ( .A(n1740), .B(n1739), .Z(n1764) );
  AND U1869 ( .A(b[2]), .B(a[70]), .Z(n1770) );
  AND U1870 ( .A(a[71]), .B(b[1]), .Z(n1768) );
  AND U1871 ( .A(a[69]), .B(b[3]), .Z(n1767) );
  XOR U1872 ( .A(n1768), .B(n1767), .Z(n1769) );
  XOR U1873 ( .A(n1770), .B(n1769), .Z(n1773) );
  NAND U1874 ( .A(b[0]), .B(a[72]), .Z(n1774) );
  XOR U1875 ( .A(n1773), .B(n1774), .Z(n1776) );
  OR U1876 ( .A(n1742), .B(n1741), .Z(n1746) );
  NANDN U1877 ( .A(n1744), .B(n1743), .Z(n1745) );
  NAND U1878 ( .A(n1746), .B(n1745), .Z(n1775) );
  XNOR U1879 ( .A(n1776), .B(n1775), .Z(n1761) );
  NANDN U1880 ( .A(n1748), .B(n1747), .Z(n1752) );
  OR U1881 ( .A(n1750), .B(n1749), .Z(n1751) );
  NAND U1882 ( .A(n1752), .B(n1751), .Z(n1762) );
  XNOR U1883 ( .A(n1761), .B(n1762), .Z(n1763) );
  XOR U1884 ( .A(n1764), .B(n1763), .Z(n1760) );
  NAND U1885 ( .A(n1753), .B(sreg[195]), .Z(n1757) );
  NANDN U1886 ( .A(n1755), .B(n1754), .Z(n1756) );
  NAND U1887 ( .A(n1757), .B(n1756), .Z(n1759) );
  XNOR U1888 ( .A(sreg[196]), .B(n1759), .Z(n1758) );
  XOR U1889 ( .A(n1760), .B(n1758), .Z(c[196]) );
  NANDN U1890 ( .A(n1762), .B(n1761), .Z(n1766) );
  NAND U1891 ( .A(n1764), .B(n1763), .Z(n1765) );
  NAND U1892 ( .A(n1766), .B(n1765), .Z(n1782) );
  AND U1893 ( .A(b[2]), .B(a[71]), .Z(n1788) );
  AND U1894 ( .A(a[72]), .B(b[1]), .Z(n1786) );
  AND U1895 ( .A(a[70]), .B(b[3]), .Z(n1785) );
  XOR U1896 ( .A(n1786), .B(n1785), .Z(n1787) );
  XOR U1897 ( .A(n1788), .B(n1787), .Z(n1791) );
  NAND U1898 ( .A(b[0]), .B(a[73]), .Z(n1792) );
  XOR U1899 ( .A(n1791), .B(n1792), .Z(n1794) );
  OR U1900 ( .A(n1768), .B(n1767), .Z(n1772) );
  NANDN U1901 ( .A(n1770), .B(n1769), .Z(n1771) );
  NAND U1902 ( .A(n1772), .B(n1771), .Z(n1793) );
  XNOR U1903 ( .A(n1794), .B(n1793), .Z(n1779) );
  NANDN U1904 ( .A(n1774), .B(n1773), .Z(n1778) );
  OR U1905 ( .A(n1776), .B(n1775), .Z(n1777) );
  NAND U1906 ( .A(n1778), .B(n1777), .Z(n1780) );
  XNOR U1907 ( .A(n1779), .B(n1780), .Z(n1781) );
  XNOR U1908 ( .A(n1782), .B(n1781), .Z(n1797) );
  XNOR U1909 ( .A(n1797), .B(sreg[197]), .Z(n1798) );
  XOR U1910 ( .A(n1799), .B(n1798), .Z(c[197]) );
  NANDN U1911 ( .A(n1780), .B(n1779), .Z(n1784) );
  NAND U1912 ( .A(n1782), .B(n1781), .Z(n1783) );
  NAND U1913 ( .A(n1784), .B(n1783), .Z(n1805) );
  AND U1914 ( .A(b[2]), .B(a[72]), .Z(n1811) );
  AND U1915 ( .A(a[73]), .B(b[1]), .Z(n1809) );
  AND U1916 ( .A(a[71]), .B(b[3]), .Z(n1808) );
  XOR U1917 ( .A(n1809), .B(n1808), .Z(n1810) );
  XOR U1918 ( .A(n1811), .B(n1810), .Z(n1814) );
  NAND U1919 ( .A(b[0]), .B(a[74]), .Z(n1815) );
  XOR U1920 ( .A(n1814), .B(n1815), .Z(n1817) );
  OR U1921 ( .A(n1786), .B(n1785), .Z(n1790) );
  NANDN U1922 ( .A(n1788), .B(n1787), .Z(n1789) );
  NAND U1923 ( .A(n1790), .B(n1789), .Z(n1816) );
  XNOR U1924 ( .A(n1817), .B(n1816), .Z(n1802) );
  NANDN U1925 ( .A(n1792), .B(n1791), .Z(n1796) );
  OR U1926 ( .A(n1794), .B(n1793), .Z(n1795) );
  NAND U1927 ( .A(n1796), .B(n1795), .Z(n1803) );
  XNOR U1928 ( .A(n1802), .B(n1803), .Z(n1804) );
  XNOR U1929 ( .A(n1805), .B(n1804), .Z(n1820) );
  XOR U1930 ( .A(sreg[198]), .B(n1820), .Z(n1821) );
  NAND U1931 ( .A(n1797), .B(sreg[197]), .Z(n1801) );
  OR U1932 ( .A(n1799), .B(n1798), .Z(n1800) );
  NAND U1933 ( .A(n1801), .B(n1800), .Z(n1822) );
  XOR U1934 ( .A(n1821), .B(n1822), .Z(c[198]) );
  NANDN U1935 ( .A(n1803), .B(n1802), .Z(n1807) );
  NAND U1936 ( .A(n1805), .B(n1804), .Z(n1806) );
  NAND U1937 ( .A(n1807), .B(n1806), .Z(n1829) );
  AND U1938 ( .A(b[2]), .B(a[73]), .Z(n1835) );
  AND U1939 ( .A(a[74]), .B(b[1]), .Z(n1833) );
  AND U1940 ( .A(a[72]), .B(b[3]), .Z(n1832) );
  XOR U1941 ( .A(n1833), .B(n1832), .Z(n1834) );
  XOR U1942 ( .A(n1835), .B(n1834), .Z(n1838) );
  NAND U1943 ( .A(b[0]), .B(a[75]), .Z(n1839) );
  XOR U1944 ( .A(n1838), .B(n1839), .Z(n1841) );
  OR U1945 ( .A(n1809), .B(n1808), .Z(n1813) );
  NANDN U1946 ( .A(n1811), .B(n1810), .Z(n1812) );
  NAND U1947 ( .A(n1813), .B(n1812), .Z(n1840) );
  XNOR U1948 ( .A(n1841), .B(n1840), .Z(n1826) );
  NANDN U1949 ( .A(n1815), .B(n1814), .Z(n1819) );
  OR U1950 ( .A(n1817), .B(n1816), .Z(n1818) );
  NAND U1951 ( .A(n1819), .B(n1818), .Z(n1827) );
  XNOR U1952 ( .A(n1826), .B(n1827), .Z(n1828) );
  XOR U1953 ( .A(n1829), .B(n1828), .Z(n1845) );
  OR U1954 ( .A(n1820), .B(sreg[198]), .Z(n1824) );
  NANDN U1955 ( .A(n1822), .B(n1821), .Z(n1823) );
  AND U1956 ( .A(n1824), .B(n1823), .Z(n1844) );
  XNOR U1957 ( .A(sreg[199]), .B(n1844), .Z(n1825) );
  XOR U1958 ( .A(n1845), .B(n1825), .Z(c[199]) );
  NANDN U1959 ( .A(n1827), .B(n1826), .Z(n1831) );
  NAND U1960 ( .A(n1829), .B(n1828), .Z(n1830) );
  NAND U1961 ( .A(n1831), .B(n1830), .Z(n1852) );
  AND U1962 ( .A(b[2]), .B(a[74]), .Z(n1858) );
  AND U1963 ( .A(a[75]), .B(b[1]), .Z(n1856) );
  AND U1964 ( .A(a[73]), .B(b[3]), .Z(n1855) );
  XOR U1965 ( .A(n1856), .B(n1855), .Z(n1857) );
  XOR U1966 ( .A(n1858), .B(n1857), .Z(n1861) );
  NAND U1967 ( .A(b[0]), .B(a[76]), .Z(n1862) );
  XOR U1968 ( .A(n1861), .B(n1862), .Z(n1864) );
  OR U1969 ( .A(n1833), .B(n1832), .Z(n1837) );
  NANDN U1970 ( .A(n1835), .B(n1834), .Z(n1836) );
  NAND U1971 ( .A(n1837), .B(n1836), .Z(n1863) );
  XNOR U1972 ( .A(n1864), .B(n1863), .Z(n1849) );
  NANDN U1973 ( .A(n1839), .B(n1838), .Z(n1843) );
  OR U1974 ( .A(n1841), .B(n1840), .Z(n1842) );
  NAND U1975 ( .A(n1843), .B(n1842), .Z(n1850) );
  XNOR U1976 ( .A(n1849), .B(n1850), .Z(n1851) );
  XOR U1977 ( .A(n1852), .B(n1851), .Z(n1848) );
  XNOR U1978 ( .A(sreg[200]), .B(n1847), .Z(n1846) );
  XOR U1979 ( .A(n1848), .B(n1846), .Z(c[200]) );
  NANDN U1980 ( .A(n1850), .B(n1849), .Z(n1854) );
  NAND U1981 ( .A(n1852), .B(n1851), .Z(n1853) );
  NAND U1982 ( .A(n1854), .B(n1853), .Z(n1870) );
  AND U1983 ( .A(b[2]), .B(a[75]), .Z(n1876) );
  AND U1984 ( .A(a[76]), .B(b[1]), .Z(n1874) );
  AND U1985 ( .A(a[74]), .B(b[3]), .Z(n1873) );
  XOR U1986 ( .A(n1874), .B(n1873), .Z(n1875) );
  XOR U1987 ( .A(n1876), .B(n1875), .Z(n1879) );
  NAND U1988 ( .A(b[0]), .B(a[77]), .Z(n1880) );
  XOR U1989 ( .A(n1879), .B(n1880), .Z(n1882) );
  OR U1990 ( .A(n1856), .B(n1855), .Z(n1860) );
  NANDN U1991 ( .A(n1858), .B(n1857), .Z(n1859) );
  NAND U1992 ( .A(n1860), .B(n1859), .Z(n1881) );
  XNOR U1993 ( .A(n1882), .B(n1881), .Z(n1867) );
  NANDN U1994 ( .A(n1862), .B(n1861), .Z(n1866) );
  OR U1995 ( .A(n1864), .B(n1863), .Z(n1865) );
  NAND U1996 ( .A(n1866), .B(n1865), .Z(n1868) );
  XNOR U1997 ( .A(n1867), .B(n1868), .Z(n1869) );
  XNOR U1998 ( .A(n1870), .B(n1869), .Z(n1885) );
  XNOR U1999 ( .A(n1885), .B(sreg[201]), .Z(n1886) );
  XOR U2000 ( .A(n1887), .B(n1886), .Z(c[201]) );
  NANDN U2001 ( .A(n1868), .B(n1867), .Z(n1872) );
  NAND U2002 ( .A(n1870), .B(n1869), .Z(n1871) );
  NAND U2003 ( .A(n1872), .B(n1871), .Z(n1893) );
  AND U2004 ( .A(b[2]), .B(a[76]), .Z(n1899) );
  AND U2005 ( .A(a[77]), .B(b[1]), .Z(n1897) );
  AND U2006 ( .A(a[75]), .B(b[3]), .Z(n1896) );
  XOR U2007 ( .A(n1897), .B(n1896), .Z(n1898) );
  XOR U2008 ( .A(n1899), .B(n1898), .Z(n1902) );
  NAND U2009 ( .A(b[0]), .B(a[78]), .Z(n1903) );
  XOR U2010 ( .A(n1902), .B(n1903), .Z(n1905) );
  OR U2011 ( .A(n1874), .B(n1873), .Z(n1878) );
  NANDN U2012 ( .A(n1876), .B(n1875), .Z(n1877) );
  NAND U2013 ( .A(n1878), .B(n1877), .Z(n1904) );
  XNOR U2014 ( .A(n1905), .B(n1904), .Z(n1890) );
  NANDN U2015 ( .A(n1880), .B(n1879), .Z(n1884) );
  OR U2016 ( .A(n1882), .B(n1881), .Z(n1883) );
  NAND U2017 ( .A(n1884), .B(n1883), .Z(n1891) );
  XNOR U2018 ( .A(n1890), .B(n1891), .Z(n1892) );
  XNOR U2019 ( .A(n1893), .B(n1892), .Z(n1908) );
  XNOR U2020 ( .A(n1908), .B(sreg[202]), .Z(n1910) );
  NAND U2021 ( .A(n1885), .B(sreg[201]), .Z(n1889) );
  OR U2022 ( .A(n1887), .B(n1886), .Z(n1888) );
  AND U2023 ( .A(n1889), .B(n1888), .Z(n1909) );
  XOR U2024 ( .A(n1910), .B(n1909), .Z(c[202]) );
  NANDN U2025 ( .A(n1891), .B(n1890), .Z(n1895) );
  NAND U2026 ( .A(n1893), .B(n1892), .Z(n1894) );
  NAND U2027 ( .A(n1895), .B(n1894), .Z(n1919) );
  AND U2028 ( .A(b[2]), .B(a[77]), .Z(n1925) );
  AND U2029 ( .A(a[78]), .B(b[1]), .Z(n1923) );
  AND U2030 ( .A(a[76]), .B(b[3]), .Z(n1922) );
  XOR U2031 ( .A(n1923), .B(n1922), .Z(n1924) );
  XOR U2032 ( .A(n1925), .B(n1924), .Z(n1928) );
  NAND U2033 ( .A(b[0]), .B(a[79]), .Z(n1929) );
  XOR U2034 ( .A(n1928), .B(n1929), .Z(n1931) );
  OR U2035 ( .A(n1897), .B(n1896), .Z(n1901) );
  NANDN U2036 ( .A(n1899), .B(n1898), .Z(n1900) );
  NAND U2037 ( .A(n1901), .B(n1900), .Z(n1930) );
  XNOR U2038 ( .A(n1931), .B(n1930), .Z(n1916) );
  NANDN U2039 ( .A(n1903), .B(n1902), .Z(n1907) );
  OR U2040 ( .A(n1905), .B(n1904), .Z(n1906) );
  NAND U2041 ( .A(n1907), .B(n1906), .Z(n1917) );
  XNOR U2042 ( .A(n1916), .B(n1917), .Z(n1918) );
  XNOR U2043 ( .A(n1919), .B(n1918), .Z(n1915) );
  NAND U2044 ( .A(n1908), .B(sreg[202]), .Z(n1912) );
  OR U2045 ( .A(n1910), .B(n1909), .Z(n1911) );
  AND U2046 ( .A(n1912), .B(n1911), .Z(n1914) );
  XNOR U2047 ( .A(n1914), .B(sreg[203]), .Z(n1913) );
  XOR U2048 ( .A(n1915), .B(n1913), .Z(c[203]) );
  NANDN U2049 ( .A(n1917), .B(n1916), .Z(n1921) );
  NAND U2050 ( .A(n1919), .B(n1918), .Z(n1920) );
  NAND U2051 ( .A(n1921), .B(n1920), .Z(n1937) );
  AND U2052 ( .A(b[2]), .B(a[78]), .Z(n1943) );
  AND U2053 ( .A(a[79]), .B(b[1]), .Z(n1941) );
  AND U2054 ( .A(a[77]), .B(b[3]), .Z(n1940) );
  XOR U2055 ( .A(n1941), .B(n1940), .Z(n1942) );
  XOR U2056 ( .A(n1943), .B(n1942), .Z(n1946) );
  NAND U2057 ( .A(b[0]), .B(a[80]), .Z(n1947) );
  XOR U2058 ( .A(n1946), .B(n1947), .Z(n1949) );
  OR U2059 ( .A(n1923), .B(n1922), .Z(n1927) );
  NANDN U2060 ( .A(n1925), .B(n1924), .Z(n1926) );
  NAND U2061 ( .A(n1927), .B(n1926), .Z(n1948) );
  XNOR U2062 ( .A(n1949), .B(n1948), .Z(n1934) );
  NANDN U2063 ( .A(n1929), .B(n1928), .Z(n1933) );
  OR U2064 ( .A(n1931), .B(n1930), .Z(n1932) );
  NAND U2065 ( .A(n1933), .B(n1932), .Z(n1935) );
  XNOR U2066 ( .A(n1934), .B(n1935), .Z(n1936) );
  XOR U2067 ( .A(n1937), .B(n1936), .Z(n1952) );
  XOR U2068 ( .A(sreg[204]), .B(n1952), .Z(n1954) );
  XNOR U2069 ( .A(n1953), .B(n1954), .Z(c[204]) );
  NANDN U2070 ( .A(n1935), .B(n1934), .Z(n1939) );
  NAND U2071 ( .A(n1937), .B(n1936), .Z(n1938) );
  NAND U2072 ( .A(n1939), .B(n1938), .Z(n1960) );
  AND U2073 ( .A(b[2]), .B(a[79]), .Z(n1966) );
  AND U2074 ( .A(a[80]), .B(b[1]), .Z(n1964) );
  AND U2075 ( .A(a[78]), .B(b[3]), .Z(n1963) );
  XOR U2076 ( .A(n1964), .B(n1963), .Z(n1965) );
  XOR U2077 ( .A(n1966), .B(n1965), .Z(n1969) );
  NAND U2078 ( .A(b[0]), .B(a[81]), .Z(n1970) );
  XOR U2079 ( .A(n1969), .B(n1970), .Z(n1972) );
  OR U2080 ( .A(n1941), .B(n1940), .Z(n1945) );
  NANDN U2081 ( .A(n1943), .B(n1942), .Z(n1944) );
  NAND U2082 ( .A(n1945), .B(n1944), .Z(n1971) );
  XNOR U2083 ( .A(n1972), .B(n1971), .Z(n1957) );
  NANDN U2084 ( .A(n1947), .B(n1946), .Z(n1951) );
  OR U2085 ( .A(n1949), .B(n1948), .Z(n1950) );
  NAND U2086 ( .A(n1951), .B(n1950), .Z(n1958) );
  XNOR U2087 ( .A(n1957), .B(n1958), .Z(n1959) );
  XNOR U2088 ( .A(n1960), .B(n1959), .Z(n1975) );
  XOR U2089 ( .A(sreg[205]), .B(n1975), .Z(n1976) );
  NANDN U2090 ( .A(n1952), .B(sreg[204]), .Z(n1956) );
  NANDN U2091 ( .A(n1954), .B(n1953), .Z(n1955) );
  NAND U2092 ( .A(n1956), .B(n1955), .Z(n1977) );
  XOR U2093 ( .A(n1976), .B(n1977), .Z(c[205]) );
  NANDN U2094 ( .A(n1958), .B(n1957), .Z(n1962) );
  NAND U2095 ( .A(n1960), .B(n1959), .Z(n1961) );
  NAND U2096 ( .A(n1962), .B(n1961), .Z(n1983) );
  AND U2097 ( .A(b[2]), .B(a[80]), .Z(n1989) );
  AND U2098 ( .A(a[81]), .B(b[1]), .Z(n1987) );
  AND U2099 ( .A(a[79]), .B(b[3]), .Z(n1986) );
  XOR U2100 ( .A(n1987), .B(n1986), .Z(n1988) );
  XOR U2101 ( .A(n1989), .B(n1988), .Z(n1992) );
  NAND U2102 ( .A(b[0]), .B(a[82]), .Z(n1993) );
  XOR U2103 ( .A(n1992), .B(n1993), .Z(n1995) );
  OR U2104 ( .A(n1964), .B(n1963), .Z(n1968) );
  NANDN U2105 ( .A(n1966), .B(n1965), .Z(n1967) );
  NAND U2106 ( .A(n1968), .B(n1967), .Z(n1994) );
  XNOR U2107 ( .A(n1995), .B(n1994), .Z(n1980) );
  NANDN U2108 ( .A(n1970), .B(n1969), .Z(n1974) );
  OR U2109 ( .A(n1972), .B(n1971), .Z(n1973) );
  NAND U2110 ( .A(n1974), .B(n1973), .Z(n1981) );
  XNOR U2111 ( .A(n1980), .B(n1981), .Z(n1982) );
  XNOR U2112 ( .A(n1983), .B(n1982), .Z(n1998) );
  XOR U2113 ( .A(sreg[206]), .B(n1998), .Z(n1999) );
  OR U2114 ( .A(n1975), .B(sreg[205]), .Z(n1979) );
  NANDN U2115 ( .A(n1977), .B(n1976), .Z(n1978) );
  AND U2116 ( .A(n1979), .B(n1978), .Z(n2000) );
  XOR U2117 ( .A(n1999), .B(n2000), .Z(c[206]) );
  NANDN U2118 ( .A(n1981), .B(n1980), .Z(n1985) );
  NAND U2119 ( .A(n1983), .B(n1982), .Z(n1984) );
  NAND U2120 ( .A(n1985), .B(n1984), .Z(n2009) );
  AND U2121 ( .A(b[2]), .B(a[81]), .Z(n2015) );
  AND U2122 ( .A(a[82]), .B(b[1]), .Z(n2013) );
  AND U2123 ( .A(a[80]), .B(b[3]), .Z(n2012) );
  XOR U2124 ( .A(n2013), .B(n2012), .Z(n2014) );
  XOR U2125 ( .A(n2015), .B(n2014), .Z(n2018) );
  NAND U2126 ( .A(b[0]), .B(a[83]), .Z(n2019) );
  XOR U2127 ( .A(n2018), .B(n2019), .Z(n2021) );
  OR U2128 ( .A(n1987), .B(n1986), .Z(n1991) );
  NANDN U2129 ( .A(n1989), .B(n1988), .Z(n1990) );
  NAND U2130 ( .A(n1991), .B(n1990), .Z(n2020) );
  XNOR U2131 ( .A(n2021), .B(n2020), .Z(n2006) );
  NANDN U2132 ( .A(n1993), .B(n1992), .Z(n1997) );
  OR U2133 ( .A(n1995), .B(n1994), .Z(n1996) );
  NAND U2134 ( .A(n1997), .B(n1996), .Z(n2007) );
  XNOR U2135 ( .A(n2006), .B(n2007), .Z(n2008) );
  XOR U2136 ( .A(n2009), .B(n2008), .Z(n2005) );
  OR U2137 ( .A(n1998), .B(sreg[206]), .Z(n2002) );
  NANDN U2138 ( .A(n2000), .B(n1999), .Z(n2001) );
  AND U2139 ( .A(n2002), .B(n2001), .Z(n2004) );
  XNOR U2140 ( .A(sreg[207]), .B(n2004), .Z(n2003) );
  XOR U2141 ( .A(n2005), .B(n2003), .Z(c[207]) );
  NANDN U2142 ( .A(n2007), .B(n2006), .Z(n2011) );
  NAND U2143 ( .A(n2009), .B(n2008), .Z(n2010) );
  NAND U2144 ( .A(n2011), .B(n2010), .Z(n2027) );
  AND U2145 ( .A(b[2]), .B(a[82]), .Z(n2039) );
  AND U2146 ( .A(a[83]), .B(b[1]), .Z(n2037) );
  AND U2147 ( .A(a[81]), .B(b[3]), .Z(n2036) );
  XOR U2148 ( .A(n2037), .B(n2036), .Z(n2038) );
  XOR U2149 ( .A(n2039), .B(n2038), .Z(n2030) );
  NAND U2150 ( .A(b[0]), .B(a[84]), .Z(n2031) );
  XOR U2151 ( .A(n2030), .B(n2031), .Z(n2033) );
  OR U2152 ( .A(n2013), .B(n2012), .Z(n2017) );
  NANDN U2153 ( .A(n2015), .B(n2014), .Z(n2016) );
  NAND U2154 ( .A(n2017), .B(n2016), .Z(n2032) );
  XNOR U2155 ( .A(n2033), .B(n2032), .Z(n2024) );
  NANDN U2156 ( .A(n2019), .B(n2018), .Z(n2023) );
  OR U2157 ( .A(n2021), .B(n2020), .Z(n2022) );
  NAND U2158 ( .A(n2023), .B(n2022), .Z(n2025) );
  XNOR U2159 ( .A(n2024), .B(n2025), .Z(n2026) );
  XNOR U2160 ( .A(n2027), .B(n2026), .Z(n2042) );
  XNOR U2161 ( .A(n2042), .B(sreg[208]), .Z(n2043) );
  XOR U2162 ( .A(n2044), .B(n2043), .Z(c[208]) );
  NANDN U2163 ( .A(n2025), .B(n2024), .Z(n2029) );
  NAND U2164 ( .A(n2027), .B(n2026), .Z(n2028) );
  NAND U2165 ( .A(n2029), .B(n2028), .Z(n2062) );
  NANDN U2166 ( .A(n2031), .B(n2030), .Z(n2035) );
  OR U2167 ( .A(n2033), .B(n2032), .Z(n2034) );
  NAND U2168 ( .A(n2035), .B(n2034), .Z(n2059) );
  AND U2169 ( .A(b[2]), .B(a[83]), .Z(n2050) );
  AND U2170 ( .A(a[84]), .B(b[1]), .Z(n2048) );
  AND U2171 ( .A(a[82]), .B(b[3]), .Z(n2047) );
  XOR U2172 ( .A(n2048), .B(n2047), .Z(n2049) );
  XOR U2173 ( .A(n2050), .B(n2049), .Z(n2053) );
  NAND U2174 ( .A(b[0]), .B(a[85]), .Z(n2054) );
  XNOR U2175 ( .A(n2053), .B(n2054), .Z(n2055) );
  OR U2176 ( .A(n2037), .B(n2036), .Z(n2041) );
  NANDN U2177 ( .A(n2039), .B(n2038), .Z(n2040) );
  AND U2178 ( .A(n2041), .B(n2040), .Z(n2056) );
  XNOR U2179 ( .A(n2055), .B(n2056), .Z(n2060) );
  XNOR U2180 ( .A(n2059), .B(n2060), .Z(n2061) );
  XNOR U2181 ( .A(n2062), .B(n2061), .Z(n2065) );
  XOR U2182 ( .A(sreg[209]), .B(n2065), .Z(n2066) );
  NAND U2183 ( .A(n2042), .B(sreg[208]), .Z(n2046) );
  OR U2184 ( .A(n2044), .B(n2043), .Z(n2045) );
  NAND U2185 ( .A(n2046), .B(n2045), .Z(n2067) );
  XOR U2186 ( .A(n2066), .B(n2067), .Z(c[209]) );
  AND U2187 ( .A(b[2]), .B(a[84]), .Z(n2082) );
  AND U2188 ( .A(a[85]), .B(b[1]), .Z(n2080) );
  AND U2189 ( .A(a[83]), .B(b[3]), .Z(n2079) );
  XOR U2190 ( .A(n2080), .B(n2079), .Z(n2081) );
  XOR U2191 ( .A(n2082), .B(n2081), .Z(n2085) );
  NAND U2192 ( .A(b[0]), .B(a[86]), .Z(n2086) );
  XOR U2193 ( .A(n2085), .B(n2086), .Z(n2088) );
  OR U2194 ( .A(n2048), .B(n2047), .Z(n2052) );
  NANDN U2195 ( .A(n2050), .B(n2049), .Z(n2051) );
  NAND U2196 ( .A(n2052), .B(n2051), .Z(n2087) );
  XNOR U2197 ( .A(n2088), .B(n2087), .Z(n2073) );
  NANDN U2198 ( .A(n2054), .B(n2053), .Z(n2058) );
  NAND U2199 ( .A(n2056), .B(n2055), .Z(n2057) );
  NAND U2200 ( .A(n2058), .B(n2057), .Z(n2074) );
  XNOR U2201 ( .A(n2073), .B(n2074), .Z(n2075) );
  NANDN U2202 ( .A(n2060), .B(n2059), .Z(n2064) );
  NANDN U2203 ( .A(n2062), .B(n2061), .Z(n2063) );
  NAND U2204 ( .A(n2064), .B(n2063), .Z(n2076) );
  XOR U2205 ( .A(n2075), .B(n2076), .Z(n2072) );
  OR U2206 ( .A(n2065), .B(sreg[209]), .Z(n2069) );
  NANDN U2207 ( .A(n2067), .B(n2066), .Z(n2068) );
  AND U2208 ( .A(n2069), .B(n2068), .Z(n2071) );
  XNOR U2209 ( .A(sreg[210]), .B(n2071), .Z(n2070) );
  XNOR U2210 ( .A(n2072), .B(n2070), .Z(c[210]) );
  NANDN U2211 ( .A(n2074), .B(n2073), .Z(n2078) );
  NANDN U2212 ( .A(n2076), .B(n2075), .Z(n2077) );
  NAND U2213 ( .A(n2078), .B(n2077), .Z(n2106) );
  AND U2214 ( .A(b[2]), .B(a[85]), .Z(n2100) );
  AND U2215 ( .A(a[86]), .B(b[1]), .Z(n2098) );
  AND U2216 ( .A(a[84]), .B(b[3]), .Z(n2097) );
  XOR U2217 ( .A(n2098), .B(n2097), .Z(n2099) );
  XOR U2218 ( .A(n2100), .B(n2099), .Z(n2091) );
  NAND U2219 ( .A(b[0]), .B(a[87]), .Z(n2092) );
  XOR U2220 ( .A(n2091), .B(n2092), .Z(n2094) );
  OR U2221 ( .A(n2080), .B(n2079), .Z(n2084) );
  NANDN U2222 ( .A(n2082), .B(n2081), .Z(n2083) );
  NAND U2223 ( .A(n2084), .B(n2083), .Z(n2093) );
  XNOR U2224 ( .A(n2094), .B(n2093), .Z(n2103) );
  NANDN U2225 ( .A(n2086), .B(n2085), .Z(n2090) );
  OR U2226 ( .A(n2088), .B(n2087), .Z(n2089) );
  NAND U2227 ( .A(n2090), .B(n2089), .Z(n2104) );
  XNOR U2228 ( .A(n2103), .B(n2104), .Z(n2105) );
  XNOR U2229 ( .A(n2106), .B(n2105), .Z(n2109) );
  XNOR U2230 ( .A(n2109), .B(sreg[211]), .Z(n2110) );
  XOR U2231 ( .A(n2111), .B(n2110), .Z(c[211]) );
  NANDN U2232 ( .A(n2092), .B(n2091), .Z(n2096) );
  OR U2233 ( .A(n2094), .B(n2093), .Z(n2095) );
  NAND U2234 ( .A(n2096), .B(n2095), .Z(n2127) );
  AND U2235 ( .A(b[2]), .B(a[86]), .Z(n2118) );
  AND U2236 ( .A(a[87]), .B(b[1]), .Z(n2116) );
  AND U2237 ( .A(a[85]), .B(b[3]), .Z(n2115) );
  XOR U2238 ( .A(n2116), .B(n2115), .Z(n2117) );
  XOR U2239 ( .A(n2118), .B(n2117), .Z(n2121) );
  NAND U2240 ( .A(b[0]), .B(a[88]), .Z(n2122) );
  XNOR U2241 ( .A(n2121), .B(n2122), .Z(n2123) );
  OR U2242 ( .A(n2098), .B(n2097), .Z(n2102) );
  NANDN U2243 ( .A(n2100), .B(n2099), .Z(n2101) );
  AND U2244 ( .A(n2102), .B(n2101), .Z(n2124) );
  XNOR U2245 ( .A(n2123), .B(n2124), .Z(n2128) );
  XNOR U2246 ( .A(n2127), .B(n2128), .Z(n2129) );
  NANDN U2247 ( .A(n2104), .B(n2103), .Z(n2108) );
  NAND U2248 ( .A(n2106), .B(n2105), .Z(n2107) );
  NAND U2249 ( .A(n2108), .B(n2107), .Z(n2130) );
  XOR U2250 ( .A(n2129), .B(n2130), .Z(n2134) );
  NAND U2251 ( .A(n2109), .B(sreg[211]), .Z(n2113) );
  OR U2252 ( .A(n2111), .B(n2110), .Z(n2112) );
  AND U2253 ( .A(n2113), .B(n2112), .Z(n2133) );
  XNOR U2254 ( .A(n2133), .B(sreg[212]), .Z(n2114) );
  XNOR U2255 ( .A(n2134), .B(n2114), .Z(c[212]) );
  AND U2256 ( .A(b[2]), .B(a[87]), .Z(n2147) );
  AND U2257 ( .A(a[88]), .B(b[1]), .Z(n2145) );
  AND U2258 ( .A(a[86]), .B(b[3]), .Z(n2144) );
  XOR U2259 ( .A(n2145), .B(n2144), .Z(n2146) );
  XOR U2260 ( .A(n2147), .B(n2146), .Z(n2150) );
  NAND U2261 ( .A(b[0]), .B(a[89]), .Z(n2151) );
  XOR U2262 ( .A(n2150), .B(n2151), .Z(n2153) );
  OR U2263 ( .A(n2116), .B(n2115), .Z(n2120) );
  NANDN U2264 ( .A(n2118), .B(n2117), .Z(n2119) );
  NAND U2265 ( .A(n2120), .B(n2119), .Z(n2152) );
  XNOR U2266 ( .A(n2153), .B(n2152), .Z(n2138) );
  NANDN U2267 ( .A(n2122), .B(n2121), .Z(n2126) );
  NAND U2268 ( .A(n2124), .B(n2123), .Z(n2125) );
  NAND U2269 ( .A(n2126), .B(n2125), .Z(n2139) );
  XNOR U2270 ( .A(n2138), .B(n2139), .Z(n2140) );
  NANDN U2271 ( .A(n2128), .B(n2127), .Z(n2132) );
  NANDN U2272 ( .A(n2130), .B(n2129), .Z(n2131) );
  AND U2273 ( .A(n2132), .B(n2131), .Z(n2141) );
  XNOR U2274 ( .A(n2140), .B(n2141), .Z(n2137) );
  XOR U2275 ( .A(n2136), .B(sreg[213]), .Z(n2135) );
  XOR U2276 ( .A(n2137), .B(n2135), .Z(c[213]) );
  NANDN U2277 ( .A(n2139), .B(n2138), .Z(n2143) );
  NAND U2278 ( .A(n2141), .B(n2140), .Z(n2142) );
  NAND U2279 ( .A(n2143), .B(n2142), .Z(n2171) );
  AND U2280 ( .A(b[2]), .B(a[88]), .Z(n2165) );
  AND U2281 ( .A(a[89]), .B(b[1]), .Z(n2163) );
  AND U2282 ( .A(a[87]), .B(b[3]), .Z(n2162) );
  XOR U2283 ( .A(n2163), .B(n2162), .Z(n2164) );
  XOR U2284 ( .A(n2165), .B(n2164), .Z(n2156) );
  NAND U2285 ( .A(b[0]), .B(a[90]), .Z(n2157) );
  XOR U2286 ( .A(n2156), .B(n2157), .Z(n2159) );
  OR U2287 ( .A(n2145), .B(n2144), .Z(n2149) );
  NANDN U2288 ( .A(n2147), .B(n2146), .Z(n2148) );
  NAND U2289 ( .A(n2149), .B(n2148), .Z(n2158) );
  XNOR U2290 ( .A(n2159), .B(n2158), .Z(n2168) );
  NANDN U2291 ( .A(n2151), .B(n2150), .Z(n2155) );
  OR U2292 ( .A(n2153), .B(n2152), .Z(n2154) );
  NAND U2293 ( .A(n2155), .B(n2154), .Z(n2169) );
  XNOR U2294 ( .A(n2168), .B(n2169), .Z(n2170) );
  XNOR U2295 ( .A(n2171), .B(n2170), .Z(n2174) );
  XNOR U2296 ( .A(n2174), .B(sreg[214]), .Z(n2176) );
  XNOR U2297 ( .A(n2175), .B(n2176), .Z(c[214]) );
  NANDN U2298 ( .A(n2157), .B(n2156), .Z(n2161) );
  OR U2299 ( .A(n2159), .B(n2158), .Z(n2160) );
  NAND U2300 ( .A(n2161), .B(n2160), .Z(n2191) );
  AND U2301 ( .A(b[2]), .B(a[89]), .Z(n2182) );
  AND U2302 ( .A(a[90]), .B(b[1]), .Z(n2180) );
  AND U2303 ( .A(a[88]), .B(b[3]), .Z(n2179) );
  XOR U2304 ( .A(n2180), .B(n2179), .Z(n2181) );
  XOR U2305 ( .A(n2182), .B(n2181), .Z(n2185) );
  NAND U2306 ( .A(b[0]), .B(a[91]), .Z(n2186) );
  XNOR U2307 ( .A(n2185), .B(n2186), .Z(n2187) );
  OR U2308 ( .A(n2163), .B(n2162), .Z(n2167) );
  NANDN U2309 ( .A(n2165), .B(n2164), .Z(n2166) );
  AND U2310 ( .A(n2167), .B(n2166), .Z(n2188) );
  XNOR U2311 ( .A(n2187), .B(n2188), .Z(n2192) );
  XNOR U2312 ( .A(n2191), .B(n2192), .Z(n2193) );
  NANDN U2313 ( .A(n2169), .B(n2168), .Z(n2173) );
  NAND U2314 ( .A(n2171), .B(n2170), .Z(n2172) );
  NAND U2315 ( .A(n2173), .B(n2172), .Z(n2194) );
  XNOR U2316 ( .A(n2193), .B(n2194), .Z(n2197) );
  XOR U2317 ( .A(sreg[215]), .B(n2197), .Z(n2198) );
  NAND U2318 ( .A(n2174), .B(sreg[214]), .Z(n2178) );
  NANDN U2319 ( .A(n2176), .B(n2175), .Z(n2177) );
  NAND U2320 ( .A(n2178), .B(n2177), .Z(n2199) );
  XOR U2321 ( .A(n2198), .B(n2199), .Z(c[215]) );
  AND U2322 ( .A(b[2]), .B(a[90]), .Z(n2212) );
  AND U2323 ( .A(a[91]), .B(b[1]), .Z(n2210) );
  AND U2324 ( .A(a[89]), .B(b[3]), .Z(n2209) );
  XOR U2325 ( .A(n2210), .B(n2209), .Z(n2211) );
  XOR U2326 ( .A(n2212), .B(n2211), .Z(n2215) );
  NAND U2327 ( .A(b[0]), .B(a[92]), .Z(n2216) );
  XOR U2328 ( .A(n2215), .B(n2216), .Z(n2218) );
  OR U2329 ( .A(n2180), .B(n2179), .Z(n2184) );
  NANDN U2330 ( .A(n2182), .B(n2181), .Z(n2183) );
  NAND U2331 ( .A(n2184), .B(n2183), .Z(n2217) );
  XNOR U2332 ( .A(n2218), .B(n2217), .Z(n2203) );
  NANDN U2333 ( .A(n2186), .B(n2185), .Z(n2190) );
  NAND U2334 ( .A(n2188), .B(n2187), .Z(n2189) );
  NAND U2335 ( .A(n2190), .B(n2189), .Z(n2204) );
  XNOR U2336 ( .A(n2203), .B(n2204), .Z(n2205) );
  NANDN U2337 ( .A(n2192), .B(n2191), .Z(n2196) );
  NANDN U2338 ( .A(n2194), .B(n2193), .Z(n2195) );
  NAND U2339 ( .A(n2196), .B(n2195), .Z(n2206) );
  XOR U2340 ( .A(n2205), .B(n2206), .Z(n2222) );
  OR U2341 ( .A(n2197), .B(sreg[215]), .Z(n2201) );
  NANDN U2342 ( .A(n2199), .B(n2198), .Z(n2200) );
  AND U2343 ( .A(n2201), .B(n2200), .Z(n2221) );
  XNOR U2344 ( .A(sreg[216]), .B(n2221), .Z(n2202) );
  XNOR U2345 ( .A(n2222), .B(n2202), .Z(c[216]) );
  NANDN U2346 ( .A(n2204), .B(n2203), .Z(n2208) );
  NANDN U2347 ( .A(n2206), .B(n2205), .Z(n2207) );
  NAND U2348 ( .A(n2208), .B(n2207), .Z(n2239) );
  AND U2349 ( .A(b[2]), .B(a[91]), .Z(n2233) );
  AND U2350 ( .A(a[92]), .B(b[1]), .Z(n2231) );
  AND U2351 ( .A(a[90]), .B(b[3]), .Z(n2230) );
  XOR U2352 ( .A(n2231), .B(n2230), .Z(n2232) );
  XOR U2353 ( .A(n2233), .B(n2232), .Z(n2224) );
  NAND U2354 ( .A(b[0]), .B(a[93]), .Z(n2225) );
  XOR U2355 ( .A(n2224), .B(n2225), .Z(n2227) );
  OR U2356 ( .A(n2210), .B(n2209), .Z(n2214) );
  NANDN U2357 ( .A(n2212), .B(n2211), .Z(n2213) );
  NAND U2358 ( .A(n2214), .B(n2213), .Z(n2226) );
  XNOR U2359 ( .A(n2227), .B(n2226), .Z(n2236) );
  NANDN U2360 ( .A(n2216), .B(n2215), .Z(n2220) );
  OR U2361 ( .A(n2218), .B(n2217), .Z(n2219) );
  NAND U2362 ( .A(n2220), .B(n2219), .Z(n2237) );
  XNOR U2363 ( .A(n2236), .B(n2237), .Z(n2238) );
  XOR U2364 ( .A(n2239), .B(n2238), .Z(n2243) );
  XNOR U2365 ( .A(sreg[217]), .B(n2242), .Z(n2223) );
  XOR U2366 ( .A(n2243), .B(n2223), .Z(c[217]) );
  NANDN U2367 ( .A(n2225), .B(n2224), .Z(n2229) );
  OR U2368 ( .A(n2227), .B(n2226), .Z(n2228) );
  NAND U2369 ( .A(n2229), .B(n2228), .Z(n2257) );
  AND U2370 ( .A(b[2]), .B(a[92]), .Z(n2248) );
  AND U2371 ( .A(a[93]), .B(b[1]), .Z(n2246) );
  AND U2372 ( .A(a[91]), .B(b[3]), .Z(n2245) );
  XOR U2373 ( .A(n2246), .B(n2245), .Z(n2247) );
  XOR U2374 ( .A(n2248), .B(n2247), .Z(n2251) );
  NAND U2375 ( .A(b[0]), .B(a[94]), .Z(n2252) );
  XNOR U2376 ( .A(n2251), .B(n2252), .Z(n2253) );
  OR U2377 ( .A(n2231), .B(n2230), .Z(n2235) );
  NANDN U2378 ( .A(n2233), .B(n2232), .Z(n2234) );
  AND U2379 ( .A(n2235), .B(n2234), .Z(n2254) );
  XNOR U2380 ( .A(n2253), .B(n2254), .Z(n2258) );
  XNOR U2381 ( .A(n2257), .B(n2258), .Z(n2259) );
  NANDN U2382 ( .A(n2237), .B(n2236), .Z(n2241) );
  NAND U2383 ( .A(n2239), .B(n2238), .Z(n2240) );
  AND U2384 ( .A(n2241), .B(n2240), .Z(n2260) );
  XNOR U2385 ( .A(n2259), .B(n2260), .Z(n2266) );
  IV U2386 ( .A(n2264), .Z(n2263) );
  XNOR U2387 ( .A(n2263), .B(sreg[218]), .Z(n2244) );
  XOR U2388 ( .A(n2266), .B(n2244), .Z(c[218]) );
  AND U2389 ( .A(b[2]), .B(a[93]), .Z(n2278) );
  AND U2390 ( .A(a[94]), .B(b[1]), .Z(n2276) );
  AND U2391 ( .A(a[92]), .B(b[3]), .Z(n2275) );
  XOR U2392 ( .A(n2276), .B(n2275), .Z(n2277) );
  XOR U2393 ( .A(n2278), .B(n2277), .Z(n2281) );
  NAND U2394 ( .A(b[0]), .B(a[95]), .Z(n2282) );
  XOR U2395 ( .A(n2281), .B(n2282), .Z(n2284) );
  OR U2396 ( .A(n2246), .B(n2245), .Z(n2250) );
  NANDN U2397 ( .A(n2248), .B(n2247), .Z(n2249) );
  NAND U2398 ( .A(n2250), .B(n2249), .Z(n2283) );
  XNOR U2399 ( .A(n2284), .B(n2283), .Z(n2269) );
  NANDN U2400 ( .A(n2252), .B(n2251), .Z(n2256) );
  NAND U2401 ( .A(n2254), .B(n2253), .Z(n2255) );
  NAND U2402 ( .A(n2256), .B(n2255), .Z(n2270) );
  XNOR U2403 ( .A(n2269), .B(n2270), .Z(n2271) );
  NANDN U2404 ( .A(n2258), .B(n2257), .Z(n2262) );
  NAND U2405 ( .A(n2260), .B(n2259), .Z(n2261) );
  NAND U2406 ( .A(n2262), .B(n2261), .Z(n2272) );
  XOR U2407 ( .A(n2271), .B(n2272), .Z(n2287) );
  XNOR U2408 ( .A(n2287), .B(sreg[219]), .Z(n2289) );
  NAND U2409 ( .A(n2263), .B(sreg[218]), .Z(n2268) );
  NANDN U2410 ( .A(sreg[218]), .B(n2264), .Z(n2265) );
  NANDN U2411 ( .A(n2266), .B(n2265), .Z(n2267) );
  AND U2412 ( .A(n2268), .B(n2267), .Z(n2288) );
  XOR U2413 ( .A(n2289), .B(n2288), .Z(c[219]) );
  NANDN U2414 ( .A(n2270), .B(n2269), .Z(n2274) );
  NANDN U2415 ( .A(n2272), .B(n2271), .Z(n2273) );
  NAND U2416 ( .A(n2274), .B(n2273), .Z(n2307) );
  AND U2417 ( .A(b[2]), .B(a[94]), .Z(n2301) );
  AND U2418 ( .A(a[95]), .B(b[1]), .Z(n2299) );
  AND U2419 ( .A(a[93]), .B(b[3]), .Z(n2298) );
  XOR U2420 ( .A(n2299), .B(n2298), .Z(n2300) );
  XOR U2421 ( .A(n2301), .B(n2300), .Z(n2292) );
  NAND U2422 ( .A(b[0]), .B(a[96]), .Z(n2293) );
  XOR U2423 ( .A(n2292), .B(n2293), .Z(n2295) );
  OR U2424 ( .A(n2276), .B(n2275), .Z(n2280) );
  NANDN U2425 ( .A(n2278), .B(n2277), .Z(n2279) );
  NAND U2426 ( .A(n2280), .B(n2279), .Z(n2294) );
  XNOR U2427 ( .A(n2295), .B(n2294), .Z(n2304) );
  NANDN U2428 ( .A(n2282), .B(n2281), .Z(n2286) );
  OR U2429 ( .A(n2284), .B(n2283), .Z(n2285) );
  NAND U2430 ( .A(n2286), .B(n2285), .Z(n2305) );
  XNOR U2431 ( .A(n2304), .B(n2305), .Z(n2306) );
  XNOR U2432 ( .A(n2307), .B(n2306), .Z(n2310) );
  XOR U2433 ( .A(sreg[220]), .B(n2310), .Z(n2311) );
  NAND U2434 ( .A(n2287), .B(sreg[219]), .Z(n2291) );
  OR U2435 ( .A(n2289), .B(n2288), .Z(n2290) );
  NAND U2436 ( .A(n2291), .B(n2290), .Z(n2312) );
  XOR U2437 ( .A(n2311), .B(n2312), .Z(c[220]) );
  NANDN U2438 ( .A(n2293), .B(n2292), .Z(n2297) );
  OR U2439 ( .A(n2295), .B(n2294), .Z(n2296) );
  NAND U2440 ( .A(n2297), .B(n2296), .Z(n2316) );
  AND U2441 ( .A(b[2]), .B(a[95]), .Z(n2331) );
  AND U2442 ( .A(a[96]), .B(b[1]), .Z(n2329) );
  AND U2443 ( .A(a[94]), .B(b[3]), .Z(n2328) );
  XOR U2444 ( .A(n2329), .B(n2328), .Z(n2330) );
  XOR U2445 ( .A(n2331), .B(n2330), .Z(n2322) );
  NAND U2446 ( .A(b[0]), .B(a[97]), .Z(n2323) );
  XNOR U2447 ( .A(n2322), .B(n2323), .Z(n2324) );
  OR U2448 ( .A(n2299), .B(n2298), .Z(n2303) );
  NANDN U2449 ( .A(n2301), .B(n2300), .Z(n2302) );
  AND U2450 ( .A(n2303), .B(n2302), .Z(n2325) );
  XNOR U2451 ( .A(n2324), .B(n2325), .Z(n2317) );
  XNOR U2452 ( .A(n2316), .B(n2317), .Z(n2318) );
  NANDN U2453 ( .A(n2305), .B(n2304), .Z(n2309) );
  NAND U2454 ( .A(n2307), .B(n2306), .Z(n2308) );
  AND U2455 ( .A(n2309), .B(n2308), .Z(n2319) );
  XNOR U2456 ( .A(n2318), .B(n2319), .Z(n2336) );
  OR U2457 ( .A(n2310), .B(sreg[220]), .Z(n2314) );
  NANDN U2458 ( .A(n2312), .B(n2311), .Z(n2313) );
  AND U2459 ( .A(n2314), .B(n2313), .Z(n2335) );
  XNOR U2460 ( .A(sreg[221]), .B(n2335), .Z(n2315) );
  XOR U2461 ( .A(n2336), .B(n2315), .Z(c[221]) );
  NANDN U2462 ( .A(n2317), .B(n2316), .Z(n2321) );
  NAND U2463 ( .A(n2319), .B(n2318), .Z(n2320) );
  NAND U2464 ( .A(n2321), .B(n2320), .Z(n2340) );
  NANDN U2465 ( .A(n2323), .B(n2322), .Z(n2327) );
  NAND U2466 ( .A(n2325), .B(n2324), .Z(n2326) );
  AND U2467 ( .A(n2327), .B(n2326), .Z(n2339) );
  AND U2468 ( .A(b[2]), .B(a[96]), .Z(n2344) );
  AND U2469 ( .A(a[97]), .B(b[1]), .Z(n2342) );
  AND U2470 ( .A(a[95]), .B(b[3]), .Z(n2341) );
  XOR U2471 ( .A(n2342), .B(n2341), .Z(n2343) );
  XOR U2472 ( .A(n2344), .B(n2343), .Z(n2347) );
  NAND U2473 ( .A(b[0]), .B(a[98]), .Z(n2348) );
  XOR U2474 ( .A(n2347), .B(n2348), .Z(n2350) );
  OR U2475 ( .A(n2329), .B(n2328), .Z(n2333) );
  NANDN U2476 ( .A(n2331), .B(n2330), .Z(n2332) );
  NAND U2477 ( .A(n2333), .B(n2332), .Z(n2349) );
  XOR U2478 ( .A(n2350), .B(n2349), .Z(n2338) );
  XNOR U2479 ( .A(n2339), .B(n2338), .Z(n2334) );
  XOR U2480 ( .A(n2340), .B(n2334), .Z(n2354) );
  XNOR U2481 ( .A(sreg[222]), .B(n2353), .Z(n2337) );
  XNOR U2482 ( .A(n2354), .B(n2337), .Z(c[222]) );
  AND U2483 ( .A(b[2]), .B(a[97]), .Z(n2365) );
  AND U2484 ( .A(a[98]), .B(b[1]), .Z(n2363) );
  AND U2485 ( .A(a[96]), .B(b[3]), .Z(n2362) );
  XOR U2486 ( .A(n2363), .B(n2362), .Z(n2364) );
  XOR U2487 ( .A(n2365), .B(n2364), .Z(n2368) );
  NAND U2488 ( .A(b[0]), .B(a[99]), .Z(n2369) );
  XOR U2489 ( .A(n2368), .B(n2369), .Z(n2371) );
  OR U2490 ( .A(n2342), .B(n2341), .Z(n2346) );
  NANDN U2491 ( .A(n2344), .B(n2343), .Z(n2345) );
  NAND U2492 ( .A(n2346), .B(n2345), .Z(n2370) );
  XNOR U2493 ( .A(n2371), .B(n2370), .Z(n2356) );
  NANDN U2494 ( .A(n2348), .B(n2347), .Z(n2352) );
  OR U2495 ( .A(n2350), .B(n2349), .Z(n2351) );
  NAND U2496 ( .A(n2352), .B(n2351), .Z(n2357) );
  XNOR U2497 ( .A(n2356), .B(n2357), .Z(n2358) );
  XOR U2498 ( .A(n2359), .B(n2358), .Z(n2376) );
  XNOR U2499 ( .A(sreg[223]), .B(n2375), .Z(n2355) );
  XNOR U2500 ( .A(n2376), .B(n2355), .Z(c[223]) );
  NANDN U2501 ( .A(n2357), .B(n2356), .Z(n2361) );
  NANDN U2502 ( .A(n2359), .B(n2358), .Z(n2360) );
  AND U2503 ( .A(n2361), .B(n2360), .Z(n2392) );
  AND U2504 ( .A(b[2]), .B(a[98]), .Z(n2387) );
  AND U2505 ( .A(a[99]), .B(b[1]), .Z(n2385) );
  AND U2506 ( .A(a[97]), .B(b[3]), .Z(n2384) );
  XOR U2507 ( .A(n2385), .B(n2384), .Z(n2386) );
  XOR U2508 ( .A(n2387), .B(n2386), .Z(n2380) );
  NAND U2509 ( .A(b[0]), .B(a[100]), .Z(n2381) );
  XOR U2510 ( .A(n2380), .B(n2381), .Z(n2382) );
  OR U2511 ( .A(n2363), .B(n2362), .Z(n2367) );
  NANDN U2512 ( .A(n2365), .B(n2364), .Z(n2366) );
  AND U2513 ( .A(n2367), .B(n2366), .Z(n2383) );
  XOR U2514 ( .A(n2382), .B(n2383), .Z(n2390) );
  NANDN U2515 ( .A(n2369), .B(n2368), .Z(n2373) );
  OR U2516 ( .A(n2371), .B(n2370), .Z(n2372) );
  AND U2517 ( .A(n2373), .B(n2372), .Z(n2391) );
  XOR U2518 ( .A(n2390), .B(n2391), .Z(n2374) );
  XNOR U2519 ( .A(n2392), .B(n2374), .Z(n2379) );
  XNOR U2520 ( .A(sreg[224]), .B(n2378), .Z(n2377) );
  XOR U2521 ( .A(n2379), .B(n2377), .Z(c[224]) );
  AND U2522 ( .A(b[2]), .B(a[99]), .Z(n2400) );
  AND U2523 ( .A(a[100]), .B(b[1]), .Z(n2398) );
  AND U2524 ( .A(a[98]), .B(b[3]), .Z(n2397) );
  XOR U2525 ( .A(n2398), .B(n2397), .Z(n2399) );
  XOR U2526 ( .A(n2400), .B(n2399), .Z(n2403) );
  NAND U2527 ( .A(b[0]), .B(a[101]), .Z(n2404) );
  XOR U2528 ( .A(n2403), .B(n2404), .Z(n2405) );
  OR U2529 ( .A(n2385), .B(n2384), .Z(n2389) );
  NANDN U2530 ( .A(n2387), .B(n2386), .Z(n2388) );
  AND U2531 ( .A(n2389), .B(n2388), .Z(n2406) );
  XOR U2532 ( .A(n2405), .B(n2406), .Z(n2395) );
  XNOR U2533 ( .A(n2395), .B(n2396), .Z(n2393) );
  XOR U2534 ( .A(n2394), .B(n2393), .Z(n2407) );
  XNOR U2535 ( .A(sreg[225]), .B(n2407), .Z(n2408) );
  XOR U2536 ( .A(n2409), .B(n2408), .Z(c[225]) );
  AND U2537 ( .A(b[2]), .B(a[100]), .Z(n2426) );
  AND U2538 ( .A(a[101]), .B(b[1]), .Z(n2424) );
  AND U2539 ( .A(a[99]), .B(b[3]), .Z(n2423) );
  XOR U2540 ( .A(n2424), .B(n2423), .Z(n2425) );
  XOR U2541 ( .A(n2426), .B(n2425), .Z(n2429) );
  NAND U2542 ( .A(b[0]), .B(a[102]), .Z(n2430) );
  XOR U2543 ( .A(n2429), .B(n2430), .Z(n2432) );
  OR U2544 ( .A(n2398), .B(n2397), .Z(n2402) );
  NANDN U2545 ( .A(n2400), .B(n2399), .Z(n2401) );
  NAND U2546 ( .A(n2402), .B(n2401), .Z(n2431) );
  XNOR U2547 ( .A(n2432), .B(n2431), .Z(n2417) );
  XNOR U2548 ( .A(n2417), .B(n2418), .Z(n2420) );
  XOR U2549 ( .A(n2419), .B(n2420), .Z(n2412) );
  XOR U2550 ( .A(sreg[226]), .B(n2412), .Z(n2414) );
  NAND U2551 ( .A(sreg[225]), .B(n2407), .Z(n2411) );
  OR U2552 ( .A(n2409), .B(n2408), .Z(n2410) );
  NAND U2553 ( .A(n2411), .B(n2410), .Z(n2413) );
  XNOR U2554 ( .A(n2414), .B(n2413), .Z(c[226]) );
  NANDN U2555 ( .A(sreg[226]), .B(n2412), .Z(n2416) );
  OR U2556 ( .A(n2414), .B(n2413), .Z(n2415) );
  AND U2557 ( .A(n2416), .B(n2415), .Z(n2454) );
  NANDN U2558 ( .A(n2418), .B(n2417), .Z(n2422) );
  NAND U2559 ( .A(n2420), .B(n2419), .Z(n2421) );
  NAND U2560 ( .A(n2422), .B(n2421), .Z(n2439) );
  AND U2561 ( .A(b[2]), .B(a[101]), .Z(n2445) );
  AND U2562 ( .A(a[102]), .B(b[1]), .Z(n2443) );
  AND U2563 ( .A(a[100]), .B(b[3]), .Z(n2442) );
  XOR U2564 ( .A(n2443), .B(n2442), .Z(n2444) );
  XOR U2565 ( .A(n2445), .B(n2444), .Z(n2448) );
  NAND U2566 ( .A(b[0]), .B(a[103]), .Z(n2449) );
  XOR U2567 ( .A(n2448), .B(n2449), .Z(n2451) );
  OR U2568 ( .A(n2424), .B(n2423), .Z(n2428) );
  NANDN U2569 ( .A(n2426), .B(n2425), .Z(n2427) );
  NAND U2570 ( .A(n2428), .B(n2427), .Z(n2450) );
  XNOR U2571 ( .A(n2451), .B(n2450), .Z(n2436) );
  NANDN U2572 ( .A(n2430), .B(n2429), .Z(n2434) );
  OR U2573 ( .A(n2432), .B(n2431), .Z(n2433) );
  NAND U2574 ( .A(n2434), .B(n2433), .Z(n2437) );
  XNOR U2575 ( .A(n2436), .B(n2437), .Z(n2438) );
  XNOR U2576 ( .A(n2439), .B(n2438), .Z(n2455) );
  XOR U2577 ( .A(sreg[227]), .B(n2455), .Z(n2435) );
  XOR U2578 ( .A(n2454), .B(n2435), .Z(c[227]) );
  NANDN U2579 ( .A(n2437), .B(n2436), .Z(n2441) );
  NAND U2580 ( .A(n2439), .B(n2438), .Z(n2440) );
  NAND U2581 ( .A(n2441), .B(n2440), .Z(n2462) );
  AND U2582 ( .A(b[2]), .B(a[102]), .Z(n2468) );
  AND U2583 ( .A(a[103]), .B(b[1]), .Z(n2466) );
  AND U2584 ( .A(a[101]), .B(b[3]), .Z(n2465) );
  XOR U2585 ( .A(n2466), .B(n2465), .Z(n2467) );
  XOR U2586 ( .A(n2468), .B(n2467), .Z(n2471) );
  NAND U2587 ( .A(b[0]), .B(a[104]), .Z(n2472) );
  XOR U2588 ( .A(n2471), .B(n2472), .Z(n2474) );
  OR U2589 ( .A(n2443), .B(n2442), .Z(n2447) );
  NANDN U2590 ( .A(n2445), .B(n2444), .Z(n2446) );
  NAND U2591 ( .A(n2447), .B(n2446), .Z(n2473) );
  XNOR U2592 ( .A(n2474), .B(n2473), .Z(n2459) );
  NANDN U2593 ( .A(n2449), .B(n2448), .Z(n2453) );
  OR U2594 ( .A(n2451), .B(n2450), .Z(n2452) );
  NAND U2595 ( .A(n2453), .B(n2452), .Z(n2460) );
  XNOR U2596 ( .A(n2459), .B(n2460), .Z(n2461) );
  XNOR U2597 ( .A(n2462), .B(n2461), .Z(n2458) );
  XOR U2598 ( .A(n2457), .B(sreg[228]), .Z(n2456) );
  XOR U2599 ( .A(n2458), .B(n2456), .Z(c[228]) );
  NANDN U2600 ( .A(n2460), .B(n2459), .Z(n2464) );
  NAND U2601 ( .A(n2462), .B(n2461), .Z(n2463) );
  NAND U2602 ( .A(n2464), .B(n2463), .Z(n2485) );
  AND U2603 ( .A(b[2]), .B(a[103]), .Z(n2491) );
  AND U2604 ( .A(a[104]), .B(b[1]), .Z(n2489) );
  AND U2605 ( .A(a[102]), .B(b[3]), .Z(n2488) );
  XOR U2606 ( .A(n2489), .B(n2488), .Z(n2490) );
  XOR U2607 ( .A(n2491), .B(n2490), .Z(n2494) );
  NAND U2608 ( .A(b[0]), .B(a[105]), .Z(n2495) );
  XOR U2609 ( .A(n2494), .B(n2495), .Z(n2497) );
  OR U2610 ( .A(n2466), .B(n2465), .Z(n2470) );
  NANDN U2611 ( .A(n2468), .B(n2467), .Z(n2469) );
  NAND U2612 ( .A(n2470), .B(n2469), .Z(n2496) );
  XNOR U2613 ( .A(n2497), .B(n2496), .Z(n2482) );
  NANDN U2614 ( .A(n2472), .B(n2471), .Z(n2476) );
  OR U2615 ( .A(n2474), .B(n2473), .Z(n2475) );
  NAND U2616 ( .A(n2476), .B(n2475), .Z(n2483) );
  XNOR U2617 ( .A(n2482), .B(n2483), .Z(n2484) );
  XNOR U2618 ( .A(n2485), .B(n2484), .Z(n2477) );
  XNOR U2619 ( .A(n2477), .B(sreg[229]), .Z(n2479) );
  XNOR U2620 ( .A(n2478), .B(n2479), .Z(c[229]) );
  NAND U2621 ( .A(n2477), .B(sreg[229]), .Z(n2481) );
  NANDN U2622 ( .A(n2479), .B(n2478), .Z(n2480) );
  AND U2623 ( .A(n2481), .B(n2480), .Z(n2502) );
  NANDN U2624 ( .A(n2483), .B(n2482), .Z(n2487) );
  NAND U2625 ( .A(n2485), .B(n2484), .Z(n2486) );
  NAND U2626 ( .A(n2487), .B(n2486), .Z(n2506) );
  AND U2627 ( .A(b[2]), .B(a[104]), .Z(n2512) );
  AND U2628 ( .A(a[105]), .B(b[1]), .Z(n2510) );
  AND U2629 ( .A(a[103]), .B(b[3]), .Z(n2509) );
  XOR U2630 ( .A(n2510), .B(n2509), .Z(n2511) );
  XOR U2631 ( .A(n2512), .B(n2511), .Z(n2515) );
  NAND U2632 ( .A(b[0]), .B(a[106]), .Z(n2516) );
  XOR U2633 ( .A(n2515), .B(n2516), .Z(n2518) );
  OR U2634 ( .A(n2489), .B(n2488), .Z(n2493) );
  NANDN U2635 ( .A(n2491), .B(n2490), .Z(n2492) );
  NAND U2636 ( .A(n2493), .B(n2492), .Z(n2517) );
  XNOR U2637 ( .A(n2518), .B(n2517), .Z(n2503) );
  NANDN U2638 ( .A(n2495), .B(n2494), .Z(n2499) );
  OR U2639 ( .A(n2497), .B(n2496), .Z(n2498) );
  NAND U2640 ( .A(n2499), .B(n2498), .Z(n2504) );
  XNOR U2641 ( .A(n2503), .B(n2504), .Z(n2505) );
  XNOR U2642 ( .A(n2506), .B(n2505), .Z(n2501) );
  XNOR U2643 ( .A(sreg[230]), .B(n2501), .Z(n2500) );
  XOR U2644 ( .A(n2502), .B(n2500), .Z(c[230]) );
  NANDN U2645 ( .A(n2504), .B(n2503), .Z(n2508) );
  NAND U2646 ( .A(n2506), .B(n2505), .Z(n2507) );
  NAND U2647 ( .A(n2508), .B(n2507), .Z(n2524) );
  AND U2648 ( .A(b[2]), .B(a[105]), .Z(n2530) );
  AND U2649 ( .A(a[106]), .B(b[1]), .Z(n2528) );
  AND U2650 ( .A(a[104]), .B(b[3]), .Z(n2527) );
  XOR U2651 ( .A(n2528), .B(n2527), .Z(n2529) );
  XOR U2652 ( .A(n2530), .B(n2529), .Z(n2533) );
  NAND U2653 ( .A(b[0]), .B(a[107]), .Z(n2534) );
  XOR U2654 ( .A(n2533), .B(n2534), .Z(n2536) );
  OR U2655 ( .A(n2510), .B(n2509), .Z(n2514) );
  NANDN U2656 ( .A(n2512), .B(n2511), .Z(n2513) );
  NAND U2657 ( .A(n2514), .B(n2513), .Z(n2535) );
  XNOR U2658 ( .A(n2536), .B(n2535), .Z(n2521) );
  NANDN U2659 ( .A(n2516), .B(n2515), .Z(n2520) );
  OR U2660 ( .A(n2518), .B(n2517), .Z(n2519) );
  NAND U2661 ( .A(n2520), .B(n2519), .Z(n2522) );
  XNOR U2662 ( .A(n2521), .B(n2522), .Z(n2523) );
  XNOR U2663 ( .A(n2524), .B(n2523), .Z(n2539) );
  XNOR U2664 ( .A(n2539), .B(sreg[231]), .Z(n2540) );
  XOR U2665 ( .A(n2541), .B(n2540), .Z(c[231]) );
  NANDN U2666 ( .A(n2522), .B(n2521), .Z(n2526) );
  NAND U2667 ( .A(n2524), .B(n2523), .Z(n2525) );
  NAND U2668 ( .A(n2526), .B(n2525), .Z(n2548) );
  AND U2669 ( .A(b[2]), .B(a[106]), .Z(n2554) );
  AND U2670 ( .A(a[107]), .B(b[1]), .Z(n2552) );
  AND U2671 ( .A(a[105]), .B(b[3]), .Z(n2551) );
  XOR U2672 ( .A(n2552), .B(n2551), .Z(n2553) );
  XOR U2673 ( .A(n2554), .B(n2553), .Z(n2557) );
  NAND U2674 ( .A(b[0]), .B(a[108]), .Z(n2558) );
  XOR U2675 ( .A(n2557), .B(n2558), .Z(n2560) );
  OR U2676 ( .A(n2528), .B(n2527), .Z(n2532) );
  NANDN U2677 ( .A(n2530), .B(n2529), .Z(n2531) );
  NAND U2678 ( .A(n2532), .B(n2531), .Z(n2559) );
  XNOR U2679 ( .A(n2560), .B(n2559), .Z(n2545) );
  NANDN U2680 ( .A(n2534), .B(n2533), .Z(n2538) );
  OR U2681 ( .A(n2536), .B(n2535), .Z(n2537) );
  NAND U2682 ( .A(n2538), .B(n2537), .Z(n2546) );
  XNOR U2683 ( .A(n2545), .B(n2546), .Z(n2547) );
  XOR U2684 ( .A(n2548), .B(n2547), .Z(n2564) );
  NAND U2685 ( .A(n2539), .B(sreg[231]), .Z(n2543) );
  OR U2686 ( .A(n2541), .B(n2540), .Z(n2542) );
  NAND U2687 ( .A(n2543), .B(n2542), .Z(n2563) );
  XNOR U2688 ( .A(sreg[232]), .B(n2563), .Z(n2544) );
  XOR U2689 ( .A(n2564), .B(n2544), .Z(c[232]) );
  NANDN U2690 ( .A(n2546), .B(n2545), .Z(n2550) );
  NAND U2691 ( .A(n2548), .B(n2547), .Z(n2549) );
  NAND U2692 ( .A(n2550), .B(n2549), .Z(n2571) );
  AND U2693 ( .A(b[2]), .B(a[107]), .Z(n2577) );
  AND U2694 ( .A(a[108]), .B(b[1]), .Z(n2575) );
  AND U2695 ( .A(a[106]), .B(b[3]), .Z(n2574) );
  XOR U2696 ( .A(n2575), .B(n2574), .Z(n2576) );
  XOR U2697 ( .A(n2577), .B(n2576), .Z(n2580) );
  NAND U2698 ( .A(b[0]), .B(a[109]), .Z(n2581) );
  XOR U2699 ( .A(n2580), .B(n2581), .Z(n2583) );
  OR U2700 ( .A(n2552), .B(n2551), .Z(n2556) );
  NANDN U2701 ( .A(n2554), .B(n2553), .Z(n2555) );
  NAND U2702 ( .A(n2556), .B(n2555), .Z(n2582) );
  XNOR U2703 ( .A(n2583), .B(n2582), .Z(n2568) );
  NANDN U2704 ( .A(n2558), .B(n2557), .Z(n2562) );
  OR U2705 ( .A(n2560), .B(n2559), .Z(n2561) );
  NAND U2706 ( .A(n2562), .B(n2561), .Z(n2569) );
  XNOR U2707 ( .A(n2568), .B(n2569), .Z(n2570) );
  XNOR U2708 ( .A(n2571), .B(n2570), .Z(n2567) );
  XOR U2709 ( .A(n2566), .B(sreg[233]), .Z(n2565) );
  XOR U2710 ( .A(n2567), .B(n2565), .Z(c[233]) );
  NANDN U2711 ( .A(n2569), .B(n2568), .Z(n2573) );
  NAND U2712 ( .A(n2571), .B(n2570), .Z(n2572) );
  NAND U2713 ( .A(n2573), .B(n2572), .Z(n2589) );
  AND U2714 ( .A(b[2]), .B(a[108]), .Z(n2595) );
  AND U2715 ( .A(a[109]), .B(b[1]), .Z(n2593) );
  AND U2716 ( .A(a[107]), .B(b[3]), .Z(n2592) );
  XOR U2717 ( .A(n2593), .B(n2592), .Z(n2594) );
  XOR U2718 ( .A(n2595), .B(n2594), .Z(n2598) );
  NAND U2719 ( .A(b[0]), .B(a[110]), .Z(n2599) );
  XOR U2720 ( .A(n2598), .B(n2599), .Z(n2601) );
  OR U2721 ( .A(n2575), .B(n2574), .Z(n2579) );
  NANDN U2722 ( .A(n2577), .B(n2576), .Z(n2578) );
  NAND U2723 ( .A(n2579), .B(n2578), .Z(n2600) );
  XNOR U2724 ( .A(n2601), .B(n2600), .Z(n2586) );
  NANDN U2725 ( .A(n2581), .B(n2580), .Z(n2585) );
  OR U2726 ( .A(n2583), .B(n2582), .Z(n2584) );
  NAND U2727 ( .A(n2585), .B(n2584), .Z(n2587) );
  XNOR U2728 ( .A(n2586), .B(n2587), .Z(n2588) );
  XNOR U2729 ( .A(n2589), .B(n2588), .Z(n2604) );
  XNOR U2730 ( .A(n2604), .B(sreg[234]), .Z(n2606) );
  XNOR U2731 ( .A(n2605), .B(n2606), .Z(c[234]) );
  NANDN U2732 ( .A(n2587), .B(n2586), .Z(n2591) );
  NAND U2733 ( .A(n2589), .B(n2588), .Z(n2590) );
  NAND U2734 ( .A(n2591), .B(n2590), .Z(n2612) );
  AND U2735 ( .A(b[2]), .B(a[109]), .Z(n2618) );
  AND U2736 ( .A(a[110]), .B(b[1]), .Z(n2616) );
  AND U2737 ( .A(a[108]), .B(b[3]), .Z(n2615) );
  XOR U2738 ( .A(n2616), .B(n2615), .Z(n2617) );
  XOR U2739 ( .A(n2618), .B(n2617), .Z(n2621) );
  NAND U2740 ( .A(b[0]), .B(a[111]), .Z(n2622) );
  XOR U2741 ( .A(n2621), .B(n2622), .Z(n2624) );
  OR U2742 ( .A(n2593), .B(n2592), .Z(n2597) );
  NANDN U2743 ( .A(n2595), .B(n2594), .Z(n2596) );
  NAND U2744 ( .A(n2597), .B(n2596), .Z(n2623) );
  XNOR U2745 ( .A(n2624), .B(n2623), .Z(n2609) );
  NANDN U2746 ( .A(n2599), .B(n2598), .Z(n2603) );
  OR U2747 ( .A(n2601), .B(n2600), .Z(n2602) );
  NAND U2748 ( .A(n2603), .B(n2602), .Z(n2610) );
  XNOR U2749 ( .A(n2609), .B(n2610), .Z(n2611) );
  XNOR U2750 ( .A(n2612), .B(n2611), .Z(n2627) );
  XNOR U2751 ( .A(n2627), .B(sreg[235]), .Z(n2629) );
  NAND U2752 ( .A(n2604), .B(sreg[234]), .Z(n2608) );
  NANDN U2753 ( .A(n2606), .B(n2605), .Z(n2607) );
  AND U2754 ( .A(n2608), .B(n2607), .Z(n2628) );
  XOR U2755 ( .A(n2629), .B(n2628), .Z(c[235]) );
  NANDN U2756 ( .A(n2610), .B(n2609), .Z(n2614) );
  NAND U2757 ( .A(n2612), .B(n2611), .Z(n2613) );
  NAND U2758 ( .A(n2614), .B(n2613), .Z(n2638) );
  AND U2759 ( .A(b[2]), .B(a[110]), .Z(n2644) );
  AND U2760 ( .A(a[111]), .B(b[1]), .Z(n2642) );
  AND U2761 ( .A(a[109]), .B(b[3]), .Z(n2641) );
  XOR U2762 ( .A(n2642), .B(n2641), .Z(n2643) );
  XOR U2763 ( .A(n2644), .B(n2643), .Z(n2647) );
  NAND U2764 ( .A(b[0]), .B(a[112]), .Z(n2648) );
  XOR U2765 ( .A(n2647), .B(n2648), .Z(n2650) );
  OR U2766 ( .A(n2616), .B(n2615), .Z(n2620) );
  NANDN U2767 ( .A(n2618), .B(n2617), .Z(n2619) );
  NAND U2768 ( .A(n2620), .B(n2619), .Z(n2649) );
  XNOR U2769 ( .A(n2650), .B(n2649), .Z(n2635) );
  NANDN U2770 ( .A(n2622), .B(n2621), .Z(n2626) );
  OR U2771 ( .A(n2624), .B(n2623), .Z(n2625) );
  NAND U2772 ( .A(n2626), .B(n2625), .Z(n2636) );
  XNOR U2773 ( .A(n2635), .B(n2636), .Z(n2637) );
  XOR U2774 ( .A(n2638), .B(n2637), .Z(n2634) );
  NAND U2775 ( .A(n2627), .B(sreg[235]), .Z(n2631) );
  OR U2776 ( .A(n2629), .B(n2628), .Z(n2630) );
  NAND U2777 ( .A(n2631), .B(n2630), .Z(n2633) );
  XNOR U2778 ( .A(sreg[236]), .B(n2633), .Z(n2632) );
  XOR U2779 ( .A(n2634), .B(n2632), .Z(c[236]) );
  NANDN U2780 ( .A(n2636), .B(n2635), .Z(n2640) );
  NAND U2781 ( .A(n2638), .B(n2637), .Z(n2639) );
  NAND U2782 ( .A(n2640), .B(n2639), .Z(n2656) );
  AND U2783 ( .A(b[2]), .B(a[111]), .Z(n2662) );
  AND U2784 ( .A(a[112]), .B(b[1]), .Z(n2660) );
  AND U2785 ( .A(a[110]), .B(b[3]), .Z(n2659) );
  XOR U2786 ( .A(n2660), .B(n2659), .Z(n2661) );
  XOR U2787 ( .A(n2662), .B(n2661), .Z(n2665) );
  NAND U2788 ( .A(b[0]), .B(a[113]), .Z(n2666) );
  XOR U2789 ( .A(n2665), .B(n2666), .Z(n2668) );
  OR U2790 ( .A(n2642), .B(n2641), .Z(n2646) );
  NANDN U2791 ( .A(n2644), .B(n2643), .Z(n2645) );
  NAND U2792 ( .A(n2646), .B(n2645), .Z(n2667) );
  XNOR U2793 ( .A(n2668), .B(n2667), .Z(n2653) );
  NANDN U2794 ( .A(n2648), .B(n2647), .Z(n2652) );
  OR U2795 ( .A(n2650), .B(n2649), .Z(n2651) );
  NAND U2796 ( .A(n2652), .B(n2651), .Z(n2654) );
  XNOR U2797 ( .A(n2653), .B(n2654), .Z(n2655) );
  XNOR U2798 ( .A(n2656), .B(n2655), .Z(n2671) );
  XNOR U2799 ( .A(n2671), .B(sreg[237]), .Z(n2672) );
  XOR U2800 ( .A(n2673), .B(n2672), .Z(c[237]) );
  NANDN U2801 ( .A(n2654), .B(n2653), .Z(n2658) );
  NAND U2802 ( .A(n2656), .B(n2655), .Z(n2657) );
  NAND U2803 ( .A(n2658), .B(n2657), .Z(n2679) );
  AND U2804 ( .A(b[2]), .B(a[112]), .Z(n2685) );
  AND U2805 ( .A(a[113]), .B(b[1]), .Z(n2683) );
  AND U2806 ( .A(a[111]), .B(b[3]), .Z(n2682) );
  XOR U2807 ( .A(n2683), .B(n2682), .Z(n2684) );
  XOR U2808 ( .A(n2685), .B(n2684), .Z(n2688) );
  NAND U2809 ( .A(b[0]), .B(a[114]), .Z(n2689) );
  XOR U2810 ( .A(n2688), .B(n2689), .Z(n2691) );
  OR U2811 ( .A(n2660), .B(n2659), .Z(n2664) );
  NANDN U2812 ( .A(n2662), .B(n2661), .Z(n2663) );
  NAND U2813 ( .A(n2664), .B(n2663), .Z(n2690) );
  XNOR U2814 ( .A(n2691), .B(n2690), .Z(n2676) );
  NANDN U2815 ( .A(n2666), .B(n2665), .Z(n2670) );
  OR U2816 ( .A(n2668), .B(n2667), .Z(n2669) );
  NAND U2817 ( .A(n2670), .B(n2669), .Z(n2677) );
  XNOR U2818 ( .A(n2676), .B(n2677), .Z(n2678) );
  XNOR U2819 ( .A(n2679), .B(n2678), .Z(n2694) );
  XNOR U2820 ( .A(n2694), .B(sreg[238]), .Z(n2696) );
  NAND U2821 ( .A(n2671), .B(sreg[237]), .Z(n2675) );
  OR U2822 ( .A(n2673), .B(n2672), .Z(n2674) );
  AND U2823 ( .A(n2675), .B(n2674), .Z(n2695) );
  XOR U2824 ( .A(n2696), .B(n2695), .Z(c[238]) );
  NANDN U2825 ( .A(n2677), .B(n2676), .Z(n2681) );
  NAND U2826 ( .A(n2679), .B(n2678), .Z(n2680) );
  NAND U2827 ( .A(n2681), .B(n2680), .Z(n2703) );
  AND U2828 ( .A(b[2]), .B(a[113]), .Z(n2709) );
  AND U2829 ( .A(a[114]), .B(b[1]), .Z(n2707) );
  AND U2830 ( .A(a[112]), .B(b[3]), .Z(n2706) );
  XOR U2831 ( .A(n2707), .B(n2706), .Z(n2708) );
  XOR U2832 ( .A(n2709), .B(n2708), .Z(n2712) );
  NAND U2833 ( .A(b[0]), .B(a[115]), .Z(n2713) );
  XOR U2834 ( .A(n2712), .B(n2713), .Z(n2715) );
  OR U2835 ( .A(n2683), .B(n2682), .Z(n2687) );
  NANDN U2836 ( .A(n2685), .B(n2684), .Z(n2686) );
  NAND U2837 ( .A(n2687), .B(n2686), .Z(n2714) );
  XNOR U2838 ( .A(n2715), .B(n2714), .Z(n2700) );
  NANDN U2839 ( .A(n2689), .B(n2688), .Z(n2693) );
  OR U2840 ( .A(n2691), .B(n2690), .Z(n2692) );
  NAND U2841 ( .A(n2693), .B(n2692), .Z(n2701) );
  XNOR U2842 ( .A(n2700), .B(n2701), .Z(n2702) );
  XOR U2843 ( .A(n2703), .B(n2702), .Z(n2719) );
  NAND U2844 ( .A(n2694), .B(sreg[238]), .Z(n2698) );
  OR U2845 ( .A(n2696), .B(n2695), .Z(n2697) );
  NAND U2846 ( .A(n2698), .B(n2697), .Z(n2718) );
  XNOR U2847 ( .A(sreg[239]), .B(n2718), .Z(n2699) );
  XOR U2848 ( .A(n2719), .B(n2699), .Z(c[239]) );
  NANDN U2849 ( .A(n2701), .B(n2700), .Z(n2705) );
  NAND U2850 ( .A(n2703), .B(n2702), .Z(n2704) );
  NAND U2851 ( .A(n2705), .B(n2704), .Z(n2724) );
  AND U2852 ( .A(b[2]), .B(a[114]), .Z(n2736) );
  AND U2853 ( .A(a[115]), .B(b[1]), .Z(n2734) );
  AND U2854 ( .A(a[113]), .B(b[3]), .Z(n2733) );
  XOR U2855 ( .A(n2734), .B(n2733), .Z(n2735) );
  XOR U2856 ( .A(n2736), .B(n2735), .Z(n2727) );
  NAND U2857 ( .A(b[0]), .B(a[116]), .Z(n2728) );
  XOR U2858 ( .A(n2727), .B(n2728), .Z(n2730) );
  OR U2859 ( .A(n2707), .B(n2706), .Z(n2711) );
  NANDN U2860 ( .A(n2709), .B(n2708), .Z(n2710) );
  NAND U2861 ( .A(n2711), .B(n2710), .Z(n2729) );
  XNOR U2862 ( .A(n2730), .B(n2729), .Z(n2721) );
  NANDN U2863 ( .A(n2713), .B(n2712), .Z(n2717) );
  OR U2864 ( .A(n2715), .B(n2714), .Z(n2716) );
  NAND U2865 ( .A(n2717), .B(n2716), .Z(n2722) );
  XNOR U2866 ( .A(n2721), .B(n2722), .Z(n2723) );
  XNOR U2867 ( .A(n2724), .B(n2723), .Z(n2740) );
  XOR U2868 ( .A(n2739), .B(sreg[240]), .Z(n2720) );
  XOR U2869 ( .A(n2740), .B(n2720), .Z(c[240]) );
  NANDN U2870 ( .A(n2722), .B(n2721), .Z(n2726) );
  NAND U2871 ( .A(n2724), .B(n2723), .Z(n2725) );
  NAND U2872 ( .A(n2726), .B(n2725), .Z(n2757) );
  NANDN U2873 ( .A(n2728), .B(n2727), .Z(n2732) );
  OR U2874 ( .A(n2730), .B(n2729), .Z(n2731) );
  NAND U2875 ( .A(n2732), .B(n2731), .Z(n2754) );
  AND U2876 ( .A(b[2]), .B(a[115]), .Z(n2745) );
  AND U2877 ( .A(a[116]), .B(b[1]), .Z(n2743) );
  AND U2878 ( .A(a[114]), .B(b[3]), .Z(n2742) );
  XOR U2879 ( .A(n2743), .B(n2742), .Z(n2744) );
  XOR U2880 ( .A(n2745), .B(n2744), .Z(n2748) );
  NAND U2881 ( .A(b[0]), .B(a[117]), .Z(n2749) );
  XNOR U2882 ( .A(n2748), .B(n2749), .Z(n2750) );
  OR U2883 ( .A(n2734), .B(n2733), .Z(n2738) );
  NANDN U2884 ( .A(n2736), .B(n2735), .Z(n2737) );
  AND U2885 ( .A(n2738), .B(n2737), .Z(n2751) );
  XNOR U2886 ( .A(n2750), .B(n2751), .Z(n2755) );
  XNOR U2887 ( .A(n2754), .B(n2755), .Z(n2756) );
  XOR U2888 ( .A(n2757), .B(n2756), .Z(n2761) );
  XOR U2889 ( .A(n2760), .B(sreg[241]), .Z(n2741) );
  XNOR U2890 ( .A(n2761), .B(n2741), .Z(c[241]) );
  AND U2891 ( .A(b[2]), .B(a[116]), .Z(n2774) );
  AND U2892 ( .A(a[117]), .B(b[1]), .Z(n2772) );
  AND U2893 ( .A(a[115]), .B(b[3]), .Z(n2771) );
  XOR U2894 ( .A(n2772), .B(n2771), .Z(n2773) );
  XOR U2895 ( .A(n2774), .B(n2773), .Z(n2777) );
  NAND U2896 ( .A(b[0]), .B(a[118]), .Z(n2778) );
  XOR U2897 ( .A(n2777), .B(n2778), .Z(n2780) );
  OR U2898 ( .A(n2743), .B(n2742), .Z(n2747) );
  NANDN U2899 ( .A(n2745), .B(n2744), .Z(n2746) );
  NAND U2900 ( .A(n2747), .B(n2746), .Z(n2779) );
  XNOR U2901 ( .A(n2780), .B(n2779), .Z(n2765) );
  NANDN U2902 ( .A(n2749), .B(n2748), .Z(n2753) );
  NAND U2903 ( .A(n2751), .B(n2750), .Z(n2752) );
  NAND U2904 ( .A(n2753), .B(n2752), .Z(n2766) );
  XNOR U2905 ( .A(n2765), .B(n2766), .Z(n2767) );
  NANDN U2906 ( .A(n2755), .B(n2754), .Z(n2759) );
  NANDN U2907 ( .A(n2757), .B(n2756), .Z(n2758) );
  NAND U2908 ( .A(n2759), .B(n2758), .Z(n2768) );
  XOR U2909 ( .A(n2767), .B(n2768), .Z(n2764) );
  XOR U2910 ( .A(sreg[242]), .B(n2763), .Z(n2762) );
  XNOR U2911 ( .A(n2764), .B(n2762), .Z(c[242]) );
  NANDN U2912 ( .A(n2766), .B(n2765), .Z(n2770) );
  NANDN U2913 ( .A(n2768), .B(n2767), .Z(n2769) );
  NAND U2914 ( .A(n2770), .B(n2769), .Z(n2798) );
  AND U2915 ( .A(b[2]), .B(a[117]), .Z(n2792) );
  AND U2916 ( .A(a[118]), .B(b[1]), .Z(n2790) );
  AND U2917 ( .A(a[116]), .B(b[3]), .Z(n2789) );
  XOR U2918 ( .A(n2790), .B(n2789), .Z(n2791) );
  XOR U2919 ( .A(n2792), .B(n2791), .Z(n2783) );
  NAND U2920 ( .A(b[0]), .B(a[119]), .Z(n2784) );
  XOR U2921 ( .A(n2783), .B(n2784), .Z(n2786) );
  OR U2922 ( .A(n2772), .B(n2771), .Z(n2776) );
  NANDN U2923 ( .A(n2774), .B(n2773), .Z(n2775) );
  NAND U2924 ( .A(n2776), .B(n2775), .Z(n2785) );
  XNOR U2925 ( .A(n2786), .B(n2785), .Z(n2795) );
  NANDN U2926 ( .A(n2778), .B(n2777), .Z(n2782) );
  OR U2927 ( .A(n2780), .B(n2779), .Z(n2781) );
  NAND U2928 ( .A(n2782), .B(n2781), .Z(n2796) );
  XNOR U2929 ( .A(n2795), .B(n2796), .Z(n2797) );
  XNOR U2930 ( .A(n2798), .B(n2797), .Z(n2801) );
  XNOR U2931 ( .A(n2801), .B(sreg[243]), .Z(n2802) );
  XOR U2932 ( .A(n2803), .B(n2802), .Z(c[243]) );
  NANDN U2933 ( .A(n2784), .B(n2783), .Z(n2788) );
  OR U2934 ( .A(n2786), .B(n2785), .Z(n2787) );
  NAND U2935 ( .A(n2788), .B(n2787), .Z(n2821) );
  AND U2936 ( .A(b[2]), .B(a[118]), .Z(n2812) );
  AND U2937 ( .A(a[119]), .B(b[1]), .Z(n2810) );
  AND U2938 ( .A(a[117]), .B(b[3]), .Z(n2809) );
  XOR U2939 ( .A(n2810), .B(n2809), .Z(n2811) );
  XOR U2940 ( .A(n2812), .B(n2811), .Z(n2815) );
  NAND U2941 ( .A(b[0]), .B(a[120]), .Z(n2816) );
  XNOR U2942 ( .A(n2815), .B(n2816), .Z(n2817) );
  OR U2943 ( .A(n2790), .B(n2789), .Z(n2794) );
  NANDN U2944 ( .A(n2792), .B(n2791), .Z(n2793) );
  AND U2945 ( .A(n2794), .B(n2793), .Z(n2818) );
  XNOR U2946 ( .A(n2817), .B(n2818), .Z(n2822) );
  XNOR U2947 ( .A(n2821), .B(n2822), .Z(n2823) );
  NANDN U2948 ( .A(n2796), .B(n2795), .Z(n2800) );
  NAND U2949 ( .A(n2798), .B(n2797), .Z(n2799) );
  NAND U2950 ( .A(n2800), .B(n2799), .Z(n2824) );
  XOR U2951 ( .A(n2823), .B(n2824), .Z(n2808) );
  NAND U2952 ( .A(n2801), .B(sreg[243]), .Z(n2805) );
  OR U2953 ( .A(n2803), .B(n2802), .Z(n2804) );
  AND U2954 ( .A(n2805), .B(n2804), .Z(n2807) );
  XNOR U2955 ( .A(n2807), .B(sreg[244]), .Z(n2806) );
  XNOR U2956 ( .A(n2808), .B(n2806), .Z(c[244]) );
  AND U2957 ( .A(b[2]), .B(a[119]), .Z(n2836) );
  AND U2958 ( .A(a[120]), .B(b[1]), .Z(n2834) );
  AND U2959 ( .A(a[118]), .B(b[3]), .Z(n2833) );
  XOR U2960 ( .A(n2834), .B(n2833), .Z(n2835) );
  XOR U2961 ( .A(n2836), .B(n2835), .Z(n2839) );
  NAND U2962 ( .A(b[0]), .B(a[121]), .Z(n2840) );
  XOR U2963 ( .A(n2839), .B(n2840), .Z(n2842) );
  OR U2964 ( .A(n2810), .B(n2809), .Z(n2814) );
  NANDN U2965 ( .A(n2812), .B(n2811), .Z(n2813) );
  NAND U2966 ( .A(n2814), .B(n2813), .Z(n2841) );
  XNOR U2967 ( .A(n2842), .B(n2841), .Z(n2827) );
  NANDN U2968 ( .A(n2816), .B(n2815), .Z(n2820) );
  NAND U2969 ( .A(n2818), .B(n2817), .Z(n2819) );
  NAND U2970 ( .A(n2820), .B(n2819), .Z(n2828) );
  XNOR U2971 ( .A(n2827), .B(n2828), .Z(n2829) );
  NANDN U2972 ( .A(n2822), .B(n2821), .Z(n2826) );
  NANDN U2973 ( .A(n2824), .B(n2823), .Z(n2825) );
  NAND U2974 ( .A(n2826), .B(n2825), .Z(n2830) );
  XOR U2975 ( .A(n2829), .B(n2830), .Z(n2845) );
  XNOR U2976 ( .A(n2845), .B(sreg[245]), .Z(n2847) );
  XNOR U2977 ( .A(n2846), .B(n2847), .Z(c[245]) );
  NANDN U2978 ( .A(n2828), .B(n2827), .Z(n2832) );
  NANDN U2979 ( .A(n2830), .B(n2829), .Z(n2831) );
  NAND U2980 ( .A(n2832), .B(n2831), .Z(n2853) );
  AND U2981 ( .A(b[2]), .B(a[120]), .Z(n2859) );
  AND U2982 ( .A(a[121]), .B(b[1]), .Z(n2857) );
  AND U2983 ( .A(a[119]), .B(b[3]), .Z(n2856) );
  XOR U2984 ( .A(n2857), .B(n2856), .Z(n2858) );
  XOR U2985 ( .A(n2859), .B(n2858), .Z(n2862) );
  NAND U2986 ( .A(b[0]), .B(a[122]), .Z(n2863) );
  XOR U2987 ( .A(n2862), .B(n2863), .Z(n2865) );
  OR U2988 ( .A(n2834), .B(n2833), .Z(n2838) );
  NANDN U2989 ( .A(n2836), .B(n2835), .Z(n2837) );
  NAND U2990 ( .A(n2838), .B(n2837), .Z(n2864) );
  XNOR U2991 ( .A(n2865), .B(n2864), .Z(n2850) );
  NANDN U2992 ( .A(n2840), .B(n2839), .Z(n2844) );
  OR U2993 ( .A(n2842), .B(n2841), .Z(n2843) );
  NAND U2994 ( .A(n2844), .B(n2843), .Z(n2851) );
  XNOR U2995 ( .A(n2850), .B(n2851), .Z(n2852) );
  XNOR U2996 ( .A(n2853), .B(n2852), .Z(n2868) );
  XOR U2997 ( .A(sreg[246]), .B(n2868), .Z(n2869) );
  NAND U2998 ( .A(n2845), .B(sreg[245]), .Z(n2849) );
  NANDN U2999 ( .A(n2847), .B(n2846), .Z(n2848) );
  NAND U3000 ( .A(n2849), .B(n2848), .Z(n2870) );
  XOR U3001 ( .A(n2869), .B(n2870), .Z(c[246]) );
  NANDN U3002 ( .A(n2851), .B(n2850), .Z(n2855) );
  NAND U3003 ( .A(n2853), .B(n2852), .Z(n2854) );
  NAND U3004 ( .A(n2855), .B(n2854), .Z(n2891) );
  AND U3005 ( .A(b[2]), .B(a[121]), .Z(n2885) );
  AND U3006 ( .A(a[122]), .B(b[1]), .Z(n2883) );
  AND U3007 ( .A(a[120]), .B(b[3]), .Z(n2882) );
  XOR U3008 ( .A(n2883), .B(n2882), .Z(n2884) );
  XOR U3009 ( .A(n2885), .B(n2884), .Z(n2876) );
  NAND U3010 ( .A(b[0]), .B(a[123]), .Z(n2877) );
  XOR U3011 ( .A(n2876), .B(n2877), .Z(n2879) );
  OR U3012 ( .A(n2857), .B(n2856), .Z(n2861) );
  NANDN U3013 ( .A(n2859), .B(n2858), .Z(n2860) );
  NAND U3014 ( .A(n2861), .B(n2860), .Z(n2878) );
  XNOR U3015 ( .A(n2879), .B(n2878), .Z(n2888) );
  NANDN U3016 ( .A(n2863), .B(n2862), .Z(n2867) );
  OR U3017 ( .A(n2865), .B(n2864), .Z(n2866) );
  NAND U3018 ( .A(n2867), .B(n2866), .Z(n2889) );
  XNOR U3019 ( .A(n2888), .B(n2889), .Z(n2890) );
  XOR U3020 ( .A(n2891), .B(n2890), .Z(n2875) );
  OR U3021 ( .A(n2868), .B(sreg[246]), .Z(n2872) );
  NANDN U3022 ( .A(n2870), .B(n2869), .Z(n2871) );
  AND U3023 ( .A(n2872), .B(n2871), .Z(n2874) );
  XNOR U3024 ( .A(sreg[247]), .B(n2874), .Z(n2873) );
  XOR U3025 ( .A(n2875), .B(n2873), .Z(c[247]) );
  NANDN U3026 ( .A(n2877), .B(n2876), .Z(n2881) );
  OR U3027 ( .A(n2879), .B(n2878), .Z(n2880) );
  NAND U3028 ( .A(n2881), .B(n2880), .Z(n2894) );
  AND U3029 ( .A(b[2]), .B(a[122]), .Z(n2903) );
  AND U3030 ( .A(a[123]), .B(b[1]), .Z(n2901) );
  AND U3031 ( .A(a[121]), .B(b[3]), .Z(n2900) );
  XOR U3032 ( .A(n2901), .B(n2900), .Z(n2902) );
  XOR U3033 ( .A(n2903), .B(n2902), .Z(n2906) );
  NAND U3034 ( .A(b[0]), .B(a[124]), .Z(n2907) );
  XNOR U3035 ( .A(n2906), .B(n2907), .Z(n2908) );
  OR U3036 ( .A(n2883), .B(n2882), .Z(n2887) );
  NANDN U3037 ( .A(n2885), .B(n2884), .Z(n2886) );
  AND U3038 ( .A(n2887), .B(n2886), .Z(n2909) );
  XNOR U3039 ( .A(n2908), .B(n2909), .Z(n2895) );
  XNOR U3040 ( .A(n2894), .B(n2895), .Z(n2896) );
  NANDN U3041 ( .A(n2889), .B(n2888), .Z(n2893) );
  NAND U3042 ( .A(n2891), .B(n2890), .Z(n2892) );
  AND U3043 ( .A(n2893), .B(n2892), .Z(n2897) );
  XOR U3044 ( .A(n2896), .B(n2897), .Z(n2912) );
  XNOR U3045 ( .A(sreg[248]), .B(n2912), .Z(n2913) );
  XOR U3046 ( .A(n2914), .B(n2913), .Z(c[248]) );
  NANDN U3047 ( .A(n2895), .B(n2894), .Z(n2899) );
  NAND U3048 ( .A(n2897), .B(n2896), .Z(n2898) );
  NAND U3049 ( .A(n2899), .B(n2898), .Z(n2923) );
  AND U3050 ( .A(b[2]), .B(a[123]), .Z(n2928) );
  AND U3051 ( .A(a[124]), .B(b[1]), .Z(n2966) );
  ANDN U3052 ( .B(a[122]), .A(n233), .Z(n2926) );
  XOR U3053 ( .A(n2966), .B(n2926), .Z(n2927) );
  XOR U3054 ( .A(n2928), .B(n2927), .Z(n2929) );
  NAND U3055 ( .A(a[125]), .B(b[0]), .Z(n2930) );
  XNOR U3056 ( .A(n2929), .B(n2930), .Z(n2931) );
  OR U3057 ( .A(n2901), .B(n2900), .Z(n2905) );
  NANDN U3058 ( .A(n2903), .B(n2902), .Z(n2904) );
  NAND U3059 ( .A(n2905), .B(n2904), .Z(n2932) );
  XOR U3060 ( .A(n2931), .B(n2932), .Z(n2920) );
  NANDN U3061 ( .A(n2907), .B(n2906), .Z(n2911) );
  NAND U3062 ( .A(n2909), .B(n2908), .Z(n2910) );
  NAND U3063 ( .A(n2911), .B(n2910), .Z(n2921) );
  XNOR U3064 ( .A(n2920), .B(n2921), .Z(n2922) );
  XOR U3065 ( .A(n2923), .B(n2922), .Z(n2919) );
  NAND U3066 ( .A(sreg[248]), .B(n2912), .Z(n2916) );
  OR U3067 ( .A(n2914), .B(n2913), .Z(n2915) );
  NAND U3068 ( .A(n2916), .B(n2915), .Z(n2918) );
  XNOR U3069 ( .A(sreg[249]), .B(n2918), .Z(n2917) );
  XNOR U3070 ( .A(n2919), .B(n2917), .Z(c[249]) );
  NANDN U3071 ( .A(n2921), .B(n2920), .Z(n2925) );
  NANDN U3072 ( .A(n2923), .B(n2922), .Z(n2924) );
  NAND U3073 ( .A(n2925), .B(n2924), .Z(n2943) );
  AND U3074 ( .A(b[2]), .B(a[124]), .Z(n2947) );
  NANDN U3075 ( .A(n233), .B(a[123]), .Z(n2945) );
  XNOR U3076 ( .A(n2946), .B(n2945), .Z(n2948) );
  XOR U3077 ( .A(n2947), .B(n2948), .Z(n2951) );
  NAND U3078 ( .A(b[0]), .B(a[126]), .Z(n2952) );
  XOR U3079 ( .A(n2951), .B(n2952), .Z(n2953) );
  XOR U3080 ( .A(n2953), .B(n2954), .Z(n2940) );
  NANDN U3081 ( .A(n2930), .B(n2929), .Z(n2934) );
  NANDN U3082 ( .A(n2932), .B(n2931), .Z(n2933) );
  AND U3083 ( .A(n2934), .B(n2933), .Z(n2941) );
  XOR U3084 ( .A(n2940), .B(n2941), .Z(n2942) );
  XOR U3085 ( .A(n2943), .B(n2942), .Z(n2935) );
  XNOR U3086 ( .A(n2935), .B(sreg[250]), .Z(n2936) );
  XOR U3087 ( .A(n2937), .B(n2936), .Z(c[250]) );
  NAND U3088 ( .A(n2935), .B(sreg[250]), .Z(n2939) );
  OR U3089 ( .A(n2937), .B(n2936), .Z(n2938) );
  NAND U3090 ( .A(n2939), .B(n2938), .Z(n2955) );
  XNOR U3091 ( .A(n2955), .B(sreg[251]), .Z(n2957) );
  AND U3092 ( .A(a[124]), .B(b[3]), .Z(n2944) );
  NAND U3093 ( .A(b[1]), .B(a[126]), .Z(n2987) );
  XOR U3094 ( .A(n2944), .B(n2987), .Z(n2968) );
  NAND U3095 ( .A(a[125]), .B(b[2]), .Z(n2967) );
  XOR U3096 ( .A(n2968), .B(n2967), .Z(n2971) );
  NAND U3097 ( .A(b[0]), .B(a[127]), .Z(n2972) );
  XOR U3098 ( .A(n2971), .B(n2972), .Z(n2973) );
  NAND U3099 ( .A(n2946), .B(n2945), .Z(n2950) );
  OR U3100 ( .A(n2948), .B(n2947), .Z(n2949) );
  AND U3101 ( .A(n2950), .B(n2949), .Z(n2974) );
  XNOR U3102 ( .A(n2973), .B(n2974), .Z(n2961) );
  XNOR U3103 ( .A(n2961), .B(n2960), .Z(n2963) );
  XOR U3104 ( .A(n2962), .B(n2963), .Z(n2956) );
  XOR U3105 ( .A(n2957), .B(n2956), .Z(c[251]) );
  NAND U3106 ( .A(n2955), .B(sreg[251]), .Z(n2959) );
  OR U3107 ( .A(n2957), .B(n2956), .Z(n2958) );
  AND U3108 ( .A(n2959), .B(n2958), .Z(n2976) );
  NANDN U3109 ( .A(n2961), .B(n2960), .Z(n2965) );
  NAND U3110 ( .A(n2963), .B(n2962), .Z(n2964) );
  NAND U3111 ( .A(n2965), .B(n2964), .Z(n2979) );
  AND U3112 ( .A(a[126]), .B(b[3]), .Z(n2997) );
  NAND U3113 ( .A(n2966), .B(n2997), .Z(n2970) );
  OR U3114 ( .A(n2968), .B(n2967), .Z(n2969) );
  NAND U3115 ( .A(n2970), .B(n2969), .Z(n2986) );
  NAND U3116 ( .A(b[1]), .B(a[127]), .Z(n2996) );
  AND U3117 ( .A(b[2]), .B(a[126]), .Z(n2995) );
  XNOR U3118 ( .A(n2996), .B(n2995), .Z(n2983) );
  NAND U3119 ( .A(a[125]), .B(b[3]), .Z(n2984) );
  XOR U3120 ( .A(n2983), .B(n2984), .Z(n2985) );
  XNOR U3121 ( .A(n2986), .B(n2985), .Z(n2978) );
  XNOR U3122 ( .A(n2978), .B(n2977), .Z(n2980) );
  XOR U3123 ( .A(n2979), .B(n2980), .Z(n2975) );
  XOR U3124 ( .A(n2976), .B(n2975), .Z(c[252]) );
  OR U3125 ( .A(n2976), .B(n2975), .Z(n3001) );
  NANDN U3126 ( .A(n2978), .B(n2977), .Z(n2982) );
  NAND U3127 ( .A(n2980), .B(n2979), .Z(n2981) );
  NAND U3128 ( .A(n2982), .B(n2981), .Z(n2992) );
  AND U3129 ( .A(n2987), .B(b[2]), .Z(n2988) );
  NAND U3130 ( .A(n2988), .B(a[127]), .Z(n2998) );
  XNOR U3131 ( .A(n2997), .B(n2998), .Z(n2990) );
  XOR U3132 ( .A(n2989), .B(n2990), .Z(n2991) );
  XOR U3133 ( .A(n2992), .B(n2991), .Z(n3002) );
  XOR U3134 ( .A(n3001), .B(n3002), .Z(c[253]) );
  NAND U3135 ( .A(n2990), .B(n2989), .Z(n2994) );
  NANDN U3136 ( .A(n2992), .B(n2991), .Z(n2993) );
  NAND U3137 ( .A(n2994), .B(n2993), .Z(n3009) );
  NAND U3138 ( .A(b[3]), .B(a[127]), .Z(n3006) );
  XOR U3139 ( .A(n3009), .B(n3006), .Z(n3004) );
  NANDN U3140 ( .A(n2996), .B(n2995), .Z(n3000) );
  NANDN U3141 ( .A(n2998), .B(n2997), .Z(n2999) );
  NAND U3142 ( .A(n3000), .B(n2999), .Z(n3007) );
  NOR U3143 ( .A(n3002), .B(n3001), .Z(n3008) );
  XOR U3144 ( .A(n3007), .B(n3008), .Z(n3003) );
  XNOR U3145 ( .A(n3004), .B(n3003), .Z(c[254]) );
  XNOR U3146 ( .A(n3008), .B(n3007), .Z(n3010) );
  XNOR U3147 ( .A(n3009), .B(n3010), .Z(n3005) );
  NANDN U3148 ( .A(n3006), .B(n3005), .Z(n3014) );
  OR U3149 ( .A(n3008), .B(n3007), .Z(n3012) );
  OR U3150 ( .A(n3010), .B(n3009), .Z(n3011) );
  NAND U3151 ( .A(n3012), .B(n3011), .Z(n3013) );
  NAND U3152 ( .A(n3014), .B(n3013), .Z(c[255]) );
endmodule

