
module modmult_step_N256_2_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279;

  IV U1 ( .A(n1278), .Z(n1) );
  IV U2 ( .A(A[1]), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(DIFF[9]) );
  XOR U4 ( .A(B[9]), .B(A[9]), .Z(n4) );
  XNOR U5 ( .A(n5), .B(n6), .Z(DIFF[99]) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(DIFF[98]) );
  XOR U8 ( .A(B[98]), .B(A[98]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(DIFF[97]) );
  XOR U10 ( .A(B[97]), .B(A[97]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(DIFF[96]) );
  XOR U12 ( .A(B[96]), .B(A[96]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(DIFF[95]) );
  XOR U14 ( .A(B[95]), .B(A[95]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(DIFF[94]) );
  XOR U16 ( .A(B[94]), .B(A[94]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(DIFF[93]) );
  XOR U18 ( .A(B[93]), .B(A[93]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(DIFF[92]) );
  XOR U20 ( .A(B[92]), .B(A[92]), .Z(n20) );
  XOR U21 ( .A(n21), .B(n22), .Z(DIFF[91]) );
  XOR U22 ( .A(B[91]), .B(A[91]), .Z(n22) );
  XOR U23 ( .A(n23), .B(n24), .Z(DIFF[90]) );
  XOR U24 ( .A(B[90]), .B(A[90]), .Z(n24) );
  XOR U25 ( .A(n25), .B(n26), .Z(DIFF[8]) );
  XOR U26 ( .A(B[8]), .B(A[8]), .Z(n26) );
  XOR U27 ( .A(n27), .B(n28), .Z(DIFF[89]) );
  XOR U28 ( .A(B[89]), .B(A[89]), .Z(n28) );
  XOR U29 ( .A(n29), .B(n30), .Z(DIFF[88]) );
  XOR U30 ( .A(B[88]), .B(A[88]), .Z(n30) );
  XOR U31 ( .A(n31), .B(n32), .Z(DIFF[87]) );
  XOR U32 ( .A(B[87]), .B(A[87]), .Z(n32) );
  XOR U33 ( .A(n33), .B(n34), .Z(DIFF[86]) );
  XOR U34 ( .A(B[86]), .B(A[86]), .Z(n34) );
  XOR U35 ( .A(n35), .B(n36), .Z(DIFF[85]) );
  XOR U36 ( .A(B[85]), .B(A[85]), .Z(n36) );
  XOR U37 ( .A(n37), .B(n38), .Z(DIFF[84]) );
  XOR U38 ( .A(B[84]), .B(A[84]), .Z(n38) );
  XOR U39 ( .A(n39), .B(n40), .Z(DIFF[83]) );
  XOR U40 ( .A(B[83]), .B(A[83]), .Z(n40) );
  XOR U41 ( .A(n41), .B(n42), .Z(DIFF[82]) );
  XOR U42 ( .A(B[82]), .B(A[82]), .Z(n42) );
  XOR U43 ( .A(n43), .B(n44), .Z(DIFF[81]) );
  XOR U44 ( .A(B[81]), .B(A[81]), .Z(n44) );
  XOR U45 ( .A(n45), .B(n46), .Z(DIFF[80]) );
  XOR U46 ( .A(B[80]), .B(A[80]), .Z(n46) );
  XOR U47 ( .A(n47), .B(n48), .Z(DIFF[7]) );
  XOR U48 ( .A(B[7]), .B(A[7]), .Z(n48) );
  XOR U49 ( .A(n49), .B(n50), .Z(DIFF[79]) );
  XOR U50 ( .A(B[79]), .B(A[79]), .Z(n50) );
  XOR U51 ( .A(n51), .B(n52), .Z(DIFF[78]) );
  XOR U52 ( .A(B[78]), .B(A[78]), .Z(n52) );
  XOR U53 ( .A(n53), .B(n54), .Z(DIFF[77]) );
  XOR U54 ( .A(B[77]), .B(A[77]), .Z(n54) );
  XOR U55 ( .A(n55), .B(n56), .Z(DIFF[76]) );
  XOR U56 ( .A(B[76]), .B(A[76]), .Z(n56) );
  XOR U57 ( .A(n57), .B(n58), .Z(DIFF[75]) );
  XOR U58 ( .A(B[75]), .B(A[75]), .Z(n58) );
  XOR U59 ( .A(n59), .B(n60), .Z(DIFF[74]) );
  XOR U60 ( .A(B[74]), .B(A[74]), .Z(n60) );
  XOR U61 ( .A(n61), .B(n62), .Z(DIFF[73]) );
  XOR U62 ( .A(B[73]), .B(A[73]), .Z(n62) );
  XOR U63 ( .A(n63), .B(n64), .Z(DIFF[72]) );
  XOR U64 ( .A(B[72]), .B(A[72]), .Z(n64) );
  XOR U65 ( .A(n65), .B(n66), .Z(DIFF[71]) );
  XOR U66 ( .A(B[71]), .B(A[71]), .Z(n66) );
  XOR U67 ( .A(n67), .B(n68), .Z(DIFF[70]) );
  XOR U68 ( .A(B[70]), .B(A[70]), .Z(n68) );
  XOR U69 ( .A(n69), .B(n70), .Z(DIFF[6]) );
  XOR U70 ( .A(B[6]), .B(A[6]), .Z(n70) );
  XOR U71 ( .A(n71), .B(n72), .Z(DIFF[69]) );
  XOR U72 ( .A(B[69]), .B(A[69]), .Z(n72) );
  XOR U73 ( .A(n73), .B(n74), .Z(DIFF[68]) );
  XOR U74 ( .A(B[68]), .B(A[68]), .Z(n74) );
  XOR U75 ( .A(n75), .B(n76), .Z(DIFF[67]) );
  XOR U76 ( .A(B[67]), .B(A[67]), .Z(n76) );
  XOR U77 ( .A(n77), .B(n78), .Z(DIFF[66]) );
  XOR U78 ( .A(B[66]), .B(A[66]), .Z(n78) );
  XOR U79 ( .A(n79), .B(n80), .Z(DIFF[65]) );
  XOR U80 ( .A(B[65]), .B(A[65]), .Z(n80) );
  XOR U81 ( .A(n81), .B(n82), .Z(DIFF[64]) );
  XOR U82 ( .A(B[64]), .B(A[64]), .Z(n82) );
  XOR U83 ( .A(n83), .B(n84), .Z(DIFF[63]) );
  XOR U84 ( .A(B[63]), .B(A[63]), .Z(n84) );
  XOR U85 ( .A(n85), .B(n86), .Z(DIFF[62]) );
  XOR U86 ( .A(B[62]), .B(A[62]), .Z(n86) );
  XOR U87 ( .A(n87), .B(n88), .Z(DIFF[61]) );
  XOR U88 ( .A(B[61]), .B(A[61]), .Z(n88) );
  XOR U89 ( .A(n89), .B(n90), .Z(DIFF[60]) );
  XOR U90 ( .A(B[60]), .B(A[60]), .Z(n90) );
  XOR U91 ( .A(n91), .B(n92), .Z(DIFF[5]) );
  XOR U92 ( .A(B[5]), .B(A[5]), .Z(n92) );
  XOR U93 ( .A(n93), .B(n94), .Z(DIFF[59]) );
  XOR U94 ( .A(B[59]), .B(A[59]), .Z(n94) );
  XOR U95 ( .A(n95), .B(n96), .Z(DIFF[58]) );
  XOR U96 ( .A(B[58]), .B(A[58]), .Z(n96) );
  XOR U97 ( .A(n97), .B(n98), .Z(DIFF[57]) );
  XOR U98 ( .A(B[57]), .B(A[57]), .Z(n98) );
  XOR U99 ( .A(n99), .B(n100), .Z(DIFF[56]) );
  XOR U100 ( .A(B[56]), .B(A[56]), .Z(n100) );
  XOR U101 ( .A(n101), .B(n102), .Z(DIFF[55]) );
  XOR U102 ( .A(B[55]), .B(A[55]), .Z(n102) );
  XOR U103 ( .A(n103), .B(n104), .Z(DIFF[54]) );
  XOR U104 ( .A(B[54]), .B(A[54]), .Z(n104) );
  XOR U105 ( .A(n105), .B(n106), .Z(DIFF[53]) );
  XOR U106 ( .A(B[53]), .B(A[53]), .Z(n106) );
  XOR U107 ( .A(n107), .B(n108), .Z(DIFF[52]) );
  XOR U108 ( .A(B[52]), .B(A[52]), .Z(n108) );
  XOR U109 ( .A(n109), .B(n110), .Z(DIFF[51]) );
  XOR U110 ( .A(B[51]), .B(A[51]), .Z(n110) );
  XOR U111 ( .A(n111), .B(n112), .Z(DIFF[50]) );
  XOR U112 ( .A(B[50]), .B(A[50]), .Z(n112) );
  XOR U113 ( .A(n113), .B(n114), .Z(DIFF[4]) );
  XOR U114 ( .A(B[4]), .B(A[4]), .Z(n114) );
  XOR U115 ( .A(n115), .B(n116), .Z(DIFF[49]) );
  XOR U116 ( .A(B[49]), .B(A[49]), .Z(n116) );
  XOR U117 ( .A(n117), .B(n118), .Z(DIFF[48]) );
  XOR U118 ( .A(B[48]), .B(A[48]), .Z(n118) );
  XOR U119 ( .A(n119), .B(n120), .Z(DIFF[47]) );
  XOR U120 ( .A(B[47]), .B(A[47]), .Z(n120) );
  XOR U121 ( .A(n121), .B(n122), .Z(DIFF[46]) );
  XOR U122 ( .A(B[46]), .B(A[46]), .Z(n122) );
  XOR U123 ( .A(n123), .B(n124), .Z(DIFF[45]) );
  XOR U124 ( .A(B[45]), .B(A[45]), .Z(n124) );
  XOR U125 ( .A(n125), .B(n126), .Z(DIFF[44]) );
  XOR U126 ( .A(B[44]), .B(A[44]), .Z(n126) );
  XOR U127 ( .A(n127), .B(n128), .Z(DIFF[43]) );
  XOR U128 ( .A(B[43]), .B(A[43]), .Z(n128) );
  XOR U129 ( .A(n129), .B(n130), .Z(DIFF[42]) );
  XOR U130 ( .A(B[42]), .B(A[42]), .Z(n130) );
  XOR U131 ( .A(n131), .B(n132), .Z(DIFF[41]) );
  XOR U132 ( .A(B[41]), .B(A[41]), .Z(n132) );
  XOR U133 ( .A(n133), .B(n134), .Z(DIFF[40]) );
  XOR U134 ( .A(B[40]), .B(A[40]), .Z(n134) );
  XOR U135 ( .A(n135), .B(n136), .Z(DIFF[3]) );
  XOR U136 ( .A(B[3]), .B(A[3]), .Z(n136) );
  XOR U137 ( .A(n137), .B(n138), .Z(DIFF[39]) );
  XOR U138 ( .A(B[39]), .B(A[39]), .Z(n138) );
  XOR U139 ( .A(n139), .B(n140), .Z(DIFF[38]) );
  XOR U140 ( .A(B[38]), .B(A[38]), .Z(n140) );
  XOR U141 ( .A(n141), .B(n142), .Z(DIFF[37]) );
  XOR U142 ( .A(B[37]), .B(A[37]), .Z(n142) );
  XOR U143 ( .A(n143), .B(n144), .Z(DIFF[36]) );
  XOR U144 ( .A(B[36]), .B(A[36]), .Z(n144) );
  XOR U145 ( .A(n145), .B(n146), .Z(DIFF[35]) );
  XOR U146 ( .A(B[35]), .B(A[35]), .Z(n146) );
  XOR U147 ( .A(n147), .B(n148), .Z(DIFF[34]) );
  XOR U148 ( .A(B[34]), .B(A[34]), .Z(n148) );
  XOR U149 ( .A(n149), .B(n150), .Z(DIFF[33]) );
  XOR U150 ( .A(B[33]), .B(A[33]), .Z(n150) );
  XOR U151 ( .A(n151), .B(n152), .Z(DIFF[32]) );
  XOR U152 ( .A(B[32]), .B(A[32]), .Z(n152) );
  XOR U153 ( .A(n153), .B(n154), .Z(DIFF[31]) );
  XOR U154 ( .A(B[31]), .B(A[31]), .Z(n154) );
  XOR U155 ( .A(n155), .B(n156), .Z(DIFF[30]) );
  XOR U156 ( .A(B[30]), .B(A[30]), .Z(n156) );
  XOR U157 ( .A(n157), .B(n158), .Z(DIFF[2]) );
  XOR U158 ( .A(B[2]), .B(A[2]), .Z(n158) );
  XOR U159 ( .A(n159), .B(n160), .Z(DIFF[29]) );
  XOR U160 ( .A(B[29]), .B(A[29]), .Z(n160) );
  XOR U161 ( .A(n161), .B(n162), .Z(DIFF[28]) );
  XOR U162 ( .A(B[28]), .B(A[28]), .Z(n162) );
  XOR U163 ( .A(n163), .B(n164), .Z(DIFF[27]) );
  XOR U164 ( .A(B[27]), .B(A[27]), .Z(n164) );
  XOR U165 ( .A(n165), .B(n166), .Z(DIFF[26]) );
  XOR U166 ( .A(B[26]), .B(A[26]), .Z(n166) );
  XOR U167 ( .A(n167), .B(n168), .Z(DIFF[25]) );
  XOR U168 ( .A(B[25]), .B(A[25]), .Z(n168) );
  XOR U169 ( .A(A[256]), .B(n169), .Z(DIFF[256]) );
  AND U170 ( .A(n170), .B(n171), .Z(n169) );
  NANDN U171 ( .A(B[255]), .B(n172), .Z(n171) );
  NANDN U172 ( .A(A[255]), .B(n173), .Z(n172) );
  NANDN U173 ( .A(n173), .B(A[255]), .Z(n170) );
  XOR U174 ( .A(n173), .B(n174), .Z(DIFF[255]) );
  XOR U175 ( .A(B[255]), .B(A[255]), .Z(n174) );
  AND U176 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U177 ( .A(B[254]), .B(n177), .Z(n176) );
  NANDN U178 ( .A(A[254]), .B(n178), .Z(n177) );
  NANDN U179 ( .A(n178), .B(A[254]), .Z(n175) );
  XOR U180 ( .A(n178), .B(n179), .Z(DIFF[254]) );
  XOR U181 ( .A(B[254]), .B(A[254]), .Z(n179) );
  AND U182 ( .A(n180), .B(n181), .Z(n178) );
  NANDN U183 ( .A(B[253]), .B(n182), .Z(n181) );
  NANDN U184 ( .A(A[253]), .B(n183), .Z(n182) );
  NANDN U185 ( .A(n183), .B(A[253]), .Z(n180) );
  XOR U186 ( .A(n183), .B(n184), .Z(DIFF[253]) );
  XOR U187 ( .A(B[253]), .B(A[253]), .Z(n184) );
  AND U188 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U189 ( .A(B[252]), .B(n187), .Z(n186) );
  NANDN U190 ( .A(A[252]), .B(n188), .Z(n187) );
  NANDN U191 ( .A(n188), .B(A[252]), .Z(n185) );
  XOR U192 ( .A(n188), .B(n189), .Z(DIFF[252]) );
  XOR U193 ( .A(B[252]), .B(A[252]), .Z(n189) );
  AND U194 ( .A(n190), .B(n191), .Z(n188) );
  NANDN U195 ( .A(B[251]), .B(n192), .Z(n191) );
  NANDN U196 ( .A(A[251]), .B(n193), .Z(n192) );
  NANDN U197 ( .A(n193), .B(A[251]), .Z(n190) );
  XOR U198 ( .A(n193), .B(n194), .Z(DIFF[251]) );
  XOR U199 ( .A(B[251]), .B(A[251]), .Z(n194) );
  AND U200 ( .A(n195), .B(n196), .Z(n193) );
  NANDN U201 ( .A(B[250]), .B(n197), .Z(n196) );
  NANDN U202 ( .A(A[250]), .B(n198), .Z(n197) );
  NANDN U203 ( .A(n198), .B(A[250]), .Z(n195) );
  XOR U204 ( .A(n198), .B(n199), .Z(DIFF[250]) );
  XOR U205 ( .A(B[250]), .B(A[250]), .Z(n199) );
  AND U206 ( .A(n200), .B(n201), .Z(n198) );
  NANDN U207 ( .A(B[249]), .B(n202), .Z(n201) );
  NANDN U208 ( .A(A[249]), .B(n203), .Z(n202) );
  NANDN U209 ( .A(n203), .B(A[249]), .Z(n200) );
  XOR U210 ( .A(n204), .B(n205), .Z(DIFF[24]) );
  XOR U211 ( .A(B[24]), .B(A[24]), .Z(n205) );
  XOR U212 ( .A(n203), .B(n206), .Z(DIFF[249]) );
  XOR U213 ( .A(B[249]), .B(A[249]), .Z(n206) );
  AND U214 ( .A(n207), .B(n208), .Z(n203) );
  NANDN U215 ( .A(B[248]), .B(n209), .Z(n208) );
  NANDN U216 ( .A(A[248]), .B(n210), .Z(n209) );
  NANDN U217 ( .A(n210), .B(A[248]), .Z(n207) );
  XOR U218 ( .A(n210), .B(n211), .Z(DIFF[248]) );
  XOR U219 ( .A(B[248]), .B(A[248]), .Z(n211) );
  AND U220 ( .A(n212), .B(n213), .Z(n210) );
  NANDN U221 ( .A(B[247]), .B(n214), .Z(n213) );
  NANDN U222 ( .A(A[247]), .B(n215), .Z(n214) );
  NANDN U223 ( .A(n215), .B(A[247]), .Z(n212) );
  XOR U224 ( .A(n215), .B(n216), .Z(DIFF[247]) );
  XOR U225 ( .A(B[247]), .B(A[247]), .Z(n216) );
  AND U226 ( .A(n217), .B(n218), .Z(n215) );
  NANDN U227 ( .A(B[246]), .B(n219), .Z(n218) );
  NANDN U228 ( .A(A[246]), .B(n220), .Z(n219) );
  NANDN U229 ( .A(n220), .B(A[246]), .Z(n217) );
  XOR U230 ( .A(n220), .B(n221), .Z(DIFF[246]) );
  XOR U231 ( .A(B[246]), .B(A[246]), .Z(n221) );
  AND U232 ( .A(n222), .B(n223), .Z(n220) );
  NANDN U233 ( .A(B[245]), .B(n224), .Z(n223) );
  NANDN U234 ( .A(A[245]), .B(n225), .Z(n224) );
  NANDN U235 ( .A(n225), .B(A[245]), .Z(n222) );
  XOR U236 ( .A(n225), .B(n226), .Z(DIFF[245]) );
  XOR U237 ( .A(B[245]), .B(A[245]), .Z(n226) );
  AND U238 ( .A(n227), .B(n228), .Z(n225) );
  NANDN U239 ( .A(B[244]), .B(n229), .Z(n228) );
  NANDN U240 ( .A(A[244]), .B(n230), .Z(n229) );
  NANDN U241 ( .A(n230), .B(A[244]), .Z(n227) );
  XOR U242 ( .A(n230), .B(n231), .Z(DIFF[244]) );
  XOR U243 ( .A(B[244]), .B(A[244]), .Z(n231) );
  AND U244 ( .A(n232), .B(n233), .Z(n230) );
  NANDN U245 ( .A(B[243]), .B(n234), .Z(n233) );
  NANDN U246 ( .A(A[243]), .B(n235), .Z(n234) );
  NANDN U247 ( .A(n235), .B(A[243]), .Z(n232) );
  XOR U248 ( .A(n235), .B(n236), .Z(DIFF[243]) );
  XOR U249 ( .A(B[243]), .B(A[243]), .Z(n236) );
  AND U250 ( .A(n237), .B(n238), .Z(n235) );
  NANDN U251 ( .A(B[242]), .B(n239), .Z(n238) );
  NANDN U252 ( .A(A[242]), .B(n240), .Z(n239) );
  NANDN U253 ( .A(n240), .B(A[242]), .Z(n237) );
  XOR U254 ( .A(n240), .B(n241), .Z(DIFF[242]) );
  XOR U255 ( .A(B[242]), .B(A[242]), .Z(n241) );
  AND U256 ( .A(n242), .B(n243), .Z(n240) );
  NANDN U257 ( .A(B[241]), .B(n244), .Z(n243) );
  NANDN U258 ( .A(A[241]), .B(n245), .Z(n244) );
  NANDN U259 ( .A(n245), .B(A[241]), .Z(n242) );
  XOR U260 ( .A(n245), .B(n246), .Z(DIFF[241]) );
  XOR U261 ( .A(B[241]), .B(A[241]), .Z(n246) );
  AND U262 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U263 ( .A(B[240]), .B(n249), .Z(n248) );
  NANDN U264 ( .A(A[240]), .B(n250), .Z(n249) );
  NANDN U265 ( .A(n250), .B(A[240]), .Z(n247) );
  XOR U266 ( .A(n250), .B(n251), .Z(DIFF[240]) );
  XOR U267 ( .A(B[240]), .B(A[240]), .Z(n251) );
  AND U268 ( .A(n252), .B(n253), .Z(n250) );
  NANDN U269 ( .A(B[239]), .B(n254), .Z(n253) );
  NANDN U270 ( .A(A[239]), .B(n255), .Z(n254) );
  NANDN U271 ( .A(n255), .B(A[239]), .Z(n252) );
  XOR U272 ( .A(n256), .B(n257), .Z(DIFF[23]) );
  XOR U273 ( .A(B[23]), .B(A[23]), .Z(n257) );
  XOR U274 ( .A(n255), .B(n258), .Z(DIFF[239]) );
  XOR U275 ( .A(B[239]), .B(A[239]), .Z(n258) );
  AND U276 ( .A(n259), .B(n260), .Z(n255) );
  NANDN U277 ( .A(B[238]), .B(n261), .Z(n260) );
  NANDN U278 ( .A(A[238]), .B(n262), .Z(n261) );
  NANDN U279 ( .A(n262), .B(A[238]), .Z(n259) );
  XOR U280 ( .A(n262), .B(n263), .Z(DIFF[238]) );
  XOR U281 ( .A(B[238]), .B(A[238]), .Z(n263) );
  AND U282 ( .A(n264), .B(n265), .Z(n262) );
  NANDN U283 ( .A(B[237]), .B(n266), .Z(n265) );
  NANDN U284 ( .A(A[237]), .B(n267), .Z(n266) );
  NANDN U285 ( .A(n267), .B(A[237]), .Z(n264) );
  XOR U286 ( .A(n267), .B(n268), .Z(DIFF[237]) );
  XOR U287 ( .A(B[237]), .B(A[237]), .Z(n268) );
  AND U288 ( .A(n269), .B(n270), .Z(n267) );
  NANDN U289 ( .A(B[236]), .B(n271), .Z(n270) );
  NANDN U290 ( .A(A[236]), .B(n272), .Z(n271) );
  NANDN U291 ( .A(n272), .B(A[236]), .Z(n269) );
  XOR U292 ( .A(n272), .B(n273), .Z(DIFF[236]) );
  XOR U293 ( .A(B[236]), .B(A[236]), .Z(n273) );
  AND U294 ( .A(n274), .B(n275), .Z(n272) );
  NANDN U295 ( .A(B[235]), .B(n276), .Z(n275) );
  NANDN U296 ( .A(A[235]), .B(n277), .Z(n276) );
  NANDN U297 ( .A(n277), .B(A[235]), .Z(n274) );
  XOR U298 ( .A(n277), .B(n278), .Z(DIFF[235]) );
  XOR U299 ( .A(B[235]), .B(A[235]), .Z(n278) );
  AND U300 ( .A(n279), .B(n280), .Z(n277) );
  NANDN U301 ( .A(B[234]), .B(n281), .Z(n280) );
  NANDN U302 ( .A(A[234]), .B(n282), .Z(n281) );
  NANDN U303 ( .A(n282), .B(A[234]), .Z(n279) );
  XOR U304 ( .A(n282), .B(n283), .Z(DIFF[234]) );
  XOR U305 ( .A(B[234]), .B(A[234]), .Z(n283) );
  AND U306 ( .A(n284), .B(n285), .Z(n282) );
  NANDN U307 ( .A(B[233]), .B(n286), .Z(n285) );
  NANDN U308 ( .A(A[233]), .B(n287), .Z(n286) );
  NANDN U309 ( .A(n287), .B(A[233]), .Z(n284) );
  XOR U310 ( .A(n287), .B(n288), .Z(DIFF[233]) );
  XOR U311 ( .A(B[233]), .B(A[233]), .Z(n288) );
  AND U312 ( .A(n289), .B(n290), .Z(n287) );
  NANDN U313 ( .A(B[232]), .B(n291), .Z(n290) );
  NANDN U314 ( .A(A[232]), .B(n292), .Z(n291) );
  NANDN U315 ( .A(n292), .B(A[232]), .Z(n289) );
  XOR U316 ( .A(n292), .B(n293), .Z(DIFF[232]) );
  XOR U317 ( .A(B[232]), .B(A[232]), .Z(n293) );
  AND U318 ( .A(n294), .B(n295), .Z(n292) );
  NANDN U319 ( .A(B[231]), .B(n296), .Z(n295) );
  NANDN U320 ( .A(A[231]), .B(n297), .Z(n296) );
  NANDN U321 ( .A(n297), .B(A[231]), .Z(n294) );
  XOR U322 ( .A(n297), .B(n298), .Z(DIFF[231]) );
  XOR U323 ( .A(B[231]), .B(A[231]), .Z(n298) );
  AND U324 ( .A(n299), .B(n300), .Z(n297) );
  NANDN U325 ( .A(B[230]), .B(n301), .Z(n300) );
  NANDN U326 ( .A(A[230]), .B(n302), .Z(n301) );
  NANDN U327 ( .A(n302), .B(A[230]), .Z(n299) );
  XOR U328 ( .A(n302), .B(n303), .Z(DIFF[230]) );
  XOR U329 ( .A(B[230]), .B(A[230]), .Z(n303) );
  AND U330 ( .A(n304), .B(n305), .Z(n302) );
  NANDN U331 ( .A(B[229]), .B(n306), .Z(n305) );
  NANDN U332 ( .A(A[229]), .B(n307), .Z(n306) );
  NANDN U333 ( .A(n307), .B(A[229]), .Z(n304) );
  XOR U334 ( .A(n308), .B(n309), .Z(DIFF[22]) );
  XOR U335 ( .A(B[22]), .B(A[22]), .Z(n309) );
  XOR U336 ( .A(n307), .B(n310), .Z(DIFF[229]) );
  XOR U337 ( .A(B[229]), .B(A[229]), .Z(n310) );
  AND U338 ( .A(n311), .B(n312), .Z(n307) );
  NANDN U339 ( .A(B[228]), .B(n313), .Z(n312) );
  NANDN U340 ( .A(A[228]), .B(n314), .Z(n313) );
  NANDN U341 ( .A(n314), .B(A[228]), .Z(n311) );
  XOR U342 ( .A(n314), .B(n315), .Z(DIFF[228]) );
  XOR U343 ( .A(B[228]), .B(A[228]), .Z(n315) );
  AND U344 ( .A(n316), .B(n317), .Z(n314) );
  NANDN U345 ( .A(B[227]), .B(n318), .Z(n317) );
  NANDN U346 ( .A(A[227]), .B(n319), .Z(n318) );
  NANDN U347 ( .A(n319), .B(A[227]), .Z(n316) );
  XOR U348 ( .A(n319), .B(n320), .Z(DIFF[227]) );
  XOR U349 ( .A(B[227]), .B(A[227]), .Z(n320) );
  AND U350 ( .A(n321), .B(n322), .Z(n319) );
  NANDN U351 ( .A(B[226]), .B(n323), .Z(n322) );
  NANDN U352 ( .A(A[226]), .B(n324), .Z(n323) );
  NANDN U353 ( .A(n324), .B(A[226]), .Z(n321) );
  XOR U354 ( .A(n324), .B(n325), .Z(DIFF[226]) );
  XOR U355 ( .A(B[226]), .B(A[226]), .Z(n325) );
  AND U356 ( .A(n326), .B(n327), .Z(n324) );
  NANDN U357 ( .A(B[225]), .B(n328), .Z(n327) );
  NANDN U358 ( .A(A[225]), .B(n329), .Z(n328) );
  NANDN U359 ( .A(n329), .B(A[225]), .Z(n326) );
  XOR U360 ( .A(n329), .B(n330), .Z(DIFF[225]) );
  XOR U361 ( .A(B[225]), .B(A[225]), .Z(n330) );
  AND U362 ( .A(n331), .B(n332), .Z(n329) );
  NANDN U363 ( .A(B[224]), .B(n333), .Z(n332) );
  NANDN U364 ( .A(A[224]), .B(n334), .Z(n333) );
  NANDN U365 ( .A(n334), .B(A[224]), .Z(n331) );
  XOR U366 ( .A(n334), .B(n335), .Z(DIFF[224]) );
  XOR U367 ( .A(B[224]), .B(A[224]), .Z(n335) );
  AND U368 ( .A(n336), .B(n337), .Z(n334) );
  NANDN U369 ( .A(B[223]), .B(n338), .Z(n337) );
  NANDN U370 ( .A(A[223]), .B(n339), .Z(n338) );
  NANDN U371 ( .A(n339), .B(A[223]), .Z(n336) );
  XOR U372 ( .A(n339), .B(n340), .Z(DIFF[223]) );
  XOR U373 ( .A(B[223]), .B(A[223]), .Z(n340) );
  AND U374 ( .A(n341), .B(n342), .Z(n339) );
  NANDN U375 ( .A(B[222]), .B(n343), .Z(n342) );
  NANDN U376 ( .A(A[222]), .B(n344), .Z(n343) );
  NANDN U377 ( .A(n344), .B(A[222]), .Z(n341) );
  XOR U378 ( .A(n344), .B(n345), .Z(DIFF[222]) );
  XOR U379 ( .A(B[222]), .B(A[222]), .Z(n345) );
  AND U380 ( .A(n346), .B(n347), .Z(n344) );
  NANDN U381 ( .A(B[221]), .B(n348), .Z(n347) );
  NANDN U382 ( .A(A[221]), .B(n349), .Z(n348) );
  NANDN U383 ( .A(n349), .B(A[221]), .Z(n346) );
  XOR U384 ( .A(n349), .B(n350), .Z(DIFF[221]) );
  XOR U385 ( .A(B[221]), .B(A[221]), .Z(n350) );
  AND U386 ( .A(n351), .B(n352), .Z(n349) );
  NANDN U387 ( .A(B[220]), .B(n353), .Z(n352) );
  NANDN U388 ( .A(A[220]), .B(n354), .Z(n353) );
  NANDN U389 ( .A(n354), .B(A[220]), .Z(n351) );
  XOR U390 ( .A(n354), .B(n355), .Z(DIFF[220]) );
  XOR U391 ( .A(B[220]), .B(A[220]), .Z(n355) );
  AND U392 ( .A(n356), .B(n357), .Z(n354) );
  NANDN U393 ( .A(B[219]), .B(n358), .Z(n357) );
  NANDN U394 ( .A(A[219]), .B(n359), .Z(n358) );
  NANDN U395 ( .A(n359), .B(A[219]), .Z(n356) );
  XOR U396 ( .A(n360), .B(n361), .Z(DIFF[21]) );
  XOR U397 ( .A(B[21]), .B(A[21]), .Z(n361) );
  XOR U398 ( .A(n359), .B(n362), .Z(DIFF[219]) );
  XOR U399 ( .A(B[219]), .B(A[219]), .Z(n362) );
  AND U400 ( .A(n363), .B(n364), .Z(n359) );
  NANDN U401 ( .A(B[218]), .B(n365), .Z(n364) );
  NANDN U402 ( .A(A[218]), .B(n366), .Z(n365) );
  NANDN U403 ( .A(n366), .B(A[218]), .Z(n363) );
  XOR U404 ( .A(n366), .B(n367), .Z(DIFF[218]) );
  XOR U405 ( .A(B[218]), .B(A[218]), .Z(n367) );
  AND U406 ( .A(n368), .B(n369), .Z(n366) );
  NANDN U407 ( .A(B[217]), .B(n370), .Z(n369) );
  NANDN U408 ( .A(A[217]), .B(n371), .Z(n370) );
  NANDN U409 ( .A(n371), .B(A[217]), .Z(n368) );
  XOR U410 ( .A(n371), .B(n372), .Z(DIFF[217]) );
  XOR U411 ( .A(B[217]), .B(A[217]), .Z(n372) );
  AND U412 ( .A(n373), .B(n374), .Z(n371) );
  NANDN U413 ( .A(B[216]), .B(n375), .Z(n374) );
  NANDN U414 ( .A(A[216]), .B(n376), .Z(n375) );
  NANDN U415 ( .A(n376), .B(A[216]), .Z(n373) );
  XOR U416 ( .A(n376), .B(n377), .Z(DIFF[216]) );
  XOR U417 ( .A(B[216]), .B(A[216]), .Z(n377) );
  AND U418 ( .A(n378), .B(n379), .Z(n376) );
  NANDN U419 ( .A(B[215]), .B(n380), .Z(n379) );
  NANDN U420 ( .A(A[215]), .B(n381), .Z(n380) );
  NANDN U421 ( .A(n381), .B(A[215]), .Z(n378) );
  XOR U422 ( .A(n381), .B(n382), .Z(DIFF[215]) );
  XOR U423 ( .A(B[215]), .B(A[215]), .Z(n382) );
  AND U424 ( .A(n383), .B(n384), .Z(n381) );
  NANDN U425 ( .A(B[214]), .B(n385), .Z(n384) );
  NANDN U426 ( .A(A[214]), .B(n386), .Z(n385) );
  NANDN U427 ( .A(n386), .B(A[214]), .Z(n383) );
  XOR U428 ( .A(n386), .B(n387), .Z(DIFF[214]) );
  XOR U429 ( .A(B[214]), .B(A[214]), .Z(n387) );
  AND U430 ( .A(n388), .B(n389), .Z(n386) );
  NANDN U431 ( .A(B[213]), .B(n390), .Z(n389) );
  NANDN U432 ( .A(A[213]), .B(n391), .Z(n390) );
  NANDN U433 ( .A(n391), .B(A[213]), .Z(n388) );
  XOR U434 ( .A(n391), .B(n392), .Z(DIFF[213]) );
  XOR U435 ( .A(B[213]), .B(A[213]), .Z(n392) );
  AND U436 ( .A(n393), .B(n394), .Z(n391) );
  NANDN U437 ( .A(B[212]), .B(n395), .Z(n394) );
  NANDN U438 ( .A(A[212]), .B(n396), .Z(n395) );
  NANDN U439 ( .A(n396), .B(A[212]), .Z(n393) );
  XOR U440 ( .A(n396), .B(n397), .Z(DIFF[212]) );
  XOR U441 ( .A(B[212]), .B(A[212]), .Z(n397) );
  AND U442 ( .A(n398), .B(n399), .Z(n396) );
  NANDN U443 ( .A(B[211]), .B(n400), .Z(n399) );
  NANDN U444 ( .A(A[211]), .B(n401), .Z(n400) );
  NANDN U445 ( .A(n401), .B(A[211]), .Z(n398) );
  XOR U446 ( .A(n401), .B(n402), .Z(DIFF[211]) );
  XOR U447 ( .A(B[211]), .B(A[211]), .Z(n402) );
  AND U448 ( .A(n403), .B(n404), .Z(n401) );
  NANDN U449 ( .A(B[210]), .B(n405), .Z(n404) );
  NANDN U450 ( .A(A[210]), .B(n406), .Z(n405) );
  NANDN U451 ( .A(n406), .B(A[210]), .Z(n403) );
  XOR U452 ( .A(n406), .B(n407), .Z(DIFF[210]) );
  XOR U453 ( .A(B[210]), .B(A[210]), .Z(n407) );
  AND U454 ( .A(n408), .B(n409), .Z(n406) );
  NANDN U455 ( .A(B[209]), .B(n410), .Z(n409) );
  NANDN U456 ( .A(A[209]), .B(n411), .Z(n410) );
  NANDN U457 ( .A(n411), .B(A[209]), .Z(n408) );
  XOR U458 ( .A(n412), .B(n413), .Z(DIFF[20]) );
  XOR U459 ( .A(B[20]), .B(A[20]), .Z(n413) );
  XOR U460 ( .A(n411), .B(n414), .Z(DIFF[209]) );
  XOR U461 ( .A(B[209]), .B(A[209]), .Z(n414) );
  AND U462 ( .A(n415), .B(n416), .Z(n411) );
  NANDN U463 ( .A(B[208]), .B(n417), .Z(n416) );
  NANDN U464 ( .A(A[208]), .B(n418), .Z(n417) );
  NANDN U465 ( .A(n418), .B(A[208]), .Z(n415) );
  XOR U466 ( .A(n418), .B(n419), .Z(DIFF[208]) );
  XOR U467 ( .A(B[208]), .B(A[208]), .Z(n419) );
  AND U468 ( .A(n420), .B(n421), .Z(n418) );
  NANDN U469 ( .A(B[207]), .B(n422), .Z(n421) );
  NANDN U470 ( .A(A[207]), .B(n423), .Z(n422) );
  NANDN U471 ( .A(n423), .B(A[207]), .Z(n420) );
  XOR U472 ( .A(n423), .B(n424), .Z(DIFF[207]) );
  XOR U473 ( .A(B[207]), .B(A[207]), .Z(n424) );
  AND U474 ( .A(n425), .B(n426), .Z(n423) );
  NANDN U475 ( .A(B[206]), .B(n427), .Z(n426) );
  NANDN U476 ( .A(A[206]), .B(n428), .Z(n427) );
  NANDN U477 ( .A(n428), .B(A[206]), .Z(n425) );
  XOR U478 ( .A(n428), .B(n429), .Z(DIFF[206]) );
  XOR U479 ( .A(B[206]), .B(A[206]), .Z(n429) );
  AND U480 ( .A(n430), .B(n431), .Z(n428) );
  NANDN U481 ( .A(B[205]), .B(n432), .Z(n431) );
  NANDN U482 ( .A(A[205]), .B(n433), .Z(n432) );
  NANDN U483 ( .A(n433), .B(A[205]), .Z(n430) );
  XOR U484 ( .A(n433), .B(n434), .Z(DIFF[205]) );
  XOR U485 ( .A(B[205]), .B(A[205]), .Z(n434) );
  AND U486 ( .A(n435), .B(n436), .Z(n433) );
  NANDN U487 ( .A(B[204]), .B(n437), .Z(n436) );
  NANDN U488 ( .A(A[204]), .B(n438), .Z(n437) );
  NANDN U489 ( .A(n438), .B(A[204]), .Z(n435) );
  XOR U490 ( .A(n438), .B(n439), .Z(DIFF[204]) );
  XOR U491 ( .A(B[204]), .B(A[204]), .Z(n439) );
  AND U492 ( .A(n440), .B(n441), .Z(n438) );
  NANDN U493 ( .A(B[203]), .B(n442), .Z(n441) );
  NANDN U494 ( .A(A[203]), .B(n443), .Z(n442) );
  NANDN U495 ( .A(n443), .B(A[203]), .Z(n440) );
  XOR U496 ( .A(n443), .B(n444), .Z(DIFF[203]) );
  XOR U497 ( .A(B[203]), .B(A[203]), .Z(n444) );
  AND U498 ( .A(n445), .B(n446), .Z(n443) );
  NANDN U499 ( .A(B[202]), .B(n447), .Z(n446) );
  NANDN U500 ( .A(A[202]), .B(n448), .Z(n447) );
  NANDN U501 ( .A(n448), .B(A[202]), .Z(n445) );
  XOR U502 ( .A(n448), .B(n449), .Z(DIFF[202]) );
  XOR U503 ( .A(B[202]), .B(A[202]), .Z(n449) );
  AND U504 ( .A(n450), .B(n451), .Z(n448) );
  NANDN U505 ( .A(B[201]), .B(n452), .Z(n451) );
  NANDN U506 ( .A(A[201]), .B(n453), .Z(n452) );
  NANDN U507 ( .A(n453), .B(A[201]), .Z(n450) );
  XOR U508 ( .A(n453), .B(n454), .Z(DIFF[201]) );
  XOR U509 ( .A(B[201]), .B(A[201]), .Z(n454) );
  AND U510 ( .A(n455), .B(n456), .Z(n453) );
  NANDN U511 ( .A(B[200]), .B(n457), .Z(n456) );
  NANDN U512 ( .A(A[200]), .B(n458), .Z(n457) );
  NANDN U513 ( .A(n458), .B(A[200]), .Z(n455) );
  XOR U514 ( .A(n458), .B(n459), .Z(DIFF[200]) );
  XOR U515 ( .A(B[200]), .B(A[200]), .Z(n459) );
  AND U516 ( .A(n460), .B(n461), .Z(n458) );
  NANDN U517 ( .A(B[199]), .B(n462), .Z(n461) );
  NANDN U518 ( .A(A[199]), .B(n463), .Z(n462) );
  NANDN U519 ( .A(n463), .B(A[199]), .Z(n460) );
  XOR U520 ( .A(n1), .B(n464), .Z(DIFF[1]) );
  XOR U521 ( .A(B[1]), .B(A[1]), .Z(n464) );
  XOR U522 ( .A(n465), .B(n466), .Z(DIFF[19]) );
  XOR U523 ( .A(B[19]), .B(A[19]), .Z(n466) );
  XOR U524 ( .A(n463), .B(n467), .Z(DIFF[199]) );
  XOR U525 ( .A(B[199]), .B(A[199]), .Z(n467) );
  AND U526 ( .A(n468), .B(n469), .Z(n463) );
  NANDN U527 ( .A(B[198]), .B(n470), .Z(n469) );
  NANDN U528 ( .A(A[198]), .B(n471), .Z(n470) );
  NANDN U529 ( .A(n471), .B(A[198]), .Z(n468) );
  XOR U530 ( .A(n471), .B(n472), .Z(DIFF[198]) );
  XOR U531 ( .A(B[198]), .B(A[198]), .Z(n472) );
  AND U532 ( .A(n473), .B(n474), .Z(n471) );
  NANDN U533 ( .A(B[197]), .B(n475), .Z(n474) );
  NANDN U534 ( .A(A[197]), .B(n476), .Z(n475) );
  NANDN U535 ( .A(n476), .B(A[197]), .Z(n473) );
  XOR U536 ( .A(n476), .B(n477), .Z(DIFF[197]) );
  XOR U537 ( .A(B[197]), .B(A[197]), .Z(n477) );
  AND U538 ( .A(n478), .B(n479), .Z(n476) );
  NANDN U539 ( .A(B[196]), .B(n480), .Z(n479) );
  NANDN U540 ( .A(A[196]), .B(n481), .Z(n480) );
  NANDN U541 ( .A(n481), .B(A[196]), .Z(n478) );
  XOR U542 ( .A(n481), .B(n482), .Z(DIFF[196]) );
  XOR U543 ( .A(B[196]), .B(A[196]), .Z(n482) );
  AND U544 ( .A(n483), .B(n484), .Z(n481) );
  NANDN U545 ( .A(B[195]), .B(n485), .Z(n484) );
  NANDN U546 ( .A(A[195]), .B(n486), .Z(n485) );
  NANDN U547 ( .A(n486), .B(A[195]), .Z(n483) );
  XOR U548 ( .A(n486), .B(n487), .Z(DIFF[195]) );
  XOR U549 ( .A(B[195]), .B(A[195]), .Z(n487) );
  AND U550 ( .A(n488), .B(n489), .Z(n486) );
  NANDN U551 ( .A(B[194]), .B(n490), .Z(n489) );
  NANDN U552 ( .A(A[194]), .B(n491), .Z(n490) );
  NANDN U553 ( .A(n491), .B(A[194]), .Z(n488) );
  XOR U554 ( .A(n491), .B(n492), .Z(DIFF[194]) );
  XOR U555 ( .A(B[194]), .B(A[194]), .Z(n492) );
  AND U556 ( .A(n493), .B(n494), .Z(n491) );
  NANDN U557 ( .A(B[193]), .B(n495), .Z(n494) );
  NANDN U558 ( .A(A[193]), .B(n496), .Z(n495) );
  NANDN U559 ( .A(n496), .B(A[193]), .Z(n493) );
  XOR U560 ( .A(n496), .B(n497), .Z(DIFF[193]) );
  XOR U561 ( .A(B[193]), .B(A[193]), .Z(n497) );
  AND U562 ( .A(n498), .B(n499), .Z(n496) );
  NANDN U563 ( .A(B[192]), .B(n500), .Z(n499) );
  NANDN U564 ( .A(A[192]), .B(n501), .Z(n500) );
  NANDN U565 ( .A(n501), .B(A[192]), .Z(n498) );
  XOR U566 ( .A(n501), .B(n502), .Z(DIFF[192]) );
  XOR U567 ( .A(B[192]), .B(A[192]), .Z(n502) );
  AND U568 ( .A(n503), .B(n504), .Z(n501) );
  NANDN U569 ( .A(B[191]), .B(n505), .Z(n504) );
  NANDN U570 ( .A(A[191]), .B(n506), .Z(n505) );
  NANDN U571 ( .A(n506), .B(A[191]), .Z(n503) );
  XOR U572 ( .A(n506), .B(n507), .Z(DIFF[191]) );
  XOR U573 ( .A(B[191]), .B(A[191]), .Z(n507) );
  AND U574 ( .A(n508), .B(n509), .Z(n506) );
  NANDN U575 ( .A(B[190]), .B(n510), .Z(n509) );
  NANDN U576 ( .A(A[190]), .B(n511), .Z(n510) );
  NANDN U577 ( .A(n511), .B(A[190]), .Z(n508) );
  XOR U578 ( .A(n511), .B(n512), .Z(DIFF[190]) );
  XOR U579 ( .A(B[190]), .B(A[190]), .Z(n512) );
  AND U580 ( .A(n513), .B(n514), .Z(n511) );
  NANDN U581 ( .A(B[189]), .B(n515), .Z(n514) );
  NANDN U582 ( .A(A[189]), .B(n516), .Z(n515) );
  NANDN U583 ( .A(n516), .B(A[189]), .Z(n513) );
  XOR U584 ( .A(n517), .B(n518), .Z(DIFF[18]) );
  XOR U585 ( .A(B[18]), .B(A[18]), .Z(n518) );
  XOR U586 ( .A(n516), .B(n519), .Z(DIFF[189]) );
  XOR U587 ( .A(B[189]), .B(A[189]), .Z(n519) );
  AND U588 ( .A(n520), .B(n521), .Z(n516) );
  NANDN U589 ( .A(B[188]), .B(n522), .Z(n521) );
  NANDN U590 ( .A(A[188]), .B(n523), .Z(n522) );
  NANDN U591 ( .A(n523), .B(A[188]), .Z(n520) );
  XOR U592 ( .A(n523), .B(n524), .Z(DIFF[188]) );
  XOR U593 ( .A(B[188]), .B(A[188]), .Z(n524) );
  AND U594 ( .A(n525), .B(n526), .Z(n523) );
  NANDN U595 ( .A(B[187]), .B(n527), .Z(n526) );
  NANDN U596 ( .A(A[187]), .B(n528), .Z(n527) );
  NANDN U597 ( .A(n528), .B(A[187]), .Z(n525) );
  XOR U598 ( .A(n528), .B(n529), .Z(DIFF[187]) );
  XOR U599 ( .A(B[187]), .B(A[187]), .Z(n529) );
  AND U600 ( .A(n530), .B(n531), .Z(n528) );
  NANDN U601 ( .A(B[186]), .B(n532), .Z(n531) );
  NANDN U602 ( .A(A[186]), .B(n533), .Z(n532) );
  NANDN U603 ( .A(n533), .B(A[186]), .Z(n530) );
  XOR U604 ( .A(n533), .B(n534), .Z(DIFF[186]) );
  XOR U605 ( .A(B[186]), .B(A[186]), .Z(n534) );
  AND U606 ( .A(n535), .B(n536), .Z(n533) );
  NANDN U607 ( .A(B[185]), .B(n537), .Z(n536) );
  NANDN U608 ( .A(A[185]), .B(n538), .Z(n537) );
  NANDN U609 ( .A(n538), .B(A[185]), .Z(n535) );
  XOR U610 ( .A(n538), .B(n539), .Z(DIFF[185]) );
  XOR U611 ( .A(B[185]), .B(A[185]), .Z(n539) );
  AND U612 ( .A(n540), .B(n541), .Z(n538) );
  NANDN U613 ( .A(B[184]), .B(n542), .Z(n541) );
  NANDN U614 ( .A(A[184]), .B(n543), .Z(n542) );
  NANDN U615 ( .A(n543), .B(A[184]), .Z(n540) );
  XOR U616 ( .A(n543), .B(n544), .Z(DIFF[184]) );
  XOR U617 ( .A(B[184]), .B(A[184]), .Z(n544) );
  AND U618 ( .A(n545), .B(n546), .Z(n543) );
  NANDN U619 ( .A(B[183]), .B(n547), .Z(n546) );
  NANDN U620 ( .A(A[183]), .B(n548), .Z(n547) );
  NANDN U621 ( .A(n548), .B(A[183]), .Z(n545) );
  XOR U622 ( .A(n548), .B(n549), .Z(DIFF[183]) );
  XOR U623 ( .A(B[183]), .B(A[183]), .Z(n549) );
  AND U624 ( .A(n550), .B(n551), .Z(n548) );
  NANDN U625 ( .A(B[182]), .B(n552), .Z(n551) );
  NANDN U626 ( .A(A[182]), .B(n553), .Z(n552) );
  NANDN U627 ( .A(n553), .B(A[182]), .Z(n550) );
  XOR U628 ( .A(n553), .B(n554), .Z(DIFF[182]) );
  XOR U629 ( .A(B[182]), .B(A[182]), .Z(n554) );
  AND U630 ( .A(n555), .B(n556), .Z(n553) );
  NANDN U631 ( .A(B[181]), .B(n557), .Z(n556) );
  NANDN U632 ( .A(A[181]), .B(n558), .Z(n557) );
  NANDN U633 ( .A(n558), .B(A[181]), .Z(n555) );
  XOR U634 ( .A(n558), .B(n559), .Z(DIFF[181]) );
  XOR U635 ( .A(B[181]), .B(A[181]), .Z(n559) );
  AND U636 ( .A(n560), .B(n561), .Z(n558) );
  NANDN U637 ( .A(B[180]), .B(n562), .Z(n561) );
  NANDN U638 ( .A(A[180]), .B(n563), .Z(n562) );
  NANDN U639 ( .A(n563), .B(A[180]), .Z(n560) );
  XOR U640 ( .A(n563), .B(n564), .Z(DIFF[180]) );
  XOR U641 ( .A(B[180]), .B(A[180]), .Z(n564) );
  AND U642 ( .A(n565), .B(n566), .Z(n563) );
  NANDN U643 ( .A(B[179]), .B(n567), .Z(n566) );
  NANDN U644 ( .A(A[179]), .B(n568), .Z(n567) );
  NANDN U645 ( .A(n568), .B(A[179]), .Z(n565) );
  XOR U646 ( .A(n569), .B(n570), .Z(DIFF[17]) );
  XOR U647 ( .A(B[17]), .B(A[17]), .Z(n570) );
  XOR U648 ( .A(n568), .B(n571), .Z(DIFF[179]) );
  XOR U649 ( .A(B[179]), .B(A[179]), .Z(n571) );
  AND U650 ( .A(n572), .B(n573), .Z(n568) );
  NANDN U651 ( .A(B[178]), .B(n574), .Z(n573) );
  NANDN U652 ( .A(A[178]), .B(n575), .Z(n574) );
  NANDN U653 ( .A(n575), .B(A[178]), .Z(n572) );
  XOR U654 ( .A(n575), .B(n576), .Z(DIFF[178]) );
  XOR U655 ( .A(B[178]), .B(A[178]), .Z(n576) );
  AND U656 ( .A(n577), .B(n578), .Z(n575) );
  NANDN U657 ( .A(B[177]), .B(n579), .Z(n578) );
  NANDN U658 ( .A(A[177]), .B(n580), .Z(n579) );
  NANDN U659 ( .A(n580), .B(A[177]), .Z(n577) );
  XOR U660 ( .A(n580), .B(n581), .Z(DIFF[177]) );
  XOR U661 ( .A(B[177]), .B(A[177]), .Z(n581) );
  AND U662 ( .A(n582), .B(n583), .Z(n580) );
  NANDN U663 ( .A(B[176]), .B(n584), .Z(n583) );
  NANDN U664 ( .A(A[176]), .B(n585), .Z(n584) );
  NANDN U665 ( .A(n585), .B(A[176]), .Z(n582) );
  XOR U666 ( .A(n585), .B(n586), .Z(DIFF[176]) );
  XOR U667 ( .A(B[176]), .B(A[176]), .Z(n586) );
  AND U668 ( .A(n587), .B(n588), .Z(n585) );
  NANDN U669 ( .A(B[175]), .B(n589), .Z(n588) );
  NANDN U670 ( .A(A[175]), .B(n590), .Z(n589) );
  NANDN U671 ( .A(n590), .B(A[175]), .Z(n587) );
  XOR U672 ( .A(n590), .B(n591), .Z(DIFF[175]) );
  XOR U673 ( .A(B[175]), .B(A[175]), .Z(n591) );
  AND U674 ( .A(n592), .B(n593), .Z(n590) );
  NANDN U675 ( .A(B[174]), .B(n594), .Z(n593) );
  NANDN U676 ( .A(A[174]), .B(n595), .Z(n594) );
  NANDN U677 ( .A(n595), .B(A[174]), .Z(n592) );
  XOR U678 ( .A(n595), .B(n596), .Z(DIFF[174]) );
  XOR U679 ( .A(B[174]), .B(A[174]), .Z(n596) );
  AND U680 ( .A(n597), .B(n598), .Z(n595) );
  NANDN U681 ( .A(B[173]), .B(n599), .Z(n598) );
  NANDN U682 ( .A(A[173]), .B(n600), .Z(n599) );
  NANDN U683 ( .A(n600), .B(A[173]), .Z(n597) );
  XOR U684 ( .A(n600), .B(n601), .Z(DIFF[173]) );
  XOR U685 ( .A(B[173]), .B(A[173]), .Z(n601) );
  AND U686 ( .A(n602), .B(n603), .Z(n600) );
  NANDN U687 ( .A(B[172]), .B(n604), .Z(n603) );
  NANDN U688 ( .A(A[172]), .B(n605), .Z(n604) );
  NANDN U689 ( .A(n605), .B(A[172]), .Z(n602) );
  XOR U690 ( .A(n605), .B(n606), .Z(DIFF[172]) );
  XOR U691 ( .A(B[172]), .B(A[172]), .Z(n606) );
  AND U692 ( .A(n607), .B(n608), .Z(n605) );
  NANDN U693 ( .A(B[171]), .B(n609), .Z(n608) );
  NANDN U694 ( .A(A[171]), .B(n610), .Z(n609) );
  NANDN U695 ( .A(n610), .B(A[171]), .Z(n607) );
  XOR U696 ( .A(n610), .B(n611), .Z(DIFF[171]) );
  XOR U697 ( .A(B[171]), .B(A[171]), .Z(n611) );
  AND U698 ( .A(n612), .B(n613), .Z(n610) );
  NANDN U699 ( .A(B[170]), .B(n614), .Z(n613) );
  NANDN U700 ( .A(A[170]), .B(n615), .Z(n614) );
  NANDN U701 ( .A(n615), .B(A[170]), .Z(n612) );
  XOR U702 ( .A(n615), .B(n616), .Z(DIFF[170]) );
  XOR U703 ( .A(B[170]), .B(A[170]), .Z(n616) );
  AND U704 ( .A(n617), .B(n618), .Z(n615) );
  NANDN U705 ( .A(B[169]), .B(n619), .Z(n618) );
  NANDN U706 ( .A(A[169]), .B(n620), .Z(n619) );
  NANDN U707 ( .A(n620), .B(A[169]), .Z(n617) );
  XOR U708 ( .A(n621), .B(n622), .Z(DIFF[16]) );
  XOR U709 ( .A(B[16]), .B(A[16]), .Z(n622) );
  XOR U710 ( .A(n620), .B(n623), .Z(DIFF[169]) );
  XOR U711 ( .A(B[169]), .B(A[169]), .Z(n623) );
  AND U712 ( .A(n624), .B(n625), .Z(n620) );
  NANDN U713 ( .A(B[168]), .B(n626), .Z(n625) );
  NANDN U714 ( .A(A[168]), .B(n627), .Z(n626) );
  NANDN U715 ( .A(n627), .B(A[168]), .Z(n624) );
  XOR U716 ( .A(n627), .B(n628), .Z(DIFF[168]) );
  XOR U717 ( .A(B[168]), .B(A[168]), .Z(n628) );
  AND U718 ( .A(n629), .B(n630), .Z(n627) );
  NANDN U719 ( .A(B[167]), .B(n631), .Z(n630) );
  NANDN U720 ( .A(A[167]), .B(n632), .Z(n631) );
  NANDN U721 ( .A(n632), .B(A[167]), .Z(n629) );
  XOR U722 ( .A(n632), .B(n633), .Z(DIFF[167]) );
  XOR U723 ( .A(B[167]), .B(A[167]), .Z(n633) );
  AND U724 ( .A(n634), .B(n635), .Z(n632) );
  NANDN U725 ( .A(B[166]), .B(n636), .Z(n635) );
  NANDN U726 ( .A(A[166]), .B(n637), .Z(n636) );
  NANDN U727 ( .A(n637), .B(A[166]), .Z(n634) );
  XOR U728 ( .A(n637), .B(n638), .Z(DIFF[166]) );
  XOR U729 ( .A(B[166]), .B(A[166]), .Z(n638) );
  AND U730 ( .A(n639), .B(n640), .Z(n637) );
  NANDN U731 ( .A(B[165]), .B(n641), .Z(n640) );
  NANDN U732 ( .A(A[165]), .B(n642), .Z(n641) );
  NANDN U733 ( .A(n642), .B(A[165]), .Z(n639) );
  XOR U734 ( .A(n642), .B(n643), .Z(DIFF[165]) );
  XOR U735 ( .A(B[165]), .B(A[165]), .Z(n643) );
  AND U736 ( .A(n644), .B(n645), .Z(n642) );
  NANDN U737 ( .A(B[164]), .B(n646), .Z(n645) );
  NANDN U738 ( .A(A[164]), .B(n647), .Z(n646) );
  NANDN U739 ( .A(n647), .B(A[164]), .Z(n644) );
  XOR U740 ( .A(n647), .B(n648), .Z(DIFF[164]) );
  XOR U741 ( .A(B[164]), .B(A[164]), .Z(n648) );
  AND U742 ( .A(n649), .B(n650), .Z(n647) );
  NANDN U743 ( .A(B[163]), .B(n651), .Z(n650) );
  NANDN U744 ( .A(A[163]), .B(n652), .Z(n651) );
  NANDN U745 ( .A(n652), .B(A[163]), .Z(n649) );
  XOR U746 ( .A(n652), .B(n653), .Z(DIFF[163]) );
  XOR U747 ( .A(B[163]), .B(A[163]), .Z(n653) );
  AND U748 ( .A(n654), .B(n655), .Z(n652) );
  NANDN U749 ( .A(B[162]), .B(n656), .Z(n655) );
  NANDN U750 ( .A(A[162]), .B(n657), .Z(n656) );
  NANDN U751 ( .A(n657), .B(A[162]), .Z(n654) );
  XOR U752 ( .A(n657), .B(n658), .Z(DIFF[162]) );
  XOR U753 ( .A(B[162]), .B(A[162]), .Z(n658) );
  AND U754 ( .A(n659), .B(n660), .Z(n657) );
  NANDN U755 ( .A(B[161]), .B(n661), .Z(n660) );
  NANDN U756 ( .A(A[161]), .B(n662), .Z(n661) );
  NANDN U757 ( .A(n662), .B(A[161]), .Z(n659) );
  XOR U758 ( .A(n662), .B(n663), .Z(DIFF[161]) );
  XOR U759 ( .A(B[161]), .B(A[161]), .Z(n663) );
  AND U760 ( .A(n664), .B(n665), .Z(n662) );
  NANDN U761 ( .A(B[160]), .B(n666), .Z(n665) );
  NANDN U762 ( .A(A[160]), .B(n667), .Z(n666) );
  NANDN U763 ( .A(n667), .B(A[160]), .Z(n664) );
  XOR U764 ( .A(n667), .B(n668), .Z(DIFF[160]) );
  XOR U765 ( .A(B[160]), .B(A[160]), .Z(n668) );
  AND U766 ( .A(n669), .B(n670), .Z(n667) );
  NANDN U767 ( .A(B[159]), .B(n671), .Z(n670) );
  NANDN U768 ( .A(A[159]), .B(n672), .Z(n671) );
  NANDN U769 ( .A(n672), .B(A[159]), .Z(n669) );
  XOR U770 ( .A(n673), .B(n674), .Z(DIFF[15]) );
  XOR U771 ( .A(B[15]), .B(A[15]), .Z(n674) );
  XOR U772 ( .A(n672), .B(n675), .Z(DIFF[159]) );
  XOR U773 ( .A(B[159]), .B(A[159]), .Z(n675) );
  AND U774 ( .A(n676), .B(n677), .Z(n672) );
  NANDN U775 ( .A(B[158]), .B(n678), .Z(n677) );
  NANDN U776 ( .A(A[158]), .B(n679), .Z(n678) );
  NANDN U777 ( .A(n679), .B(A[158]), .Z(n676) );
  XOR U778 ( .A(n679), .B(n680), .Z(DIFF[158]) );
  XOR U779 ( .A(B[158]), .B(A[158]), .Z(n680) );
  AND U780 ( .A(n681), .B(n682), .Z(n679) );
  NANDN U781 ( .A(B[157]), .B(n683), .Z(n682) );
  NANDN U782 ( .A(A[157]), .B(n684), .Z(n683) );
  NANDN U783 ( .A(n684), .B(A[157]), .Z(n681) );
  XOR U784 ( .A(n684), .B(n685), .Z(DIFF[157]) );
  XOR U785 ( .A(B[157]), .B(A[157]), .Z(n685) );
  AND U786 ( .A(n686), .B(n687), .Z(n684) );
  NANDN U787 ( .A(B[156]), .B(n688), .Z(n687) );
  NANDN U788 ( .A(A[156]), .B(n689), .Z(n688) );
  NANDN U789 ( .A(n689), .B(A[156]), .Z(n686) );
  XOR U790 ( .A(n689), .B(n690), .Z(DIFF[156]) );
  XOR U791 ( .A(B[156]), .B(A[156]), .Z(n690) );
  AND U792 ( .A(n691), .B(n692), .Z(n689) );
  NANDN U793 ( .A(B[155]), .B(n693), .Z(n692) );
  NANDN U794 ( .A(A[155]), .B(n694), .Z(n693) );
  NANDN U795 ( .A(n694), .B(A[155]), .Z(n691) );
  XOR U796 ( .A(n694), .B(n695), .Z(DIFF[155]) );
  XOR U797 ( .A(B[155]), .B(A[155]), .Z(n695) );
  AND U798 ( .A(n696), .B(n697), .Z(n694) );
  NANDN U799 ( .A(B[154]), .B(n698), .Z(n697) );
  NANDN U800 ( .A(A[154]), .B(n699), .Z(n698) );
  NANDN U801 ( .A(n699), .B(A[154]), .Z(n696) );
  XOR U802 ( .A(n699), .B(n700), .Z(DIFF[154]) );
  XOR U803 ( .A(B[154]), .B(A[154]), .Z(n700) );
  AND U804 ( .A(n701), .B(n702), .Z(n699) );
  NANDN U805 ( .A(B[153]), .B(n703), .Z(n702) );
  NANDN U806 ( .A(A[153]), .B(n704), .Z(n703) );
  NANDN U807 ( .A(n704), .B(A[153]), .Z(n701) );
  XOR U808 ( .A(n704), .B(n705), .Z(DIFF[153]) );
  XOR U809 ( .A(B[153]), .B(A[153]), .Z(n705) );
  AND U810 ( .A(n706), .B(n707), .Z(n704) );
  NANDN U811 ( .A(B[152]), .B(n708), .Z(n707) );
  NANDN U812 ( .A(A[152]), .B(n709), .Z(n708) );
  NANDN U813 ( .A(n709), .B(A[152]), .Z(n706) );
  XOR U814 ( .A(n709), .B(n710), .Z(DIFF[152]) );
  XOR U815 ( .A(B[152]), .B(A[152]), .Z(n710) );
  AND U816 ( .A(n711), .B(n712), .Z(n709) );
  NANDN U817 ( .A(B[151]), .B(n713), .Z(n712) );
  NANDN U818 ( .A(A[151]), .B(n714), .Z(n713) );
  NANDN U819 ( .A(n714), .B(A[151]), .Z(n711) );
  XOR U820 ( .A(n714), .B(n715), .Z(DIFF[151]) );
  XOR U821 ( .A(B[151]), .B(A[151]), .Z(n715) );
  AND U822 ( .A(n716), .B(n717), .Z(n714) );
  NANDN U823 ( .A(B[150]), .B(n718), .Z(n717) );
  NANDN U824 ( .A(A[150]), .B(n719), .Z(n718) );
  NANDN U825 ( .A(n719), .B(A[150]), .Z(n716) );
  XOR U826 ( .A(n719), .B(n720), .Z(DIFF[150]) );
  XOR U827 ( .A(B[150]), .B(A[150]), .Z(n720) );
  AND U828 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U829 ( .A(B[149]), .B(n723), .Z(n722) );
  NANDN U830 ( .A(A[149]), .B(n724), .Z(n723) );
  NANDN U831 ( .A(n724), .B(A[149]), .Z(n721) );
  XOR U832 ( .A(n725), .B(n726), .Z(DIFF[14]) );
  XOR U833 ( .A(B[14]), .B(A[14]), .Z(n726) );
  XOR U834 ( .A(n724), .B(n727), .Z(DIFF[149]) );
  XOR U835 ( .A(B[149]), .B(A[149]), .Z(n727) );
  AND U836 ( .A(n728), .B(n729), .Z(n724) );
  NANDN U837 ( .A(B[148]), .B(n730), .Z(n729) );
  NANDN U838 ( .A(A[148]), .B(n731), .Z(n730) );
  NANDN U839 ( .A(n731), .B(A[148]), .Z(n728) );
  XOR U840 ( .A(n731), .B(n732), .Z(DIFF[148]) );
  XOR U841 ( .A(B[148]), .B(A[148]), .Z(n732) );
  AND U842 ( .A(n733), .B(n734), .Z(n731) );
  NANDN U843 ( .A(B[147]), .B(n735), .Z(n734) );
  NANDN U844 ( .A(A[147]), .B(n736), .Z(n735) );
  NANDN U845 ( .A(n736), .B(A[147]), .Z(n733) );
  XOR U846 ( .A(n736), .B(n737), .Z(DIFF[147]) );
  XOR U847 ( .A(B[147]), .B(A[147]), .Z(n737) );
  AND U848 ( .A(n738), .B(n739), .Z(n736) );
  NANDN U849 ( .A(B[146]), .B(n740), .Z(n739) );
  NANDN U850 ( .A(A[146]), .B(n741), .Z(n740) );
  NANDN U851 ( .A(n741), .B(A[146]), .Z(n738) );
  XOR U852 ( .A(n741), .B(n742), .Z(DIFF[146]) );
  XOR U853 ( .A(B[146]), .B(A[146]), .Z(n742) );
  AND U854 ( .A(n743), .B(n744), .Z(n741) );
  NANDN U855 ( .A(B[145]), .B(n745), .Z(n744) );
  NANDN U856 ( .A(A[145]), .B(n746), .Z(n745) );
  NANDN U857 ( .A(n746), .B(A[145]), .Z(n743) );
  XOR U858 ( .A(n746), .B(n747), .Z(DIFF[145]) );
  XOR U859 ( .A(B[145]), .B(A[145]), .Z(n747) );
  AND U860 ( .A(n748), .B(n749), .Z(n746) );
  NANDN U861 ( .A(B[144]), .B(n750), .Z(n749) );
  NANDN U862 ( .A(A[144]), .B(n751), .Z(n750) );
  NANDN U863 ( .A(n751), .B(A[144]), .Z(n748) );
  XOR U864 ( .A(n751), .B(n752), .Z(DIFF[144]) );
  XOR U865 ( .A(B[144]), .B(A[144]), .Z(n752) );
  AND U866 ( .A(n753), .B(n754), .Z(n751) );
  NANDN U867 ( .A(B[143]), .B(n755), .Z(n754) );
  NANDN U868 ( .A(A[143]), .B(n756), .Z(n755) );
  NANDN U869 ( .A(n756), .B(A[143]), .Z(n753) );
  XOR U870 ( .A(n756), .B(n757), .Z(DIFF[143]) );
  XOR U871 ( .A(B[143]), .B(A[143]), .Z(n757) );
  AND U872 ( .A(n758), .B(n759), .Z(n756) );
  NANDN U873 ( .A(B[142]), .B(n760), .Z(n759) );
  NANDN U874 ( .A(A[142]), .B(n761), .Z(n760) );
  NANDN U875 ( .A(n761), .B(A[142]), .Z(n758) );
  XOR U876 ( .A(n761), .B(n762), .Z(DIFF[142]) );
  XOR U877 ( .A(B[142]), .B(A[142]), .Z(n762) );
  AND U878 ( .A(n763), .B(n764), .Z(n761) );
  NANDN U879 ( .A(B[141]), .B(n765), .Z(n764) );
  NANDN U880 ( .A(A[141]), .B(n766), .Z(n765) );
  NANDN U881 ( .A(n766), .B(A[141]), .Z(n763) );
  XOR U882 ( .A(n766), .B(n767), .Z(DIFF[141]) );
  XOR U883 ( .A(B[141]), .B(A[141]), .Z(n767) );
  AND U884 ( .A(n768), .B(n769), .Z(n766) );
  NANDN U885 ( .A(B[140]), .B(n770), .Z(n769) );
  NANDN U886 ( .A(A[140]), .B(n771), .Z(n770) );
  NANDN U887 ( .A(n771), .B(A[140]), .Z(n768) );
  XOR U888 ( .A(n771), .B(n772), .Z(DIFF[140]) );
  XOR U889 ( .A(B[140]), .B(A[140]), .Z(n772) );
  AND U890 ( .A(n773), .B(n774), .Z(n771) );
  NANDN U891 ( .A(B[139]), .B(n775), .Z(n774) );
  NANDN U892 ( .A(A[139]), .B(n776), .Z(n775) );
  NANDN U893 ( .A(n776), .B(A[139]), .Z(n773) );
  XOR U894 ( .A(n777), .B(n778), .Z(DIFF[13]) );
  XOR U895 ( .A(B[13]), .B(A[13]), .Z(n778) );
  XOR U896 ( .A(n776), .B(n779), .Z(DIFF[139]) );
  XOR U897 ( .A(B[139]), .B(A[139]), .Z(n779) );
  AND U898 ( .A(n780), .B(n781), .Z(n776) );
  NANDN U899 ( .A(B[138]), .B(n782), .Z(n781) );
  NANDN U900 ( .A(A[138]), .B(n783), .Z(n782) );
  NANDN U901 ( .A(n783), .B(A[138]), .Z(n780) );
  XOR U902 ( .A(n783), .B(n784), .Z(DIFF[138]) );
  XOR U903 ( .A(B[138]), .B(A[138]), .Z(n784) );
  AND U904 ( .A(n785), .B(n786), .Z(n783) );
  NANDN U905 ( .A(B[137]), .B(n787), .Z(n786) );
  NANDN U906 ( .A(A[137]), .B(n788), .Z(n787) );
  NANDN U907 ( .A(n788), .B(A[137]), .Z(n785) );
  XOR U908 ( .A(n788), .B(n789), .Z(DIFF[137]) );
  XOR U909 ( .A(B[137]), .B(A[137]), .Z(n789) );
  AND U910 ( .A(n790), .B(n791), .Z(n788) );
  NANDN U911 ( .A(B[136]), .B(n792), .Z(n791) );
  NANDN U912 ( .A(A[136]), .B(n793), .Z(n792) );
  NANDN U913 ( .A(n793), .B(A[136]), .Z(n790) );
  XOR U914 ( .A(n793), .B(n794), .Z(DIFF[136]) );
  XOR U915 ( .A(B[136]), .B(A[136]), .Z(n794) );
  AND U916 ( .A(n795), .B(n796), .Z(n793) );
  NANDN U917 ( .A(B[135]), .B(n797), .Z(n796) );
  NANDN U918 ( .A(A[135]), .B(n798), .Z(n797) );
  NANDN U919 ( .A(n798), .B(A[135]), .Z(n795) );
  XOR U920 ( .A(n798), .B(n799), .Z(DIFF[135]) );
  XOR U921 ( .A(B[135]), .B(A[135]), .Z(n799) );
  AND U922 ( .A(n800), .B(n801), .Z(n798) );
  NANDN U923 ( .A(B[134]), .B(n802), .Z(n801) );
  NANDN U924 ( .A(A[134]), .B(n803), .Z(n802) );
  NANDN U925 ( .A(n803), .B(A[134]), .Z(n800) );
  XOR U926 ( .A(n803), .B(n804), .Z(DIFF[134]) );
  XOR U927 ( .A(B[134]), .B(A[134]), .Z(n804) );
  AND U928 ( .A(n805), .B(n806), .Z(n803) );
  NANDN U929 ( .A(B[133]), .B(n807), .Z(n806) );
  NANDN U930 ( .A(A[133]), .B(n808), .Z(n807) );
  NANDN U931 ( .A(n808), .B(A[133]), .Z(n805) );
  XOR U932 ( .A(n808), .B(n809), .Z(DIFF[133]) );
  XOR U933 ( .A(B[133]), .B(A[133]), .Z(n809) );
  AND U934 ( .A(n810), .B(n811), .Z(n808) );
  NANDN U935 ( .A(B[132]), .B(n812), .Z(n811) );
  NANDN U936 ( .A(A[132]), .B(n813), .Z(n812) );
  NANDN U937 ( .A(n813), .B(A[132]), .Z(n810) );
  XOR U938 ( .A(n813), .B(n814), .Z(DIFF[132]) );
  XOR U939 ( .A(B[132]), .B(A[132]), .Z(n814) );
  AND U940 ( .A(n815), .B(n816), .Z(n813) );
  NANDN U941 ( .A(B[131]), .B(n817), .Z(n816) );
  NANDN U942 ( .A(A[131]), .B(n818), .Z(n817) );
  NANDN U943 ( .A(n818), .B(A[131]), .Z(n815) );
  XOR U944 ( .A(n818), .B(n819), .Z(DIFF[131]) );
  XOR U945 ( .A(B[131]), .B(A[131]), .Z(n819) );
  AND U946 ( .A(n820), .B(n821), .Z(n818) );
  NANDN U947 ( .A(B[130]), .B(n822), .Z(n821) );
  NANDN U948 ( .A(A[130]), .B(n823), .Z(n822) );
  NANDN U949 ( .A(n823), .B(A[130]), .Z(n820) );
  XOR U950 ( .A(n823), .B(n824), .Z(DIFF[130]) );
  XOR U951 ( .A(B[130]), .B(A[130]), .Z(n824) );
  AND U952 ( .A(n825), .B(n826), .Z(n823) );
  NANDN U953 ( .A(B[129]), .B(n827), .Z(n826) );
  NANDN U954 ( .A(A[129]), .B(n828), .Z(n827) );
  NANDN U955 ( .A(n828), .B(A[129]), .Z(n825) );
  XOR U956 ( .A(n829), .B(n830), .Z(DIFF[12]) );
  XOR U957 ( .A(B[12]), .B(A[12]), .Z(n830) );
  XOR U958 ( .A(n828), .B(n831), .Z(DIFF[129]) );
  XOR U959 ( .A(B[129]), .B(A[129]), .Z(n831) );
  AND U960 ( .A(n832), .B(n833), .Z(n828) );
  NANDN U961 ( .A(B[128]), .B(n834), .Z(n833) );
  NANDN U962 ( .A(A[128]), .B(n835), .Z(n834) );
  NANDN U963 ( .A(n835), .B(A[128]), .Z(n832) );
  XOR U964 ( .A(n835), .B(n836), .Z(DIFF[128]) );
  XOR U965 ( .A(B[128]), .B(A[128]), .Z(n836) );
  AND U966 ( .A(n837), .B(n838), .Z(n835) );
  NANDN U967 ( .A(B[127]), .B(n839), .Z(n838) );
  NANDN U968 ( .A(A[127]), .B(n840), .Z(n839) );
  NANDN U969 ( .A(n840), .B(A[127]), .Z(n837) );
  XOR U970 ( .A(n840), .B(n841), .Z(DIFF[127]) );
  XOR U971 ( .A(B[127]), .B(A[127]), .Z(n841) );
  AND U972 ( .A(n842), .B(n843), .Z(n840) );
  NANDN U973 ( .A(B[126]), .B(n844), .Z(n843) );
  NANDN U974 ( .A(A[126]), .B(n845), .Z(n844) );
  NANDN U975 ( .A(n845), .B(A[126]), .Z(n842) );
  XOR U976 ( .A(n845), .B(n846), .Z(DIFF[126]) );
  XOR U977 ( .A(B[126]), .B(A[126]), .Z(n846) );
  AND U978 ( .A(n847), .B(n848), .Z(n845) );
  NANDN U979 ( .A(B[125]), .B(n849), .Z(n848) );
  NANDN U980 ( .A(A[125]), .B(n850), .Z(n849) );
  NANDN U981 ( .A(n850), .B(A[125]), .Z(n847) );
  XOR U982 ( .A(n850), .B(n851), .Z(DIFF[125]) );
  XOR U983 ( .A(B[125]), .B(A[125]), .Z(n851) );
  AND U984 ( .A(n852), .B(n853), .Z(n850) );
  NANDN U985 ( .A(B[124]), .B(n854), .Z(n853) );
  NANDN U986 ( .A(A[124]), .B(n855), .Z(n854) );
  NANDN U987 ( .A(n855), .B(A[124]), .Z(n852) );
  XOR U988 ( .A(n855), .B(n856), .Z(DIFF[124]) );
  XOR U989 ( .A(B[124]), .B(A[124]), .Z(n856) );
  AND U990 ( .A(n857), .B(n858), .Z(n855) );
  NANDN U991 ( .A(B[123]), .B(n859), .Z(n858) );
  NANDN U992 ( .A(A[123]), .B(n860), .Z(n859) );
  NANDN U993 ( .A(n860), .B(A[123]), .Z(n857) );
  XOR U994 ( .A(n860), .B(n861), .Z(DIFF[123]) );
  XOR U995 ( .A(B[123]), .B(A[123]), .Z(n861) );
  AND U996 ( .A(n862), .B(n863), .Z(n860) );
  NANDN U997 ( .A(B[122]), .B(n864), .Z(n863) );
  NANDN U998 ( .A(A[122]), .B(n865), .Z(n864) );
  NANDN U999 ( .A(n865), .B(A[122]), .Z(n862) );
  XOR U1000 ( .A(n865), .B(n866), .Z(DIFF[122]) );
  XOR U1001 ( .A(B[122]), .B(A[122]), .Z(n866) );
  AND U1002 ( .A(n867), .B(n868), .Z(n865) );
  NANDN U1003 ( .A(B[121]), .B(n869), .Z(n868) );
  NANDN U1004 ( .A(A[121]), .B(n870), .Z(n869) );
  NANDN U1005 ( .A(n870), .B(A[121]), .Z(n867) );
  XOR U1006 ( .A(n870), .B(n871), .Z(DIFF[121]) );
  XOR U1007 ( .A(B[121]), .B(A[121]), .Z(n871) );
  AND U1008 ( .A(n872), .B(n873), .Z(n870) );
  NANDN U1009 ( .A(B[120]), .B(n874), .Z(n873) );
  NANDN U1010 ( .A(A[120]), .B(n875), .Z(n874) );
  NANDN U1011 ( .A(n875), .B(A[120]), .Z(n872) );
  XOR U1012 ( .A(n875), .B(n876), .Z(DIFF[120]) );
  XOR U1013 ( .A(B[120]), .B(A[120]), .Z(n876) );
  AND U1014 ( .A(n877), .B(n878), .Z(n875) );
  NANDN U1015 ( .A(B[119]), .B(n879), .Z(n878) );
  NANDN U1016 ( .A(A[119]), .B(n880), .Z(n879) );
  NANDN U1017 ( .A(n880), .B(A[119]), .Z(n877) );
  XOR U1018 ( .A(n881), .B(n882), .Z(DIFF[11]) );
  XOR U1019 ( .A(B[11]), .B(A[11]), .Z(n882) );
  XOR U1020 ( .A(n880), .B(n883), .Z(DIFF[119]) );
  XOR U1021 ( .A(B[119]), .B(A[119]), .Z(n883) );
  AND U1022 ( .A(n884), .B(n885), .Z(n880) );
  NANDN U1023 ( .A(B[118]), .B(n886), .Z(n885) );
  NANDN U1024 ( .A(A[118]), .B(n887), .Z(n886) );
  NANDN U1025 ( .A(n887), .B(A[118]), .Z(n884) );
  XOR U1026 ( .A(n887), .B(n888), .Z(DIFF[118]) );
  XOR U1027 ( .A(B[118]), .B(A[118]), .Z(n888) );
  AND U1028 ( .A(n889), .B(n890), .Z(n887) );
  NANDN U1029 ( .A(B[117]), .B(n891), .Z(n890) );
  NANDN U1030 ( .A(A[117]), .B(n892), .Z(n891) );
  NANDN U1031 ( .A(n892), .B(A[117]), .Z(n889) );
  XOR U1032 ( .A(n892), .B(n893), .Z(DIFF[117]) );
  XOR U1033 ( .A(B[117]), .B(A[117]), .Z(n893) );
  AND U1034 ( .A(n894), .B(n895), .Z(n892) );
  NANDN U1035 ( .A(B[116]), .B(n896), .Z(n895) );
  NANDN U1036 ( .A(A[116]), .B(n897), .Z(n896) );
  NANDN U1037 ( .A(n897), .B(A[116]), .Z(n894) );
  XOR U1038 ( .A(n897), .B(n898), .Z(DIFF[116]) );
  XOR U1039 ( .A(B[116]), .B(A[116]), .Z(n898) );
  AND U1040 ( .A(n899), .B(n900), .Z(n897) );
  NANDN U1041 ( .A(B[115]), .B(n901), .Z(n900) );
  NANDN U1042 ( .A(A[115]), .B(n902), .Z(n901) );
  NANDN U1043 ( .A(n902), .B(A[115]), .Z(n899) );
  XOR U1044 ( .A(n902), .B(n903), .Z(DIFF[115]) );
  XOR U1045 ( .A(B[115]), .B(A[115]), .Z(n903) );
  AND U1046 ( .A(n904), .B(n905), .Z(n902) );
  NANDN U1047 ( .A(B[114]), .B(n906), .Z(n905) );
  NANDN U1048 ( .A(A[114]), .B(n907), .Z(n906) );
  NANDN U1049 ( .A(n907), .B(A[114]), .Z(n904) );
  XOR U1050 ( .A(n907), .B(n908), .Z(DIFF[114]) );
  XOR U1051 ( .A(B[114]), .B(A[114]), .Z(n908) );
  AND U1052 ( .A(n909), .B(n910), .Z(n907) );
  NANDN U1053 ( .A(B[113]), .B(n911), .Z(n910) );
  NANDN U1054 ( .A(A[113]), .B(n912), .Z(n911) );
  NANDN U1055 ( .A(n912), .B(A[113]), .Z(n909) );
  XOR U1056 ( .A(n912), .B(n913), .Z(DIFF[113]) );
  XOR U1057 ( .A(B[113]), .B(A[113]), .Z(n913) );
  AND U1058 ( .A(n914), .B(n915), .Z(n912) );
  NANDN U1059 ( .A(B[112]), .B(n916), .Z(n915) );
  NANDN U1060 ( .A(A[112]), .B(n917), .Z(n916) );
  NANDN U1061 ( .A(n917), .B(A[112]), .Z(n914) );
  XOR U1062 ( .A(n917), .B(n918), .Z(DIFF[112]) );
  XOR U1063 ( .A(B[112]), .B(A[112]), .Z(n918) );
  AND U1064 ( .A(n919), .B(n920), .Z(n917) );
  NANDN U1065 ( .A(B[111]), .B(n921), .Z(n920) );
  NANDN U1066 ( .A(A[111]), .B(n922), .Z(n921) );
  NANDN U1067 ( .A(n922), .B(A[111]), .Z(n919) );
  XOR U1068 ( .A(n922), .B(n923), .Z(DIFF[111]) );
  XOR U1069 ( .A(B[111]), .B(A[111]), .Z(n923) );
  AND U1070 ( .A(n924), .B(n925), .Z(n922) );
  NANDN U1071 ( .A(B[110]), .B(n926), .Z(n925) );
  NANDN U1072 ( .A(A[110]), .B(n927), .Z(n926) );
  NANDN U1073 ( .A(n927), .B(A[110]), .Z(n924) );
  XOR U1074 ( .A(n927), .B(n928), .Z(DIFF[110]) );
  XOR U1075 ( .A(B[110]), .B(A[110]), .Z(n928) );
  AND U1076 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U1077 ( .A(B[109]), .B(n931), .Z(n930) );
  NANDN U1078 ( .A(A[109]), .B(n932), .Z(n931) );
  NANDN U1079 ( .A(n932), .B(A[109]), .Z(n929) );
  XOR U1080 ( .A(n933), .B(n934), .Z(DIFF[10]) );
  XOR U1081 ( .A(B[10]), .B(A[10]), .Z(n934) );
  XOR U1082 ( .A(n932), .B(n935), .Z(DIFF[109]) );
  XOR U1083 ( .A(B[109]), .B(A[109]), .Z(n935) );
  AND U1084 ( .A(n936), .B(n937), .Z(n932) );
  NANDN U1085 ( .A(B[108]), .B(n938), .Z(n937) );
  NANDN U1086 ( .A(A[108]), .B(n939), .Z(n938) );
  NANDN U1087 ( .A(n939), .B(A[108]), .Z(n936) );
  XOR U1088 ( .A(n939), .B(n940), .Z(DIFF[108]) );
  XOR U1089 ( .A(B[108]), .B(A[108]), .Z(n940) );
  AND U1090 ( .A(n941), .B(n942), .Z(n939) );
  NANDN U1091 ( .A(B[107]), .B(n943), .Z(n942) );
  NANDN U1092 ( .A(A[107]), .B(n944), .Z(n943) );
  NANDN U1093 ( .A(n944), .B(A[107]), .Z(n941) );
  XOR U1094 ( .A(n944), .B(n945), .Z(DIFF[107]) );
  XOR U1095 ( .A(B[107]), .B(A[107]), .Z(n945) );
  AND U1096 ( .A(n946), .B(n947), .Z(n944) );
  NANDN U1097 ( .A(B[106]), .B(n948), .Z(n947) );
  NANDN U1098 ( .A(A[106]), .B(n949), .Z(n948) );
  NANDN U1099 ( .A(n949), .B(A[106]), .Z(n946) );
  XOR U1100 ( .A(n949), .B(n950), .Z(DIFF[106]) );
  XOR U1101 ( .A(B[106]), .B(A[106]), .Z(n950) );
  AND U1102 ( .A(n951), .B(n952), .Z(n949) );
  NANDN U1103 ( .A(B[105]), .B(n953), .Z(n952) );
  NANDN U1104 ( .A(A[105]), .B(n954), .Z(n953) );
  NANDN U1105 ( .A(n954), .B(A[105]), .Z(n951) );
  XOR U1106 ( .A(n954), .B(n955), .Z(DIFF[105]) );
  XOR U1107 ( .A(B[105]), .B(A[105]), .Z(n955) );
  AND U1108 ( .A(n956), .B(n957), .Z(n954) );
  NANDN U1109 ( .A(B[104]), .B(n958), .Z(n957) );
  NANDN U1110 ( .A(A[104]), .B(n959), .Z(n958) );
  NANDN U1111 ( .A(n959), .B(A[104]), .Z(n956) );
  XOR U1112 ( .A(n959), .B(n960), .Z(DIFF[104]) );
  XOR U1113 ( .A(B[104]), .B(A[104]), .Z(n960) );
  AND U1114 ( .A(n961), .B(n962), .Z(n959) );
  NANDN U1115 ( .A(B[103]), .B(n963), .Z(n962) );
  NANDN U1116 ( .A(A[103]), .B(n964), .Z(n963) );
  NANDN U1117 ( .A(n964), .B(A[103]), .Z(n961) );
  XOR U1118 ( .A(n964), .B(n965), .Z(DIFF[103]) );
  XOR U1119 ( .A(B[103]), .B(A[103]), .Z(n965) );
  AND U1120 ( .A(n966), .B(n967), .Z(n964) );
  NANDN U1121 ( .A(B[102]), .B(n968), .Z(n967) );
  NANDN U1122 ( .A(A[102]), .B(n969), .Z(n968) );
  NANDN U1123 ( .A(n969), .B(A[102]), .Z(n966) );
  XOR U1124 ( .A(n969), .B(n970), .Z(DIFF[102]) );
  XOR U1125 ( .A(B[102]), .B(A[102]), .Z(n970) );
  AND U1126 ( .A(n971), .B(n972), .Z(n969) );
  NANDN U1127 ( .A(B[101]), .B(n973), .Z(n972) );
  NANDN U1128 ( .A(A[101]), .B(n974), .Z(n973) );
  NANDN U1129 ( .A(n974), .B(A[101]), .Z(n971) );
  XOR U1130 ( .A(n974), .B(n975), .Z(DIFF[101]) );
  XOR U1131 ( .A(B[101]), .B(A[101]), .Z(n975) );
  AND U1132 ( .A(n976), .B(n977), .Z(n974) );
  NANDN U1133 ( .A(B[100]), .B(n978), .Z(n977) );
  NANDN U1134 ( .A(A[100]), .B(n979), .Z(n978) );
  NANDN U1135 ( .A(n979), .B(A[100]), .Z(n976) );
  XOR U1136 ( .A(n979), .B(n980), .Z(DIFF[100]) );
  XOR U1137 ( .A(B[100]), .B(A[100]), .Z(n980) );
  AND U1138 ( .A(n981), .B(n982), .Z(n979) );
  NANDN U1139 ( .A(B[99]), .B(n983), .Z(n982) );
  OR U1140 ( .A(n5), .B(A[99]), .Z(n983) );
  NAND U1141 ( .A(A[99]), .B(n5), .Z(n981) );
  NAND U1142 ( .A(n984), .B(n985), .Z(n5) );
  NANDN U1143 ( .A(B[98]), .B(n986), .Z(n985) );
  NANDN U1144 ( .A(A[98]), .B(n7), .Z(n986) );
  NANDN U1145 ( .A(n7), .B(A[98]), .Z(n984) );
  AND U1146 ( .A(n987), .B(n988), .Z(n7) );
  NANDN U1147 ( .A(B[97]), .B(n989), .Z(n988) );
  NANDN U1148 ( .A(A[97]), .B(n9), .Z(n989) );
  NANDN U1149 ( .A(n9), .B(A[97]), .Z(n987) );
  AND U1150 ( .A(n990), .B(n991), .Z(n9) );
  NANDN U1151 ( .A(B[96]), .B(n992), .Z(n991) );
  NANDN U1152 ( .A(A[96]), .B(n11), .Z(n992) );
  NANDN U1153 ( .A(n11), .B(A[96]), .Z(n990) );
  AND U1154 ( .A(n993), .B(n994), .Z(n11) );
  NANDN U1155 ( .A(B[95]), .B(n995), .Z(n994) );
  NANDN U1156 ( .A(A[95]), .B(n13), .Z(n995) );
  NANDN U1157 ( .A(n13), .B(A[95]), .Z(n993) );
  AND U1158 ( .A(n996), .B(n997), .Z(n13) );
  NANDN U1159 ( .A(B[94]), .B(n998), .Z(n997) );
  NANDN U1160 ( .A(A[94]), .B(n15), .Z(n998) );
  NANDN U1161 ( .A(n15), .B(A[94]), .Z(n996) );
  AND U1162 ( .A(n999), .B(n1000), .Z(n15) );
  NANDN U1163 ( .A(B[93]), .B(n1001), .Z(n1000) );
  NANDN U1164 ( .A(A[93]), .B(n17), .Z(n1001) );
  NANDN U1165 ( .A(n17), .B(A[93]), .Z(n999) );
  AND U1166 ( .A(n1002), .B(n1003), .Z(n17) );
  NANDN U1167 ( .A(B[92]), .B(n1004), .Z(n1003) );
  NANDN U1168 ( .A(A[92]), .B(n19), .Z(n1004) );
  NANDN U1169 ( .A(n19), .B(A[92]), .Z(n1002) );
  AND U1170 ( .A(n1005), .B(n1006), .Z(n19) );
  NANDN U1171 ( .A(B[91]), .B(n1007), .Z(n1006) );
  NANDN U1172 ( .A(A[91]), .B(n21), .Z(n1007) );
  NANDN U1173 ( .A(n21), .B(A[91]), .Z(n1005) );
  AND U1174 ( .A(n1008), .B(n1009), .Z(n21) );
  NANDN U1175 ( .A(B[90]), .B(n1010), .Z(n1009) );
  NANDN U1176 ( .A(A[90]), .B(n23), .Z(n1010) );
  NANDN U1177 ( .A(n23), .B(A[90]), .Z(n1008) );
  AND U1178 ( .A(n1011), .B(n1012), .Z(n23) );
  NANDN U1179 ( .A(B[89]), .B(n1013), .Z(n1012) );
  NANDN U1180 ( .A(A[89]), .B(n27), .Z(n1013) );
  NANDN U1181 ( .A(n27), .B(A[89]), .Z(n1011) );
  AND U1182 ( .A(n1014), .B(n1015), .Z(n27) );
  NANDN U1183 ( .A(B[88]), .B(n1016), .Z(n1015) );
  NANDN U1184 ( .A(A[88]), .B(n29), .Z(n1016) );
  NANDN U1185 ( .A(n29), .B(A[88]), .Z(n1014) );
  AND U1186 ( .A(n1017), .B(n1018), .Z(n29) );
  NANDN U1187 ( .A(B[87]), .B(n1019), .Z(n1018) );
  NANDN U1188 ( .A(A[87]), .B(n31), .Z(n1019) );
  NANDN U1189 ( .A(n31), .B(A[87]), .Z(n1017) );
  AND U1190 ( .A(n1020), .B(n1021), .Z(n31) );
  NANDN U1191 ( .A(B[86]), .B(n1022), .Z(n1021) );
  NANDN U1192 ( .A(A[86]), .B(n33), .Z(n1022) );
  NANDN U1193 ( .A(n33), .B(A[86]), .Z(n1020) );
  AND U1194 ( .A(n1023), .B(n1024), .Z(n33) );
  NANDN U1195 ( .A(B[85]), .B(n1025), .Z(n1024) );
  NANDN U1196 ( .A(A[85]), .B(n35), .Z(n1025) );
  NANDN U1197 ( .A(n35), .B(A[85]), .Z(n1023) );
  AND U1198 ( .A(n1026), .B(n1027), .Z(n35) );
  NANDN U1199 ( .A(B[84]), .B(n1028), .Z(n1027) );
  NANDN U1200 ( .A(A[84]), .B(n37), .Z(n1028) );
  NANDN U1201 ( .A(n37), .B(A[84]), .Z(n1026) );
  AND U1202 ( .A(n1029), .B(n1030), .Z(n37) );
  NANDN U1203 ( .A(B[83]), .B(n1031), .Z(n1030) );
  NANDN U1204 ( .A(A[83]), .B(n39), .Z(n1031) );
  NANDN U1205 ( .A(n39), .B(A[83]), .Z(n1029) );
  AND U1206 ( .A(n1032), .B(n1033), .Z(n39) );
  NANDN U1207 ( .A(B[82]), .B(n1034), .Z(n1033) );
  NANDN U1208 ( .A(A[82]), .B(n41), .Z(n1034) );
  NANDN U1209 ( .A(n41), .B(A[82]), .Z(n1032) );
  AND U1210 ( .A(n1035), .B(n1036), .Z(n41) );
  NANDN U1211 ( .A(B[81]), .B(n1037), .Z(n1036) );
  NANDN U1212 ( .A(A[81]), .B(n43), .Z(n1037) );
  NANDN U1213 ( .A(n43), .B(A[81]), .Z(n1035) );
  AND U1214 ( .A(n1038), .B(n1039), .Z(n43) );
  NANDN U1215 ( .A(B[80]), .B(n1040), .Z(n1039) );
  NANDN U1216 ( .A(A[80]), .B(n45), .Z(n1040) );
  NANDN U1217 ( .A(n45), .B(A[80]), .Z(n1038) );
  AND U1218 ( .A(n1041), .B(n1042), .Z(n45) );
  NANDN U1219 ( .A(B[79]), .B(n1043), .Z(n1042) );
  NANDN U1220 ( .A(A[79]), .B(n49), .Z(n1043) );
  NANDN U1221 ( .A(n49), .B(A[79]), .Z(n1041) );
  AND U1222 ( .A(n1044), .B(n1045), .Z(n49) );
  NANDN U1223 ( .A(B[78]), .B(n1046), .Z(n1045) );
  NANDN U1224 ( .A(A[78]), .B(n51), .Z(n1046) );
  NANDN U1225 ( .A(n51), .B(A[78]), .Z(n1044) );
  AND U1226 ( .A(n1047), .B(n1048), .Z(n51) );
  NANDN U1227 ( .A(B[77]), .B(n1049), .Z(n1048) );
  NANDN U1228 ( .A(A[77]), .B(n53), .Z(n1049) );
  NANDN U1229 ( .A(n53), .B(A[77]), .Z(n1047) );
  AND U1230 ( .A(n1050), .B(n1051), .Z(n53) );
  NANDN U1231 ( .A(B[76]), .B(n1052), .Z(n1051) );
  NANDN U1232 ( .A(A[76]), .B(n55), .Z(n1052) );
  NANDN U1233 ( .A(n55), .B(A[76]), .Z(n1050) );
  AND U1234 ( .A(n1053), .B(n1054), .Z(n55) );
  NANDN U1235 ( .A(B[75]), .B(n1055), .Z(n1054) );
  NANDN U1236 ( .A(A[75]), .B(n57), .Z(n1055) );
  NANDN U1237 ( .A(n57), .B(A[75]), .Z(n1053) );
  AND U1238 ( .A(n1056), .B(n1057), .Z(n57) );
  NANDN U1239 ( .A(B[74]), .B(n1058), .Z(n1057) );
  NANDN U1240 ( .A(A[74]), .B(n59), .Z(n1058) );
  NANDN U1241 ( .A(n59), .B(A[74]), .Z(n1056) );
  AND U1242 ( .A(n1059), .B(n1060), .Z(n59) );
  NANDN U1243 ( .A(B[73]), .B(n1061), .Z(n1060) );
  NANDN U1244 ( .A(A[73]), .B(n61), .Z(n1061) );
  NANDN U1245 ( .A(n61), .B(A[73]), .Z(n1059) );
  AND U1246 ( .A(n1062), .B(n1063), .Z(n61) );
  NANDN U1247 ( .A(B[72]), .B(n1064), .Z(n1063) );
  NANDN U1248 ( .A(A[72]), .B(n63), .Z(n1064) );
  NANDN U1249 ( .A(n63), .B(A[72]), .Z(n1062) );
  AND U1250 ( .A(n1065), .B(n1066), .Z(n63) );
  NANDN U1251 ( .A(B[71]), .B(n1067), .Z(n1066) );
  NANDN U1252 ( .A(A[71]), .B(n65), .Z(n1067) );
  NANDN U1253 ( .A(n65), .B(A[71]), .Z(n1065) );
  AND U1254 ( .A(n1068), .B(n1069), .Z(n65) );
  NANDN U1255 ( .A(B[70]), .B(n1070), .Z(n1069) );
  NANDN U1256 ( .A(A[70]), .B(n67), .Z(n1070) );
  NANDN U1257 ( .A(n67), .B(A[70]), .Z(n1068) );
  AND U1258 ( .A(n1071), .B(n1072), .Z(n67) );
  NANDN U1259 ( .A(B[69]), .B(n1073), .Z(n1072) );
  NANDN U1260 ( .A(A[69]), .B(n71), .Z(n1073) );
  NANDN U1261 ( .A(n71), .B(A[69]), .Z(n1071) );
  AND U1262 ( .A(n1074), .B(n1075), .Z(n71) );
  NANDN U1263 ( .A(B[68]), .B(n1076), .Z(n1075) );
  NANDN U1264 ( .A(A[68]), .B(n73), .Z(n1076) );
  NANDN U1265 ( .A(n73), .B(A[68]), .Z(n1074) );
  AND U1266 ( .A(n1077), .B(n1078), .Z(n73) );
  NANDN U1267 ( .A(B[67]), .B(n1079), .Z(n1078) );
  NANDN U1268 ( .A(A[67]), .B(n75), .Z(n1079) );
  NANDN U1269 ( .A(n75), .B(A[67]), .Z(n1077) );
  AND U1270 ( .A(n1080), .B(n1081), .Z(n75) );
  NANDN U1271 ( .A(B[66]), .B(n1082), .Z(n1081) );
  NANDN U1272 ( .A(A[66]), .B(n77), .Z(n1082) );
  NANDN U1273 ( .A(n77), .B(A[66]), .Z(n1080) );
  AND U1274 ( .A(n1083), .B(n1084), .Z(n77) );
  NANDN U1275 ( .A(B[65]), .B(n1085), .Z(n1084) );
  NANDN U1276 ( .A(A[65]), .B(n79), .Z(n1085) );
  NANDN U1277 ( .A(n79), .B(A[65]), .Z(n1083) );
  AND U1278 ( .A(n1086), .B(n1087), .Z(n79) );
  NANDN U1279 ( .A(B[64]), .B(n1088), .Z(n1087) );
  NANDN U1280 ( .A(A[64]), .B(n81), .Z(n1088) );
  NANDN U1281 ( .A(n81), .B(A[64]), .Z(n1086) );
  AND U1282 ( .A(n1089), .B(n1090), .Z(n81) );
  NANDN U1283 ( .A(B[63]), .B(n1091), .Z(n1090) );
  NANDN U1284 ( .A(A[63]), .B(n83), .Z(n1091) );
  NANDN U1285 ( .A(n83), .B(A[63]), .Z(n1089) );
  AND U1286 ( .A(n1092), .B(n1093), .Z(n83) );
  NANDN U1287 ( .A(B[62]), .B(n1094), .Z(n1093) );
  NANDN U1288 ( .A(A[62]), .B(n85), .Z(n1094) );
  NANDN U1289 ( .A(n85), .B(A[62]), .Z(n1092) );
  AND U1290 ( .A(n1095), .B(n1096), .Z(n85) );
  NANDN U1291 ( .A(B[61]), .B(n1097), .Z(n1096) );
  NANDN U1292 ( .A(A[61]), .B(n87), .Z(n1097) );
  NANDN U1293 ( .A(n87), .B(A[61]), .Z(n1095) );
  AND U1294 ( .A(n1098), .B(n1099), .Z(n87) );
  NANDN U1295 ( .A(B[60]), .B(n1100), .Z(n1099) );
  NANDN U1296 ( .A(A[60]), .B(n89), .Z(n1100) );
  NANDN U1297 ( .A(n89), .B(A[60]), .Z(n1098) );
  AND U1298 ( .A(n1101), .B(n1102), .Z(n89) );
  NANDN U1299 ( .A(B[59]), .B(n1103), .Z(n1102) );
  NANDN U1300 ( .A(A[59]), .B(n93), .Z(n1103) );
  NANDN U1301 ( .A(n93), .B(A[59]), .Z(n1101) );
  AND U1302 ( .A(n1104), .B(n1105), .Z(n93) );
  NANDN U1303 ( .A(B[58]), .B(n1106), .Z(n1105) );
  NANDN U1304 ( .A(A[58]), .B(n95), .Z(n1106) );
  NANDN U1305 ( .A(n95), .B(A[58]), .Z(n1104) );
  AND U1306 ( .A(n1107), .B(n1108), .Z(n95) );
  NANDN U1307 ( .A(B[57]), .B(n1109), .Z(n1108) );
  NANDN U1308 ( .A(A[57]), .B(n97), .Z(n1109) );
  NANDN U1309 ( .A(n97), .B(A[57]), .Z(n1107) );
  AND U1310 ( .A(n1110), .B(n1111), .Z(n97) );
  NANDN U1311 ( .A(B[56]), .B(n1112), .Z(n1111) );
  NANDN U1312 ( .A(A[56]), .B(n99), .Z(n1112) );
  NANDN U1313 ( .A(n99), .B(A[56]), .Z(n1110) );
  AND U1314 ( .A(n1113), .B(n1114), .Z(n99) );
  NANDN U1315 ( .A(B[55]), .B(n1115), .Z(n1114) );
  NANDN U1316 ( .A(A[55]), .B(n101), .Z(n1115) );
  NANDN U1317 ( .A(n101), .B(A[55]), .Z(n1113) );
  AND U1318 ( .A(n1116), .B(n1117), .Z(n101) );
  NANDN U1319 ( .A(B[54]), .B(n1118), .Z(n1117) );
  NANDN U1320 ( .A(A[54]), .B(n103), .Z(n1118) );
  NANDN U1321 ( .A(n103), .B(A[54]), .Z(n1116) );
  AND U1322 ( .A(n1119), .B(n1120), .Z(n103) );
  NANDN U1323 ( .A(B[53]), .B(n1121), .Z(n1120) );
  NANDN U1324 ( .A(A[53]), .B(n105), .Z(n1121) );
  NANDN U1325 ( .A(n105), .B(A[53]), .Z(n1119) );
  AND U1326 ( .A(n1122), .B(n1123), .Z(n105) );
  NANDN U1327 ( .A(B[52]), .B(n1124), .Z(n1123) );
  NANDN U1328 ( .A(A[52]), .B(n107), .Z(n1124) );
  NANDN U1329 ( .A(n107), .B(A[52]), .Z(n1122) );
  AND U1330 ( .A(n1125), .B(n1126), .Z(n107) );
  NANDN U1331 ( .A(B[51]), .B(n1127), .Z(n1126) );
  NANDN U1332 ( .A(A[51]), .B(n109), .Z(n1127) );
  NANDN U1333 ( .A(n109), .B(A[51]), .Z(n1125) );
  AND U1334 ( .A(n1128), .B(n1129), .Z(n109) );
  NANDN U1335 ( .A(B[50]), .B(n1130), .Z(n1129) );
  NANDN U1336 ( .A(A[50]), .B(n111), .Z(n1130) );
  NANDN U1337 ( .A(n111), .B(A[50]), .Z(n1128) );
  AND U1338 ( .A(n1131), .B(n1132), .Z(n111) );
  NANDN U1339 ( .A(B[49]), .B(n1133), .Z(n1132) );
  NANDN U1340 ( .A(A[49]), .B(n115), .Z(n1133) );
  NANDN U1341 ( .A(n115), .B(A[49]), .Z(n1131) );
  AND U1342 ( .A(n1134), .B(n1135), .Z(n115) );
  NANDN U1343 ( .A(B[48]), .B(n1136), .Z(n1135) );
  NANDN U1344 ( .A(A[48]), .B(n117), .Z(n1136) );
  NANDN U1345 ( .A(n117), .B(A[48]), .Z(n1134) );
  AND U1346 ( .A(n1137), .B(n1138), .Z(n117) );
  NANDN U1347 ( .A(B[47]), .B(n1139), .Z(n1138) );
  NANDN U1348 ( .A(A[47]), .B(n119), .Z(n1139) );
  NANDN U1349 ( .A(n119), .B(A[47]), .Z(n1137) );
  AND U1350 ( .A(n1140), .B(n1141), .Z(n119) );
  NANDN U1351 ( .A(B[46]), .B(n1142), .Z(n1141) );
  NANDN U1352 ( .A(A[46]), .B(n121), .Z(n1142) );
  NANDN U1353 ( .A(n121), .B(A[46]), .Z(n1140) );
  AND U1354 ( .A(n1143), .B(n1144), .Z(n121) );
  NANDN U1355 ( .A(B[45]), .B(n1145), .Z(n1144) );
  NANDN U1356 ( .A(A[45]), .B(n123), .Z(n1145) );
  NANDN U1357 ( .A(n123), .B(A[45]), .Z(n1143) );
  AND U1358 ( .A(n1146), .B(n1147), .Z(n123) );
  NANDN U1359 ( .A(B[44]), .B(n1148), .Z(n1147) );
  NANDN U1360 ( .A(A[44]), .B(n125), .Z(n1148) );
  NANDN U1361 ( .A(n125), .B(A[44]), .Z(n1146) );
  AND U1362 ( .A(n1149), .B(n1150), .Z(n125) );
  NANDN U1363 ( .A(B[43]), .B(n1151), .Z(n1150) );
  NANDN U1364 ( .A(A[43]), .B(n127), .Z(n1151) );
  NANDN U1365 ( .A(n127), .B(A[43]), .Z(n1149) );
  AND U1366 ( .A(n1152), .B(n1153), .Z(n127) );
  NANDN U1367 ( .A(B[42]), .B(n1154), .Z(n1153) );
  NANDN U1368 ( .A(A[42]), .B(n129), .Z(n1154) );
  NANDN U1369 ( .A(n129), .B(A[42]), .Z(n1152) );
  AND U1370 ( .A(n1155), .B(n1156), .Z(n129) );
  NANDN U1371 ( .A(B[41]), .B(n1157), .Z(n1156) );
  NANDN U1372 ( .A(A[41]), .B(n131), .Z(n1157) );
  NANDN U1373 ( .A(n131), .B(A[41]), .Z(n1155) );
  AND U1374 ( .A(n1158), .B(n1159), .Z(n131) );
  NANDN U1375 ( .A(B[40]), .B(n1160), .Z(n1159) );
  NANDN U1376 ( .A(A[40]), .B(n133), .Z(n1160) );
  NANDN U1377 ( .A(n133), .B(A[40]), .Z(n1158) );
  AND U1378 ( .A(n1161), .B(n1162), .Z(n133) );
  NANDN U1379 ( .A(B[39]), .B(n1163), .Z(n1162) );
  NANDN U1380 ( .A(A[39]), .B(n137), .Z(n1163) );
  NANDN U1381 ( .A(n137), .B(A[39]), .Z(n1161) );
  AND U1382 ( .A(n1164), .B(n1165), .Z(n137) );
  NANDN U1383 ( .A(B[38]), .B(n1166), .Z(n1165) );
  NANDN U1384 ( .A(A[38]), .B(n139), .Z(n1166) );
  NANDN U1385 ( .A(n139), .B(A[38]), .Z(n1164) );
  AND U1386 ( .A(n1167), .B(n1168), .Z(n139) );
  NANDN U1387 ( .A(B[37]), .B(n1169), .Z(n1168) );
  NANDN U1388 ( .A(A[37]), .B(n141), .Z(n1169) );
  NANDN U1389 ( .A(n141), .B(A[37]), .Z(n1167) );
  AND U1390 ( .A(n1170), .B(n1171), .Z(n141) );
  NANDN U1391 ( .A(B[36]), .B(n1172), .Z(n1171) );
  NANDN U1392 ( .A(A[36]), .B(n143), .Z(n1172) );
  NANDN U1393 ( .A(n143), .B(A[36]), .Z(n1170) );
  AND U1394 ( .A(n1173), .B(n1174), .Z(n143) );
  NANDN U1395 ( .A(B[35]), .B(n1175), .Z(n1174) );
  NANDN U1396 ( .A(A[35]), .B(n145), .Z(n1175) );
  NANDN U1397 ( .A(n145), .B(A[35]), .Z(n1173) );
  AND U1398 ( .A(n1176), .B(n1177), .Z(n145) );
  NANDN U1399 ( .A(B[34]), .B(n1178), .Z(n1177) );
  NANDN U1400 ( .A(A[34]), .B(n147), .Z(n1178) );
  NANDN U1401 ( .A(n147), .B(A[34]), .Z(n1176) );
  AND U1402 ( .A(n1179), .B(n1180), .Z(n147) );
  NANDN U1403 ( .A(B[33]), .B(n1181), .Z(n1180) );
  NANDN U1404 ( .A(A[33]), .B(n149), .Z(n1181) );
  NANDN U1405 ( .A(n149), .B(A[33]), .Z(n1179) );
  AND U1406 ( .A(n1182), .B(n1183), .Z(n149) );
  NANDN U1407 ( .A(B[32]), .B(n1184), .Z(n1183) );
  NANDN U1408 ( .A(A[32]), .B(n151), .Z(n1184) );
  NANDN U1409 ( .A(n151), .B(A[32]), .Z(n1182) );
  AND U1410 ( .A(n1185), .B(n1186), .Z(n151) );
  NANDN U1411 ( .A(B[31]), .B(n1187), .Z(n1186) );
  NANDN U1412 ( .A(A[31]), .B(n153), .Z(n1187) );
  NANDN U1413 ( .A(n153), .B(A[31]), .Z(n1185) );
  AND U1414 ( .A(n1188), .B(n1189), .Z(n153) );
  NANDN U1415 ( .A(B[30]), .B(n1190), .Z(n1189) );
  NANDN U1416 ( .A(A[30]), .B(n155), .Z(n1190) );
  NANDN U1417 ( .A(n155), .B(A[30]), .Z(n1188) );
  AND U1418 ( .A(n1191), .B(n1192), .Z(n155) );
  NANDN U1419 ( .A(B[29]), .B(n1193), .Z(n1192) );
  NANDN U1420 ( .A(A[29]), .B(n159), .Z(n1193) );
  NANDN U1421 ( .A(n159), .B(A[29]), .Z(n1191) );
  AND U1422 ( .A(n1194), .B(n1195), .Z(n159) );
  NANDN U1423 ( .A(B[28]), .B(n1196), .Z(n1195) );
  NANDN U1424 ( .A(A[28]), .B(n161), .Z(n1196) );
  NANDN U1425 ( .A(n161), .B(A[28]), .Z(n1194) );
  AND U1426 ( .A(n1197), .B(n1198), .Z(n161) );
  NANDN U1427 ( .A(B[27]), .B(n1199), .Z(n1198) );
  NANDN U1428 ( .A(A[27]), .B(n163), .Z(n1199) );
  NANDN U1429 ( .A(n163), .B(A[27]), .Z(n1197) );
  AND U1430 ( .A(n1200), .B(n1201), .Z(n163) );
  NANDN U1431 ( .A(B[26]), .B(n1202), .Z(n1201) );
  NANDN U1432 ( .A(A[26]), .B(n165), .Z(n1202) );
  NANDN U1433 ( .A(n165), .B(A[26]), .Z(n1200) );
  AND U1434 ( .A(n1203), .B(n1204), .Z(n165) );
  NANDN U1435 ( .A(B[25]), .B(n1205), .Z(n1204) );
  NANDN U1436 ( .A(A[25]), .B(n167), .Z(n1205) );
  NANDN U1437 ( .A(n167), .B(A[25]), .Z(n1203) );
  AND U1438 ( .A(n1206), .B(n1207), .Z(n167) );
  NANDN U1439 ( .A(B[24]), .B(n1208), .Z(n1207) );
  NANDN U1440 ( .A(A[24]), .B(n204), .Z(n1208) );
  NANDN U1441 ( .A(n204), .B(A[24]), .Z(n1206) );
  AND U1442 ( .A(n1209), .B(n1210), .Z(n204) );
  NANDN U1443 ( .A(B[23]), .B(n1211), .Z(n1210) );
  NANDN U1444 ( .A(A[23]), .B(n256), .Z(n1211) );
  NANDN U1445 ( .A(n256), .B(A[23]), .Z(n1209) );
  AND U1446 ( .A(n1212), .B(n1213), .Z(n256) );
  NANDN U1447 ( .A(B[22]), .B(n1214), .Z(n1213) );
  NANDN U1448 ( .A(A[22]), .B(n308), .Z(n1214) );
  NANDN U1449 ( .A(n308), .B(A[22]), .Z(n1212) );
  AND U1450 ( .A(n1215), .B(n1216), .Z(n308) );
  NANDN U1451 ( .A(B[21]), .B(n1217), .Z(n1216) );
  NANDN U1452 ( .A(A[21]), .B(n360), .Z(n1217) );
  NANDN U1453 ( .A(n360), .B(A[21]), .Z(n1215) );
  AND U1454 ( .A(n1218), .B(n1219), .Z(n360) );
  NANDN U1455 ( .A(B[20]), .B(n1220), .Z(n1219) );
  NANDN U1456 ( .A(A[20]), .B(n412), .Z(n1220) );
  NANDN U1457 ( .A(n412), .B(A[20]), .Z(n1218) );
  AND U1458 ( .A(n1221), .B(n1222), .Z(n412) );
  NANDN U1459 ( .A(B[19]), .B(n1223), .Z(n1222) );
  NANDN U1460 ( .A(A[19]), .B(n465), .Z(n1223) );
  NANDN U1461 ( .A(n465), .B(A[19]), .Z(n1221) );
  AND U1462 ( .A(n1224), .B(n1225), .Z(n465) );
  NANDN U1463 ( .A(B[18]), .B(n1226), .Z(n1225) );
  NANDN U1464 ( .A(A[18]), .B(n517), .Z(n1226) );
  NANDN U1465 ( .A(n517), .B(A[18]), .Z(n1224) );
  AND U1466 ( .A(n1227), .B(n1228), .Z(n517) );
  NANDN U1467 ( .A(B[17]), .B(n1229), .Z(n1228) );
  NANDN U1468 ( .A(A[17]), .B(n569), .Z(n1229) );
  NANDN U1469 ( .A(n569), .B(A[17]), .Z(n1227) );
  AND U1470 ( .A(n1230), .B(n1231), .Z(n569) );
  NANDN U1471 ( .A(B[16]), .B(n1232), .Z(n1231) );
  NANDN U1472 ( .A(A[16]), .B(n621), .Z(n1232) );
  NANDN U1473 ( .A(n621), .B(A[16]), .Z(n1230) );
  AND U1474 ( .A(n1233), .B(n1234), .Z(n621) );
  NANDN U1475 ( .A(B[15]), .B(n1235), .Z(n1234) );
  NANDN U1476 ( .A(A[15]), .B(n673), .Z(n1235) );
  NANDN U1477 ( .A(n673), .B(A[15]), .Z(n1233) );
  AND U1478 ( .A(n1236), .B(n1237), .Z(n673) );
  NANDN U1479 ( .A(B[14]), .B(n1238), .Z(n1237) );
  NANDN U1480 ( .A(A[14]), .B(n725), .Z(n1238) );
  NANDN U1481 ( .A(n725), .B(A[14]), .Z(n1236) );
  AND U1482 ( .A(n1239), .B(n1240), .Z(n725) );
  NANDN U1483 ( .A(B[13]), .B(n1241), .Z(n1240) );
  NANDN U1484 ( .A(A[13]), .B(n777), .Z(n1241) );
  NANDN U1485 ( .A(n777), .B(A[13]), .Z(n1239) );
  AND U1486 ( .A(n1242), .B(n1243), .Z(n777) );
  NANDN U1487 ( .A(B[12]), .B(n1244), .Z(n1243) );
  NANDN U1488 ( .A(A[12]), .B(n829), .Z(n1244) );
  NANDN U1489 ( .A(n829), .B(A[12]), .Z(n1242) );
  AND U1490 ( .A(n1245), .B(n1246), .Z(n829) );
  NANDN U1491 ( .A(B[11]), .B(n1247), .Z(n1246) );
  NANDN U1492 ( .A(A[11]), .B(n881), .Z(n1247) );
  NANDN U1493 ( .A(n881), .B(A[11]), .Z(n1245) );
  AND U1494 ( .A(n1248), .B(n1249), .Z(n881) );
  NANDN U1495 ( .A(B[10]), .B(n1250), .Z(n1249) );
  NANDN U1496 ( .A(A[10]), .B(n933), .Z(n1250) );
  NANDN U1497 ( .A(n933), .B(A[10]), .Z(n1248) );
  AND U1498 ( .A(n1251), .B(n1252), .Z(n933) );
  NANDN U1499 ( .A(B[9]), .B(n1253), .Z(n1252) );
  OR U1500 ( .A(n3), .B(A[9]), .Z(n1253) );
  NAND U1501 ( .A(A[9]), .B(n3), .Z(n1251) );
  NAND U1502 ( .A(n1254), .B(n1255), .Z(n3) );
  NANDN U1503 ( .A(B[8]), .B(n1256), .Z(n1255) );
  NANDN U1504 ( .A(A[8]), .B(n25), .Z(n1256) );
  NANDN U1505 ( .A(n25), .B(A[8]), .Z(n1254) );
  AND U1506 ( .A(n1257), .B(n1258), .Z(n25) );
  NANDN U1507 ( .A(B[7]), .B(n1259), .Z(n1258) );
  NANDN U1508 ( .A(A[7]), .B(n47), .Z(n1259) );
  NANDN U1509 ( .A(n47), .B(A[7]), .Z(n1257) );
  AND U1510 ( .A(n1260), .B(n1261), .Z(n47) );
  NANDN U1511 ( .A(B[6]), .B(n1262), .Z(n1261) );
  NANDN U1512 ( .A(A[6]), .B(n69), .Z(n1262) );
  NANDN U1513 ( .A(n69), .B(A[6]), .Z(n1260) );
  AND U1514 ( .A(n1263), .B(n1264), .Z(n69) );
  NANDN U1515 ( .A(B[5]), .B(n1265), .Z(n1264) );
  NANDN U1516 ( .A(A[5]), .B(n91), .Z(n1265) );
  NANDN U1517 ( .A(n91), .B(A[5]), .Z(n1263) );
  AND U1518 ( .A(n1266), .B(n1267), .Z(n91) );
  NANDN U1519 ( .A(B[4]), .B(n1268), .Z(n1267) );
  NANDN U1520 ( .A(A[4]), .B(n113), .Z(n1268) );
  NANDN U1521 ( .A(n113), .B(A[4]), .Z(n1266) );
  AND U1522 ( .A(n1269), .B(n1270), .Z(n113) );
  NANDN U1523 ( .A(B[3]), .B(n1271), .Z(n1270) );
  NANDN U1524 ( .A(A[3]), .B(n135), .Z(n1271) );
  NANDN U1525 ( .A(n135), .B(A[3]), .Z(n1269) );
  AND U1526 ( .A(n1272), .B(n1273), .Z(n135) );
  NANDN U1527 ( .A(B[2]), .B(n1274), .Z(n1273) );
  NANDN U1528 ( .A(A[2]), .B(n157), .Z(n1274) );
  NANDN U1529 ( .A(n157), .B(A[2]), .Z(n1272) );
  AND U1530 ( .A(n1275), .B(n1276), .Z(n157) );
  NANDN U1531 ( .A(B[1]), .B(n1277), .Z(n1276) );
  NAND U1532 ( .A(n1), .B(n2), .Z(n1277) );
  NAND U1533 ( .A(A[1]), .B(n1278), .Z(n1275) );
  NAND U1534 ( .A(n1278), .B(n1279), .Z(DIFF[0]) );
  NANDN U1535 ( .A(B[0]), .B(A[0]), .Z(n1279) );
  NANDN U1536 ( .A(A[0]), .B(B[0]), .Z(n1278) );
endmodule


module modmult_step_N256_2_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [255:0] A;
  input [0:0] B;
  output [256:0] PRODUCT;
  input TC;


  AND U2 ( .A(A[255]), .B(B[0]), .Z(PRODUCT[255]) );
  AND U3 ( .A(A[254]), .B(B[0]), .Z(PRODUCT[254]) );
  AND U4 ( .A(A[253]), .B(B[0]), .Z(PRODUCT[253]) );
  AND U5 ( .A(A[252]), .B(B[0]), .Z(PRODUCT[252]) );
  AND U6 ( .A(A[251]), .B(B[0]), .Z(PRODUCT[251]) );
  AND U7 ( .A(A[250]), .B(B[0]), .Z(PRODUCT[250]) );
  AND U8 ( .A(A[249]), .B(B[0]), .Z(PRODUCT[249]) );
  AND U9 ( .A(A[248]), .B(B[0]), .Z(PRODUCT[248]) );
  AND U10 ( .A(A[247]), .B(B[0]), .Z(PRODUCT[247]) );
  AND U11 ( .A(A[246]), .B(B[0]), .Z(PRODUCT[246]) );
  AND U12 ( .A(A[245]), .B(B[0]), .Z(PRODUCT[245]) );
  AND U13 ( .A(A[244]), .B(B[0]), .Z(PRODUCT[244]) );
  AND U14 ( .A(A[243]), .B(B[0]), .Z(PRODUCT[243]) );
  AND U15 ( .A(A[242]), .B(B[0]), .Z(PRODUCT[242]) );
  AND U16 ( .A(A[241]), .B(B[0]), .Z(PRODUCT[241]) );
  AND U17 ( .A(A[240]), .B(B[0]), .Z(PRODUCT[240]) );
  AND U18 ( .A(A[239]), .B(B[0]), .Z(PRODUCT[239]) );
  AND U19 ( .A(A[238]), .B(B[0]), .Z(PRODUCT[238]) );
  AND U20 ( .A(A[237]), .B(B[0]), .Z(PRODUCT[237]) );
  AND U21 ( .A(A[236]), .B(B[0]), .Z(PRODUCT[236]) );
  AND U22 ( .A(A[235]), .B(B[0]), .Z(PRODUCT[235]) );
  AND U23 ( .A(A[234]), .B(B[0]), .Z(PRODUCT[234]) );
  AND U24 ( .A(A[233]), .B(B[0]), .Z(PRODUCT[233]) );
  AND U25 ( .A(A[232]), .B(B[0]), .Z(PRODUCT[232]) );
  AND U26 ( .A(A[231]), .B(B[0]), .Z(PRODUCT[231]) );
  AND U27 ( .A(A[230]), .B(B[0]), .Z(PRODUCT[230]) );
  AND U28 ( .A(A[229]), .B(B[0]), .Z(PRODUCT[229]) );
  AND U29 ( .A(A[228]), .B(B[0]), .Z(PRODUCT[228]) );
  AND U30 ( .A(A[227]), .B(B[0]), .Z(PRODUCT[227]) );
  AND U31 ( .A(A[226]), .B(B[0]), .Z(PRODUCT[226]) );
  AND U32 ( .A(A[225]), .B(B[0]), .Z(PRODUCT[225]) );
  AND U33 ( .A(A[224]), .B(B[0]), .Z(PRODUCT[224]) );
  AND U34 ( .A(A[223]), .B(B[0]), .Z(PRODUCT[223]) );
  AND U35 ( .A(A[222]), .B(B[0]), .Z(PRODUCT[222]) );
  AND U36 ( .A(A[221]), .B(B[0]), .Z(PRODUCT[221]) );
  AND U37 ( .A(A[220]), .B(B[0]), .Z(PRODUCT[220]) );
  AND U38 ( .A(A[219]), .B(B[0]), .Z(PRODUCT[219]) );
  AND U39 ( .A(A[218]), .B(B[0]), .Z(PRODUCT[218]) );
  AND U40 ( .A(A[217]), .B(B[0]), .Z(PRODUCT[217]) );
  AND U41 ( .A(A[216]), .B(B[0]), .Z(PRODUCT[216]) );
  AND U42 ( .A(A[215]), .B(B[0]), .Z(PRODUCT[215]) );
  AND U43 ( .A(A[214]), .B(B[0]), .Z(PRODUCT[214]) );
  AND U44 ( .A(A[213]), .B(B[0]), .Z(PRODUCT[213]) );
  AND U45 ( .A(A[212]), .B(B[0]), .Z(PRODUCT[212]) );
  AND U46 ( .A(A[211]), .B(B[0]), .Z(PRODUCT[211]) );
  AND U47 ( .A(A[210]), .B(B[0]), .Z(PRODUCT[210]) );
  AND U48 ( .A(A[209]), .B(B[0]), .Z(PRODUCT[209]) );
  AND U49 ( .A(A[208]), .B(B[0]), .Z(PRODUCT[208]) );
  AND U50 ( .A(A[207]), .B(B[0]), .Z(PRODUCT[207]) );
  AND U51 ( .A(A[206]), .B(B[0]), .Z(PRODUCT[206]) );
  AND U52 ( .A(A[205]), .B(B[0]), .Z(PRODUCT[205]) );
  AND U53 ( .A(A[204]), .B(B[0]), .Z(PRODUCT[204]) );
  AND U54 ( .A(A[203]), .B(B[0]), .Z(PRODUCT[203]) );
  AND U55 ( .A(A[202]), .B(B[0]), .Z(PRODUCT[202]) );
  AND U56 ( .A(A[201]), .B(B[0]), .Z(PRODUCT[201]) );
  AND U57 ( .A(A[200]), .B(B[0]), .Z(PRODUCT[200]) );
  AND U58 ( .A(A[199]), .B(B[0]), .Z(PRODUCT[199]) );
  AND U59 ( .A(A[198]), .B(B[0]), .Z(PRODUCT[198]) );
  AND U60 ( .A(A[197]), .B(B[0]), .Z(PRODUCT[197]) );
  AND U61 ( .A(A[196]), .B(B[0]), .Z(PRODUCT[196]) );
  AND U62 ( .A(A[195]), .B(B[0]), .Z(PRODUCT[195]) );
  AND U63 ( .A(A[194]), .B(B[0]), .Z(PRODUCT[194]) );
  AND U64 ( .A(A[193]), .B(B[0]), .Z(PRODUCT[193]) );
  AND U65 ( .A(A[192]), .B(B[0]), .Z(PRODUCT[192]) );
  AND U66 ( .A(A[191]), .B(B[0]), .Z(PRODUCT[191]) );
  AND U67 ( .A(A[190]), .B(B[0]), .Z(PRODUCT[190]) );
  AND U68 ( .A(A[189]), .B(B[0]), .Z(PRODUCT[189]) );
  AND U69 ( .A(A[188]), .B(B[0]), .Z(PRODUCT[188]) );
  AND U70 ( .A(A[187]), .B(B[0]), .Z(PRODUCT[187]) );
  AND U71 ( .A(A[186]), .B(B[0]), .Z(PRODUCT[186]) );
  AND U72 ( .A(A[185]), .B(B[0]), .Z(PRODUCT[185]) );
  AND U73 ( .A(A[184]), .B(B[0]), .Z(PRODUCT[184]) );
  AND U74 ( .A(A[183]), .B(B[0]), .Z(PRODUCT[183]) );
  AND U75 ( .A(A[182]), .B(B[0]), .Z(PRODUCT[182]) );
  AND U76 ( .A(A[181]), .B(B[0]), .Z(PRODUCT[181]) );
  AND U77 ( .A(A[180]), .B(B[0]), .Z(PRODUCT[180]) );
  AND U78 ( .A(A[179]), .B(B[0]), .Z(PRODUCT[179]) );
  AND U79 ( .A(A[178]), .B(B[0]), .Z(PRODUCT[178]) );
  AND U80 ( .A(A[177]), .B(B[0]), .Z(PRODUCT[177]) );
  AND U81 ( .A(A[176]), .B(B[0]), .Z(PRODUCT[176]) );
  AND U82 ( .A(A[175]), .B(B[0]), .Z(PRODUCT[175]) );
  AND U83 ( .A(A[174]), .B(B[0]), .Z(PRODUCT[174]) );
  AND U84 ( .A(A[173]), .B(B[0]), .Z(PRODUCT[173]) );
  AND U85 ( .A(A[172]), .B(B[0]), .Z(PRODUCT[172]) );
  AND U86 ( .A(A[171]), .B(B[0]), .Z(PRODUCT[171]) );
  AND U87 ( .A(A[170]), .B(B[0]), .Z(PRODUCT[170]) );
  AND U88 ( .A(A[169]), .B(B[0]), .Z(PRODUCT[169]) );
  AND U89 ( .A(A[168]), .B(B[0]), .Z(PRODUCT[168]) );
  AND U90 ( .A(A[167]), .B(B[0]), .Z(PRODUCT[167]) );
  AND U91 ( .A(A[166]), .B(B[0]), .Z(PRODUCT[166]) );
  AND U92 ( .A(A[165]), .B(B[0]), .Z(PRODUCT[165]) );
  AND U93 ( .A(A[164]), .B(B[0]), .Z(PRODUCT[164]) );
  AND U94 ( .A(A[163]), .B(B[0]), .Z(PRODUCT[163]) );
  AND U95 ( .A(A[162]), .B(B[0]), .Z(PRODUCT[162]) );
  AND U96 ( .A(A[161]), .B(B[0]), .Z(PRODUCT[161]) );
  AND U97 ( .A(A[160]), .B(B[0]), .Z(PRODUCT[160]) );
  AND U98 ( .A(A[159]), .B(B[0]), .Z(PRODUCT[159]) );
  AND U99 ( .A(A[158]), .B(B[0]), .Z(PRODUCT[158]) );
  AND U100 ( .A(A[157]), .B(B[0]), .Z(PRODUCT[157]) );
  AND U101 ( .A(A[156]), .B(B[0]), .Z(PRODUCT[156]) );
  AND U102 ( .A(A[155]), .B(B[0]), .Z(PRODUCT[155]) );
  AND U103 ( .A(A[154]), .B(B[0]), .Z(PRODUCT[154]) );
  AND U104 ( .A(A[153]), .B(B[0]), .Z(PRODUCT[153]) );
  AND U105 ( .A(A[152]), .B(B[0]), .Z(PRODUCT[152]) );
  AND U106 ( .A(A[151]), .B(B[0]), .Z(PRODUCT[151]) );
  AND U107 ( .A(A[150]), .B(B[0]), .Z(PRODUCT[150]) );
  AND U108 ( .A(A[149]), .B(B[0]), .Z(PRODUCT[149]) );
  AND U109 ( .A(A[148]), .B(B[0]), .Z(PRODUCT[148]) );
  AND U110 ( .A(A[147]), .B(B[0]), .Z(PRODUCT[147]) );
  AND U111 ( .A(A[146]), .B(B[0]), .Z(PRODUCT[146]) );
  AND U112 ( .A(A[145]), .B(B[0]), .Z(PRODUCT[145]) );
  AND U113 ( .A(A[144]), .B(B[0]), .Z(PRODUCT[144]) );
  AND U114 ( .A(A[143]), .B(B[0]), .Z(PRODUCT[143]) );
  AND U115 ( .A(A[142]), .B(B[0]), .Z(PRODUCT[142]) );
  AND U116 ( .A(A[141]), .B(B[0]), .Z(PRODUCT[141]) );
  AND U117 ( .A(A[140]), .B(B[0]), .Z(PRODUCT[140]) );
  AND U118 ( .A(A[139]), .B(B[0]), .Z(PRODUCT[139]) );
  AND U119 ( .A(A[138]), .B(B[0]), .Z(PRODUCT[138]) );
  AND U120 ( .A(A[137]), .B(B[0]), .Z(PRODUCT[137]) );
  AND U121 ( .A(A[136]), .B(B[0]), .Z(PRODUCT[136]) );
  AND U122 ( .A(A[135]), .B(B[0]), .Z(PRODUCT[135]) );
  AND U123 ( .A(A[134]), .B(B[0]), .Z(PRODUCT[134]) );
  AND U124 ( .A(A[133]), .B(B[0]), .Z(PRODUCT[133]) );
  AND U125 ( .A(A[132]), .B(B[0]), .Z(PRODUCT[132]) );
  AND U126 ( .A(A[131]), .B(B[0]), .Z(PRODUCT[131]) );
  AND U127 ( .A(A[130]), .B(B[0]), .Z(PRODUCT[130]) );
  AND U128 ( .A(A[129]), .B(B[0]), .Z(PRODUCT[129]) );
  AND U129 ( .A(A[128]), .B(B[0]), .Z(PRODUCT[128]) );
  AND U130 ( .A(A[127]), .B(B[0]), .Z(PRODUCT[127]) );
  AND U131 ( .A(A[126]), .B(B[0]), .Z(PRODUCT[126]) );
  AND U132 ( .A(A[125]), .B(B[0]), .Z(PRODUCT[125]) );
  AND U133 ( .A(A[124]), .B(B[0]), .Z(PRODUCT[124]) );
  AND U134 ( .A(A[123]), .B(B[0]), .Z(PRODUCT[123]) );
  AND U135 ( .A(A[122]), .B(B[0]), .Z(PRODUCT[122]) );
  AND U136 ( .A(A[121]), .B(B[0]), .Z(PRODUCT[121]) );
  AND U137 ( .A(A[120]), .B(B[0]), .Z(PRODUCT[120]) );
  AND U138 ( .A(A[119]), .B(B[0]), .Z(PRODUCT[119]) );
  AND U139 ( .A(A[118]), .B(B[0]), .Z(PRODUCT[118]) );
  AND U140 ( .A(A[117]), .B(B[0]), .Z(PRODUCT[117]) );
  AND U141 ( .A(A[116]), .B(B[0]), .Z(PRODUCT[116]) );
  AND U142 ( .A(A[115]), .B(B[0]), .Z(PRODUCT[115]) );
  AND U143 ( .A(A[114]), .B(B[0]), .Z(PRODUCT[114]) );
  AND U144 ( .A(A[113]), .B(B[0]), .Z(PRODUCT[113]) );
  AND U145 ( .A(A[112]), .B(B[0]), .Z(PRODUCT[112]) );
  AND U146 ( .A(A[111]), .B(B[0]), .Z(PRODUCT[111]) );
  AND U147 ( .A(A[110]), .B(B[0]), .Z(PRODUCT[110]) );
  AND U148 ( .A(A[109]), .B(B[0]), .Z(PRODUCT[109]) );
  AND U149 ( .A(A[108]), .B(B[0]), .Z(PRODUCT[108]) );
  AND U150 ( .A(A[107]), .B(B[0]), .Z(PRODUCT[107]) );
  AND U151 ( .A(A[106]), .B(B[0]), .Z(PRODUCT[106]) );
  AND U152 ( .A(A[105]), .B(B[0]), .Z(PRODUCT[105]) );
  AND U153 ( .A(A[104]), .B(B[0]), .Z(PRODUCT[104]) );
  AND U154 ( .A(A[103]), .B(B[0]), .Z(PRODUCT[103]) );
  AND U155 ( .A(A[102]), .B(B[0]), .Z(PRODUCT[102]) );
  AND U156 ( .A(A[101]), .B(B[0]), .Z(PRODUCT[101]) );
  AND U157 ( .A(A[100]), .B(B[0]), .Z(PRODUCT[100]) );
  AND U158 ( .A(A[99]), .B(B[0]), .Z(PRODUCT[99]) );
  AND U159 ( .A(A[98]), .B(B[0]), .Z(PRODUCT[98]) );
  AND U160 ( .A(A[97]), .B(B[0]), .Z(PRODUCT[97]) );
  AND U161 ( .A(A[96]), .B(B[0]), .Z(PRODUCT[96]) );
  AND U162 ( .A(A[95]), .B(B[0]), .Z(PRODUCT[95]) );
  AND U163 ( .A(A[94]), .B(B[0]), .Z(PRODUCT[94]) );
  AND U164 ( .A(A[93]), .B(B[0]), .Z(PRODUCT[93]) );
  AND U165 ( .A(A[92]), .B(B[0]), .Z(PRODUCT[92]) );
  AND U166 ( .A(A[91]), .B(B[0]), .Z(PRODUCT[91]) );
  AND U167 ( .A(A[90]), .B(B[0]), .Z(PRODUCT[90]) );
  AND U168 ( .A(A[89]), .B(B[0]), .Z(PRODUCT[89]) );
  AND U169 ( .A(A[88]), .B(B[0]), .Z(PRODUCT[88]) );
  AND U170 ( .A(A[87]), .B(B[0]), .Z(PRODUCT[87]) );
  AND U171 ( .A(A[86]), .B(B[0]), .Z(PRODUCT[86]) );
  AND U172 ( .A(A[85]), .B(B[0]), .Z(PRODUCT[85]) );
  AND U173 ( .A(A[84]), .B(B[0]), .Z(PRODUCT[84]) );
  AND U174 ( .A(A[83]), .B(B[0]), .Z(PRODUCT[83]) );
  AND U175 ( .A(A[82]), .B(B[0]), .Z(PRODUCT[82]) );
  AND U176 ( .A(A[81]), .B(B[0]), .Z(PRODUCT[81]) );
  AND U177 ( .A(A[80]), .B(B[0]), .Z(PRODUCT[80]) );
  AND U178 ( .A(A[79]), .B(B[0]), .Z(PRODUCT[79]) );
  AND U179 ( .A(A[78]), .B(B[0]), .Z(PRODUCT[78]) );
  AND U180 ( .A(A[77]), .B(B[0]), .Z(PRODUCT[77]) );
  AND U181 ( .A(A[76]), .B(B[0]), .Z(PRODUCT[76]) );
  AND U182 ( .A(A[75]), .B(B[0]), .Z(PRODUCT[75]) );
  AND U183 ( .A(A[74]), .B(B[0]), .Z(PRODUCT[74]) );
  AND U184 ( .A(A[73]), .B(B[0]), .Z(PRODUCT[73]) );
  AND U185 ( .A(A[72]), .B(B[0]), .Z(PRODUCT[72]) );
  AND U186 ( .A(A[71]), .B(B[0]), .Z(PRODUCT[71]) );
  AND U187 ( .A(A[70]), .B(B[0]), .Z(PRODUCT[70]) );
  AND U188 ( .A(A[69]), .B(B[0]), .Z(PRODUCT[69]) );
  AND U189 ( .A(A[68]), .B(B[0]), .Z(PRODUCT[68]) );
  AND U190 ( .A(A[67]), .B(B[0]), .Z(PRODUCT[67]) );
  AND U191 ( .A(A[66]), .B(B[0]), .Z(PRODUCT[66]) );
  AND U192 ( .A(A[65]), .B(B[0]), .Z(PRODUCT[65]) );
  AND U193 ( .A(A[64]), .B(B[0]), .Z(PRODUCT[64]) );
  AND U194 ( .A(A[63]), .B(B[0]), .Z(PRODUCT[63]) );
  AND U195 ( .A(A[62]), .B(B[0]), .Z(PRODUCT[62]) );
  AND U196 ( .A(A[61]), .B(B[0]), .Z(PRODUCT[61]) );
  AND U197 ( .A(A[60]), .B(B[0]), .Z(PRODUCT[60]) );
  AND U198 ( .A(A[59]), .B(B[0]), .Z(PRODUCT[59]) );
  AND U199 ( .A(A[58]), .B(B[0]), .Z(PRODUCT[58]) );
  AND U200 ( .A(A[57]), .B(B[0]), .Z(PRODUCT[57]) );
  AND U201 ( .A(A[56]), .B(B[0]), .Z(PRODUCT[56]) );
  AND U202 ( .A(A[55]), .B(B[0]), .Z(PRODUCT[55]) );
  AND U203 ( .A(A[54]), .B(B[0]), .Z(PRODUCT[54]) );
  AND U204 ( .A(A[53]), .B(B[0]), .Z(PRODUCT[53]) );
  AND U205 ( .A(A[52]), .B(B[0]), .Z(PRODUCT[52]) );
  AND U206 ( .A(A[51]), .B(B[0]), .Z(PRODUCT[51]) );
  AND U207 ( .A(A[50]), .B(B[0]), .Z(PRODUCT[50]) );
  AND U208 ( .A(A[49]), .B(B[0]), .Z(PRODUCT[49]) );
  AND U209 ( .A(A[48]), .B(B[0]), .Z(PRODUCT[48]) );
  AND U210 ( .A(A[47]), .B(B[0]), .Z(PRODUCT[47]) );
  AND U211 ( .A(A[46]), .B(B[0]), .Z(PRODUCT[46]) );
  AND U212 ( .A(A[45]), .B(B[0]), .Z(PRODUCT[45]) );
  AND U213 ( .A(A[44]), .B(B[0]), .Z(PRODUCT[44]) );
  AND U214 ( .A(A[43]), .B(B[0]), .Z(PRODUCT[43]) );
  AND U215 ( .A(A[42]), .B(B[0]), .Z(PRODUCT[42]) );
  AND U216 ( .A(A[41]), .B(B[0]), .Z(PRODUCT[41]) );
  AND U217 ( .A(A[40]), .B(B[0]), .Z(PRODUCT[40]) );
  AND U218 ( .A(A[39]), .B(B[0]), .Z(PRODUCT[39]) );
  AND U219 ( .A(A[38]), .B(B[0]), .Z(PRODUCT[38]) );
  AND U220 ( .A(A[37]), .B(B[0]), .Z(PRODUCT[37]) );
  AND U221 ( .A(A[36]), .B(B[0]), .Z(PRODUCT[36]) );
  AND U222 ( .A(A[35]), .B(B[0]), .Z(PRODUCT[35]) );
  AND U223 ( .A(A[34]), .B(B[0]), .Z(PRODUCT[34]) );
  AND U224 ( .A(A[33]), .B(B[0]), .Z(PRODUCT[33]) );
  AND U225 ( .A(A[32]), .B(B[0]), .Z(PRODUCT[32]) );
  AND U226 ( .A(A[31]), .B(B[0]), .Z(PRODUCT[31]) );
  AND U227 ( .A(A[30]), .B(B[0]), .Z(PRODUCT[30]) );
  AND U228 ( .A(A[29]), .B(B[0]), .Z(PRODUCT[29]) );
  AND U229 ( .A(A[28]), .B(B[0]), .Z(PRODUCT[28]) );
  AND U230 ( .A(A[27]), .B(B[0]), .Z(PRODUCT[27]) );
  AND U231 ( .A(A[26]), .B(B[0]), .Z(PRODUCT[26]) );
  AND U232 ( .A(A[25]), .B(B[0]), .Z(PRODUCT[25]) );
  AND U233 ( .A(A[24]), .B(B[0]), .Z(PRODUCT[24]) );
  AND U234 ( .A(A[23]), .B(B[0]), .Z(PRODUCT[23]) );
  AND U235 ( .A(A[22]), .B(B[0]), .Z(PRODUCT[22]) );
  AND U236 ( .A(A[21]), .B(B[0]), .Z(PRODUCT[21]) );
  AND U237 ( .A(A[20]), .B(B[0]), .Z(PRODUCT[20]) );
  AND U238 ( .A(A[19]), .B(B[0]), .Z(PRODUCT[19]) );
  AND U239 ( .A(A[18]), .B(B[0]), .Z(PRODUCT[18]) );
  AND U240 ( .A(A[17]), .B(B[0]), .Z(PRODUCT[17]) );
  AND U241 ( .A(A[16]), .B(B[0]), .Z(PRODUCT[16]) );
  AND U242 ( .A(A[15]), .B(B[0]), .Z(PRODUCT[15]) );
  AND U243 ( .A(A[14]), .B(B[0]), .Z(PRODUCT[14]) );
  AND U244 ( .A(A[13]), .B(B[0]), .Z(PRODUCT[13]) );
  AND U245 ( .A(A[12]), .B(B[0]), .Z(PRODUCT[12]) );
  AND U246 ( .A(A[11]), .B(B[0]), .Z(PRODUCT[11]) );
  AND U247 ( .A(A[10]), .B(B[0]), .Z(PRODUCT[10]) );
  AND U248 ( .A(B[0]), .B(A[9]), .Z(PRODUCT[9]) );
  AND U249 ( .A(A[8]), .B(B[0]), .Z(PRODUCT[8]) );
  AND U250 ( .A(A[7]), .B(B[0]), .Z(PRODUCT[7]) );
  AND U251 ( .A(A[6]), .B(B[0]), .Z(PRODUCT[6]) );
  AND U252 ( .A(A[5]), .B(B[0]), .Z(PRODUCT[5]) );
  AND U253 ( .A(A[4]), .B(B[0]), .Z(PRODUCT[4]) );
  AND U254 ( .A(A[3]), .B(B[0]), .Z(PRODUCT[3]) );
  AND U255 ( .A(A[2]), .B(B[0]), .Z(PRODUCT[2]) );
  AND U256 ( .A(A[1]), .B(B[0]), .Z(PRODUCT[1]) );
  AND U257 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
endmodule


module modmult_step_N256_2_DW01_cmp2_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [257:0] A;
  input [257:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;

  NAND U1 ( .A(n1), .B(n2), .Z(LT_LE) );
  NOR U2 ( .A(B[257]), .B(B[256]), .Z(n2) );
  AND U3 ( .A(n3), .B(n4), .Z(n1) );
  NAND U4 ( .A(n5), .B(n6), .Z(n4) );
  NANDN U5 ( .A(B[255]), .B(A[255]), .Z(n6) );
  NAND U6 ( .A(n7), .B(n8), .Z(n5) );
  NANDN U7 ( .A(A[254]), .B(B[254]), .Z(n8) );
  NAND U8 ( .A(n9), .B(n10), .Z(n7) );
  NANDN U9 ( .A(B[254]), .B(A[254]), .Z(n10) );
  AND U10 ( .A(n11), .B(n12), .Z(n9) );
  NAND U11 ( .A(n13), .B(n14), .Z(n12) );
  NANDN U12 ( .A(A[253]), .B(B[253]), .Z(n14) );
  AND U13 ( .A(n15), .B(n16), .Z(n13) );
  NANDN U14 ( .A(A[252]), .B(B[252]), .Z(n16) );
  NAND U15 ( .A(n17), .B(n18), .Z(n15) );
  NANDN U16 ( .A(B[252]), .B(A[252]), .Z(n18) );
  AND U17 ( .A(n19), .B(n20), .Z(n17) );
  NAND U18 ( .A(n21), .B(n22), .Z(n20) );
  NANDN U19 ( .A(A[251]), .B(B[251]), .Z(n22) );
  AND U20 ( .A(n23), .B(n24), .Z(n21) );
  NANDN U21 ( .A(A[250]), .B(B[250]), .Z(n24) );
  NAND U22 ( .A(n25), .B(n26), .Z(n23) );
  NANDN U23 ( .A(B[250]), .B(A[250]), .Z(n26) );
  AND U24 ( .A(n27), .B(n28), .Z(n25) );
  NAND U25 ( .A(n29), .B(n30), .Z(n28) );
  NANDN U26 ( .A(A[249]), .B(B[249]), .Z(n30) );
  AND U27 ( .A(n31), .B(n32), .Z(n29) );
  NANDN U28 ( .A(A[248]), .B(B[248]), .Z(n32) );
  NAND U29 ( .A(n33), .B(n34), .Z(n31) );
  NANDN U30 ( .A(B[248]), .B(A[248]), .Z(n34) );
  AND U31 ( .A(n35), .B(n36), .Z(n33) );
  NAND U32 ( .A(n37), .B(n38), .Z(n36) );
  NANDN U33 ( .A(A[247]), .B(B[247]), .Z(n38) );
  AND U34 ( .A(n39), .B(n40), .Z(n37) );
  NANDN U35 ( .A(A[246]), .B(B[246]), .Z(n40) );
  NAND U36 ( .A(n41), .B(n42), .Z(n39) );
  NANDN U37 ( .A(B[246]), .B(A[246]), .Z(n42) );
  AND U38 ( .A(n43), .B(n44), .Z(n41) );
  NAND U39 ( .A(n45), .B(n46), .Z(n44) );
  NANDN U40 ( .A(A[245]), .B(B[245]), .Z(n46) );
  AND U41 ( .A(n47), .B(n48), .Z(n45) );
  NANDN U42 ( .A(A[244]), .B(B[244]), .Z(n48) );
  NAND U43 ( .A(n49), .B(n50), .Z(n47) );
  NANDN U44 ( .A(B[244]), .B(A[244]), .Z(n50) );
  AND U45 ( .A(n51), .B(n52), .Z(n49) );
  NAND U46 ( .A(n53), .B(n54), .Z(n52) );
  NANDN U47 ( .A(A[243]), .B(B[243]), .Z(n54) );
  AND U48 ( .A(n55), .B(n56), .Z(n53) );
  NANDN U49 ( .A(A[242]), .B(B[242]), .Z(n56) );
  NAND U50 ( .A(n57), .B(n58), .Z(n55) );
  NANDN U51 ( .A(B[242]), .B(A[242]), .Z(n58) );
  AND U52 ( .A(n59), .B(n60), .Z(n57) );
  NAND U53 ( .A(n61), .B(n62), .Z(n60) );
  NANDN U54 ( .A(A[241]), .B(B[241]), .Z(n62) );
  AND U55 ( .A(n63), .B(n64), .Z(n61) );
  NANDN U56 ( .A(A[240]), .B(B[240]), .Z(n64) );
  NAND U57 ( .A(n65), .B(n66), .Z(n63) );
  NANDN U58 ( .A(B[240]), .B(A[240]), .Z(n66) );
  AND U59 ( .A(n67), .B(n68), .Z(n65) );
  NAND U60 ( .A(n69), .B(n70), .Z(n68) );
  NANDN U61 ( .A(A[239]), .B(B[239]), .Z(n70) );
  AND U62 ( .A(n71), .B(n72), .Z(n69) );
  NANDN U63 ( .A(A[238]), .B(B[238]), .Z(n72) );
  NAND U64 ( .A(n73), .B(n74), .Z(n71) );
  NANDN U65 ( .A(B[238]), .B(A[238]), .Z(n74) );
  AND U66 ( .A(n75), .B(n76), .Z(n73) );
  NAND U67 ( .A(n77), .B(n78), .Z(n76) );
  NANDN U68 ( .A(A[237]), .B(B[237]), .Z(n78) );
  AND U69 ( .A(n79), .B(n80), .Z(n77) );
  NANDN U70 ( .A(A[236]), .B(B[236]), .Z(n80) );
  NAND U71 ( .A(n81), .B(n82), .Z(n79) );
  NANDN U72 ( .A(B[236]), .B(A[236]), .Z(n82) );
  AND U73 ( .A(n83), .B(n84), .Z(n81) );
  NAND U74 ( .A(n85), .B(n86), .Z(n84) );
  NANDN U75 ( .A(A[235]), .B(B[235]), .Z(n86) );
  AND U76 ( .A(n87), .B(n88), .Z(n85) );
  NANDN U77 ( .A(A[234]), .B(B[234]), .Z(n88) );
  NAND U78 ( .A(n89), .B(n90), .Z(n87) );
  NANDN U79 ( .A(B[234]), .B(A[234]), .Z(n90) );
  AND U80 ( .A(n91), .B(n92), .Z(n89) );
  NAND U81 ( .A(n93), .B(n94), .Z(n92) );
  NANDN U82 ( .A(A[233]), .B(B[233]), .Z(n94) );
  AND U83 ( .A(n95), .B(n96), .Z(n93) );
  NANDN U84 ( .A(A[232]), .B(B[232]), .Z(n96) );
  NAND U85 ( .A(n97), .B(n98), .Z(n95) );
  NANDN U86 ( .A(B[232]), .B(A[232]), .Z(n98) );
  AND U87 ( .A(n99), .B(n100), .Z(n97) );
  NAND U88 ( .A(n101), .B(n102), .Z(n100) );
  NANDN U89 ( .A(A[231]), .B(B[231]), .Z(n102) );
  AND U90 ( .A(n103), .B(n104), .Z(n101) );
  NANDN U91 ( .A(A[230]), .B(B[230]), .Z(n104) );
  NAND U92 ( .A(n105), .B(n106), .Z(n103) );
  NANDN U93 ( .A(B[230]), .B(A[230]), .Z(n106) );
  AND U94 ( .A(n107), .B(n108), .Z(n105) );
  NAND U95 ( .A(n109), .B(n110), .Z(n108) );
  NANDN U96 ( .A(A[229]), .B(B[229]), .Z(n110) );
  AND U97 ( .A(n111), .B(n112), .Z(n109) );
  NANDN U98 ( .A(A[228]), .B(B[228]), .Z(n112) );
  NAND U99 ( .A(n113), .B(n114), .Z(n111) );
  NANDN U100 ( .A(B[228]), .B(A[228]), .Z(n114) );
  AND U101 ( .A(n115), .B(n116), .Z(n113) );
  NAND U102 ( .A(n117), .B(n118), .Z(n116) );
  NANDN U103 ( .A(A[227]), .B(B[227]), .Z(n118) );
  AND U104 ( .A(n119), .B(n120), .Z(n117) );
  NANDN U105 ( .A(A[226]), .B(B[226]), .Z(n120) );
  NAND U106 ( .A(n121), .B(n122), .Z(n119) );
  NANDN U107 ( .A(B[226]), .B(A[226]), .Z(n122) );
  AND U108 ( .A(n123), .B(n124), .Z(n121) );
  NAND U109 ( .A(n125), .B(n126), .Z(n124) );
  NANDN U110 ( .A(A[225]), .B(B[225]), .Z(n126) );
  AND U111 ( .A(n127), .B(n128), .Z(n125) );
  NANDN U112 ( .A(A[224]), .B(B[224]), .Z(n128) );
  NAND U113 ( .A(n129), .B(n130), .Z(n127) );
  NANDN U114 ( .A(B[224]), .B(A[224]), .Z(n130) );
  AND U115 ( .A(n131), .B(n132), .Z(n129) );
  NAND U116 ( .A(n133), .B(n134), .Z(n132) );
  NANDN U117 ( .A(A[223]), .B(B[223]), .Z(n134) );
  AND U118 ( .A(n135), .B(n136), .Z(n133) );
  NANDN U119 ( .A(A[222]), .B(B[222]), .Z(n136) );
  NAND U120 ( .A(n137), .B(n138), .Z(n135) );
  NANDN U121 ( .A(B[222]), .B(A[222]), .Z(n138) );
  AND U122 ( .A(n139), .B(n140), .Z(n137) );
  NAND U123 ( .A(n141), .B(n142), .Z(n140) );
  NANDN U124 ( .A(A[221]), .B(B[221]), .Z(n142) );
  AND U125 ( .A(n143), .B(n144), .Z(n141) );
  NANDN U126 ( .A(A[220]), .B(B[220]), .Z(n144) );
  NAND U127 ( .A(n145), .B(n146), .Z(n143) );
  NANDN U128 ( .A(B[220]), .B(A[220]), .Z(n146) );
  AND U129 ( .A(n147), .B(n148), .Z(n145) );
  NAND U130 ( .A(n149), .B(n150), .Z(n148) );
  NANDN U131 ( .A(A[219]), .B(B[219]), .Z(n150) );
  AND U132 ( .A(n151), .B(n152), .Z(n149) );
  NANDN U133 ( .A(A[218]), .B(B[218]), .Z(n152) );
  NAND U134 ( .A(n153), .B(n154), .Z(n151) );
  NANDN U135 ( .A(B[218]), .B(A[218]), .Z(n154) );
  AND U136 ( .A(n155), .B(n156), .Z(n153) );
  NAND U137 ( .A(n157), .B(n158), .Z(n156) );
  NANDN U138 ( .A(A[217]), .B(B[217]), .Z(n158) );
  AND U139 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U140 ( .A(A[216]), .B(B[216]), .Z(n160) );
  NAND U141 ( .A(n161), .B(n162), .Z(n159) );
  NANDN U142 ( .A(B[216]), .B(A[216]), .Z(n162) );
  AND U143 ( .A(n163), .B(n164), .Z(n161) );
  NAND U144 ( .A(n165), .B(n166), .Z(n164) );
  NANDN U145 ( .A(A[215]), .B(B[215]), .Z(n166) );
  AND U146 ( .A(n167), .B(n168), .Z(n165) );
  NANDN U147 ( .A(A[214]), .B(B[214]), .Z(n168) );
  NAND U148 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U149 ( .A(B[214]), .B(A[214]), .Z(n170) );
  AND U150 ( .A(n171), .B(n172), .Z(n169) );
  NAND U151 ( .A(n173), .B(n174), .Z(n172) );
  NANDN U152 ( .A(A[213]), .B(B[213]), .Z(n174) );
  AND U153 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U154 ( .A(A[212]), .B(B[212]), .Z(n176) );
  NAND U155 ( .A(n177), .B(n178), .Z(n175) );
  NANDN U156 ( .A(B[212]), .B(A[212]), .Z(n178) );
  AND U157 ( .A(n179), .B(n180), .Z(n177) );
  NAND U158 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U159 ( .A(A[211]), .B(B[211]), .Z(n182) );
  AND U160 ( .A(n183), .B(n184), .Z(n181) );
  NANDN U161 ( .A(A[210]), .B(B[210]), .Z(n184) );
  NAND U162 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U163 ( .A(B[210]), .B(A[210]), .Z(n186) );
  AND U164 ( .A(n187), .B(n188), .Z(n185) );
  NAND U165 ( .A(n189), .B(n190), .Z(n188) );
  NANDN U166 ( .A(A[209]), .B(B[209]), .Z(n190) );
  AND U167 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U168 ( .A(A[208]), .B(B[208]), .Z(n192) );
  NAND U169 ( .A(n193), .B(n194), .Z(n191) );
  NANDN U170 ( .A(B[208]), .B(A[208]), .Z(n194) );
  AND U171 ( .A(n195), .B(n196), .Z(n193) );
  NAND U172 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U173 ( .A(A[207]), .B(B[207]), .Z(n198) );
  AND U174 ( .A(n199), .B(n200), .Z(n197) );
  NANDN U175 ( .A(A[206]), .B(B[206]), .Z(n200) );
  NAND U176 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U177 ( .A(B[206]), .B(A[206]), .Z(n202) );
  AND U178 ( .A(n203), .B(n204), .Z(n201) );
  NAND U179 ( .A(n205), .B(n206), .Z(n204) );
  NANDN U180 ( .A(A[205]), .B(B[205]), .Z(n206) );
  AND U181 ( .A(n207), .B(n208), .Z(n205) );
  NANDN U182 ( .A(A[204]), .B(B[204]), .Z(n208) );
  NAND U183 ( .A(n209), .B(n210), .Z(n207) );
  NANDN U184 ( .A(B[204]), .B(A[204]), .Z(n210) );
  AND U185 ( .A(n211), .B(n212), .Z(n209) );
  NAND U186 ( .A(n213), .B(n214), .Z(n212) );
  NANDN U187 ( .A(A[203]), .B(B[203]), .Z(n214) );
  AND U188 ( .A(n215), .B(n216), .Z(n213) );
  NANDN U189 ( .A(A[202]), .B(B[202]), .Z(n216) );
  NAND U190 ( .A(n217), .B(n218), .Z(n215) );
  NANDN U191 ( .A(B[202]), .B(A[202]), .Z(n218) );
  AND U192 ( .A(n219), .B(n220), .Z(n217) );
  NAND U193 ( .A(n221), .B(n222), .Z(n220) );
  NANDN U194 ( .A(A[201]), .B(B[201]), .Z(n222) );
  AND U195 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U196 ( .A(A[200]), .B(B[200]), .Z(n224) );
  NAND U197 ( .A(n225), .B(n226), .Z(n223) );
  NANDN U198 ( .A(B[200]), .B(A[200]), .Z(n226) );
  AND U199 ( .A(n227), .B(n228), .Z(n225) );
  NAND U200 ( .A(n229), .B(n230), .Z(n228) );
  NANDN U201 ( .A(A[199]), .B(B[199]), .Z(n230) );
  AND U202 ( .A(n231), .B(n232), .Z(n229) );
  NANDN U203 ( .A(A[198]), .B(B[198]), .Z(n232) );
  NAND U204 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U205 ( .A(B[198]), .B(A[198]), .Z(n234) );
  AND U206 ( .A(n235), .B(n236), .Z(n233) );
  NAND U207 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U208 ( .A(A[197]), .B(B[197]), .Z(n238) );
  AND U209 ( .A(n239), .B(n240), .Z(n237) );
  NANDN U210 ( .A(A[196]), .B(B[196]), .Z(n240) );
  NAND U211 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U212 ( .A(B[196]), .B(A[196]), .Z(n242) );
  AND U213 ( .A(n243), .B(n244), .Z(n241) );
  NAND U214 ( .A(n245), .B(n246), .Z(n244) );
  NANDN U215 ( .A(A[195]), .B(B[195]), .Z(n246) );
  AND U216 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U217 ( .A(A[194]), .B(B[194]), .Z(n248) );
  NAND U218 ( .A(n249), .B(n250), .Z(n247) );
  NANDN U219 ( .A(B[194]), .B(A[194]), .Z(n250) );
  AND U220 ( .A(n251), .B(n252), .Z(n249) );
  NAND U221 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U222 ( .A(A[193]), .B(B[193]), .Z(n254) );
  AND U223 ( .A(n255), .B(n256), .Z(n253) );
  NANDN U224 ( .A(A[192]), .B(B[192]), .Z(n256) );
  NAND U225 ( .A(n257), .B(n258), .Z(n255) );
  NANDN U226 ( .A(B[192]), .B(A[192]), .Z(n258) );
  AND U227 ( .A(n259), .B(n260), .Z(n257) );
  NAND U228 ( .A(n261), .B(n262), .Z(n260) );
  NANDN U229 ( .A(A[191]), .B(B[191]), .Z(n262) );
  AND U230 ( .A(n263), .B(n264), .Z(n261) );
  NANDN U231 ( .A(A[190]), .B(B[190]), .Z(n264) );
  NAND U232 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U233 ( .A(B[190]), .B(A[190]), .Z(n266) );
  AND U234 ( .A(n267), .B(n268), .Z(n265) );
  NAND U235 ( .A(n269), .B(n270), .Z(n268) );
  NANDN U236 ( .A(A[189]), .B(B[189]), .Z(n270) );
  AND U237 ( .A(n271), .B(n272), .Z(n269) );
  NANDN U238 ( .A(A[188]), .B(B[188]), .Z(n272) );
  NAND U239 ( .A(n273), .B(n274), .Z(n271) );
  NANDN U240 ( .A(B[188]), .B(A[188]), .Z(n274) );
  AND U241 ( .A(n275), .B(n276), .Z(n273) );
  NAND U242 ( .A(n277), .B(n278), .Z(n276) );
  NANDN U243 ( .A(A[187]), .B(B[187]), .Z(n278) );
  AND U244 ( .A(n279), .B(n280), .Z(n277) );
  NANDN U245 ( .A(A[186]), .B(B[186]), .Z(n280) );
  NAND U246 ( .A(n281), .B(n282), .Z(n279) );
  NANDN U247 ( .A(B[186]), .B(A[186]), .Z(n282) );
  AND U248 ( .A(n283), .B(n284), .Z(n281) );
  NAND U249 ( .A(n285), .B(n286), .Z(n284) );
  NANDN U250 ( .A(A[185]), .B(B[185]), .Z(n286) );
  AND U251 ( .A(n287), .B(n288), .Z(n285) );
  NANDN U252 ( .A(A[184]), .B(B[184]), .Z(n288) );
  NAND U253 ( .A(n289), .B(n290), .Z(n287) );
  NANDN U254 ( .A(B[184]), .B(A[184]), .Z(n290) );
  AND U255 ( .A(n291), .B(n292), .Z(n289) );
  NAND U256 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U257 ( .A(A[183]), .B(B[183]), .Z(n294) );
  AND U258 ( .A(n295), .B(n296), .Z(n293) );
  NANDN U259 ( .A(A[182]), .B(B[182]), .Z(n296) );
  NAND U260 ( .A(n297), .B(n298), .Z(n295) );
  NANDN U261 ( .A(B[182]), .B(A[182]), .Z(n298) );
  AND U262 ( .A(n299), .B(n300), .Z(n297) );
  NAND U263 ( .A(n301), .B(n302), .Z(n300) );
  NANDN U264 ( .A(A[181]), .B(B[181]), .Z(n302) );
  AND U265 ( .A(n303), .B(n304), .Z(n301) );
  NANDN U266 ( .A(A[180]), .B(B[180]), .Z(n304) );
  NAND U267 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U268 ( .A(B[180]), .B(A[180]), .Z(n306) );
  AND U269 ( .A(n307), .B(n308), .Z(n305) );
  NAND U270 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U271 ( .A(A[179]), .B(B[179]), .Z(n310) );
  AND U272 ( .A(n311), .B(n312), .Z(n309) );
  NANDN U273 ( .A(A[178]), .B(B[178]), .Z(n312) );
  NAND U274 ( .A(n313), .B(n314), .Z(n311) );
  NANDN U275 ( .A(B[178]), .B(A[178]), .Z(n314) );
  AND U276 ( .A(n315), .B(n316), .Z(n313) );
  NAND U277 ( .A(n317), .B(n318), .Z(n316) );
  NANDN U278 ( .A(A[177]), .B(B[177]), .Z(n318) );
  AND U279 ( .A(n319), .B(n320), .Z(n317) );
  NANDN U280 ( .A(A[176]), .B(B[176]), .Z(n320) );
  NAND U281 ( .A(n321), .B(n322), .Z(n319) );
  NANDN U282 ( .A(B[176]), .B(A[176]), .Z(n322) );
  AND U283 ( .A(n323), .B(n324), .Z(n321) );
  NAND U284 ( .A(n325), .B(n326), .Z(n324) );
  NANDN U285 ( .A(A[175]), .B(B[175]), .Z(n326) );
  AND U286 ( .A(n327), .B(n328), .Z(n325) );
  NANDN U287 ( .A(A[174]), .B(B[174]), .Z(n328) );
  NAND U288 ( .A(n329), .B(n330), .Z(n327) );
  NANDN U289 ( .A(B[174]), .B(A[174]), .Z(n330) );
  AND U290 ( .A(n331), .B(n332), .Z(n329) );
  NAND U291 ( .A(n333), .B(n334), .Z(n332) );
  NANDN U292 ( .A(A[173]), .B(B[173]), .Z(n334) );
  AND U293 ( .A(n335), .B(n336), .Z(n333) );
  NANDN U294 ( .A(A[172]), .B(B[172]), .Z(n336) );
  NAND U295 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U296 ( .A(B[172]), .B(A[172]), .Z(n338) );
  AND U297 ( .A(n339), .B(n340), .Z(n337) );
  NAND U298 ( .A(n341), .B(n342), .Z(n340) );
  NANDN U299 ( .A(A[171]), .B(B[171]), .Z(n342) );
  AND U300 ( .A(n343), .B(n344), .Z(n341) );
  NANDN U301 ( .A(A[170]), .B(B[170]), .Z(n344) );
  NAND U302 ( .A(n345), .B(n346), .Z(n343) );
  NANDN U303 ( .A(B[170]), .B(A[170]), .Z(n346) );
  AND U304 ( .A(n347), .B(n348), .Z(n345) );
  NAND U305 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U306 ( .A(A[169]), .B(B[169]), .Z(n350) );
  AND U307 ( .A(n351), .B(n352), .Z(n349) );
  NANDN U308 ( .A(A[168]), .B(B[168]), .Z(n352) );
  NAND U309 ( .A(n353), .B(n354), .Z(n351) );
  NANDN U310 ( .A(B[168]), .B(A[168]), .Z(n354) );
  AND U311 ( .A(n355), .B(n356), .Z(n353) );
  NAND U312 ( .A(n357), .B(n358), .Z(n356) );
  NANDN U313 ( .A(A[167]), .B(B[167]), .Z(n358) );
  AND U314 ( .A(n359), .B(n360), .Z(n357) );
  NANDN U315 ( .A(A[166]), .B(B[166]), .Z(n360) );
  NAND U316 ( .A(n361), .B(n362), .Z(n359) );
  NANDN U317 ( .A(B[166]), .B(A[166]), .Z(n362) );
  AND U318 ( .A(n363), .B(n364), .Z(n361) );
  NAND U319 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U320 ( .A(A[165]), .B(B[165]), .Z(n366) );
  AND U321 ( .A(n367), .B(n368), .Z(n365) );
  NANDN U322 ( .A(A[164]), .B(B[164]), .Z(n368) );
  NAND U323 ( .A(n369), .B(n370), .Z(n367) );
  NANDN U324 ( .A(B[164]), .B(A[164]), .Z(n370) );
  AND U325 ( .A(n371), .B(n372), .Z(n369) );
  NAND U326 ( .A(n373), .B(n374), .Z(n372) );
  NANDN U327 ( .A(A[163]), .B(B[163]), .Z(n374) );
  AND U328 ( .A(n375), .B(n376), .Z(n373) );
  NANDN U329 ( .A(A[162]), .B(B[162]), .Z(n376) );
  NAND U330 ( .A(n377), .B(n378), .Z(n375) );
  NANDN U331 ( .A(B[162]), .B(A[162]), .Z(n378) );
  AND U332 ( .A(n379), .B(n380), .Z(n377) );
  NAND U333 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U334 ( .A(A[161]), .B(B[161]), .Z(n382) );
  AND U335 ( .A(n383), .B(n384), .Z(n381) );
  NANDN U336 ( .A(A[160]), .B(B[160]), .Z(n384) );
  NAND U337 ( .A(n385), .B(n386), .Z(n383) );
  NANDN U338 ( .A(B[160]), .B(A[160]), .Z(n386) );
  AND U339 ( .A(n387), .B(n388), .Z(n385) );
  NAND U340 ( .A(n389), .B(n390), .Z(n388) );
  NANDN U341 ( .A(A[159]), .B(B[159]), .Z(n390) );
  AND U342 ( .A(n391), .B(n392), .Z(n389) );
  NANDN U343 ( .A(A[158]), .B(B[158]), .Z(n392) );
  NAND U344 ( .A(n393), .B(n394), .Z(n391) );
  NANDN U345 ( .A(B[158]), .B(A[158]), .Z(n394) );
  AND U346 ( .A(n395), .B(n396), .Z(n393) );
  NAND U347 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U348 ( .A(A[157]), .B(B[157]), .Z(n398) );
  AND U349 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U350 ( .A(A[156]), .B(B[156]), .Z(n400) );
  NAND U351 ( .A(n401), .B(n402), .Z(n399) );
  NANDN U352 ( .A(B[156]), .B(A[156]), .Z(n402) );
  AND U353 ( .A(n403), .B(n404), .Z(n401) );
  NAND U354 ( .A(n405), .B(n406), .Z(n404) );
  NANDN U355 ( .A(A[155]), .B(B[155]), .Z(n406) );
  AND U356 ( .A(n407), .B(n408), .Z(n405) );
  NANDN U357 ( .A(A[154]), .B(B[154]), .Z(n408) );
  NAND U358 ( .A(n409), .B(n410), .Z(n407) );
  NANDN U359 ( .A(B[154]), .B(A[154]), .Z(n410) );
  AND U360 ( .A(n411), .B(n412), .Z(n409) );
  NAND U361 ( .A(n413), .B(n414), .Z(n412) );
  NANDN U362 ( .A(A[153]), .B(B[153]), .Z(n414) );
  AND U363 ( .A(n415), .B(n416), .Z(n413) );
  NANDN U364 ( .A(A[152]), .B(B[152]), .Z(n416) );
  NAND U365 ( .A(n417), .B(n418), .Z(n415) );
  NANDN U366 ( .A(B[152]), .B(A[152]), .Z(n418) );
  AND U367 ( .A(n419), .B(n420), .Z(n417) );
  NAND U368 ( .A(n421), .B(n422), .Z(n420) );
  NANDN U369 ( .A(A[151]), .B(B[151]), .Z(n422) );
  AND U370 ( .A(n423), .B(n424), .Z(n421) );
  NANDN U371 ( .A(A[150]), .B(B[150]), .Z(n424) );
  NAND U372 ( .A(n425), .B(n426), .Z(n423) );
  NANDN U373 ( .A(B[150]), .B(A[150]), .Z(n426) );
  AND U374 ( .A(n427), .B(n428), .Z(n425) );
  NAND U375 ( .A(n429), .B(n430), .Z(n428) );
  NANDN U376 ( .A(A[149]), .B(B[149]), .Z(n430) );
  AND U377 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U378 ( .A(A[148]), .B(B[148]), .Z(n432) );
  NAND U379 ( .A(n433), .B(n434), .Z(n431) );
  NANDN U380 ( .A(B[148]), .B(A[148]), .Z(n434) );
  AND U381 ( .A(n435), .B(n436), .Z(n433) );
  NAND U382 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U383 ( .A(A[147]), .B(B[147]), .Z(n438) );
  AND U384 ( .A(n439), .B(n440), .Z(n437) );
  NANDN U385 ( .A(A[146]), .B(B[146]), .Z(n440) );
  NAND U386 ( .A(n441), .B(n442), .Z(n439) );
  NANDN U387 ( .A(B[146]), .B(A[146]), .Z(n442) );
  AND U388 ( .A(n443), .B(n444), .Z(n441) );
  NAND U389 ( .A(n445), .B(n446), .Z(n444) );
  NANDN U390 ( .A(A[145]), .B(B[145]), .Z(n446) );
  AND U391 ( .A(n447), .B(n448), .Z(n445) );
  NANDN U392 ( .A(A[144]), .B(B[144]), .Z(n448) );
  NAND U393 ( .A(n449), .B(n450), .Z(n447) );
  NANDN U394 ( .A(B[144]), .B(A[144]), .Z(n450) );
  AND U395 ( .A(n451), .B(n452), .Z(n449) );
  NAND U396 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U397 ( .A(A[143]), .B(B[143]), .Z(n454) );
  AND U398 ( .A(n455), .B(n456), .Z(n453) );
  NANDN U399 ( .A(A[142]), .B(B[142]), .Z(n456) );
  NAND U400 ( .A(n457), .B(n458), .Z(n455) );
  NANDN U401 ( .A(B[142]), .B(A[142]), .Z(n458) );
  AND U402 ( .A(n459), .B(n460), .Z(n457) );
  NAND U403 ( .A(n461), .B(n462), .Z(n460) );
  NANDN U404 ( .A(A[141]), .B(B[141]), .Z(n462) );
  AND U405 ( .A(n463), .B(n464), .Z(n461) );
  NANDN U406 ( .A(A[140]), .B(B[140]), .Z(n464) );
  NAND U407 ( .A(n465), .B(n466), .Z(n463) );
  NANDN U408 ( .A(B[140]), .B(A[140]), .Z(n466) );
  AND U409 ( .A(n467), .B(n468), .Z(n465) );
  NAND U410 ( .A(n469), .B(n470), .Z(n468) );
  NANDN U411 ( .A(A[139]), .B(B[139]), .Z(n470) );
  AND U412 ( .A(n471), .B(n472), .Z(n469) );
  NANDN U413 ( .A(A[138]), .B(B[138]), .Z(n472) );
  NAND U414 ( .A(n473), .B(n474), .Z(n471) );
  NANDN U415 ( .A(B[138]), .B(A[138]), .Z(n474) );
  AND U416 ( .A(n475), .B(n476), .Z(n473) );
  NAND U417 ( .A(n477), .B(n478), .Z(n476) );
  NANDN U418 ( .A(A[137]), .B(B[137]), .Z(n478) );
  AND U419 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U420 ( .A(A[136]), .B(B[136]), .Z(n480) );
  NAND U421 ( .A(n481), .B(n482), .Z(n479) );
  NANDN U422 ( .A(B[136]), .B(A[136]), .Z(n482) );
  AND U423 ( .A(n483), .B(n484), .Z(n481) );
  NAND U424 ( .A(n485), .B(n486), .Z(n484) );
  NANDN U425 ( .A(A[135]), .B(B[135]), .Z(n486) );
  AND U426 ( .A(n487), .B(n488), .Z(n485) );
  NANDN U427 ( .A(A[134]), .B(B[134]), .Z(n488) );
  NAND U428 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U429 ( .A(B[134]), .B(A[134]), .Z(n490) );
  AND U430 ( .A(n491), .B(n492), .Z(n489) );
  NAND U431 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U432 ( .A(A[133]), .B(B[133]), .Z(n494) );
  AND U433 ( .A(n495), .B(n496), .Z(n493) );
  NANDN U434 ( .A(A[132]), .B(B[132]), .Z(n496) );
  NAND U435 ( .A(n497), .B(n498), .Z(n495) );
  NANDN U436 ( .A(B[132]), .B(A[132]), .Z(n498) );
  AND U437 ( .A(n499), .B(n500), .Z(n497) );
  NAND U438 ( .A(n501), .B(n502), .Z(n500) );
  NANDN U439 ( .A(A[131]), .B(B[131]), .Z(n502) );
  AND U440 ( .A(n503), .B(n504), .Z(n501) );
  NANDN U441 ( .A(A[130]), .B(B[130]), .Z(n504) );
  NAND U442 ( .A(n505), .B(n506), .Z(n503) );
  NANDN U443 ( .A(B[130]), .B(A[130]), .Z(n506) );
  AND U444 ( .A(n507), .B(n508), .Z(n505) );
  NAND U445 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U446 ( .A(A[129]), .B(B[129]), .Z(n510) );
  AND U447 ( .A(n511), .B(n512), .Z(n509) );
  NANDN U448 ( .A(A[128]), .B(B[128]), .Z(n512) );
  NAND U449 ( .A(n513), .B(n514), .Z(n511) );
  NANDN U450 ( .A(B[128]), .B(A[128]), .Z(n514) );
  AND U451 ( .A(n515), .B(n516), .Z(n513) );
  NAND U452 ( .A(n517), .B(n518), .Z(n516) );
  NANDN U453 ( .A(A[127]), .B(B[127]), .Z(n518) );
  AND U454 ( .A(n519), .B(n520), .Z(n517) );
  NANDN U455 ( .A(A[126]), .B(B[126]), .Z(n520) );
  NAND U456 ( .A(n521), .B(n522), .Z(n519) );
  NANDN U457 ( .A(B[126]), .B(A[126]), .Z(n522) );
  AND U458 ( .A(n523), .B(n524), .Z(n521) );
  NAND U459 ( .A(n525), .B(n526), .Z(n524) );
  NANDN U460 ( .A(A[125]), .B(B[125]), .Z(n526) );
  AND U461 ( .A(n527), .B(n528), .Z(n525) );
  NANDN U462 ( .A(A[124]), .B(B[124]), .Z(n528) );
  NAND U463 ( .A(n529), .B(n530), .Z(n527) );
  NANDN U464 ( .A(B[124]), .B(A[124]), .Z(n530) );
  AND U465 ( .A(n531), .B(n532), .Z(n529) );
  NAND U466 ( .A(n533), .B(n534), .Z(n532) );
  NANDN U467 ( .A(A[123]), .B(B[123]), .Z(n534) );
  AND U468 ( .A(n535), .B(n536), .Z(n533) );
  NANDN U469 ( .A(A[122]), .B(B[122]), .Z(n536) );
  NAND U470 ( .A(n537), .B(n538), .Z(n535) );
  NANDN U471 ( .A(B[122]), .B(A[122]), .Z(n538) );
  AND U472 ( .A(n539), .B(n540), .Z(n537) );
  NAND U473 ( .A(n541), .B(n542), .Z(n540) );
  NANDN U474 ( .A(A[121]), .B(B[121]), .Z(n542) );
  AND U475 ( .A(n543), .B(n544), .Z(n541) );
  NANDN U476 ( .A(A[120]), .B(B[120]), .Z(n544) );
  NAND U477 ( .A(n545), .B(n546), .Z(n543) );
  NANDN U478 ( .A(B[120]), .B(A[120]), .Z(n546) );
  AND U479 ( .A(n547), .B(n548), .Z(n545) );
  NAND U480 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U481 ( .A(A[119]), .B(B[119]), .Z(n550) );
  AND U482 ( .A(n551), .B(n552), .Z(n549) );
  NANDN U483 ( .A(A[118]), .B(B[118]), .Z(n552) );
  NAND U484 ( .A(n553), .B(n554), .Z(n551) );
  NANDN U485 ( .A(B[118]), .B(A[118]), .Z(n554) );
  AND U486 ( .A(n555), .B(n556), .Z(n553) );
  NAND U487 ( .A(n557), .B(n558), .Z(n556) );
  NANDN U488 ( .A(A[117]), .B(B[117]), .Z(n558) );
  AND U489 ( .A(n559), .B(n560), .Z(n557) );
  NANDN U490 ( .A(A[116]), .B(B[116]), .Z(n560) );
  NAND U491 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U492 ( .A(B[116]), .B(A[116]), .Z(n562) );
  AND U493 ( .A(n563), .B(n564), .Z(n561) );
  NAND U494 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U495 ( .A(A[115]), .B(B[115]), .Z(n566) );
  AND U496 ( .A(n567), .B(n568), .Z(n565) );
  NANDN U497 ( .A(A[114]), .B(B[114]), .Z(n568) );
  NAND U498 ( .A(n569), .B(n570), .Z(n567) );
  NANDN U499 ( .A(B[114]), .B(A[114]), .Z(n570) );
  AND U500 ( .A(n571), .B(n572), .Z(n569) );
  NAND U501 ( .A(n573), .B(n574), .Z(n572) );
  NANDN U502 ( .A(A[113]), .B(B[113]), .Z(n574) );
  AND U503 ( .A(n575), .B(n576), .Z(n573) );
  NANDN U504 ( .A(A[112]), .B(B[112]), .Z(n576) );
  NAND U505 ( .A(n577), .B(n578), .Z(n575) );
  NANDN U506 ( .A(B[112]), .B(A[112]), .Z(n578) );
  AND U507 ( .A(n579), .B(n580), .Z(n577) );
  NAND U508 ( .A(n581), .B(n582), .Z(n580) );
  NANDN U509 ( .A(A[111]), .B(B[111]), .Z(n582) );
  AND U510 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U511 ( .A(A[110]), .B(B[110]), .Z(n584) );
  NAND U512 ( .A(n585), .B(n586), .Z(n583) );
  NANDN U513 ( .A(B[110]), .B(A[110]), .Z(n586) );
  AND U514 ( .A(n587), .B(n588), .Z(n585) );
  NAND U515 ( .A(n589), .B(n590), .Z(n588) );
  NANDN U516 ( .A(A[109]), .B(B[109]), .Z(n590) );
  AND U517 ( .A(n591), .B(n592), .Z(n589) );
  NANDN U518 ( .A(A[108]), .B(B[108]), .Z(n592) );
  NAND U519 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U520 ( .A(B[108]), .B(A[108]), .Z(n594) );
  AND U521 ( .A(n595), .B(n596), .Z(n593) );
  NAND U522 ( .A(n597), .B(n598), .Z(n596) );
  NANDN U523 ( .A(A[107]), .B(B[107]), .Z(n598) );
  AND U524 ( .A(n599), .B(n600), .Z(n597) );
  NANDN U525 ( .A(A[106]), .B(B[106]), .Z(n600) );
  NAND U526 ( .A(n601), .B(n602), .Z(n599) );
  NANDN U527 ( .A(B[106]), .B(A[106]), .Z(n602) );
  AND U528 ( .A(n603), .B(n604), .Z(n601) );
  NAND U529 ( .A(n605), .B(n606), .Z(n604) );
  NANDN U530 ( .A(A[105]), .B(B[105]), .Z(n606) );
  AND U531 ( .A(n607), .B(n608), .Z(n605) );
  NANDN U532 ( .A(A[104]), .B(B[104]), .Z(n608) );
  NAND U533 ( .A(n609), .B(n610), .Z(n607) );
  NANDN U534 ( .A(B[104]), .B(A[104]), .Z(n610) );
  AND U535 ( .A(n611), .B(n612), .Z(n609) );
  NAND U536 ( .A(n613), .B(n614), .Z(n612) );
  NANDN U537 ( .A(A[103]), .B(B[103]), .Z(n614) );
  AND U538 ( .A(n615), .B(n616), .Z(n613) );
  NANDN U539 ( .A(A[102]), .B(B[102]), .Z(n616) );
  NAND U540 ( .A(n617), .B(n618), .Z(n615) );
  NANDN U541 ( .A(B[102]), .B(A[102]), .Z(n618) );
  AND U542 ( .A(n619), .B(n620), .Z(n617) );
  NAND U543 ( .A(n621), .B(n622), .Z(n620) );
  NANDN U544 ( .A(A[101]), .B(B[101]), .Z(n622) );
  AND U545 ( .A(n623), .B(n624), .Z(n621) );
  NANDN U546 ( .A(A[100]), .B(B[100]), .Z(n624) );
  NAND U547 ( .A(n625), .B(n626), .Z(n623) );
  NANDN U548 ( .A(B[99]), .B(A[99]), .Z(n626) );
  AND U549 ( .A(n627), .B(n628), .Z(n625) );
  NAND U550 ( .A(n629), .B(n630), .Z(n628) );
  NANDN U551 ( .A(A[99]), .B(B[99]), .Z(n630) );
  AND U552 ( .A(n631), .B(n632), .Z(n629) );
  NANDN U553 ( .A(A[98]), .B(B[98]), .Z(n632) );
  NAND U554 ( .A(n633), .B(n634), .Z(n631) );
  NANDN U555 ( .A(B[98]), .B(A[98]), .Z(n634) );
  AND U556 ( .A(n635), .B(n636), .Z(n633) );
  NAND U557 ( .A(n637), .B(n638), .Z(n636) );
  NANDN U558 ( .A(A[97]), .B(B[97]), .Z(n638) );
  AND U559 ( .A(n639), .B(n640), .Z(n637) );
  NANDN U560 ( .A(A[96]), .B(B[96]), .Z(n640) );
  NAND U561 ( .A(n641), .B(n642), .Z(n639) );
  NANDN U562 ( .A(B[96]), .B(A[96]), .Z(n642) );
  AND U563 ( .A(n643), .B(n644), .Z(n641) );
  NAND U564 ( .A(n645), .B(n646), .Z(n644) );
  NANDN U565 ( .A(A[95]), .B(B[95]), .Z(n646) );
  AND U566 ( .A(n647), .B(n648), .Z(n645) );
  NANDN U567 ( .A(A[94]), .B(B[94]), .Z(n648) );
  NAND U568 ( .A(n649), .B(n650), .Z(n647) );
  NANDN U569 ( .A(B[94]), .B(A[94]), .Z(n650) );
  AND U570 ( .A(n651), .B(n652), .Z(n649) );
  NAND U571 ( .A(n653), .B(n654), .Z(n652) );
  NANDN U572 ( .A(A[93]), .B(B[93]), .Z(n654) );
  AND U573 ( .A(n655), .B(n656), .Z(n653) );
  NANDN U574 ( .A(A[92]), .B(B[92]), .Z(n656) );
  NAND U575 ( .A(n657), .B(n658), .Z(n655) );
  NANDN U576 ( .A(B[92]), .B(A[92]), .Z(n658) );
  AND U577 ( .A(n659), .B(n660), .Z(n657) );
  NAND U578 ( .A(n661), .B(n662), .Z(n660) );
  NANDN U579 ( .A(A[91]), .B(B[91]), .Z(n662) );
  AND U580 ( .A(n663), .B(n664), .Z(n661) );
  NANDN U581 ( .A(A[90]), .B(B[90]), .Z(n664) );
  NAND U582 ( .A(n665), .B(n666), .Z(n663) );
  NANDN U583 ( .A(B[90]), .B(A[90]), .Z(n666) );
  AND U584 ( .A(n667), .B(n668), .Z(n665) );
  NAND U585 ( .A(n669), .B(n670), .Z(n668) );
  NANDN U586 ( .A(A[89]), .B(B[89]), .Z(n670) );
  AND U587 ( .A(n671), .B(n672), .Z(n669) );
  NANDN U588 ( .A(A[88]), .B(B[88]), .Z(n672) );
  NAND U589 ( .A(n673), .B(n674), .Z(n671) );
  NANDN U590 ( .A(B[88]), .B(A[88]), .Z(n674) );
  AND U591 ( .A(n675), .B(n676), .Z(n673) );
  NAND U592 ( .A(n677), .B(n678), .Z(n676) );
  NANDN U593 ( .A(A[87]), .B(B[87]), .Z(n678) );
  AND U594 ( .A(n679), .B(n680), .Z(n677) );
  NANDN U595 ( .A(A[86]), .B(B[86]), .Z(n680) );
  NAND U596 ( .A(n681), .B(n682), .Z(n679) );
  NANDN U597 ( .A(B[86]), .B(A[86]), .Z(n682) );
  AND U598 ( .A(n683), .B(n684), .Z(n681) );
  NAND U599 ( .A(n685), .B(n686), .Z(n684) );
  NANDN U600 ( .A(A[85]), .B(B[85]), .Z(n686) );
  AND U601 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U602 ( .A(A[84]), .B(B[84]), .Z(n688) );
  NAND U603 ( .A(n689), .B(n690), .Z(n687) );
  NANDN U604 ( .A(B[84]), .B(A[84]), .Z(n690) );
  AND U605 ( .A(n691), .B(n692), .Z(n689) );
  NAND U606 ( .A(n693), .B(n694), .Z(n692) );
  NANDN U607 ( .A(A[83]), .B(B[83]), .Z(n694) );
  AND U608 ( .A(n695), .B(n696), .Z(n693) );
  NANDN U609 ( .A(A[82]), .B(B[82]), .Z(n696) );
  NAND U610 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U611 ( .A(B[82]), .B(A[82]), .Z(n698) );
  AND U612 ( .A(n699), .B(n700), .Z(n697) );
  NAND U613 ( .A(n701), .B(n702), .Z(n700) );
  NANDN U614 ( .A(A[81]), .B(B[81]), .Z(n702) );
  AND U615 ( .A(n703), .B(n704), .Z(n701) );
  NANDN U616 ( .A(A[80]), .B(B[80]), .Z(n704) );
  NAND U617 ( .A(n705), .B(n706), .Z(n703) );
  NANDN U618 ( .A(B[80]), .B(A[80]), .Z(n706) );
  AND U619 ( .A(n707), .B(n708), .Z(n705) );
  NAND U620 ( .A(n709), .B(n710), .Z(n708) );
  NANDN U621 ( .A(A[79]), .B(B[79]), .Z(n710) );
  AND U622 ( .A(n711), .B(n712), .Z(n709) );
  NANDN U623 ( .A(A[78]), .B(B[78]), .Z(n712) );
  NAND U624 ( .A(n713), .B(n714), .Z(n711) );
  NANDN U625 ( .A(B[78]), .B(A[78]), .Z(n714) );
  AND U626 ( .A(n715), .B(n716), .Z(n713) );
  NAND U627 ( .A(n717), .B(n718), .Z(n716) );
  NANDN U628 ( .A(A[77]), .B(B[77]), .Z(n718) );
  AND U629 ( .A(n719), .B(n720), .Z(n717) );
  NANDN U630 ( .A(A[76]), .B(B[76]), .Z(n720) );
  NAND U631 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U632 ( .A(B[76]), .B(A[76]), .Z(n722) );
  AND U633 ( .A(n723), .B(n724), .Z(n721) );
  NAND U634 ( .A(n725), .B(n726), .Z(n724) );
  NANDN U635 ( .A(A[75]), .B(B[75]), .Z(n726) );
  AND U636 ( .A(n727), .B(n728), .Z(n725) );
  NANDN U637 ( .A(A[74]), .B(B[74]), .Z(n728) );
  NAND U638 ( .A(n729), .B(n730), .Z(n727) );
  NANDN U639 ( .A(B[74]), .B(A[74]), .Z(n730) );
  AND U640 ( .A(n731), .B(n732), .Z(n729) );
  NAND U641 ( .A(n733), .B(n734), .Z(n732) );
  NANDN U642 ( .A(A[73]), .B(B[73]), .Z(n734) );
  AND U643 ( .A(n735), .B(n736), .Z(n733) );
  NANDN U644 ( .A(A[72]), .B(B[72]), .Z(n736) );
  NAND U645 ( .A(n737), .B(n738), .Z(n735) );
  NANDN U646 ( .A(B[72]), .B(A[72]), .Z(n738) );
  AND U647 ( .A(n739), .B(n740), .Z(n737) );
  NAND U648 ( .A(n741), .B(n742), .Z(n740) );
  NANDN U649 ( .A(A[71]), .B(B[71]), .Z(n742) );
  AND U650 ( .A(n743), .B(n744), .Z(n741) );
  NANDN U651 ( .A(A[70]), .B(B[70]), .Z(n744) );
  NAND U652 ( .A(n745), .B(n746), .Z(n743) );
  NANDN U653 ( .A(B[70]), .B(A[70]), .Z(n746) );
  AND U654 ( .A(n747), .B(n748), .Z(n745) );
  NAND U655 ( .A(n749), .B(n750), .Z(n748) );
  NANDN U656 ( .A(A[69]), .B(B[69]), .Z(n750) );
  AND U657 ( .A(n751), .B(n752), .Z(n749) );
  NANDN U658 ( .A(A[68]), .B(B[68]), .Z(n752) );
  NAND U659 ( .A(n753), .B(n754), .Z(n751) );
  NANDN U660 ( .A(B[68]), .B(A[68]), .Z(n754) );
  AND U661 ( .A(n755), .B(n756), .Z(n753) );
  NAND U662 ( .A(n757), .B(n758), .Z(n756) );
  NANDN U663 ( .A(A[67]), .B(B[67]), .Z(n758) );
  AND U664 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U665 ( .A(A[66]), .B(B[66]), .Z(n760) );
  NAND U666 ( .A(n761), .B(n762), .Z(n759) );
  NANDN U667 ( .A(B[66]), .B(A[66]), .Z(n762) );
  AND U668 ( .A(n763), .B(n764), .Z(n761) );
  NAND U669 ( .A(n765), .B(n766), .Z(n764) );
  NANDN U670 ( .A(A[65]), .B(B[65]), .Z(n766) );
  AND U671 ( .A(n767), .B(n768), .Z(n765) );
  NANDN U672 ( .A(A[64]), .B(B[64]), .Z(n768) );
  NAND U673 ( .A(n769), .B(n770), .Z(n767) );
  NANDN U674 ( .A(B[64]), .B(A[64]), .Z(n770) );
  AND U675 ( .A(n771), .B(n772), .Z(n769) );
  NAND U676 ( .A(n773), .B(n774), .Z(n772) );
  NANDN U677 ( .A(A[63]), .B(B[63]), .Z(n774) );
  AND U678 ( .A(n775), .B(n776), .Z(n773) );
  NANDN U679 ( .A(A[62]), .B(B[62]), .Z(n776) );
  NAND U680 ( .A(n777), .B(n778), .Z(n775) );
  NANDN U681 ( .A(B[62]), .B(A[62]), .Z(n778) );
  AND U682 ( .A(n779), .B(n780), .Z(n777) );
  NAND U683 ( .A(n781), .B(n782), .Z(n780) );
  NANDN U684 ( .A(A[61]), .B(B[61]), .Z(n782) );
  AND U685 ( .A(n783), .B(n784), .Z(n781) );
  NANDN U686 ( .A(A[60]), .B(B[60]), .Z(n784) );
  NAND U687 ( .A(n785), .B(n786), .Z(n783) );
  NANDN U688 ( .A(B[60]), .B(A[60]), .Z(n786) );
  AND U689 ( .A(n787), .B(n788), .Z(n785) );
  NAND U690 ( .A(n789), .B(n790), .Z(n788) );
  NANDN U691 ( .A(A[59]), .B(B[59]), .Z(n790) );
  AND U692 ( .A(n791), .B(n792), .Z(n789) );
  NANDN U693 ( .A(A[58]), .B(B[58]), .Z(n792) );
  NAND U694 ( .A(n793), .B(n794), .Z(n791) );
  NANDN U695 ( .A(B[58]), .B(A[58]), .Z(n794) );
  AND U696 ( .A(n795), .B(n796), .Z(n793) );
  NAND U697 ( .A(n797), .B(n798), .Z(n796) );
  NANDN U698 ( .A(A[57]), .B(B[57]), .Z(n798) );
  AND U699 ( .A(n799), .B(n800), .Z(n797) );
  NANDN U700 ( .A(A[56]), .B(B[56]), .Z(n800) );
  NAND U701 ( .A(n801), .B(n802), .Z(n799) );
  NANDN U702 ( .A(B[56]), .B(A[56]), .Z(n802) );
  AND U703 ( .A(n803), .B(n804), .Z(n801) );
  NAND U704 ( .A(n805), .B(n806), .Z(n804) );
  NANDN U705 ( .A(A[55]), .B(B[55]), .Z(n806) );
  AND U706 ( .A(n807), .B(n808), .Z(n805) );
  NANDN U707 ( .A(A[54]), .B(B[54]), .Z(n808) );
  NAND U708 ( .A(n809), .B(n810), .Z(n807) );
  NANDN U709 ( .A(B[54]), .B(A[54]), .Z(n810) );
  AND U710 ( .A(n811), .B(n812), .Z(n809) );
  NAND U711 ( .A(n813), .B(n814), .Z(n812) );
  NANDN U712 ( .A(A[53]), .B(B[53]), .Z(n814) );
  AND U713 ( .A(n815), .B(n816), .Z(n813) );
  NANDN U714 ( .A(A[52]), .B(B[52]), .Z(n816) );
  NAND U715 ( .A(n817), .B(n818), .Z(n815) );
  NANDN U716 ( .A(B[52]), .B(A[52]), .Z(n818) );
  AND U717 ( .A(n819), .B(n820), .Z(n817) );
  NAND U718 ( .A(n821), .B(n822), .Z(n820) );
  NANDN U719 ( .A(A[51]), .B(B[51]), .Z(n822) );
  AND U720 ( .A(n823), .B(n824), .Z(n821) );
  NANDN U721 ( .A(A[50]), .B(B[50]), .Z(n824) );
  NAND U722 ( .A(n825), .B(n826), .Z(n823) );
  NANDN U723 ( .A(B[50]), .B(A[50]), .Z(n826) );
  AND U724 ( .A(n827), .B(n828), .Z(n825) );
  NAND U725 ( .A(n829), .B(n830), .Z(n828) );
  NANDN U726 ( .A(A[49]), .B(B[49]), .Z(n830) );
  AND U727 ( .A(n831), .B(n832), .Z(n829) );
  NANDN U728 ( .A(A[48]), .B(B[48]), .Z(n832) );
  NAND U729 ( .A(n833), .B(n834), .Z(n831) );
  NANDN U730 ( .A(B[48]), .B(A[48]), .Z(n834) );
  AND U731 ( .A(n835), .B(n836), .Z(n833) );
  NAND U732 ( .A(n837), .B(n838), .Z(n836) );
  NANDN U733 ( .A(A[47]), .B(B[47]), .Z(n838) );
  AND U734 ( .A(n839), .B(n840), .Z(n837) );
  NANDN U735 ( .A(A[46]), .B(B[46]), .Z(n840) );
  NAND U736 ( .A(n841), .B(n842), .Z(n839) );
  NANDN U737 ( .A(B[46]), .B(A[46]), .Z(n842) );
  AND U738 ( .A(n843), .B(n844), .Z(n841) );
  NAND U739 ( .A(n845), .B(n846), .Z(n844) );
  NANDN U740 ( .A(A[45]), .B(B[45]), .Z(n846) );
  AND U741 ( .A(n847), .B(n848), .Z(n845) );
  NANDN U742 ( .A(A[44]), .B(B[44]), .Z(n848) );
  NAND U743 ( .A(n849), .B(n850), .Z(n847) );
  NANDN U744 ( .A(B[44]), .B(A[44]), .Z(n850) );
  AND U745 ( .A(n851), .B(n852), .Z(n849) );
  NAND U746 ( .A(n853), .B(n854), .Z(n852) );
  NANDN U747 ( .A(A[43]), .B(B[43]), .Z(n854) );
  AND U748 ( .A(n855), .B(n856), .Z(n853) );
  NANDN U749 ( .A(A[42]), .B(B[42]), .Z(n856) );
  NAND U750 ( .A(n857), .B(n858), .Z(n855) );
  NANDN U751 ( .A(B[42]), .B(A[42]), .Z(n858) );
  AND U752 ( .A(n859), .B(n860), .Z(n857) );
  NAND U753 ( .A(n861), .B(n862), .Z(n860) );
  NANDN U754 ( .A(A[41]), .B(B[41]), .Z(n862) );
  AND U755 ( .A(n863), .B(n864), .Z(n861) );
  NANDN U756 ( .A(A[40]), .B(B[40]), .Z(n864) );
  NAND U757 ( .A(n865), .B(n866), .Z(n863) );
  NANDN U758 ( .A(B[40]), .B(A[40]), .Z(n866) );
  AND U759 ( .A(n867), .B(n868), .Z(n865) );
  NAND U760 ( .A(n869), .B(n870), .Z(n868) );
  NANDN U761 ( .A(A[39]), .B(B[39]), .Z(n870) );
  AND U762 ( .A(n871), .B(n872), .Z(n869) );
  NANDN U763 ( .A(A[38]), .B(B[38]), .Z(n872) );
  NAND U764 ( .A(n873), .B(n874), .Z(n871) );
  NANDN U765 ( .A(B[38]), .B(A[38]), .Z(n874) );
  AND U766 ( .A(n875), .B(n876), .Z(n873) );
  NAND U767 ( .A(n877), .B(n878), .Z(n876) );
  NANDN U768 ( .A(A[37]), .B(B[37]), .Z(n878) );
  AND U769 ( .A(n879), .B(n880), .Z(n877) );
  NANDN U770 ( .A(A[36]), .B(B[36]), .Z(n880) );
  NAND U771 ( .A(n881), .B(n882), .Z(n879) );
  NANDN U772 ( .A(B[36]), .B(A[36]), .Z(n882) );
  AND U773 ( .A(n883), .B(n884), .Z(n881) );
  NAND U774 ( .A(n885), .B(n886), .Z(n884) );
  NANDN U775 ( .A(A[35]), .B(B[35]), .Z(n886) );
  AND U776 ( .A(n887), .B(n888), .Z(n885) );
  NANDN U777 ( .A(A[34]), .B(B[34]), .Z(n888) );
  NAND U778 ( .A(n889), .B(n890), .Z(n887) );
  NANDN U779 ( .A(B[34]), .B(A[34]), .Z(n890) );
  AND U780 ( .A(n891), .B(n892), .Z(n889) );
  NAND U781 ( .A(n893), .B(n894), .Z(n892) );
  NANDN U782 ( .A(A[33]), .B(B[33]), .Z(n894) );
  AND U783 ( .A(n895), .B(n896), .Z(n893) );
  NANDN U784 ( .A(A[32]), .B(B[32]), .Z(n896) );
  NAND U785 ( .A(n897), .B(n898), .Z(n895) );
  NANDN U786 ( .A(B[32]), .B(A[32]), .Z(n898) );
  AND U787 ( .A(n899), .B(n900), .Z(n897) );
  NAND U788 ( .A(n901), .B(n902), .Z(n900) );
  NANDN U789 ( .A(A[31]), .B(B[31]), .Z(n902) );
  AND U790 ( .A(n903), .B(n904), .Z(n901) );
  NANDN U791 ( .A(A[30]), .B(B[30]), .Z(n904) );
  NAND U792 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U793 ( .A(B[30]), .B(A[30]), .Z(n906) );
  AND U794 ( .A(n907), .B(n908), .Z(n905) );
  NAND U795 ( .A(n909), .B(n910), .Z(n908) );
  NANDN U796 ( .A(A[29]), .B(B[29]), .Z(n910) );
  AND U797 ( .A(n911), .B(n912), .Z(n909) );
  NANDN U798 ( .A(A[28]), .B(B[28]), .Z(n912) );
  NAND U799 ( .A(n913), .B(n914), .Z(n911) );
  NANDN U800 ( .A(B[28]), .B(A[28]), .Z(n914) );
  AND U801 ( .A(n915), .B(n916), .Z(n913) );
  NAND U802 ( .A(n917), .B(n918), .Z(n916) );
  NANDN U803 ( .A(A[27]), .B(B[27]), .Z(n918) );
  AND U804 ( .A(n919), .B(n920), .Z(n917) );
  NANDN U805 ( .A(A[26]), .B(B[26]), .Z(n920) );
  NAND U806 ( .A(n921), .B(n922), .Z(n919) );
  NANDN U807 ( .A(B[26]), .B(A[26]), .Z(n922) );
  AND U808 ( .A(n923), .B(n924), .Z(n921) );
  NAND U809 ( .A(n925), .B(n926), .Z(n924) );
  NANDN U810 ( .A(A[25]), .B(B[25]), .Z(n926) );
  AND U811 ( .A(n927), .B(n928), .Z(n925) );
  NANDN U812 ( .A(A[24]), .B(B[24]), .Z(n928) );
  NAND U813 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U814 ( .A(B[24]), .B(A[24]), .Z(n930) );
  AND U815 ( .A(n931), .B(n932), .Z(n929) );
  NAND U816 ( .A(n933), .B(n934), .Z(n932) );
  NANDN U817 ( .A(A[23]), .B(B[23]), .Z(n934) );
  AND U818 ( .A(n935), .B(n936), .Z(n933) );
  NANDN U819 ( .A(A[22]), .B(B[22]), .Z(n936) );
  NAND U820 ( .A(n937), .B(n938), .Z(n935) );
  NANDN U821 ( .A(B[22]), .B(A[22]), .Z(n938) );
  AND U822 ( .A(n939), .B(n940), .Z(n937) );
  NAND U823 ( .A(n941), .B(n942), .Z(n940) );
  NANDN U824 ( .A(A[21]), .B(B[21]), .Z(n942) );
  AND U825 ( .A(n943), .B(n944), .Z(n941) );
  NANDN U826 ( .A(A[20]), .B(B[20]), .Z(n944) );
  NAND U827 ( .A(n945), .B(n946), .Z(n943) );
  NANDN U828 ( .A(B[20]), .B(A[20]), .Z(n946) );
  AND U829 ( .A(n947), .B(n948), .Z(n945) );
  NAND U830 ( .A(n949), .B(n950), .Z(n948) );
  NANDN U831 ( .A(A[19]), .B(B[19]), .Z(n950) );
  AND U832 ( .A(n951), .B(n952), .Z(n949) );
  NANDN U833 ( .A(A[18]), .B(B[18]), .Z(n952) );
  NAND U834 ( .A(n953), .B(n954), .Z(n951) );
  NANDN U835 ( .A(B[18]), .B(A[18]), .Z(n954) );
  AND U836 ( .A(n955), .B(n956), .Z(n953) );
  NAND U837 ( .A(n957), .B(n958), .Z(n956) );
  NANDN U838 ( .A(A[17]), .B(B[17]), .Z(n958) );
  AND U839 ( .A(n959), .B(n960), .Z(n957) );
  NANDN U840 ( .A(A[16]), .B(B[16]), .Z(n960) );
  NAND U841 ( .A(n961), .B(n962), .Z(n959) );
  NANDN U842 ( .A(B[16]), .B(A[16]), .Z(n962) );
  AND U843 ( .A(n963), .B(n964), .Z(n961) );
  NAND U844 ( .A(n965), .B(n966), .Z(n964) );
  NANDN U845 ( .A(A[15]), .B(B[15]), .Z(n966) );
  AND U846 ( .A(n967), .B(n968), .Z(n965) );
  NANDN U847 ( .A(A[14]), .B(B[14]), .Z(n968) );
  NAND U848 ( .A(n969), .B(n970), .Z(n967) );
  NANDN U849 ( .A(B[14]), .B(A[14]), .Z(n970) );
  AND U850 ( .A(n971), .B(n972), .Z(n969) );
  NAND U851 ( .A(n973), .B(n974), .Z(n972) );
  NANDN U852 ( .A(A[13]), .B(B[13]), .Z(n974) );
  AND U853 ( .A(n975), .B(n976), .Z(n973) );
  NANDN U854 ( .A(A[12]), .B(B[12]), .Z(n976) );
  NAND U855 ( .A(n977), .B(n978), .Z(n975) );
  NANDN U856 ( .A(B[12]), .B(A[12]), .Z(n978) );
  AND U857 ( .A(n979), .B(n980), .Z(n977) );
  NAND U858 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U859 ( .A(A[11]), .B(B[11]), .Z(n982) );
  AND U860 ( .A(n983), .B(n984), .Z(n981) );
  NANDN U861 ( .A(A[10]), .B(B[10]), .Z(n984) );
  NAND U862 ( .A(n985), .B(n986), .Z(n983) );
  NANDN U863 ( .A(B[9]), .B(A[9]), .Z(n986) );
  AND U864 ( .A(n987), .B(n988), .Z(n985) );
  NAND U865 ( .A(n989), .B(n990), .Z(n988) );
  NANDN U866 ( .A(A[9]), .B(B[9]), .Z(n990) );
  AND U867 ( .A(n991), .B(n992), .Z(n989) );
  NANDN U868 ( .A(A[8]), .B(B[8]), .Z(n992) );
  NAND U869 ( .A(n993), .B(n994), .Z(n991) );
  NANDN U870 ( .A(B[8]), .B(A[8]), .Z(n994) );
  AND U871 ( .A(n995), .B(n996), .Z(n993) );
  NAND U872 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U873 ( .A(A[7]), .B(B[7]), .Z(n998) );
  AND U874 ( .A(n999), .B(n1000), .Z(n997) );
  NANDN U875 ( .A(A[6]), .B(B[6]), .Z(n1000) );
  NAND U876 ( .A(n1001), .B(n1002), .Z(n999) );
  NANDN U877 ( .A(B[6]), .B(A[6]), .Z(n1002) );
  AND U878 ( .A(n1003), .B(n1004), .Z(n1001) );
  NAND U879 ( .A(n1005), .B(n1006), .Z(n1004) );
  NANDN U880 ( .A(A[5]), .B(B[5]), .Z(n1006) );
  AND U881 ( .A(n1007), .B(n1008), .Z(n1005) );
  NANDN U882 ( .A(A[4]), .B(B[4]), .Z(n1008) );
  NAND U883 ( .A(n1009), .B(n1010), .Z(n1007) );
  NANDN U884 ( .A(B[4]), .B(A[4]), .Z(n1010) );
  AND U885 ( .A(n1011), .B(n1012), .Z(n1009) );
  NAND U886 ( .A(n1013), .B(n1014), .Z(n1012) );
  NANDN U887 ( .A(A[3]), .B(B[3]), .Z(n1014) );
  AND U888 ( .A(n1015), .B(n1016), .Z(n1013) );
  NANDN U889 ( .A(A[2]), .B(B[2]), .Z(n1016) );
  NAND U890 ( .A(n1017), .B(n1018), .Z(n1015) );
  NANDN U891 ( .A(B[2]), .B(A[2]), .Z(n1018) );
  AND U892 ( .A(n1019), .B(n1020), .Z(n1017) );
  NAND U893 ( .A(n1021), .B(A[0]), .Z(n1020) );
  ANDN U894 ( .B(n1022), .A(B[0]), .Z(n1021) );
  NANDN U895 ( .A(A[1]), .B(B[1]), .Z(n1022) );
  NANDN U896 ( .A(B[1]), .B(A[1]), .Z(n1019) );
  NANDN U897 ( .A(B[3]), .B(A[3]), .Z(n1011) );
  NANDN U898 ( .A(B[5]), .B(A[5]), .Z(n1003) );
  NANDN U899 ( .A(B[7]), .B(A[7]), .Z(n995) );
  NANDN U900 ( .A(B[10]), .B(A[10]), .Z(n987) );
  NANDN U901 ( .A(B[11]), .B(A[11]), .Z(n979) );
  NANDN U902 ( .A(B[13]), .B(A[13]), .Z(n971) );
  NANDN U903 ( .A(B[15]), .B(A[15]), .Z(n963) );
  NANDN U904 ( .A(B[17]), .B(A[17]), .Z(n955) );
  NANDN U905 ( .A(B[19]), .B(A[19]), .Z(n947) );
  NANDN U906 ( .A(B[21]), .B(A[21]), .Z(n939) );
  NANDN U907 ( .A(B[23]), .B(A[23]), .Z(n931) );
  NANDN U908 ( .A(B[25]), .B(A[25]), .Z(n923) );
  NANDN U909 ( .A(B[27]), .B(A[27]), .Z(n915) );
  NANDN U910 ( .A(B[29]), .B(A[29]), .Z(n907) );
  NANDN U911 ( .A(B[31]), .B(A[31]), .Z(n899) );
  NANDN U912 ( .A(B[33]), .B(A[33]), .Z(n891) );
  NANDN U913 ( .A(B[35]), .B(A[35]), .Z(n883) );
  NANDN U914 ( .A(B[37]), .B(A[37]), .Z(n875) );
  NANDN U915 ( .A(B[39]), .B(A[39]), .Z(n867) );
  NANDN U916 ( .A(B[41]), .B(A[41]), .Z(n859) );
  NANDN U917 ( .A(B[43]), .B(A[43]), .Z(n851) );
  NANDN U918 ( .A(B[45]), .B(A[45]), .Z(n843) );
  NANDN U919 ( .A(B[47]), .B(A[47]), .Z(n835) );
  NANDN U920 ( .A(B[49]), .B(A[49]), .Z(n827) );
  NANDN U921 ( .A(B[51]), .B(A[51]), .Z(n819) );
  NANDN U922 ( .A(B[53]), .B(A[53]), .Z(n811) );
  NANDN U923 ( .A(B[55]), .B(A[55]), .Z(n803) );
  NANDN U924 ( .A(B[57]), .B(A[57]), .Z(n795) );
  NANDN U925 ( .A(B[59]), .B(A[59]), .Z(n787) );
  NANDN U926 ( .A(B[61]), .B(A[61]), .Z(n779) );
  NANDN U927 ( .A(B[63]), .B(A[63]), .Z(n771) );
  NANDN U928 ( .A(B[65]), .B(A[65]), .Z(n763) );
  NANDN U929 ( .A(B[67]), .B(A[67]), .Z(n755) );
  NANDN U930 ( .A(B[69]), .B(A[69]), .Z(n747) );
  NANDN U931 ( .A(B[71]), .B(A[71]), .Z(n739) );
  NANDN U932 ( .A(B[73]), .B(A[73]), .Z(n731) );
  NANDN U933 ( .A(B[75]), .B(A[75]), .Z(n723) );
  NANDN U934 ( .A(B[77]), .B(A[77]), .Z(n715) );
  NANDN U935 ( .A(B[79]), .B(A[79]), .Z(n707) );
  NANDN U936 ( .A(B[81]), .B(A[81]), .Z(n699) );
  NANDN U937 ( .A(B[83]), .B(A[83]), .Z(n691) );
  NANDN U938 ( .A(B[85]), .B(A[85]), .Z(n683) );
  NANDN U939 ( .A(B[87]), .B(A[87]), .Z(n675) );
  NANDN U940 ( .A(B[89]), .B(A[89]), .Z(n667) );
  NANDN U941 ( .A(B[91]), .B(A[91]), .Z(n659) );
  NANDN U942 ( .A(B[93]), .B(A[93]), .Z(n651) );
  NANDN U943 ( .A(B[95]), .B(A[95]), .Z(n643) );
  NANDN U944 ( .A(B[97]), .B(A[97]), .Z(n635) );
  NANDN U945 ( .A(B[100]), .B(A[100]), .Z(n627) );
  NANDN U946 ( .A(B[101]), .B(A[101]), .Z(n619) );
  NANDN U947 ( .A(B[103]), .B(A[103]), .Z(n611) );
  NANDN U948 ( .A(B[105]), .B(A[105]), .Z(n603) );
  NANDN U949 ( .A(B[107]), .B(A[107]), .Z(n595) );
  NANDN U950 ( .A(B[109]), .B(A[109]), .Z(n587) );
  NANDN U951 ( .A(B[111]), .B(A[111]), .Z(n579) );
  NANDN U952 ( .A(B[113]), .B(A[113]), .Z(n571) );
  NANDN U953 ( .A(B[115]), .B(A[115]), .Z(n563) );
  NANDN U954 ( .A(B[117]), .B(A[117]), .Z(n555) );
  NANDN U955 ( .A(B[119]), .B(A[119]), .Z(n547) );
  NANDN U956 ( .A(B[121]), .B(A[121]), .Z(n539) );
  NANDN U957 ( .A(B[123]), .B(A[123]), .Z(n531) );
  NANDN U958 ( .A(B[125]), .B(A[125]), .Z(n523) );
  NANDN U959 ( .A(B[127]), .B(A[127]), .Z(n515) );
  NANDN U960 ( .A(B[129]), .B(A[129]), .Z(n507) );
  NANDN U961 ( .A(B[131]), .B(A[131]), .Z(n499) );
  NANDN U962 ( .A(B[133]), .B(A[133]), .Z(n491) );
  NANDN U963 ( .A(B[135]), .B(A[135]), .Z(n483) );
  NANDN U964 ( .A(B[137]), .B(A[137]), .Z(n475) );
  NANDN U965 ( .A(B[139]), .B(A[139]), .Z(n467) );
  NANDN U966 ( .A(B[141]), .B(A[141]), .Z(n459) );
  NANDN U967 ( .A(B[143]), .B(A[143]), .Z(n451) );
  NANDN U968 ( .A(B[145]), .B(A[145]), .Z(n443) );
  NANDN U969 ( .A(B[147]), .B(A[147]), .Z(n435) );
  NANDN U970 ( .A(B[149]), .B(A[149]), .Z(n427) );
  NANDN U971 ( .A(B[151]), .B(A[151]), .Z(n419) );
  NANDN U972 ( .A(B[153]), .B(A[153]), .Z(n411) );
  NANDN U973 ( .A(B[155]), .B(A[155]), .Z(n403) );
  NANDN U974 ( .A(B[157]), .B(A[157]), .Z(n395) );
  NANDN U975 ( .A(B[159]), .B(A[159]), .Z(n387) );
  NANDN U976 ( .A(B[161]), .B(A[161]), .Z(n379) );
  NANDN U977 ( .A(B[163]), .B(A[163]), .Z(n371) );
  NANDN U978 ( .A(B[165]), .B(A[165]), .Z(n363) );
  NANDN U979 ( .A(B[167]), .B(A[167]), .Z(n355) );
  NANDN U980 ( .A(B[169]), .B(A[169]), .Z(n347) );
  NANDN U981 ( .A(B[171]), .B(A[171]), .Z(n339) );
  NANDN U982 ( .A(B[173]), .B(A[173]), .Z(n331) );
  NANDN U983 ( .A(B[175]), .B(A[175]), .Z(n323) );
  NANDN U984 ( .A(B[177]), .B(A[177]), .Z(n315) );
  NANDN U985 ( .A(B[179]), .B(A[179]), .Z(n307) );
  NANDN U986 ( .A(B[181]), .B(A[181]), .Z(n299) );
  NANDN U987 ( .A(B[183]), .B(A[183]), .Z(n291) );
  NANDN U988 ( .A(B[185]), .B(A[185]), .Z(n283) );
  NANDN U989 ( .A(B[187]), .B(A[187]), .Z(n275) );
  NANDN U990 ( .A(B[189]), .B(A[189]), .Z(n267) );
  NANDN U991 ( .A(B[191]), .B(A[191]), .Z(n259) );
  NANDN U992 ( .A(B[193]), .B(A[193]), .Z(n251) );
  NANDN U993 ( .A(B[195]), .B(A[195]), .Z(n243) );
  NANDN U994 ( .A(B[197]), .B(A[197]), .Z(n235) );
  NANDN U995 ( .A(B[199]), .B(A[199]), .Z(n227) );
  NANDN U996 ( .A(B[201]), .B(A[201]), .Z(n219) );
  NANDN U997 ( .A(B[203]), .B(A[203]), .Z(n211) );
  NANDN U998 ( .A(B[205]), .B(A[205]), .Z(n203) );
  NANDN U999 ( .A(B[207]), .B(A[207]), .Z(n195) );
  NANDN U1000 ( .A(B[209]), .B(A[209]), .Z(n187) );
  NANDN U1001 ( .A(B[211]), .B(A[211]), .Z(n179) );
  NANDN U1002 ( .A(B[213]), .B(A[213]), .Z(n171) );
  NANDN U1003 ( .A(B[215]), .B(A[215]), .Z(n163) );
  NANDN U1004 ( .A(B[217]), .B(A[217]), .Z(n155) );
  NANDN U1005 ( .A(B[219]), .B(A[219]), .Z(n147) );
  NANDN U1006 ( .A(B[221]), .B(A[221]), .Z(n139) );
  NANDN U1007 ( .A(B[223]), .B(A[223]), .Z(n131) );
  NANDN U1008 ( .A(B[225]), .B(A[225]), .Z(n123) );
  NANDN U1009 ( .A(B[227]), .B(A[227]), .Z(n115) );
  NANDN U1010 ( .A(B[229]), .B(A[229]), .Z(n107) );
  NANDN U1011 ( .A(B[231]), .B(A[231]), .Z(n99) );
  NANDN U1012 ( .A(B[233]), .B(A[233]), .Z(n91) );
  NANDN U1013 ( .A(B[235]), .B(A[235]), .Z(n83) );
  NANDN U1014 ( .A(B[237]), .B(A[237]), .Z(n75) );
  NANDN U1015 ( .A(B[239]), .B(A[239]), .Z(n67) );
  NANDN U1016 ( .A(B[241]), .B(A[241]), .Z(n59) );
  NANDN U1017 ( .A(B[243]), .B(A[243]), .Z(n51) );
  NANDN U1018 ( .A(B[245]), .B(A[245]), .Z(n43) );
  NANDN U1019 ( .A(B[247]), .B(A[247]), .Z(n35) );
  NANDN U1020 ( .A(B[249]), .B(A[249]), .Z(n27) );
  NANDN U1021 ( .A(B[251]), .B(A[251]), .Z(n19) );
  NANDN U1022 ( .A(B[253]), .B(A[253]), .Z(n11) );
  NANDN U1023 ( .A(A[255]), .B(B[255]), .Z(n3) );
endmodule


module modmult_step_N256_2_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280;

  IV U1 ( .A(A[1]), .Z(n1) );
  IV U2 ( .A(n1279), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(DIFF[9]) );
  XOR U4 ( .A(B[9]), .B(A[9]), .Z(n4) );
  XNOR U5 ( .A(n5), .B(n6), .Z(DIFF[99]) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(DIFF[98]) );
  XOR U8 ( .A(B[98]), .B(A[98]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(DIFF[97]) );
  XOR U10 ( .A(B[97]), .B(A[97]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(DIFF[96]) );
  XOR U12 ( .A(B[96]), .B(A[96]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(DIFF[95]) );
  XOR U14 ( .A(B[95]), .B(A[95]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(DIFF[94]) );
  XOR U16 ( .A(B[94]), .B(A[94]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(DIFF[93]) );
  XOR U18 ( .A(B[93]), .B(A[93]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(DIFF[92]) );
  XOR U20 ( .A(B[92]), .B(A[92]), .Z(n20) );
  XOR U21 ( .A(n21), .B(n22), .Z(DIFF[91]) );
  XOR U22 ( .A(B[91]), .B(A[91]), .Z(n22) );
  XOR U23 ( .A(n23), .B(n24), .Z(DIFF[90]) );
  XOR U24 ( .A(B[90]), .B(A[90]), .Z(n24) );
  XOR U25 ( .A(n25), .B(n26), .Z(DIFF[8]) );
  XOR U26 ( .A(B[8]), .B(A[8]), .Z(n26) );
  XOR U27 ( .A(n27), .B(n28), .Z(DIFF[89]) );
  XOR U28 ( .A(B[89]), .B(A[89]), .Z(n28) );
  XOR U29 ( .A(n29), .B(n30), .Z(DIFF[88]) );
  XOR U30 ( .A(B[88]), .B(A[88]), .Z(n30) );
  XOR U31 ( .A(n31), .B(n32), .Z(DIFF[87]) );
  XOR U32 ( .A(B[87]), .B(A[87]), .Z(n32) );
  XOR U33 ( .A(n33), .B(n34), .Z(DIFF[86]) );
  XOR U34 ( .A(B[86]), .B(A[86]), .Z(n34) );
  XOR U35 ( .A(n35), .B(n36), .Z(DIFF[85]) );
  XOR U36 ( .A(B[85]), .B(A[85]), .Z(n36) );
  XOR U37 ( .A(n37), .B(n38), .Z(DIFF[84]) );
  XOR U38 ( .A(B[84]), .B(A[84]), .Z(n38) );
  XOR U39 ( .A(n39), .B(n40), .Z(DIFF[83]) );
  XOR U40 ( .A(B[83]), .B(A[83]), .Z(n40) );
  XOR U41 ( .A(n41), .B(n42), .Z(DIFF[82]) );
  XOR U42 ( .A(B[82]), .B(A[82]), .Z(n42) );
  XOR U43 ( .A(n43), .B(n44), .Z(DIFF[81]) );
  XOR U44 ( .A(B[81]), .B(A[81]), .Z(n44) );
  XOR U45 ( .A(n45), .B(n46), .Z(DIFF[80]) );
  XOR U46 ( .A(B[80]), .B(A[80]), .Z(n46) );
  XOR U47 ( .A(n47), .B(n48), .Z(DIFF[7]) );
  XOR U48 ( .A(B[7]), .B(A[7]), .Z(n48) );
  XOR U49 ( .A(n49), .B(n50), .Z(DIFF[79]) );
  XOR U50 ( .A(B[79]), .B(A[79]), .Z(n50) );
  XOR U51 ( .A(n51), .B(n52), .Z(DIFF[78]) );
  XOR U52 ( .A(B[78]), .B(A[78]), .Z(n52) );
  XOR U53 ( .A(n53), .B(n54), .Z(DIFF[77]) );
  XOR U54 ( .A(B[77]), .B(A[77]), .Z(n54) );
  XOR U55 ( .A(n55), .B(n56), .Z(DIFF[76]) );
  XOR U56 ( .A(B[76]), .B(A[76]), .Z(n56) );
  XOR U57 ( .A(n57), .B(n58), .Z(DIFF[75]) );
  XOR U58 ( .A(B[75]), .B(A[75]), .Z(n58) );
  XOR U59 ( .A(n59), .B(n60), .Z(DIFF[74]) );
  XOR U60 ( .A(B[74]), .B(A[74]), .Z(n60) );
  XOR U61 ( .A(n61), .B(n62), .Z(DIFF[73]) );
  XOR U62 ( .A(B[73]), .B(A[73]), .Z(n62) );
  XOR U63 ( .A(n63), .B(n64), .Z(DIFF[72]) );
  XOR U64 ( .A(B[72]), .B(A[72]), .Z(n64) );
  XOR U65 ( .A(n65), .B(n66), .Z(DIFF[71]) );
  XOR U66 ( .A(B[71]), .B(A[71]), .Z(n66) );
  XOR U67 ( .A(n67), .B(n68), .Z(DIFF[70]) );
  XOR U68 ( .A(B[70]), .B(A[70]), .Z(n68) );
  XOR U69 ( .A(n69), .B(n70), .Z(DIFF[6]) );
  XOR U70 ( .A(B[6]), .B(A[6]), .Z(n70) );
  XOR U71 ( .A(n71), .B(n72), .Z(DIFF[69]) );
  XOR U72 ( .A(B[69]), .B(A[69]), .Z(n72) );
  XOR U73 ( .A(n73), .B(n74), .Z(DIFF[68]) );
  XOR U74 ( .A(B[68]), .B(A[68]), .Z(n74) );
  XOR U75 ( .A(n75), .B(n76), .Z(DIFF[67]) );
  XOR U76 ( .A(B[67]), .B(A[67]), .Z(n76) );
  XOR U77 ( .A(n77), .B(n78), .Z(DIFF[66]) );
  XOR U78 ( .A(B[66]), .B(A[66]), .Z(n78) );
  XOR U79 ( .A(n79), .B(n80), .Z(DIFF[65]) );
  XOR U80 ( .A(B[65]), .B(A[65]), .Z(n80) );
  XOR U81 ( .A(n81), .B(n82), .Z(DIFF[64]) );
  XOR U82 ( .A(B[64]), .B(A[64]), .Z(n82) );
  XOR U83 ( .A(n83), .B(n84), .Z(DIFF[63]) );
  XOR U84 ( .A(B[63]), .B(A[63]), .Z(n84) );
  XOR U85 ( .A(n85), .B(n86), .Z(DIFF[62]) );
  XOR U86 ( .A(B[62]), .B(A[62]), .Z(n86) );
  XOR U87 ( .A(n87), .B(n88), .Z(DIFF[61]) );
  XOR U88 ( .A(B[61]), .B(A[61]), .Z(n88) );
  XOR U89 ( .A(n89), .B(n90), .Z(DIFF[60]) );
  XOR U90 ( .A(B[60]), .B(A[60]), .Z(n90) );
  XOR U91 ( .A(n91), .B(n92), .Z(DIFF[5]) );
  XOR U92 ( .A(B[5]), .B(A[5]), .Z(n92) );
  XOR U93 ( .A(n93), .B(n94), .Z(DIFF[59]) );
  XOR U94 ( .A(B[59]), .B(A[59]), .Z(n94) );
  XOR U95 ( .A(n95), .B(n96), .Z(DIFF[58]) );
  XOR U96 ( .A(B[58]), .B(A[58]), .Z(n96) );
  XOR U97 ( .A(n97), .B(n98), .Z(DIFF[57]) );
  XOR U98 ( .A(B[57]), .B(A[57]), .Z(n98) );
  XOR U99 ( .A(n99), .B(n100), .Z(DIFF[56]) );
  XOR U100 ( .A(B[56]), .B(A[56]), .Z(n100) );
  XOR U101 ( .A(n101), .B(n102), .Z(DIFF[55]) );
  XOR U102 ( .A(B[55]), .B(A[55]), .Z(n102) );
  XOR U103 ( .A(n103), .B(n104), .Z(DIFF[54]) );
  XOR U104 ( .A(B[54]), .B(A[54]), .Z(n104) );
  XOR U105 ( .A(n105), .B(n106), .Z(DIFF[53]) );
  XOR U106 ( .A(B[53]), .B(A[53]), .Z(n106) );
  XOR U107 ( .A(n107), .B(n108), .Z(DIFF[52]) );
  XOR U108 ( .A(B[52]), .B(A[52]), .Z(n108) );
  XOR U109 ( .A(n109), .B(n110), .Z(DIFF[51]) );
  XOR U110 ( .A(B[51]), .B(A[51]), .Z(n110) );
  XOR U111 ( .A(n111), .B(n112), .Z(DIFF[50]) );
  XOR U112 ( .A(B[50]), .B(A[50]), .Z(n112) );
  XOR U113 ( .A(n113), .B(n114), .Z(DIFF[4]) );
  XOR U114 ( .A(B[4]), .B(A[4]), .Z(n114) );
  XOR U115 ( .A(n115), .B(n116), .Z(DIFF[49]) );
  XOR U116 ( .A(B[49]), .B(A[49]), .Z(n116) );
  XOR U117 ( .A(n117), .B(n118), .Z(DIFF[48]) );
  XOR U118 ( .A(B[48]), .B(A[48]), .Z(n118) );
  XOR U119 ( .A(n119), .B(n120), .Z(DIFF[47]) );
  XOR U120 ( .A(B[47]), .B(A[47]), .Z(n120) );
  XOR U121 ( .A(n121), .B(n122), .Z(DIFF[46]) );
  XOR U122 ( .A(B[46]), .B(A[46]), .Z(n122) );
  XOR U123 ( .A(n123), .B(n124), .Z(DIFF[45]) );
  XOR U124 ( .A(B[45]), .B(A[45]), .Z(n124) );
  XOR U125 ( .A(n125), .B(n126), .Z(DIFF[44]) );
  XOR U126 ( .A(B[44]), .B(A[44]), .Z(n126) );
  XOR U127 ( .A(n127), .B(n128), .Z(DIFF[43]) );
  XOR U128 ( .A(B[43]), .B(A[43]), .Z(n128) );
  XOR U129 ( .A(n129), .B(n130), .Z(DIFF[42]) );
  XOR U130 ( .A(B[42]), .B(A[42]), .Z(n130) );
  XOR U131 ( .A(n131), .B(n132), .Z(DIFF[41]) );
  XOR U132 ( .A(B[41]), .B(A[41]), .Z(n132) );
  XOR U133 ( .A(n133), .B(n134), .Z(DIFF[40]) );
  XOR U134 ( .A(B[40]), .B(A[40]), .Z(n134) );
  XOR U135 ( .A(n135), .B(n136), .Z(DIFF[3]) );
  XOR U136 ( .A(B[3]), .B(A[3]), .Z(n136) );
  XOR U137 ( .A(n137), .B(n138), .Z(DIFF[39]) );
  XOR U138 ( .A(B[39]), .B(A[39]), .Z(n138) );
  XOR U139 ( .A(n139), .B(n140), .Z(DIFF[38]) );
  XOR U140 ( .A(B[38]), .B(A[38]), .Z(n140) );
  XOR U141 ( .A(n141), .B(n142), .Z(DIFF[37]) );
  XOR U142 ( .A(B[37]), .B(A[37]), .Z(n142) );
  XOR U143 ( .A(n143), .B(n144), .Z(DIFF[36]) );
  XOR U144 ( .A(B[36]), .B(A[36]), .Z(n144) );
  XOR U145 ( .A(n145), .B(n146), .Z(DIFF[35]) );
  XOR U146 ( .A(B[35]), .B(A[35]), .Z(n146) );
  XOR U147 ( .A(n147), .B(n148), .Z(DIFF[34]) );
  XOR U148 ( .A(B[34]), .B(A[34]), .Z(n148) );
  XOR U149 ( .A(n149), .B(n150), .Z(DIFF[33]) );
  XOR U150 ( .A(B[33]), .B(A[33]), .Z(n150) );
  XOR U151 ( .A(n151), .B(n152), .Z(DIFF[32]) );
  XOR U152 ( .A(B[32]), .B(A[32]), .Z(n152) );
  XOR U153 ( .A(n153), .B(n154), .Z(DIFF[31]) );
  XOR U154 ( .A(B[31]), .B(A[31]), .Z(n154) );
  XOR U155 ( .A(n155), .B(n156), .Z(DIFF[30]) );
  XOR U156 ( .A(B[30]), .B(A[30]), .Z(n156) );
  XOR U157 ( .A(n157), .B(n158), .Z(DIFF[2]) );
  XOR U158 ( .A(B[2]), .B(A[2]), .Z(n158) );
  XOR U159 ( .A(n159), .B(n160), .Z(DIFF[29]) );
  XOR U160 ( .A(B[29]), .B(A[29]), .Z(n160) );
  XOR U161 ( .A(n161), .B(n162), .Z(DIFF[28]) );
  XOR U162 ( .A(B[28]), .B(A[28]), .Z(n162) );
  XOR U163 ( .A(n163), .B(n164), .Z(DIFF[27]) );
  XOR U164 ( .A(B[27]), .B(A[27]), .Z(n164) );
  XOR U165 ( .A(n165), .B(n166), .Z(DIFF[26]) );
  XOR U166 ( .A(B[26]), .B(A[26]), .Z(n166) );
  XOR U167 ( .A(n167), .B(n168), .Z(DIFF[25]) );
  XOR U168 ( .A(B[25]), .B(A[25]), .Z(n168) );
  XOR U169 ( .A(A[257]), .B(n169), .Z(DIFF[257]) );
  ANDN U170 ( .B(n170), .A(A[256]), .Z(n169) );
  XOR U171 ( .A(A[256]), .B(n170), .Z(DIFF[256]) );
  AND U172 ( .A(n171), .B(n172), .Z(n170) );
  NANDN U173 ( .A(B[255]), .B(n173), .Z(n172) );
  NANDN U174 ( .A(A[255]), .B(n174), .Z(n173) );
  NANDN U175 ( .A(n174), .B(A[255]), .Z(n171) );
  XOR U176 ( .A(n174), .B(n175), .Z(DIFF[255]) );
  XOR U177 ( .A(B[255]), .B(A[255]), .Z(n175) );
  AND U178 ( .A(n176), .B(n177), .Z(n174) );
  NANDN U179 ( .A(B[254]), .B(n178), .Z(n177) );
  NANDN U180 ( .A(A[254]), .B(n179), .Z(n178) );
  NANDN U181 ( .A(n179), .B(A[254]), .Z(n176) );
  XOR U182 ( .A(n179), .B(n180), .Z(DIFF[254]) );
  XOR U183 ( .A(B[254]), .B(A[254]), .Z(n180) );
  AND U184 ( .A(n181), .B(n182), .Z(n179) );
  NANDN U185 ( .A(B[253]), .B(n183), .Z(n182) );
  NANDN U186 ( .A(A[253]), .B(n184), .Z(n183) );
  NANDN U187 ( .A(n184), .B(A[253]), .Z(n181) );
  XOR U188 ( .A(n184), .B(n185), .Z(DIFF[253]) );
  XOR U189 ( .A(B[253]), .B(A[253]), .Z(n185) );
  AND U190 ( .A(n186), .B(n187), .Z(n184) );
  NANDN U191 ( .A(B[252]), .B(n188), .Z(n187) );
  NANDN U192 ( .A(A[252]), .B(n189), .Z(n188) );
  NANDN U193 ( .A(n189), .B(A[252]), .Z(n186) );
  XOR U194 ( .A(n189), .B(n190), .Z(DIFF[252]) );
  XOR U195 ( .A(B[252]), .B(A[252]), .Z(n190) );
  AND U196 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U197 ( .A(B[251]), .B(n193), .Z(n192) );
  NANDN U198 ( .A(A[251]), .B(n194), .Z(n193) );
  NANDN U199 ( .A(n194), .B(A[251]), .Z(n191) );
  XOR U200 ( .A(n194), .B(n195), .Z(DIFF[251]) );
  XOR U201 ( .A(B[251]), .B(A[251]), .Z(n195) );
  AND U202 ( .A(n196), .B(n197), .Z(n194) );
  NANDN U203 ( .A(B[250]), .B(n198), .Z(n197) );
  NANDN U204 ( .A(A[250]), .B(n199), .Z(n198) );
  NANDN U205 ( .A(n199), .B(A[250]), .Z(n196) );
  XOR U206 ( .A(n199), .B(n200), .Z(DIFF[250]) );
  XOR U207 ( .A(B[250]), .B(A[250]), .Z(n200) );
  AND U208 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U209 ( .A(B[249]), .B(n203), .Z(n202) );
  NANDN U210 ( .A(A[249]), .B(n204), .Z(n203) );
  NANDN U211 ( .A(n204), .B(A[249]), .Z(n201) );
  XOR U212 ( .A(n205), .B(n206), .Z(DIFF[24]) );
  XOR U213 ( .A(B[24]), .B(A[24]), .Z(n206) );
  XOR U214 ( .A(n204), .B(n207), .Z(DIFF[249]) );
  XOR U215 ( .A(B[249]), .B(A[249]), .Z(n207) );
  AND U216 ( .A(n208), .B(n209), .Z(n204) );
  NANDN U217 ( .A(B[248]), .B(n210), .Z(n209) );
  NANDN U218 ( .A(A[248]), .B(n211), .Z(n210) );
  NANDN U219 ( .A(n211), .B(A[248]), .Z(n208) );
  XOR U220 ( .A(n211), .B(n212), .Z(DIFF[248]) );
  XOR U221 ( .A(B[248]), .B(A[248]), .Z(n212) );
  AND U222 ( .A(n213), .B(n214), .Z(n211) );
  NANDN U223 ( .A(B[247]), .B(n215), .Z(n214) );
  NANDN U224 ( .A(A[247]), .B(n216), .Z(n215) );
  NANDN U225 ( .A(n216), .B(A[247]), .Z(n213) );
  XOR U226 ( .A(n216), .B(n217), .Z(DIFF[247]) );
  XOR U227 ( .A(B[247]), .B(A[247]), .Z(n217) );
  AND U228 ( .A(n218), .B(n219), .Z(n216) );
  NANDN U229 ( .A(B[246]), .B(n220), .Z(n219) );
  NANDN U230 ( .A(A[246]), .B(n221), .Z(n220) );
  NANDN U231 ( .A(n221), .B(A[246]), .Z(n218) );
  XOR U232 ( .A(n221), .B(n222), .Z(DIFF[246]) );
  XOR U233 ( .A(B[246]), .B(A[246]), .Z(n222) );
  AND U234 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U235 ( .A(B[245]), .B(n225), .Z(n224) );
  NANDN U236 ( .A(A[245]), .B(n226), .Z(n225) );
  NANDN U237 ( .A(n226), .B(A[245]), .Z(n223) );
  XOR U238 ( .A(n226), .B(n227), .Z(DIFF[245]) );
  XOR U239 ( .A(B[245]), .B(A[245]), .Z(n227) );
  AND U240 ( .A(n228), .B(n229), .Z(n226) );
  NANDN U241 ( .A(B[244]), .B(n230), .Z(n229) );
  NANDN U242 ( .A(A[244]), .B(n231), .Z(n230) );
  NANDN U243 ( .A(n231), .B(A[244]), .Z(n228) );
  XOR U244 ( .A(n231), .B(n232), .Z(DIFF[244]) );
  XOR U245 ( .A(B[244]), .B(A[244]), .Z(n232) );
  AND U246 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U247 ( .A(B[243]), .B(n235), .Z(n234) );
  NANDN U248 ( .A(A[243]), .B(n236), .Z(n235) );
  NANDN U249 ( .A(n236), .B(A[243]), .Z(n233) );
  XOR U250 ( .A(n236), .B(n237), .Z(DIFF[243]) );
  XOR U251 ( .A(B[243]), .B(A[243]), .Z(n237) );
  AND U252 ( .A(n238), .B(n239), .Z(n236) );
  NANDN U253 ( .A(B[242]), .B(n240), .Z(n239) );
  NANDN U254 ( .A(A[242]), .B(n241), .Z(n240) );
  NANDN U255 ( .A(n241), .B(A[242]), .Z(n238) );
  XOR U256 ( .A(n241), .B(n242), .Z(DIFF[242]) );
  XOR U257 ( .A(B[242]), .B(A[242]), .Z(n242) );
  AND U258 ( .A(n243), .B(n244), .Z(n241) );
  NANDN U259 ( .A(B[241]), .B(n245), .Z(n244) );
  NANDN U260 ( .A(A[241]), .B(n246), .Z(n245) );
  NANDN U261 ( .A(n246), .B(A[241]), .Z(n243) );
  XOR U262 ( .A(n246), .B(n247), .Z(DIFF[241]) );
  XOR U263 ( .A(B[241]), .B(A[241]), .Z(n247) );
  AND U264 ( .A(n248), .B(n249), .Z(n246) );
  NANDN U265 ( .A(B[240]), .B(n250), .Z(n249) );
  NANDN U266 ( .A(A[240]), .B(n251), .Z(n250) );
  NANDN U267 ( .A(n251), .B(A[240]), .Z(n248) );
  XOR U268 ( .A(n251), .B(n252), .Z(DIFF[240]) );
  XOR U269 ( .A(B[240]), .B(A[240]), .Z(n252) );
  AND U270 ( .A(n253), .B(n254), .Z(n251) );
  NANDN U271 ( .A(B[239]), .B(n255), .Z(n254) );
  NANDN U272 ( .A(A[239]), .B(n256), .Z(n255) );
  NANDN U273 ( .A(n256), .B(A[239]), .Z(n253) );
  XOR U274 ( .A(n257), .B(n258), .Z(DIFF[23]) );
  XOR U275 ( .A(B[23]), .B(A[23]), .Z(n258) );
  XOR U276 ( .A(n256), .B(n259), .Z(DIFF[239]) );
  XOR U277 ( .A(B[239]), .B(A[239]), .Z(n259) );
  AND U278 ( .A(n260), .B(n261), .Z(n256) );
  NANDN U279 ( .A(B[238]), .B(n262), .Z(n261) );
  NANDN U280 ( .A(A[238]), .B(n263), .Z(n262) );
  NANDN U281 ( .A(n263), .B(A[238]), .Z(n260) );
  XOR U282 ( .A(n263), .B(n264), .Z(DIFF[238]) );
  XOR U283 ( .A(B[238]), .B(A[238]), .Z(n264) );
  AND U284 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U285 ( .A(B[237]), .B(n267), .Z(n266) );
  NANDN U286 ( .A(A[237]), .B(n268), .Z(n267) );
  NANDN U287 ( .A(n268), .B(A[237]), .Z(n265) );
  XOR U288 ( .A(n268), .B(n269), .Z(DIFF[237]) );
  XOR U289 ( .A(B[237]), .B(A[237]), .Z(n269) );
  AND U290 ( .A(n270), .B(n271), .Z(n268) );
  NANDN U291 ( .A(B[236]), .B(n272), .Z(n271) );
  NANDN U292 ( .A(A[236]), .B(n273), .Z(n272) );
  NANDN U293 ( .A(n273), .B(A[236]), .Z(n270) );
  XOR U294 ( .A(n273), .B(n274), .Z(DIFF[236]) );
  XOR U295 ( .A(B[236]), .B(A[236]), .Z(n274) );
  AND U296 ( .A(n275), .B(n276), .Z(n273) );
  NANDN U297 ( .A(B[235]), .B(n277), .Z(n276) );
  NANDN U298 ( .A(A[235]), .B(n278), .Z(n277) );
  NANDN U299 ( .A(n278), .B(A[235]), .Z(n275) );
  XOR U300 ( .A(n278), .B(n279), .Z(DIFF[235]) );
  XOR U301 ( .A(B[235]), .B(A[235]), .Z(n279) );
  AND U302 ( .A(n280), .B(n281), .Z(n278) );
  NANDN U303 ( .A(B[234]), .B(n282), .Z(n281) );
  NANDN U304 ( .A(A[234]), .B(n283), .Z(n282) );
  NANDN U305 ( .A(n283), .B(A[234]), .Z(n280) );
  XOR U306 ( .A(n283), .B(n284), .Z(DIFF[234]) );
  XOR U307 ( .A(B[234]), .B(A[234]), .Z(n284) );
  AND U308 ( .A(n285), .B(n286), .Z(n283) );
  NANDN U309 ( .A(B[233]), .B(n287), .Z(n286) );
  NANDN U310 ( .A(A[233]), .B(n288), .Z(n287) );
  NANDN U311 ( .A(n288), .B(A[233]), .Z(n285) );
  XOR U312 ( .A(n288), .B(n289), .Z(DIFF[233]) );
  XOR U313 ( .A(B[233]), .B(A[233]), .Z(n289) );
  AND U314 ( .A(n290), .B(n291), .Z(n288) );
  NANDN U315 ( .A(B[232]), .B(n292), .Z(n291) );
  NANDN U316 ( .A(A[232]), .B(n293), .Z(n292) );
  NANDN U317 ( .A(n293), .B(A[232]), .Z(n290) );
  XOR U318 ( .A(n293), .B(n294), .Z(DIFF[232]) );
  XOR U319 ( .A(B[232]), .B(A[232]), .Z(n294) );
  AND U320 ( .A(n295), .B(n296), .Z(n293) );
  NANDN U321 ( .A(B[231]), .B(n297), .Z(n296) );
  NANDN U322 ( .A(A[231]), .B(n298), .Z(n297) );
  NANDN U323 ( .A(n298), .B(A[231]), .Z(n295) );
  XOR U324 ( .A(n298), .B(n299), .Z(DIFF[231]) );
  XOR U325 ( .A(B[231]), .B(A[231]), .Z(n299) );
  AND U326 ( .A(n300), .B(n301), .Z(n298) );
  NANDN U327 ( .A(B[230]), .B(n302), .Z(n301) );
  NANDN U328 ( .A(A[230]), .B(n303), .Z(n302) );
  NANDN U329 ( .A(n303), .B(A[230]), .Z(n300) );
  XOR U330 ( .A(n303), .B(n304), .Z(DIFF[230]) );
  XOR U331 ( .A(B[230]), .B(A[230]), .Z(n304) );
  AND U332 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U333 ( .A(B[229]), .B(n307), .Z(n306) );
  NANDN U334 ( .A(A[229]), .B(n308), .Z(n307) );
  NANDN U335 ( .A(n308), .B(A[229]), .Z(n305) );
  XOR U336 ( .A(n309), .B(n310), .Z(DIFF[22]) );
  XOR U337 ( .A(B[22]), .B(A[22]), .Z(n310) );
  XOR U338 ( .A(n308), .B(n311), .Z(DIFF[229]) );
  XOR U339 ( .A(B[229]), .B(A[229]), .Z(n311) );
  AND U340 ( .A(n312), .B(n313), .Z(n308) );
  NANDN U341 ( .A(B[228]), .B(n314), .Z(n313) );
  NANDN U342 ( .A(A[228]), .B(n315), .Z(n314) );
  NANDN U343 ( .A(n315), .B(A[228]), .Z(n312) );
  XOR U344 ( .A(n315), .B(n316), .Z(DIFF[228]) );
  XOR U345 ( .A(B[228]), .B(A[228]), .Z(n316) );
  AND U346 ( .A(n317), .B(n318), .Z(n315) );
  NANDN U347 ( .A(B[227]), .B(n319), .Z(n318) );
  NANDN U348 ( .A(A[227]), .B(n320), .Z(n319) );
  NANDN U349 ( .A(n320), .B(A[227]), .Z(n317) );
  XOR U350 ( .A(n320), .B(n321), .Z(DIFF[227]) );
  XOR U351 ( .A(B[227]), .B(A[227]), .Z(n321) );
  AND U352 ( .A(n322), .B(n323), .Z(n320) );
  NANDN U353 ( .A(B[226]), .B(n324), .Z(n323) );
  NANDN U354 ( .A(A[226]), .B(n325), .Z(n324) );
  NANDN U355 ( .A(n325), .B(A[226]), .Z(n322) );
  XOR U356 ( .A(n325), .B(n326), .Z(DIFF[226]) );
  XOR U357 ( .A(B[226]), .B(A[226]), .Z(n326) );
  AND U358 ( .A(n327), .B(n328), .Z(n325) );
  NANDN U359 ( .A(B[225]), .B(n329), .Z(n328) );
  NANDN U360 ( .A(A[225]), .B(n330), .Z(n329) );
  NANDN U361 ( .A(n330), .B(A[225]), .Z(n327) );
  XOR U362 ( .A(n330), .B(n331), .Z(DIFF[225]) );
  XOR U363 ( .A(B[225]), .B(A[225]), .Z(n331) );
  AND U364 ( .A(n332), .B(n333), .Z(n330) );
  NANDN U365 ( .A(B[224]), .B(n334), .Z(n333) );
  NANDN U366 ( .A(A[224]), .B(n335), .Z(n334) );
  NANDN U367 ( .A(n335), .B(A[224]), .Z(n332) );
  XOR U368 ( .A(n335), .B(n336), .Z(DIFF[224]) );
  XOR U369 ( .A(B[224]), .B(A[224]), .Z(n336) );
  AND U370 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U371 ( .A(B[223]), .B(n339), .Z(n338) );
  NANDN U372 ( .A(A[223]), .B(n340), .Z(n339) );
  NANDN U373 ( .A(n340), .B(A[223]), .Z(n337) );
  XOR U374 ( .A(n340), .B(n341), .Z(DIFF[223]) );
  XOR U375 ( .A(B[223]), .B(A[223]), .Z(n341) );
  AND U376 ( .A(n342), .B(n343), .Z(n340) );
  NANDN U377 ( .A(B[222]), .B(n344), .Z(n343) );
  NANDN U378 ( .A(A[222]), .B(n345), .Z(n344) );
  NANDN U379 ( .A(n345), .B(A[222]), .Z(n342) );
  XOR U380 ( .A(n345), .B(n346), .Z(DIFF[222]) );
  XOR U381 ( .A(B[222]), .B(A[222]), .Z(n346) );
  AND U382 ( .A(n347), .B(n348), .Z(n345) );
  NANDN U383 ( .A(B[221]), .B(n349), .Z(n348) );
  NANDN U384 ( .A(A[221]), .B(n350), .Z(n349) );
  NANDN U385 ( .A(n350), .B(A[221]), .Z(n347) );
  XOR U386 ( .A(n350), .B(n351), .Z(DIFF[221]) );
  XOR U387 ( .A(B[221]), .B(A[221]), .Z(n351) );
  AND U388 ( .A(n352), .B(n353), .Z(n350) );
  NANDN U389 ( .A(B[220]), .B(n354), .Z(n353) );
  NANDN U390 ( .A(A[220]), .B(n355), .Z(n354) );
  NANDN U391 ( .A(n355), .B(A[220]), .Z(n352) );
  XOR U392 ( .A(n355), .B(n356), .Z(DIFF[220]) );
  XOR U393 ( .A(B[220]), .B(A[220]), .Z(n356) );
  AND U394 ( .A(n357), .B(n358), .Z(n355) );
  NANDN U395 ( .A(B[219]), .B(n359), .Z(n358) );
  NANDN U396 ( .A(A[219]), .B(n360), .Z(n359) );
  NANDN U397 ( .A(n360), .B(A[219]), .Z(n357) );
  XOR U398 ( .A(n361), .B(n362), .Z(DIFF[21]) );
  XOR U399 ( .A(B[21]), .B(A[21]), .Z(n362) );
  XOR U400 ( .A(n360), .B(n363), .Z(DIFF[219]) );
  XOR U401 ( .A(B[219]), .B(A[219]), .Z(n363) );
  AND U402 ( .A(n364), .B(n365), .Z(n360) );
  NANDN U403 ( .A(B[218]), .B(n366), .Z(n365) );
  NANDN U404 ( .A(A[218]), .B(n367), .Z(n366) );
  NANDN U405 ( .A(n367), .B(A[218]), .Z(n364) );
  XOR U406 ( .A(n367), .B(n368), .Z(DIFF[218]) );
  XOR U407 ( .A(B[218]), .B(A[218]), .Z(n368) );
  AND U408 ( .A(n369), .B(n370), .Z(n367) );
  NANDN U409 ( .A(B[217]), .B(n371), .Z(n370) );
  NANDN U410 ( .A(A[217]), .B(n372), .Z(n371) );
  NANDN U411 ( .A(n372), .B(A[217]), .Z(n369) );
  XOR U412 ( .A(n372), .B(n373), .Z(DIFF[217]) );
  XOR U413 ( .A(B[217]), .B(A[217]), .Z(n373) );
  AND U414 ( .A(n374), .B(n375), .Z(n372) );
  NANDN U415 ( .A(B[216]), .B(n376), .Z(n375) );
  NANDN U416 ( .A(A[216]), .B(n377), .Z(n376) );
  NANDN U417 ( .A(n377), .B(A[216]), .Z(n374) );
  XOR U418 ( .A(n377), .B(n378), .Z(DIFF[216]) );
  XOR U419 ( .A(B[216]), .B(A[216]), .Z(n378) );
  AND U420 ( .A(n379), .B(n380), .Z(n377) );
  NANDN U421 ( .A(B[215]), .B(n381), .Z(n380) );
  NANDN U422 ( .A(A[215]), .B(n382), .Z(n381) );
  NANDN U423 ( .A(n382), .B(A[215]), .Z(n379) );
  XOR U424 ( .A(n382), .B(n383), .Z(DIFF[215]) );
  XOR U425 ( .A(B[215]), .B(A[215]), .Z(n383) );
  AND U426 ( .A(n384), .B(n385), .Z(n382) );
  NANDN U427 ( .A(B[214]), .B(n386), .Z(n385) );
  NANDN U428 ( .A(A[214]), .B(n387), .Z(n386) );
  NANDN U429 ( .A(n387), .B(A[214]), .Z(n384) );
  XOR U430 ( .A(n387), .B(n388), .Z(DIFF[214]) );
  XOR U431 ( .A(B[214]), .B(A[214]), .Z(n388) );
  AND U432 ( .A(n389), .B(n390), .Z(n387) );
  NANDN U433 ( .A(B[213]), .B(n391), .Z(n390) );
  NANDN U434 ( .A(A[213]), .B(n392), .Z(n391) );
  NANDN U435 ( .A(n392), .B(A[213]), .Z(n389) );
  XOR U436 ( .A(n392), .B(n393), .Z(DIFF[213]) );
  XOR U437 ( .A(B[213]), .B(A[213]), .Z(n393) );
  AND U438 ( .A(n394), .B(n395), .Z(n392) );
  NANDN U439 ( .A(B[212]), .B(n396), .Z(n395) );
  NANDN U440 ( .A(A[212]), .B(n397), .Z(n396) );
  NANDN U441 ( .A(n397), .B(A[212]), .Z(n394) );
  XOR U442 ( .A(n397), .B(n398), .Z(DIFF[212]) );
  XOR U443 ( .A(B[212]), .B(A[212]), .Z(n398) );
  AND U444 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U445 ( .A(B[211]), .B(n401), .Z(n400) );
  NANDN U446 ( .A(A[211]), .B(n402), .Z(n401) );
  NANDN U447 ( .A(n402), .B(A[211]), .Z(n399) );
  XOR U448 ( .A(n402), .B(n403), .Z(DIFF[211]) );
  XOR U449 ( .A(B[211]), .B(A[211]), .Z(n403) );
  AND U450 ( .A(n404), .B(n405), .Z(n402) );
  NANDN U451 ( .A(B[210]), .B(n406), .Z(n405) );
  NANDN U452 ( .A(A[210]), .B(n407), .Z(n406) );
  NANDN U453 ( .A(n407), .B(A[210]), .Z(n404) );
  XOR U454 ( .A(n407), .B(n408), .Z(DIFF[210]) );
  XOR U455 ( .A(B[210]), .B(A[210]), .Z(n408) );
  AND U456 ( .A(n409), .B(n410), .Z(n407) );
  NANDN U457 ( .A(B[209]), .B(n411), .Z(n410) );
  NANDN U458 ( .A(A[209]), .B(n412), .Z(n411) );
  NANDN U459 ( .A(n412), .B(A[209]), .Z(n409) );
  XOR U460 ( .A(n413), .B(n414), .Z(DIFF[20]) );
  XOR U461 ( .A(B[20]), .B(A[20]), .Z(n414) );
  XOR U462 ( .A(n412), .B(n415), .Z(DIFF[209]) );
  XOR U463 ( .A(B[209]), .B(A[209]), .Z(n415) );
  AND U464 ( .A(n416), .B(n417), .Z(n412) );
  NANDN U465 ( .A(B[208]), .B(n418), .Z(n417) );
  NANDN U466 ( .A(A[208]), .B(n419), .Z(n418) );
  NANDN U467 ( .A(n419), .B(A[208]), .Z(n416) );
  XOR U468 ( .A(n419), .B(n420), .Z(DIFF[208]) );
  XOR U469 ( .A(B[208]), .B(A[208]), .Z(n420) );
  AND U470 ( .A(n421), .B(n422), .Z(n419) );
  NANDN U471 ( .A(B[207]), .B(n423), .Z(n422) );
  NANDN U472 ( .A(A[207]), .B(n424), .Z(n423) );
  NANDN U473 ( .A(n424), .B(A[207]), .Z(n421) );
  XOR U474 ( .A(n424), .B(n425), .Z(DIFF[207]) );
  XOR U475 ( .A(B[207]), .B(A[207]), .Z(n425) );
  AND U476 ( .A(n426), .B(n427), .Z(n424) );
  NANDN U477 ( .A(B[206]), .B(n428), .Z(n427) );
  NANDN U478 ( .A(A[206]), .B(n429), .Z(n428) );
  NANDN U479 ( .A(n429), .B(A[206]), .Z(n426) );
  XOR U480 ( .A(n429), .B(n430), .Z(DIFF[206]) );
  XOR U481 ( .A(B[206]), .B(A[206]), .Z(n430) );
  AND U482 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U483 ( .A(B[205]), .B(n433), .Z(n432) );
  NANDN U484 ( .A(A[205]), .B(n434), .Z(n433) );
  NANDN U485 ( .A(n434), .B(A[205]), .Z(n431) );
  XOR U486 ( .A(n434), .B(n435), .Z(DIFF[205]) );
  XOR U487 ( .A(B[205]), .B(A[205]), .Z(n435) );
  AND U488 ( .A(n436), .B(n437), .Z(n434) );
  NANDN U489 ( .A(B[204]), .B(n438), .Z(n437) );
  NANDN U490 ( .A(A[204]), .B(n439), .Z(n438) );
  NANDN U491 ( .A(n439), .B(A[204]), .Z(n436) );
  XOR U492 ( .A(n439), .B(n440), .Z(DIFF[204]) );
  XOR U493 ( .A(B[204]), .B(A[204]), .Z(n440) );
  AND U494 ( .A(n441), .B(n442), .Z(n439) );
  NANDN U495 ( .A(B[203]), .B(n443), .Z(n442) );
  NANDN U496 ( .A(A[203]), .B(n444), .Z(n443) );
  NANDN U497 ( .A(n444), .B(A[203]), .Z(n441) );
  XOR U498 ( .A(n444), .B(n445), .Z(DIFF[203]) );
  XOR U499 ( .A(B[203]), .B(A[203]), .Z(n445) );
  AND U500 ( .A(n446), .B(n447), .Z(n444) );
  NANDN U501 ( .A(B[202]), .B(n448), .Z(n447) );
  NANDN U502 ( .A(A[202]), .B(n449), .Z(n448) );
  NANDN U503 ( .A(n449), .B(A[202]), .Z(n446) );
  XOR U504 ( .A(n449), .B(n450), .Z(DIFF[202]) );
  XOR U505 ( .A(B[202]), .B(A[202]), .Z(n450) );
  AND U506 ( .A(n451), .B(n452), .Z(n449) );
  NANDN U507 ( .A(B[201]), .B(n453), .Z(n452) );
  NANDN U508 ( .A(A[201]), .B(n454), .Z(n453) );
  NANDN U509 ( .A(n454), .B(A[201]), .Z(n451) );
  XOR U510 ( .A(n454), .B(n455), .Z(DIFF[201]) );
  XOR U511 ( .A(B[201]), .B(A[201]), .Z(n455) );
  AND U512 ( .A(n456), .B(n457), .Z(n454) );
  NANDN U513 ( .A(B[200]), .B(n458), .Z(n457) );
  NANDN U514 ( .A(A[200]), .B(n459), .Z(n458) );
  NANDN U515 ( .A(n459), .B(A[200]), .Z(n456) );
  XOR U516 ( .A(n459), .B(n460), .Z(DIFF[200]) );
  XOR U517 ( .A(B[200]), .B(A[200]), .Z(n460) );
  AND U518 ( .A(n461), .B(n462), .Z(n459) );
  NANDN U519 ( .A(B[199]), .B(n463), .Z(n462) );
  NANDN U520 ( .A(A[199]), .B(n464), .Z(n463) );
  NANDN U521 ( .A(n464), .B(A[199]), .Z(n461) );
  XOR U522 ( .A(n2), .B(n465), .Z(DIFF[1]) );
  XOR U523 ( .A(B[1]), .B(A[1]), .Z(n465) );
  XOR U524 ( .A(n466), .B(n467), .Z(DIFF[19]) );
  XOR U525 ( .A(B[19]), .B(A[19]), .Z(n467) );
  XOR U526 ( .A(n464), .B(n468), .Z(DIFF[199]) );
  XOR U527 ( .A(B[199]), .B(A[199]), .Z(n468) );
  AND U528 ( .A(n469), .B(n470), .Z(n464) );
  NANDN U529 ( .A(B[198]), .B(n471), .Z(n470) );
  NANDN U530 ( .A(A[198]), .B(n472), .Z(n471) );
  NANDN U531 ( .A(n472), .B(A[198]), .Z(n469) );
  XOR U532 ( .A(n472), .B(n473), .Z(DIFF[198]) );
  XOR U533 ( .A(B[198]), .B(A[198]), .Z(n473) );
  AND U534 ( .A(n474), .B(n475), .Z(n472) );
  NANDN U535 ( .A(B[197]), .B(n476), .Z(n475) );
  NANDN U536 ( .A(A[197]), .B(n477), .Z(n476) );
  NANDN U537 ( .A(n477), .B(A[197]), .Z(n474) );
  XOR U538 ( .A(n477), .B(n478), .Z(DIFF[197]) );
  XOR U539 ( .A(B[197]), .B(A[197]), .Z(n478) );
  AND U540 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U541 ( .A(B[196]), .B(n481), .Z(n480) );
  NANDN U542 ( .A(A[196]), .B(n482), .Z(n481) );
  NANDN U543 ( .A(n482), .B(A[196]), .Z(n479) );
  XOR U544 ( .A(n482), .B(n483), .Z(DIFF[196]) );
  XOR U545 ( .A(B[196]), .B(A[196]), .Z(n483) );
  AND U546 ( .A(n484), .B(n485), .Z(n482) );
  NANDN U547 ( .A(B[195]), .B(n486), .Z(n485) );
  NANDN U548 ( .A(A[195]), .B(n487), .Z(n486) );
  NANDN U549 ( .A(n487), .B(A[195]), .Z(n484) );
  XOR U550 ( .A(n487), .B(n488), .Z(DIFF[195]) );
  XOR U551 ( .A(B[195]), .B(A[195]), .Z(n488) );
  AND U552 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U553 ( .A(B[194]), .B(n491), .Z(n490) );
  NANDN U554 ( .A(A[194]), .B(n492), .Z(n491) );
  NANDN U555 ( .A(n492), .B(A[194]), .Z(n489) );
  XOR U556 ( .A(n492), .B(n493), .Z(DIFF[194]) );
  XOR U557 ( .A(B[194]), .B(A[194]), .Z(n493) );
  AND U558 ( .A(n494), .B(n495), .Z(n492) );
  NANDN U559 ( .A(B[193]), .B(n496), .Z(n495) );
  NANDN U560 ( .A(A[193]), .B(n497), .Z(n496) );
  NANDN U561 ( .A(n497), .B(A[193]), .Z(n494) );
  XOR U562 ( .A(n497), .B(n498), .Z(DIFF[193]) );
  XOR U563 ( .A(B[193]), .B(A[193]), .Z(n498) );
  AND U564 ( .A(n499), .B(n500), .Z(n497) );
  NANDN U565 ( .A(B[192]), .B(n501), .Z(n500) );
  NANDN U566 ( .A(A[192]), .B(n502), .Z(n501) );
  NANDN U567 ( .A(n502), .B(A[192]), .Z(n499) );
  XOR U568 ( .A(n502), .B(n503), .Z(DIFF[192]) );
  XOR U569 ( .A(B[192]), .B(A[192]), .Z(n503) );
  AND U570 ( .A(n504), .B(n505), .Z(n502) );
  NANDN U571 ( .A(B[191]), .B(n506), .Z(n505) );
  NANDN U572 ( .A(A[191]), .B(n507), .Z(n506) );
  NANDN U573 ( .A(n507), .B(A[191]), .Z(n504) );
  XOR U574 ( .A(n507), .B(n508), .Z(DIFF[191]) );
  XOR U575 ( .A(B[191]), .B(A[191]), .Z(n508) );
  AND U576 ( .A(n509), .B(n510), .Z(n507) );
  NANDN U577 ( .A(B[190]), .B(n511), .Z(n510) );
  NANDN U578 ( .A(A[190]), .B(n512), .Z(n511) );
  NANDN U579 ( .A(n512), .B(A[190]), .Z(n509) );
  XOR U580 ( .A(n512), .B(n513), .Z(DIFF[190]) );
  XOR U581 ( .A(B[190]), .B(A[190]), .Z(n513) );
  AND U582 ( .A(n514), .B(n515), .Z(n512) );
  NANDN U583 ( .A(B[189]), .B(n516), .Z(n515) );
  NANDN U584 ( .A(A[189]), .B(n517), .Z(n516) );
  NANDN U585 ( .A(n517), .B(A[189]), .Z(n514) );
  XOR U586 ( .A(n518), .B(n519), .Z(DIFF[18]) );
  XOR U587 ( .A(B[18]), .B(A[18]), .Z(n519) );
  XOR U588 ( .A(n517), .B(n520), .Z(DIFF[189]) );
  XOR U589 ( .A(B[189]), .B(A[189]), .Z(n520) );
  AND U590 ( .A(n521), .B(n522), .Z(n517) );
  NANDN U591 ( .A(B[188]), .B(n523), .Z(n522) );
  NANDN U592 ( .A(A[188]), .B(n524), .Z(n523) );
  NANDN U593 ( .A(n524), .B(A[188]), .Z(n521) );
  XOR U594 ( .A(n524), .B(n525), .Z(DIFF[188]) );
  XOR U595 ( .A(B[188]), .B(A[188]), .Z(n525) );
  AND U596 ( .A(n526), .B(n527), .Z(n524) );
  NANDN U597 ( .A(B[187]), .B(n528), .Z(n527) );
  NANDN U598 ( .A(A[187]), .B(n529), .Z(n528) );
  NANDN U599 ( .A(n529), .B(A[187]), .Z(n526) );
  XOR U600 ( .A(n529), .B(n530), .Z(DIFF[187]) );
  XOR U601 ( .A(B[187]), .B(A[187]), .Z(n530) );
  AND U602 ( .A(n531), .B(n532), .Z(n529) );
  NANDN U603 ( .A(B[186]), .B(n533), .Z(n532) );
  NANDN U604 ( .A(A[186]), .B(n534), .Z(n533) );
  NANDN U605 ( .A(n534), .B(A[186]), .Z(n531) );
  XOR U606 ( .A(n534), .B(n535), .Z(DIFF[186]) );
  XOR U607 ( .A(B[186]), .B(A[186]), .Z(n535) );
  AND U608 ( .A(n536), .B(n537), .Z(n534) );
  NANDN U609 ( .A(B[185]), .B(n538), .Z(n537) );
  NANDN U610 ( .A(A[185]), .B(n539), .Z(n538) );
  NANDN U611 ( .A(n539), .B(A[185]), .Z(n536) );
  XOR U612 ( .A(n539), .B(n540), .Z(DIFF[185]) );
  XOR U613 ( .A(B[185]), .B(A[185]), .Z(n540) );
  AND U614 ( .A(n541), .B(n542), .Z(n539) );
  NANDN U615 ( .A(B[184]), .B(n543), .Z(n542) );
  NANDN U616 ( .A(A[184]), .B(n544), .Z(n543) );
  NANDN U617 ( .A(n544), .B(A[184]), .Z(n541) );
  XOR U618 ( .A(n544), .B(n545), .Z(DIFF[184]) );
  XOR U619 ( .A(B[184]), .B(A[184]), .Z(n545) );
  AND U620 ( .A(n546), .B(n547), .Z(n544) );
  NANDN U621 ( .A(B[183]), .B(n548), .Z(n547) );
  NANDN U622 ( .A(A[183]), .B(n549), .Z(n548) );
  NANDN U623 ( .A(n549), .B(A[183]), .Z(n546) );
  XOR U624 ( .A(n549), .B(n550), .Z(DIFF[183]) );
  XOR U625 ( .A(B[183]), .B(A[183]), .Z(n550) );
  AND U626 ( .A(n551), .B(n552), .Z(n549) );
  NANDN U627 ( .A(B[182]), .B(n553), .Z(n552) );
  NANDN U628 ( .A(A[182]), .B(n554), .Z(n553) );
  NANDN U629 ( .A(n554), .B(A[182]), .Z(n551) );
  XOR U630 ( .A(n554), .B(n555), .Z(DIFF[182]) );
  XOR U631 ( .A(B[182]), .B(A[182]), .Z(n555) );
  AND U632 ( .A(n556), .B(n557), .Z(n554) );
  NANDN U633 ( .A(B[181]), .B(n558), .Z(n557) );
  NANDN U634 ( .A(A[181]), .B(n559), .Z(n558) );
  NANDN U635 ( .A(n559), .B(A[181]), .Z(n556) );
  XOR U636 ( .A(n559), .B(n560), .Z(DIFF[181]) );
  XOR U637 ( .A(B[181]), .B(A[181]), .Z(n560) );
  AND U638 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U639 ( .A(B[180]), .B(n563), .Z(n562) );
  NANDN U640 ( .A(A[180]), .B(n564), .Z(n563) );
  NANDN U641 ( .A(n564), .B(A[180]), .Z(n561) );
  XOR U642 ( .A(n564), .B(n565), .Z(DIFF[180]) );
  XOR U643 ( .A(B[180]), .B(A[180]), .Z(n565) );
  AND U644 ( .A(n566), .B(n567), .Z(n564) );
  NANDN U645 ( .A(B[179]), .B(n568), .Z(n567) );
  NANDN U646 ( .A(A[179]), .B(n569), .Z(n568) );
  NANDN U647 ( .A(n569), .B(A[179]), .Z(n566) );
  XOR U648 ( .A(n570), .B(n571), .Z(DIFF[17]) );
  XOR U649 ( .A(B[17]), .B(A[17]), .Z(n571) );
  XOR U650 ( .A(n569), .B(n572), .Z(DIFF[179]) );
  XOR U651 ( .A(B[179]), .B(A[179]), .Z(n572) );
  AND U652 ( .A(n573), .B(n574), .Z(n569) );
  NANDN U653 ( .A(B[178]), .B(n575), .Z(n574) );
  NANDN U654 ( .A(A[178]), .B(n576), .Z(n575) );
  NANDN U655 ( .A(n576), .B(A[178]), .Z(n573) );
  XOR U656 ( .A(n576), .B(n577), .Z(DIFF[178]) );
  XOR U657 ( .A(B[178]), .B(A[178]), .Z(n577) );
  AND U658 ( .A(n578), .B(n579), .Z(n576) );
  NANDN U659 ( .A(B[177]), .B(n580), .Z(n579) );
  NANDN U660 ( .A(A[177]), .B(n581), .Z(n580) );
  NANDN U661 ( .A(n581), .B(A[177]), .Z(n578) );
  XOR U662 ( .A(n581), .B(n582), .Z(DIFF[177]) );
  XOR U663 ( .A(B[177]), .B(A[177]), .Z(n582) );
  AND U664 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U665 ( .A(B[176]), .B(n585), .Z(n584) );
  NANDN U666 ( .A(A[176]), .B(n586), .Z(n585) );
  NANDN U667 ( .A(n586), .B(A[176]), .Z(n583) );
  XOR U668 ( .A(n586), .B(n587), .Z(DIFF[176]) );
  XOR U669 ( .A(B[176]), .B(A[176]), .Z(n587) );
  AND U670 ( .A(n588), .B(n589), .Z(n586) );
  NANDN U671 ( .A(B[175]), .B(n590), .Z(n589) );
  NANDN U672 ( .A(A[175]), .B(n591), .Z(n590) );
  NANDN U673 ( .A(n591), .B(A[175]), .Z(n588) );
  XOR U674 ( .A(n591), .B(n592), .Z(DIFF[175]) );
  XOR U675 ( .A(B[175]), .B(A[175]), .Z(n592) );
  AND U676 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U677 ( .A(B[174]), .B(n595), .Z(n594) );
  NANDN U678 ( .A(A[174]), .B(n596), .Z(n595) );
  NANDN U679 ( .A(n596), .B(A[174]), .Z(n593) );
  XOR U680 ( .A(n596), .B(n597), .Z(DIFF[174]) );
  XOR U681 ( .A(B[174]), .B(A[174]), .Z(n597) );
  AND U682 ( .A(n598), .B(n599), .Z(n596) );
  NANDN U683 ( .A(B[173]), .B(n600), .Z(n599) );
  NANDN U684 ( .A(A[173]), .B(n601), .Z(n600) );
  NANDN U685 ( .A(n601), .B(A[173]), .Z(n598) );
  XOR U686 ( .A(n601), .B(n602), .Z(DIFF[173]) );
  XOR U687 ( .A(B[173]), .B(A[173]), .Z(n602) );
  AND U688 ( .A(n603), .B(n604), .Z(n601) );
  NANDN U689 ( .A(B[172]), .B(n605), .Z(n604) );
  NANDN U690 ( .A(A[172]), .B(n606), .Z(n605) );
  NANDN U691 ( .A(n606), .B(A[172]), .Z(n603) );
  XOR U692 ( .A(n606), .B(n607), .Z(DIFF[172]) );
  XOR U693 ( .A(B[172]), .B(A[172]), .Z(n607) );
  AND U694 ( .A(n608), .B(n609), .Z(n606) );
  NANDN U695 ( .A(B[171]), .B(n610), .Z(n609) );
  NANDN U696 ( .A(A[171]), .B(n611), .Z(n610) );
  NANDN U697 ( .A(n611), .B(A[171]), .Z(n608) );
  XOR U698 ( .A(n611), .B(n612), .Z(DIFF[171]) );
  XOR U699 ( .A(B[171]), .B(A[171]), .Z(n612) );
  AND U700 ( .A(n613), .B(n614), .Z(n611) );
  NANDN U701 ( .A(B[170]), .B(n615), .Z(n614) );
  NANDN U702 ( .A(A[170]), .B(n616), .Z(n615) );
  NANDN U703 ( .A(n616), .B(A[170]), .Z(n613) );
  XOR U704 ( .A(n616), .B(n617), .Z(DIFF[170]) );
  XOR U705 ( .A(B[170]), .B(A[170]), .Z(n617) );
  AND U706 ( .A(n618), .B(n619), .Z(n616) );
  NANDN U707 ( .A(B[169]), .B(n620), .Z(n619) );
  NANDN U708 ( .A(A[169]), .B(n621), .Z(n620) );
  NANDN U709 ( .A(n621), .B(A[169]), .Z(n618) );
  XOR U710 ( .A(n622), .B(n623), .Z(DIFF[16]) );
  XOR U711 ( .A(B[16]), .B(A[16]), .Z(n623) );
  XOR U712 ( .A(n621), .B(n624), .Z(DIFF[169]) );
  XOR U713 ( .A(B[169]), .B(A[169]), .Z(n624) );
  AND U714 ( .A(n625), .B(n626), .Z(n621) );
  NANDN U715 ( .A(B[168]), .B(n627), .Z(n626) );
  NANDN U716 ( .A(A[168]), .B(n628), .Z(n627) );
  NANDN U717 ( .A(n628), .B(A[168]), .Z(n625) );
  XOR U718 ( .A(n628), .B(n629), .Z(DIFF[168]) );
  XOR U719 ( .A(B[168]), .B(A[168]), .Z(n629) );
  AND U720 ( .A(n630), .B(n631), .Z(n628) );
  NANDN U721 ( .A(B[167]), .B(n632), .Z(n631) );
  NANDN U722 ( .A(A[167]), .B(n633), .Z(n632) );
  NANDN U723 ( .A(n633), .B(A[167]), .Z(n630) );
  XOR U724 ( .A(n633), .B(n634), .Z(DIFF[167]) );
  XOR U725 ( .A(B[167]), .B(A[167]), .Z(n634) );
  AND U726 ( .A(n635), .B(n636), .Z(n633) );
  NANDN U727 ( .A(B[166]), .B(n637), .Z(n636) );
  NANDN U728 ( .A(A[166]), .B(n638), .Z(n637) );
  NANDN U729 ( .A(n638), .B(A[166]), .Z(n635) );
  XOR U730 ( .A(n638), .B(n639), .Z(DIFF[166]) );
  XOR U731 ( .A(B[166]), .B(A[166]), .Z(n639) );
  AND U732 ( .A(n640), .B(n641), .Z(n638) );
  NANDN U733 ( .A(B[165]), .B(n642), .Z(n641) );
  NANDN U734 ( .A(A[165]), .B(n643), .Z(n642) );
  NANDN U735 ( .A(n643), .B(A[165]), .Z(n640) );
  XOR U736 ( .A(n643), .B(n644), .Z(DIFF[165]) );
  XOR U737 ( .A(B[165]), .B(A[165]), .Z(n644) );
  AND U738 ( .A(n645), .B(n646), .Z(n643) );
  NANDN U739 ( .A(B[164]), .B(n647), .Z(n646) );
  NANDN U740 ( .A(A[164]), .B(n648), .Z(n647) );
  NANDN U741 ( .A(n648), .B(A[164]), .Z(n645) );
  XOR U742 ( .A(n648), .B(n649), .Z(DIFF[164]) );
  XOR U743 ( .A(B[164]), .B(A[164]), .Z(n649) );
  AND U744 ( .A(n650), .B(n651), .Z(n648) );
  NANDN U745 ( .A(B[163]), .B(n652), .Z(n651) );
  NANDN U746 ( .A(A[163]), .B(n653), .Z(n652) );
  NANDN U747 ( .A(n653), .B(A[163]), .Z(n650) );
  XOR U748 ( .A(n653), .B(n654), .Z(DIFF[163]) );
  XOR U749 ( .A(B[163]), .B(A[163]), .Z(n654) );
  AND U750 ( .A(n655), .B(n656), .Z(n653) );
  NANDN U751 ( .A(B[162]), .B(n657), .Z(n656) );
  NANDN U752 ( .A(A[162]), .B(n658), .Z(n657) );
  NANDN U753 ( .A(n658), .B(A[162]), .Z(n655) );
  XOR U754 ( .A(n658), .B(n659), .Z(DIFF[162]) );
  XOR U755 ( .A(B[162]), .B(A[162]), .Z(n659) );
  AND U756 ( .A(n660), .B(n661), .Z(n658) );
  NANDN U757 ( .A(B[161]), .B(n662), .Z(n661) );
  NANDN U758 ( .A(A[161]), .B(n663), .Z(n662) );
  NANDN U759 ( .A(n663), .B(A[161]), .Z(n660) );
  XOR U760 ( .A(n663), .B(n664), .Z(DIFF[161]) );
  XOR U761 ( .A(B[161]), .B(A[161]), .Z(n664) );
  AND U762 ( .A(n665), .B(n666), .Z(n663) );
  NANDN U763 ( .A(B[160]), .B(n667), .Z(n666) );
  NANDN U764 ( .A(A[160]), .B(n668), .Z(n667) );
  NANDN U765 ( .A(n668), .B(A[160]), .Z(n665) );
  XOR U766 ( .A(n668), .B(n669), .Z(DIFF[160]) );
  XOR U767 ( .A(B[160]), .B(A[160]), .Z(n669) );
  AND U768 ( .A(n670), .B(n671), .Z(n668) );
  NANDN U769 ( .A(B[159]), .B(n672), .Z(n671) );
  NANDN U770 ( .A(A[159]), .B(n673), .Z(n672) );
  NANDN U771 ( .A(n673), .B(A[159]), .Z(n670) );
  XOR U772 ( .A(n674), .B(n675), .Z(DIFF[15]) );
  XOR U773 ( .A(B[15]), .B(A[15]), .Z(n675) );
  XOR U774 ( .A(n673), .B(n676), .Z(DIFF[159]) );
  XOR U775 ( .A(B[159]), .B(A[159]), .Z(n676) );
  AND U776 ( .A(n677), .B(n678), .Z(n673) );
  NANDN U777 ( .A(B[158]), .B(n679), .Z(n678) );
  NANDN U778 ( .A(A[158]), .B(n680), .Z(n679) );
  NANDN U779 ( .A(n680), .B(A[158]), .Z(n677) );
  XOR U780 ( .A(n680), .B(n681), .Z(DIFF[158]) );
  XOR U781 ( .A(B[158]), .B(A[158]), .Z(n681) );
  AND U782 ( .A(n682), .B(n683), .Z(n680) );
  NANDN U783 ( .A(B[157]), .B(n684), .Z(n683) );
  NANDN U784 ( .A(A[157]), .B(n685), .Z(n684) );
  NANDN U785 ( .A(n685), .B(A[157]), .Z(n682) );
  XOR U786 ( .A(n685), .B(n686), .Z(DIFF[157]) );
  XOR U787 ( .A(B[157]), .B(A[157]), .Z(n686) );
  AND U788 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U789 ( .A(B[156]), .B(n689), .Z(n688) );
  NANDN U790 ( .A(A[156]), .B(n690), .Z(n689) );
  NANDN U791 ( .A(n690), .B(A[156]), .Z(n687) );
  XOR U792 ( .A(n690), .B(n691), .Z(DIFF[156]) );
  XOR U793 ( .A(B[156]), .B(A[156]), .Z(n691) );
  AND U794 ( .A(n692), .B(n693), .Z(n690) );
  NANDN U795 ( .A(B[155]), .B(n694), .Z(n693) );
  NANDN U796 ( .A(A[155]), .B(n695), .Z(n694) );
  NANDN U797 ( .A(n695), .B(A[155]), .Z(n692) );
  XOR U798 ( .A(n695), .B(n696), .Z(DIFF[155]) );
  XOR U799 ( .A(B[155]), .B(A[155]), .Z(n696) );
  AND U800 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U801 ( .A(B[154]), .B(n699), .Z(n698) );
  NANDN U802 ( .A(A[154]), .B(n700), .Z(n699) );
  NANDN U803 ( .A(n700), .B(A[154]), .Z(n697) );
  XOR U804 ( .A(n700), .B(n701), .Z(DIFF[154]) );
  XOR U805 ( .A(B[154]), .B(A[154]), .Z(n701) );
  AND U806 ( .A(n702), .B(n703), .Z(n700) );
  NANDN U807 ( .A(B[153]), .B(n704), .Z(n703) );
  NANDN U808 ( .A(A[153]), .B(n705), .Z(n704) );
  NANDN U809 ( .A(n705), .B(A[153]), .Z(n702) );
  XOR U810 ( .A(n705), .B(n706), .Z(DIFF[153]) );
  XOR U811 ( .A(B[153]), .B(A[153]), .Z(n706) );
  AND U812 ( .A(n707), .B(n708), .Z(n705) );
  NANDN U813 ( .A(B[152]), .B(n709), .Z(n708) );
  NANDN U814 ( .A(A[152]), .B(n710), .Z(n709) );
  NANDN U815 ( .A(n710), .B(A[152]), .Z(n707) );
  XOR U816 ( .A(n710), .B(n711), .Z(DIFF[152]) );
  XOR U817 ( .A(B[152]), .B(A[152]), .Z(n711) );
  AND U818 ( .A(n712), .B(n713), .Z(n710) );
  NANDN U819 ( .A(B[151]), .B(n714), .Z(n713) );
  NANDN U820 ( .A(A[151]), .B(n715), .Z(n714) );
  NANDN U821 ( .A(n715), .B(A[151]), .Z(n712) );
  XOR U822 ( .A(n715), .B(n716), .Z(DIFF[151]) );
  XOR U823 ( .A(B[151]), .B(A[151]), .Z(n716) );
  AND U824 ( .A(n717), .B(n718), .Z(n715) );
  NANDN U825 ( .A(B[150]), .B(n719), .Z(n718) );
  NANDN U826 ( .A(A[150]), .B(n720), .Z(n719) );
  NANDN U827 ( .A(n720), .B(A[150]), .Z(n717) );
  XOR U828 ( .A(n720), .B(n721), .Z(DIFF[150]) );
  XOR U829 ( .A(B[150]), .B(A[150]), .Z(n721) );
  AND U830 ( .A(n722), .B(n723), .Z(n720) );
  NANDN U831 ( .A(B[149]), .B(n724), .Z(n723) );
  NANDN U832 ( .A(A[149]), .B(n725), .Z(n724) );
  NANDN U833 ( .A(n725), .B(A[149]), .Z(n722) );
  XOR U834 ( .A(n726), .B(n727), .Z(DIFF[14]) );
  XOR U835 ( .A(B[14]), .B(A[14]), .Z(n727) );
  XOR U836 ( .A(n725), .B(n728), .Z(DIFF[149]) );
  XOR U837 ( .A(B[149]), .B(A[149]), .Z(n728) );
  AND U838 ( .A(n729), .B(n730), .Z(n725) );
  NANDN U839 ( .A(B[148]), .B(n731), .Z(n730) );
  NANDN U840 ( .A(A[148]), .B(n732), .Z(n731) );
  NANDN U841 ( .A(n732), .B(A[148]), .Z(n729) );
  XOR U842 ( .A(n732), .B(n733), .Z(DIFF[148]) );
  XOR U843 ( .A(B[148]), .B(A[148]), .Z(n733) );
  AND U844 ( .A(n734), .B(n735), .Z(n732) );
  NANDN U845 ( .A(B[147]), .B(n736), .Z(n735) );
  NANDN U846 ( .A(A[147]), .B(n737), .Z(n736) );
  NANDN U847 ( .A(n737), .B(A[147]), .Z(n734) );
  XOR U848 ( .A(n737), .B(n738), .Z(DIFF[147]) );
  XOR U849 ( .A(B[147]), .B(A[147]), .Z(n738) );
  AND U850 ( .A(n739), .B(n740), .Z(n737) );
  NANDN U851 ( .A(B[146]), .B(n741), .Z(n740) );
  NANDN U852 ( .A(A[146]), .B(n742), .Z(n741) );
  NANDN U853 ( .A(n742), .B(A[146]), .Z(n739) );
  XOR U854 ( .A(n742), .B(n743), .Z(DIFF[146]) );
  XOR U855 ( .A(B[146]), .B(A[146]), .Z(n743) );
  AND U856 ( .A(n744), .B(n745), .Z(n742) );
  NANDN U857 ( .A(B[145]), .B(n746), .Z(n745) );
  NANDN U858 ( .A(A[145]), .B(n747), .Z(n746) );
  NANDN U859 ( .A(n747), .B(A[145]), .Z(n744) );
  XOR U860 ( .A(n747), .B(n748), .Z(DIFF[145]) );
  XOR U861 ( .A(B[145]), .B(A[145]), .Z(n748) );
  AND U862 ( .A(n749), .B(n750), .Z(n747) );
  NANDN U863 ( .A(B[144]), .B(n751), .Z(n750) );
  NANDN U864 ( .A(A[144]), .B(n752), .Z(n751) );
  NANDN U865 ( .A(n752), .B(A[144]), .Z(n749) );
  XOR U866 ( .A(n752), .B(n753), .Z(DIFF[144]) );
  XOR U867 ( .A(B[144]), .B(A[144]), .Z(n753) );
  AND U868 ( .A(n754), .B(n755), .Z(n752) );
  NANDN U869 ( .A(B[143]), .B(n756), .Z(n755) );
  NANDN U870 ( .A(A[143]), .B(n757), .Z(n756) );
  NANDN U871 ( .A(n757), .B(A[143]), .Z(n754) );
  XOR U872 ( .A(n757), .B(n758), .Z(DIFF[143]) );
  XOR U873 ( .A(B[143]), .B(A[143]), .Z(n758) );
  AND U874 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U875 ( .A(B[142]), .B(n761), .Z(n760) );
  NANDN U876 ( .A(A[142]), .B(n762), .Z(n761) );
  NANDN U877 ( .A(n762), .B(A[142]), .Z(n759) );
  XOR U878 ( .A(n762), .B(n763), .Z(DIFF[142]) );
  XOR U879 ( .A(B[142]), .B(A[142]), .Z(n763) );
  AND U880 ( .A(n764), .B(n765), .Z(n762) );
  NANDN U881 ( .A(B[141]), .B(n766), .Z(n765) );
  NANDN U882 ( .A(A[141]), .B(n767), .Z(n766) );
  NANDN U883 ( .A(n767), .B(A[141]), .Z(n764) );
  XOR U884 ( .A(n767), .B(n768), .Z(DIFF[141]) );
  XOR U885 ( .A(B[141]), .B(A[141]), .Z(n768) );
  AND U886 ( .A(n769), .B(n770), .Z(n767) );
  NANDN U887 ( .A(B[140]), .B(n771), .Z(n770) );
  NANDN U888 ( .A(A[140]), .B(n772), .Z(n771) );
  NANDN U889 ( .A(n772), .B(A[140]), .Z(n769) );
  XOR U890 ( .A(n772), .B(n773), .Z(DIFF[140]) );
  XOR U891 ( .A(B[140]), .B(A[140]), .Z(n773) );
  AND U892 ( .A(n774), .B(n775), .Z(n772) );
  NANDN U893 ( .A(B[139]), .B(n776), .Z(n775) );
  NANDN U894 ( .A(A[139]), .B(n777), .Z(n776) );
  NANDN U895 ( .A(n777), .B(A[139]), .Z(n774) );
  XOR U896 ( .A(n778), .B(n779), .Z(DIFF[13]) );
  XOR U897 ( .A(B[13]), .B(A[13]), .Z(n779) );
  XOR U898 ( .A(n777), .B(n780), .Z(DIFF[139]) );
  XOR U899 ( .A(B[139]), .B(A[139]), .Z(n780) );
  AND U900 ( .A(n781), .B(n782), .Z(n777) );
  NANDN U901 ( .A(B[138]), .B(n783), .Z(n782) );
  NANDN U902 ( .A(A[138]), .B(n784), .Z(n783) );
  NANDN U903 ( .A(n784), .B(A[138]), .Z(n781) );
  XOR U904 ( .A(n784), .B(n785), .Z(DIFF[138]) );
  XOR U905 ( .A(B[138]), .B(A[138]), .Z(n785) );
  AND U906 ( .A(n786), .B(n787), .Z(n784) );
  NANDN U907 ( .A(B[137]), .B(n788), .Z(n787) );
  NANDN U908 ( .A(A[137]), .B(n789), .Z(n788) );
  NANDN U909 ( .A(n789), .B(A[137]), .Z(n786) );
  XOR U910 ( .A(n789), .B(n790), .Z(DIFF[137]) );
  XOR U911 ( .A(B[137]), .B(A[137]), .Z(n790) );
  AND U912 ( .A(n791), .B(n792), .Z(n789) );
  NANDN U913 ( .A(B[136]), .B(n793), .Z(n792) );
  NANDN U914 ( .A(A[136]), .B(n794), .Z(n793) );
  NANDN U915 ( .A(n794), .B(A[136]), .Z(n791) );
  XOR U916 ( .A(n794), .B(n795), .Z(DIFF[136]) );
  XOR U917 ( .A(B[136]), .B(A[136]), .Z(n795) );
  AND U918 ( .A(n796), .B(n797), .Z(n794) );
  NANDN U919 ( .A(B[135]), .B(n798), .Z(n797) );
  NANDN U920 ( .A(A[135]), .B(n799), .Z(n798) );
  NANDN U921 ( .A(n799), .B(A[135]), .Z(n796) );
  XOR U922 ( .A(n799), .B(n800), .Z(DIFF[135]) );
  XOR U923 ( .A(B[135]), .B(A[135]), .Z(n800) );
  AND U924 ( .A(n801), .B(n802), .Z(n799) );
  NANDN U925 ( .A(B[134]), .B(n803), .Z(n802) );
  NANDN U926 ( .A(A[134]), .B(n804), .Z(n803) );
  NANDN U927 ( .A(n804), .B(A[134]), .Z(n801) );
  XOR U928 ( .A(n804), .B(n805), .Z(DIFF[134]) );
  XOR U929 ( .A(B[134]), .B(A[134]), .Z(n805) );
  AND U930 ( .A(n806), .B(n807), .Z(n804) );
  NANDN U931 ( .A(B[133]), .B(n808), .Z(n807) );
  NANDN U932 ( .A(A[133]), .B(n809), .Z(n808) );
  NANDN U933 ( .A(n809), .B(A[133]), .Z(n806) );
  XOR U934 ( .A(n809), .B(n810), .Z(DIFF[133]) );
  XOR U935 ( .A(B[133]), .B(A[133]), .Z(n810) );
  AND U936 ( .A(n811), .B(n812), .Z(n809) );
  NANDN U937 ( .A(B[132]), .B(n813), .Z(n812) );
  NANDN U938 ( .A(A[132]), .B(n814), .Z(n813) );
  NANDN U939 ( .A(n814), .B(A[132]), .Z(n811) );
  XOR U940 ( .A(n814), .B(n815), .Z(DIFF[132]) );
  XOR U941 ( .A(B[132]), .B(A[132]), .Z(n815) );
  AND U942 ( .A(n816), .B(n817), .Z(n814) );
  NANDN U943 ( .A(B[131]), .B(n818), .Z(n817) );
  NANDN U944 ( .A(A[131]), .B(n819), .Z(n818) );
  NANDN U945 ( .A(n819), .B(A[131]), .Z(n816) );
  XOR U946 ( .A(n819), .B(n820), .Z(DIFF[131]) );
  XOR U947 ( .A(B[131]), .B(A[131]), .Z(n820) );
  AND U948 ( .A(n821), .B(n822), .Z(n819) );
  NANDN U949 ( .A(B[130]), .B(n823), .Z(n822) );
  NANDN U950 ( .A(A[130]), .B(n824), .Z(n823) );
  NANDN U951 ( .A(n824), .B(A[130]), .Z(n821) );
  XOR U952 ( .A(n824), .B(n825), .Z(DIFF[130]) );
  XOR U953 ( .A(B[130]), .B(A[130]), .Z(n825) );
  AND U954 ( .A(n826), .B(n827), .Z(n824) );
  NANDN U955 ( .A(B[129]), .B(n828), .Z(n827) );
  NANDN U956 ( .A(A[129]), .B(n829), .Z(n828) );
  NANDN U957 ( .A(n829), .B(A[129]), .Z(n826) );
  XOR U958 ( .A(n830), .B(n831), .Z(DIFF[12]) );
  XOR U959 ( .A(B[12]), .B(A[12]), .Z(n831) );
  XOR U960 ( .A(n829), .B(n832), .Z(DIFF[129]) );
  XOR U961 ( .A(B[129]), .B(A[129]), .Z(n832) );
  AND U962 ( .A(n833), .B(n834), .Z(n829) );
  NANDN U963 ( .A(B[128]), .B(n835), .Z(n834) );
  NANDN U964 ( .A(A[128]), .B(n836), .Z(n835) );
  NANDN U965 ( .A(n836), .B(A[128]), .Z(n833) );
  XOR U966 ( .A(n836), .B(n837), .Z(DIFF[128]) );
  XOR U967 ( .A(B[128]), .B(A[128]), .Z(n837) );
  AND U968 ( .A(n838), .B(n839), .Z(n836) );
  NANDN U969 ( .A(B[127]), .B(n840), .Z(n839) );
  NANDN U970 ( .A(A[127]), .B(n841), .Z(n840) );
  NANDN U971 ( .A(n841), .B(A[127]), .Z(n838) );
  XOR U972 ( .A(n841), .B(n842), .Z(DIFF[127]) );
  XOR U973 ( .A(B[127]), .B(A[127]), .Z(n842) );
  AND U974 ( .A(n843), .B(n844), .Z(n841) );
  NANDN U975 ( .A(B[126]), .B(n845), .Z(n844) );
  NANDN U976 ( .A(A[126]), .B(n846), .Z(n845) );
  NANDN U977 ( .A(n846), .B(A[126]), .Z(n843) );
  XOR U978 ( .A(n846), .B(n847), .Z(DIFF[126]) );
  XOR U979 ( .A(B[126]), .B(A[126]), .Z(n847) );
  AND U980 ( .A(n848), .B(n849), .Z(n846) );
  NANDN U981 ( .A(B[125]), .B(n850), .Z(n849) );
  NANDN U982 ( .A(A[125]), .B(n851), .Z(n850) );
  NANDN U983 ( .A(n851), .B(A[125]), .Z(n848) );
  XOR U984 ( .A(n851), .B(n852), .Z(DIFF[125]) );
  XOR U985 ( .A(B[125]), .B(A[125]), .Z(n852) );
  AND U986 ( .A(n853), .B(n854), .Z(n851) );
  NANDN U987 ( .A(B[124]), .B(n855), .Z(n854) );
  NANDN U988 ( .A(A[124]), .B(n856), .Z(n855) );
  NANDN U989 ( .A(n856), .B(A[124]), .Z(n853) );
  XOR U990 ( .A(n856), .B(n857), .Z(DIFF[124]) );
  XOR U991 ( .A(B[124]), .B(A[124]), .Z(n857) );
  AND U992 ( .A(n858), .B(n859), .Z(n856) );
  NANDN U993 ( .A(B[123]), .B(n860), .Z(n859) );
  NANDN U994 ( .A(A[123]), .B(n861), .Z(n860) );
  NANDN U995 ( .A(n861), .B(A[123]), .Z(n858) );
  XOR U996 ( .A(n861), .B(n862), .Z(DIFF[123]) );
  XOR U997 ( .A(B[123]), .B(A[123]), .Z(n862) );
  AND U998 ( .A(n863), .B(n864), .Z(n861) );
  NANDN U999 ( .A(B[122]), .B(n865), .Z(n864) );
  NANDN U1000 ( .A(A[122]), .B(n866), .Z(n865) );
  NANDN U1001 ( .A(n866), .B(A[122]), .Z(n863) );
  XOR U1002 ( .A(n866), .B(n867), .Z(DIFF[122]) );
  XOR U1003 ( .A(B[122]), .B(A[122]), .Z(n867) );
  AND U1004 ( .A(n868), .B(n869), .Z(n866) );
  NANDN U1005 ( .A(B[121]), .B(n870), .Z(n869) );
  NANDN U1006 ( .A(A[121]), .B(n871), .Z(n870) );
  NANDN U1007 ( .A(n871), .B(A[121]), .Z(n868) );
  XOR U1008 ( .A(n871), .B(n872), .Z(DIFF[121]) );
  XOR U1009 ( .A(B[121]), .B(A[121]), .Z(n872) );
  AND U1010 ( .A(n873), .B(n874), .Z(n871) );
  NANDN U1011 ( .A(B[120]), .B(n875), .Z(n874) );
  NANDN U1012 ( .A(A[120]), .B(n876), .Z(n875) );
  NANDN U1013 ( .A(n876), .B(A[120]), .Z(n873) );
  XOR U1014 ( .A(n876), .B(n877), .Z(DIFF[120]) );
  XOR U1015 ( .A(B[120]), .B(A[120]), .Z(n877) );
  AND U1016 ( .A(n878), .B(n879), .Z(n876) );
  NANDN U1017 ( .A(B[119]), .B(n880), .Z(n879) );
  NANDN U1018 ( .A(A[119]), .B(n881), .Z(n880) );
  NANDN U1019 ( .A(n881), .B(A[119]), .Z(n878) );
  XOR U1020 ( .A(n882), .B(n883), .Z(DIFF[11]) );
  XOR U1021 ( .A(B[11]), .B(A[11]), .Z(n883) );
  XOR U1022 ( .A(n881), .B(n884), .Z(DIFF[119]) );
  XOR U1023 ( .A(B[119]), .B(A[119]), .Z(n884) );
  AND U1024 ( .A(n885), .B(n886), .Z(n881) );
  NANDN U1025 ( .A(B[118]), .B(n887), .Z(n886) );
  NANDN U1026 ( .A(A[118]), .B(n888), .Z(n887) );
  NANDN U1027 ( .A(n888), .B(A[118]), .Z(n885) );
  XOR U1028 ( .A(n888), .B(n889), .Z(DIFF[118]) );
  XOR U1029 ( .A(B[118]), .B(A[118]), .Z(n889) );
  AND U1030 ( .A(n890), .B(n891), .Z(n888) );
  NANDN U1031 ( .A(B[117]), .B(n892), .Z(n891) );
  NANDN U1032 ( .A(A[117]), .B(n893), .Z(n892) );
  NANDN U1033 ( .A(n893), .B(A[117]), .Z(n890) );
  XOR U1034 ( .A(n893), .B(n894), .Z(DIFF[117]) );
  XOR U1035 ( .A(B[117]), .B(A[117]), .Z(n894) );
  AND U1036 ( .A(n895), .B(n896), .Z(n893) );
  NANDN U1037 ( .A(B[116]), .B(n897), .Z(n896) );
  NANDN U1038 ( .A(A[116]), .B(n898), .Z(n897) );
  NANDN U1039 ( .A(n898), .B(A[116]), .Z(n895) );
  XOR U1040 ( .A(n898), .B(n899), .Z(DIFF[116]) );
  XOR U1041 ( .A(B[116]), .B(A[116]), .Z(n899) );
  AND U1042 ( .A(n900), .B(n901), .Z(n898) );
  NANDN U1043 ( .A(B[115]), .B(n902), .Z(n901) );
  NANDN U1044 ( .A(A[115]), .B(n903), .Z(n902) );
  NANDN U1045 ( .A(n903), .B(A[115]), .Z(n900) );
  XOR U1046 ( .A(n903), .B(n904), .Z(DIFF[115]) );
  XOR U1047 ( .A(B[115]), .B(A[115]), .Z(n904) );
  AND U1048 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U1049 ( .A(B[114]), .B(n907), .Z(n906) );
  NANDN U1050 ( .A(A[114]), .B(n908), .Z(n907) );
  NANDN U1051 ( .A(n908), .B(A[114]), .Z(n905) );
  XOR U1052 ( .A(n908), .B(n909), .Z(DIFF[114]) );
  XOR U1053 ( .A(B[114]), .B(A[114]), .Z(n909) );
  AND U1054 ( .A(n910), .B(n911), .Z(n908) );
  NANDN U1055 ( .A(B[113]), .B(n912), .Z(n911) );
  NANDN U1056 ( .A(A[113]), .B(n913), .Z(n912) );
  NANDN U1057 ( .A(n913), .B(A[113]), .Z(n910) );
  XOR U1058 ( .A(n913), .B(n914), .Z(DIFF[113]) );
  XOR U1059 ( .A(B[113]), .B(A[113]), .Z(n914) );
  AND U1060 ( .A(n915), .B(n916), .Z(n913) );
  NANDN U1061 ( .A(B[112]), .B(n917), .Z(n916) );
  NANDN U1062 ( .A(A[112]), .B(n918), .Z(n917) );
  NANDN U1063 ( .A(n918), .B(A[112]), .Z(n915) );
  XOR U1064 ( .A(n918), .B(n919), .Z(DIFF[112]) );
  XOR U1065 ( .A(B[112]), .B(A[112]), .Z(n919) );
  AND U1066 ( .A(n920), .B(n921), .Z(n918) );
  NANDN U1067 ( .A(B[111]), .B(n922), .Z(n921) );
  NANDN U1068 ( .A(A[111]), .B(n923), .Z(n922) );
  NANDN U1069 ( .A(n923), .B(A[111]), .Z(n920) );
  XOR U1070 ( .A(n923), .B(n924), .Z(DIFF[111]) );
  XOR U1071 ( .A(B[111]), .B(A[111]), .Z(n924) );
  AND U1072 ( .A(n925), .B(n926), .Z(n923) );
  NANDN U1073 ( .A(B[110]), .B(n927), .Z(n926) );
  NANDN U1074 ( .A(A[110]), .B(n928), .Z(n927) );
  NANDN U1075 ( .A(n928), .B(A[110]), .Z(n925) );
  XOR U1076 ( .A(n928), .B(n929), .Z(DIFF[110]) );
  XOR U1077 ( .A(B[110]), .B(A[110]), .Z(n929) );
  AND U1078 ( .A(n930), .B(n931), .Z(n928) );
  NANDN U1079 ( .A(B[109]), .B(n932), .Z(n931) );
  NANDN U1080 ( .A(A[109]), .B(n933), .Z(n932) );
  NANDN U1081 ( .A(n933), .B(A[109]), .Z(n930) );
  XOR U1082 ( .A(n934), .B(n935), .Z(DIFF[10]) );
  XOR U1083 ( .A(B[10]), .B(A[10]), .Z(n935) );
  XOR U1084 ( .A(n933), .B(n936), .Z(DIFF[109]) );
  XOR U1085 ( .A(B[109]), .B(A[109]), .Z(n936) );
  AND U1086 ( .A(n937), .B(n938), .Z(n933) );
  NANDN U1087 ( .A(B[108]), .B(n939), .Z(n938) );
  NANDN U1088 ( .A(A[108]), .B(n940), .Z(n939) );
  NANDN U1089 ( .A(n940), .B(A[108]), .Z(n937) );
  XOR U1090 ( .A(n940), .B(n941), .Z(DIFF[108]) );
  XOR U1091 ( .A(B[108]), .B(A[108]), .Z(n941) );
  AND U1092 ( .A(n942), .B(n943), .Z(n940) );
  NANDN U1093 ( .A(B[107]), .B(n944), .Z(n943) );
  NANDN U1094 ( .A(A[107]), .B(n945), .Z(n944) );
  NANDN U1095 ( .A(n945), .B(A[107]), .Z(n942) );
  XOR U1096 ( .A(n945), .B(n946), .Z(DIFF[107]) );
  XOR U1097 ( .A(B[107]), .B(A[107]), .Z(n946) );
  AND U1098 ( .A(n947), .B(n948), .Z(n945) );
  NANDN U1099 ( .A(B[106]), .B(n949), .Z(n948) );
  NANDN U1100 ( .A(A[106]), .B(n950), .Z(n949) );
  NANDN U1101 ( .A(n950), .B(A[106]), .Z(n947) );
  XOR U1102 ( .A(n950), .B(n951), .Z(DIFF[106]) );
  XOR U1103 ( .A(B[106]), .B(A[106]), .Z(n951) );
  AND U1104 ( .A(n952), .B(n953), .Z(n950) );
  NANDN U1105 ( .A(B[105]), .B(n954), .Z(n953) );
  NANDN U1106 ( .A(A[105]), .B(n955), .Z(n954) );
  NANDN U1107 ( .A(n955), .B(A[105]), .Z(n952) );
  XOR U1108 ( .A(n955), .B(n956), .Z(DIFF[105]) );
  XOR U1109 ( .A(B[105]), .B(A[105]), .Z(n956) );
  AND U1110 ( .A(n957), .B(n958), .Z(n955) );
  NANDN U1111 ( .A(B[104]), .B(n959), .Z(n958) );
  NANDN U1112 ( .A(A[104]), .B(n960), .Z(n959) );
  NANDN U1113 ( .A(n960), .B(A[104]), .Z(n957) );
  XOR U1114 ( .A(n960), .B(n961), .Z(DIFF[104]) );
  XOR U1115 ( .A(B[104]), .B(A[104]), .Z(n961) );
  AND U1116 ( .A(n962), .B(n963), .Z(n960) );
  NANDN U1117 ( .A(B[103]), .B(n964), .Z(n963) );
  NANDN U1118 ( .A(A[103]), .B(n965), .Z(n964) );
  NANDN U1119 ( .A(n965), .B(A[103]), .Z(n962) );
  XOR U1120 ( .A(n965), .B(n966), .Z(DIFF[103]) );
  XOR U1121 ( .A(B[103]), .B(A[103]), .Z(n966) );
  AND U1122 ( .A(n967), .B(n968), .Z(n965) );
  NANDN U1123 ( .A(B[102]), .B(n969), .Z(n968) );
  NANDN U1124 ( .A(A[102]), .B(n970), .Z(n969) );
  NANDN U1125 ( .A(n970), .B(A[102]), .Z(n967) );
  XOR U1126 ( .A(n970), .B(n971), .Z(DIFF[102]) );
  XOR U1127 ( .A(B[102]), .B(A[102]), .Z(n971) );
  AND U1128 ( .A(n972), .B(n973), .Z(n970) );
  NANDN U1129 ( .A(B[101]), .B(n974), .Z(n973) );
  NANDN U1130 ( .A(A[101]), .B(n975), .Z(n974) );
  NANDN U1131 ( .A(n975), .B(A[101]), .Z(n972) );
  XOR U1132 ( .A(n975), .B(n976), .Z(DIFF[101]) );
  XOR U1133 ( .A(B[101]), .B(A[101]), .Z(n976) );
  AND U1134 ( .A(n977), .B(n978), .Z(n975) );
  NANDN U1135 ( .A(B[100]), .B(n979), .Z(n978) );
  NANDN U1136 ( .A(A[100]), .B(n980), .Z(n979) );
  NANDN U1137 ( .A(n980), .B(A[100]), .Z(n977) );
  XOR U1138 ( .A(n980), .B(n981), .Z(DIFF[100]) );
  XOR U1139 ( .A(B[100]), .B(A[100]), .Z(n981) );
  AND U1140 ( .A(n982), .B(n983), .Z(n980) );
  NANDN U1141 ( .A(B[99]), .B(n984), .Z(n983) );
  OR U1142 ( .A(n5), .B(A[99]), .Z(n984) );
  NAND U1143 ( .A(A[99]), .B(n5), .Z(n982) );
  NAND U1144 ( .A(n985), .B(n986), .Z(n5) );
  NANDN U1145 ( .A(B[98]), .B(n987), .Z(n986) );
  NANDN U1146 ( .A(A[98]), .B(n7), .Z(n987) );
  NANDN U1147 ( .A(n7), .B(A[98]), .Z(n985) );
  AND U1148 ( .A(n988), .B(n989), .Z(n7) );
  NANDN U1149 ( .A(B[97]), .B(n990), .Z(n989) );
  NANDN U1150 ( .A(A[97]), .B(n9), .Z(n990) );
  NANDN U1151 ( .A(n9), .B(A[97]), .Z(n988) );
  AND U1152 ( .A(n991), .B(n992), .Z(n9) );
  NANDN U1153 ( .A(B[96]), .B(n993), .Z(n992) );
  NANDN U1154 ( .A(A[96]), .B(n11), .Z(n993) );
  NANDN U1155 ( .A(n11), .B(A[96]), .Z(n991) );
  AND U1156 ( .A(n994), .B(n995), .Z(n11) );
  NANDN U1157 ( .A(B[95]), .B(n996), .Z(n995) );
  NANDN U1158 ( .A(A[95]), .B(n13), .Z(n996) );
  NANDN U1159 ( .A(n13), .B(A[95]), .Z(n994) );
  AND U1160 ( .A(n997), .B(n998), .Z(n13) );
  NANDN U1161 ( .A(B[94]), .B(n999), .Z(n998) );
  NANDN U1162 ( .A(A[94]), .B(n15), .Z(n999) );
  NANDN U1163 ( .A(n15), .B(A[94]), .Z(n997) );
  AND U1164 ( .A(n1000), .B(n1001), .Z(n15) );
  NANDN U1165 ( .A(B[93]), .B(n1002), .Z(n1001) );
  NANDN U1166 ( .A(A[93]), .B(n17), .Z(n1002) );
  NANDN U1167 ( .A(n17), .B(A[93]), .Z(n1000) );
  AND U1168 ( .A(n1003), .B(n1004), .Z(n17) );
  NANDN U1169 ( .A(B[92]), .B(n1005), .Z(n1004) );
  NANDN U1170 ( .A(A[92]), .B(n19), .Z(n1005) );
  NANDN U1171 ( .A(n19), .B(A[92]), .Z(n1003) );
  AND U1172 ( .A(n1006), .B(n1007), .Z(n19) );
  NANDN U1173 ( .A(B[91]), .B(n1008), .Z(n1007) );
  NANDN U1174 ( .A(A[91]), .B(n21), .Z(n1008) );
  NANDN U1175 ( .A(n21), .B(A[91]), .Z(n1006) );
  AND U1176 ( .A(n1009), .B(n1010), .Z(n21) );
  NANDN U1177 ( .A(B[90]), .B(n1011), .Z(n1010) );
  NANDN U1178 ( .A(A[90]), .B(n23), .Z(n1011) );
  NANDN U1179 ( .A(n23), .B(A[90]), .Z(n1009) );
  AND U1180 ( .A(n1012), .B(n1013), .Z(n23) );
  NANDN U1181 ( .A(B[89]), .B(n1014), .Z(n1013) );
  NANDN U1182 ( .A(A[89]), .B(n27), .Z(n1014) );
  NANDN U1183 ( .A(n27), .B(A[89]), .Z(n1012) );
  AND U1184 ( .A(n1015), .B(n1016), .Z(n27) );
  NANDN U1185 ( .A(B[88]), .B(n1017), .Z(n1016) );
  NANDN U1186 ( .A(A[88]), .B(n29), .Z(n1017) );
  NANDN U1187 ( .A(n29), .B(A[88]), .Z(n1015) );
  AND U1188 ( .A(n1018), .B(n1019), .Z(n29) );
  NANDN U1189 ( .A(B[87]), .B(n1020), .Z(n1019) );
  NANDN U1190 ( .A(A[87]), .B(n31), .Z(n1020) );
  NANDN U1191 ( .A(n31), .B(A[87]), .Z(n1018) );
  AND U1192 ( .A(n1021), .B(n1022), .Z(n31) );
  NANDN U1193 ( .A(B[86]), .B(n1023), .Z(n1022) );
  NANDN U1194 ( .A(A[86]), .B(n33), .Z(n1023) );
  NANDN U1195 ( .A(n33), .B(A[86]), .Z(n1021) );
  AND U1196 ( .A(n1024), .B(n1025), .Z(n33) );
  NANDN U1197 ( .A(B[85]), .B(n1026), .Z(n1025) );
  NANDN U1198 ( .A(A[85]), .B(n35), .Z(n1026) );
  NANDN U1199 ( .A(n35), .B(A[85]), .Z(n1024) );
  AND U1200 ( .A(n1027), .B(n1028), .Z(n35) );
  NANDN U1201 ( .A(B[84]), .B(n1029), .Z(n1028) );
  NANDN U1202 ( .A(A[84]), .B(n37), .Z(n1029) );
  NANDN U1203 ( .A(n37), .B(A[84]), .Z(n1027) );
  AND U1204 ( .A(n1030), .B(n1031), .Z(n37) );
  NANDN U1205 ( .A(B[83]), .B(n1032), .Z(n1031) );
  NANDN U1206 ( .A(A[83]), .B(n39), .Z(n1032) );
  NANDN U1207 ( .A(n39), .B(A[83]), .Z(n1030) );
  AND U1208 ( .A(n1033), .B(n1034), .Z(n39) );
  NANDN U1209 ( .A(B[82]), .B(n1035), .Z(n1034) );
  NANDN U1210 ( .A(A[82]), .B(n41), .Z(n1035) );
  NANDN U1211 ( .A(n41), .B(A[82]), .Z(n1033) );
  AND U1212 ( .A(n1036), .B(n1037), .Z(n41) );
  NANDN U1213 ( .A(B[81]), .B(n1038), .Z(n1037) );
  NANDN U1214 ( .A(A[81]), .B(n43), .Z(n1038) );
  NANDN U1215 ( .A(n43), .B(A[81]), .Z(n1036) );
  AND U1216 ( .A(n1039), .B(n1040), .Z(n43) );
  NANDN U1217 ( .A(B[80]), .B(n1041), .Z(n1040) );
  NANDN U1218 ( .A(A[80]), .B(n45), .Z(n1041) );
  NANDN U1219 ( .A(n45), .B(A[80]), .Z(n1039) );
  AND U1220 ( .A(n1042), .B(n1043), .Z(n45) );
  NANDN U1221 ( .A(B[79]), .B(n1044), .Z(n1043) );
  NANDN U1222 ( .A(A[79]), .B(n49), .Z(n1044) );
  NANDN U1223 ( .A(n49), .B(A[79]), .Z(n1042) );
  AND U1224 ( .A(n1045), .B(n1046), .Z(n49) );
  NANDN U1225 ( .A(B[78]), .B(n1047), .Z(n1046) );
  NANDN U1226 ( .A(A[78]), .B(n51), .Z(n1047) );
  NANDN U1227 ( .A(n51), .B(A[78]), .Z(n1045) );
  AND U1228 ( .A(n1048), .B(n1049), .Z(n51) );
  NANDN U1229 ( .A(B[77]), .B(n1050), .Z(n1049) );
  NANDN U1230 ( .A(A[77]), .B(n53), .Z(n1050) );
  NANDN U1231 ( .A(n53), .B(A[77]), .Z(n1048) );
  AND U1232 ( .A(n1051), .B(n1052), .Z(n53) );
  NANDN U1233 ( .A(B[76]), .B(n1053), .Z(n1052) );
  NANDN U1234 ( .A(A[76]), .B(n55), .Z(n1053) );
  NANDN U1235 ( .A(n55), .B(A[76]), .Z(n1051) );
  AND U1236 ( .A(n1054), .B(n1055), .Z(n55) );
  NANDN U1237 ( .A(B[75]), .B(n1056), .Z(n1055) );
  NANDN U1238 ( .A(A[75]), .B(n57), .Z(n1056) );
  NANDN U1239 ( .A(n57), .B(A[75]), .Z(n1054) );
  AND U1240 ( .A(n1057), .B(n1058), .Z(n57) );
  NANDN U1241 ( .A(B[74]), .B(n1059), .Z(n1058) );
  NANDN U1242 ( .A(A[74]), .B(n59), .Z(n1059) );
  NANDN U1243 ( .A(n59), .B(A[74]), .Z(n1057) );
  AND U1244 ( .A(n1060), .B(n1061), .Z(n59) );
  NANDN U1245 ( .A(B[73]), .B(n1062), .Z(n1061) );
  NANDN U1246 ( .A(A[73]), .B(n61), .Z(n1062) );
  NANDN U1247 ( .A(n61), .B(A[73]), .Z(n1060) );
  AND U1248 ( .A(n1063), .B(n1064), .Z(n61) );
  NANDN U1249 ( .A(B[72]), .B(n1065), .Z(n1064) );
  NANDN U1250 ( .A(A[72]), .B(n63), .Z(n1065) );
  NANDN U1251 ( .A(n63), .B(A[72]), .Z(n1063) );
  AND U1252 ( .A(n1066), .B(n1067), .Z(n63) );
  NANDN U1253 ( .A(B[71]), .B(n1068), .Z(n1067) );
  NANDN U1254 ( .A(A[71]), .B(n65), .Z(n1068) );
  NANDN U1255 ( .A(n65), .B(A[71]), .Z(n1066) );
  AND U1256 ( .A(n1069), .B(n1070), .Z(n65) );
  NANDN U1257 ( .A(B[70]), .B(n1071), .Z(n1070) );
  NANDN U1258 ( .A(A[70]), .B(n67), .Z(n1071) );
  NANDN U1259 ( .A(n67), .B(A[70]), .Z(n1069) );
  AND U1260 ( .A(n1072), .B(n1073), .Z(n67) );
  NANDN U1261 ( .A(B[69]), .B(n1074), .Z(n1073) );
  NANDN U1262 ( .A(A[69]), .B(n71), .Z(n1074) );
  NANDN U1263 ( .A(n71), .B(A[69]), .Z(n1072) );
  AND U1264 ( .A(n1075), .B(n1076), .Z(n71) );
  NANDN U1265 ( .A(B[68]), .B(n1077), .Z(n1076) );
  NANDN U1266 ( .A(A[68]), .B(n73), .Z(n1077) );
  NANDN U1267 ( .A(n73), .B(A[68]), .Z(n1075) );
  AND U1268 ( .A(n1078), .B(n1079), .Z(n73) );
  NANDN U1269 ( .A(B[67]), .B(n1080), .Z(n1079) );
  NANDN U1270 ( .A(A[67]), .B(n75), .Z(n1080) );
  NANDN U1271 ( .A(n75), .B(A[67]), .Z(n1078) );
  AND U1272 ( .A(n1081), .B(n1082), .Z(n75) );
  NANDN U1273 ( .A(B[66]), .B(n1083), .Z(n1082) );
  NANDN U1274 ( .A(A[66]), .B(n77), .Z(n1083) );
  NANDN U1275 ( .A(n77), .B(A[66]), .Z(n1081) );
  AND U1276 ( .A(n1084), .B(n1085), .Z(n77) );
  NANDN U1277 ( .A(B[65]), .B(n1086), .Z(n1085) );
  NANDN U1278 ( .A(A[65]), .B(n79), .Z(n1086) );
  NANDN U1279 ( .A(n79), .B(A[65]), .Z(n1084) );
  AND U1280 ( .A(n1087), .B(n1088), .Z(n79) );
  NANDN U1281 ( .A(B[64]), .B(n1089), .Z(n1088) );
  NANDN U1282 ( .A(A[64]), .B(n81), .Z(n1089) );
  NANDN U1283 ( .A(n81), .B(A[64]), .Z(n1087) );
  AND U1284 ( .A(n1090), .B(n1091), .Z(n81) );
  NANDN U1285 ( .A(B[63]), .B(n1092), .Z(n1091) );
  NANDN U1286 ( .A(A[63]), .B(n83), .Z(n1092) );
  NANDN U1287 ( .A(n83), .B(A[63]), .Z(n1090) );
  AND U1288 ( .A(n1093), .B(n1094), .Z(n83) );
  NANDN U1289 ( .A(B[62]), .B(n1095), .Z(n1094) );
  NANDN U1290 ( .A(A[62]), .B(n85), .Z(n1095) );
  NANDN U1291 ( .A(n85), .B(A[62]), .Z(n1093) );
  AND U1292 ( .A(n1096), .B(n1097), .Z(n85) );
  NANDN U1293 ( .A(B[61]), .B(n1098), .Z(n1097) );
  NANDN U1294 ( .A(A[61]), .B(n87), .Z(n1098) );
  NANDN U1295 ( .A(n87), .B(A[61]), .Z(n1096) );
  AND U1296 ( .A(n1099), .B(n1100), .Z(n87) );
  NANDN U1297 ( .A(B[60]), .B(n1101), .Z(n1100) );
  NANDN U1298 ( .A(A[60]), .B(n89), .Z(n1101) );
  NANDN U1299 ( .A(n89), .B(A[60]), .Z(n1099) );
  AND U1300 ( .A(n1102), .B(n1103), .Z(n89) );
  NANDN U1301 ( .A(B[59]), .B(n1104), .Z(n1103) );
  NANDN U1302 ( .A(A[59]), .B(n93), .Z(n1104) );
  NANDN U1303 ( .A(n93), .B(A[59]), .Z(n1102) );
  AND U1304 ( .A(n1105), .B(n1106), .Z(n93) );
  NANDN U1305 ( .A(B[58]), .B(n1107), .Z(n1106) );
  NANDN U1306 ( .A(A[58]), .B(n95), .Z(n1107) );
  NANDN U1307 ( .A(n95), .B(A[58]), .Z(n1105) );
  AND U1308 ( .A(n1108), .B(n1109), .Z(n95) );
  NANDN U1309 ( .A(B[57]), .B(n1110), .Z(n1109) );
  NANDN U1310 ( .A(A[57]), .B(n97), .Z(n1110) );
  NANDN U1311 ( .A(n97), .B(A[57]), .Z(n1108) );
  AND U1312 ( .A(n1111), .B(n1112), .Z(n97) );
  NANDN U1313 ( .A(B[56]), .B(n1113), .Z(n1112) );
  NANDN U1314 ( .A(A[56]), .B(n99), .Z(n1113) );
  NANDN U1315 ( .A(n99), .B(A[56]), .Z(n1111) );
  AND U1316 ( .A(n1114), .B(n1115), .Z(n99) );
  NANDN U1317 ( .A(B[55]), .B(n1116), .Z(n1115) );
  NANDN U1318 ( .A(A[55]), .B(n101), .Z(n1116) );
  NANDN U1319 ( .A(n101), .B(A[55]), .Z(n1114) );
  AND U1320 ( .A(n1117), .B(n1118), .Z(n101) );
  NANDN U1321 ( .A(B[54]), .B(n1119), .Z(n1118) );
  NANDN U1322 ( .A(A[54]), .B(n103), .Z(n1119) );
  NANDN U1323 ( .A(n103), .B(A[54]), .Z(n1117) );
  AND U1324 ( .A(n1120), .B(n1121), .Z(n103) );
  NANDN U1325 ( .A(B[53]), .B(n1122), .Z(n1121) );
  NANDN U1326 ( .A(A[53]), .B(n105), .Z(n1122) );
  NANDN U1327 ( .A(n105), .B(A[53]), .Z(n1120) );
  AND U1328 ( .A(n1123), .B(n1124), .Z(n105) );
  NANDN U1329 ( .A(B[52]), .B(n1125), .Z(n1124) );
  NANDN U1330 ( .A(A[52]), .B(n107), .Z(n1125) );
  NANDN U1331 ( .A(n107), .B(A[52]), .Z(n1123) );
  AND U1332 ( .A(n1126), .B(n1127), .Z(n107) );
  NANDN U1333 ( .A(B[51]), .B(n1128), .Z(n1127) );
  NANDN U1334 ( .A(A[51]), .B(n109), .Z(n1128) );
  NANDN U1335 ( .A(n109), .B(A[51]), .Z(n1126) );
  AND U1336 ( .A(n1129), .B(n1130), .Z(n109) );
  NANDN U1337 ( .A(B[50]), .B(n1131), .Z(n1130) );
  NANDN U1338 ( .A(A[50]), .B(n111), .Z(n1131) );
  NANDN U1339 ( .A(n111), .B(A[50]), .Z(n1129) );
  AND U1340 ( .A(n1132), .B(n1133), .Z(n111) );
  NANDN U1341 ( .A(B[49]), .B(n1134), .Z(n1133) );
  NANDN U1342 ( .A(A[49]), .B(n115), .Z(n1134) );
  NANDN U1343 ( .A(n115), .B(A[49]), .Z(n1132) );
  AND U1344 ( .A(n1135), .B(n1136), .Z(n115) );
  NANDN U1345 ( .A(B[48]), .B(n1137), .Z(n1136) );
  NANDN U1346 ( .A(A[48]), .B(n117), .Z(n1137) );
  NANDN U1347 ( .A(n117), .B(A[48]), .Z(n1135) );
  AND U1348 ( .A(n1138), .B(n1139), .Z(n117) );
  NANDN U1349 ( .A(B[47]), .B(n1140), .Z(n1139) );
  NANDN U1350 ( .A(A[47]), .B(n119), .Z(n1140) );
  NANDN U1351 ( .A(n119), .B(A[47]), .Z(n1138) );
  AND U1352 ( .A(n1141), .B(n1142), .Z(n119) );
  NANDN U1353 ( .A(B[46]), .B(n1143), .Z(n1142) );
  NANDN U1354 ( .A(A[46]), .B(n121), .Z(n1143) );
  NANDN U1355 ( .A(n121), .B(A[46]), .Z(n1141) );
  AND U1356 ( .A(n1144), .B(n1145), .Z(n121) );
  NANDN U1357 ( .A(B[45]), .B(n1146), .Z(n1145) );
  NANDN U1358 ( .A(A[45]), .B(n123), .Z(n1146) );
  NANDN U1359 ( .A(n123), .B(A[45]), .Z(n1144) );
  AND U1360 ( .A(n1147), .B(n1148), .Z(n123) );
  NANDN U1361 ( .A(B[44]), .B(n1149), .Z(n1148) );
  NANDN U1362 ( .A(A[44]), .B(n125), .Z(n1149) );
  NANDN U1363 ( .A(n125), .B(A[44]), .Z(n1147) );
  AND U1364 ( .A(n1150), .B(n1151), .Z(n125) );
  NANDN U1365 ( .A(B[43]), .B(n1152), .Z(n1151) );
  NANDN U1366 ( .A(A[43]), .B(n127), .Z(n1152) );
  NANDN U1367 ( .A(n127), .B(A[43]), .Z(n1150) );
  AND U1368 ( .A(n1153), .B(n1154), .Z(n127) );
  NANDN U1369 ( .A(B[42]), .B(n1155), .Z(n1154) );
  NANDN U1370 ( .A(A[42]), .B(n129), .Z(n1155) );
  NANDN U1371 ( .A(n129), .B(A[42]), .Z(n1153) );
  AND U1372 ( .A(n1156), .B(n1157), .Z(n129) );
  NANDN U1373 ( .A(B[41]), .B(n1158), .Z(n1157) );
  NANDN U1374 ( .A(A[41]), .B(n131), .Z(n1158) );
  NANDN U1375 ( .A(n131), .B(A[41]), .Z(n1156) );
  AND U1376 ( .A(n1159), .B(n1160), .Z(n131) );
  NANDN U1377 ( .A(B[40]), .B(n1161), .Z(n1160) );
  NANDN U1378 ( .A(A[40]), .B(n133), .Z(n1161) );
  NANDN U1379 ( .A(n133), .B(A[40]), .Z(n1159) );
  AND U1380 ( .A(n1162), .B(n1163), .Z(n133) );
  NANDN U1381 ( .A(B[39]), .B(n1164), .Z(n1163) );
  NANDN U1382 ( .A(A[39]), .B(n137), .Z(n1164) );
  NANDN U1383 ( .A(n137), .B(A[39]), .Z(n1162) );
  AND U1384 ( .A(n1165), .B(n1166), .Z(n137) );
  NANDN U1385 ( .A(B[38]), .B(n1167), .Z(n1166) );
  NANDN U1386 ( .A(A[38]), .B(n139), .Z(n1167) );
  NANDN U1387 ( .A(n139), .B(A[38]), .Z(n1165) );
  AND U1388 ( .A(n1168), .B(n1169), .Z(n139) );
  NANDN U1389 ( .A(B[37]), .B(n1170), .Z(n1169) );
  NANDN U1390 ( .A(A[37]), .B(n141), .Z(n1170) );
  NANDN U1391 ( .A(n141), .B(A[37]), .Z(n1168) );
  AND U1392 ( .A(n1171), .B(n1172), .Z(n141) );
  NANDN U1393 ( .A(B[36]), .B(n1173), .Z(n1172) );
  NANDN U1394 ( .A(A[36]), .B(n143), .Z(n1173) );
  NANDN U1395 ( .A(n143), .B(A[36]), .Z(n1171) );
  AND U1396 ( .A(n1174), .B(n1175), .Z(n143) );
  NANDN U1397 ( .A(B[35]), .B(n1176), .Z(n1175) );
  NANDN U1398 ( .A(A[35]), .B(n145), .Z(n1176) );
  NANDN U1399 ( .A(n145), .B(A[35]), .Z(n1174) );
  AND U1400 ( .A(n1177), .B(n1178), .Z(n145) );
  NANDN U1401 ( .A(B[34]), .B(n1179), .Z(n1178) );
  NANDN U1402 ( .A(A[34]), .B(n147), .Z(n1179) );
  NANDN U1403 ( .A(n147), .B(A[34]), .Z(n1177) );
  AND U1404 ( .A(n1180), .B(n1181), .Z(n147) );
  NANDN U1405 ( .A(B[33]), .B(n1182), .Z(n1181) );
  NANDN U1406 ( .A(A[33]), .B(n149), .Z(n1182) );
  NANDN U1407 ( .A(n149), .B(A[33]), .Z(n1180) );
  AND U1408 ( .A(n1183), .B(n1184), .Z(n149) );
  NANDN U1409 ( .A(B[32]), .B(n1185), .Z(n1184) );
  NANDN U1410 ( .A(A[32]), .B(n151), .Z(n1185) );
  NANDN U1411 ( .A(n151), .B(A[32]), .Z(n1183) );
  AND U1412 ( .A(n1186), .B(n1187), .Z(n151) );
  NANDN U1413 ( .A(B[31]), .B(n1188), .Z(n1187) );
  NANDN U1414 ( .A(A[31]), .B(n153), .Z(n1188) );
  NANDN U1415 ( .A(n153), .B(A[31]), .Z(n1186) );
  AND U1416 ( .A(n1189), .B(n1190), .Z(n153) );
  NANDN U1417 ( .A(B[30]), .B(n1191), .Z(n1190) );
  NANDN U1418 ( .A(A[30]), .B(n155), .Z(n1191) );
  NANDN U1419 ( .A(n155), .B(A[30]), .Z(n1189) );
  AND U1420 ( .A(n1192), .B(n1193), .Z(n155) );
  NANDN U1421 ( .A(B[29]), .B(n1194), .Z(n1193) );
  NANDN U1422 ( .A(A[29]), .B(n159), .Z(n1194) );
  NANDN U1423 ( .A(n159), .B(A[29]), .Z(n1192) );
  AND U1424 ( .A(n1195), .B(n1196), .Z(n159) );
  NANDN U1425 ( .A(B[28]), .B(n1197), .Z(n1196) );
  NANDN U1426 ( .A(A[28]), .B(n161), .Z(n1197) );
  NANDN U1427 ( .A(n161), .B(A[28]), .Z(n1195) );
  AND U1428 ( .A(n1198), .B(n1199), .Z(n161) );
  NANDN U1429 ( .A(B[27]), .B(n1200), .Z(n1199) );
  NANDN U1430 ( .A(A[27]), .B(n163), .Z(n1200) );
  NANDN U1431 ( .A(n163), .B(A[27]), .Z(n1198) );
  AND U1432 ( .A(n1201), .B(n1202), .Z(n163) );
  NANDN U1433 ( .A(B[26]), .B(n1203), .Z(n1202) );
  NANDN U1434 ( .A(A[26]), .B(n165), .Z(n1203) );
  NANDN U1435 ( .A(n165), .B(A[26]), .Z(n1201) );
  AND U1436 ( .A(n1204), .B(n1205), .Z(n165) );
  NANDN U1437 ( .A(B[25]), .B(n1206), .Z(n1205) );
  NANDN U1438 ( .A(A[25]), .B(n167), .Z(n1206) );
  NANDN U1439 ( .A(n167), .B(A[25]), .Z(n1204) );
  AND U1440 ( .A(n1207), .B(n1208), .Z(n167) );
  NANDN U1441 ( .A(B[24]), .B(n1209), .Z(n1208) );
  NANDN U1442 ( .A(A[24]), .B(n205), .Z(n1209) );
  NANDN U1443 ( .A(n205), .B(A[24]), .Z(n1207) );
  AND U1444 ( .A(n1210), .B(n1211), .Z(n205) );
  NANDN U1445 ( .A(B[23]), .B(n1212), .Z(n1211) );
  NANDN U1446 ( .A(A[23]), .B(n257), .Z(n1212) );
  NANDN U1447 ( .A(n257), .B(A[23]), .Z(n1210) );
  AND U1448 ( .A(n1213), .B(n1214), .Z(n257) );
  NANDN U1449 ( .A(B[22]), .B(n1215), .Z(n1214) );
  NANDN U1450 ( .A(A[22]), .B(n309), .Z(n1215) );
  NANDN U1451 ( .A(n309), .B(A[22]), .Z(n1213) );
  AND U1452 ( .A(n1216), .B(n1217), .Z(n309) );
  NANDN U1453 ( .A(B[21]), .B(n1218), .Z(n1217) );
  NANDN U1454 ( .A(A[21]), .B(n361), .Z(n1218) );
  NANDN U1455 ( .A(n361), .B(A[21]), .Z(n1216) );
  AND U1456 ( .A(n1219), .B(n1220), .Z(n361) );
  NANDN U1457 ( .A(B[20]), .B(n1221), .Z(n1220) );
  NANDN U1458 ( .A(A[20]), .B(n413), .Z(n1221) );
  NANDN U1459 ( .A(n413), .B(A[20]), .Z(n1219) );
  AND U1460 ( .A(n1222), .B(n1223), .Z(n413) );
  NANDN U1461 ( .A(B[19]), .B(n1224), .Z(n1223) );
  NANDN U1462 ( .A(A[19]), .B(n466), .Z(n1224) );
  NANDN U1463 ( .A(n466), .B(A[19]), .Z(n1222) );
  AND U1464 ( .A(n1225), .B(n1226), .Z(n466) );
  NANDN U1465 ( .A(B[18]), .B(n1227), .Z(n1226) );
  NANDN U1466 ( .A(A[18]), .B(n518), .Z(n1227) );
  NANDN U1467 ( .A(n518), .B(A[18]), .Z(n1225) );
  AND U1468 ( .A(n1228), .B(n1229), .Z(n518) );
  NANDN U1469 ( .A(B[17]), .B(n1230), .Z(n1229) );
  NANDN U1470 ( .A(A[17]), .B(n570), .Z(n1230) );
  NANDN U1471 ( .A(n570), .B(A[17]), .Z(n1228) );
  AND U1472 ( .A(n1231), .B(n1232), .Z(n570) );
  NANDN U1473 ( .A(B[16]), .B(n1233), .Z(n1232) );
  NANDN U1474 ( .A(A[16]), .B(n622), .Z(n1233) );
  NANDN U1475 ( .A(n622), .B(A[16]), .Z(n1231) );
  AND U1476 ( .A(n1234), .B(n1235), .Z(n622) );
  NANDN U1477 ( .A(B[15]), .B(n1236), .Z(n1235) );
  NANDN U1478 ( .A(A[15]), .B(n674), .Z(n1236) );
  NANDN U1479 ( .A(n674), .B(A[15]), .Z(n1234) );
  AND U1480 ( .A(n1237), .B(n1238), .Z(n674) );
  NANDN U1481 ( .A(B[14]), .B(n1239), .Z(n1238) );
  NANDN U1482 ( .A(A[14]), .B(n726), .Z(n1239) );
  NANDN U1483 ( .A(n726), .B(A[14]), .Z(n1237) );
  AND U1484 ( .A(n1240), .B(n1241), .Z(n726) );
  NANDN U1485 ( .A(B[13]), .B(n1242), .Z(n1241) );
  NANDN U1486 ( .A(A[13]), .B(n778), .Z(n1242) );
  NANDN U1487 ( .A(n778), .B(A[13]), .Z(n1240) );
  AND U1488 ( .A(n1243), .B(n1244), .Z(n778) );
  NANDN U1489 ( .A(B[12]), .B(n1245), .Z(n1244) );
  NANDN U1490 ( .A(A[12]), .B(n830), .Z(n1245) );
  NANDN U1491 ( .A(n830), .B(A[12]), .Z(n1243) );
  AND U1492 ( .A(n1246), .B(n1247), .Z(n830) );
  NANDN U1493 ( .A(B[11]), .B(n1248), .Z(n1247) );
  NANDN U1494 ( .A(A[11]), .B(n882), .Z(n1248) );
  NANDN U1495 ( .A(n882), .B(A[11]), .Z(n1246) );
  AND U1496 ( .A(n1249), .B(n1250), .Z(n882) );
  NANDN U1497 ( .A(B[10]), .B(n1251), .Z(n1250) );
  NANDN U1498 ( .A(A[10]), .B(n934), .Z(n1251) );
  NANDN U1499 ( .A(n934), .B(A[10]), .Z(n1249) );
  AND U1500 ( .A(n1252), .B(n1253), .Z(n934) );
  NANDN U1501 ( .A(B[9]), .B(n1254), .Z(n1253) );
  OR U1502 ( .A(n3), .B(A[9]), .Z(n1254) );
  NAND U1503 ( .A(A[9]), .B(n3), .Z(n1252) );
  NAND U1504 ( .A(n1255), .B(n1256), .Z(n3) );
  NANDN U1505 ( .A(B[8]), .B(n1257), .Z(n1256) );
  NANDN U1506 ( .A(A[8]), .B(n25), .Z(n1257) );
  NANDN U1507 ( .A(n25), .B(A[8]), .Z(n1255) );
  AND U1508 ( .A(n1258), .B(n1259), .Z(n25) );
  NANDN U1509 ( .A(B[7]), .B(n1260), .Z(n1259) );
  NANDN U1510 ( .A(A[7]), .B(n47), .Z(n1260) );
  NANDN U1511 ( .A(n47), .B(A[7]), .Z(n1258) );
  AND U1512 ( .A(n1261), .B(n1262), .Z(n47) );
  NANDN U1513 ( .A(B[6]), .B(n1263), .Z(n1262) );
  NANDN U1514 ( .A(A[6]), .B(n69), .Z(n1263) );
  NANDN U1515 ( .A(n69), .B(A[6]), .Z(n1261) );
  AND U1516 ( .A(n1264), .B(n1265), .Z(n69) );
  NANDN U1517 ( .A(B[5]), .B(n1266), .Z(n1265) );
  NANDN U1518 ( .A(A[5]), .B(n91), .Z(n1266) );
  NANDN U1519 ( .A(n91), .B(A[5]), .Z(n1264) );
  AND U1520 ( .A(n1267), .B(n1268), .Z(n91) );
  NANDN U1521 ( .A(B[4]), .B(n1269), .Z(n1268) );
  NANDN U1522 ( .A(A[4]), .B(n113), .Z(n1269) );
  NANDN U1523 ( .A(n113), .B(A[4]), .Z(n1267) );
  AND U1524 ( .A(n1270), .B(n1271), .Z(n113) );
  NANDN U1525 ( .A(B[3]), .B(n1272), .Z(n1271) );
  NANDN U1526 ( .A(A[3]), .B(n135), .Z(n1272) );
  NANDN U1527 ( .A(n135), .B(A[3]), .Z(n1270) );
  AND U1528 ( .A(n1273), .B(n1274), .Z(n135) );
  NANDN U1529 ( .A(B[2]), .B(n1275), .Z(n1274) );
  NANDN U1530 ( .A(A[2]), .B(n157), .Z(n1275) );
  NANDN U1531 ( .A(n157), .B(A[2]), .Z(n1273) );
  AND U1532 ( .A(n1276), .B(n1277), .Z(n157) );
  NANDN U1533 ( .A(B[1]), .B(n1278), .Z(n1277) );
  NAND U1534 ( .A(n2), .B(n1), .Z(n1278) );
  NAND U1535 ( .A(A[1]), .B(n1279), .Z(n1276) );
  NAND U1536 ( .A(n1279), .B(n1280), .Z(DIFF[0]) );
  NANDN U1537 ( .A(B[0]), .B(A[0]), .Z(n1280) );
  NANDN U1538 ( .A(A[0]), .B(B[0]), .Z(n1279) );
endmodule


module modmult_step_N256_2_DW01_cmp2_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [257:0] A;
  input [257:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;

  NAND U1 ( .A(n1), .B(n2), .Z(LT_LE) );
  NOR U2 ( .A(B[257]), .B(B[256]), .Z(n2) );
  AND U3 ( .A(n3), .B(n4), .Z(n1) );
  NAND U4 ( .A(n5), .B(n6), .Z(n4) );
  NANDN U5 ( .A(B[255]), .B(A[255]), .Z(n6) );
  NAND U6 ( .A(n7), .B(n8), .Z(n5) );
  NANDN U7 ( .A(A[254]), .B(B[254]), .Z(n8) );
  NAND U8 ( .A(n9), .B(n10), .Z(n7) );
  NANDN U9 ( .A(B[254]), .B(A[254]), .Z(n10) );
  AND U10 ( .A(n11), .B(n12), .Z(n9) );
  NAND U11 ( .A(n13), .B(n14), .Z(n12) );
  NANDN U12 ( .A(A[253]), .B(B[253]), .Z(n14) );
  AND U13 ( .A(n15), .B(n16), .Z(n13) );
  NANDN U14 ( .A(A[252]), .B(B[252]), .Z(n16) );
  NAND U15 ( .A(n17), .B(n18), .Z(n15) );
  NANDN U16 ( .A(B[252]), .B(A[252]), .Z(n18) );
  AND U17 ( .A(n19), .B(n20), .Z(n17) );
  NAND U18 ( .A(n21), .B(n22), .Z(n20) );
  NANDN U19 ( .A(A[251]), .B(B[251]), .Z(n22) );
  AND U20 ( .A(n23), .B(n24), .Z(n21) );
  NANDN U21 ( .A(A[250]), .B(B[250]), .Z(n24) );
  NAND U22 ( .A(n25), .B(n26), .Z(n23) );
  NANDN U23 ( .A(B[250]), .B(A[250]), .Z(n26) );
  AND U24 ( .A(n27), .B(n28), .Z(n25) );
  NAND U25 ( .A(n29), .B(n30), .Z(n28) );
  NANDN U26 ( .A(A[249]), .B(B[249]), .Z(n30) );
  AND U27 ( .A(n31), .B(n32), .Z(n29) );
  NANDN U28 ( .A(A[248]), .B(B[248]), .Z(n32) );
  NAND U29 ( .A(n33), .B(n34), .Z(n31) );
  NANDN U30 ( .A(B[248]), .B(A[248]), .Z(n34) );
  AND U31 ( .A(n35), .B(n36), .Z(n33) );
  NAND U32 ( .A(n37), .B(n38), .Z(n36) );
  NANDN U33 ( .A(A[247]), .B(B[247]), .Z(n38) );
  AND U34 ( .A(n39), .B(n40), .Z(n37) );
  NANDN U35 ( .A(A[246]), .B(B[246]), .Z(n40) );
  NAND U36 ( .A(n41), .B(n42), .Z(n39) );
  NANDN U37 ( .A(B[246]), .B(A[246]), .Z(n42) );
  AND U38 ( .A(n43), .B(n44), .Z(n41) );
  NAND U39 ( .A(n45), .B(n46), .Z(n44) );
  NANDN U40 ( .A(A[245]), .B(B[245]), .Z(n46) );
  AND U41 ( .A(n47), .B(n48), .Z(n45) );
  NANDN U42 ( .A(A[244]), .B(B[244]), .Z(n48) );
  NAND U43 ( .A(n49), .B(n50), .Z(n47) );
  NANDN U44 ( .A(B[244]), .B(A[244]), .Z(n50) );
  AND U45 ( .A(n51), .B(n52), .Z(n49) );
  NAND U46 ( .A(n53), .B(n54), .Z(n52) );
  NANDN U47 ( .A(A[243]), .B(B[243]), .Z(n54) );
  AND U48 ( .A(n55), .B(n56), .Z(n53) );
  NANDN U49 ( .A(A[242]), .B(B[242]), .Z(n56) );
  NAND U50 ( .A(n57), .B(n58), .Z(n55) );
  NANDN U51 ( .A(B[242]), .B(A[242]), .Z(n58) );
  AND U52 ( .A(n59), .B(n60), .Z(n57) );
  NAND U53 ( .A(n61), .B(n62), .Z(n60) );
  NANDN U54 ( .A(A[241]), .B(B[241]), .Z(n62) );
  AND U55 ( .A(n63), .B(n64), .Z(n61) );
  NANDN U56 ( .A(A[240]), .B(B[240]), .Z(n64) );
  NAND U57 ( .A(n65), .B(n66), .Z(n63) );
  NANDN U58 ( .A(B[240]), .B(A[240]), .Z(n66) );
  AND U59 ( .A(n67), .B(n68), .Z(n65) );
  NAND U60 ( .A(n69), .B(n70), .Z(n68) );
  NANDN U61 ( .A(A[239]), .B(B[239]), .Z(n70) );
  AND U62 ( .A(n71), .B(n72), .Z(n69) );
  NANDN U63 ( .A(A[238]), .B(B[238]), .Z(n72) );
  NAND U64 ( .A(n73), .B(n74), .Z(n71) );
  NANDN U65 ( .A(B[238]), .B(A[238]), .Z(n74) );
  AND U66 ( .A(n75), .B(n76), .Z(n73) );
  NAND U67 ( .A(n77), .B(n78), .Z(n76) );
  NANDN U68 ( .A(A[237]), .B(B[237]), .Z(n78) );
  AND U69 ( .A(n79), .B(n80), .Z(n77) );
  NANDN U70 ( .A(A[236]), .B(B[236]), .Z(n80) );
  NAND U71 ( .A(n81), .B(n82), .Z(n79) );
  NANDN U72 ( .A(B[236]), .B(A[236]), .Z(n82) );
  AND U73 ( .A(n83), .B(n84), .Z(n81) );
  NAND U74 ( .A(n85), .B(n86), .Z(n84) );
  NANDN U75 ( .A(A[235]), .B(B[235]), .Z(n86) );
  AND U76 ( .A(n87), .B(n88), .Z(n85) );
  NANDN U77 ( .A(A[234]), .B(B[234]), .Z(n88) );
  NAND U78 ( .A(n89), .B(n90), .Z(n87) );
  NANDN U79 ( .A(B[234]), .B(A[234]), .Z(n90) );
  AND U80 ( .A(n91), .B(n92), .Z(n89) );
  NAND U81 ( .A(n93), .B(n94), .Z(n92) );
  NANDN U82 ( .A(A[233]), .B(B[233]), .Z(n94) );
  AND U83 ( .A(n95), .B(n96), .Z(n93) );
  NANDN U84 ( .A(A[232]), .B(B[232]), .Z(n96) );
  NAND U85 ( .A(n97), .B(n98), .Z(n95) );
  NANDN U86 ( .A(B[232]), .B(A[232]), .Z(n98) );
  AND U87 ( .A(n99), .B(n100), .Z(n97) );
  NAND U88 ( .A(n101), .B(n102), .Z(n100) );
  NANDN U89 ( .A(A[231]), .B(B[231]), .Z(n102) );
  AND U90 ( .A(n103), .B(n104), .Z(n101) );
  NANDN U91 ( .A(A[230]), .B(B[230]), .Z(n104) );
  NAND U92 ( .A(n105), .B(n106), .Z(n103) );
  NANDN U93 ( .A(B[230]), .B(A[230]), .Z(n106) );
  AND U94 ( .A(n107), .B(n108), .Z(n105) );
  NAND U95 ( .A(n109), .B(n110), .Z(n108) );
  NANDN U96 ( .A(A[229]), .B(B[229]), .Z(n110) );
  AND U97 ( .A(n111), .B(n112), .Z(n109) );
  NANDN U98 ( .A(A[228]), .B(B[228]), .Z(n112) );
  NAND U99 ( .A(n113), .B(n114), .Z(n111) );
  NANDN U100 ( .A(B[228]), .B(A[228]), .Z(n114) );
  AND U101 ( .A(n115), .B(n116), .Z(n113) );
  NAND U102 ( .A(n117), .B(n118), .Z(n116) );
  NANDN U103 ( .A(A[227]), .B(B[227]), .Z(n118) );
  AND U104 ( .A(n119), .B(n120), .Z(n117) );
  NANDN U105 ( .A(A[226]), .B(B[226]), .Z(n120) );
  NAND U106 ( .A(n121), .B(n122), .Z(n119) );
  NANDN U107 ( .A(B[226]), .B(A[226]), .Z(n122) );
  AND U108 ( .A(n123), .B(n124), .Z(n121) );
  NAND U109 ( .A(n125), .B(n126), .Z(n124) );
  NANDN U110 ( .A(A[225]), .B(B[225]), .Z(n126) );
  AND U111 ( .A(n127), .B(n128), .Z(n125) );
  NANDN U112 ( .A(A[224]), .B(B[224]), .Z(n128) );
  NAND U113 ( .A(n129), .B(n130), .Z(n127) );
  NANDN U114 ( .A(B[224]), .B(A[224]), .Z(n130) );
  AND U115 ( .A(n131), .B(n132), .Z(n129) );
  NAND U116 ( .A(n133), .B(n134), .Z(n132) );
  NANDN U117 ( .A(A[223]), .B(B[223]), .Z(n134) );
  AND U118 ( .A(n135), .B(n136), .Z(n133) );
  NANDN U119 ( .A(A[222]), .B(B[222]), .Z(n136) );
  NAND U120 ( .A(n137), .B(n138), .Z(n135) );
  NANDN U121 ( .A(B[222]), .B(A[222]), .Z(n138) );
  AND U122 ( .A(n139), .B(n140), .Z(n137) );
  NAND U123 ( .A(n141), .B(n142), .Z(n140) );
  NANDN U124 ( .A(A[221]), .B(B[221]), .Z(n142) );
  AND U125 ( .A(n143), .B(n144), .Z(n141) );
  NANDN U126 ( .A(A[220]), .B(B[220]), .Z(n144) );
  NAND U127 ( .A(n145), .B(n146), .Z(n143) );
  NANDN U128 ( .A(B[220]), .B(A[220]), .Z(n146) );
  AND U129 ( .A(n147), .B(n148), .Z(n145) );
  NAND U130 ( .A(n149), .B(n150), .Z(n148) );
  NANDN U131 ( .A(A[219]), .B(B[219]), .Z(n150) );
  AND U132 ( .A(n151), .B(n152), .Z(n149) );
  NANDN U133 ( .A(A[218]), .B(B[218]), .Z(n152) );
  NAND U134 ( .A(n153), .B(n154), .Z(n151) );
  NANDN U135 ( .A(B[218]), .B(A[218]), .Z(n154) );
  AND U136 ( .A(n155), .B(n156), .Z(n153) );
  NAND U137 ( .A(n157), .B(n158), .Z(n156) );
  NANDN U138 ( .A(A[217]), .B(B[217]), .Z(n158) );
  AND U139 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U140 ( .A(A[216]), .B(B[216]), .Z(n160) );
  NAND U141 ( .A(n161), .B(n162), .Z(n159) );
  NANDN U142 ( .A(B[216]), .B(A[216]), .Z(n162) );
  AND U143 ( .A(n163), .B(n164), .Z(n161) );
  NAND U144 ( .A(n165), .B(n166), .Z(n164) );
  NANDN U145 ( .A(A[215]), .B(B[215]), .Z(n166) );
  AND U146 ( .A(n167), .B(n168), .Z(n165) );
  NANDN U147 ( .A(A[214]), .B(B[214]), .Z(n168) );
  NAND U148 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U149 ( .A(B[214]), .B(A[214]), .Z(n170) );
  AND U150 ( .A(n171), .B(n172), .Z(n169) );
  NAND U151 ( .A(n173), .B(n174), .Z(n172) );
  NANDN U152 ( .A(A[213]), .B(B[213]), .Z(n174) );
  AND U153 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U154 ( .A(A[212]), .B(B[212]), .Z(n176) );
  NAND U155 ( .A(n177), .B(n178), .Z(n175) );
  NANDN U156 ( .A(B[212]), .B(A[212]), .Z(n178) );
  AND U157 ( .A(n179), .B(n180), .Z(n177) );
  NAND U158 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U159 ( .A(A[211]), .B(B[211]), .Z(n182) );
  AND U160 ( .A(n183), .B(n184), .Z(n181) );
  NANDN U161 ( .A(A[210]), .B(B[210]), .Z(n184) );
  NAND U162 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U163 ( .A(B[210]), .B(A[210]), .Z(n186) );
  AND U164 ( .A(n187), .B(n188), .Z(n185) );
  NAND U165 ( .A(n189), .B(n190), .Z(n188) );
  NANDN U166 ( .A(A[209]), .B(B[209]), .Z(n190) );
  AND U167 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U168 ( .A(A[208]), .B(B[208]), .Z(n192) );
  NAND U169 ( .A(n193), .B(n194), .Z(n191) );
  NANDN U170 ( .A(B[208]), .B(A[208]), .Z(n194) );
  AND U171 ( .A(n195), .B(n196), .Z(n193) );
  NAND U172 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U173 ( .A(A[207]), .B(B[207]), .Z(n198) );
  AND U174 ( .A(n199), .B(n200), .Z(n197) );
  NANDN U175 ( .A(A[206]), .B(B[206]), .Z(n200) );
  NAND U176 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U177 ( .A(B[206]), .B(A[206]), .Z(n202) );
  AND U178 ( .A(n203), .B(n204), .Z(n201) );
  NAND U179 ( .A(n205), .B(n206), .Z(n204) );
  NANDN U180 ( .A(A[205]), .B(B[205]), .Z(n206) );
  AND U181 ( .A(n207), .B(n208), .Z(n205) );
  NANDN U182 ( .A(A[204]), .B(B[204]), .Z(n208) );
  NAND U183 ( .A(n209), .B(n210), .Z(n207) );
  NANDN U184 ( .A(B[204]), .B(A[204]), .Z(n210) );
  AND U185 ( .A(n211), .B(n212), .Z(n209) );
  NAND U186 ( .A(n213), .B(n214), .Z(n212) );
  NANDN U187 ( .A(A[203]), .B(B[203]), .Z(n214) );
  AND U188 ( .A(n215), .B(n216), .Z(n213) );
  NANDN U189 ( .A(A[202]), .B(B[202]), .Z(n216) );
  NAND U190 ( .A(n217), .B(n218), .Z(n215) );
  NANDN U191 ( .A(B[202]), .B(A[202]), .Z(n218) );
  AND U192 ( .A(n219), .B(n220), .Z(n217) );
  NAND U193 ( .A(n221), .B(n222), .Z(n220) );
  NANDN U194 ( .A(A[201]), .B(B[201]), .Z(n222) );
  AND U195 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U196 ( .A(A[200]), .B(B[200]), .Z(n224) );
  NAND U197 ( .A(n225), .B(n226), .Z(n223) );
  NANDN U198 ( .A(B[200]), .B(A[200]), .Z(n226) );
  AND U199 ( .A(n227), .B(n228), .Z(n225) );
  NAND U200 ( .A(n229), .B(n230), .Z(n228) );
  NANDN U201 ( .A(A[199]), .B(B[199]), .Z(n230) );
  AND U202 ( .A(n231), .B(n232), .Z(n229) );
  NANDN U203 ( .A(A[198]), .B(B[198]), .Z(n232) );
  NAND U204 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U205 ( .A(B[198]), .B(A[198]), .Z(n234) );
  AND U206 ( .A(n235), .B(n236), .Z(n233) );
  NAND U207 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U208 ( .A(A[197]), .B(B[197]), .Z(n238) );
  AND U209 ( .A(n239), .B(n240), .Z(n237) );
  NANDN U210 ( .A(A[196]), .B(B[196]), .Z(n240) );
  NAND U211 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U212 ( .A(B[196]), .B(A[196]), .Z(n242) );
  AND U213 ( .A(n243), .B(n244), .Z(n241) );
  NAND U214 ( .A(n245), .B(n246), .Z(n244) );
  NANDN U215 ( .A(A[195]), .B(B[195]), .Z(n246) );
  AND U216 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U217 ( .A(A[194]), .B(B[194]), .Z(n248) );
  NAND U218 ( .A(n249), .B(n250), .Z(n247) );
  NANDN U219 ( .A(B[194]), .B(A[194]), .Z(n250) );
  AND U220 ( .A(n251), .B(n252), .Z(n249) );
  NAND U221 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U222 ( .A(A[193]), .B(B[193]), .Z(n254) );
  AND U223 ( .A(n255), .B(n256), .Z(n253) );
  NANDN U224 ( .A(A[192]), .B(B[192]), .Z(n256) );
  NAND U225 ( .A(n257), .B(n258), .Z(n255) );
  NANDN U226 ( .A(B[192]), .B(A[192]), .Z(n258) );
  AND U227 ( .A(n259), .B(n260), .Z(n257) );
  NAND U228 ( .A(n261), .B(n262), .Z(n260) );
  NANDN U229 ( .A(A[191]), .B(B[191]), .Z(n262) );
  AND U230 ( .A(n263), .B(n264), .Z(n261) );
  NANDN U231 ( .A(A[190]), .B(B[190]), .Z(n264) );
  NAND U232 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U233 ( .A(B[190]), .B(A[190]), .Z(n266) );
  AND U234 ( .A(n267), .B(n268), .Z(n265) );
  NAND U235 ( .A(n269), .B(n270), .Z(n268) );
  NANDN U236 ( .A(A[189]), .B(B[189]), .Z(n270) );
  AND U237 ( .A(n271), .B(n272), .Z(n269) );
  NANDN U238 ( .A(A[188]), .B(B[188]), .Z(n272) );
  NAND U239 ( .A(n273), .B(n274), .Z(n271) );
  NANDN U240 ( .A(B[188]), .B(A[188]), .Z(n274) );
  AND U241 ( .A(n275), .B(n276), .Z(n273) );
  NAND U242 ( .A(n277), .B(n278), .Z(n276) );
  NANDN U243 ( .A(A[187]), .B(B[187]), .Z(n278) );
  AND U244 ( .A(n279), .B(n280), .Z(n277) );
  NANDN U245 ( .A(A[186]), .B(B[186]), .Z(n280) );
  NAND U246 ( .A(n281), .B(n282), .Z(n279) );
  NANDN U247 ( .A(B[186]), .B(A[186]), .Z(n282) );
  AND U248 ( .A(n283), .B(n284), .Z(n281) );
  NAND U249 ( .A(n285), .B(n286), .Z(n284) );
  NANDN U250 ( .A(A[185]), .B(B[185]), .Z(n286) );
  AND U251 ( .A(n287), .B(n288), .Z(n285) );
  NANDN U252 ( .A(A[184]), .B(B[184]), .Z(n288) );
  NAND U253 ( .A(n289), .B(n290), .Z(n287) );
  NANDN U254 ( .A(B[184]), .B(A[184]), .Z(n290) );
  AND U255 ( .A(n291), .B(n292), .Z(n289) );
  NAND U256 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U257 ( .A(A[183]), .B(B[183]), .Z(n294) );
  AND U258 ( .A(n295), .B(n296), .Z(n293) );
  NANDN U259 ( .A(A[182]), .B(B[182]), .Z(n296) );
  NAND U260 ( .A(n297), .B(n298), .Z(n295) );
  NANDN U261 ( .A(B[182]), .B(A[182]), .Z(n298) );
  AND U262 ( .A(n299), .B(n300), .Z(n297) );
  NAND U263 ( .A(n301), .B(n302), .Z(n300) );
  NANDN U264 ( .A(A[181]), .B(B[181]), .Z(n302) );
  AND U265 ( .A(n303), .B(n304), .Z(n301) );
  NANDN U266 ( .A(A[180]), .B(B[180]), .Z(n304) );
  NAND U267 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U268 ( .A(B[180]), .B(A[180]), .Z(n306) );
  AND U269 ( .A(n307), .B(n308), .Z(n305) );
  NAND U270 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U271 ( .A(A[179]), .B(B[179]), .Z(n310) );
  AND U272 ( .A(n311), .B(n312), .Z(n309) );
  NANDN U273 ( .A(A[178]), .B(B[178]), .Z(n312) );
  NAND U274 ( .A(n313), .B(n314), .Z(n311) );
  NANDN U275 ( .A(B[178]), .B(A[178]), .Z(n314) );
  AND U276 ( .A(n315), .B(n316), .Z(n313) );
  NAND U277 ( .A(n317), .B(n318), .Z(n316) );
  NANDN U278 ( .A(A[177]), .B(B[177]), .Z(n318) );
  AND U279 ( .A(n319), .B(n320), .Z(n317) );
  NANDN U280 ( .A(A[176]), .B(B[176]), .Z(n320) );
  NAND U281 ( .A(n321), .B(n322), .Z(n319) );
  NANDN U282 ( .A(B[176]), .B(A[176]), .Z(n322) );
  AND U283 ( .A(n323), .B(n324), .Z(n321) );
  NAND U284 ( .A(n325), .B(n326), .Z(n324) );
  NANDN U285 ( .A(A[175]), .B(B[175]), .Z(n326) );
  AND U286 ( .A(n327), .B(n328), .Z(n325) );
  NANDN U287 ( .A(A[174]), .B(B[174]), .Z(n328) );
  NAND U288 ( .A(n329), .B(n330), .Z(n327) );
  NANDN U289 ( .A(B[174]), .B(A[174]), .Z(n330) );
  AND U290 ( .A(n331), .B(n332), .Z(n329) );
  NAND U291 ( .A(n333), .B(n334), .Z(n332) );
  NANDN U292 ( .A(A[173]), .B(B[173]), .Z(n334) );
  AND U293 ( .A(n335), .B(n336), .Z(n333) );
  NANDN U294 ( .A(A[172]), .B(B[172]), .Z(n336) );
  NAND U295 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U296 ( .A(B[172]), .B(A[172]), .Z(n338) );
  AND U297 ( .A(n339), .B(n340), .Z(n337) );
  NAND U298 ( .A(n341), .B(n342), .Z(n340) );
  NANDN U299 ( .A(A[171]), .B(B[171]), .Z(n342) );
  AND U300 ( .A(n343), .B(n344), .Z(n341) );
  NANDN U301 ( .A(A[170]), .B(B[170]), .Z(n344) );
  NAND U302 ( .A(n345), .B(n346), .Z(n343) );
  NANDN U303 ( .A(B[170]), .B(A[170]), .Z(n346) );
  AND U304 ( .A(n347), .B(n348), .Z(n345) );
  NAND U305 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U306 ( .A(A[169]), .B(B[169]), .Z(n350) );
  AND U307 ( .A(n351), .B(n352), .Z(n349) );
  NANDN U308 ( .A(A[168]), .B(B[168]), .Z(n352) );
  NAND U309 ( .A(n353), .B(n354), .Z(n351) );
  NANDN U310 ( .A(B[168]), .B(A[168]), .Z(n354) );
  AND U311 ( .A(n355), .B(n356), .Z(n353) );
  NAND U312 ( .A(n357), .B(n358), .Z(n356) );
  NANDN U313 ( .A(A[167]), .B(B[167]), .Z(n358) );
  AND U314 ( .A(n359), .B(n360), .Z(n357) );
  NANDN U315 ( .A(A[166]), .B(B[166]), .Z(n360) );
  NAND U316 ( .A(n361), .B(n362), .Z(n359) );
  NANDN U317 ( .A(B[166]), .B(A[166]), .Z(n362) );
  AND U318 ( .A(n363), .B(n364), .Z(n361) );
  NAND U319 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U320 ( .A(A[165]), .B(B[165]), .Z(n366) );
  AND U321 ( .A(n367), .B(n368), .Z(n365) );
  NANDN U322 ( .A(A[164]), .B(B[164]), .Z(n368) );
  NAND U323 ( .A(n369), .B(n370), .Z(n367) );
  NANDN U324 ( .A(B[164]), .B(A[164]), .Z(n370) );
  AND U325 ( .A(n371), .B(n372), .Z(n369) );
  NAND U326 ( .A(n373), .B(n374), .Z(n372) );
  NANDN U327 ( .A(A[163]), .B(B[163]), .Z(n374) );
  AND U328 ( .A(n375), .B(n376), .Z(n373) );
  NANDN U329 ( .A(A[162]), .B(B[162]), .Z(n376) );
  NAND U330 ( .A(n377), .B(n378), .Z(n375) );
  NANDN U331 ( .A(B[162]), .B(A[162]), .Z(n378) );
  AND U332 ( .A(n379), .B(n380), .Z(n377) );
  NAND U333 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U334 ( .A(A[161]), .B(B[161]), .Z(n382) );
  AND U335 ( .A(n383), .B(n384), .Z(n381) );
  NANDN U336 ( .A(A[160]), .B(B[160]), .Z(n384) );
  NAND U337 ( .A(n385), .B(n386), .Z(n383) );
  NANDN U338 ( .A(B[160]), .B(A[160]), .Z(n386) );
  AND U339 ( .A(n387), .B(n388), .Z(n385) );
  NAND U340 ( .A(n389), .B(n390), .Z(n388) );
  NANDN U341 ( .A(A[159]), .B(B[159]), .Z(n390) );
  AND U342 ( .A(n391), .B(n392), .Z(n389) );
  NANDN U343 ( .A(A[158]), .B(B[158]), .Z(n392) );
  NAND U344 ( .A(n393), .B(n394), .Z(n391) );
  NANDN U345 ( .A(B[158]), .B(A[158]), .Z(n394) );
  AND U346 ( .A(n395), .B(n396), .Z(n393) );
  NAND U347 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U348 ( .A(A[157]), .B(B[157]), .Z(n398) );
  AND U349 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U350 ( .A(A[156]), .B(B[156]), .Z(n400) );
  NAND U351 ( .A(n401), .B(n402), .Z(n399) );
  NANDN U352 ( .A(B[156]), .B(A[156]), .Z(n402) );
  AND U353 ( .A(n403), .B(n404), .Z(n401) );
  NAND U354 ( .A(n405), .B(n406), .Z(n404) );
  NANDN U355 ( .A(A[155]), .B(B[155]), .Z(n406) );
  AND U356 ( .A(n407), .B(n408), .Z(n405) );
  NANDN U357 ( .A(A[154]), .B(B[154]), .Z(n408) );
  NAND U358 ( .A(n409), .B(n410), .Z(n407) );
  NANDN U359 ( .A(B[154]), .B(A[154]), .Z(n410) );
  AND U360 ( .A(n411), .B(n412), .Z(n409) );
  NAND U361 ( .A(n413), .B(n414), .Z(n412) );
  NANDN U362 ( .A(A[153]), .B(B[153]), .Z(n414) );
  AND U363 ( .A(n415), .B(n416), .Z(n413) );
  NANDN U364 ( .A(A[152]), .B(B[152]), .Z(n416) );
  NAND U365 ( .A(n417), .B(n418), .Z(n415) );
  NANDN U366 ( .A(B[152]), .B(A[152]), .Z(n418) );
  AND U367 ( .A(n419), .B(n420), .Z(n417) );
  NAND U368 ( .A(n421), .B(n422), .Z(n420) );
  NANDN U369 ( .A(A[151]), .B(B[151]), .Z(n422) );
  AND U370 ( .A(n423), .B(n424), .Z(n421) );
  NANDN U371 ( .A(A[150]), .B(B[150]), .Z(n424) );
  NAND U372 ( .A(n425), .B(n426), .Z(n423) );
  NANDN U373 ( .A(B[150]), .B(A[150]), .Z(n426) );
  AND U374 ( .A(n427), .B(n428), .Z(n425) );
  NAND U375 ( .A(n429), .B(n430), .Z(n428) );
  NANDN U376 ( .A(A[149]), .B(B[149]), .Z(n430) );
  AND U377 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U378 ( .A(A[148]), .B(B[148]), .Z(n432) );
  NAND U379 ( .A(n433), .B(n434), .Z(n431) );
  NANDN U380 ( .A(B[148]), .B(A[148]), .Z(n434) );
  AND U381 ( .A(n435), .B(n436), .Z(n433) );
  NAND U382 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U383 ( .A(A[147]), .B(B[147]), .Z(n438) );
  AND U384 ( .A(n439), .B(n440), .Z(n437) );
  NANDN U385 ( .A(A[146]), .B(B[146]), .Z(n440) );
  NAND U386 ( .A(n441), .B(n442), .Z(n439) );
  NANDN U387 ( .A(B[146]), .B(A[146]), .Z(n442) );
  AND U388 ( .A(n443), .B(n444), .Z(n441) );
  NAND U389 ( .A(n445), .B(n446), .Z(n444) );
  NANDN U390 ( .A(A[145]), .B(B[145]), .Z(n446) );
  AND U391 ( .A(n447), .B(n448), .Z(n445) );
  NANDN U392 ( .A(A[144]), .B(B[144]), .Z(n448) );
  NAND U393 ( .A(n449), .B(n450), .Z(n447) );
  NANDN U394 ( .A(B[144]), .B(A[144]), .Z(n450) );
  AND U395 ( .A(n451), .B(n452), .Z(n449) );
  NAND U396 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U397 ( .A(A[143]), .B(B[143]), .Z(n454) );
  AND U398 ( .A(n455), .B(n456), .Z(n453) );
  NANDN U399 ( .A(A[142]), .B(B[142]), .Z(n456) );
  NAND U400 ( .A(n457), .B(n458), .Z(n455) );
  NANDN U401 ( .A(B[142]), .B(A[142]), .Z(n458) );
  AND U402 ( .A(n459), .B(n460), .Z(n457) );
  NAND U403 ( .A(n461), .B(n462), .Z(n460) );
  NANDN U404 ( .A(A[141]), .B(B[141]), .Z(n462) );
  AND U405 ( .A(n463), .B(n464), .Z(n461) );
  NANDN U406 ( .A(A[140]), .B(B[140]), .Z(n464) );
  NAND U407 ( .A(n465), .B(n466), .Z(n463) );
  NANDN U408 ( .A(B[140]), .B(A[140]), .Z(n466) );
  AND U409 ( .A(n467), .B(n468), .Z(n465) );
  NAND U410 ( .A(n469), .B(n470), .Z(n468) );
  NANDN U411 ( .A(A[139]), .B(B[139]), .Z(n470) );
  AND U412 ( .A(n471), .B(n472), .Z(n469) );
  NANDN U413 ( .A(A[138]), .B(B[138]), .Z(n472) );
  NAND U414 ( .A(n473), .B(n474), .Z(n471) );
  NANDN U415 ( .A(B[138]), .B(A[138]), .Z(n474) );
  AND U416 ( .A(n475), .B(n476), .Z(n473) );
  NAND U417 ( .A(n477), .B(n478), .Z(n476) );
  NANDN U418 ( .A(A[137]), .B(B[137]), .Z(n478) );
  AND U419 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U420 ( .A(A[136]), .B(B[136]), .Z(n480) );
  NAND U421 ( .A(n481), .B(n482), .Z(n479) );
  NANDN U422 ( .A(B[136]), .B(A[136]), .Z(n482) );
  AND U423 ( .A(n483), .B(n484), .Z(n481) );
  NAND U424 ( .A(n485), .B(n486), .Z(n484) );
  NANDN U425 ( .A(A[135]), .B(B[135]), .Z(n486) );
  AND U426 ( .A(n487), .B(n488), .Z(n485) );
  NANDN U427 ( .A(A[134]), .B(B[134]), .Z(n488) );
  NAND U428 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U429 ( .A(B[134]), .B(A[134]), .Z(n490) );
  AND U430 ( .A(n491), .B(n492), .Z(n489) );
  NAND U431 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U432 ( .A(A[133]), .B(B[133]), .Z(n494) );
  AND U433 ( .A(n495), .B(n496), .Z(n493) );
  NANDN U434 ( .A(A[132]), .B(B[132]), .Z(n496) );
  NAND U435 ( .A(n497), .B(n498), .Z(n495) );
  NANDN U436 ( .A(B[132]), .B(A[132]), .Z(n498) );
  AND U437 ( .A(n499), .B(n500), .Z(n497) );
  NAND U438 ( .A(n501), .B(n502), .Z(n500) );
  NANDN U439 ( .A(A[131]), .B(B[131]), .Z(n502) );
  AND U440 ( .A(n503), .B(n504), .Z(n501) );
  NANDN U441 ( .A(A[130]), .B(B[130]), .Z(n504) );
  NAND U442 ( .A(n505), .B(n506), .Z(n503) );
  NANDN U443 ( .A(B[130]), .B(A[130]), .Z(n506) );
  AND U444 ( .A(n507), .B(n508), .Z(n505) );
  NAND U445 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U446 ( .A(A[129]), .B(B[129]), .Z(n510) );
  AND U447 ( .A(n511), .B(n512), .Z(n509) );
  NANDN U448 ( .A(A[128]), .B(B[128]), .Z(n512) );
  NAND U449 ( .A(n513), .B(n514), .Z(n511) );
  NANDN U450 ( .A(B[128]), .B(A[128]), .Z(n514) );
  AND U451 ( .A(n515), .B(n516), .Z(n513) );
  NAND U452 ( .A(n517), .B(n518), .Z(n516) );
  NANDN U453 ( .A(A[127]), .B(B[127]), .Z(n518) );
  AND U454 ( .A(n519), .B(n520), .Z(n517) );
  NANDN U455 ( .A(A[126]), .B(B[126]), .Z(n520) );
  NAND U456 ( .A(n521), .B(n522), .Z(n519) );
  NANDN U457 ( .A(B[126]), .B(A[126]), .Z(n522) );
  AND U458 ( .A(n523), .B(n524), .Z(n521) );
  NAND U459 ( .A(n525), .B(n526), .Z(n524) );
  NANDN U460 ( .A(A[125]), .B(B[125]), .Z(n526) );
  AND U461 ( .A(n527), .B(n528), .Z(n525) );
  NANDN U462 ( .A(A[124]), .B(B[124]), .Z(n528) );
  NAND U463 ( .A(n529), .B(n530), .Z(n527) );
  NANDN U464 ( .A(B[124]), .B(A[124]), .Z(n530) );
  AND U465 ( .A(n531), .B(n532), .Z(n529) );
  NAND U466 ( .A(n533), .B(n534), .Z(n532) );
  NANDN U467 ( .A(A[123]), .B(B[123]), .Z(n534) );
  AND U468 ( .A(n535), .B(n536), .Z(n533) );
  NANDN U469 ( .A(A[122]), .B(B[122]), .Z(n536) );
  NAND U470 ( .A(n537), .B(n538), .Z(n535) );
  NANDN U471 ( .A(B[122]), .B(A[122]), .Z(n538) );
  AND U472 ( .A(n539), .B(n540), .Z(n537) );
  NAND U473 ( .A(n541), .B(n542), .Z(n540) );
  NANDN U474 ( .A(A[121]), .B(B[121]), .Z(n542) );
  AND U475 ( .A(n543), .B(n544), .Z(n541) );
  NANDN U476 ( .A(A[120]), .B(B[120]), .Z(n544) );
  NAND U477 ( .A(n545), .B(n546), .Z(n543) );
  NANDN U478 ( .A(B[120]), .B(A[120]), .Z(n546) );
  AND U479 ( .A(n547), .B(n548), .Z(n545) );
  NAND U480 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U481 ( .A(A[119]), .B(B[119]), .Z(n550) );
  AND U482 ( .A(n551), .B(n552), .Z(n549) );
  NANDN U483 ( .A(A[118]), .B(B[118]), .Z(n552) );
  NAND U484 ( .A(n553), .B(n554), .Z(n551) );
  NANDN U485 ( .A(B[118]), .B(A[118]), .Z(n554) );
  AND U486 ( .A(n555), .B(n556), .Z(n553) );
  NAND U487 ( .A(n557), .B(n558), .Z(n556) );
  NANDN U488 ( .A(A[117]), .B(B[117]), .Z(n558) );
  AND U489 ( .A(n559), .B(n560), .Z(n557) );
  NANDN U490 ( .A(A[116]), .B(B[116]), .Z(n560) );
  NAND U491 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U492 ( .A(B[116]), .B(A[116]), .Z(n562) );
  AND U493 ( .A(n563), .B(n564), .Z(n561) );
  NAND U494 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U495 ( .A(A[115]), .B(B[115]), .Z(n566) );
  AND U496 ( .A(n567), .B(n568), .Z(n565) );
  NANDN U497 ( .A(A[114]), .B(B[114]), .Z(n568) );
  NAND U498 ( .A(n569), .B(n570), .Z(n567) );
  NANDN U499 ( .A(B[114]), .B(A[114]), .Z(n570) );
  AND U500 ( .A(n571), .B(n572), .Z(n569) );
  NAND U501 ( .A(n573), .B(n574), .Z(n572) );
  NANDN U502 ( .A(A[113]), .B(B[113]), .Z(n574) );
  AND U503 ( .A(n575), .B(n576), .Z(n573) );
  NANDN U504 ( .A(A[112]), .B(B[112]), .Z(n576) );
  NAND U505 ( .A(n577), .B(n578), .Z(n575) );
  NANDN U506 ( .A(B[112]), .B(A[112]), .Z(n578) );
  AND U507 ( .A(n579), .B(n580), .Z(n577) );
  NAND U508 ( .A(n581), .B(n582), .Z(n580) );
  NANDN U509 ( .A(A[111]), .B(B[111]), .Z(n582) );
  AND U510 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U511 ( .A(A[110]), .B(B[110]), .Z(n584) );
  NAND U512 ( .A(n585), .B(n586), .Z(n583) );
  NANDN U513 ( .A(B[110]), .B(A[110]), .Z(n586) );
  AND U514 ( .A(n587), .B(n588), .Z(n585) );
  NAND U515 ( .A(n589), .B(n590), .Z(n588) );
  NANDN U516 ( .A(A[109]), .B(B[109]), .Z(n590) );
  AND U517 ( .A(n591), .B(n592), .Z(n589) );
  NANDN U518 ( .A(A[108]), .B(B[108]), .Z(n592) );
  NAND U519 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U520 ( .A(B[108]), .B(A[108]), .Z(n594) );
  AND U521 ( .A(n595), .B(n596), .Z(n593) );
  NAND U522 ( .A(n597), .B(n598), .Z(n596) );
  NANDN U523 ( .A(A[107]), .B(B[107]), .Z(n598) );
  AND U524 ( .A(n599), .B(n600), .Z(n597) );
  NANDN U525 ( .A(A[106]), .B(B[106]), .Z(n600) );
  NAND U526 ( .A(n601), .B(n602), .Z(n599) );
  NANDN U527 ( .A(B[106]), .B(A[106]), .Z(n602) );
  AND U528 ( .A(n603), .B(n604), .Z(n601) );
  NAND U529 ( .A(n605), .B(n606), .Z(n604) );
  NANDN U530 ( .A(A[105]), .B(B[105]), .Z(n606) );
  AND U531 ( .A(n607), .B(n608), .Z(n605) );
  NANDN U532 ( .A(A[104]), .B(B[104]), .Z(n608) );
  NAND U533 ( .A(n609), .B(n610), .Z(n607) );
  NANDN U534 ( .A(B[104]), .B(A[104]), .Z(n610) );
  AND U535 ( .A(n611), .B(n612), .Z(n609) );
  NAND U536 ( .A(n613), .B(n614), .Z(n612) );
  NANDN U537 ( .A(A[103]), .B(B[103]), .Z(n614) );
  AND U538 ( .A(n615), .B(n616), .Z(n613) );
  NANDN U539 ( .A(A[102]), .B(B[102]), .Z(n616) );
  NAND U540 ( .A(n617), .B(n618), .Z(n615) );
  NANDN U541 ( .A(B[102]), .B(A[102]), .Z(n618) );
  AND U542 ( .A(n619), .B(n620), .Z(n617) );
  NAND U543 ( .A(n621), .B(n622), .Z(n620) );
  NANDN U544 ( .A(A[101]), .B(B[101]), .Z(n622) );
  AND U545 ( .A(n623), .B(n624), .Z(n621) );
  NANDN U546 ( .A(A[100]), .B(B[100]), .Z(n624) );
  NAND U547 ( .A(n625), .B(n626), .Z(n623) );
  NANDN U548 ( .A(B[99]), .B(A[99]), .Z(n626) );
  AND U549 ( .A(n627), .B(n628), .Z(n625) );
  NAND U550 ( .A(n629), .B(n630), .Z(n628) );
  NANDN U551 ( .A(A[99]), .B(B[99]), .Z(n630) );
  AND U552 ( .A(n631), .B(n632), .Z(n629) );
  NANDN U553 ( .A(A[98]), .B(B[98]), .Z(n632) );
  NAND U554 ( .A(n633), .B(n634), .Z(n631) );
  NANDN U555 ( .A(B[98]), .B(A[98]), .Z(n634) );
  AND U556 ( .A(n635), .B(n636), .Z(n633) );
  NAND U557 ( .A(n637), .B(n638), .Z(n636) );
  NANDN U558 ( .A(A[97]), .B(B[97]), .Z(n638) );
  AND U559 ( .A(n639), .B(n640), .Z(n637) );
  NANDN U560 ( .A(A[96]), .B(B[96]), .Z(n640) );
  NAND U561 ( .A(n641), .B(n642), .Z(n639) );
  NANDN U562 ( .A(B[96]), .B(A[96]), .Z(n642) );
  AND U563 ( .A(n643), .B(n644), .Z(n641) );
  NAND U564 ( .A(n645), .B(n646), .Z(n644) );
  NANDN U565 ( .A(A[95]), .B(B[95]), .Z(n646) );
  AND U566 ( .A(n647), .B(n648), .Z(n645) );
  NANDN U567 ( .A(A[94]), .B(B[94]), .Z(n648) );
  NAND U568 ( .A(n649), .B(n650), .Z(n647) );
  NANDN U569 ( .A(B[94]), .B(A[94]), .Z(n650) );
  AND U570 ( .A(n651), .B(n652), .Z(n649) );
  NAND U571 ( .A(n653), .B(n654), .Z(n652) );
  NANDN U572 ( .A(A[93]), .B(B[93]), .Z(n654) );
  AND U573 ( .A(n655), .B(n656), .Z(n653) );
  NANDN U574 ( .A(A[92]), .B(B[92]), .Z(n656) );
  NAND U575 ( .A(n657), .B(n658), .Z(n655) );
  NANDN U576 ( .A(B[92]), .B(A[92]), .Z(n658) );
  AND U577 ( .A(n659), .B(n660), .Z(n657) );
  NAND U578 ( .A(n661), .B(n662), .Z(n660) );
  NANDN U579 ( .A(A[91]), .B(B[91]), .Z(n662) );
  AND U580 ( .A(n663), .B(n664), .Z(n661) );
  NANDN U581 ( .A(A[90]), .B(B[90]), .Z(n664) );
  NAND U582 ( .A(n665), .B(n666), .Z(n663) );
  NANDN U583 ( .A(B[90]), .B(A[90]), .Z(n666) );
  AND U584 ( .A(n667), .B(n668), .Z(n665) );
  NAND U585 ( .A(n669), .B(n670), .Z(n668) );
  NANDN U586 ( .A(A[89]), .B(B[89]), .Z(n670) );
  AND U587 ( .A(n671), .B(n672), .Z(n669) );
  NANDN U588 ( .A(A[88]), .B(B[88]), .Z(n672) );
  NAND U589 ( .A(n673), .B(n674), .Z(n671) );
  NANDN U590 ( .A(B[88]), .B(A[88]), .Z(n674) );
  AND U591 ( .A(n675), .B(n676), .Z(n673) );
  NAND U592 ( .A(n677), .B(n678), .Z(n676) );
  NANDN U593 ( .A(A[87]), .B(B[87]), .Z(n678) );
  AND U594 ( .A(n679), .B(n680), .Z(n677) );
  NANDN U595 ( .A(A[86]), .B(B[86]), .Z(n680) );
  NAND U596 ( .A(n681), .B(n682), .Z(n679) );
  NANDN U597 ( .A(B[86]), .B(A[86]), .Z(n682) );
  AND U598 ( .A(n683), .B(n684), .Z(n681) );
  NAND U599 ( .A(n685), .B(n686), .Z(n684) );
  NANDN U600 ( .A(A[85]), .B(B[85]), .Z(n686) );
  AND U601 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U602 ( .A(A[84]), .B(B[84]), .Z(n688) );
  NAND U603 ( .A(n689), .B(n690), .Z(n687) );
  NANDN U604 ( .A(B[84]), .B(A[84]), .Z(n690) );
  AND U605 ( .A(n691), .B(n692), .Z(n689) );
  NAND U606 ( .A(n693), .B(n694), .Z(n692) );
  NANDN U607 ( .A(A[83]), .B(B[83]), .Z(n694) );
  AND U608 ( .A(n695), .B(n696), .Z(n693) );
  NANDN U609 ( .A(A[82]), .B(B[82]), .Z(n696) );
  NAND U610 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U611 ( .A(B[82]), .B(A[82]), .Z(n698) );
  AND U612 ( .A(n699), .B(n700), .Z(n697) );
  NAND U613 ( .A(n701), .B(n702), .Z(n700) );
  NANDN U614 ( .A(A[81]), .B(B[81]), .Z(n702) );
  AND U615 ( .A(n703), .B(n704), .Z(n701) );
  NANDN U616 ( .A(A[80]), .B(B[80]), .Z(n704) );
  NAND U617 ( .A(n705), .B(n706), .Z(n703) );
  NANDN U618 ( .A(B[80]), .B(A[80]), .Z(n706) );
  AND U619 ( .A(n707), .B(n708), .Z(n705) );
  NAND U620 ( .A(n709), .B(n710), .Z(n708) );
  NANDN U621 ( .A(A[79]), .B(B[79]), .Z(n710) );
  AND U622 ( .A(n711), .B(n712), .Z(n709) );
  NANDN U623 ( .A(A[78]), .B(B[78]), .Z(n712) );
  NAND U624 ( .A(n713), .B(n714), .Z(n711) );
  NANDN U625 ( .A(B[78]), .B(A[78]), .Z(n714) );
  AND U626 ( .A(n715), .B(n716), .Z(n713) );
  NAND U627 ( .A(n717), .B(n718), .Z(n716) );
  NANDN U628 ( .A(A[77]), .B(B[77]), .Z(n718) );
  AND U629 ( .A(n719), .B(n720), .Z(n717) );
  NANDN U630 ( .A(A[76]), .B(B[76]), .Z(n720) );
  NAND U631 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U632 ( .A(B[76]), .B(A[76]), .Z(n722) );
  AND U633 ( .A(n723), .B(n724), .Z(n721) );
  NAND U634 ( .A(n725), .B(n726), .Z(n724) );
  NANDN U635 ( .A(A[75]), .B(B[75]), .Z(n726) );
  AND U636 ( .A(n727), .B(n728), .Z(n725) );
  NANDN U637 ( .A(A[74]), .B(B[74]), .Z(n728) );
  NAND U638 ( .A(n729), .B(n730), .Z(n727) );
  NANDN U639 ( .A(B[74]), .B(A[74]), .Z(n730) );
  AND U640 ( .A(n731), .B(n732), .Z(n729) );
  NAND U641 ( .A(n733), .B(n734), .Z(n732) );
  NANDN U642 ( .A(A[73]), .B(B[73]), .Z(n734) );
  AND U643 ( .A(n735), .B(n736), .Z(n733) );
  NANDN U644 ( .A(A[72]), .B(B[72]), .Z(n736) );
  NAND U645 ( .A(n737), .B(n738), .Z(n735) );
  NANDN U646 ( .A(B[72]), .B(A[72]), .Z(n738) );
  AND U647 ( .A(n739), .B(n740), .Z(n737) );
  NAND U648 ( .A(n741), .B(n742), .Z(n740) );
  NANDN U649 ( .A(A[71]), .B(B[71]), .Z(n742) );
  AND U650 ( .A(n743), .B(n744), .Z(n741) );
  NANDN U651 ( .A(A[70]), .B(B[70]), .Z(n744) );
  NAND U652 ( .A(n745), .B(n746), .Z(n743) );
  NANDN U653 ( .A(B[70]), .B(A[70]), .Z(n746) );
  AND U654 ( .A(n747), .B(n748), .Z(n745) );
  NAND U655 ( .A(n749), .B(n750), .Z(n748) );
  NANDN U656 ( .A(A[69]), .B(B[69]), .Z(n750) );
  AND U657 ( .A(n751), .B(n752), .Z(n749) );
  NANDN U658 ( .A(A[68]), .B(B[68]), .Z(n752) );
  NAND U659 ( .A(n753), .B(n754), .Z(n751) );
  NANDN U660 ( .A(B[68]), .B(A[68]), .Z(n754) );
  AND U661 ( .A(n755), .B(n756), .Z(n753) );
  NAND U662 ( .A(n757), .B(n758), .Z(n756) );
  NANDN U663 ( .A(A[67]), .B(B[67]), .Z(n758) );
  AND U664 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U665 ( .A(A[66]), .B(B[66]), .Z(n760) );
  NAND U666 ( .A(n761), .B(n762), .Z(n759) );
  NANDN U667 ( .A(B[66]), .B(A[66]), .Z(n762) );
  AND U668 ( .A(n763), .B(n764), .Z(n761) );
  NAND U669 ( .A(n765), .B(n766), .Z(n764) );
  NANDN U670 ( .A(A[65]), .B(B[65]), .Z(n766) );
  AND U671 ( .A(n767), .B(n768), .Z(n765) );
  NANDN U672 ( .A(A[64]), .B(B[64]), .Z(n768) );
  NAND U673 ( .A(n769), .B(n770), .Z(n767) );
  NANDN U674 ( .A(B[64]), .B(A[64]), .Z(n770) );
  AND U675 ( .A(n771), .B(n772), .Z(n769) );
  NAND U676 ( .A(n773), .B(n774), .Z(n772) );
  NANDN U677 ( .A(A[63]), .B(B[63]), .Z(n774) );
  AND U678 ( .A(n775), .B(n776), .Z(n773) );
  NANDN U679 ( .A(A[62]), .B(B[62]), .Z(n776) );
  NAND U680 ( .A(n777), .B(n778), .Z(n775) );
  NANDN U681 ( .A(B[62]), .B(A[62]), .Z(n778) );
  AND U682 ( .A(n779), .B(n780), .Z(n777) );
  NAND U683 ( .A(n781), .B(n782), .Z(n780) );
  NANDN U684 ( .A(A[61]), .B(B[61]), .Z(n782) );
  AND U685 ( .A(n783), .B(n784), .Z(n781) );
  NANDN U686 ( .A(A[60]), .B(B[60]), .Z(n784) );
  NAND U687 ( .A(n785), .B(n786), .Z(n783) );
  NANDN U688 ( .A(B[60]), .B(A[60]), .Z(n786) );
  AND U689 ( .A(n787), .B(n788), .Z(n785) );
  NAND U690 ( .A(n789), .B(n790), .Z(n788) );
  NANDN U691 ( .A(A[59]), .B(B[59]), .Z(n790) );
  AND U692 ( .A(n791), .B(n792), .Z(n789) );
  NANDN U693 ( .A(A[58]), .B(B[58]), .Z(n792) );
  NAND U694 ( .A(n793), .B(n794), .Z(n791) );
  NANDN U695 ( .A(B[58]), .B(A[58]), .Z(n794) );
  AND U696 ( .A(n795), .B(n796), .Z(n793) );
  NAND U697 ( .A(n797), .B(n798), .Z(n796) );
  NANDN U698 ( .A(A[57]), .B(B[57]), .Z(n798) );
  AND U699 ( .A(n799), .B(n800), .Z(n797) );
  NANDN U700 ( .A(A[56]), .B(B[56]), .Z(n800) );
  NAND U701 ( .A(n801), .B(n802), .Z(n799) );
  NANDN U702 ( .A(B[56]), .B(A[56]), .Z(n802) );
  AND U703 ( .A(n803), .B(n804), .Z(n801) );
  NAND U704 ( .A(n805), .B(n806), .Z(n804) );
  NANDN U705 ( .A(A[55]), .B(B[55]), .Z(n806) );
  AND U706 ( .A(n807), .B(n808), .Z(n805) );
  NANDN U707 ( .A(A[54]), .B(B[54]), .Z(n808) );
  NAND U708 ( .A(n809), .B(n810), .Z(n807) );
  NANDN U709 ( .A(B[54]), .B(A[54]), .Z(n810) );
  AND U710 ( .A(n811), .B(n812), .Z(n809) );
  NAND U711 ( .A(n813), .B(n814), .Z(n812) );
  NANDN U712 ( .A(A[53]), .B(B[53]), .Z(n814) );
  AND U713 ( .A(n815), .B(n816), .Z(n813) );
  NANDN U714 ( .A(A[52]), .B(B[52]), .Z(n816) );
  NAND U715 ( .A(n817), .B(n818), .Z(n815) );
  NANDN U716 ( .A(B[52]), .B(A[52]), .Z(n818) );
  AND U717 ( .A(n819), .B(n820), .Z(n817) );
  NAND U718 ( .A(n821), .B(n822), .Z(n820) );
  NANDN U719 ( .A(A[51]), .B(B[51]), .Z(n822) );
  AND U720 ( .A(n823), .B(n824), .Z(n821) );
  NANDN U721 ( .A(A[50]), .B(B[50]), .Z(n824) );
  NAND U722 ( .A(n825), .B(n826), .Z(n823) );
  NANDN U723 ( .A(B[50]), .B(A[50]), .Z(n826) );
  AND U724 ( .A(n827), .B(n828), .Z(n825) );
  NAND U725 ( .A(n829), .B(n830), .Z(n828) );
  NANDN U726 ( .A(A[49]), .B(B[49]), .Z(n830) );
  AND U727 ( .A(n831), .B(n832), .Z(n829) );
  NANDN U728 ( .A(A[48]), .B(B[48]), .Z(n832) );
  NAND U729 ( .A(n833), .B(n834), .Z(n831) );
  NANDN U730 ( .A(B[48]), .B(A[48]), .Z(n834) );
  AND U731 ( .A(n835), .B(n836), .Z(n833) );
  NAND U732 ( .A(n837), .B(n838), .Z(n836) );
  NANDN U733 ( .A(A[47]), .B(B[47]), .Z(n838) );
  AND U734 ( .A(n839), .B(n840), .Z(n837) );
  NANDN U735 ( .A(A[46]), .B(B[46]), .Z(n840) );
  NAND U736 ( .A(n841), .B(n842), .Z(n839) );
  NANDN U737 ( .A(B[46]), .B(A[46]), .Z(n842) );
  AND U738 ( .A(n843), .B(n844), .Z(n841) );
  NAND U739 ( .A(n845), .B(n846), .Z(n844) );
  NANDN U740 ( .A(A[45]), .B(B[45]), .Z(n846) );
  AND U741 ( .A(n847), .B(n848), .Z(n845) );
  NANDN U742 ( .A(A[44]), .B(B[44]), .Z(n848) );
  NAND U743 ( .A(n849), .B(n850), .Z(n847) );
  NANDN U744 ( .A(B[44]), .B(A[44]), .Z(n850) );
  AND U745 ( .A(n851), .B(n852), .Z(n849) );
  NAND U746 ( .A(n853), .B(n854), .Z(n852) );
  NANDN U747 ( .A(A[43]), .B(B[43]), .Z(n854) );
  AND U748 ( .A(n855), .B(n856), .Z(n853) );
  NANDN U749 ( .A(A[42]), .B(B[42]), .Z(n856) );
  NAND U750 ( .A(n857), .B(n858), .Z(n855) );
  NANDN U751 ( .A(B[42]), .B(A[42]), .Z(n858) );
  AND U752 ( .A(n859), .B(n860), .Z(n857) );
  NAND U753 ( .A(n861), .B(n862), .Z(n860) );
  NANDN U754 ( .A(A[41]), .B(B[41]), .Z(n862) );
  AND U755 ( .A(n863), .B(n864), .Z(n861) );
  NANDN U756 ( .A(A[40]), .B(B[40]), .Z(n864) );
  NAND U757 ( .A(n865), .B(n866), .Z(n863) );
  NANDN U758 ( .A(B[40]), .B(A[40]), .Z(n866) );
  AND U759 ( .A(n867), .B(n868), .Z(n865) );
  NAND U760 ( .A(n869), .B(n870), .Z(n868) );
  NANDN U761 ( .A(A[39]), .B(B[39]), .Z(n870) );
  AND U762 ( .A(n871), .B(n872), .Z(n869) );
  NANDN U763 ( .A(A[38]), .B(B[38]), .Z(n872) );
  NAND U764 ( .A(n873), .B(n874), .Z(n871) );
  NANDN U765 ( .A(B[38]), .B(A[38]), .Z(n874) );
  AND U766 ( .A(n875), .B(n876), .Z(n873) );
  NAND U767 ( .A(n877), .B(n878), .Z(n876) );
  NANDN U768 ( .A(A[37]), .B(B[37]), .Z(n878) );
  AND U769 ( .A(n879), .B(n880), .Z(n877) );
  NANDN U770 ( .A(A[36]), .B(B[36]), .Z(n880) );
  NAND U771 ( .A(n881), .B(n882), .Z(n879) );
  NANDN U772 ( .A(B[36]), .B(A[36]), .Z(n882) );
  AND U773 ( .A(n883), .B(n884), .Z(n881) );
  NAND U774 ( .A(n885), .B(n886), .Z(n884) );
  NANDN U775 ( .A(A[35]), .B(B[35]), .Z(n886) );
  AND U776 ( .A(n887), .B(n888), .Z(n885) );
  NANDN U777 ( .A(A[34]), .B(B[34]), .Z(n888) );
  NAND U778 ( .A(n889), .B(n890), .Z(n887) );
  NANDN U779 ( .A(B[34]), .B(A[34]), .Z(n890) );
  AND U780 ( .A(n891), .B(n892), .Z(n889) );
  NAND U781 ( .A(n893), .B(n894), .Z(n892) );
  NANDN U782 ( .A(A[33]), .B(B[33]), .Z(n894) );
  AND U783 ( .A(n895), .B(n896), .Z(n893) );
  NANDN U784 ( .A(A[32]), .B(B[32]), .Z(n896) );
  NAND U785 ( .A(n897), .B(n898), .Z(n895) );
  NANDN U786 ( .A(B[32]), .B(A[32]), .Z(n898) );
  AND U787 ( .A(n899), .B(n900), .Z(n897) );
  NAND U788 ( .A(n901), .B(n902), .Z(n900) );
  NANDN U789 ( .A(A[31]), .B(B[31]), .Z(n902) );
  AND U790 ( .A(n903), .B(n904), .Z(n901) );
  NANDN U791 ( .A(A[30]), .B(B[30]), .Z(n904) );
  NAND U792 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U793 ( .A(B[30]), .B(A[30]), .Z(n906) );
  AND U794 ( .A(n907), .B(n908), .Z(n905) );
  NAND U795 ( .A(n909), .B(n910), .Z(n908) );
  NANDN U796 ( .A(A[29]), .B(B[29]), .Z(n910) );
  AND U797 ( .A(n911), .B(n912), .Z(n909) );
  NANDN U798 ( .A(A[28]), .B(B[28]), .Z(n912) );
  NAND U799 ( .A(n913), .B(n914), .Z(n911) );
  NANDN U800 ( .A(B[28]), .B(A[28]), .Z(n914) );
  AND U801 ( .A(n915), .B(n916), .Z(n913) );
  NAND U802 ( .A(n917), .B(n918), .Z(n916) );
  NANDN U803 ( .A(A[27]), .B(B[27]), .Z(n918) );
  AND U804 ( .A(n919), .B(n920), .Z(n917) );
  NANDN U805 ( .A(A[26]), .B(B[26]), .Z(n920) );
  NAND U806 ( .A(n921), .B(n922), .Z(n919) );
  NANDN U807 ( .A(B[26]), .B(A[26]), .Z(n922) );
  AND U808 ( .A(n923), .B(n924), .Z(n921) );
  NAND U809 ( .A(n925), .B(n926), .Z(n924) );
  NANDN U810 ( .A(A[25]), .B(B[25]), .Z(n926) );
  AND U811 ( .A(n927), .B(n928), .Z(n925) );
  NANDN U812 ( .A(A[24]), .B(B[24]), .Z(n928) );
  NAND U813 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U814 ( .A(B[24]), .B(A[24]), .Z(n930) );
  AND U815 ( .A(n931), .B(n932), .Z(n929) );
  NAND U816 ( .A(n933), .B(n934), .Z(n932) );
  NANDN U817 ( .A(A[23]), .B(B[23]), .Z(n934) );
  AND U818 ( .A(n935), .B(n936), .Z(n933) );
  NANDN U819 ( .A(A[22]), .B(B[22]), .Z(n936) );
  NAND U820 ( .A(n937), .B(n938), .Z(n935) );
  NANDN U821 ( .A(B[22]), .B(A[22]), .Z(n938) );
  AND U822 ( .A(n939), .B(n940), .Z(n937) );
  NAND U823 ( .A(n941), .B(n942), .Z(n940) );
  NANDN U824 ( .A(A[21]), .B(B[21]), .Z(n942) );
  AND U825 ( .A(n943), .B(n944), .Z(n941) );
  NANDN U826 ( .A(A[20]), .B(B[20]), .Z(n944) );
  NAND U827 ( .A(n945), .B(n946), .Z(n943) );
  NANDN U828 ( .A(B[20]), .B(A[20]), .Z(n946) );
  AND U829 ( .A(n947), .B(n948), .Z(n945) );
  NAND U830 ( .A(n949), .B(n950), .Z(n948) );
  NANDN U831 ( .A(A[19]), .B(B[19]), .Z(n950) );
  AND U832 ( .A(n951), .B(n952), .Z(n949) );
  NANDN U833 ( .A(A[18]), .B(B[18]), .Z(n952) );
  NAND U834 ( .A(n953), .B(n954), .Z(n951) );
  NANDN U835 ( .A(B[18]), .B(A[18]), .Z(n954) );
  AND U836 ( .A(n955), .B(n956), .Z(n953) );
  NAND U837 ( .A(n957), .B(n958), .Z(n956) );
  NANDN U838 ( .A(A[17]), .B(B[17]), .Z(n958) );
  AND U839 ( .A(n959), .B(n960), .Z(n957) );
  NANDN U840 ( .A(A[16]), .B(B[16]), .Z(n960) );
  NAND U841 ( .A(n961), .B(n962), .Z(n959) );
  NANDN U842 ( .A(B[16]), .B(A[16]), .Z(n962) );
  AND U843 ( .A(n963), .B(n964), .Z(n961) );
  NAND U844 ( .A(n965), .B(n966), .Z(n964) );
  NANDN U845 ( .A(A[15]), .B(B[15]), .Z(n966) );
  AND U846 ( .A(n967), .B(n968), .Z(n965) );
  NANDN U847 ( .A(A[14]), .B(B[14]), .Z(n968) );
  NAND U848 ( .A(n969), .B(n970), .Z(n967) );
  NANDN U849 ( .A(B[14]), .B(A[14]), .Z(n970) );
  AND U850 ( .A(n971), .B(n972), .Z(n969) );
  NAND U851 ( .A(n973), .B(n974), .Z(n972) );
  NANDN U852 ( .A(A[13]), .B(B[13]), .Z(n974) );
  AND U853 ( .A(n975), .B(n976), .Z(n973) );
  NANDN U854 ( .A(A[12]), .B(B[12]), .Z(n976) );
  NAND U855 ( .A(n977), .B(n978), .Z(n975) );
  NANDN U856 ( .A(B[12]), .B(A[12]), .Z(n978) );
  AND U857 ( .A(n979), .B(n980), .Z(n977) );
  NAND U858 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U859 ( .A(A[11]), .B(B[11]), .Z(n982) );
  AND U860 ( .A(n983), .B(n984), .Z(n981) );
  NANDN U861 ( .A(A[10]), .B(B[10]), .Z(n984) );
  NAND U862 ( .A(n985), .B(n986), .Z(n983) );
  NANDN U863 ( .A(B[9]), .B(A[9]), .Z(n986) );
  AND U864 ( .A(n987), .B(n988), .Z(n985) );
  NAND U865 ( .A(n989), .B(n990), .Z(n988) );
  NANDN U866 ( .A(A[9]), .B(B[9]), .Z(n990) );
  AND U867 ( .A(n991), .B(n992), .Z(n989) );
  NANDN U868 ( .A(A[8]), .B(B[8]), .Z(n992) );
  NAND U869 ( .A(n993), .B(n994), .Z(n991) );
  NANDN U870 ( .A(B[8]), .B(A[8]), .Z(n994) );
  AND U871 ( .A(n995), .B(n996), .Z(n993) );
  NAND U872 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U873 ( .A(A[7]), .B(B[7]), .Z(n998) );
  AND U874 ( .A(n999), .B(n1000), .Z(n997) );
  NANDN U875 ( .A(A[6]), .B(B[6]), .Z(n1000) );
  NAND U876 ( .A(n1001), .B(n1002), .Z(n999) );
  NANDN U877 ( .A(B[6]), .B(A[6]), .Z(n1002) );
  AND U878 ( .A(n1003), .B(n1004), .Z(n1001) );
  NAND U879 ( .A(n1005), .B(n1006), .Z(n1004) );
  NANDN U880 ( .A(A[5]), .B(B[5]), .Z(n1006) );
  AND U881 ( .A(n1007), .B(n1008), .Z(n1005) );
  NANDN U882 ( .A(A[4]), .B(B[4]), .Z(n1008) );
  NAND U883 ( .A(n1009), .B(n1010), .Z(n1007) );
  NANDN U884 ( .A(B[4]), .B(A[4]), .Z(n1010) );
  AND U885 ( .A(n1011), .B(n1012), .Z(n1009) );
  NAND U886 ( .A(n1013), .B(n1014), .Z(n1012) );
  NANDN U887 ( .A(A[3]), .B(B[3]), .Z(n1014) );
  AND U888 ( .A(n1015), .B(n1016), .Z(n1013) );
  NANDN U889 ( .A(A[2]), .B(B[2]), .Z(n1016) );
  NAND U890 ( .A(n1017), .B(n1018), .Z(n1015) );
  NANDN U891 ( .A(B[2]), .B(A[2]), .Z(n1018) );
  AND U892 ( .A(n1019), .B(n1020), .Z(n1017) );
  NANDN U893 ( .A(B[1]), .B(n1021), .Z(n1020) );
  NANDN U894 ( .A(A[1]), .B(n1022), .Z(n1021) );
  NANDN U895 ( .A(n1022), .B(A[1]), .Z(n1019) );
  ANDN U896 ( .B(B[0]), .A(A[0]), .Z(n1022) );
  NANDN U897 ( .A(B[3]), .B(A[3]), .Z(n1011) );
  NANDN U898 ( .A(B[5]), .B(A[5]), .Z(n1003) );
  NANDN U899 ( .A(B[7]), .B(A[7]), .Z(n995) );
  NANDN U900 ( .A(B[10]), .B(A[10]), .Z(n987) );
  NANDN U901 ( .A(B[11]), .B(A[11]), .Z(n979) );
  NANDN U902 ( .A(B[13]), .B(A[13]), .Z(n971) );
  NANDN U903 ( .A(B[15]), .B(A[15]), .Z(n963) );
  NANDN U904 ( .A(B[17]), .B(A[17]), .Z(n955) );
  NANDN U905 ( .A(B[19]), .B(A[19]), .Z(n947) );
  NANDN U906 ( .A(B[21]), .B(A[21]), .Z(n939) );
  NANDN U907 ( .A(B[23]), .B(A[23]), .Z(n931) );
  NANDN U908 ( .A(B[25]), .B(A[25]), .Z(n923) );
  NANDN U909 ( .A(B[27]), .B(A[27]), .Z(n915) );
  NANDN U910 ( .A(B[29]), .B(A[29]), .Z(n907) );
  NANDN U911 ( .A(B[31]), .B(A[31]), .Z(n899) );
  NANDN U912 ( .A(B[33]), .B(A[33]), .Z(n891) );
  NANDN U913 ( .A(B[35]), .B(A[35]), .Z(n883) );
  NANDN U914 ( .A(B[37]), .B(A[37]), .Z(n875) );
  NANDN U915 ( .A(B[39]), .B(A[39]), .Z(n867) );
  NANDN U916 ( .A(B[41]), .B(A[41]), .Z(n859) );
  NANDN U917 ( .A(B[43]), .B(A[43]), .Z(n851) );
  NANDN U918 ( .A(B[45]), .B(A[45]), .Z(n843) );
  NANDN U919 ( .A(B[47]), .B(A[47]), .Z(n835) );
  NANDN U920 ( .A(B[49]), .B(A[49]), .Z(n827) );
  NANDN U921 ( .A(B[51]), .B(A[51]), .Z(n819) );
  NANDN U922 ( .A(B[53]), .B(A[53]), .Z(n811) );
  NANDN U923 ( .A(B[55]), .B(A[55]), .Z(n803) );
  NANDN U924 ( .A(B[57]), .B(A[57]), .Z(n795) );
  NANDN U925 ( .A(B[59]), .B(A[59]), .Z(n787) );
  NANDN U926 ( .A(B[61]), .B(A[61]), .Z(n779) );
  NANDN U927 ( .A(B[63]), .B(A[63]), .Z(n771) );
  NANDN U928 ( .A(B[65]), .B(A[65]), .Z(n763) );
  NANDN U929 ( .A(B[67]), .B(A[67]), .Z(n755) );
  NANDN U930 ( .A(B[69]), .B(A[69]), .Z(n747) );
  NANDN U931 ( .A(B[71]), .B(A[71]), .Z(n739) );
  NANDN U932 ( .A(B[73]), .B(A[73]), .Z(n731) );
  NANDN U933 ( .A(B[75]), .B(A[75]), .Z(n723) );
  NANDN U934 ( .A(B[77]), .B(A[77]), .Z(n715) );
  NANDN U935 ( .A(B[79]), .B(A[79]), .Z(n707) );
  NANDN U936 ( .A(B[81]), .B(A[81]), .Z(n699) );
  NANDN U937 ( .A(B[83]), .B(A[83]), .Z(n691) );
  NANDN U938 ( .A(B[85]), .B(A[85]), .Z(n683) );
  NANDN U939 ( .A(B[87]), .B(A[87]), .Z(n675) );
  NANDN U940 ( .A(B[89]), .B(A[89]), .Z(n667) );
  NANDN U941 ( .A(B[91]), .B(A[91]), .Z(n659) );
  NANDN U942 ( .A(B[93]), .B(A[93]), .Z(n651) );
  NANDN U943 ( .A(B[95]), .B(A[95]), .Z(n643) );
  NANDN U944 ( .A(B[97]), .B(A[97]), .Z(n635) );
  NANDN U945 ( .A(B[100]), .B(A[100]), .Z(n627) );
  NANDN U946 ( .A(B[101]), .B(A[101]), .Z(n619) );
  NANDN U947 ( .A(B[103]), .B(A[103]), .Z(n611) );
  NANDN U948 ( .A(B[105]), .B(A[105]), .Z(n603) );
  NANDN U949 ( .A(B[107]), .B(A[107]), .Z(n595) );
  NANDN U950 ( .A(B[109]), .B(A[109]), .Z(n587) );
  NANDN U951 ( .A(B[111]), .B(A[111]), .Z(n579) );
  NANDN U952 ( .A(B[113]), .B(A[113]), .Z(n571) );
  NANDN U953 ( .A(B[115]), .B(A[115]), .Z(n563) );
  NANDN U954 ( .A(B[117]), .B(A[117]), .Z(n555) );
  NANDN U955 ( .A(B[119]), .B(A[119]), .Z(n547) );
  NANDN U956 ( .A(B[121]), .B(A[121]), .Z(n539) );
  NANDN U957 ( .A(B[123]), .B(A[123]), .Z(n531) );
  NANDN U958 ( .A(B[125]), .B(A[125]), .Z(n523) );
  NANDN U959 ( .A(B[127]), .B(A[127]), .Z(n515) );
  NANDN U960 ( .A(B[129]), .B(A[129]), .Z(n507) );
  NANDN U961 ( .A(B[131]), .B(A[131]), .Z(n499) );
  NANDN U962 ( .A(B[133]), .B(A[133]), .Z(n491) );
  NANDN U963 ( .A(B[135]), .B(A[135]), .Z(n483) );
  NANDN U964 ( .A(B[137]), .B(A[137]), .Z(n475) );
  NANDN U965 ( .A(B[139]), .B(A[139]), .Z(n467) );
  NANDN U966 ( .A(B[141]), .B(A[141]), .Z(n459) );
  NANDN U967 ( .A(B[143]), .B(A[143]), .Z(n451) );
  NANDN U968 ( .A(B[145]), .B(A[145]), .Z(n443) );
  NANDN U969 ( .A(B[147]), .B(A[147]), .Z(n435) );
  NANDN U970 ( .A(B[149]), .B(A[149]), .Z(n427) );
  NANDN U971 ( .A(B[151]), .B(A[151]), .Z(n419) );
  NANDN U972 ( .A(B[153]), .B(A[153]), .Z(n411) );
  NANDN U973 ( .A(B[155]), .B(A[155]), .Z(n403) );
  NANDN U974 ( .A(B[157]), .B(A[157]), .Z(n395) );
  NANDN U975 ( .A(B[159]), .B(A[159]), .Z(n387) );
  NANDN U976 ( .A(B[161]), .B(A[161]), .Z(n379) );
  NANDN U977 ( .A(B[163]), .B(A[163]), .Z(n371) );
  NANDN U978 ( .A(B[165]), .B(A[165]), .Z(n363) );
  NANDN U979 ( .A(B[167]), .B(A[167]), .Z(n355) );
  NANDN U980 ( .A(B[169]), .B(A[169]), .Z(n347) );
  NANDN U981 ( .A(B[171]), .B(A[171]), .Z(n339) );
  NANDN U982 ( .A(B[173]), .B(A[173]), .Z(n331) );
  NANDN U983 ( .A(B[175]), .B(A[175]), .Z(n323) );
  NANDN U984 ( .A(B[177]), .B(A[177]), .Z(n315) );
  NANDN U985 ( .A(B[179]), .B(A[179]), .Z(n307) );
  NANDN U986 ( .A(B[181]), .B(A[181]), .Z(n299) );
  NANDN U987 ( .A(B[183]), .B(A[183]), .Z(n291) );
  NANDN U988 ( .A(B[185]), .B(A[185]), .Z(n283) );
  NANDN U989 ( .A(B[187]), .B(A[187]), .Z(n275) );
  NANDN U990 ( .A(B[189]), .B(A[189]), .Z(n267) );
  NANDN U991 ( .A(B[191]), .B(A[191]), .Z(n259) );
  NANDN U992 ( .A(B[193]), .B(A[193]), .Z(n251) );
  NANDN U993 ( .A(B[195]), .B(A[195]), .Z(n243) );
  NANDN U994 ( .A(B[197]), .B(A[197]), .Z(n235) );
  NANDN U995 ( .A(B[199]), .B(A[199]), .Z(n227) );
  NANDN U996 ( .A(B[201]), .B(A[201]), .Z(n219) );
  NANDN U997 ( .A(B[203]), .B(A[203]), .Z(n211) );
  NANDN U998 ( .A(B[205]), .B(A[205]), .Z(n203) );
  NANDN U999 ( .A(B[207]), .B(A[207]), .Z(n195) );
  NANDN U1000 ( .A(B[209]), .B(A[209]), .Z(n187) );
  NANDN U1001 ( .A(B[211]), .B(A[211]), .Z(n179) );
  NANDN U1002 ( .A(B[213]), .B(A[213]), .Z(n171) );
  NANDN U1003 ( .A(B[215]), .B(A[215]), .Z(n163) );
  NANDN U1004 ( .A(B[217]), .B(A[217]), .Z(n155) );
  NANDN U1005 ( .A(B[219]), .B(A[219]), .Z(n147) );
  NANDN U1006 ( .A(B[221]), .B(A[221]), .Z(n139) );
  NANDN U1007 ( .A(B[223]), .B(A[223]), .Z(n131) );
  NANDN U1008 ( .A(B[225]), .B(A[225]), .Z(n123) );
  NANDN U1009 ( .A(B[227]), .B(A[227]), .Z(n115) );
  NANDN U1010 ( .A(B[229]), .B(A[229]), .Z(n107) );
  NANDN U1011 ( .A(B[231]), .B(A[231]), .Z(n99) );
  NANDN U1012 ( .A(B[233]), .B(A[233]), .Z(n91) );
  NANDN U1013 ( .A(B[235]), .B(A[235]), .Z(n83) );
  NANDN U1014 ( .A(B[237]), .B(A[237]), .Z(n75) );
  NANDN U1015 ( .A(B[239]), .B(A[239]), .Z(n67) );
  NANDN U1016 ( .A(B[241]), .B(A[241]), .Z(n59) );
  NANDN U1017 ( .A(B[243]), .B(A[243]), .Z(n51) );
  NANDN U1018 ( .A(B[245]), .B(A[245]), .Z(n43) );
  NANDN U1019 ( .A(B[247]), .B(A[247]), .Z(n35) );
  NANDN U1020 ( .A(B[249]), .B(A[249]), .Z(n27) );
  NANDN U1021 ( .A(B[251]), .B(A[251]), .Z(n19) );
  NANDN U1022 ( .A(B[253]), .B(A[253]), .Z(n11) );
  NANDN U1023 ( .A(A[255]), .B(B[255]), .Z(n3) );
endmodule


module modmult_step_N256_2_DW01_add_0 ( A, B, CI, SUM, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] SUM;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272;
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];

  XNOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(SUM[99]) );
  XNOR U4 ( .A(B[99]), .B(A[99]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[98]) );
  XNOR U6 ( .A(B[98]), .B(A[98]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[97]) );
  XNOR U8 ( .A(B[97]), .B(A[97]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[96]) );
  XNOR U10 ( .A(B[96]), .B(A[96]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[95]) );
  XNOR U12 ( .A(B[95]), .B(A[95]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[94]) );
  XNOR U14 ( .A(B[94]), .B(A[94]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[93]) );
  XNOR U16 ( .A(B[93]), .B(A[93]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(SUM[92]) );
  XNOR U18 ( .A(B[92]), .B(A[92]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(SUM[91]) );
  XNOR U20 ( .A(B[91]), .B(A[91]), .Z(n20) );
  XOR U21 ( .A(n21), .B(n22), .Z(SUM[90]) );
  XNOR U22 ( .A(B[90]), .B(A[90]), .Z(n22) );
  XOR U23 ( .A(n23), .B(n24), .Z(SUM[8]) );
  XNOR U24 ( .A(B[8]), .B(A[8]), .Z(n24) );
  XOR U25 ( .A(n25), .B(n26), .Z(SUM[89]) );
  XNOR U26 ( .A(B[89]), .B(A[89]), .Z(n26) );
  XOR U27 ( .A(n27), .B(n28), .Z(SUM[88]) );
  XNOR U28 ( .A(B[88]), .B(A[88]), .Z(n28) );
  XOR U29 ( .A(n29), .B(n30), .Z(SUM[87]) );
  XNOR U30 ( .A(B[87]), .B(A[87]), .Z(n30) );
  XOR U31 ( .A(n31), .B(n32), .Z(SUM[86]) );
  XNOR U32 ( .A(B[86]), .B(A[86]), .Z(n32) );
  XOR U33 ( .A(n33), .B(n34), .Z(SUM[85]) );
  XNOR U34 ( .A(B[85]), .B(A[85]), .Z(n34) );
  XOR U35 ( .A(n35), .B(n36), .Z(SUM[84]) );
  XNOR U36 ( .A(B[84]), .B(A[84]), .Z(n36) );
  XOR U37 ( .A(n37), .B(n38), .Z(SUM[83]) );
  XNOR U38 ( .A(B[83]), .B(A[83]), .Z(n38) );
  XOR U39 ( .A(n39), .B(n40), .Z(SUM[82]) );
  XNOR U40 ( .A(B[82]), .B(A[82]), .Z(n40) );
  XOR U41 ( .A(n41), .B(n42), .Z(SUM[81]) );
  XNOR U42 ( .A(B[81]), .B(A[81]), .Z(n42) );
  XOR U43 ( .A(n43), .B(n44), .Z(SUM[80]) );
  XNOR U44 ( .A(B[80]), .B(A[80]), .Z(n44) );
  XOR U45 ( .A(n45), .B(n46), .Z(SUM[7]) );
  XNOR U46 ( .A(B[7]), .B(A[7]), .Z(n46) );
  XOR U47 ( .A(n47), .B(n48), .Z(SUM[79]) );
  XNOR U48 ( .A(B[79]), .B(A[79]), .Z(n48) );
  XOR U49 ( .A(n49), .B(n50), .Z(SUM[78]) );
  XNOR U50 ( .A(B[78]), .B(A[78]), .Z(n50) );
  XOR U51 ( .A(n51), .B(n52), .Z(SUM[77]) );
  XNOR U52 ( .A(B[77]), .B(A[77]), .Z(n52) );
  XOR U53 ( .A(n53), .B(n54), .Z(SUM[76]) );
  XNOR U54 ( .A(B[76]), .B(A[76]), .Z(n54) );
  XOR U55 ( .A(n55), .B(n56), .Z(SUM[75]) );
  XNOR U56 ( .A(B[75]), .B(A[75]), .Z(n56) );
  XOR U57 ( .A(n57), .B(n58), .Z(SUM[74]) );
  XNOR U58 ( .A(B[74]), .B(A[74]), .Z(n58) );
  XOR U59 ( .A(n59), .B(n60), .Z(SUM[73]) );
  XNOR U60 ( .A(B[73]), .B(A[73]), .Z(n60) );
  XOR U61 ( .A(n61), .B(n62), .Z(SUM[72]) );
  XNOR U62 ( .A(B[72]), .B(A[72]), .Z(n62) );
  XOR U63 ( .A(n63), .B(n64), .Z(SUM[71]) );
  XNOR U64 ( .A(B[71]), .B(A[71]), .Z(n64) );
  XOR U65 ( .A(n65), .B(n66), .Z(SUM[70]) );
  XNOR U66 ( .A(B[70]), .B(A[70]), .Z(n66) );
  XOR U67 ( .A(n67), .B(n68), .Z(SUM[6]) );
  XNOR U68 ( .A(B[6]), .B(A[6]), .Z(n68) );
  XOR U69 ( .A(n69), .B(n70), .Z(SUM[69]) );
  XNOR U70 ( .A(B[69]), .B(A[69]), .Z(n70) );
  XOR U71 ( .A(n71), .B(n72), .Z(SUM[68]) );
  XNOR U72 ( .A(B[68]), .B(A[68]), .Z(n72) );
  XOR U73 ( .A(n73), .B(n74), .Z(SUM[67]) );
  XNOR U74 ( .A(B[67]), .B(A[67]), .Z(n74) );
  XOR U75 ( .A(n75), .B(n76), .Z(SUM[66]) );
  XNOR U76 ( .A(B[66]), .B(A[66]), .Z(n76) );
  XOR U77 ( .A(n77), .B(n78), .Z(SUM[65]) );
  XNOR U78 ( .A(B[65]), .B(A[65]), .Z(n78) );
  XOR U79 ( .A(n79), .B(n80), .Z(SUM[64]) );
  XNOR U80 ( .A(B[64]), .B(A[64]), .Z(n80) );
  XOR U81 ( .A(n81), .B(n82), .Z(SUM[63]) );
  XNOR U82 ( .A(B[63]), .B(A[63]), .Z(n82) );
  XOR U83 ( .A(n83), .B(n84), .Z(SUM[62]) );
  XNOR U84 ( .A(B[62]), .B(A[62]), .Z(n84) );
  XOR U85 ( .A(n85), .B(n86), .Z(SUM[61]) );
  XNOR U86 ( .A(B[61]), .B(A[61]), .Z(n86) );
  XOR U87 ( .A(n87), .B(n88), .Z(SUM[60]) );
  XNOR U88 ( .A(B[60]), .B(A[60]), .Z(n88) );
  XOR U89 ( .A(n89), .B(n90), .Z(SUM[5]) );
  XNOR U90 ( .A(B[5]), .B(A[5]), .Z(n90) );
  XOR U91 ( .A(n91), .B(n92), .Z(SUM[59]) );
  XNOR U92 ( .A(B[59]), .B(A[59]), .Z(n92) );
  XOR U93 ( .A(n93), .B(n94), .Z(SUM[58]) );
  XNOR U94 ( .A(B[58]), .B(A[58]), .Z(n94) );
  XOR U95 ( .A(n95), .B(n96), .Z(SUM[57]) );
  XNOR U96 ( .A(B[57]), .B(A[57]), .Z(n96) );
  XOR U97 ( .A(n97), .B(n98), .Z(SUM[56]) );
  XNOR U98 ( .A(B[56]), .B(A[56]), .Z(n98) );
  XOR U99 ( .A(n99), .B(n100), .Z(SUM[55]) );
  XNOR U100 ( .A(B[55]), .B(A[55]), .Z(n100) );
  XOR U101 ( .A(n101), .B(n102), .Z(SUM[54]) );
  XNOR U102 ( .A(B[54]), .B(A[54]), .Z(n102) );
  XOR U103 ( .A(n103), .B(n104), .Z(SUM[53]) );
  XNOR U104 ( .A(B[53]), .B(A[53]), .Z(n104) );
  XOR U105 ( .A(n105), .B(n106), .Z(SUM[52]) );
  XNOR U106 ( .A(B[52]), .B(A[52]), .Z(n106) );
  XOR U107 ( .A(n107), .B(n108), .Z(SUM[51]) );
  XNOR U108 ( .A(B[51]), .B(A[51]), .Z(n108) );
  XOR U109 ( .A(n109), .B(n110), .Z(SUM[50]) );
  XNOR U110 ( .A(B[50]), .B(A[50]), .Z(n110) );
  XOR U111 ( .A(n111), .B(n112), .Z(SUM[4]) );
  XNOR U112 ( .A(B[4]), .B(A[4]), .Z(n112) );
  XOR U113 ( .A(n113), .B(n114), .Z(SUM[49]) );
  XNOR U114 ( .A(B[49]), .B(A[49]), .Z(n114) );
  XOR U115 ( .A(n115), .B(n116), .Z(SUM[48]) );
  XNOR U116 ( .A(B[48]), .B(A[48]), .Z(n116) );
  XOR U117 ( .A(n117), .B(n118), .Z(SUM[47]) );
  XNOR U118 ( .A(B[47]), .B(A[47]), .Z(n118) );
  XOR U119 ( .A(n119), .B(n120), .Z(SUM[46]) );
  XNOR U120 ( .A(B[46]), .B(A[46]), .Z(n120) );
  XOR U121 ( .A(n121), .B(n122), .Z(SUM[45]) );
  XNOR U122 ( .A(B[45]), .B(A[45]), .Z(n122) );
  XOR U123 ( .A(n123), .B(n124), .Z(SUM[44]) );
  XNOR U124 ( .A(B[44]), .B(A[44]), .Z(n124) );
  XOR U125 ( .A(n125), .B(n126), .Z(SUM[43]) );
  XNOR U126 ( .A(B[43]), .B(A[43]), .Z(n126) );
  XOR U127 ( .A(n127), .B(n128), .Z(SUM[42]) );
  XNOR U128 ( .A(B[42]), .B(A[42]), .Z(n128) );
  XOR U129 ( .A(n129), .B(n130), .Z(SUM[41]) );
  XNOR U130 ( .A(B[41]), .B(A[41]), .Z(n130) );
  XOR U131 ( .A(n131), .B(n132), .Z(SUM[40]) );
  XNOR U132 ( .A(B[40]), .B(A[40]), .Z(n132) );
  XOR U133 ( .A(n133), .B(n134), .Z(SUM[3]) );
  XNOR U134 ( .A(B[3]), .B(A[3]), .Z(n134) );
  XOR U135 ( .A(n135), .B(n136), .Z(SUM[39]) );
  XNOR U136 ( .A(B[39]), .B(A[39]), .Z(n136) );
  XOR U137 ( .A(n137), .B(n138), .Z(SUM[38]) );
  XNOR U138 ( .A(B[38]), .B(A[38]), .Z(n138) );
  XOR U139 ( .A(n139), .B(n140), .Z(SUM[37]) );
  XNOR U140 ( .A(B[37]), .B(A[37]), .Z(n140) );
  XOR U141 ( .A(n141), .B(n142), .Z(SUM[36]) );
  XNOR U142 ( .A(B[36]), .B(A[36]), .Z(n142) );
  XOR U143 ( .A(n143), .B(n144), .Z(SUM[35]) );
  XNOR U144 ( .A(B[35]), .B(A[35]), .Z(n144) );
  XOR U145 ( .A(n145), .B(n146), .Z(SUM[34]) );
  XNOR U146 ( .A(B[34]), .B(A[34]), .Z(n146) );
  XOR U147 ( .A(n147), .B(n148), .Z(SUM[33]) );
  XNOR U148 ( .A(B[33]), .B(A[33]), .Z(n148) );
  XOR U149 ( .A(n149), .B(n150), .Z(SUM[32]) );
  XNOR U150 ( .A(B[32]), .B(A[32]), .Z(n150) );
  XOR U151 ( .A(n151), .B(n152), .Z(SUM[31]) );
  XNOR U152 ( .A(B[31]), .B(A[31]), .Z(n152) );
  XOR U153 ( .A(n153), .B(n154), .Z(SUM[30]) );
  XNOR U154 ( .A(B[30]), .B(A[30]), .Z(n154) );
  XOR U155 ( .A(n155), .B(n156), .Z(SUM[2]) );
  XOR U156 ( .A(B[2]), .B(A[2]), .Z(n156) );
  XOR U157 ( .A(n157), .B(n158), .Z(SUM[29]) );
  XNOR U158 ( .A(B[29]), .B(A[29]), .Z(n158) );
  XOR U159 ( .A(n159), .B(n160), .Z(SUM[28]) );
  XNOR U160 ( .A(B[28]), .B(A[28]), .Z(n160) );
  XOR U161 ( .A(n161), .B(n162), .Z(SUM[27]) );
  XNOR U162 ( .A(B[27]), .B(A[27]), .Z(n162) );
  XOR U163 ( .A(n163), .B(n164), .Z(SUM[26]) );
  XNOR U164 ( .A(B[26]), .B(A[26]), .Z(n164) );
  XOR U165 ( .A(n165), .B(n166), .Z(SUM[25]) );
  XNOR U166 ( .A(B[25]), .B(A[25]), .Z(n166) );
  XOR U167 ( .A(A[257]), .B(n167), .Z(SUM[257]) );
  AND U168 ( .A(A[256]), .B(n168), .Z(n167) );
  XOR U169 ( .A(A[256]), .B(n168), .Z(SUM[256]) );
  NAND U170 ( .A(n169), .B(n170), .Z(n168) );
  NAND U171 ( .A(B[255]), .B(n171), .Z(n170) );
  NANDN U172 ( .A(A[255]), .B(n172), .Z(n171) );
  NANDN U173 ( .A(n172), .B(A[255]), .Z(n169) );
  XOR U174 ( .A(n172), .B(n173), .Z(SUM[255]) );
  XNOR U175 ( .A(B[255]), .B(A[255]), .Z(n173) );
  AND U176 ( .A(n174), .B(n175), .Z(n172) );
  NAND U177 ( .A(B[254]), .B(n176), .Z(n175) );
  NANDN U178 ( .A(A[254]), .B(n177), .Z(n176) );
  NANDN U179 ( .A(n177), .B(A[254]), .Z(n174) );
  XOR U180 ( .A(n177), .B(n178), .Z(SUM[254]) );
  XNOR U181 ( .A(B[254]), .B(A[254]), .Z(n178) );
  AND U182 ( .A(n179), .B(n180), .Z(n177) );
  NAND U183 ( .A(B[253]), .B(n181), .Z(n180) );
  NANDN U184 ( .A(A[253]), .B(n182), .Z(n181) );
  NANDN U185 ( .A(n182), .B(A[253]), .Z(n179) );
  XOR U186 ( .A(n182), .B(n183), .Z(SUM[253]) );
  XNOR U187 ( .A(B[253]), .B(A[253]), .Z(n183) );
  AND U188 ( .A(n184), .B(n185), .Z(n182) );
  NAND U189 ( .A(B[252]), .B(n186), .Z(n185) );
  NANDN U190 ( .A(A[252]), .B(n187), .Z(n186) );
  NANDN U191 ( .A(n187), .B(A[252]), .Z(n184) );
  XOR U192 ( .A(n187), .B(n188), .Z(SUM[252]) );
  XNOR U193 ( .A(B[252]), .B(A[252]), .Z(n188) );
  AND U194 ( .A(n189), .B(n190), .Z(n187) );
  NAND U195 ( .A(B[251]), .B(n191), .Z(n190) );
  NANDN U196 ( .A(A[251]), .B(n192), .Z(n191) );
  NANDN U197 ( .A(n192), .B(A[251]), .Z(n189) );
  XOR U198 ( .A(n192), .B(n193), .Z(SUM[251]) );
  XNOR U199 ( .A(B[251]), .B(A[251]), .Z(n193) );
  AND U200 ( .A(n194), .B(n195), .Z(n192) );
  NAND U201 ( .A(B[250]), .B(n196), .Z(n195) );
  NANDN U202 ( .A(A[250]), .B(n197), .Z(n196) );
  NANDN U203 ( .A(n197), .B(A[250]), .Z(n194) );
  XOR U204 ( .A(n197), .B(n198), .Z(SUM[250]) );
  XNOR U205 ( .A(B[250]), .B(A[250]), .Z(n198) );
  AND U206 ( .A(n199), .B(n200), .Z(n197) );
  NAND U207 ( .A(B[249]), .B(n201), .Z(n200) );
  NANDN U208 ( .A(A[249]), .B(n202), .Z(n201) );
  NANDN U209 ( .A(n202), .B(A[249]), .Z(n199) );
  XOR U210 ( .A(n203), .B(n204), .Z(SUM[24]) );
  XNOR U211 ( .A(B[24]), .B(A[24]), .Z(n204) );
  XOR U212 ( .A(n202), .B(n205), .Z(SUM[249]) );
  XNOR U213 ( .A(B[249]), .B(A[249]), .Z(n205) );
  AND U214 ( .A(n206), .B(n207), .Z(n202) );
  NAND U215 ( .A(B[248]), .B(n208), .Z(n207) );
  NANDN U216 ( .A(A[248]), .B(n209), .Z(n208) );
  NANDN U217 ( .A(n209), .B(A[248]), .Z(n206) );
  XOR U218 ( .A(n209), .B(n210), .Z(SUM[248]) );
  XNOR U219 ( .A(B[248]), .B(A[248]), .Z(n210) );
  AND U220 ( .A(n211), .B(n212), .Z(n209) );
  NAND U221 ( .A(B[247]), .B(n213), .Z(n212) );
  NANDN U222 ( .A(A[247]), .B(n214), .Z(n213) );
  NANDN U223 ( .A(n214), .B(A[247]), .Z(n211) );
  XOR U224 ( .A(n214), .B(n215), .Z(SUM[247]) );
  XNOR U225 ( .A(B[247]), .B(A[247]), .Z(n215) );
  AND U226 ( .A(n216), .B(n217), .Z(n214) );
  NAND U227 ( .A(B[246]), .B(n218), .Z(n217) );
  NANDN U228 ( .A(A[246]), .B(n219), .Z(n218) );
  NANDN U229 ( .A(n219), .B(A[246]), .Z(n216) );
  XOR U230 ( .A(n219), .B(n220), .Z(SUM[246]) );
  XNOR U231 ( .A(B[246]), .B(A[246]), .Z(n220) );
  AND U232 ( .A(n221), .B(n222), .Z(n219) );
  NAND U233 ( .A(B[245]), .B(n223), .Z(n222) );
  NANDN U234 ( .A(A[245]), .B(n224), .Z(n223) );
  NANDN U235 ( .A(n224), .B(A[245]), .Z(n221) );
  XOR U236 ( .A(n224), .B(n225), .Z(SUM[245]) );
  XNOR U237 ( .A(B[245]), .B(A[245]), .Z(n225) );
  AND U238 ( .A(n226), .B(n227), .Z(n224) );
  NAND U239 ( .A(B[244]), .B(n228), .Z(n227) );
  NANDN U240 ( .A(A[244]), .B(n229), .Z(n228) );
  NANDN U241 ( .A(n229), .B(A[244]), .Z(n226) );
  XOR U242 ( .A(n229), .B(n230), .Z(SUM[244]) );
  XNOR U243 ( .A(B[244]), .B(A[244]), .Z(n230) );
  AND U244 ( .A(n231), .B(n232), .Z(n229) );
  NAND U245 ( .A(B[243]), .B(n233), .Z(n232) );
  NANDN U246 ( .A(A[243]), .B(n234), .Z(n233) );
  NANDN U247 ( .A(n234), .B(A[243]), .Z(n231) );
  XOR U248 ( .A(n234), .B(n235), .Z(SUM[243]) );
  XNOR U249 ( .A(B[243]), .B(A[243]), .Z(n235) );
  AND U250 ( .A(n236), .B(n237), .Z(n234) );
  NAND U251 ( .A(B[242]), .B(n238), .Z(n237) );
  NANDN U252 ( .A(A[242]), .B(n239), .Z(n238) );
  NANDN U253 ( .A(n239), .B(A[242]), .Z(n236) );
  XOR U254 ( .A(n239), .B(n240), .Z(SUM[242]) );
  XNOR U255 ( .A(B[242]), .B(A[242]), .Z(n240) );
  AND U256 ( .A(n241), .B(n242), .Z(n239) );
  NAND U257 ( .A(B[241]), .B(n243), .Z(n242) );
  NANDN U258 ( .A(A[241]), .B(n244), .Z(n243) );
  NANDN U259 ( .A(n244), .B(A[241]), .Z(n241) );
  XOR U260 ( .A(n244), .B(n245), .Z(SUM[241]) );
  XNOR U261 ( .A(B[241]), .B(A[241]), .Z(n245) );
  AND U262 ( .A(n246), .B(n247), .Z(n244) );
  NAND U263 ( .A(B[240]), .B(n248), .Z(n247) );
  NANDN U264 ( .A(A[240]), .B(n249), .Z(n248) );
  NANDN U265 ( .A(n249), .B(A[240]), .Z(n246) );
  XOR U266 ( .A(n249), .B(n250), .Z(SUM[240]) );
  XNOR U267 ( .A(B[240]), .B(A[240]), .Z(n250) );
  AND U268 ( .A(n251), .B(n252), .Z(n249) );
  NAND U269 ( .A(B[239]), .B(n253), .Z(n252) );
  NANDN U270 ( .A(A[239]), .B(n254), .Z(n253) );
  NANDN U271 ( .A(n254), .B(A[239]), .Z(n251) );
  XOR U272 ( .A(n255), .B(n256), .Z(SUM[23]) );
  XNOR U273 ( .A(B[23]), .B(A[23]), .Z(n256) );
  XOR U274 ( .A(n254), .B(n257), .Z(SUM[239]) );
  XNOR U275 ( .A(B[239]), .B(A[239]), .Z(n257) );
  AND U276 ( .A(n258), .B(n259), .Z(n254) );
  NAND U277 ( .A(B[238]), .B(n260), .Z(n259) );
  NANDN U278 ( .A(A[238]), .B(n261), .Z(n260) );
  NANDN U279 ( .A(n261), .B(A[238]), .Z(n258) );
  XOR U280 ( .A(n261), .B(n262), .Z(SUM[238]) );
  XNOR U281 ( .A(B[238]), .B(A[238]), .Z(n262) );
  AND U282 ( .A(n263), .B(n264), .Z(n261) );
  NAND U283 ( .A(B[237]), .B(n265), .Z(n264) );
  NANDN U284 ( .A(A[237]), .B(n266), .Z(n265) );
  NANDN U285 ( .A(n266), .B(A[237]), .Z(n263) );
  XOR U286 ( .A(n266), .B(n267), .Z(SUM[237]) );
  XNOR U287 ( .A(B[237]), .B(A[237]), .Z(n267) );
  AND U288 ( .A(n268), .B(n269), .Z(n266) );
  NAND U289 ( .A(B[236]), .B(n270), .Z(n269) );
  NANDN U290 ( .A(A[236]), .B(n271), .Z(n270) );
  NANDN U291 ( .A(n271), .B(A[236]), .Z(n268) );
  XOR U292 ( .A(n271), .B(n272), .Z(SUM[236]) );
  XNOR U293 ( .A(B[236]), .B(A[236]), .Z(n272) );
  AND U294 ( .A(n273), .B(n274), .Z(n271) );
  NAND U295 ( .A(B[235]), .B(n275), .Z(n274) );
  NANDN U296 ( .A(A[235]), .B(n276), .Z(n275) );
  NANDN U297 ( .A(n276), .B(A[235]), .Z(n273) );
  XOR U298 ( .A(n276), .B(n277), .Z(SUM[235]) );
  XNOR U299 ( .A(B[235]), .B(A[235]), .Z(n277) );
  AND U300 ( .A(n278), .B(n279), .Z(n276) );
  NAND U301 ( .A(B[234]), .B(n280), .Z(n279) );
  NANDN U302 ( .A(A[234]), .B(n281), .Z(n280) );
  NANDN U303 ( .A(n281), .B(A[234]), .Z(n278) );
  XOR U304 ( .A(n281), .B(n282), .Z(SUM[234]) );
  XNOR U305 ( .A(B[234]), .B(A[234]), .Z(n282) );
  AND U306 ( .A(n283), .B(n284), .Z(n281) );
  NAND U307 ( .A(B[233]), .B(n285), .Z(n284) );
  NANDN U308 ( .A(A[233]), .B(n286), .Z(n285) );
  NANDN U309 ( .A(n286), .B(A[233]), .Z(n283) );
  XOR U310 ( .A(n286), .B(n287), .Z(SUM[233]) );
  XNOR U311 ( .A(B[233]), .B(A[233]), .Z(n287) );
  AND U312 ( .A(n288), .B(n289), .Z(n286) );
  NAND U313 ( .A(B[232]), .B(n290), .Z(n289) );
  NANDN U314 ( .A(A[232]), .B(n291), .Z(n290) );
  NANDN U315 ( .A(n291), .B(A[232]), .Z(n288) );
  XOR U316 ( .A(n291), .B(n292), .Z(SUM[232]) );
  XNOR U317 ( .A(B[232]), .B(A[232]), .Z(n292) );
  AND U318 ( .A(n293), .B(n294), .Z(n291) );
  NAND U319 ( .A(B[231]), .B(n295), .Z(n294) );
  NANDN U320 ( .A(A[231]), .B(n296), .Z(n295) );
  NANDN U321 ( .A(n296), .B(A[231]), .Z(n293) );
  XOR U322 ( .A(n296), .B(n297), .Z(SUM[231]) );
  XNOR U323 ( .A(B[231]), .B(A[231]), .Z(n297) );
  AND U324 ( .A(n298), .B(n299), .Z(n296) );
  NAND U325 ( .A(B[230]), .B(n300), .Z(n299) );
  NANDN U326 ( .A(A[230]), .B(n301), .Z(n300) );
  NANDN U327 ( .A(n301), .B(A[230]), .Z(n298) );
  XOR U328 ( .A(n301), .B(n302), .Z(SUM[230]) );
  XNOR U329 ( .A(B[230]), .B(A[230]), .Z(n302) );
  AND U330 ( .A(n303), .B(n304), .Z(n301) );
  NAND U331 ( .A(B[229]), .B(n305), .Z(n304) );
  NANDN U332 ( .A(A[229]), .B(n306), .Z(n305) );
  NANDN U333 ( .A(n306), .B(A[229]), .Z(n303) );
  XOR U334 ( .A(n307), .B(n308), .Z(SUM[22]) );
  XNOR U335 ( .A(B[22]), .B(A[22]), .Z(n308) );
  XOR U336 ( .A(n306), .B(n309), .Z(SUM[229]) );
  XNOR U337 ( .A(B[229]), .B(A[229]), .Z(n309) );
  AND U338 ( .A(n310), .B(n311), .Z(n306) );
  NAND U339 ( .A(B[228]), .B(n312), .Z(n311) );
  NANDN U340 ( .A(A[228]), .B(n313), .Z(n312) );
  NANDN U341 ( .A(n313), .B(A[228]), .Z(n310) );
  XOR U342 ( .A(n313), .B(n314), .Z(SUM[228]) );
  XNOR U343 ( .A(B[228]), .B(A[228]), .Z(n314) );
  AND U344 ( .A(n315), .B(n316), .Z(n313) );
  NAND U345 ( .A(B[227]), .B(n317), .Z(n316) );
  NANDN U346 ( .A(A[227]), .B(n318), .Z(n317) );
  NANDN U347 ( .A(n318), .B(A[227]), .Z(n315) );
  XOR U348 ( .A(n318), .B(n319), .Z(SUM[227]) );
  XNOR U349 ( .A(B[227]), .B(A[227]), .Z(n319) );
  AND U350 ( .A(n320), .B(n321), .Z(n318) );
  NAND U351 ( .A(B[226]), .B(n322), .Z(n321) );
  NANDN U352 ( .A(A[226]), .B(n323), .Z(n322) );
  NANDN U353 ( .A(n323), .B(A[226]), .Z(n320) );
  XOR U354 ( .A(n323), .B(n324), .Z(SUM[226]) );
  XNOR U355 ( .A(B[226]), .B(A[226]), .Z(n324) );
  AND U356 ( .A(n325), .B(n326), .Z(n323) );
  NAND U357 ( .A(B[225]), .B(n327), .Z(n326) );
  NANDN U358 ( .A(A[225]), .B(n328), .Z(n327) );
  NANDN U359 ( .A(n328), .B(A[225]), .Z(n325) );
  XOR U360 ( .A(n328), .B(n329), .Z(SUM[225]) );
  XNOR U361 ( .A(B[225]), .B(A[225]), .Z(n329) );
  AND U362 ( .A(n330), .B(n331), .Z(n328) );
  NAND U363 ( .A(B[224]), .B(n332), .Z(n331) );
  NANDN U364 ( .A(A[224]), .B(n333), .Z(n332) );
  NANDN U365 ( .A(n333), .B(A[224]), .Z(n330) );
  XOR U366 ( .A(n333), .B(n334), .Z(SUM[224]) );
  XNOR U367 ( .A(B[224]), .B(A[224]), .Z(n334) );
  AND U368 ( .A(n335), .B(n336), .Z(n333) );
  NAND U369 ( .A(B[223]), .B(n337), .Z(n336) );
  NANDN U370 ( .A(A[223]), .B(n338), .Z(n337) );
  NANDN U371 ( .A(n338), .B(A[223]), .Z(n335) );
  XOR U372 ( .A(n338), .B(n339), .Z(SUM[223]) );
  XNOR U373 ( .A(B[223]), .B(A[223]), .Z(n339) );
  AND U374 ( .A(n340), .B(n341), .Z(n338) );
  NAND U375 ( .A(B[222]), .B(n342), .Z(n341) );
  NANDN U376 ( .A(A[222]), .B(n343), .Z(n342) );
  NANDN U377 ( .A(n343), .B(A[222]), .Z(n340) );
  XOR U378 ( .A(n343), .B(n344), .Z(SUM[222]) );
  XNOR U379 ( .A(B[222]), .B(A[222]), .Z(n344) );
  AND U380 ( .A(n345), .B(n346), .Z(n343) );
  NAND U381 ( .A(B[221]), .B(n347), .Z(n346) );
  NANDN U382 ( .A(A[221]), .B(n348), .Z(n347) );
  NANDN U383 ( .A(n348), .B(A[221]), .Z(n345) );
  XOR U384 ( .A(n348), .B(n349), .Z(SUM[221]) );
  XNOR U385 ( .A(B[221]), .B(A[221]), .Z(n349) );
  AND U386 ( .A(n350), .B(n351), .Z(n348) );
  NAND U387 ( .A(B[220]), .B(n352), .Z(n351) );
  NANDN U388 ( .A(A[220]), .B(n353), .Z(n352) );
  NANDN U389 ( .A(n353), .B(A[220]), .Z(n350) );
  XOR U390 ( .A(n353), .B(n354), .Z(SUM[220]) );
  XNOR U391 ( .A(B[220]), .B(A[220]), .Z(n354) );
  AND U392 ( .A(n355), .B(n356), .Z(n353) );
  NAND U393 ( .A(B[219]), .B(n357), .Z(n356) );
  NANDN U394 ( .A(A[219]), .B(n358), .Z(n357) );
  NANDN U395 ( .A(n358), .B(A[219]), .Z(n355) );
  XOR U396 ( .A(n359), .B(n360), .Z(SUM[21]) );
  XNOR U397 ( .A(B[21]), .B(A[21]), .Z(n360) );
  XOR U398 ( .A(n358), .B(n361), .Z(SUM[219]) );
  XNOR U399 ( .A(B[219]), .B(A[219]), .Z(n361) );
  AND U400 ( .A(n362), .B(n363), .Z(n358) );
  NAND U401 ( .A(B[218]), .B(n364), .Z(n363) );
  NANDN U402 ( .A(A[218]), .B(n365), .Z(n364) );
  NANDN U403 ( .A(n365), .B(A[218]), .Z(n362) );
  XOR U404 ( .A(n365), .B(n366), .Z(SUM[218]) );
  XNOR U405 ( .A(B[218]), .B(A[218]), .Z(n366) );
  AND U406 ( .A(n367), .B(n368), .Z(n365) );
  NAND U407 ( .A(B[217]), .B(n369), .Z(n368) );
  NANDN U408 ( .A(A[217]), .B(n370), .Z(n369) );
  NANDN U409 ( .A(n370), .B(A[217]), .Z(n367) );
  XOR U410 ( .A(n370), .B(n371), .Z(SUM[217]) );
  XNOR U411 ( .A(B[217]), .B(A[217]), .Z(n371) );
  AND U412 ( .A(n372), .B(n373), .Z(n370) );
  NAND U413 ( .A(B[216]), .B(n374), .Z(n373) );
  NANDN U414 ( .A(A[216]), .B(n375), .Z(n374) );
  NANDN U415 ( .A(n375), .B(A[216]), .Z(n372) );
  XOR U416 ( .A(n375), .B(n376), .Z(SUM[216]) );
  XNOR U417 ( .A(B[216]), .B(A[216]), .Z(n376) );
  AND U418 ( .A(n377), .B(n378), .Z(n375) );
  NAND U419 ( .A(B[215]), .B(n379), .Z(n378) );
  NANDN U420 ( .A(A[215]), .B(n380), .Z(n379) );
  NANDN U421 ( .A(n380), .B(A[215]), .Z(n377) );
  XOR U422 ( .A(n380), .B(n381), .Z(SUM[215]) );
  XNOR U423 ( .A(B[215]), .B(A[215]), .Z(n381) );
  AND U424 ( .A(n382), .B(n383), .Z(n380) );
  NAND U425 ( .A(B[214]), .B(n384), .Z(n383) );
  NANDN U426 ( .A(A[214]), .B(n385), .Z(n384) );
  NANDN U427 ( .A(n385), .B(A[214]), .Z(n382) );
  XOR U428 ( .A(n385), .B(n386), .Z(SUM[214]) );
  XNOR U429 ( .A(B[214]), .B(A[214]), .Z(n386) );
  AND U430 ( .A(n387), .B(n388), .Z(n385) );
  NAND U431 ( .A(B[213]), .B(n389), .Z(n388) );
  NANDN U432 ( .A(A[213]), .B(n390), .Z(n389) );
  NANDN U433 ( .A(n390), .B(A[213]), .Z(n387) );
  XOR U434 ( .A(n390), .B(n391), .Z(SUM[213]) );
  XNOR U435 ( .A(B[213]), .B(A[213]), .Z(n391) );
  AND U436 ( .A(n392), .B(n393), .Z(n390) );
  NAND U437 ( .A(B[212]), .B(n394), .Z(n393) );
  NANDN U438 ( .A(A[212]), .B(n395), .Z(n394) );
  NANDN U439 ( .A(n395), .B(A[212]), .Z(n392) );
  XOR U440 ( .A(n395), .B(n396), .Z(SUM[212]) );
  XNOR U441 ( .A(B[212]), .B(A[212]), .Z(n396) );
  AND U442 ( .A(n397), .B(n398), .Z(n395) );
  NAND U443 ( .A(B[211]), .B(n399), .Z(n398) );
  NANDN U444 ( .A(A[211]), .B(n400), .Z(n399) );
  NANDN U445 ( .A(n400), .B(A[211]), .Z(n397) );
  XOR U446 ( .A(n400), .B(n401), .Z(SUM[211]) );
  XNOR U447 ( .A(B[211]), .B(A[211]), .Z(n401) );
  AND U448 ( .A(n402), .B(n403), .Z(n400) );
  NAND U449 ( .A(B[210]), .B(n404), .Z(n403) );
  NANDN U450 ( .A(A[210]), .B(n405), .Z(n404) );
  NANDN U451 ( .A(n405), .B(A[210]), .Z(n402) );
  XOR U452 ( .A(n405), .B(n406), .Z(SUM[210]) );
  XNOR U453 ( .A(B[210]), .B(A[210]), .Z(n406) );
  AND U454 ( .A(n407), .B(n408), .Z(n405) );
  NAND U455 ( .A(B[209]), .B(n409), .Z(n408) );
  NANDN U456 ( .A(A[209]), .B(n410), .Z(n409) );
  NANDN U457 ( .A(n410), .B(A[209]), .Z(n407) );
  XOR U458 ( .A(n411), .B(n412), .Z(SUM[20]) );
  XNOR U459 ( .A(B[20]), .B(A[20]), .Z(n412) );
  XOR U460 ( .A(n410), .B(n413), .Z(SUM[209]) );
  XNOR U461 ( .A(B[209]), .B(A[209]), .Z(n413) );
  AND U462 ( .A(n414), .B(n415), .Z(n410) );
  NAND U463 ( .A(B[208]), .B(n416), .Z(n415) );
  NANDN U464 ( .A(A[208]), .B(n417), .Z(n416) );
  NANDN U465 ( .A(n417), .B(A[208]), .Z(n414) );
  XOR U466 ( .A(n417), .B(n418), .Z(SUM[208]) );
  XNOR U467 ( .A(B[208]), .B(A[208]), .Z(n418) );
  AND U468 ( .A(n419), .B(n420), .Z(n417) );
  NAND U469 ( .A(B[207]), .B(n421), .Z(n420) );
  NANDN U470 ( .A(A[207]), .B(n422), .Z(n421) );
  NANDN U471 ( .A(n422), .B(A[207]), .Z(n419) );
  XOR U472 ( .A(n422), .B(n423), .Z(SUM[207]) );
  XNOR U473 ( .A(B[207]), .B(A[207]), .Z(n423) );
  AND U474 ( .A(n424), .B(n425), .Z(n422) );
  NAND U475 ( .A(B[206]), .B(n426), .Z(n425) );
  NANDN U476 ( .A(A[206]), .B(n427), .Z(n426) );
  NANDN U477 ( .A(n427), .B(A[206]), .Z(n424) );
  XOR U478 ( .A(n427), .B(n428), .Z(SUM[206]) );
  XNOR U479 ( .A(B[206]), .B(A[206]), .Z(n428) );
  AND U480 ( .A(n429), .B(n430), .Z(n427) );
  NAND U481 ( .A(B[205]), .B(n431), .Z(n430) );
  NANDN U482 ( .A(A[205]), .B(n432), .Z(n431) );
  NANDN U483 ( .A(n432), .B(A[205]), .Z(n429) );
  XOR U484 ( .A(n432), .B(n433), .Z(SUM[205]) );
  XNOR U485 ( .A(B[205]), .B(A[205]), .Z(n433) );
  AND U486 ( .A(n434), .B(n435), .Z(n432) );
  NAND U487 ( .A(B[204]), .B(n436), .Z(n435) );
  NANDN U488 ( .A(A[204]), .B(n437), .Z(n436) );
  NANDN U489 ( .A(n437), .B(A[204]), .Z(n434) );
  XOR U490 ( .A(n437), .B(n438), .Z(SUM[204]) );
  XNOR U491 ( .A(B[204]), .B(A[204]), .Z(n438) );
  AND U492 ( .A(n439), .B(n440), .Z(n437) );
  NAND U493 ( .A(B[203]), .B(n441), .Z(n440) );
  NANDN U494 ( .A(A[203]), .B(n442), .Z(n441) );
  NANDN U495 ( .A(n442), .B(A[203]), .Z(n439) );
  XOR U496 ( .A(n442), .B(n443), .Z(SUM[203]) );
  XNOR U497 ( .A(B[203]), .B(A[203]), .Z(n443) );
  AND U498 ( .A(n444), .B(n445), .Z(n442) );
  NAND U499 ( .A(B[202]), .B(n446), .Z(n445) );
  NANDN U500 ( .A(A[202]), .B(n447), .Z(n446) );
  NANDN U501 ( .A(n447), .B(A[202]), .Z(n444) );
  XOR U502 ( .A(n447), .B(n448), .Z(SUM[202]) );
  XNOR U503 ( .A(B[202]), .B(A[202]), .Z(n448) );
  AND U504 ( .A(n449), .B(n450), .Z(n447) );
  NAND U505 ( .A(B[201]), .B(n451), .Z(n450) );
  NANDN U506 ( .A(A[201]), .B(n452), .Z(n451) );
  NANDN U507 ( .A(n452), .B(A[201]), .Z(n449) );
  XOR U508 ( .A(n452), .B(n453), .Z(SUM[201]) );
  XNOR U509 ( .A(B[201]), .B(A[201]), .Z(n453) );
  AND U510 ( .A(n454), .B(n455), .Z(n452) );
  NAND U511 ( .A(B[200]), .B(n456), .Z(n455) );
  NANDN U512 ( .A(A[200]), .B(n457), .Z(n456) );
  NANDN U513 ( .A(n457), .B(A[200]), .Z(n454) );
  XOR U514 ( .A(n457), .B(n458), .Z(SUM[200]) );
  XNOR U515 ( .A(B[200]), .B(A[200]), .Z(n458) );
  AND U516 ( .A(n459), .B(n460), .Z(n457) );
  NAND U517 ( .A(B[199]), .B(n461), .Z(n460) );
  NANDN U518 ( .A(A[199]), .B(n462), .Z(n461) );
  NANDN U519 ( .A(n462), .B(A[199]), .Z(n459) );
  XOR U520 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  XOR U521 ( .A(n463), .B(n464), .Z(SUM[19]) );
  XNOR U522 ( .A(B[19]), .B(A[19]), .Z(n464) );
  XOR U523 ( .A(n462), .B(n465), .Z(SUM[199]) );
  XNOR U524 ( .A(B[199]), .B(A[199]), .Z(n465) );
  AND U525 ( .A(n466), .B(n467), .Z(n462) );
  NAND U526 ( .A(B[198]), .B(n468), .Z(n467) );
  NANDN U527 ( .A(A[198]), .B(n469), .Z(n468) );
  NANDN U528 ( .A(n469), .B(A[198]), .Z(n466) );
  XOR U529 ( .A(n469), .B(n470), .Z(SUM[198]) );
  XNOR U530 ( .A(B[198]), .B(A[198]), .Z(n470) );
  AND U531 ( .A(n471), .B(n472), .Z(n469) );
  NAND U532 ( .A(B[197]), .B(n473), .Z(n472) );
  NANDN U533 ( .A(A[197]), .B(n474), .Z(n473) );
  NANDN U534 ( .A(n474), .B(A[197]), .Z(n471) );
  XOR U535 ( .A(n474), .B(n475), .Z(SUM[197]) );
  XNOR U536 ( .A(B[197]), .B(A[197]), .Z(n475) );
  AND U537 ( .A(n476), .B(n477), .Z(n474) );
  NAND U538 ( .A(B[196]), .B(n478), .Z(n477) );
  NANDN U539 ( .A(A[196]), .B(n479), .Z(n478) );
  NANDN U540 ( .A(n479), .B(A[196]), .Z(n476) );
  XOR U541 ( .A(n479), .B(n480), .Z(SUM[196]) );
  XNOR U542 ( .A(B[196]), .B(A[196]), .Z(n480) );
  AND U543 ( .A(n481), .B(n482), .Z(n479) );
  NAND U544 ( .A(B[195]), .B(n483), .Z(n482) );
  NANDN U545 ( .A(A[195]), .B(n484), .Z(n483) );
  NANDN U546 ( .A(n484), .B(A[195]), .Z(n481) );
  XOR U547 ( .A(n484), .B(n485), .Z(SUM[195]) );
  XNOR U548 ( .A(B[195]), .B(A[195]), .Z(n485) );
  AND U549 ( .A(n486), .B(n487), .Z(n484) );
  NAND U550 ( .A(B[194]), .B(n488), .Z(n487) );
  NANDN U551 ( .A(A[194]), .B(n489), .Z(n488) );
  NANDN U552 ( .A(n489), .B(A[194]), .Z(n486) );
  XOR U553 ( .A(n489), .B(n490), .Z(SUM[194]) );
  XNOR U554 ( .A(B[194]), .B(A[194]), .Z(n490) );
  AND U555 ( .A(n491), .B(n492), .Z(n489) );
  NAND U556 ( .A(B[193]), .B(n493), .Z(n492) );
  NANDN U557 ( .A(A[193]), .B(n494), .Z(n493) );
  NANDN U558 ( .A(n494), .B(A[193]), .Z(n491) );
  XOR U559 ( .A(n494), .B(n495), .Z(SUM[193]) );
  XNOR U560 ( .A(B[193]), .B(A[193]), .Z(n495) );
  AND U561 ( .A(n496), .B(n497), .Z(n494) );
  NAND U562 ( .A(B[192]), .B(n498), .Z(n497) );
  NANDN U563 ( .A(A[192]), .B(n499), .Z(n498) );
  NANDN U564 ( .A(n499), .B(A[192]), .Z(n496) );
  XOR U565 ( .A(n499), .B(n500), .Z(SUM[192]) );
  XNOR U566 ( .A(B[192]), .B(A[192]), .Z(n500) );
  AND U567 ( .A(n501), .B(n502), .Z(n499) );
  NAND U568 ( .A(B[191]), .B(n503), .Z(n502) );
  NANDN U569 ( .A(A[191]), .B(n504), .Z(n503) );
  NANDN U570 ( .A(n504), .B(A[191]), .Z(n501) );
  XOR U571 ( .A(n504), .B(n505), .Z(SUM[191]) );
  XNOR U572 ( .A(B[191]), .B(A[191]), .Z(n505) );
  AND U573 ( .A(n506), .B(n507), .Z(n504) );
  NAND U574 ( .A(B[190]), .B(n508), .Z(n507) );
  NANDN U575 ( .A(A[190]), .B(n509), .Z(n508) );
  NANDN U576 ( .A(n509), .B(A[190]), .Z(n506) );
  XOR U577 ( .A(n509), .B(n510), .Z(SUM[190]) );
  XNOR U578 ( .A(B[190]), .B(A[190]), .Z(n510) );
  AND U579 ( .A(n511), .B(n512), .Z(n509) );
  NAND U580 ( .A(B[189]), .B(n513), .Z(n512) );
  NANDN U581 ( .A(A[189]), .B(n514), .Z(n513) );
  NANDN U582 ( .A(n514), .B(A[189]), .Z(n511) );
  XOR U583 ( .A(n515), .B(n516), .Z(SUM[18]) );
  XNOR U584 ( .A(B[18]), .B(A[18]), .Z(n516) );
  XOR U585 ( .A(n514), .B(n517), .Z(SUM[189]) );
  XNOR U586 ( .A(B[189]), .B(A[189]), .Z(n517) );
  AND U587 ( .A(n518), .B(n519), .Z(n514) );
  NAND U588 ( .A(B[188]), .B(n520), .Z(n519) );
  NANDN U589 ( .A(A[188]), .B(n521), .Z(n520) );
  NANDN U590 ( .A(n521), .B(A[188]), .Z(n518) );
  XOR U591 ( .A(n521), .B(n522), .Z(SUM[188]) );
  XNOR U592 ( .A(B[188]), .B(A[188]), .Z(n522) );
  AND U593 ( .A(n523), .B(n524), .Z(n521) );
  NAND U594 ( .A(B[187]), .B(n525), .Z(n524) );
  NANDN U595 ( .A(A[187]), .B(n526), .Z(n525) );
  NANDN U596 ( .A(n526), .B(A[187]), .Z(n523) );
  XOR U597 ( .A(n526), .B(n527), .Z(SUM[187]) );
  XNOR U598 ( .A(B[187]), .B(A[187]), .Z(n527) );
  AND U599 ( .A(n528), .B(n529), .Z(n526) );
  NAND U600 ( .A(B[186]), .B(n530), .Z(n529) );
  NANDN U601 ( .A(A[186]), .B(n531), .Z(n530) );
  NANDN U602 ( .A(n531), .B(A[186]), .Z(n528) );
  XOR U603 ( .A(n531), .B(n532), .Z(SUM[186]) );
  XNOR U604 ( .A(B[186]), .B(A[186]), .Z(n532) );
  AND U605 ( .A(n533), .B(n534), .Z(n531) );
  NAND U606 ( .A(B[185]), .B(n535), .Z(n534) );
  NANDN U607 ( .A(A[185]), .B(n536), .Z(n535) );
  NANDN U608 ( .A(n536), .B(A[185]), .Z(n533) );
  XOR U609 ( .A(n536), .B(n537), .Z(SUM[185]) );
  XNOR U610 ( .A(B[185]), .B(A[185]), .Z(n537) );
  AND U611 ( .A(n538), .B(n539), .Z(n536) );
  NAND U612 ( .A(B[184]), .B(n540), .Z(n539) );
  NANDN U613 ( .A(A[184]), .B(n541), .Z(n540) );
  NANDN U614 ( .A(n541), .B(A[184]), .Z(n538) );
  XOR U615 ( .A(n541), .B(n542), .Z(SUM[184]) );
  XNOR U616 ( .A(B[184]), .B(A[184]), .Z(n542) );
  AND U617 ( .A(n543), .B(n544), .Z(n541) );
  NAND U618 ( .A(B[183]), .B(n545), .Z(n544) );
  NANDN U619 ( .A(A[183]), .B(n546), .Z(n545) );
  NANDN U620 ( .A(n546), .B(A[183]), .Z(n543) );
  XOR U621 ( .A(n546), .B(n547), .Z(SUM[183]) );
  XNOR U622 ( .A(B[183]), .B(A[183]), .Z(n547) );
  AND U623 ( .A(n548), .B(n549), .Z(n546) );
  NAND U624 ( .A(B[182]), .B(n550), .Z(n549) );
  NANDN U625 ( .A(A[182]), .B(n551), .Z(n550) );
  NANDN U626 ( .A(n551), .B(A[182]), .Z(n548) );
  XOR U627 ( .A(n551), .B(n552), .Z(SUM[182]) );
  XNOR U628 ( .A(B[182]), .B(A[182]), .Z(n552) );
  AND U629 ( .A(n553), .B(n554), .Z(n551) );
  NAND U630 ( .A(B[181]), .B(n555), .Z(n554) );
  NANDN U631 ( .A(A[181]), .B(n556), .Z(n555) );
  NANDN U632 ( .A(n556), .B(A[181]), .Z(n553) );
  XOR U633 ( .A(n556), .B(n557), .Z(SUM[181]) );
  XNOR U634 ( .A(B[181]), .B(A[181]), .Z(n557) );
  AND U635 ( .A(n558), .B(n559), .Z(n556) );
  NAND U636 ( .A(B[180]), .B(n560), .Z(n559) );
  NANDN U637 ( .A(A[180]), .B(n561), .Z(n560) );
  NANDN U638 ( .A(n561), .B(A[180]), .Z(n558) );
  XOR U639 ( .A(n561), .B(n562), .Z(SUM[180]) );
  XNOR U640 ( .A(B[180]), .B(A[180]), .Z(n562) );
  AND U641 ( .A(n563), .B(n564), .Z(n561) );
  NAND U642 ( .A(B[179]), .B(n565), .Z(n564) );
  NANDN U643 ( .A(A[179]), .B(n566), .Z(n565) );
  NANDN U644 ( .A(n566), .B(A[179]), .Z(n563) );
  XOR U645 ( .A(n567), .B(n568), .Z(SUM[17]) );
  XNOR U646 ( .A(B[17]), .B(A[17]), .Z(n568) );
  XOR U647 ( .A(n566), .B(n569), .Z(SUM[179]) );
  XNOR U648 ( .A(B[179]), .B(A[179]), .Z(n569) );
  AND U649 ( .A(n570), .B(n571), .Z(n566) );
  NAND U650 ( .A(B[178]), .B(n572), .Z(n571) );
  NANDN U651 ( .A(A[178]), .B(n573), .Z(n572) );
  NANDN U652 ( .A(n573), .B(A[178]), .Z(n570) );
  XOR U653 ( .A(n573), .B(n574), .Z(SUM[178]) );
  XNOR U654 ( .A(B[178]), .B(A[178]), .Z(n574) );
  AND U655 ( .A(n575), .B(n576), .Z(n573) );
  NAND U656 ( .A(B[177]), .B(n577), .Z(n576) );
  NANDN U657 ( .A(A[177]), .B(n578), .Z(n577) );
  NANDN U658 ( .A(n578), .B(A[177]), .Z(n575) );
  XOR U659 ( .A(n578), .B(n579), .Z(SUM[177]) );
  XNOR U660 ( .A(B[177]), .B(A[177]), .Z(n579) );
  AND U661 ( .A(n580), .B(n581), .Z(n578) );
  NAND U662 ( .A(B[176]), .B(n582), .Z(n581) );
  NANDN U663 ( .A(A[176]), .B(n583), .Z(n582) );
  NANDN U664 ( .A(n583), .B(A[176]), .Z(n580) );
  XOR U665 ( .A(n583), .B(n584), .Z(SUM[176]) );
  XNOR U666 ( .A(B[176]), .B(A[176]), .Z(n584) );
  AND U667 ( .A(n585), .B(n586), .Z(n583) );
  NAND U668 ( .A(B[175]), .B(n587), .Z(n586) );
  NANDN U669 ( .A(A[175]), .B(n588), .Z(n587) );
  NANDN U670 ( .A(n588), .B(A[175]), .Z(n585) );
  XOR U671 ( .A(n588), .B(n589), .Z(SUM[175]) );
  XNOR U672 ( .A(B[175]), .B(A[175]), .Z(n589) );
  AND U673 ( .A(n590), .B(n591), .Z(n588) );
  NAND U674 ( .A(B[174]), .B(n592), .Z(n591) );
  NANDN U675 ( .A(A[174]), .B(n593), .Z(n592) );
  NANDN U676 ( .A(n593), .B(A[174]), .Z(n590) );
  XOR U677 ( .A(n593), .B(n594), .Z(SUM[174]) );
  XNOR U678 ( .A(B[174]), .B(A[174]), .Z(n594) );
  AND U679 ( .A(n595), .B(n596), .Z(n593) );
  NAND U680 ( .A(B[173]), .B(n597), .Z(n596) );
  NANDN U681 ( .A(A[173]), .B(n598), .Z(n597) );
  NANDN U682 ( .A(n598), .B(A[173]), .Z(n595) );
  XOR U683 ( .A(n598), .B(n599), .Z(SUM[173]) );
  XNOR U684 ( .A(B[173]), .B(A[173]), .Z(n599) );
  AND U685 ( .A(n600), .B(n601), .Z(n598) );
  NAND U686 ( .A(B[172]), .B(n602), .Z(n601) );
  NANDN U687 ( .A(A[172]), .B(n603), .Z(n602) );
  NANDN U688 ( .A(n603), .B(A[172]), .Z(n600) );
  XOR U689 ( .A(n603), .B(n604), .Z(SUM[172]) );
  XNOR U690 ( .A(B[172]), .B(A[172]), .Z(n604) );
  AND U691 ( .A(n605), .B(n606), .Z(n603) );
  NAND U692 ( .A(B[171]), .B(n607), .Z(n606) );
  NANDN U693 ( .A(A[171]), .B(n608), .Z(n607) );
  NANDN U694 ( .A(n608), .B(A[171]), .Z(n605) );
  XOR U695 ( .A(n608), .B(n609), .Z(SUM[171]) );
  XNOR U696 ( .A(B[171]), .B(A[171]), .Z(n609) );
  AND U697 ( .A(n610), .B(n611), .Z(n608) );
  NAND U698 ( .A(B[170]), .B(n612), .Z(n611) );
  NANDN U699 ( .A(A[170]), .B(n613), .Z(n612) );
  NANDN U700 ( .A(n613), .B(A[170]), .Z(n610) );
  XOR U701 ( .A(n613), .B(n614), .Z(SUM[170]) );
  XNOR U702 ( .A(B[170]), .B(A[170]), .Z(n614) );
  AND U703 ( .A(n615), .B(n616), .Z(n613) );
  NAND U704 ( .A(B[169]), .B(n617), .Z(n616) );
  NANDN U705 ( .A(A[169]), .B(n618), .Z(n617) );
  NANDN U706 ( .A(n618), .B(A[169]), .Z(n615) );
  XOR U707 ( .A(n619), .B(n620), .Z(SUM[16]) );
  XNOR U708 ( .A(B[16]), .B(A[16]), .Z(n620) );
  XOR U709 ( .A(n618), .B(n621), .Z(SUM[169]) );
  XNOR U710 ( .A(B[169]), .B(A[169]), .Z(n621) );
  AND U711 ( .A(n622), .B(n623), .Z(n618) );
  NAND U712 ( .A(B[168]), .B(n624), .Z(n623) );
  NANDN U713 ( .A(A[168]), .B(n625), .Z(n624) );
  NANDN U714 ( .A(n625), .B(A[168]), .Z(n622) );
  XOR U715 ( .A(n625), .B(n626), .Z(SUM[168]) );
  XNOR U716 ( .A(B[168]), .B(A[168]), .Z(n626) );
  AND U717 ( .A(n627), .B(n628), .Z(n625) );
  NAND U718 ( .A(B[167]), .B(n629), .Z(n628) );
  NANDN U719 ( .A(A[167]), .B(n630), .Z(n629) );
  NANDN U720 ( .A(n630), .B(A[167]), .Z(n627) );
  XOR U721 ( .A(n630), .B(n631), .Z(SUM[167]) );
  XNOR U722 ( .A(B[167]), .B(A[167]), .Z(n631) );
  AND U723 ( .A(n632), .B(n633), .Z(n630) );
  NAND U724 ( .A(B[166]), .B(n634), .Z(n633) );
  NANDN U725 ( .A(A[166]), .B(n635), .Z(n634) );
  NANDN U726 ( .A(n635), .B(A[166]), .Z(n632) );
  XOR U727 ( .A(n635), .B(n636), .Z(SUM[166]) );
  XNOR U728 ( .A(B[166]), .B(A[166]), .Z(n636) );
  AND U729 ( .A(n637), .B(n638), .Z(n635) );
  NAND U730 ( .A(B[165]), .B(n639), .Z(n638) );
  NANDN U731 ( .A(A[165]), .B(n640), .Z(n639) );
  NANDN U732 ( .A(n640), .B(A[165]), .Z(n637) );
  XOR U733 ( .A(n640), .B(n641), .Z(SUM[165]) );
  XNOR U734 ( .A(B[165]), .B(A[165]), .Z(n641) );
  AND U735 ( .A(n642), .B(n643), .Z(n640) );
  NAND U736 ( .A(B[164]), .B(n644), .Z(n643) );
  NANDN U737 ( .A(A[164]), .B(n645), .Z(n644) );
  NANDN U738 ( .A(n645), .B(A[164]), .Z(n642) );
  XOR U739 ( .A(n645), .B(n646), .Z(SUM[164]) );
  XNOR U740 ( .A(B[164]), .B(A[164]), .Z(n646) );
  AND U741 ( .A(n647), .B(n648), .Z(n645) );
  NAND U742 ( .A(B[163]), .B(n649), .Z(n648) );
  NANDN U743 ( .A(A[163]), .B(n650), .Z(n649) );
  NANDN U744 ( .A(n650), .B(A[163]), .Z(n647) );
  XOR U745 ( .A(n650), .B(n651), .Z(SUM[163]) );
  XNOR U746 ( .A(B[163]), .B(A[163]), .Z(n651) );
  AND U747 ( .A(n652), .B(n653), .Z(n650) );
  NAND U748 ( .A(B[162]), .B(n654), .Z(n653) );
  NANDN U749 ( .A(A[162]), .B(n655), .Z(n654) );
  NANDN U750 ( .A(n655), .B(A[162]), .Z(n652) );
  XOR U751 ( .A(n655), .B(n656), .Z(SUM[162]) );
  XNOR U752 ( .A(B[162]), .B(A[162]), .Z(n656) );
  AND U753 ( .A(n657), .B(n658), .Z(n655) );
  NAND U754 ( .A(B[161]), .B(n659), .Z(n658) );
  NANDN U755 ( .A(A[161]), .B(n660), .Z(n659) );
  NANDN U756 ( .A(n660), .B(A[161]), .Z(n657) );
  XOR U757 ( .A(n660), .B(n661), .Z(SUM[161]) );
  XNOR U758 ( .A(B[161]), .B(A[161]), .Z(n661) );
  AND U759 ( .A(n662), .B(n663), .Z(n660) );
  NAND U760 ( .A(B[160]), .B(n664), .Z(n663) );
  NANDN U761 ( .A(A[160]), .B(n665), .Z(n664) );
  NANDN U762 ( .A(n665), .B(A[160]), .Z(n662) );
  XOR U763 ( .A(n665), .B(n666), .Z(SUM[160]) );
  XNOR U764 ( .A(B[160]), .B(A[160]), .Z(n666) );
  AND U765 ( .A(n667), .B(n668), .Z(n665) );
  NAND U766 ( .A(B[159]), .B(n669), .Z(n668) );
  NANDN U767 ( .A(A[159]), .B(n670), .Z(n669) );
  NANDN U768 ( .A(n670), .B(A[159]), .Z(n667) );
  XOR U769 ( .A(n671), .B(n672), .Z(SUM[15]) );
  XNOR U770 ( .A(B[15]), .B(A[15]), .Z(n672) );
  XOR U771 ( .A(n670), .B(n673), .Z(SUM[159]) );
  XNOR U772 ( .A(B[159]), .B(A[159]), .Z(n673) );
  AND U773 ( .A(n674), .B(n675), .Z(n670) );
  NAND U774 ( .A(B[158]), .B(n676), .Z(n675) );
  NANDN U775 ( .A(A[158]), .B(n677), .Z(n676) );
  NANDN U776 ( .A(n677), .B(A[158]), .Z(n674) );
  XOR U777 ( .A(n677), .B(n678), .Z(SUM[158]) );
  XNOR U778 ( .A(B[158]), .B(A[158]), .Z(n678) );
  AND U779 ( .A(n679), .B(n680), .Z(n677) );
  NAND U780 ( .A(B[157]), .B(n681), .Z(n680) );
  NANDN U781 ( .A(A[157]), .B(n682), .Z(n681) );
  NANDN U782 ( .A(n682), .B(A[157]), .Z(n679) );
  XOR U783 ( .A(n682), .B(n683), .Z(SUM[157]) );
  XNOR U784 ( .A(B[157]), .B(A[157]), .Z(n683) );
  AND U785 ( .A(n684), .B(n685), .Z(n682) );
  NAND U786 ( .A(B[156]), .B(n686), .Z(n685) );
  NANDN U787 ( .A(A[156]), .B(n687), .Z(n686) );
  NANDN U788 ( .A(n687), .B(A[156]), .Z(n684) );
  XOR U789 ( .A(n687), .B(n688), .Z(SUM[156]) );
  XNOR U790 ( .A(B[156]), .B(A[156]), .Z(n688) );
  AND U791 ( .A(n689), .B(n690), .Z(n687) );
  NAND U792 ( .A(B[155]), .B(n691), .Z(n690) );
  NANDN U793 ( .A(A[155]), .B(n692), .Z(n691) );
  NANDN U794 ( .A(n692), .B(A[155]), .Z(n689) );
  XOR U795 ( .A(n692), .B(n693), .Z(SUM[155]) );
  XNOR U796 ( .A(B[155]), .B(A[155]), .Z(n693) );
  AND U797 ( .A(n694), .B(n695), .Z(n692) );
  NAND U798 ( .A(B[154]), .B(n696), .Z(n695) );
  NANDN U799 ( .A(A[154]), .B(n697), .Z(n696) );
  NANDN U800 ( .A(n697), .B(A[154]), .Z(n694) );
  XOR U801 ( .A(n697), .B(n698), .Z(SUM[154]) );
  XNOR U802 ( .A(B[154]), .B(A[154]), .Z(n698) );
  AND U803 ( .A(n699), .B(n700), .Z(n697) );
  NAND U804 ( .A(B[153]), .B(n701), .Z(n700) );
  NANDN U805 ( .A(A[153]), .B(n702), .Z(n701) );
  NANDN U806 ( .A(n702), .B(A[153]), .Z(n699) );
  XOR U807 ( .A(n702), .B(n703), .Z(SUM[153]) );
  XNOR U808 ( .A(B[153]), .B(A[153]), .Z(n703) );
  AND U809 ( .A(n704), .B(n705), .Z(n702) );
  NAND U810 ( .A(B[152]), .B(n706), .Z(n705) );
  NANDN U811 ( .A(A[152]), .B(n707), .Z(n706) );
  NANDN U812 ( .A(n707), .B(A[152]), .Z(n704) );
  XOR U813 ( .A(n707), .B(n708), .Z(SUM[152]) );
  XNOR U814 ( .A(B[152]), .B(A[152]), .Z(n708) );
  AND U815 ( .A(n709), .B(n710), .Z(n707) );
  NAND U816 ( .A(B[151]), .B(n711), .Z(n710) );
  NANDN U817 ( .A(A[151]), .B(n712), .Z(n711) );
  NANDN U818 ( .A(n712), .B(A[151]), .Z(n709) );
  XOR U819 ( .A(n712), .B(n713), .Z(SUM[151]) );
  XNOR U820 ( .A(B[151]), .B(A[151]), .Z(n713) );
  AND U821 ( .A(n714), .B(n715), .Z(n712) );
  NAND U822 ( .A(B[150]), .B(n716), .Z(n715) );
  NANDN U823 ( .A(A[150]), .B(n717), .Z(n716) );
  NANDN U824 ( .A(n717), .B(A[150]), .Z(n714) );
  XOR U825 ( .A(n717), .B(n718), .Z(SUM[150]) );
  XNOR U826 ( .A(B[150]), .B(A[150]), .Z(n718) );
  AND U827 ( .A(n719), .B(n720), .Z(n717) );
  NAND U828 ( .A(B[149]), .B(n721), .Z(n720) );
  NANDN U829 ( .A(A[149]), .B(n722), .Z(n721) );
  NANDN U830 ( .A(n722), .B(A[149]), .Z(n719) );
  XOR U831 ( .A(n723), .B(n724), .Z(SUM[14]) );
  XNOR U832 ( .A(B[14]), .B(A[14]), .Z(n724) );
  XOR U833 ( .A(n722), .B(n725), .Z(SUM[149]) );
  XNOR U834 ( .A(B[149]), .B(A[149]), .Z(n725) );
  AND U835 ( .A(n726), .B(n727), .Z(n722) );
  NAND U836 ( .A(B[148]), .B(n728), .Z(n727) );
  NANDN U837 ( .A(A[148]), .B(n729), .Z(n728) );
  NANDN U838 ( .A(n729), .B(A[148]), .Z(n726) );
  XOR U839 ( .A(n729), .B(n730), .Z(SUM[148]) );
  XNOR U840 ( .A(B[148]), .B(A[148]), .Z(n730) );
  AND U841 ( .A(n731), .B(n732), .Z(n729) );
  NAND U842 ( .A(B[147]), .B(n733), .Z(n732) );
  NANDN U843 ( .A(A[147]), .B(n734), .Z(n733) );
  NANDN U844 ( .A(n734), .B(A[147]), .Z(n731) );
  XOR U845 ( .A(n734), .B(n735), .Z(SUM[147]) );
  XNOR U846 ( .A(B[147]), .B(A[147]), .Z(n735) );
  AND U847 ( .A(n736), .B(n737), .Z(n734) );
  NAND U848 ( .A(B[146]), .B(n738), .Z(n737) );
  NANDN U849 ( .A(A[146]), .B(n739), .Z(n738) );
  NANDN U850 ( .A(n739), .B(A[146]), .Z(n736) );
  XOR U851 ( .A(n739), .B(n740), .Z(SUM[146]) );
  XNOR U852 ( .A(B[146]), .B(A[146]), .Z(n740) );
  AND U853 ( .A(n741), .B(n742), .Z(n739) );
  NAND U854 ( .A(B[145]), .B(n743), .Z(n742) );
  NANDN U855 ( .A(A[145]), .B(n744), .Z(n743) );
  NANDN U856 ( .A(n744), .B(A[145]), .Z(n741) );
  XOR U857 ( .A(n744), .B(n745), .Z(SUM[145]) );
  XNOR U858 ( .A(B[145]), .B(A[145]), .Z(n745) );
  AND U859 ( .A(n746), .B(n747), .Z(n744) );
  NAND U860 ( .A(B[144]), .B(n748), .Z(n747) );
  NANDN U861 ( .A(A[144]), .B(n749), .Z(n748) );
  NANDN U862 ( .A(n749), .B(A[144]), .Z(n746) );
  XOR U863 ( .A(n749), .B(n750), .Z(SUM[144]) );
  XNOR U864 ( .A(B[144]), .B(A[144]), .Z(n750) );
  AND U865 ( .A(n751), .B(n752), .Z(n749) );
  NAND U866 ( .A(B[143]), .B(n753), .Z(n752) );
  NANDN U867 ( .A(A[143]), .B(n754), .Z(n753) );
  NANDN U868 ( .A(n754), .B(A[143]), .Z(n751) );
  XOR U869 ( .A(n754), .B(n755), .Z(SUM[143]) );
  XNOR U870 ( .A(B[143]), .B(A[143]), .Z(n755) );
  AND U871 ( .A(n756), .B(n757), .Z(n754) );
  NAND U872 ( .A(B[142]), .B(n758), .Z(n757) );
  NANDN U873 ( .A(A[142]), .B(n759), .Z(n758) );
  NANDN U874 ( .A(n759), .B(A[142]), .Z(n756) );
  XOR U875 ( .A(n759), .B(n760), .Z(SUM[142]) );
  XNOR U876 ( .A(B[142]), .B(A[142]), .Z(n760) );
  AND U877 ( .A(n761), .B(n762), .Z(n759) );
  NAND U878 ( .A(B[141]), .B(n763), .Z(n762) );
  NANDN U879 ( .A(A[141]), .B(n764), .Z(n763) );
  NANDN U880 ( .A(n764), .B(A[141]), .Z(n761) );
  XOR U881 ( .A(n764), .B(n765), .Z(SUM[141]) );
  XNOR U882 ( .A(B[141]), .B(A[141]), .Z(n765) );
  AND U883 ( .A(n766), .B(n767), .Z(n764) );
  NAND U884 ( .A(B[140]), .B(n768), .Z(n767) );
  NANDN U885 ( .A(A[140]), .B(n769), .Z(n768) );
  NANDN U886 ( .A(n769), .B(A[140]), .Z(n766) );
  XOR U887 ( .A(n769), .B(n770), .Z(SUM[140]) );
  XNOR U888 ( .A(B[140]), .B(A[140]), .Z(n770) );
  AND U889 ( .A(n771), .B(n772), .Z(n769) );
  NAND U890 ( .A(B[139]), .B(n773), .Z(n772) );
  NANDN U891 ( .A(A[139]), .B(n774), .Z(n773) );
  NANDN U892 ( .A(n774), .B(A[139]), .Z(n771) );
  XOR U893 ( .A(n775), .B(n776), .Z(SUM[13]) );
  XNOR U894 ( .A(B[13]), .B(A[13]), .Z(n776) );
  XOR U895 ( .A(n774), .B(n777), .Z(SUM[139]) );
  XNOR U896 ( .A(B[139]), .B(A[139]), .Z(n777) );
  AND U897 ( .A(n778), .B(n779), .Z(n774) );
  NAND U898 ( .A(B[138]), .B(n780), .Z(n779) );
  NANDN U899 ( .A(A[138]), .B(n781), .Z(n780) );
  NANDN U900 ( .A(n781), .B(A[138]), .Z(n778) );
  XOR U901 ( .A(n781), .B(n782), .Z(SUM[138]) );
  XNOR U902 ( .A(B[138]), .B(A[138]), .Z(n782) );
  AND U903 ( .A(n783), .B(n784), .Z(n781) );
  NAND U904 ( .A(B[137]), .B(n785), .Z(n784) );
  NANDN U905 ( .A(A[137]), .B(n786), .Z(n785) );
  NANDN U906 ( .A(n786), .B(A[137]), .Z(n783) );
  XOR U907 ( .A(n786), .B(n787), .Z(SUM[137]) );
  XNOR U908 ( .A(B[137]), .B(A[137]), .Z(n787) );
  AND U909 ( .A(n788), .B(n789), .Z(n786) );
  NAND U910 ( .A(B[136]), .B(n790), .Z(n789) );
  NANDN U911 ( .A(A[136]), .B(n791), .Z(n790) );
  NANDN U912 ( .A(n791), .B(A[136]), .Z(n788) );
  XOR U913 ( .A(n791), .B(n792), .Z(SUM[136]) );
  XNOR U914 ( .A(B[136]), .B(A[136]), .Z(n792) );
  AND U915 ( .A(n793), .B(n794), .Z(n791) );
  NAND U916 ( .A(B[135]), .B(n795), .Z(n794) );
  NANDN U917 ( .A(A[135]), .B(n796), .Z(n795) );
  NANDN U918 ( .A(n796), .B(A[135]), .Z(n793) );
  XOR U919 ( .A(n796), .B(n797), .Z(SUM[135]) );
  XNOR U920 ( .A(B[135]), .B(A[135]), .Z(n797) );
  AND U921 ( .A(n798), .B(n799), .Z(n796) );
  NAND U922 ( .A(B[134]), .B(n800), .Z(n799) );
  NANDN U923 ( .A(A[134]), .B(n801), .Z(n800) );
  NANDN U924 ( .A(n801), .B(A[134]), .Z(n798) );
  XOR U925 ( .A(n801), .B(n802), .Z(SUM[134]) );
  XNOR U926 ( .A(B[134]), .B(A[134]), .Z(n802) );
  AND U927 ( .A(n803), .B(n804), .Z(n801) );
  NAND U928 ( .A(B[133]), .B(n805), .Z(n804) );
  NANDN U929 ( .A(A[133]), .B(n806), .Z(n805) );
  NANDN U930 ( .A(n806), .B(A[133]), .Z(n803) );
  XOR U931 ( .A(n806), .B(n807), .Z(SUM[133]) );
  XNOR U932 ( .A(B[133]), .B(A[133]), .Z(n807) );
  AND U933 ( .A(n808), .B(n809), .Z(n806) );
  NAND U934 ( .A(B[132]), .B(n810), .Z(n809) );
  NANDN U935 ( .A(A[132]), .B(n811), .Z(n810) );
  NANDN U936 ( .A(n811), .B(A[132]), .Z(n808) );
  XOR U937 ( .A(n811), .B(n812), .Z(SUM[132]) );
  XNOR U938 ( .A(B[132]), .B(A[132]), .Z(n812) );
  AND U939 ( .A(n813), .B(n814), .Z(n811) );
  NAND U940 ( .A(B[131]), .B(n815), .Z(n814) );
  NANDN U941 ( .A(A[131]), .B(n816), .Z(n815) );
  NANDN U942 ( .A(n816), .B(A[131]), .Z(n813) );
  XOR U943 ( .A(n816), .B(n817), .Z(SUM[131]) );
  XNOR U944 ( .A(B[131]), .B(A[131]), .Z(n817) );
  AND U945 ( .A(n818), .B(n819), .Z(n816) );
  NAND U946 ( .A(B[130]), .B(n820), .Z(n819) );
  NANDN U947 ( .A(A[130]), .B(n821), .Z(n820) );
  NANDN U948 ( .A(n821), .B(A[130]), .Z(n818) );
  XOR U949 ( .A(n821), .B(n822), .Z(SUM[130]) );
  XNOR U950 ( .A(B[130]), .B(A[130]), .Z(n822) );
  AND U951 ( .A(n823), .B(n824), .Z(n821) );
  NAND U952 ( .A(B[129]), .B(n825), .Z(n824) );
  NANDN U953 ( .A(A[129]), .B(n826), .Z(n825) );
  NANDN U954 ( .A(n826), .B(A[129]), .Z(n823) );
  XOR U955 ( .A(n827), .B(n828), .Z(SUM[12]) );
  XNOR U956 ( .A(B[12]), .B(A[12]), .Z(n828) );
  XOR U957 ( .A(n826), .B(n829), .Z(SUM[129]) );
  XNOR U958 ( .A(B[129]), .B(A[129]), .Z(n829) );
  AND U959 ( .A(n830), .B(n831), .Z(n826) );
  NAND U960 ( .A(B[128]), .B(n832), .Z(n831) );
  NANDN U961 ( .A(A[128]), .B(n833), .Z(n832) );
  NANDN U962 ( .A(n833), .B(A[128]), .Z(n830) );
  XOR U963 ( .A(n833), .B(n834), .Z(SUM[128]) );
  XNOR U964 ( .A(B[128]), .B(A[128]), .Z(n834) );
  AND U965 ( .A(n835), .B(n836), .Z(n833) );
  NAND U966 ( .A(B[127]), .B(n837), .Z(n836) );
  NANDN U967 ( .A(A[127]), .B(n838), .Z(n837) );
  NANDN U968 ( .A(n838), .B(A[127]), .Z(n835) );
  XOR U969 ( .A(n838), .B(n839), .Z(SUM[127]) );
  XNOR U970 ( .A(B[127]), .B(A[127]), .Z(n839) );
  AND U971 ( .A(n840), .B(n841), .Z(n838) );
  NAND U972 ( .A(B[126]), .B(n842), .Z(n841) );
  NANDN U973 ( .A(A[126]), .B(n843), .Z(n842) );
  NANDN U974 ( .A(n843), .B(A[126]), .Z(n840) );
  XOR U975 ( .A(n843), .B(n844), .Z(SUM[126]) );
  XNOR U976 ( .A(B[126]), .B(A[126]), .Z(n844) );
  AND U977 ( .A(n845), .B(n846), .Z(n843) );
  NAND U978 ( .A(B[125]), .B(n847), .Z(n846) );
  NANDN U979 ( .A(A[125]), .B(n848), .Z(n847) );
  NANDN U980 ( .A(n848), .B(A[125]), .Z(n845) );
  XOR U981 ( .A(n848), .B(n849), .Z(SUM[125]) );
  XNOR U982 ( .A(B[125]), .B(A[125]), .Z(n849) );
  AND U983 ( .A(n850), .B(n851), .Z(n848) );
  NAND U984 ( .A(B[124]), .B(n852), .Z(n851) );
  NANDN U985 ( .A(A[124]), .B(n853), .Z(n852) );
  NANDN U986 ( .A(n853), .B(A[124]), .Z(n850) );
  XOR U987 ( .A(n853), .B(n854), .Z(SUM[124]) );
  XNOR U988 ( .A(B[124]), .B(A[124]), .Z(n854) );
  AND U989 ( .A(n855), .B(n856), .Z(n853) );
  NAND U990 ( .A(B[123]), .B(n857), .Z(n856) );
  NANDN U991 ( .A(A[123]), .B(n858), .Z(n857) );
  NANDN U992 ( .A(n858), .B(A[123]), .Z(n855) );
  XOR U993 ( .A(n858), .B(n859), .Z(SUM[123]) );
  XNOR U994 ( .A(B[123]), .B(A[123]), .Z(n859) );
  AND U995 ( .A(n860), .B(n861), .Z(n858) );
  NAND U996 ( .A(B[122]), .B(n862), .Z(n861) );
  NANDN U997 ( .A(A[122]), .B(n863), .Z(n862) );
  NANDN U998 ( .A(n863), .B(A[122]), .Z(n860) );
  XOR U999 ( .A(n863), .B(n864), .Z(SUM[122]) );
  XNOR U1000 ( .A(B[122]), .B(A[122]), .Z(n864) );
  AND U1001 ( .A(n865), .B(n866), .Z(n863) );
  NAND U1002 ( .A(B[121]), .B(n867), .Z(n866) );
  NANDN U1003 ( .A(A[121]), .B(n868), .Z(n867) );
  NANDN U1004 ( .A(n868), .B(A[121]), .Z(n865) );
  XOR U1005 ( .A(n868), .B(n869), .Z(SUM[121]) );
  XNOR U1006 ( .A(B[121]), .B(A[121]), .Z(n869) );
  AND U1007 ( .A(n870), .B(n871), .Z(n868) );
  NAND U1008 ( .A(B[120]), .B(n872), .Z(n871) );
  NANDN U1009 ( .A(A[120]), .B(n873), .Z(n872) );
  NANDN U1010 ( .A(n873), .B(A[120]), .Z(n870) );
  XOR U1011 ( .A(n873), .B(n874), .Z(SUM[120]) );
  XNOR U1012 ( .A(B[120]), .B(A[120]), .Z(n874) );
  AND U1013 ( .A(n875), .B(n876), .Z(n873) );
  NAND U1014 ( .A(B[119]), .B(n877), .Z(n876) );
  NANDN U1015 ( .A(A[119]), .B(n878), .Z(n877) );
  NANDN U1016 ( .A(n878), .B(A[119]), .Z(n875) );
  XOR U1017 ( .A(n879), .B(n880), .Z(SUM[11]) );
  XNOR U1018 ( .A(B[11]), .B(A[11]), .Z(n880) );
  XOR U1019 ( .A(n878), .B(n881), .Z(SUM[119]) );
  XNOR U1020 ( .A(B[119]), .B(A[119]), .Z(n881) );
  AND U1021 ( .A(n882), .B(n883), .Z(n878) );
  NAND U1022 ( .A(B[118]), .B(n884), .Z(n883) );
  NANDN U1023 ( .A(A[118]), .B(n885), .Z(n884) );
  NANDN U1024 ( .A(n885), .B(A[118]), .Z(n882) );
  XOR U1025 ( .A(n885), .B(n886), .Z(SUM[118]) );
  XNOR U1026 ( .A(B[118]), .B(A[118]), .Z(n886) );
  AND U1027 ( .A(n887), .B(n888), .Z(n885) );
  NAND U1028 ( .A(B[117]), .B(n889), .Z(n888) );
  NANDN U1029 ( .A(A[117]), .B(n890), .Z(n889) );
  NANDN U1030 ( .A(n890), .B(A[117]), .Z(n887) );
  XOR U1031 ( .A(n890), .B(n891), .Z(SUM[117]) );
  XNOR U1032 ( .A(B[117]), .B(A[117]), .Z(n891) );
  AND U1033 ( .A(n892), .B(n893), .Z(n890) );
  NAND U1034 ( .A(B[116]), .B(n894), .Z(n893) );
  NANDN U1035 ( .A(A[116]), .B(n895), .Z(n894) );
  NANDN U1036 ( .A(n895), .B(A[116]), .Z(n892) );
  XOR U1037 ( .A(n895), .B(n896), .Z(SUM[116]) );
  XNOR U1038 ( .A(B[116]), .B(A[116]), .Z(n896) );
  AND U1039 ( .A(n897), .B(n898), .Z(n895) );
  NAND U1040 ( .A(B[115]), .B(n899), .Z(n898) );
  NANDN U1041 ( .A(A[115]), .B(n900), .Z(n899) );
  NANDN U1042 ( .A(n900), .B(A[115]), .Z(n897) );
  XOR U1043 ( .A(n900), .B(n901), .Z(SUM[115]) );
  XNOR U1044 ( .A(B[115]), .B(A[115]), .Z(n901) );
  AND U1045 ( .A(n902), .B(n903), .Z(n900) );
  NAND U1046 ( .A(B[114]), .B(n904), .Z(n903) );
  NANDN U1047 ( .A(A[114]), .B(n905), .Z(n904) );
  NANDN U1048 ( .A(n905), .B(A[114]), .Z(n902) );
  XOR U1049 ( .A(n905), .B(n906), .Z(SUM[114]) );
  XNOR U1050 ( .A(B[114]), .B(A[114]), .Z(n906) );
  AND U1051 ( .A(n907), .B(n908), .Z(n905) );
  NAND U1052 ( .A(B[113]), .B(n909), .Z(n908) );
  NANDN U1053 ( .A(A[113]), .B(n910), .Z(n909) );
  NANDN U1054 ( .A(n910), .B(A[113]), .Z(n907) );
  XOR U1055 ( .A(n910), .B(n911), .Z(SUM[113]) );
  XNOR U1056 ( .A(B[113]), .B(A[113]), .Z(n911) );
  AND U1057 ( .A(n912), .B(n913), .Z(n910) );
  NAND U1058 ( .A(B[112]), .B(n914), .Z(n913) );
  NANDN U1059 ( .A(A[112]), .B(n915), .Z(n914) );
  NANDN U1060 ( .A(n915), .B(A[112]), .Z(n912) );
  XOR U1061 ( .A(n915), .B(n916), .Z(SUM[112]) );
  XNOR U1062 ( .A(B[112]), .B(A[112]), .Z(n916) );
  AND U1063 ( .A(n917), .B(n918), .Z(n915) );
  NAND U1064 ( .A(B[111]), .B(n919), .Z(n918) );
  NANDN U1065 ( .A(A[111]), .B(n920), .Z(n919) );
  NANDN U1066 ( .A(n920), .B(A[111]), .Z(n917) );
  XOR U1067 ( .A(n920), .B(n921), .Z(SUM[111]) );
  XNOR U1068 ( .A(B[111]), .B(A[111]), .Z(n921) );
  AND U1069 ( .A(n922), .B(n923), .Z(n920) );
  NAND U1070 ( .A(B[110]), .B(n924), .Z(n923) );
  NANDN U1071 ( .A(A[110]), .B(n925), .Z(n924) );
  NANDN U1072 ( .A(n925), .B(A[110]), .Z(n922) );
  XOR U1073 ( .A(n925), .B(n926), .Z(SUM[110]) );
  XNOR U1074 ( .A(B[110]), .B(A[110]), .Z(n926) );
  AND U1075 ( .A(n927), .B(n928), .Z(n925) );
  NAND U1076 ( .A(B[109]), .B(n929), .Z(n928) );
  NANDN U1077 ( .A(A[109]), .B(n930), .Z(n929) );
  NANDN U1078 ( .A(n930), .B(A[109]), .Z(n927) );
  XOR U1079 ( .A(n931), .B(n932), .Z(SUM[10]) );
  XNOR U1080 ( .A(B[10]), .B(A[10]), .Z(n932) );
  XOR U1081 ( .A(n930), .B(n933), .Z(SUM[109]) );
  XNOR U1082 ( .A(B[109]), .B(A[109]), .Z(n933) );
  AND U1083 ( .A(n934), .B(n935), .Z(n930) );
  NAND U1084 ( .A(B[108]), .B(n936), .Z(n935) );
  NANDN U1085 ( .A(A[108]), .B(n937), .Z(n936) );
  NANDN U1086 ( .A(n937), .B(A[108]), .Z(n934) );
  XOR U1087 ( .A(n937), .B(n938), .Z(SUM[108]) );
  XNOR U1088 ( .A(B[108]), .B(A[108]), .Z(n938) );
  AND U1089 ( .A(n939), .B(n940), .Z(n937) );
  NAND U1090 ( .A(B[107]), .B(n941), .Z(n940) );
  NANDN U1091 ( .A(A[107]), .B(n942), .Z(n941) );
  NANDN U1092 ( .A(n942), .B(A[107]), .Z(n939) );
  XOR U1093 ( .A(n942), .B(n943), .Z(SUM[107]) );
  XNOR U1094 ( .A(B[107]), .B(A[107]), .Z(n943) );
  AND U1095 ( .A(n944), .B(n945), .Z(n942) );
  NAND U1096 ( .A(B[106]), .B(n946), .Z(n945) );
  NANDN U1097 ( .A(A[106]), .B(n947), .Z(n946) );
  NANDN U1098 ( .A(n947), .B(A[106]), .Z(n944) );
  XOR U1099 ( .A(n947), .B(n948), .Z(SUM[106]) );
  XNOR U1100 ( .A(B[106]), .B(A[106]), .Z(n948) );
  AND U1101 ( .A(n949), .B(n950), .Z(n947) );
  NAND U1102 ( .A(B[105]), .B(n951), .Z(n950) );
  NANDN U1103 ( .A(A[105]), .B(n952), .Z(n951) );
  NANDN U1104 ( .A(n952), .B(A[105]), .Z(n949) );
  XOR U1105 ( .A(n952), .B(n953), .Z(SUM[105]) );
  XNOR U1106 ( .A(B[105]), .B(A[105]), .Z(n953) );
  AND U1107 ( .A(n954), .B(n955), .Z(n952) );
  NAND U1108 ( .A(B[104]), .B(n956), .Z(n955) );
  NANDN U1109 ( .A(A[104]), .B(n957), .Z(n956) );
  NANDN U1110 ( .A(n957), .B(A[104]), .Z(n954) );
  XOR U1111 ( .A(n957), .B(n958), .Z(SUM[104]) );
  XNOR U1112 ( .A(B[104]), .B(A[104]), .Z(n958) );
  AND U1113 ( .A(n959), .B(n960), .Z(n957) );
  NAND U1114 ( .A(B[103]), .B(n961), .Z(n960) );
  NANDN U1115 ( .A(A[103]), .B(n962), .Z(n961) );
  NANDN U1116 ( .A(n962), .B(A[103]), .Z(n959) );
  XOR U1117 ( .A(n962), .B(n963), .Z(SUM[103]) );
  XNOR U1118 ( .A(B[103]), .B(A[103]), .Z(n963) );
  AND U1119 ( .A(n964), .B(n965), .Z(n962) );
  NAND U1120 ( .A(B[102]), .B(n966), .Z(n965) );
  NANDN U1121 ( .A(A[102]), .B(n967), .Z(n966) );
  NANDN U1122 ( .A(n967), .B(A[102]), .Z(n964) );
  XOR U1123 ( .A(n967), .B(n968), .Z(SUM[102]) );
  XNOR U1124 ( .A(B[102]), .B(A[102]), .Z(n968) );
  AND U1125 ( .A(n969), .B(n970), .Z(n967) );
  NAND U1126 ( .A(B[101]), .B(n971), .Z(n970) );
  NANDN U1127 ( .A(A[101]), .B(n972), .Z(n971) );
  NANDN U1128 ( .A(n972), .B(A[101]), .Z(n969) );
  XOR U1129 ( .A(n972), .B(n973), .Z(SUM[101]) );
  XNOR U1130 ( .A(B[101]), .B(A[101]), .Z(n973) );
  AND U1131 ( .A(n974), .B(n975), .Z(n972) );
  NAND U1132 ( .A(B[100]), .B(n976), .Z(n975) );
  NANDN U1133 ( .A(A[100]), .B(n977), .Z(n976) );
  NANDN U1134 ( .A(n977), .B(A[100]), .Z(n974) );
  XOR U1135 ( .A(n977), .B(n978), .Z(SUM[100]) );
  XNOR U1136 ( .A(B[100]), .B(A[100]), .Z(n978) );
  AND U1137 ( .A(n979), .B(n980), .Z(n977) );
  NAND U1138 ( .A(B[99]), .B(n981), .Z(n980) );
  OR U1139 ( .A(n3), .B(A[99]), .Z(n981) );
  NAND U1140 ( .A(A[99]), .B(n3), .Z(n979) );
  NAND U1141 ( .A(n982), .B(n983), .Z(n3) );
  NAND U1142 ( .A(B[98]), .B(n984), .Z(n983) );
  NANDN U1143 ( .A(A[98]), .B(n5), .Z(n984) );
  NANDN U1144 ( .A(n5), .B(A[98]), .Z(n982) );
  AND U1145 ( .A(n985), .B(n986), .Z(n5) );
  NAND U1146 ( .A(B[97]), .B(n987), .Z(n986) );
  NANDN U1147 ( .A(A[97]), .B(n7), .Z(n987) );
  NANDN U1148 ( .A(n7), .B(A[97]), .Z(n985) );
  AND U1149 ( .A(n988), .B(n989), .Z(n7) );
  NAND U1150 ( .A(B[96]), .B(n990), .Z(n989) );
  NANDN U1151 ( .A(A[96]), .B(n9), .Z(n990) );
  NANDN U1152 ( .A(n9), .B(A[96]), .Z(n988) );
  AND U1153 ( .A(n991), .B(n992), .Z(n9) );
  NAND U1154 ( .A(B[95]), .B(n993), .Z(n992) );
  NANDN U1155 ( .A(A[95]), .B(n11), .Z(n993) );
  NANDN U1156 ( .A(n11), .B(A[95]), .Z(n991) );
  AND U1157 ( .A(n994), .B(n995), .Z(n11) );
  NAND U1158 ( .A(B[94]), .B(n996), .Z(n995) );
  NANDN U1159 ( .A(A[94]), .B(n13), .Z(n996) );
  NANDN U1160 ( .A(n13), .B(A[94]), .Z(n994) );
  AND U1161 ( .A(n997), .B(n998), .Z(n13) );
  NAND U1162 ( .A(B[93]), .B(n999), .Z(n998) );
  NANDN U1163 ( .A(A[93]), .B(n15), .Z(n999) );
  NANDN U1164 ( .A(n15), .B(A[93]), .Z(n997) );
  AND U1165 ( .A(n1000), .B(n1001), .Z(n15) );
  NAND U1166 ( .A(B[92]), .B(n1002), .Z(n1001) );
  NANDN U1167 ( .A(A[92]), .B(n17), .Z(n1002) );
  NANDN U1168 ( .A(n17), .B(A[92]), .Z(n1000) );
  AND U1169 ( .A(n1003), .B(n1004), .Z(n17) );
  NAND U1170 ( .A(B[91]), .B(n1005), .Z(n1004) );
  NANDN U1171 ( .A(A[91]), .B(n19), .Z(n1005) );
  NANDN U1172 ( .A(n19), .B(A[91]), .Z(n1003) );
  AND U1173 ( .A(n1006), .B(n1007), .Z(n19) );
  NAND U1174 ( .A(B[90]), .B(n1008), .Z(n1007) );
  NANDN U1175 ( .A(A[90]), .B(n21), .Z(n1008) );
  NANDN U1176 ( .A(n21), .B(A[90]), .Z(n1006) );
  AND U1177 ( .A(n1009), .B(n1010), .Z(n21) );
  NAND U1178 ( .A(B[89]), .B(n1011), .Z(n1010) );
  NANDN U1179 ( .A(A[89]), .B(n25), .Z(n1011) );
  NANDN U1180 ( .A(n25), .B(A[89]), .Z(n1009) );
  AND U1181 ( .A(n1012), .B(n1013), .Z(n25) );
  NAND U1182 ( .A(B[88]), .B(n1014), .Z(n1013) );
  NANDN U1183 ( .A(A[88]), .B(n27), .Z(n1014) );
  NANDN U1184 ( .A(n27), .B(A[88]), .Z(n1012) );
  AND U1185 ( .A(n1015), .B(n1016), .Z(n27) );
  NAND U1186 ( .A(B[87]), .B(n1017), .Z(n1016) );
  NANDN U1187 ( .A(A[87]), .B(n29), .Z(n1017) );
  NANDN U1188 ( .A(n29), .B(A[87]), .Z(n1015) );
  AND U1189 ( .A(n1018), .B(n1019), .Z(n29) );
  NAND U1190 ( .A(B[86]), .B(n1020), .Z(n1019) );
  NANDN U1191 ( .A(A[86]), .B(n31), .Z(n1020) );
  NANDN U1192 ( .A(n31), .B(A[86]), .Z(n1018) );
  AND U1193 ( .A(n1021), .B(n1022), .Z(n31) );
  NAND U1194 ( .A(B[85]), .B(n1023), .Z(n1022) );
  NANDN U1195 ( .A(A[85]), .B(n33), .Z(n1023) );
  NANDN U1196 ( .A(n33), .B(A[85]), .Z(n1021) );
  AND U1197 ( .A(n1024), .B(n1025), .Z(n33) );
  NAND U1198 ( .A(B[84]), .B(n1026), .Z(n1025) );
  NANDN U1199 ( .A(A[84]), .B(n35), .Z(n1026) );
  NANDN U1200 ( .A(n35), .B(A[84]), .Z(n1024) );
  AND U1201 ( .A(n1027), .B(n1028), .Z(n35) );
  NAND U1202 ( .A(B[83]), .B(n1029), .Z(n1028) );
  NANDN U1203 ( .A(A[83]), .B(n37), .Z(n1029) );
  NANDN U1204 ( .A(n37), .B(A[83]), .Z(n1027) );
  AND U1205 ( .A(n1030), .B(n1031), .Z(n37) );
  NAND U1206 ( .A(B[82]), .B(n1032), .Z(n1031) );
  NANDN U1207 ( .A(A[82]), .B(n39), .Z(n1032) );
  NANDN U1208 ( .A(n39), .B(A[82]), .Z(n1030) );
  AND U1209 ( .A(n1033), .B(n1034), .Z(n39) );
  NAND U1210 ( .A(B[81]), .B(n1035), .Z(n1034) );
  NANDN U1211 ( .A(A[81]), .B(n41), .Z(n1035) );
  NANDN U1212 ( .A(n41), .B(A[81]), .Z(n1033) );
  AND U1213 ( .A(n1036), .B(n1037), .Z(n41) );
  NAND U1214 ( .A(B[80]), .B(n1038), .Z(n1037) );
  NANDN U1215 ( .A(A[80]), .B(n43), .Z(n1038) );
  NANDN U1216 ( .A(n43), .B(A[80]), .Z(n1036) );
  AND U1217 ( .A(n1039), .B(n1040), .Z(n43) );
  NAND U1218 ( .A(B[79]), .B(n1041), .Z(n1040) );
  NANDN U1219 ( .A(A[79]), .B(n47), .Z(n1041) );
  NANDN U1220 ( .A(n47), .B(A[79]), .Z(n1039) );
  AND U1221 ( .A(n1042), .B(n1043), .Z(n47) );
  NAND U1222 ( .A(B[78]), .B(n1044), .Z(n1043) );
  NANDN U1223 ( .A(A[78]), .B(n49), .Z(n1044) );
  NANDN U1224 ( .A(n49), .B(A[78]), .Z(n1042) );
  AND U1225 ( .A(n1045), .B(n1046), .Z(n49) );
  NAND U1226 ( .A(B[77]), .B(n1047), .Z(n1046) );
  NANDN U1227 ( .A(A[77]), .B(n51), .Z(n1047) );
  NANDN U1228 ( .A(n51), .B(A[77]), .Z(n1045) );
  AND U1229 ( .A(n1048), .B(n1049), .Z(n51) );
  NAND U1230 ( .A(B[76]), .B(n1050), .Z(n1049) );
  NANDN U1231 ( .A(A[76]), .B(n53), .Z(n1050) );
  NANDN U1232 ( .A(n53), .B(A[76]), .Z(n1048) );
  AND U1233 ( .A(n1051), .B(n1052), .Z(n53) );
  NAND U1234 ( .A(B[75]), .B(n1053), .Z(n1052) );
  NANDN U1235 ( .A(A[75]), .B(n55), .Z(n1053) );
  NANDN U1236 ( .A(n55), .B(A[75]), .Z(n1051) );
  AND U1237 ( .A(n1054), .B(n1055), .Z(n55) );
  NAND U1238 ( .A(B[74]), .B(n1056), .Z(n1055) );
  NANDN U1239 ( .A(A[74]), .B(n57), .Z(n1056) );
  NANDN U1240 ( .A(n57), .B(A[74]), .Z(n1054) );
  AND U1241 ( .A(n1057), .B(n1058), .Z(n57) );
  NAND U1242 ( .A(B[73]), .B(n1059), .Z(n1058) );
  NANDN U1243 ( .A(A[73]), .B(n59), .Z(n1059) );
  NANDN U1244 ( .A(n59), .B(A[73]), .Z(n1057) );
  AND U1245 ( .A(n1060), .B(n1061), .Z(n59) );
  NAND U1246 ( .A(B[72]), .B(n1062), .Z(n1061) );
  NANDN U1247 ( .A(A[72]), .B(n61), .Z(n1062) );
  NANDN U1248 ( .A(n61), .B(A[72]), .Z(n1060) );
  AND U1249 ( .A(n1063), .B(n1064), .Z(n61) );
  NAND U1250 ( .A(B[71]), .B(n1065), .Z(n1064) );
  NANDN U1251 ( .A(A[71]), .B(n63), .Z(n1065) );
  NANDN U1252 ( .A(n63), .B(A[71]), .Z(n1063) );
  AND U1253 ( .A(n1066), .B(n1067), .Z(n63) );
  NAND U1254 ( .A(B[70]), .B(n1068), .Z(n1067) );
  NANDN U1255 ( .A(A[70]), .B(n65), .Z(n1068) );
  NANDN U1256 ( .A(n65), .B(A[70]), .Z(n1066) );
  AND U1257 ( .A(n1069), .B(n1070), .Z(n65) );
  NAND U1258 ( .A(B[69]), .B(n1071), .Z(n1070) );
  NANDN U1259 ( .A(A[69]), .B(n69), .Z(n1071) );
  NANDN U1260 ( .A(n69), .B(A[69]), .Z(n1069) );
  AND U1261 ( .A(n1072), .B(n1073), .Z(n69) );
  NAND U1262 ( .A(B[68]), .B(n1074), .Z(n1073) );
  NANDN U1263 ( .A(A[68]), .B(n71), .Z(n1074) );
  NANDN U1264 ( .A(n71), .B(A[68]), .Z(n1072) );
  AND U1265 ( .A(n1075), .B(n1076), .Z(n71) );
  NAND U1266 ( .A(B[67]), .B(n1077), .Z(n1076) );
  NANDN U1267 ( .A(A[67]), .B(n73), .Z(n1077) );
  NANDN U1268 ( .A(n73), .B(A[67]), .Z(n1075) );
  AND U1269 ( .A(n1078), .B(n1079), .Z(n73) );
  NAND U1270 ( .A(B[66]), .B(n1080), .Z(n1079) );
  NANDN U1271 ( .A(A[66]), .B(n75), .Z(n1080) );
  NANDN U1272 ( .A(n75), .B(A[66]), .Z(n1078) );
  AND U1273 ( .A(n1081), .B(n1082), .Z(n75) );
  NAND U1274 ( .A(B[65]), .B(n1083), .Z(n1082) );
  NANDN U1275 ( .A(A[65]), .B(n77), .Z(n1083) );
  NANDN U1276 ( .A(n77), .B(A[65]), .Z(n1081) );
  AND U1277 ( .A(n1084), .B(n1085), .Z(n77) );
  NAND U1278 ( .A(B[64]), .B(n1086), .Z(n1085) );
  NANDN U1279 ( .A(A[64]), .B(n79), .Z(n1086) );
  NANDN U1280 ( .A(n79), .B(A[64]), .Z(n1084) );
  AND U1281 ( .A(n1087), .B(n1088), .Z(n79) );
  NAND U1282 ( .A(B[63]), .B(n1089), .Z(n1088) );
  NANDN U1283 ( .A(A[63]), .B(n81), .Z(n1089) );
  NANDN U1284 ( .A(n81), .B(A[63]), .Z(n1087) );
  AND U1285 ( .A(n1090), .B(n1091), .Z(n81) );
  NAND U1286 ( .A(B[62]), .B(n1092), .Z(n1091) );
  NANDN U1287 ( .A(A[62]), .B(n83), .Z(n1092) );
  NANDN U1288 ( .A(n83), .B(A[62]), .Z(n1090) );
  AND U1289 ( .A(n1093), .B(n1094), .Z(n83) );
  NAND U1290 ( .A(B[61]), .B(n1095), .Z(n1094) );
  NANDN U1291 ( .A(A[61]), .B(n85), .Z(n1095) );
  NANDN U1292 ( .A(n85), .B(A[61]), .Z(n1093) );
  AND U1293 ( .A(n1096), .B(n1097), .Z(n85) );
  NAND U1294 ( .A(B[60]), .B(n1098), .Z(n1097) );
  NANDN U1295 ( .A(A[60]), .B(n87), .Z(n1098) );
  NANDN U1296 ( .A(n87), .B(A[60]), .Z(n1096) );
  AND U1297 ( .A(n1099), .B(n1100), .Z(n87) );
  NAND U1298 ( .A(B[59]), .B(n1101), .Z(n1100) );
  NANDN U1299 ( .A(A[59]), .B(n91), .Z(n1101) );
  NANDN U1300 ( .A(n91), .B(A[59]), .Z(n1099) );
  AND U1301 ( .A(n1102), .B(n1103), .Z(n91) );
  NAND U1302 ( .A(B[58]), .B(n1104), .Z(n1103) );
  NANDN U1303 ( .A(A[58]), .B(n93), .Z(n1104) );
  NANDN U1304 ( .A(n93), .B(A[58]), .Z(n1102) );
  AND U1305 ( .A(n1105), .B(n1106), .Z(n93) );
  NAND U1306 ( .A(B[57]), .B(n1107), .Z(n1106) );
  NANDN U1307 ( .A(A[57]), .B(n95), .Z(n1107) );
  NANDN U1308 ( .A(n95), .B(A[57]), .Z(n1105) );
  AND U1309 ( .A(n1108), .B(n1109), .Z(n95) );
  NAND U1310 ( .A(B[56]), .B(n1110), .Z(n1109) );
  NANDN U1311 ( .A(A[56]), .B(n97), .Z(n1110) );
  NANDN U1312 ( .A(n97), .B(A[56]), .Z(n1108) );
  AND U1313 ( .A(n1111), .B(n1112), .Z(n97) );
  NAND U1314 ( .A(B[55]), .B(n1113), .Z(n1112) );
  NANDN U1315 ( .A(A[55]), .B(n99), .Z(n1113) );
  NANDN U1316 ( .A(n99), .B(A[55]), .Z(n1111) );
  AND U1317 ( .A(n1114), .B(n1115), .Z(n99) );
  NAND U1318 ( .A(B[54]), .B(n1116), .Z(n1115) );
  NANDN U1319 ( .A(A[54]), .B(n101), .Z(n1116) );
  NANDN U1320 ( .A(n101), .B(A[54]), .Z(n1114) );
  AND U1321 ( .A(n1117), .B(n1118), .Z(n101) );
  NAND U1322 ( .A(B[53]), .B(n1119), .Z(n1118) );
  NANDN U1323 ( .A(A[53]), .B(n103), .Z(n1119) );
  NANDN U1324 ( .A(n103), .B(A[53]), .Z(n1117) );
  AND U1325 ( .A(n1120), .B(n1121), .Z(n103) );
  NAND U1326 ( .A(B[52]), .B(n1122), .Z(n1121) );
  NANDN U1327 ( .A(A[52]), .B(n105), .Z(n1122) );
  NANDN U1328 ( .A(n105), .B(A[52]), .Z(n1120) );
  AND U1329 ( .A(n1123), .B(n1124), .Z(n105) );
  NAND U1330 ( .A(B[51]), .B(n1125), .Z(n1124) );
  NANDN U1331 ( .A(A[51]), .B(n107), .Z(n1125) );
  NANDN U1332 ( .A(n107), .B(A[51]), .Z(n1123) );
  AND U1333 ( .A(n1126), .B(n1127), .Z(n107) );
  NAND U1334 ( .A(B[50]), .B(n1128), .Z(n1127) );
  NANDN U1335 ( .A(A[50]), .B(n109), .Z(n1128) );
  NANDN U1336 ( .A(n109), .B(A[50]), .Z(n1126) );
  AND U1337 ( .A(n1129), .B(n1130), .Z(n109) );
  NAND U1338 ( .A(B[49]), .B(n1131), .Z(n1130) );
  NANDN U1339 ( .A(A[49]), .B(n113), .Z(n1131) );
  NANDN U1340 ( .A(n113), .B(A[49]), .Z(n1129) );
  AND U1341 ( .A(n1132), .B(n1133), .Z(n113) );
  NAND U1342 ( .A(B[48]), .B(n1134), .Z(n1133) );
  NANDN U1343 ( .A(A[48]), .B(n115), .Z(n1134) );
  NANDN U1344 ( .A(n115), .B(A[48]), .Z(n1132) );
  AND U1345 ( .A(n1135), .B(n1136), .Z(n115) );
  NAND U1346 ( .A(B[47]), .B(n1137), .Z(n1136) );
  NANDN U1347 ( .A(A[47]), .B(n117), .Z(n1137) );
  NANDN U1348 ( .A(n117), .B(A[47]), .Z(n1135) );
  AND U1349 ( .A(n1138), .B(n1139), .Z(n117) );
  NAND U1350 ( .A(B[46]), .B(n1140), .Z(n1139) );
  NANDN U1351 ( .A(A[46]), .B(n119), .Z(n1140) );
  NANDN U1352 ( .A(n119), .B(A[46]), .Z(n1138) );
  AND U1353 ( .A(n1141), .B(n1142), .Z(n119) );
  NAND U1354 ( .A(B[45]), .B(n1143), .Z(n1142) );
  NANDN U1355 ( .A(A[45]), .B(n121), .Z(n1143) );
  NANDN U1356 ( .A(n121), .B(A[45]), .Z(n1141) );
  AND U1357 ( .A(n1144), .B(n1145), .Z(n121) );
  NAND U1358 ( .A(B[44]), .B(n1146), .Z(n1145) );
  NANDN U1359 ( .A(A[44]), .B(n123), .Z(n1146) );
  NANDN U1360 ( .A(n123), .B(A[44]), .Z(n1144) );
  AND U1361 ( .A(n1147), .B(n1148), .Z(n123) );
  NAND U1362 ( .A(B[43]), .B(n1149), .Z(n1148) );
  NANDN U1363 ( .A(A[43]), .B(n125), .Z(n1149) );
  NANDN U1364 ( .A(n125), .B(A[43]), .Z(n1147) );
  AND U1365 ( .A(n1150), .B(n1151), .Z(n125) );
  NAND U1366 ( .A(B[42]), .B(n1152), .Z(n1151) );
  NANDN U1367 ( .A(A[42]), .B(n127), .Z(n1152) );
  NANDN U1368 ( .A(n127), .B(A[42]), .Z(n1150) );
  AND U1369 ( .A(n1153), .B(n1154), .Z(n127) );
  NAND U1370 ( .A(B[41]), .B(n1155), .Z(n1154) );
  NANDN U1371 ( .A(A[41]), .B(n129), .Z(n1155) );
  NANDN U1372 ( .A(n129), .B(A[41]), .Z(n1153) );
  AND U1373 ( .A(n1156), .B(n1157), .Z(n129) );
  NAND U1374 ( .A(B[40]), .B(n1158), .Z(n1157) );
  NANDN U1375 ( .A(A[40]), .B(n131), .Z(n1158) );
  NANDN U1376 ( .A(n131), .B(A[40]), .Z(n1156) );
  AND U1377 ( .A(n1159), .B(n1160), .Z(n131) );
  NAND U1378 ( .A(B[39]), .B(n1161), .Z(n1160) );
  NANDN U1379 ( .A(A[39]), .B(n135), .Z(n1161) );
  NANDN U1380 ( .A(n135), .B(A[39]), .Z(n1159) );
  AND U1381 ( .A(n1162), .B(n1163), .Z(n135) );
  NAND U1382 ( .A(B[38]), .B(n1164), .Z(n1163) );
  NANDN U1383 ( .A(A[38]), .B(n137), .Z(n1164) );
  NANDN U1384 ( .A(n137), .B(A[38]), .Z(n1162) );
  AND U1385 ( .A(n1165), .B(n1166), .Z(n137) );
  NAND U1386 ( .A(B[37]), .B(n1167), .Z(n1166) );
  NANDN U1387 ( .A(A[37]), .B(n139), .Z(n1167) );
  NANDN U1388 ( .A(n139), .B(A[37]), .Z(n1165) );
  AND U1389 ( .A(n1168), .B(n1169), .Z(n139) );
  NAND U1390 ( .A(B[36]), .B(n1170), .Z(n1169) );
  NANDN U1391 ( .A(A[36]), .B(n141), .Z(n1170) );
  NANDN U1392 ( .A(n141), .B(A[36]), .Z(n1168) );
  AND U1393 ( .A(n1171), .B(n1172), .Z(n141) );
  NAND U1394 ( .A(B[35]), .B(n1173), .Z(n1172) );
  NANDN U1395 ( .A(A[35]), .B(n143), .Z(n1173) );
  NANDN U1396 ( .A(n143), .B(A[35]), .Z(n1171) );
  AND U1397 ( .A(n1174), .B(n1175), .Z(n143) );
  NAND U1398 ( .A(B[34]), .B(n1176), .Z(n1175) );
  NANDN U1399 ( .A(A[34]), .B(n145), .Z(n1176) );
  NANDN U1400 ( .A(n145), .B(A[34]), .Z(n1174) );
  AND U1401 ( .A(n1177), .B(n1178), .Z(n145) );
  NAND U1402 ( .A(B[33]), .B(n1179), .Z(n1178) );
  NANDN U1403 ( .A(A[33]), .B(n147), .Z(n1179) );
  NANDN U1404 ( .A(n147), .B(A[33]), .Z(n1177) );
  AND U1405 ( .A(n1180), .B(n1181), .Z(n147) );
  NAND U1406 ( .A(B[32]), .B(n1182), .Z(n1181) );
  NANDN U1407 ( .A(A[32]), .B(n149), .Z(n1182) );
  NANDN U1408 ( .A(n149), .B(A[32]), .Z(n1180) );
  AND U1409 ( .A(n1183), .B(n1184), .Z(n149) );
  NAND U1410 ( .A(B[31]), .B(n1185), .Z(n1184) );
  NANDN U1411 ( .A(A[31]), .B(n151), .Z(n1185) );
  NANDN U1412 ( .A(n151), .B(A[31]), .Z(n1183) );
  AND U1413 ( .A(n1186), .B(n1187), .Z(n151) );
  NAND U1414 ( .A(B[30]), .B(n1188), .Z(n1187) );
  NANDN U1415 ( .A(A[30]), .B(n153), .Z(n1188) );
  NANDN U1416 ( .A(n153), .B(A[30]), .Z(n1186) );
  AND U1417 ( .A(n1189), .B(n1190), .Z(n153) );
  NAND U1418 ( .A(B[29]), .B(n1191), .Z(n1190) );
  NANDN U1419 ( .A(A[29]), .B(n157), .Z(n1191) );
  NANDN U1420 ( .A(n157), .B(A[29]), .Z(n1189) );
  AND U1421 ( .A(n1192), .B(n1193), .Z(n157) );
  NAND U1422 ( .A(B[28]), .B(n1194), .Z(n1193) );
  NANDN U1423 ( .A(A[28]), .B(n159), .Z(n1194) );
  NANDN U1424 ( .A(n159), .B(A[28]), .Z(n1192) );
  AND U1425 ( .A(n1195), .B(n1196), .Z(n159) );
  NAND U1426 ( .A(B[27]), .B(n1197), .Z(n1196) );
  NANDN U1427 ( .A(A[27]), .B(n161), .Z(n1197) );
  NANDN U1428 ( .A(n161), .B(A[27]), .Z(n1195) );
  AND U1429 ( .A(n1198), .B(n1199), .Z(n161) );
  NAND U1430 ( .A(B[26]), .B(n1200), .Z(n1199) );
  NANDN U1431 ( .A(A[26]), .B(n163), .Z(n1200) );
  NANDN U1432 ( .A(n163), .B(A[26]), .Z(n1198) );
  AND U1433 ( .A(n1201), .B(n1202), .Z(n163) );
  NAND U1434 ( .A(B[25]), .B(n1203), .Z(n1202) );
  NANDN U1435 ( .A(A[25]), .B(n165), .Z(n1203) );
  NANDN U1436 ( .A(n165), .B(A[25]), .Z(n1201) );
  AND U1437 ( .A(n1204), .B(n1205), .Z(n165) );
  NAND U1438 ( .A(B[24]), .B(n1206), .Z(n1205) );
  NANDN U1439 ( .A(A[24]), .B(n203), .Z(n1206) );
  NANDN U1440 ( .A(n203), .B(A[24]), .Z(n1204) );
  AND U1441 ( .A(n1207), .B(n1208), .Z(n203) );
  NAND U1442 ( .A(B[23]), .B(n1209), .Z(n1208) );
  NANDN U1443 ( .A(A[23]), .B(n255), .Z(n1209) );
  NANDN U1444 ( .A(n255), .B(A[23]), .Z(n1207) );
  AND U1445 ( .A(n1210), .B(n1211), .Z(n255) );
  NAND U1446 ( .A(B[22]), .B(n1212), .Z(n1211) );
  NANDN U1447 ( .A(A[22]), .B(n307), .Z(n1212) );
  NANDN U1448 ( .A(n307), .B(A[22]), .Z(n1210) );
  AND U1449 ( .A(n1213), .B(n1214), .Z(n307) );
  NAND U1450 ( .A(B[21]), .B(n1215), .Z(n1214) );
  NANDN U1451 ( .A(A[21]), .B(n359), .Z(n1215) );
  NANDN U1452 ( .A(n359), .B(A[21]), .Z(n1213) );
  AND U1453 ( .A(n1216), .B(n1217), .Z(n359) );
  NAND U1454 ( .A(B[20]), .B(n1218), .Z(n1217) );
  NANDN U1455 ( .A(A[20]), .B(n411), .Z(n1218) );
  NANDN U1456 ( .A(n411), .B(A[20]), .Z(n1216) );
  AND U1457 ( .A(n1219), .B(n1220), .Z(n411) );
  NAND U1458 ( .A(B[19]), .B(n1221), .Z(n1220) );
  NANDN U1459 ( .A(A[19]), .B(n463), .Z(n1221) );
  NANDN U1460 ( .A(n463), .B(A[19]), .Z(n1219) );
  AND U1461 ( .A(n1222), .B(n1223), .Z(n463) );
  NAND U1462 ( .A(B[18]), .B(n1224), .Z(n1223) );
  NANDN U1463 ( .A(A[18]), .B(n515), .Z(n1224) );
  NANDN U1464 ( .A(n515), .B(A[18]), .Z(n1222) );
  AND U1465 ( .A(n1225), .B(n1226), .Z(n515) );
  NAND U1466 ( .A(B[17]), .B(n1227), .Z(n1226) );
  NANDN U1467 ( .A(A[17]), .B(n567), .Z(n1227) );
  NANDN U1468 ( .A(n567), .B(A[17]), .Z(n1225) );
  AND U1469 ( .A(n1228), .B(n1229), .Z(n567) );
  NAND U1470 ( .A(B[16]), .B(n1230), .Z(n1229) );
  NANDN U1471 ( .A(A[16]), .B(n619), .Z(n1230) );
  NANDN U1472 ( .A(n619), .B(A[16]), .Z(n1228) );
  AND U1473 ( .A(n1231), .B(n1232), .Z(n619) );
  NAND U1474 ( .A(B[15]), .B(n1233), .Z(n1232) );
  NANDN U1475 ( .A(A[15]), .B(n671), .Z(n1233) );
  NANDN U1476 ( .A(n671), .B(A[15]), .Z(n1231) );
  AND U1477 ( .A(n1234), .B(n1235), .Z(n671) );
  NAND U1478 ( .A(B[14]), .B(n1236), .Z(n1235) );
  NANDN U1479 ( .A(A[14]), .B(n723), .Z(n1236) );
  NANDN U1480 ( .A(n723), .B(A[14]), .Z(n1234) );
  AND U1481 ( .A(n1237), .B(n1238), .Z(n723) );
  NAND U1482 ( .A(B[13]), .B(n1239), .Z(n1238) );
  NANDN U1483 ( .A(A[13]), .B(n775), .Z(n1239) );
  NANDN U1484 ( .A(n775), .B(A[13]), .Z(n1237) );
  AND U1485 ( .A(n1240), .B(n1241), .Z(n775) );
  NAND U1486 ( .A(B[12]), .B(n1242), .Z(n1241) );
  NANDN U1487 ( .A(A[12]), .B(n827), .Z(n1242) );
  NANDN U1488 ( .A(n827), .B(A[12]), .Z(n1240) );
  AND U1489 ( .A(n1243), .B(n1244), .Z(n827) );
  NAND U1490 ( .A(B[11]), .B(n1245), .Z(n1244) );
  NANDN U1491 ( .A(A[11]), .B(n879), .Z(n1245) );
  NANDN U1492 ( .A(n879), .B(A[11]), .Z(n1243) );
  AND U1493 ( .A(n1246), .B(n1247), .Z(n879) );
  NAND U1494 ( .A(B[10]), .B(n1248), .Z(n1247) );
  NANDN U1495 ( .A(A[10]), .B(n931), .Z(n1248) );
  NANDN U1496 ( .A(n931), .B(A[10]), .Z(n1246) );
  AND U1497 ( .A(n1249), .B(n1250), .Z(n931) );
  NAND U1498 ( .A(B[9]), .B(n1251), .Z(n1250) );
  OR U1499 ( .A(n1), .B(A[9]), .Z(n1251) );
  NAND U1500 ( .A(A[9]), .B(n1), .Z(n1249) );
  NAND U1501 ( .A(n1252), .B(n1253), .Z(n1) );
  NAND U1502 ( .A(B[8]), .B(n1254), .Z(n1253) );
  NANDN U1503 ( .A(A[8]), .B(n23), .Z(n1254) );
  NANDN U1504 ( .A(n23), .B(A[8]), .Z(n1252) );
  AND U1505 ( .A(n1255), .B(n1256), .Z(n23) );
  NAND U1506 ( .A(B[7]), .B(n1257), .Z(n1256) );
  NANDN U1507 ( .A(A[7]), .B(n45), .Z(n1257) );
  NANDN U1508 ( .A(n45), .B(A[7]), .Z(n1255) );
  AND U1509 ( .A(n1258), .B(n1259), .Z(n45) );
  NAND U1510 ( .A(B[6]), .B(n1260), .Z(n1259) );
  NANDN U1511 ( .A(A[6]), .B(n67), .Z(n1260) );
  NANDN U1512 ( .A(n67), .B(A[6]), .Z(n1258) );
  AND U1513 ( .A(n1261), .B(n1262), .Z(n67) );
  NAND U1514 ( .A(B[5]), .B(n1263), .Z(n1262) );
  NANDN U1515 ( .A(A[5]), .B(n89), .Z(n1263) );
  NANDN U1516 ( .A(n89), .B(A[5]), .Z(n1261) );
  AND U1517 ( .A(n1264), .B(n1265), .Z(n89) );
  NAND U1518 ( .A(B[4]), .B(n1266), .Z(n1265) );
  NANDN U1519 ( .A(A[4]), .B(n111), .Z(n1266) );
  NANDN U1520 ( .A(n111), .B(A[4]), .Z(n1264) );
  AND U1521 ( .A(n1267), .B(n1268), .Z(n111) );
  NAND U1522 ( .A(B[3]), .B(n1269), .Z(n1268) );
  NANDN U1523 ( .A(A[3]), .B(n133), .Z(n1269) );
  NANDN U1524 ( .A(n133), .B(A[3]), .Z(n1267) );
  AND U1525 ( .A(n1270), .B(n1271), .Z(n133) );
  NAND U1526 ( .A(B[2]), .B(n1272), .Z(n1271) );
  OR U1527 ( .A(n155), .B(A[2]), .Z(n1272) );
  NAND U1528 ( .A(A[2]), .B(n155), .Z(n1270) );
  AND U1529 ( .A(B[1]), .B(A[1]), .Z(n155) );
endmodule


module modmult_step_N256_2 ( xregN_1, y, n, zin, zout );
  input [255:0] y;
  input [255:0] n;
  input [257:0] zin;
  output [257:0] zout;
  input xregN_1;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123,
         N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200,
         N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211,
         N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222,
         N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233,
         N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244,
         N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255,
         N256, N257, N258, N259, N260, N261, N262, N264, N265, N266, N267,
         N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278,
         N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289,
         N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300,
         N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311,
         N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322,
         N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333,
         N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344,
         N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366,
         N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377,
         N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410,
         N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421,
         N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432,
         N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443,
         N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454,
         N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465,
         N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476,
         N477, N478, N479, N480, N481, N482, N483, N484, N485, N486, N487,
         N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, N498,
         N499, N500, N501, N502, N503, N504, N505, N506, N507, N508, N509,
         N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, N520,
         N521, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771,
         N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760,
         N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749,
         N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738,
         N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727,
         N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716,
         N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705,
         N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694,
         N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683,
         N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672,
         N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661,
         N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650,
         N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639,
         N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628,
         N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617,
         N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606,
         N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595,
         N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584,
         N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573,
         N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562,
         N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551,
         N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540,
         N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529,
         N528, N527, N526, N525, N522, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039;
  wire   [257:0] z2;
  wire   [257:0] z3;
  wire   SYNOPSYS_UNCONNECTED__0;

  modmult_step_N256_2_DW01_sub_0 sub_129_aco ( .A(z3), .B({1'b0, 1'b0, N780, 
        N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, 
        N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, 
        N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, 
        N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, 
        N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, 
        N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, 
        N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, 
        N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, 
        N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, 
        N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, 
        N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, 
        N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, 
        N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, 
        N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, 
        N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, 
        N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, 
        N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, 
        N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, 
        N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, 
        N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, 
        N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, 
        N527, N526, N525}), .CI(1'b0), .DIFF(zout) );
  modmult_step_N256_2_DW02_mult_0 mult_sub_129_aco ( .A(n), .B(N522), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__0, N780, N779, N778, N777, N776, N775, N774, 
        N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, 
        N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, 
        N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, 
        N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, 
        N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, 
        N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, 
        N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, 
        N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, 
        N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, 
        N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, 
        N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, 
        N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, 
        N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, 
        N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, 
        N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, 
        N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, 
        N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, 
        N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, 
        N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, 
        N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, 
        N533, N532, N531, N530, N529, N528, N527, N526, N525}) );
  modmult_step_N256_2_DW01_cmp2_0 gte_128 ( .A({1'b0, 1'b0, n}), .B(z3), .LEQ(
        1'b1), .TC(1'b0), .LT_LE(N522) );
  modmult_step_N256_2_DW01_sub_1 sub_124 ( .A(z2), .B({1'b0, 1'b0, n}), .CI(
        1'b0), .DIFF({N521, N520, N519, N518, N517, N516, N515, N514, N513, 
        N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, 
        N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, 
        N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, 
        N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, 
        N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, 
        N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, 
        N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, 
        N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, 
        N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, 
        N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, 
        N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, 
        N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, 
        N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, 
        N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, 
        N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, 
        N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, 
        N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, 
        N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, 
        N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, 
        N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, 
        N272, N271, N270, N269, N268, N267, N266, N265, N264}) );
  modmult_step_N256_2_DW01_cmp2_1 gt_123 ( .A({1'b0, 1'b0, n}), .B(z2), .LEQ(
        1'b0), .TC(1'b0), .LT_LE(N262) );
  modmult_step_N256_2_DW01_add_0 add_119 ( .A({zin[256:0], 1'b0}), .B({1'b0, 
        1'b0, y}), .CI(1'b0), .SUM({N261, N260, N259, N258, N257, N256, N255, 
        N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, 
        N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, 
        N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, 
        N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, 
        N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, 
        N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, 
        N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, 
        N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, 
        N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, 
        N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, 
        N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, 
        N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, 
        N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, 
        N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, 
        N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4}) );
  NAND U5 ( .A(n1), .B(n2), .Z(z3[9]) );
  NANDN U6 ( .A(N262), .B(z2[9]), .Z(n2) );
  NANDN U7 ( .A(n3), .B(N273), .Z(n1) );
  NAND U8 ( .A(n4), .B(n5), .Z(z3[99]) );
  NANDN U9 ( .A(N262), .B(z2[99]), .Z(n5) );
  NANDN U10 ( .A(n3), .B(N363), .Z(n4) );
  NAND U11 ( .A(n6), .B(n7), .Z(z3[98]) );
  NANDN U17 ( .A(N262), .B(z2[98]), .Z(n7) );
  NANDN U18 ( .A(n3), .B(N362), .Z(n6) );
  NAND U19 ( .A(n8), .B(n9), .Z(z3[97]) );
  NANDN U20 ( .A(N262), .B(z2[97]), .Z(n9) );
  NANDN U21 ( .A(n3), .B(N361), .Z(n8) );
  NAND U22 ( .A(n10), .B(n11), .Z(z3[96]) );
  NANDN U23 ( .A(N262), .B(z2[96]), .Z(n11) );
  NANDN U24 ( .A(n3), .B(N360), .Z(n10) );
  NAND U25 ( .A(n12), .B(n13), .Z(z3[95]) );
  NANDN U26 ( .A(N262), .B(z2[95]), .Z(n13) );
  NANDN U27 ( .A(n3), .B(N359), .Z(n12) );
  NAND U28 ( .A(n14), .B(n23), .Z(z3[94]) );
  NANDN U29 ( .A(N262), .B(z2[94]), .Z(n23) );
  NANDN U30 ( .A(n3), .B(N358), .Z(n14) );
  NAND U31 ( .A(n24), .B(n25), .Z(z3[93]) );
  NANDN U32 ( .A(N262), .B(z2[93]), .Z(n25) );
  NANDN U33 ( .A(n3), .B(N357), .Z(n24) );
  NAND U34 ( .A(n26), .B(n27), .Z(z3[92]) );
  NANDN U35 ( .A(N262), .B(z2[92]), .Z(n27) );
  NANDN U36 ( .A(n3), .B(N356), .Z(n26) );
  NAND U37 ( .A(n28), .B(n29), .Z(z3[91]) );
  NANDN U38 ( .A(N262), .B(z2[91]), .Z(n29) );
  NANDN U39 ( .A(n3), .B(N355), .Z(n28) );
  NAND U40 ( .A(n30), .B(n31), .Z(z3[90]) );
  NANDN U41 ( .A(N262), .B(z2[90]), .Z(n31) );
  NANDN U42 ( .A(n3), .B(N354), .Z(n30) );
  NAND U43 ( .A(n32), .B(n33), .Z(z3[8]) );
  NANDN U44 ( .A(N262), .B(z2[8]), .Z(n33) );
  NANDN U45 ( .A(n3), .B(N272), .Z(n32) );
  NAND U46 ( .A(n34), .B(n35), .Z(z3[89]) );
  NANDN U47 ( .A(N262), .B(z2[89]), .Z(n35) );
  NANDN U48 ( .A(n3), .B(N353), .Z(n34) );
  NAND U49 ( .A(n36), .B(n37), .Z(z3[88]) );
  NANDN U50 ( .A(N262), .B(z2[88]), .Z(n37) );
  NANDN U51 ( .A(n3), .B(N352), .Z(n36) );
  NAND U52 ( .A(n38), .B(n39), .Z(z3[87]) );
  NANDN U53 ( .A(N262), .B(z2[87]), .Z(n39) );
  NANDN U54 ( .A(n3), .B(N351), .Z(n38) );
  NAND U55 ( .A(n40), .B(n41), .Z(z3[86]) );
  NANDN U56 ( .A(N262), .B(z2[86]), .Z(n41) );
  NANDN U57 ( .A(n3), .B(N350), .Z(n40) );
  NAND U58 ( .A(n42), .B(n43), .Z(z3[85]) );
  NANDN U59 ( .A(N262), .B(z2[85]), .Z(n43) );
  NANDN U60 ( .A(n3), .B(N349), .Z(n42) );
  NAND U61 ( .A(n44), .B(n45), .Z(z3[84]) );
  NANDN U62 ( .A(N262), .B(z2[84]), .Z(n45) );
  NANDN U63 ( .A(n3), .B(N348), .Z(n44) );
  NAND U64 ( .A(n46), .B(n47), .Z(z3[83]) );
  NANDN U65 ( .A(N262), .B(z2[83]), .Z(n47) );
  NANDN U66 ( .A(n3), .B(N347), .Z(n46) );
  NAND U67 ( .A(n48), .B(n49), .Z(z3[82]) );
  NANDN U68 ( .A(N262), .B(z2[82]), .Z(n49) );
  NANDN U69 ( .A(n3), .B(N346), .Z(n48) );
  NAND U70 ( .A(n50), .B(n51), .Z(z3[81]) );
  NANDN U71 ( .A(N262), .B(z2[81]), .Z(n51) );
  NANDN U72 ( .A(n3), .B(N345), .Z(n50) );
  NAND U73 ( .A(n52), .B(n53), .Z(z3[80]) );
  NANDN U74 ( .A(N262), .B(z2[80]), .Z(n53) );
  NANDN U75 ( .A(n3), .B(N344), .Z(n52) );
  NAND U76 ( .A(n54), .B(n55), .Z(z3[7]) );
  NANDN U77 ( .A(N262), .B(z2[7]), .Z(n55) );
  NANDN U78 ( .A(n3), .B(N271), .Z(n54) );
  NAND U79 ( .A(n56), .B(n57), .Z(z3[79]) );
  NANDN U80 ( .A(N262), .B(z2[79]), .Z(n57) );
  NANDN U81 ( .A(n3), .B(N343), .Z(n56) );
  NAND U82 ( .A(n58), .B(n59), .Z(z3[78]) );
  NANDN U83 ( .A(N262), .B(z2[78]), .Z(n59) );
  NANDN U84 ( .A(n3), .B(N342), .Z(n58) );
  NAND U85 ( .A(n60), .B(n61), .Z(z3[77]) );
  NANDN U86 ( .A(N262), .B(z2[77]), .Z(n61) );
  NANDN U87 ( .A(n3), .B(N341), .Z(n60) );
  NAND U88 ( .A(n62), .B(n63), .Z(z3[76]) );
  NANDN U89 ( .A(N262), .B(z2[76]), .Z(n63) );
  NANDN U90 ( .A(n3), .B(N340), .Z(n62) );
  NAND U91 ( .A(n64), .B(n65), .Z(z3[75]) );
  NANDN U92 ( .A(N262), .B(z2[75]), .Z(n65) );
  NANDN U93 ( .A(n3), .B(N339), .Z(n64) );
  NAND U94 ( .A(n66), .B(n67), .Z(z3[74]) );
  NANDN U95 ( .A(N262), .B(z2[74]), .Z(n67) );
  NANDN U96 ( .A(n3), .B(N338), .Z(n66) );
  NAND U97 ( .A(n68), .B(n69), .Z(z3[73]) );
  NANDN U98 ( .A(N262), .B(z2[73]), .Z(n69) );
  NANDN U99 ( .A(n3), .B(N337), .Z(n68) );
  NAND U100 ( .A(n70), .B(n71), .Z(z3[72]) );
  NANDN U101 ( .A(N262), .B(z2[72]), .Z(n71) );
  NANDN U102 ( .A(n3), .B(N336), .Z(n70) );
  NAND U103 ( .A(n72), .B(n73), .Z(z3[71]) );
  NANDN U104 ( .A(N262), .B(z2[71]), .Z(n73) );
  NANDN U105 ( .A(n3), .B(N335), .Z(n72) );
  NAND U106 ( .A(n74), .B(n75), .Z(z3[70]) );
  NANDN U107 ( .A(N262), .B(z2[70]), .Z(n75) );
  NANDN U108 ( .A(n3), .B(N334), .Z(n74) );
  NAND U109 ( .A(n76), .B(n77), .Z(z3[6]) );
  NANDN U110 ( .A(N262), .B(z2[6]), .Z(n77) );
  NANDN U111 ( .A(n3), .B(N270), .Z(n76) );
  NAND U112 ( .A(n78), .B(n79), .Z(z3[69]) );
  NANDN U113 ( .A(N262), .B(z2[69]), .Z(n79) );
  NANDN U114 ( .A(n3), .B(N333), .Z(n78) );
  NAND U115 ( .A(n80), .B(n81), .Z(z3[68]) );
  NANDN U116 ( .A(N262), .B(z2[68]), .Z(n81) );
  NANDN U117 ( .A(n3), .B(N332), .Z(n80) );
  NAND U118 ( .A(n82), .B(n83), .Z(z3[67]) );
  NANDN U119 ( .A(N262), .B(z2[67]), .Z(n83) );
  NANDN U120 ( .A(n3), .B(N331), .Z(n82) );
  NAND U121 ( .A(n84), .B(n85), .Z(z3[66]) );
  NANDN U122 ( .A(N262), .B(z2[66]), .Z(n85) );
  NANDN U123 ( .A(n3), .B(N330), .Z(n84) );
  NAND U124 ( .A(n86), .B(n87), .Z(z3[65]) );
  NANDN U125 ( .A(N262), .B(z2[65]), .Z(n87) );
  NANDN U126 ( .A(n3), .B(N329), .Z(n86) );
  NAND U127 ( .A(n88), .B(n89), .Z(z3[64]) );
  NANDN U128 ( .A(N262), .B(z2[64]), .Z(n89) );
  NANDN U129 ( .A(n3), .B(N328), .Z(n88) );
  NAND U130 ( .A(n90), .B(n91), .Z(z3[63]) );
  NANDN U131 ( .A(N262), .B(z2[63]), .Z(n91) );
  NANDN U132 ( .A(n3), .B(N327), .Z(n90) );
  NAND U133 ( .A(n92), .B(n93), .Z(z3[62]) );
  NANDN U134 ( .A(N262), .B(z2[62]), .Z(n93) );
  NANDN U135 ( .A(n3), .B(N326), .Z(n92) );
  NAND U136 ( .A(n94), .B(n95), .Z(z3[61]) );
  NANDN U137 ( .A(N262), .B(z2[61]), .Z(n95) );
  NANDN U138 ( .A(n3), .B(N325), .Z(n94) );
  NAND U139 ( .A(n96), .B(n97), .Z(z3[60]) );
  NANDN U140 ( .A(N262), .B(z2[60]), .Z(n97) );
  NANDN U141 ( .A(n3), .B(N324), .Z(n96) );
  NAND U142 ( .A(n98), .B(n99), .Z(z3[5]) );
  NANDN U143 ( .A(N262), .B(z2[5]), .Z(n99) );
  NANDN U144 ( .A(n3), .B(N269), .Z(n98) );
  NAND U145 ( .A(n100), .B(n101), .Z(z3[59]) );
  NANDN U146 ( .A(N262), .B(z2[59]), .Z(n101) );
  NANDN U147 ( .A(n3), .B(N323), .Z(n100) );
  NAND U148 ( .A(n102), .B(n103), .Z(z3[58]) );
  NANDN U149 ( .A(N262), .B(z2[58]), .Z(n103) );
  NANDN U150 ( .A(n3), .B(N322), .Z(n102) );
  NAND U151 ( .A(n104), .B(n105), .Z(z3[57]) );
  NANDN U152 ( .A(N262), .B(z2[57]), .Z(n105) );
  NANDN U153 ( .A(n3), .B(N321), .Z(n104) );
  NAND U154 ( .A(n106), .B(n107), .Z(z3[56]) );
  NANDN U155 ( .A(N262), .B(z2[56]), .Z(n107) );
  NANDN U156 ( .A(n3), .B(N320), .Z(n106) );
  NAND U157 ( .A(n108), .B(n109), .Z(z3[55]) );
  NANDN U158 ( .A(N262), .B(z2[55]), .Z(n109) );
  NANDN U159 ( .A(n3), .B(N319), .Z(n108) );
  NAND U160 ( .A(n110), .B(n111), .Z(z3[54]) );
  NANDN U161 ( .A(N262), .B(z2[54]), .Z(n111) );
  NANDN U162 ( .A(n3), .B(N318), .Z(n110) );
  NAND U163 ( .A(n112), .B(n113), .Z(z3[53]) );
  NANDN U164 ( .A(N262), .B(z2[53]), .Z(n113) );
  NANDN U165 ( .A(n3), .B(N317), .Z(n112) );
  NAND U166 ( .A(n114), .B(n115), .Z(z3[52]) );
  NANDN U167 ( .A(N262), .B(z2[52]), .Z(n115) );
  NANDN U168 ( .A(n3), .B(N316), .Z(n114) );
  NAND U169 ( .A(n116), .B(n117), .Z(z3[51]) );
  NANDN U170 ( .A(N262), .B(z2[51]), .Z(n117) );
  NANDN U171 ( .A(n3), .B(N315), .Z(n116) );
  NAND U172 ( .A(n118), .B(n119), .Z(z3[50]) );
  NANDN U173 ( .A(N262), .B(z2[50]), .Z(n119) );
  NANDN U174 ( .A(n3), .B(N314), .Z(n118) );
  NAND U175 ( .A(n120), .B(n121), .Z(z3[4]) );
  NANDN U176 ( .A(N262), .B(z2[4]), .Z(n121) );
  NANDN U177 ( .A(n3), .B(N268), .Z(n120) );
  NAND U178 ( .A(n122), .B(n123), .Z(z3[49]) );
  NANDN U179 ( .A(N262), .B(z2[49]), .Z(n123) );
  NANDN U180 ( .A(n3), .B(N313), .Z(n122) );
  NAND U181 ( .A(n124), .B(n125), .Z(z3[48]) );
  NANDN U182 ( .A(N262), .B(z2[48]), .Z(n125) );
  NANDN U183 ( .A(n3), .B(N312), .Z(n124) );
  NAND U184 ( .A(n126), .B(n127), .Z(z3[47]) );
  NANDN U185 ( .A(N262), .B(z2[47]), .Z(n127) );
  NANDN U186 ( .A(n3), .B(N311), .Z(n126) );
  NAND U187 ( .A(n128), .B(n129), .Z(z3[46]) );
  NANDN U188 ( .A(N262), .B(z2[46]), .Z(n129) );
  NANDN U189 ( .A(n3), .B(N310), .Z(n128) );
  NAND U190 ( .A(n130), .B(n131), .Z(z3[45]) );
  NANDN U191 ( .A(N262), .B(z2[45]), .Z(n131) );
  NANDN U192 ( .A(n3), .B(N309), .Z(n130) );
  NAND U193 ( .A(n132), .B(n133), .Z(z3[44]) );
  NANDN U194 ( .A(N262), .B(z2[44]), .Z(n133) );
  NANDN U195 ( .A(n3), .B(N308), .Z(n132) );
  NAND U196 ( .A(n134), .B(n135), .Z(z3[43]) );
  NANDN U197 ( .A(N262), .B(z2[43]), .Z(n135) );
  NANDN U198 ( .A(n3), .B(N307), .Z(n134) );
  NAND U199 ( .A(n136), .B(n137), .Z(z3[42]) );
  NANDN U200 ( .A(N262), .B(z2[42]), .Z(n137) );
  NANDN U201 ( .A(n3), .B(N306), .Z(n136) );
  NAND U202 ( .A(n138), .B(n139), .Z(z3[41]) );
  NANDN U203 ( .A(N262), .B(z2[41]), .Z(n139) );
  NANDN U204 ( .A(n3), .B(N305), .Z(n138) );
  NAND U205 ( .A(n140), .B(n141), .Z(z3[40]) );
  NANDN U206 ( .A(N262), .B(z2[40]), .Z(n141) );
  NANDN U207 ( .A(n3), .B(N304), .Z(n140) );
  NAND U208 ( .A(n142), .B(n143), .Z(z3[3]) );
  NANDN U209 ( .A(N262), .B(z2[3]), .Z(n143) );
  NANDN U210 ( .A(n3), .B(N267), .Z(n142) );
  NAND U211 ( .A(n144), .B(n145), .Z(z3[39]) );
  NANDN U212 ( .A(N262), .B(z2[39]), .Z(n145) );
  NANDN U213 ( .A(n3), .B(N303), .Z(n144) );
  NAND U214 ( .A(n146), .B(n147), .Z(z3[38]) );
  NANDN U215 ( .A(N262), .B(z2[38]), .Z(n147) );
  NANDN U216 ( .A(n3), .B(N302), .Z(n146) );
  NAND U217 ( .A(n148), .B(n149), .Z(z3[37]) );
  NANDN U218 ( .A(N262), .B(z2[37]), .Z(n149) );
  NANDN U219 ( .A(n3), .B(N301), .Z(n148) );
  NAND U220 ( .A(n150), .B(n151), .Z(z3[36]) );
  NANDN U221 ( .A(N262), .B(z2[36]), .Z(n151) );
  NANDN U222 ( .A(n3), .B(N300), .Z(n150) );
  NAND U223 ( .A(n152), .B(n153), .Z(z3[35]) );
  NANDN U224 ( .A(N262), .B(z2[35]), .Z(n153) );
  NANDN U225 ( .A(n3), .B(N299), .Z(n152) );
  NAND U226 ( .A(n154), .B(n155), .Z(z3[34]) );
  NANDN U227 ( .A(N262), .B(z2[34]), .Z(n155) );
  NANDN U228 ( .A(n3), .B(N298), .Z(n154) );
  NAND U229 ( .A(n156), .B(n157), .Z(z3[33]) );
  NANDN U230 ( .A(N262), .B(z2[33]), .Z(n157) );
  NANDN U231 ( .A(n3), .B(N297), .Z(n156) );
  NAND U232 ( .A(n158), .B(n159), .Z(z3[32]) );
  NANDN U233 ( .A(N262), .B(z2[32]), .Z(n159) );
  NANDN U234 ( .A(n3), .B(N296), .Z(n158) );
  NAND U235 ( .A(n160), .B(n161), .Z(z3[31]) );
  NANDN U236 ( .A(N262), .B(z2[31]), .Z(n161) );
  NANDN U237 ( .A(n3), .B(N295), .Z(n160) );
  NAND U238 ( .A(n162), .B(n163), .Z(z3[30]) );
  NANDN U239 ( .A(N262), .B(z2[30]), .Z(n163) );
  NANDN U240 ( .A(n3), .B(N294), .Z(n162) );
  NAND U241 ( .A(n164), .B(n165), .Z(z3[2]) );
  NANDN U242 ( .A(N262), .B(z2[2]), .Z(n165) );
  NANDN U243 ( .A(n3), .B(N266), .Z(n164) );
  NAND U244 ( .A(n166), .B(n167), .Z(z3[29]) );
  NANDN U245 ( .A(N262), .B(z2[29]), .Z(n167) );
  NANDN U246 ( .A(n3), .B(N293), .Z(n166) );
  NAND U247 ( .A(n168), .B(n169), .Z(z3[28]) );
  NANDN U248 ( .A(N262), .B(z2[28]), .Z(n169) );
  NANDN U249 ( .A(n3), .B(N292), .Z(n168) );
  NAND U250 ( .A(n170), .B(n171), .Z(z3[27]) );
  NANDN U251 ( .A(N262), .B(z2[27]), .Z(n171) );
  NANDN U252 ( .A(n3), .B(N291), .Z(n170) );
  NAND U253 ( .A(n172), .B(n173), .Z(z3[26]) );
  NANDN U254 ( .A(N262), .B(z2[26]), .Z(n173) );
  NANDN U255 ( .A(n3), .B(N290), .Z(n172) );
  NAND U256 ( .A(n174), .B(n175), .Z(z3[25]) );
  NANDN U257 ( .A(N262), .B(z2[25]), .Z(n175) );
  NANDN U258 ( .A(n3), .B(N289), .Z(n174) );
  NAND U259 ( .A(n176), .B(n177), .Z(z3[257]) );
  NANDN U260 ( .A(N262), .B(z2[257]), .Z(n177) );
  NANDN U261 ( .A(n3), .B(N521), .Z(n176) );
  NAND U262 ( .A(n178), .B(n179), .Z(z3[256]) );
  NANDN U263 ( .A(N262), .B(z2[256]), .Z(n179) );
  NANDN U264 ( .A(n3), .B(N520), .Z(n178) );
  NAND U265 ( .A(n180), .B(n181), .Z(z3[255]) );
  NANDN U266 ( .A(N262), .B(z2[255]), .Z(n181) );
  NANDN U267 ( .A(n3), .B(N519), .Z(n180) );
  NAND U268 ( .A(n182), .B(n183), .Z(z3[254]) );
  NANDN U269 ( .A(N262), .B(z2[254]), .Z(n183) );
  NANDN U270 ( .A(n3), .B(N518), .Z(n182) );
  NAND U271 ( .A(n184), .B(n185), .Z(z3[253]) );
  NANDN U272 ( .A(N262), .B(z2[253]), .Z(n185) );
  NANDN U273 ( .A(n3), .B(N517), .Z(n184) );
  NAND U274 ( .A(n186), .B(n187), .Z(z3[252]) );
  NANDN U275 ( .A(N262), .B(z2[252]), .Z(n187) );
  NANDN U276 ( .A(n3), .B(N516), .Z(n186) );
  NAND U277 ( .A(n188), .B(n189), .Z(z3[251]) );
  NANDN U278 ( .A(N262), .B(z2[251]), .Z(n189) );
  NANDN U279 ( .A(n3), .B(N515), .Z(n188) );
  NAND U280 ( .A(n190), .B(n191), .Z(z3[250]) );
  NANDN U281 ( .A(N262), .B(z2[250]), .Z(n191) );
  NANDN U282 ( .A(n3), .B(N514), .Z(n190) );
  NAND U283 ( .A(n192), .B(n193), .Z(z3[24]) );
  NANDN U284 ( .A(N262), .B(z2[24]), .Z(n193) );
  NANDN U285 ( .A(n3), .B(N288), .Z(n192) );
  NAND U286 ( .A(n194), .B(n195), .Z(z3[249]) );
  NANDN U287 ( .A(N262), .B(z2[249]), .Z(n195) );
  NANDN U288 ( .A(n3), .B(N513), .Z(n194) );
  NAND U289 ( .A(n196), .B(n197), .Z(z3[248]) );
  NANDN U290 ( .A(N262), .B(z2[248]), .Z(n197) );
  NANDN U291 ( .A(n3), .B(N512), .Z(n196) );
  NAND U292 ( .A(n198), .B(n199), .Z(z3[247]) );
  NANDN U293 ( .A(N262), .B(z2[247]), .Z(n199) );
  NANDN U294 ( .A(n3), .B(N511), .Z(n198) );
  NAND U295 ( .A(n200), .B(n201), .Z(z3[246]) );
  NANDN U296 ( .A(N262), .B(z2[246]), .Z(n201) );
  NANDN U297 ( .A(n3), .B(N510), .Z(n200) );
  NAND U298 ( .A(n202), .B(n203), .Z(z3[245]) );
  NANDN U299 ( .A(N262), .B(z2[245]), .Z(n203) );
  NANDN U300 ( .A(n3), .B(N509), .Z(n202) );
  NAND U301 ( .A(n204), .B(n205), .Z(z3[244]) );
  NANDN U302 ( .A(N262), .B(z2[244]), .Z(n205) );
  NANDN U303 ( .A(n3), .B(N508), .Z(n204) );
  NAND U304 ( .A(n206), .B(n207), .Z(z3[243]) );
  NANDN U305 ( .A(N262), .B(z2[243]), .Z(n207) );
  NANDN U306 ( .A(n3), .B(N507), .Z(n206) );
  NAND U307 ( .A(n208), .B(n209), .Z(z3[242]) );
  NANDN U308 ( .A(N262), .B(z2[242]), .Z(n209) );
  NANDN U309 ( .A(n3), .B(N506), .Z(n208) );
  NAND U310 ( .A(n210), .B(n211), .Z(z3[241]) );
  NANDN U311 ( .A(N262), .B(z2[241]), .Z(n211) );
  NANDN U312 ( .A(n3), .B(N505), .Z(n210) );
  NAND U313 ( .A(n212), .B(n213), .Z(z3[240]) );
  NANDN U314 ( .A(N262), .B(z2[240]), .Z(n213) );
  NANDN U315 ( .A(n3), .B(N504), .Z(n212) );
  NAND U316 ( .A(n214), .B(n215), .Z(z3[23]) );
  NANDN U317 ( .A(N262), .B(z2[23]), .Z(n215) );
  NANDN U318 ( .A(n3), .B(N287), .Z(n214) );
  NAND U319 ( .A(n216), .B(n217), .Z(z3[239]) );
  NANDN U320 ( .A(N262), .B(z2[239]), .Z(n217) );
  NANDN U321 ( .A(n3), .B(N503), .Z(n216) );
  NAND U322 ( .A(n218), .B(n219), .Z(z3[238]) );
  NANDN U323 ( .A(N262), .B(z2[238]), .Z(n219) );
  NANDN U324 ( .A(n3), .B(N502), .Z(n218) );
  NAND U325 ( .A(n220), .B(n221), .Z(z3[237]) );
  NANDN U326 ( .A(N262), .B(z2[237]), .Z(n221) );
  NANDN U327 ( .A(n3), .B(N501), .Z(n220) );
  NAND U328 ( .A(n222), .B(n223), .Z(z3[236]) );
  NANDN U329 ( .A(N262), .B(z2[236]), .Z(n223) );
  NANDN U330 ( .A(n3), .B(N500), .Z(n222) );
  NAND U331 ( .A(n224), .B(n225), .Z(z3[235]) );
  NANDN U332 ( .A(N262), .B(z2[235]), .Z(n225) );
  NANDN U333 ( .A(n3), .B(N499), .Z(n224) );
  NAND U334 ( .A(n226), .B(n227), .Z(z3[234]) );
  NANDN U335 ( .A(N262), .B(z2[234]), .Z(n227) );
  NANDN U336 ( .A(n3), .B(N498), .Z(n226) );
  NAND U337 ( .A(n228), .B(n229), .Z(z3[233]) );
  NANDN U338 ( .A(N262), .B(z2[233]), .Z(n229) );
  NANDN U339 ( .A(n3), .B(N497), .Z(n228) );
  NAND U340 ( .A(n230), .B(n231), .Z(z3[232]) );
  NANDN U341 ( .A(N262), .B(z2[232]), .Z(n231) );
  NANDN U342 ( .A(n3), .B(N496), .Z(n230) );
  NAND U343 ( .A(n232), .B(n233), .Z(z3[231]) );
  NANDN U344 ( .A(N262), .B(z2[231]), .Z(n233) );
  NANDN U345 ( .A(n3), .B(N495), .Z(n232) );
  NAND U346 ( .A(n234), .B(n235), .Z(z3[230]) );
  NANDN U347 ( .A(N262), .B(z2[230]), .Z(n235) );
  NANDN U348 ( .A(n3), .B(N494), .Z(n234) );
  NAND U349 ( .A(n236), .B(n237), .Z(z3[22]) );
  NANDN U350 ( .A(N262), .B(z2[22]), .Z(n237) );
  NANDN U351 ( .A(n3), .B(N286), .Z(n236) );
  NAND U352 ( .A(n238), .B(n239), .Z(z3[229]) );
  NANDN U353 ( .A(N262), .B(z2[229]), .Z(n239) );
  NANDN U354 ( .A(n3), .B(N493), .Z(n238) );
  NAND U355 ( .A(n240), .B(n241), .Z(z3[228]) );
  NANDN U356 ( .A(N262), .B(z2[228]), .Z(n241) );
  NANDN U357 ( .A(n3), .B(N492), .Z(n240) );
  NAND U358 ( .A(n242), .B(n243), .Z(z3[227]) );
  NANDN U359 ( .A(N262), .B(z2[227]), .Z(n243) );
  NANDN U360 ( .A(n3), .B(N491), .Z(n242) );
  NAND U361 ( .A(n244), .B(n245), .Z(z3[226]) );
  NANDN U362 ( .A(N262), .B(z2[226]), .Z(n245) );
  NANDN U363 ( .A(n3), .B(N490), .Z(n244) );
  NAND U364 ( .A(n246), .B(n247), .Z(z3[225]) );
  NANDN U365 ( .A(N262), .B(z2[225]), .Z(n247) );
  NANDN U366 ( .A(n3), .B(N489), .Z(n246) );
  NAND U367 ( .A(n248), .B(n249), .Z(z3[224]) );
  NANDN U368 ( .A(N262), .B(z2[224]), .Z(n249) );
  NANDN U369 ( .A(n3), .B(N488), .Z(n248) );
  NAND U370 ( .A(n250), .B(n251), .Z(z3[223]) );
  NANDN U371 ( .A(N262), .B(z2[223]), .Z(n251) );
  NANDN U372 ( .A(n3), .B(N487), .Z(n250) );
  NAND U373 ( .A(n252), .B(n253), .Z(z3[222]) );
  NANDN U374 ( .A(N262), .B(z2[222]), .Z(n253) );
  NANDN U375 ( .A(n3), .B(N486), .Z(n252) );
  NAND U376 ( .A(n254), .B(n255), .Z(z3[221]) );
  NANDN U377 ( .A(N262), .B(z2[221]), .Z(n255) );
  NANDN U378 ( .A(n3), .B(N485), .Z(n254) );
  NAND U379 ( .A(n256), .B(n257), .Z(z3[220]) );
  NANDN U380 ( .A(N262), .B(z2[220]), .Z(n257) );
  NANDN U381 ( .A(n3), .B(N484), .Z(n256) );
  NAND U382 ( .A(n258), .B(n259), .Z(z3[21]) );
  NANDN U383 ( .A(N262), .B(z2[21]), .Z(n259) );
  NANDN U384 ( .A(n3), .B(N285), .Z(n258) );
  NAND U385 ( .A(n260), .B(n261), .Z(z3[219]) );
  NANDN U386 ( .A(N262), .B(z2[219]), .Z(n261) );
  NANDN U387 ( .A(n3), .B(N483), .Z(n260) );
  NAND U388 ( .A(n262), .B(n263), .Z(z3[218]) );
  NANDN U389 ( .A(N262), .B(z2[218]), .Z(n263) );
  NANDN U390 ( .A(n3), .B(N482), .Z(n262) );
  NAND U391 ( .A(n264), .B(n265), .Z(z3[217]) );
  NANDN U392 ( .A(N262), .B(z2[217]), .Z(n265) );
  NANDN U393 ( .A(n3), .B(N481), .Z(n264) );
  NAND U394 ( .A(n266), .B(n267), .Z(z3[216]) );
  NANDN U395 ( .A(N262), .B(z2[216]), .Z(n267) );
  NANDN U396 ( .A(n3), .B(N480), .Z(n266) );
  NAND U397 ( .A(n268), .B(n269), .Z(z3[215]) );
  NANDN U398 ( .A(N262), .B(z2[215]), .Z(n269) );
  NANDN U399 ( .A(n3), .B(N479), .Z(n268) );
  NAND U400 ( .A(n270), .B(n271), .Z(z3[214]) );
  NANDN U401 ( .A(N262), .B(z2[214]), .Z(n271) );
  NANDN U402 ( .A(n3), .B(N478), .Z(n270) );
  NAND U403 ( .A(n272), .B(n273), .Z(z3[213]) );
  NANDN U404 ( .A(N262), .B(z2[213]), .Z(n273) );
  NANDN U405 ( .A(n3), .B(N477), .Z(n272) );
  NAND U406 ( .A(n274), .B(n275), .Z(z3[212]) );
  NANDN U407 ( .A(N262), .B(z2[212]), .Z(n275) );
  NANDN U408 ( .A(n3), .B(N476), .Z(n274) );
  NAND U409 ( .A(n276), .B(n277), .Z(z3[211]) );
  NANDN U410 ( .A(N262), .B(z2[211]), .Z(n277) );
  NANDN U411 ( .A(n3), .B(N475), .Z(n276) );
  NAND U412 ( .A(n278), .B(n279), .Z(z3[210]) );
  NANDN U413 ( .A(N262), .B(z2[210]), .Z(n279) );
  NANDN U414 ( .A(n3), .B(N474), .Z(n278) );
  NAND U415 ( .A(n280), .B(n281), .Z(z3[20]) );
  NANDN U416 ( .A(N262), .B(z2[20]), .Z(n281) );
  NANDN U417 ( .A(n3), .B(N284), .Z(n280) );
  NAND U418 ( .A(n282), .B(n283), .Z(z3[209]) );
  NANDN U419 ( .A(N262), .B(z2[209]), .Z(n283) );
  NANDN U420 ( .A(n3), .B(N473), .Z(n282) );
  NAND U421 ( .A(n284), .B(n285), .Z(z3[208]) );
  NANDN U422 ( .A(N262), .B(z2[208]), .Z(n285) );
  NANDN U423 ( .A(n3), .B(N472), .Z(n284) );
  NAND U424 ( .A(n286), .B(n287), .Z(z3[207]) );
  NANDN U425 ( .A(N262), .B(z2[207]), .Z(n287) );
  NANDN U426 ( .A(n3), .B(N471), .Z(n286) );
  NAND U427 ( .A(n288), .B(n289), .Z(z3[206]) );
  NANDN U428 ( .A(N262), .B(z2[206]), .Z(n289) );
  NANDN U429 ( .A(n3), .B(N470), .Z(n288) );
  NAND U430 ( .A(n290), .B(n291), .Z(z3[205]) );
  NANDN U431 ( .A(N262), .B(z2[205]), .Z(n291) );
  NANDN U432 ( .A(n3), .B(N469), .Z(n290) );
  NAND U433 ( .A(n292), .B(n293), .Z(z3[204]) );
  NANDN U434 ( .A(N262), .B(z2[204]), .Z(n293) );
  NANDN U435 ( .A(n3), .B(N468), .Z(n292) );
  NAND U436 ( .A(n294), .B(n295), .Z(z3[203]) );
  NANDN U437 ( .A(N262), .B(z2[203]), .Z(n295) );
  NANDN U438 ( .A(n3), .B(N467), .Z(n294) );
  NAND U439 ( .A(n296), .B(n297), .Z(z3[202]) );
  NANDN U440 ( .A(N262), .B(z2[202]), .Z(n297) );
  NANDN U441 ( .A(n3), .B(N466), .Z(n296) );
  NAND U442 ( .A(n298), .B(n299), .Z(z3[201]) );
  NANDN U443 ( .A(N262), .B(z2[201]), .Z(n299) );
  NANDN U444 ( .A(n3), .B(N465), .Z(n298) );
  NAND U445 ( .A(n300), .B(n301), .Z(z3[200]) );
  NANDN U446 ( .A(N262), .B(z2[200]), .Z(n301) );
  NANDN U447 ( .A(n3), .B(N464), .Z(n300) );
  NAND U448 ( .A(n302), .B(n303), .Z(z3[1]) );
  NANDN U449 ( .A(N262), .B(z2[1]), .Z(n303) );
  NANDN U450 ( .A(n3), .B(N265), .Z(n302) );
  NAND U451 ( .A(n304), .B(n305), .Z(z3[19]) );
  NANDN U452 ( .A(N262), .B(z2[19]), .Z(n305) );
  NANDN U453 ( .A(n3), .B(N283), .Z(n304) );
  NAND U454 ( .A(n306), .B(n307), .Z(z3[199]) );
  NANDN U455 ( .A(N262), .B(z2[199]), .Z(n307) );
  NANDN U456 ( .A(n3), .B(N463), .Z(n306) );
  NAND U457 ( .A(n308), .B(n309), .Z(z3[198]) );
  NANDN U458 ( .A(N262), .B(z2[198]), .Z(n309) );
  NANDN U459 ( .A(n3), .B(N462), .Z(n308) );
  NAND U460 ( .A(n310), .B(n311), .Z(z3[197]) );
  NANDN U461 ( .A(N262), .B(z2[197]), .Z(n311) );
  NANDN U462 ( .A(n3), .B(N461), .Z(n310) );
  NAND U463 ( .A(n312), .B(n313), .Z(z3[196]) );
  NANDN U464 ( .A(N262), .B(z2[196]), .Z(n313) );
  NANDN U465 ( .A(n3), .B(N460), .Z(n312) );
  NAND U466 ( .A(n314), .B(n315), .Z(z3[195]) );
  NANDN U467 ( .A(N262), .B(z2[195]), .Z(n315) );
  NANDN U468 ( .A(n3), .B(N459), .Z(n314) );
  NAND U469 ( .A(n316), .B(n317), .Z(z3[194]) );
  NANDN U470 ( .A(N262), .B(z2[194]), .Z(n317) );
  NANDN U471 ( .A(n3), .B(N458), .Z(n316) );
  NAND U472 ( .A(n318), .B(n319), .Z(z3[193]) );
  NANDN U473 ( .A(N262), .B(z2[193]), .Z(n319) );
  NANDN U474 ( .A(n3), .B(N457), .Z(n318) );
  NAND U475 ( .A(n320), .B(n321), .Z(z3[192]) );
  NANDN U476 ( .A(N262), .B(z2[192]), .Z(n321) );
  NANDN U477 ( .A(n3), .B(N456), .Z(n320) );
  NAND U478 ( .A(n322), .B(n323), .Z(z3[191]) );
  NANDN U479 ( .A(N262), .B(z2[191]), .Z(n323) );
  NANDN U480 ( .A(n3), .B(N455), .Z(n322) );
  NAND U481 ( .A(n324), .B(n325), .Z(z3[190]) );
  NANDN U482 ( .A(N262), .B(z2[190]), .Z(n325) );
  NANDN U483 ( .A(n3), .B(N454), .Z(n324) );
  NAND U484 ( .A(n326), .B(n327), .Z(z3[18]) );
  NANDN U485 ( .A(N262), .B(z2[18]), .Z(n327) );
  NANDN U486 ( .A(n3), .B(N282), .Z(n326) );
  NAND U487 ( .A(n328), .B(n329), .Z(z3[189]) );
  NANDN U488 ( .A(N262), .B(z2[189]), .Z(n329) );
  NANDN U489 ( .A(n3), .B(N453), .Z(n328) );
  NAND U490 ( .A(n330), .B(n331), .Z(z3[188]) );
  NANDN U491 ( .A(N262), .B(z2[188]), .Z(n331) );
  NANDN U492 ( .A(n3), .B(N452), .Z(n330) );
  NAND U493 ( .A(n332), .B(n333), .Z(z3[187]) );
  NANDN U494 ( .A(N262), .B(z2[187]), .Z(n333) );
  NANDN U495 ( .A(n3), .B(N451), .Z(n332) );
  NAND U496 ( .A(n334), .B(n335), .Z(z3[186]) );
  NANDN U497 ( .A(N262), .B(z2[186]), .Z(n335) );
  NANDN U498 ( .A(n3), .B(N450), .Z(n334) );
  NAND U499 ( .A(n336), .B(n337), .Z(z3[185]) );
  NANDN U500 ( .A(N262), .B(z2[185]), .Z(n337) );
  NANDN U501 ( .A(n3), .B(N449), .Z(n336) );
  NAND U502 ( .A(n338), .B(n339), .Z(z3[184]) );
  NANDN U503 ( .A(N262), .B(z2[184]), .Z(n339) );
  NANDN U504 ( .A(n3), .B(N448), .Z(n338) );
  NAND U505 ( .A(n340), .B(n341), .Z(z3[183]) );
  NANDN U506 ( .A(N262), .B(z2[183]), .Z(n341) );
  NANDN U507 ( .A(n3), .B(N447), .Z(n340) );
  NAND U508 ( .A(n342), .B(n343), .Z(z3[182]) );
  NANDN U509 ( .A(N262), .B(z2[182]), .Z(n343) );
  NANDN U510 ( .A(n3), .B(N446), .Z(n342) );
  NAND U511 ( .A(n344), .B(n345), .Z(z3[181]) );
  NANDN U512 ( .A(N262), .B(z2[181]), .Z(n345) );
  NANDN U513 ( .A(n3), .B(N445), .Z(n344) );
  NAND U514 ( .A(n346), .B(n347), .Z(z3[180]) );
  NANDN U515 ( .A(N262), .B(z2[180]), .Z(n347) );
  NANDN U516 ( .A(n3), .B(N444), .Z(n346) );
  NAND U517 ( .A(n348), .B(n349), .Z(z3[17]) );
  NANDN U518 ( .A(N262), .B(z2[17]), .Z(n349) );
  NANDN U519 ( .A(n3), .B(N281), .Z(n348) );
  NAND U520 ( .A(n350), .B(n351), .Z(z3[179]) );
  NANDN U521 ( .A(N262), .B(z2[179]), .Z(n351) );
  NANDN U522 ( .A(n3), .B(N443), .Z(n350) );
  NAND U523 ( .A(n352), .B(n353), .Z(z3[178]) );
  NANDN U524 ( .A(N262), .B(z2[178]), .Z(n353) );
  NANDN U525 ( .A(n3), .B(N442), .Z(n352) );
  NAND U526 ( .A(n354), .B(n355), .Z(z3[177]) );
  NANDN U527 ( .A(N262), .B(z2[177]), .Z(n355) );
  NANDN U528 ( .A(n3), .B(N441), .Z(n354) );
  NAND U529 ( .A(n356), .B(n357), .Z(z3[176]) );
  NANDN U530 ( .A(N262), .B(z2[176]), .Z(n357) );
  NANDN U531 ( .A(n3), .B(N440), .Z(n356) );
  NAND U532 ( .A(n358), .B(n359), .Z(z3[175]) );
  NANDN U533 ( .A(N262), .B(z2[175]), .Z(n359) );
  NANDN U534 ( .A(n3), .B(N439), .Z(n358) );
  NAND U535 ( .A(n360), .B(n361), .Z(z3[174]) );
  NANDN U536 ( .A(N262), .B(z2[174]), .Z(n361) );
  NANDN U537 ( .A(n3), .B(N438), .Z(n360) );
  NAND U538 ( .A(n362), .B(n363), .Z(z3[173]) );
  NANDN U539 ( .A(N262), .B(z2[173]), .Z(n363) );
  NANDN U540 ( .A(n3), .B(N437), .Z(n362) );
  NAND U541 ( .A(n364), .B(n365), .Z(z3[172]) );
  NANDN U542 ( .A(N262), .B(z2[172]), .Z(n365) );
  NANDN U543 ( .A(n3), .B(N436), .Z(n364) );
  NAND U544 ( .A(n366), .B(n367), .Z(z3[171]) );
  NANDN U545 ( .A(N262), .B(z2[171]), .Z(n367) );
  NANDN U546 ( .A(n3), .B(N435), .Z(n366) );
  NAND U547 ( .A(n368), .B(n369), .Z(z3[170]) );
  NANDN U548 ( .A(N262), .B(z2[170]), .Z(n369) );
  NANDN U549 ( .A(n3), .B(N434), .Z(n368) );
  NAND U550 ( .A(n370), .B(n371), .Z(z3[16]) );
  NANDN U551 ( .A(N262), .B(z2[16]), .Z(n371) );
  NANDN U552 ( .A(n3), .B(N280), .Z(n370) );
  NAND U553 ( .A(n372), .B(n373), .Z(z3[169]) );
  NANDN U554 ( .A(N262), .B(z2[169]), .Z(n373) );
  NANDN U555 ( .A(n3), .B(N433), .Z(n372) );
  NAND U556 ( .A(n374), .B(n375), .Z(z3[168]) );
  NANDN U557 ( .A(N262), .B(z2[168]), .Z(n375) );
  NANDN U558 ( .A(n3), .B(N432), .Z(n374) );
  NAND U559 ( .A(n376), .B(n377), .Z(z3[167]) );
  NANDN U560 ( .A(N262), .B(z2[167]), .Z(n377) );
  NANDN U561 ( .A(n3), .B(N431), .Z(n376) );
  NAND U562 ( .A(n378), .B(n379), .Z(z3[166]) );
  NANDN U563 ( .A(N262), .B(z2[166]), .Z(n379) );
  NANDN U564 ( .A(n3), .B(N430), .Z(n378) );
  NAND U565 ( .A(n380), .B(n381), .Z(z3[165]) );
  NANDN U566 ( .A(N262), .B(z2[165]), .Z(n381) );
  NANDN U567 ( .A(n3), .B(N429), .Z(n380) );
  NAND U568 ( .A(n382), .B(n383), .Z(z3[164]) );
  NANDN U569 ( .A(N262), .B(z2[164]), .Z(n383) );
  NANDN U570 ( .A(n3), .B(N428), .Z(n382) );
  NAND U571 ( .A(n384), .B(n385), .Z(z3[163]) );
  NANDN U572 ( .A(N262), .B(z2[163]), .Z(n385) );
  NANDN U573 ( .A(n3), .B(N427), .Z(n384) );
  NAND U574 ( .A(n386), .B(n387), .Z(z3[162]) );
  NANDN U575 ( .A(N262), .B(z2[162]), .Z(n387) );
  NANDN U576 ( .A(n3), .B(N426), .Z(n386) );
  NAND U577 ( .A(n388), .B(n389), .Z(z3[161]) );
  NANDN U578 ( .A(N262), .B(z2[161]), .Z(n389) );
  NANDN U579 ( .A(n3), .B(N425), .Z(n388) );
  NAND U580 ( .A(n390), .B(n391), .Z(z3[160]) );
  NANDN U581 ( .A(N262), .B(z2[160]), .Z(n391) );
  NANDN U582 ( .A(n3), .B(N424), .Z(n390) );
  NAND U583 ( .A(n392), .B(n393), .Z(z3[15]) );
  NANDN U584 ( .A(N262), .B(z2[15]), .Z(n393) );
  NANDN U585 ( .A(n3), .B(N279), .Z(n392) );
  NAND U586 ( .A(n394), .B(n395), .Z(z3[159]) );
  NANDN U587 ( .A(N262), .B(z2[159]), .Z(n395) );
  NANDN U588 ( .A(n3), .B(N423), .Z(n394) );
  NAND U589 ( .A(n396), .B(n397), .Z(z3[158]) );
  NANDN U590 ( .A(N262), .B(z2[158]), .Z(n397) );
  NANDN U591 ( .A(n3), .B(N422), .Z(n396) );
  NAND U592 ( .A(n398), .B(n399), .Z(z3[157]) );
  NANDN U593 ( .A(N262), .B(z2[157]), .Z(n399) );
  NANDN U594 ( .A(n3), .B(N421), .Z(n398) );
  NAND U595 ( .A(n400), .B(n401), .Z(z3[156]) );
  NANDN U596 ( .A(N262), .B(z2[156]), .Z(n401) );
  NANDN U597 ( .A(n3), .B(N420), .Z(n400) );
  NAND U598 ( .A(n402), .B(n403), .Z(z3[155]) );
  NANDN U599 ( .A(N262), .B(z2[155]), .Z(n403) );
  NANDN U600 ( .A(n3), .B(N419), .Z(n402) );
  NAND U601 ( .A(n404), .B(n405), .Z(z3[154]) );
  NANDN U602 ( .A(N262), .B(z2[154]), .Z(n405) );
  NANDN U603 ( .A(n3), .B(N418), .Z(n404) );
  NAND U604 ( .A(n406), .B(n407), .Z(z3[153]) );
  NANDN U605 ( .A(N262), .B(z2[153]), .Z(n407) );
  NANDN U606 ( .A(n3), .B(N417), .Z(n406) );
  NAND U607 ( .A(n408), .B(n409), .Z(z3[152]) );
  NANDN U608 ( .A(N262), .B(z2[152]), .Z(n409) );
  NANDN U609 ( .A(n3), .B(N416), .Z(n408) );
  NAND U610 ( .A(n410), .B(n411), .Z(z3[151]) );
  NANDN U611 ( .A(N262), .B(z2[151]), .Z(n411) );
  NANDN U612 ( .A(n3), .B(N415), .Z(n410) );
  NAND U613 ( .A(n412), .B(n413), .Z(z3[150]) );
  NANDN U614 ( .A(N262), .B(z2[150]), .Z(n413) );
  NANDN U615 ( .A(n3), .B(N414), .Z(n412) );
  NAND U616 ( .A(n414), .B(n415), .Z(z3[14]) );
  NANDN U617 ( .A(N262), .B(z2[14]), .Z(n415) );
  NANDN U618 ( .A(n3), .B(N278), .Z(n414) );
  NAND U619 ( .A(n416), .B(n417), .Z(z3[149]) );
  NANDN U620 ( .A(N262), .B(z2[149]), .Z(n417) );
  NANDN U621 ( .A(n3), .B(N413), .Z(n416) );
  NAND U622 ( .A(n418), .B(n419), .Z(z3[148]) );
  NANDN U623 ( .A(N262), .B(z2[148]), .Z(n419) );
  NANDN U624 ( .A(n3), .B(N412), .Z(n418) );
  NAND U625 ( .A(n420), .B(n421), .Z(z3[147]) );
  NANDN U626 ( .A(N262), .B(z2[147]), .Z(n421) );
  NANDN U627 ( .A(n3), .B(N411), .Z(n420) );
  NAND U628 ( .A(n422), .B(n423), .Z(z3[146]) );
  NANDN U629 ( .A(N262), .B(z2[146]), .Z(n423) );
  NANDN U630 ( .A(n3), .B(N410), .Z(n422) );
  NAND U631 ( .A(n424), .B(n425), .Z(z3[145]) );
  NANDN U632 ( .A(N262), .B(z2[145]), .Z(n425) );
  NANDN U633 ( .A(n3), .B(N409), .Z(n424) );
  NAND U634 ( .A(n426), .B(n427), .Z(z3[144]) );
  NANDN U635 ( .A(N262), .B(z2[144]), .Z(n427) );
  NANDN U636 ( .A(n3), .B(N408), .Z(n426) );
  NAND U637 ( .A(n428), .B(n429), .Z(z3[143]) );
  NANDN U638 ( .A(N262), .B(z2[143]), .Z(n429) );
  NANDN U639 ( .A(n3), .B(N407), .Z(n428) );
  NAND U640 ( .A(n430), .B(n431), .Z(z3[142]) );
  NANDN U641 ( .A(N262), .B(z2[142]), .Z(n431) );
  NANDN U642 ( .A(n3), .B(N406), .Z(n430) );
  NAND U643 ( .A(n432), .B(n433), .Z(z3[141]) );
  NANDN U644 ( .A(N262), .B(z2[141]), .Z(n433) );
  NANDN U645 ( .A(n3), .B(N405), .Z(n432) );
  NAND U646 ( .A(n434), .B(n435), .Z(z3[140]) );
  NANDN U647 ( .A(N262), .B(z2[140]), .Z(n435) );
  NANDN U648 ( .A(n3), .B(N404), .Z(n434) );
  NAND U649 ( .A(n436), .B(n437), .Z(z3[13]) );
  NANDN U650 ( .A(N262), .B(z2[13]), .Z(n437) );
  NANDN U651 ( .A(n3), .B(N277), .Z(n436) );
  NAND U652 ( .A(n438), .B(n439), .Z(z3[139]) );
  NANDN U653 ( .A(N262), .B(z2[139]), .Z(n439) );
  NANDN U654 ( .A(n3), .B(N403), .Z(n438) );
  NAND U655 ( .A(n440), .B(n441), .Z(z3[138]) );
  NANDN U656 ( .A(N262), .B(z2[138]), .Z(n441) );
  NANDN U657 ( .A(n3), .B(N402), .Z(n440) );
  NAND U658 ( .A(n442), .B(n443), .Z(z3[137]) );
  NANDN U659 ( .A(N262), .B(z2[137]), .Z(n443) );
  NANDN U660 ( .A(n3), .B(N401), .Z(n442) );
  NAND U661 ( .A(n444), .B(n445), .Z(z3[136]) );
  NANDN U662 ( .A(N262), .B(z2[136]), .Z(n445) );
  NANDN U663 ( .A(n3), .B(N400), .Z(n444) );
  NAND U664 ( .A(n446), .B(n447), .Z(z3[135]) );
  NANDN U665 ( .A(N262), .B(z2[135]), .Z(n447) );
  NANDN U666 ( .A(n3), .B(N399), .Z(n446) );
  NAND U667 ( .A(n448), .B(n449), .Z(z3[134]) );
  NANDN U668 ( .A(N262), .B(z2[134]), .Z(n449) );
  NANDN U669 ( .A(n3), .B(N398), .Z(n448) );
  NAND U670 ( .A(n450), .B(n451), .Z(z3[133]) );
  NANDN U671 ( .A(N262), .B(z2[133]), .Z(n451) );
  NANDN U672 ( .A(n3), .B(N397), .Z(n450) );
  NAND U673 ( .A(n452), .B(n453), .Z(z3[132]) );
  NANDN U674 ( .A(N262), .B(z2[132]), .Z(n453) );
  NANDN U675 ( .A(n3), .B(N396), .Z(n452) );
  NAND U676 ( .A(n454), .B(n455), .Z(z3[131]) );
  NANDN U677 ( .A(N262), .B(z2[131]), .Z(n455) );
  NANDN U678 ( .A(n3), .B(N395), .Z(n454) );
  NAND U679 ( .A(n456), .B(n457), .Z(z3[130]) );
  NANDN U680 ( .A(N262), .B(z2[130]), .Z(n457) );
  NANDN U681 ( .A(n3), .B(N394), .Z(n456) );
  NAND U682 ( .A(n458), .B(n459), .Z(z3[12]) );
  NANDN U683 ( .A(N262), .B(z2[12]), .Z(n459) );
  NANDN U684 ( .A(n3), .B(N276), .Z(n458) );
  NAND U685 ( .A(n460), .B(n461), .Z(z3[129]) );
  NANDN U686 ( .A(N262), .B(z2[129]), .Z(n461) );
  NANDN U687 ( .A(n3), .B(N393), .Z(n460) );
  NAND U688 ( .A(n462), .B(n463), .Z(z3[128]) );
  NANDN U689 ( .A(N262), .B(z2[128]), .Z(n463) );
  NANDN U690 ( .A(n3), .B(N392), .Z(n462) );
  NAND U691 ( .A(n464), .B(n465), .Z(z3[127]) );
  NANDN U692 ( .A(N262), .B(z2[127]), .Z(n465) );
  NANDN U693 ( .A(n3), .B(N391), .Z(n464) );
  NAND U694 ( .A(n466), .B(n467), .Z(z3[126]) );
  NANDN U695 ( .A(N262), .B(z2[126]), .Z(n467) );
  NANDN U696 ( .A(n3), .B(N390), .Z(n466) );
  NAND U697 ( .A(n468), .B(n469), .Z(z3[125]) );
  NANDN U698 ( .A(N262), .B(z2[125]), .Z(n469) );
  NANDN U699 ( .A(n3), .B(N389), .Z(n468) );
  NAND U700 ( .A(n470), .B(n471), .Z(z3[124]) );
  NANDN U701 ( .A(N262), .B(z2[124]), .Z(n471) );
  NANDN U702 ( .A(n3), .B(N388), .Z(n470) );
  NAND U703 ( .A(n472), .B(n473), .Z(z3[123]) );
  NANDN U704 ( .A(N262), .B(z2[123]), .Z(n473) );
  NANDN U705 ( .A(n3), .B(N387), .Z(n472) );
  NAND U706 ( .A(n474), .B(n475), .Z(z3[122]) );
  NANDN U707 ( .A(N262), .B(z2[122]), .Z(n475) );
  NANDN U708 ( .A(n3), .B(N386), .Z(n474) );
  NAND U709 ( .A(n476), .B(n477), .Z(z3[121]) );
  NANDN U710 ( .A(N262), .B(z2[121]), .Z(n477) );
  NANDN U711 ( .A(n3), .B(N385), .Z(n476) );
  NAND U712 ( .A(n478), .B(n479), .Z(z3[120]) );
  NANDN U713 ( .A(N262), .B(z2[120]), .Z(n479) );
  NANDN U714 ( .A(n3), .B(N384), .Z(n478) );
  NAND U715 ( .A(n480), .B(n481), .Z(z3[11]) );
  NANDN U716 ( .A(N262), .B(z2[11]), .Z(n481) );
  NANDN U717 ( .A(n3), .B(N275), .Z(n480) );
  NAND U718 ( .A(n482), .B(n483), .Z(z3[119]) );
  NANDN U719 ( .A(N262), .B(z2[119]), .Z(n483) );
  NANDN U720 ( .A(n3), .B(N383), .Z(n482) );
  NAND U721 ( .A(n484), .B(n485), .Z(z3[118]) );
  NANDN U722 ( .A(N262), .B(z2[118]), .Z(n485) );
  NANDN U723 ( .A(n3), .B(N382), .Z(n484) );
  NAND U724 ( .A(n486), .B(n487), .Z(z3[117]) );
  NANDN U725 ( .A(N262), .B(z2[117]), .Z(n487) );
  NANDN U726 ( .A(n3), .B(N381), .Z(n486) );
  NAND U727 ( .A(n488), .B(n489), .Z(z3[116]) );
  NANDN U728 ( .A(N262), .B(z2[116]), .Z(n489) );
  NANDN U729 ( .A(n3), .B(N380), .Z(n488) );
  NAND U730 ( .A(n490), .B(n491), .Z(z3[115]) );
  NANDN U731 ( .A(N262), .B(z2[115]), .Z(n491) );
  NANDN U732 ( .A(n3), .B(N379), .Z(n490) );
  NAND U733 ( .A(n492), .B(n493), .Z(z3[114]) );
  NANDN U734 ( .A(N262), .B(z2[114]), .Z(n493) );
  NANDN U735 ( .A(n3), .B(N378), .Z(n492) );
  NAND U736 ( .A(n494), .B(n495), .Z(z3[113]) );
  NANDN U737 ( .A(N262), .B(z2[113]), .Z(n495) );
  NANDN U738 ( .A(n3), .B(N377), .Z(n494) );
  NAND U739 ( .A(n496), .B(n497), .Z(z3[112]) );
  NANDN U740 ( .A(N262), .B(z2[112]), .Z(n497) );
  NANDN U741 ( .A(n3), .B(N376), .Z(n496) );
  NAND U742 ( .A(n498), .B(n499), .Z(z3[111]) );
  NANDN U743 ( .A(N262), .B(z2[111]), .Z(n499) );
  NANDN U744 ( .A(n3), .B(N375), .Z(n498) );
  NAND U745 ( .A(n500), .B(n501), .Z(z3[110]) );
  NANDN U746 ( .A(N262), .B(z2[110]), .Z(n501) );
  NANDN U747 ( .A(n3), .B(N374), .Z(n500) );
  NAND U748 ( .A(n502), .B(n503), .Z(z3[10]) );
  NANDN U749 ( .A(N262), .B(z2[10]), .Z(n503) );
  NANDN U750 ( .A(n3), .B(N274), .Z(n502) );
  NAND U751 ( .A(n504), .B(n505), .Z(z3[109]) );
  NANDN U752 ( .A(N262), .B(z2[109]), .Z(n505) );
  NANDN U753 ( .A(n3), .B(N373), .Z(n504) );
  NAND U754 ( .A(n506), .B(n507), .Z(z3[108]) );
  NANDN U755 ( .A(N262), .B(z2[108]), .Z(n507) );
  NANDN U756 ( .A(n3), .B(N372), .Z(n506) );
  NAND U757 ( .A(n508), .B(n509), .Z(z3[107]) );
  NANDN U758 ( .A(N262), .B(z2[107]), .Z(n509) );
  NANDN U759 ( .A(n3), .B(N371), .Z(n508) );
  NAND U760 ( .A(n510), .B(n511), .Z(z3[106]) );
  NANDN U761 ( .A(N262), .B(z2[106]), .Z(n511) );
  NANDN U762 ( .A(n3), .B(N370), .Z(n510) );
  NAND U763 ( .A(n512), .B(n513), .Z(z3[105]) );
  NANDN U764 ( .A(N262), .B(z2[105]), .Z(n513) );
  NANDN U765 ( .A(n3), .B(N369), .Z(n512) );
  NAND U766 ( .A(n514), .B(n515), .Z(z3[104]) );
  NANDN U767 ( .A(N262), .B(z2[104]), .Z(n515) );
  NANDN U768 ( .A(n3), .B(N368), .Z(n514) );
  NAND U769 ( .A(n516), .B(n517), .Z(z3[103]) );
  NANDN U770 ( .A(N262), .B(z2[103]), .Z(n517) );
  NANDN U771 ( .A(n3), .B(N367), .Z(n516) );
  NAND U772 ( .A(n518), .B(n519), .Z(z3[102]) );
  NANDN U773 ( .A(N262), .B(z2[102]), .Z(n519) );
  NANDN U774 ( .A(n3), .B(N366), .Z(n518) );
  NAND U775 ( .A(n520), .B(n521), .Z(z3[101]) );
  NANDN U776 ( .A(N262), .B(z2[101]), .Z(n521) );
  NANDN U777 ( .A(n3), .B(N365), .Z(n520) );
  NAND U778 ( .A(n522), .B(n523), .Z(z3[100]) );
  NANDN U779 ( .A(N262), .B(z2[100]), .Z(n523) );
  NANDN U780 ( .A(n3), .B(N364), .Z(n522) );
  NAND U781 ( .A(n524), .B(n525), .Z(z3[0]) );
  NANDN U782 ( .A(N262), .B(z2[0]), .Z(n525) );
  NANDN U783 ( .A(n3), .B(N264), .Z(n524) );
  IV U784 ( .A(N262), .Z(n3) );
  NAND U785 ( .A(n526), .B(n527), .Z(z2[9]) );
  NANDN U786 ( .A(xregN_1), .B(zin[8]), .Z(n527) );
  NAND U787 ( .A(N13), .B(xregN_1), .Z(n526) );
  NAND U788 ( .A(n528), .B(n529), .Z(z2[99]) );
  NANDN U789 ( .A(xregN_1), .B(zin[98]), .Z(n529) );
  NAND U790 ( .A(N103), .B(xregN_1), .Z(n528) );
  NAND U791 ( .A(n530), .B(n531), .Z(z2[98]) );
  NANDN U792 ( .A(xregN_1), .B(zin[97]), .Z(n531) );
  NAND U793 ( .A(N102), .B(xregN_1), .Z(n530) );
  NAND U794 ( .A(n532), .B(n533), .Z(z2[97]) );
  NANDN U795 ( .A(xregN_1), .B(zin[96]), .Z(n533) );
  NAND U796 ( .A(N101), .B(xregN_1), .Z(n532) );
  NAND U797 ( .A(n534), .B(n535), .Z(z2[96]) );
  NANDN U798 ( .A(xregN_1), .B(zin[95]), .Z(n535) );
  NAND U799 ( .A(N100), .B(xregN_1), .Z(n534) );
  NAND U800 ( .A(n536), .B(n537), .Z(z2[95]) );
  NANDN U801 ( .A(xregN_1), .B(zin[94]), .Z(n537) );
  NAND U802 ( .A(N99), .B(xregN_1), .Z(n536) );
  NAND U803 ( .A(n538), .B(n539), .Z(z2[94]) );
  NANDN U804 ( .A(xregN_1), .B(zin[93]), .Z(n539) );
  NAND U805 ( .A(N98), .B(xregN_1), .Z(n538) );
  NAND U806 ( .A(n540), .B(n541), .Z(z2[93]) );
  NANDN U807 ( .A(xregN_1), .B(zin[92]), .Z(n541) );
  NAND U808 ( .A(N97), .B(xregN_1), .Z(n540) );
  NAND U809 ( .A(n542), .B(n543), .Z(z2[92]) );
  NANDN U810 ( .A(xregN_1), .B(zin[91]), .Z(n543) );
  NAND U811 ( .A(N96), .B(xregN_1), .Z(n542) );
  NAND U812 ( .A(n544), .B(n545), .Z(z2[91]) );
  NANDN U813 ( .A(xregN_1), .B(zin[90]), .Z(n545) );
  NAND U814 ( .A(N95), .B(xregN_1), .Z(n544) );
  NAND U815 ( .A(n546), .B(n547), .Z(z2[90]) );
  NANDN U816 ( .A(xregN_1), .B(zin[89]), .Z(n547) );
  NAND U817 ( .A(N94), .B(xregN_1), .Z(n546) );
  NAND U818 ( .A(n548), .B(n549), .Z(z2[8]) );
  NANDN U819 ( .A(xregN_1), .B(zin[7]), .Z(n549) );
  NAND U820 ( .A(N12), .B(xregN_1), .Z(n548) );
  NAND U821 ( .A(n550), .B(n551), .Z(z2[89]) );
  NANDN U822 ( .A(xregN_1), .B(zin[88]), .Z(n551) );
  NAND U823 ( .A(N93), .B(xregN_1), .Z(n550) );
  NAND U824 ( .A(n552), .B(n553), .Z(z2[88]) );
  NANDN U825 ( .A(xregN_1), .B(zin[87]), .Z(n553) );
  NAND U826 ( .A(N92), .B(xregN_1), .Z(n552) );
  NAND U827 ( .A(n554), .B(n555), .Z(z2[87]) );
  NANDN U828 ( .A(xregN_1), .B(zin[86]), .Z(n555) );
  NAND U829 ( .A(N91), .B(xregN_1), .Z(n554) );
  NAND U830 ( .A(n556), .B(n557), .Z(z2[86]) );
  NANDN U831 ( .A(xregN_1), .B(zin[85]), .Z(n557) );
  NAND U832 ( .A(N90), .B(xregN_1), .Z(n556) );
  NAND U833 ( .A(n558), .B(n559), .Z(z2[85]) );
  NANDN U834 ( .A(xregN_1), .B(zin[84]), .Z(n559) );
  NAND U835 ( .A(N89), .B(xregN_1), .Z(n558) );
  NAND U836 ( .A(n560), .B(n561), .Z(z2[84]) );
  NANDN U837 ( .A(xregN_1), .B(zin[83]), .Z(n561) );
  NAND U838 ( .A(N88), .B(xregN_1), .Z(n560) );
  NAND U839 ( .A(n562), .B(n563), .Z(z2[83]) );
  NANDN U840 ( .A(xregN_1), .B(zin[82]), .Z(n563) );
  NAND U841 ( .A(N87), .B(xregN_1), .Z(n562) );
  NAND U842 ( .A(n564), .B(n565), .Z(z2[82]) );
  NANDN U843 ( .A(xregN_1), .B(zin[81]), .Z(n565) );
  NAND U844 ( .A(N86), .B(xregN_1), .Z(n564) );
  NAND U845 ( .A(n566), .B(n567), .Z(z2[81]) );
  NANDN U846 ( .A(xregN_1), .B(zin[80]), .Z(n567) );
  NAND U847 ( .A(N85), .B(xregN_1), .Z(n566) );
  NAND U848 ( .A(n568), .B(n569), .Z(z2[80]) );
  NANDN U849 ( .A(xregN_1), .B(zin[79]), .Z(n569) );
  NAND U850 ( .A(N84), .B(xregN_1), .Z(n568) );
  NAND U851 ( .A(n570), .B(n571), .Z(z2[7]) );
  NANDN U852 ( .A(xregN_1), .B(zin[6]), .Z(n571) );
  NAND U853 ( .A(N11), .B(xregN_1), .Z(n570) );
  NAND U854 ( .A(n572), .B(n573), .Z(z2[79]) );
  NANDN U855 ( .A(xregN_1), .B(zin[78]), .Z(n573) );
  NAND U856 ( .A(N83), .B(xregN_1), .Z(n572) );
  NAND U857 ( .A(n574), .B(n575), .Z(z2[78]) );
  NANDN U858 ( .A(xregN_1), .B(zin[77]), .Z(n575) );
  NAND U859 ( .A(N82), .B(xregN_1), .Z(n574) );
  NAND U860 ( .A(n576), .B(n577), .Z(z2[77]) );
  NANDN U861 ( .A(xregN_1), .B(zin[76]), .Z(n577) );
  NAND U862 ( .A(N81), .B(xregN_1), .Z(n576) );
  NAND U863 ( .A(n578), .B(n579), .Z(z2[76]) );
  NANDN U864 ( .A(xregN_1), .B(zin[75]), .Z(n579) );
  NAND U865 ( .A(N80), .B(xregN_1), .Z(n578) );
  NAND U866 ( .A(n580), .B(n581), .Z(z2[75]) );
  NANDN U867 ( .A(xregN_1), .B(zin[74]), .Z(n581) );
  NAND U868 ( .A(N79), .B(xregN_1), .Z(n580) );
  NAND U869 ( .A(n582), .B(n583), .Z(z2[74]) );
  NANDN U870 ( .A(xregN_1), .B(zin[73]), .Z(n583) );
  NAND U871 ( .A(N78), .B(xregN_1), .Z(n582) );
  NAND U872 ( .A(n584), .B(n585), .Z(z2[73]) );
  NANDN U873 ( .A(xregN_1), .B(zin[72]), .Z(n585) );
  NAND U874 ( .A(N77), .B(xregN_1), .Z(n584) );
  NAND U875 ( .A(n586), .B(n587), .Z(z2[72]) );
  NANDN U876 ( .A(xregN_1), .B(zin[71]), .Z(n587) );
  NAND U877 ( .A(N76), .B(xregN_1), .Z(n586) );
  NAND U878 ( .A(n588), .B(n589), .Z(z2[71]) );
  NANDN U879 ( .A(xregN_1), .B(zin[70]), .Z(n589) );
  NAND U880 ( .A(N75), .B(xregN_1), .Z(n588) );
  NAND U881 ( .A(n590), .B(n591), .Z(z2[70]) );
  NANDN U882 ( .A(xregN_1), .B(zin[69]), .Z(n591) );
  NAND U883 ( .A(N74), .B(xregN_1), .Z(n590) );
  NAND U884 ( .A(n592), .B(n593), .Z(z2[6]) );
  NANDN U885 ( .A(xregN_1), .B(zin[5]), .Z(n593) );
  NAND U886 ( .A(N10), .B(xregN_1), .Z(n592) );
  NAND U887 ( .A(n594), .B(n595), .Z(z2[69]) );
  NANDN U888 ( .A(xregN_1), .B(zin[68]), .Z(n595) );
  NAND U889 ( .A(N73), .B(xregN_1), .Z(n594) );
  NAND U890 ( .A(n596), .B(n597), .Z(z2[68]) );
  NANDN U891 ( .A(xregN_1), .B(zin[67]), .Z(n597) );
  NAND U892 ( .A(N72), .B(xregN_1), .Z(n596) );
  NAND U893 ( .A(n598), .B(n599), .Z(z2[67]) );
  NANDN U894 ( .A(xregN_1), .B(zin[66]), .Z(n599) );
  NAND U895 ( .A(N71), .B(xregN_1), .Z(n598) );
  NAND U896 ( .A(n600), .B(n601), .Z(z2[66]) );
  NANDN U897 ( .A(xregN_1), .B(zin[65]), .Z(n601) );
  NAND U898 ( .A(N70), .B(xregN_1), .Z(n600) );
  NAND U899 ( .A(n602), .B(n603), .Z(z2[65]) );
  NANDN U900 ( .A(xregN_1), .B(zin[64]), .Z(n603) );
  NAND U901 ( .A(N69), .B(xregN_1), .Z(n602) );
  NAND U902 ( .A(n604), .B(n605), .Z(z2[64]) );
  NANDN U903 ( .A(xregN_1), .B(zin[63]), .Z(n605) );
  NAND U904 ( .A(N68), .B(xregN_1), .Z(n604) );
  NAND U905 ( .A(n606), .B(n607), .Z(z2[63]) );
  NANDN U906 ( .A(xregN_1), .B(zin[62]), .Z(n607) );
  NAND U907 ( .A(N67), .B(xregN_1), .Z(n606) );
  NAND U908 ( .A(n608), .B(n609), .Z(z2[62]) );
  NANDN U909 ( .A(xregN_1), .B(zin[61]), .Z(n609) );
  NAND U910 ( .A(N66), .B(xregN_1), .Z(n608) );
  NAND U911 ( .A(n610), .B(n611), .Z(z2[61]) );
  NANDN U912 ( .A(xregN_1), .B(zin[60]), .Z(n611) );
  NAND U913 ( .A(N65), .B(xregN_1), .Z(n610) );
  NAND U914 ( .A(n612), .B(n613), .Z(z2[60]) );
  NANDN U915 ( .A(xregN_1), .B(zin[59]), .Z(n613) );
  NAND U916 ( .A(N64), .B(xregN_1), .Z(n612) );
  NAND U917 ( .A(n614), .B(n615), .Z(z2[5]) );
  NANDN U918 ( .A(xregN_1), .B(zin[4]), .Z(n615) );
  NAND U919 ( .A(N9), .B(xregN_1), .Z(n614) );
  NAND U920 ( .A(n616), .B(n617), .Z(z2[59]) );
  NANDN U921 ( .A(xregN_1), .B(zin[58]), .Z(n617) );
  NAND U922 ( .A(N63), .B(xregN_1), .Z(n616) );
  NAND U923 ( .A(n618), .B(n619), .Z(z2[58]) );
  NANDN U924 ( .A(xregN_1), .B(zin[57]), .Z(n619) );
  NAND U925 ( .A(N62), .B(xregN_1), .Z(n618) );
  NAND U926 ( .A(n620), .B(n621), .Z(z2[57]) );
  NANDN U927 ( .A(xregN_1), .B(zin[56]), .Z(n621) );
  NAND U928 ( .A(N61), .B(xregN_1), .Z(n620) );
  NAND U929 ( .A(n622), .B(n623), .Z(z2[56]) );
  NANDN U930 ( .A(xregN_1), .B(zin[55]), .Z(n623) );
  NAND U931 ( .A(N60), .B(xregN_1), .Z(n622) );
  NAND U932 ( .A(n624), .B(n625), .Z(z2[55]) );
  NANDN U933 ( .A(xregN_1), .B(zin[54]), .Z(n625) );
  NAND U934 ( .A(N59), .B(xregN_1), .Z(n624) );
  NAND U935 ( .A(n626), .B(n627), .Z(z2[54]) );
  NANDN U936 ( .A(xregN_1), .B(zin[53]), .Z(n627) );
  NAND U937 ( .A(N58), .B(xregN_1), .Z(n626) );
  NAND U938 ( .A(n628), .B(n629), .Z(z2[53]) );
  NANDN U939 ( .A(xregN_1), .B(zin[52]), .Z(n629) );
  NAND U940 ( .A(N57), .B(xregN_1), .Z(n628) );
  NAND U941 ( .A(n630), .B(n631), .Z(z2[52]) );
  NANDN U942 ( .A(xregN_1), .B(zin[51]), .Z(n631) );
  NAND U943 ( .A(N56), .B(xregN_1), .Z(n630) );
  NAND U944 ( .A(n632), .B(n633), .Z(z2[51]) );
  NANDN U945 ( .A(xregN_1), .B(zin[50]), .Z(n633) );
  NAND U946 ( .A(N55), .B(xregN_1), .Z(n632) );
  NAND U947 ( .A(n634), .B(n635), .Z(z2[50]) );
  NANDN U948 ( .A(xregN_1), .B(zin[49]), .Z(n635) );
  NAND U949 ( .A(N54), .B(xregN_1), .Z(n634) );
  NAND U950 ( .A(n636), .B(n637), .Z(z2[4]) );
  NANDN U951 ( .A(xregN_1), .B(zin[3]), .Z(n637) );
  NAND U952 ( .A(N8), .B(xregN_1), .Z(n636) );
  NAND U953 ( .A(n638), .B(n639), .Z(z2[49]) );
  NANDN U954 ( .A(xregN_1), .B(zin[48]), .Z(n639) );
  NAND U955 ( .A(N53), .B(xregN_1), .Z(n638) );
  NAND U956 ( .A(n640), .B(n641), .Z(z2[48]) );
  NANDN U957 ( .A(xregN_1), .B(zin[47]), .Z(n641) );
  NAND U958 ( .A(N52), .B(xregN_1), .Z(n640) );
  NAND U959 ( .A(n642), .B(n643), .Z(z2[47]) );
  NANDN U960 ( .A(xregN_1), .B(zin[46]), .Z(n643) );
  NAND U961 ( .A(N51), .B(xregN_1), .Z(n642) );
  NAND U962 ( .A(n644), .B(n645), .Z(z2[46]) );
  NANDN U963 ( .A(xregN_1), .B(zin[45]), .Z(n645) );
  NAND U964 ( .A(N50), .B(xregN_1), .Z(n644) );
  NAND U965 ( .A(n646), .B(n647), .Z(z2[45]) );
  NANDN U966 ( .A(xregN_1), .B(zin[44]), .Z(n647) );
  NAND U967 ( .A(N49), .B(xregN_1), .Z(n646) );
  NAND U968 ( .A(n648), .B(n649), .Z(z2[44]) );
  NANDN U969 ( .A(xregN_1), .B(zin[43]), .Z(n649) );
  NAND U970 ( .A(N48), .B(xregN_1), .Z(n648) );
  NAND U971 ( .A(n650), .B(n651), .Z(z2[43]) );
  NANDN U972 ( .A(xregN_1), .B(zin[42]), .Z(n651) );
  NAND U973 ( .A(N47), .B(xregN_1), .Z(n650) );
  NAND U974 ( .A(n652), .B(n653), .Z(z2[42]) );
  NANDN U975 ( .A(xregN_1), .B(zin[41]), .Z(n653) );
  NAND U976 ( .A(N46), .B(xregN_1), .Z(n652) );
  NAND U977 ( .A(n654), .B(n655), .Z(z2[41]) );
  NANDN U978 ( .A(xregN_1), .B(zin[40]), .Z(n655) );
  NAND U979 ( .A(N45), .B(xregN_1), .Z(n654) );
  NAND U980 ( .A(n656), .B(n657), .Z(z2[40]) );
  NANDN U981 ( .A(xregN_1), .B(zin[39]), .Z(n657) );
  NAND U982 ( .A(N44), .B(xregN_1), .Z(n656) );
  NAND U983 ( .A(n658), .B(n659), .Z(z2[3]) );
  NANDN U984 ( .A(xregN_1), .B(zin[2]), .Z(n659) );
  NAND U985 ( .A(N7), .B(xregN_1), .Z(n658) );
  NAND U986 ( .A(n660), .B(n661), .Z(z2[39]) );
  NANDN U987 ( .A(xregN_1), .B(zin[38]), .Z(n661) );
  NAND U988 ( .A(N43), .B(xregN_1), .Z(n660) );
  NAND U989 ( .A(n662), .B(n663), .Z(z2[38]) );
  NANDN U990 ( .A(xregN_1), .B(zin[37]), .Z(n663) );
  NAND U991 ( .A(N42), .B(xregN_1), .Z(n662) );
  NAND U992 ( .A(n664), .B(n665), .Z(z2[37]) );
  NANDN U993 ( .A(xregN_1), .B(zin[36]), .Z(n665) );
  NAND U994 ( .A(N41), .B(xregN_1), .Z(n664) );
  NAND U995 ( .A(n666), .B(n667), .Z(z2[36]) );
  NANDN U996 ( .A(xregN_1), .B(zin[35]), .Z(n667) );
  NAND U997 ( .A(N40), .B(xregN_1), .Z(n666) );
  NAND U998 ( .A(n668), .B(n669), .Z(z2[35]) );
  NANDN U999 ( .A(xregN_1), .B(zin[34]), .Z(n669) );
  NAND U1000 ( .A(N39), .B(xregN_1), .Z(n668) );
  NAND U1001 ( .A(n670), .B(n671), .Z(z2[34]) );
  NANDN U1002 ( .A(xregN_1), .B(zin[33]), .Z(n671) );
  NAND U1003 ( .A(N38), .B(xregN_1), .Z(n670) );
  NAND U1004 ( .A(n672), .B(n673), .Z(z2[33]) );
  NANDN U1005 ( .A(xregN_1), .B(zin[32]), .Z(n673) );
  NAND U1006 ( .A(N37), .B(xregN_1), .Z(n672) );
  NAND U1007 ( .A(n674), .B(n675), .Z(z2[32]) );
  NANDN U1008 ( .A(xregN_1), .B(zin[31]), .Z(n675) );
  NAND U1009 ( .A(N36), .B(xregN_1), .Z(n674) );
  NAND U1010 ( .A(n676), .B(n677), .Z(z2[31]) );
  NANDN U1011 ( .A(xregN_1), .B(zin[30]), .Z(n677) );
  NAND U1012 ( .A(N35), .B(xregN_1), .Z(n676) );
  NAND U1013 ( .A(n678), .B(n679), .Z(z2[30]) );
  NANDN U1014 ( .A(xregN_1), .B(zin[29]), .Z(n679) );
  NAND U1015 ( .A(N34), .B(xregN_1), .Z(n678) );
  NAND U1016 ( .A(n680), .B(n681), .Z(z2[2]) );
  NANDN U1017 ( .A(xregN_1), .B(zin[1]), .Z(n681) );
  NAND U1018 ( .A(N6), .B(xregN_1), .Z(n680) );
  NAND U1019 ( .A(n682), .B(n683), .Z(z2[29]) );
  NANDN U1020 ( .A(xregN_1), .B(zin[28]), .Z(n683) );
  NAND U1021 ( .A(N33), .B(xregN_1), .Z(n682) );
  NAND U1022 ( .A(n684), .B(n685), .Z(z2[28]) );
  NANDN U1023 ( .A(xregN_1), .B(zin[27]), .Z(n685) );
  NAND U1024 ( .A(N32), .B(xregN_1), .Z(n684) );
  NAND U1025 ( .A(n686), .B(n687), .Z(z2[27]) );
  NANDN U1026 ( .A(xregN_1), .B(zin[26]), .Z(n687) );
  NAND U1027 ( .A(N31), .B(xregN_1), .Z(n686) );
  NAND U1028 ( .A(n688), .B(n689), .Z(z2[26]) );
  NANDN U1029 ( .A(xregN_1), .B(zin[25]), .Z(n689) );
  NAND U1030 ( .A(N30), .B(xregN_1), .Z(n688) );
  NAND U1031 ( .A(n690), .B(n691), .Z(z2[25]) );
  NANDN U1032 ( .A(xregN_1), .B(zin[24]), .Z(n691) );
  NAND U1033 ( .A(N29), .B(xregN_1), .Z(n690) );
  NAND U1034 ( .A(n692), .B(n693), .Z(z2[257]) );
  NANDN U1035 ( .A(xregN_1), .B(zin[256]), .Z(n693) );
  NAND U1036 ( .A(N261), .B(xregN_1), .Z(n692) );
  NAND U1037 ( .A(n694), .B(n695), .Z(z2[256]) );
  NANDN U1038 ( .A(xregN_1), .B(zin[255]), .Z(n695) );
  NAND U1039 ( .A(N260), .B(xregN_1), .Z(n694) );
  NAND U1040 ( .A(n696), .B(n697), .Z(z2[255]) );
  NANDN U1041 ( .A(xregN_1), .B(zin[254]), .Z(n697) );
  NAND U1042 ( .A(N259), .B(xregN_1), .Z(n696) );
  NAND U1043 ( .A(n698), .B(n699), .Z(z2[254]) );
  NANDN U1044 ( .A(xregN_1), .B(zin[253]), .Z(n699) );
  NAND U1045 ( .A(N258), .B(xregN_1), .Z(n698) );
  NAND U1046 ( .A(n700), .B(n701), .Z(z2[253]) );
  NANDN U1047 ( .A(xregN_1), .B(zin[252]), .Z(n701) );
  NAND U1048 ( .A(N257), .B(xregN_1), .Z(n700) );
  NAND U1049 ( .A(n702), .B(n703), .Z(z2[252]) );
  NANDN U1050 ( .A(xregN_1), .B(zin[251]), .Z(n703) );
  NAND U1051 ( .A(N256), .B(xregN_1), .Z(n702) );
  NAND U1052 ( .A(n704), .B(n705), .Z(z2[251]) );
  NANDN U1053 ( .A(xregN_1), .B(zin[250]), .Z(n705) );
  NAND U1054 ( .A(N255), .B(xregN_1), .Z(n704) );
  NAND U1055 ( .A(n706), .B(n707), .Z(z2[250]) );
  NANDN U1056 ( .A(xregN_1), .B(zin[249]), .Z(n707) );
  NAND U1057 ( .A(N254), .B(xregN_1), .Z(n706) );
  NAND U1058 ( .A(n708), .B(n709), .Z(z2[24]) );
  NANDN U1059 ( .A(xregN_1), .B(zin[23]), .Z(n709) );
  NAND U1060 ( .A(N28), .B(xregN_1), .Z(n708) );
  NAND U1061 ( .A(n710), .B(n711), .Z(z2[249]) );
  NANDN U1062 ( .A(xregN_1), .B(zin[248]), .Z(n711) );
  NAND U1063 ( .A(N253), .B(xregN_1), .Z(n710) );
  NAND U1064 ( .A(n712), .B(n713), .Z(z2[248]) );
  NANDN U1065 ( .A(xregN_1), .B(zin[247]), .Z(n713) );
  NAND U1066 ( .A(N252), .B(xregN_1), .Z(n712) );
  NAND U1067 ( .A(n714), .B(n715), .Z(z2[247]) );
  NANDN U1068 ( .A(xregN_1), .B(zin[246]), .Z(n715) );
  NAND U1069 ( .A(N251), .B(xregN_1), .Z(n714) );
  NAND U1070 ( .A(n716), .B(n717), .Z(z2[246]) );
  NANDN U1071 ( .A(xregN_1), .B(zin[245]), .Z(n717) );
  NAND U1072 ( .A(N250), .B(xregN_1), .Z(n716) );
  NAND U1073 ( .A(n718), .B(n719), .Z(z2[245]) );
  NANDN U1074 ( .A(xregN_1), .B(zin[244]), .Z(n719) );
  NAND U1075 ( .A(N249), .B(xregN_1), .Z(n718) );
  NAND U1076 ( .A(n720), .B(n721), .Z(z2[244]) );
  NANDN U1077 ( .A(xregN_1), .B(zin[243]), .Z(n721) );
  NAND U1078 ( .A(N248), .B(xregN_1), .Z(n720) );
  NAND U1079 ( .A(n722), .B(n723), .Z(z2[243]) );
  NANDN U1080 ( .A(xregN_1), .B(zin[242]), .Z(n723) );
  NAND U1081 ( .A(N247), .B(xregN_1), .Z(n722) );
  NAND U1082 ( .A(n724), .B(n725), .Z(z2[242]) );
  NANDN U1083 ( .A(xregN_1), .B(zin[241]), .Z(n725) );
  NAND U1084 ( .A(N246), .B(xregN_1), .Z(n724) );
  NAND U1085 ( .A(n726), .B(n727), .Z(z2[241]) );
  NANDN U1086 ( .A(xregN_1), .B(zin[240]), .Z(n727) );
  NAND U1087 ( .A(N245), .B(xregN_1), .Z(n726) );
  NAND U1088 ( .A(n728), .B(n729), .Z(z2[240]) );
  NANDN U1089 ( .A(xregN_1), .B(zin[239]), .Z(n729) );
  NAND U1090 ( .A(N244), .B(xregN_1), .Z(n728) );
  NAND U1091 ( .A(n730), .B(n731), .Z(z2[23]) );
  NANDN U1092 ( .A(xregN_1), .B(zin[22]), .Z(n731) );
  NAND U1093 ( .A(N27), .B(xregN_1), .Z(n730) );
  NAND U1094 ( .A(n732), .B(n733), .Z(z2[239]) );
  NANDN U1095 ( .A(xregN_1), .B(zin[238]), .Z(n733) );
  NAND U1096 ( .A(N243), .B(xregN_1), .Z(n732) );
  NAND U1097 ( .A(n734), .B(n735), .Z(z2[238]) );
  NANDN U1098 ( .A(xregN_1), .B(zin[237]), .Z(n735) );
  NAND U1099 ( .A(N242), .B(xregN_1), .Z(n734) );
  NAND U1100 ( .A(n736), .B(n737), .Z(z2[237]) );
  NANDN U1101 ( .A(xregN_1), .B(zin[236]), .Z(n737) );
  NAND U1102 ( .A(N241), .B(xregN_1), .Z(n736) );
  NAND U1103 ( .A(n738), .B(n739), .Z(z2[236]) );
  NANDN U1104 ( .A(xregN_1), .B(zin[235]), .Z(n739) );
  NAND U1105 ( .A(N240), .B(xregN_1), .Z(n738) );
  NAND U1106 ( .A(n740), .B(n741), .Z(z2[235]) );
  NANDN U1107 ( .A(xregN_1), .B(zin[234]), .Z(n741) );
  NAND U1108 ( .A(N239), .B(xregN_1), .Z(n740) );
  NAND U1109 ( .A(n742), .B(n743), .Z(z2[234]) );
  NANDN U1110 ( .A(xregN_1), .B(zin[233]), .Z(n743) );
  NAND U1111 ( .A(N238), .B(xregN_1), .Z(n742) );
  NAND U1112 ( .A(n744), .B(n745), .Z(z2[233]) );
  NANDN U1113 ( .A(xregN_1), .B(zin[232]), .Z(n745) );
  NAND U1114 ( .A(N237), .B(xregN_1), .Z(n744) );
  NAND U1115 ( .A(n746), .B(n747), .Z(z2[232]) );
  NANDN U1116 ( .A(xregN_1), .B(zin[231]), .Z(n747) );
  NAND U1117 ( .A(N236), .B(xregN_1), .Z(n746) );
  NAND U1118 ( .A(n748), .B(n749), .Z(z2[231]) );
  NANDN U1119 ( .A(xregN_1), .B(zin[230]), .Z(n749) );
  NAND U1120 ( .A(N235), .B(xregN_1), .Z(n748) );
  NAND U1121 ( .A(n750), .B(n751), .Z(z2[230]) );
  NANDN U1122 ( .A(xregN_1), .B(zin[229]), .Z(n751) );
  NAND U1123 ( .A(N234), .B(xregN_1), .Z(n750) );
  NAND U1124 ( .A(n752), .B(n753), .Z(z2[22]) );
  NANDN U1125 ( .A(xregN_1), .B(zin[21]), .Z(n753) );
  NAND U1126 ( .A(N26), .B(xregN_1), .Z(n752) );
  NAND U1127 ( .A(n754), .B(n755), .Z(z2[229]) );
  NANDN U1128 ( .A(xregN_1), .B(zin[228]), .Z(n755) );
  NAND U1129 ( .A(N233), .B(xregN_1), .Z(n754) );
  NAND U1130 ( .A(n756), .B(n757), .Z(z2[228]) );
  NANDN U1131 ( .A(xregN_1), .B(zin[227]), .Z(n757) );
  NAND U1132 ( .A(N232), .B(xregN_1), .Z(n756) );
  NAND U1133 ( .A(n758), .B(n759), .Z(z2[227]) );
  NANDN U1134 ( .A(xregN_1), .B(zin[226]), .Z(n759) );
  NAND U1135 ( .A(N231), .B(xregN_1), .Z(n758) );
  NAND U1136 ( .A(n760), .B(n761), .Z(z2[226]) );
  NANDN U1137 ( .A(xregN_1), .B(zin[225]), .Z(n761) );
  NAND U1138 ( .A(N230), .B(xregN_1), .Z(n760) );
  NAND U1139 ( .A(n762), .B(n763), .Z(z2[225]) );
  NANDN U1140 ( .A(xregN_1), .B(zin[224]), .Z(n763) );
  NAND U1141 ( .A(N229), .B(xregN_1), .Z(n762) );
  NAND U1142 ( .A(n764), .B(n765), .Z(z2[224]) );
  NANDN U1143 ( .A(xregN_1), .B(zin[223]), .Z(n765) );
  NAND U1144 ( .A(N228), .B(xregN_1), .Z(n764) );
  NAND U1145 ( .A(n766), .B(n767), .Z(z2[223]) );
  NANDN U1146 ( .A(xregN_1), .B(zin[222]), .Z(n767) );
  NAND U1147 ( .A(N227), .B(xregN_1), .Z(n766) );
  NAND U1148 ( .A(n768), .B(n769), .Z(z2[222]) );
  NANDN U1149 ( .A(xregN_1), .B(zin[221]), .Z(n769) );
  NAND U1150 ( .A(N226), .B(xregN_1), .Z(n768) );
  NAND U1151 ( .A(n770), .B(n771), .Z(z2[221]) );
  NANDN U1152 ( .A(xregN_1), .B(zin[220]), .Z(n771) );
  NAND U1153 ( .A(N225), .B(xregN_1), .Z(n770) );
  NAND U1154 ( .A(n772), .B(n773), .Z(z2[220]) );
  NANDN U1155 ( .A(xregN_1), .B(zin[219]), .Z(n773) );
  NAND U1156 ( .A(N224), .B(xregN_1), .Z(n772) );
  NAND U1157 ( .A(n774), .B(n775), .Z(z2[21]) );
  NANDN U1158 ( .A(xregN_1), .B(zin[20]), .Z(n775) );
  NAND U1159 ( .A(N25), .B(xregN_1), .Z(n774) );
  NAND U1160 ( .A(n776), .B(n777), .Z(z2[219]) );
  NANDN U1161 ( .A(xregN_1), .B(zin[218]), .Z(n777) );
  NAND U1162 ( .A(N223), .B(xregN_1), .Z(n776) );
  NAND U1163 ( .A(n778), .B(n779), .Z(z2[218]) );
  NANDN U1164 ( .A(xregN_1), .B(zin[217]), .Z(n779) );
  NAND U1165 ( .A(N222), .B(xregN_1), .Z(n778) );
  NAND U1166 ( .A(n780), .B(n781), .Z(z2[217]) );
  NANDN U1167 ( .A(xregN_1), .B(zin[216]), .Z(n781) );
  NAND U1168 ( .A(N221), .B(xregN_1), .Z(n780) );
  NAND U1169 ( .A(n782), .B(n783), .Z(z2[216]) );
  NANDN U1170 ( .A(xregN_1), .B(zin[215]), .Z(n783) );
  NAND U1171 ( .A(N220), .B(xregN_1), .Z(n782) );
  NAND U1172 ( .A(n784), .B(n785), .Z(z2[215]) );
  NANDN U1173 ( .A(xregN_1), .B(zin[214]), .Z(n785) );
  NAND U1174 ( .A(N219), .B(xregN_1), .Z(n784) );
  NAND U1175 ( .A(n786), .B(n787), .Z(z2[214]) );
  NANDN U1176 ( .A(xregN_1), .B(zin[213]), .Z(n787) );
  NAND U1177 ( .A(N218), .B(xregN_1), .Z(n786) );
  NAND U1178 ( .A(n788), .B(n789), .Z(z2[213]) );
  NANDN U1179 ( .A(xregN_1), .B(zin[212]), .Z(n789) );
  NAND U1180 ( .A(N217), .B(xregN_1), .Z(n788) );
  NAND U1181 ( .A(n790), .B(n791), .Z(z2[212]) );
  NANDN U1182 ( .A(xregN_1), .B(zin[211]), .Z(n791) );
  NAND U1183 ( .A(N216), .B(xregN_1), .Z(n790) );
  NAND U1184 ( .A(n792), .B(n793), .Z(z2[211]) );
  NANDN U1185 ( .A(xregN_1), .B(zin[210]), .Z(n793) );
  NAND U1186 ( .A(N215), .B(xregN_1), .Z(n792) );
  NAND U1187 ( .A(n794), .B(n795), .Z(z2[210]) );
  NANDN U1188 ( .A(xregN_1), .B(zin[209]), .Z(n795) );
  NAND U1189 ( .A(N214), .B(xregN_1), .Z(n794) );
  NAND U1190 ( .A(n796), .B(n797), .Z(z2[20]) );
  NANDN U1191 ( .A(xregN_1), .B(zin[19]), .Z(n797) );
  NAND U1192 ( .A(N24), .B(xregN_1), .Z(n796) );
  NAND U1193 ( .A(n798), .B(n799), .Z(z2[209]) );
  NANDN U1194 ( .A(xregN_1), .B(zin[208]), .Z(n799) );
  NAND U1195 ( .A(N213), .B(xregN_1), .Z(n798) );
  NAND U1196 ( .A(n800), .B(n801), .Z(z2[208]) );
  NANDN U1197 ( .A(xregN_1), .B(zin[207]), .Z(n801) );
  NAND U1198 ( .A(N212), .B(xregN_1), .Z(n800) );
  NAND U1199 ( .A(n802), .B(n803), .Z(z2[207]) );
  NANDN U1200 ( .A(xregN_1), .B(zin[206]), .Z(n803) );
  NAND U1201 ( .A(N211), .B(xregN_1), .Z(n802) );
  NAND U1202 ( .A(n804), .B(n805), .Z(z2[206]) );
  NANDN U1203 ( .A(xregN_1), .B(zin[205]), .Z(n805) );
  NAND U1204 ( .A(N210), .B(xregN_1), .Z(n804) );
  NAND U1205 ( .A(n806), .B(n807), .Z(z2[205]) );
  NANDN U1206 ( .A(xregN_1), .B(zin[204]), .Z(n807) );
  NAND U1207 ( .A(N209), .B(xregN_1), .Z(n806) );
  NAND U1208 ( .A(n808), .B(n809), .Z(z2[204]) );
  NANDN U1209 ( .A(xregN_1), .B(zin[203]), .Z(n809) );
  NAND U1210 ( .A(N208), .B(xregN_1), .Z(n808) );
  NAND U1211 ( .A(n810), .B(n811), .Z(z2[203]) );
  NANDN U1212 ( .A(xregN_1), .B(zin[202]), .Z(n811) );
  NAND U1213 ( .A(N207), .B(xregN_1), .Z(n810) );
  NAND U1214 ( .A(n812), .B(n813), .Z(z2[202]) );
  NANDN U1215 ( .A(xregN_1), .B(zin[201]), .Z(n813) );
  NAND U1216 ( .A(N206), .B(xregN_1), .Z(n812) );
  NAND U1217 ( .A(n814), .B(n815), .Z(z2[201]) );
  NANDN U1218 ( .A(xregN_1), .B(zin[200]), .Z(n815) );
  NAND U1219 ( .A(N205), .B(xregN_1), .Z(n814) );
  NAND U1220 ( .A(n816), .B(n817), .Z(z2[200]) );
  NANDN U1221 ( .A(xregN_1), .B(zin[199]), .Z(n817) );
  NAND U1222 ( .A(N204), .B(xregN_1), .Z(n816) );
  NAND U1223 ( .A(n818), .B(n819), .Z(z2[1]) );
  NANDN U1224 ( .A(xregN_1), .B(zin[0]), .Z(n819) );
  NAND U1225 ( .A(N5), .B(xregN_1), .Z(n818) );
  NAND U1226 ( .A(n820), .B(n821), .Z(z2[19]) );
  NANDN U1227 ( .A(xregN_1), .B(zin[18]), .Z(n821) );
  NAND U1228 ( .A(N23), .B(xregN_1), .Z(n820) );
  NAND U1229 ( .A(n822), .B(n823), .Z(z2[199]) );
  NANDN U1230 ( .A(xregN_1), .B(zin[198]), .Z(n823) );
  NAND U1231 ( .A(N203), .B(xregN_1), .Z(n822) );
  NAND U1232 ( .A(n824), .B(n825), .Z(z2[198]) );
  NANDN U1233 ( .A(xregN_1), .B(zin[197]), .Z(n825) );
  NAND U1234 ( .A(N202), .B(xregN_1), .Z(n824) );
  NAND U1235 ( .A(n826), .B(n827), .Z(z2[197]) );
  NANDN U1236 ( .A(xregN_1), .B(zin[196]), .Z(n827) );
  NAND U1237 ( .A(N201), .B(xregN_1), .Z(n826) );
  NAND U1238 ( .A(n828), .B(n829), .Z(z2[196]) );
  NANDN U1239 ( .A(xregN_1), .B(zin[195]), .Z(n829) );
  NAND U1240 ( .A(N200), .B(xregN_1), .Z(n828) );
  NAND U1241 ( .A(n830), .B(n831), .Z(z2[195]) );
  NANDN U1242 ( .A(xregN_1), .B(zin[194]), .Z(n831) );
  NAND U1243 ( .A(N199), .B(xregN_1), .Z(n830) );
  NAND U1244 ( .A(n832), .B(n833), .Z(z2[194]) );
  NANDN U1245 ( .A(xregN_1), .B(zin[193]), .Z(n833) );
  NAND U1246 ( .A(N198), .B(xregN_1), .Z(n832) );
  NAND U1247 ( .A(n834), .B(n835), .Z(z2[193]) );
  NANDN U1248 ( .A(xregN_1), .B(zin[192]), .Z(n835) );
  NAND U1249 ( .A(N197), .B(xregN_1), .Z(n834) );
  NAND U1250 ( .A(n836), .B(n837), .Z(z2[192]) );
  NANDN U1251 ( .A(xregN_1), .B(zin[191]), .Z(n837) );
  NAND U1252 ( .A(N196), .B(xregN_1), .Z(n836) );
  NAND U1253 ( .A(n838), .B(n839), .Z(z2[191]) );
  NANDN U1254 ( .A(xregN_1), .B(zin[190]), .Z(n839) );
  NAND U1255 ( .A(N195), .B(xregN_1), .Z(n838) );
  NAND U1256 ( .A(n840), .B(n841), .Z(z2[190]) );
  NANDN U1257 ( .A(xregN_1), .B(zin[189]), .Z(n841) );
  NAND U1258 ( .A(N194), .B(xregN_1), .Z(n840) );
  NAND U1259 ( .A(n842), .B(n843), .Z(z2[18]) );
  NANDN U1260 ( .A(xregN_1), .B(zin[17]), .Z(n843) );
  NAND U1261 ( .A(N22), .B(xregN_1), .Z(n842) );
  NAND U1262 ( .A(n844), .B(n845), .Z(z2[189]) );
  NANDN U1263 ( .A(xregN_1), .B(zin[188]), .Z(n845) );
  NAND U1264 ( .A(N193), .B(xregN_1), .Z(n844) );
  NAND U1265 ( .A(n846), .B(n847), .Z(z2[188]) );
  NANDN U1266 ( .A(xregN_1), .B(zin[187]), .Z(n847) );
  NAND U1267 ( .A(N192), .B(xregN_1), .Z(n846) );
  NAND U1268 ( .A(n848), .B(n849), .Z(z2[187]) );
  NANDN U1269 ( .A(xregN_1), .B(zin[186]), .Z(n849) );
  NAND U1270 ( .A(N191), .B(xregN_1), .Z(n848) );
  NAND U1271 ( .A(n850), .B(n851), .Z(z2[186]) );
  NANDN U1272 ( .A(xregN_1), .B(zin[185]), .Z(n851) );
  NAND U1273 ( .A(N190), .B(xregN_1), .Z(n850) );
  NAND U1274 ( .A(n852), .B(n853), .Z(z2[185]) );
  NANDN U1275 ( .A(xregN_1), .B(zin[184]), .Z(n853) );
  NAND U1276 ( .A(N189), .B(xregN_1), .Z(n852) );
  NAND U1277 ( .A(n854), .B(n855), .Z(z2[184]) );
  NANDN U1278 ( .A(xregN_1), .B(zin[183]), .Z(n855) );
  NAND U1279 ( .A(N188), .B(xregN_1), .Z(n854) );
  NAND U1280 ( .A(n856), .B(n857), .Z(z2[183]) );
  NANDN U1281 ( .A(xregN_1), .B(zin[182]), .Z(n857) );
  NAND U1282 ( .A(N187), .B(xregN_1), .Z(n856) );
  NAND U1283 ( .A(n858), .B(n859), .Z(z2[182]) );
  NANDN U1284 ( .A(xregN_1), .B(zin[181]), .Z(n859) );
  NAND U1285 ( .A(N186), .B(xregN_1), .Z(n858) );
  NAND U1286 ( .A(n860), .B(n861), .Z(z2[181]) );
  NANDN U1287 ( .A(xregN_1), .B(zin[180]), .Z(n861) );
  NAND U1288 ( .A(N185), .B(xregN_1), .Z(n860) );
  NAND U1289 ( .A(n862), .B(n863), .Z(z2[180]) );
  NANDN U1290 ( .A(xregN_1), .B(zin[179]), .Z(n863) );
  NAND U1291 ( .A(N184), .B(xregN_1), .Z(n862) );
  NAND U1292 ( .A(n864), .B(n865), .Z(z2[17]) );
  NANDN U1293 ( .A(xregN_1), .B(zin[16]), .Z(n865) );
  NAND U1294 ( .A(N21), .B(xregN_1), .Z(n864) );
  NAND U1295 ( .A(n866), .B(n867), .Z(z2[179]) );
  NANDN U1296 ( .A(xregN_1), .B(zin[178]), .Z(n867) );
  NAND U1297 ( .A(N183), .B(xregN_1), .Z(n866) );
  NAND U1298 ( .A(n868), .B(n869), .Z(z2[178]) );
  NANDN U1299 ( .A(xregN_1), .B(zin[177]), .Z(n869) );
  NAND U1300 ( .A(N182), .B(xregN_1), .Z(n868) );
  NAND U1301 ( .A(n870), .B(n871), .Z(z2[177]) );
  NANDN U1302 ( .A(xregN_1), .B(zin[176]), .Z(n871) );
  NAND U1303 ( .A(N181), .B(xregN_1), .Z(n870) );
  NAND U1304 ( .A(n872), .B(n873), .Z(z2[176]) );
  NANDN U1305 ( .A(xregN_1), .B(zin[175]), .Z(n873) );
  NAND U1306 ( .A(N180), .B(xregN_1), .Z(n872) );
  NAND U1307 ( .A(n874), .B(n875), .Z(z2[175]) );
  NANDN U1308 ( .A(xregN_1), .B(zin[174]), .Z(n875) );
  NAND U1309 ( .A(N179), .B(xregN_1), .Z(n874) );
  NAND U1310 ( .A(n876), .B(n877), .Z(z2[174]) );
  NANDN U1311 ( .A(xregN_1), .B(zin[173]), .Z(n877) );
  NAND U1312 ( .A(N178), .B(xregN_1), .Z(n876) );
  NAND U1313 ( .A(n878), .B(n879), .Z(z2[173]) );
  NANDN U1314 ( .A(xregN_1), .B(zin[172]), .Z(n879) );
  NAND U1315 ( .A(N177), .B(xregN_1), .Z(n878) );
  NAND U1316 ( .A(n880), .B(n881), .Z(z2[172]) );
  NANDN U1317 ( .A(xregN_1), .B(zin[171]), .Z(n881) );
  NAND U1318 ( .A(N176), .B(xregN_1), .Z(n880) );
  NAND U1319 ( .A(n882), .B(n883), .Z(z2[171]) );
  NANDN U1320 ( .A(xregN_1), .B(zin[170]), .Z(n883) );
  NAND U1321 ( .A(N175), .B(xregN_1), .Z(n882) );
  NAND U1322 ( .A(n884), .B(n885), .Z(z2[170]) );
  NANDN U1323 ( .A(xregN_1), .B(zin[169]), .Z(n885) );
  NAND U1324 ( .A(N174), .B(xregN_1), .Z(n884) );
  NAND U1325 ( .A(n886), .B(n887), .Z(z2[16]) );
  NANDN U1326 ( .A(xregN_1), .B(zin[15]), .Z(n887) );
  NAND U1327 ( .A(N20), .B(xregN_1), .Z(n886) );
  NAND U1328 ( .A(n888), .B(n889), .Z(z2[169]) );
  NANDN U1329 ( .A(xregN_1), .B(zin[168]), .Z(n889) );
  NAND U1330 ( .A(N173), .B(xregN_1), .Z(n888) );
  NAND U1331 ( .A(n890), .B(n891), .Z(z2[168]) );
  NANDN U1332 ( .A(xregN_1), .B(zin[167]), .Z(n891) );
  NAND U1333 ( .A(N172), .B(xregN_1), .Z(n890) );
  NAND U1334 ( .A(n892), .B(n893), .Z(z2[167]) );
  NANDN U1335 ( .A(xregN_1), .B(zin[166]), .Z(n893) );
  NAND U1336 ( .A(N171), .B(xregN_1), .Z(n892) );
  NAND U1337 ( .A(n894), .B(n895), .Z(z2[166]) );
  NANDN U1338 ( .A(xregN_1), .B(zin[165]), .Z(n895) );
  NAND U1339 ( .A(N170), .B(xregN_1), .Z(n894) );
  NAND U1340 ( .A(n896), .B(n897), .Z(z2[165]) );
  NANDN U1341 ( .A(xregN_1), .B(zin[164]), .Z(n897) );
  NAND U1342 ( .A(N169), .B(xregN_1), .Z(n896) );
  NAND U1343 ( .A(n898), .B(n899), .Z(z2[164]) );
  NANDN U1344 ( .A(xregN_1), .B(zin[163]), .Z(n899) );
  NAND U1345 ( .A(N168), .B(xregN_1), .Z(n898) );
  NAND U1346 ( .A(n900), .B(n901), .Z(z2[163]) );
  NANDN U1347 ( .A(xregN_1), .B(zin[162]), .Z(n901) );
  NAND U1348 ( .A(N167), .B(xregN_1), .Z(n900) );
  NAND U1349 ( .A(n902), .B(n903), .Z(z2[162]) );
  NANDN U1350 ( .A(xregN_1), .B(zin[161]), .Z(n903) );
  NAND U1351 ( .A(N166), .B(xregN_1), .Z(n902) );
  NAND U1352 ( .A(n904), .B(n905), .Z(z2[161]) );
  NANDN U1353 ( .A(xregN_1), .B(zin[160]), .Z(n905) );
  NAND U1354 ( .A(N165), .B(xregN_1), .Z(n904) );
  NAND U1355 ( .A(n906), .B(n907), .Z(z2[160]) );
  NANDN U1356 ( .A(xregN_1), .B(zin[159]), .Z(n907) );
  NAND U1357 ( .A(N164), .B(xregN_1), .Z(n906) );
  NAND U1358 ( .A(n908), .B(n909), .Z(z2[15]) );
  NANDN U1359 ( .A(xregN_1), .B(zin[14]), .Z(n909) );
  NAND U1360 ( .A(N19), .B(xregN_1), .Z(n908) );
  NAND U1361 ( .A(n910), .B(n911), .Z(z2[159]) );
  NANDN U1362 ( .A(xregN_1), .B(zin[158]), .Z(n911) );
  NAND U1363 ( .A(N163), .B(xregN_1), .Z(n910) );
  NAND U1364 ( .A(n912), .B(n913), .Z(z2[158]) );
  NANDN U1365 ( .A(xregN_1), .B(zin[157]), .Z(n913) );
  NAND U1366 ( .A(N162), .B(xregN_1), .Z(n912) );
  NAND U1367 ( .A(n914), .B(n915), .Z(z2[157]) );
  NANDN U1368 ( .A(xregN_1), .B(zin[156]), .Z(n915) );
  NAND U1369 ( .A(N161), .B(xregN_1), .Z(n914) );
  NAND U1370 ( .A(n916), .B(n917), .Z(z2[156]) );
  NANDN U1371 ( .A(xregN_1), .B(zin[155]), .Z(n917) );
  NAND U1372 ( .A(N160), .B(xregN_1), .Z(n916) );
  NAND U1373 ( .A(n918), .B(n919), .Z(z2[155]) );
  NANDN U1374 ( .A(xregN_1), .B(zin[154]), .Z(n919) );
  NAND U1375 ( .A(N159), .B(xregN_1), .Z(n918) );
  NAND U1376 ( .A(n920), .B(n921), .Z(z2[154]) );
  NANDN U1377 ( .A(xregN_1), .B(zin[153]), .Z(n921) );
  NAND U1378 ( .A(N158), .B(xregN_1), .Z(n920) );
  NAND U1379 ( .A(n922), .B(n923), .Z(z2[153]) );
  NANDN U1380 ( .A(xregN_1), .B(zin[152]), .Z(n923) );
  NAND U1381 ( .A(N157), .B(xregN_1), .Z(n922) );
  NAND U1382 ( .A(n924), .B(n925), .Z(z2[152]) );
  NANDN U1383 ( .A(xregN_1), .B(zin[151]), .Z(n925) );
  NAND U1384 ( .A(N156), .B(xregN_1), .Z(n924) );
  NAND U1385 ( .A(n926), .B(n927), .Z(z2[151]) );
  NANDN U1386 ( .A(xregN_1), .B(zin[150]), .Z(n927) );
  NAND U1387 ( .A(N155), .B(xregN_1), .Z(n926) );
  NAND U1388 ( .A(n928), .B(n929), .Z(z2[150]) );
  NANDN U1389 ( .A(xregN_1), .B(zin[149]), .Z(n929) );
  NAND U1390 ( .A(N154), .B(xregN_1), .Z(n928) );
  NAND U1391 ( .A(n930), .B(n931), .Z(z2[14]) );
  NANDN U1392 ( .A(xregN_1), .B(zin[13]), .Z(n931) );
  NAND U1393 ( .A(N18), .B(xregN_1), .Z(n930) );
  NAND U1394 ( .A(n932), .B(n933), .Z(z2[149]) );
  NANDN U1395 ( .A(xregN_1), .B(zin[148]), .Z(n933) );
  NAND U1396 ( .A(N153), .B(xregN_1), .Z(n932) );
  NAND U1397 ( .A(n934), .B(n935), .Z(z2[148]) );
  NANDN U1398 ( .A(xregN_1), .B(zin[147]), .Z(n935) );
  NAND U1399 ( .A(N152), .B(xregN_1), .Z(n934) );
  NAND U1400 ( .A(n936), .B(n937), .Z(z2[147]) );
  NANDN U1401 ( .A(xregN_1), .B(zin[146]), .Z(n937) );
  NAND U1402 ( .A(N151), .B(xregN_1), .Z(n936) );
  NAND U1403 ( .A(n938), .B(n939), .Z(z2[146]) );
  NANDN U1404 ( .A(xregN_1), .B(zin[145]), .Z(n939) );
  NAND U1405 ( .A(N150), .B(xregN_1), .Z(n938) );
  NAND U1406 ( .A(n940), .B(n941), .Z(z2[145]) );
  NANDN U1407 ( .A(xregN_1), .B(zin[144]), .Z(n941) );
  NAND U1408 ( .A(N149), .B(xregN_1), .Z(n940) );
  NAND U1409 ( .A(n942), .B(n943), .Z(z2[144]) );
  NANDN U1410 ( .A(xregN_1), .B(zin[143]), .Z(n943) );
  NAND U1411 ( .A(N148), .B(xregN_1), .Z(n942) );
  NAND U1412 ( .A(n944), .B(n945), .Z(z2[143]) );
  NANDN U1413 ( .A(xregN_1), .B(zin[142]), .Z(n945) );
  NAND U1414 ( .A(N147), .B(xregN_1), .Z(n944) );
  NAND U1415 ( .A(n946), .B(n947), .Z(z2[142]) );
  NANDN U1416 ( .A(xregN_1), .B(zin[141]), .Z(n947) );
  NAND U1417 ( .A(N146), .B(xregN_1), .Z(n946) );
  NAND U1418 ( .A(n948), .B(n949), .Z(z2[141]) );
  NANDN U1419 ( .A(xregN_1), .B(zin[140]), .Z(n949) );
  NAND U1420 ( .A(N145), .B(xregN_1), .Z(n948) );
  NAND U1421 ( .A(n950), .B(n951), .Z(z2[140]) );
  NANDN U1422 ( .A(xregN_1), .B(zin[139]), .Z(n951) );
  NAND U1423 ( .A(N144), .B(xregN_1), .Z(n950) );
  NAND U1424 ( .A(n952), .B(n953), .Z(z2[13]) );
  NANDN U1425 ( .A(xregN_1), .B(zin[12]), .Z(n953) );
  NAND U1426 ( .A(N17), .B(xregN_1), .Z(n952) );
  NAND U1427 ( .A(n954), .B(n955), .Z(z2[139]) );
  NANDN U1428 ( .A(xregN_1), .B(zin[138]), .Z(n955) );
  NAND U1429 ( .A(N143), .B(xregN_1), .Z(n954) );
  NAND U1430 ( .A(n956), .B(n957), .Z(z2[138]) );
  NANDN U1431 ( .A(xregN_1), .B(zin[137]), .Z(n957) );
  NAND U1432 ( .A(N142), .B(xregN_1), .Z(n956) );
  NAND U1433 ( .A(n958), .B(n959), .Z(z2[137]) );
  NANDN U1434 ( .A(xregN_1), .B(zin[136]), .Z(n959) );
  NAND U1435 ( .A(N141), .B(xregN_1), .Z(n958) );
  NAND U1436 ( .A(n960), .B(n961), .Z(z2[136]) );
  NANDN U1437 ( .A(xregN_1), .B(zin[135]), .Z(n961) );
  NAND U1438 ( .A(N140), .B(xregN_1), .Z(n960) );
  NAND U1439 ( .A(n962), .B(n963), .Z(z2[135]) );
  NANDN U1440 ( .A(xregN_1), .B(zin[134]), .Z(n963) );
  NAND U1441 ( .A(N139), .B(xregN_1), .Z(n962) );
  NAND U1442 ( .A(n964), .B(n965), .Z(z2[134]) );
  NANDN U1443 ( .A(xregN_1), .B(zin[133]), .Z(n965) );
  NAND U1444 ( .A(N138), .B(xregN_1), .Z(n964) );
  NAND U1445 ( .A(n966), .B(n967), .Z(z2[133]) );
  NANDN U1446 ( .A(xregN_1), .B(zin[132]), .Z(n967) );
  NAND U1447 ( .A(N137), .B(xregN_1), .Z(n966) );
  NAND U1448 ( .A(n968), .B(n969), .Z(z2[132]) );
  NANDN U1449 ( .A(xregN_1), .B(zin[131]), .Z(n969) );
  NAND U1450 ( .A(N136), .B(xregN_1), .Z(n968) );
  NAND U1451 ( .A(n970), .B(n971), .Z(z2[131]) );
  NANDN U1452 ( .A(xregN_1), .B(zin[130]), .Z(n971) );
  NAND U1453 ( .A(N135), .B(xregN_1), .Z(n970) );
  NAND U1454 ( .A(n972), .B(n973), .Z(z2[130]) );
  NANDN U1455 ( .A(xregN_1), .B(zin[129]), .Z(n973) );
  NAND U1456 ( .A(N134), .B(xregN_1), .Z(n972) );
  NAND U1457 ( .A(n974), .B(n975), .Z(z2[12]) );
  NANDN U1458 ( .A(xregN_1), .B(zin[11]), .Z(n975) );
  NAND U1459 ( .A(N16), .B(xregN_1), .Z(n974) );
  NAND U1460 ( .A(n976), .B(n977), .Z(z2[129]) );
  NANDN U1461 ( .A(xregN_1), .B(zin[128]), .Z(n977) );
  NAND U1462 ( .A(N133), .B(xregN_1), .Z(n976) );
  NAND U1463 ( .A(n978), .B(n979), .Z(z2[128]) );
  NANDN U1464 ( .A(xregN_1), .B(zin[127]), .Z(n979) );
  NAND U1465 ( .A(N132), .B(xregN_1), .Z(n978) );
  NAND U1466 ( .A(n980), .B(n981), .Z(z2[127]) );
  NANDN U1467 ( .A(xregN_1), .B(zin[126]), .Z(n981) );
  NAND U1468 ( .A(N131), .B(xregN_1), .Z(n980) );
  NAND U1469 ( .A(n982), .B(n983), .Z(z2[126]) );
  NANDN U1470 ( .A(xregN_1), .B(zin[125]), .Z(n983) );
  NAND U1471 ( .A(N130), .B(xregN_1), .Z(n982) );
  NAND U1472 ( .A(n984), .B(n985), .Z(z2[125]) );
  NANDN U1473 ( .A(xregN_1), .B(zin[124]), .Z(n985) );
  NAND U1474 ( .A(N129), .B(xregN_1), .Z(n984) );
  NAND U1475 ( .A(n986), .B(n987), .Z(z2[124]) );
  NANDN U1476 ( .A(xregN_1), .B(zin[123]), .Z(n987) );
  NAND U1477 ( .A(N128), .B(xregN_1), .Z(n986) );
  NAND U1478 ( .A(n988), .B(n989), .Z(z2[123]) );
  NANDN U1479 ( .A(xregN_1), .B(zin[122]), .Z(n989) );
  NAND U1480 ( .A(N127), .B(xregN_1), .Z(n988) );
  NAND U1481 ( .A(n990), .B(n991), .Z(z2[122]) );
  NANDN U1482 ( .A(xregN_1), .B(zin[121]), .Z(n991) );
  NAND U1483 ( .A(N126), .B(xregN_1), .Z(n990) );
  NAND U1484 ( .A(n992), .B(n993), .Z(z2[121]) );
  NANDN U1485 ( .A(xregN_1), .B(zin[120]), .Z(n993) );
  NAND U1486 ( .A(N125), .B(xregN_1), .Z(n992) );
  NAND U1487 ( .A(n994), .B(n995), .Z(z2[120]) );
  NANDN U1488 ( .A(xregN_1), .B(zin[119]), .Z(n995) );
  NAND U1489 ( .A(N124), .B(xregN_1), .Z(n994) );
  NAND U1490 ( .A(n996), .B(n997), .Z(z2[11]) );
  NANDN U1491 ( .A(xregN_1), .B(zin[10]), .Z(n997) );
  NAND U1492 ( .A(N15), .B(xregN_1), .Z(n996) );
  NAND U1493 ( .A(n998), .B(n999), .Z(z2[119]) );
  NANDN U1494 ( .A(xregN_1), .B(zin[118]), .Z(n999) );
  NAND U1495 ( .A(N123), .B(xregN_1), .Z(n998) );
  NAND U1496 ( .A(n1000), .B(n1001), .Z(z2[118]) );
  NANDN U1497 ( .A(xregN_1), .B(zin[117]), .Z(n1001) );
  NAND U1498 ( .A(N122), .B(xregN_1), .Z(n1000) );
  NAND U1499 ( .A(n1002), .B(n1003), .Z(z2[117]) );
  NANDN U1500 ( .A(xregN_1), .B(zin[116]), .Z(n1003) );
  NAND U1501 ( .A(N121), .B(xregN_1), .Z(n1002) );
  NAND U1502 ( .A(n1004), .B(n1005), .Z(z2[116]) );
  NANDN U1503 ( .A(xregN_1), .B(zin[115]), .Z(n1005) );
  NAND U1504 ( .A(N120), .B(xregN_1), .Z(n1004) );
  NAND U1505 ( .A(n1006), .B(n1007), .Z(z2[115]) );
  NANDN U1506 ( .A(xregN_1), .B(zin[114]), .Z(n1007) );
  NAND U1507 ( .A(N119), .B(xregN_1), .Z(n1006) );
  NAND U1508 ( .A(n1008), .B(n1009), .Z(z2[114]) );
  NANDN U1509 ( .A(xregN_1), .B(zin[113]), .Z(n1009) );
  NAND U1510 ( .A(N118), .B(xregN_1), .Z(n1008) );
  NAND U1511 ( .A(n1010), .B(n1011), .Z(z2[113]) );
  NANDN U1512 ( .A(xregN_1), .B(zin[112]), .Z(n1011) );
  NAND U1513 ( .A(N117), .B(xregN_1), .Z(n1010) );
  NAND U1514 ( .A(n1012), .B(n1013), .Z(z2[112]) );
  NANDN U1515 ( .A(xregN_1), .B(zin[111]), .Z(n1013) );
  NAND U1516 ( .A(N116), .B(xregN_1), .Z(n1012) );
  NAND U1517 ( .A(n1014), .B(n1015), .Z(z2[111]) );
  NANDN U1518 ( .A(xregN_1), .B(zin[110]), .Z(n1015) );
  NAND U1519 ( .A(N115), .B(xregN_1), .Z(n1014) );
  NAND U1520 ( .A(n1016), .B(n1017), .Z(z2[110]) );
  NANDN U1521 ( .A(xregN_1), .B(zin[109]), .Z(n1017) );
  NAND U1522 ( .A(N114), .B(xregN_1), .Z(n1016) );
  NAND U1523 ( .A(n1018), .B(n1019), .Z(z2[10]) );
  NANDN U1524 ( .A(xregN_1), .B(zin[9]), .Z(n1019) );
  NAND U1525 ( .A(N14), .B(xregN_1), .Z(n1018) );
  NAND U1526 ( .A(n1020), .B(n1021), .Z(z2[109]) );
  NANDN U1527 ( .A(xregN_1), .B(zin[108]), .Z(n1021) );
  NAND U1528 ( .A(N113), .B(xregN_1), .Z(n1020) );
  NAND U1529 ( .A(n1022), .B(n1023), .Z(z2[108]) );
  NANDN U1530 ( .A(xregN_1), .B(zin[107]), .Z(n1023) );
  NAND U1531 ( .A(N112), .B(xregN_1), .Z(n1022) );
  NAND U1532 ( .A(n1024), .B(n1025), .Z(z2[107]) );
  NANDN U1533 ( .A(xregN_1), .B(zin[106]), .Z(n1025) );
  NAND U1534 ( .A(N111), .B(xregN_1), .Z(n1024) );
  NAND U1535 ( .A(n1026), .B(n1027), .Z(z2[106]) );
  NANDN U1536 ( .A(xregN_1), .B(zin[105]), .Z(n1027) );
  NAND U1537 ( .A(N110), .B(xregN_1), .Z(n1026) );
  NAND U1538 ( .A(n1028), .B(n1029), .Z(z2[105]) );
  NANDN U1539 ( .A(xregN_1), .B(zin[104]), .Z(n1029) );
  NAND U1540 ( .A(N109), .B(xregN_1), .Z(n1028) );
  NAND U1541 ( .A(n1030), .B(n1031), .Z(z2[104]) );
  NANDN U1542 ( .A(xregN_1), .B(zin[103]), .Z(n1031) );
  NAND U1543 ( .A(N108), .B(xregN_1), .Z(n1030) );
  NAND U1544 ( .A(n1032), .B(n1033), .Z(z2[103]) );
  NANDN U1545 ( .A(xregN_1), .B(zin[102]), .Z(n1033) );
  NAND U1546 ( .A(N107), .B(xregN_1), .Z(n1032) );
  NAND U1547 ( .A(n1034), .B(n1035), .Z(z2[102]) );
  NANDN U1548 ( .A(xregN_1), .B(zin[101]), .Z(n1035) );
  NAND U1549 ( .A(N106), .B(xregN_1), .Z(n1034) );
  NAND U1550 ( .A(n1036), .B(n1037), .Z(z2[101]) );
  NANDN U1551 ( .A(xregN_1), .B(zin[100]), .Z(n1037) );
  NAND U1552 ( .A(N105), .B(xregN_1), .Z(n1036) );
  NAND U1553 ( .A(n1038), .B(n1039), .Z(z2[100]) );
  NANDN U1554 ( .A(xregN_1), .B(zin[99]), .Z(n1039) );
  NAND U1555 ( .A(N104), .B(xregN_1), .Z(n1038) );
  AND U1556 ( .A(N4), .B(xregN_1), .Z(z2[0]) );
endmodule


module modmult_step_N256_5_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279;

  IV U1 ( .A(n1278), .Z(n1) );
  IV U2 ( .A(A[1]), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(DIFF[9]) );
  XOR U4 ( .A(B[9]), .B(A[9]), .Z(n4) );
  XNOR U5 ( .A(n5), .B(n6), .Z(DIFF[99]) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(DIFF[98]) );
  XOR U8 ( .A(B[98]), .B(A[98]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(DIFF[97]) );
  XOR U10 ( .A(B[97]), .B(A[97]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(DIFF[96]) );
  XOR U12 ( .A(B[96]), .B(A[96]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(DIFF[95]) );
  XOR U14 ( .A(B[95]), .B(A[95]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(DIFF[94]) );
  XOR U16 ( .A(B[94]), .B(A[94]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(DIFF[93]) );
  XOR U18 ( .A(B[93]), .B(A[93]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(DIFF[92]) );
  XOR U20 ( .A(B[92]), .B(A[92]), .Z(n20) );
  XOR U21 ( .A(n21), .B(n22), .Z(DIFF[91]) );
  XOR U22 ( .A(B[91]), .B(A[91]), .Z(n22) );
  XOR U23 ( .A(n23), .B(n24), .Z(DIFF[90]) );
  XOR U24 ( .A(B[90]), .B(A[90]), .Z(n24) );
  XOR U25 ( .A(n25), .B(n26), .Z(DIFF[8]) );
  XOR U26 ( .A(B[8]), .B(A[8]), .Z(n26) );
  XOR U27 ( .A(n27), .B(n28), .Z(DIFF[89]) );
  XOR U28 ( .A(B[89]), .B(A[89]), .Z(n28) );
  XOR U29 ( .A(n29), .B(n30), .Z(DIFF[88]) );
  XOR U30 ( .A(B[88]), .B(A[88]), .Z(n30) );
  XOR U31 ( .A(n31), .B(n32), .Z(DIFF[87]) );
  XOR U32 ( .A(B[87]), .B(A[87]), .Z(n32) );
  XOR U33 ( .A(n33), .B(n34), .Z(DIFF[86]) );
  XOR U34 ( .A(B[86]), .B(A[86]), .Z(n34) );
  XOR U35 ( .A(n35), .B(n36), .Z(DIFF[85]) );
  XOR U36 ( .A(B[85]), .B(A[85]), .Z(n36) );
  XOR U37 ( .A(n37), .B(n38), .Z(DIFF[84]) );
  XOR U38 ( .A(B[84]), .B(A[84]), .Z(n38) );
  XOR U39 ( .A(n39), .B(n40), .Z(DIFF[83]) );
  XOR U40 ( .A(B[83]), .B(A[83]), .Z(n40) );
  XOR U41 ( .A(n41), .B(n42), .Z(DIFF[82]) );
  XOR U42 ( .A(B[82]), .B(A[82]), .Z(n42) );
  XOR U43 ( .A(n43), .B(n44), .Z(DIFF[81]) );
  XOR U44 ( .A(B[81]), .B(A[81]), .Z(n44) );
  XOR U45 ( .A(n45), .B(n46), .Z(DIFF[80]) );
  XOR U46 ( .A(B[80]), .B(A[80]), .Z(n46) );
  XOR U47 ( .A(n47), .B(n48), .Z(DIFF[7]) );
  XOR U48 ( .A(B[7]), .B(A[7]), .Z(n48) );
  XOR U49 ( .A(n49), .B(n50), .Z(DIFF[79]) );
  XOR U50 ( .A(B[79]), .B(A[79]), .Z(n50) );
  XOR U51 ( .A(n51), .B(n52), .Z(DIFF[78]) );
  XOR U52 ( .A(B[78]), .B(A[78]), .Z(n52) );
  XOR U53 ( .A(n53), .B(n54), .Z(DIFF[77]) );
  XOR U54 ( .A(B[77]), .B(A[77]), .Z(n54) );
  XOR U55 ( .A(n55), .B(n56), .Z(DIFF[76]) );
  XOR U56 ( .A(B[76]), .B(A[76]), .Z(n56) );
  XOR U57 ( .A(n57), .B(n58), .Z(DIFF[75]) );
  XOR U58 ( .A(B[75]), .B(A[75]), .Z(n58) );
  XOR U59 ( .A(n59), .B(n60), .Z(DIFF[74]) );
  XOR U60 ( .A(B[74]), .B(A[74]), .Z(n60) );
  XOR U61 ( .A(n61), .B(n62), .Z(DIFF[73]) );
  XOR U62 ( .A(B[73]), .B(A[73]), .Z(n62) );
  XOR U63 ( .A(n63), .B(n64), .Z(DIFF[72]) );
  XOR U64 ( .A(B[72]), .B(A[72]), .Z(n64) );
  XOR U65 ( .A(n65), .B(n66), .Z(DIFF[71]) );
  XOR U66 ( .A(B[71]), .B(A[71]), .Z(n66) );
  XOR U67 ( .A(n67), .B(n68), .Z(DIFF[70]) );
  XOR U68 ( .A(B[70]), .B(A[70]), .Z(n68) );
  XOR U69 ( .A(n69), .B(n70), .Z(DIFF[6]) );
  XOR U70 ( .A(B[6]), .B(A[6]), .Z(n70) );
  XOR U71 ( .A(n71), .B(n72), .Z(DIFF[69]) );
  XOR U72 ( .A(B[69]), .B(A[69]), .Z(n72) );
  XOR U73 ( .A(n73), .B(n74), .Z(DIFF[68]) );
  XOR U74 ( .A(B[68]), .B(A[68]), .Z(n74) );
  XOR U75 ( .A(n75), .B(n76), .Z(DIFF[67]) );
  XOR U76 ( .A(B[67]), .B(A[67]), .Z(n76) );
  XOR U77 ( .A(n77), .B(n78), .Z(DIFF[66]) );
  XOR U78 ( .A(B[66]), .B(A[66]), .Z(n78) );
  XOR U79 ( .A(n79), .B(n80), .Z(DIFF[65]) );
  XOR U80 ( .A(B[65]), .B(A[65]), .Z(n80) );
  XOR U81 ( .A(n81), .B(n82), .Z(DIFF[64]) );
  XOR U82 ( .A(B[64]), .B(A[64]), .Z(n82) );
  XOR U83 ( .A(n83), .B(n84), .Z(DIFF[63]) );
  XOR U84 ( .A(B[63]), .B(A[63]), .Z(n84) );
  XOR U85 ( .A(n85), .B(n86), .Z(DIFF[62]) );
  XOR U86 ( .A(B[62]), .B(A[62]), .Z(n86) );
  XOR U87 ( .A(n87), .B(n88), .Z(DIFF[61]) );
  XOR U88 ( .A(B[61]), .B(A[61]), .Z(n88) );
  XOR U89 ( .A(n89), .B(n90), .Z(DIFF[60]) );
  XOR U90 ( .A(B[60]), .B(A[60]), .Z(n90) );
  XOR U91 ( .A(n91), .B(n92), .Z(DIFF[5]) );
  XOR U92 ( .A(B[5]), .B(A[5]), .Z(n92) );
  XOR U93 ( .A(n93), .B(n94), .Z(DIFF[59]) );
  XOR U94 ( .A(B[59]), .B(A[59]), .Z(n94) );
  XOR U95 ( .A(n95), .B(n96), .Z(DIFF[58]) );
  XOR U96 ( .A(B[58]), .B(A[58]), .Z(n96) );
  XOR U97 ( .A(n97), .B(n98), .Z(DIFF[57]) );
  XOR U98 ( .A(B[57]), .B(A[57]), .Z(n98) );
  XOR U99 ( .A(n99), .B(n100), .Z(DIFF[56]) );
  XOR U100 ( .A(B[56]), .B(A[56]), .Z(n100) );
  XOR U101 ( .A(n101), .B(n102), .Z(DIFF[55]) );
  XOR U102 ( .A(B[55]), .B(A[55]), .Z(n102) );
  XOR U103 ( .A(n103), .B(n104), .Z(DIFF[54]) );
  XOR U104 ( .A(B[54]), .B(A[54]), .Z(n104) );
  XOR U105 ( .A(n105), .B(n106), .Z(DIFF[53]) );
  XOR U106 ( .A(B[53]), .B(A[53]), .Z(n106) );
  XOR U107 ( .A(n107), .B(n108), .Z(DIFF[52]) );
  XOR U108 ( .A(B[52]), .B(A[52]), .Z(n108) );
  XOR U109 ( .A(n109), .B(n110), .Z(DIFF[51]) );
  XOR U110 ( .A(B[51]), .B(A[51]), .Z(n110) );
  XOR U111 ( .A(n111), .B(n112), .Z(DIFF[50]) );
  XOR U112 ( .A(B[50]), .B(A[50]), .Z(n112) );
  XOR U113 ( .A(n113), .B(n114), .Z(DIFF[4]) );
  XOR U114 ( .A(B[4]), .B(A[4]), .Z(n114) );
  XOR U115 ( .A(n115), .B(n116), .Z(DIFF[49]) );
  XOR U116 ( .A(B[49]), .B(A[49]), .Z(n116) );
  XOR U117 ( .A(n117), .B(n118), .Z(DIFF[48]) );
  XOR U118 ( .A(B[48]), .B(A[48]), .Z(n118) );
  XOR U119 ( .A(n119), .B(n120), .Z(DIFF[47]) );
  XOR U120 ( .A(B[47]), .B(A[47]), .Z(n120) );
  XOR U121 ( .A(n121), .B(n122), .Z(DIFF[46]) );
  XOR U122 ( .A(B[46]), .B(A[46]), .Z(n122) );
  XOR U123 ( .A(n123), .B(n124), .Z(DIFF[45]) );
  XOR U124 ( .A(B[45]), .B(A[45]), .Z(n124) );
  XOR U125 ( .A(n125), .B(n126), .Z(DIFF[44]) );
  XOR U126 ( .A(B[44]), .B(A[44]), .Z(n126) );
  XOR U127 ( .A(n127), .B(n128), .Z(DIFF[43]) );
  XOR U128 ( .A(B[43]), .B(A[43]), .Z(n128) );
  XOR U129 ( .A(n129), .B(n130), .Z(DIFF[42]) );
  XOR U130 ( .A(B[42]), .B(A[42]), .Z(n130) );
  XOR U131 ( .A(n131), .B(n132), .Z(DIFF[41]) );
  XOR U132 ( .A(B[41]), .B(A[41]), .Z(n132) );
  XOR U133 ( .A(n133), .B(n134), .Z(DIFF[40]) );
  XOR U134 ( .A(B[40]), .B(A[40]), .Z(n134) );
  XOR U135 ( .A(n135), .B(n136), .Z(DIFF[3]) );
  XOR U136 ( .A(B[3]), .B(A[3]), .Z(n136) );
  XOR U137 ( .A(n137), .B(n138), .Z(DIFF[39]) );
  XOR U138 ( .A(B[39]), .B(A[39]), .Z(n138) );
  XOR U139 ( .A(n139), .B(n140), .Z(DIFF[38]) );
  XOR U140 ( .A(B[38]), .B(A[38]), .Z(n140) );
  XOR U141 ( .A(n141), .B(n142), .Z(DIFF[37]) );
  XOR U142 ( .A(B[37]), .B(A[37]), .Z(n142) );
  XOR U143 ( .A(n143), .B(n144), .Z(DIFF[36]) );
  XOR U144 ( .A(B[36]), .B(A[36]), .Z(n144) );
  XOR U145 ( .A(n145), .B(n146), .Z(DIFF[35]) );
  XOR U146 ( .A(B[35]), .B(A[35]), .Z(n146) );
  XOR U147 ( .A(n147), .B(n148), .Z(DIFF[34]) );
  XOR U148 ( .A(B[34]), .B(A[34]), .Z(n148) );
  XOR U149 ( .A(n149), .B(n150), .Z(DIFF[33]) );
  XOR U150 ( .A(B[33]), .B(A[33]), .Z(n150) );
  XOR U151 ( .A(n151), .B(n152), .Z(DIFF[32]) );
  XOR U152 ( .A(B[32]), .B(A[32]), .Z(n152) );
  XOR U153 ( .A(n153), .B(n154), .Z(DIFF[31]) );
  XOR U154 ( .A(B[31]), .B(A[31]), .Z(n154) );
  XOR U155 ( .A(n155), .B(n156), .Z(DIFF[30]) );
  XOR U156 ( .A(B[30]), .B(A[30]), .Z(n156) );
  XOR U157 ( .A(n157), .B(n158), .Z(DIFF[2]) );
  XOR U158 ( .A(B[2]), .B(A[2]), .Z(n158) );
  XOR U159 ( .A(n159), .B(n160), .Z(DIFF[29]) );
  XOR U160 ( .A(B[29]), .B(A[29]), .Z(n160) );
  XOR U161 ( .A(n161), .B(n162), .Z(DIFF[28]) );
  XOR U162 ( .A(B[28]), .B(A[28]), .Z(n162) );
  XOR U163 ( .A(n163), .B(n164), .Z(DIFF[27]) );
  XOR U164 ( .A(B[27]), .B(A[27]), .Z(n164) );
  XOR U165 ( .A(n165), .B(n166), .Z(DIFF[26]) );
  XOR U166 ( .A(B[26]), .B(A[26]), .Z(n166) );
  XOR U167 ( .A(n167), .B(n168), .Z(DIFF[25]) );
  XOR U168 ( .A(B[25]), .B(A[25]), .Z(n168) );
  XOR U169 ( .A(A[256]), .B(n169), .Z(DIFF[256]) );
  AND U170 ( .A(n170), .B(n171), .Z(n169) );
  NANDN U171 ( .A(B[255]), .B(n172), .Z(n171) );
  NANDN U172 ( .A(A[255]), .B(n173), .Z(n172) );
  NANDN U173 ( .A(n173), .B(A[255]), .Z(n170) );
  XOR U174 ( .A(n173), .B(n174), .Z(DIFF[255]) );
  XOR U175 ( .A(B[255]), .B(A[255]), .Z(n174) );
  AND U176 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U177 ( .A(B[254]), .B(n177), .Z(n176) );
  NANDN U178 ( .A(A[254]), .B(n178), .Z(n177) );
  NANDN U179 ( .A(n178), .B(A[254]), .Z(n175) );
  XOR U180 ( .A(n178), .B(n179), .Z(DIFF[254]) );
  XOR U181 ( .A(B[254]), .B(A[254]), .Z(n179) );
  AND U182 ( .A(n180), .B(n181), .Z(n178) );
  NANDN U183 ( .A(B[253]), .B(n182), .Z(n181) );
  NANDN U184 ( .A(A[253]), .B(n183), .Z(n182) );
  NANDN U185 ( .A(n183), .B(A[253]), .Z(n180) );
  XOR U186 ( .A(n183), .B(n184), .Z(DIFF[253]) );
  XOR U187 ( .A(B[253]), .B(A[253]), .Z(n184) );
  AND U188 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U189 ( .A(B[252]), .B(n187), .Z(n186) );
  NANDN U190 ( .A(A[252]), .B(n188), .Z(n187) );
  NANDN U191 ( .A(n188), .B(A[252]), .Z(n185) );
  XOR U192 ( .A(n188), .B(n189), .Z(DIFF[252]) );
  XOR U193 ( .A(B[252]), .B(A[252]), .Z(n189) );
  AND U194 ( .A(n190), .B(n191), .Z(n188) );
  NANDN U195 ( .A(B[251]), .B(n192), .Z(n191) );
  NANDN U196 ( .A(A[251]), .B(n193), .Z(n192) );
  NANDN U197 ( .A(n193), .B(A[251]), .Z(n190) );
  XOR U198 ( .A(n193), .B(n194), .Z(DIFF[251]) );
  XOR U199 ( .A(B[251]), .B(A[251]), .Z(n194) );
  AND U200 ( .A(n195), .B(n196), .Z(n193) );
  NANDN U201 ( .A(B[250]), .B(n197), .Z(n196) );
  NANDN U202 ( .A(A[250]), .B(n198), .Z(n197) );
  NANDN U203 ( .A(n198), .B(A[250]), .Z(n195) );
  XOR U204 ( .A(n198), .B(n199), .Z(DIFF[250]) );
  XOR U205 ( .A(B[250]), .B(A[250]), .Z(n199) );
  AND U206 ( .A(n200), .B(n201), .Z(n198) );
  NANDN U207 ( .A(B[249]), .B(n202), .Z(n201) );
  NANDN U208 ( .A(A[249]), .B(n203), .Z(n202) );
  NANDN U209 ( .A(n203), .B(A[249]), .Z(n200) );
  XOR U210 ( .A(n204), .B(n205), .Z(DIFF[24]) );
  XOR U211 ( .A(B[24]), .B(A[24]), .Z(n205) );
  XOR U212 ( .A(n203), .B(n206), .Z(DIFF[249]) );
  XOR U213 ( .A(B[249]), .B(A[249]), .Z(n206) );
  AND U214 ( .A(n207), .B(n208), .Z(n203) );
  NANDN U215 ( .A(B[248]), .B(n209), .Z(n208) );
  NANDN U216 ( .A(A[248]), .B(n210), .Z(n209) );
  NANDN U217 ( .A(n210), .B(A[248]), .Z(n207) );
  XOR U218 ( .A(n210), .B(n211), .Z(DIFF[248]) );
  XOR U219 ( .A(B[248]), .B(A[248]), .Z(n211) );
  AND U220 ( .A(n212), .B(n213), .Z(n210) );
  NANDN U221 ( .A(B[247]), .B(n214), .Z(n213) );
  NANDN U222 ( .A(A[247]), .B(n215), .Z(n214) );
  NANDN U223 ( .A(n215), .B(A[247]), .Z(n212) );
  XOR U224 ( .A(n215), .B(n216), .Z(DIFF[247]) );
  XOR U225 ( .A(B[247]), .B(A[247]), .Z(n216) );
  AND U226 ( .A(n217), .B(n218), .Z(n215) );
  NANDN U227 ( .A(B[246]), .B(n219), .Z(n218) );
  NANDN U228 ( .A(A[246]), .B(n220), .Z(n219) );
  NANDN U229 ( .A(n220), .B(A[246]), .Z(n217) );
  XOR U230 ( .A(n220), .B(n221), .Z(DIFF[246]) );
  XOR U231 ( .A(B[246]), .B(A[246]), .Z(n221) );
  AND U232 ( .A(n222), .B(n223), .Z(n220) );
  NANDN U233 ( .A(B[245]), .B(n224), .Z(n223) );
  NANDN U234 ( .A(A[245]), .B(n225), .Z(n224) );
  NANDN U235 ( .A(n225), .B(A[245]), .Z(n222) );
  XOR U236 ( .A(n225), .B(n226), .Z(DIFF[245]) );
  XOR U237 ( .A(B[245]), .B(A[245]), .Z(n226) );
  AND U238 ( .A(n227), .B(n228), .Z(n225) );
  NANDN U239 ( .A(B[244]), .B(n229), .Z(n228) );
  NANDN U240 ( .A(A[244]), .B(n230), .Z(n229) );
  NANDN U241 ( .A(n230), .B(A[244]), .Z(n227) );
  XOR U242 ( .A(n230), .B(n231), .Z(DIFF[244]) );
  XOR U243 ( .A(B[244]), .B(A[244]), .Z(n231) );
  AND U244 ( .A(n232), .B(n233), .Z(n230) );
  NANDN U245 ( .A(B[243]), .B(n234), .Z(n233) );
  NANDN U246 ( .A(A[243]), .B(n235), .Z(n234) );
  NANDN U247 ( .A(n235), .B(A[243]), .Z(n232) );
  XOR U248 ( .A(n235), .B(n236), .Z(DIFF[243]) );
  XOR U249 ( .A(B[243]), .B(A[243]), .Z(n236) );
  AND U250 ( .A(n237), .B(n238), .Z(n235) );
  NANDN U251 ( .A(B[242]), .B(n239), .Z(n238) );
  NANDN U252 ( .A(A[242]), .B(n240), .Z(n239) );
  NANDN U253 ( .A(n240), .B(A[242]), .Z(n237) );
  XOR U254 ( .A(n240), .B(n241), .Z(DIFF[242]) );
  XOR U255 ( .A(B[242]), .B(A[242]), .Z(n241) );
  AND U256 ( .A(n242), .B(n243), .Z(n240) );
  NANDN U257 ( .A(B[241]), .B(n244), .Z(n243) );
  NANDN U258 ( .A(A[241]), .B(n245), .Z(n244) );
  NANDN U259 ( .A(n245), .B(A[241]), .Z(n242) );
  XOR U260 ( .A(n245), .B(n246), .Z(DIFF[241]) );
  XOR U261 ( .A(B[241]), .B(A[241]), .Z(n246) );
  AND U262 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U263 ( .A(B[240]), .B(n249), .Z(n248) );
  NANDN U264 ( .A(A[240]), .B(n250), .Z(n249) );
  NANDN U265 ( .A(n250), .B(A[240]), .Z(n247) );
  XOR U266 ( .A(n250), .B(n251), .Z(DIFF[240]) );
  XOR U267 ( .A(B[240]), .B(A[240]), .Z(n251) );
  AND U268 ( .A(n252), .B(n253), .Z(n250) );
  NANDN U269 ( .A(B[239]), .B(n254), .Z(n253) );
  NANDN U270 ( .A(A[239]), .B(n255), .Z(n254) );
  NANDN U271 ( .A(n255), .B(A[239]), .Z(n252) );
  XOR U272 ( .A(n256), .B(n257), .Z(DIFF[23]) );
  XOR U273 ( .A(B[23]), .B(A[23]), .Z(n257) );
  XOR U274 ( .A(n255), .B(n258), .Z(DIFF[239]) );
  XOR U275 ( .A(B[239]), .B(A[239]), .Z(n258) );
  AND U276 ( .A(n259), .B(n260), .Z(n255) );
  NANDN U277 ( .A(B[238]), .B(n261), .Z(n260) );
  NANDN U278 ( .A(A[238]), .B(n262), .Z(n261) );
  NANDN U279 ( .A(n262), .B(A[238]), .Z(n259) );
  XOR U280 ( .A(n262), .B(n263), .Z(DIFF[238]) );
  XOR U281 ( .A(B[238]), .B(A[238]), .Z(n263) );
  AND U282 ( .A(n264), .B(n265), .Z(n262) );
  NANDN U283 ( .A(B[237]), .B(n266), .Z(n265) );
  NANDN U284 ( .A(A[237]), .B(n267), .Z(n266) );
  NANDN U285 ( .A(n267), .B(A[237]), .Z(n264) );
  XOR U286 ( .A(n267), .B(n268), .Z(DIFF[237]) );
  XOR U287 ( .A(B[237]), .B(A[237]), .Z(n268) );
  AND U288 ( .A(n269), .B(n270), .Z(n267) );
  NANDN U289 ( .A(B[236]), .B(n271), .Z(n270) );
  NANDN U290 ( .A(A[236]), .B(n272), .Z(n271) );
  NANDN U291 ( .A(n272), .B(A[236]), .Z(n269) );
  XOR U292 ( .A(n272), .B(n273), .Z(DIFF[236]) );
  XOR U293 ( .A(B[236]), .B(A[236]), .Z(n273) );
  AND U294 ( .A(n274), .B(n275), .Z(n272) );
  NANDN U295 ( .A(B[235]), .B(n276), .Z(n275) );
  NANDN U296 ( .A(A[235]), .B(n277), .Z(n276) );
  NANDN U297 ( .A(n277), .B(A[235]), .Z(n274) );
  XOR U298 ( .A(n277), .B(n278), .Z(DIFF[235]) );
  XOR U299 ( .A(B[235]), .B(A[235]), .Z(n278) );
  AND U300 ( .A(n279), .B(n280), .Z(n277) );
  NANDN U301 ( .A(B[234]), .B(n281), .Z(n280) );
  NANDN U302 ( .A(A[234]), .B(n282), .Z(n281) );
  NANDN U303 ( .A(n282), .B(A[234]), .Z(n279) );
  XOR U304 ( .A(n282), .B(n283), .Z(DIFF[234]) );
  XOR U305 ( .A(B[234]), .B(A[234]), .Z(n283) );
  AND U306 ( .A(n284), .B(n285), .Z(n282) );
  NANDN U307 ( .A(B[233]), .B(n286), .Z(n285) );
  NANDN U308 ( .A(A[233]), .B(n287), .Z(n286) );
  NANDN U309 ( .A(n287), .B(A[233]), .Z(n284) );
  XOR U310 ( .A(n287), .B(n288), .Z(DIFF[233]) );
  XOR U311 ( .A(B[233]), .B(A[233]), .Z(n288) );
  AND U312 ( .A(n289), .B(n290), .Z(n287) );
  NANDN U313 ( .A(B[232]), .B(n291), .Z(n290) );
  NANDN U314 ( .A(A[232]), .B(n292), .Z(n291) );
  NANDN U315 ( .A(n292), .B(A[232]), .Z(n289) );
  XOR U316 ( .A(n292), .B(n293), .Z(DIFF[232]) );
  XOR U317 ( .A(B[232]), .B(A[232]), .Z(n293) );
  AND U318 ( .A(n294), .B(n295), .Z(n292) );
  NANDN U319 ( .A(B[231]), .B(n296), .Z(n295) );
  NANDN U320 ( .A(A[231]), .B(n297), .Z(n296) );
  NANDN U321 ( .A(n297), .B(A[231]), .Z(n294) );
  XOR U322 ( .A(n297), .B(n298), .Z(DIFF[231]) );
  XOR U323 ( .A(B[231]), .B(A[231]), .Z(n298) );
  AND U324 ( .A(n299), .B(n300), .Z(n297) );
  NANDN U325 ( .A(B[230]), .B(n301), .Z(n300) );
  NANDN U326 ( .A(A[230]), .B(n302), .Z(n301) );
  NANDN U327 ( .A(n302), .B(A[230]), .Z(n299) );
  XOR U328 ( .A(n302), .B(n303), .Z(DIFF[230]) );
  XOR U329 ( .A(B[230]), .B(A[230]), .Z(n303) );
  AND U330 ( .A(n304), .B(n305), .Z(n302) );
  NANDN U331 ( .A(B[229]), .B(n306), .Z(n305) );
  NANDN U332 ( .A(A[229]), .B(n307), .Z(n306) );
  NANDN U333 ( .A(n307), .B(A[229]), .Z(n304) );
  XOR U334 ( .A(n308), .B(n309), .Z(DIFF[22]) );
  XOR U335 ( .A(B[22]), .B(A[22]), .Z(n309) );
  XOR U336 ( .A(n307), .B(n310), .Z(DIFF[229]) );
  XOR U337 ( .A(B[229]), .B(A[229]), .Z(n310) );
  AND U338 ( .A(n311), .B(n312), .Z(n307) );
  NANDN U339 ( .A(B[228]), .B(n313), .Z(n312) );
  NANDN U340 ( .A(A[228]), .B(n314), .Z(n313) );
  NANDN U341 ( .A(n314), .B(A[228]), .Z(n311) );
  XOR U342 ( .A(n314), .B(n315), .Z(DIFF[228]) );
  XOR U343 ( .A(B[228]), .B(A[228]), .Z(n315) );
  AND U344 ( .A(n316), .B(n317), .Z(n314) );
  NANDN U345 ( .A(B[227]), .B(n318), .Z(n317) );
  NANDN U346 ( .A(A[227]), .B(n319), .Z(n318) );
  NANDN U347 ( .A(n319), .B(A[227]), .Z(n316) );
  XOR U348 ( .A(n319), .B(n320), .Z(DIFF[227]) );
  XOR U349 ( .A(B[227]), .B(A[227]), .Z(n320) );
  AND U350 ( .A(n321), .B(n322), .Z(n319) );
  NANDN U351 ( .A(B[226]), .B(n323), .Z(n322) );
  NANDN U352 ( .A(A[226]), .B(n324), .Z(n323) );
  NANDN U353 ( .A(n324), .B(A[226]), .Z(n321) );
  XOR U354 ( .A(n324), .B(n325), .Z(DIFF[226]) );
  XOR U355 ( .A(B[226]), .B(A[226]), .Z(n325) );
  AND U356 ( .A(n326), .B(n327), .Z(n324) );
  NANDN U357 ( .A(B[225]), .B(n328), .Z(n327) );
  NANDN U358 ( .A(A[225]), .B(n329), .Z(n328) );
  NANDN U359 ( .A(n329), .B(A[225]), .Z(n326) );
  XOR U360 ( .A(n329), .B(n330), .Z(DIFF[225]) );
  XOR U361 ( .A(B[225]), .B(A[225]), .Z(n330) );
  AND U362 ( .A(n331), .B(n332), .Z(n329) );
  NANDN U363 ( .A(B[224]), .B(n333), .Z(n332) );
  NANDN U364 ( .A(A[224]), .B(n334), .Z(n333) );
  NANDN U365 ( .A(n334), .B(A[224]), .Z(n331) );
  XOR U366 ( .A(n334), .B(n335), .Z(DIFF[224]) );
  XOR U367 ( .A(B[224]), .B(A[224]), .Z(n335) );
  AND U368 ( .A(n336), .B(n337), .Z(n334) );
  NANDN U369 ( .A(B[223]), .B(n338), .Z(n337) );
  NANDN U370 ( .A(A[223]), .B(n339), .Z(n338) );
  NANDN U371 ( .A(n339), .B(A[223]), .Z(n336) );
  XOR U372 ( .A(n339), .B(n340), .Z(DIFF[223]) );
  XOR U373 ( .A(B[223]), .B(A[223]), .Z(n340) );
  AND U374 ( .A(n341), .B(n342), .Z(n339) );
  NANDN U375 ( .A(B[222]), .B(n343), .Z(n342) );
  NANDN U376 ( .A(A[222]), .B(n344), .Z(n343) );
  NANDN U377 ( .A(n344), .B(A[222]), .Z(n341) );
  XOR U378 ( .A(n344), .B(n345), .Z(DIFF[222]) );
  XOR U379 ( .A(B[222]), .B(A[222]), .Z(n345) );
  AND U380 ( .A(n346), .B(n347), .Z(n344) );
  NANDN U381 ( .A(B[221]), .B(n348), .Z(n347) );
  NANDN U382 ( .A(A[221]), .B(n349), .Z(n348) );
  NANDN U383 ( .A(n349), .B(A[221]), .Z(n346) );
  XOR U384 ( .A(n349), .B(n350), .Z(DIFF[221]) );
  XOR U385 ( .A(B[221]), .B(A[221]), .Z(n350) );
  AND U386 ( .A(n351), .B(n352), .Z(n349) );
  NANDN U387 ( .A(B[220]), .B(n353), .Z(n352) );
  NANDN U388 ( .A(A[220]), .B(n354), .Z(n353) );
  NANDN U389 ( .A(n354), .B(A[220]), .Z(n351) );
  XOR U390 ( .A(n354), .B(n355), .Z(DIFF[220]) );
  XOR U391 ( .A(B[220]), .B(A[220]), .Z(n355) );
  AND U392 ( .A(n356), .B(n357), .Z(n354) );
  NANDN U393 ( .A(B[219]), .B(n358), .Z(n357) );
  NANDN U394 ( .A(A[219]), .B(n359), .Z(n358) );
  NANDN U395 ( .A(n359), .B(A[219]), .Z(n356) );
  XOR U396 ( .A(n360), .B(n361), .Z(DIFF[21]) );
  XOR U397 ( .A(B[21]), .B(A[21]), .Z(n361) );
  XOR U398 ( .A(n359), .B(n362), .Z(DIFF[219]) );
  XOR U399 ( .A(B[219]), .B(A[219]), .Z(n362) );
  AND U400 ( .A(n363), .B(n364), .Z(n359) );
  NANDN U401 ( .A(B[218]), .B(n365), .Z(n364) );
  NANDN U402 ( .A(A[218]), .B(n366), .Z(n365) );
  NANDN U403 ( .A(n366), .B(A[218]), .Z(n363) );
  XOR U404 ( .A(n366), .B(n367), .Z(DIFF[218]) );
  XOR U405 ( .A(B[218]), .B(A[218]), .Z(n367) );
  AND U406 ( .A(n368), .B(n369), .Z(n366) );
  NANDN U407 ( .A(B[217]), .B(n370), .Z(n369) );
  NANDN U408 ( .A(A[217]), .B(n371), .Z(n370) );
  NANDN U409 ( .A(n371), .B(A[217]), .Z(n368) );
  XOR U410 ( .A(n371), .B(n372), .Z(DIFF[217]) );
  XOR U411 ( .A(B[217]), .B(A[217]), .Z(n372) );
  AND U412 ( .A(n373), .B(n374), .Z(n371) );
  NANDN U413 ( .A(B[216]), .B(n375), .Z(n374) );
  NANDN U414 ( .A(A[216]), .B(n376), .Z(n375) );
  NANDN U415 ( .A(n376), .B(A[216]), .Z(n373) );
  XOR U416 ( .A(n376), .B(n377), .Z(DIFF[216]) );
  XOR U417 ( .A(B[216]), .B(A[216]), .Z(n377) );
  AND U418 ( .A(n378), .B(n379), .Z(n376) );
  NANDN U419 ( .A(B[215]), .B(n380), .Z(n379) );
  NANDN U420 ( .A(A[215]), .B(n381), .Z(n380) );
  NANDN U421 ( .A(n381), .B(A[215]), .Z(n378) );
  XOR U422 ( .A(n381), .B(n382), .Z(DIFF[215]) );
  XOR U423 ( .A(B[215]), .B(A[215]), .Z(n382) );
  AND U424 ( .A(n383), .B(n384), .Z(n381) );
  NANDN U425 ( .A(B[214]), .B(n385), .Z(n384) );
  NANDN U426 ( .A(A[214]), .B(n386), .Z(n385) );
  NANDN U427 ( .A(n386), .B(A[214]), .Z(n383) );
  XOR U428 ( .A(n386), .B(n387), .Z(DIFF[214]) );
  XOR U429 ( .A(B[214]), .B(A[214]), .Z(n387) );
  AND U430 ( .A(n388), .B(n389), .Z(n386) );
  NANDN U431 ( .A(B[213]), .B(n390), .Z(n389) );
  NANDN U432 ( .A(A[213]), .B(n391), .Z(n390) );
  NANDN U433 ( .A(n391), .B(A[213]), .Z(n388) );
  XOR U434 ( .A(n391), .B(n392), .Z(DIFF[213]) );
  XOR U435 ( .A(B[213]), .B(A[213]), .Z(n392) );
  AND U436 ( .A(n393), .B(n394), .Z(n391) );
  NANDN U437 ( .A(B[212]), .B(n395), .Z(n394) );
  NANDN U438 ( .A(A[212]), .B(n396), .Z(n395) );
  NANDN U439 ( .A(n396), .B(A[212]), .Z(n393) );
  XOR U440 ( .A(n396), .B(n397), .Z(DIFF[212]) );
  XOR U441 ( .A(B[212]), .B(A[212]), .Z(n397) );
  AND U442 ( .A(n398), .B(n399), .Z(n396) );
  NANDN U443 ( .A(B[211]), .B(n400), .Z(n399) );
  NANDN U444 ( .A(A[211]), .B(n401), .Z(n400) );
  NANDN U445 ( .A(n401), .B(A[211]), .Z(n398) );
  XOR U446 ( .A(n401), .B(n402), .Z(DIFF[211]) );
  XOR U447 ( .A(B[211]), .B(A[211]), .Z(n402) );
  AND U448 ( .A(n403), .B(n404), .Z(n401) );
  NANDN U449 ( .A(B[210]), .B(n405), .Z(n404) );
  NANDN U450 ( .A(A[210]), .B(n406), .Z(n405) );
  NANDN U451 ( .A(n406), .B(A[210]), .Z(n403) );
  XOR U452 ( .A(n406), .B(n407), .Z(DIFF[210]) );
  XOR U453 ( .A(B[210]), .B(A[210]), .Z(n407) );
  AND U454 ( .A(n408), .B(n409), .Z(n406) );
  NANDN U455 ( .A(B[209]), .B(n410), .Z(n409) );
  NANDN U456 ( .A(A[209]), .B(n411), .Z(n410) );
  NANDN U457 ( .A(n411), .B(A[209]), .Z(n408) );
  XOR U458 ( .A(n412), .B(n413), .Z(DIFF[20]) );
  XOR U459 ( .A(B[20]), .B(A[20]), .Z(n413) );
  XOR U460 ( .A(n411), .B(n414), .Z(DIFF[209]) );
  XOR U461 ( .A(B[209]), .B(A[209]), .Z(n414) );
  AND U462 ( .A(n415), .B(n416), .Z(n411) );
  NANDN U463 ( .A(B[208]), .B(n417), .Z(n416) );
  NANDN U464 ( .A(A[208]), .B(n418), .Z(n417) );
  NANDN U465 ( .A(n418), .B(A[208]), .Z(n415) );
  XOR U466 ( .A(n418), .B(n419), .Z(DIFF[208]) );
  XOR U467 ( .A(B[208]), .B(A[208]), .Z(n419) );
  AND U468 ( .A(n420), .B(n421), .Z(n418) );
  NANDN U469 ( .A(B[207]), .B(n422), .Z(n421) );
  NANDN U470 ( .A(A[207]), .B(n423), .Z(n422) );
  NANDN U471 ( .A(n423), .B(A[207]), .Z(n420) );
  XOR U472 ( .A(n423), .B(n424), .Z(DIFF[207]) );
  XOR U473 ( .A(B[207]), .B(A[207]), .Z(n424) );
  AND U474 ( .A(n425), .B(n426), .Z(n423) );
  NANDN U475 ( .A(B[206]), .B(n427), .Z(n426) );
  NANDN U476 ( .A(A[206]), .B(n428), .Z(n427) );
  NANDN U477 ( .A(n428), .B(A[206]), .Z(n425) );
  XOR U478 ( .A(n428), .B(n429), .Z(DIFF[206]) );
  XOR U479 ( .A(B[206]), .B(A[206]), .Z(n429) );
  AND U480 ( .A(n430), .B(n431), .Z(n428) );
  NANDN U481 ( .A(B[205]), .B(n432), .Z(n431) );
  NANDN U482 ( .A(A[205]), .B(n433), .Z(n432) );
  NANDN U483 ( .A(n433), .B(A[205]), .Z(n430) );
  XOR U484 ( .A(n433), .B(n434), .Z(DIFF[205]) );
  XOR U485 ( .A(B[205]), .B(A[205]), .Z(n434) );
  AND U486 ( .A(n435), .B(n436), .Z(n433) );
  NANDN U487 ( .A(B[204]), .B(n437), .Z(n436) );
  NANDN U488 ( .A(A[204]), .B(n438), .Z(n437) );
  NANDN U489 ( .A(n438), .B(A[204]), .Z(n435) );
  XOR U490 ( .A(n438), .B(n439), .Z(DIFF[204]) );
  XOR U491 ( .A(B[204]), .B(A[204]), .Z(n439) );
  AND U492 ( .A(n440), .B(n441), .Z(n438) );
  NANDN U493 ( .A(B[203]), .B(n442), .Z(n441) );
  NANDN U494 ( .A(A[203]), .B(n443), .Z(n442) );
  NANDN U495 ( .A(n443), .B(A[203]), .Z(n440) );
  XOR U496 ( .A(n443), .B(n444), .Z(DIFF[203]) );
  XOR U497 ( .A(B[203]), .B(A[203]), .Z(n444) );
  AND U498 ( .A(n445), .B(n446), .Z(n443) );
  NANDN U499 ( .A(B[202]), .B(n447), .Z(n446) );
  NANDN U500 ( .A(A[202]), .B(n448), .Z(n447) );
  NANDN U501 ( .A(n448), .B(A[202]), .Z(n445) );
  XOR U502 ( .A(n448), .B(n449), .Z(DIFF[202]) );
  XOR U503 ( .A(B[202]), .B(A[202]), .Z(n449) );
  AND U504 ( .A(n450), .B(n451), .Z(n448) );
  NANDN U505 ( .A(B[201]), .B(n452), .Z(n451) );
  NANDN U506 ( .A(A[201]), .B(n453), .Z(n452) );
  NANDN U507 ( .A(n453), .B(A[201]), .Z(n450) );
  XOR U508 ( .A(n453), .B(n454), .Z(DIFF[201]) );
  XOR U509 ( .A(B[201]), .B(A[201]), .Z(n454) );
  AND U510 ( .A(n455), .B(n456), .Z(n453) );
  NANDN U511 ( .A(B[200]), .B(n457), .Z(n456) );
  NANDN U512 ( .A(A[200]), .B(n458), .Z(n457) );
  NANDN U513 ( .A(n458), .B(A[200]), .Z(n455) );
  XOR U514 ( .A(n458), .B(n459), .Z(DIFF[200]) );
  XOR U515 ( .A(B[200]), .B(A[200]), .Z(n459) );
  AND U516 ( .A(n460), .B(n461), .Z(n458) );
  NANDN U517 ( .A(B[199]), .B(n462), .Z(n461) );
  NANDN U518 ( .A(A[199]), .B(n463), .Z(n462) );
  NANDN U519 ( .A(n463), .B(A[199]), .Z(n460) );
  XOR U520 ( .A(n1), .B(n464), .Z(DIFF[1]) );
  XOR U521 ( .A(B[1]), .B(A[1]), .Z(n464) );
  XOR U522 ( .A(n465), .B(n466), .Z(DIFF[19]) );
  XOR U523 ( .A(B[19]), .B(A[19]), .Z(n466) );
  XOR U524 ( .A(n463), .B(n467), .Z(DIFF[199]) );
  XOR U525 ( .A(B[199]), .B(A[199]), .Z(n467) );
  AND U526 ( .A(n468), .B(n469), .Z(n463) );
  NANDN U527 ( .A(B[198]), .B(n470), .Z(n469) );
  NANDN U528 ( .A(A[198]), .B(n471), .Z(n470) );
  NANDN U529 ( .A(n471), .B(A[198]), .Z(n468) );
  XOR U530 ( .A(n471), .B(n472), .Z(DIFF[198]) );
  XOR U531 ( .A(B[198]), .B(A[198]), .Z(n472) );
  AND U532 ( .A(n473), .B(n474), .Z(n471) );
  NANDN U533 ( .A(B[197]), .B(n475), .Z(n474) );
  NANDN U534 ( .A(A[197]), .B(n476), .Z(n475) );
  NANDN U535 ( .A(n476), .B(A[197]), .Z(n473) );
  XOR U536 ( .A(n476), .B(n477), .Z(DIFF[197]) );
  XOR U537 ( .A(B[197]), .B(A[197]), .Z(n477) );
  AND U538 ( .A(n478), .B(n479), .Z(n476) );
  NANDN U539 ( .A(B[196]), .B(n480), .Z(n479) );
  NANDN U540 ( .A(A[196]), .B(n481), .Z(n480) );
  NANDN U541 ( .A(n481), .B(A[196]), .Z(n478) );
  XOR U542 ( .A(n481), .B(n482), .Z(DIFF[196]) );
  XOR U543 ( .A(B[196]), .B(A[196]), .Z(n482) );
  AND U544 ( .A(n483), .B(n484), .Z(n481) );
  NANDN U545 ( .A(B[195]), .B(n485), .Z(n484) );
  NANDN U546 ( .A(A[195]), .B(n486), .Z(n485) );
  NANDN U547 ( .A(n486), .B(A[195]), .Z(n483) );
  XOR U548 ( .A(n486), .B(n487), .Z(DIFF[195]) );
  XOR U549 ( .A(B[195]), .B(A[195]), .Z(n487) );
  AND U550 ( .A(n488), .B(n489), .Z(n486) );
  NANDN U551 ( .A(B[194]), .B(n490), .Z(n489) );
  NANDN U552 ( .A(A[194]), .B(n491), .Z(n490) );
  NANDN U553 ( .A(n491), .B(A[194]), .Z(n488) );
  XOR U554 ( .A(n491), .B(n492), .Z(DIFF[194]) );
  XOR U555 ( .A(B[194]), .B(A[194]), .Z(n492) );
  AND U556 ( .A(n493), .B(n494), .Z(n491) );
  NANDN U557 ( .A(B[193]), .B(n495), .Z(n494) );
  NANDN U558 ( .A(A[193]), .B(n496), .Z(n495) );
  NANDN U559 ( .A(n496), .B(A[193]), .Z(n493) );
  XOR U560 ( .A(n496), .B(n497), .Z(DIFF[193]) );
  XOR U561 ( .A(B[193]), .B(A[193]), .Z(n497) );
  AND U562 ( .A(n498), .B(n499), .Z(n496) );
  NANDN U563 ( .A(B[192]), .B(n500), .Z(n499) );
  NANDN U564 ( .A(A[192]), .B(n501), .Z(n500) );
  NANDN U565 ( .A(n501), .B(A[192]), .Z(n498) );
  XOR U566 ( .A(n501), .B(n502), .Z(DIFF[192]) );
  XOR U567 ( .A(B[192]), .B(A[192]), .Z(n502) );
  AND U568 ( .A(n503), .B(n504), .Z(n501) );
  NANDN U569 ( .A(B[191]), .B(n505), .Z(n504) );
  NANDN U570 ( .A(A[191]), .B(n506), .Z(n505) );
  NANDN U571 ( .A(n506), .B(A[191]), .Z(n503) );
  XOR U572 ( .A(n506), .B(n507), .Z(DIFF[191]) );
  XOR U573 ( .A(B[191]), .B(A[191]), .Z(n507) );
  AND U574 ( .A(n508), .B(n509), .Z(n506) );
  NANDN U575 ( .A(B[190]), .B(n510), .Z(n509) );
  NANDN U576 ( .A(A[190]), .B(n511), .Z(n510) );
  NANDN U577 ( .A(n511), .B(A[190]), .Z(n508) );
  XOR U578 ( .A(n511), .B(n512), .Z(DIFF[190]) );
  XOR U579 ( .A(B[190]), .B(A[190]), .Z(n512) );
  AND U580 ( .A(n513), .B(n514), .Z(n511) );
  NANDN U581 ( .A(B[189]), .B(n515), .Z(n514) );
  NANDN U582 ( .A(A[189]), .B(n516), .Z(n515) );
  NANDN U583 ( .A(n516), .B(A[189]), .Z(n513) );
  XOR U584 ( .A(n517), .B(n518), .Z(DIFF[18]) );
  XOR U585 ( .A(B[18]), .B(A[18]), .Z(n518) );
  XOR U586 ( .A(n516), .B(n519), .Z(DIFF[189]) );
  XOR U587 ( .A(B[189]), .B(A[189]), .Z(n519) );
  AND U588 ( .A(n520), .B(n521), .Z(n516) );
  NANDN U589 ( .A(B[188]), .B(n522), .Z(n521) );
  NANDN U590 ( .A(A[188]), .B(n523), .Z(n522) );
  NANDN U591 ( .A(n523), .B(A[188]), .Z(n520) );
  XOR U592 ( .A(n523), .B(n524), .Z(DIFF[188]) );
  XOR U593 ( .A(B[188]), .B(A[188]), .Z(n524) );
  AND U594 ( .A(n525), .B(n526), .Z(n523) );
  NANDN U595 ( .A(B[187]), .B(n527), .Z(n526) );
  NANDN U596 ( .A(A[187]), .B(n528), .Z(n527) );
  NANDN U597 ( .A(n528), .B(A[187]), .Z(n525) );
  XOR U598 ( .A(n528), .B(n529), .Z(DIFF[187]) );
  XOR U599 ( .A(B[187]), .B(A[187]), .Z(n529) );
  AND U600 ( .A(n530), .B(n531), .Z(n528) );
  NANDN U601 ( .A(B[186]), .B(n532), .Z(n531) );
  NANDN U602 ( .A(A[186]), .B(n533), .Z(n532) );
  NANDN U603 ( .A(n533), .B(A[186]), .Z(n530) );
  XOR U604 ( .A(n533), .B(n534), .Z(DIFF[186]) );
  XOR U605 ( .A(B[186]), .B(A[186]), .Z(n534) );
  AND U606 ( .A(n535), .B(n536), .Z(n533) );
  NANDN U607 ( .A(B[185]), .B(n537), .Z(n536) );
  NANDN U608 ( .A(A[185]), .B(n538), .Z(n537) );
  NANDN U609 ( .A(n538), .B(A[185]), .Z(n535) );
  XOR U610 ( .A(n538), .B(n539), .Z(DIFF[185]) );
  XOR U611 ( .A(B[185]), .B(A[185]), .Z(n539) );
  AND U612 ( .A(n540), .B(n541), .Z(n538) );
  NANDN U613 ( .A(B[184]), .B(n542), .Z(n541) );
  NANDN U614 ( .A(A[184]), .B(n543), .Z(n542) );
  NANDN U615 ( .A(n543), .B(A[184]), .Z(n540) );
  XOR U616 ( .A(n543), .B(n544), .Z(DIFF[184]) );
  XOR U617 ( .A(B[184]), .B(A[184]), .Z(n544) );
  AND U618 ( .A(n545), .B(n546), .Z(n543) );
  NANDN U619 ( .A(B[183]), .B(n547), .Z(n546) );
  NANDN U620 ( .A(A[183]), .B(n548), .Z(n547) );
  NANDN U621 ( .A(n548), .B(A[183]), .Z(n545) );
  XOR U622 ( .A(n548), .B(n549), .Z(DIFF[183]) );
  XOR U623 ( .A(B[183]), .B(A[183]), .Z(n549) );
  AND U624 ( .A(n550), .B(n551), .Z(n548) );
  NANDN U625 ( .A(B[182]), .B(n552), .Z(n551) );
  NANDN U626 ( .A(A[182]), .B(n553), .Z(n552) );
  NANDN U627 ( .A(n553), .B(A[182]), .Z(n550) );
  XOR U628 ( .A(n553), .B(n554), .Z(DIFF[182]) );
  XOR U629 ( .A(B[182]), .B(A[182]), .Z(n554) );
  AND U630 ( .A(n555), .B(n556), .Z(n553) );
  NANDN U631 ( .A(B[181]), .B(n557), .Z(n556) );
  NANDN U632 ( .A(A[181]), .B(n558), .Z(n557) );
  NANDN U633 ( .A(n558), .B(A[181]), .Z(n555) );
  XOR U634 ( .A(n558), .B(n559), .Z(DIFF[181]) );
  XOR U635 ( .A(B[181]), .B(A[181]), .Z(n559) );
  AND U636 ( .A(n560), .B(n561), .Z(n558) );
  NANDN U637 ( .A(B[180]), .B(n562), .Z(n561) );
  NANDN U638 ( .A(A[180]), .B(n563), .Z(n562) );
  NANDN U639 ( .A(n563), .B(A[180]), .Z(n560) );
  XOR U640 ( .A(n563), .B(n564), .Z(DIFF[180]) );
  XOR U641 ( .A(B[180]), .B(A[180]), .Z(n564) );
  AND U642 ( .A(n565), .B(n566), .Z(n563) );
  NANDN U643 ( .A(B[179]), .B(n567), .Z(n566) );
  NANDN U644 ( .A(A[179]), .B(n568), .Z(n567) );
  NANDN U645 ( .A(n568), .B(A[179]), .Z(n565) );
  XOR U646 ( .A(n569), .B(n570), .Z(DIFF[17]) );
  XOR U647 ( .A(B[17]), .B(A[17]), .Z(n570) );
  XOR U648 ( .A(n568), .B(n571), .Z(DIFF[179]) );
  XOR U649 ( .A(B[179]), .B(A[179]), .Z(n571) );
  AND U650 ( .A(n572), .B(n573), .Z(n568) );
  NANDN U651 ( .A(B[178]), .B(n574), .Z(n573) );
  NANDN U652 ( .A(A[178]), .B(n575), .Z(n574) );
  NANDN U653 ( .A(n575), .B(A[178]), .Z(n572) );
  XOR U654 ( .A(n575), .B(n576), .Z(DIFF[178]) );
  XOR U655 ( .A(B[178]), .B(A[178]), .Z(n576) );
  AND U656 ( .A(n577), .B(n578), .Z(n575) );
  NANDN U657 ( .A(B[177]), .B(n579), .Z(n578) );
  NANDN U658 ( .A(A[177]), .B(n580), .Z(n579) );
  NANDN U659 ( .A(n580), .B(A[177]), .Z(n577) );
  XOR U660 ( .A(n580), .B(n581), .Z(DIFF[177]) );
  XOR U661 ( .A(B[177]), .B(A[177]), .Z(n581) );
  AND U662 ( .A(n582), .B(n583), .Z(n580) );
  NANDN U663 ( .A(B[176]), .B(n584), .Z(n583) );
  NANDN U664 ( .A(A[176]), .B(n585), .Z(n584) );
  NANDN U665 ( .A(n585), .B(A[176]), .Z(n582) );
  XOR U666 ( .A(n585), .B(n586), .Z(DIFF[176]) );
  XOR U667 ( .A(B[176]), .B(A[176]), .Z(n586) );
  AND U668 ( .A(n587), .B(n588), .Z(n585) );
  NANDN U669 ( .A(B[175]), .B(n589), .Z(n588) );
  NANDN U670 ( .A(A[175]), .B(n590), .Z(n589) );
  NANDN U671 ( .A(n590), .B(A[175]), .Z(n587) );
  XOR U672 ( .A(n590), .B(n591), .Z(DIFF[175]) );
  XOR U673 ( .A(B[175]), .B(A[175]), .Z(n591) );
  AND U674 ( .A(n592), .B(n593), .Z(n590) );
  NANDN U675 ( .A(B[174]), .B(n594), .Z(n593) );
  NANDN U676 ( .A(A[174]), .B(n595), .Z(n594) );
  NANDN U677 ( .A(n595), .B(A[174]), .Z(n592) );
  XOR U678 ( .A(n595), .B(n596), .Z(DIFF[174]) );
  XOR U679 ( .A(B[174]), .B(A[174]), .Z(n596) );
  AND U680 ( .A(n597), .B(n598), .Z(n595) );
  NANDN U681 ( .A(B[173]), .B(n599), .Z(n598) );
  NANDN U682 ( .A(A[173]), .B(n600), .Z(n599) );
  NANDN U683 ( .A(n600), .B(A[173]), .Z(n597) );
  XOR U684 ( .A(n600), .B(n601), .Z(DIFF[173]) );
  XOR U685 ( .A(B[173]), .B(A[173]), .Z(n601) );
  AND U686 ( .A(n602), .B(n603), .Z(n600) );
  NANDN U687 ( .A(B[172]), .B(n604), .Z(n603) );
  NANDN U688 ( .A(A[172]), .B(n605), .Z(n604) );
  NANDN U689 ( .A(n605), .B(A[172]), .Z(n602) );
  XOR U690 ( .A(n605), .B(n606), .Z(DIFF[172]) );
  XOR U691 ( .A(B[172]), .B(A[172]), .Z(n606) );
  AND U692 ( .A(n607), .B(n608), .Z(n605) );
  NANDN U693 ( .A(B[171]), .B(n609), .Z(n608) );
  NANDN U694 ( .A(A[171]), .B(n610), .Z(n609) );
  NANDN U695 ( .A(n610), .B(A[171]), .Z(n607) );
  XOR U696 ( .A(n610), .B(n611), .Z(DIFF[171]) );
  XOR U697 ( .A(B[171]), .B(A[171]), .Z(n611) );
  AND U698 ( .A(n612), .B(n613), .Z(n610) );
  NANDN U699 ( .A(B[170]), .B(n614), .Z(n613) );
  NANDN U700 ( .A(A[170]), .B(n615), .Z(n614) );
  NANDN U701 ( .A(n615), .B(A[170]), .Z(n612) );
  XOR U702 ( .A(n615), .B(n616), .Z(DIFF[170]) );
  XOR U703 ( .A(B[170]), .B(A[170]), .Z(n616) );
  AND U704 ( .A(n617), .B(n618), .Z(n615) );
  NANDN U705 ( .A(B[169]), .B(n619), .Z(n618) );
  NANDN U706 ( .A(A[169]), .B(n620), .Z(n619) );
  NANDN U707 ( .A(n620), .B(A[169]), .Z(n617) );
  XOR U708 ( .A(n621), .B(n622), .Z(DIFF[16]) );
  XOR U709 ( .A(B[16]), .B(A[16]), .Z(n622) );
  XOR U710 ( .A(n620), .B(n623), .Z(DIFF[169]) );
  XOR U711 ( .A(B[169]), .B(A[169]), .Z(n623) );
  AND U712 ( .A(n624), .B(n625), .Z(n620) );
  NANDN U713 ( .A(B[168]), .B(n626), .Z(n625) );
  NANDN U714 ( .A(A[168]), .B(n627), .Z(n626) );
  NANDN U715 ( .A(n627), .B(A[168]), .Z(n624) );
  XOR U716 ( .A(n627), .B(n628), .Z(DIFF[168]) );
  XOR U717 ( .A(B[168]), .B(A[168]), .Z(n628) );
  AND U718 ( .A(n629), .B(n630), .Z(n627) );
  NANDN U719 ( .A(B[167]), .B(n631), .Z(n630) );
  NANDN U720 ( .A(A[167]), .B(n632), .Z(n631) );
  NANDN U721 ( .A(n632), .B(A[167]), .Z(n629) );
  XOR U722 ( .A(n632), .B(n633), .Z(DIFF[167]) );
  XOR U723 ( .A(B[167]), .B(A[167]), .Z(n633) );
  AND U724 ( .A(n634), .B(n635), .Z(n632) );
  NANDN U725 ( .A(B[166]), .B(n636), .Z(n635) );
  NANDN U726 ( .A(A[166]), .B(n637), .Z(n636) );
  NANDN U727 ( .A(n637), .B(A[166]), .Z(n634) );
  XOR U728 ( .A(n637), .B(n638), .Z(DIFF[166]) );
  XOR U729 ( .A(B[166]), .B(A[166]), .Z(n638) );
  AND U730 ( .A(n639), .B(n640), .Z(n637) );
  NANDN U731 ( .A(B[165]), .B(n641), .Z(n640) );
  NANDN U732 ( .A(A[165]), .B(n642), .Z(n641) );
  NANDN U733 ( .A(n642), .B(A[165]), .Z(n639) );
  XOR U734 ( .A(n642), .B(n643), .Z(DIFF[165]) );
  XOR U735 ( .A(B[165]), .B(A[165]), .Z(n643) );
  AND U736 ( .A(n644), .B(n645), .Z(n642) );
  NANDN U737 ( .A(B[164]), .B(n646), .Z(n645) );
  NANDN U738 ( .A(A[164]), .B(n647), .Z(n646) );
  NANDN U739 ( .A(n647), .B(A[164]), .Z(n644) );
  XOR U740 ( .A(n647), .B(n648), .Z(DIFF[164]) );
  XOR U741 ( .A(B[164]), .B(A[164]), .Z(n648) );
  AND U742 ( .A(n649), .B(n650), .Z(n647) );
  NANDN U743 ( .A(B[163]), .B(n651), .Z(n650) );
  NANDN U744 ( .A(A[163]), .B(n652), .Z(n651) );
  NANDN U745 ( .A(n652), .B(A[163]), .Z(n649) );
  XOR U746 ( .A(n652), .B(n653), .Z(DIFF[163]) );
  XOR U747 ( .A(B[163]), .B(A[163]), .Z(n653) );
  AND U748 ( .A(n654), .B(n655), .Z(n652) );
  NANDN U749 ( .A(B[162]), .B(n656), .Z(n655) );
  NANDN U750 ( .A(A[162]), .B(n657), .Z(n656) );
  NANDN U751 ( .A(n657), .B(A[162]), .Z(n654) );
  XOR U752 ( .A(n657), .B(n658), .Z(DIFF[162]) );
  XOR U753 ( .A(B[162]), .B(A[162]), .Z(n658) );
  AND U754 ( .A(n659), .B(n660), .Z(n657) );
  NANDN U755 ( .A(B[161]), .B(n661), .Z(n660) );
  NANDN U756 ( .A(A[161]), .B(n662), .Z(n661) );
  NANDN U757 ( .A(n662), .B(A[161]), .Z(n659) );
  XOR U758 ( .A(n662), .B(n663), .Z(DIFF[161]) );
  XOR U759 ( .A(B[161]), .B(A[161]), .Z(n663) );
  AND U760 ( .A(n664), .B(n665), .Z(n662) );
  NANDN U761 ( .A(B[160]), .B(n666), .Z(n665) );
  NANDN U762 ( .A(A[160]), .B(n667), .Z(n666) );
  NANDN U763 ( .A(n667), .B(A[160]), .Z(n664) );
  XOR U764 ( .A(n667), .B(n668), .Z(DIFF[160]) );
  XOR U765 ( .A(B[160]), .B(A[160]), .Z(n668) );
  AND U766 ( .A(n669), .B(n670), .Z(n667) );
  NANDN U767 ( .A(B[159]), .B(n671), .Z(n670) );
  NANDN U768 ( .A(A[159]), .B(n672), .Z(n671) );
  NANDN U769 ( .A(n672), .B(A[159]), .Z(n669) );
  XOR U770 ( .A(n673), .B(n674), .Z(DIFF[15]) );
  XOR U771 ( .A(B[15]), .B(A[15]), .Z(n674) );
  XOR U772 ( .A(n672), .B(n675), .Z(DIFF[159]) );
  XOR U773 ( .A(B[159]), .B(A[159]), .Z(n675) );
  AND U774 ( .A(n676), .B(n677), .Z(n672) );
  NANDN U775 ( .A(B[158]), .B(n678), .Z(n677) );
  NANDN U776 ( .A(A[158]), .B(n679), .Z(n678) );
  NANDN U777 ( .A(n679), .B(A[158]), .Z(n676) );
  XOR U778 ( .A(n679), .B(n680), .Z(DIFF[158]) );
  XOR U779 ( .A(B[158]), .B(A[158]), .Z(n680) );
  AND U780 ( .A(n681), .B(n682), .Z(n679) );
  NANDN U781 ( .A(B[157]), .B(n683), .Z(n682) );
  NANDN U782 ( .A(A[157]), .B(n684), .Z(n683) );
  NANDN U783 ( .A(n684), .B(A[157]), .Z(n681) );
  XOR U784 ( .A(n684), .B(n685), .Z(DIFF[157]) );
  XOR U785 ( .A(B[157]), .B(A[157]), .Z(n685) );
  AND U786 ( .A(n686), .B(n687), .Z(n684) );
  NANDN U787 ( .A(B[156]), .B(n688), .Z(n687) );
  NANDN U788 ( .A(A[156]), .B(n689), .Z(n688) );
  NANDN U789 ( .A(n689), .B(A[156]), .Z(n686) );
  XOR U790 ( .A(n689), .B(n690), .Z(DIFF[156]) );
  XOR U791 ( .A(B[156]), .B(A[156]), .Z(n690) );
  AND U792 ( .A(n691), .B(n692), .Z(n689) );
  NANDN U793 ( .A(B[155]), .B(n693), .Z(n692) );
  NANDN U794 ( .A(A[155]), .B(n694), .Z(n693) );
  NANDN U795 ( .A(n694), .B(A[155]), .Z(n691) );
  XOR U796 ( .A(n694), .B(n695), .Z(DIFF[155]) );
  XOR U797 ( .A(B[155]), .B(A[155]), .Z(n695) );
  AND U798 ( .A(n696), .B(n697), .Z(n694) );
  NANDN U799 ( .A(B[154]), .B(n698), .Z(n697) );
  NANDN U800 ( .A(A[154]), .B(n699), .Z(n698) );
  NANDN U801 ( .A(n699), .B(A[154]), .Z(n696) );
  XOR U802 ( .A(n699), .B(n700), .Z(DIFF[154]) );
  XOR U803 ( .A(B[154]), .B(A[154]), .Z(n700) );
  AND U804 ( .A(n701), .B(n702), .Z(n699) );
  NANDN U805 ( .A(B[153]), .B(n703), .Z(n702) );
  NANDN U806 ( .A(A[153]), .B(n704), .Z(n703) );
  NANDN U807 ( .A(n704), .B(A[153]), .Z(n701) );
  XOR U808 ( .A(n704), .B(n705), .Z(DIFF[153]) );
  XOR U809 ( .A(B[153]), .B(A[153]), .Z(n705) );
  AND U810 ( .A(n706), .B(n707), .Z(n704) );
  NANDN U811 ( .A(B[152]), .B(n708), .Z(n707) );
  NANDN U812 ( .A(A[152]), .B(n709), .Z(n708) );
  NANDN U813 ( .A(n709), .B(A[152]), .Z(n706) );
  XOR U814 ( .A(n709), .B(n710), .Z(DIFF[152]) );
  XOR U815 ( .A(B[152]), .B(A[152]), .Z(n710) );
  AND U816 ( .A(n711), .B(n712), .Z(n709) );
  NANDN U817 ( .A(B[151]), .B(n713), .Z(n712) );
  NANDN U818 ( .A(A[151]), .B(n714), .Z(n713) );
  NANDN U819 ( .A(n714), .B(A[151]), .Z(n711) );
  XOR U820 ( .A(n714), .B(n715), .Z(DIFF[151]) );
  XOR U821 ( .A(B[151]), .B(A[151]), .Z(n715) );
  AND U822 ( .A(n716), .B(n717), .Z(n714) );
  NANDN U823 ( .A(B[150]), .B(n718), .Z(n717) );
  NANDN U824 ( .A(A[150]), .B(n719), .Z(n718) );
  NANDN U825 ( .A(n719), .B(A[150]), .Z(n716) );
  XOR U826 ( .A(n719), .B(n720), .Z(DIFF[150]) );
  XOR U827 ( .A(B[150]), .B(A[150]), .Z(n720) );
  AND U828 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U829 ( .A(B[149]), .B(n723), .Z(n722) );
  NANDN U830 ( .A(A[149]), .B(n724), .Z(n723) );
  NANDN U831 ( .A(n724), .B(A[149]), .Z(n721) );
  XOR U832 ( .A(n725), .B(n726), .Z(DIFF[14]) );
  XOR U833 ( .A(B[14]), .B(A[14]), .Z(n726) );
  XOR U834 ( .A(n724), .B(n727), .Z(DIFF[149]) );
  XOR U835 ( .A(B[149]), .B(A[149]), .Z(n727) );
  AND U836 ( .A(n728), .B(n729), .Z(n724) );
  NANDN U837 ( .A(B[148]), .B(n730), .Z(n729) );
  NANDN U838 ( .A(A[148]), .B(n731), .Z(n730) );
  NANDN U839 ( .A(n731), .B(A[148]), .Z(n728) );
  XOR U840 ( .A(n731), .B(n732), .Z(DIFF[148]) );
  XOR U841 ( .A(B[148]), .B(A[148]), .Z(n732) );
  AND U842 ( .A(n733), .B(n734), .Z(n731) );
  NANDN U843 ( .A(B[147]), .B(n735), .Z(n734) );
  NANDN U844 ( .A(A[147]), .B(n736), .Z(n735) );
  NANDN U845 ( .A(n736), .B(A[147]), .Z(n733) );
  XOR U846 ( .A(n736), .B(n737), .Z(DIFF[147]) );
  XOR U847 ( .A(B[147]), .B(A[147]), .Z(n737) );
  AND U848 ( .A(n738), .B(n739), .Z(n736) );
  NANDN U849 ( .A(B[146]), .B(n740), .Z(n739) );
  NANDN U850 ( .A(A[146]), .B(n741), .Z(n740) );
  NANDN U851 ( .A(n741), .B(A[146]), .Z(n738) );
  XOR U852 ( .A(n741), .B(n742), .Z(DIFF[146]) );
  XOR U853 ( .A(B[146]), .B(A[146]), .Z(n742) );
  AND U854 ( .A(n743), .B(n744), .Z(n741) );
  NANDN U855 ( .A(B[145]), .B(n745), .Z(n744) );
  NANDN U856 ( .A(A[145]), .B(n746), .Z(n745) );
  NANDN U857 ( .A(n746), .B(A[145]), .Z(n743) );
  XOR U858 ( .A(n746), .B(n747), .Z(DIFF[145]) );
  XOR U859 ( .A(B[145]), .B(A[145]), .Z(n747) );
  AND U860 ( .A(n748), .B(n749), .Z(n746) );
  NANDN U861 ( .A(B[144]), .B(n750), .Z(n749) );
  NANDN U862 ( .A(A[144]), .B(n751), .Z(n750) );
  NANDN U863 ( .A(n751), .B(A[144]), .Z(n748) );
  XOR U864 ( .A(n751), .B(n752), .Z(DIFF[144]) );
  XOR U865 ( .A(B[144]), .B(A[144]), .Z(n752) );
  AND U866 ( .A(n753), .B(n754), .Z(n751) );
  NANDN U867 ( .A(B[143]), .B(n755), .Z(n754) );
  NANDN U868 ( .A(A[143]), .B(n756), .Z(n755) );
  NANDN U869 ( .A(n756), .B(A[143]), .Z(n753) );
  XOR U870 ( .A(n756), .B(n757), .Z(DIFF[143]) );
  XOR U871 ( .A(B[143]), .B(A[143]), .Z(n757) );
  AND U872 ( .A(n758), .B(n759), .Z(n756) );
  NANDN U873 ( .A(B[142]), .B(n760), .Z(n759) );
  NANDN U874 ( .A(A[142]), .B(n761), .Z(n760) );
  NANDN U875 ( .A(n761), .B(A[142]), .Z(n758) );
  XOR U876 ( .A(n761), .B(n762), .Z(DIFF[142]) );
  XOR U877 ( .A(B[142]), .B(A[142]), .Z(n762) );
  AND U878 ( .A(n763), .B(n764), .Z(n761) );
  NANDN U879 ( .A(B[141]), .B(n765), .Z(n764) );
  NANDN U880 ( .A(A[141]), .B(n766), .Z(n765) );
  NANDN U881 ( .A(n766), .B(A[141]), .Z(n763) );
  XOR U882 ( .A(n766), .B(n767), .Z(DIFF[141]) );
  XOR U883 ( .A(B[141]), .B(A[141]), .Z(n767) );
  AND U884 ( .A(n768), .B(n769), .Z(n766) );
  NANDN U885 ( .A(B[140]), .B(n770), .Z(n769) );
  NANDN U886 ( .A(A[140]), .B(n771), .Z(n770) );
  NANDN U887 ( .A(n771), .B(A[140]), .Z(n768) );
  XOR U888 ( .A(n771), .B(n772), .Z(DIFF[140]) );
  XOR U889 ( .A(B[140]), .B(A[140]), .Z(n772) );
  AND U890 ( .A(n773), .B(n774), .Z(n771) );
  NANDN U891 ( .A(B[139]), .B(n775), .Z(n774) );
  NANDN U892 ( .A(A[139]), .B(n776), .Z(n775) );
  NANDN U893 ( .A(n776), .B(A[139]), .Z(n773) );
  XOR U894 ( .A(n777), .B(n778), .Z(DIFF[13]) );
  XOR U895 ( .A(B[13]), .B(A[13]), .Z(n778) );
  XOR U896 ( .A(n776), .B(n779), .Z(DIFF[139]) );
  XOR U897 ( .A(B[139]), .B(A[139]), .Z(n779) );
  AND U898 ( .A(n780), .B(n781), .Z(n776) );
  NANDN U899 ( .A(B[138]), .B(n782), .Z(n781) );
  NANDN U900 ( .A(A[138]), .B(n783), .Z(n782) );
  NANDN U901 ( .A(n783), .B(A[138]), .Z(n780) );
  XOR U902 ( .A(n783), .B(n784), .Z(DIFF[138]) );
  XOR U903 ( .A(B[138]), .B(A[138]), .Z(n784) );
  AND U904 ( .A(n785), .B(n786), .Z(n783) );
  NANDN U905 ( .A(B[137]), .B(n787), .Z(n786) );
  NANDN U906 ( .A(A[137]), .B(n788), .Z(n787) );
  NANDN U907 ( .A(n788), .B(A[137]), .Z(n785) );
  XOR U908 ( .A(n788), .B(n789), .Z(DIFF[137]) );
  XOR U909 ( .A(B[137]), .B(A[137]), .Z(n789) );
  AND U910 ( .A(n790), .B(n791), .Z(n788) );
  NANDN U911 ( .A(B[136]), .B(n792), .Z(n791) );
  NANDN U912 ( .A(A[136]), .B(n793), .Z(n792) );
  NANDN U913 ( .A(n793), .B(A[136]), .Z(n790) );
  XOR U914 ( .A(n793), .B(n794), .Z(DIFF[136]) );
  XOR U915 ( .A(B[136]), .B(A[136]), .Z(n794) );
  AND U916 ( .A(n795), .B(n796), .Z(n793) );
  NANDN U917 ( .A(B[135]), .B(n797), .Z(n796) );
  NANDN U918 ( .A(A[135]), .B(n798), .Z(n797) );
  NANDN U919 ( .A(n798), .B(A[135]), .Z(n795) );
  XOR U920 ( .A(n798), .B(n799), .Z(DIFF[135]) );
  XOR U921 ( .A(B[135]), .B(A[135]), .Z(n799) );
  AND U922 ( .A(n800), .B(n801), .Z(n798) );
  NANDN U923 ( .A(B[134]), .B(n802), .Z(n801) );
  NANDN U924 ( .A(A[134]), .B(n803), .Z(n802) );
  NANDN U925 ( .A(n803), .B(A[134]), .Z(n800) );
  XOR U926 ( .A(n803), .B(n804), .Z(DIFF[134]) );
  XOR U927 ( .A(B[134]), .B(A[134]), .Z(n804) );
  AND U928 ( .A(n805), .B(n806), .Z(n803) );
  NANDN U929 ( .A(B[133]), .B(n807), .Z(n806) );
  NANDN U930 ( .A(A[133]), .B(n808), .Z(n807) );
  NANDN U931 ( .A(n808), .B(A[133]), .Z(n805) );
  XOR U932 ( .A(n808), .B(n809), .Z(DIFF[133]) );
  XOR U933 ( .A(B[133]), .B(A[133]), .Z(n809) );
  AND U934 ( .A(n810), .B(n811), .Z(n808) );
  NANDN U935 ( .A(B[132]), .B(n812), .Z(n811) );
  NANDN U936 ( .A(A[132]), .B(n813), .Z(n812) );
  NANDN U937 ( .A(n813), .B(A[132]), .Z(n810) );
  XOR U938 ( .A(n813), .B(n814), .Z(DIFF[132]) );
  XOR U939 ( .A(B[132]), .B(A[132]), .Z(n814) );
  AND U940 ( .A(n815), .B(n816), .Z(n813) );
  NANDN U941 ( .A(B[131]), .B(n817), .Z(n816) );
  NANDN U942 ( .A(A[131]), .B(n818), .Z(n817) );
  NANDN U943 ( .A(n818), .B(A[131]), .Z(n815) );
  XOR U944 ( .A(n818), .B(n819), .Z(DIFF[131]) );
  XOR U945 ( .A(B[131]), .B(A[131]), .Z(n819) );
  AND U946 ( .A(n820), .B(n821), .Z(n818) );
  NANDN U947 ( .A(B[130]), .B(n822), .Z(n821) );
  NANDN U948 ( .A(A[130]), .B(n823), .Z(n822) );
  NANDN U949 ( .A(n823), .B(A[130]), .Z(n820) );
  XOR U950 ( .A(n823), .B(n824), .Z(DIFF[130]) );
  XOR U951 ( .A(B[130]), .B(A[130]), .Z(n824) );
  AND U952 ( .A(n825), .B(n826), .Z(n823) );
  NANDN U953 ( .A(B[129]), .B(n827), .Z(n826) );
  NANDN U954 ( .A(A[129]), .B(n828), .Z(n827) );
  NANDN U955 ( .A(n828), .B(A[129]), .Z(n825) );
  XOR U956 ( .A(n829), .B(n830), .Z(DIFF[12]) );
  XOR U957 ( .A(B[12]), .B(A[12]), .Z(n830) );
  XOR U958 ( .A(n828), .B(n831), .Z(DIFF[129]) );
  XOR U959 ( .A(B[129]), .B(A[129]), .Z(n831) );
  AND U960 ( .A(n832), .B(n833), .Z(n828) );
  NANDN U961 ( .A(B[128]), .B(n834), .Z(n833) );
  NANDN U962 ( .A(A[128]), .B(n835), .Z(n834) );
  NANDN U963 ( .A(n835), .B(A[128]), .Z(n832) );
  XOR U964 ( .A(n835), .B(n836), .Z(DIFF[128]) );
  XOR U965 ( .A(B[128]), .B(A[128]), .Z(n836) );
  AND U966 ( .A(n837), .B(n838), .Z(n835) );
  NANDN U967 ( .A(B[127]), .B(n839), .Z(n838) );
  NANDN U968 ( .A(A[127]), .B(n840), .Z(n839) );
  NANDN U969 ( .A(n840), .B(A[127]), .Z(n837) );
  XOR U970 ( .A(n840), .B(n841), .Z(DIFF[127]) );
  XOR U971 ( .A(B[127]), .B(A[127]), .Z(n841) );
  AND U972 ( .A(n842), .B(n843), .Z(n840) );
  NANDN U973 ( .A(B[126]), .B(n844), .Z(n843) );
  NANDN U974 ( .A(A[126]), .B(n845), .Z(n844) );
  NANDN U975 ( .A(n845), .B(A[126]), .Z(n842) );
  XOR U976 ( .A(n845), .B(n846), .Z(DIFF[126]) );
  XOR U977 ( .A(B[126]), .B(A[126]), .Z(n846) );
  AND U978 ( .A(n847), .B(n848), .Z(n845) );
  NANDN U979 ( .A(B[125]), .B(n849), .Z(n848) );
  NANDN U980 ( .A(A[125]), .B(n850), .Z(n849) );
  NANDN U981 ( .A(n850), .B(A[125]), .Z(n847) );
  XOR U982 ( .A(n850), .B(n851), .Z(DIFF[125]) );
  XOR U983 ( .A(B[125]), .B(A[125]), .Z(n851) );
  AND U984 ( .A(n852), .B(n853), .Z(n850) );
  NANDN U985 ( .A(B[124]), .B(n854), .Z(n853) );
  NANDN U986 ( .A(A[124]), .B(n855), .Z(n854) );
  NANDN U987 ( .A(n855), .B(A[124]), .Z(n852) );
  XOR U988 ( .A(n855), .B(n856), .Z(DIFF[124]) );
  XOR U989 ( .A(B[124]), .B(A[124]), .Z(n856) );
  AND U990 ( .A(n857), .B(n858), .Z(n855) );
  NANDN U991 ( .A(B[123]), .B(n859), .Z(n858) );
  NANDN U992 ( .A(A[123]), .B(n860), .Z(n859) );
  NANDN U993 ( .A(n860), .B(A[123]), .Z(n857) );
  XOR U994 ( .A(n860), .B(n861), .Z(DIFF[123]) );
  XOR U995 ( .A(B[123]), .B(A[123]), .Z(n861) );
  AND U996 ( .A(n862), .B(n863), .Z(n860) );
  NANDN U997 ( .A(B[122]), .B(n864), .Z(n863) );
  NANDN U998 ( .A(A[122]), .B(n865), .Z(n864) );
  NANDN U999 ( .A(n865), .B(A[122]), .Z(n862) );
  XOR U1000 ( .A(n865), .B(n866), .Z(DIFF[122]) );
  XOR U1001 ( .A(B[122]), .B(A[122]), .Z(n866) );
  AND U1002 ( .A(n867), .B(n868), .Z(n865) );
  NANDN U1003 ( .A(B[121]), .B(n869), .Z(n868) );
  NANDN U1004 ( .A(A[121]), .B(n870), .Z(n869) );
  NANDN U1005 ( .A(n870), .B(A[121]), .Z(n867) );
  XOR U1006 ( .A(n870), .B(n871), .Z(DIFF[121]) );
  XOR U1007 ( .A(B[121]), .B(A[121]), .Z(n871) );
  AND U1008 ( .A(n872), .B(n873), .Z(n870) );
  NANDN U1009 ( .A(B[120]), .B(n874), .Z(n873) );
  NANDN U1010 ( .A(A[120]), .B(n875), .Z(n874) );
  NANDN U1011 ( .A(n875), .B(A[120]), .Z(n872) );
  XOR U1012 ( .A(n875), .B(n876), .Z(DIFF[120]) );
  XOR U1013 ( .A(B[120]), .B(A[120]), .Z(n876) );
  AND U1014 ( .A(n877), .B(n878), .Z(n875) );
  NANDN U1015 ( .A(B[119]), .B(n879), .Z(n878) );
  NANDN U1016 ( .A(A[119]), .B(n880), .Z(n879) );
  NANDN U1017 ( .A(n880), .B(A[119]), .Z(n877) );
  XOR U1018 ( .A(n881), .B(n882), .Z(DIFF[11]) );
  XOR U1019 ( .A(B[11]), .B(A[11]), .Z(n882) );
  XOR U1020 ( .A(n880), .B(n883), .Z(DIFF[119]) );
  XOR U1021 ( .A(B[119]), .B(A[119]), .Z(n883) );
  AND U1022 ( .A(n884), .B(n885), .Z(n880) );
  NANDN U1023 ( .A(B[118]), .B(n886), .Z(n885) );
  NANDN U1024 ( .A(A[118]), .B(n887), .Z(n886) );
  NANDN U1025 ( .A(n887), .B(A[118]), .Z(n884) );
  XOR U1026 ( .A(n887), .B(n888), .Z(DIFF[118]) );
  XOR U1027 ( .A(B[118]), .B(A[118]), .Z(n888) );
  AND U1028 ( .A(n889), .B(n890), .Z(n887) );
  NANDN U1029 ( .A(B[117]), .B(n891), .Z(n890) );
  NANDN U1030 ( .A(A[117]), .B(n892), .Z(n891) );
  NANDN U1031 ( .A(n892), .B(A[117]), .Z(n889) );
  XOR U1032 ( .A(n892), .B(n893), .Z(DIFF[117]) );
  XOR U1033 ( .A(B[117]), .B(A[117]), .Z(n893) );
  AND U1034 ( .A(n894), .B(n895), .Z(n892) );
  NANDN U1035 ( .A(B[116]), .B(n896), .Z(n895) );
  NANDN U1036 ( .A(A[116]), .B(n897), .Z(n896) );
  NANDN U1037 ( .A(n897), .B(A[116]), .Z(n894) );
  XOR U1038 ( .A(n897), .B(n898), .Z(DIFF[116]) );
  XOR U1039 ( .A(B[116]), .B(A[116]), .Z(n898) );
  AND U1040 ( .A(n899), .B(n900), .Z(n897) );
  NANDN U1041 ( .A(B[115]), .B(n901), .Z(n900) );
  NANDN U1042 ( .A(A[115]), .B(n902), .Z(n901) );
  NANDN U1043 ( .A(n902), .B(A[115]), .Z(n899) );
  XOR U1044 ( .A(n902), .B(n903), .Z(DIFF[115]) );
  XOR U1045 ( .A(B[115]), .B(A[115]), .Z(n903) );
  AND U1046 ( .A(n904), .B(n905), .Z(n902) );
  NANDN U1047 ( .A(B[114]), .B(n906), .Z(n905) );
  NANDN U1048 ( .A(A[114]), .B(n907), .Z(n906) );
  NANDN U1049 ( .A(n907), .B(A[114]), .Z(n904) );
  XOR U1050 ( .A(n907), .B(n908), .Z(DIFF[114]) );
  XOR U1051 ( .A(B[114]), .B(A[114]), .Z(n908) );
  AND U1052 ( .A(n909), .B(n910), .Z(n907) );
  NANDN U1053 ( .A(B[113]), .B(n911), .Z(n910) );
  NANDN U1054 ( .A(A[113]), .B(n912), .Z(n911) );
  NANDN U1055 ( .A(n912), .B(A[113]), .Z(n909) );
  XOR U1056 ( .A(n912), .B(n913), .Z(DIFF[113]) );
  XOR U1057 ( .A(B[113]), .B(A[113]), .Z(n913) );
  AND U1058 ( .A(n914), .B(n915), .Z(n912) );
  NANDN U1059 ( .A(B[112]), .B(n916), .Z(n915) );
  NANDN U1060 ( .A(A[112]), .B(n917), .Z(n916) );
  NANDN U1061 ( .A(n917), .B(A[112]), .Z(n914) );
  XOR U1062 ( .A(n917), .B(n918), .Z(DIFF[112]) );
  XOR U1063 ( .A(B[112]), .B(A[112]), .Z(n918) );
  AND U1064 ( .A(n919), .B(n920), .Z(n917) );
  NANDN U1065 ( .A(B[111]), .B(n921), .Z(n920) );
  NANDN U1066 ( .A(A[111]), .B(n922), .Z(n921) );
  NANDN U1067 ( .A(n922), .B(A[111]), .Z(n919) );
  XOR U1068 ( .A(n922), .B(n923), .Z(DIFF[111]) );
  XOR U1069 ( .A(B[111]), .B(A[111]), .Z(n923) );
  AND U1070 ( .A(n924), .B(n925), .Z(n922) );
  NANDN U1071 ( .A(B[110]), .B(n926), .Z(n925) );
  NANDN U1072 ( .A(A[110]), .B(n927), .Z(n926) );
  NANDN U1073 ( .A(n927), .B(A[110]), .Z(n924) );
  XOR U1074 ( .A(n927), .B(n928), .Z(DIFF[110]) );
  XOR U1075 ( .A(B[110]), .B(A[110]), .Z(n928) );
  AND U1076 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U1077 ( .A(B[109]), .B(n931), .Z(n930) );
  NANDN U1078 ( .A(A[109]), .B(n932), .Z(n931) );
  NANDN U1079 ( .A(n932), .B(A[109]), .Z(n929) );
  XOR U1080 ( .A(n933), .B(n934), .Z(DIFF[10]) );
  XOR U1081 ( .A(B[10]), .B(A[10]), .Z(n934) );
  XOR U1082 ( .A(n932), .B(n935), .Z(DIFF[109]) );
  XOR U1083 ( .A(B[109]), .B(A[109]), .Z(n935) );
  AND U1084 ( .A(n936), .B(n937), .Z(n932) );
  NANDN U1085 ( .A(B[108]), .B(n938), .Z(n937) );
  NANDN U1086 ( .A(A[108]), .B(n939), .Z(n938) );
  NANDN U1087 ( .A(n939), .B(A[108]), .Z(n936) );
  XOR U1088 ( .A(n939), .B(n940), .Z(DIFF[108]) );
  XOR U1089 ( .A(B[108]), .B(A[108]), .Z(n940) );
  AND U1090 ( .A(n941), .B(n942), .Z(n939) );
  NANDN U1091 ( .A(B[107]), .B(n943), .Z(n942) );
  NANDN U1092 ( .A(A[107]), .B(n944), .Z(n943) );
  NANDN U1093 ( .A(n944), .B(A[107]), .Z(n941) );
  XOR U1094 ( .A(n944), .B(n945), .Z(DIFF[107]) );
  XOR U1095 ( .A(B[107]), .B(A[107]), .Z(n945) );
  AND U1096 ( .A(n946), .B(n947), .Z(n944) );
  NANDN U1097 ( .A(B[106]), .B(n948), .Z(n947) );
  NANDN U1098 ( .A(A[106]), .B(n949), .Z(n948) );
  NANDN U1099 ( .A(n949), .B(A[106]), .Z(n946) );
  XOR U1100 ( .A(n949), .B(n950), .Z(DIFF[106]) );
  XOR U1101 ( .A(B[106]), .B(A[106]), .Z(n950) );
  AND U1102 ( .A(n951), .B(n952), .Z(n949) );
  NANDN U1103 ( .A(B[105]), .B(n953), .Z(n952) );
  NANDN U1104 ( .A(A[105]), .B(n954), .Z(n953) );
  NANDN U1105 ( .A(n954), .B(A[105]), .Z(n951) );
  XOR U1106 ( .A(n954), .B(n955), .Z(DIFF[105]) );
  XOR U1107 ( .A(B[105]), .B(A[105]), .Z(n955) );
  AND U1108 ( .A(n956), .B(n957), .Z(n954) );
  NANDN U1109 ( .A(B[104]), .B(n958), .Z(n957) );
  NANDN U1110 ( .A(A[104]), .B(n959), .Z(n958) );
  NANDN U1111 ( .A(n959), .B(A[104]), .Z(n956) );
  XOR U1112 ( .A(n959), .B(n960), .Z(DIFF[104]) );
  XOR U1113 ( .A(B[104]), .B(A[104]), .Z(n960) );
  AND U1114 ( .A(n961), .B(n962), .Z(n959) );
  NANDN U1115 ( .A(B[103]), .B(n963), .Z(n962) );
  NANDN U1116 ( .A(A[103]), .B(n964), .Z(n963) );
  NANDN U1117 ( .A(n964), .B(A[103]), .Z(n961) );
  XOR U1118 ( .A(n964), .B(n965), .Z(DIFF[103]) );
  XOR U1119 ( .A(B[103]), .B(A[103]), .Z(n965) );
  AND U1120 ( .A(n966), .B(n967), .Z(n964) );
  NANDN U1121 ( .A(B[102]), .B(n968), .Z(n967) );
  NANDN U1122 ( .A(A[102]), .B(n969), .Z(n968) );
  NANDN U1123 ( .A(n969), .B(A[102]), .Z(n966) );
  XOR U1124 ( .A(n969), .B(n970), .Z(DIFF[102]) );
  XOR U1125 ( .A(B[102]), .B(A[102]), .Z(n970) );
  AND U1126 ( .A(n971), .B(n972), .Z(n969) );
  NANDN U1127 ( .A(B[101]), .B(n973), .Z(n972) );
  NANDN U1128 ( .A(A[101]), .B(n974), .Z(n973) );
  NANDN U1129 ( .A(n974), .B(A[101]), .Z(n971) );
  XOR U1130 ( .A(n974), .B(n975), .Z(DIFF[101]) );
  XOR U1131 ( .A(B[101]), .B(A[101]), .Z(n975) );
  AND U1132 ( .A(n976), .B(n977), .Z(n974) );
  NANDN U1133 ( .A(B[100]), .B(n978), .Z(n977) );
  NANDN U1134 ( .A(A[100]), .B(n979), .Z(n978) );
  NANDN U1135 ( .A(n979), .B(A[100]), .Z(n976) );
  XOR U1136 ( .A(n979), .B(n980), .Z(DIFF[100]) );
  XOR U1137 ( .A(B[100]), .B(A[100]), .Z(n980) );
  AND U1138 ( .A(n981), .B(n982), .Z(n979) );
  NANDN U1139 ( .A(B[99]), .B(n983), .Z(n982) );
  OR U1140 ( .A(n5), .B(A[99]), .Z(n983) );
  NAND U1141 ( .A(A[99]), .B(n5), .Z(n981) );
  NAND U1142 ( .A(n984), .B(n985), .Z(n5) );
  NANDN U1143 ( .A(B[98]), .B(n986), .Z(n985) );
  NANDN U1144 ( .A(A[98]), .B(n7), .Z(n986) );
  NANDN U1145 ( .A(n7), .B(A[98]), .Z(n984) );
  AND U1146 ( .A(n987), .B(n988), .Z(n7) );
  NANDN U1147 ( .A(B[97]), .B(n989), .Z(n988) );
  NANDN U1148 ( .A(A[97]), .B(n9), .Z(n989) );
  NANDN U1149 ( .A(n9), .B(A[97]), .Z(n987) );
  AND U1150 ( .A(n990), .B(n991), .Z(n9) );
  NANDN U1151 ( .A(B[96]), .B(n992), .Z(n991) );
  NANDN U1152 ( .A(A[96]), .B(n11), .Z(n992) );
  NANDN U1153 ( .A(n11), .B(A[96]), .Z(n990) );
  AND U1154 ( .A(n993), .B(n994), .Z(n11) );
  NANDN U1155 ( .A(B[95]), .B(n995), .Z(n994) );
  NANDN U1156 ( .A(A[95]), .B(n13), .Z(n995) );
  NANDN U1157 ( .A(n13), .B(A[95]), .Z(n993) );
  AND U1158 ( .A(n996), .B(n997), .Z(n13) );
  NANDN U1159 ( .A(B[94]), .B(n998), .Z(n997) );
  NANDN U1160 ( .A(A[94]), .B(n15), .Z(n998) );
  NANDN U1161 ( .A(n15), .B(A[94]), .Z(n996) );
  AND U1162 ( .A(n999), .B(n1000), .Z(n15) );
  NANDN U1163 ( .A(B[93]), .B(n1001), .Z(n1000) );
  NANDN U1164 ( .A(A[93]), .B(n17), .Z(n1001) );
  NANDN U1165 ( .A(n17), .B(A[93]), .Z(n999) );
  AND U1166 ( .A(n1002), .B(n1003), .Z(n17) );
  NANDN U1167 ( .A(B[92]), .B(n1004), .Z(n1003) );
  NANDN U1168 ( .A(A[92]), .B(n19), .Z(n1004) );
  NANDN U1169 ( .A(n19), .B(A[92]), .Z(n1002) );
  AND U1170 ( .A(n1005), .B(n1006), .Z(n19) );
  NANDN U1171 ( .A(B[91]), .B(n1007), .Z(n1006) );
  NANDN U1172 ( .A(A[91]), .B(n21), .Z(n1007) );
  NANDN U1173 ( .A(n21), .B(A[91]), .Z(n1005) );
  AND U1174 ( .A(n1008), .B(n1009), .Z(n21) );
  NANDN U1175 ( .A(B[90]), .B(n1010), .Z(n1009) );
  NANDN U1176 ( .A(A[90]), .B(n23), .Z(n1010) );
  NANDN U1177 ( .A(n23), .B(A[90]), .Z(n1008) );
  AND U1178 ( .A(n1011), .B(n1012), .Z(n23) );
  NANDN U1179 ( .A(B[89]), .B(n1013), .Z(n1012) );
  NANDN U1180 ( .A(A[89]), .B(n27), .Z(n1013) );
  NANDN U1181 ( .A(n27), .B(A[89]), .Z(n1011) );
  AND U1182 ( .A(n1014), .B(n1015), .Z(n27) );
  NANDN U1183 ( .A(B[88]), .B(n1016), .Z(n1015) );
  NANDN U1184 ( .A(A[88]), .B(n29), .Z(n1016) );
  NANDN U1185 ( .A(n29), .B(A[88]), .Z(n1014) );
  AND U1186 ( .A(n1017), .B(n1018), .Z(n29) );
  NANDN U1187 ( .A(B[87]), .B(n1019), .Z(n1018) );
  NANDN U1188 ( .A(A[87]), .B(n31), .Z(n1019) );
  NANDN U1189 ( .A(n31), .B(A[87]), .Z(n1017) );
  AND U1190 ( .A(n1020), .B(n1021), .Z(n31) );
  NANDN U1191 ( .A(B[86]), .B(n1022), .Z(n1021) );
  NANDN U1192 ( .A(A[86]), .B(n33), .Z(n1022) );
  NANDN U1193 ( .A(n33), .B(A[86]), .Z(n1020) );
  AND U1194 ( .A(n1023), .B(n1024), .Z(n33) );
  NANDN U1195 ( .A(B[85]), .B(n1025), .Z(n1024) );
  NANDN U1196 ( .A(A[85]), .B(n35), .Z(n1025) );
  NANDN U1197 ( .A(n35), .B(A[85]), .Z(n1023) );
  AND U1198 ( .A(n1026), .B(n1027), .Z(n35) );
  NANDN U1199 ( .A(B[84]), .B(n1028), .Z(n1027) );
  NANDN U1200 ( .A(A[84]), .B(n37), .Z(n1028) );
  NANDN U1201 ( .A(n37), .B(A[84]), .Z(n1026) );
  AND U1202 ( .A(n1029), .B(n1030), .Z(n37) );
  NANDN U1203 ( .A(B[83]), .B(n1031), .Z(n1030) );
  NANDN U1204 ( .A(A[83]), .B(n39), .Z(n1031) );
  NANDN U1205 ( .A(n39), .B(A[83]), .Z(n1029) );
  AND U1206 ( .A(n1032), .B(n1033), .Z(n39) );
  NANDN U1207 ( .A(B[82]), .B(n1034), .Z(n1033) );
  NANDN U1208 ( .A(A[82]), .B(n41), .Z(n1034) );
  NANDN U1209 ( .A(n41), .B(A[82]), .Z(n1032) );
  AND U1210 ( .A(n1035), .B(n1036), .Z(n41) );
  NANDN U1211 ( .A(B[81]), .B(n1037), .Z(n1036) );
  NANDN U1212 ( .A(A[81]), .B(n43), .Z(n1037) );
  NANDN U1213 ( .A(n43), .B(A[81]), .Z(n1035) );
  AND U1214 ( .A(n1038), .B(n1039), .Z(n43) );
  NANDN U1215 ( .A(B[80]), .B(n1040), .Z(n1039) );
  NANDN U1216 ( .A(A[80]), .B(n45), .Z(n1040) );
  NANDN U1217 ( .A(n45), .B(A[80]), .Z(n1038) );
  AND U1218 ( .A(n1041), .B(n1042), .Z(n45) );
  NANDN U1219 ( .A(B[79]), .B(n1043), .Z(n1042) );
  NANDN U1220 ( .A(A[79]), .B(n49), .Z(n1043) );
  NANDN U1221 ( .A(n49), .B(A[79]), .Z(n1041) );
  AND U1222 ( .A(n1044), .B(n1045), .Z(n49) );
  NANDN U1223 ( .A(B[78]), .B(n1046), .Z(n1045) );
  NANDN U1224 ( .A(A[78]), .B(n51), .Z(n1046) );
  NANDN U1225 ( .A(n51), .B(A[78]), .Z(n1044) );
  AND U1226 ( .A(n1047), .B(n1048), .Z(n51) );
  NANDN U1227 ( .A(B[77]), .B(n1049), .Z(n1048) );
  NANDN U1228 ( .A(A[77]), .B(n53), .Z(n1049) );
  NANDN U1229 ( .A(n53), .B(A[77]), .Z(n1047) );
  AND U1230 ( .A(n1050), .B(n1051), .Z(n53) );
  NANDN U1231 ( .A(B[76]), .B(n1052), .Z(n1051) );
  NANDN U1232 ( .A(A[76]), .B(n55), .Z(n1052) );
  NANDN U1233 ( .A(n55), .B(A[76]), .Z(n1050) );
  AND U1234 ( .A(n1053), .B(n1054), .Z(n55) );
  NANDN U1235 ( .A(B[75]), .B(n1055), .Z(n1054) );
  NANDN U1236 ( .A(A[75]), .B(n57), .Z(n1055) );
  NANDN U1237 ( .A(n57), .B(A[75]), .Z(n1053) );
  AND U1238 ( .A(n1056), .B(n1057), .Z(n57) );
  NANDN U1239 ( .A(B[74]), .B(n1058), .Z(n1057) );
  NANDN U1240 ( .A(A[74]), .B(n59), .Z(n1058) );
  NANDN U1241 ( .A(n59), .B(A[74]), .Z(n1056) );
  AND U1242 ( .A(n1059), .B(n1060), .Z(n59) );
  NANDN U1243 ( .A(B[73]), .B(n1061), .Z(n1060) );
  NANDN U1244 ( .A(A[73]), .B(n61), .Z(n1061) );
  NANDN U1245 ( .A(n61), .B(A[73]), .Z(n1059) );
  AND U1246 ( .A(n1062), .B(n1063), .Z(n61) );
  NANDN U1247 ( .A(B[72]), .B(n1064), .Z(n1063) );
  NANDN U1248 ( .A(A[72]), .B(n63), .Z(n1064) );
  NANDN U1249 ( .A(n63), .B(A[72]), .Z(n1062) );
  AND U1250 ( .A(n1065), .B(n1066), .Z(n63) );
  NANDN U1251 ( .A(B[71]), .B(n1067), .Z(n1066) );
  NANDN U1252 ( .A(A[71]), .B(n65), .Z(n1067) );
  NANDN U1253 ( .A(n65), .B(A[71]), .Z(n1065) );
  AND U1254 ( .A(n1068), .B(n1069), .Z(n65) );
  NANDN U1255 ( .A(B[70]), .B(n1070), .Z(n1069) );
  NANDN U1256 ( .A(A[70]), .B(n67), .Z(n1070) );
  NANDN U1257 ( .A(n67), .B(A[70]), .Z(n1068) );
  AND U1258 ( .A(n1071), .B(n1072), .Z(n67) );
  NANDN U1259 ( .A(B[69]), .B(n1073), .Z(n1072) );
  NANDN U1260 ( .A(A[69]), .B(n71), .Z(n1073) );
  NANDN U1261 ( .A(n71), .B(A[69]), .Z(n1071) );
  AND U1262 ( .A(n1074), .B(n1075), .Z(n71) );
  NANDN U1263 ( .A(B[68]), .B(n1076), .Z(n1075) );
  NANDN U1264 ( .A(A[68]), .B(n73), .Z(n1076) );
  NANDN U1265 ( .A(n73), .B(A[68]), .Z(n1074) );
  AND U1266 ( .A(n1077), .B(n1078), .Z(n73) );
  NANDN U1267 ( .A(B[67]), .B(n1079), .Z(n1078) );
  NANDN U1268 ( .A(A[67]), .B(n75), .Z(n1079) );
  NANDN U1269 ( .A(n75), .B(A[67]), .Z(n1077) );
  AND U1270 ( .A(n1080), .B(n1081), .Z(n75) );
  NANDN U1271 ( .A(B[66]), .B(n1082), .Z(n1081) );
  NANDN U1272 ( .A(A[66]), .B(n77), .Z(n1082) );
  NANDN U1273 ( .A(n77), .B(A[66]), .Z(n1080) );
  AND U1274 ( .A(n1083), .B(n1084), .Z(n77) );
  NANDN U1275 ( .A(B[65]), .B(n1085), .Z(n1084) );
  NANDN U1276 ( .A(A[65]), .B(n79), .Z(n1085) );
  NANDN U1277 ( .A(n79), .B(A[65]), .Z(n1083) );
  AND U1278 ( .A(n1086), .B(n1087), .Z(n79) );
  NANDN U1279 ( .A(B[64]), .B(n1088), .Z(n1087) );
  NANDN U1280 ( .A(A[64]), .B(n81), .Z(n1088) );
  NANDN U1281 ( .A(n81), .B(A[64]), .Z(n1086) );
  AND U1282 ( .A(n1089), .B(n1090), .Z(n81) );
  NANDN U1283 ( .A(B[63]), .B(n1091), .Z(n1090) );
  NANDN U1284 ( .A(A[63]), .B(n83), .Z(n1091) );
  NANDN U1285 ( .A(n83), .B(A[63]), .Z(n1089) );
  AND U1286 ( .A(n1092), .B(n1093), .Z(n83) );
  NANDN U1287 ( .A(B[62]), .B(n1094), .Z(n1093) );
  NANDN U1288 ( .A(A[62]), .B(n85), .Z(n1094) );
  NANDN U1289 ( .A(n85), .B(A[62]), .Z(n1092) );
  AND U1290 ( .A(n1095), .B(n1096), .Z(n85) );
  NANDN U1291 ( .A(B[61]), .B(n1097), .Z(n1096) );
  NANDN U1292 ( .A(A[61]), .B(n87), .Z(n1097) );
  NANDN U1293 ( .A(n87), .B(A[61]), .Z(n1095) );
  AND U1294 ( .A(n1098), .B(n1099), .Z(n87) );
  NANDN U1295 ( .A(B[60]), .B(n1100), .Z(n1099) );
  NANDN U1296 ( .A(A[60]), .B(n89), .Z(n1100) );
  NANDN U1297 ( .A(n89), .B(A[60]), .Z(n1098) );
  AND U1298 ( .A(n1101), .B(n1102), .Z(n89) );
  NANDN U1299 ( .A(B[59]), .B(n1103), .Z(n1102) );
  NANDN U1300 ( .A(A[59]), .B(n93), .Z(n1103) );
  NANDN U1301 ( .A(n93), .B(A[59]), .Z(n1101) );
  AND U1302 ( .A(n1104), .B(n1105), .Z(n93) );
  NANDN U1303 ( .A(B[58]), .B(n1106), .Z(n1105) );
  NANDN U1304 ( .A(A[58]), .B(n95), .Z(n1106) );
  NANDN U1305 ( .A(n95), .B(A[58]), .Z(n1104) );
  AND U1306 ( .A(n1107), .B(n1108), .Z(n95) );
  NANDN U1307 ( .A(B[57]), .B(n1109), .Z(n1108) );
  NANDN U1308 ( .A(A[57]), .B(n97), .Z(n1109) );
  NANDN U1309 ( .A(n97), .B(A[57]), .Z(n1107) );
  AND U1310 ( .A(n1110), .B(n1111), .Z(n97) );
  NANDN U1311 ( .A(B[56]), .B(n1112), .Z(n1111) );
  NANDN U1312 ( .A(A[56]), .B(n99), .Z(n1112) );
  NANDN U1313 ( .A(n99), .B(A[56]), .Z(n1110) );
  AND U1314 ( .A(n1113), .B(n1114), .Z(n99) );
  NANDN U1315 ( .A(B[55]), .B(n1115), .Z(n1114) );
  NANDN U1316 ( .A(A[55]), .B(n101), .Z(n1115) );
  NANDN U1317 ( .A(n101), .B(A[55]), .Z(n1113) );
  AND U1318 ( .A(n1116), .B(n1117), .Z(n101) );
  NANDN U1319 ( .A(B[54]), .B(n1118), .Z(n1117) );
  NANDN U1320 ( .A(A[54]), .B(n103), .Z(n1118) );
  NANDN U1321 ( .A(n103), .B(A[54]), .Z(n1116) );
  AND U1322 ( .A(n1119), .B(n1120), .Z(n103) );
  NANDN U1323 ( .A(B[53]), .B(n1121), .Z(n1120) );
  NANDN U1324 ( .A(A[53]), .B(n105), .Z(n1121) );
  NANDN U1325 ( .A(n105), .B(A[53]), .Z(n1119) );
  AND U1326 ( .A(n1122), .B(n1123), .Z(n105) );
  NANDN U1327 ( .A(B[52]), .B(n1124), .Z(n1123) );
  NANDN U1328 ( .A(A[52]), .B(n107), .Z(n1124) );
  NANDN U1329 ( .A(n107), .B(A[52]), .Z(n1122) );
  AND U1330 ( .A(n1125), .B(n1126), .Z(n107) );
  NANDN U1331 ( .A(B[51]), .B(n1127), .Z(n1126) );
  NANDN U1332 ( .A(A[51]), .B(n109), .Z(n1127) );
  NANDN U1333 ( .A(n109), .B(A[51]), .Z(n1125) );
  AND U1334 ( .A(n1128), .B(n1129), .Z(n109) );
  NANDN U1335 ( .A(B[50]), .B(n1130), .Z(n1129) );
  NANDN U1336 ( .A(A[50]), .B(n111), .Z(n1130) );
  NANDN U1337 ( .A(n111), .B(A[50]), .Z(n1128) );
  AND U1338 ( .A(n1131), .B(n1132), .Z(n111) );
  NANDN U1339 ( .A(B[49]), .B(n1133), .Z(n1132) );
  NANDN U1340 ( .A(A[49]), .B(n115), .Z(n1133) );
  NANDN U1341 ( .A(n115), .B(A[49]), .Z(n1131) );
  AND U1342 ( .A(n1134), .B(n1135), .Z(n115) );
  NANDN U1343 ( .A(B[48]), .B(n1136), .Z(n1135) );
  NANDN U1344 ( .A(A[48]), .B(n117), .Z(n1136) );
  NANDN U1345 ( .A(n117), .B(A[48]), .Z(n1134) );
  AND U1346 ( .A(n1137), .B(n1138), .Z(n117) );
  NANDN U1347 ( .A(B[47]), .B(n1139), .Z(n1138) );
  NANDN U1348 ( .A(A[47]), .B(n119), .Z(n1139) );
  NANDN U1349 ( .A(n119), .B(A[47]), .Z(n1137) );
  AND U1350 ( .A(n1140), .B(n1141), .Z(n119) );
  NANDN U1351 ( .A(B[46]), .B(n1142), .Z(n1141) );
  NANDN U1352 ( .A(A[46]), .B(n121), .Z(n1142) );
  NANDN U1353 ( .A(n121), .B(A[46]), .Z(n1140) );
  AND U1354 ( .A(n1143), .B(n1144), .Z(n121) );
  NANDN U1355 ( .A(B[45]), .B(n1145), .Z(n1144) );
  NANDN U1356 ( .A(A[45]), .B(n123), .Z(n1145) );
  NANDN U1357 ( .A(n123), .B(A[45]), .Z(n1143) );
  AND U1358 ( .A(n1146), .B(n1147), .Z(n123) );
  NANDN U1359 ( .A(B[44]), .B(n1148), .Z(n1147) );
  NANDN U1360 ( .A(A[44]), .B(n125), .Z(n1148) );
  NANDN U1361 ( .A(n125), .B(A[44]), .Z(n1146) );
  AND U1362 ( .A(n1149), .B(n1150), .Z(n125) );
  NANDN U1363 ( .A(B[43]), .B(n1151), .Z(n1150) );
  NANDN U1364 ( .A(A[43]), .B(n127), .Z(n1151) );
  NANDN U1365 ( .A(n127), .B(A[43]), .Z(n1149) );
  AND U1366 ( .A(n1152), .B(n1153), .Z(n127) );
  NANDN U1367 ( .A(B[42]), .B(n1154), .Z(n1153) );
  NANDN U1368 ( .A(A[42]), .B(n129), .Z(n1154) );
  NANDN U1369 ( .A(n129), .B(A[42]), .Z(n1152) );
  AND U1370 ( .A(n1155), .B(n1156), .Z(n129) );
  NANDN U1371 ( .A(B[41]), .B(n1157), .Z(n1156) );
  NANDN U1372 ( .A(A[41]), .B(n131), .Z(n1157) );
  NANDN U1373 ( .A(n131), .B(A[41]), .Z(n1155) );
  AND U1374 ( .A(n1158), .B(n1159), .Z(n131) );
  NANDN U1375 ( .A(B[40]), .B(n1160), .Z(n1159) );
  NANDN U1376 ( .A(A[40]), .B(n133), .Z(n1160) );
  NANDN U1377 ( .A(n133), .B(A[40]), .Z(n1158) );
  AND U1378 ( .A(n1161), .B(n1162), .Z(n133) );
  NANDN U1379 ( .A(B[39]), .B(n1163), .Z(n1162) );
  NANDN U1380 ( .A(A[39]), .B(n137), .Z(n1163) );
  NANDN U1381 ( .A(n137), .B(A[39]), .Z(n1161) );
  AND U1382 ( .A(n1164), .B(n1165), .Z(n137) );
  NANDN U1383 ( .A(B[38]), .B(n1166), .Z(n1165) );
  NANDN U1384 ( .A(A[38]), .B(n139), .Z(n1166) );
  NANDN U1385 ( .A(n139), .B(A[38]), .Z(n1164) );
  AND U1386 ( .A(n1167), .B(n1168), .Z(n139) );
  NANDN U1387 ( .A(B[37]), .B(n1169), .Z(n1168) );
  NANDN U1388 ( .A(A[37]), .B(n141), .Z(n1169) );
  NANDN U1389 ( .A(n141), .B(A[37]), .Z(n1167) );
  AND U1390 ( .A(n1170), .B(n1171), .Z(n141) );
  NANDN U1391 ( .A(B[36]), .B(n1172), .Z(n1171) );
  NANDN U1392 ( .A(A[36]), .B(n143), .Z(n1172) );
  NANDN U1393 ( .A(n143), .B(A[36]), .Z(n1170) );
  AND U1394 ( .A(n1173), .B(n1174), .Z(n143) );
  NANDN U1395 ( .A(B[35]), .B(n1175), .Z(n1174) );
  NANDN U1396 ( .A(A[35]), .B(n145), .Z(n1175) );
  NANDN U1397 ( .A(n145), .B(A[35]), .Z(n1173) );
  AND U1398 ( .A(n1176), .B(n1177), .Z(n145) );
  NANDN U1399 ( .A(B[34]), .B(n1178), .Z(n1177) );
  NANDN U1400 ( .A(A[34]), .B(n147), .Z(n1178) );
  NANDN U1401 ( .A(n147), .B(A[34]), .Z(n1176) );
  AND U1402 ( .A(n1179), .B(n1180), .Z(n147) );
  NANDN U1403 ( .A(B[33]), .B(n1181), .Z(n1180) );
  NANDN U1404 ( .A(A[33]), .B(n149), .Z(n1181) );
  NANDN U1405 ( .A(n149), .B(A[33]), .Z(n1179) );
  AND U1406 ( .A(n1182), .B(n1183), .Z(n149) );
  NANDN U1407 ( .A(B[32]), .B(n1184), .Z(n1183) );
  NANDN U1408 ( .A(A[32]), .B(n151), .Z(n1184) );
  NANDN U1409 ( .A(n151), .B(A[32]), .Z(n1182) );
  AND U1410 ( .A(n1185), .B(n1186), .Z(n151) );
  NANDN U1411 ( .A(B[31]), .B(n1187), .Z(n1186) );
  NANDN U1412 ( .A(A[31]), .B(n153), .Z(n1187) );
  NANDN U1413 ( .A(n153), .B(A[31]), .Z(n1185) );
  AND U1414 ( .A(n1188), .B(n1189), .Z(n153) );
  NANDN U1415 ( .A(B[30]), .B(n1190), .Z(n1189) );
  NANDN U1416 ( .A(A[30]), .B(n155), .Z(n1190) );
  NANDN U1417 ( .A(n155), .B(A[30]), .Z(n1188) );
  AND U1418 ( .A(n1191), .B(n1192), .Z(n155) );
  NANDN U1419 ( .A(B[29]), .B(n1193), .Z(n1192) );
  NANDN U1420 ( .A(A[29]), .B(n159), .Z(n1193) );
  NANDN U1421 ( .A(n159), .B(A[29]), .Z(n1191) );
  AND U1422 ( .A(n1194), .B(n1195), .Z(n159) );
  NANDN U1423 ( .A(B[28]), .B(n1196), .Z(n1195) );
  NANDN U1424 ( .A(A[28]), .B(n161), .Z(n1196) );
  NANDN U1425 ( .A(n161), .B(A[28]), .Z(n1194) );
  AND U1426 ( .A(n1197), .B(n1198), .Z(n161) );
  NANDN U1427 ( .A(B[27]), .B(n1199), .Z(n1198) );
  NANDN U1428 ( .A(A[27]), .B(n163), .Z(n1199) );
  NANDN U1429 ( .A(n163), .B(A[27]), .Z(n1197) );
  AND U1430 ( .A(n1200), .B(n1201), .Z(n163) );
  NANDN U1431 ( .A(B[26]), .B(n1202), .Z(n1201) );
  NANDN U1432 ( .A(A[26]), .B(n165), .Z(n1202) );
  NANDN U1433 ( .A(n165), .B(A[26]), .Z(n1200) );
  AND U1434 ( .A(n1203), .B(n1204), .Z(n165) );
  NANDN U1435 ( .A(B[25]), .B(n1205), .Z(n1204) );
  NANDN U1436 ( .A(A[25]), .B(n167), .Z(n1205) );
  NANDN U1437 ( .A(n167), .B(A[25]), .Z(n1203) );
  AND U1438 ( .A(n1206), .B(n1207), .Z(n167) );
  NANDN U1439 ( .A(B[24]), .B(n1208), .Z(n1207) );
  NANDN U1440 ( .A(A[24]), .B(n204), .Z(n1208) );
  NANDN U1441 ( .A(n204), .B(A[24]), .Z(n1206) );
  AND U1442 ( .A(n1209), .B(n1210), .Z(n204) );
  NANDN U1443 ( .A(B[23]), .B(n1211), .Z(n1210) );
  NANDN U1444 ( .A(A[23]), .B(n256), .Z(n1211) );
  NANDN U1445 ( .A(n256), .B(A[23]), .Z(n1209) );
  AND U1446 ( .A(n1212), .B(n1213), .Z(n256) );
  NANDN U1447 ( .A(B[22]), .B(n1214), .Z(n1213) );
  NANDN U1448 ( .A(A[22]), .B(n308), .Z(n1214) );
  NANDN U1449 ( .A(n308), .B(A[22]), .Z(n1212) );
  AND U1450 ( .A(n1215), .B(n1216), .Z(n308) );
  NANDN U1451 ( .A(B[21]), .B(n1217), .Z(n1216) );
  NANDN U1452 ( .A(A[21]), .B(n360), .Z(n1217) );
  NANDN U1453 ( .A(n360), .B(A[21]), .Z(n1215) );
  AND U1454 ( .A(n1218), .B(n1219), .Z(n360) );
  NANDN U1455 ( .A(B[20]), .B(n1220), .Z(n1219) );
  NANDN U1456 ( .A(A[20]), .B(n412), .Z(n1220) );
  NANDN U1457 ( .A(n412), .B(A[20]), .Z(n1218) );
  AND U1458 ( .A(n1221), .B(n1222), .Z(n412) );
  NANDN U1459 ( .A(B[19]), .B(n1223), .Z(n1222) );
  NANDN U1460 ( .A(A[19]), .B(n465), .Z(n1223) );
  NANDN U1461 ( .A(n465), .B(A[19]), .Z(n1221) );
  AND U1462 ( .A(n1224), .B(n1225), .Z(n465) );
  NANDN U1463 ( .A(B[18]), .B(n1226), .Z(n1225) );
  NANDN U1464 ( .A(A[18]), .B(n517), .Z(n1226) );
  NANDN U1465 ( .A(n517), .B(A[18]), .Z(n1224) );
  AND U1466 ( .A(n1227), .B(n1228), .Z(n517) );
  NANDN U1467 ( .A(B[17]), .B(n1229), .Z(n1228) );
  NANDN U1468 ( .A(A[17]), .B(n569), .Z(n1229) );
  NANDN U1469 ( .A(n569), .B(A[17]), .Z(n1227) );
  AND U1470 ( .A(n1230), .B(n1231), .Z(n569) );
  NANDN U1471 ( .A(B[16]), .B(n1232), .Z(n1231) );
  NANDN U1472 ( .A(A[16]), .B(n621), .Z(n1232) );
  NANDN U1473 ( .A(n621), .B(A[16]), .Z(n1230) );
  AND U1474 ( .A(n1233), .B(n1234), .Z(n621) );
  NANDN U1475 ( .A(B[15]), .B(n1235), .Z(n1234) );
  NANDN U1476 ( .A(A[15]), .B(n673), .Z(n1235) );
  NANDN U1477 ( .A(n673), .B(A[15]), .Z(n1233) );
  AND U1478 ( .A(n1236), .B(n1237), .Z(n673) );
  NANDN U1479 ( .A(B[14]), .B(n1238), .Z(n1237) );
  NANDN U1480 ( .A(A[14]), .B(n725), .Z(n1238) );
  NANDN U1481 ( .A(n725), .B(A[14]), .Z(n1236) );
  AND U1482 ( .A(n1239), .B(n1240), .Z(n725) );
  NANDN U1483 ( .A(B[13]), .B(n1241), .Z(n1240) );
  NANDN U1484 ( .A(A[13]), .B(n777), .Z(n1241) );
  NANDN U1485 ( .A(n777), .B(A[13]), .Z(n1239) );
  AND U1486 ( .A(n1242), .B(n1243), .Z(n777) );
  NANDN U1487 ( .A(B[12]), .B(n1244), .Z(n1243) );
  NANDN U1488 ( .A(A[12]), .B(n829), .Z(n1244) );
  NANDN U1489 ( .A(n829), .B(A[12]), .Z(n1242) );
  AND U1490 ( .A(n1245), .B(n1246), .Z(n829) );
  NANDN U1491 ( .A(B[11]), .B(n1247), .Z(n1246) );
  NANDN U1492 ( .A(A[11]), .B(n881), .Z(n1247) );
  NANDN U1493 ( .A(n881), .B(A[11]), .Z(n1245) );
  AND U1494 ( .A(n1248), .B(n1249), .Z(n881) );
  NANDN U1495 ( .A(B[10]), .B(n1250), .Z(n1249) );
  NANDN U1496 ( .A(A[10]), .B(n933), .Z(n1250) );
  NANDN U1497 ( .A(n933), .B(A[10]), .Z(n1248) );
  AND U1498 ( .A(n1251), .B(n1252), .Z(n933) );
  NANDN U1499 ( .A(B[9]), .B(n1253), .Z(n1252) );
  OR U1500 ( .A(n3), .B(A[9]), .Z(n1253) );
  NAND U1501 ( .A(A[9]), .B(n3), .Z(n1251) );
  NAND U1502 ( .A(n1254), .B(n1255), .Z(n3) );
  NANDN U1503 ( .A(B[8]), .B(n1256), .Z(n1255) );
  NANDN U1504 ( .A(A[8]), .B(n25), .Z(n1256) );
  NANDN U1505 ( .A(n25), .B(A[8]), .Z(n1254) );
  AND U1506 ( .A(n1257), .B(n1258), .Z(n25) );
  NANDN U1507 ( .A(B[7]), .B(n1259), .Z(n1258) );
  NANDN U1508 ( .A(A[7]), .B(n47), .Z(n1259) );
  NANDN U1509 ( .A(n47), .B(A[7]), .Z(n1257) );
  AND U1510 ( .A(n1260), .B(n1261), .Z(n47) );
  NANDN U1511 ( .A(B[6]), .B(n1262), .Z(n1261) );
  NANDN U1512 ( .A(A[6]), .B(n69), .Z(n1262) );
  NANDN U1513 ( .A(n69), .B(A[6]), .Z(n1260) );
  AND U1514 ( .A(n1263), .B(n1264), .Z(n69) );
  NANDN U1515 ( .A(B[5]), .B(n1265), .Z(n1264) );
  NANDN U1516 ( .A(A[5]), .B(n91), .Z(n1265) );
  NANDN U1517 ( .A(n91), .B(A[5]), .Z(n1263) );
  AND U1518 ( .A(n1266), .B(n1267), .Z(n91) );
  NANDN U1519 ( .A(B[4]), .B(n1268), .Z(n1267) );
  NANDN U1520 ( .A(A[4]), .B(n113), .Z(n1268) );
  NANDN U1521 ( .A(n113), .B(A[4]), .Z(n1266) );
  AND U1522 ( .A(n1269), .B(n1270), .Z(n113) );
  NANDN U1523 ( .A(B[3]), .B(n1271), .Z(n1270) );
  NANDN U1524 ( .A(A[3]), .B(n135), .Z(n1271) );
  NANDN U1525 ( .A(n135), .B(A[3]), .Z(n1269) );
  AND U1526 ( .A(n1272), .B(n1273), .Z(n135) );
  NANDN U1527 ( .A(B[2]), .B(n1274), .Z(n1273) );
  NANDN U1528 ( .A(A[2]), .B(n157), .Z(n1274) );
  NANDN U1529 ( .A(n157), .B(A[2]), .Z(n1272) );
  AND U1530 ( .A(n1275), .B(n1276), .Z(n157) );
  NANDN U1531 ( .A(B[1]), .B(n1277), .Z(n1276) );
  NAND U1532 ( .A(n1), .B(n2), .Z(n1277) );
  NAND U1533 ( .A(A[1]), .B(n1278), .Z(n1275) );
  NAND U1534 ( .A(n1278), .B(n1279), .Z(DIFF[0]) );
  NANDN U1535 ( .A(B[0]), .B(A[0]), .Z(n1279) );
  NANDN U1536 ( .A(A[0]), .B(B[0]), .Z(n1278) );
endmodule


module modmult_step_N256_5_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [255:0] A;
  input [0:0] B;
  output [256:0] PRODUCT;
  input TC;


  AND U2 ( .A(A[255]), .B(B[0]), .Z(PRODUCT[255]) );
  AND U3 ( .A(A[254]), .B(B[0]), .Z(PRODUCT[254]) );
  AND U4 ( .A(A[253]), .B(B[0]), .Z(PRODUCT[253]) );
  AND U5 ( .A(A[252]), .B(B[0]), .Z(PRODUCT[252]) );
  AND U6 ( .A(A[251]), .B(B[0]), .Z(PRODUCT[251]) );
  AND U7 ( .A(A[250]), .B(B[0]), .Z(PRODUCT[250]) );
  AND U8 ( .A(A[249]), .B(B[0]), .Z(PRODUCT[249]) );
  AND U9 ( .A(A[248]), .B(B[0]), .Z(PRODUCT[248]) );
  AND U10 ( .A(A[247]), .B(B[0]), .Z(PRODUCT[247]) );
  AND U11 ( .A(A[246]), .B(B[0]), .Z(PRODUCT[246]) );
  AND U12 ( .A(A[245]), .B(B[0]), .Z(PRODUCT[245]) );
  AND U13 ( .A(A[244]), .B(B[0]), .Z(PRODUCT[244]) );
  AND U14 ( .A(A[243]), .B(B[0]), .Z(PRODUCT[243]) );
  AND U15 ( .A(A[242]), .B(B[0]), .Z(PRODUCT[242]) );
  AND U16 ( .A(A[241]), .B(B[0]), .Z(PRODUCT[241]) );
  AND U17 ( .A(A[240]), .B(B[0]), .Z(PRODUCT[240]) );
  AND U18 ( .A(A[239]), .B(B[0]), .Z(PRODUCT[239]) );
  AND U19 ( .A(A[238]), .B(B[0]), .Z(PRODUCT[238]) );
  AND U20 ( .A(A[237]), .B(B[0]), .Z(PRODUCT[237]) );
  AND U21 ( .A(A[236]), .B(B[0]), .Z(PRODUCT[236]) );
  AND U22 ( .A(A[235]), .B(B[0]), .Z(PRODUCT[235]) );
  AND U23 ( .A(A[234]), .B(B[0]), .Z(PRODUCT[234]) );
  AND U24 ( .A(A[233]), .B(B[0]), .Z(PRODUCT[233]) );
  AND U25 ( .A(A[232]), .B(B[0]), .Z(PRODUCT[232]) );
  AND U26 ( .A(A[231]), .B(B[0]), .Z(PRODUCT[231]) );
  AND U27 ( .A(A[230]), .B(B[0]), .Z(PRODUCT[230]) );
  AND U28 ( .A(A[229]), .B(B[0]), .Z(PRODUCT[229]) );
  AND U29 ( .A(A[228]), .B(B[0]), .Z(PRODUCT[228]) );
  AND U30 ( .A(A[227]), .B(B[0]), .Z(PRODUCT[227]) );
  AND U31 ( .A(A[226]), .B(B[0]), .Z(PRODUCT[226]) );
  AND U32 ( .A(A[225]), .B(B[0]), .Z(PRODUCT[225]) );
  AND U33 ( .A(A[224]), .B(B[0]), .Z(PRODUCT[224]) );
  AND U34 ( .A(A[223]), .B(B[0]), .Z(PRODUCT[223]) );
  AND U35 ( .A(A[222]), .B(B[0]), .Z(PRODUCT[222]) );
  AND U36 ( .A(A[221]), .B(B[0]), .Z(PRODUCT[221]) );
  AND U37 ( .A(A[220]), .B(B[0]), .Z(PRODUCT[220]) );
  AND U38 ( .A(A[219]), .B(B[0]), .Z(PRODUCT[219]) );
  AND U39 ( .A(A[218]), .B(B[0]), .Z(PRODUCT[218]) );
  AND U40 ( .A(A[217]), .B(B[0]), .Z(PRODUCT[217]) );
  AND U41 ( .A(A[216]), .B(B[0]), .Z(PRODUCT[216]) );
  AND U42 ( .A(A[215]), .B(B[0]), .Z(PRODUCT[215]) );
  AND U43 ( .A(A[214]), .B(B[0]), .Z(PRODUCT[214]) );
  AND U44 ( .A(A[213]), .B(B[0]), .Z(PRODUCT[213]) );
  AND U45 ( .A(A[212]), .B(B[0]), .Z(PRODUCT[212]) );
  AND U46 ( .A(A[211]), .B(B[0]), .Z(PRODUCT[211]) );
  AND U47 ( .A(A[210]), .B(B[0]), .Z(PRODUCT[210]) );
  AND U48 ( .A(A[209]), .B(B[0]), .Z(PRODUCT[209]) );
  AND U49 ( .A(A[208]), .B(B[0]), .Z(PRODUCT[208]) );
  AND U50 ( .A(A[207]), .B(B[0]), .Z(PRODUCT[207]) );
  AND U51 ( .A(A[206]), .B(B[0]), .Z(PRODUCT[206]) );
  AND U52 ( .A(A[205]), .B(B[0]), .Z(PRODUCT[205]) );
  AND U53 ( .A(A[204]), .B(B[0]), .Z(PRODUCT[204]) );
  AND U54 ( .A(A[203]), .B(B[0]), .Z(PRODUCT[203]) );
  AND U55 ( .A(A[202]), .B(B[0]), .Z(PRODUCT[202]) );
  AND U56 ( .A(A[201]), .B(B[0]), .Z(PRODUCT[201]) );
  AND U57 ( .A(A[200]), .B(B[0]), .Z(PRODUCT[200]) );
  AND U58 ( .A(A[199]), .B(B[0]), .Z(PRODUCT[199]) );
  AND U59 ( .A(A[198]), .B(B[0]), .Z(PRODUCT[198]) );
  AND U60 ( .A(A[197]), .B(B[0]), .Z(PRODUCT[197]) );
  AND U61 ( .A(A[196]), .B(B[0]), .Z(PRODUCT[196]) );
  AND U62 ( .A(A[195]), .B(B[0]), .Z(PRODUCT[195]) );
  AND U63 ( .A(A[194]), .B(B[0]), .Z(PRODUCT[194]) );
  AND U64 ( .A(A[193]), .B(B[0]), .Z(PRODUCT[193]) );
  AND U65 ( .A(A[192]), .B(B[0]), .Z(PRODUCT[192]) );
  AND U66 ( .A(A[191]), .B(B[0]), .Z(PRODUCT[191]) );
  AND U67 ( .A(A[190]), .B(B[0]), .Z(PRODUCT[190]) );
  AND U68 ( .A(A[189]), .B(B[0]), .Z(PRODUCT[189]) );
  AND U69 ( .A(A[188]), .B(B[0]), .Z(PRODUCT[188]) );
  AND U70 ( .A(A[187]), .B(B[0]), .Z(PRODUCT[187]) );
  AND U71 ( .A(A[186]), .B(B[0]), .Z(PRODUCT[186]) );
  AND U72 ( .A(A[185]), .B(B[0]), .Z(PRODUCT[185]) );
  AND U73 ( .A(A[184]), .B(B[0]), .Z(PRODUCT[184]) );
  AND U74 ( .A(A[183]), .B(B[0]), .Z(PRODUCT[183]) );
  AND U75 ( .A(A[182]), .B(B[0]), .Z(PRODUCT[182]) );
  AND U76 ( .A(A[181]), .B(B[0]), .Z(PRODUCT[181]) );
  AND U77 ( .A(A[180]), .B(B[0]), .Z(PRODUCT[180]) );
  AND U78 ( .A(A[179]), .B(B[0]), .Z(PRODUCT[179]) );
  AND U79 ( .A(A[178]), .B(B[0]), .Z(PRODUCT[178]) );
  AND U80 ( .A(A[177]), .B(B[0]), .Z(PRODUCT[177]) );
  AND U81 ( .A(A[176]), .B(B[0]), .Z(PRODUCT[176]) );
  AND U82 ( .A(A[175]), .B(B[0]), .Z(PRODUCT[175]) );
  AND U83 ( .A(A[174]), .B(B[0]), .Z(PRODUCT[174]) );
  AND U84 ( .A(A[173]), .B(B[0]), .Z(PRODUCT[173]) );
  AND U85 ( .A(A[172]), .B(B[0]), .Z(PRODUCT[172]) );
  AND U86 ( .A(A[171]), .B(B[0]), .Z(PRODUCT[171]) );
  AND U87 ( .A(A[170]), .B(B[0]), .Z(PRODUCT[170]) );
  AND U88 ( .A(A[169]), .B(B[0]), .Z(PRODUCT[169]) );
  AND U89 ( .A(A[168]), .B(B[0]), .Z(PRODUCT[168]) );
  AND U90 ( .A(A[167]), .B(B[0]), .Z(PRODUCT[167]) );
  AND U91 ( .A(A[166]), .B(B[0]), .Z(PRODUCT[166]) );
  AND U92 ( .A(A[165]), .B(B[0]), .Z(PRODUCT[165]) );
  AND U93 ( .A(A[164]), .B(B[0]), .Z(PRODUCT[164]) );
  AND U94 ( .A(A[163]), .B(B[0]), .Z(PRODUCT[163]) );
  AND U95 ( .A(A[162]), .B(B[0]), .Z(PRODUCT[162]) );
  AND U96 ( .A(A[161]), .B(B[0]), .Z(PRODUCT[161]) );
  AND U97 ( .A(A[160]), .B(B[0]), .Z(PRODUCT[160]) );
  AND U98 ( .A(A[159]), .B(B[0]), .Z(PRODUCT[159]) );
  AND U99 ( .A(A[158]), .B(B[0]), .Z(PRODUCT[158]) );
  AND U100 ( .A(A[157]), .B(B[0]), .Z(PRODUCT[157]) );
  AND U101 ( .A(A[156]), .B(B[0]), .Z(PRODUCT[156]) );
  AND U102 ( .A(A[155]), .B(B[0]), .Z(PRODUCT[155]) );
  AND U103 ( .A(A[154]), .B(B[0]), .Z(PRODUCT[154]) );
  AND U104 ( .A(A[153]), .B(B[0]), .Z(PRODUCT[153]) );
  AND U105 ( .A(A[152]), .B(B[0]), .Z(PRODUCT[152]) );
  AND U106 ( .A(A[151]), .B(B[0]), .Z(PRODUCT[151]) );
  AND U107 ( .A(A[150]), .B(B[0]), .Z(PRODUCT[150]) );
  AND U108 ( .A(A[149]), .B(B[0]), .Z(PRODUCT[149]) );
  AND U109 ( .A(A[148]), .B(B[0]), .Z(PRODUCT[148]) );
  AND U110 ( .A(A[147]), .B(B[0]), .Z(PRODUCT[147]) );
  AND U111 ( .A(A[146]), .B(B[0]), .Z(PRODUCT[146]) );
  AND U112 ( .A(A[145]), .B(B[0]), .Z(PRODUCT[145]) );
  AND U113 ( .A(A[144]), .B(B[0]), .Z(PRODUCT[144]) );
  AND U114 ( .A(A[143]), .B(B[0]), .Z(PRODUCT[143]) );
  AND U115 ( .A(A[142]), .B(B[0]), .Z(PRODUCT[142]) );
  AND U116 ( .A(A[141]), .B(B[0]), .Z(PRODUCT[141]) );
  AND U117 ( .A(A[140]), .B(B[0]), .Z(PRODUCT[140]) );
  AND U118 ( .A(A[139]), .B(B[0]), .Z(PRODUCT[139]) );
  AND U119 ( .A(A[138]), .B(B[0]), .Z(PRODUCT[138]) );
  AND U120 ( .A(A[137]), .B(B[0]), .Z(PRODUCT[137]) );
  AND U121 ( .A(A[136]), .B(B[0]), .Z(PRODUCT[136]) );
  AND U122 ( .A(A[135]), .B(B[0]), .Z(PRODUCT[135]) );
  AND U123 ( .A(A[134]), .B(B[0]), .Z(PRODUCT[134]) );
  AND U124 ( .A(A[133]), .B(B[0]), .Z(PRODUCT[133]) );
  AND U125 ( .A(A[132]), .B(B[0]), .Z(PRODUCT[132]) );
  AND U126 ( .A(A[131]), .B(B[0]), .Z(PRODUCT[131]) );
  AND U127 ( .A(A[130]), .B(B[0]), .Z(PRODUCT[130]) );
  AND U128 ( .A(A[129]), .B(B[0]), .Z(PRODUCT[129]) );
  AND U129 ( .A(A[128]), .B(B[0]), .Z(PRODUCT[128]) );
  AND U130 ( .A(A[127]), .B(B[0]), .Z(PRODUCT[127]) );
  AND U131 ( .A(A[126]), .B(B[0]), .Z(PRODUCT[126]) );
  AND U132 ( .A(A[125]), .B(B[0]), .Z(PRODUCT[125]) );
  AND U133 ( .A(A[124]), .B(B[0]), .Z(PRODUCT[124]) );
  AND U134 ( .A(A[123]), .B(B[0]), .Z(PRODUCT[123]) );
  AND U135 ( .A(A[122]), .B(B[0]), .Z(PRODUCT[122]) );
  AND U136 ( .A(A[121]), .B(B[0]), .Z(PRODUCT[121]) );
  AND U137 ( .A(A[120]), .B(B[0]), .Z(PRODUCT[120]) );
  AND U138 ( .A(A[119]), .B(B[0]), .Z(PRODUCT[119]) );
  AND U139 ( .A(A[118]), .B(B[0]), .Z(PRODUCT[118]) );
  AND U140 ( .A(A[117]), .B(B[0]), .Z(PRODUCT[117]) );
  AND U141 ( .A(A[116]), .B(B[0]), .Z(PRODUCT[116]) );
  AND U142 ( .A(A[115]), .B(B[0]), .Z(PRODUCT[115]) );
  AND U143 ( .A(A[114]), .B(B[0]), .Z(PRODUCT[114]) );
  AND U144 ( .A(A[113]), .B(B[0]), .Z(PRODUCT[113]) );
  AND U145 ( .A(A[112]), .B(B[0]), .Z(PRODUCT[112]) );
  AND U146 ( .A(A[111]), .B(B[0]), .Z(PRODUCT[111]) );
  AND U147 ( .A(A[110]), .B(B[0]), .Z(PRODUCT[110]) );
  AND U148 ( .A(A[109]), .B(B[0]), .Z(PRODUCT[109]) );
  AND U149 ( .A(A[108]), .B(B[0]), .Z(PRODUCT[108]) );
  AND U150 ( .A(A[107]), .B(B[0]), .Z(PRODUCT[107]) );
  AND U151 ( .A(A[106]), .B(B[0]), .Z(PRODUCT[106]) );
  AND U152 ( .A(A[105]), .B(B[0]), .Z(PRODUCT[105]) );
  AND U153 ( .A(A[104]), .B(B[0]), .Z(PRODUCT[104]) );
  AND U154 ( .A(A[103]), .B(B[0]), .Z(PRODUCT[103]) );
  AND U155 ( .A(A[102]), .B(B[0]), .Z(PRODUCT[102]) );
  AND U156 ( .A(A[101]), .B(B[0]), .Z(PRODUCT[101]) );
  AND U157 ( .A(A[100]), .B(B[0]), .Z(PRODUCT[100]) );
  AND U158 ( .A(A[99]), .B(B[0]), .Z(PRODUCT[99]) );
  AND U159 ( .A(A[98]), .B(B[0]), .Z(PRODUCT[98]) );
  AND U160 ( .A(A[97]), .B(B[0]), .Z(PRODUCT[97]) );
  AND U161 ( .A(A[96]), .B(B[0]), .Z(PRODUCT[96]) );
  AND U162 ( .A(A[95]), .B(B[0]), .Z(PRODUCT[95]) );
  AND U163 ( .A(A[94]), .B(B[0]), .Z(PRODUCT[94]) );
  AND U164 ( .A(A[93]), .B(B[0]), .Z(PRODUCT[93]) );
  AND U165 ( .A(A[92]), .B(B[0]), .Z(PRODUCT[92]) );
  AND U166 ( .A(A[91]), .B(B[0]), .Z(PRODUCT[91]) );
  AND U167 ( .A(A[90]), .B(B[0]), .Z(PRODUCT[90]) );
  AND U168 ( .A(A[89]), .B(B[0]), .Z(PRODUCT[89]) );
  AND U169 ( .A(A[88]), .B(B[0]), .Z(PRODUCT[88]) );
  AND U170 ( .A(A[87]), .B(B[0]), .Z(PRODUCT[87]) );
  AND U171 ( .A(A[86]), .B(B[0]), .Z(PRODUCT[86]) );
  AND U172 ( .A(A[85]), .B(B[0]), .Z(PRODUCT[85]) );
  AND U173 ( .A(A[84]), .B(B[0]), .Z(PRODUCT[84]) );
  AND U174 ( .A(A[83]), .B(B[0]), .Z(PRODUCT[83]) );
  AND U175 ( .A(A[82]), .B(B[0]), .Z(PRODUCT[82]) );
  AND U176 ( .A(A[81]), .B(B[0]), .Z(PRODUCT[81]) );
  AND U177 ( .A(A[80]), .B(B[0]), .Z(PRODUCT[80]) );
  AND U178 ( .A(A[79]), .B(B[0]), .Z(PRODUCT[79]) );
  AND U179 ( .A(A[78]), .B(B[0]), .Z(PRODUCT[78]) );
  AND U180 ( .A(A[77]), .B(B[0]), .Z(PRODUCT[77]) );
  AND U181 ( .A(A[76]), .B(B[0]), .Z(PRODUCT[76]) );
  AND U182 ( .A(A[75]), .B(B[0]), .Z(PRODUCT[75]) );
  AND U183 ( .A(A[74]), .B(B[0]), .Z(PRODUCT[74]) );
  AND U184 ( .A(A[73]), .B(B[0]), .Z(PRODUCT[73]) );
  AND U185 ( .A(A[72]), .B(B[0]), .Z(PRODUCT[72]) );
  AND U186 ( .A(A[71]), .B(B[0]), .Z(PRODUCT[71]) );
  AND U187 ( .A(A[70]), .B(B[0]), .Z(PRODUCT[70]) );
  AND U188 ( .A(A[69]), .B(B[0]), .Z(PRODUCT[69]) );
  AND U189 ( .A(A[68]), .B(B[0]), .Z(PRODUCT[68]) );
  AND U190 ( .A(A[67]), .B(B[0]), .Z(PRODUCT[67]) );
  AND U191 ( .A(A[66]), .B(B[0]), .Z(PRODUCT[66]) );
  AND U192 ( .A(A[65]), .B(B[0]), .Z(PRODUCT[65]) );
  AND U193 ( .A(A[64]), .B(B[0]), .Z(PRODUCT[64]) );
  AND U194 ( .A(A[63]), .B(B[0]), .Z(PRODUCT[63]) );
  AND U195 ( .A(A[62]), .B(B[0]), .Z(PRODUCT[62]) );
  AND U196 ( .A(A[61]), .B(B[0]), .Z(PRODUCT[61]) );
  AND U197 ( .A(A[60]), .B(B[0]), .Z(PRODUCT[60]) );
  AND U198 ( .A(A[59]), .B(B[0]), .Z(PRODUCT[59]) );
  AND U199 ( .A(A[58]), .B(B[0]), .Z(PRODUCT[58]) );
  AND U200 ( .A(A[57]), .B(B[0]), .Z(PRODUCT[57]) );
  AND U201 ( .A(A[56]), .B(B[0]), .Z(PRODUCT[56]) );
  AND U202 ( .A(A[55]), .B(B[0]), .Z(PRODUCT[55]) );
  AND U203 ( .A(A[54]), .B(B[0]), .Z(PRODUCT[54]) );
  AND U204 ( .A(A[53]), .B(B[0]), .Z(PRODUCT[53]) );
  AND U205 ( .A(A[52]), .B(B[0]), .Z(PRODUCT[52]) );
  AND U206 ( .A(A[51]), .B(B[0]), .Z(PRODUCT[51]) );
  AND U207 ( .A(A[50]), .B(B[0]), .Z(PRODUCT[50]) );
  AND U208 ( .A(A[49]), .B(B[0]), .Z(PRODUCT[49]) );
  AND U209 ( .A(A[48]), .B(B[0]), .Z(PRODUCT[48]) );
  AND U210 ( .A(A[47]), .B(B[0]), .Z(PRODUCT[47]) );
  AND U211 ( .A(A[46]), .B(B[0]), .Z(PRODUCT[46]) );
  AND U212 ( .A(A[45]), .B(B[0]), .Z(PRODUCT[45]) );
  AND U213 ( .A(A[44]), .B(B[0]), .Z(PRODUCT[44]) );
  AND U214 ( .A(A[43]), .B(B[0]), .Z(PRODUCT[43]) );
  AND U215 ( .A(A[42]), .B(B[0]), .Z(PRODUCT[42]) );
  AND U216 ( .A(A[41]), .B(B[0]), .Z(PRODUCT[41]) );
  AND U217 ( .A(A[40]), .B(B[0]), .Z(PRODUCT[40]) );
  AND U218 ( .A(A[39]), .B(B[0]), .Z(PRODUCT[39]) );
  AND U219 ( .A(A[38]), .B(B[0]), .Z(PRODUCT[38]) );
  AND U220 ( .A(A[37]), .B(B[0]), .Z(PRODUCT[37]) );
  AND U221 ( .A(A[36]), .B(B[0]), .Z(PRODUCT[36]) );
  AND U222 ( .A(A[35]), .B(B[0]), .Z(PRODUCT[35]) );
  AND U223 ( .A(A[34]), .B(B[0]), .Z(PRODUCT[34]) );
  AND U224 ( .A(A[33]), .B(B[0]), .Z(PRODUCT[33]) );
  AND U225 ( .A(A[32]), .B(B[0]), .Z(PRODUCT[32]) );
  AND U226 ( .A(A[31]), .B(B[0]), .Z(PRODUCT[31]) );
  AND U227 ( .A(A[30]), .B(B[0]), .Z(PRODUCT[30]) );
  AND U228 ( .A(A[29]), .B(B[0]), .Z(PRODUCT[29]) );
  AND U229 ( .A(A[28]), .B(B[0]), .Z(PRODUCT[28]) );
  AND U230 ( .A(A[27]), .B(B[0]), .Z(PRODUCT[27]) );
  AND U231 ( .A(A[26]), .B(B[0]), .Z(PRODUCT[26]) );
  AND U232 ( .A(A[25]), .B(B[0]), .Z(PRODUCT[25]) );
  AND U233 ( .A(A[24]), .B(B[0]), .Z(PRODUCT[24]) );
  AND U234 ( .A(A[23]), .B(B[0]), .Z(PRODUCT[23]) );
  AND U235 ( .A(A[22]), .B(B[0]), .Z(PRODUCT[22]) );
  AND U236 ( .A(A[21]), .B(B[0]), .Z(PRODUCT[21]) );
  AND U237 ( .A(A[20]), .B(B[0]), .Z(PRODUCT[20]) );
  AND U238 ( .A(A[19]), .B(B[0]), .Z(PRODUCT[19]) );
  AND U239 ( .A(A[18]), .B(B[0]), .Z(PRODUCT[18]) );
  AND U240 ( .A(A[17]), .B(B[0]), .Z(PRODUCT[17]) );
  AND U241 ( .A(A[16]), .B(B[0]), .Z(PRODUCT[16]) );
  AND U242 ( .A(A[15]), .B(B[0]), .Z(PRODUCT[15]) );
  AND U243 ( .A(A[14]), .B(B[0]), .Z(PRODUCT[14]) );
  AND U244 ( .A(A[13]), .B(B[0]), .Z(PRODUCT[13]) );
  AND U245 ( .A(A[12]), .B(B[0]), .Z(PRODUCT[12]) );
  AND U246 ( .A(A[11]), .B(B[0]), .Z(PRODUCT[11]) );
  AND U247 ( .A(A[10]), .B(B[0]), .Z(PRODUCT[10]) );
  AND U248 ( .A(B[0]), .B(A[9]), .Z(PRODUCT[9]) );
  AND U249 ( .A(A[8]), .B(B[0]), .Z(PRODUCT[8]) );
  AND U250 ( .A(A[7]), .B(B[0]), .Z(PRODUCT[7]) );
  AND U251 ( .A(A[6]), .B(B[0]), .Z(PRODUCT[6]) );
  AND U252 ( .A(A[5]), .B(B[0]), .Z(PRODUCT[5]) );
  AND U253 ( .A(A[4]), .B(B[0]), .Z(PRODUCT[4]) );
  AND U254 ( .A(A[3]), .B(B[0]), .Z(PRODUCT[3]) );
  AND U255 ( .A(A[2]), .B(B[0]), .Z(PRODUCT[2]) );
  AND U256 ( .A(A[1]), .B(B[0]), .Z(PRODUCT[1]) );
  AND U257 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
endmodule


module modmult_step_N256_5_DW01_cmp2_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [257:0] A;
  input [257:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;

  NAND U1 ( .A(n1), .B(n2), .Z(LT_LE) );
  NOR U2 ( .A(B[257]), .B(B[256]), .Z(n2) );
  AND U3 ( .A(n3), .B(n4), .Z(n1) );
  NAND U4 ( .A(n5), .B(n6), .Z(n4) );
  NANDN U5 ( .A(B[255]), .B(A[255]), .Z(n6) );
  NAND U6 ( .A(n7), .B(n8), .Z(n5) );
  NANDN U7 ( .A(A[254]), .B(B[254]), .Z(n8) );
  NAND U8 ( .A(n9), .B(n10), .Z(n7) );
  NANDN U9 ( .A(B[254]), .B(A[254]), .Z(n10) );
  AND U10 ( .A(n11), .B(n12), .Z(n9) );
  NAND U11 ( .A(n13), .B(n14), .Z(n12) );
  NANDN U12 ( .A(A[253]), .B(B[253]), .Z(n14) );
  AND U13 ( .A(n15), .B(n16), .Z(n13) );
  NANDN U14 ( .A(A[252]), .B(B[252]), .Z(n16) );
  NAND U15 ( .A(n17), .B(n18), .Z(n15) );
  NANDN U16 ( .A(B[252]), .B(A[252]), .Z(n18) );
  AND U17 ( .A(n19), .B(n20), .Z(n17) );
  NAND U18 ( .A(n21), .B(n22), .Z(n20) );
  NANDN U19 ( .A(A[251]), .B(B[251]), .Z(n22) );
  AND U20 ( .A(n23), .B(n24), .Z(n21) );
  NANDN U21 ( .A(A[250]), .B(B[250]), .Z(n24) );
  NAND U22 ( .A(n25), .B(n26), .Z(n23) );
  NANDN U23 ( .A(B[250]), .B(A[250]), .Z(n26) );
  AND U24 ( .A(n27), .B(n28), .Z(n25) );
  NAND U25 ( .A(n29), .B(n30), .Z(n28) );
  NANDN U26 ( .A(A[249]), .B(B[249]), .Z(n30) );
  AND U27 ( .A(n31), .B(n32), .Z(n29) );
  NANDN U28 ( .A(A[248]), .B(B[248]), .Z(n32) );
  NAND U29 ( .A(n33), .B(n34), .Z(n31) );
  NANDN U30 ( .A(B[248]), .B(A[248]), .Z(n34) );
  AND U31 ( .A(n35), .B(n36), .Z(n33) );
  NAND U32 ( .A(n37), .B(n38), .Z(n36) );
  NANDN U33 ( .A(A[247]), .B(B[247]), .Z(n38) );
  AND U34 ( .A(n39), .B(n40), .Z(n37) );
  NANDN U35 ( .A(A[246]), .B(B[246]), .Z(n40) );
  NAND U36 ( .A(n41), .B(n42), .Z(n39) );
  NANDN U37 ( .A(B[246]), .B(A[246]), .Z(n42) );
  AND U38 ( .A(n43), .B(n44), .Z(n41) );
  NAND U39 ( .A(n45), .B(n46), .Z(n44) );
  NANDN U40 ( .A(A[245]), .B(B[245]), .Z(n46) );
  AND U41 ( .A(n47), .B(n48), .Z(n45) );
  NANDN U42 ( .A(A[244]), .B(B[244]), .Z(n48) );
  NAND U43 ( .A(n49), .B(n50), .Z(n47) );
  NANDN U44 ( .A(B[244]), .B(A[244]), .Z(n50) );
  AND U45 ( .A(n51), .B(n52), .Z(n49) );
  NAND U46 ( .A(n53), .B(n54), .Z(n52) );
  NANDN U47 ( .A(A[243]), .B(B[243]), .Z(n54) );
  AND U48 ( .A(n55), .B(n56), .Z(n53) );
  NANDN U49 ( .A(A[242]), .B(B[242]), .Z(n56) );
  NAND U50 ( .A(n57), .B(n58), .Z(n55) );
  NANDN U51 ( .A(B[242]), .B(A[242]), .Z(n58) );
  AND U52 ( .A(n59), .B(n60), .Z(n57) );
  NAND U53 ( .A(n61), .B(n62), .Z(n60) );
  NANDN U54 ( .A(A[241]), .B(B[241]), .Z(n62) );
  AND U55 ( .A(n63), .B(n64), .Z(n61) );
  NANDN U56 ( .A(A[240]), .B(B[240]), .Z(n64) );
  NAND U57 ( .A(n65), .B(n66), .Z(n63) );
  NANDN U58 ( .A(B[240]), .B(A[240]), .Z(n66) );
  AND U59 ( .A(n67), .B(n68), .Z(n65) );
  NAND U60 ( .A(n69), .B(n70), .Z(n68) );
  NANDN U61 ( .A(A[239]), .B(B[239]), .Z(n70) );
  AND U62 ( .A(n71), .B(n72), .Z(n69) );
  NANDN U63 ( .A(A[238]), .B(B[238]), .Z(n72) );
  NAND U64 ( .A(n73), .B(n74), .Z(n71) );
  NANDN U65 ( .A(B[238]), .B(A[238]), .Z(n74) );
  AND U66 ( .A(n75), .B(n76), .Z(n73) );
  NAND U67 ( .A(n77), .B(n78), .Z(n76) );
  NANDN U68 ( .A(A[237]), .B(B[237]), .Z(n78) );
  AND U69 ( .A(n79), .B(n80), .Z(n77) );
  NANDN U70 ( .A(A[236]), .B(B[236]), .Z(n80) );
  NAND U71 ( .A(n81), .B(n82), .Z(n79) );
  NANDN U72 ( .A(B[236]), .B(A[236]), .Z(n82) );
  AND U73 ( .A(n83), .B(n84), .Z(n81) );
  NAND U74 ( .A(n85), .B(n86), .Z(n84) );
  NANDN U75 ( .A(A[235]), .B(B[235]), .Z(n86) );
  AND U76 ( .A(n87), .B(n88), .Z(n85) );
  NANDN U77 ( .A(A[234]), .B(B[234]), .Z(n88) );
  NAND U78 ( .A(n89), .B(n90), .Z(n87) );
  NANDN U79 ( .A(B[234]), .B(A[234]), .Z(n90) );
  AND U80 ( .A(n91), .B(n92), .Z(n89) );
  NAND U81 ( .A(n93), .B(n94), .Z(n92) );
  NANDN U82 ( .A(A[233]), .B(B[233]), .Z(n94) );
  AND U83 ( .A(n95), .B(n96), .Z(n93) );
  NANDN U84 ( .A(A[232]), .B(B[232]), .Z(n96) );
  NAND U85 ( .A(n97), .B(n98), .Z(n95) );
  NANDN U86 ( .A(B[232]), .B(A[232]), .Z(n98) );
  AND U87 ( .A(n99), .B(n100), .Z(n97) );
  NAND U88 ( .A(n101), .B(n102), .Z(n100) );
  NANDN U89 ( .A(A[231]), .B(B[231]), .Z(n102) );
  AND U90 ( .A(n103), .B(n104), .Z(n101) );
  NANDN U91 ( .A(A[230]), .B(B[230]), .Z(n104) );
  NAND U92 ( .A(n105), .B(n106), .Z(n103) );
  NANDN U93 ( .A(B[230]), .B(A[230]), .Z(n106) );
  AND U94 ( .A(n107), .B(n108), .Z(n105) );
  NAND U95 ( .A(n109), .B(n110), .Z(n108) );
  NANDN U96 ( .A(A[229]), .B(B[229]), .Z(n110) );
  AND U97 ( .A(n111), .B(n112), .Z(n109) );
  NANDN U98 ( .A(A[228]), .B(B[228]), .Z(n112) );
  NAND U99 ( .A(n113), .B(n114), .Z(n111) );
  NANDN U100 ( .A(B[228]), .B(A[228]), .Z(n114) );
  AND U101 ( .A(n115), .B(n116), .Z(n113) );
  NAND U102 ( .A(n117), .B(n118), .Z(n116) );
  NANDN U103 ( .A(A[227]), .B(B[227]), .Z(n118) );
  AND U104 ( .A(n119), .B(n120), .Z(n117) );
  NANDN U105 ( .A(A[226]), .B(B[226]), .Z(n120) );
  NAND U106 ( .A(n121), .B(n122), .Z(n119) );
  NANDN U107 ( .A(B[226]), .B(A[226]), .Z(n122) );
  AND U108 ( .A(n123), .B(n124), .Z(n121) );
  NAND U109 ( .A(n125), .B(n126), .Z(n124) );
  NANDN U110 ( .A(A[225]), .B(B[225]), .Z(n126) );
  AND U111 ( .A(n127), .B(n128), .Z(n125) );
  NANDN U112 ( .A(A[224]), .B(B[224]), .Z(n128) );
  NAND U113 ( .A(n129), .B(n130), .Z(n127) );
  NANDN U114 ( .A(B[224]), .B(A[224]), .Z(n130) );
  AND U115 ( .A(n131), .B(n132), .Z(n129) );
  NAND U116 ( .A(n133), .B(n134), .Z(n132) );
  NANDN U117 ( .A(A[223]), .B(B[223]), .Z(n134) );
  AND U118 ( .A(n135), .B(n136), .Z(n133) );
  NANDN U119 ( .A(A[222]), .B(B[222]), .Z(n136) );
  NAND U120 ( .A(n137), .B(n138), .Z(n135) );
  NANDN U121 ( .A(B[222]), .B(A[222]), .Z(n138) );
  AND U122 ( .A(n139), .B(n140), .Z(n137) );
  NAND U123 ( .A(n141), .B(n142), .Z(n140) );
  NANDN U124 ( .A(A[221]), .B(B[221]), .Z(n142) );
  AND U125 ( .A(n143), .B(n144), .Z(n141) );
  NANDN U126 ( .A(A[220]), .B(B[220]), .Z(n144) );
  NAND U127 ( .A(n145), .B(n146), .Z(n143) );
  NANDN U128 ( .A(B[220]), .B(A[220]), .Z(n146) );
  AND U129 ( .A(n147), .B(n148), .Z(n145) );
  NAND U130 ( .A(n149), .B(n150), .Z(n148) );
  NANDN U131 ( .A(A[219]), .B(B[219]), .Z(n150) );
  AND U132 ( .A(n151), .B(n152), .Z(n149) );
  NANDN U133 ( .A(A[218]), .B(B[218]), .Z(n152) );
  NAND U134 ( .A(n153), .B(n154), .Z(n151) );
  NANDN U135 ( .A(B[218]), .B(A[218]), .Z(n154) );
  AND U136 ( .A(n155), .B(n156), .Z(n153) );
  NAND U137 ( .A(n157), .B(n158), .Z(n156) );
  NANDN U138 ( .A(A[217]), .B(B[217]), .Z(n158) );
  AND U139 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U140 ( .A(A[216]), .B(B[216]), .Z(n160) );
  NAND U141 ( .A(n161), .B(n162), .Z(n159) );
  NANDN U142 ( .A(B[216]), .B(A[216]), .Z(n162) );
  AND U143 ( .A(n163), .B(n164), .Z(n161) );
  NAND U144 ( .A(n165), .B(n166), .Z(n164) );
  NANDN U145 ( .A(A[215]), .B(B[215]), .Z(n166) );
  AND U146 ( .A(n167), .B(n168), .Z(n165) );
  NANDN U147 ( .A(A[214]), .B(B[214]), .Z(n168) );
  NAND U148 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U149 ( .A(B[214]), .B(A[214]), .Z(n170) );
  AND U150 ( .A(n171), .B(n172), .Z(n169) );
  NAND U151 ( .A(n173), .B(n174), .Z(n172) );
  NANDN U152 ( .A(A[213]), .B(B[213]), .Z(n174) );
  AND U153 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U154 ( .A(A[212]), .B(B[212]), .Z(n176) );
  NAND U155 ( .A(n177), .B(n178), .Z(n175) );
  NANDN U156 ( .A(B[212]), .B(A[212]), .Z(n178) );
  AND U157 ( .A(n179), .B(n180), .Z(n177) );
  NAND U158 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U159 ( .A(A[211]), .B(B[211]), .Z(n182) );
  AND U160 ( .A(n183), .B(n184), .Z(n181) );
  NANDN U161 ( .A(A[210]), .B(B[210]), .Z(n184) );
  NAND U162 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U163 ( .A(B[210]), .B(A[210]), .Z(n186) );
  AND U164 ( .A(n187), .B(n188), .Z(n185) );
  NAND U165 ( .A(n189), .B(n190), .Z(n188) );
  NANDN U166 ( .A(A[209]), .B(B[209]), .Z(n190) );
  AND U167 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U168 ( .A(A[208]), .B(B[208]), .Z(n192) );
  NAND U169 ( .A(n193), .B(n194), .Z(n191) );
  NANDN U170 ( .A(B[208]), .B(A[208]), .Z(n194) );
  AND U171 ( .A(n195), .B(n196), .Z(n193) );
  NAND U172 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U173 ( .A(A[207]), .B(B[207]), .Z(n198) );
  AND U174 ( .A(n199), .B(n200), .Z(n197) );
  NANDN U175 ( .A(A[206]), .B(B[206]), .Z(n200) );
  NAND U176 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U177 ( .A(B[206]), .B(A[206]), .Z(n202) );
  AND U178 ( .A(n203), .B(n204), .Z(n201) );
  NAND U179 ( .A(n205), .B(n206), .Z(n204) );
  NANDN U180 ( .A(A[205]), .B(B[205]), .Z(n206) );
  AND U181 ( .A(n207), .B(n208), .Z(n205) );
  NANDN U182 ( .A(A[204]), .B(B[204]), .Z(n208) );
  NAND U183 ( .A(n209), .B(n210), .Z(n207) );
  NANDN U184 ( .A(B[204]), .B(A[204]), .Z(n210) );
  AND U185 ( .A(n211), .B(n212), .Z(n209) );
  NAND U186 ( .A(n213), .B(n214), .Z(n212) );
  NANDN U187 ( .A(A[203]), .B(B[203]), .Z(n214) );
  AND U188 ( .A(n215), .B(n216), .Z(n213) );
  NANDN U189 ( .A(A[202]), .B(B[202]), .Z(n216) );
  NAND U190 ( .A(n217), .B(n218), .Z(n215) );
  NANDN U191 ( .A(B[202]), .B(A[202]), .Z(n218) );
  AND U192 ( .A(n219), .B(n220), .Z(n217) );
  NAND U193 ( .A(n221), .B(n222), .Z(n220) );
  NANDN U194 ( .A(A[201]), .B(B[201]), .Z(n222) );
  AND U195 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U196 ( .A(A[200]), .B(B[200]), .Z(n224) );
  NAND U197 ( .A(n225), .B(n226), .Z(n223) );
  NANDN U198 ( .A(B[200]), .B(A[200]), .Z(n226) );
  AND U199 ( .A(n227), .B(n228), .Z(n225) );
  NAND U200 ( .A(n229), .B(n230), .Z(n228) );
  NANDN U201 ( .A(A[199]), .B(B[199]), .Z(n230) );
  AND U202 ( .A(n231), .B(n232), .Z(n229) );
  NANDN U203 ( .A(A[198]), .B(B[198]), .Z(n232) );
  NAND U204 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U205 ( .A(B[198]), .B(A[198]), .Z(n234) );
  AND U206 ( .A(n235), .B(n236), .Z(n233) );
  NAND U207 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U208 ( .A(A[197]), .B(B[197]), .Z(n238) );
  AND U209 ( .A(n239), .B(n240), .Z(n237) );
  NANDN U210 ( .A(A[196]), .B(B[196]), .Z(n240) );
  NAND U211 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U212 ( .A(B[196]), .B(A[196]), .Z(n242) );
  AND U213 ( .A(n243), .B(n244), .Z(n241) );
  NAND U214 ( .A(n245), .B(n246), .Z(n244) );
  NANDN U215 ( .A(A[195]), .B(B[195]), .Z(n246) );
  AND U216 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U217 ( .A(A[194]), .B(B[194]), .Z(n248) );
  NAND U218 ( .A(n249), .B(n250), .Z(n247) );
  NANDN U219 ( .A(B[194]), .B(A[194]), .Z(n250) );
  AND U220 ( .A(n251), .B(n252), .Z(n249) );
  NAND U221 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U222 ( .A(A[193]), .B(B[193]), .Z(n254) );
  AND U223 ( .A(n255), .B(n256), .Z(n253) );
  NANDN U224 ( .A(A[192]), .B(B[192]), .Z(n256) );
  NAND U225 ( .A(n257), .B(n258), .Z(n255) );
  NANDN U226 ( .A(B[192]), .B(A[192]), .Z(n258) );
  AND U227 ( .A(n259), .B(n260), .Z(n257) );
  NAND U228 ( .A(n261), .B(n262), .Z(n260) );
  NANDN U229 ( .A(A[191]), .B(B[191]), .Z(n262) );
  AND U230 ( .A(n263), .B(n264), .Z(n261) );
  NANDN U231 ( .A(A[190]), .B(B[190]), .Z(n264) );
  NAND U232 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U233 ( .A(B[190]), .B(A[190]), .Z(n266) );
  AND U234 ( .A(n267), .B(n268), .Z(n265) );
  NAND U235 ( .A(n269), .B(n270), .Z(n268) );
  NANDN U236 ( .A(A[189]), .B(B[189]), .Z(n270) );
  AND U237 ( .A(n271), .B(n272), .Z(n269) );
  NANDN U238 ( .A(A[188]), .B(B[188]), .Z(n272) );
  NAND U239 ( .A(n273), .B(n274), .Z(n271) );
  NANDN U240 ( .A(B[188]), .B(A[188]), .Z(n274) );
  AND U241 ( .A(n275), .B(n276), .Z(n273) );
  NAND U242 ( .A(n277), .B(n278), .Z(n276) );
  NANDN U243 ( .A(A[187]), .B(B[187]), .Z(n278) );
  AND U244 ( .A(n279), .B(n280), .Z(n277) );
  NANDN U245 ( .A(A[186]), .B(B[186]), .Z(n280) );
  NAND U246 ( .A(n281), .B(n282), .Z(n279) );
  NANDN U247 ( .A(B[186]), .B(A[186]), .Z(n282) );
  AND U248 ( .A(n283), .B(n284), .Z(n281) );
  NAND U249 ( .A(n285), .B(n286), .Z(n284) );
  NANDN U250 ( .A(A[185]), .B(B[185]), .Z(n286) );
  AND U251 ( .A(n287), .B(n288), .Z(n285) );
  NANDN U252 ( .A(A[184]), .B(B[184]), .Z(n288) );
  NAND U253 ( .A(n289), .B(n290), .Z(n287) );
  NANDN U254 ( .A(B[184]), .B(A[184]), .Z(n290) );
  AND U255 ( .A(n291), .B(n292), .Z(n289) );
  NAND U256 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U257 ( .A(A[183]), .B(B[183]), .Z(n294) );
  AND U258 ( .A(n295), .B(n296), .Z(n293) );
  NANDN U259 ( .A(A[182]), .B(B[182]), .Z(n296) );
  NAND U260 ( .A(n297), .B(n298), .Z(n295) );
  NANDN U261 ( .A(B[182]), .B(A[182]), .Z(n298) );
  AND U262 ( .A(n299), .B(n300), .Z(n297) );
  NAND U263 ( .A(n301), .B(n302), .Z(n300) );
  NANDN U264 ( .A(A[181]), .B(B[181]), .Z(n302) );
  AND U265 ( .A(n303), .B(n304), .Z(n301) );
  NANDN U266 ( .A(A[180]), .B(B[180]), .Z(n304) );
  NAND U267 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U268 ( .A(B[180]), .B(A[180]), .Z(n306) );
  AND U269 ( .A(n307), .B(n308), .Z(n305) );
  NAND U270 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U271 ( .A(A[179]), .B(B[179]), .Z(n310) );
  AND U272 ( .A(n311), .B(n312), .Z(n309) );
  NANDN U273 ( .A(A[178]), .B(B[178]), .Z(n312) );
  NAND U274 ( .A(n313), .B(n314), .Z(n311) );
  NANDN U275 ( .A(B[178]), .B(A[178]), .Z(n314) );
  AND U276 ( .A(n315), .B(n316), .Z(n313) );
  NAND U277 ( .A(n317), .B(n318), .Z(n316) );
  NANDN U278 ( .A(A[177]), .B(B[177]), .Z(n318) );
  AND U279 ( .A(n319), .B(n320), .Z(n317) );
  NANDN U280 ( .A(A[176]), .B(B[176]), .Z(n320) );
  NAND U281 ( .A(n321), .B(n322), .Z(n319) );
  NANDN U282 ( .A(B[176]), .B(A[176]), .Z(n322) );
  AND U283 ( .A(n323), .B(n324), .Z(n321) );
  NAND U284 ( .A(n325), .B(n326), .Z(n324) );
  NANDN U285 ( .A(A[175]), .B(B[175]), .Z(n326) );
  AND U286 ( .A(n327), .B(n328), .Z(n325) );
  NANDN U287 ( .A(A[174]), .B(B[174]), .Z(n328) );
  NAND U288 ( .A(n329), .B(n330), .Z(n327) );
  NANDN U289 ( .A(B[174]), .B(A[174]), .Z(n330) );
  AND U290 ( .A(n331), .B(n332), .Z(n329) );
  NAND U291 ( .A(n333), .B(n334), .Z(n332) );
  NANDN U292 ( .A(A[173]), .B(B[173]), .Z(n334) );
  AND U293 ( .A(n335), .B(n336), .Z(n333) );
  NANDN U294 ( .A(A[172]), .B(B[172]), .Z(n336) );
  NAND U295 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U296 ( .A(B[172]), .B(A[172]), .Z(n338) );
  AND U297 ( .A(n339), .B(n340), .Z(n337) );
  NAND U298 ( .A(n341), .B(n342), .Z(n340) );
  NANDN U299 ( .A(A[171]), .B(B[171]), .Z(n342) );
  AND U300 ( .A(n343), .B(n344), .Z(n341) );
  NANDN U301 ( .A(A[170]), .B(B[170]), .Z(n344) );
  NAND U302 ( .A(n345), .B(n346), .Z(n343) );
  NANDN U303 ( .A(B[170]), .B(A[170]), .Z(n346) );
  AND U304 ( .A(n347), .B(n348), .Z(n345) );
  NAND U305 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U306 ( .A(A[169]), .B(B[169]), .Z(n350) );
  AND U307 ( .A(n351), .B(n352), .Z(n349) );
  NANDN U308 ( .A(A[168]), .B(B[168]), .Z(n352) );
  NAND U309 ( .A(n353), .B(n354), .Z(n351) );
  NANDN U310 ( .A(B[168]), .B(A[168]), .Z(n354) );
  AND U311 ( .A(n355), .B(n356), .Z(n353) );
  NAND U312 ( .A(n357), .B(n358), .Z(n356) );
  NANDN U313 ( .A(A[167]), .B(B[167]), .Z(n358) );
  AND U314 ( .A(n359), .B(n360), .Z(n357) );
  NANDN U315 ( .A(A[166]), .B(B[166]), .Z(n360) );
  NAND U316 ( .A(n361), .B(n362), .Z(n359) );
  NANDN U317 ( .A(B[166]), .B(A[166]), .Z(n362) );
  AND U318 ( .A(n363), .B(n364), .Z(n361) );
  NAND U319 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U320 ( .A(A[165]), .B(B[165]), .Z(n366) );
  AND U321 ( .A(n367), .B(n368), .Z(n365) );
  NANDN U322 ( .A(A[164]), .B(B[164]), .Z(n368) );
  NAND U323 ( .A(n369), .B(n370), .Z(n367) );
  NANDN U324 ( .A(B[164]), .B(A[164]), .Z(n370) );
  AND U325 ( .A(n371), .B(n372), .Z(n369) );
  NAND U326 ( .A(n373), .B(n374), .Z(n372) );
  NANDN U327 ( .A(A[163]), .B(B[163]), .Z(n374) );
  AND U328 ( .A(n375), .B(n376), .Z(n373) );
  NANDN U329 ( .A(A[162]), .B(B[162]), .Z(n376) );
  NAND U330 ( .A(n377), .B(n378), .Z(n375) );
  NANDN U331 ( .A(B[162]), .B(A[162]), .Z(n378) );
  AND U332 ( .A(n379), .B(n380), .Z(n377) );
  NAND U333 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U334 ( .A(A[161]), .B(B[161]), .Z(n382) );
  AND U335 ( .A(n383), .B(n384), .Z(n381) );
  NANDN U336 ( .A(A[160]), .B(B[160]), .Z(n384) );
  NAND U337 ( .A(n385), .B(n386), .Z(n383) );
  NANDN U338 ( .A(B[160]), .B(A[160]), .Z(n386) );
  AND U339 ( .A(n387), .B(n388), .Z(n385) );
  NAND U340 ( .A(n389), .B(n390), .Z(n388) );
  NANDN U341 ( .A(A[159]), .B(B[159]), .Z(n390) );
  AND U342 ( .A(n391), .B(n392), .Z(n389) );
  NANDN U343 ( .A(A[158]), .B(B[158]), .Z(n392) );
  NAND U344 ( .A(n393), .B(n394), .Z(n391) );
  NANDN U345 ( .A(B[158]), .B(A[158]), .Z(n394) );
  AND U346 ( .A(n395), .B(n396), .Z(n393) );
  NAND U347 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U348 ( .A(A[157]), .B(B[157]), .Z(n398) );
  AND U349 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U350 ( .A(A[156]), .B(B[156]), .Z(n400) );
  NAND U351 ( .A(n401), .B(n402), .Z(n399) );
  NANDN U352 ( .A(B[156]), .B(A[156]), .Z(n402) );
  AND U353 ( .A(n403), .B(n404), .Z(n401) );
  NAND U354 ( .A(n405), .B(n406), .Z(n404) );
  NANDN U355 ( .A(A[155]), .B(B[155]), .Z(n406) );
  AND U356 ( .A(n407), .B(n408), .Z(n405) );
  NANDN U357 ( .A(A[154]), .B(B[154]), .Z(n408) );
  NAND U358 ( .A(n409), .B(n410), .Z(n407) );
  NANDN U359 ( .A(B[154]), .B(A[154]), .Z(n410) );
  AND U360 ( .A(n411), .B(n412), .Z(n409) );
  NAND U361 ( .A(n413), .B(n414), .Z(n412) );
  NANDN U362 ( .A(A[153]), .B(B[153]), .Z(n414) );
  AND U363 ( .A(n415), .B(n416), .Z(n413) );
  NANDN U364 ( .A(A[152]), .B(B[152]), .Z(n416) );
  NAND U365 ( .A(n417), .B(n418), .Z(n415) );
  NANDN U366 ( .A(B[152]), .B(A[152]), .Z(n418) );
  AND U367 ( .A(n419), .B(n420), .Z(n417) );
  NAND U368 ( .A(n421), .B(n422), .Z(n420) );
  NANDN U369 ( .A(A[151]), .B(B[151]), .Z(n422) );
  AND U370 ( .A(n423), .B(n424), .Z(n421) );
  NANDN U371 ( .A(A[150]), .B(B[150]), .Z(n424) );
  NAND U372 ( .A(n425), .B(n426), .Z(n423) );
  NANDN U373 ( .A(B[150]), .B(A[150]), .Z(n426) );
  AND U374 ( .A(n427), .B(n428), .Z(n425) );
  NAND U375 ( .A(n429), .B(n430), .Z(n428) );
  NANDN U376 ( .A(A[149]), .B(B[149]), .Z(n430) );
  AND U377 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U378 ( .A(A[148]), .B(B[148]), .Z(n432) );
  NAND U379 ( .A(n433), .B(n434), .Z(n431) );
  NANDN U380 ( .A(B[148]), .B(A[148]), .Z(n434) );
  AND U381 ( .A(n435), .B(n436), .Z(n433) );
  NAND U382 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U383 ( .A(A[147]), .B(B[147]), .Z(n438) );
  AND U384 ( .A(n439), .B(n440), .Z(n437) );
  NANDN U385 ( .A(A[146]), .B(B[146]), .Z(n440) );
  NAND U386 ( .A(n441), .B(n442), .Z(n439) );
  NANDN U387 ( .A(B[146]), .B(A[146]), .Z(n442) );
  AND U388 ( .A(n443), .B(n444), .Z(n441) );
  NAND U389 ( .A(n445), .B(n446), .Z(n444) );
  NANDN U390 ( .A(A[145]), .B(B[145]), .Z(n446) );
  AND U391 ( .A(n447), .B(n448), .Z(n445) );
  NANDN U392 ( .A(A[144]), .B(B[144]), .Z(n448) );
  NAND U393 ( .A(n449), .B(n450), .Z(n447) );
  NANDN U394 ( .A(B[144]), .B(A[144]), .Z(n450) );
  AND U395 ( .A(n451), .B(n452), .Z(n449) );
  NAND U396 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U397 ( .A(A[143]), .B(B[143]), .Z(n454) );
  AND U398 ( .A(n455), .B(n456), .Z(n453) );
  NANDN U399 ( .A(A[142]), .B(B[142]), .Z(n456) );
  NAND U400 ( .A(n457), .B(n458), .Z(n455) );
  NANDN U401 ( .A(B[142]), .B(A[142]), .Z(n458) );
  AND U402 ( .A(n459), .B(n460), .Z(n457) );
  NAND U403 ( .A(n461), .B(n462), .Z(n460) );
  NANDN U404 ( .A(A[141]), .B(B[141]), .Z(n462) );
  AND U405 ( .A(n463), .B(n464), .Z(n461) );
  NANDN U406 ( .A(A[140]), .B(B[140]), .Z(n464) );
  NAND U407 ( .A(n465), .B(n466), .Z(n463) );
  NANDN U408 ( .A(B[140]), .B(A[140]), .Z(n466) );
  AND U409 ( .A(n467), .B(n468), .Z(n465) );
  NAND U410 ( .A(n469), .B(n470), .Z(n468) );
  NANDN U411 ( .A(A[139]), .B(B[139]), .Z(n470) );
  AND U412 ( .A(n471), .B(n472), .Z(n469) );
  NANDN U413 ( .A(A[138]), .B(B[138]), .Z(n472) );
  NAND U414 ( .A(n473), .B(n474), .Z(n471) );
  NANDN U415 ( .A(B[138]), .B(A[138]), .Z(n474) );
  AND U416 ( .A(n475), .B(n476), .Z(n473) );
  NAND U417 ( .A(n477), .B(n478), .Z(n476) );
  NANDN U418 ( .A(A[137]), .B(B[137]), .Z(n478) );
  AND U419 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U420 ( .A(A[136]), .B(B[136]), .Z(n480) );
  NAND U421 ( .A(n481), .B(n482), .Z(n479) );
  NANDN U422 ( .A(B[136]), .B(A[136]), .Z(n482) );
  AND U423 ( .A(n483), .B(n484), .Z(n481) );
  NAND U424 ( .A(n485), .B(n486), .Z(n484) );
  NANDN U425 ( .A(A[135]), .B(B[135]), .Z(n486) );
  AND U426 ( .A(n487), .B(n488), .Z(n485) );
  NANDN U427 ( .A(A[134]), .B(B[134]), .Z(n488) );
  NAND U428 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U429 ( .A(B[134]), .B(A[134]), .Z(n490) );
  AND U430 ( .A(n491), .B(n492), .Z(n489) );
  NAND U431 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U432 ( .A(A[133]), .B(B[133]), .Z(n494) );
  AND U433 ( .A(n495), .B(n496), .Z(n493) );
  NANDN U434 ( .A(A[132]), .B(B[132]), .Z(n496) );
  NAND U435 ( .A(n497), .B(n498), .Z(n495) );
  NANDN U436 ( .A(B[132]), .B(A[132]), .Z(n498) );
  AND U437 ( .A(n499), .B(n500), .Z(n497) );
  NAND U438 ( .A(n501), .B(n502), .Z(n500) );
  NANDN U439 ( .A(A[131]), .B(B[131]), .Z(n502) );
  AND U440 ( .A(n503), .B(n504), .Z(n501) );
  NANDN U441 ( .A(A[130]), .B(B[130]), .Z(n504) );
  NAND U442 ( .A(n505), .B(n506), .Z(n503) );
  NANDN U443 ( .A(B[130]), .B(A[130]), .Z(n506) );
  AND U444 ( .A(n507), .B(n508), .Z(n505) );
  NAND U445 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U446 ( .A(A[129]), .B(B[129]), .Z(n510) );
  AND U447 ( .A(n511), .B(n512), .Z(n509) );
  NANDN U448 ( .A(A[128]), .B(B[128]), .Z(n512) );
  NAND U449 ( .A(n513), .B(n514), .Z(n511) );
  NANDN U450 ( .A(B[128]), .B(A[128]), .Z(n514) );
  AND U451 ( .A(n515), .B(n516), .Z(n513) );
  NAND U452 ( .A(n517), .B(n518), .Z(n516) );
  NANDN U453 ( .A(A[127]), .B(B[127]), .Z(n518) );
  AND U454 ( .A(n519), .B(n520), .Z(n517) );
  NANDN U455 ( .A(A[126]), .B(B[126]), .Z(n520) );
  NAND U456 ( .A(n521), .B(n522), .Z(n519) );
  NANDN U457 ( .A(B[126]), .B(A[126]), .Z(n522) );
  AND U458 ( .A(n523), .B(n524), .Z(n521) );
  NAND U459 ( .A(n525), .B(n526), .Z(n524) );
  NANDN U460 ( .A(A[125]), .B(B[125]), .Z(n526) );
  AND U461 ( .A(n527), .B(n528), .Z(n525) );
  NANDN U462 ( .A(A[124]), .B(B[124]), .Z(n528) );
  NAND U463 ( .A(n529), .B(n530), .Z(n527) );
  NANDN U464 ( .A(B[124]), .B(A[124]), .Z(n530) );
  AND U465 ( .A(n531), .B(n532), .Z(n529) );
  NAND U466 ( .A(n533), .B(n534), .Z(n532) );
  NANDN U467 ( .A(A[123]), .B(B[123]), .Z(n534) );
  AND U468 ( .A(n535), .B(n536), .Z(n533) );
  NANDN U469 ( .A(A[122]), .B(B[122]), .Z(n536) );
  NAND U470 ( .A(n537), .B(n538), .Z(n535) );
  NANDN U471 ( .A(B[122]), .B(A[122]), .Z(n538) );
  AND U472 ( .A(n539), .B(n540), .Z(n537) );
  NAND U473 ( .A(n541), .B(n542), .Z(n540) );
  NANDN U474 ( .A(A[121]), .B(B[121]), .Z(n542) );
  AND U475 ( .A(n543), .B(n544), .Z(n541) );
  NANDN U476 ( .A(A[120]), .B(B[120]), .Z(n544) );
  NAND U477 ( .A(n545), .B(n546), .Z(n543) );
  NANDN U478 ( .A(B[120]), .B(A[120]), .Z(n546) );
  AND U479 ( .A(n547), .B(n548), .Z(n545) );
  NAND U480 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U481 ( .A(A[119]), .B(B[119]), .Z(n550) );
  AND U482 ( .A(n551), .B(n552), .Z(n549) );
  NANDN U483 ( .A(A[118]), .B(B[118]), .Z(n552) );
  NAND U484 ( .A(n553), .B(n554), .Z(n551) );
  NANDN U485 ( .A(B[118]), .B(A[118]), .Z(n554) );
  AND U486 ( .A(n555), .B(n556), .Z(n553) );
  NAND U487 ( .A(n557), .B(n558), .Z(n556) );
  NANDN U488 ( .A(A[117]), .B(B[117]), .Z(n558) );
  AND U489 ( .A(n559), .B(n560), .Z(n557) );
  NANDN U490 ( .A(A[116]), .B(B[116]), .Z(n560) );
  NAND U491 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U492 ( .A(B[116]), .B(A[116]), .Z(n562) );
  AND U493 ( .A(n563), .B(n564), .Z(n561) );
  NAND U494 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U495 ( .A(A[115]), .B(B[115]), .Z(n566) );
  AND U496 ( .A(n567), .B(n568), .Z(n565) );
  NANDN U497 ( .A(A[114]), .B(B[114]), .Z(n568) );
  NAND U498 ( .A(n569), .B(n570), .Z(n567) );
  NANDN U499 ( .A(B[114]), .B(A[114]), .Z(n570) );
  AND U500 ( .A(n571), .B(n572), .Z(n569) );
  NAND U501 ( .A(n573), .B(n574), .Z(n572) );
  NANDN U502 ( .A(A[113]), .B(B[113]), .Z(n574) );
  AND U503 ( .A(n575), .B(n576), .Z(n573) );
  NANDN U504 ( .A(A[112]), .B(B[112]), .Z(n576) );
  NAND U505 ( .A(n577), .B(n578), .Z(n575) );
  NANDN U506 ( .A(B[112]), .B(A[112]), .Z(n578) );
  AND U507 ( .A(n579), .B(n580), .Z(n577) );
  NAND U508 ( .A(n581), .B(n582), .Z(n580) );
  NANDN U509 ( .A(A[111]), .B(B[111]), .Z(n582) );
  AND U510 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U511 ( .A(A[110]), .B(B[110]), .Z(n584) );
  NAND U512 ( .A(n585), .B(n586), .Z(n583) );
  NANDN U513 ( .A(B[110]), .B(A[110]), .Z(n586) );
  AND U514 ( .A(n587), .B(n588), .Z(n585) );
  NAND U515 ( .A(n589), .B(n590), .Z(n588) );
  NANDN U516 ( .A(A[109]), .B(B[109]), .Z(n590) );
  AND U517 ( .A(n591), .B(n592), .Z(n589) );
  NANDN U518 ( .A(A[108]), .B(B[108]), .Z(n592) );
  NAND U519 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U520 ( .A(B[108]), .B(A[108]), .Z(n594) );
  AND U521 ( .A(n595), .B(n596), .Z(n593) );
  NAND U522 ( .A(n597), .B(n598), .Z(n596) );
  NANDN U523 ( .A(A[107]), .B(B[107]), .Z(n598) );
  AND U524 ( .A(n599), .B(n600), .Z(n597) );
  NANDN U525 ( .A(A[106]), .B(B[106]), .Z(n600) );
  NAND U526 ( .A(n601), .B(n602), .Z(n599) );
  NANDN U527 ( .A(B[106]), .B(A[106]), .Z(n602) );
  AND U528 ( .A(n603), .B(n604), .Z(n601) );
  NAND U529 ( .A(n605), .B(n606), .Z(n604) );
  NANDN U530 ( .A(A[105]), .B(B[105]), .Z(n606) );
  AND U531 ( .A(n607), .B(n608), .Z(n605) );
  NANDN U532 ( .A(A[104]), .B(B[104]), .Z(n608) );
  NAND U533 ( .A(n609), .B(n610), .Z(n607) );
  NANDN U534 ( .A(B[104]), .B(A[104]), .Z(n610) );
  AND U535 ( .A(n611), .B(n612), .Z(n609) );
  NAND U536 ( .A(n613), .B(n614), .Z(n612) );
  NANDN U537 ( .A(A[103]), .B(B[103]), .Z(n614) );
  AND U538 ( .A(n615), .B(n616), .Z(n613) );
  NANDN U539 ( .A(A[102]), .B(B[102]), .Z(n616) );
  NAND U540 ( .A(n617), .B(n618), .Z(n615) );
  NANDN U541 ( .A(B[102]), .B(A[102]), .Z(n618) );
  AND U542 ( .A(n619), .B(n620), .Z(n617) );
  NAND U543 ( .A(n621), .B(n622), .Z(n620) );
  NANDN U544 ( .A(A[101]), .B(B[101]), .Z(n622) );
  AND U545 ( .A(n623), .B(n624), .Z(n621) );
  NANDN U546 ( .A(A[100]), .B(B[100]), .Z(n624) );
  NAND U547 ( .A(n625), .B(n626), .Z(n623) );
  NANDN U548 ( .A(B[99]), .B(A[99]), .Z(n626) );
  AND U549 ( .A(n627), .B(n628), .Z(n625) );
  NAND U550 ( .A(n629), .B(n630), .Z(n628) );
  NANDN U551 ( .A(A[99]), .B(B[99]), .Z(n630) );
  AND U552 ( .A(n631), .B(n632), .Z(n629) );
  NANDN U553 ( .A(A[98]), .B(B[98]), .Z(n632) );
  NAND U554 ( .A(n633), .B(n634), .Z(n631) );
  NANDN U555 ( .A(B[98]), .B(A[98]), .Z(n634) );
  AND U556 ( .A(n635), .B(n636), .Z(n633) );
  NAND U557 ( .A(n637), .B(n638), .Z(n636) );
  NANDN U558 ( .A(A[97]), .B(B[97]), .Z(n638) );
  AND U559 ( .A(n639), .B(n640), .Z(n637) );
  NANDN U560 ( .A(A[96]), .B(B[96]), .Z(n640) );
  NAND U561 ( .A(n641), .B(n642), .Z(n639) );
  NANDN U562 ( .A(B[96]), .B(A[96]), .Z(n642) );
  AND U563 ( .A(n643), .B(n644), .Z(n641) );
  NAND U564 ( .A(n645), .B(n646), .Z(n644) );
  NANDN U565 ( .A(A[95]), .B(B[95]), .Z(n646) );
  AND U566 ( .A(n647), .B(n648), .Z(n645) );
  NANDN U567 ( .A(A[94]), .B(B[94]), .Z(n648) );
  NAND U568 ( .A(n649), .B(n650), .Z(n647) );
  NANDN U569 ( .A(B[94]), .B(A[94]), .Z(n650) );
  AND U570 ( .A(n651), .B(n652), .Z(n649) );
  NAND U571 ( .A(n653), .B(n654), .Z(n652) );
  NANDN U572 ( .A(A[93]), .B(B[93]), .Z(n654) );
  AND U573 ( .A(n655), .B(n656), .Z(n653) );
  NANDN U574 ( .A(A[92]), .B(B[92]), .Z(n656) );
  NAND U575 ( .A(n657), .B(n658), .Z(n655) );
  NANDN U576 ( .A(B[92]), .B(A[92]), .Z(n658) );
  AND U577 ( .A(n659), .B(n660), .Z(n657) );
  NAND U578 ( .A(n661), .B(n662), .Z(n660) );
  NANDN U579 ( .A(A[91]), .B(B[91]), .Z(n662) );
  AND U580 ( .A(n663), .B(n664), .Z(n661) );
  NANDN U581 ( .A(A[90]), .B(B[90]), .Z(n664) );
  NAND U582 ( .A(n665), .B(n666), .Z(n663) );
  NANDN U583 ( .A(B[90]), .B(A[90]), .Z(n666) );
  AND U584 ( .A(n667), .B(n668), .Z(n665) );
  NAND U585 ( .A(n669), .B(n670), .Z(n668) );
  NANDN U586 ( .A(A[89]), .B(B[89]), .Z(n670) );
  AND U587 ( .A(n671), .B(n672), .Z(n669) );
  NANDN U588 ( .A(A[88]), .B(B[88]), .Z(n672) );
  NAND U589 ( .A(n673), .B(n674), .Z(n671) );
  NANDN U590 ( .A(B[88]), .B(A[88]), .Z(n674) );
  AND U591 ( .A(n675), .B(n676), .Z(n673) );
  NAND U592 ( .A(n677), .B(n678), .Z(n676) );
  NANDN U593 ( .A(A[87]), .B(B[87]), .Z(n678) );
  AND U594 ( .A(n679), .B(n680), .Z(n677) );
  NANDN U595 ( .A(A[86]), .B(B[86]), .Z(n680) );
  NAND U596 ( .A(n681), .B(n682), .Z(n679) );
  NANDN U597 ( .A(B[86]), .B(A[86]), .Z(n682) );
  AND U598 ( .A(n683), .B(n684), .Z(n681) );
  NAND U599 ( .A(n685), .B(n686), .Z(n684) );
  NANDN U600 ( .A(A[85]), .B(B[85]), .Z(n686) );
  AND U601 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U602 ( .A(A[84]), .B(B[84]), .Z(n688) );
  NAND U603 ( .A(n689), .B(n690), .Z(n687) );
  NANDN U604 ( .A(B[84]), .B(A[84]), .Z(n690) );
  AND U605 ( .A(n691), .B(n692), .Z(n689) );
  NAND U606 ( .A(n693), .B(n694), .Z(n692) );
  NANDN U607 ( .A(A[83]), .B(B[83]), .Z(n694) );
  AND U608 ( .A(n695), .B(n696), .Z(n693) );
  NANDN U609 ( .A(A[82]), .B(B[82]), .Z(n696) );
  NAND U610 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U611 ( .A(B[82]), .B(A[82]), .Z(n698) );
  AND U612 ( .A(n699), .B(n700), .Z(n697) );
  NAND U613 ( .A(n701), .B(n702), .Z(n700) );
  NANDN U614 ( .A(A[81]), .B(B[81]), .Z(n702) );
  AND U615 ( .A(n703), .B(n704), .Z(n701) );
  NANDN U616 ( .A(A[80]), .B(B[80]), .Z(n704) );
  NAND U617 ( .A(n705), .B(n706), .Z(n703) );
  NANDN U618 ( .A(B[80]), .B(A[80]), .Z(n706) );
  AND U619 ( .A(n707), .B(n708), .Z(n705) );
  NAND U620 ( .A(n709), .B(n710), .Z(n708) );
  NANDN U621 ( .A(A[79]), .B(B[79]), .Z(n710) );
  AND U622 ( .A(n711), .B(n712), .Z(n709) );
  NANDN U623 ( .A(A[78]), .B(B[78]), .Z(n712) );
  NAND U624 ( .A(n713), .B(n714), .Z(n711) );
  NANDN U625 ( .A(B[78]), .B(A[78]), .Z(n714) );
  AND U626 ( .A(n715), .B(n716), .Z(n713) );
  NAND U627 ( .A(n717), .B(n718), .Z(n716) );
  NANDN U628 ( .A(A[77]), .B(B[77]), .Z(n718) );
  AND U629 ( .A(n719), .B(n720), .Z(n717) );
  NANDN U630 ( .A(A[76]), .B(B[76]), .Z(n720) );
  NAND U631 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U632 ( .A(B[76]), .B(A[76]), .Z(n722) );
  AND U633 ( .A(n723), .B(n724), .Z(n721) );
  NAND U634 ( .A(n725), .B(n726), .Z(n724) );
  NANDN U635 ( .A(A[75]), .B(B[75]), .Z(n726) );
  AND U636 ( .A(n727), .B(n728), .Z(n725) );
  NANDN U637 ( .A(A[74]), .B(B[74]), .Z(n728) );
  NAND U638 ( .A(n729), .B(n730), .Z(n727) );
  NANDN U639 ( .A(B[74]), .B(A[74]), .Z(n730) );
  AND U640 ( .A(n731), .B(n732), .Z(n729) );
  NAND U641 ( .A(n733), .B(n734), .Z(n732) );
  NANDN U642 ( .A(A[73]), .B(B[73]), .Z(n734) );
  AND U643 ( .A(n735), .B(n736), .Z(n733) );
  NANDN U644 ( .A(A[72]), .B(B[72]), .Z(n736) );
  NAND U645 ( .A(n737), .B(n738), .Z(n735) );
  NANDN U646 ( .A(B[72]), .B(A[72]), .Z(n738) );
  AND U647 ( .A(n739), .B(n740), .Z(n737) );
  NAND U648 ( .A(n741), .B(n742), .Z(n740) );
  NANDN U649 ( .A(A[71]), .B(B[71]), .Z(n742) );
  AND U650 ( .A(n743), .B(n744), .Z(n741) );
  NANDN U651 ( .A(A[70]), .B(B[70]), .Z(n744) );
  NAND U652 ( .A(n745), .B(n746), .Z(n743) );
  NANDN U653 ( .A(B[70]), .B(A[70]), .Z(n746) );
  AND U654 ( .A(n747), .B(n748), .Z(n745) );
  NAND U655 ( .A(n749), .B(n750), .Z(n748) );
  NANDN U656 ( .A(A[69]), .B(B[69]), .Z(n750) );
  AND U657 ( .A(n751), .B(n752), .Z(n749) );
  NANDN U658 ( .A(A[68]), .B(B[68]), .Z(n752) );
  NAND U659 ( .A(n753), .B(n754), .Z(n751) );
  NANDN U660 ( .A(B[68]), .B(A[68]), .Z(n754) );
  AND U661 ( .A(n755), .B(n756), .Z(n753) );
  NAND U662 ( .A(n757), .B(n758), .Z(n756) );
  NANDN U663 ( .A(A[67]), .B(B[67]), .Z(n758) );
  AND U664 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U665 ( .A(A[66]), .B(B[66]), .Z(n760) );
  NAND U666 ( .A(n761), .B(n762), .Z(n759) );
  NANDN U667 ( .A(B[66]), .B(A[66]), .Z(n762) );
  AND U668 ( .A(n763), .B(n764), .Z(n761) );
  NAND U669 ( .A(n765), .B(n766), .Z(n764) );
  NANDN U670 ( .A(A[65]), .B(B[65]), .Z(n766) );
  AND U671 ( .A(n767), .B(n768), .Z(n765) );
  NANDN U672 ( .A(A[64]), .B(B[64]), .Z(n768) );
  NAND U673 ( .A(n769), .B(n770), .Z(n767) );
  NANDN U674 ( .A(B[64]), .B(A[64]), .Z(n770) );
  AND U675 ( .A(n771), .B(n772), .Z(n769) );
  NAND U676 ( .A(n773), .B(n774), .Z(n772) );
  NANDN U677 ( .A(A[63]), .B(B[63]), .Z(n774) );
  AND U678 ( .A(n775), .B(n776), .Z(n773) );
  NANDN U679 ( .A(A[62]), .B(B[62]), .Z(n776) );
  NAND U680 ( .A(n777), .B(n778), .Z(n775) );
  NANDN U681 ( .A(B[62]), .B(A[62]), .Z(n778) );
  AND U682 ( .A(n779), .B(n780), .Z(n777) );
  NAND U683 ( .A(n781), .B(n782), .Z(n780) );
  NANDN U684 ( .A(A[61]), .B(B[61]), .Z(n782) );
  AND U685 ( .A(n783), .B(n784), .Z(n781) );
  NANDN U686 ( .A(A[60]), .B(B[60]), .Z(n784) );
  NAND U687 ( .A(n785), .B(n786), .Z(n783) );
  NANDN U688 ( .A(B[60]), .B(A[60]), .Z(n786) );
  AND U689 ( .A(n787), .B(n788), .Z(n785) );
  NAND U690 ( .A(n789), .B(n790), .Z(n788) );
  NANDN U691 ( .A(A[59]), .B(B[59]), .Z(n790) );
  AND U692 ( .A(n791), .B(n792), .Z(n789) );
  NANDN U693 ( .A(A[58]), .B(B[58]), .Z(n792) );
  NAND U694 ( .A(n793), .B(n794), .Z(n791) );
  NANDN U695 ( .A(B[58]), .B(A[58]), .Z(n794) );
  AND U696 ( .A(n795), .B(n796), .Z(n793) );
  NAND U697 ( .A(n797), .B(n798), .Z(n796) );
  NANDN U698 ( .A(A[57]), .B(B[57]), .Z(n798) );
  AND U699 ( .A(n799), .B(n800), .Z(n797) );
  NANDN U700 ( .A(A[56]), .B(B[56]), .Z(n800) );
  NAND U701 ( .A(n801), .B(n802), .Z(n799) );
  NANDN U702 ( .A(B[56]), .B(A[56]), .Z(n802) );
  AND U703 ( .A(n803), .B(n804), .Z(n801) );
  NAND U704 ( .A(n805), .B(n806), .Z(n804) );
  NANDN U705 ( .A(A[55]), .B(B[55]), .Z(n806) );
  AND U706 ( .A(n807), .B(n808), .Z(n805) );
  NANDN U707 ( .A(A[54]), .B(B[54]), .Z(n808) );
  NAND U708 ( .A(n809), .B(n810), .Z(n807) );
  NANDN U709 ( .A(B[54]), .B(A[54]), .Z(n810) );
  AND U710 ( .A(n811), .B(n812), .Z(n809) );
  NAND U711 ( .A(n813), .B(n814), .Z(n812) );
  NANDN U712 ( .A(A[53]), .B(B[53]), .Z(n814) );
  AND U713 ( .A(n815), .B(n816), .Z(n813) );
  NANDN U714 ( .A(A[52]), .B(B[52]), .Z(n816) );
  NAND U715 ( .A(n817), .B(n818), .Z(n815) );
  NANDN U716 ( .A(B[52]), .B(A[52]), .Z(n818) );
  AND U717 ( .A(n819), .B(n820), .Z(n817) );
  NAND U718 ( .A(n821), .B(n822), .Z(n820) );
  NANDN U719 ( .A(A[51]), .B(B[51]), .Z(n822) );
  AND U720 ( .A(n823), .B(n824), .Z(n821) );
  NANDN U721 ( .A(A[50]), .B(B[50]), .Z(n824) );
  NAND U722 ( .A(n825), .B(n826), .Z(n823) );
  NANDN U723 ( .A(B[50]), .B(A[50]), .Z(n826) );
  AND U724 ( .A(n827), .B(n828), .Z(n825) );
  NAND U725 ( .A(n829), .B(n830), .Z(n828) );
  NANDN U726 ( .A(A[49]), .B(B[49]), .Z(n830) );
  AND U727 ( .A(n831), .B(n832), .Z(n829) );
  NANDN U728 ( .A(A[48]), .B(B[48]), .Z(n832) );
  NAND U729 ( .A(n833), .B(n834), .Z(n831) );
  NANDN U730 ( .A(B[48]), .B(A[48]), .Z(n834) );
  AND U731 ( .A(n835), .B(n836), .Z(n833) );
  NAND U732 ( .A(n837), .B(n838), .Z(n836) );
  NANDN U733 ( .A(A[47]), .B(B[47]), .Z(n838) );
  AND U734 ( .A(n839), .B(n840), .Z(n837) );
  NANDN U735 ( .A(A[46]), .B(B[46]), .Z(n840) );
  NAND U736 ( .A(n841), .B(n842), .Z(n839) );
  NANDN U737 ( .A(B[46]), .B(A[46]), .Z(n842) );
  AND U738 ( .A(n843), .B(n844), .Z(n841) );
  NAND U739 ( .A(n845), .B(n846), .Z(n844) );
  NANDN U740 ( .A(A[45]), .B(B[45]), .Z(n846) );
  AND U741 ( .A(n847), .B(n848), .Z(n845) );
  NANDN U742 ( .A(A[44]), .B(B[44]), .Z(n848) );
  NAND U743 ( .A(n849), .B(n850), .Z(n847) );
  NANDN U744 ( .A(B[44]), .B(A[44]), .Z(n850) );
  AND U745 ( .A(n851), .B(n852), .Z(n849) );
  NAND U746 ( .A(n853), .B(n854), .Z(n852) );
  NANDN U747 ( .A(A[43]), .B(B[43]), .Z(n854) );
  AND U748 ( .A(n855), .B(n856), .Z(n853) );
  NANDN U749 ( .A(A[42]), .B(B[42]), .Z(n856) );
  NAND U750 ( .A(n857), .B(n858), .Z(n855) );
  NANDN U751 ( .A(B[42]), .B(A[42]), .Z(n858) );
  AND U752 ( .A(n859), .B(n860), .Z(n857) );
  NAND U753 ( .A(n861), .B(n862), .Z(n860) );
  NANDN U754 ( .A(A[41]), .B(B[41]), .Z(n862) );
  AND U755 ( .A(n863), .B(n864), .Z(n861) );
  NANDN U756 ( .A(A[40]), .B(B[40]), .Z(n864) );
  NAND U757 ( .A(n865), .B(n866), .Z(n863) );
  NANDN U758 ( .A(B[40]), .B(A[40]), .Z(n866) );
  AND U759 ( .A(n867), .B(n868), .Z(n865) );
  NAND U760 ( .A(n869), .B(n870), .Z(n868) );
  NANDN U761 ( .A(A[39]), .B(B[39]), .Z(n870) );
  AND U762 ( .A(n871), .B(n872), .Z(n869) );
  NANDN U763 ( .A(A[38]), .B(B[38]), .Z(n872) );
  NAND U764 ( .A(n873), .B(n874), .Z(n871) );
  NANDN U765 ( .A(B[38]), .B(A[38]), .Z(n874) );
  AND U766 ( .A(n875), .B(n876), .Z(n873) );
  NAND U767 ( .A(n877), .B(n878), .Z(n876) );
  NANDN U768 ( .A(A[37]), .B(B[37]), .Z(n878) );
  AND U769 ( .A(n879), .B(n880), .Z(n877) );
  NANDN U770 ( .A(A[36]), .B(B[36]), .Z(n880) );
  NAND U771 ( .A(n881), .B(n882), .Z(n879) );
  NANDN U772 ( .A(B[36]), .B(A[36]), .Z(n882) );
  AND U773 ( .A(n883), .B(n884), .Z(n881) );
  NAND U774 ( .A(n885), .B(n886), .Z(n884) );
  NANDN U775 ( .A(A[35]), .B(B[35]), .Z(n886) );
  AND U776 ( .A(n887), .B(n888), .Z(n885) );
  NANDN U777 ( .A(A[34]), .B(B[34]), .Z(n888) );
  NAND U778 ( .A(n889), .B(n890), .Z(n887) );
  NANDN U779 ( .A(B[34]), .B(A[34]), .Z(n890) );
  AND U780 ( .A(n891), .B(n892), .Z(n889) );
  NAND U781 ( .A(n893), .B(n894), .Z(n892) );
  NANDN U782 ( .A(A[33]), .B(B[33]), .Z(n894) );
  AND U783 ( .A(n895), .B(n896), .Z(n893) );
  NANDN U784 ( .A(A[32]), .B(B[32]), .Z(n896) );
  NAND U785 ( .A(n897), .B(n898), .Z(n895) );
  NANDN U786 ( .A(B[32]), .B(A[32]), .Z(n898) );
  AND U787 ( .A(n899), .B(n900), .Z(n897) );
  NAND U788 ( .A(n901), .B(n902), .Z(n900) );
  NANDN U789 ( .A(A[31]), .B(B[31]), .Z(n902) );
  AND U790 ( .A(n903), .B(n904), .Z(n901) );
  NANDN U791 ( .A(A[30]), .B(B[30]), .Z(n904) );
  NAND U792 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U793 ( .A(B[30]), .B(A[30]), .Z(n906) );
  AND U794 ( .A(n907), .B(n908), .Z(n905) );
  NAND U795 ( .A(n909), .B(n910), .Z(n908) );
  NANDN U796 ( .A(A[29]), .B(B[29]), .Z(n910) );
  AND U797 ( .A(n911), .B(n912), .Z(n909) );
  NANDN U798 ( .A(A[28]), .B(B[28]), .Z(n912) );
  NAND U799 ( .A(n913), .B(n914), .Z(n911) );
  NANDN U800 ( .A(B[28]), .B(A[28]), .Z(n914) );
  AND U801 ( .A(n915), .B(n916), .Z(n913) );
  NAND U802 ( .A(n917), .B(n918), .Z(n916) );
  NANDN U803 ( .A(A[27]), .B(B[27]), .Z(n918) );
  AND U804 ( .A(n919), .B(n920), .Z(n917) );
  NANDN U805 ( .A(A[26]), .B(B[26]), .Z(n920) );
  NAND U806 ( .A(n921), .B(n922), .Z(n919) );
  NANDN U807 ( .A(B[26]), .B(A[26]), .Z(n922) );
  AND U808 ( .A(n923), .B(n924), .Z(n921) );
  NAND U809 ( .A(n925), .B(n926), .Z(n924) );
  NANDN U810 ( .A(A[25]), .B(B[25]), .Z(n926) );
  AND U811 ( .A(n927), .B(n928), .Z(n925) );
  NANDN U812 ( .A(A[24]), .B(B[24]), .Z(n928) );
  NAND U813 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U814 ( .A(B[24]), .B(A[24]), .Z(n930) );
  AND U815 ( .A(n931), .B(n932), .Z(n929) );
  NAND U816 ( .A(n933), .B(n934), .Z(n932) );
  NANDN U817 ( .A(A[23]), .B(B[23]), .Z(n934) );
  AND U818 ( .A(n935), .B(n936), .Z(n933) );
  NANDN U819 ( .A(A[22]), .B(B[22]), .Z(n936) );
  NAND U820 ( .A(n937), .B(n938), .Z(n935) );
  NANDN U821 ( .A(B[22]), .B(A[22]), .Z(n938) );
  AND U822 ( .A(n939), .B(n940), .Z(n937) );
  NAND U823 ( .A(n941), .B(n942), .Z(n940) );
  NANDN U824 ( .A(A[21]), .B(B[21]), .Z(n942) );
  AND U825 ( .A(n943), .B(n944), .Z(n941) );
  NANDN U826 ( .A(A[20]), .B(B[20]), .Z(n944) );
  NAND U827 ( .A(n945), .B(n946), .Z(n943) );
  NANDN U828 ( .A(B[20]), .B(A[20]), .Z(n946) );
  AND U829 ( .A(n947), .B(n948), .Z(n945) );
  NAND U830 ( .A(n949), .B(n950), .Z(n948) );
  NANDN U831 ( .A(A[19]), .B(B[19]), .Z(n950) );
  AND U832 ( .A(n951), .B(n952), .Z(n949) );
  NANDN U833 ( .A(A[18]), .B(B[18]), .Z(n952) );
  NAND U834 ( .A(n953), .B(n954), .Z(n951) );
  NANDN U835 ( .A(B[18]), .B(A[18]), .Z(n954) );
  AND U836 ( .A(n955), .B(n956), .Z(n953) );
  NAND U837 ( .A(n957), .B(n958), .Z(n956) );
  NANDN U838 ( .A(A[17]), .B(B[17]), .Z(n958) );
  AND U839 ( .A(n959), .B(n960), .Z(n957) );
  NANDN U840 ( .A(A[16]), .B(B[16]), .Z(n960) );
  NAND U841 ( .A(n961), .B(n962), .Z(n959) );
  NANDN U842 ( .A(B[16]), .B(A[16]), .Z(n962) );
  AND U843 ( .A(n963), .B(n964), .Z(n961) );
  NAND U844 ( .A(n965), .B(n966), .Z(n964) );
  NANDN U845 ( .A(A[15]), .B(B[15]), .Z(n966) );
  AND U846 ( .A(n967), .B(n968), .Z(n965) );
  NANDN U847 ( .A(A[14]), .B(B[14]), .Z(n968) );
  NAND U848 ( .A(n969), .B(n970), .Z(n967) );
  NANDN U849 ( .A(B[14]), .B(A[14]), .Z(n970) );
  AND U850 ( .A(n971), .B(n972), .Z(n969) );
  NAND U851 ( .A(n973), .B(n974), .Z(n972) );
  NANDN U852 ( .A(A[13]), .B(B[13]), .Z(n974) );
  AND U853 ( .A(n975), .B(n976), .Z(n973) );
  NANDN U854 ( .A(A[12]), .B(B[12]), .Z(n976) );
  NAND U855 ( .A(n977), .B(n978), .Z(n975) );
  NANDN U856 ( .A(B[12]), .B(A[12]), .Z(n978) );
  AND U857 ( .A(n979), .B(n980), .Z(n977) );
  NAND U858 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U859 ( .A(A[11]), .B(B[11]), .Z(n982) );
  AND U860 ( .A(n983), .B(n984), .Z(n981) );
  NANDN U861 ( .A(A[10]), .B(B[10]), .Z(n984) );
  NAND U862 ( .A(n985), .B(n986), .Z(n983) );
  NANDN U863 ( .A(B[9]), .B(A[9]), .Z(n986) );
  AND U864 ( .A(n987), .B(n988), .Z(n985) );
  NAND U865 ( .A(n989), .B(n990), .Z(n988) );
  NANDN U866 ( .A(A[9]), .B(B[9]), .Z(n990) );
  AND U867 ( .A(n991), .B(n992), .Z(n989) );
  NANDN U868 ( .A(A[8]), .B(B[8]), .Z(n992) );
  NAND U869 ( .A(n993), .B(n994), .Z(n991) );
  NANDN U870 ( .A(B[8]), .B(A[8]), .Z(n994) );
  AND U871 ( .A(n995), .B(n996), .Z(n993) );
  NAND U872 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U873 ( .A(A[7]), .B(B[7]), .Z(n998) );
  AND U874 ( .A(n999), .B(n1000), .Z(n997) );
  NANDN U875 ( .A(A[6]), .B(B[6]), .Z(n1000) );
  NAND U876 ( .A(n1001), .B(n1002), .Z(n999) );
  NANDN U877 ( .A(B[6]), .B(A[6]), .Z(n1002) );
  AND U878 ( .A(n1003), .B(n1004), .Z(n1001) );
  NAND U879 ( .A(n1005), .B(n1006), .Z(n1004) );
  NANDN U880 ( .A(A[5]), .B(B[5]), .Z(n1006) );
  AND U881 ( .A(n1007), .B(n1008), .Z(n1005) );
  NANDN U882 ( .A(A[4]), .B(B[4]), .Z(n1008) );
  NAND U883 ( .A(n1009), .B(n1010), .Z(n1007) );
  NANDN U884 ( .A(B[4]), .B(A[4]), .Z(n1010) );
  AND U885 ( .A(n1011), .B(n1012), .Z(n1009) );
  NAND U886 ( .A(n1013), .B(n1014), .Z(n1012) );
  NANDN U887 ( .A(A[3]), .B(B[3]), .Z(n1014) );
  AND U888 ( .A(n1015), .B(n1016), .Z(n1013) );
  NANDN U889 ( .A(A[2]), .B(B[2]), .Z(n1016) );
  NAND U890 ( .A(n1017), .B(n1018), .Z(n1015) );
  NANDN U891 ( .A(B[2]), .B(A[2]), .Z(n1018) );
  AND U892 ( .A(n1019), .B(n1020), .Z(n1017) );
  NAND U893 ( .A(n1021), .B(A[0]), .Z(n1020) );
  ANDN U894 ( .B(n1022), .A(B[0]), .Z(n1021) );
  NANDN U895 ( .A(A[1]), .B(B[1]), .Z(n1022) );
  NANDN U896 ( .A(B[1]), .B(A[1]), .Z(n1019) );
  NANDN U897 ( .A(B[3]), .B(A[3]), .Z(n1011) );
  NANDN U898 ( .A(B[5]), .B(A[5]), .Z(n1003) );
  NANDN U899 ( .A(B[7]), .B(A[7]), .Z(n995) );
  NANDN U900 ( .A(B[10]), .B(A[10]), .Z(n987) );
  NANDN U901 ( .A(B[11]), .B(A[11]), .Z(n979) );
  NANDN U902 ( .A(B[13]), .B(A[13]), .Z(n971) );
  NANDN U903 ( .A(B[15]), .B(A[15]), .Z(n963) );
  NANDN U904 ( .A(B[17]), .B(A[17]), .Z(n955) );
  NANDN U905 ( .A(B[19]), .B(A[19]), .Z(n947) );
  NANDN U906 ( .A(B[21]), .B(A[21]), .Z(n939) );
  NANDN U907 ( .A(B[23]), .B(A[23]), .Z(n931) );
  NANDN U908 ( .A(B[25]), .B(A[25]), .Z(n923) );
  NANDN U909 ( .A(B[27]), .B(A[27]), .Z(n915) );
  NANDN U910 ( .A(B[29]), .B(A[29]), .Z(n907) );
  NANDN U911 ( .A(B[31]), .B(A[31]), .Z(n899) );
  NANDN U912 ( .A(B[33]), .B(A[33]), .Z(n891) );
  NANDN U913 ( .A(B[35]), .B(A[35]), .Z(n883) );
  NANDN U914 ( .A(B[37]), .B(A[37]), .Z(n875) );
  NANDN U915 ( .A(B[39]), .B(A[39]), .Z(n867) );
  NANDN U916 ( .A(B[41]), .B(A[41]), .Z(n859) );
  NANDN U917 ( .A(B[43]), .B(A[43]), .Z(n851) );
  NANDN U918 ( .A(B[45]), .B(A[45]), .Z(n843) );
  NANDN U919 ( .A(B[47]), .B(A[47]), .Z(n835) );
  NANDN U920 ( .A(B[49]), .B(A[49]), .Z(n827) );
  NANDN U921 ( .A(B[51]), .B(A[51]), .Z(n819) );
  NANDN U922 ( .A(B[53]), .B(A[53]), .Z(n811) );
  NANDN U923 ( .A(B[55]), .B(A[55]), .Z(n803) );
  NANDN U924 ( .A(B[57]), .B(A[57]), .Z(n795) );
  NANDN U925 ( .A(B[59]), .B(A[59]), .Z(n787) );
  NANDN U926 ( .A(B[61]), .B(A[61]), .Z(n779) );
  NANDN U927 ( .A(B[63]), .B(A[63]), .Z(n771) );
  NANDN U928 ( .A(B[65]), .B(A[65]), .Z(n763) );
  NANDN U929 ( .A(B[67]), .B(A[67]), .Z(n755) );
  NANDN U930 ( .A(B[69]), .B(A[69]), .Z(n747) );
  NANDN U931 ( .A(B[71]), .B(A[71]), .Z(n739) );
  NANDN U932 ( .A(B[73]), .B(A[73]), .Z(n731) );
  NANDN U933 ( .A(B[75]), .B(A[75]), .Z(n723) );
  NANDN U934 ( .A(B[77]), .B(A[77]), .Z(n715) );
  NANDN U935 ( .A(B[79]), .B(A[79]), .Z(n707) );
  NANDN U936 ( .A(B[81]), .B(A[81]), .Z(n699) );
  NANDN U937 ( .A(B[83]), .B(A[83]), .Z(n691) );
  NANDN U938 ( .A(B[85]), .B(A[85]), .Z(n683) );
  NANDN U939 ( .A(B[87]), .B(A[87]), .Z(n675) );
  NANDN U940 ( .A(B[89]), .B(A[89]), .Z(n667) );
  NANDN U941 ( .A(B[91]), .B(A[91]), .Z(n659) );
  NANDN U942 ( .A(B[93]), .B(A[93]), .Z(n651) );
  NANDN U943 ( .A(B[95]), .B(A[95]), .Z(n643) );
  NANDN U944 ( .A(B[97]), .B(A[97]), .Z(n635) );
  NANDN U945 ( .A(B[100]), .B(A[100]), .Z(n627) );
  NANDN U946 ( .A(B[101]), .B(A[101]), .Z(n619) );
  NANDN U947 ( .A(B[103]), .B(A[103]), .Z(n611) );
  NANDN U948 ( .A(B[105]), .B(A[105]), .Z(n603) );
  NANDN U949 ( .A(B[107]), .B(A[107]), .Z(n595) );
  NANDN U950 ( .A(B[109]), .B(A[109]), .Z(n587) );
  NANDN U951 ( .A(B[111]), .B(A[111]), .Z(n579) );
  NANDN U952 ( .A(B[113]), .B(A[113]), .Z(n571) );
  NANDN U953 ( .A(B[115]), .B(A[115]), .Z(n563) );
  NANDN U954 ( .A(B[117]), .B(A[117]), .Z(n555) );
  NANDN U955 ( .A(B[119]), .B(A[119]), .Z(n547) );
  NANDN U956 ( .A(B[121]), .B(A[121]), .Z(n539) );
  NANDN U957 ( .A(B[123]), .B(A[123]), .Z(n531) );
  NANDN U958 ( .A(B[125]), .B(A[125]), .Z(n523) );
  NANDN U959 ( .A(B[127]), .B(A[127]), .Z(n515) );
  NANDN U960 ( .A(B[129]), .B(A[129]), .Z(n507) );
  NANDN U961 ( .A(B[131]), .B(A[131]), .Z(n499) );
  NANDN U962 ( .A(B[133]), .B(A[133]), .Z(n491) );
  NANDN U963 ( .A(B[135]), .B(A[135]), .Z(n483) );
  NANDN U964 ( .A(B[137]), .B(A[137]), .Z(n475) );
  NANDN U965 ( .A(B[139]), .B(A[139]), .Z(n467) );
  NANDN U966 ( .A(B[141]), .B(A[141]), .Z(n459) );
  NANDN U967 ( .A(B[143]), .B(A[143]), .Z(n451) );
  NANDN U968 ( .A(B[145]), .B(A[145]), .Z(n443) );
  NANDN U969 ( .A(B[147]), .B(A[147]), .Z(n435) );
  NANDN U970 ( .A(B[149]), .B(A[149]), .Z(n427) );
  NANDN U971 ( .A(B[151]), .B(A[151]), .Z(n419) );
  NANDN U972 ( .A(B[153]), .B(A[153]), .Z(n411) );
  NANDN U973 ( .A(B[155]), .B(A[155]), .Z(n403) );
  NANDN U974 ( .A(B[157]), .B(A[157]), .Z(n395) );
  NANDN U975 ( .A(B[159]), .B(A[159]), .Z(n387) );
  NANDN U976 ( .A(B[161]), .B(A[161]), .Z(n379) );
  NANDN U977 ( .A(B[163]), .B(A[163]), .Z(n371) );
  NANDN U978 ( .A(B[165]), .B(A[165]), .Z(n363) );
  NANDN U979 ( .A(B[167]), .B(A[167]), .Z(n355) );
  NANDN U980 ( .A(B[169]), .B(A[169]), .Z(n347) );
  NANDN U981 ( .A(B[171]), .B(A[171]), .Z(n339) );
  NANDN U982 ( .A(B[173]), .B(A[173]), .Z(n331) );
  NANDN U983 ( .A(B[175]), .B(A[175]), .Z(n323) );
  NANDN U984 ( .A(B[177]), .B(A[177]), .Z(n315) );
  NANDN U985 ( .A(B[179]), .B(A[179]), .Z(n307) );
  NANDN U986 ( .A(B[181]), .B(A[181]), .Z(n299) );
  NANDN U987 ( .A(B[183]), .B(A[183]), .Z(n291) );
  NANDN U988 ( .A(B[185]), .B(A[185]), .Z(n283) );
  NANDN U989 ( .A(B[187]), .B(A[187]), .Z(n275) );
  NANDN U990 ( .A(B[189]), .B(A[189]), .Z(n267) );
  NANDN U991 ( .A(B[191]), .B(A[191]), .Z(n259) );
  NANDN U992 ( .A(B[193]), .B(A[193]), .Z(n251) );
  NANDN U993 ( .A(B[195]), .B(A[195]), .Z(n243) );
  NANDN U994 ( .A(B[197]), .B(A[197]), .Z(n235) );
  NANDN U995 ( .A(B[199]), .B(A[199]), .Z(n227) );
  NANDN U996 ( .A(B[201]), .B(A[201]), .Z(n219) );
  NANDN U997 ( .A(B[203]), .B(A[203]), .Z(n211) );
  NANDN U998 ( .A(B[205]), .B(A[205]), .Z(n203) );
  NANDN U999 ( .A(B[207]), .B(A[207]), .Z(n195) );
  NANDN U1000 ( .A(B[209]), .B(A[209]), .Z(n187) );
  NANDN U1001 ( .A(B[211]), .B(A[211]), .Z(n179) );
  NANDN U1002 ( .A(B[213]), .B(A[213]), .Z(n171) );
  NANDN U1003 ( .A(B[215]), .B(A[215]), .Z(n163) );
  NANDN U1004 ( .A(B[217]), .B(A[217]), .Z(n155) );
  NANDN U1005 ( .A(B[219]), .B(A[219]), .Z(n147) );
  NANDN U1006 ( .A(B[221]), .B(A[221]), .Z(n139) );
  NANDN U1007 ( .A(B[223]), .B(A[223]), .Z(n131) );
  NANDN U1008 ( .A(B[225]), .B(A[225]), .Z(n123) );
  NANDN U1009 ( .A(B[227]), .B(A[227]), .Z(n115) );
  NANDN U1010 ( .A(B[229]), .B(A[229]), .Z(n107) );
  NANDN U1011 ( .A(B[231]), .B(A[231]), .Z(n99) );
  NANDN U1012 ( .A(B[233]), .B(A[233]), .Z(n91) );
  NANDN U1013 ( .A(B[235]), .B(A[235]), .Z(n83) );
  NANDN U1014 ( .A(B[237]), .B(A[237]), .Z(n75) );
  NANDN U1015 ( .A(B[239]), .B(A[239]), .Z(n67) );
  NANDN U1016 ( .A(B[241]), .B(A[241]), .Z(n59) );
  NANDN U1017 ( .A(B[243]), .B(A[243]), .Z(n51) );
  NANDN U1018 ( .A(B[245]), .B(A[245]), .Z(n43) );
  NANDN U1019 ( .A(B[247]), .B(A[247]), .Z(n35) );
  NANDN U1020 ( .A(B[249]), .B(A[249]), .Z(n27) );
  NANDN U1021 ( .A(B[251]), .B(A[251]), .Z(n19) );
  NANDN U1022 ( .A(B[253]), .B(A[253]), .Z(n11) );
  NANDN U1023 ( .A(A[255]), .B(B[255]), .Z(n3) );
endmodule


module modmult_step_N256_5_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280;

  IV U1 ( .A(A[1]), .Z(n1) );
  IV U2 ( .A(n1279), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(DIFF[9]) );
  XOR U4 ( .A(B[9]), .B(A[9]), .Z(n4) );
  XNOR U5 ( .A(n5), .B(n6), .Z(DIFF[99]) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(DIFF[98]) );
  XOR U8 ( .A(B[98]), .B(A[98]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(DIFF[97]) );
  XOR U10 ( .A(B[97]), .B(A[97]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(DIFF[96]) );
  XOR U12 ( .A(B[96]), .B(A[96]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(DIFF[95]) );
  XOR U14 ( .A(B[95]), .B(A[95]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(DIFF[94]) );
  XOR U16 ( .A(B[94]), .B(A[94]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(DIFF[93]) );
  XOR U18 ( .A(B[93]), .B(A[93]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(DIFF[92]) );
  XOR U20 ( .A(B[92]), .B(A[92]), .Z(n20) );
  XOR U21 ( .A(n21), .B(n22), .Z(DIFF[91]) );
  XOR U22 ( .A(B[91]), .B(A[91]), .Z(n22) );
  XOR U23 ( .A(n23), .B(n24), .Z(DIFF[90]) );
  XOR U24 ( .A(B[90]), .B(A[90]), .Z(n24) );
  XOR U25 ( .A(n25), .B(n26), .Z(DIFF[8]) );
  XOR U26 ( .A(B[8]), .B(A[8]), .Z(n26) );
  XOR U27 ( .A(n27), .B(n28), .Z(DIFF[89]) );
  XOR U28 ( .A(B[89]), .B(A[89]), .Z(n28) );
  XOR U29 ( .A(n29), .B(n30), .Z(DIFF[88]) );
  XOR U30 ( .A(B[88]), .B(A[88]), .Z(n30) );
  XOR U31 ( .A(n31), .B(n32), .Z(DIFF[87]) );
  XOR U32 ( .A(B[87]), .B(A[87]), .Z(n32) );
  XOR U33 ( .A(n33), .B(n34), .Z(DIFF[86]) );
  XOR U34 ( .A(B[86]), .B(A[86]), .Z(n34) );
  XOR U35 ( .A(n35), .B(n36), .Z(DIFF[85]) );
  XOR U36 ( .A(B[85]), .B(A[85]), .Z(n36) );
  XOR U37 ( .A(n37), .B(n38), .Z(DIFF[84]) );
  XOR U38 ( .A(B[84]), .B(A[84]), .Z(n38) );
  XOR U39 ( .A(n39), .B(n40), .Z(DIFF[83]) );
  XOR U40 ( .A(B[83]), .B(A[83]), .Z(n40) );
  XOR U41 ( .A(n41), .B(n42), .Z(DIFF[82]) );
  XOR U42 ( .A(B[82]), .B(A[82]), .Z(n42) );
  XOR U43 ( .A(n43), .B(n44), .Z(DIFF[81]) );
  XOR U44 ( .A(B[81]), .B(A[81]), .Z(n44) );
  XOR U45 ( .A(n45), .B(n46), .Z(DIFF[80]) );
  XOR U46 ( .A(B[80]), .B(A[80]), .Z(n46) );
  XOR U47 ( .A(n47), .B(n48), .Z(DIFF[7]) );
  XOR U48 ( .A(B[7]), .B(A[7]), .Z(n48) );
  XOR U49 ( .A(n49), .B(n50), .Z(DIFF[79]) );
  XOR U50 ( .A(B[79]), .B(A[79]), .Z(n50) );
  XOR U51 ( .A(n51), .B(n52), .Z(DIFF[78]) );
  XOR U52 ( .A(B[78]), .B(A[78]), .Z(n52) );
  XOR U53 ( .A(n53), .B(n54), .Z(DIFF[77]) );
  XOR U54 ( .A(B[77]), .B(A[77]), .Z(n54) );
  XOR U55 ( .A(n55), .B(n56), .Z(DIFF[76]) );
  XOR U56 ( .A(B[76]), .B(A[76]), .Z(n56) );
  XOR U57 ( .A(n57), .B(n58), .Z(DIFF[75]) );
  XOR U58 ( .A(B[75]), .B(A[75]), .Z(n58) );
  XOR U59 ( .A(n59), .B(n60), .Z(DIFF[74]) );
  XOR U60 ( .A(B[74]), .B(A[74]), .Z(n60) );
  XOR U61 ( .A(n61), .B(n62), .Z(DIFF[73]) );
  XOR U62 ( .A(B[73]), .B(A[73]), .Z(n62) );
  XOR U63 ( .A(n63), .B(n64), .Z(DIFF[72]) );
  XOR U64 ( .A(B[72]), .B(A[72]), .Z(n64) );
  XOR U65 ( .A(n65), .B(n66), .Z(DIFF[71]) );
  XOR U66 ( .A(B[71]), .B(A[71]), .Z(n66) );
  XOR U67 ( .A(n67), .B(n68), .Z(DIFF[70]) );
  XOR U68 ( .A(B[70]), .B(A[70]), .Z(n68) );
  XOR U69 ( .A(n69), .B(n70), .Z(DIFF[6]) );
  XOR U70 ( .A(B[6]), .B(A[6]), .Z(n70) );
  XOR U71 ( .A(n71), .B(n72), .Z(DIFF[69]) );
  XOR U72 ( .A(B[69]), .B(A[69]), .Z(n72) );
  XOR U73 ( .A(n73), .B(n74), .Z(DIFF[68]) );
  XOR U74 ( .A(B[68]), .B(A[68]), .Z(n74) );
  XOR U75 ( .A(n75), .B(n76), .Z(DIFF[67]) );
  XOR U76 ( .A(B[67]), .B(A[67]), .Z(n76) );
  XOR U77 ( .A(n77), .B(n78), .Z(DIFF[66]) );
  XOR U78 ( .A(B[66]), .B(A[66]), .Z(n78) );
  XOR U79 ( .A(n79), .B(n80), .Z(DIFF[65]) );
  XOR U80 ( .A(B[65]), .B(A[65]), .Z(n80) );
  XOR U81 ( .A(n81), .B(n82), .Z(DIFF[64]) );
  XOR U82 ( .A(B[64]), .B(A[64]), .Z(n82) );
  XOR U83 ( .A(n83), .B(n84), .Z(DIFF[63]) );
  XOR U84 ( .A(B[63]), .B(A[63]), .Z(n84) );
  XOR U85 ( .A(n85), .B(n86), .Z(DIFF[62]) );
  XOR U86 ( .A(B[62]), .B(A[62]), .Z(n86) );
  XOR U87 ( .A(n87), .B(n88), .Z(DIFF[61]) );
  XOR U88 ( .A(B[61]), .B(A[61]), .Z(n88) );
  XOR U89 ( .A(n89), .B(n90), .Z(DIFF[60]) );
  XOR U90 ( .A(B[60]), .B(A[60]), .Z(n90) );
  XOR U91 ( .A(n91), .B(n92), .Z(DIFF[5]) );
  XOR U92 ( .A(B[5]), .B(A[5]), .Z(n92) );
  XOR U93 ( .A(n93), .B(n94), .Z(DIFF[59]) );
  XOR U94 ( .A(B[59]), .B(A[59]), .Z(n94) );
  XOR U95 ( .A(n95), .B(n96), .Z(DIFF[58]) );
  XOR U96 ( .A(B[58]), .B(A[58]), .Z(n96) );
  XOR U97 ( .A(n97), .B(n98), .Z(DIFF[57]) );
  XOR U98 ( .A(B[57]), .B(A[57]), .Z(n98) );
  XOR U99 ( .A(n99), .B(n100), .Z(DIFF[56]) );
  XOR U100 ( .A(B[56]), .B(A[56]), .Z(n100) );
  XOR U101 ( .A(n101), .B(n102), .Z(DIFF[55]) );
  XOR U102 ( .A(B[55]), .B(A[55]), .Z(n102) );
  XOR U103 ( .A(n103), .B(n104), .Z(DIFF[54]) );
  XOR U104 ( .A(B[54]), .B(A[54]), .Z(n104) );
  XOR U105 ( .A(n105), .B(n106), .Z(DIFF[53]) );
  XOR U106 ( .A(B[53]), .B(A[53]), .Z(n106) );
  XOR U107 ( .A(n107), .B(n108), .Z(DIFF[52]) );
  XOR U108 ( .A(B[52]), .B(A[52]), .Z(n108) );
  XOR U109 ( .A(n109), .B(n110), .Z(DIFF[51]) );
  XOR U110 ( .A(B[51]), .B(A[51]), .Z(n110) );
  XOR U111 ( .A(n111), .B(n112), .Z(DIFF[50]) );
  XOR U112 ( .A(B[50]), .B(A[50]), .Z(n112) );
  XOR U113 ( .A(n113), .B(n114), .Z(DIFF[4]) );
  XOR U114 ( .A(B[4]), .B(A[4]), .Z(n114) );
  XOR U115 ( .A(n115), .B(n116), .Z(DIFF[49]) );
  XOR U116 ( .A(B[49]), .B(A[49]), .Z(n116) );
  XOR U117 ( .A(n117), .B(n118), .Z(DIFF[48]) );
  XOR U118 ( .A(B[48]), .B(A[48]), .Z(n118) );
  XOR U119 ( .A(n119), .B(n120), .Z(DIFF[47]) );
  XOR U120 ( .A(B[47]), .B(A[47]), .Z(n120) );
  XOR U121 ( .A(n121), .B(n122), .Z(DIFF[46]) );
  XOR U122 ( .A(B[46]), .B(A[46]), .Z(n122) );
  XOR U123 ( .A(n123), .B(n124), .Z(DIFF[45]) );
  XOR U124 ( .A(B[45]), .B(A[45]), .Z(n124) );
  XOR U125 ( .A(n125), .B(n126), .Z(DIFF[44]) );
  XOR U126 ( .A(B[44]), .B(A[44]), .Z(n126) );
  XOR U127 ( .A(n127), .B(n128), .Z(DIFF[43]) );
  XOR U128 ( .A(B[43]), .B(A[43]), .Z(n128) );
  XOR U129 ( .A(n129), .B(n130), .Z(DIFF[42]) );
  XOR U130 ( .A(B[42]), .B(A[42]), .Z(n130) );
  XOR U131 ( .A(n131), .B(n132), .Z(DIFF[41]) );
  XOR U132 ( .A(B[41]), .B(A[41]), .Z(n132) );
  XOR U133 ( .A(n133), .B(n134), .Z(DIFF[40]) );
  XOR U134 ( .A(B[40]), .B(A[40]), .Z(n134) );
  XOR U135 ( .A(n135), .B(n136), .Z(DIFF[3]) );
  XOR U136 ( .A(B[3]), .B(A[3]), .Z(n136) );
  XOR U137 ( .A(n137), .B(n138), .Z(DIFF[39]) );
  XOR U138 ( .A(B[39]), .B(A[39]), .Z(n138) );
  XOR U139 ( .A(n139), .B(n140), .Z(DIFF[38]) );
  XOR U140 ( .A(B[38]), .B(A[38]), .Z(n140) );
  XOR U141 ( .A(n141), .B(n142), .Z(DIFF[37]) );
  XOR U142 ( .A(B[37]), .B(A[37]), .Z(n142) );
  XOR U143 ( .A(n143), .B(n144), .Z(DIFF[36]) );
  XOR U144 ( .A(B[36]), .B(A[36]), .Z(n144) );
  XOR U145 ( .A(n145), .B(n146), .Z(DIFF[35]) );
  XOR U146 ( .A(B[35]), .B(A[35]), .Z(n146) );
  XOR U147 ( .A(n147), .B(n148), .Z(DIFF[34]) );
  XOR U148 ( .A(B[34]), .B(A[34]), .Z(n148) );
  XOR U149 ( .A(n149), .B(n150), .Z(DIFF[33]) );
  XOR U150 ( .A(B[33]), .B(A[33]), .Z(n150) );
  XOR U151 ( .A(n151), .B(n152), .Z(DIFF[32]) );
  XOR U152 ( .A(B[32]), .B(A[32]), .Z(n152) );
  XOR U153 ( .A(n153), .B(n154), .Z(DIFF[31]) );
  XOR U154 ( .A(B[31]), .B(A[31]), .Z(n154) );
  XOR U155 ( .A(n155), .B(n156), .Z(DIFF[30]) );
  XOR U156 ( .A(B[30]), .B(A[30]), .Z(n156) );
  XOR U157 ( .A(n157), .B(n158), .Z(DIFF[2]) );
  XOR U158 ( .A(B[2]), .B(A[2]), .Z(n158) );
  XOR U159 ( .A(n159), .B(n160), .Z(DIFF[29]) );
  XOR U160 ( .A(B[29]), .B(A[29]), .Z(n160) );
  XOR U161 ( .A(n161), .B(n162), .Z(DIFF[28]) );
  XOR U162 ( .A(B[28]), .B(A[28]), .Z(n162) );
  XOR U163 ( .A(n163), .B(n164), .Z(DIFF[27]) );
  XOR U164 ( .A(B[27]), .B(A[27]), .Z(n164) );
  XOR U165 ( .A(n165), .B(n166), .Z(DIFF[26]) );
  XOR U166 ( .A(B[26]), .B(A[26]), .Z(n166) );
  XOR U167 ( .A(n167), .B(n168), .Z(DIFF[25]) );
  XOR U168 ( .A(B[25]), .B(A[25]), .Z(n168) );
  XOR U169 ( .A(A[257]), .B(n169), .Z(DIFF[257]) );
  ANDN U170 ( .B(n170), .A(A[256]), .Z(n169) );
  XOR U171 ( .A(A[256]), .B(n170), .Z(DIFF[256]) );
  AND U172 ( .A(n171), .B(n172), .Z(n170) );
  NANDN U173 ( .A(B[255]), .B(n173), .Z(n172) );
  NANDN U174 ( .A(A[255]), .B(n174), .Z(n173) );
  NANDN U175 ( .A(n174), .B(A[255]), .Z(n171) );
  XOR U176 ( .A(n174), .B(n175), .Z(DIFF[255]) );
  XOR U177 ( .A(B[255]), .B(A[255]), .Z(n175) );
  AND U178 ( .A(n176), .B(n177), .Z(n174) );
  NANDN U179 ( .A(B[254]), .B(n178), .Z(n177) );
  NANDN U180 ( .A(A[254]), .B(n179), .Z(n178) );
  NANDN U181 ( .A(n179), .B(A[254]), .Z(n176) );
  XOR U182 ( .A(n179), .B(n180), .Z(DIFF[254]) );
  XOR U183 ( .A(B[254]), .B(A[254]), .Z(n180) );
  AND U184 ( .A(n181), .B(n182), .Z(n179) );
  NANDN U185 ( .A(B[253]), .B(n183), .Z(n182) );
  NANDN U186 ( .A(A[253]), .B(n184), .Z(n183) );
  NANDN U187 ( .A(n184), .B(A[253]), .Z(n181) );
  XOR U188 ( .A(n184), .B(n185), .Z(DIFF[253]) );
  XOR U189 ( .A(B[253]), .B(A[253]), .Z(n185) );
  AND U190 ( .A(n186), .B(n187), .Z(n184) );
  NANDN U191 ( .A(B[252]), .B(n188), .Z(n187) );
  NANDN U192 ( .A(A[252]), .B(n189), .Z(n188) );
  NANDN U193 ( .A(n189), .B(A[252]), .Z(n186) );
  XOR U194 ( .A(n189), .B(n190), .Z(DIFF[252]) );
  XOR U195 ( .A(B[252]), .B(A[252]), .Z(n190) );
  AND U196 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U197 ( .A(B[251]), .B(n193), .Z(n192) );
  NANDN U198 ( .A(A[251]), .B(n194), .Z(n193) );
  NANDN U199 ( .A(n194), .B(A[251]), .Z(n191) );
  XOR U200 ( .A(n194), .B(n195), .Z(DIFF[251]) );
  XOR U201 ( .A(B[251]), .B(A[251]), .Z(n195) );
  AND U202 ( .A(n196), .B(n197), .Z(n194) );
  NANDN U203 ( .A(B[250]), .B(n198), .Z(n197) );
  NANDN U204 ( .A(A[250]), .B(n199), .Z(n198) );
  NANDN U205 ( .A(n199), .B(A[250]), .Z(n196) );
  XOR U206 ( .A(n199), .B(n200), .Z(DIFF[250]) );
  XOR U207 ( .A(B[250]), .B(A[250]), .Z(n200) );
  AND U208 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U209 ( .A(B[249]), .B(n203), .Z(n202) );
  NANDN U210 ( .A(A[249]), .B(n204), .Z(n203) );
  NANDN U211 ( .A(n204), .B(A[249]), .Z(n201) );
  XOR U212 ( .A(n205), .B(n206), .Z(DIFF[24]) );
  XOR U213 ( .A(B[24]), .B(A[24]), .Z(n206) );
  XOR U214 ( .A(n204), .B(n207), .Z(DIFF[249]) );
  XOR U215 ( .A(B[249]), .B(A[249]), .Z(n207) );
  AND U216 ( .A(n208), .B(n209), .Z(n204) );
  NANDN U217 ( .A(B[248]), .B(n210), .Z(n209) );
  NANDN U218 ( .A(A[248]), .B(n211), .Z(n210) );
  NANDN U219 ( .A(n211), .B(A[248]), .Z(n208) );
  XOR U220 ( .A(n211), .B(n212), .Z(DIFF[248]) );
  XOR U221 ( .A(B[248]), .B(A[248]), .Z(n212) );
  AND U222 ( .A(n213), .B(n214), .Z(n211) );
  NANDN U223 ( .A(B[247]), .B(n215), .Z(n214) );
  NANDN U224 ( .A(A[247]), .B(n216), .Z(n215) );
  NANDN U225 ( .A(n216), .B(A[247]), .Z(n213) );
  XOR U226 ( .A(n216), .B(n217), .Z(DIFF[247]) );
  XOR U227 ( .A(B[247]), .B(A[247]), .Z(n217) );
  AND U228 ( .A(n218), .B(n219), .Z(n216) );
  NANDN U229 ( .A(B[246]), .B(n220), .Z(n219) );
  NANDN U230 ( .A(A[246]), .B(n221), .Z(n220) );
  NANDN U231 ( .A(n221), .B(A[246]), .Z(n218) );
  XOR U232 ( .A(n221), .B(n222), .Z(DIFF[246]) );
  XOR U233 ( .A(B[246]), .B(A[246]), .Z(n222) );
  AND U234 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U235 ( .A(B[245]), .B(n225), .Z(n224) );
  NANDN U236 ( .A(A[245]), .B(n226), .Z(n225) );
  NANDN U237 ( .A(n226), .B(A[245]), .Z(n223) );
  XOR U238 ( .A(n226), .B(n227), .Z(DIFF[245]) );
  XOR U239 ( .A(B[245]), .B(A[245]), .Z(n227) );
  AND U240 ( .A(n228), .B(n229), .Z(n226) );
  NANDN U241 ( .A(B[244]), .B(n230), .Z(n229) );
  NANDN U242 ( .A(A[244]), .B(n231), .Z(n230) );
  NANDN U243 ( .A(n231), .B(A[244]), .Z(n228) );
  XOR U244 ( .A(n231), .B(n232), .Z(DIFF[244]) );
  XOR U245 ( .A(B[244]), .B(A[244]), .Z(n232) );
  AND U246 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U247 ( .A(B[243]), .B(n235), .Z(n234) );
  NANDN U248 ( .A(A[243]), .B(n236), .Z(n235) );
  NANDN U249 ( .A(n236), .B(A[243]), .Z(n233) );
  XOR U250 ( .A(n236), .B(n237), .Z(DIFF[243]) );
  XOR U251 ( .A(B[243]), .B(A[243]), .Z(n237) );
  AND U252 ( .A(n238), .B(n239), .Z(n236) );
  NANDN U253 ( .A(B[242]), .B(n240), .Z(n239) );
  NANDN U254 ( .A(A[242]), .B(n241), .Z(n240) );
  NANDN U255 ( .A(n241), .B(A[242]), .Z(n238) );
  XOR U256 ( .A(n241), .B(n242), .Z(DIFF[242]) );
  XOR U257 ( .A(B[242]), .B(A[242]), .Z(n242) );
  AND U258 ( .A(n243), .B(n244), .Z(n241) );
  NANDN U259 ( .A(B[241]), .B(n245), .Z(n244) );
  NANDN U260 ( .A(A[241]), .B(n246), .Z(n245) );
  NANDN U261 ( .A(n246), .B(A[241]), .Z(n243) );
  XOR U262 ( .A(n246), .B(n247), .Z(DIFF[241]) );
  XOR U263 ( .A(B[241]), .B(A[241]), .Z(n247) );
  AND U264 ( .A(n248), .B(n249), .Z(n246) );
  NANDN U265 ( .A(B[240]), .B(n250), .Z(n249) );
  NANDN U266 ( .A(A[240]), .B(n251), .Z(n250) );
  NANDN U267 ( .A(n251), .B(A[240]), .Z(n248) );
  XOR U268 ( .A(n251), .B(n252), .Z(DIFF[240]) );
  XOR U269 ( .A(B[240]), .B(A[240]), .Z(n252) );
  AND U270 ( .A(n253), .B(n254), .Z(n251) );
  NANDN U271 ( .A(B[239]), .B(n255), .Z(n254) );
  NANDN U272 ( .A(A[239]), .B(n256), .Z(n255) );
  NANDN U273 ( .A(n256), .B(A[239]), .Z(n253) );
  XOR U274 ( .A(n257), .B(n258), .Z(DIFF[23]) );
  XOR U275 ( .A(B[23]), .B(A[23]), .Z(n258) );
  XOR U276 ( .A(n256), .B(n259), .Z(DIFF[239]) );
  XOR U277 ( .A(B[239]), .B(A[239]), .Z(n259) );
  AND U278 ( .A(n260), .B(n261), .Z(n256) );
  NANDN U279 ( .A(B[238]), .B(n262), .Z(n261) );
  NANDN U280 ( .A(A[238]), .B(n263), .Z(n262) );
  NANDN U281 ( .A(n263), .B(A[238]), .Z(n260) );
  XOR U282 ( .A(n263), .B(n264), .Z(DIFF[238]) );
  XOR U283 ( .A(B[238]), .B(A[238]), .Z(n264) );
  AND U284 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U285 ( .A(B[237]), .B(n267), .Z(n266) );
  NANDN U286 ( .A(A[237]), .B(n268), .Z(n267) );
  NANDN U287 ( .A(n268), .B(A[237]), .Z(n265) );
  XOR U288 ( .A(n268), .B(n269), .Z(DIFF[237]) );
  XOR U289 ( .A(B[237]), .B(A[237]), .Z(n269) );
  AND U290 ( .A(n270), .B(n271), .Z(n268) );
  NANDN U291 ( .A(B[236]), .B(n272), .Z(n271) );
  NANDN U292 ( .A(A[236]), .B(n273), .Z(n272) );
  NANDN U293 ( .A(n273), .B(A[236]), .Z(n270) );
  XOR U294 ( .A(n273), .B(n274), .Z(DIFF[236]) );
  XOR U295 ( .A(B[236]), .B(A[236]), .Z(n274) );
  AND U296 ( .A(n275), .B(n276), .Z(n273) );
  NANDN U297 ( .A(B[235]), .B(n277), .Z(n276) );
  NANDN U298 ( .A(A[235]), .B(n278), .Z(n277) );
  NANDN U299 ( .A(n278), .B(A[235]), .Z(n275) );
  XOR U300 ( .A(n278), .B(n279), .Z(DIFF[235]) );
  XOR U301 ( .A(B[235]), .B(A[235]), .Z(n279) );
  AND U302 ( .A(n280), .B(n281), .Z(n278) );
  NANDN U303 ( .A(B[234]), .B(n282), .Z(n281) );
  NANDN U304 ( .A(A[234]), .B(n283), .Z(n282) );
  NANDN U305 ( .A(n283), .B(A[234]), .Z(n280) );
  XOR U306 ( .A(n283), .B(n284), .Z(DIFF[234]) );
  XOR U307 ( .A(B[234]), .B(A[234]), .Z(n284) );
  AND U308 ( .A(n285), .B(n286), .Z(n283) );
  NANDN U309 ( .A(B[233]), .B(n287), .Z(n286) );
  NANDN U310 ( .A(A[233]), .B(n288), .Z(n287) );
  NANDN U311 ( .A(n288), .B(A[233]), .Z(n285) );
  XOR U312 ( .A(n288), .B(n289), .Z(DIFF[233]) );
  XOR U313 ( .A(B[233]), .B(A[233]), .Z(n289) );
  AND U314 ( .A(n290), .B(n291), .Z(n288) );
  NANDN U315 ( .A(B[232]), .B(n292), .Z(n291) );
  NANDN U316 ( .A(A[232]), .B(n293), .Z(n292) );
  NANDN U317 ( .A(n293), .B(A[232]), .Z(n290) );
  XOR U318 ( .A(n293), .B(n294), .Z(DIFF[232]) );
  XOR U319 ( .A(B[232]), .B(A[232]), .Z(n294) );
  AND U320 ( .A(n295), .B(n296), .Z(n293) );
  NANDN U321 ( .A(B[231]), .B(n297), .Z(n296) );
  NANDN U322 ( .A(A[231]), .B(n298), .Z(n297) );
  NANDN U323 ( .A(n298), .B(A[231]), .Z(n295) );
  XOR U324 ( .A(n298), .B(n299), .Z(DIFF[231]) );
  XOR U325 ( .A(B[231]), .B(A[231]), .Z(n299) );
  AND U326 ( .A(n300), .B(n301), .Z(n298) );
  NANDN U327 ( .A(B[230]), .B(n302), .Z(n301) );
  NANDN U328 ( .A(A[230]), .B(n303), .Z(n302) );
  NANDN U329 ( .A(n303), .B(A[230]), .Z(n300) );
  XOR U330 ( .A(n303), .B(n304), .Z(DIFF[230]) );
  XOR U331 ( .A(B[230]), .B(A[230]), .Z(n304) );
  AND U332 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U333 ( .A(B[229]), .B(n307), .Z(n306) );
  NANDN U334 ( .A(A[229]), .B(n308), .Z(n307) );
  NANDN U335 ( .A(n308), .B(A[229]), .Z(n305) );
  XOR U336 ( .A(n309), .B(n310), .Z(DIFF[22]) );
  XOR U337 ( .A(B[22]), .B(A[22]), .Z(n310) );
  XOR U338 ( .A(n308), .B(n311), .Z(DIFF[229]) );
  XOR U339 ( .A(B[229]), .B(A[229]), .Z(n311) );
  AND U340 ( .A(n312), .B(n313), .Z(n308) );
  NANDN U341 ( .A(B[228]), .B(n314), .Z(n313) );
  NANDN U342 ( .A(A[228]), .B(n315), .Z(n314) );
  NANDN U343 ( .A(n315), .B(A[228]), .Z(n312) );
  XOR U344 ( .A(n315), .B(n316), .Z(DIFF[228]) );
  XOR U345 ( .A(B[228]), .B(A[228]), .Z(n316) );
  AND U346 ( .A(n317), .B(n318), .Z(n315) );
  NANDN U347 ( .A(B[227]), .B(n319), .Z(n318) );
  NANDN U348 ( .A(A[227]), .B(n320), .Z(n319) );
  NANDN U349 ( .A(n320), .B(A[227]), .Z(n317) );
  XOR U350 ( .A(n320), .B(n321), .Z(DIFF[227]) );
  XOR U351 ( .A(B[227]), .B(A[227]), .Z(n321) );
  AND U352 ( .A(n322), .B(n323), .Z(n320) );
  NANDN U353 ( .A(B[226]), .B(n324), .Z(n323) );
  NANDN U354 ( .A(A[226]), .B(n325), .Z(n324) );
  NANDN U355 ( .A(n325), .B(A[226]), .Z(n322) );
  XOR U356 ( .A(n325), .B(n326), .Z(DIFF[226]) );
  XOR U357 ( .A(B[226]), .B(A[226]), .Z(n326) );
  AND U358 ( .A(n327), .B(n328), .Z(n325) );
  NANDN U359 ( .A(B[225]), .B(n329), .Z(n328) );
  NANDN U360 ( .A(A[225]), .B(n330), .Z(n329) );
  NANDN U361 ( .A(n330), .B(A[225]), .Z(n327) );
  XOR U362 ( .A(n330), .B(n331), .Z(DIFF[225]) );
  XOR U363 ( .A(B[225]), .B(A[225]), .Z(n331) );
  AND U364 ( .A(n332), .B(n333), .Z(n330) );
  NANDN U365 ( .A(B[224]), .B(n334), .Z(n333) );
  NANDN U366 ( .A(A[224]), .B(n335), .Z(n334) );
  NANDN U367 ( .A(n335), .B(A[224]), .Z(n332) );
  XOR U368 ( .A(n335), .B(n336), .Z(DIFF[224]) );
  XOR U369 ( .A(B[224]), .B(A[224]), .Z(n336) );
  AND U370 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U371 ( .A(B[223]), .B(n339), .Z(n338) );
  NANDN U372 ( .A(A[223]), .B(n340), .Z(n339) );
  NANDN U373 ( .A(n340), .B(A[223]), .Z(n337) );
  XOR U374 ( .A(n340), .B(n341), .Z(DIFF[223]) );
  XOR U375 ( .A(B[223]), .B(A[223]), .Z(n341) );
  AND U376 ( .A(n342), .B(n343), .Z(n340) );
  NANDN U377 ( .A(B[222]), .B(n344), .Z(n343) );
  NANDN U378 ( .A(A[222]), .B(n345), .Z(n344) );
  NANDN U379 ( .A(n345), .B(A[222]), .Z(n342) );
  XOR U380 ( .A(n345), .B(n346), .Z(DIFF[222]) );
  XOR U381 ( .A(B[222]), .B(A[222]), .Z(n346) );
  AND U382 ( .A(n347), .B(n348), .Z(n345) );
  NANDN U383 ( .A(B[221]), .B(n349), .Z(n348) );
  NANDN U384 ( .A(A[221]), .B(n350), .Z(n349) );
  NANDN U385 ( .A(n350), .B(A[221]), .Z(n347) );
  XOR U386 ( .A(n350), .B(n351), .Z(DIFF[221]) );
  XOR U387 ( .A(B[221]), .B(A[221]), .Z(n351) );
  AND U388 ( .A(n352), .B(n353), .Z(n350) );
  NANDN U389 ( .A(B[220]), .B(n354), .Z(n353) );
  NANDN U390 ( .A(A[220]), .B(n355), .Z(n354) );
  NANDN U391 ( .A(n355), .B(A[220]), .Z(n352) );
  XOR U392 ( .A(n355), .B(n356), .Z(DIFF[220]) );
  XOR U393 ( .A(B[220]), .B(A[220]), .Z(n356) );
  AND U394 ( .A(n357), .B(n358), .Z(n355) );
  NANDN U395 ( .A(B[219]), .B(n359), .Z(n358) );
  NANDN U396 ( .A(A[219]), .B(n360), .Z(n359) );
  NANDN U397 ( .A(n360), .B(A[219]), .Z(n357) );
  XOR U398 ( .A(n361), .B(n362), .Z(DIFF[21]) );
  XOR U399 ( .A(B[21]), .B(A[21]), .Z(n362) );
  XOR U400 ( .A(n360), .B(n363), .Z(DIFF[219]) );
  XOR U401 ( .A(B[219]), .B(A[219]), .Z(n363) );
  AND U402 ( .A(n364), .B(n365), .Z(n360) );
  NANDN U403 ( .A(B[218]), .B(n366), .Z(n365) );
  NANDN U404 ( .A(A[218]), .B(n367), .Z(n366) );
  NANDN U405 ( .A(n367), .B(A[218]), .Z(n364) );
  XOR U406 ( .A(n367), .B(n368), .Z(DIFF[218]) );
  XOR U407 ( .A(B[218]), .B(A[218]), .Z(n368) );
  AND U408 ( .A(n369), .B(n370), .Z(n367) );
  NANDN U409 ( .A(B[217]), .B(n371), .Z(n370) );
  NANDN U410 ( .A(A[217]), .B(n372), .Z(n371) );
  NANDN U411 ( .A(n372), .B(A[217]), .Z(n369) );
  XOR U412 ( .A(n372), .B(n373), .Z(DIFF[217]) );
  XOR U413 ( .A(B[217]), .B(A[217]), .Z(n373) );
  AND U414 ( .A(n374), .B(n375), .Z(n372) );
  NANDN U415 ( .A(B[216]), .B(n376), .Z(n375) );
  NANDN U416 ( .A(A[216]), .B(n377), .Z(n376) );
  NANDN U417 ( .A(n377), .B(A[216]), .Z(n374) );
  XOR U418 ( .A(n377), .B(n378), .Z(DIFF[216]) );
  XOR U419 ( .A(B[216]), .B(A[216]), .Z(n378) );
  AND U420 ( .A(n379), .B(n380), .Z(n377) );
  NANDN U421 ( .A(B[215]), .B(n381), .Z(n380) );
  NANDN U422 ( .A(A[215]), .B(n382), .Z(n381) );
  NANDN U423 ( .A(n382), .B(A[215]), .Z(n379) );
  XOR U424 ( .A(n382), .B(n383), .Z(DIFF[215]) );
  XOR U425 ( .A(B[215]), .B(A[215]), .Z(n383) );
  AND U426 ( .A(n384), .B(n385), .Z(n382) );
  NANDN U427 ( .A(B[214]), .B(n386), .Z(n385) );
  NANDN U428 ( .A(A[214]), .B(n387), .Z(n386) );
  NANDN U429 ( .A(n387), .B(A[214]), .Z(n384) );
  XOR U430 ( .A(n387), .B(n388), .Z(DIFF[214]) );
  XOR U431 ( .A(B[214]), .B(A[214]), .Z(n388) );
  AND U432 ( .A(n389), .B(n390), .Z(n387) );
  NANDN U433 ( .A(B[213]), .B(n391), .Z(n390) );
  NANDN U434 ( .A(A[213]), .B(n392), .Z(n391) );
  NANDN U435 ( .A(n392), .B(A[213]), .Z(n389) );
  XOR U436 ( .A(n392), .B(n393), .Z(DIFF[213]) );
  XOR U437 ( .A(B[213]), .B(A[213]), .Z(n393) );
  AND U438 ( .A(n394), .B(n395), .Z(n392) );
  NANDN U439 ( .A(B[212]), .B(n396), .Z(n395) );
  NANDN U440 ( .A(A[212]), .B(n397), .Z(n396) );
  NANDN U441 ( .A(n397), .B(A[212]), .Z(n394) );
  XOR U442 ( .A(n397), .B(n398), .Z(DIFF[212]) );
  XOR U443 ( .A(B[212]), .B(A[212]), .Z(n398) );
  AND U444 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U445 ( .A(B[211]), .B(n401), .Z(n400) );
  NANDN U446 ( .A(A[211]), .B(n402), .Z(n401) );
  NANDN U447 ( .A(n402), .B(A[211]), .Z(n399) );
  XOR U448 ( .A(n402), .B(n403), .Z(DIFF[211]) );
  XOR U449 ( .A(B[211]), .B(A[211]), .Z(n403) );
  AND U450 ( .A(n404), .B(n405), .Z(n402) );
  NANDN U451 ( .A(B[210]), .B(n406), .Z(n405) );
  NANDN U452 ( .A(A[210]), .B(n407), .Z(n406) );
  NANDN U453 ( .A(n407), .B(A[210]), .Z(n404) );
  XOR U454 ( .A(n407), .B(n408), .Z(DIFF[210]) );
  XOR U455 ( .A(B[210]), .B(A[210]), .Z(n408) );
  AND U456 ( .A(n409), .B(n410), .Z(n407) );
  NANDN U457 ( .A(B[209]), .B(n411), .Z(n410) );
  NANDN U458 ( .A(A[209]), .B(n412), .Z(n411) );
  NANDN U459 ( .A(n412), .B(A[209]), .Z(n409) );
  XOR U460 ( .A(n413), .B(n414), .Z(DIFF[20]) );
  XOR U461 ( .A(B[20]), .B(A[20]), .Z(n414) );
  XOR U462 ( .A(n412), .B(n415), .Z(DIFF[209]) );
  XOR U463 ( .A(B[209]), .B(A[209]), .Z(n415) );
  AND U464 ( .A(n416), .B(n417), .Z(n412) );
  NANDN U465 ( .A(B[208]), .B(n418), .Z(n417) );
  NANDN U466 ( .A(A[208]), .B(n419), .Z(n418) );
  NANDN U467 ( .A(n419), .B(A[208]), .Z(n416) );
  XOR U468 ( .A(n419), .B(n420), .Z(DIFF[208]) );
  XOR U469 ( .A(B[208]), .B(A[208]), .Z(n420) );
  AND U470 ( .A(n421), .B(n422), .Z(n419) );
  NANDN U471 ( .A(B[207]), .B(n423), .Z(n422) );
  NANDN U472 ( .A(A[207]), .B(n424), .Z(n423) );
  NANDN U473 ( .A(n424), .B(A[207]), .Z(n421) );
  XOR U474 ( .A(n424), .B(n425), .Z(DIFF[207]) );
  XOR U475 ( .A(B[207]), .B(A[207]), .Z(n425) );
  AND U476 ( .A(n426), .B(n427), .Z(n424) );
  NANDN U477 ( .A(B[206]), .B(n428), .Z(n427) );
  NANDN U478 ( .A(A[206]), .B(n429), .Z(n428) );
  NANDN U479 ( .A(n429), .B(A[206]), .Z(n426) );
  XOR U480 ( .A(n429), .B(n430), .Z(DIFF[206]) );
  XOR U481 ( .A(B[206]), .B(A[206]), .Z(n430) );
  AND U482 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U483 ( .A(B[205]), .B(n433), .Z(n432) );
  NANDN U484 ( .A(A[205]), .B(n434), .Z(n433) );
  NANDN U485 ( .A(n434), .B(A[205]), .Z(n431) );
  XOR U486 ( .A(n434), .B(n435), .Z(DIFF[205]) );
  XOR U487 ( .A(B[205]), .B(A[205]), .Z(n435) );
  AND U488 ( .A(n436), .B(n437), .Z(n434) );
  NANDN U489 ( .A(B[204]), .B(n438), .Z(n437) );
  NANDN U490 ( .A(A[204]), .B(n439), .Z(n438) );
  NANDN U491 ( .A(n439), .B(A[204]), .Z(n436) );
  XOR U492 ( .A(n439), .B(n440), .Z(DIFF[204]) );
  XOR U493 ( .A(B[204]), .B(A[204]), .Z(n440) );
  AND U494 ( .A(n441), .B(n442), .Z(n439) );
  NANDN U495 ( .A(B[203]), .B(n443), .Z(n442) );
  NANDN U496 ( .A(A[203]), .B(n444), .Z(n443) );
  NANDN U497 ( .A(n444), .B(A[203]), .Z(n441) );
  XOR U498 ( .A(n444), .B(n445), .Z(DIFF[203]) );
  XOR U499 ( .A(B[203]), .B(A[203]), .Z(n445) );
  AND U500 ( .A(n446), .B(n447), .Z(n444) );
  NANDN U501 ( .A(B[202]), .B(n448), .Z(n447) );
  NANDN U502 ( .A(A[202]), .B(n449), .Z(n448) );
  NANDN U503 ( .A(n449), .B(A[202]), .Z(n446) );
  XOR U504 ( .A(n449), .B(n450), .Z(DIFF[202]) );
  XOR U505 ( .A(B[202]), .B(A[202]), .Z(n450) );
  AND U506 ( .A(n451), .B(n452), .Z(n449) );
  NANDN U507 ( .A(B[201]), .B(n453), .Z(n452) );
  NANDN U508 ( .A(A[201]), .B(n454), .Z(n453) );
  NANDN U509 ( .A(n454), .B(A[201]), .Z(n451) );
  XOR U510 ( .A(n454), .B(n455), .Z(DIFF[201]) );
  XOR U511 ( .A(B[201]), .B(A[201]), .Z(n455) );
  AND U512 ( .A(n456), .B(n457), .Z(n454) );
  NANDN U513 ( .A(B[200]), .B(n458), .Z(n457) );
  NANDN U514 ( .A(A[200]), .B(n459), .Z(n458) );
  NANDN U515 ( .A(n459), .B(A[200]), .Z(n456) );
  XOR U516 ( .A(n459), .B(n460), .Z(DIFF[200]) );
  XOR U517 ( .A(B[200]), .B(A[200]), .Z(n460) );
  AND U518 ( .A(n461), .B(n462), .Z(n459) );
  NANDN U519 ( .A(B[199]), .B(n463), .Z(n462) );
  NANDN U520 ( .A(A[199]), .B(n464), .Z(n463) );
  NANDN U521 ( .A(n464), .B(A[199]), .Z(n461) );
  XOR U522 ( .A(n2), .B(n465), .Z(DIFF[1]) );
  XOR U523 ( .A(B[1]), .B(A[1]), .Z(n465) );
  XOR U524 ( .A(n466), .B(n467), .Z(DIFF[19]) );
  XOR U525 ( .A(B[19]), .B(A[19]), .Z(n467) );
  XOR U526 ( .A(n464), .B(n468), .Z(DIFF[199]) );
  XOR U527 ( .A(B[199]), .B(A[199]), .Z(n468) );
  AND U528 ( .A(n469), .B(n470), .Z(n464) );
  NANDN U529 ( .A(B[198]), .B(n471), .Z(n470) );
  NANDN U530 ( .A(A[198]), .B(n472), .Z(n471) );
  NANDN U531 ( .A(n472), .B(A[198]), .Z(n469) );
  XOR U532 ( .A(n472), .B(n473), .Z(DIFF[198]) );
  XOR U533 ( .A(B[198]), .B(A[198]), .Z(n473) );
  AND U534 ( .A(n474), .B(n475), .Z(n472) );
  NANDN U535 ( .A(B[197]), .B(n476), .Z(n475) );
  NANDN U536 ( .A(A[197]), .B(n477), .Z(n476) );
  NANDN U537 ( .A(n477), .B(A[197]), .Z(n474) );
  XOR U538 ( .A(n477), .B(n478), .Z(DIFF[197]) );
  XOR U539 ( .A(B[197]), .B(A[197]), .Z(n478) );
  AND U540 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U541 ( .A(B[196]), .B(n481), .Z(n480) );
  NANDN U542 ( .A(A[196]), .B(n482), .Z(n481) );
  NANDN U543 ( .A(n482), .B(A[196]), .Z(n479) );
  XOR U544 ( .A(n482), .B(n483), .Z(DIFF[196]) );
  XOR U545 ( .A(B[196]), .B(A[196]), .Z(n483) );
  AND U546 ( .A(n484), .B(n485), .Z(n482) );
  NANDN U547 ( .A(B[195]), .B(n486), .Z(n485) );
  NANDN U548 ( .A(A[195]), .B(n487), .Z(n486) );
  NANDN U549 ( .A(n487), .B(A[195]), .Z(n484) );
  XOR U550 ( .A(n487), .B(n488), .Z(DIFF[195]) );
  XOR U551 ( .A(B[195]), .B(A[195]), .Z(n488) );
  AND U552 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U553 ( .A(B[194]), .B(n491), .Z(n490) );
  NANDN U554 ( .A(A[194]), .B(n492), .Z(n491) );
  NANDN U555 ( .A(n492), .B(A[194]), .Z(n489) );
  XOR U556 ( .A(n492), .B(n493), .Z(DIFF[194]) );
  XOR U557 ( .A(B[194]), .B(A[194]), .Z(n493) );
  AND U558 ( .A(n494), .B(n495), .Z(n492) );
  NANDN U559 ( .A(B[193]), .B(n496), .Z(n495) );
  NANDN U560 ( .A(A[193]), .B(n497), .Z(n496) );
  NANDN U561 ( .A(n497), .B(A[193]), .Z(n494) );
  XOR U562 ( .A(n497), .B(n498), .Z(DIFF[193]) );
  XOR U563 ( .A(B[193]), .B(A[193]), .Z(n498) );
  AND U564 ( .A(n499), .B(n500), .Z(n497) );
  NANDN U565 ( .A(B[192]), .B(n501), .Z(n500) );
  NANDN U566 ( .A(A[192]), .B(n502), .Z(n501) );
  NANDN U567 ( .A(n502), .B(A[192]), .Z(n499) );
  XOR U568 ( .A(n502), .B(n503), .Z(DIFF[192]) );
  XOR U569 ( .A(B[192]), .B(A[192]), .Z(n503) );
  AND U570 ( .A(n504), .B(n505), .Z(n502) );
  NANDN U571 ( .A(B[191]), .B(n506), .Z(n505) );
  NANDN U572 ( .A(A[191]), .B(n507), .Z(n506) );
  NANDN U573 ( .A(n507), .B(A[191]), .Z(n504) );
  XOR U574 ( .A(n507), .B(n508), .Z(DIFF[191]) );
  XOR U575 ( .A(B[191]), .B(A[191]), .Z(n508) );
  AND U576 ( .A(n509), .B(n510), .Z(n507) );
  NANDN U577 ( .A(B[190]), .B(n511), .Z(n510) );
  NANDN U578 ( .A(A[190]), .B(n512), .Z(n511) );
  NANDN U579 ( .A(n512), .B(A[190]), .Z(n509) );
  XOR U580 ( .A(n512), .B(n513), .Z(DIFF[190]) );
  XOR U581 ( .A(B[190]), .B(A[190]), .Z(n513) );
  AND U582 ( .A(n514), .B(n515), .Z(n512) );
  NANDN U583 ( .A(B[189]), .B(n516), .Z(n515) );
  NANDN U584 ( .A(A[189]), .B(n517), .Z(n516) );
  NANDN U585 ( .A(n517), .B(A[189]), .Z(n514) );
  XOR U586 ( .A(n518), .B(n519), .Z(DIFF[18]) );
  XOR U587 ( .A(B[18]), .B(A[18]), .Z(n519) );
  XOR U588 ( .A(n517), .B(n520), .Z(DIFF[189]) );
  XOR U589 ( .A(B[189]), .B(A[189]), .Z(n520) );
  AND U590 ( .A(n521), .B(n522), .Z(n517) );
  NANDN U591 ( .A(B[188]), .B(n523), .Z(n522) );
  NANDN U592 ( .A(A[188]), .B(n524), .Z(n523) );
  NANDN U593 ( .A(n524), .B(A[188]), .Z(n521) );
  XOR U594 ( .A(n524), .B(n525), .Z(DIFF[188]) );
  XOR U595 ( .A(B[188]), .B(A[188]), .Z(n525) );
  AND U596 ( .A(n526), .B(n527), .Z(n524) );
  NANDN U597 ( .A(B[187]), .B(n528), .Z(n527) );
  NANDN U598 ( .A(A[187]), .B(n529), .Z(n528) );
  NANDN U599 ( .A(n529), .B(A[187]), .Z(n526) );
  XOR U600 ( .A(n529), .B(n530), .Z(DIFF[187]) );
  XOR U601 ( .A(B[187]), .B(A[187]), .Z(n530) );
  AND U602 ( .A(n531), .B(n532), .Z(n529) );
  NANDN U603 ( .A(B[186]), .B(n533), .Z(n532) );
  NANDN U604 ( .A(A[186]), .B(n534), .Z(n533) );
  NANDN U605 ( .A(n534), .B(A[186]), .Z(n531) );
  XOR U606 ( .A(n534), .B(n535), .Z(DIFF[186]) );
  XOR U607 ( .A(B[186]), .B(A[186]), .Z(n535) );
  AND U608 ( .A(n536), .B(n537), .Z(n534) );
  NANDN U609 ( .A(B[185]), .B(n538), .Z(n537) );
  NANDN U610 ( .A(A[185]), .B(n539), .Z(n538) );
  NANDN U611 ( .A(n539), .B(A[185]), .Z(n536) );
  XOR U612 ( .A(n539), .B(n540), .Z(DIFF[185]) );
  XOR U613 ( .A(B[185]), .B(A[185]), .Z(n540) );
  AND U614 ( .A(n541), .B(n542), .Z(n539) );
  NANDN U615 ( .A(B[184]), .B(n543), .Z(n542) );
  NANDN U616 ( .A(A[184]), .B(n544), .Z(n543) );
  NANDN U617 ( .A(n544), .B(A[184]), .Z(n541) );
  XOR U618 ( .A(n544), .B(n545), .Z(DIFF[184]) );
  XOR U619 ( .A(B[184]), .B(A[184]), .Z(n545) );
  AND U620 ( .A(n546), .B(n547), .Z(n544) );
  NANDN U621 ( .A(B[183]), .B(n548), .Z(n547) );
  NANDN U622 ( .A(A[183]), .B(n549), .Z(n548) );
  NANDN U623 ( .A(n549), .B(A[183]), .Z(n546) );
  XOR U624 ( .A(n549), .B(n550), .Z(DIFF[183]) );
  XOR U625 ( .A(B[183]), .B(A[183]), .Z(n550) );
  AND U626 ( .A(n551), .B(n552), .Z(n549) );
  NANDN U627 ( .A(B[182]), .B(n553), .Z(n552) );
  NANDN U628 ( .A(A[182]), .B(n554), .Z(n553) );
  NANDN U629 ( .A(n554), .B(A[182]), .Z(n551) );
  XOR U630 ( .A(n554), .B(n555), .Z(DIFF[182]) );
  XOR U631 ( .A(B[182]), .B(A[182]), .Z(n555) );
  AND U632 ( .A(n556), .B(n557), .Z(n554) );
  NANDN U633 ( .A(B[181]), .B(n558), .Z(n557) );
  NANDN U634 ( .A(A[181]), .B(n559), .Z(n558) );
  NANDN U635 ( .A(n559), .B(A[181]), .Z(n556) );
  XOR U636 ( .A(n559), .B(n560), .Z(DIFF[181]) );
  XOR U637 ( .A(B[181]), .B(A[181]), .Z(n560) );
  AND U638 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U639 ( .A(B[180]), .B(n563), .Z(n562) );
  NANDN U640 ( .A(A[180]), .B(n564), .Z(n563) );
  NANDN U641 ( .A(n564), .B(A[180]), .Z(n561) );
  XOR U642 ( .A(n564), .B(n565), .Z(DIFF[180]) );
  XOR U643 ( .A(B[180]), .B(A[180]), .Z(n565) );
  AND U644 ( .A(n566), .B(n567), .Z(n564) );
  NANDN U645 ( .A(B[179]), .B(n568), .Z(n567) );
  NANDN U646 ( .A(A[179]), .B(n569), .Z(n568) );
  NANDN U647 ( .A(n569), .B(A[179]), .Z(n566) );
  XOR U648 ( .A(n570), .B(n571), .Z(DIFF[17]) );
  XOR U649 ( .A(B[17]), .B(A[17]), .Z(n571) );
  XOR U650 ( .A(n569), .B(n572), .Z(DIFF[179]) );
  XOR U651 ( .A(B[179]), .B(A[179]), .Z(n572) );
  AND U652 ( .A(n573), .B(n574), .Z(n569) );
  NANDN U653 ( .A(B[178]), .B(n575), .Z(n574) );
  NANDN U654 ( .A(A[178]), .B(n576), .Z(n575) );
  NANDN U655 ( .A(n576), .B(A[178]), .Z(n573) );
  XOR U656 ( .A(n576), .B(n577), .Z(DIFF[178]) );
  XOR U657 ( .A(B[178]), .B(A[178]), .Z(n577) );
  AND U658 ( .A(n578), .B(n579), .Z(n576) );
  NANDN U659 ( .A(B[177]), .B(n580), .Z(n579) );
  NANDN U660 ( .A(A[177]), .B(n581), .Z(n580) );
  NANDN U661 ( .A(n581), .B(A[177]), .Z(n578) );
  XOR U662 ( .A(n581), .B(n582), .Z(DIFF[177]) );
  XOR U663 ( .A(B[177]), .B(A[177]), .Z(n582) );
  AND U664 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U665 ( .A(B[176]), .B(n585), .Z(n584) );
  NANDN U666 ( .A(A[176]), .B(n586), .Z(n585) );
  NANDN U667 ( .A(n586), .B(A[176]), .Z(n583) );
  XOR U668 ( .A(n586), .B(n587), .Z(DIFF[176]) );
  XOR U669 ( .A(B[176]), .B(A[176]), .Z(n587) );
  AND U670 ( .A(n588), .B(n589), .Z(n586) );
  NANDN U671 ( .A(B[175]), .B(n590), .Z(n589) );
  NANDN U672 ( .A(A[175]), .B(n591), .Z(n590) );
  NANDN U673 ( .A(n591), .B(A[175]), .Z(n588) );
  XOR U674 ( .A(n591), .B(n592), .Z(DIFF[175]) );
  XOR U675 ( .A(B[175]), .B(A[175]), .Z(n592) );
  AND U676 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U677 ( .A(B[174]), .B(n595), .Z(n594) );
  NANDN U678 ( .A(A[174]), .B(n596), .Z(n595) );
  NANDN U679 ( .A(n596), .B(A[174]), .Z(n593) );
  XOR U680 ( .A(n596), .B(n597), .Z(DIFF[174]) );
  XOR U681 ( .A(B[174]), .B(A[174]), .Z(n597) );
  AND U682 ( .A(n598), .B(n599), .Z(n596) );
  NANDN U683 ( .A(B[173]), .B(n600), .Z(n599) );
  NANDN U684 ( .A(A[173]), .B(n601), .Z(n600) );
  NANDN U685 ( .A(n601), .B(A[173]), .Z(n598) );
  XOR U686 ( .A(n601), .B(n602), .Z(DIFF[173]) );
  XOR U687 ( .A(B[173]), .B(A[173]), .Z(n602) );
  AND U688 ( .A(n603), .B(n604), .Z(n601) );
  NANDN U689 ( .A(B[172]), .B(n605), .Z(n604) );
  NANDN U690 ( .A(A[172]), .B(n606), .Z(n605) );
  NANDN U691 ( .A(n606), .B(A[172]), .Z(n603) );
  XOR U692 ( .A(n606), .B(n607), .Z(DIFF[172]) );
  XOR U693 ( .A(B[172]), .B(A[172]), .Z(n607) );
  AND U694 ( .A(n608), .B(n609), .Z(n606) );
  NANDN U695 ( .A(B[171]), .B(n610), .Z(n609) );
  NANDN U696 ( .A(A[171]), .B(n611), .Z(n610) );
  NANDN U697 ( .A(n611), .B(A[171]), .Z(n608) );
  XOR U698 ( .A(n611), .B(n612), .Z(DIFF[171]) );
  XOR U699 ( .A(B[171]), .B(A[171]), .Z(n612) );
  AND U700 ( .A(n613), .B(n614), .Z(n611) );
  NANDN U701 ( .A(B[170]), .B(n615), .Z(n614) );
  NANDN U702 ( .A(A[170]), .B(n616), .Z(n615) );
  NANDN U703 ( .A(n616), .B(A[170]), .Z(n613) );
  XOR U704 ( .A(n616), .B(n617), .Z(DIFF[170]) );
  XOR U705 ( .A(B[170]), .B(A[170]), .Z(n617) );
  AND U706 ( .A(n618), .B(n619), .Z(n616) );
  NANDN U707 ( .A(B[169]), .B(n620), .Z(n619) );
  NANDN U708 ( .A(A[169]), .B(n621), .Z(n620) );
  NANDN U709 ( .A(n621), .B(A[169]), .Z(n618) );
  XOR U710 ( .A(n622), .B(n623), .Z(DIFF[16]) );
  XOR U711 ( .A(B[16]), .B(A[16]), .Z(n623) );
  XOR U712 ( .A(n621), .B(n624), .Z(DIFF[169]) );
  XOR U713 ( .A(B[169]), .B(A[169]), .Z(n624) );
  AND U714 ( .A(n625), .B(n626), .Z(n621) );
  NANDN U715 ( .A(B[168]), .B(n627), .Z(n626) );
  NANDN U716 ( .A(A[168]), .B(n628), .Z(n627) );
  NANDN U717 ( .A(n628), .B(A[168]), .Z(n625) );
  XOR U718 ( .A(n628), .B(n629), .Z(DIFF[168]) );
  XOR U719 ( .A(B[168]), .B(A[168]), .Z(n629) );
  AND U720 ( .A(n630), .B(n631), .Z(n628) );
  NANDN U721 ( .A(B[167]), .B(n632), .Z(n631) );
  NANDN U722 ( .A(A[167]), .B(n633), .Z(n632) );
  NANDN U723 ( .A(n633), .B(A[167]), .Z(n630) );
  XOR U724 ( .A(n633), .B(n634), .Z(DIFF[167]) );
  XOR U725 ( .A(B[167]), .B(A[167]), .Z(n634) );
  AND U726 ( .A(n635), .B(n636), .Z(n633) );
  NANDN U727 ( .A(B[166]), .B(n637), .Z(n636) );
  NANDN U728 ( .A(A[166]), .B(n638), .Z(n637) );
  NANDN U729 ( .A(n638), .B(A[166]), .Z(n635) );
  XOR U730 ( .A(n638), .B(n639), .Z(DIFF[166]) );
  XOR U731 ( .A(B[166]), .B(A[166]), .Z(n639) );
  AND U732 ( .A(n640), .B(n641), .Z(n638) );
  NANDN U733 ( .A(B[165]), .B(n642), .Z(n641) );
  NANDN U734 ( .A(A[165]), .B(n643), .Z(n642) );
  NANDN U735 ( .A(n643), .B(A[165]), .Z(n640) );
  XOR U736 ( .A(n643), .B(n644), .Z(DIFF[165]) );
  XOR U737 ( .A(B[165]), .B(A[165]), .Z(n644) );
  AND U738 ( .A(n645), .B(n646), .Z(n643) );
  NANDN U739 ( .A(B[164]), .B(n647), .Z(n646) );
  NANDN U740 ( .A(A[164]), .B(n648), .Z(n647) );
  NANDN U741 ( .A(n648), .B(A[164]), .Z(n645) );
  XOR U742 ( .A(n648), .B(n649), .Z(DIFF[164]) );
  XOR U743 ( .A(B[164]), .B(A[164]), .Z(n649) );
  AND U744 ( .A(n650), .B(n651), .Z(n648) );
  NANDN U745 ( .A(B[163]), .B(n652), .Z(n651) );
  NANDN U746 ( .A(A[163]), .B(n653), .Z(n652) );
  NANDN U747 ( .A(n653), .B(A[163]), .Z(n650) );
  XOR U748 ( .A(n653), .B(n654), .Z(DIFF[163]) );
  XOR U749 ( .A(B[163]), .B(A[163]), .Z(n654) );
  AND U750 ( .A(n655), .B(n656), .Z(n653) );
  NANDN U751 ( .A(B[162]), .B(n657), .Z(n656) );
  NANDN U752 ( .A(A[162]), .B(n658), .Z(n657) );
  NANDN U753 ( .A(n658), .B(A[162]), .Z(n655) );
  XOR U754 ( .A(n658), .B(n659), .Z(DIFF[162]) );
  XOR U755 ( .A(B[162]), .B(A[162]), .Z(n659) );
  AND U756 ( .A(n660), .B(n661), .Z(n658) );
  NANDN U757 ( .A(B[161]), .B(n662), .Z(n661) );
  NANDN U758 ( .A(A[161]), .B(n663), .Z(n662) );
  NANDN U759 ( .A(n663), .B(A[161]), .Z(n660) );
  XOR U760 ( .A(n663), .B(n664), .Z(DIFF[161]) );
  XOR U761 ( .A(B[161]), .B(A[161]), .Z(n664) );
  AND U762 ( .A(n665), .B(n666), .Z(n663) );
  NANDN U763 ( .A(B[160]), .B(n667), .Z(n666) );
  NANDN U764 ( .A(A[160]), .B(n668), .Z(n667) );
  NANDN U765 ( .A(n668), .B(A[160]), .Z(n665) );
  XOR U766 ( .A(n668), .B(n669), .Z(DIFF[160]) );
  XOR U767 ( .A(B[160]), .B(A[160]), .Z(n669) );
  AND U768 ( .A(n670), .B(n671), .Z(n668) );
  NANDN U769 ( .A(B[159]), .B(n672), .Z(n671) );
  NANDN U770 ( .A(A[159]), .B(n673), .Z(n672) );
  NANDN U771 ( .A(n673), .B(A[159]), .Z(n670) );
  XOR U772 ( .A(n674), .B(n675), .Z(DIFF[15]) );
  XOR U773 ( .A(B[15]), .B(A[15]), .Z(n675) );
  XOR U774 ( .A(n673), .B(n676), .Z(DIFF[159]) );
  XOR U775 ( .A(B[159]), .B(A[159]), .Z(n676) );
  AND U776 ( .A(n677), .B(n678), .Z(n673) );
  NANDN U777 ( .A(B[158]), .B(n679), .Z(n678) );
  NANDN U778 ( .A(A[158]), .B(n680), .Z(n679) );
  NANDN U779 ( .A(n680), .B(A[158]), .Z(n677) );
  XOR U780 ( .A(n680), .B(n681), .Z(DIFF[158]) );
  XOR U781 ( .A(B[158]), .B(A[158]), .Z(n681) );
  AND U782 ( .A(n682), .B(n683), .Z(n680) );
  NANDN U783 ( .A(B[157]), .B(n684), .Z(n683) );
  NANDN U784 ( .A(A[157]), .B(n685), .Z(n684) );
  NANDN U785 ( .A(n685), .B(A[157]), .Z(n682) );
  XOR U786 ( .A(n685), .B(n686), .Z(DIFF[157]) );
  XOR U787 ( .A(B[157]), .B(A[157]), .Z(n686) );
  AND U788 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U789 ( .A(B[156]), .B(n689), .Z(n688) );
  NANDN U790 ( .A(A[156]), .B(n690), .Z(n689) );
  NANDN U791 ( .A(n690), .B(A[156]), .Z(n687) );
  XOR U792 ( .A(n690), .B(n691), .Z(DIFF[156]) );
  XOR U793 ( .A(B[156]), .B(A[156]), .Z(n691) );
  AND U794 ( .A(n692), .B(n693), .Z(n690) );
  NANDN U795 ( .A(B[155]), .B(n694), .Z(n693) );
  NANDN U796 ( .A(A[155]), .B(n695), .Z(n694) );
  NANDN U797 ( .A(n695), .B(A[155]), .Z(n692) );
  XOR U798 ( .A(n695), .B(n696), .Z(DIFF[155]) );
  XOR U799 ( .A(B[155]), .B(A[155]), .Z(n696) );
  AND U800 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U801 ( .A(B[154]), .B(n699), .Z(n698) );
  NANDN U802 ( .A(A[154]), .B(n700), .Z(n699) );
  NANDN U803 ( .A(n700), .B(A[154]), .Z(n697) );
  XOR U804 ( .A(n700), .B(n701), .Z(DIFF[154]) );
  XOR U805 ( .A(B[154]), .B(A[154]), .Z(n701) );
  AND U806 ( .A(n702), .B(n703), .Z(n700) );
  NANDN U807 ( .A(B[153]), .B(n704), .Z(n703) );
  NANDN U808 ( .A(A[153]), .B(n705), .Z(n704) );
  NANDN U809 ( .A(n705), .B(A[153]), .Z(n702) );
  XOR U810 ( .A(n705), .B(n706), .Z(DIFF[153]) );
  XOR U811 ( .A(B[153]), .B(A[153]), .Z(n706) );
  AND U812 ( .A(n707), .B(n708), .Z(n705) );
  NANDN U813 ( .A(B[152]), .B(n709), .Z(n708) );
  NANDN U814 ( .A(A[152]), .B(n710), .Z(n709) );
  NANDN U815 ( .A(n710), .B(A[152]), .Z(n707) );
  XOR U816 ( .A(n710), .B(n711), .Z(DIFF[152]) );
  XOR U817 ( .A(B[152]), .B(A[152]), .Z(n711) );
  AND U818 ( .A(n712), .B(n713), .Z(n710) );
  NANDN U819 ( .A(B[151]), .B(n714), .Z(n713) );
  NANDN U820 ( .A(A[151]), .B(n715), .Z(n714) );
  NANDN U821 ( .A(n715), .B(A[151]), .Z(n712) );
  XOR U822 ( .A(n715), .B(n716), .Z(DIFF[151]) );
  XOR U823 ( .A(B[151]), .B(A[151]), .Z(n716) );
  AND U824 ( .A(n717), .B(n718), .Z(n715) );
  NANDN U825 ( .A(B[150]), .B(n719), .Z(n718) );
  NANDN U826 ( .A(A[150]), .B(n720), .Z(n719) );
  NANDN U827 ( .A(n720), .B(A[150]), .Z(n717) );
  XOR U828 ( .A(n720), .B(n721), .Z(DIFF[150]) );
  XOR U829 ( .A(B[150]), .B(A[150]), .Z(n721) );
  AND U830 ( .A(n722), .B(n723), .Z(n720) );
  NANDN U831 ( .A(B[149]), .B(n724), .Z(n723) );
  NANDN U832 ( .A(A[149]), .B(n725), .Z(n724) );
  NANDN U833 ( .A(n725), .B(A[149]), .Z(n722) );
  XOR U834 ( .A(n726), .B(n727), .Z(DIFF[14]) );
  XOR U835 ( .A(B[14]), .B(A[14]), .Z(n727) );
  XOR U836 ( .A(n725), .B(n728), .Z(DIFF[149]) );
  XOR U837 ( .A(B[149]), .B(A[149]), .Z(n728) );
  AND U838 ( .A(n729), .B(n730), .Z(n725) );
  NANDN U839 ( .A(B[148]), .B(n731), .Z(n730) );
  NANDN U840 ( .A(A[148]), .B(n732), .Z(n731) );
  NANDN U841 ( .A(n732), .B(A[148]), .Z(n729) );
  XOR U842 ( .A(n732), .B(n733), .Z(DIFF[148]) );
  XOR U843 ( .A(B[148]), .B(A[148]), .Z(n733) );
  AND U844 ( .A(n734), .B(n735), .Z(n732) );
  NANDN U845 ( .A(B[147]), .B(n736), .Z(n735) );
  NANDN U846 ( .A(A[147]), .B(n737), .Z(n736) );
  NANDN U847 ( .A(n737), .B(A[147]), .Z(n734) );
  XOR U848 ( .A(n737), .B(n738), .Z(DIFF[147]) );
  XOR U849 ( .A(B[147]), .B(A[147]), .Z(n738) );
  AND U850 ( .A(n739), .B(n740), .Z(n737) );
  NANDN U851 ( .A(B[146]), .B(n741), .Z(n740) );
  NANDN U852 ( .A(A[146]), .B(n742), .Z(n741) );
  NANDN U853 ( .A(n742), .B(A[146]), .Z(n739) );
  XOR U854 ( .A(n742), .B(n743), .Z(DIFF[146]) );
  XOR U855 ( .A(B[146]), .B(A[146]), .Z(n743) );
  AND U856 ( .A(n744), .B(n745), .Z(n742) );
  NANDN U857 ( .A(B[145]), .B(n746), .Z(n745) );
  NANDN U858 ( .A(A[145]), .B(n747), .Z(n746) );
  NANDN U859 ( .A(n747), .B(A[145]), .Z(n744) );
  XOR U860 ( .A(n747), .B(n748), .Z(DIFF[145]) );
  XOR U861 ( .A(B[145]), .B(A[145]), .Z(n748) );
  AND U862 ( .A(n749), .B(n750), .Z(n747) );
  NANDN U863 ( .A(B[144]), .B(n751), .Z(n750) );
  NANDN U864 ( .A(A[144]), .B(n752), .Z(n751) );
  NANDN U865 ( .A(n752), .B(A[144]), .Z(n749) );
  XOR U866 ( .A(n752), .B(n753), .Z(DIFF[144]) );
  XOR U867 ( .A(B[144]), .B(A[144]), .Z(n753) );
  AND U868 ( .A(n754), .B(n755), .Z(n752) );
  NANDN U869 ( .A(B[143]), .B(n756), .Z(n755) );
  NANDN U870 ( .A(A[143]), .B(n757), .Z(n756) );
  NANDN U871 ( .A(n757), .B(A[143]), .Z(n754) );
  XOR U872 ( .A(n757), .B(n758), .Z(DIFF[143]) );
  XOR U873 ( .A(B[143]), .B(A[143]), .Z(n758) );
  AND U874 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U875 ( .A(B[142]), .B(n761), .Z(n760) );
  NANDN U876 ( .A(A[142]), .B(n762), .Z(n761) );
  NANDN U877 ( .A(n762), .B(A[142]), .Z(n759) );
  XOR U878 ( .A(n762), .B(n763), .Z(DIFF[142]) );
  XOR U879 ( .A(B[142]), .B(A[142]), .Z(n763) );
  AND U880 ( .A(n764), .B(n765), .Z(n762) );
  NANDN U881 ( .A(B[141]), .B(n766), .Z(n765) );
  NANDN U882 ( .A(A[141]), .B(n767), .Z(n766) );
  NANDN U883 ( .A(n767), .B(A[141]), .Z(n764) );
  XOR U884 ( .A(n767), .B(n768), .Z(DIFF[141]) );
  XOR U885 ( .A(B[141]), .B(A[141]), .Z(n768) );
  AND U886 ( .A(n769), .B(n770), .Z(n767) );
  NANDN U887 ( .A(B[140]), .B(n771), .Z(n770) );
  NANDN U888 ( .A(A[140]), .B(n772), .Z(n771) );
  NANDN U889 ( .A(n772), .B(A[140]), .Z(n769) );
  XOR U890 ( .A(n772), .B(n773), .Z(DIFF[140]) );
  XOR U891 ( .A(B[140]), .B(A[140]), .Z(n773) );
  AND U892 ( .A(n774), .B(n775), .Z(n772) );
  NANDN U893 ( .A(B[139]), .B(n776), .Z(n775) );
  NANDN U894 ( .A(A[139]), .B(n777), .Z(n776) );
  NANDN U895 ( .A(n777), .B(A[139]), .Z(n774) );
  XOR U896 ( .A(n778), .B(n779), .Z(DIFF[13]) );
  XOR U897 ( .A(B[13]), .B(A[13]), .Z(n779) );
  XOR U898 ( .A(n777), .B(n780), .Z(DIFF[139]) );
  XOR U899 ( .A(B[139]), .B(A[139]), .Z(n780) );
  AND U900 ( .A(n781), .B(n782), .Z(n777) );
  NANDN U901 ( .A(B[138]), .B(n783), .Z(n782) );
  NANDN U902 ( .A(A[138]), .B(n784), .Z(n783) );
  NANDN U903 ( .A(n784), .B(A[138]), .Z(n781) );
  XOR U904 ( .A(n784), .B(n785), .Z(DIFF[138]) );
  XOR U905 ( .A(B[138]), .B(A[138]), .Z(n785) );
  AND U906 ( .A(n786), .B(n787), .Z(n784) );
  NANDN U907 ( .A(B[137]), .B(n788), .Z(n787) );
  NANDN U908 ( .A(A[137]), .B(n789), .Z(n788) );
  NANDN U909 ( .A(n789), .B(A[137]), .Z(n786) );
  XOR U910 ( .A(n789), .B(n790), .Z(DIFF[137]) );
  XOR U911 ( .A(B[137]), .B(A[137]), .Z(n790) );
  AND U912 ( .A(n791), .B(n792), .Z(n789) );
  NANDN U913 ( .A(B[136]), .B(n793), .Z(n792) );
  NANDN U914 ( .A(A[136]), .B(n794), .Z(n793) );
  NANDN U915 ( .A(n794), .B(A[136]), .Z(n791) );
  XOR U916 ( .A(n794), .B(n795), .Z(DIFF[136]) );
  XOR U917 ( .A(B[136]), .B(A[136]), .Z(n795) );
  AND U918 ( .A(n796), .B(n797), .Z(n794) );
  NANDN U919 ( .A(B[135]), .B(n798), .Z(n797) );
  NANDN U920 ( .A(A[135]), .B(n799), .Z(n798) );
  NANDN U921 ( .A(n799), .B(A[135]), .Z(n796) );
  XOR U922 ( .A(n799), .B(n800), .Z(DIFF[135]) );
  XOR U923 ( .A(B[135]), .B(A[135]), .Z(n800) );
  AND U924 ( .A(n801), .B(n802), .Z(n799) );
  NANDN U925 ( .A(B[134]), .B(n803), .Z(n802) );
  NANDN U926 ( .A(A[134]), .B(n804), .Z(n803) );
  NANDN U927 ( .A(n804), .B(A[134]), .Z(n801) );
  XOR U928 ( .A(n804), .B(n805), .Z(DIFF[134]) );
  XOR U929 ( .A(B[134]), .B(A[134]), .Z(n805) );
  AND U930 ( .A(n806), .B(n807), .Z(n804) );
  NANDN U931 ( .A(B[133]), .B(n808), .Z(n807) );
  NANDN U932 ( .A(A[133]), .B(n809), .Z(n808) );
  NANDN U933 ( .A(n809), .B(A[133]), .Z(n806) );
  XOR U934 ( .A(n809), .B(n810), .Z(DIFF[133]) );
  XOR U935 ( .A(B[133]), .B(A[133]), .Z(n810) );
  AND U936 ( .A(n811), .B(n812), .Z(n809) );
  NANDN U937 ( .A(B[132]), .B(n813), .Z(n812) );
  NANDN U938 ( .A(A[132]), .B(n814), .Z(n813) );
  NANDN U939 ( .A(n814), .B(A[132]), .Z(n811) );
  XOR U940 ( .A(n814), .B(n815), .Z(DIFF[132]) );
  XOR U941 ( .A(B[132]), .B(A[132]), .Z(n815) );
  AND U942 ( .A(n816), .B(n817), .Z(n814) );
  NANDN U943 ( .A(B[131]), .B(n818), .Z(n817) );
  NANDN U944 ( .A(A[131]), .B(n819), .Z(n818) );
  NANDN U945 ( .A(n819), .B(A[131]), .Z(n816) );
  XOR U946 ( .A(n819), .B(n820), .Z(DIFF[131]) );
  XOR U947 ( .A(B[131]), .B(A[131]), .Z(n820) );
  AND U948 ( .A(n821), .B(n822), .Z(n819) );
  NANDN U949 ( .A(B[130]), .B(n823), .Z(n822) );
  NANDN U950 ( .A(A[130]), .B(n824), .Z(n823) );
  NANDN U951 ( .A(n824), .B(A[130]), .Z(n821) );
  XOR U952 ( .A(n824), .B(n825), .Z(DIFF[130]) );
  XOR U953 ( .A(B[130]), .B(A[130]), .Z(n825) );
  AND U954 ( .A(n826), .B(n827), .Z(n824) );
  NANDN U955 ( .A(B[129]), .B(n828), .Z(n827) );
  NANDN U956 ( .A(A[129]), .B(n829), .Z(n828) );
  NANDN U957 ( .A(n829), .B(A[129]), .Z(n826) );
  XOR U958 ( .A(n830), .B(n831), .Z(DIFF[12]) );
  XOR U959 ( .A(B[12]), .B(A[12]), .Z(n831) );
  XOR U960 ( .A(n829), .B(n832), .Z(DIFF[129]) );
  XOR U961 ( .A(B[129]), .B(A[129]), .Z(n832) );
  AND U962 ( .A(n833), .B(n834), .Z(n829) );
  NANDN U963 ( .A(B[128]), .B(n835), .Z(n834) );
  NANDN U964 ( .A(A[128]), .B(n836), .Z(n835) );
  NANDN U965 ( .A(n836), .B(A[128]), .Z(n833) );
  XOR U966 ( .A(n836), .B(n837), .Z(DIFF[128]) );
  XOR U967 ( .A(B[128]), .B(A[128]), .Z(n837) );
  AND U968 ( .A(n838), .B(n839), .Z(n836) );
  NANDN U969 ( .A(B[127]), .B(n840), .Z(n839) );
  NANDN U970 ( .A(A[127]), .B(n841), .Z(n840) );
  NANDN U971 ( .A(n841), .B(A[127]), .Z(n838) );
  XOR U972 ( .A(n841), .B(n842), .Z(DIFF[127]) );
  XOR U973 ( .A(B[127]), .B(A[127]), .Z(n842) );
  AND U974 ( .A(n843), .B(n844), .Z(n841) );
  NANDN U975 ( .A(B[126]), .B(n845), .Z(n844) );
  NANDN U976 ( .A(A[126]), .B(n846), .Z(n845) );
  NANDN U977 ( .A(n846), .B(A[126]), .Z(n843) );
  XOR U978 ( .A(n846), .B(n847), .Z(DIFF[126]) );
  XOR U979 ( .A(B[126]), .B(A[126]), .Z(n847) );
  AND U980 ( .A(n848), .B(n849), .Z(n846) );
  NANDN U981 ( .A(B[125]), .B(n850), .Z(n849) );
  NANDN U982 ( .A(A[125]), .B(n851), .Z(n850) );
  NANDN U983 ( .A(n851), .B(A[125]), .Z(n848) );
  XOR U984 ( .A(n851), .B(n852), .Z(DIFF[125]) );
  XOR U985 ( .A(B[125]), .B(A[125]), .Z(n852) );
  AND U986 ( .A(n853), .B(n854), .Z(n851) );
  NANDN U987 ( .A(B[124]), .B(n855), .Z(n854) );
  NANDN U988 ( .A(A[124]), .B(n856), .Z(n855) );
  NANDN U989 ( .A(n856), .B(A[124]), .Z(n853) );
  XOR U990 ( .A(n856), .B(n857), .Z(DIFF[124]) );
  XOR U991 ( .A(B[124]), .B(A[124]), .Z(n857) );
  AND U992 ( .A(n858), .B(n859), .Z(n856) );
  NANDN U993 ( .A(B[123]), .B(n860), .Z(n859) );
  NANDN U994 ( .A(A[123]), .B(n861), .Z(n860) );
  NANDN U995 ( .A(n861), .B(A[123]), .Z(n858) );
  XOR U996 ( .A(n861), .B(n862), .Z(DIFF[123]) );
  XOR U997 ( .A(B[123]), .B(A[123]), .Z(n862) );
  AND U998 ( .A(n863), .B(n864), .Z(n861) );
  NANDN U999 ( .A(B[122]), .B(n865), .Z(n864) );
  NANDN U1000 ( .A(A[122]), .B(n866), .Z(n865) );
  NANDN U1001 ( .A(n866), .B(A[122]), .Z(n863) );
  XOR U1002 ( .A(n866), .B(n867), .Z(DIFF[122]) );
  XOR U1003 ( .A(B[122]), .B(A[122]), .Z(n867) );
  AND U1004 ( .A(n868), .B(n869), .Z(n866) );
  NANDN U1005 ( .A(B[121]), .B(n870), .Z(n869) );
  NANDN U1006 ( .A(A[121]), .B(n871), .Z(n870) );
  NANDN U1007 ( .A(n871), .B(A[121]), .Z(n868) );
  XOR U1008 ( .A(n871), .B(n872), .Z(DIFF[121]) );
  XOR U1009 ( .A(B[121]), .B(A[121]), .Z(n872) );
  AND U1010 ( .A(n873), .B(n874), .Z(n871) );
  NANDN U1011 ( .A(B[120]), .B(n875), .Z(n874) );
  NANDN U1012 ( .A(A[120]), .B(n876), .Z(n875) );
  NANDN U1013 ( .A(n876), .B(A[120]), .Z(n873) );
  XOR U1014 ( .A(n876), .B(n877), .Z(DIFF[120]) );
  XOR U1015 ( .A(B[120]), .B(A[120]), .Z(n877) );
  AND U1016 ( .A(n878), .B(n879), .Z(n876) );
  NANDN U1017 ( .A(B[119]), .B(n880), .Z(n879) );
  NANDN U1018 ( .A(A[119]), .B(n881), .Z(n880) );
  NANDN U1019 ( .A(n881), .B(A[119]), .Z(n878) );
  XOR U1020 ( .A(n882), .B(n883), .Z(DIFF[11]) );
  XOR U1021 ( .A(B[11]), .B(A[11]), .Z(n883) );
  XOR U1022 ( .A(n881), .B(n884), .Z(DIFF[119]) );
  XOR U1023 ( .A(B[119]), .B(A[119]), .Z(n884) );
  AND U1024 ( .A(n885), .B(n886), .Z(n881) );
  NANDN U1025 ( .A(B[118]), .B(n887), .Z(n886) );
  NANDN U1026 ( .A(A[118]), .B(n888), .Z(n887) );
  NANDN U1027 ( .A(n888), .B(A[118]), .Z(n885) );
  XOR U1028 ( .A(n888), .B(n889), .Z(DIFF[118]) );
  XOR U1029 ( .A(B[118]), .B(A[118]), .Z(n889) );
  AND U1030 ( .A(n890), .B(n891), .Z(n888) );
  NANDN U1031 ( .A(B[117]), .B(n892), .Z(n891) );
  NANDN U1032 ( .A(A[117]), .B(n893), .Z(n892) );
  NANDN U1033 ( .A(n893), .B(A[117]), .Z(n890) );
  XOR U1034 ( .A(n893), .B(n894), .Z(DIFF[117]) );
  XOR U1035 ( .A(B[117]), .B(A[117]), .Z(n894) );
  AND U1036 ( .A(n895), .B(n896), .Z(n893) );
  NANDN U1037 ( .A(B[116]), .B(n897), .Z(n896) );
  NANDN U1038 ( .A(A[116]), .B(n898), .Z(n897) );
  NANDN U1039 ( .A(n898), .B(A[116]), .Z(n895) );
  XOR U1040 ( .A(n898), .B(n899), .Z(DIFF[116]) );
  XOR U1041 ( .A(B[116]), .B(A[116]), .Z(n899) );
  AND U1042 ( .A(n900), .B(n901), .Z(n898) );
  NANDN U1043 ( .A(B[115]), .B(n902), .Z(n901) );
  NANDN U1044 ( .A(A[115]), .B(n903), .Z(n902) );
  NANDN U1045 ( .A(n903), .B(A[115]), .Z(n900) );
  XOR U1046 ( .A(n903), .B(n904), .Z(DIFF[115]) );
  XOR U1047 ( .A(B[115]), .B(A[115]), .Z(n904) );
  AND U1048 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U1049 ( .A(B[114]), .B(n907), .Z(n906) );
  NANDN U1050 ( .A(A[114]), .B(n908), .Z(n907) );
  NANDN U1051 ( .A(n908), .B(A[114]), .Z(n905) );
  XOR U1052 ( .A(n908), .B(n909), .Z(DIFF[114]) );
  XOR U1053 ( .A(B[114]), .B(A[114]), .Z(n909) );
  AND U1054 ( .A(n910), .B(n911), .Z(n908) );
  NANDN U1055 ( .A(B[113]), .B(n912), .Z(n911) );
  NANDN U1056 ( .A(A[113]), .B(n913), .Z(n912) );
  NANDN U1057 ( .A(n913), .B(A[113]), .Z(n910) );
  XOR U1058 ( .A(n913), .B(n914), .Z(DIFF[113]) );
  XOR U1059 ( .A(B[113]), .B(A[113]), .Z(n914) );
  AND U1060 ( .A(n915), .B(n916), .Z(n913) );
  NANDN U1061 ( .A(B[112]), .B(n917), .Z(n916) );
  NANDN U1062 ( .A(A[112]), .B(n918), .Z(n917) );
  NANDN U1063 ( .A(n918), .B(A[112]), .Z(n915) );
  XOR U1064 ( .A(n918), .B(n919), .Z(DIFF[112]) );
  XOR U1065 ( .A(B[112]), .B(A[112]), .Z(n919) );
  AND U1066 ( .A(n920), .B(n921), .Z(n918) );
  NANDN U1067 ( .A(B[111]), .B(n922), .Z(n921) );
  NANDN U1068 ( .A(A[111]), .B(n923), .Z(n922) );
  NANDN U1069 ( .A(n923), .B(A[111]), .Z(n920) );
  XOR U1070 ( .A(n923), .B(n924), .Z(DIFF[111]) );
  XOR U1071 ( .A(B[111]), .B(A[111]), .Z(n924) );
  AND U1072 ( .A(n925), .B(n926), .Z(n923) );
  NANDN U1073 ( .A(B[110]), .B(n927), .Z(n926) );
  NANDN U1074 ( .A(A[110]), .B(n928), .Z(n927) );
  NANDN U1075 ( .A(n928), .B(A[110]), .Z(n925) );
  XOR U1076 ( .A(n928), .B(n929), .Z(DIFF[110]) );
  XOR U1077 ( .A(B[110]), .B(A[110]), .Z(n929) );
  AND U1078 ( .A(n930), .B(n931), .Z(n928) );
  NANDN U1079 ( .A(B[109]), .B(n932), .Z(n931) );
  NANDN U1080 ( .A(A[109]), .B(n933), .Z(n932) );
  NANDN U1081 ( .A(n933), .B(A[109]), .Z(n930) );
  XOR U1082 ( .A(n934), .B(n935), .Z(DIFF[10]) );
  XOR U1083 ( .A(B[10]), .B(A[10]), .Z(n935) );
  XOR U1084 ( .A(n933), .B(n936), .Z(DIFF[109]) );
  XOR U1085 ( .A(B[109]), .B(A[109]), .Z(n936) );
  AND U1086 ( .A(n937), .B(n938), .Z(n933) );
  NANDN U1087 ( .A(B[108]), .B(n939), .Z(n938) );
  NANDN U1088 ( .A(A[108]), .B(n940), .Z(n939) );
  NANDN U1089 ( .A(n940), .B(A[108]), .Z(n937) );
  XOR U1090 ( .A(n940), .B(n941), .Z(DIFF[108]) );
  XOR U1091 ( .A(B[108]), .B(A[108]), .Z(n941) );
  AND U1092 ( .A(n942), .B(n943), .Z(n940) );
  NANDN U1093 ( .A(B[107]), .B(n944), .Z(n943) );
  NANDN U1094 ( .A(A[107]), .B(n945), .Z(n944) );
  NANDN U1095 ( .A(n945), .B(A[107]), .Z(n942) );
  XOR U1096 ( .A(n945), .B(n946), .Z(DIFF[107]) );
  XOR U1097 ( .A(B[107]), .B(A[107]), .Z(n946) );
  AND U1098 ( .A(n947), .B(n948), .Z(n945) );
  NANDN U1099 ( .A(B[106]), .B(n949), .Z(n948) );
  NANDN U1100 ( .A(A[106]), .B(n950), .Z(n949) );
  NANDN U1101 ( .A(n950), .B(A[106]), .Z(n947) );
  XOR U1102 ( .A(n950), .B(n951), .Z(DIFF[106]) );
  XOR U1103 ( .A(B[106]), .B(A[106]), .Z(n951) );
  AND U1104 ( .A(n952), .B(n953), .Z(n950) );
  NANDN U1105 ( .A(B[105]), .B(n954), .Z(n953) );
  NANDN U1106 ( .A(A[105]), .B(n955), .Z(n954) );
  NANDN U1107 ( .A(n955), .B(A[105]), .Z(n952) );
  XOR U1108 ( .A(n955), .B(n956), .Z(DIFF[105]) );
  XOR U1109 ( .A(B[105]), .B(A[105]), .Z(n956) );
  AND U1110 ( .A(n957), .B(n958), .Z(n955) );
  NANDN U1111 ( .A(B[104]), .B(n959), .Z(n958) );
  NANDN U1112 ( .A(A[104]), .B(n960), .Z(n959) );
  NANDN U1113 ( .A(n960), .B(A[104]), .Z(n957) );
  XOR U1114 ( .A(n960), .B(n961), .Z(DIFF[104]) );
  XOR U1115 ( .A(B[104]), .B(A[104]), .Z(n961) );
  AND U1116 ( .A(n962), .B(n963), .Z(n960) );
  NANDN U1117 ( .A(B[103]), .B(n964), .Z(n963) );
  NANDN U1118 ( .A(A[103]), .B(n965), .Z(n964) );
  NANDN U1119 ( .A(n965), .B(A[103]), .Z(n962) );
  XOR U1120 ( .A(n965), .B(n966), .Z(DIFF[103]) );
  XOR U1121 ( .A(B[103]), .B(A[103]), .Z(n966) );
  AND U1122 ( .A(n967), .B(n968), .Z(n965) );
  NANDN U1123 ( .A(B[102]), .B(n969), .Z(n968) );
  NANDN U1124 ( .A(A[102]), .B(n970), .Z(n969) );
  NANDN U1125 ( .A(n970), .B(A[102]), .Z(n967) );
  XOR U1126 ( .A(n970), .B(n971), .Z(DIFF[102]) );
  XOR U1127 ( .A(B[102]), .B(A[102]), .Z(n971) );
  AND U1128 ( .A(n972), .B(n973), .Z(n970) );
  NANDN U1129 ( .A(B[101]), .B(n974), .Z(n973) );
  NANDN U1130 ( .A(A[101]), .B(n975), .Z(n974) );
  NANDN U1131 ( .A(n975), .B(A[101]), .Z(n972) );
  XOR U1132 ( .A(n975), .B(n976), .Z(DIFF[101]) );
  XOR U1133 ( .A(B[101]), .B(A[101]), .Z(n976) );
  AND U1134 ( .A(n977), .B(n978), .Z(n975) );
  NANDN U1135 ( .A(B[100]), .B(n979), .Z(n978) );
  NANDN U1136 ( .A(A[100]), .B(n980), .Z(n979) );
  NANDN U1137 ( .A(n980), .B(A[100]), .Z(n977) );
  XOR U1138 ( .A(n980), .B(n981), .Z(DIFF[100]) );
  XOR U1139 ( .A(B[100]), .B(A[100]), .Z(n981) );
  AND U1140 ( .A(n982), .B(n983), .Z(n980) );
  NANDN U1141 ( .A(B[99]), .B(n984), .Z(n983) );
  OR U1142 ( .A(n5), .B(A[99]), .Z(n984) );
  NAND U1143 ( .A(A[99]), .B(n5), .Z(n982) );
  NAND U1144 ( .A(n985), .B(n986), .Z(n5) );
  NANDN U1145 ( .A(B[98]), .B(n987), .Z(n986) );
  NANDN U1146 ( .A(A[98]), .B(n7), .Z(n987) );
  NANDN U1147 ( .A(n7), .B(A[98]), .Z(n985) );
  AND U1148 ( .A(n988), .B(n989), .Z(n7) );
  NANDN U1149 ( .A(B[97]), .B(n990), .Z(n989) );
  NANDN U1150 ( .A(A[97]), .B(n9), .Z(n990) );
  NANDN U1151 ( .A(n9), .B(A[97]), .Z(n988) );
  AND U1152 ( .A(n991), .B(n992), .Z(n9) );
  NANDN U1153 ( .A(B[96]), .B(n993), .Z(n992) );
  NANDN U1154 ( .A(A[96]), .B(n11), .Z(n993) );
  NANDN U1155 ( .A(n11), .B(A[96]), .Z(n991) );
  AND U1156 ( .A(n994), .B(n995), .Z(n11) );
  NANDN U1157 ( .A(B[95]), .B(n996), .Z(n995) );
  NANDN U1158 ( .A(A[95]), .B(n13), .Z(n996) );
  NANDN U1159 ( .A(n13), .B(A[95]), .Z(n994) );
  AND U1160 ( .A(n997), .B(n998), .Z(n13) );
  NANDN U1161 ( .A(B[94]), .B(n999), .Z(n998) );
  NANDN U1162 ( .A(A[94]), .B(n15), .Z(n999) );
  NANDN U1163 ( .A(n15), .B(A[94]), .Z(n997) );
  AND U1164 ( .A(n1000), .B(n1001), .Z(n15) );
  NANDN U1165 ( .A(B[93]), .B(n1002), .Z(n1001) );
  NANDN U1166 ( .A(A[93]), .B(n17), .Z(n1002) );
  NANDN U1167 ( .A(n17), .B(A[93]), .Z(n1000) );
  AND U1168 ( .A(n1003), .B(n1004), .Z(n17) );
  NANDN U1169 ( .A(B[92]), .B(n1005), .Z(n1004) );
  NANDN U1170 ( .A(A[92]), .B(n19), .Z(n1005) );
  NANDN U1171 ( .A(n19), .B(A[92]), .Z(n1003) );
  AND U1172 ( .A(n1006), .B(n1007), .Z(n19) );
  NANDN U1173 ( .A(B[91]), .B(n1008), .Z(n1007) );
  NANDN U1174 ( .A(A[91]), .B(n21), .Z(n1008) );
  NANDN U1175 ( .A(n21), .B(A[91]), .Z(n1006) );
  AND U1176 ( .A(n1009), .B(n1010), .Z(n21) );
  NANDN U1177 ( .A(B[90]), .B(n1011), .Z(n1010) );
  NANDN U1178 ( .A(A[90]), .B(n23), .Z(n1011) );
  NANDN U1179 ( .A(n23), .B(A[90]), .Z(n1009) );
  AND U1180 ( .A(n1012), .B(n1013), .Z(n23) );
  NANDN U1181 ( .A(B[89]), .B(n1014), .Z(n1013) );
  NANDN U1182 ( .A(A[89]), .B(n27), .Z(n1014) );
  NANDN U1183 ( .A(n27), .B(A[89]), .Z(n1012) );
  AND U1184 ( .A(n1015), .B(n1016), .Z(n27) );
  NANDN U1185 ( .A(B[88]), .B(n1017), .Z(n1016) );
  NANDN U1186 ( .A(A[88]), .B(n29), .Z(n1017) );
  NANDN U1187 ( .A(n29), .B(A[88]), .Z(n1015) );
  AND U1188 ( .A(n1018), .B(n1019), .Z(n29) );
  NANDN U1189 ( .A(B[87]), .B(n1020), .Z(n1019) );
  NANDN U1190 ( .A(A[87]), .B(n31), .Z(n1020) );
  NANDN U1191 ( .A(n31), .B(A[87]), .Z(n1018) );
  AND U1192 ( .A(n1021), .B(n1022), .Z(n31) );
  NANDN U1193 ( .A(B[86]), .B(n1023), .Z(n1022) );
  NANDN U1194 ( .A(A[86]), .B(n33), .Z(n1023) );
  NANDN U1195 ( .A(n33), .B(A[86]), .Z(n1021) );
  AND U1196 ( .A(n1024), .B(n1025), .Z(n33) );
  NANDN U1197 ( .A(B[85]), .B(n1026), .Z(n1025) );
  NANDN U1198 ( .A(A[85]), .B(n35), .Z(n1026) );
  NANDN U1199 ( .A(n35), .B(A[85]), .Z(n1024) );
  AND U1200 ( .A(n1027), .B(n1028), .Z(n35) );
  NANDN U1201 ( .A(B[84]), .B(n1029), .Z(n1028) );
  NANDN U1202 ( .A(A[84]), .B(n37), .Z(n1029) );
  NANDN U1203 ( .A(n37), .B(A[84]), .Z(n1027) );
  AND U1204 ( .A(n1030), .B(n1031), .Z(n37) );
  NANDN U1205 ( .A(B[83]), .B(n1032), .Z(n1031) );
  NANDN U1206 ( .A(A[83]), .B(n39), .Z(n1032) );
  NANDN U1207 ( .A(n39), .B(A[83]), .Z(n1030) );
  AND U1208 ( .A(n1033), .B(n1034), .Z(n39) );
  NANDN U1209 ( .A(B[82]), .B(n1035), .Z(n1034) );
  NANDN U1210 ( .A(A[82]), .B(n41), .Z(n1035) );
  NANDN U1211 ( .A(n41), .B(A[82]), .Z(n1033) );
  AND U1212 ( .A(n1036), .B(n1037), .Z(n41) );
  NANDN U1213 ( .A(B[81]), .B(n1038), .Z(n1037) );
  NANDN U1214 ( .A(A[81]), .B(n43), .Z(n1038) );
  NANDN U1215 ( .A(n43), .B(A[81]), .Z(n1036) );
  AND U1216 ( .A(n1039), .B(n1040), .Z(n43) );
  NANDN U1217 ( .A(B[80]), .B(n1041), .Z(n1040) );
  NANDN U1218 ( .A(A[80]), .B(n45), .Z(n1041) );
  NANDN U1219 ( .A(n45), .B(A[80]), .Z(n1039) );
  AND U1220 ( .A(n1042), .B(n1043), .Z(n45) );
  NANDN U1221 ( .A(B[79]), .B(n1044), .Z(n1043) );
  NANDN U1222 ( .A(A[79]), .B(n49), .Z(n1044) );
  NANDN U1223 ( .A(n49), .B(A[79]), .Z(n1042) );
  AND U1224 ( .A(n1045), .B(n1046), .Z(n49) );
  NANDN U1225 ( .A(B[78]), .B(n1047), .Z(n1046) );
  NANDN U1226 ( .A(A[78]), .B(n51), .Z(n1047) );
  NANDN U1227 ( .A(n51), .B(A[78]), .Z(n1045) );
  AND U1228 ( .A(n1048), .B(n1049), .Z(n51) );
  NANDN U1229 ( .A(B[77]), .B(n1050), .Z(n1049) );
  NANDN U1230 ( .A(A[77]), .B(n53), .Z(n1050) );
  NANDN U1231 ( .A(n53), .B(A[77]), .Z(n1048) );
  AND U1232 ( .A(n1051), .B(n1052), .Z(n53) );
  NANDN U1233 ( .A(B[76]), .B(n1053), .Z(n1052) );
  NANDN U1234 ( .A(A[76]), .B(n55), .Z(n1053) );
  NANDN U1235 ( .A(n55), .B(A[76]), .Z(n1051) );
  AND U1236 ( .A(n1054), .B(n1055), .Z(n55) );
  NANDN U1237 ( .A(B[75]), .B(n1056), .Z(n1055) );
  NANDN U1238 ( .A(A[75]), .B(n57), .Z(n1056) );
  NANDN U1239 ( .A(n57), .B(A[75]), .Z(n1054) );
  AND U1240 ( .A(n1057), .B(n1058), .Z(n57) );
  NANDN U1241 ( .A(B[74]), .B(n1059), .Z(n1058) );
  NANDN U1242 ( .A(A[74]), .B(n59), .Z(n1059) );
  NANDN U1243 ( .A(n59), .B(A[74]), .Z(n1057) );
  AND U1244 ( .A(n1060), .B(n1061), .Z(n59) );
  NANDN U1245 ( .A(B[73]), .B(n1062), .Z(n1061) );
  NANDN U1246 ( .A(A[73]), .B(n61), .Z(n1062) );
  NANDN U1247 ( .A(n61), .B(A[73]), .Z(n1060) );
  AND U1248 ( .A(n1063), .B(n1064), .Z(n61) );
  NANDN U1249 ( .A(B[72]), .B(n1065), .Z(n1064) );
  NANDN U1250 ( .A(A[72]), .B(n63), .Z(n1065) );
  NANDN U1251 ( .A(n63), .B(A[72]), .Z(n1063) );
  AND U1252 ( .A(n1066), .B(n1067), .Z(n63) );
  NANDN U1253 ( .A(B[71]), .B(n1068), .Z(n1067) );
  NANDN U1254 ( .A(A[71]), .B(n65), .Z(n1068) );
  NANDN U1255 ( .A(n65), .B(A[71]), .Z(n1066) );
  AND U1256 ( .A(n1069), .B(n1070), .Z(n65) );
  NANDN U1257 ( .A(B[70]), .B(n1071), .Z(n1070) );
  NANDN U1258 ( .A(A[70]), .B(n67), .Z(n1071) );
  NANDN U1259 ( .A(n67), .B(A[70]), .Z(n1069) );
  AND U1260 ( .A(n1072), .B(n1073), .Z(n67) );
  NANDN U1261 ( .A(B[69]), .B(n1074), .Z(n1073) );
  NANDN U1262 ( .A(A[69]), .B(n71), .Z(n1074) );
  NANDN U1263 ( .A(n71), .B(A[69]), .Z(n1072) );
  AND U1264 ( .A(n1075), .B(n1076), .Z(n71) );
  NANDN U1265 ( .A(B[68]), .B(n1077), .Z(n1076) );
  NANDN U1266 ( .A(A[68]), .B(n73), .Z(n1077) );
  NANDN U1267 ( .A(n73), .B(A[68]), .Z(n1075) );
  AND U1268 ( .A(n1078), .B(n1079), .Z(n73) );
  NANDN U1269 ( .A(B[67]), .B(n1080), .Z(n1079) );
  NANDN U1270 ( .A(A[67]), .B(n75), .Z(n1080) );
  NANDN U1271 ( .A(n75), .B(A[67]), .Z(n1078) );
  AND U1272 ( .A(n1081), .B(n1082), .Z(n75) );
  NANDN U1273 ( .A(B[66]), .B(n1083), .Z(n1082) );
  NANDN U1274 ( .A(A[66]), .B(n77), .Z(n1083) );
  NANDN U1275 ( .A(n77), .B(A[66]), .Z(n1081) );
  AND U1276 ( .A(n1084), .B(n1085), .Z(n77) );
  NANDN U1277 ( .A(B[65]), .B(n1086), .Z(n1085) );
  NANDN U1278 ( .A(A[65]), .B(n79), .Z(n1086) );
  NANDN U1279 ( .A(n79), .B(A[65]), .Z(n1084) );
  AND U1280 ( .A(n1087), .B(n1088), .Z(n79) );
  NANDN U1281 ( .A(B[64]), .B(n1089), .Z(n1088) );
  NANDN U1282 ( .A(A[64]), .B(n81), .Z(n1089) );
  NANDN U1283 ( .A(n81), .B(A[64]), .Z(n1087) );
  AND U1284 ( .A(n1090), .B(n1091), .Z(n81) );
  NANDN U1285 ( .A(B[63]), .B(n1092), .Z(n1091) );
  NANDN U1286 ( .A(A[63]), .B(n83), .Z(n1092) );
  NANDN U1287 ( .A(n83), .B(A[63]), .Z(n1090) );
  AND U1288 ( .A(n1093), .B(n1094), .Z(n83) );
  NANDN U1289 ( .A(B[62]), .B(n1095), .Z(n1094) );
  NANDN U1290 ( .A(A[62]), .B(n85), .Z(n1095) );
  NANDN U1291 ( .A(n85), .B(A[62]), .Z(n1093) );
  AND U1292 ( .A(n1096), .B(n1097), .Z(n85) );
  NANDN U1293 ( .A(B[61]), .B(n1098), .Z(n1097) );
  NANDN U1294 ( .A(A[61]), .B(n87), .Z(n1098) );
  NANDN U1295 ( .A(n87), .B(A[61]), .Z(n1096) );
  AND U1296 ( .A(n1099), .B(n1100), .Z(n87) );
  NANDN U1297 ( .A(B[60]), .B(n1101), .Z(n1100) );
  NANDN U1298 ( .A(A[60]), .B(n89), .Z(n1101) );
  NANDN U1299 ( .A(n89), .B(A[60]), .Z(n1099) );
  AND U1300 ( .A(n1102), .B(n1103), .Z(n89) );
  NANDN U1301 ( .A(B[59]), .B(n1104), .Z(n1103) );
  NANDN U1302 ( .A(A[59]), .B(n93), .Z(n1104) );
  NANDN U1303 ( .A(n93), .B(A[59]), .Z(n1102) );
  AND U1304 ( .A(n1105), .B(n1106), .Z(n93) );
  NANDN U1305 ( .A(B[58]), .B(n1107), .Z(n1106) );
  NANDN U1306 ( .A(A[58]), .B(n95), .Z(n1107) );
  NANDN U1307 ( .A(n95), .B(A[58]), .Z(n1105) );
  AND U1308 ( .A(n1108), .B(n1109), .Z(n95) );
  NANDN U1309 ( .A(B[57]), .B(n1110), .Z(n1109) );
  NANDN U1310 ( .A(A[57]), .B(n97), .Z(n1110) );
  NANDN U1311 ( .A(n97), .B(A[57]), .Z(n1108) );
  AND U1312 ( .A(n1111), .B(n1112), .Z(n97) );
  NANDN U1313 ( .A(B[56]), .B(n1113), .Z(n1112) );
  NANDN U1314 ( .A(A[56]), .B(n99), .Z(n1113) );
  NANDN U1315 ( .A(n99), .B(A[56]), .Z(n1111) );
  AND U1316 ( .A(n1114), .B(n1115), .Z(n99) );
  NANDN U1317 ( .A(B[55]), .B(n1116), .Z(n1115) );
  NANDN U1318 ( .A(A[55]), .B(n101), .Z(n1116) );
  NANDN U1319 ( .A(n101), .B(A[55]), .Z(n1114) );
  AND U1320 ( .A(n1117), .B(n1118), .Z(n101) );
  NANDN U1321 ( .A(B[54]), .B(n1119), .Z(n1118) );
  NANDN U1322 ( .A(A[54]), .B(n103), .Z(n1119) );
  NANDN U1323 ( .A(n103), .B(A[54]), .Z(n1117) );
  AND U1324 ( .A(n1120), .B(n1121), .Z(n103) );
  NANDN U1325 ( .A(B[53]), .B(n1122), .Z(n1121) );
  NANDN U1326 ( .A(A[53]), .B(n105), .Z(n1122) );
  NANDN U1327 ( .A(n105), .B(A[53]), .Z(n1120) );
  AND U1328 ( .A(n1123), .B(n1124), .Z(n105) );
  NANDN U1329 ( .A(B[52]), .B(n1125), .Z(n1124) );
  NANDN U1330 ( .A(A[52]), .B(n107), .Z(n1125) );
  NANDN U1331 ( .A(n107), .B(A[52]), .Z(n1123) );
  AND U1332 ( .A(n1126), .B(n1127), .Z(n107) );
  NANDN U1333 ( .A(B[51]), .B(n1128), .Z(n1127) );
  NANDN U1334 ( .A(A[51]), .B(n109), .Z(n1128) );
  NANDN U1335 ( .A(n109), .B(A[51]), .Z(n1126) );
  AND U1336 ( .A(n1129), .B(n1130), .Z(n109) );
  NANDN U1337 ( .A(B[50]), .B(n1131), .Z(n1130) );
  NANDN U1338 ( .A(A[50]), .B(n111), .Z(n1131) );
  NANDN U1339 ( .A(n111), .B(A[50]), .Z(n1129) );
  AND U1340 ( .A(n1132), .B(n1133), .Z(n111) );
  NANDN U1341 ( .A(B[49]), .B(n1134), .Z(n1133) );
  NANDN U1342 ( .A(A[49]), .B(n115), .Z(n1134) );
  NANDN U1343 ( .A(n115), .B(A[49]), .Z(n1132) );
  AND U1344 ( .A(n1135), .B(n1136), .Z(n115) );
  NANDN U1345 ( .A(B[48]), .B(n1137), .Z(n1136) );
  NANDN U1346 ( .A(A[48]), .B(n117), .Z(n1137) );
  NANDN U1347 ( .A(n117), .B(A[48]), .Z(n1135) );
  AND U1348 ( .A(n1138), .B(n1139), .Z(n117) );
  NANDN U1349 ( .A(B[47]), .B(n1140), .Z(n1139) );
  NANDN U1350 ( .A(A[47]), .B(n119), .Z(n1140) );
  NANDN U1351 ( .A(n119), .B(A[47]), .Z(n1138) );
  AND U1352 ( .A(n1141), .B(n1142), .Z(n119) );
  NANDN U1353 ( .A(B[46]), .B(n1143), .Z(n1142) );
  NANDN U1354 ( .A(A[46]), .B(n121), .Z(n1143) );
  NANDN U1355 ( .A(n121), .B(A[46]), .Z(n1141) );
  AND U1356 ( .A(n1144), .B(n1145), .Z(n121) );
  NANDN U1357 ( .A(B[45]), .B(n1146), .Z(n1145) );
  NANDN U1358 ( .A(A[45]), .B(n123), .Z(n1146) );
  NANDN U1359 ( .A(n123), .B(A[45]), .Z(n1144) );
  AND U1360 ( .A(n1147), .B(n1148), .Z(n123) );
  NANDN U1361 ( .A(B[44]), .B(n1149), .Z(n1148) );
  NANDN U1362 ( .A(A[44]), .B(n125), .Z(n1149) );
  NANDN U1363 ( .A(n125), .B(A[44]), .Z(n1147) );
  AND U1364 ( .A(n1150), .B(n1151), .Z(n125) );
  NANDN U1365 ( .A(B[43]), .B(n1152), .Z(n1151) );
  NANDN U1366 ( .A(A[43]), .B(n127), .Z(n1152) );
  NANDN U1367 ( .A(n127), .B(A[43]), .Z(n1150) );
  AND U1368 ( .A(n1153), .B(n1154), .Z(n127) );
  NANDN U1369 ( .A(B[42]), .B(n1155), .Z(n1154) );
  NANDN U1370 ( .A(A[42]), .B(n129), .Z(n1155) );
  NANDN U1371 ( .A(n129), .B(A[42]), .Z(n1153) );
  AND U1372 ( .A(n1156), .B(n1157), .Z(n129) );
  NANDN U1373 ( .A(B[41]), .B(n1158), .Z(n1157) );
  NANDN U1374 ( .A(A[41]), .B(n131), .Z(n1158) );
  NANDN U1375 ( .A(n131), .B(A[41]), .Z(n1156) );
  AND U1376 ( .A(n1159), .B(n1160), .Z(n131) );
  NANDN U1377 ( .A(B[40]), .B(n1161), .Z(n1160) );
  NANDN U1378 ( .A(A[40]), .B(n133), .Z(n1161) );
  NANDN U1379 ( .A(n133), .B(A[40]), .Z(n1159) );
  AND U1380 ( .A(n1162), .B(n1163), .Z(n133) );
  NANDN U1381 ( .A(B[39]), .B(n1164), .Z(n1163) );
  NANDN U1382 ( .A(A[39]), .B(n137), .Z(n1164) );
  NANDN U1383 ( .A(n137), .B(A[39]), .Z(n1162) );
  AND U1384 ( .A(n1165), .B(n1166), .Z(n137) );
  NANDN U1385 ( .A(B[38]), .B(n1167), .Z(n1166) );
  NANDN U1386 ( .A(A[38]), .B(n139), .Z(n1167) );
  NANDN U1387 ( .A(n139), .B(A[38]), .Z(n1165) );
  AND U1388 ( .A(n1168), .B(n1169), .Z(n139) );
  NANDN U1389 ( .A(B[37]), .B(n1170), .Z(n1169) );
  NANDN U1390 ( .A(A[37]), .B(n141), .Z(n1170) );
  NANDN U1391 ( .A(n141), .B(A[37]), .Z(n1168) );
  AND U1392 ( .A(n1171), .B(n1172), .Z(n141) );
  NANDN U1393 ( .A(B[36]), .B(n1173), .Z(n1172) );
  NANDN U1394 ( .A(A[36]), .B(n143), .Z(n1173) );
  NANDN U1395 ( .A(n143), .B(A[36]), .Z(n1171) );
  AND U1396 ( .A(n1174), .B(n1175), .Z(n143) );
  NANDN U1397 ( .A(B[35]), .B(n1176), .Z(n1175) );
  NANDN U1398 ( .A(A[35]), .B(n145), .Z(n1176) );
  NANDN U1399 ( .A(n145), .B(A[35]), .Z(n1174) );
  AND U1400 ( .A(n1177), .B(n1178), .Z(n145) );
  NANDN U1401 ( .A(B[34]), .B(n1179), .Z(n1178) );
  NANDN U1402 ( .A(A[34]), .B(n147), .Z(n1179) );
  NANDN U1403 ( .A(n147), .B(A[34]), .Z(n1177) );
  AND U1404 ( .A(n1180), .B(n1181), .Z(n147) );
  NANDN U1405 ( .A(B[33]), .B(n1182), .Z(n1181) );
  NANDN U1406 ( .A(A[33]), .B(n149), .Z(n1182) );
  NANDN U1407 ( .A(n149), .B(A[33]), .Z(n1180) );
  AND U1408 ( .A(n1183), .B(n1184), .Z(n149) );
  NANDN U1409 ( .A(B[32]), .B(n1185), .Z(n1184) );
  NANDN U1410 ( .A(A[32]), .B(n151), .Z(n1185) );
  NANDN U1411 ( .A(n151), .B(A[32]), .Z(n1183) );
  AND U1412 ( .A(n1186), .B(n1187), .Z(n151) );
  NANDN U1413 ( .A(B[31]), .B(n1188), .Z(n1187) );
  NANDN U1414 ( .A(A[31]), .B(n153), .Z(n1188) );
  NANDN U1415 ( .A(n153), .B(A[31]), .Z(n1186) );
  AND U1416 ( .A(n1189), .B(n1190), .Z(n153) );
  NANDN U1417 ( .A(B[30]), .B(n1191), .Z(n1190) );
  NANDN U1418 ( .A(A[30]), .B(n155), .Z(n1191) );
  NANDN U1419 ( .A(n155), .B(A[30]), .Z(n1189) );
  AND U1420 ( .A(n1192), .B(n1193), .Z(n155) );
  NANDN U1421 ( .A(B[29]), .B(n1194), .Z(n1193) );
  NANDN U1422 ( .A(A[29]), .B(n159), .Z(n1194) );
  NANDN U1423 ( .A(n159), .B(A[29]), .Z(n1192) );
  AND U1424 ( .A(n1195), .B(n1196), .Z(n159) );
  NANDN U1425 ( .A(B[28]), .B(n1197), .Z(n1196) );
  NANDN U1426 ( .A(A[28]), .B(n161), .Z(n1197) );
  NANDN U1427 ( .A(n161), .B(A[28]), .Z(n1195) );
  AND U1428 ( .A(n1198), .B(n1199), .Z(n161) );
  NANDN U1429 ( .A(B[27]), .B(n1200), .Z(n1199) );
  NANDN U1430 ( .A(A[27]), .B(n163), .Z(n1200) );
  NANDN U1431 ( .A(n163), .B(A[27]), .Z(n1198) );
  AND U1432 ( .A(n1201), .B(n1202), .Z(n163) );
  NANDN U1433 ( .A(B[26]), .B(n1203), .Z(n1202) );
  NANDN U1434 ( .A(A[26]), .B(n165), .Z(n1203) );
  NANDN U1435 ( .A(n165), .B(A[26]), .Z(n1201) );
  AND U1436 ( .A(n1204), .B(n1205), .Z(n165) );
  NANDN U1437 ( .A(B[25]), .B(n1206), .Z(n1205) );
  NANDN U1438 ( .A(A[25]), .B(n167), .Z(n1206) );
  NANDN U1439 ( .A(n167), .B(A[25]), .Z(n1204) );
  AND U1440 ( .A(n1207), .B(n1208), .Z(n167) );
  NANDN U1441 ( .A(B[24]), .B(n1209), .Z(n1208) );
  NANDN U1442 ( .A(A[24]), .B(n205), .Z(n1209) );
  NANDN U1443 ( .A(n205), .B(A[24]), .Z(n1207) );
  AND U1444 ( .A(n1210), .B(n1211), .Z(n205) );
  NANDN U1445 ( .A(B[23]), .B(n1212), .Z(n1211) );
  NANDN U1446 ( .A(A[23]), .B(n257), .Z(n1212) );
  NANDN U1447 ( .A(n257), .B(A[23]), .Z(n1210) );
  AND U1448 ( .A(n1213), .B(n1214), .Z(n257) );
  NANDN U1449 ( .A(B[22]), .B(n1215), .Z(n1214) );
  NANDN U1450 ( .A(A[22]), .B(n309), .Z(n1215) );
  NANDN U1451 ( .A(n309), .B(A[22]), .Z(n1213) );
  AND U1452 ( .A(n1216), .B(n1217), .Z(n309) );
  NANDN U1453 ( .A(B[21]), .B(n1218), .Z(n1217) );
  NANDN U1454 ( .A(A[21]), .B(n361), .Z(n1218) );
  NANDN U1455 ( .A(n361), .B(A[21]), .Z(n1216) );
  AND U1456 ( .A(n1219), .B(n1220), .Z(n361) );
  NANDN U1457 ( .A(B[20]), .B(n1221), .Z(n1220) );
  NANDN U1458 ( .A(A[20]), .B(n413), .Z(n1221) );
  NANDN U1459 ( .A(n413), .B(A[20]), .Z(n1219) );
  AND U1460 ( .A(n1222), .B(n1223), .Z(n413) );
  NANDN U1461 ( .A(B[19]), .B(n1224), .Z(n1223) );
  NANDN U1462 ( .A(A[19]), .B(n466), .Z(n1224) );
  NANDN U1463 ( .A(n466), .B(A[19]), .Z(n1222) );
  AND U1464 ( .A(n1225), .B(n1226), .Z(n466) );
  NANDN U1465 ( .A(B[18]), .B(n1227), .Z(n1226) );
  NANDN U1466 ( .A(A[18]), .B(n518), .Z(n1227) );
  NANDN U1467 ( .A(n518), .B(A[18]), .Z(n1225) );
  AND U1468 ( .A(n1228), .B(n1229), .Z(n518) );
  NANDN U1469 ( .A(B[17]), .B(n1230), .Z(n1229) );
  NANDN U1470 ( .A(A[17]), .B(n570), .Z(n1230) );
  NANDN U1471 ( .A(n570), .B(A[17]), .Z(n1228) );
  AND U1472 ( .A(n1231), .B(n1232), .Z(n570) );
  NANDN U1473 ( .A(B[16]), .B(n1233), .Z(n1232) );
  NANDN U1474 ( .A(A[16]), .B(n622), .Z(n1233) );
  NANDN U1475 ( .A(n622), .B(A[16]), .Z(n1231) );
  AND U1476 ( .A(n1234), .B(n1235), .Z(n622) );
  NANDN U1477 ( .A(B[15]), .B(n1236), .Z(n1235) );
  NANDN U1478 ( .A(A[15]), .B(n674), .Z(n1236) );
  NANDN U1479 ( .A(n674), .B(A[15]), .Z(n1234) );
  AND U1480 ( .A(n1237), .B(n1238), .Z(n674) );
  NANDN U1481 ( .A(B[14]), .B(n1239), .Z(n1238) );
  NANDN U1482 ( .A(A[14]), .B(n726), .Z(n1239) );
  NANDN U1483 ( .A(n726), .B(A[14]), .Z(n1237) );
  AND U1484 ( .A(n1240), .B(n1241), .Z(n726) );
  NANDN U1485 ( .A(B[13]), .B(n1242), .Z(n1241) );
  NANDN U1486 ( .A(A[13]), .B(n778), .Z(n1242) );
  NANDN U1487 ( .A(n778), .B(A[13]), .Z(n1240) );
  AND U1488 ( .A(n1243), .B(n1244), .Z(n778) );
  NANDN U1489 ( .A(B[12]), .B(n1245), .Z(n1244) );
  NANDN U1490 ( .A(A[12]), .B(n830), .Z(n1245) );
  NANDN U1491 ( .A(n830), .B(A[12]), .Z(n1243) );
  AND U1492 ( .A(n1246), .B(n1247), .Z(n830) );
  NANDN U1493 ( .A(B[11]), .B(n1248), .Z(n1247) );
  NANDN U1494 ( .A(A[11]), .B(n882), .Z(n1248) );
  NANDN U1495 ( .A(n882), .B(A[11]), .Z(n1246) );
  AND U1496 ( .A(n1249), .B(n1250), .Z(n882) );
  NANDN U1497 ( .A(B[10]), .B(n1251), .Z(n1250) );
  NANDN U1498 ( .A(A[10]), .B(n934), .Z(n1251) );
  NANDN U1499 ( .A(n934), .B(A[10]), .Z(n1249) );
  AND U1500 ( .A(n1252), .B(n1253), .Z(n934) );
  NANDN U1501 ( .A(B[9]), .B(n1254), .Z(n1253) );
  OR U1502 ( .A(n3), .B(A[9]), .Z(n1254) );
  NAND U1503 ( .A(A[9]), .B(n3), .Z(n1252) );
  NAND U1504 ( .A(n1255), .B(n1256), .Z(n3) );
  NANDN U1505 ( .A(B[8]), .B(n1257), .Z(n1256) );
  NANDN U1506 ( .A(A[8]), .B(n25), .Z(n1257) );
  NANDN U1507 ( .A(n25), .B(A[8]), .Z(n1255) );
  AND U1508 ( .A(n1258), .B(n1259), .Z(n25) );
  NANDN U1509 ( .A(B[7]), .B(n1260), .Z(n1259) );
  NANDN U1510 ( .A(A[7]), .B(n47), .Z(n1260) );
  NANDN U1511 ( .A(n47), .B(A[7]), .Z(n1258) );
  AND U1512 ( .A(n1261), .B(n1262), .Z(n47) );
  NANDN U1513 ( .A(B[6]), .B(n1263), .Z(n1262) );
  NANDN U1514 ( .A(A[6]), .B(n69), .Z(n1263) );
  NANDN U1515 ( .A(n69), .B(A[6]), .Z(n1261) );
  AND U1516 ( .A(n1264), .B(n1265), .Z(n69) );
  NANDN U1517 ( .A(B[5]), .B(n1266), .Z(n1265) );
  NANDN U1518 ( .A(A[5]), .B(n91), .Z(n1266) );
  NANDN U1519 ( .A(n91), .B(A[5]), .Z(n1264) );
  AND U1520 ( .A(n1267), .B(n1268), .Z(n91) );
  NANDN U1521 ( .A(B[4]), .B(n1269), .Z(n1268) );
  NANDN U1522 ( .A(A[4]), .B(n113), .Z(n1269) );
  NANDN U1523 ( .A(n113), .B(A[4]), .Z(n1267) );
  AND U1524 ( .A(n1270), .B(n1271), .Z(n113) );
  NANDN U1525 ( .A(B[3]), .B(n1272), .Z(n1271) );
  NANDN U1526 ( .A(A[3]), .B(n135), .Z(n1272) );
  NANDN U1527 ( .A(n135), .B(A[3]), .Z(n1270) );
  AND U1528 ( .A(n1273), .B(n1274), .Z(n135) );
  NANDN U1529 ( .A(B[2]), .B(n1275), .Z(n1274) );
  NANDN U1530 ( .A(A[2]), .B(n157), .Z(n1275) );
  NANDN U1531 ( .A(n157), .B(A[2]), .Z(n1273) );
  AND U1532 ( .A(n1276), .B(n1277), .Z(n157) );
  NANDN U1533 ( .A(B[1]), .B(n1278), .Z(n1277) );
  NAND U1534 ( .A(n2), .B(n1), .Z(n1278) );
  NAND U1535 ( .A(A[1]), .B(n1279), .Z(n1276) );
  NAND U1536 ( .A(n1279), .B(n1280), .Z(DIFF[0]) );
  NANDN U1537 ( .A(B[0]), .B(A[0]), .Z(n1280) );
  NANDN U1538 ( .A(A[0]), .B(B[0]), .Z(n1279) );
endmodule


module modmult_step_N256_5_DW01_cmp2_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [257:0] A;
  input [257:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;

  NAND U1 ( .A(n1), .B(n2), .Z(LT_LE) );
  NOR U2 ( .A(B[257]), .B(B[256]), .Z(n2) );
  AND U3 ( .A(n3), .B(n4), .Z(n1) );
  NAND U4 ( .A(n5), .B(n6), .Z(n4) );
  NANDN U5 ( .A(B[255]), .B(A[255]), .Z(n6) );
  NAND U6 ( .A(n7), .B(n8), .Z(n5) );
  NANDN U7 ( .A(A[254]), .B(B[254]), .Z(n8) );
  NAND U8 ( .A(n9), .B(n10), .Z(n7) );
  NANDN U9 ( .A(B[254]), .B(A[254]), .Z(n10) );
  AND U10 ( .A(n11), .B(n12), .Z(n9) );
  NAND U11 ( .A(n13), .B(n14), .Z(n12) );
  NANDN U12 ( .A(A[253]), .B(B[253]), .Z(n14) );
  AND U13 ( .A(n15), .B(n16), .Z(n13) );
  NANDN U14 ( .A(A[252]), .B(B[252]), .Z(n16) );
  NAND U15 ( .A(n17), .B(n18), .Z(n15) );
  NANDN U16 ( .A(B[252]), .B(A[252]), .Z(n18) );
  AND U17 ( .A(n19), .B(n20), .Z(n17) );
  NAND U18 ( .A(n21), .B(n22), .Z(n20) );
  NANDN U19 ( .A(A[251]), .B(B[251]), .Z(n22) );
  AND U20 ( .A(n23), .B(n24), .Z(n21) );
  NANDN U21 ( .A(A[250]), .B(B[250]), .Z(n24) );
  NAND U22 ( .A(n25), .B(n26), .Z(n23) );
  NANDN U23 ( .A(B[250]), .B(A[250]), .Z(n26) );
  AND U24 ( .A(n27), .B(n28), .Z(n25) );
  NAND U25 ( .A(n29), .B(n30), .Z(n28) );
  NANDN U26 ( .A(A[249]), .B(B[249]), .Z(n30) );
  AND U27 ( .A(n31), .B(n32), .Z(n29) );
  NANDN U28 ( .A(A[248]), .B(B[248]), .Z(n32) );
  NAND U29 ( .A(n33), .B(n34), .Z(n31) );
  NANDN U30 ( .A(B[248]), .B(A[248]), .Z(n34) );
  AND U31 ( .A(n35), .B(n36), .Z(n33) );
  NAND U32 ( .A(n37), .B(n38), .Z(n36) );
  NANDN U33 ( .A(A[247]), .B(B[247]), .Z(n38) );
  AND U34 ( .A(n39), .B(n40), .Z(n37) );
  NANDN U35 ( .A(A[246]), .B(B[246]), .Z(n40) );
  NAND U36 ( .A(n41), .B(n42), .Z(n39) );
  NANDN U37 ( .A(B[246]), .B(A[246]), .Z(n42) );
  AND U38 ( .A(n43), .B(n44), .Z(n41) );
  NAND U39 ( .A(n45), .B(n46), .Z(n44) );
  NANDN U40 ( .A(A[245]), .B(B[245]), .Z(n46) );
  AND U41 ( .A(n47), .B(n48), .Z(n45) );
  NANDN U42 ( .A(A[244]), .B(B[244]), .Z(n48) );
  NAND U43 ( .A(n49), .B(n50), .Z(n47) );
  NANDN U44 ( .A(B[244]), .B(A[244]), .Z(n50) );
  AND U45 ( .A(n51), .B(n52), .Z(n49) );
  NAND U46 ( .A(n53), .B(n54), .Z(n52) );
  NANDN U47 ( .A(A[243]), .B(B[243]), .Z(n54) );
  AND U48 ( .A(n55), .B(n56), .Z(n53) );
  NANDN U49 ( .A(A[242]), .B(B[242]), .Z(n56) );
  NAND U50 ( .A(n57), .B(n58), .Z(n55) );
  NANDN U51 ( .A(B[242]), .B(A[242]), .Z(n58) );
  AND U52 ( .A(n59), .B(n60), .Z(n57) );
  NAND U53 ( .A(n61), .B(n62), .Z(n60) );
  NANDN U54 ( .A(A[241]), .B(B[241]), .Z(n62) );
  AND U55 ( .A(n63), .B(n64), .Z(n61) );
  NANDN U56 ( .A(A[240]), .B(B[240]), .Z(n64) );
  NAND U57 ( .A(n65), .B(n66), .Z(n63) );
  NANDN U58 ( .A(B[240]), .B(A[240]), .Z(n66) );
  AND U59 ( .A(n67), .B(n68), .Z(n65) );
  NAND U60 ( .A(n69), .B(n70), .Z(n68) );
  NANDN U61 ( .A(A[239]), .B(B[239]), .Z(n70) );
  AND U62 ( .A(n71), .B(n72), .Z(n69) );
  NANDN U63 ( .A(A[238]), .B(B[238]), .Z(n72) );
  NAND U64 ( .A(n73), .B(n74), .Z(n71) );
  NANDN U65 ( .A(B[238]), .B(A[238]), .Z(n74) );
  AND U66 ( .A(n75), .B(n76), .Z(n73) );
  NAND U67 ( .A(n77), .B(n78), .Z(n76) );
  NANDN U68 ( .A(A[237]), .B(B[237]), .Z(n78) );
  AND U69 ( .A(n79), .B(n80), .Z(n77) );
  NANDN U70 ( .A(A[236]), .B(B[236]), .Z(n80) );
  NAND U71 ( .A(n81), .B(n82), .Z(n79) );
  NANDN U72 ( .A(B[236]), .B(A[236]), .Z(n82) );
  AND U73 ( .A(n83), .B(n84), .Z(n81) );
  NAND U74 ( .A(n85), .B(n86), .Z(n84) );
  NANDN U75 ( .A(A[235]), .B(B[235]), .Z(n86) );
  AND U76 ( .A(n87), .B(n88), .Z(n85) );
  NANDN U77 ( .A(A[234]), .B(B[234]), .Z(n88) );
  NAND U78 ( .A(n89), .B(n90), .Z(n87) );
  NANDN U79 ( .A(B[234]), .B(A[234]), .Z(n90) );
  AND U80 ( .A(n91), .B(n92), .Z(n89) );
  NAND U81 ( .A(n93), .B(n94), .Z(n92) );
  NANDN U82 ( .A(A[233]), .B(B[233]), .Z(n94) );
  AND U83 ( .A(n95), .B(n96), .Z(n93) );
  NANDN U84 ( .A(A[232]), .B(B[232]), .Z(n96) );
  NAND U85 ( .A(n97), .B(n98), .Z(n95) );
  NANDN U86 ( .A(B[232]), .B(A[232]), .Z(n98) );
  AND U87 ( .A(n99), .B(n100), .Z(n97) );
  NAND U88 ( .A(n101), .B(n102), .Z(n100) );
  NANDN U89 ( .A(A[231]), .B(B[231]), .Z(n102) );
  AND U90 ( .A(n103), .B(n104), .Z(n101) );
  NANDN U91 ( .A(A[230]), .B(B[230]), .Z(n104) );
  NAND U92 ( .A(n105), .B(n106), .Z(n103) );
  NANDN U93 ( .A(B[230]), .B(A[230]), .Z(n106) );
  AND U94 ( .A(n107), .B(n108), .Z(n105) );
  NAND U95 ( .A(n109), .B(n110), .Z(n108) );
  NANDN U96 ( .A(A[229]), .B(B[229]), .Z(n110) );
  AND U97 ( .A(n111), .B(n112), .Z(n109) );
  NANDN U98 ( .A(A[228]), .B(B[228]), .Z(n112) );
  NAND U99 ( .A(n113), .B(n114), .Z(n111) );
  NANDN U100 ( .A(B[228]), .B(A[228]), .Z(n114) );
  AND U101 ( .A(n115), .B(n116), .Z(n113) );
  NAND U102 ( .A(n117), .B(n118), .Z(n116) );
  NANDN U103 ( .A(A[227]), .B(B[227]), .Z(n118) );
  AND U104 ( .A(n119), .B(n120), .Z(n117) );
  NANDN U105 ( .A(A[226]), .B(B[226]), .Z(n120) );
  NAND U106 ( .A(n121), .B(n122), .Z(n119) );
  NANDN U107 ( .A(B[226]), .B(A[226]), .Z(n122) );
  AND U108 ( .A(n123), .B(n124), .Z(n121) );
  NAND U109 ( .A(n125), .B(n126), .Z(n124) );
  NANDN U110 ( .A(A[225]), .B(B[225]), .Z(n126) );
  AND U111 ( .A(n127), .B(n128), .Z(n125) );
  NANDN U112 ( .A(A[224]), .B(B[224]), .Z(n128) );
  NAND U113 ( .A(n129), .B(n130), .Z(n127) );
  NANDN U114 ( .A(B[224]), .B(A[224]), .Z(n130) );
  AND U115 ( .A(n131), .B(n132), .Z(n129) );
  NAND U116 ( .A(n133), .B(n134), .Z(n132) );
  NANDN U117 ( .A(A[223]), .B(B[223]), .Z(n134) );
  AND U118 ( .A(n135), .B(n136), .Z(n133) );
  NANDN U119 ( .A(A[222]), .B(B[222]), .Z(n136) );
  NAND U120 ( .A(n137), .B(n138), .Z(n135) );
  NANDN U121 ( .A(B[222]), .B(A[222]), .Z(n138) );
  AND U122 ( .A(n139), .B(n140), .Z(n137) );
  NAND U123 ( .A(n141), .B(n142), .Z(n140) );
  NANDN U124 ( .A(A[221]), .B(B[221]), .Z(n142) );
  AND U125 ( .A(n143), .B(n144), .Z(n141) );
  NANDN U126 ( .A(A[220]), .B(B[220]), .Z(n144) );
  NAND U127 ( .A(n145), .B(n146), .Z(n143) );
  NANDN U128 ( .A(B[220]), .B(A[220]), .Z(n146) );
  AND U129 ( .A(n147), .B(n148), .Z(n145) );
  NAND U130 ( .A(n149), .B(n150), .Z(n148) );
  NANDN U131 ( .A(A[219]), .B(B[219]), .Z(n150) );
  AND U132 ( .A(n151), .B(n152), .Z(n149) );
  NANDN U133 ( .A(A[218]), .B(B[218]), .Z(n152) );
  NAND U134 ( .A(n153), .B(n154), .Z(n151) );
  NANDN U135 ( .A(B[218]), .B(A[218]), .Z(n154) );
  AND U136 ( .A(n155), .B(n156), .Z(n153) );
  NAND U137 ( .A(n157), .B(n158), .Z(n156) );
  NANDN U138 ( .A(A[217]), .B(B[217]), .Z(n158) );
  AND U139 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U140 ( .A(A[216]), .B(B[216]), .Z(n160) );
  NAND U141 ( .A(n161), .B(n162), .Z(n159) );
  NANDN U142 ( .A(B[216]), .B(A[216]), .Z(n162) );
  AND U143 ( .A(n163), .B(n164), .Z(n161) );
  NAND U144 ( .A(n165), .B(n166), .Z(n164) );
  NANDN U145 ( .A(A[215]), .B(B[215]), .Z(n166) );
  AND U146 ( .A(n167), .B(n168), .Z(n165) );
  NANDN U147 ( .A(A[214]), .B(B[214]), .Z(n168) );
  NAND U148 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U149 ( .A(B[214]), .B(A[214]), .Z(n170) );
  AND U150 ( .A(n171), .B(n172), .Z(n169) );
  NAND U151 ( .A(n173), .B(n174), .Z(n172) );
  NANDN U152 ( .A(A[213]), .B(B[213]), .Z(n174) );
  AND U153 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U154 ( .A(A[212]), .B(B[212]), .Z(n176) );
  NAND U155 ( .A(n177), .B(n178), .Z(n175) );
  NANDN U156 ( .A(B[212]), .B(A[212]), .Z(n178) );
  AND U157 ( .A(n179), .B(n180), .Z(n177) );
  NAND U158 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U159 ( .A(A[211]), .B(B[211]), .Z(n182) );
  AND U160 ( .A(n183), .B(n184), .Z(n181) );
  NANDN U161 ( .A(A[210]), .B(B[210]), .Z(n184) );
  NAND U162 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U163 ( .A(B[210]), .B(A[210]), .Z(n186) );
  AND U164 ( .A(n187), .B(n188), .Z(n185) );
  NAND U165 ( .A(n189), .B(n190), .Z(n188) );
  NANDN U166 ( .A(A[209]), .B(B[209]), .Z(n190) );
  AND U167 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U168 ( .A(A[208]), .B(B[208]), .Z(n192) );
  NAND U169 ( .A(n193), .B(n194), .Z(n191) );
  NANDN U170 ( .A(B[208]), .B(A[208]), .Z(n194) );
  AND U171 ( .A(n195), .B(n196), .Z(n193) );
  NAND U172 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U173 ( .A(A[207]), .B(B[207]), .Z(n198) );
  AND U174 ( .A(n199), .B(n200), .Z(n197) );
  NANDN U175 ( .A(A[206]), .B(B[206]), .Z(n200) );
  NAND U176 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U177 ( .A(B[206]), .B(A[206]), .Z(n202) );
  AND U178 ( .A(n203), .B(n204), .Z(n201) );
  NAND U179 ( .A(n205), .B(n206), .Z(n204) );
  NANDN U180 ( .A(A[205]), .B(B[205]), .Z(n206) );
  AND U181 ( .A(n207), .B(n208), .Z(n205) );
  NANDN U182 ( .A(A[204]), .B(B[204]), .Z(n208) );
  NAND U183 ( .A(n209), .B(n210), .Z(n207) );
  NANDN U184 ( .A(B[204]), .B(A[204]), .Z(n210) );
  AND U185 ( .A(n211), .B(n212), .Z(n209) );
  NAND U186 ( .A(n213), .B(n214), .Z(n212) );
  NANDN U187 ( .A(A[203]), .B(B[203]), .Z(n214) );
  AND U188 ( .A(n215), .B(n216), .Z(n213) );
  NANDN U189 ( .A(A[202]), .B(B[202]), .Z(n216) );
  NAND U190 ( .A(n217), .B(n218), .Z(n215) );
  NANDN U191 ( .A(B[202]), .B(A[202]), .Z(n218) );
  AND U192 ( .A(n219), .B(n220), .Z(n217) );
  NAND U193 ( .A(n221), .B(n222), .Z(n220) );
  NANDN U194 ( .A(A[201]), .B(B[201]), .Z(n222) );
  AND U195 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U196 ( .A(A[200]), .B(B[200]), .Z(n224) );
  NAND U197 ( .A(n225), .B(n226), .Z(n223) );
  NANDN U198 ( .A(B[200]), .B(A[200]), .Z(n226) );
  AND U199 ( .A(n227), .B(n228), .Z(n225) );
  NAND U200 ( .A(n229), .B(n230), .Z(n228) );
  NANDN U201 ( .A(A[199]), .B(B[199]), .Z(n230) );
  AND U202 ( .A(n231), .B(n232), .Z(n229) );
  NANDN U203 ( .A(A[198]), .B(B[198]), .Z(n232) );
  NAND U204 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U205 ( .A(B[198]), .B(A[198]), .Z(n234) );
  AND U206 ( .A(n235), .B(n236), .Z(n233) );
  NAND U207 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U208 ( .A(A[197]), .B(B[197]), .Z(n238) );
  AND U209 ( .A(n239), .B(n240), .Z(n237) );
  NANDN U210 ( .A(A[196]), .B(B[196]), .Z(n240) );
  NAND U211 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U212 ( .A(B[196]), .B(A[196]), .Z(n242) );
  AND U213 ( .A(n243), .B(n244), .Z(n241) );
  NAND U214 ( .A(n245), .B(n246), .Z(n244) );
  NANDN U215 ( .A(A[195]), .B(B[195]), .Z(n246) );
  AND U216 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U217 ( .A(A[194]), .B(B[194]), .Z(n248) );
  NAND U218 ( .A(n249), .B(n250), .Z(n247) );
  NANDN U219 ( .A(B[194]), .B(A[194]), .Z(n250) );
  AND U220 ( .A(n251), .B(n252), .Z(n249) );
  NAND U221 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U222 ( .A(A[193]), .B(B[193]), .Z(n254) );
  AND U223 ( .A(n255), .B(n256), .Z(n253) );
  NANDN U224 ( .A(A[192]), .B(B[192]), .Z(n256) );
  NAND U225 ( .A(n257), .B(n258), .Z(n255) );
  NANDN U226 ( .A(B[192]), .B(A[192]), .Z(n258) );
  AND U227 ( .A(n259), .B(n260), .Z(n257) );
  NAND U228 ( .A(n261), .B(n262), .Z(n260) );
  NANDN U229 ( .A(A[191]), .B(B[191]), .Z(n262) );
  AND U230 ( .A(n263), .B(n264), .Z(n261) );
  NANDN U231 ( .A(A[190]), .B(B[190]), .Z(n264) );
  NAND U232 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U233 ( .A(B[190]), .B(A[190]), .Z(n266) );
  AND U234 ( .A(n267), .B(n268), .Z(n265) );
  NAND U235 ( .A(n269), .B(n270), .Z(n268) );
  NANDN U236 ( .A(A[189]), .B(B[189]), .Z(n270) );
  AND U237 ( .A(n271), .B(n272), .Z(n269) );
  NANDN U238 ( .A(A[188]), .B(B[188]), .Z(n272) );
  NAND U239 ( .A(n273), .B(n274), .Z(n271) );
  NANDN U240 ( .A(B[188]), .B(A[188]), .Z(n274) );
  AND U241 ( .A(n275), .B(n276), .Z(n273) );
  NAND U242 ( .A(n277), .B(n278), .Z(n276) );
  NANDN U243 ( .A(A[187]), .B(B[187]), .Z(n278) );
  AND U244 ( .A(n279), .B(n280), .Z(n277) );
  NANDN U245 ( .A(A[186]), .B(B[186]), .Z(n280) );
  NAND U246 ( .A(n281), .B(n282), .Z(n279) );
  NANDN U247 ( .A(B[186]), .B(A[186]), .Z(n282) );
  AND U248 ( .A(n283), .B(n284), .Z(n281) );
  NAND U249 ( .A(n285), .B(n286), .Z(n284) );
  NANDN U250 ( .A(A[185]), .B(B[185]), .Z(n286) );
  AND U251 ( .A(n287), .B(n288), .Z(n285) );
  NANDN U252 ( .A(A[184]), .B(B[184]), .Z(n288) );
  NAND U253 ( .A(n289), .B(n290), .Z(n287) );
  NANDN U254 ( .A(B[184]), .B(A[184]), .Z(n290) );
  AND U255 ( .A(n291), .B(n292), .Z(n289) );
  NAND U256 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U257 ( .A(A[183]), .B(B[183]), .Z(n294) );
  AND U258 ( .A(n295), .B(n296), .Z(n293) );
  NANDN U259 ( .A(A[182]), .B(B[182]), .Z(n296) );
  NAND U260 ( .A(n297), .B(n298), .Z(n295) );
  NANDN U261 ( .A(B[182]), .B(A[182]), .Z(n298) );
  AND U262 ( .A(n299), .B(n300), .Z(n297) );
  NAND U263 ( .A(n301), .B(n302), .Z(n300) );
  NANDN U264 ( .A(A[181]), .B(B[181]), .Z(n302) );
  AND U265 ( .A(n303), .B(n304), .Z(n301) );
  NANDN U266 ( .A(A[180]), .B(B[180]), .Z(n304) );
  NAND U267 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U268 ( .A(B[180]), .B(A[180]), .Z(n306) );
  AND U269 ( .A(n307), .B(n308), .Z(n305) );
  NAND U270 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U271 ( .A(A[179]), .B(B[179]), .Z(n310) );
  AND U272 ( .A(n311), .B(n312), .Z(n309) );
  NANDN U273 ( .A(A[178]), .B(B[178]), .Z(n312) );
  NAND U274 ( .A(n313), .B(n314), .Z(n311) );
  NANDN U275 ( .A(B[178]), .B(A[178]), .Z(n314) );
  AND U276 ( .A(n315), .B(n316), .Z(n313) );
  NAND U277 ( .A(n317), .B(n318), .Z(n316) );
  NANDN U278 ( .A(A[177]), .B(B[177]), .Z(n318) );
  AND U279 ( .A(n319), .B(n320), .Z(n317) );
  NANDN U280 ( .A(A[176]), .B(B[176]), .Z(n320) );
  NAND U281 ( .A(n321), .B(n322), .Z(n319) );
  NANDN U282 ( .A(B[176]), .B(A[176]), .Z(n322) );
  AND U283 ( .A(n323), .B(n324), .Z(n321) );
  NAND U284 ( .A(n325), .B(n326), .Z(n324) );
  NANDN U285 ( .A(A[175]), .B(B[175]), .Z(n326) );
  AND U286 ( .A(n327), .B(n328), .Z(n325) );
  NANDN U287 ( .A(A[174]), .B(B[174]), .Z(n328) );
  NAND U288 ( .A(n329), .B(n330), .Z(n327) );
  NANDN U289 ( .A(B[174]), .B(A[174]), .Z(n330) );
  AND U290 ( .A(n331), .B(n332), .Z(n329) );
  NAND U291 ( .A(n333), .B(n334), .Z(n332) );
  NANDN U292 ( .A(A[173]), .B(B[173]), .Z(n334) );
  AND U293 ( .A(n335), .B(n336), .Z(n333) );
  NANDN U294 ( .A(A[172]), .B(B[172]), .Z(n336) );
  NAND U295 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U296 ( .A(B[172]), .B(A[172]), .Z(n338) );
  AND U297 ( .A(n339), .B(n340), .Z(n337) );
  NAND U298 ( .A(n341), .B(n342), .Z(n340) );
  NANDN U299 ( .A(A[171]), .B(B[171]), .Z(n342) );
  AND U300 ( .A(n343), .B(n344), .Z(n341) );
  NANDN U301 ( .A(A[170]), .B(B[170]), .Z(n344) );
  NAND U302 ( .A(n345), .B(n346), .Z(n343) );
  NANDN U303 ( .A(B[170]), .B(A[170]), .Z(n346) );
  AND U304 ( .A(n347), .B(n348), .Z(n345) );
  NAND U305 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U306 ( .A(A[169]), .B(B[169]), .Z(n350) );
  AND U307 ( .A(n351), .B(n352), .Z(n349) );
  NANDN U308 ( .A(A[168]), .B(B[168]), .Z(n352) );
  NAND U309 ( .A(n353), .B(n354), .Z(n351) );
  NANDN U310 ( .A(B[168]), .B(A[168]), .Z(n354) );
  AND U311 ( .A(n355), .B(n356), .Z(n353) );
  NAND U312 ( .A(n357), .B(n358), .Z(n356) );
  NANDN U313 ( .A(A[167]), .B(B[167]), .Z(n358) );
  AND U314 ( .A(n359), .B(n360), .Z(n357) );
  NANDN U315 ( .A(A[166]), .B(B[166]), .Z(n360) );
  NAND U316 ( .A(n361), .B(n362), .Z(n359) );
  NANDN U317 ( .A(B[166]), .B(A[166]), .Z(n362) );
  AND U318 ( .A(n363), .B(n364), .Z(n361) );
  NAND U319 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U320 ( .A(A[165]), .B(B[165]), .Z(n366) );
  AND U321 ( .A(n367), .B(n368), .Z(n365) );
  NANDN U322 ( .A(A[164]), .B(B[164]), .Z(n368) );
  NAND U323 ( .A(n369), .B(n370), .Z(n367) );
  NANDN U324 ( .A(B[164]), .B(A[164]), .Z(n370) );
  AND U325 ( .A(n371), .B(n372), .Z(n369) );
  NAND U326 ( .A(n373), .B(n374), .Z(n372) );
  NANDN U327 ( .A(A[163]), .B(B[163]), .Z(n374) );
  AND U328 ( .A(n375), .B(n376), .Z(n373) );
  NANDN U329 ( .A(A[162]), .B(B[162]), .Z(n376) );
  NAND U330 ( .A(n377), .B(n378), .Z(n375) );
  NANDN U331 ( .A(B[162]), .B(A[162]), .Z(n378) );
  AND U332 ( .A(n379), .B(n380), .Z(n377) );
  NAND U333 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U334 ( .A(A[161]), .B(B[161]), .Z(n382) );
  AND U335 ( .A(n383), .B(n384), .Z(n381) );
  NANDN U336 ( .A(A[160]), .B(B[160]), .Z(n384) );
  NAND U337 ( .A(n385), .B(n386), .Z(n383) );
  NANDN U338 ( .A(B[160]), .B(A[160]), .Z(n386) );
  AND U339 ( .A(n387), .B(n388), .Z(n385) );
  NAND U340 ( .A(n389), .B(n390), .Z(n388) );
  NANDN U341 ( .A(A[159]), .B(B[159]), .Z(n390) );
  AND U342 ( .A(n391), .B(n392), .Z(n389) );
  NANDN U343 ( .A(A[158]), .B(B[158]), .Z(n392) );
  NAND U344 ( .A(n393), .B(n394), .Z(n391) );
  NANDN U345 ( .A(B[158]), .B(A[158]), .Z(n394) );
  AND U346 ( .A(n395), .B(n396), .Z(n393) );
  NAND U347 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U348 ( .A(A[157]), .B(B[157]), .Z(n398) );
  AND U349 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U350 ( .A(A[156]), .B(B[156]), .Z(n400) );
  NAND U351 ( .A(n401), .B(n402), .Z(n399) );
  NANDN U352 ( .A(B[156]), .B(A[156]), .Z(n402) );
  AND U353 ( .A(n403), .B(n404), .Z(n401) );
  NAND U354 ( .A(n405), .B(n406), .Z(n404) );
  NANDN U355 ( .A(A[155]), .B(B[155]), .Z(n406) );
  AND U356 ( .A(n407), .B(n408), .Z(n405) );
  NANDN U357 ( .A(A[154]), .B(B[154]), .Z(n408) );
  NAND U358 ( .A(n409), .B(n410), .Z(n407) );
  NANDN U359 ( .A(B[154]), .B(A[154]), .Z(n410) );
  AND U360 ( .A(n411), .B(n412), .Z(n409) );
  NAND U361 ( .A(n413), .B(n414), .Z(n412) );
  NANDN U362 ( .A(A[153]), .B(B[153]), .Z(n414) );
  AND U363 ( .A(n415), .B(n416), .Z(n413) );
  NANDN U364 ( .A(A[152]), .B(B[152]), .Z(n416) );
  NAND U365 ( .A(n417), .B(n418), .Z(n415) );
  NANDN U366 ( .A(B[152]), .B(A[152]), .Z(n418) );
  AND U367 ( .A(n419), .B(n420), .Z(n417) );
  NAND U368 ( .A(n421), .B(n422), .Z(n420) );
  NANDN U369 ( .A(A[151]), .B(B[151]), .Z(n422) );
  AND U370 ( .A(n423), .B(n424), .Z(n421) );
  NANDN U371 ( .A(A[150]), .B(B[150]), .Z(n424) );
  NAND U372 ( .A(n425), .B(n426), .Z(n423) );
  NANDN U373 ( .A(B[150]), .B(A[150]), .Z(n426) );
  AND U374 ( .A(n427), .B(n428), .Z(n425) );
  NAND U375 ( .A(n429), .B(n430), .Z(n428) );
  NANDN U376 ( .A(A[149]), .B(B[149]), .Z(n430) );
  AND U377 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U378 ( .A(A[148]), .B(B[148]), .Z(n432) );
  NAND U379 ( .A(n433), .B(n434), .Z(n431) );
  NANDN U380 ( .A(B[148]), .B(A[148]), .Z(n434) );
  AND U381 ( .A(n435), .B(n436), .Z(n433) );
  NAND U382 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U383 ( .A(A[147]), .B(B[147]), .Z(n438) );
  AND U384 ( .A(n439), .B(n440), .Z(n437) );
  NANDN U385 ( .A(A[146]), .B(B[146]), .Z(n440) );
  NAND U386 ( .A(n441), .B(n442), .Z(n439) );
  NANDN U387 ( .A(B[146]), .B(A[146]), .Z(n442) );
  AND U388 ( .A(n443), .B(n444), .Z(n441) );
  NAND U389 ( .A(n445), .B(n446), .Z(n444) );
  NANDN U390 ( .A(A[145]), .B(B[145]), .Z(n446) );
  AND U391 ( .A(n447), .B(n448), .Z(n445) );
  NANDN U392 ( .A(A[144]), .B(B[144]), .Z(n448) );
  NAND U393 ( .A(n449), .B(n450), .Z(n447) );
  NANDN U394 ( .A(B[144]), .B(A[144]), .Z(n450) );
  AND U395 ( .A(n451), .B(n452), .Z(n449) );
  NAND U396 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U397 ( .A(A[143]), .B(B[143]), .Z(n454) );
  AND U398 ( .A(n455), .B(n456), .Z(n453) );
  NANDN U399 ( .A(A[142]), .B(B[142]), .Z(n456) );
  NAND U400 ( .A(n457), .B(n458), .Z(n455) );
  NANDN U401 ( .A(B[142]), .B(A[142]), .Z(n458) );
  AND U402 ( .A(n459), .B(n460), .Z(n457) );
  NAND U403 ( .A(n461), .B(n462), .Z(n460) );
  NANDN U404 ( .A(A[141]), .B(B[141]), .Z(n462) );
  AND U405 ( .A(n463), .B(n464), .Z(n461) );
  NANDN U406 ( .A(A[140]), .B(B[140]), .Z(n464) );
  NAND U407 ( .A(n465), .B(n466), .Z(n463) );
  NANDN U408 ( .A(B[140]), .B(A[140]), .Z(n466) );
  AND U409 ( .A(n467), .B(n468), .Z(n465) );
  NAND U410 ( .A(n469), .B(n470), .Z(n468) );
  NANDN U411 ( .A(A[139]), .B(B[139]), .Z(n470) );
  AND U412 ( .A(n471), .B(n472), .Z(n469) );
  NANDN U413 ( .A(A[138]), .B(B[138]), .Z(n472) );
  NAND U414 ( .A(n473), .B(n474), .Z(n471) );
  NANDN U415 ( .A(B[138]), .B(A[138]), .Z(n474) );
  AND U416 ( .A(n475), .B(n476), .Z(n473) );
  NAND U417 ( .A(n477), .B(n478), .Z(n476) );
  NANDN U418 ( .A(A[137]), .B(B[137]), .Z(n478) );
  AND U419 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U420 ( .A(A[136]), .B(B[136]), .Z(n480) );
  NAND U421 ( .A(n481), .B(n482), .Z(n479) );
  NANDN U422 ( .A(B[136]), .B(A[136]), .Z(n482) );
  AND U423 ( .A(n483), .B(n484), .Z(n481) );
  NAND U424 ( .A(n485), .B(n486), .Z(n484) );
  NANDN U425 ( .A(A[135]), .B(B[135]), .Z(n486) );
  AND U426 ( .A(n487), .B(n488), .Z(n485) );
  NANDN U427 ( .A(A[134]), .B(B[134]), .Z(n488) );
  NAND U428 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U429 ( .A(B[134]), .B(A[134]), .Z(n490) );
  AND U430 ( .A(n491), .B(n492), .Z(n489) );
  NAND U431 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U432 ( .A(A[133]), .B(B[133]), .Z(n494) );
  AND U433 ( .A(n495), .B(n496), .Z(n493) );
  NANDN U434 ( .A(A[132]), .B(B[132]), .Z(n496) );
  NAND U435 ( .A(n497), .B(n498), .Z(n495) );
  NANDN U436 ( .A(B[132]), .B(A[132]), .Z(n498) );
  AND U437 ( .A(n499), .B(n500), .Z(n497) );
  NAND U438 ( .A(n501), .B(n502), .Z(n500) );
  NANDN U439 ( .A(A[131]), .B(B[131]), .Z(n502) );
  AND U440 ( .A(n503), .B(n504), .Z(n501) );
  NANDN U441 ( .A(A[130]), .B(B[130]), .Z(n504) );
  NAND U442 ( .A(n505), .B(n506), .Z(n503) );
  NANDN U443 ( .A(B[130]), .B(A[130]), .Z(n506) );
  AND U444 ( .A(n507), .B(n508), .Z(n505) );
  NAND U445 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U446 ( .A(A[129]), .B(B[129]), .Z(n510) );
  AND U447 ( .A(n511), .B(n512), .Z(n509) );
  NANDN U448 ( .A(A[128]), .B(B[128]), .Z(n512) );
  NAND U449 ( .A(n513), .B(n514), .Z(n511) );
  NANDN U450 ( .A(B[128]), .B(A[128]), .Z(n514) );
  AND U451 ( .A(n515), .B(n516), .Z(n513) );
  NAND U452 ( .A(n517), .B(n518), .Z(n516) );
  NANDN U453 ( .A(A[127]), .B(B[127]), .Z(n518) );
  AND U454 ( .A(n519), .B(n520), .Z(n517) );
  NANDN U455 ( .A(A[126]), .B(B[126]), .Z(n520) );
  NAND U456 ( .A(n521), .B(n522), .Z(n519) );
  NANDN U457 ( .A(B[126]), .B(A[126]), .Z(n522) );
  AND U458 ( .A(n523), .B(n524), .Z(n521) );
  NAND U459 ( .A(n525), .B(n526), .Z(n524) );
  NANDN U460 ( .A(A[125]), .B(B[125]), .Z(n526) );
  AND U461 ( .A(n527), .B(n528), .Z(n525) );
  NANDN U462 ( .A(A[124]), .B(B[124]), .Z(n528) );
  NAND U463 ( .A(n529), .B(n530), .Z(n527) );
  NANDN U464 ( .A(B[124]), .B(A[124]), .Z(n530) );
  AND U465 ( .A(n531), .B(n532), .Z(n529) );
  NAND U466 ( .A(n533), .B(n534), .Z(n532) );
  NANDN U467 ( .A(A[123]), .B(B[123]), .Z(n534) );
  AND U468 ( .A(n535), .B(n536), .Z(n533) );
  NANDN U469 ( .A(A[122]), .B(B[122]), .Z(n536) );
  NAND U470 ( .A(n537), .B(n538), .Z(n535) );
  NANDN U471 ( .A(B[122]), .B(A[122]), .Z(n538) );
  AND U472 ( .A(n539), .B(n540), .Z(n537) );
  NAND U473 ( .A(n541), .B(n542), .Z(n540) );
  NANDN U474 ( .A(A[121]), .B(B[121]), .Z(n542) );
  AND U475 ( .A(n543), .B(n544), .Z(n541) );
  NANDN U476 ( .A(A[120]), .B(B[120]), .Z(n544) );
  NAND U477 ( .A(n545), .B(n546), .Z(n543) );
  NANDN U478 ( .A(B[120]), .B(A[120]), .Z(n546) );
  AND U479 ( .A(n547), .B(n548), .Z(n545) );
  NAND U480 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U481 ( .A(A[119]), .B(B[119]), .Z(n550) );
  AND U482 ( .A(n551), .B(n552), .Z(n549) );
  NANDN U483 ( .A(A[118]), .B(B[118]), .Z(n552) );
  NAND U484 ( .A(n553), .B(n554), .Z(n551) );
  NANDN U485 ( .A(B[118]), .B(A[118]), .Z(n554) );
  AND U486 ( .A(n555), .B(n556), .Z(n553) );
  NAND U487 ( .A(n557), .B(n558), .Z(n556) );
  NANDN U488 ( .A(A[117]), .B(B[117]), .Z(n558) );
  AND U489 ( .A(n559), .B(n560), .Z(n557) );
  NANDN U490 ( .A(A[116]), .B(B[116]), .Z(n560) );
  NAND U491 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U492 ( .A(B[116]), .B(A[116]), .Z(n562) );
  AND U493 ( .A(n563), .B(n564), .Z(n561) );
  NAND U494 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U495 ( .A(A[115]), .B(B[115]), .Z(n566) );
  AND U496 ( .A(n567), .B(n568), .Z(n565) );
  NANDN U497 ( .A(A[114]), .B(B[114]), .Z(n568) );
  NAND U498 ( .A(n569), .B(n570), .Z(n567) );
  NANDN U499 ( .A(B[114]), .B(A[114]), .Z(n570) );
  AND U500 ( .A(n571), .B(n572), .Z(n569) );
  NAND U501 ( .A(n573), .B(n574), .Z(n572) );
  NANDN U502 ( .A(A[113]), .B(B[113]), .Z(n574) );
  AND U503 ( .A(n575), .B(n576), .Z(n573) );
  NANDN U504 ( .A(A[112]), .B(B[112]), .Z(n576) );
  NAND U505 ( .A(n577), .B(n578), .Z(n575) );
  NANDN U506 ( .A(B[112]), .B(A[112]), .Z(n578) );
  AND U507 ( .A(n579), .B(n580), .Z(n577) );
  NAND U508 ( .A(n581), .B(n582), .Z(n580) );
  NANDN U509 ( .A(A[111]), .B(B[111]), .Z(n582) );
  AND U510 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U511 ( .A(A[110]), .B(B[110]), .Z(n584) );
  NAND U512 ( .A(n585), .B(n586), .Z(n583) );
  NANDN U513 ( .A(B[110]), .B(A[110]), .Z(n586) );
  AND U514 ( .A(n587), .B(n588), .Z(n585) );
  NAND U515 ( .A(n589), .B(n590), .Z(n588) );
  NANDN U516 ( .A(A[109]), .B(B[109]), .Z(n590) );
  AND U517 ( .A(n591), .B(n592), .Z(n589) );
  NANDN U518 ( .A(A[108]), .B(B[108]), .Z(n592) );
  NAND U519 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U520 ( .A(B[108]), .B(A[108]), .Z(n594) );
  AND U521 ( .A(n595), .B(n596), .Z(n593) );
  NAND U522 ( .A(n597), .B(n598), .Z(n596) );
  NANDN U523 ( .A(A[107]), .B(B[107]), .Z(n598) );
  AND U524 ( .A(n599), .B(n600), .Z(n597) );
  NANDN U525 ( .A(A[106]), .B(B[106]), .Z(n600) );
  NAND U526 ( .A(n601), .B(n602), .Z(n599) );
  NANDN U527 ( .A(B[106]), .B(A[106]), .Z(n602) );
  AND U528 ( .A(n603), .B(n604), .Z(n601) );
  NAND U529 ( .A(n605), .B(n606), .Z(n604) );
  NANDN U530 ( .A(A[105]), .B(B[105]), .Z(n606) );
  AND U531 ( .A(n607), .B(n608), .Z(n605) );
  NANDN U532 ( .A(A[104]), .B(B[104]), .Z(n608) );
  NAND U533 ( .A(n609), .B(n610), .Z(n607) );
  NANDN U534 ( .A(B[104]), .B(A[104]), .Z(n610) );
  AND U535 ( .A(n611), .B(n612), .Z(n609) );
  NAND U536 ( .A(n613), .B(n614), .Z(n612) );
  NANDN U537 ( .A(A[103]), .B(B[103]), .Z(n614) );
  AND U538 ( .A(n615), .B(n616), .Z(n613) );
  NANDN U539 ( .A(A[102]), .B(B[102]), .Z(n616) );
  NAND U540 ( .A(n617), .B(n618), .Z(n615) );
  NANDN U541 ( .A(B[102]), .B(A[102]), .Z(n618) );
  AND U542 ( .A(n619), .B(n620), .Z(n617) );
  NAND U543 ( .A(n621), .B(n622), .Z(n620) );
  NANDN U544 ( .A(A[101]), .B(B[101]), .Z(n622) );
  AND U545 ( .A(n623), .B(n624), .Z(n621) );
  NANDN U546 ( .A(A[100]), .B(B[100]), .Z(n624) );
  NAND U547 ( .A(n625), .B(n626), .Z(n623) );
  NANDN U548 ( .A(B[99]), .B(A[99]), .Z(n626) );
  AND U549 ( .A(n627), .B(n628), .Z(n625) );
  NAND U550 ( .A(n629), .B(n630), .Z(n628) );
  NANDN U551 ( .A(A[99]), .B(B[99]), .Z(n630) );
  AND U552 ( .A(n631), .B(n632), .Z(n629) );
  NANDN U553 ( .A(A[98]), .B(B[98]), .Z(n632) );
  NAND U554 ( .A(n633), .B(n634), .Z(n631) );
  NANDN U555 ( .A(B[98]), .B(A[98]), .Z(n634) );
  AND U556 ( .A(n635), .B(n636), .Z(n633) );
  NAND U557 ( .A(n637), .B(n638), .Z(n636) );
  NANDN U558 ( .A(A[97]), .B(B[97]), .Z(n638) );
  AND U559 ( .A(n639), .B(n640), .Z(n637) );
  NANDN U560 ( .A(A[96]), .B(B[96]), .Z(n640) );
  NAND U561 ( .A(n641), .B(n642), .Z(n639) );
  NANDN U562 ( .A(B[96]), .B(A[96]), .Z(n642) );
  AND U563 ( .A(n643), .B(n644), .Z(n641) );
  NAND U564 ( .A(n645), .B(n646), .Z(n644) );
  NANDN U565 ( .A(A[95]), .B(B[95]), .Z(n646) );
  AND U566 ( .A(n647), .B(n648), .Z(n645) );
  NANDN U567 ( .A(A[94]), .B(B[94]), .Z(n648) );
  NAND U568 ( .A(n649), .B(n650), .Z(n647) );
  NANDN U569 ( .A(B[94]), .B(A[94]), .Z(n650) );
  AND U570 ( .A(n651), .B(n652), .Z(n649) );
  NAND U571 ( .A(n653), .B(n654), .Z(n652) );
  NANDN U572 ( .A(A[93]), .B(B[93]), .Z(n654) );
  AND U573 ( .A(n655), .B(n656), .Z(n653) );
  NANDN U574 ( .A(A[92]), .B(B[92]), .Z(n656) );
  NAND U575 ( .A(n657), .B(n658), .Z(n655) );
  NANDN U576 ( .A(B[92]), .B(A[92]), .Z(n658) );
  AND U577 ( .A(n659), .B(n660), .Z(n657) );
  NAND U578 ( .A(n661), .B(n662), .Z(n660) );
  NANDN U579 ( .A(A[91]), .B(B[91]), .Z(n662) );
  AND U580 ( .A(n663), .B(n664), .Z(n661) );
  NANDN U581 ( .A(A[90]), .B(B[90]), .Z(n664) );
  NAND U582 ( .A(n665), .B(n666), .Z(n663) );
  NANDN U583 ( .A(B[90]), .B(A[90]), .Z(n666) );
  AND U584 ( .A(n667), .B(n668), .Z(n665) );
  NAND U585 ( .A(n669), .B(n670), .Z(n668) );
  NANDN U586 ( .A(A[89]), .B(B[89]), .Z(n670) );
  AND U587 ( .A(n671), .B(n672), .Z(n669) );
  NANDN U588 ( .A(A[88]), .B(B[88]), .Z(n672) );
  NAND U589 ( .A(n673), .B(n674), .Z(n671) );
  NANDN U590 ( .A(B[88]), .B(A[88]), .Z(n674) );
  AND U591 ( .A(n675), .B(n676), .Z(n673) );
  NAND U592 ( .A(n677), .B(n678), .Z(n676) );
  NANDN U593 ( .A(A[87]), .B(B[87]), .Z(n678) );
  AND U594 ( .A(n679), .B(n680), .Z(n677) );
  NANDN U595 ( .A(A[86]), .B(B[86]), .Z(n680) );
  NAND U596 ( .A(n681), .B(n682), .Z(n679) );
  NANDN U597 ( .A(B[86]), .B(A[86]), .Z(n682) );
  AND U598 ( .A(n683), .B(n684), .Z(n681) );
  NAND U599 ( .A(n685), .B(n686), .Z(n684) );
  NANDN U600 ( .A(A[85]), .B(B[85]), .Z(n686) );
  AND U601 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U602 ( .A(A[84]), .B(B[84]), .Z(n688) );
  NAND U603 ( .A(n689), .B(n690), .Z(n687) );
  NANDN U604 ( .A(B[84]), .B(A[84]), .Z(n690) );
  AND U605 ( .A(n691), .B(n692), .Z(n689) );
  NAND U606 ( .A(n693), .B(n694), .Z(n692) );
  NANDN U607 ( .A(A[83]), .B(B[83]), .Z(n694) );
  AND U608 ( .A(n695), .B(n696), .Z(n693) );
  NANDN U609 ( .A(A[82]), .B(B[82]), .Z(n696) );
  NAND U610 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U611 ( .A(B[82]), .B(A[82]), .Z(n698) );
  AND U612 ( .A(n699), .B(n700), .Z(n697) );
  NAND U613 ( .A(n701), .B(n702), .Z(n700) );
  NANDN U614 ( .A(A[81]), .B(B[81]), .Z(n702) );
  AND U615 ( .A(n703), .B(n704), .Z(n701) );
  NANDN U616 ( .A(A[80]), .B(B[80]), .Z(n704) );
  NAND U617 ( .A(n705), .B(n706), .Z(n703) );
  NANDN U618 ( .A(B[80]), .B(A[80]), .Z(n706) );
  AND U619 ( .A(n707), .B(n708), .Z(n705) );
  NAND U620 ( .A(n709), .B(n710), .Z(n708) );
  NANDN U621 ( .A(A[79]), .B(B[79]), .Z(n710) );
  AND U622 ( .A(n711), .B(n712), .Z(n709) );
  NANDN U623 ( .A(A[78]), .B(B[78]), .Z(n712) );
  NAND U624 ( .A(n713), .B(n714), .Z(n711) );
  NANDN U625 ( .A(B[78]), .B(A[78]), .Z(n714) );
  AND U626 ( .A(n715), .B(n716), .Z(n713) );
  NAND U627 ( .A(n717), .B(n718), .Z(n716) );
  NANDN U628 ( .A(A[77]), .B(B[77]), .Z(n718) );
  AND U629 ( .A(n719), .B(n720), .Z(n717) );
  NANDN U630 ( .A(A[76]), .B(B[76]), .Z(n720) );
  NAND U631 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U632 ( .A(B[76]), .B(A[76]), .Z(n722) );
  AND U633 ( .A(n723), .B(n724), .Z(n721) );
  NAND U634 ( .A(n725), .B(n726), .Z(n724) );
  NANDN U635 ( .A(A[75]), .B(B[75]), .Z(n726) );
  AND U636 ( .A(n727), .B(n728), .Z(n725) );
  NANDN U637 ( .A(A[74]), .B(B[74]), .Z(n728) );
  NAND U638 ( .A(n729), .B(n730), .Z(n727) );
  NANDN U639 ( .A(B[74]), .B(A[74]), .Z(n730) );
  AND U640 ( .A(n731), .B(n732), .Z(n729) );
  NAND U641 ( .A(n733), .B(n734), .Z(n732) );
  NANDN U642 ( .A(A[73]), .B(B[73]), .Z(n734) );
  AND U643 ( .A(n735), .B(n736), .Z(n733) );
  NANDN U644 ( .A(A[72]), .B(B[72]), .Z(n736) );
  NAND U645 ( .A(n737), .B(n738), .Z(n735) );
  NANDN U646 ( .A(B[72]), .B(A[72]), .Z(n738) );
  AND U647 ( .A(n739), .B(n740), .Z(n737) );
  NAND U648 ( .A(n741), .B(n742), .Z(n740) );
  NANDN U649 ( .A(A[71]), .B(B[71]), .Z(n742) );
  AND U650 ( .A(n743), .B(n744), .Z(n741) );
  NANDN U651 ( .A(A[70]), .B(B[70]), .Z(n744) );
  NAND U652 ( .A(n745), .B(n746), .Z(n743) );
  NANDN U653 ( .A(B[70]), .B(A[70]), .Z(n746) );
  AND U654 ( .A(n747), .B(n748), .Z(n745) );
  NAND U655 ( .A(n749), .B(n750), .Z(n748) );
  NANDN U656 ( .A(A[69]), .B(B[69]), .Z(n750) );
  AND U657 ( .A(n751), .B(n752), .Z(n749) );
  NANDN U658 ( .A(A[68]), .B(B[68]), .Z(n752) );
  NAND U659 ( .A(n753), .B(n754), .Z(n751) );
  NANDN U660 ( .A(B[68]), .B(A[68]), .Z(n754) );
  AND U661 ( .A(n755), .B(n756), .Z(n753) );
  NAND U662 ( .A(n757), .B(n758), .Z(n756) );
  NANDN U663 ( .A(A[67]), .B(B[67]), .Z(n758) );
  AND U664 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U665 ( .A(A[66]), .B(B[66]), .Z(n760) );
  NAND U666 ( .A(n761), .B(n762), .Z(n759) );
  NANDN U667 ( .A(B[66]), .B(A[66]), .Z(n762) );
  AND U668 ( .A(n763), .B(n764), .Z(n761) );
  NAND U669 ( .A(n765), .B(n766), .Z(n764) );
  NANDN U670 ( .A(A[65]), .B(B[65]), .Z(n766) );
  AND U671 ( .A(n767), .B(n768), .Z(n765) );
  NANDN U672 ( .A(A[64]), .B(B[64]), .Z(n768) );
  NAND U673 ( .A(n769), .B(n770), .Z(n767) );
  NANDN U674 ( .A(B[64]), .B(A[64]), .Z(n770) );
  AND U675 ( .A(n771), .B(n772), .Z(n769) );
  NAND U676 ( .A(n773), .B(n774), .Z(n772) );
  NANDN U677 ( .A(A[63]), .B(B[63]), .Z(n774) );
  AND U678 ( .A(n775), .B(n776), .Z(n773) );
  NANDN U679 ( .A(A[62]), .B(B[62]), .Z(n776) );
  NAND U680 ( .A(n777), .B(n778), .Z(n775) );
  NANDN U681 ( .A(B[62]), .B(A[62]), .Z(n778) );
  AND U682 ( .A(n779), .B(n780), .Z(n777) );
  NAND U683 ( .A(n781), .B(n782), .Z(n780) );
  NANDN U684 ( .A(A[61]), .B(B[61]), .Z(n782) );
  AND U685 ( .A(n783), .B(n784), .Z(n781) );
  NANDN U686 ( .A(A[60]), .B(B[60]), .Z(n784) );
  NAND U687 ( .A(n785), .B(n786), .Z(n783) );
  NANDN U688 ( .A(B[60]), .B(A[60]), .Z(n786) );
  AND U689 ( .A(n787), .B(n788), .Z(n785) );
  NAND U690 ( .A(n789), .B(n790), .Z(n788) );
  NANDN U691 ( .A(A[59]), .B(B[59]), .Z(n790) );
  AND U692 ( .A(n791), .B(n792), .Z(n789) );
  NANDN U693 ( .A(A[58]), .B(B[58]), .Z(n792) );
  NAND U694 ( .A(n793), .B(n794), .Z(n791) );
  NANDN U695 ( .A(B[58]), .B(A[58]), .Z(n794) );
  AND U696 ( .A(n795), .B(n796), .Z(n793) );
  NAND U697 ( .A(n797), .B(n798), .Z(n796) );
  NANDN U698 ( .A(A[57]), .B(B[57]), .Z(n798) );
  AND U699 ( .A(n799), .B(n800), .Z(n797) );
  NANDN U700 ( .A(A[56]), .B(B[56]), .Z(n800) );
  NAND U701 ( .A(n801), .B(n802), .Z(n799) );
  NANDN U702 ( .A(B[56]), .B(A[56]), .Z(n802) );
  AND U703 ( .A(n803), .B(n804), .Z(n801) );
  NAND U704 ( .A(n805), .B(n806), .Z(n804) );
  NANDN U705 ( .A(A[55]), .B(B[55]), .Z(n806) );
  AND U706 ( .A(n807), .B(n808), .Z(n805) );
  NANDN U707 ( .A(A[54]), .B(B[54]), .Z(n808) );
  NAND U708 ( .A(n809), .B(n810), .Z(n807) );
  NANDN U709 ( .A(B[54]), .B(A[54]), .Z(n810) );
  AND U710 ( .A(n811), .B(n812), .Z(n809) );
  NAND U711 ( .A(n813), .B(n814), .Z(n812) );
  NANDN U712 ( .A(A[53]), .B(B[53]), .Z(n814) );
  AND U713 ( .A(n815), .B(n816), .Z(n813) );
  NANDN U714 ( .A(A[52]), .B(B[52]), .Z(n816) );
  NAND U715 ( .A(n817), .B(n818), .Z(n815) );
  NANDN U716 ( .A(B[52]), .B(A[52]), .Z(n818) );
  AND U717 ( .A(n819), .B(n820), .Z(n817) );
  NAND U718 ( .A(n821), .B(n822), .Z(n820) );
  NANDN U719 ( .A(A[51]), .B(B[51]), .Z(n822) );
  AND U720 ( .A(n823), .B(n824), .Z(n821) );
  NANDN U721 ( .A(A[50]), .B(B[50]), .Z(n824) );
  NAND U722 ( .A(n825), .B(n826), .Z(n823) );
  NANDN U723 ( .A(B[50]), .B(A[50]), .Z(n826) );
  AND U724 ( .A(n827), .B(n828), .Z(n825) );
  NAND U725 ( .A(n829), .B(n830), .Z(n828) );
  NANDN U726 ( .A(A[49]), .B(B[49]), .Z(n830) );
  AND U727 ( .A(n831), .B(n832), .Z(n829) );
  NANDN U728 ( .A(A[48]), .B(B[48]), .Z(n832) );
  NAND U729 ( .A(n833), .B(n834), .Z(n831) );
  NANDN U730 ( .A(B[48]), .B(A[48]), .Z(n834) );
  AND U731 ( .A(n835), .B(n836), .Z(n833) );
  NAND U732 ( .A(n837), .B(n838), .Z(n836) );
  NANDN U733 ( .A(A[47]), .B(B[47]), .Z(n838) );
  AND U734 ( .A(n839), .B(n840), .Z(n837) );
  NANDN U735 ( .A(A[46]), .B(B[46]), .Z(n840) );
  NAND U736 ( .A(n841), .B(n842), .Z(n839) );
  NANDN U737 ( .A(B[46]), .B(A[46]), .Z(n842) );
  AND U738 ( .A(n843), .B(n844), .Z(n841) );
  NAND U739 ( .A(n845), .B(n846), .Z(n844) );
  NANDN U740 ( .A(A[45]), .B(B[45]), .Z(n846) );
  AND U741 ( .A(n847), .B(n848), .Z(n845) );
  NANDN U742 ( .A(A[44]), .B(B[44]), .Z(n848) );
  NAND U743 ( .A(n849), .B(n850), .Z(n847) );
  NANDN U744 ( .A(B[44]), .B(A[44]), .Z(n850) );
  AND U745 ( .A(n851), .B(n852), .Z(n849) );
  NAND U746 ( .A(n853), .B(n854), .Z(n852) );
  NANDN U747 ( .A(A[43]), .B(B[43]), .Z(n854) );
  AND U748 ( .A(n855), .B(n856), .Z(n853) );
  NANDN U749 ( .A(A[42]), .B(B[42]), .Z(n856) );
  NAND U750 ( .A(n857), .B(n858), .Z(n855) );
  NANDN U751 ( .A(B[42]), .B(A[42]), .Z(n858) );
  AND U752 ( .A(n859), .B(n860), .Z(n857) );
  NAND U753 ( .A(n861), .B(n862), .Z(n860) );
  NANDN U754 ( .A(A[41]), .B(B[41]), .Z(n862) );
  AND U755 ( .A(n863), .B(n864), .Z(n861) );
  NANDN U756 ( .A(A[40]), .B(B[40]), .Z(n864) );
  NAND U757 ( .A(n865), .B(n866), .Z(n863) );
  NANDN U758 ( .A(B[40]), .B(A[40]), .Z(n866) );
  AND U759 ( .A(n867), .B(n868), .Z(n865) );
  NAND U760 ( .A(n869), .B(n870), .Z(n868) );
  NANDN U761 ( .A(A[39]), .B(B[39]), .Z(n870) );
  AND U762 ( .A(n871), .B(n872), .Z(n869) );
  NANDN U763 ( .A(A[38]), .B(B[38]), .Z(n872) );
  NAND U764 ( .A(n873), .B(n874), .Z(n871) );
  NANDN U765 ( .A(B[38]), .B(A[38]), .Z(n874) );
  AND U766 ( .A(n875), .B(n876), .Z(n873) );
  NAND U767 ( .A(n877), .B(n878), .Z(n876) );
  NANDN U768 ( .A(A[37]), .B(B[37]), .Z(n878) );
  AND U769 ( .A(n879), .B(n880), .Z(n877) );
  NANDN U770 ( .A(A[36]), .B(B[36]), .Z(n880) );
  NAND U771 ( .A(n881), .B(n882), .Z(n879) );
  NANDN U772 ( .A(B[36]), .B(A[36]), .Z(n882) );
  AND U773 ( .A(n883), .B(n884), .Z(n881) );
  NAND U774 ( .A(n885), .B(n886), .Z(n884) );
  NANDN U775 ( .A(A[35]), .B(B[35]), .Z(n886) );
  AND U776 ( .A(n887), .B(n888), .Z(n885) );
  NANDN U777 ( .A(A[34]), .B(B[34]), .Z(n888) );
  NAND U778 ( .A(n889), .B(n890), .Z(n887) );
  NANDN U779 ( .A(B[34]), .B(A[34]), .Z(n890) );
  AND U780 ( .A(n891), .B(n892), .Z(n889) );
  NAND U781 ( .A(n893), .B(n894), .Z(n892) );
  NANDN U782 ( .A(A[33]), .B(B[33]), .Z(n894) );
  AND U783 ( .A(n895), .B(n896), .Z(n893) );
  NANDN U784 ( .A(A[32]), .B(B[32]), .Z(n896) );
  NAND U785 ( .A(n897), .B(n898), .Z(n895) );
  NANDN U786 ( .A(B[32]), .B(A[32]), .Z(n898) );
  AND U787 ( .A(n899), .B(n900), .Z(n897) );
  NAND U788 ( .A(n901), .B(n902), .Z(n900) );
  NANDN U789 ( .A(A[31]), .B(B[31]), .Z(n902) );
  AND U790 ( .A(n903), .B(n904), .Z(n901) );
  NANDN U791 ( .A(A[30]), .B(B[30]), .Z(n904) );
  NAND U792 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U793 ( .A(B[30]), .B(A[30]), .Z(n906) );
  AND U794 ( .A(n907), .B(n908), .Z(n905) );
  NAND U795 ( .A(n909), .B(n910), .Z(n908) );
  NANDN U796 ( .A(A[29]), .B(B[29]), .Z(n910) );
  AND U797 ( .A(n911), .B(n912), .Z(n909) );
  NANDN U798 ( .A(A[28]), .B(B[28]), .Z(n912) );
  NAND U799 ( .A(n913), .B(n914), .Z(n911) );
  NANDN U800 ( .A(B[28]), .B(A[28]), .Z(n914) );
  AND U801 ( .A(n915), .B(n916), .Z(n913) );
  NAND U802 ( .A(n917), .B(n918), .Z(n916) );
  NANDN U803 ( .A(A[27]), .B(B[27]), .Z(n918) );
  AND U804 ( .A(n919), .B(n920), .Z(n917) );
  NANDN U805 ( .A(A[26]), .B(B[26]), .Z(n920) );
  NAND U806 ( .A(n921), .B(n922), .Z(n919) );
  NANDN U807 ( .A(B[26]), .B(A[26]), .Z(n922) );
  AND U808 ( .A(n923), .B(n924), .Z(n921) );
  NAND U809 ( .A(n925), .B(n926), .Z(n924) );
  NANDN U810 ( .A(A[25]), .B(B[25]), .Z(n926) );
  AND U811 ( .A(n927), .B(n928), .Z(n925) );
  NANDN U812 ( .A(A[24]), .B(B[24]), .Z(n928) );
  NAND U813 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U814 ( .A(B[24]), .B(A[24]), .Z(n930) );
  AND U815 ( .A(n931), .B(n932), .Z(n929) );
  NAND U816 ( .A(n933), .B(n934), .Z(n932) );
  NANDN U817 ( .A(A[23]), .B(B[23]), .Z(n934) );
  AND U818 ( .A(n935), .B(n936), .Z(n933) );
  NANDN U819 ( .A(A[22]), .B(B[22]), .Z(n936) );
  NAND U820 ( .A(n937), .B(n938), .Z(n935) );
  NANDN U821 ( .A(B[22]), .B(A[22]), .Z(n938) );
  AND U822 ( .A(n939), .B(n940), .Z(n937) );
  NAND U823 ( .A(n941), .B(n942), .Z(n940) );
  NANDN U824 ( .A(A[21]), .B(B[21]), .Z(n942) );
  AND U825 ( .A(n943), .B(n944), .Z(n941) );
  NANDN U826 ( .A(A[20]), .B(B[20]), .Z(n944) );
  NAND U827 ( .A(n945), .B(n946), .Z(n943) );
  NANDN U828 ( .A(B[20]), .B(A[20]), .Z(n946) );
  AND U829 ( .A(n947), .B(n948), .Z(n945) );
  NAND U830 ( .A(n949), .B(n950), .Z(n948) );
  NANDN U831 ( .A(A[19]), .B(B[19]), .Z(n950) );
  AND U832 ( .A(n951), .B(n952), .Z(n949) );
  NANDN U833 ( .A(A[18]), .B(B[18]), .Z(n952) );
  NAND U834 ( .A(n953), .B(n954), .Z(n951) );
  NANDN U835 ( .A(B[18]), .B(A[18]), .Z(n954) );
  AND U836 ( .A(n955), .B(n956), .Z(n953) );
  NAND U837 ( .A(n957), .B(n958), .Z(n956) );
  NANDN U838 ( .A(A[17]), .B(B[17]), .Z(n958) );
  AND U839 ( .A(n959), .B(n960), .Z(n957) );
  NANDN U840 ( .A(A[16]), .B(B[16]), .Z(n960) );
  NAND U841 ( .A(n961), .B(n962), .Z(n959) );
  NANDN U842 ( .A(B[16]), .B(A[16]), .Z(n962) );
  AND U843 ( .A(n963), .B(n964), .Z(n961) );
  NAND U844 ( .A(n965), .B(n966), .Z(n964) );
  NANDN U845 ( .A(A[15]), .B(B[15]), .Z(n966) );
  AND U846 ( .A(n967), .B(n968), .Z(n965) );
  NANDN U847 ( .A(A[14]), .B(B[14]), .Z(n968) );
  NAND U848 ( .A(n969), .B(n970), .Z(n967) );
  NANDN U849 ( .A(B[14]), .B(A[14]), .Z(n970) );
  AND U850 ( .A(n971), .B(n972), .Z(n969) );
  NAND U851 ( .A(n973), .B(n974), .Z(n972) );
  NANDN U852 ( .A(A[13]), .B(B[13]), .Z(n974) );
  AND U853 ( .A(n975), .B(n976), .Z(n973) );
  NANDN U854 ( .A(A[12]), .B(B[12]), .Z(n976) );
  NAND U855 ( .A(n977), .B(n978), .Z(n975) );
  NANDN U856 ( .A(B[12]), .B(A[12]), .Z(n978) );
  AND U857 ( .A(n979), .B(n980), .Z(n977) );
  NAND U858 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U859 ( .A(A[11]), .B(B[11]), .Z(n982) );
  AND U860 ( .A(n983), .B(n984), .Z(n981) );
  NANDN U861 ( .A(A[10]), .B(B[10]), .Z(n984) );
  NAND U862 ( .A(n985), .B(n986), .Z(n983) );
  NANDN U863 ( .A(B[9]), .B(A[9]), .Z(n986) );
  AND U864 ( .A(n987), .B(n988), .Z(n985) );
  NAND U865 ( .A(n989), .B(n990), .Z(n988) );
  NANDN U866 ( .A(A[9]), .B(B[9]), .Z(n990) );
  AND U867 ( .A(n991), .B(n992), .Z(n989) );
  NANDN U868 ( .A(A[8]), .B(B[8]), .Z(n992) );
  NAND U869 ( .A(n993), .B(n994), .Z(n991) );
  NANDN U870 ( .A(B[8]), .B(A[8]), .Z(n994) );
  AND U871 ( .A(n995), .B(n996), .Z(n993) );
  NAND U872 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U873 ( .A(A[7]), .B(B[7]), .Z(n998) );
  AND U874 ( .A(n999), .B(n1000), .Z(n997) );
  NANDN U875 ( .A(A[6]), .B(B[6]), .Z(n1000) );
  NAND U876 ( .A(n1001), .B(n1002), .Z(n999) );
  NANDN U877 ( .A(B[6]), .B(A[6]), .Z(n1002) );
  AND U878 ( .A(n1003), .B(n1004), .Z(n1001) );
  NAND U879 ( .A(n1005), .B(n1006), .Z(n1004) );
  NANDN U880 ( .A(A[5]), .B(B[5]), .Z(n1006) );
  AND U881 ( .A(n1007), .B(n1008), .Z(n1005) );
  NANDN U882 ( .A(A[4]), .B(B[4]), .Z(n1008) );
  NAND U883 ( .A(n1009), .B(n1010), .Z(n1007) );
  NANDN U884 ( .A(B[4]), .B(A[4]), .Z(n1010) );
  AND U885 ( .A(n1011), .B(n1012), .Z(n1009) );
  NAND U886 ( .A(n1013), .B(n1014), .Z(n1012) );
  NANDN U887 ( .A(A[3]), .B(B[3]), .Z(n1014) );
  AND U888 ( .A(n1015), .B(n1016), .Z(n1013) );
  NANDN U889 ( .A(A[2]), .B(B[2]), .Z(n1016) );
  NAND U890 ( .A(n1017), .B(n1018), .Z(n1015) );
  NANDN U891 ( .A(B[2]), .B(A[2]), .Z(n1018) );
  AND U892 ( .A(n1019), .B(n1020), .Z(n1017) );
  NANDN U893 ( .A(B[1]), .B(n1021), .Z(n1020) );
  NANDN U894 ( .A(A[1]), .B(n1022), .Z(n1021) );
  NANDN U895 ( .A(n1022), .B(A[1]), .Z(n1019) );
  ANDN U896 ( .B(B[0]), .A(A[0]), .Z(n1022) );
  NANDN U897 ( .A(B[3]), .B(A[3]), .Z(n1011) );
  NANDN U898 ( .A(B[5]), .B(A[5]), .Z(n1003) );
  NANDN U899 ( .A(B[7]), .B(A[7]), .Z(n995) );
  NANDN U900 ( .A(B[10]), .B(A[10]), .Z(n987) );
  NANDN U901 ( .A(B[11]), .B(A[11]), .Z(n979) );
  NANDN U902 ( .A(B[13]), .B(A[13]), .Z(n971) );
  NANDN U903 ( .A(B[15]), .B(A[15]), .Z(n963) );
  NANDN U904 ( .A(B[17]), .B(A[17]), .Z(n955) );
  NANDN U905 ( .A(B[19]), .B(A[19]), .Z(n947) );
  NANDN U906 ( .A(B[21]), .B(A[21]), .Z(n939) );
  NANDN U907 ( .A(B[23]), .B(A[23]), .Z(n931) );
  NANDN U908 ( .A(B[25]), .B(A[25]), .Z(n923) );
  NANDN U909 ( .A(B[27]), .B(A[27]), .Z(n915) );
  NANDN U910 ( .A(B[29]), .B(A[29]), .Z(n907) );
  NANDN U911 ( .A(B[31]), .B(A[31]), .Z(n899) );
  NANDN U912 ( .A(B[33]), .B(A[33]), .Z(n891) );
  NANDN U913 ( .A(B[35]), .B(A[35]), .Z(n883) );
  NANDN U914 ( .A(B[37]), .B(A[37]), .Z(n875) );
  NANDN U915 ( .A(B[39]), .B(A[39]), .Z(n867) );
  NANDN U916 ( .A(B[41]), .B(A[41]), .Z(n859) );
  NANDN U917 ( .A(B[43]), .B(A[43]), .Z(n851) );
  NANDN U918 ( .A(B[45]), .B(A[45]), .Z(n843) );
  NANDN U919 ( .A(B[47]), .B(A[47]), .Z(n835) );
  NANDN U920 ( .A(B[49]), .B(A[49]), .Z(n827) );
  NANDN U921 ( .A(B[51]), .B(A[51]), .Z(n819) );
  NANDN U922 ( .A(B[53]), .B(A[53]), .Z(n811) );
  NANDN U923 ( .A(B[55]), .B(A[55]), .Z(n803) );
  NANDN U924 ( .A(B[57]), .B(A[57]), .Z(n795) );
  NANDN U925 ( .A(B[59]), .B(A[59]), .Z(n787) );
  NANDN U926 ( .A(B[61]), .B(A[61]), .Z(n779) );
  NANDN U927 ( .A(B[63]), .B(A[63]), .Z(n771) );
  NANDN U928 ( .A(B[65]), .B(A[65]), .Z(n763) );
  NANDN U929 ( .A(B[67]), .B(A[67]), .Z(n755) );
  NANDN U930 ( .A(B[69]), .B(A[69]), .Z(n747) );
  NANDN U931 ( .A(B[71]), .B(A[71]), .Z(n739) );
  NANDN U932 ( .A(B[73]), .B(A[73]), .Z(n731) );
  NANDN U933 ( .A(B[75]), .B(A[75]), .Z(n723) );
  NANDN U934 ( .A(B[77]), .B(A[77]), .Z(n715) );
  NANDN U935 ( .A(B[79]), .B(A[79]), .Z(n707) );
  NANDN U936 ( .A(B[81]), .B(A[81]), .Z(n699) );
  NANDN U937 ( .A(B[83]), .B(A[83]), .Z(n691) );
  NANDN U938 ( .A(B[85]), .B(A[85]), .Z(n683) );
  NANDN U939 ( .A(B[87]), .B(A[87]), .Z(n675) );
  NANDN U940 ( .A(B[89]), .B(A[89]), .Z(n667) );
  NANDN U941 ( .A(B[91]), .B(A[91]), .Z(n659) );
  NANDN U942 ( .A(B[93]), .B(A[93]), .Z(n651) );
  NANDN U943 ( .A(B[95]), .B(A[95]), .Z(n643) );
  NANDN U944 ( .A(B[97]), .B(A[97]), .Z(n635) );
  NANDN U945 ( .A(B[100]), .B(A[100]), .Z(n627) );
  NANDN U946 ( .A(B[101]), .B(A[101]), .Z(n619) );
  NANDN U947 ( .A(B[103]), .B(A[103]), .Z(n611) );
  NANDN U948 ( .A(B[105]), .B(A[105]), .Z(n603) );
  NANDN U949 ( .A(B[107]), .B(A[107]), .Z(n595) );
  NANDN U950 ( .A(B[109]), .B(A[109]), .Z(n587) );
  NANDN U951 ( .A(B[111]), .B(A[111]), .Z(n579) );
  NANDN U952 ( .A(B[113]), .B(A[113]), .Z(n571) );
  NANDN U953 ( .A(B[115]), .B(A[115]), .Z(n563) );
  NANDN U954 ( .A(B[117]), .B(A[117]), .Z(n555) );
  NANDN U955 ( .A(B[119]), .B(A[119]), .Z(n547) );
  NANDN U956 ( .A(B[121]), .B(A[121]), .Z(n539) );
  NANDN U957 ( .A(B[123]), .B(A[123]), .Z(n531) );
  NANDN U958 ( .A(B[125]), .B(A[125]), .Z(n523) );
  NANDN U959 ( .A(B[127]), .B(A[127]), .Z(n515) );
  NANDN U960 ( .A(B[129]), .B(A[129]), .Z(n507) );
  NANDN U961 ( .A(B[131]), .B(A[131]), .Z(n499) );
  NANDN U962 ( .A(B[133]), .B(A[133]), .Z(n491) );
  NANDN U963 ( .A(B[135]), .B(A[135]), .Z(n483) );
  NANDN U964 ( .A(B[137]), .B(A[137]), .Z(n475) );
  NANDN U965 ( .A(B[139]), .B(A[139]), .Z(n467) );
  NANDN U966 ( .A(B[141]), .B(A[141]), .Z(n459) );
  NANDN U967 ( .A(B[143]), .B(A[143]), .Z(n451) );
  NANDN U968 ( .A(B[145]), .B(A[145]), .Z(n443) );
  NANDN U969 ( .A(B[147]), .B(A[147]), .Z(n435) );
  NANDN U970 ( .A(B[149]), .B(A[149]), .Z(n427) );
  NANDN U971 ( .A(B[151]), .B(A[151]), .Z(n419) );
  NANDN U972 ( .A(B[153]), .B(A[153]), .Z(n411) );
  NANDN U973 ( .A(B[155]), .B(A[155]), .Z(n403) );
  NANDN U974 ( .A(B[157]), .B(A[157]), .Z(n395) );
  NANDN U975 ( .A(B[159]), .B(A[159]), .Z(n387) );
  NANDN U976 ( .A(B[161]), .B(A[161]), .Z(n379) );
  NANDN U977 ( .A(B[163]), .B(A[163]), .Z(n371) );
  NANDN U978 ( .A(B[165]), .B(A[165]), .Z(n363) );
  NANDN U979 ( .A(B[167]), .B(A[167]), .Z(n355) );
  NANDN U980 ( .A(B[169]), .B(A[169]), .Z(n347) );
  NANDN U981 ( .A(B[171]), .B(A[171]), .Z(n339) );
  NANDN U982 ( .A(B[173]), .B(A[173]), .Z(n331) );
  NANDN U983 ( .A(B[175]), .B(A[175]), .Z(n323) );
  NANDN U984 ( .A(B[177]), .B(A[177]), .Z(n315) );
  NANDN U985 ( .A(B[179]), .B(A[179]), .Z(n307) );
  NANDN U986 ( .A(B[181]), .B(A[181]), .Z(n299) );
  NANDN U987 ( .A(B[183]), .B(A[183]), .Z(n291) );
  NANDN U988 ( .A(B[185]), .B(A[185]), .Z(n283) );
  NANDN U989 ( .A(B[187]), .B(A[187]), .Z(n275) );
  NANDN U990 ( .A(B[189]), .B(A[189]), .Z(n267) );
  NANDN U991 ( .A(B[191]), .B(A[191]), .Z(n259) );
  NANDN U992 ( .A(B[193]), .B(A[193]), .Z(n251) );
  NANDN U993 ( .A(B[195]), .B(A[195]), .Z(n243) );
  NANDN U994 ( .A(B[197]), .B(A[197]), .Z(n235) );
  NANDN U995 ( .A(B[199]), .B(A[199]), .Z(n227) );
  NANDN U996 ( .A(B[201]), .B(A[201]), .Z(n219) );
  NANDN U997 ( .A(B[203]), .B(A[203]), .Z(n211) );
  NANDN U998 ( .A(B[205]), .B(A[205]), .Z(n203) );
  NANDN U999 ( .A(B[207]), .B(A[207]), .Z(n195) );
  NANDN U1000 ( .A(B[209]), .B(A[209]), .Z(n187) );
  NANDN U1001 ( .A(B[211]), .B(A[211]), .Z(n179) );
  NANDN U1002 ( .A(B[213]), .B(A[213]), .Z(n171) );
  NANDN U1003 ( .A(B[215]), .B(A[215]), .Z(n163) );
  NANDN U1004 ( .A(B[217]), .B(A[217]), .Z(n155) );
  NANDN U1005 ( .A(B[219]), .B(A[219]), .Z(n147) );
  NANDN U1006 ( .A(B[221]), .B(A[221]), .Z(n139) );
  NANDN U1007 ( .A(B[223]), .B(A[223]), .Z(n131) );
  NANDN U1008 ( .A(B[225]), .B(A[225]), .Z(n123) );
  NANDN U1009 ( .A(B[227]), .B(A[227]), .Z(n115) );
  NANDN U1010 ( .A(B[229]), .B(A[229]), .Z(n107) );
  NANDN U1011 ( .A(B[231]), .B(A[231]), .Z(n99) );
  NANDN U1012 ( .A(B[233]), .B(A[233]), .Z(n91) );
  NANDN U1013 ( .A(B[235]), .B(A[235]), .Z(n83) );
  NANDN U1014 ( .A(B[237]), .B(A[237]), .Z(n75) );
  NANDN U1015 ( .A(B[239]), .B(A[239]), .Z(n67) );
  NANDN U1016 ( .A(B[241]), .B(A[241]), .Z(n59) );
  NANDN U1017 ( .A(B[243]), .B(A[243]), .Z(n51) );
  NANDN U1018 ( .A(B[245]), .B(A[245]), .Z(n43) );
  NANDN U1019 ( .A(B[247]), .B(A[247]), .Z(n35) );
  NANDN U1020 ( .A(B[249]), .B(A[249]), .Z(n27) );
  NANDN U1021 ( .A(B[251]), .B(A[251]), .Z(n19) );
  NANDN U1022 ( .A(B[253]), .B(A[253]), .Z(n11) );
  NANDN U1023 ( .A(A[255]), .B(B[255]), .Z(n3) );
endmodule


module modmult_step_N256_5_DW01_add_0 ( A, B, CI, SUM, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] SUM;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272;
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];

  XNOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(SUM[99]) );
  XNOR U4 ( .A(B[99]), .B(A[99]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[98]) );
  XNOR U6 ( .A(B[98]), .B(A[98]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[97]) );
  XNOR U8 ( .A(B[97]), .B(A[97]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[96]) );
  XNOR U10 ( .A(B[96]), .B(A[96]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[95]) );
  XNOR U12 ( .A(B[95]), .B(A[95]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[94]) );
  XNOR U14 ( .A(B[94]), .B(A[94]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[93]) );
  XNOR U16 ( .A(B[93]), .B(A[93]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(SUM[92]) );
  XNOR U18 ( .A(B[92]), .B(A[92]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(SUM[91]) );
  XNOR U20 ( .A(B[91]), .B(A[91]), .Z(n20) );
  XOR U21 ( .A(n21), .B(n22), .Z(SUM[90]) );
  XNOR U22 ( .A(B[90]), .B(A[90]), .Z(n22) );
  XOR U23 ( .A(n23), .B(n24), .Z(SUM[8]) );
  XNOR U24 ( .A(B[8]), .B(A[8]), .Z(n24) );
  XOR U25 ( .A(n25), .B(n26), .Z(SUM[89]) );
  XNOR U26 ( .A(B[89]), .B(A[89]), .Z(n26) );
  XOR U27 ( .A(n27), .B(n28), .Z(SUM[88]) );
  XNOR U28 ( .A(B[88]), .B(A[88]), .Z(n28) );
  XOR U29 ( .A(n29), .B(n30), .Z(SUM[87]) );
  XNOR U30 ( .A(B[87]), .B(A[87]), .Z(n30) );
  XOR U31 ( .A(n31), .B(n32), .Z(SUM[86]) );
  XNOR U32 ( .A(B[86]), .B(A[86]), .Z(n32) );
  XOR U33 ( .A(n33), .B(n34), .Z(SUM[85]) );
  XNOR U34 ( .A(B[85]), .B(A[85]), .Z(n34) );
  XOR U35 ( .A(n35), .B(n36), .Z(SUM[84]) );
  XNOR U36 ( .A(B[84]), .B(A[84]), .Z(n36) );
  XOR U37 ( .A(n37), .B(n38), .Z(SUM[83]) );
  XNOR U38 ( .A(B[83]), .B(A[83]), .Z(n38) );
  XOR U39 ( .A(n39), .B(n40), .Z(SUM[82]) );
  XNOR U40 ( .A(B[82]), .B(A[82]), .Z(n40) );
  XOR U41 ( .A(n41), .B(n42), .Z(SUM[81]) );
  XNOR U42 ( .A(B[81]), .B(A[81]), .Z(n42) );
  XOR U43 ( .A(n43), .B(n44), .Z(SUM[80]) );
  XNOR U44 ( .A(B[80]), .B(A[80]), .Z(n44) );
  XOR U45 ( .A(n45), .B(n46), .Z(SUM[7]) );
  XNOR U46 ( .A(B[7]), .B(A[7]), .Z(n46) );
  XOR U47 ( .A(n47), .B(n48), .Z(SUM[79]) );
  XNOR U48 ( .A(B[79]), .B(A[79]), .Z(n48) );
  XOR U49 ( .A(n49), .B(n50), .Z(SUM[78]) );
  XNOR U50 ( .A(B[78]), .B(A[78]), .Z(n50) );
  XOR U51 ( .A(n51), .B(n52), .Z(SUM[77]) );
  XNOR U52 ( .A(B[77]), .B(A[77]), .Z(n52) );
  XOR U53 ( .A(n53), .B(n54), .Z(SUM[76]) );
  XNOR U54 ( .A(B[76]), .B(A[76]), .Z(n54) );
  XOR U55 ( .A(n55), .B(n56), .Z(SUM[75]) );
  XNOR U56 ( .A(B[75]), .B(A[75]), .Z(n56) );
  XOR U57 ( .A(n57), .B(n58), .Z(SUM[74]) );
  XNOR U58 ( .A(B[74]), .B(A[74]), .Z(n58) );
  XOR U59 ( .A(n59), .B(n60), .Z(SUM[73]) );
  XNOR U60 ( .A(B[73]), .B(A[73]), .Z(n60) );
  XOR U61 ( .A(n61), .B(n62), .Z(SUM[72]) );
  XNOR U62 ( .A(B[72]), .B(A[72]), .Z(n62) );
  XOR U63 ( .A(n63), .B(n64), .Z(SUM[71]) );
  XNOR U64 ( .A(B[71]), .B(A[71]), .Z(n64) );
  XOR U65 ( .A(n65), .B(n66), .Z(SUM[70]) );
  XNOR U66 ( .A(B[70]), .B(A[70]), .Z(n66) );
  XOR U67 ( .A(n67), .B(n68), .Z(SUM[6]) );
  XNOR U68 ( .A(B[6]), .B(A[6]), .Z(n68) );
  XOR U69 ( .A(n69), .B(n70), .Z(SUM[69]) );
  XNOR U70 ( .A(B[69]), .B(A[69]), .Z(n70) );
  XOR U71 ( .A(n71), .B(n72), .Z(SUM[68]) );
  XNOR U72 ( .A(B[68]), .B(A[68]), .Z(n72) );
  XOR U73 ( .A(n73), .B(n74), .Z(SUM[67]) );
  XNOR U74 ( .A(B[67]), .B(A[67]), .Z(n74) );
  XOR U75 ( .A(n75), .B(n76), .Z(SUM[66]) );
  XNOR U76 ( .A(B[66]), .B(A[66]), .Z(n76) );
  XOR U77 ( .A(n77), .B(n78), .Z(SUM[65]) );
  XNOR U78 ( .A(B[65]), .B(A[65]), .Z(n78) );
  XOR U79 ( .A(n79), .B(n80), .Z(SUM[64]) );
  XNOR U80 ( .A(B[64]), .B(A[64]), .Z(n80) );
  XOR U81 ( .A(n81), .B(n82), .Z(SUM[63]) );
  XNOR U82 ( .A(B[63]), .B(A[63]), .Z(n82) );
  XOR U83 ( .A(n83), .B(n84), .Z(SUM[62]) );
  XNOR U84 ( .A(B[62]), .B(A[62]), .Z(n84) );
  XOR U85 ( .A(n85), .B(n86), .Z(SUM[61]) );
  XNOR U86 ( .A(B[61]), .B(A[61]), .Z(n86) );
  XOR U87 ( .A(n87), .B(n88), .Z(SUM[60]) );
  XNOR U88 ( .A(B[60]), .B(A[60]), .Z(n88) );
  XOR U89 ( .A(n89), .B(n90), .Z(SUM[5]) );
  XNOR U90 ( .A(B[5]), .B(A[5]), .Z(n90) );
  XOR U91 ( .A(n91), .B(n92), .Z(SUM[59]) );
  XNOR U92 ( .A(B[59]), .B(A[59]), .Z(n92) );
  XOR U93 ( .A(n93), .B(n94), .Z(SUM[58]) );
  XNOR U94 ( .A(B[58]), .B(A[58]), .Z(n94) );
  XOR U95 ( .A(n95), .B(n96), .Z(SUM[57]) );
  XNOR U96 ( .A(B[57]), .B(A[57]), .Z(n96) );
  XOR U97 ( .A(n97), .B(n98), .Z(SUM[56]) );
  XNOR U98 ( .A(B[56]), .B(A[56]), .Z(n98) );
  XOR U99 ( .A(n99), .B(n100), .Z(SUM[55]) );
  XNOR U100 ( .A(B[55]), .B(A[55]), .Z(n100) );
  XOR U101 ( .A(n101), .B(n102), .Z(SUM[54]) );
  XNOR U102 ( .A(B[54]), .B(A[54]), .Z(n102) );
  XOR U103 ( .A(n103), .B(n104), .Z(SUM[53]) );
  XNOR U104 ( .A(B[53]), .B(A[53]), .Z(n104) );
  XOR U105 ( .A(n105), .B(n106), .Z(SUM[52]) );
  XNOR U106 ( .A(B[52]), .B(A[52]), .Z(n106) );
  XOR U107 ( .A(n107), .B(n108), .Z(SUM[51]) );
  XNOR U108 ( .A(B[51]), .B(A[51]), .Z(n108) );
  XOR U109 ( .A(n109), .B(n110), .Z(SUM[50]) );
  XNOR U110 ( .A(B[50]), .B(A[50]), .Z(n110) );
  XOR U111 ( .A(n111), .B(n112), .Z(SUM[4]) );
  XNOR U112 ( .A(B[4]), .B(A[4]), .Z(n112) );
  XOR U113 ( .A(n113), .B(n114), .Z(SUM[49]) );
  XNOR U114 ( .A(B[49]), .B(A[49]), .Z(n114) );
  XOR U115 ( .A(n115), .B(n116), .Z(SUM[48]) );
  XNOR U116 ( .A(B[48]), .B(A[48]), .Z(n116) );
  XOR U117 ( .A(n117), .B(n118), .Z(SUM[47]) );
  XNOR U118 ( .A(B[47]), .B(A[47]), .Z(n118) );
  XOR U119 ( .A(n119), .B(n120), .Z(SUM[46]) );
  XNOR U120 ( .A(B[46]), .B(A[46]), .Z(n120) );
  XOR U121 ( .A(n121), .B(n122), .Z(SUM[45]) );
  XNOR U122 ( .A(B[45]), .B(A[45]), .Z(n122) );
  XOR U123 ( .A(n123), .B(n124), .Z(SUM[44]) );
  XNOR U124 ( .A(B[44]), .B(A[44]), .Z(n124) );
  XOR U125 ( .A(n125), .B(n126), .Z(SUM[43]) );
  XNOR U126 ( .A(B[43]), .B(A[43]), .Z(n126) );
  XOR U127 ( .A(n127), .B(n128), .Z(SUM[42]) );
  XNOR U128 ( .A(B[42]), .B(A[42]), .Z(n128) );
  XOR U129 ( .A(n129), .B(n130), .Z(SUM[41]) );
  XNOR U130 ( .A(B[41]), .B(A[41]), .Z(n130) );
  XOR U131 ( .A(n131), .B(n132), .Z(SUM[40]) );
  XNOR U132 ( .A(B[40]), .B(A[40]), .Z(n132) );
  XOR U133 ( .A(n133), .B(n134), .Z(SUM[3]) );
  XNOR U134 ( .A(B[3]), .B(A[3]), .Z(n134) );
  XOR U135 ( .A(n135), .B(n136), .Z(SUM[39]) );
  XNOR U136 ( .A(B[39]), .B(A[39]), .Z(n136) );
  XOR U137 ( .A(n137), .B(n138), .Z(SUM[38]) );
  XNOR U138 ( .A(B[38]), .B(A[38]), .Z(n138) );
  XOR U139 ( .A(n139), .B(n140), .Z(SUM[37]) );
  XNOR U140 ( .A(B[37]), .B(A[37]), .Z(n140) );
  XOR U141 ( .A(n141), .B(n142), .Z(SUM[36]) );
  XNOR U142 ( .A(B[36]), .B(A[36]), .Z(n142) );
  XOR U143 ( .A(n143), .B(n144), .Z(SUM[35]) );
  XNOR U144 ( .A(B[35]), .B(A[35]), .Z(n144) );
  XOR U145 ( .A(n145), .B(n146), .Z(SUM[34]) );
  XNOR U146 ( .A(B[34]), .B(A[34]), .Z(n146) );
  XOR U147 ( .A(n147), .B(n148), .Z(SUM[33]) );
  XNOR U148 ( .A(B[33]), .B(A[33]), .Z(n148) );
  XOR U149 ( .A(n149), .B(n150), .Z(SUM[32]) );
  XNOR U150 ( .A(B[32]), .B(A[32]), .Z(n150) );
  XOR U151 ( .A(n151), .B(n152), .Z(SUM[31]) );
  XNOR U152 ( .A(B[31]), .B(A[31]), .Z(n152) );
  XOR U153 ( .A(n153), .B(n154), .Z(SUM[30]) );
  XNOR U154 ( .A(B[30]), .B(A[30]), .Z(n154) );
  XOR U155 ( .A(n155), .B(n156), .Z(SUM[2]) );
  XOR U156 ( .A(B[2]), .B(A[2]), .Z(n156) );
  XOR U157 ( .A(n157), .B(n158), .Z(SUM[29]) );
  XNOR U158 ( .A(B[29]), .B(A[29]), .Z(n158) );
  XOR U159 ( .A(n159), .B(n160), .Z(SUM[28]) );
  XNOR U160 ( .A(B[28]), .B(A[28]), .Z(n160) );
  XOR U161 ( .A(n161), .B(n162), .Z(SUM[27]) );
  XNOR U162 ( .A(B[27]), .B(A[27]), .Z(n162) );
  XOR U163 ( .A(n163), .B(n164), .Z(SUM[26]) );
  XNOR U164 ( .A(B[26]), .B(A[26]), .Z(n164) );
  XOR U165 ( .A(n165), .B(n166), .Z(SUM[25]) );
  XNOR U166 ( .A(B[25]), .B(A[25]), .Z(n166) );
  XOR U167 ( .A(A[257]), .B(n167), .Z(SUM[257]) );
  AND U168 ( .A(A[256]), .B(n168), .Z(n167) );
  XOR U169 ( .A(A[256]), .B(n168), .Z(SUM[256]) );
  NAND U170 ( .A(n169), .B(n170), .Z(n168) );
  NAND U171 ( .A(B[255]), .B(n171), .Z(n170) );
  NANDN U172 ( .A(A[255]), .B(n172), .Z(n171) );
  NANDN U173 ( .A(n172), .B(A[255]), .Z(n169) );
  XOR U174 ( .A(n172), .B(n173), .Z(SUM[255]) );
  XNOR U175 ( .A(B[255]), .B(A[255]), .Z(n173) );
  AND U176 ( .A(n174), .B(n175), .Z(n172) );
  NAND U177 ( .A(B[254]), .B(n176), .Z(n175) );
  NANDN U178 ( .A(A[254]), .B(n177), .Z(n176) );
  NANDN U179 ( .A(n177), .B(A[254]), .Z(n174) );
  XOR U180 ( .A(n177), .B(n178), .Z(SUM[254]) );
  XNOR U181 ( .A(B[254]), .B(A[254]), .Z(n178) );
  AND U182 ( .A(n179), .B(n180), .Z(n177) );
  NAND U183 ( .A(B[253]), .B(n181), .Z(n180) );
  NANDN U184 ( .A(A[253]), .B(n182), .Z(n181) );
  NANDN U185 ( .A(n182), .B(A[253]), .Z(n179) );
  XOR U186 ( .A(n182), .B(n183), .Z(SUM[253]) );
  XNOR U187 ( .A(B[253]), .B(A[253]), .Z(n183) );
  AND U188 ( .A(n184), .B(n185), .Z(n182) );
  NAND U189 ( .A(B[252]), .B(n186), .Z(n185) );
  NANDN U190 ( .A(A[252]), .B(n187), .Z(n186) );
  NANDN U191 ( .A(n187), .B(A[252]), .Z(n184) );
  XOR U192 ( .A(n187), .B(n188), .Z(SUM[252]) );
  XNOR U193 ( .A(B[252]), .B(A[252]), .Z(n188) );
  AND U194 ( .A(n189), .B(n190), .Z(n187) );
  NAND U195 ( .A(B[251]), .B(n191), .Z(n190) );
  NANDN U196 ( .A(A[251]), .B(n192), .Z(n191) );
  NANDN U197 ( .A(n192), .B(A[251]), .Z(n189) );
  XOR U198 ( .A(n192), .B(n193), .Z(SUM[251]) );
  XNOR U199 ( .A(B[251]), .B(A[251]), .Z(n193) );
  AND U200 ( .A(n194), .B(n195), .Z(n192) );
  NAND U201 ( .A(B[250]), .B(n196), .Z(n195) );
  NANDN U202 ( .A(A[250]), .B(n197), .Z(n196) );
  NANDN U203 ( .A(n197), .B(A[250]), .Z(n194) );
  XOR U204 ( .A(n197), .B(n198), .Z(SUM[250]) );
  XNOR U205 ( .A(B[250]), .B(A[250]), .Z(n198) );
  AND U206 ( .A(n199), .B(n200), .Z(n197) );
  NAND U207 ( .A(B[249]), .B(n201), .Z(n200) );
  NANDN U208 ( .A(A[249]), .B(n202), .Z(n201) );
  NANDN U209 ( .A(n202), .B(A[249]), .Z(n199) );
  XOR U210 ( .A(n203), .B(n204), .Z(SUM[24]) );
  XNOR U211 ( .A(B[24]), .B(A[24]), .Z(n204) );
  XOR U212 ( .A(n202), .B(n205), .Z(SUM[249]) );
  XNOR U213 ( .A(B[249]), .B(A[249]), .Z(n205) );
  AND U214 ( .A(n206), .B(n207), .Z(n202) );
  NAND U215 ( .A(B[248]), .B(n208), .Z(n207) );
  NANDN U216 ( .A(A[248]), .B(n209), .Z(n208) );
  NANDN U217 ( .A(n209), .B(A[248]), .Z(n206) );
  XOR U218 ( .A(n209), .B(n210), .Z(SUM[248]) );
  XNOR U219 ( .A(B[248]), .B(A[248]), .Z(n210) );
  AND U220 ( .A(n211), .B(n212), .Z(n209) );
  NAND U221 ( .A(B[247]), .B(n213), .Z(n212) );
  NANDN U222 ( .A(A[247]), .B(n214), .Z(n213) );
  NANDN U223 ( .A(n214), .B(A[247]), .Z(n211) );
  XOR U224 ( .A(n214), .B(n215), .Z(SUM[247]) );
  XNOR U225 ( .A(B[247]), .B(A[247]), .Z(n215) );
  AND U226 ( .A(n216), .B(n217), .Z(n214) );
  NAND U227 ( .A(B[246]), .B(n218), .Z(n217) );
  NANDN U228 ( .A(A[246]), .B(n219), .Z(n218) );
  NANDN U229 ( .A(n219), .B(A[246]), .Z(n216) );
  XOR U230 ( .A(n219), .B(n220), .Z(SUM[246]) );
  XNOR U231 ( .A(B[246]), .B(A[246]), .Z(n220) );
  AND U232 ( .A(n221), .B(n222), .Z(n219) );
  NAND U233 ( .A(B[245]), .B(n223), .Z(n222) );
  NANDN U234 ( .A(A[245]), .B(n224), .Z(n223) );
  NANDN U235 ( .A(n224), .B(A[245]), .Z(n221) );
  XOR U236 ( .A(n224), .B(n225), .Z(SUM[245]) );
  XNOR U237 ( .A(B[245]), .B(A[245]), .Z(n225) );
  AND U238 ( .A(n226), .B(n227), .Z(n224) );
  NAND U239 ( .A(B[244]), .B(n228), .Z(n227) );
  NANDN U240 ( .A(A[244]), .B(n229), .Z(n228) );
  NANDN U241 ( .A(n229), .B(A[244]), .Z(n226) );
  XOR U242 ( .A(n229), .B(n230), .Z(SUM[244]) );
  XNOR U243 ( .A(B[244]), .B(A[244]), .Z(n230) );
  AND U244 ( .A(n231), .B(n232), .Z(n229) );
  NAND U245 ( .A(B[243]), .B(n233), .Z(n232) );
  NANDN U246 ( .A(A[243]), .B(n234), .Z(n233) );
  NANDN U247 ( .A(n234), .B(A[243]), .Z(n231) );
  XOR U248 ( .A(n234), .B(n235), .Z(SUM[243]) );
  XNOR U249 ( .A(B[243]), .B(A[243]), .Z(n235) );
  AND U250 ( .A(n236), .B(n237), .Z(n234) );
  NAND U251 ( .A(B[242]), .B(n238), .Z(n237) );
  NANDN U252 ( .A(A[242]), .B(n239), .Z(n238) );
  NANDN U253 ( .A(n239), .B(A[242]), .Z(n236) );
  XOR U254 ( .A(n239), .B(n240), .Z(SUM[242]) );
  XNOR U255 ( .A(B[242]), .B(A[242]), .Z(n240) );
  AND U256 ( .A(n241), .B(n242), .Z(n239) );
  NAND U257 ( .A(B[241]), .B(n243), .Z(n242) );
  NANDN U258 ( .A(A[241]), .B(n244), .Z(n243) );
  NANDN U259 ( .A(n244), .B(A[241]), .Z(n241) );
  XOR U260 ( .A(n244), .B(n245), .Z(SUM[241]) );
  XNOR U261 ( .A(B[241]), .B(A[241]), .Z(n245) );
  AND U262 ( .A(n246), .B(n247), .Z(n244) );
  NAND U263 ( .A(B[240]), .B(n248), .Z(n247) );
  NANDN U264 ( .A(A[240]), .B(n249), .Z(n248) );
  NANDN U265 ( .A(n249), .B(A[240]), .Z(n246) );
  XOR U266 ( .A(n249), .B(n250), .Z(SUM[240]) );
  XNOR U267 ( .A(B[240]), .B(A[240]), .Z(n250) );
  AND U268 ( .A(n251), .B(n252), .Z(n249) );
  NAND U269 ( .A(B[239]), .B(n253), .Z(n252) );
  NANDN U270 ( .A(A[239]), .B(n254), .Z(n253) );
  NANDN U271 ( .A(n254), .B(A[239]), .Z(n251) );
  XOR U272 ( .A(n255), .B(n256), .Z(SUM[23]) );
  XNOR U273 ( .A(B[23]), .B(A[23]), .Z(n256) );
  XOR U274 ( .A(n254), .B(n257), .Z(SUM[239]) );
  XNOR U275 ( .A(B[239]), .B(A[239]), .Z(n257) );
  AND U276 ( .A(n258), .B(n259), .Z(n254) );
  NAND U277 ( .A(B[238]), .B(n260), .Z(n259) );
  NANDN U278 ( .A(A[238]), .B(n261), .Z(n260) );
  NANDN U279 ( .A(n261), .B(A[238]), .Z(n258) );
  XOR U280 ( .A(n261), .B(n262), .Z(SUM[238]) );
  XNOR U281 ( .A(B[238]), .B(A[238]), .Z(n262) );
  AND U282 ( .A(n263), .B(n264), .Z(n261) );
  NAND U283 ( .A(B[237]), .B(n265), .Z(n264) );
  NANDN U284 ( .A(A[237]), .B(n266), .Z(n265) );
  NANDN U285 ( .A(n266), .B(A[237]), .Z(n263) );
  XOR U286 ( .A(n266), .B(n267), .Z(SUM[237]) );
  XNOR U287 ( .A(B[237]), .B(A[237]), .Z(n267) );
  AND U288 ( .A(n268), .B(n269), .Z(n266) );
  NAND U289 ( .A(B[236]), .B(n270), .Z(n269) );
  NANDN U290 ( .A(A[236]), .B(n271), .Z(n270) );
  NANDN U291 ( .A(n271), .B(A[236]), .Z(n268) );
  XOR U292 ( .A(n271), .B(n272), .Z(SUM[236]) );
  XNOR U293 ( .A(B[236]), .B(A[236]), .Z(n272) );
  AND U294 ( .A(n273), .B(n274), .Z(n271) );
  NAND U295 ( .A(B[235]), .B(n275), .Z(n274) );
  NANDN U296 ( .A(A[235]), .B(n276), .Z(n275) );
  NANDN U297 ( .A(n276), .B(A[235]), .Z(n273) );
  XOR U298 ( .A(n276), .B(n277), .Z(SUM[235]) );
  XNOR U299 ( .A(B[235]), .B(A[235]), .Z(n277) );
  AND U300 ( .A(n278), .B(n279), .Z(n276) );
  NAND U301 ( .A(B[234]), .B(n280), .Z(n279) );
  NANDN U302 ( .A(A[234]), .B(n281), .Z(n280) );
  NANDN U303 ( .A(n281), .B(A[234]), .Z(n278) );
  XOR U304 ( .A(n281), .B(n282), .Z(SUM[234]) );
  XNOR U305 ( .A(B[234]), .B(A[234]), .Z(n282) );
  AND U306 ( .A(n283), .B(n284), .Z(n281) );
  NAND U307 ( .A(B[233]), .B(n285), .Z(n284) );
  NANDN U308 ( .A(A[233]), .B(n286), .Z(n285) );
  NANDN U309 ( .A(n286), .B(A[233]), .Z(n283) );
  XOR U310 ( .A(n286), .B(n287), .Z(SUM[233]) );
  XNOR U311 ( .A(B[233]), .B(A[233]), .Z(n287) );
  AND U312 ( .A(n288), .B(n289), .Z(n286) );
  NAND U313 ( .A(B[232]), .B(n290), .Z(n289) );
  NANDN U314 ( .A(A[232]), .B(n291), .Z(n290) );
  NANDN U315 ( .A(n291), .B(A[232]), .Z(n288) );
  XOR U316 ( .A(n291), .B(n292), .Z(SUM[232]) );
  XNOR U317 ( .A(B[232]), .B(A[232]), .Z(n292) );
  AND U318 ( .A(n293), .B(n294), .Z(n291) );
  NAND U319 ( .A(B[231]), .B(n295), .Z(n294) );
  NANDN U320 ( .A(A[231]), .B(n296), .Z(n295) );
  NANDN U321 ( .A(n296), .B(A[231]), .Z(n293) );
  XOR U322 ( .A(n296), .B(n297), .Z(SUM[231]) );
  XNOR U323 ( .A(B[231]), .B(A[231]), .Z(n297) );
  AND U324 ( .A(n298), .B(n299), .Z(n296) );
  NAND U325 ( .A(B[230]), .B(n300), .Z(n299) );
  NANDN U326 ( .A(A[230]), .B(n301), .Z(n300) );
  NANDN U327 ( .A(n301), .B(A[230]), .Z(n298) );
  XOR U328 ( .A(n301), .B(n302), .Z(SUM[230]) );
  XNOR U329 ( .A(B[230]), .B(A[230]), .Z(n302) );
  AND U330 ( .A(n303), .B(n304), .Z(n301) );
  NAND U331 ( .A(B[229]), .B(n305), .Z(n304) );
  NANDN U332 ( .A(A[229]), .B(n306), .Z(n305) );
  NANDN U333 ( .A(n306), .B(A[229]), .Z(n303) );
  XOR U334 ( .A(n307), .B(n308), .Z(SUM[22]) );
  XNOR U335 ( .A(B[22]), .B(A[22]), .Z(n308) );
  XOR U336 ( .A(n306), .B(n309), .Z(SUM[229]) );
  XNOR U337 ( .A(B[229]), .B(A[229]), .Z(n309) );
  AND U338 ( .A(n310), .B(n311), .Z(n306) );
  NAND U339 ( .A(B[228]), .B(n312), .Z(n311) );
  NANDN U340 ( .A(A[228]), .B(n313), .Z(n312) );
  NANDN U341 ( .A(n313), .B(A[228]), .Z(n310) );
  XOR U342 ( .A(n313), .B(n314), .Z(SUM[228]) );
  XNOR U343 ( .A(B[228]), .B(A[228]), .Z(n314) );
  AND U344 ( .A(n315), .B(n316), .Z(n313) );
  NAND U345 ( .A(B[227]), .B(n317), .Z(n316) );
  NANDN U346 ( .A(A[227]), .B(n318), .Z(n317) );
  NANDN U347 ( .A(n318), .B(A[227]), .Z(n315) );
  XOR U348 ( .A(n318), .B(n319), .Z(SUM[227]) );
  XNOR U349 ( .A(B[227]), .B(A[227]), .Z(n319) );
  AND U350 ( .A(n320), .B(n321), .Z(n318) );
  NAND U351 ( .A(B[226]), .B(n322), .Z(n321) );
  NANDN U352 ( .A(A[226]), .B(n323), .Z(n322) );
  NANDN U353 ( .A(n323), .B(A[226]), .Z(n320) );
  XOR U354 ( .A(n323), .B(n324), .Z(SUM[226]) );
  XNOR U355 ( .A(B[226]), .B(A[226]), .Z(n324) );
  AND U356 ( .A(n325), .B(n326), .Z(n323) );
  NAND U357 ( .A(B[225]), .B(n327), .Z(n326) );
  NANDN U358 ( .A(A[225]), .B(n328), .Z(n327) );
  NANDN U359 ( .A(n328), .B(A[225]), .Z(n325) );
  XOR U360 ( .A(n328), .B(n329), .Z(SUM[225]) );
  XNOR U361 ( .A(B[225]), .B(A[225]), .Z(n329) );
  AND U362 ( .A(n330), .B(n331), .Z(n328) );
  NAND U363 ( .A(B[224]), .B(n332), .Z(n331) );
  NANDN U364 ( .A(A[224]), .B(n333), .Z(n332) );
  NANDN U365 ( .A(n333), .B(A[224]), .Z(n330) );
  XOR U366 ( .A(n333), .B(n334), .Z(SUM[224]) );
  XNOR U367 ( .A(B[224]), .B(A[224]), .Z(n334) );
  AND U368 ( .A(n335), .B(n336), .Z(n333) );
  NAND U369 ( .A(B[223]), .B(n337), .Z(n336) );
  NANDN U370 ( .A(A[223]), .B(n338), .Z(n337) );
  NANDN U371 ( .A(n338), .B(A[223]), .Z(n335) );
  XOR U372 ( .A(n338), .B(n339), .Z(SUM[223]) );
  XNOR U373 ( .A(B[223]), .B(A[223]), .Z(n339) );
  AND U374 ( .A(n340), .B(n341), .Z(n338) );
  NAND U375 ( .A(B[222]), .B(n342), .Z(n341) );
  NANDN U376 ( .A(A[222]), .B(n343), .Z(n342) );
  NANDN U377 ( .A(n343), .B(A[222]), .Z(n340) );
  XOR U378 ( .A(n343), .B(n344), .Z(SUM[222]) );
  XNOR U379 ( .A(B[222]), .B(A[222]), .Z(n344) );
  AND U380 ( .A(n345), .B(n346), .Z(n343) );
  NAND U381 ( .A(B[221]), .B(n347), .Z(n346) );
  NANDN U382 ( .A(A[221]), .B(n348), .Z(n347) );
  NANDN U383 ( .A(n348), .B(A[221]), .Z(n345) );
  XOR U384 ( .A(n348), .B(n349), .Z(SUM[221]) );
  XNOR U385 ( .A(B[221]), .B(A[221]), .Z(n349) );
  AND U386 ( .A(n350), .B(n351), .Z(n348) );
  NAND U387 ( .A(B[220]), .B(n352), .Z(n351) );
  NANDN U388 ( .A(A[220]), .B(n353), .Z(n352) );
  NANDN U389 ( .A(n353), .B(A[220]), .Z(n350) );
  XOR U390 ( .A(n353), .B(n354), .Z(SUM[220]) );
  XNOR U391 ( .A(B[220]), .B(A[220]), .Z(n354) );
  AND U392 ( .A(n355), .B(n356), .Z(n353) );
  NAND U393 ( .A(B[219]), .B(n357), .Z(n356) );
  NANDN U394 ( .A(A[219]), .B(n358), .Z(n357) );
  NANDN U395 ( .A(n358), .B(A[219]), .Z(n355) );
  XOR U396 ( .A(n359), .B(n360), .Z(SUM[21]) );
  XNOR U397 ( .A(B[21]), .B(A[21]), .Z(n360) );
  XOR U398 ( .A(n358), .B(n361), .Z(SUM[219]) );
  XNOR U399 ( .A(B[219]), .B(A[219]), .Z(n361) );
  AND U400 ( .A(n362), .B(n363), .Z(n358) );
  NAND U401 ( .A(B[218]), .B(n364), .Z(n363) );
  NANDN U402 ( .A(A[218]), .B(n365), .Z(n364) );
  NANDN U403 ( .A(n365), .B(A[218]), .Z(n362) );
  XOR U404 ( .A(n365), .B(n366), .Z(SUM[218]) );
  XNOR U405 ( .A(B[218]), .B(A[218]), .Z(n366) );
  AND U406 ( .A(n367), .B(n368), .Z(n365) );
  NAND U407 ( .A(B[217]), .B(n369), .Z(n368) );
  NANDN U408 ( .A(A[217]), .B(n370), .Z(n369) );
  NANDN U409 ( .A(n370), .B(A[217]), .Z(n367) );
  XOR U410 ( .A(n370), .B(n371), .Z(SUM[217]) );
  XNOR U411 ( .A(B[217]), .B(A[217]), .Z(n371) );
  AND U412 ( .A(n372), .B(n373), .Z(n370) );
  NAND U413 ( .A(B[216]), .B(n374), .Z(n373) );
  NANDN U414 ( .A(A[216]), .B(n375), .Z(n374) );
  NANDN U415 ( .A(n375), .B(A[216]), .Z(n372) );
  XOR U416 ( .A(n375), .B(n376), .Z(SUM[216]) );
  XNOR U417 ( .A(B[216]), .B(A[216]), .Z(n376) );
  AND U418 ( .A(n377), .B(n378), .Z(n375) );
  NAND U419 ( .A(B[215]), .B(n379), .Z(n378) );
  NANDN U420 ( .A(A[215]), .B(n380), .Z(n379) );
  NANDN U421 ( .A(n380), .B(A[215]), .Z(n377) );
  XOR U422 ( .A(n380), .B(n381), .Z(SUM[215]) );
  XNOR U423 ( .A(B[215]), .B(A[215]), .Z(n381) );
  AND U424 ( .A(n382), .B(n383), .Z(n380) );
  NAND U425 ( .A(B[214]), .B(n384), .Z(n383) );
  NANDN U426 ( .A(A[214]), .B(n385), .Z(n384) );
  NANDN U427 ( .A(n385), .B(A[214]), .Z(n382) );
  XOR U428 ( .A(n385), .B(n386), .Z(SUM[214]) );
  XNOR U429 ( .A(B[214]), .B(A[214]), .Z(n386) );
  AND U430 ( .A(n387), .B(n388), .Z(n385) );
  NAND U431 ( .A(B[213]), .B(n389), .Z(n388) );
  NANDN U432 ( .A(A[213]), .B(n390), .Z(n389) );
  NANDN U433 ( .A(n390), .B(A[213]), .Z(n387) );
  XOR U434 ( .A(n390), .B(n391), .Z(SUM[213]) );
  XNOR U435 ( .A(B[213]), .B(A[213]), .Z(n391) );
  AND U436 ( .A(n392), .B(n393), .Z(n390) );
  NAND U437 ( .A(B[212]), .B(n394), .Z(n393) );
  NANDN U438 ( .A(A[212]), .B(n395), .Z(n394) );
  NANDN U439 ( .A(n395), .B(A[212]), .Z(n392) );
  XOR U440 ( .A(n395), .B(n396), .Z(SUM[212]) );
  XNOR U441 ( .A(B[212]), .B(A[212]), .Z(n396) );
  AND U442 ( .A(n397), .B(n398), .Z(n395) );
  NAND U443 ( .A(B[211]), .B(n399), .Z(n398) );
  NANDN U444 ( .A(A[211]), .B(n400), .Z(n399) );
  NANDN U445 ( .A(n400), .B(A[211]), .Z(n397) );
  XOR U446 ( .A(n400), .B(n401), .Z(SUM[211]) );
  XNOR U447 ( .A(B[211]), .B(A[211]), .Z(n401) );
  AND U448 ( .A(n402), .B(n403), .Z(n400) );
  NAND U449 ( .A(B[210]), .B(n404), .Z(n403) );
  NANDN U450 ( .A(A[210]), .B(n405), .Z(n404) );
  NANDN U451 ( .A(n405), .B(A[210]), .Z(n402) );
  XOR U452 ( .A(n405), .B(n406), .Z(SUM[210]) );
  XNOR U453 ( .A(B[210]), .B(A[210]), .Z(n406) );
  AND U454 ( .A(n407), .B(n408), .Z(n405) );
  NAND U455 ( .A(B[209]), .B(n409), .Z(n408) );
  NANDN U456 ( .A(A[209]), .B(n410), .Z(n409) );
  NANDN U457 ( .A(n410), .B(A[209]), .Z(n407) );
  XOR U458 ( .A(n411), .B(n412), .Z(SUM[20]) );
  XNOR U459 ( .A(B[20]), .B(A[20]), .Z(n412) );
  XOR U460 ( .A(n410), .B(n413), .Z(SUM[209]) );
  XNOR U461 ( .A(B[209]), .B(A[209]), .Z(n413) );
  AND U462 ( .A(n414), .B(n415), .Z(n410) );
  NAND U463 ( .A(B[208]), .B(n416), .Z(n415) );
  NANDN U464 ( .A(A[208]), .B(n417), .Z(n416) );
  NANDN U465 ( .A(n417), .B(A[208]), .Z(n414) );
  XOR U466 ( .A(n417), .B(n418), .Z(SUM[208]) );
  XNOR U467 ( .A(B[208]), .B(A[208]), .Z(n418) );
  AND U468 ( .A(n419), .B(n420), .Z(n417) );
  NAND U469 ( .A(B[207]), .B(n421), .Z(n420) );
  NANDN U470 ( .A(A[207]), .B(n422), .Z(n421) );
  NANDN U471 ( .A(n422), .B(A[207]), .Z(n419) );
  XOR U472 ( .A(n422), .B(n423), .Z(SUM[207]) );
  XNOR U473 ( .A(B[207]), .B(A[207]), .Z(n423) );
  AND U474 ( .A(n424), .B(n425), .Z(n422) );
  NAND U475 ( .A(B[206]), .B(n426), .Z(n425) );
  NANDN U476 ( .A(A[206]), .B(n427), .Z(n426) );
  NANDN U477 ( .A(n427), .B(A[206]), .Z(n424) );
  XOR U478 ( .A(n427), .B(n428), .Z(SUM[206]) );
  XNOR U479 ( .A(B[206]), .B(A[206]), .Z(n428) );
  AND U480 ( .A(n429), .B(n430), .Z(n427) );
  NAND U481 ( .A(B[205]), .B(n431), .Z(n430) );
  NANDN U482 ( .A(A[205]), .B(n432), .Z(n431) );
  NANDN U483 ( .A(n432), .B(A[205]), .Z(n429) );
  XOR U484 ( .A(n432), .B(n433), .Z(SUM[205]) );
  XNOR U485 ( .A(B[205]), .B(A[205]), .Z(n433) );
  AND U486 ( .A(n434), .B(n435), .Z(n432) );
  NAND U487 ( .A(B[204]), .B(n436), .Z(n435) );
  NANDN U488 ( .A(A[204]), .B(n437), .Z(n436) );
  NANDN U489 ( .A(n437), .B(A[204]), .Z(n434) );
  XOR U490 ( .A(n437), .B(n438), .Z(SUM[204]) );
  XNOR U491 ( .A(B[204]), .B(A[204]), .Z(n438) );
  AND U492 ( .A(n439), .B(n440), .Z(n437) );
  NAND U493 ( .A(B[203]), .B(n441), .Z(n440) );
  NANDN U494 ( .A(A[203]), .B(n442), .Z(n441) );
  NANDN U495 ( .A(n442), .B(A[203]), .Z(n439) );
  XOR U496 ( .A(n442), .B(n443), .Z(SUM[203]) );
  XNOR U497 ( .A(B[203]), .B(A[203]), .Z(n443) );
  AND U498 ( .A(n444), .B(n445), .Z(n442) );
  NAND U499 ( .A(B[202]), .B(n446), .Z(n445) );
  NANDN U500 ( .A(A[202]), .B(n447), .Z(n446) );
  NANDN U501 ( .A(n447), .B(A[202]), .Z(n444) );
  XOR U502 ( .A(n447), .B(n448), .Z(SUM[202]) );
  XNOR U503 ( .A(B[202]), .B(A[202]), .Z(n448) );
  AND U504 ( .A(n449), .B(n450), .Z(n447) );
  NAND U505 ( .A(B[201]), .B(n451), .Z(n450) );
  NANDN U506 ( .A(A[201]), .B(n452), .Z(n451) );
  NANDN U507 ( .A(n452), .B(A[201]), .Z(n449) );
  XOR U508 ( .A(n452), .B(n453), .Z(SUM[201]) );
  XNOR U509 ( .A(B[201]), .B(A[201]), .Z(n453) );
  AND U510 ( .A(n454), .B(n455), .Z(n452) );
  NAND U511 ( .A(B[200]), .B(n456), .Z(n455) );
  NANDN U512 ( .A(A[200]), .B(n457), .Z(n456) );
  NANDN U513 ( .A(n457), .B(A[200]), .Z(n454) );
  XOR U514 ( .A(n457), .B(n458), .Z(SUM[200]) );
  XNOR U515 ( .A(B[200]), .B(A[200]), .Z(n458) );
  AND U516 ( .A(n459), .B(n460), .Z(n457) );
  NAND U517 ( .A(B[199]), .B(n461), .Z(n460) );
  NANDN U518 ( .A(A[199]), .B(n462), .Z(n461) );
  NANDN U519 ( .A(n462), .B(A[199]), .Z(n459) );
  XOR U520 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  XOR U521 ( .A(n463), .B(n464), .Z(SUM[19]) );
  XNOR U522 ( .A(B[19]), .B(A[19]), .Z(n464) );
  XOR U523 ( .A(n462), .B(n465), .Z(SUM[199]) );
  XNOR U524 ( .A(B[199]), .B(A[199]), .Z(n465) );
  AND U525 ( .A(n466), .B(n467), .Z(n462) );
  NAND U526 ( .A(B[198]), .B(n468), .Z(n467) );
  NANDN U527 ( .A(A[198]), .B(n469), .Z(n468) );
  NANDN U528 ( .A(n469), .B(A[198]), .Z(n466) );
  XOR U529 ( .A(n469), .B(n470), .Z(SUM[198]) );
  XNOR U530 ( .A(B[198]), .B(A[198]), .Z(n470) );
  AND U531 ( .A(n471), .B(n472), .Z(n469) );
  NAND U532 ( .A(B[197]), .B(n473), .Z(n472) );
  NANDN U533 ( .A(A[197]), .B(n474), .Z(n473) );
  NANDN U534 ( .A(n474), .B(A[197]), .Z(n471) );
  XOR U535 ( .A(n474), .B(n475), .Z(SUM[197]) );
  XNOR U536 ( .A(B[197]), .B(A[197]), .Z(n475) );
  AND U537 ( .A(n476), .B(n477), .Z(n474) );
  NAND U538 ( .A(B[196]), .B(n478), .Z(n477) );
  NANDN U539 ( .A(A[196]), .B(n479), .Z(n478) );
  NANDN U540 ( .A(n479), .B(A[196]), .Z(n476) );
  XOR U541 ( .A(n479), .B(n480), .Z(SUM[196]) );
  XNOR U542 ( .A(B[196]), .B(A[196]), .Z(n480) );
  AND U543 ( .A(n481), .B(n482), .Z(n479) );
  NAND U544 ( .A(B[195]), .B(n483), .Z(n482) );
  NANDN U545 ( .A(A[195]), .B(n484), .Z(n483) );
  NANDN U546 ( .A(n484), .B(A[195]), .Z(n481) );
  XOR U547 ( .A(n484), .B(n485), .Z(SUM[195]) );
  XNOR U548 ( .A(B[195]), .B(A[195]), .Z(n485) );
  AND U549 ( .A(n486), .B(n487), .Z(n484) );
  NAND U550 ( .A(B[194]), .B(n488), .Z(n487) );
  NANDN U551 ( .A(A[194]), .B(n489), .Z(n488) );
  NANDN U552 ( .A(n489), .B(A[194]), .Z(n486) );
  XOR U553 ( .A(n489), .B(n490), .Z(SUM[194]) );
  XNOR U554 ( .A(B[194]), .B(A[194]), .Z(n490) );
  AND U555 ( .A(n491), .B(n492), .Z(n489) );
  NAND U556 ( .A(B[193]), .B(n493), .Z(n492) );
  NANDN U557 ( .A(A[193]), .B(n494), .Z(n493) );
  NANDN U558 ( .A(n494), .B(A[193]), .Z(n491) );
  XOR U559 ( .A(n494), .B(n495), .Z(SUM[193]) );
  XNOR U560 ( .A(B[193]), .B(A[193]), .Z(n495) );
  AND U561 ( .A(n496), .B(n497), .Z(n494) );
  NAND U562 ( .A(B[192]), .B(n498), .Z(n497) );
  NANDN U563 ( .A(A[192]), .B(n499), .Z(n498) );
  NANDN U564 ( .A(n499), .B(A[192]), .Z(n496) );
  XOR U565 ( .A(n499), .B(n500), .Z(SUM[192]) );
  XNOR U566 ( .A(B[192]), .B(A[192]), .Z(n500) );
  AND U567 ( .A(n501), .B(n502), .Z(n499) );
  NAND U568 ( .A(B[191]), .B(n503), .Z(n502) );
  NANDN U569 ( .A(A[191]), .B(n504), .Z(n503) );
  NANDN U570 ( .A(n504), .B(A[191]), .Z(n501) );
  XOR U571 ( .A(n504), .B(n505), .Z(SUM[191]) );
  XNOR U572 ( .A(B[191]), .B(A[191]), .Z(n505) );
  AND U573 ( .A(n506), .B(n507), .Z(n504) );
  NAND U574 ( .A(B[190]), .B(n508), .Z(n507) );
  NANDN U575 ( .A(A[190]), .B(n509), .Z(n508) );
  NANDN U576 ( .A(n509), .B(A[190]), .Z(n506) );
  XOR U577 ( .A(n509), .B(n510), .Z(SUM[190]) );
  XNOR U578 ( .A(B[190]), .B(A[190]), .Z(n510) );
  AND U579 ( .A(n511), .B(n512), .Z(n509) );
  NAND U580 ( .A(B[189]), .B(n513), .Z(n512) );
  NANDN U581 ( .A(A[189]), .B(n514), .Z(n513) );
  NANDN U582 ( .A(n514), .B(A[189]), .Z(n511) );
  XOR U583 ( .A(n515), .B(n516), .Z(SUM[18]) );
  XNOR U584 ( .A(B[18]), .B(A[18]), .Z(n516) );
  XOR U585 ( .A(n514), .B(n517), .Z(SUM[189]) );
  XNOR U586 ( .A(B[189]), .B(A[189]), .Z(n517) );
  AND U587 ( .A(n518), .B(n519), .Z(n514) );
  NAND U588 ( .A(B[188]), .B(n520), .Z(n519) );
  NANDN U589 ( .A(A[188]), .B(n521), .Z(n520) );
  NANDN U590 ( .A(n521), .B(A[188]), .Z(n518) );
  XOR U591 ( .A(n521), .B(n522), .Z(SUM[188]) );
  XNOR U592 ( .A(B[188]), .B(A[188]), .Z(n522) );
  AND U593 ( .A(n523), .B(n524), .Z(n521) );
  NAND U594 ( .A(B[187]), .B(n525), .Z(n524) );
  NANDN U595 ( .A(A[187]), .B(n526), .Z(n525) );
  NANDN U596 ( .A(n526), .B(A[187]), .Z(n523) );
  XOR U597 ( .A(n526), .B(n527), .Z(SUM[187]) );
  XNOR U598 ( .A(B[187]), .B(A[187]), .Z(n527) );
  AND U599 ( .A(n528), .B(n529), .Z(n526) );
  NAND U600 ( .A(B[186]), .B(n530), .Z(n529) );
  NANDN U601 ( .A(A[186]), .B(n531), .Z(n530) );
  NANDN U602 ( .A(n531), .B(A[186]), .Z(n528) );
  XOR U603 ( .A(n531), .B(n532), .Z(SUM[186]) );
  XNOR U604 ( .A(B[186]), .B(A[186]), .Z(n532) );
  AND U605 ( .A(n533), .B(n534), .Z(n531) );
  NAND U606 ( .A(B[185]), .B(n535), .Z(n534) );
  NANDN U607 ( .A(A[185]), .B(n536), .Z(n535) );
  NANDN U608 ( .A(n536), .B(A[185]), .Z(n533) );
  XOR U609 ( .A(n536), .B(n537), .Z(SUM[185]) );
  XNOR U610 ( .A(B[185]), .B(A[185]), .Z(n537) );
  AND U611 ( .A(n538), .B(n539), .Z(n536) );
  NAND U612 ( .A(B[184]), .B(n540), .Z(n539) );
  NANDN U613 ( .A(A[184]), .B(n541), .Z(n540) );
  NANDN U614 ( .A(n541), .B(A[184]), .Z(n538) );
  XOR U615 ( .A(n541), .B(n542), .Z(SUM[184]) );
  XNOR U616 ( .A(B[184]), .B(A[184]), .Z(n542) );
  AND U617 ( .A(n543), .B(n544), .Z(n541) );
  NAND U618 ( .A(B[183]), .B(n545), .Z(n544) );
  NANDN U619 ( .A(A[183]), .B(n546), .Z(n545) );
  NANDN U620 ( .A(n546), .B(A[183]), .Z(n543) );
  XOR U621 ( .A(n546), .B(n547), .Z(SUM[183]) );
  XNOR U622 ( .A(B[183]), .B(A[183]), .Z(n547) );
  AND U623 ( .A(n548), .B(n549), .Z(n546) );
  NAND U624 ( .A(B[182]), .B(n550), .Z(n549) );
  NANDN U625 ( .A(A[182]), .B(n551), .Z(n550) );
  NANDN U626 ( .A(n551), .B(A[182]), .Z(n548) );
  XOR U627 ( .A(n551), .B(n552), .Z(SUM[182]) );
  XNOR U628 ( .A(B[182]), .B(A[182]), .Z(n552) );
  AND U629 ( .A(n553), .B(n554), .Z(n551) );
  NAND U630 ( .A(B[181]), .B(n555), .Z(n554) );
  NANDN U631 ( .A(A[181]), .B(n556), .Z(n555) );
  NANDN U632 ( .A(n556), .B(A[181]), .Z(n553) );
  XOR U633 ( .A(n556), .B(n557), .Z(SUM[181]) );
  XNOR U634 ( .A(B[181]), .B(A[181]), .Z(n557) );
  AND U635 ( .A(n558), .B(n559), .Z(n556) );
  NAND U636 ( .A(B[180]), .B(n560), .Z(n559) );
  NANDN U637 ( .A(A[180]), .B(n561), .Z(n560) );
  NANDN U638 ( .A(n561), .B(A[180]), .Z(n558) );
  XOR U639 ( .A(n561), .B(n562), .Z(SUM[180]) );
  XNOR U640 ( .A(B[180]), .B(A[180]), .Z(n562) );
  AND U641 ( .A(n563), .B(n564), .Z(n561) );
  NAND U642 ( .A(B[179]), .B(n565), .Z(n564) );
  NANDN U643 ( .A(A[179]), .B(n566), .Z(n565) );
  NANDN U644 ( .A(n566), .B(A[179]), .Z(n563) );
  XOR U645 ( .A(n567), .B(n568), .Z(SUM[17]) );
  XNOR U646 ( .A(B[17]), .B(A[17]), .Z(n568) );
  XOR U647 ( .A(n566), .B(n569), .Z(SUM[179]) );
  XNOR U648 ( .A(B[179]), .B(A[179]), .Z(n569) );
  AND U649 ( .A(n570), .B(n571), .Z(n566) );
  NAND U650 ( .A(B[178]), .B(n572), .Z(n571) );
  NANDN U651 ( .A(A[178]), .B(n573), .Z(n572) );
  NANDN U652 ( .A(n573), .B(A[178]), .Z(n570) );
  XOR U653 ( .A(n573), .B(n574), .Z(SUM[178]) );
  XNOR U654 ( .A(B[178]), .B(A[178]), .Z(n574) );
  AND U655 ( .A(n575), .B(n576), .Z(n573) );
  NAND U656 ( .A(B[177]), .B(n577), .Z(n576) );
  NANDN U657 ( .A(A[177]), .B(n578), .Z(n577) );
  NANDN U658 ( .A(n578), .B(A[177]), .Z(n575) );
  XOR U659 ( .A(n578), .B(n579), .Z(SUM[177]) );
  XNOR U660 ( .A(B[177]), .B(A[177]), .Z(n579) );
  AND U661 ( .A(n580), .B(n581), .Z(n578) );
  NAND U662 ( .A(B[176]), .B(n582), .Z(n581) );
  NANDN U663 ( .A(A[176]), .B(n583), .Z(n582) );
  NANDN U664 ( .A(n583), .B(A[176]), .Z(n580) );
  XOR U665 ( .A(n583), .B(n584), .Z(SUM[176]) );
  XNOR U666 ( .A(B[176]), .B(A[176]), .Z(n584) );
  AND U667 ( .A(n585), .B(n586), .Z(n583) );
  NAND U668 ( .A(B[175]), .B(n587), .Z(n586) );
  NANDN U669 ( .A(A[175]), .B(n588), .Z(n587) );
  NANDN U670 ( .A(n588), .B(A[175]), .Z(n585) );
  XOR U671 ( .A(n588), .B(n589), .Z(SUM[175]) );
  XNOR U672 ( .A(B[175]), .B(A[175]), .Z(n589) );
  AND U673 ( .A(n590), .B(n591), .Z(n588) );
  NAND U674 ( .A(B[174]), .B(n592), .Z(n591) );
  NANDN U675 ( .A(A[174]), .B(n593), .Z(n592) );
  NANDN U676 ( .A(n593), .B(A[174]), .Z(n590) );
  XOR U677 ( .A(n593), .B(n594), .Z(SUM[174]) );
  XNOR U678 ( .A(B[174]), .B(A[174]), .Z(n594) );
  AND U679 ( .A(n595), .B(n596), .Z(n593) );
  NAND U680 ( .A(B[173]), .B(n597), .Z(n596) );
  NANDN U681 ( .A(A[173]), .B(n598), .Z(n597) );
  NANDN U682 ( .A(n598), .B(A[173]), .Z(n595) );
  XOR U683 ( .A(n598), .B(n599), .Z(SUM[173]) );
  XNOR U684 ( .A(B[173]), .B(A[173]), .Z(n599) );
  AND U685 ( .A(n600), .B(n601), .Z(n598) );
  NAND U686 ( .A(B[172]), .B(n602), .Z(n601) );
  NANDN U687 ( .A(A[172]), .B(n603), .Z(n602) );
  NANDN U688 ( .A(n603), .B(A[172]), .Z(n600) );
  XOR U689 ( .A(n603), .B(n604), .Z(SUM[172]) );
  XNOR U690 ( .A(B[172]), .B(A[172]), .Z(n604) );
  AND U691 ( .A(n605), .B(n606), .Z(n603) );
  NAND U692 ( .A(B[171]), .B(n607), .Z(n606) );
  NANDN U693 ( .A(A[171]), .B(n608), .Z(n607) );
  NANDN U694 ( .A(n608), .B(A[171]), .Z(n605) );
  XOR U695 ( .A(n608), .B(n609), .Z(SUM[171]) );
  XNOR U696 ( .A(B[171]), .B(A[171]), .Z(n609) );
  AND U697 ( .A(n610), .B(n611), .Z(n608) );
  NAND U698 ( .A(B[170]), .B(n612), .Z(n611) );
  NANDN U699 ( .A(A[170]), .B(n613), .Z(n612) );
  NANDN U700 ( .A(n613), .B(A[170]), .Z(n610) );
  XOR U701 ( .A(n613), .B(n614), .Z(SUM[170]) );
  XNOR U702 ( .A(B[170]), .B(A[170]), .Z(n614) );
  AND U703 ( .A(n615), .B(n616), .Z(n613) );
  NAND U704 ( .A(B[169]), .B(n617), .Z(n616) );
  NANDN U705 ( .A(A[169]), .B(n618), .Z(n617) );
  NANDN U706 ( .A(n618), .B(A[169]), .Z(n615) );
  XOR U707 ( .A(n619), .B(n620), .Z(SUM[16]) );
  XNOR U708 ( .A(B[16]), .B(A[16]), .Z(n620) );
  XOR U709 ( .A(n618), .B(n621), .Z(SUM[169]) );
  XNOR U710 ( .A(B[169]), .B(A[169]), .Z(n621) );
  AND U711 ( .A(n622), .B(n623), .Z(n618) );
  NAND U712 ( .A(B[168]), .B(n624), .Z(n623) );
  NANDN U713 ( .A(A[168]), .B(n625), .Z(n624) );
  NANDN U714 ( .A(n625), .B(A[168]), .Z(n622) );
  XOR U715 ( .A(n625), .B(n626), .Z(SUM[168]) );
  XNOR U716 ( .A(B[168]), .B(A[168]), .Z(n626) );
  AND U717 ( .A(n627), .B(n628), .Z(n625) );
  NAND U718 ( .A(B[167]), .B(n629), .Z(n628) );
  NANDN U719 ( .A(A[167]), .B(n630), .Z(n629) );
  NANDN U720 ( .A(n630), .B(A[167]), .Z(n627) );
  XOR U721 ( .A(n630), .B(n631), .Z(SUM[167]) );
  XNOR U722 ( .A(B[167]), .B(A[167]), .Z(n631) );
  AND U723 ( .A(n632), .B(n633), .Z(n630) );
  NAND U724 ( .A(B[166]), .B(n634), .Z(n633) );
  NANDN U725 ( .A(A[166]), .B(n635), .Z(n634) );
  NANDN U726 ( .A(n635), .B(A[166]), .Z(n632) );
  XOR U727 ( .A(n635), .B(n636), .Z(SUM[166]) );
  XNOR U728 ( .A(B[166]), .B(A[166]), .Z(n636) );
  AND U729 ( .A(n637), .B(n638), .Z(n635) );
  NAND U730 ( .A(B[165]), .B(n639), .Z(n638) );
  NANDN U731 ( .A(A[165]), .B(n640), .Z(n639) );
  NANDN U732 ( .A(n640), .B(A[165]), .Z(n637) );
  XOR U733 ( .A(n640), .B(n641), .Z(SUM[165]) );
  XNOR U734 ( .A(B[165]), .B(A[165]), .Z(n641) );
  AND U735 ( .A(n642), .B(n643), .Z(n640) );
  NAND U736 ( .A(B[164]), .B(n644), .Z(n643) );
  NANDN U737 ( .A(A[164]), .B(n645), .Z(n644) );
  NANDN U738 ( .A(n645), .B(A[164]), .Z(n642) );
  XOR U739 ( .A(n645), .B(n646), .Z(SUM[164]) );
  XNOR U740 ( .A(B[164]), .B(A[164]), .Z(n646) );
  AND U741 ( .A(n647), .B(n648), .Z(n645) );
  NAND U742 ( .A(B[163]), .B(n649), .Z(n648) );
  NANDN U743 ( .A(A[163]), .B(n650), .Z(n649) );
  NANDN U744 ( .A(n650), .B(A[163]), .Z(n647) );
  XOR U745 ( .A(n650), .B(n651), .Z(SUM[163]) );
  XNOR U746 ( .A(B[163]), .B(A[163]), .Z(n651) );
  AND U747 ( .A(n652), .B(n653), .Z(n650) );
  NAND U748 ( .A(B[162]), .B(n654), .Z(n653) );
  NANDN U749 ( .A(A[162]), .B(n655), .Z(n654) );
  NANDN U750 ( .A(n655), .B(A[162]), .Z(n652) );
  XOR U751 ( .A(n655), .B(n656), .Z(SUM[162]) );
  XNOR U752 ( .A(B[162]), .B(A[162]), .Z(n656) );
  AND U753 ( .A(n657), .B(n658), .Z(n655) );
  NAND U754 ( .A(B[161]), .B(n659), .Z(n658) );
  NANDN U755 ( .A(A[161]), .B(n660), .Z(n659) );
  NANDN U756 ( .A(n660), .B(A[161]), .Z(n657) );
  XOR U757 ( .A(n660), .B(n661), .Z(SUM[161]) );
  XNOR U758 ( .A(B[161]), .B(A[161]), .Z(n661) );
  AND U759 ( .A(n662), .B(n663), .Z(n660) );
  NAND U760 ( .A(B[160]), .B(n664), .Z(n663) );
  NANDN U761 ( .A(A[160]), .B(n665), .Z(n664) );
  NANDN U762 ( .A(n665), .B(A[160]), .Z(n662) );
  XOR U763 ( .A(n665), .B(n666), .Z(SUM[160]) );
  XNOR U764 ( .A(B[160]), .B(A[160]), .Z(n666) );
  AND U765 ( .A(n667), .B(n668), .Z(n665) );
  NAND U766 ( .A(B[159]), .B(n669), .Z(n668) );
  NANDN U767 ( .A(A[159]), .B(n670), .Z(n669) );
  NANDN U768 ( .A(n670), .B(A[159]), .Z(n667) );
  XOR U769 ( .A(n671), .B(n672), .Z(SUM[15]) );
  XNOR U770 ( .A(B[15]), .B(A[15]), .Z(n672) );
  XOR U771 ( .A(n670), .B(n673), .Z(SUM[159]) );
  XNOR U772 ( .A(B[159]), .B(A[159]), .Z(n673) );
  AND U773 ( .A(n674), .B(n675), .Z(n670) );
  NAND U774 ( .A(B[158]), .B(n676), .Z(n675) );
  NANDN U775 ( .A(A[158]), .B(n677), .Z(n676) );
  NANDN U776 ( .A(n677), .B(A[158]), .Z(n674) );
  XOR U777 ( .A(n677), .B(n678), .Z(SUM[158]) );
  XNOR U778 ( .A(B[158]), .B(A[158]), .Z(n678) );
  AND U779 ( .A(n679), .B(n680), .Z(n677) );
  NAND U780 ( .A(B[157]), .B(n681), .Z(n680) );
  NANDN U781 ( .A(A[157]), .B(n682), .Z(n681) );
  NANDN U782 ( .A(n682), .B(A[157]), .Z(n679) );
  XOR U783 ( .A(n682), .B(n683), .Z(SUM[157]) );
  XNOR U784 ( .A(B[157]), .B(A[157]), .Z(n683) );
  AND U785 ( .A(n684), .B(n685), .Z(n682) );
  NAND U786 ( .A(B[156]), .B(n686), .Z(n685) );
  NANDN U787 ( .A(A[156]), .B(n687), .Z(n686) );
  NANDN U788 ( .A(n687), .B(A[156]), .Z(n684) );
  XOR U789 ( .A(n687), .B(n688), .Z(SUM[156]) );
  XNOR U790 ( .A(B[156]), .B(A[156]), .Z(n688) );
  AND U791 ( .A(n689), .B(n690), .Z(n687) );
  NAND U792 ( .A(B[155]), .B(n691), .Z(n690) );
  NANDN U793 ( .A(A[155]), .B(n692), .Z(n691) );
  NANDN U794 ( .A(n692), .B(A[155]), .Z(n689) );
  XOR U795 ( .A(n692), .B(n693), .Z(SUM[155]) );
  XNOR U796 ( .A(B[155]), .B(A[155]), .Z(n693) );
  AND U797 ( .A(n694), .B(n695), .Z(n692) );
  NAND U798 ( .A(B[154]), .B(n696), .Z(n695) );
  NANDN U799 ( .A(A[154]), .B(n697), .Z(n696) );
  NANDN U800 ( .A(n697), .B(A[154]), .Z(n694) );
  XOR U801 ( .A(n697), .B(n698), .Z(SUM[154]) );
  XNOR U802 ( .A(B[154]), .B(A[154]), .Z(n698) );
  AND U803 ( .A(n699), .B(n700), .Z(n697) );
  NAND U804 ( .A(B[153]), .B(n701), .Z(n700) );
  NANDN U805 ( .A(A[153]), .B(n702), .Z(n701) );
  NANDN U806 ( .A(n702), .B(A[153]), .Z(n699) );
  XOR U807 ( .A(n702), .B(n703), .Z(SUM[153]) );
  XNOR U808 ( .A(B[153]), .B(A[153]), .Z(n703) );
  AND U809 ( .A(n704), .B(n705), .Z(n702) );
  NAND U810 ( .A(B[152]), .B(n706), .Z(n705) );
  NANDN U811 ( .A(A[152]), .B(n707), .Z(n706) );
  NANDN U812 ( .A(n707), .B(A[152]), .Z(n704) );
  XOR U813 ( .A(n707), .B(n708), .Z(SUM[152]) );
  XNOR U814 ( .A(B[152]), .B(A[152]), .Z(n708) );
  AND U815 ( .A(n709), .B(n710), .Z(n707) );
  NAND U816 ( .A(B[151]), .B(n711), .Z(n710) );
  NANDN U817 ( .A(A[151]), .B(n712), .Z(n711) );
  NANDN U818 ( .A(n712), .B(A[151]), .Z(n709) );
  XOR U819 ( .A(n712), .B(n713), .Z(SUM[151]) );
  XNOR U820 ( .A(B[151]), .B(A[151]), .Z(n713) );
  AND U821 ( .A(n714), .B(n715), .Z(n712) );
  NAND U822 ( .A(B[150]), .B(n716), .Z(n715) );
  NANDN U823 ( .A(A[150]), .B(n717), .Z(n716) );
  NANDN U824 ( .A(n717), .B(A[150]), .Z(n714) );
  XOR U825 ( .A(n717), .B(n718), .Z(SUM[150]) );
  XNOR U826 ( .A(B[150]), .B(A[150]), .Z(n718) );
  AND U827 ( .A(n719), .B(n720), .Z(n717) );
  NAND U828 ( .A(B[149]), .B(n721), .Z(n720) );
  NANDN U829 ( .A(A[149]), .B(n722), .Z(n721) );
  NANDN U830 ( .A(n722), .B(A[149]), .Z(n719) );
  XOR U831 ( .A(n723), .B(n724), .Z(SUM[14]) );
  XNOR U832 ( .A(B[14]), .B(A[14]), .Z(n724) );
  XOR U833 ( .A(n722), .B(n725), .Z(SUM[149]) );
  XNOR U834 ( .A(B[149]), .B(A[149]), .Z(n725) );
  AND U835 ( .A(n726), .B(n727), .Z(n722) );
  NAND U836 ( .A(B[148]), .B(n728), .Z(n727) );
  NANDN U837 ( .A(A[148]), .B(n729), .Z(n728) );
  NANDN U838 ( .A(n729), .B(A[148]), .Z(n726) );
  XOR U839 ( .A(n729), .B(n730), .Z(SUM[148]) );
  XNOR U840 ( .A(B[148]), .B(A[148]), .Z(n730) );
  AND U841 ( .A(n731), .B(n732), .Z(n729) );
  NAND U842 ( .A(B[147]), .B(n733), .Z(n732) );
  NANDN U843 ( .A(A[147]), .B(n734), .Z(n733) );
  NANDN U844 ( .A(n734), .B(A[147]), .Z(n731) );
  XOR U845 ( .A(n734), .B(n735), .Z(SUM[147]) );
  XNOR U846 ( .A(B[147]), .B(A[147]), .Z(n735) );
  AND U847 ( .A(n736), .B(n737), .Z(n734) );
  NAND U848 ( .A(B[146]), .B(n738), .Z(n737) );
  NANDN U849 ( .A(A[146]), .B(n739), .Z(n738) );
  NANDN U850 ( .A(n739), .B(A[146]), .Z(n736) );
  XOR U851 ( .A(n739), .B(n740), .Z(SUM[146]) );
  XNOR U852 ( .A(B[146]), .B(A[146]), .Z(n740) );
  AND U853 ( .A(n741), .B(n742), .Z(n739) );
  NAND U854 ( .A(B[145]), .B(n743), .Z(n742) );
  NANDN U855 ( .A(A[145]), .B(n744), .Z(n743) );
  NANDN U856 ( .A(n744), .B(A[145]), .Z(n741) );
  XOR U857 ( .A(n744), .B(n745), .Z(SUM[145]) );
  XNOR U858 ( .A(B[145]), .B(A[145]), .Z(n745) );
  AND U859 ( .A(n746), .B(n747), .Z(n744) );
  NAND U860 ( .A(B[144]), .B(n748), .Z(n747) );
  NANDN U861 ( .A(A[144]), .B(n749), .Z(n748) );
  NANDN U862 ( .A(n749), .B(A[144]), .Z(n746) );
  XOR U863 ( .A(n749), .B(n750), .Z(SUM[144]) );
  XNOR U864 ( .A(B[144]), .B(A[144]), .Z(n750) );
  AND U865 ( .A(n751), .B(n752), .Z(n749) );
  NAND U866 ( .A(B[143]), .B(n753), .Z(n752) );
  NANDN U867 ( .A(A[143]), .B(n754), .Z(n753) );
  NANDN U868 ( .A(n754), .B(A[143]), .Z(n751) );
  XOR U869 ( .A(n754), .B(n755), .Z(SUM[143]) );
  XNOR U870 ( .A(B[143]), .B(A[143]), .Z(n755) );
  AND U871 ( .A(n756), .B(n757), .Z(n754) );
  NAND U872 ( .A(B[142]), .B(n758), .Z(n757) );
  NANDN U873 ( .A(A[142]), .B(n759), .Z(n758) );
  NANDN U874 ( .A(n759), .B(A[142]), .Z(n756) );
  XOR U875 ( .A(n759), .B(n760), .Z(SUM[142]) );
  XNOR U876 ( .A(B[142]), .B(A[142]), .Z(n760) );
  AND U877 ( .A(n761), .B(n762), .Z(n759) );
  NAND U878 ( .A(B[141]), .B(n763), .Z(n762) );
  NANDN U879 ( .A(A[141]), .B(n764), .Z(n763) );
  NANDN U880 ( .A(n764), .B(A[141]), .Z(n761) );
  XOR U881 ( .A(n764), .B(n765), .Z(SUM[141]) );
  XNOR U882 ( .A(B[141]), .B(A[141]), .Z(n765) );
  AND U883 ( .A(n766), .B(n767), .Z(n764) );
  NAND U884 ( .A(B[140]), .B(n768), .Z(n767) );
  NANDN U885 ( .A(A[140]), .B(n769), .Z(n768) );
  NANDN U886 ( .A(n769), .B(A[140]), .Z(n766) );
  XOR U887 ( .A(n769), .B(n770), .Z(SUM[140]) );
  XNOR U888 ( .A(B[140]), .B(A[140]), .Z(n770) );
  AND U889 ( .A(n771), .B(n772), .Z(n769) );
  NAND U890 ( .A(B[139]), .B(n773), .Z(n772) );
  NANDN U891 ( .A(A[139]), .B(n774), .Z(n773) );
  NANDN U892 ( .A(n774), .B(A[139]), .Z(n771) );
  XOR U893 ( .A(n775), .B(n776), .Z(SUM[13]) );
  XNOR U894 ( .A(B[13]), .B(A[13]), .Z(n776) );
  XOR U895 ( .A(n774), .B(n777), .Z(SUM[139]) );
  XNOR U896 ( .A(B[139]), .B(A[139]), .Z(n777) );
  AND U897 ( .A(n778), .B(n779), .Z(n774) );
  NAND U898 ( .A(B[138]), .B(n780), .Z(n779) );
  NANDN U899 ( .A(A[138]), .B(n781), .Z(n780) );
  NANDN U900 ( .A(n781), .B(A[138]), .Z(n778) );
  XOR U901 ( .A(n781), .B(n782), .Z(SUM[138]) );
  XNOR U902 ( .A(B[138]), .B(A[138]), .Z(n782) );
  AND U903 ( .A(n783), .B(n784), .Z(n781) );
  NAND U904 ( .A(B[137]), .B(n785), .Z(n784) );
  NANDN U905 ( .A(A[137]), .B(n786), .Z(n785) );
  NANDN U906 ( .A(n786), .B(A[137]), .Z(n783) );
  XOR U907 ( .A(n786), .B(n787), .Z(SUM[137]) );
  XNOR U908 ( .A(B[137]), .B(A[137]), .Z(n787) );
  AND U909 ( .A(n788), .B(n789), .Z(n786) );
  NAND U910 ( .A(B[136]), .B(n790), .Z(n789) );
  NANDN U911 ( .A(A[136]), .B(n791), .Z(n790) );
  NANDN U912 ( .A(n791), .B(A[136]), .Z(n788) );
  XOR U913 ( .A(n791), .B(n792), .Z(SUM[136]) );
  XNOR U914 ( .A(B[136]), .B(A[136]), .Z(n792) );
  AND U915 ( .A(n793), .B(n794), .Z(n791) );
  NAND U916 ( .A(B[135]), .B(n795), .Z(n794) );
  NANDN U917 ( .A(A[135]), .B(n796), .Z(n795) );
  NANDN U918 ( .A(n796), .B(A[135]), .Z(n793) );
  XOR U919 ( .A(n796), .B(n797), .Z(SUM[135]) );
  XNOR U920 ( .A(B[135]), .B(A[135]), .Z(n797) );
  AND U921 ( .A(n798), .B(n799), .Z(n796) );
  NAND U922 ( .A(B[134]), .B(n800), .Z(n799) );
  NANDN U923 ( .A(A[134]), .B(n801), .Z(n800) );
  NANDN U924 ( .A(n801), .B(A[134]), .Z(n798) );
  XOR U925 ( .A(n801), .B(n802), .Z(SUM[134]) );
  XNOR U926 ( .A(B[134]), .B(A[134]), .Z(n802) );
  AND U927 ( .A(n803), .B(n804), .Z(n801) );
  NAND U928 ( .A(B[133]), .B(n805), .Z(n804) );
  NANDN U929 ( .A(A[133]), .B(n806), .Z(n805) );
  NANDN U930 ( .A(n806), .B(A[133]), .Z(n803) );
  XOR U931 ( .A(n806), .B(n807), .Z(SUM[133]) );
  XNOR U932 ( .A(B[133]), .B(A[133]), .Z(n807) );
  AND U933 ( .A(n808), .B(n809), .Z(n806) );
  NAND U934 ( .A(B[132]), .B(n810), .Z(n809) );
  NANDN U935 ( .A(A[132]), .B(n811), .Z(n810) );
  NANDN U936 ( .A(n811), .B(A[132]), .Z(n808) );
  XOR U937 ( .A(n811), .B(n812), .Z(SUM[132]) );
  XNOR U938 ( .A(B[132]), .B(A[132]), .Z(n812) );
  AND U939 ( .A(n813), .B(n814), .Z(n811) );
  NAND U940 ( .A(B[131]), .B(n815), .Z(n814) );
  NANDN U941 ( .A(A[131]), .B(n816), .Z(n815) );
  NANDN U942 ( .A(n816), .B(A[131]), .Z(n813) );
  XOR U943 ( .A(n816), .B(n817), .Z(SUM[131]) );
  XNOR U944 ( .A(B[131]), .B(A[131]), .Z(n817) );
  AND U945 ( .A(n818), .B(n819), .Z(n816) );
  NAND U946 ( .A(B[130]), .B(n820), .Z(n819) );
  NANDN U947 ( .A(A[130]), .B(n821), .Z(n820) );
  NANDN U948 ( .A(n821), .B(A[130]), .Z(n818) );
  XOR U949 ( .A(n821), .B(n822), .Z(SUM[130]) );
  XNOR U950 ( .A(B[130]), .B(A[130]), .Z(n822) );
  AND U951 ( .A(n823), .B(n824), .Z(n821) );
  NAND U952 ( .A(B[129]), .B(n825), .Z(n824) );
  NANDN U953 ( .A(A[129]), .B(n826), .Z(n825) );
  NANDN U954 ( .A(n826), .B(A[129]), .Z(n823) );
  XOR U955 ( .A(n827), .B(n828), .Z(SUM[12]) );
  XNOR U956 ( .A(B[12]), .B(A[12]), .Z(n828) );
  XOR U957 ( .A(n826), .B(n829), .Z(SUM[129]) );
  XNOR U958 ( .A(B[129]), .B(A[129]), .Z(n829) );
  AND U959 ( .A(n830), .B(n831), .Z(n826) );
  NAND U960 ( .A(B[128]), .B(n832), .Z(n831) );
  NANDN U961 ( .A(A[128]), .B(n833), .Z(n832) );
  NANDN U962 ( .A(n833), .B(A[128]), .Z(n830) );
  XOR U963 ( .A(n833), .B(n834), .Z(SUM[128]) );
  XNOR U964 ( .A(B[128]), .B(A[128]), .Z(n834) );
  AND U965 ( .A(n835), .B(n836), .Z(n833) );
  NAND U966 ( .A(B[127]), .B(n837), .Z(n836) );
  NANDN U967 ( .A(A[127]), .B(n838), .Z(n837) );
  NANDN U968 ( .A(n838), .B(A[127]), .Z(n835) );
  XOR U969 ( .A(n838), .B(n839), .Z(SUM[127]) );
  XNOR U970 ( .A(B[127]), .B(A[127]), .Z(n839) );
  AND U971 ( .A(n840), .B(n841), .Z(n838) );
  NAND U972 ( .A(B[126]), .B(n842), .Z(n841) );
  NANDN U973 ( .A(A[126]), .B(n843), .Z(n842) );
  NANDN U974 ( .A(n843), .B(A[126]), .Z(n840) );
  XOR U975 ( .A(n843), .B(n844), .Z(SUM[126]) );
  XNOR U976 ( .A(B[126]), .B(A[126]), .Z(n844) );
  AND U977 ( .A(n845), .B(n846), .Z(n843) );
  NAND U978 ( .A(B[125]), .B(n847), .Z(n846) );
  NANDN U979 ( .A(A[125]), .B(n848), .Z(n847) );
  NANDN U980 ( .A(n848), .B(A[125]), .Z(n845) );
  XOR U981 ( .A(n848), .B(n849), .Z(SUM[125]) );
  XNOR U982 ( .A(B[125]), .B(A[125]), .Z(n849) );
  AND U983 ( .A(n850), .B(n851), .Z(n848) );
  NAND U984 ( .A(B[124]), .B(n852), .Z(n851) );
  NANDN U985 ( .A(A[124]), .B(n853), .Z(n852) );
  NANDN U986 ( .A(n853), .B(A[124]), .Z(n850) );
  XOR U987 ( .A(n853), .B(n854), .Z(SUM[124]) );
  XNOR U988 ( .A(B[124]), .B(A[124]), .Z(n854) );
  AND U989 ( .A(n855), .B(n856), .Z(n853) );
  NAND U990 ( .A(B[123]), .B(n857), .Z(n856) );
  NANDN U991 ( .A(A[123]), .B(n858), .Z(n857) );
  NANDN U992 ( .A(n858), .B(A[123]), .Z(n855) );
  XOR U993 ( .A(n858), .B(n859), .Z(SUM[123]) );
  XNOR U994 ( .A(B[123]), .B(A[123]), .Z(n859) );
  AND U995 ( .A(n860), .B(n861), .Z(n858) );
  NAND U996 ( .A(B[122]), .B(n862), .Z(n861) );
  NANDN U997 ( .A(A[122]), .B(n863), .Z(n862) );
  NANDN U998 ( .A(n863), .B(A[122]), .Z(n860) );
  XOR U999 ( .A(n863), .B(n864), .Z(SUM[122]) );
  XNOR U1000 ( .A(B[122]), .B(A[122]), .Z(n864) );
  AND U1001 ( .A(n865), .B(n866), .Z(n863) );
  NAND U1002 ( .A(B[121]), .B(n867), .Z(n866) );
  NANDN U1003 ( .A(A[121]), .B(n868), .Z(n867) );
  NANDN U1004 ( .A(n868), .B(A[121]), .Z(n865) );
  XOR U1005 ( .A(n868), .B(n869), .Z(SUM[121]) );
  XNOR U1006 ( .A(B[121]), .B(A[121]), .Z(n869) );
  AND U1007 ( .A(n870), .B(n871), .Z(n868) );
  NAND U1008 ( .A(B[120]), .B(n872), .Z(n871) );
  NANDN U1009 ( .A(A[120]), .B(n873), .Z(n872) );
  NANDN U1010 ( .A(n873), .B(A[120]), .Z(n870) );
  XOR U1011 ( .A(n873), .B(n874), .Z(SUM[120]) );
  XNOR U1012 ( .A(B[120]), .B(A[120]), .Z(n874) );
  AND U1013 ( .A(n875), .B(n876), .Z(n873) );
  NAND U1014 ( .A(B[119]), .B(n877), .Z(n876) );
  NANDN U1015 ( .A(A[119]), .B(n878), .Z(n877) );
  NANDN U1016 ( .A(n878), .B(A[119]), .Z(n875) );
  XOR U1017 ( .A(n879), .B(n880), .Z(SUM[11]) );
  XNOR U1018 ( .A(B[11]), .B(A[11]), .Z(n880) );
  XOR U1019 ( .A(n878), .B(n881), .Z(SUM[119]) );
  XNOR U1020 ( .A(B[119]), .B(A[119]), .Z(n881) );
  AND U1021 ( .A(n882), .B(n883), .Z(n878) );
  NAND U1022 ( .A(B[118]), .B(n884), .Z(n883) );
  NANDN U1023 ( .A(A[118]), .B(n885), .Z(n884) );
  NANDN U1024 ( .A(n885), .B(A[118]), .Z(n882) );
  XOR U1025 ( .A(n885), .B(n886), .Z(SUM[118]) );
  XNOR U1026 ( .A(B[118]), .B(A[118]), .Z(n886) );
  AND U1027 ( .A(n887), .B(n888), .Z(n885) );
  NAND U1028 ( .A(B[117]), .B(n889), .Z(n888) );
  NANDN U1029 ( .A(A[117]), .B(n890), .Z(n889) );
  NANDN U1030 ( .A(n890), .B(A[117]), .Z(n887) );
  XOR U1031 ( .A(n890), .B(n891), .Z(SUM[117]) );
  XNOR U1032 ( .A(B[117]), .B(A[117]), .Z(n891) );
  AND U1033 ( .A(n892), .B(n893), .Z(n890) );
  NAND U1034 ( .A(B[116]), .B(n894), .Z(n893) );
  NANDN U1035 ( .A(A[116]), .B(n895), .Z(n894) );
  NANDN U1036 ( .A(n895), .B(A[116]), .Z(n892) );
  XOR U1037 ( .A(n895), .B(n896), .Z(SUM[116]) );
  XNOR U1038 ( .A(B[116]), .B(A[116]), .Z(n896) );
  AND U1039 ( .A(n897), .B(n898), .Z(n895) );
  NAND U1040 ( .A(B[115]), .B(n899), .Z(n898) );
  NANDN U1041 ( .A(A[115]), .B(n900), .Z(n899) );
  NANDN U1042 ( .A(n900), .B(A[115]), .Z(n897) );
  XOR U1043 ( .A(n900), .B(n901), .Z(SUM[115]) );
  XNOR U1044 ( .A(B[115]), .B(A[115]), .Z(n901) );
  AND U1045 ( .A(n902), .B(n903), .Z(n900) );
  NAND U1046 ( .A(B[114]), .B(n904), .Z(n903) );
  NANDN U1047 ( .A(A[114]), .B(n905), .Z(n904) );
  NANDN U1048 ( .A(n905), .B(A[114]), .Z(n902) );
  XOR U1049 ( .A(n905), .B(n906), .Z(SUM[114]) );
  XNOR U1050 ( .A(B[114]), .B(A[114]), .Z(n906) );
  AND U1051 ( .A(n907), .B(n908), .Z(n905) );
  NAND U1052 ( .A(B[113]), .B(n909), .Z(n908) );
  NANDN U1053 ( .A(A[113]), .B(n910), .Z(n909) );
  NANDN U1054 ( .A(n910), .B(A[113]), .Z(n907) );
  XOR U1055 ( .A(n910), .B(n911), .Z(SUM[113]) );
  XNOR U1056 ( .A(B[113]), .B(A[113]), .Z(n911) );
  AND U1057 ( .A(n912), .B(n913), .Z(n910) );
  NAND U1058 ( .A(B[112]), .B(n914), .Z(n913) );
  NANDN U1059 ( .A(A[112]), .B(n915), .Z(n914) );
  NANDN U1060 ( .A(n915), .B(A[112]), .Z(n912) );
  XOR U1061 ( .A(n915), .B(n916), .Z(SUM[112]) );
  XNOR U1062 ( .A(B[112]), .B(A[112]), .Z(n916) );
  AND U1063 ( .A(n917), .B(n918), .Z(n915) );
  NAND U1064 ( .A(B[111]), .B(n919), .Z(n918) );
  NANDN U1065 ( .A(A[111]), .B(n920), .Z(n919) );
  NANDN U1066 ( .A(n920), .B(A[111]), .Z(n917) );
  XOR U1067 ( .A(n920), .B(n921), .Z(SUM[111]) );
  XNOR U1068 ( .A(B[111]), .B(A[111]), .Z(n921) );
  AND U1069 ( .A(n922), .B(n923), .Z(n920) );
  NAND U1070 ( .A(B[110]), .B(n924), .Z(n923) );
  NANDN U1071 ( .A(A[110]), .B(n925), .Z(n924) );
  NANDN U1072 ( .A(n925), .B(A[110]), .Z(n922) );
  XOR U1073 ( .A(n925), .B(n926), .Z(SUM[110]) );
  XNOR U1074 ( .A(B[110]), .B(A[110]), .Z(n926) );
  AND U1075 ( .A(n927), .B(n928), .Z(n925) );
  NAND U1076 ( .A(B[109]), .B(n929), .Z(n928) );
  NANDN U1077 ( .A(A[109]), .B(n930), .Z(n929) );
  NANDN U1078 ( .A(n930), .B(A[109]), .Z(n927) );
  XOR U1079 ( .A(n931), .B(n932), .Z(SUM[10]) );
  XNOR U1080 ( .A(B[10]), .B(A[10]), .Z(n932) );
  XOR U1081 ( .A(n930), .B(n933), .Z(SUM[109]) );
  XNOR U1082 ( .A(B[109]), .B(A[109]), .Z(n933) );
  AND U1083 ( .A(n934), .B(n935), .Z(n930) );
  NAND U1084 ( .A(B[108]), .B(n936), .Z(n935) );
  NANDN U1085 ( .A(A[108]), .B(n937), .Z(n936) );
  NANDN U1086 ( .A(n937), .B(A[108]), .Z(n934) );
  XOR U1087 ( .A(n937), .B(n938), .Z(SUM[108]) );
  XNOR U1088 ( .A(B[108]), .B(A[108]), .Z(n938) );
  AND U1089 ( .A(n939), .B(n940), .Z(n937) );
  NAND U1090 ( .A(B[107]), .B(n941), .Z(n940) );
  NANDN U1091 ( .A(A[107]), .B(n942), .Z(n941) );
  NANDN U1092 ( .A(n942), .B(A[107]), .Z(n939) );
  XOR U1093 ( .A(n942), .B(n943), .Z(SUM[107]) );
  XNOR U1094 ( .A(B[107]), .B(A[107]), .Z(n943) );
  AND U1095 ( .A(n944), .B(n945), .Z(n942) );
  NAND U1096 ( .A(B[106]), .B(n946), .Z(n945) );
  NANDN U1097 ( .A(A[106]), .B(n947), .Z(n946) );
  NANDN U1098 ( .A(n947), .B(A[106]), .Z(n944) );
  XOR U1099 ( .A(n947), .B(n948), .Z(SUM[106]) );
  XNOR U1100 ( .A(B[106]), .B(A[106]), .Z(n948) );
  AND U1101 ( .A(n949), .B(n950), .Z(n947) );
  NAND U1102 ( .A(B[105]), .B(n951), .Z(n950) );
  NANDN U1103 ( .A(A[105]), .B(n952), .Z(n951) );
  NANDN U1104 ( .A(n952), .B(A[105]), .Z(n949) );
  XOR U1105 ( .A(n952), .B(n953), .Z(SUM[105]) );
  XNOR U1106 ( .A(B[105]), .B(A[105]), .Z(n953) );
  AND U1107 ( .A(n954), .B(n955), .Z(n952) );
  NAND U1108 ( .A(B[104]), .B(n956), .Z(n955) );
  NANDN U1109 ( .A(A[104]), .B(n957), .Z(n956) );
  NANDN U1110 ( .A(n957), .B(A[104]), .Z(n954) );
  XOR U1111 ( .A(n957), .B(n958), .Z(SUM[104]) );
  XNOR U1112 ( .A(B[104]), .B(A[104]), .Z(n958) );
  AND U1113 ( .A(n959), .B(n960), .Z(n957) );
  NAND U1114 ( .A(B[103]), .B(n961), .Z(n960) );
  NANDN U1115 ( .A(A[103]), .B(n962), .Z(n961) );
  NANDN U1116 ( .A(n962), .B(A[103]), .Z(n959) );
  XOR U1117 ( .A(n962), .B(n963), .Z(SUM[103]) );
  XNOR U1118 ( .A(B[103]), .B(A[103]), .Z(n963) );
  AND U1119 ( .A(n964), .B(n965), .Z(n962) );
  NAND U1120 ( .A(B[102]), .B(n966), .Z(n965) );
  NANDN U1121 ( .A(A[102]), .B(n967), .Z(n966) );
  NANDN U1122 ( .A(n967), .B(A[102]), .Z(n964) );
  XOR U1123 ( .A(n967), .B(n968), .Z(SUM[102]) );
  XNOR U1124 ( .A(B[102]), .B(A[102]), .Z(n968) );
  AND U1125 ( .A(n969), .B(n970), .Z(n967) );
  NAND U1126 ( .A(B[101]), .B(n971), .Z(n970) );
  NANDN U1127 ( .A(A[101]), .B(n972), .Z(n971) );
  NANDN U1128 ( .A(n972), .B(A[101]), .Z(n969) );
  XOR U1129 ( .A(n972), .B(n973), .Z(SUM[101]) );
  XNOR U1130 ( .A(B[101]), .B(A[101]), .Z(n973) );
  AND U1131 ( .A(n974), .B(n975), .Z(n972) );
  NAND U1132 ( .A(B[100]), .B(n976), .Z(n975) );
  NANDN U1133 ( .A(A[100]), .B(n977), .Z(n976) );
  NANDN U1134 ( .A(n977), .B(A[100]), .Z(n974) );
  XOR U1135 ( .A(n977), .B(n978), .Z(SUM[100]) );
  XNOR U1136 ( .A(B[100]), .B(A[100]), .Z(n978) );
  AND U1137 ( .A(n979), .B(n980), .Z(n977) );
  NAND U1138 ( .A(B[99]), .B(n981), .Z(n980) );
  OR U1139 ( .A(n3), .B(A[99]), .Z(n981) );
  NAND U1140 ( .A(A[99]), .B(n3), .Z(n979) );
  NAND U1141 ( .A(n982), .B(n983), .Z(n3) );
  NAND U1142 ( .A(B[98]), .B(n984), .Z(n983) );
  NANDN U1143 ( .A(A[98]), .B(n5), .Z(n984) );
  NANDN U1144 ( .A(n5), .B(A[98]), .Z(n982) );
  AND U1145 ( .A(n985), .B(n986), .Z(n5) );
  NAND U1146 ( .A(B[97]), .B(n987), .Z(n986) );
  NANDN U1147 ( .A(A[97]), .B(n7), .Z(n987) );
  NANDN U1148 ( .A(n7), .B(A[97]), .Z(n985) );
  AND U1149 ( .A(n988), .B(n989), .Z(n7) );
  NAND U1150 ( .A(B[96]), .B(n990), .Z(n989) );
  NANDN U1151 ( .A(A[96]), .B(n9), .Z(n990) );
  NANDN U1152 ( .A(n9), .B(A[96]), .Z(n988) );
  AND U1153 ( .A(n991), .B(n992), .Z(n9) );
  NAND U1154 ( .A(B[95]), .B(n993), .Z(n992) );
  NANDN U1155 ( .A(A[95]), .B(n11), .Z(n993) );
  NANDN U1156 ( .A(n11), .B(A[95]), .Z(n991) );
  AND U1157 ( .A(n994), .B(n995), .Z(n11) );
  NAND U1158 ( .A(B[94]), .B(n996), .Z(n995) );
  NANDN U1159 ( .A(A[94]), .B(n13), .Z(n996) );
  NANDN U1160 ( .A(n13), .B(A[94]), .Z(n994) );
  AND U1161 ( .A(n997), .B(n998), .Z(n13) );
  NAND U1162 ( .A(B[93]), .B(n999), .Z(n998) );
  NANDN U1163 ( .A(A[93]), .B(n15), .Z(n999) );
  NANDN U1164 ( .A(n15), .B(A[93]), .Z(n997) );
  AND U1165 ( .A(n1000), .B(n1001), .Z(n15) );
  NAND U1166 ( .A(B[92]), .B(n1002), .Z(n1001) );
  NANDN U1167 ( .A(A[92]), .B(n17), .Z(n1002) );
  NANDN U1168 ( .A(n17), .B(A[92]), .Z(n1000) );
  AND U1169 ( .A(n1003), .B(n1004), .Z(n17) );
  NAND U1170 ( .A(B[91]), .B(n1005), .Z(n1004) );
  NANDN U1171 ( .A(A[91]), .B(n19), .Z(n1005) );
  NANDN U1172 ( .A(n19), .B(A[91]), .Z(n1003) );
  AND U1173 ( .A(n1006), .B(n1007), .Z(n19) );
  NAND U1174 ( .A(B[90]), .B(n1008), .Z(n1007) );
  NANDN U1175 ( .A(A[90]), .B(n21), .Z(n1008) );
  NANDN U1176 ( .A(n21), .B(A[90]), .Z(n1006) );
  AND U1177 ( .A(n1009), .B(n1010), .Z(n21) );
  NAND U1178 ( .A(B[89]), .B(n1011), .Z(n1010) );
  NANDN U1179 ( .A(A[89]), .B(n25), .Z(n1011) );
  NANDN U1180 ( .A(n25), .B(A[89]), .Z(n1009) );
  AND U1181 ( .A(n1012), .B(n1013), .Z(n25) );
  NAND U1182 ( .A(B[88]), .B(n1014), .Z(n1013) );
  NANDN U1183 ( .A(A[88]), .B(n27), .Z(n1014) );
  NANDN U1184 ( .A(n27), .B(A[88]), .Z(n1012) );
  AND U1185 ( .A(n1015), .B(n1016), .Z(n27) );
  NAND U1186 ( .A(B[87]), .B(n1017), .Z(n1016) );
  NANDN U1187 ( .A(A[87]), .B(n29), .Z(n1017) );
  NANDN U1188 ( .A(n29), .B(A[87]), .Z(n1015) );
  AND U1189 ( .A(n1018), .B(n1019), .Z(n29) );
  NAND U1190 ( .A(B[86]), .B(n1020), .Z(n1019) );
  NANDN U1191 ( .A(A[86]), .B(n31), .Z(n1020) );
  NANDN U1192 ( .A(n31), .B(A[86]), .Z(n1018) );
  AND U1193 ( .A(n1021), .B(n1022), .Z(n31) );
  NAND U1194 ( .A(B[85]), .B(n1023), .Z(n1022) );
  NANDN U1195 ( .A(A[85]), .B(n33), .Z(n1023) );
  NANDN U1196 ( .A(n33), .B(A[85]), .Z(n1021) );
  AND U1197 ( .A(n1024), .B(n1025), .Z(n33) );
  NAND U1198 ( .A(B[84]), .B(n1026), .Z(n1025) );
  NANDN U1199 ( .A(A[84]), .B(n35), .Z(n1026) );
  NANDN U1200 ( .A(n35), .B(A[84]), .Z(n1024) );
  AND U1201 ( .A(n1027), .B(n1028), .Z(n35) );
  NAND U1202 ( .A(B[83]), .B(n1029), .Z(n1028) );
  NANDN U1203 ( .A(A[83]), .B(n37), .Z(n1029) );
  NANDN U1204 ( .A(n37), .B(A[83]), .Z(n1027) );
  AND U1205 ( .A(n1030), .B(n1031), .Z(n37) );
  NAND U1206 ( .A(B[82]), .B(n1032), .Z(n1031) );
  NANDN U1207 ( .A(A[82]), .B(n39), .Z(n1032) );
  NANDN U1208 ( .A(n39), .B(A[82]), .Z(n1030) );
  AND U1209 ( .A(n1033), .B(n1034), .Z(n39) );
  NAND U1210 ( .A(B[81]), .B(n1035), .Z(n1034) );
  NANDN U1211 ( .A(A[81]), .B(n41), .Z(n1035) );
  NANDN U1212 ( .A(n41), .B(A[81]), .Z(n1033) );
  AND U1213 ( .A(n1036), .B(n1037), .Z(n41) );
  NAND U1214 ( .A(B[80]), .B(n1038), .Z(n1037) );
  NANDN U1215 ( .A(A[80]), .B(n43), .Z(n1038) );
  NANDN U1216 ( .A(n43), .B(A[80]), .Z(n1036) );
  AND U1217 ( .A(n1039), .B(n1040), .Z(n43) );
  NAND U1218 ( .A(B[79]), .B(n1041), .Z(n1040) );
  NANDN U1219 ( .A(A[79]), .B(n47), .Z(n1041) );
  NANDN U1220 ( .A(n47), .B(A[79]), .Z(n1039) );
  AND U1221 ( .A(n1042), .B(n1043), .Z(n47) );
  NAND U1222 ( .A(B[78]), .B(n1044), .Z(n1043) );
  NANDN U1223 ( .A(A[78]), .B(n49), .Z(n1044) );
  NANDN U1224 ( .A(n49), .B(A[78]), .Z(n1042) );
  AND U1225 ( .A(n1045), .B(n1046), .Z(n49) );
  NAND U1226 ( .A(B[77]), .B(n1047), .Z(n1046) );
  NANDN U1227 ( .A(A[77]), .B(n51), .Z(n1047) );
  NANDN U1228 ( .A(n51), .B(A[77]), .Z(n1045) );
  AND U1229 ( .A(n1048), .B(n1049), .Z(n51) );
  NAND U1230 ( .A(B[76]), .B(n1050), .Z(n1049) );
  NANDN U1231 ( .A(A[76]), .B(n53), .Z(n1050) );
  NANDN U1232 ( .A(n53), .B(A[76]), .Z(n1048) );
  AND U1233 ( .A(n1051), .B(n1052), .Z(n53) );
  NAND U1234 ( .A(B[75]), .B(n1053), .Z(n1052) );
  NANDN U1235 ( .A(A[75]), .B(n55), .Z(n1053) );
  NANDN U1236 ( .A(n55), .B(A[75]), .Z(n1051) );
  AND U1237 ( .A(n1054), .B(n1055), .Z(n55) );
  NAND U1238 ( .A(B[74]), .B(n1056), .Z(n1055) );
  NANDN U1239 ( .A(A[74]), .B(n57), .Z(n1056) );
  NANDN U1240 ( .A(n57), .B(A[74]), .Z(n1054) );
  AND U1241 ( .A(n1057), .B(n1058), .Z(n57) );
  NAND U1242 ( .A(B[73]), .B(n1059), .Z(n1058) );
  NANDN U1243 ( .A(A[73]), .B(n59), .Z(n1059) );
  NANDN U1244 ( .A(n59), .B(A[73]), .Z(n1057) );
  AND U1245 ( .A(n1060), .B(n1061), .Z(n59) );
  NAND U1246 ( .A(B[72]), .B(n1062), .Z(n1061) );
  NANDN U1247 ( .A(A[72]), .B(n61), .Z(n1062) );
  NANDN U1248 ( .A(n61), .B(A[72]), .Z(n1060) );
  AND U1249 ( .A(n1063), .B(n1064), .Z(n61) );
  NAND U1250 ( .A(B[71]), .B(n1065), .Z(n1064) );
  NANDN U1251 ( .A(A[71]), .B(n63), .Z(n1065) );
  NANDN U1252 ( .A(n63), .B(A[71]), .Z(n1063) );
  AND U1253 ( .A(n1066), .B(n1067), .Z(n63) );
  NAND U1254 ( .A(B[70]), .B(n1068), .Z(n1067) );
  NANDN U1255 ( .A(A[70]), .B(n65), .Z(n1068) );
  NANDN U1256 ( .A(n65), .B(A[70]), .Z(n1066) );
  AND U1257 ( .A(n1069), .B(n1070), .Z(n65) );
  NAND U1258 ( .A(B[69]), .B(n1071), .Z(n1070) );
  NANDN U1259 ( .A(A[69]), .B(n69), .Z(n1071) );
  NANDN U1260 ( .A(n69), .B(A[69]), .Z(n1069) );
  AND U1261 ( .A(n1072), .B(n1073), .Z(n69) );
  NAND U1262 ( .A(B[68]), .B(n1074), .Z(n1073) );
  NANDN U1263 ( .A(A[68]), .B(n71), .Z(n1074) );
  NANDN U1264 ( .A(n71), .B(A[68]), .Z(n1072) );
  AND U1265 ( .A(n1075), .B(n1076), .Z(n71) );
  NAND U1266 ( .A(B[67]), .B(n1077), .Z(n1076) );
  NANDN U1267 ( .A(A[67]), .B(n73), .Z(n1077) );
  NANDN U1268 ( .A(n73), .B(A[67]), .Z(n1075) );
  AND U1269 ( .A(n1078), .B(n1079), .Z(n73) );
  NAND U1270 ( .A(B[66]), .B(n1080), .Z(n1079) );
  NANDN U1271 ( .A(A[66]), .B(n75), .Z(n1080) );
  NANDN U1272 ( .A(n75), .B(A[66]), .Z(n1078) );
  AND U1273 ( .A(n1081), .B(n1082), .Z(n75) );
  NAND U1274 ( .A(B[65]), .B(n1083), .Z(n1082) );
  NANDN U1275 ( .A(A[65]), .B(n77), .Z(n1083) );
  NANDN U1276 ( .A(n77), .B(A[65]), .Z(n1081) );
  AND U1277 ( .A(n1084), .B(n1085), .Z(n77) );
  NAND U1278 ( .A(B[64]), .B(n1086), .Z(n1085) );
  NANDN U1279 ( .A(A[64]), .B(n79), .Z(n1086) );
  NANDN U1280 ( .A(n79), .B(A[64]), .Z(n1084) );
  AND U1281 ( .A(n1087), .B(n1088), .Z(n79) );
  NAND U1282 ( .A(B[63]), .B(n1089), .Z(n1088) );
  NANDN U1283 ( .A(A[63]), .B(n81), .Z(n1089) );
  NANDN U1284 ( .A(n81), .B(A[63]), .Z(n1087) );
  AND U1285 ( .A(n1090), .B(n1091), .Z(n81) );
  NAND U1286 ( .A(B[62]), .B(n1092), .Z(n1091) );
  NANDN U1287 ( .A(A[62]), .B(n83), .Z(n1092) );
  NANDN U1288 ( .A(n83), .B(A[62]), .Z(n1090) );
  AND U1289 ( .A(n1093), .B(n1094), .Z(n83) );
  NAND U1290 ( .A(B[61]), .B(n1095), .Z(n1094) );
  NANDN U1291 ( .A(A[61]), .B(n85), .Z(n1095) );
  NANDN U1292 ( .A(n85), .B(A[61]), .Z(n1093) );
  AND U1293 ( .A(n1096), .B(n1097), .Z(n85) );
  NAND U1294 ( .A(B[60]), .B(n1098), .Z(n1097) );
  NANDN U1295 ( .A(A[60]), .B(n87), .Z(n1098) );
  NANDN U1296 ( .A(n87), .B(A[60]), .Z(n1096) );
  AND U1297 ( .A(n1099), .B(n1100), .Z(n87) );
  NAND U1298 ( .A(B[59]), .B(n1101), .Z(n1100) );
  NANDN U1299 ( .A(A[59]), .B(n91), .Z(n1101) );
  NANDN U1300 ( .A(n91), .B(A[59]), .Z(n1099) );
  AND U1301 ( .A(n1102), .B(n1103), .Z(n91) );
  NAND U1302 ( .A(B[58]), .B(n1104), .Z(n1103) );
  NANDN U1303 ( .A(A[58]), .B(n93), .Z(n1104) );
  NANDN U1304 ( .A(n93), .B(A[58]), .Z(n1102) );
  AND U1305 ( .A(n1105), .B(n1106), .Z(n93) );
  NAND U1306 ( .A(B[57]), .B(n1107), .Z(n1106) );
  NANDN U1307 ( .A(A[57]), .B(n95), .Z(n1107) );
  NANDN U1308 ( .A(n95), .B(A[57]), .Z(n1105) );
  AND U1309 ( .A(n1108), .B(n1109), .Z(n95) );
  NAND U1310 ( .A(B[56]), .B(n1110), .Z(n1109) );
  NANDN U1311 ( .A(A[56]), .B(n97), .Z(n1110) );
  NANDN U1312 ( .A(n97), .B(A[56]), .Z(n1108) );
  AND U1313 ( .A(n1111), .B(n1112), .Z(n97) );
  NAND U1314 ( .A(B[55]), .B(n1113), .Z(n1112) );
  NANDN U1315 ( .A(A[55]), .B(n99), .Z(n1113) );
  NANDN U1316 ( .A(n99), .B(A[55]), .Z(n1111) );
  AND U1317 ( .A(n1114), .B(n1115), .Z(n99) );
  NAND U1318 ( .A(B[54]), .B(n1116), .Z(n1115) );
  NANDN U1319 ( .A(A[54]), .B(n101), .Z(n1116) );
  NANDN U1320 ( .A(n101), .B(A[54]), .Z(n1114) );
  AND U1321 ( .A(n1117), .B(n1118), .Z(n101) );
  NAND U1322 ( .A(B[53]), .B(n1119), .Z(n1118) );
  NANDN U1323 ( .A(A[53]), .B(n103), .Z(n1119) );
  NANDN U1324 ( .A(n103), .B(A[53]), .Z(n1117) );
  AND U1325 ( .A(n1120), .B(n1121), .Z(n103) );
  NAND U1326 ( .A(B[52]), .B(n1122), .Z(n1121) );
  NANDN U1327 ( .A(A[52]), .B(n105), .Z(n1122) );
  NANDN U1328 ( .A(n105), .B(A[52]), .Z(n1120) );
  AND U1329 ( .A(n1123), .B(n1124), .Z(n105) );
  NAND U1330 ( .A(B[51]), .B(n1125), .Z(n1124) );
  NANDN U1331 ( .A(A[51]), .B(n107), .Z(n1125) );
  NANDN U1332 ( .A(n107), .B(A[51]), .Z(n1123) );
  AND U1333 ( .A(n1126), .B(n1127), .Z(n107) );
  NAND U1334 ( .A(B[50]), .B(n1128), .Z(n1127) );
  NANDN U1335 ( .A(A[50]), .B(n109), .Z(n1128) );
  NANDN U1336 ( .A(n109), .B(A[50]), .Z(n1126) );
  AND U1337 ( .A(n1129), .B(n1130), .Z(n109) );
  NAND U1338 ( .A(B[49]), .B(n1131), .Z(n1130) );
  NANDN U1339 ( .A(A[49]), .B(n113), .Z(n1131) );
  NANDN U1340 ( .A(n113), .B(A[49]), .Z(n1129) );
  AND U1341 ( .A(n1132), .B(n1133), .Z(n113) );
  NAND U1342 ( .A(B[48]), .B(n1134), .Z(n1133) );
  NANDN U1343 ( .A(A[48]), .B(n115), .Z(n1134) );
  NANDN U1344 ( .A(n115), .B(A[48]), .Z(n1132) );
  AND U1345 ( .A(n1135), .B(n1136), .Z(n115) );
  NAND U1346 ( .A(B[47]), .B(n1137), .Z(n1136) );
  NANDN U1347 ( .A(A[47]), .B(n117), .Z(n1137) );
  NANDN U1348 ( .A(n117), .B(A[47]), .Z(n1135) );
  AND U1349 ( .A(n1138), .B(n1139), .Z(n117) );
  NAND U1350 ( .A(B[46]), .B(n1140), .Z(n1139) );
  NANDN U1351 ( .A(A[46]), .B(n119), .Z(n1140) );
  NANDN U1352 ( .A(n119), .B(A[46]), .Z(n1138) );
  AND U1353 ( .A(n1141), .B(n1142), .Z(n119) );
  NAND U1354 ( .A(B[45]), .B(n1143), .Z(n1142) );
  NANDN U1355 ( .A(A[45]), .B(n121), .Z(n1143) );
  NANDN U1356 ( .A(n121), .B(A[45]), .Z(n1141) );
  AND U1357 ( .A(n1144), .B(n1145), .Z(n121) );
  NAND U1358 ( .A(B[44]), .B(n1146), .Z(n1145) );
  NANDN U1359 ( .A(A[44]), .B(n123), .Z(n1146) );
  NANDN U1360 ( .A(n123), .B(A[44]), .Z(n1144) );
  AND U1361 ( .A(n1147), .B(n1148), .Z(n123) );
  NAND U1362 ( .A(B[43]), .B(n1149), .Z(n1148) );
  NANDN U1363 ( .A(A[43]), .B(n125), .Z(n1149) );
  NANDN U1364 ( .A(n125), .B(A[43]), .Z(n1147) );
  AND U1365 ( .A(n1150), .B(n1151), .Z(n125) );
  NAND U1366 ( .A(B[42]), .B(n1152), .Z(n1151) );
  NANDN U1367 ( .A(A[42]), .B(n127), .Z(n1152) );
  NANDN U1368 ( .A(n127), .B(A[42]), .Z(n1150) );
  AND U1369 ( .A(n1153), .B(n1154), .Z(n127) );
  NAND U1370 ( .A(B[41]), .B(n1155), .Z(n1154) );
  NANDN U1371 ( .A(A[41]), .B(n129), .Z(n1155) );
  NANDN U1372 ( .A(n129), .B(A[41]), .Z(n1153) );
  AND U1373 ( .A(n1156), .B(n1157), .Z(n129) );
  NAND U1374 ( .A(B[40]), .B(n1158), .Z(n1157) );
  NANDN U1375 ( .A(A[40]), .B(n131), .Z(n1158) );
  NANDN U1376 ( .A(n131), .B(A[40]), .Z(n1156) );
  AND U1377 ( .A(n1159), .B(n1160), .Z(n131) );
  NAND U1378 ( .A(B[39]), .B(n1161), .Z(n1160) );
  NANDN U1379 ( .A(A[39]), .B(n135), .Z(n1161) );
  NANDN U1380 ( .A(n135), .B(A[39]), .Z(n1159) );
  AND U1381 ( .A(n1162), .B(n1163), .Z(n135) );
  NAND U1382 ( .A(B[38]), .B(n1164), .Z(n1163) );
  NANDN U1383 ( .A(A[38]), .B(n137), .Z(n1164) );
  NANDN U1384 ( .A(n137), .B(A[38]), .Z(n1162) );
  AND U1385 ( .A(n1165), .B(n1166), .Z(n137) );
  NAND U1386 ( .A(B[37]), .B(n1167), .Z(n1166) );
  NANDN U1387 ( .A(A[37]), .B(n139), .Z(n1167) );
  NANDN U1388 ( .A(n139), .B(A[37]), .Z(n1165) );
  AND U1389 ( .A(n1168), .B(n1169), .Z(n139) );
  NAND U1390 ( .A(B[36]), .B(n1170), .Z(n1169) );
  NANDN U1391 ( .A(A[36]), .B(n141), .Z(n1170) );
  NANDN U1392 ( .A(n141), .B(A[36]), .Z(n1168) );
  AND U1393 ( .A(n1171), .B(n1172), .Z(n141) );
  NAND U1394 ( .A(B[35]), .B(n1173), .Z(n1172) );
  NANDN U1395 ( .A(A[35]), .B(n143), .Z(n1173) );
  NANDN U1396 ( .A(n143), .B(A[35]), .Z(n1171) );
  AND U1397 ( .A(n1174), .B(n1175), .Z(n143) );
  NAND U1398 ( .A(B[34]), .B(n1176), .Z(n1175) );
  NANDN U1399 ( .A(A[34]), .B(n145), .Z(n1176) );
  NANDN U1400 ( .A(n145), .B(A[34]), .Z(n1174) );
  AND U1401 ( .A(n1177), .B(n1178), .Z(n145) );
  NAND U1402 ( .A(B[33]), .B(n1179), .Z(n1178) );
  NANDN U1403 ( .A(A[33]), .B(n147), .Z(n1179) );
  NANDN U1404 ( .A(n147), .B(A[33]), .Z(n1177) );
  AND U1405 ( .A(n1180), .B(n1181), .Z(n147) );
  NAND U1406 ( .A(B[32]), .B(n1182), .Z(n1181) );
  NANDN U1407 ( .A(A[32]), .B(n149), .Z(n1182) );
  NANDN U1408 ( .A(n149), .B(A[32]), .Z(n1180) );
  AND U1409 ( .A(n1183), .B(n1184), .Z(n149) );
  NAND U1410 ( .A(B[31]), .B(n1185), .Z(n1184) );
  NANDN U1411 ( .A(A[31]), .B(n151), .Z(n1185) );
  NANDN U1412 ( .A(n151), .B(A[31]), .Z(n1183) );
  AND U1413 ( .A(n1186), .B(n1187), .Z(n151) );
  NAND U1414 ( .A(B[30]), .B(n1188), .Z(n1187) );
  NANDN U1415 ( .A(A[30]), .B(n153), .Z(n1188) );
  NANDN U1416 ( .A(n153), .B(A[30]), .Z(n1186) );
  AND U1417 ( .A(n1189), .B(n1190), .Z(n153) );
  NAND U1418 ( .A(B[29]), .B(n1191), .Z(n1190) );
  NANDN U1419 ( .A(A[29]), .B(n157), .Z(n1191) );
  NANDN U1420 ( .A(n157), .B(A[29]), .Z(n1189) );
  AND U1421 ( .A(n1192), .B(n1193), .Z(n157) );
  NAND U1422 ( .A(B[28]), .B(n1194), .Z(n1193) );
  NANDN U1423 ( .A(A[28]), .B(n159), .Z(n1194) );
  NANDN U1424 ( .A(n159), .B(A[28]), .Z(n1192) );
  AND U1425 ( .A(n1195), .B(n1196), .Z(n159) );
  NAND U1426 ( .A(B[27]), .B(n1197), .Z(n1196) );
  NANDN U1427 ( .A(A[27]), .B(n161), .Z(n1197) );
  NANDN U1428 ( .A(n161), .B(A[27]), .Z(n1195) );
  AND U1429 ( .A(n1198), .B(n1199), .Z(n161) );
  NAND U1430 ( .A(B[26]), .B(n1200), .Z(n1199) );
  NANDN U1431 ( .A(A[26]), .B(n163), .Z(n1200) );
  NANDN U1432 ( .A(n163), .B(A[26]), .Z(n1198) );
  AND U1433 ( .A(n1201), .B(n1202), .Z(n163) );
  NAND U1434 ( .A(B[25]), .B(n1203), .Z(n1202) );
  NANDN U1435 ( .A(A[25]), .B(n165), .Z(n1203) );
  NANDN U1436 ( .A(n165), .B(A[25]), .Z(n1201) );
  AND U1437 ( .A(n1204), .B(n1205), .Z(n165) );
  NAND U1438 ( .A(B[24]), .B(n1206), .Z(n1205) );
  NANDN U1439 ( .A(A[24]), .B(n203), .Z(n1206) );
  NANDN U1440 ( .A(n203), .B(A[24]), .Z(n1204) );
  AND U1441 ( .A(n1207), .B(n1208), .Z(n203) );
  NAND U1442 ( .A(B[23]), .B(n1209), .Z(n1208) );
  NANDN U1443 ( .A(A[23]), .B(n255), .Z(n1209) );
  NANDN U1444 ( .A(n255), .B(A[23]), .Z(n1207) );
  AND U1445 ( .A(n1210), .B(n1211), .Z(n255) );
  NAND U1446 ( .A(B[22]), .B(n1212), .Z(n1211) );
  NANDN U1447 ( .A(A[22]), .B(n307), .Z(n1212) );
  NANDN U1448 ( .A(n307), .B(A[22]), .Z(n1210) );
  AND U1449 ( .A(n1213), .B(n1214), .Z(n307) );
  NAND U1450 ( .A(B[21]), .B(n1215), .Z(n1214) );
  NANDN U1451 ( .A(A[21]), .B(n359), .Z(n1215) );
  NANDN U1452 ( .A(n359), .B(A[21]), .Z(n1213) );
  AND U1453 ( .A(n1216), .B(n1217), .Z(n359) );
  NAND U1454 ( .A(B[20]), .B(n1218), .Z(n1217) );
  NANDN U1455 ( .A(A[20]), .B(n411), .Z(n1218) );
  NANDN U1456 ( .A(n411), .B(A[20]), .Z(n1216) );
  AND U1457 ( .A(n1219), .B(n1220), .Z(n411) );
  NAND U1458 ( .A(B[19]), .B(n1221), .Z(n1220) );
  NANDN U1459 ( .A(A[19]), .B(n463), .Z(n1221) );
  NANDN U1460 ( .A(n463), .B(A[19]), .Z(n1219) );
  AND U1461 ( .A(n1222), .B(n1223), .Z(n463) );
  NAND U1462 ( .A(B[18]), .B(n1224), .Z(n1223) );
  NANDN U1463 ( .A(A[18]), .B(n515), .Z(n1224) );
  NANDN U1464 ( .A(n515), .B(A[18]), .Z(n1222) );
  AND U1465 ( .A(n1225), .B(n1226), .Z(n515) );
  NAND U1466 ( .A(B[17]), .B(n1227), .Z(n1226) );
  NANDN U1467 ( .A(A[17]), .B(n567), .Z(n1227) );
  NANDN U1468 ( .A(n567), .B(A[17]), .Z(n1225) );
  AND U1469 ( .A(n1228), .B(n1229), .Z(n567) );
  NAND U1470 ( .A(B[16]), .B(n1230), .Z(n1229) );
  NANDN U1471 ( .A(A[16]), .B(n619), .Z(n1230) );
  NANDN U1472 ( .A(n619), .B(A[16]), .Z(n1228) );
  AND U1473 ( .A(n1231), .B(n1232), .Z(n619) );
  NAND U1474 ( .A(B[15]), .B(n1233), .Z(n1232) );
  NANDN U1475 ( .A(A[15]), .B(n671), .Z(n1233) );
  NANDN U1476 ( .A(n671), .B(A[15]), .Z(n1231) );
  AND U1477 ( .A(n1234), .B(n1235), .Z(n671) );
  NAND U1478 ( .A(B[14]), .B(n1236), .Z(n1235) );
  NANDN U1479 ( .A(A[14]), .B(n723), .Z(n1236) );
  NANDN U1480 ( .A(n723), .B(A[14]), .Z(n1234) );
  AND U1481 ( .A(n1237), .B(n1238), .Z(n723) );
  NAND U1482 ( .A(B[13]), .B(n1239), .Z(n1238) );
  NANDN U1483 ( .A(A[13]), .B(n775), .Z(n1239) );
  NANDN U1484 ( .A(n775), .B(A[13]), .Z(n1237) );
  AND U1485 ( .A(n1240), .B(n1241), .Z(n775) );
  NAND U1486 ( .A(B[12]), .B(n1242), .Z(n1241) );
  NANDN U1487 ( .A(A[12]), .B(n827), .Z(n1242) );
  NANDN U1488 ( .A(n827), .B(A[12]), .Z(n1240) );
  AND U1489 ( .A(n1243), .B(n1244), .Z(n827) );
  NAND U1490 ( .A(B[11]), .B(n1245), .Z(n1244) );
  NANDN U1491 ( .A(A[11]), .B(n879), .Z(n1245) );
  NANDN U1492 ( .A(n879), .B(A[11]), .Z(n1243) );
  AND U1493 ( .A(n1246), .B(n1247), .Z(n879) );
  NAND U1494 ( .A(B[10]), .B(n1248), .Z(n1247) );
  NANDN U1495 ( .A(A[10]), .B(n931), .Z(n1248) );
  NANDN U1496 ( .A(n931), .B(A[10]), .Z(n1246) );
  AND U1497 ( .A(n1249), .B(n1250), .Z(n931) );
  NAND U1498 ( .A(B[9]), .B(n1251), .Z(n1250) );
  OR U1499 ( .A(n1), .B(A[9]), .Z(n1251) );
  NAND U1500 ( .A(A[9]), .B(n1), .Z(n1249) );
  NAND U1501 ( .A(n1252), .B(n1253), .Z(n1) );
  NAND U1502 ( .A(B[8]), .B(n1254), .Z(n1253) );
  NANDN U1503 ( .A(A[8]), .B(n23), .Z(n1254) );
  NANDN U1504 ( .A(n23), .B(A[8]), .Z(n1252) );
  AND U1505 ( .A(n1255), .B(n1256), .Z(n23) );
  NAND U1506 ( .A(B[7]), .B(n1257), .Z(n1256) );
  NANDN U1507 ( .A(A[7]), .B(n45), .Z(n1257) );
  NANDN U1508 ( .A(n45), .B(A[7]), .Z(n1255) );
  AND U1509 ( .A(n1258), .B(n1259), .Z(n45) );
  NAND U1510 ( .A(B[6]), .B(n1260), .Z(n1259) );
  NANDN U1511 ( .A(A[6]), .B(n67), .Z(n1260) );
  NANDN U1512 ( .A(n67), .B(A[6]), .Z(n1258) );
  AND U1513 ( .A(n1261), .B(n1262), .Z(n67) );
  NAND U1514 ( .A(B[5]), .B(n1263), .Z(n1262) );
  NANDN U1515 ( .A(A[5]), .B(n89), .Z(n1263) );
  NANDN U1516 ( .A(n89), .B(A[5]), .Z(n1261) );
  AND U1517 ( .A(n1264), .B(n1265), .Z(n89) );
  NAND U1518 ( .A(B[4]), .B(n1266), .Z(n1265) );
  NANDN U1519 ( .A(A[4]), .B(n111), .Z(n1266) );
  NANDN U1520 ( .A(n111), .B(A[4]), .Z(n1264) );
  AND U1521 ( .A(n1267), .B(n1268), .Z(n111) );
  NAND U1522 ( .A(B[3]), .B(n1269), .Z(n1268) );
  NANDN U1523 ( .A(A[3]), .B(n133), .Z(n1269) );
  NANDN U1524 ( .A(n133), .B(A[3]), .Z(n1267) );
  AND U1525 ( .A(n1270), .B(n1271), .Z(n133) );
  NAND U1526 ( .A(B[2]), .B(n1272), .Z(n1271) );
  OR U1527 ( .A(n155), .B(A[2]), .Z(n1272) );
  NAND U1528 ( .A(A[2]), .B(n155), .Z(n1270) );
  AND U1529 ( .A(B[1]), .B(A[1]), .Z(n155) );
endmodule


module modmult_step_N256_5 ( xregN_1, y, n, zin, zout );
  input [255:0] y;
  input [255:0] n;
  input [257:0] zin;
  output [257:0] zout;
  input xregN_1;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123,
         N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200,
         N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211,
         N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222,
         N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233,
         N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244,
         N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255,
         N256, N257, N258, N259, N260, N261, N262, N264, N265, N266, N267,
         N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278,
         N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289,
         N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300,
         N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311,
         N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322,
         N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333,
         N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344,
         N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366,
         N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377,
         N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410,
         N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421,
         N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432,
         N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443,
         N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454,
         N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465,
         N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476,
         N477, N478, N479, N480, N481, N482, N483, N484, N485, N486, N487,
         N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, N498,
         N499, N500, N501, N502, N503, N504, N505, N506, N507, N508, N509,
         N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, N520,
         N521, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771,
         N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760,
         N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749,
         N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738,
         N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727,
         N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716,
         N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705,
         N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694,
         N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683,
         N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672,
         N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661,
         N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650,
         N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639,
         N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628,
         N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617,
         N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606,
         N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595,
         N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584,
         N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573,
         N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562,
         N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551,
         N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540,
         N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529,
         N528, N527, N526, N525, N522, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039;
  wire   [257:0] z2;
  wire   [257:0] z3;
  wire   SYNOPSYS_UNCONNECTED__0;

  modmult_step_N256_5_DW01_sub_0 sub_129_aco ( .A(z3), .B({1'b0, 1'b0, N780, 
        N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, 
        N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, 
        N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, 
        N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, 
        N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, 
        N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, 
        N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, 
        N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, 
        N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, 
        N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, 
        N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, 
        N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, 
        N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, 
        N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, 
        N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, 
        N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, 
        N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, 
        N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, 
        N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, 
        N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, 
        N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, 
        N527, N526, N525}), .CI(1'b0), .DIFF(zout) );
  modmult_step_N256_5_DW02_mult_0 mult_sub_129_aco ( .A(n), .B(N522), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__0, N780, N779, N778, N777, N776, N775, N774, 
        N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, 
        N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, 
        N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, 
        N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, 
        N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, 
        N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, 
        N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, 
        N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, 
        N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, 
        N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, 
        N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, 
        N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, 
        N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, 
        N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, 
        N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, 
        N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, 
        N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, 
        N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, 
        N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, 
        N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, 
        N533, N532, N531, N530, N529, N528, N527, N526, N525}) );
  modmult_step_N256_5_DW01_cmp2_0 gte_128 ( .A({1'b0, 1'b0, n}), .B(z3), .LEQ(
        1'b1), .TC(1'b0), .LT_LE(N522) );
  modmult_step_N256_5_DW01_sub_1 sub_124 ( .A(z2), .B({1'b0, 1'b0, n}), .CI(
        1'b0), .DIFF({N521, N520, N519, N518, N517, N516, N515, N514, N513, 
        N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, 
        N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, 
        N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, 
        N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, 
        N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, 
        N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, 
        N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, 
        N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, 
        N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, 
        N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, 
        N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, 
        N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, 
        N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, 
        N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, 
        N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, 
        N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, 
        N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, 
        N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, 
        N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, 
        N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, 
        N272, N271, N270, N269, N268, N267, N266, N265, N264}) );
  modmult_step_N256_5_DW01_cmp2_1 gt_123 ( .A({1'b0, 1'b0, n}), .B(z2), .LEQ(
        1'b0), .TC(1'b0), .LT_LE(N262) );
  modmult_step_N256_5_DW01_add_0 add_119 ( .A({zin[256:0], 1'b0}), .B({1'b0, 
        1'b0, y}), .CI(1'b0), .SUM({N261, N260, N259, N258, N257, N256, N255, 
        N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, 
        N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, 
        N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, 
        N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, 
        N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, 
        N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, 
        N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, 
        N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, 
        N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, 
        N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, 
        N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, 
        N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, 
        N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, 
        N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, 
        N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4}) );
  NAND U5 ( .A(n1), .B(n2), .Z(z3[9]) );
  NANDN U6 ( .A(N262), .B(z2[9]), .Z(n2) );
  NANDN U7 ( .A(n3), .B(N273), .Z(n1) );
  NAND U8 ( .A(n4), .B(n5), .Z(z3[99]) );
  NANDN U9 ( .A(N262), .B(z2[99]), .Z(n5) );
  NANDN U10 ( .A(n3), .B(N363), .Z(n4) );
  NAND U11 ( .A(n6), .B(n7), .Z(z3[98]) );
  NANDN U17 ( .A(N262), .B(z2[98]), .Z(n7) );
  NANDN U18 ( .A(n3), .B(N362), .Z(n6) );
  NAND U19 ( .A(n8), .B(n9), .Z(z3[97]) );
  NANDN U20 ( .A(N262), .B(z2[97]), .Z(n9) );
  NANDN U21 ( .A(n3), .B(N361), .Z(n8) );
  NAND U22 ( .A(n10), .B(n11), .Z(z3[96]) );
  NANDN U23 ( .A(N262), .B(z2[96]), .Z(n11) );
  NANDN U24 ( .A(n3), .B(N360), .Z(n10) );
  NAND U25 ( .A(n12), .B(n13), .Z(z3[95]) );
  NANDN U26 ( .A(N262), .B(z2[95]), .Z(n13) );
  NANDN U27 ( .A(n3), .B(N359), .Z(n12) );
  NAND U28 ( .A(n14), .B(n23), .Z(z3[94]) );
  NANDN U29 ( .A(N262), .B(z2[94]), .Z(n23) );
  NANDN U30 ( .A(n3), .B(N358), .Z(n14) );
  NAND U31 ( .A(n24), .B(n25), .Z(z3[93]) );
  NANDN U32 ( .A(N262), .B(z2[93]), .Z(n25) );
  NANDN U33 ( .A(n3), .B(N357), .Z(n24) );
  NAND U34 ( .A(n26), .B(n27), .Z(z3[92]) );
  NANDN U35 ( .A(N262), .B(z2[92]), .Z(n27) );
  NANDN U36 ( .A(n3), .B(N356), .Z(n26) );
  NAND U37 ( .A(n28), .B(n29), .Z(z3[91]) );
  NANDN U38 ( .A(N262), .B(z2[91]), .Z(n29) );
  NANDN U39 ( .A(n3), .B(N355), .Z(n28) );
  NAND U40 ( .A(n30), .B(n31), .Z(z3[90]) );
  NANDN U41 ( .A(N262), .B(z2[90]), .Z(n31) );
  NANDN U42 ( .A(n3), .B(N354), .Z(n30) );
  NAND U43 ( .A(n32), .B(n33), .Z(z3[8]) );
  NANDN U44 ( .A(N262), .B(z2[8]), .Z(n33) );
  NANDN U45 ( .A(n3), .B(N272), .Z(n32) );
  NAND U46 ( .A(n34), .B(n35), .Z(z3[89]) );
  NANDN U47 ( .A(N262), .B(z2[89]), .Z(n35) );
  NANDN U48 ( .A(n3), .B(N353), .Z(n34) );
  NAND U49 ( .A(n36), .B(n37), .Z(z3[88]) );
  NANDN U50 ( .A(N262), .B(z2[88]), .Z(n37) );
  NANDN U51 ( .A(n3), .B(N352), .Z(n36) );
  NAND U52 ( .A(n38), .B(n39), .Z(z3[87]) );
  NANDN U53 ( .A(N262), .B(z2[87]), .Z(n39) );
  NANDN U54 ( .A(n3), .B(N351), .Z(n38) );
  NAND U55 ( .A(n40), .B(n41), .Z(z3[86]) );
  NANDN U56 ( .A(N262), .B(z2[86]), .Z(n41) );
  NANDN U57 ( .A(n3), .B(N350), .Z(n40) );
  NAND U58 ( .A(n42), .B(n43), .Z(z3[85]) );
  NANDN U59 ( .A(N262), .B(z2[85]), .Z(n43) );
  NANDN U60 ( .A(n3), .B(N349), .Z(n42) );
  NAND U61 ( .A(n44), .B(n45), .Z(z3[84]) );
  NANDN U62 ( .A(N262), .B(z2[84]), .Z(n45) );
  NANDN U63 ( .A(n3), .B(N348), .Z(n44) );
  NAND U64 ( .A(n46), .B(n47), .Z(z3[83]) );
  NANDN U65 ( .A(N262), .B(z2[83]), .Z(n47) );
  NANDN U66 ( .A(n3), .B(N347), .Z(n46) );
  NAND U67 ( .A(n48), .B(n49), .Z(z3[82]) );
  NANDN U68 ( .A(N262), .B(z2[82]), .Z(n49) );
  NANDN U69 ( .A(n3), .B(N346), .Z(n48) );
  NAND U70 ( .A(n50), .B(n51), .Z(z3[81]) );
  NANDN U71 ( .A(N262), .B(z2[81]), .Z(n51) );
  NANDN U72 ( .A(n3), .B(N345), .Z(n50) );
  NAND U73 ( .A(n52), .B(n53), .Z(z3[80]) );
  NANDN U74 ( .A(N262), .B(z2[80]), .Z(n53) );
  NANDN U75 ( .A(n3), .B(N344), .Z(n52) );
  NAND U76 ( .A(n54), .B(n55), .Z(z3[7]) );
  NANDN U77 ( .A(N262), .B(z2[7]), .Z(n55) );
  NANDN U78 ( .A(n3), .B(N271), .Z(n54) );
  NAND U79 ( .A(n56), .B(n57), .Z(z3[79]) );
  NANDN U80 ( .A(N262), .B(z2[79]), .Z(n57) );
  NANDN U81 ( .A(n3), .B(N343), .Z(n56) );
  NAND U82 ( .A(n58), .B(n59), .Z(z3[78]) );
  NANDN U83 ( .A(N262), .B(z2[78]), .Z(n59) );
  NANDN U84 ( .A(n3), .B(N342), .Z(n58) );
  NAND U85 ( .A(n60), .B(n61), .Z(z3[77]) );
  NANDN U86 ( .A(N262), .B(z2[77]), .Z(n61) );
  NANDN U87 ( .A(n3), .B(N341), .Z(n60) );
  NAND U88 ( .A(n62), .B(n63), .Z(z3[76]) );
  NANDN U89 ( .A(N262), .B(z2[76]), .Z(n63) );
  NANDN U90 ( .A(n3), .B(N340), .Z(n62) );
  NAND U91 ( .A(n64), .B(n65), .Z(z3[75]) );
  NANDN U92 ( .A(N262), .B(z2[75]), .Z(n65) );
  NANDN U93 ( .A(n3), .B(N339), .Z(n64) );
  NAND U94 ( .A(n66), .B(n67), .Z(z3[74]) );
  NANDN U95 ( .A(N262), .B(z2[74]), .Z(n67) );
  NANDN U96 ( .A(n3), .B(N338), .Z(n66) );
  NAND U97 ( .A(n68), .B(n69), .Z(z3[73]) );
  NANDN U98 ( .A(N262), .B(z2[73]), .Z(n69) );
  NANDN U99 ( .A(n3), .B(N337), .Z(n68) );
  NAND U100 ( .A(n70), .B(n71), .Z(z3[72]) );
  NANDN U101 ( .A(N262), .B(z2[72]), .Z(n71) );
  NANDN U102 ( .A(n3), .B(N336), .Z(n70) );
  NAND U103 ( .A(n72), .B(n73), .Z(z3[71]) );
  NANDN U104 ( .A(N262), .B(z2[71]), .Z(n73) );
  NANDN U105 ( .A(n3), .B(N335), .Z(n72) );
  NAND U106 ( .A(n74), .B(n75), .Z(z3[70]) );
  NANDN U107 ( .A(N262), .B(z2[70]), .Z(n75) );
  NANDN U108 ( .A(n3), .B(N334), .Z(n74) );
  NAND U109 ( .A(n76), .B(n77), .Z(z3[6]) );
  NANDN U110 ( .A(N262), .B(z2[6]), .Z(n77) );
  NANDN U111 ( .A(n3), .B(N270), .Z(n76) );
  NAND U112 ( .A(n78), .B(n79), .Z(z3[69]) );
  NANDN U113 ( .A(N262), .B(z2[69]), .Z(n79) );
  NANDN U114 ( .A(n3), .B(N333), .Z(n78) );
  NAND U115 ( .A(n80), .B(n81), .Z(z3[68]) );
  NANDN U116 ( .A(N262), .B(z2[68]), .Z(n81) );
  NANDN U117 ( .A(n3), .B(N332), .Z(n80) );
  NAND U118 ( .A(n82), .B(n83), .Z(z3[67]) );
  NANDN U119 ( .A(N262), .B(z2[67]), .Z(n83) );
  NANDN U120 ( .A(n3), .B(N331), .Z(n82) );
  NAND U121 ( .A(n84), .B(n85), .Z(z3[66]) );
  NANDN U122 ( .A(N262), .B(z2[66]), .Z(n85) );
  NANDN U123 ( .A(n3), .B(N330), .Z(n84) );
  NAND U124 ( .A(n86), .B(n87), .Z(z3[65]) );
  NANDN U125 ( .A(N262), .B(z2[65]), .Z(n87) );
  NANDN U126 ( .A(n3), .B(N329), .Z(n86) );
  NAND U127 ( .A(n88), .B(n89), .Z(z3[64]) );
  NANDN U128 ( .A(N262), .B(z2[64]), .Z(n89) );
  NANDN U129 ( .A(n3), .B(N328), .Z(n88) );
  NAND U130 ( .A(n90), .B(n91), .Z(z3[63]) );
  NANDN U131 ( .A(N262), .B(z2[63]), .Z(n91) );
  NANDN U132 ( .A(n3), .B(N327), .Z(n90) );
  NAND U133 ( .A(n92), .B(n93), .Z(z3[62]) );
  NANDN U134 ( .A(N262), .B(z2[62]), .Z(n93) );
  NANDN U135 ( .A(n3), .B(N326), .Z(n92) );
  NAND U136 ( .A(n94), .B(n95), .Z(z3[61]) );
  NANDN U137 ( .A(N262), .B(z2[61]), .Z(n95) );
  NANDN U138 ( .A(n3), .B(N325), .Z(n94) );
  NAND U139 ( .A(n96), .B(n97), .Z(z3[60]) );
  NANDN U140 ( .A(N262), .B(z2[60]), .Z(n97) );
  NANDN U141 ( .A(n3), .B(N324), .Z(n96) );
  NAND U142 ( .A(n98), .B(n99), .Z(z3[5]) );
  NANDN U143 ( .A(N262), .B(z2[5]), .Z(n99) );
  NANDN U144 ( .A(n3), .B(N269), .Z(n98) );
  NAND U145 ( .A(n100), .B(n101), .Z(z3[59]) );
  NANDN U146 ( .A(N262), .B(z2[59]), .Z(n101) );
  NANDN U147 ( .A(n3), .B(N323), .Z(n100) );
  NAND U148 ( .A(n102), .B(n103), .Z(z3[58]) );
  NANDN U149 ( .A(N262), .B(z2[58]), .Z(n103) );
  NANDN U150 ( .A(n3), .B(N322), .Z(n102) );
  NAND U151 ( .A(n104), .B(n105), .Z(z3[57]) );
  NANDN U152 ( .A(N262), .B(z2[57]), .Z(n105) );
  NANDN U153 ( .A(n3), .B(N321), .Z(n104) );
  NAND U154 ( .A(n106), .B(n107), .Z(z3[56]) );
  NANDN U155 ( .A(N262), .B(z2[56]), .Z(n107) );
  NANDN U156 ( .A(n3), .B(N320), .Z(n106) );
  NAND U157 ( .A(n108), .B(n109), .Z(z3[55]) );
  NANDN U158 ( .A(N262), .B(z2[55]), .Z(n109) );
  NANDN U159 ( .A(n3), .B(N319), .Z(n108) );
  NAND U160 ( .A(n110), .B(n111), .Z(z3[54]) );
  NANDN U161 ( .A(N262), .B(z2[54]), .Z(n111) );
  NANDN U162 ( .A(n3), .B(N318), .Z(n110) );
  NAND U163 ( .A(n112), .B(n113), .Z(z3[53]) );
  NANDN U164 ( .A(N262), .B(z2[53]), .Z(n113) );
  NANDN U165 ( .A(n3), .B(N317), .Z(n112) );
  NAND U166 ( .A(n114), .B(n115), .Z(z3[52]) );
  NANDN U167 ( .A(N262), .B(z2[52]), .Z(n115) );
  NANDN U168 ( .A(n3), .B(N316), .Z(n114) );
  NAND U169 ( .A(n116), .B(n117), .Z(z3[51]) );
  NANDN U170 ( .A(N262), .B(z2[51]), .Z(n117) );
  NANDN U171 ( .A(n3), .B(N315), .Z(n116) );
  NAND U172 ( .A(n118), .B(n119), .Z(z3[50]) );
  NANDN U173 ( .A(N262), .B(z2[50]), .Z(n119) );
  NANDN U174 ( .A(n3), .B(N314), .Z(n118) );
  NAND U175 ( .A(n120), .B(n121), .Z(z3[4]) );
  NANDN U176 ( .A(N262), .B(z2[4]), .Z(n121) );
  NANDN U177 ( .A(n3), .B(N268), .Z(n120) );
  NAND U178 ( .A(n122), .B(n123), .Z(z3[49]) );
  NANDN U179 ( .A(N262), .B(z2[49]), .Z(n123) );
  NANDN U180 ( .A(n3), .B(N313), .Z(n122) );
  NAND U181 ( .A(n124), .B(n125), .Z(z3[48]) );
  NANDN U182 ( .A(N262), .B(z2[48]), .Z(n125) );
  NANDN U183 ( .A(n3), .B(N312), .Z(n124) );
  NAND U184 ( .A(n126), .B(n127), .Z(z3[47]) );
  NANDN U185 ( .A(N262), .B(z2[47]), .Z(n127) );
  NANDN U186 ( .A(n3), .B(N311), .Z(n126) );
  NAND U187 ( .A(n128), .B(n129), .Z(z3[46]) );
  NANDN U188 ( .A(N262), .B(z2[46]), .Z(n129) );
  NANDN U189 ( .A(n3), .B(N310), .Z(n128) );
  NAND U190 ( .A(n130), .B(n131), .Z(z3[45]) );
  NANDN U191 ( .A(N262), .B(z2[45]), .Z(n131) );
  NANDN U192 ( .A(n3), .B(N309), .Z(n130) );
  NAND U193 ( .A(n132), .B(n133), .Z(z3[44]) );
  NANDN U194 ( .A(N262), .B(z2[44]), .Z(n133) );
  NANDN U195 ( .A(n3), .B(N308), .Z(n132) );
  NAND U196 ( .A(n134), .B(n135), .Z(z3[43]) );
  NANDN U197 ( .A(N262), .B(z2[43]), .Z(n135) );
  NANDN U198 ( .A(n3), .B(N307), .Z(n134) );
  NAND U199 ( .A(n136), .B(n137), .Z(z3[42]) );
  NANDN U200 ( .A(N262), .B(z2[42]), .Z(n137) );
  NANDN U201 ( .A(n3), .B(N306), .Z(n136) );
  NAND U202 ( .A(n138), .B(n139), .Z(z3[41]) );
  NANDN U203 ( .A(N262), .B(z2[41]), .Z(n139) );
  NANDN U204 ( .A(n3), .B(N305), .Z(n138) );
  NAND U205 ( .A(n140), .B(n141), .Z(z3[40]) );
  NANDN U206 ( .A(N262), .B(z2[40]), .Z(n141) );
  NANDN U207 ( .A(n3), .B(N304), .Z(n140) );
  NAND U208 ( .A(n142), .B(n143), .Z(z3[3]) );
  NANDN U209 ( .A(N262), .B(z2[3]), .Z(n143) );
  NANDN U210 ( .A(n3), .B(N267), .Z(n142) );
  NAND U211 ( .A(n144), .B(n145), .Z(z3[39]) );
  NANDN U212 ( .A(N262), .B(z2[39]), .Z(n145) );
  NANDN U213 ( .A(n3), .B(N303), .Z(n144) );
  NAND U214 ( .A(n146), .B(n147), .Z(z3[38]) );
  NANDN U215 ( .A(N262), .B(z2[38]), .Z(n147) );
  NANDN U216 ( .A(n3), .B(N302), .Z(n146) );
  NAND U217 ( .A(n148), .B(n149), .Z(z3[37]) );
  NANDN U218 ( .A(N262), .B(z2[37]), .Z(n149) );
  NANDN U219 ( .A(n3), .B(N301), .Z(n148) );
  NAND U220 ( .A(n150), .B(n151), .Z(z3[36]) );
  NANDN U221 ( .A(N262), .B(z2[36]), .Z(n151) );
  NANDN U222 ( .A(n3), .B(N300), .Z(n150) );
  NAND U223 ( .A(n152), .B(n153), .Z(z3[35]) );
  NANDN U224 ( .A(N262), .B(z2[35]), .Z(n153) );
  NANDN U225 ( .A(n3), .B(N299), .Z(n152) );
  NAND U226 ( .A(n154), .B(n155), .Z(z3[34]) );
  NANDN U227 ( .A(N262), .B(z2[34]), .Z(n155) );
  NANDN U228 ( .A(n3), .B(N298), .Z(n154) );
  NAND U229 ( .A(n156), .B(n157), .Z(z3[33]) );
  NANDN U230 ( .A(N262), .B(z2[33]), .Z(n157) );
  NANDN U231 ( .A(n3), .B(N297), .Z(n156) );
  NAND U232 ( .A(n158), .B(n159), .Z(z3[32]) );
  NANDN U233 ( .A(N262), .B(z2[32]), .Z(n159) );
  NANDN U234 ( .A(n3), .B(N296), .Z(n158) );
  NAND U235 ( .A(n160), .B(n161), .Z(z3[31]) );
  NANDN U236 ( .A(N262), .B(z2[31]), .Z(n161) );
  NANDN U237 ( .A(n3), .B(N295), .Z(n160) );
  NAND U238 ( .A(n162), .B(n163), .Z(z3[30]) );
  NANDN U239 ( .A(N262), .B(z2[30]), .Z(n163) );
  NANDN U240 ( .A(n3), .B(N294), .Z(n162) );
  NAND U241 ( .A(n164), .B(n165), .Z(z3[2]) );
  NANDN U242 ( .A(N262), .B(z2[2]), .Z(n165) );
  NANDN U243 ( .A(n3), .B(N266), .Z(n164) );
  NAND U244 ( .A(n166), .B(n167), .Z(z3[29]) );
  NANDN U245 ( .A(N262), .B(z2[29]), .Z(n167) );
  NANDN U246 ( .A(n3), .B(N293), .Z(n166) );
  NAND U247 ( .A(n168), .B(n169), .Z(z3[28]) );
  NANDN U248 ( .A(N262), .B(z2[28]), .Z(n169) );
  NANDN U249 ( .A(n3), .B(N292), .Z(n168) );
  NAND U250 ( .A(n170), .B(n171), .Z(z3[27]) );
  NANDN U251 ( .A(N262), .B(z2[27]), .Z(n171) );
  NANDN U252 ( .A(n3), .B(N291), .Z(n170) );
  NAND U253 ( .A(n172), .B(n173), .Z(z3[26]) );
  NANDN U254 ( .A(N262), .B(z2[26]), .Z(n173) );
  NANDN U255 ( .A(n3), .B(N290), .Z(n172) );
  NAND U256 ( .A(n174), .B(n175), .Z(z3[25]) );
  NANDN U257 ( .A(N262), .B(z2[25]), .Z(n175) );
  NANDN U258 ( .A(n3), .B(N289), .Z(n174) );
  NAND U259 ( .A(n176), .B(n177), .Z(z3[257]) );
  NANDN U260 ( .A(N262), .B(z2[257]), .Z(n177) );
  NANDN U261 ( .A(n3), .B(N521), .Z(n176) );
  NAND U262 ( .A(n178), .B(n179), .Z(z3[256]) );
  NANDN U263 ( .A(N262), .B(z2[256]), .Z(n179) );
  NANDN U264 ( .A(n3), .B(N520), .Z(n178) );
  NAND U265 ( .A(n180), .B(n181), .Z(z3[255]) );
  NANDN U266 ( .A(N262), .B(z2[255]), .Z(n181) );
  NANDN U267 ( .A(n3), .B(N519), .Z(n180) );
  NAND U268 ( .A(n182), .B(n183), .Z(z3[254]) );
  NANDN U269 ( .A(N262), .B(z2[254]), .Z(n183) );
  NANDN U270 ( .A(n3), .B(N518), .Z(n182) );
  NAND U271 ( .A(n184), .B(n185), .Z(z3[253]) );
  NANDN U272 ( .A(N262), .B(z2[253]), .Z(n185) );
  NANDN U273 ( .A(n3), .B(N517), .Z(n184) );
  NAND U274 ( .A(n186), .B(n187), .Z(z3[252]) );
  NANDN U275 ( .A(N262), .B(z2[252]), .Z(n187) );
  NANDN U276 ( .A(n3), .B(N516), .Z(n186) );
  NAND U277 ( .A(n188), .B(n189), .Z(z3[251]) );
  NANDN U278 ( .A(N262), .B(z2[251]), .Z(n189) );
  NANDN U279 ( .A(n3), .B(N515), .Z(n188) );
  NAND U280 ( .A(n190), .B(n191), .Z(z3[250]) );
  NANDN U281 ( .A(N262), .B(z2[250]), .Z(n191) );
  NANDN U282 ( .A(n3), .B(N514), .Z(n190) );
  NAND U283 ( .A(n192), .B(n193), .Z(z3[24]) );
  NANDN U284 ( .A(N262), .B(z2[24]), .Z(n193) );
  NANDN U285 ( .A(n3), .B(N288), .Z(n192) );
  NAND U286 ( .A(n194), .B(n195), .Z(z3[249]) );
  NANDN U287 ( .A(N262), .B(z2[249]), .Z(n195) );
  NANDN U288 ( .A(n3), .B(N513), .Z(n194) );
  NAND U289 ( .A(n196), .B(n197), .Z(z3[248]) );
  NANDN U290 ( .A(N262), .B(z2[248]), .Z(n197) );
  NANDN U291 ( .A(n3), .B(N512), .Z(n196) );
  NAND U292 ( .A(n198), .B(n199), .Z(z3[247]) );
  NANDN U293 ( .A(N262), .B(z2[247]), .Z(n199) );
  NANDN U294 ( .A(n3), .B(N511), .Z(n198) );
  NAND U295 ( .A(n200), .B(n201), .Z(z3[246]) );
  NANDN U296 ( .A(N262), .B(z2[246]), .Z(n201) );
  NANDN U297 ( .A(n3), .B(N510), .Z(n200) );
  NAND U298 ( .A(n202), .B(n203), .Z(z3[245]) );
  NANDN U299 ( .A(N262), .B(z2[245]), .Z(n203) );
  NANDN U300 ( .A(n3), .B(N509), .Z(n202) );
  NAND U301 ( .A(n204), .B(n205), .Z(z3[244]) );
  NANDN U302 ( .A(N262), .B(z2[244]), .Z(n205) );
  NANDN U303 ( .A(n3), .B(N508), .Z(n204) );
  NAND U304 ( .A(n206), .B(n207), .Z(z3[243]) );
  NANDN U305 ( .A(N262), .B(z2[243]), .Z(n207) );
  NANDN U306 ( .A(n3), .B(N507), .Z(n206) );
  NAND U307 ( .A(n208), .B(n209), .Z(z3[242]) );
  NANDN U308 ( .A(N262), .B(z2[242]), .Z(n209) );
  NANDN U309 ( .A(n3), .B(N506), .Z(n208) );
  NAND U310 ( .A(n210), .B(n211), .Z(z3[241]) );
  NANDN U311 ( .A(N262), .B(z2[241]), .Z(n211) );
  NANDN U312 ( .A(n3), .B(N505), .Z(n210) );
  NAND U313 ( .A(n212), .B(n213), .Z(z3[240]) );
  NANDN U314 ( .A(N262), .B(z2[240]), .Z(n213) );
  NANDN U315 ( .A(n3), .B(N504), .Z(n212) );
  NAND U316 ( .A(n214), .B(n215), .Z(z3[23]) );
  NANDN U317 ( .A(N262), .B(z2[23]), .Z(n215) );
  NANDN U318 ( .A(n3), .B(N287), .Z(n214) );
  NAND U319 ( .A(n216), .B(n217), .Z(z3[239]) );
  NANDN U320 ( .A(N262), .B(z2[239]), .Z(n217) );
  NANDN U321 ( .A(n3), .B(N503), .Z(n216) );
  NAND U322 ( .A(n218), .B(n219), .Z(z3[238]) );
  NANDN U323 ( .A(N262), .B(z2[238]), .Z(n219) );
  NANDN U324 ( .A(n3), .B(N502), .Z(n218) );
  NAND U325 ( .A(n220), .B(n221), .Z(z3[237]) );
  NANDN U326 ( .A(N262), .B(z2[237]), .Z(n221) );
  NANDN U327 ( .A(n3), .B(N501), .Z(n220) );
  NAND U328 ( .A(n222), .B(n223), .Z(z3[236]) );
  NANDN U329 ( .A(N262), .B(z2[236]), .Z(n223) );
  NANDN U330 ( .A(n3), .B(N500), .Z(n222) );
  NAND U331 ( .A(n224), .B(n225), .Z(z3[235]) );
  NANDN U332 ( .A(N262), .B(z2[235]), .Z(n225) );
  NANDN U333 ( .A(n3), .B(N499), .Z(n224) );
  NAND U334 ( .A(n226), .B(n227), .Z(z3[234]) );
  NANDN U335 ( .A(N262), .B(z2[234]), .Z(n227) );
  NANDN U336 ( .A(n3), .B(N498), .Z(n226) );
  NAND U337 ( .A(n228), .B(n229), .Z(z3[233]) );
  NANDN U338 ( .A(N262), .B(z2[233]), .Z(n229) );
  NANDN U339 ( .A(n3), .B(N497), .Z(n228) );
  NAND U340 ( .A(n230), .B(n231), .Z(z3[232]) );
  NANDN U341 ( .A(N262), .B(z2[232]), .Z(n231) );
  NANDN U342 ( .A(n3), .B(N496), .Z(n230) );
  NAND U343 ( .A(n232), .B(n233), .Z(z3[231]) );
  NANDN U344 ( .A(N262), .B(z2[231]), .Z(n233) );
  NANDN U345 ( .A(n3), .B(N495), .Z(n232) );
  NAND U346 ( .A(n234), .B(n235), .Z(z3[230]) );
  NANDN U347 ( .A(N262), .B(z2[230]), .Z(n235) );
  NANDN U348 ( .A(n3), .B(N494), .Z(n234) );
  NAND U349 ( .A(n236), .B(n237), .Z(z3[22]) );
  NANDN U350 ( .A(N262), .B(z2[22]), .Z(n237) );
  NANDN U351 ( .A(n3), .B(N286), .Z(n236) );
  NAND U352 ( .A(n238), .B(n239), .Z(z3[229]) );
  NANDN U353 ( .A(N262), .B(z2[229]), .Z(n239) );
  NANDN U354 ( .A(n3), .B(N493), .Z(n238) );
  NAND U355 ( .A(n240), .B(n241), .Z(z3[228]) );
  NANDN U356 ( .A(N262), .B(z2[228]), .Z(n241) );
  NANDN U357 ( .A(n3), .B(N492), .Z(n240) );
  NAND U358 ( .A(n242), .B(n243), .Z(z3[227]) );
  NANDN U359 ( .A(N262), .B(z2[227]), .Z(n243) );
  NANDN U360 ( .A(n3), .B(N491), .Z(n242) );
  NAND U361 ( .A(n244), .B(n245), .Z(z3[226]) );
  NANDN U362 ( .A(N262), .B(z2[226]), .Z(n245) );
  NANDN U363 ( .A(n3), .B(N490), .Z(n244) );
  NAND U364 ( .A(n246), .B(n247), .Z(z3[225]) );
  NANDN U365 ( .A(N262), .B(z2[225]), .Z(n247) );
  NANDN U366 ( .A(n3), .B(N489), .Z(n246) );
  NAND U367 ( .A(n248), .B(n249), .Z(z3[224]) );
  NANDN U368 ( .A(N262), .B(z2[224]), .Z(n249) );
  NANDN U369 ( .A(n3), .B(N488), .Z(n248) );
  NAND U370 ( .A(n250), .B(n251), .Z(z3[223]) );
  NANDN U371 ( .A(N262), .B(z2[223]), .Z(n251) );
  NANDN U372 ( .A(n3), .B(N487), .Z(n250) );
  NAND U373 ( .A(n252), .B(n253), .Z(z3[222]) );
  NANDN U374 ( .A(N262), .B(z2[222]), .Z(n253) );
  NANDN U375 ( .A(n3), .B(N486), .Z(n252) );
  NAND U376 ( .A(n254), .B(n255), .Z(z3[221]) );
  NANDN U377 ( .A(N262), .B(z2[221]), .Z(n255) );
  NANDN U378 ( .A(n3), .B(N485), .Z(n254) );
  NAND U379 ( .A(n256), .B(n257), .Z(z3[220]) );
  NANDN U380 ( .A(N262), .B(z2[220]), .Z(n257) );
  NANDN U381 ( .A(n3), .B(N484), .Z(n256) );
  NAND U382 ( .A(n258), .B(n259), .Z(z3[21]) );
  NANDN U383 ( .A(N262), .B(z2[21]), .Z(n259) );
  NANDN U384 ( .A(n3), .B(N285), .Z(n258) );
  NAND U385 ( .A(n260), .B(n261), .Z(z3[219]) );
  NANDN U386 ( .A(N262), .B(z2[219]), .Z(n261) );
  NANDN U387 ( .A(n3), .B(N483), .Z(n260) );
  NAND U388 ( .A(n262), .B(n263), .Z(z3[218]) );
  NANDN U389 ( .A(N262), .B(z2[218]), .Z(n263) );
  NANDN U390 ( .A(n3), .B(N482), .Z(n262) );
  NAND U391 ( .A(n264), .B(n265), .Z(z3[217]) );
  NANDN U392 ( .A(N262), .B(z2[217]), .Z(n265) );
  NANDN U393 ( .A(n3), .B(N481), .Z(n264) );
  NAND U394 ( .A(n266), .B(n267), .Z(z3[216]) );
  NANDN U395 ( .A(N262), .B(z2[216]), .Z(n267) );
  NANDN U396 ( .A(n3), .B(N480), .Z(n266) );
  NAND U397 ( .A(n268), .B(n269), .Z(z3[215]) );
  NANDN U398 ( .A(N262), .B(z2[215]), .Z(n269) );
  NANDN U399 ( .A(n3), .B(N479), .Z(n268) );
  NAND U400 ( .A(n270), .B(n271), .Z(z3[214]) );
  NANDN U401 ( .A(N262), .B(z2[214]), .Z(n271) );
  NANDN U402 ( .A(n3), .B(N478), .Z(n270) );
  NAND U403 ( .A(n272), .B(n273), .Z(z3[213]) );
  NANDN U404 ( .A(N262), .B(z2[213]), .Z(n273) );
  NANDN U405 ( .A(n3), .B(N477), .Z(n272) );
  NAND U406 ( .A(n274), .B(n275), .Z(z3[212]) );
  NANDN U407 ( .A(N262), .B(z2[212]), .Z(n275) );
  NANDN U408 ( .A(n3), .B(N476), .Z(n274) );
  NAND U409 ( .A(n276), .B(n277), .Z(z3[211]) );
  NANDN U410 ( .A(N262), .B(z2[211]), .Z(n277) );
  NANDN U411 ( .A(n3), .B(N475), .Z(n276) );
  NAND U412 ( .A(n278), .B(n279), .Z(z3[210]) );
  NANDN U413 ( .A(N262), .B(z2[210]), .Z(n279) );
  NANDN U414 ( .A(n3), .B(N474), .Z(n278) );
  NAND U415 ( .A(n280), .B(n281), .Z(z3[20]) );
  NANDN U416 ( .A(N262), .B(z2[20]), .Z(n281) );
  NANDN U417 ( .A(n3), .B(N284), .Z(n280) );
  NAND U418 ( .A(n282), .B(n283), .Z(z3[209]) );
  NANDN U419 ( .A(N262), .B(z2[209]), .Z(n283) );
  NANDN U420 ( .A(n3), .B(N473), .Z(n282) );
  NAND U421 ( .A(n284), .B(n285), .Z(z3[208]) );
  NANDN U422 ( .A(N262), .B(z2[208]), .Z(n285) );
  NANDN U423 ( .A(n3), .B(N472), .Z(n284) );
  NAND U424 ( .A(n286), .B(n287), .Z(z3[207]) );
  NANDN U425 ( .A(N262), .B(z2[207]), .Z(n287) );
  NANDN U426 ( .A(n3), .B(N471), .Z(n286) );
  NAND U427 ( .A(n288), .B(n289), .Z(z3[206]) );
  NANDN U428 ( .A(N262), .B(z2[206]), .Z(n289) );
  NANDN U429 ( .A(n3), .B(N470), .Z(n288) );
  NAND U430 ( .A(n290), .B(n291), .Z(z3[205]) );
  NANDN U431 ( .A(N262), .B(z2[205]), .Z(n291) );
  NANDN U432 ( .A(n3), .B(N469), .Z(n290) );
  NAND U433 ( .A(n292), .B(n293), .Z(z3[204]) );
  NANDN U434 ( .A(N262), .B(z2[204]), .Z(n293) );
  NANDN U435 ( .A(n3), .B(N468), .Z(n292) );
  NAND U436 ( .A(n294), .B(n295), .Z(z3[203]) );
  NANDN U437 ( .A(N262), .B(z2[203]), .Z(n295) );
  NANDN U438 ( .A(n3), .B(N467), .Z(n294) );
  NAND U439 ( .A(n296), .B(n297), .Z(z3[202]) );
  NANDN U440 ( .A(N262), .B(z2[202]), .Z(n297) );
  NANDN U441 ( .A(n3), .B(N466), .Z(n296) );
  NAND U442 ( .A(n298), .B(n299), .Z(z3[201]) );
  NANDN U443 ( .A(N262), .B(z2[201]), .Z(n299) );
  NANDN U444 ( .A(n3), .B(N465), .Z(n298) );
  NAND U445 ( .A(n300), .B(n301), .Z(z3[200]) );
  NANDN U446 ( .A(N262), .B(z2[200]), .Z(n301) );
  NANDN U447 ( .A(n3), .B(N464), .Z(n300) );
  NAND U448 ( .A(n302), .B(n303), .Z(z3[1]) );
  NANDN U449 ( .A(N262), .B(z2[1]), .Z(n303) );
  NANDN U450 ( .A(n3), .B(N265), .Z(n302) );
  NAND U451 ( .A(n304), .B(n305), .Z(z3[19]) );
  NANDN U452 ( .A(N262), .B(z2[19]), .Z(n305) );
  NANDN U453 ( .A(n3), .B(N283), .Z(n304) );
  NAND U454 ( .A(n306), .B(n307), .Z(z3[199]) );
  NANDN U455 ( .A(N262), .B(z2[199]), .Z(n307) );
  NANDN U456 ( .A(n3), .B(N463), .Z(n306) );
  NAND U457 ( .A(n308), .B(n309), .Z(z3[198]) );
  NANDN U458 ( .A(N262), .B(z2[198]), .Z(n309) );
  NANDN U459 ( .A(n3), .B(N462), .Z(n308) );
  NAND U460 ( .A(n310), .B(n311), .Z(z3[197]) );
  NANDN U461 ( .A(N262), .B(z2[197]), .Z(n311) );
  NANDN U462 ( .A(n3), .B(N461), .Z(n310) );
  NAND U463 ( .A(n312), .B(n313), .Z(z3[196]) );
  NANDN U464 ( .A(N262), .B(z2[196]), .Z(n313) );
  NANDN U465 ( .A(n3), .B(N460), .Z(n312) );
  NAND U466 ( .A(n314), .B(n315), .Z(z3[195]) );
  NANDN U467 ( .A(N262), .B(z2[195]), .Z(n315) );
  NANDN U468 ( .A(n3), .B(N459), .Z(n314) );
  NAND U469 ( .A(n316), .B(n317), .Z(z3[194]) );
  NANDN U470 ( .A(N262), .B(z2[194]), .Z(n317) );
  NANDN U471 ( .A(n3), .B(N458), .Z(n316) );
  NAND U472 ( .A(n318), .B(n319), .Z(z3[193]) );
  NANDN U473 ( .A(N262), .B(z2[193]), .Z(n319) );
  NANDN U474 ( .A(n3), .B(N457), .Z(n318) );
  NAND U475 ( .A(n320), .B(n321), .Z(z3[192]) );
  NANDN U476 ( .A(N262), .B(z2[192]), .Z(n321) );
  NANDN U477 ( .A(n3), .B(N456), .Z(n320) );
  NAND U478 ( .A(n322), .B(n323), .Z(z3[191]) );
  NANDN U479 ( .A(N262), .B(z2[191]), .Z(n323) );
  NANDN U480 ( .A(n3), .B(N455), .Z(n322) );
  NAND U481 ( .A(n324), .B(n325), .Z(z3[190]) );
  NANDN U482 ( .A(N262), .B(z2[190]), .Z(n325) );
  NANDN U483 ( .A(n3), .B(N454), .Z(n324) );
  NAND U484 ( .A(n326), .B(n327), .Z(z3[18]) );
  NANDN U485 ( .A(N262), .B(z2[18]), .Z(n327) );
  NANDN U486 ( .A(n3), .B(N282), .Z(n326) );
  NAND U487 ( .A(n328), .B(n329), .Z(z3[189]) );
  NANDN U488 ( .A(N262), .B(z2[189]), .Z(n329) );
  NANDN U489 ( .A(n3), .B(N453), .Z(n328) );
  NAND U490 ( .A(n330), .B(n331), .Z(z3[188]) );
  NANDN U491 ( .A(N262), .B(z2[188]), .Z(n331) );
  NANDN U492 ( .A(n3), .B(N452), .Z(n330) );
  NAND U493 ( .A(n332), .B(n333), .Z(z3[187]) );
  NANDN U494 ( .A(N262), .B(z2[187]), .Z(n333) );
  NANDN U495 ( .A(n3), .B(N451), .Z(n332) );
  NAND U496 ( .A(n334), .B(n335), .Z(z3[186]) );
  NANDN U497 ( .A(N262), .B(z2[186]), .Z(n335) );
  NANDN U498 ( .A(n3), .B(N450), .Z(n334) );
  NAND U499 ( .A(n336), .B(n337), .Z(z3[185]) );
  NANDN U500 ( .A(N262), .B(z2[185]), .Z(n337) );
  NANDN U501 ( .A(n3), .B(N449), .Z(n336) );
  NAND U502 ( .A(n338), .B(n339), .Z(z3[184]) );
  NANDN U503 ( .A(N262), .B(z2[184]), .Z(n339) );
  NANDN U504 ( .A(n3), .B(N448), .Z(n338) );
  NAND U505 ( .A(n340), .B(n341), .Z(z3[183]) );
  NANDN U506 ( .A(N262), .B(z2[183]), .Z(n341) );
  NANDN U507 ( .A(n3), .B(N447), .Z(n340) );
  NAND U508 ( .A(n342), .B(n343), .Z(z3[182]) );
  NANDN U509 ( .A(N262), .B(z2[182]), .Z(n343) );
  NANDN U510 ( .A(n3), .B(N446), .Z(n342) );
  NAND U511 ( .A(n344), .B(n345), .Z(z3[181]) );
  NANDN U512 ( .A(N262), .B(z2[181]), .Z(n345) );
  NANDN U513 ( .A(n3), .B(N445), .Z(n344) );
  NAND U514 ( .A(n346), .B(n347), .Z(z3[180]) );
  NANDN U515 ( .A(N262), .B(z2[180]), .Z(n347) );
  NANDN U516 ( .A(n3), .B(N444), .Z(n346) );
  NAND U517 ( .A(n348), .B(n349), .Z(z3[17]) );
  NANDN U518 ( .A(N262), .B(z2[17]), .Z(n349) );
  NANDN U519 ( .A(n3), .B(N281), .Z(n348) );
  NAND U520 ( .A(n350), .B(n351), .Z(z3[179]) );
  NANDN U521 ( .A(N262), .B(z2[179]), .Z(n351) );
  NANDN U522 ( .A(n3), .B(N443), .Z(n350) );
  NAND U523 ( .A(n352), .B(n353), .Z(z3[178]) );
  NANDN U524 ( .A(N262), .B(z2[178]), .Z(n353) );
  NANDN U525 ( .A(n3), .B(N442), .Z(n352) );
  NAND U526 ( .A(n354), .B(n355), .Z(z3[177]) );
  NANDN U527 ( .A(N262), .B(z2[177]), .Z(n355) );
  NANDN U528 ( .A(n3), .B(N441), .Z(n354) );
  NAND U529 ( .A(n356), .B(n357), .Z(z3[176]) );
  NANDN U530 ( .A(N262), .B(z2[176]), .Z(n357) );
  NANDN U531 ( .A(n3), .B(N440), .Z(n356) );
  NAND U532 ( .A(n358), .B(n359), .Z(z3[175]) );
  NANDN U533 ( .A(N262), .B(z2[175]), .Z(n359) );
  NANDN U534 ( .A(n3), .B(N439), .Z(n358) );
  NAND U535 ( .A(n360), .B(n361), .Z(z3[174]) );
  NANDN U536 ( .A(N262), .B(z2[174]), .Z(n361) );
  NANDN U537 ( .A(n3), .B(N438), .Z(n360) );
  NAND U538 ( .A(n362), .B(n363), .Z(z3[173]) );
  NANDN U539 ( .A(N262), .B(z2[173]), .Z(n363) );
  NANDN U540 ( .A(n3), .B(N437), .Z(n362) );
  NAND U541 ( .A(n364), .B(n365), .Z(z3[172]) );
  NANDN U542 ( .A(N262), .B(z2[172]), .Z(n365) );
  NANDN U543 ( .A(n3), .B(N436), .Z(n364) );
  NAND U544 ( .A(n366), .B(n367), .Z(z3[171]) );
  NANDN U545 ( .A(N262), .B(z2[171]), .Z(n367) );
  NANDN U546 ( .A(n3), .B(N435), .Z(n366) );
  NAND U547 ( .A(n368), .B(n369), .Z(z3[170]) );
  NANDN U548 ( .A(N262), .B(z2[170]), .Z(n369) );
  NANDN U549 ( .A(n3), .B(N434), .Z(n368) );
  NAND U550 ( .A(n370), .B(n371), .Z(z3[16]) );
  NANDN U551 ( .A(N262), .B(z2[16]), .Z(n371) );
  NANDN U552 ( .A(n3), .B(N280), .Z(n370) );
  NAND U553 ( .A(n372), .B(n373), .Z(z3[169]) );
  NANDN U554 ( .A(N262), .B(z2[169]), .Z(n373) );
  NANDN U555 ( .A(n3), .B(N433), .Z(n372) );
  NAND U556 ( .A(n374), .B(n375), .Z(z3[168]) );
  NANDN U557 ( .A(N262), .B(z2[168]), .Z(n375) );
  NANDN U558 ( .A(n3), .B(N432), .Z(n374) );
  NAND U559 ( .A(n376), .B(n377), .Z(z3[167]) );
  NANDN U560 ( .A(N262), .B(z2[167]), .Z(n377) );
  NANDN U561 ( .A(n3), .B(N431), .Z(n376) );
  NAND U562 ( .A(n378), .B(n379), .Z(z3[166]) );
  NANDN U563 ( .A(N262), .B(z2[166]), .Z(n379) );
  NANDN U564 ( .A(n3), .B(N430), .Z(n378) );
  NAND U565 ( .A(n380), .B(n381), .Z(z3[165]) );
  NANDN U566 ( .A(N262), .B(z2[165]), .Z(n381) );
  NANDN U567 ( .A(n3), .B(N429), .Z(n380) );
  NAND U568 ( .A(n382), .B(n383), .Z(z3[164]) );
  NANDN U569 ( .A(N262), .B(z2[164]), .Z(n383) );
  NANDN U570 ( .A(n3), .B(N428), .Z(n382) );
  NAND U571 ( .A(n384), .B(n385), .Z(z3[163]) );
  NANDN U572 ( .A(N262), .B(z2[163]), .Z(n385) );
  NANDN U573 ( .A(n3), .B(N427), .Z(n384) );
  NAND U574 ( .A(n386), .B(n387), .Z(z3[162]) );
  NANDN U575 ( .A(N262), .B(z2[162]), .Z(n387) );
  NANDN U576 ( .A(n3), .B(N426), .Z(n386) );
  NAND U577 ( .A(n388), .B(n389), .Z(z3[161]) );
  NANDN U578 ( .A(N262), .B(z2[161]), .Z(n389) );
  NANDN U579 ( .A(n3), .B(N425), .Z(n388) );
  NAND U580 ( .A(n390), .B(n391), .Z(z3[160]) );
  NANDN U581 ( .A(N262), .B(z2[160]), .Z(n391) );
  NANDN U582 ( .A(n3), .B(N424), .Z(n390) );
  NAND U583 ( .A(n392), .B(n393), .Z(z3[15]) );
  NANDN U584 ( .A(N262), .B(z2[15]), .Z(n393) );
  NANDN U585 ( .A(n3), .B(N279), .Z(n392) );
  NAND U586 ( .A(n394), .B(n395), .Z(z3[159]) );
  NANDN U587 ( .A(N262), .B(z2[159]), .Z(n395) );
  NANDN U588 ( .A(n3), .B(N423), .Z(n394) );
  NAND U589 ( .A(n396), .B(n397), .Z(z3[158]) );
  NANDN U590 ( .A(N262), .B(z2[158]), .Z(n397) );
  NANDN U591 ( .A(n3), .B(N422), .Z(n396) );
  NAND U592 ( .A(n398), .B(n399), .Z(z3[157]) );
  NANDN U593 ( .A(N262), .B(z2[157]), .Z(n399) );
  NANDN U594 ( .A(n3), .B(N421), .Z(n398) );
  NAND U595 ( .A(n400), .B(n401), .Z(z3[156]) );
  NANDN U596 ( .A(N262), .B(z2[156]), .Z(n401) );
  NANDN U597 ( .A(n3), .B(N420), .Z(n400) );
  NAND U598 ( .A(n402), .B(n403), .Z(z3[155]) );
  NANDN U599 ( .A(N262), .B(z2[155]), .Z(n403) );
  NANDN U600 ( .A(n3), .B(N419), .Z(n402) );
  NAND U601 ( .A(n404), .B(n405), .Z(z3[154]) );
  NANDN U602 ( .A(N262), .B(z2[154]), .Z(n405) );
  NANDN U603 ( .A(n3), .B(N418), .Z(n404) );
  NAND U604 ( .A(n406), .B(n407), .Z(z3[153]) );
  NANDN U605 ( .A(N262), .B(z2[153]), .Z(n407) );
  NANDN U606 ( .A(n3), .B(N417), .Z(n406) );
  NAND U607 ( .A(n408), .B(n409), .Z(z3[152]) );
  NANDN U608 ( .A(N262), .B(z2[152]), .Z(n409) );
  NANDN U609 ( .A(n3), .B(N416), .Z(n408) );
  NAND U610 ( .A(n410), .B(n411), .Z(z3[151]) );
  NANDN U611 ( .A(N262), .B(z2[151]), .Z(n411) );
  NANDN U612 ( .A(n3), .B(N415), .Z(n410) );
  NAND U613 ( .A(n412), .B(n413), .Z(z3[150]) );
  NANDN U614 ( .A(N262), .B(z2[150]), .Z(n413) );
  NANDN U615 ( .A(n3), .B(N414), .Z(n412) );
  NAND U616 ( .A(n414), .B(n415), .Z(z3[14]) );
  NANDN U617 ( .A(N262), .B(z2[14]), .Z(n415) );
  NANDN U618 ( .A(n3), .B(N278), .Z(n414) );
  NAND U619 ( .A(n416), .B(n417), .Z(z3[149]) );
  NANDN U620 ( .A(N262), .B(z2[149]), .Z(n417) );
  NANDN U621 ( .A(n3), .B(N413), .Z(n416) );
  NAND U622 ( .A(n418), .B(n419), .Z(z3[148]) );
  NANDN U623 ( .A(N262), .B(z2[148]), .Z(n419) );
  NANDN U624 ( .A(n3), .B(N412), .Z(n418) );
  NAND U625 ( .A(n420), .B(n421), .Z(z3[147]) );
  NANDN U626 ( .A(N262), .B(z2[147]), .Z(n421) );
  NANDN U627 ( .A(n3), .B(N411), .Z(n420) );
  NAND U628 ( .A(n422), .B(n423), .Z(z3[146]) );
  NANDN U629 ( .A(N262), .B(z2[146]), .Z(n423) );
  NANDN U630 ( .A(n3), .B(N410), .Z(n422) );
  NAND U631 ( .A(n424), .B(n425), .Z(z3[145]) );
  NANDN U632 ( .A(N262), .B(z2[145]), .Z(n425) );
  NANDN U633 ( .A(n3), .B(N409), .Z(n424) );
  NAND U634 ( .A(n426), .B(n427), .Z(z3[144]) );
  NANDN U635 ( .A(N262), .B(z2[144]), .Z(n427) );
  NANDN U636 ( .A(n3), .B(N408), .Z(n426) );
  NAND U637 ( .A(n428), .B(n429), .Z(z3[143]) );
  NANDN U638 ( .A(N262), .B(z2[143]), .Z(n429) );
  NANDN U639 ( .A(n3), .B(N407), .Z(n428) );
  NAND U640 ( .A(n430), .B(n431), .Z(z3[142]) );
  NANDN U641 ( .A(N262), .B(z2[142]), .Z(n431) );
  NANDN U642 ( .A(n3), .B(N406), .Z(n430) );
  NAND U643 ( .A(n432), .B(n433), .Z(z3[141]) );
  NANDN U644 ( .A(N262), .B(z2[141]), .Z(n433) );
  NANDN U645 ( .A(n3), .B(N405), .Z(n432) );
  NAND U646 ( .A(n434), .B(n435), .Z(z3[140]) );
  NANDN U647 ( .A(N262), .B(z2[140]), .Z(n435) );
  NANDN U648 ( .A(n3), .B(N404), .Z(n434) );
  NAND U649 ( .A(n436), .B(n437), .Z(z3[13]) );
  NANDN U650 ( .A(N262), .B(z2[13]), .Z(n437) );
  NANDN U651 ( .A(n3), .B(N277), .Z(n436) );
  NAND U652 ( .A(n438), .B(n439), .Z(z3[139]) );
  NANDN U653 ( .A(N262), .B(z2[139]), .Z(n439) );
  NANDN U654 ( .A(n3), .B(N403), .Z(n438) );
  NAND U655 ( .A(n440), .B(n441), .Z(z3[138]) );
  NANDN U656 ( .A(N262), .B(z2[138]), .Z(n441) );
  NANDN U657 ( .A(n3), .B(N402), .Z(n440) );
  NAND U658 ( .A(n442), .B(n443), .Z(z3[137]) );
  NANDN U659 ( .A(N262), .B(z2[137]), .Z(n443) );
  NANDN U660 ( .A(n3), .B(N401), .Z(n442) );
  NAND U661 ( .A(n444), .B(n445), .Z(z3[136]) );
  NANDN U662 ( .A(N262), .B(z2[136]), .Z(n445) );
  NANDN U663 ( .A(n3), .B(N400), .Z(n444) );
  NAND U664 ( .A(n446), .B(n447), .Z(z3[135]) );
  NANDN U665 ( .A(N262), .B(z2[135]), .Z(n447) );
  NANDN U666 ( .A(n3), .B(N399), .Z(n446) );
  NAND U667 ( .A(n448), .B(n449), .Z(z3[134]) );
  NANDN U668 ( .A(N262), .B(z2[134]), .Z(n449) );
  NANDN U669 ( .A(n3), .B(N398), .Z(n448) );
  NAND U670 ( .A(n450), .B(n451), .Z(z3[133]) );
  NANDN U671 ( .A(N262), .B(z2[133]), .Z(n451) );
  NANDN U672 ( .A(n3), .B(N397), .Z(n450) );
  NAND U673 ( .A(n452), .B(n453), .Z(z3[132]) );
  NANDN U674 ( .A(N262), .B(z2[132]), .Z(n453) );
  NANDN U675 ( .A(n3), .B(N396), .Z(n452) );
  NAND U676 ( .A(n454), .B(n455), .Z(z3[131]) );
  NANDN U677 ( .A(N262), .B(z2[131]), .Z(n455) );
  NANDN U678 ( .A(n3), .B(N395), .Z(n454) );
  NAND U679 ( .A(n456), .B(n457), .Z(z3[130]) );
  NANDN U680 ( .A(N262), .B(z2[130]), .Z(n457) );
  NANDN U681 ( .A(n3), .B(N394), .Z(n456) );
  NAND U682 ( .A(n458), .B(n459), .Z(z3[12]) );
  NANDN U683 ( .A(N262), .B(z2[12]), .Z(n459) );
  NANDN U684 ( .A(n3), .B(N276), .Z(n458) );
  NAND U685 ( .A(n460), .B(n461), .Z(z3[129]) );
  NANDN U686 ( .A(N262), .B(z2[129]), .Z(n461) );
  NANDN U687 ( .A(n3), .B(N393), .Z(n460) );
  NAND U688 ( .A(n462), .B(n463), .Z(z3[128]) );
  NANDN U689 ( .A(N262), .B(z2[128]), .Z(n463) );
  NANDN U690 ( .A(n3), .B(N392), .Z(n462) );
  NAND U691 ( .A(n464), .B(n465), .Z(z3[127]) );
  NANDN U692 ( .A(N262), .B(z2[127]), .Z(n465) );
  NANDN U693 ( .A(n3), .B(N391), .Z(n464) );
  NAND U694 ( .A(n466), .B(n467), .Z(z3[126]) );
  NANDN U695 ( .A(N262), .B(z2[126]), .Z(n467) );
  NANDN U696 ( .A(n3), .B(N390), .Z(n466) );
  NAND U697 ( .A(n468), .B(n469), .Z(z3[125]) );
  NANDN U698 ( .A(N262), .B(z2[125]), .Z(n469) );
  NANDN U699 ( .A(n3), .B(N389), .Z(n468) );
  NAND U700 ( .A(n470), .B(n471), .Z(z3[124]) );
  NANDN U701 ( .A(N262), .B(z2[124]), .Z(n471) );
  NANDN U702 ( .A(n3), .B(N388), .Z(n470) );
  NAND U703 ( .A(n472), .B(n473), .Z(z3[123]) );
  NANDN U704 ( .A(N262), .B(z2[123]), .Z(n473) );
  NANDN U705 ( .A(n3), .B(N387), .Z(n472) );
  NAND U706 ( .A(n474), .B(n475), .Z(z3[122]) );
  NANDN U707 ( .A(N262), .B(z2[122]), .Z(n475) );
  NANDN U708 ( .A(n3), .B(N386), .Z(n474) );
  NAND U709 ( .A(n476), .B(n477), .Z(z3[121]) );
  NANDN U710 ( .A(N262), .B(z2[121]), .Z(n477) );
  NANDN U711 ( .A(n3), .B(N385), .Z(n476) );
  NAND U712 ( .A(n478), .B(n479), .Z(z3[120]) );
  NANDN U713 ( .A(N262), .B(z2[120]), .Z(n479) );
  NANDN U714 ( .A(n3), .B(N384), .Z(n478) );
  NAND U715 ( .A(n480), .B(n481), .Z(z3[11]) );
  NANDN U716 ( .A(N262), .B(z2[11]), .Z(n481) );
  NANDN U717 ( .A(n3), .B(N275), .Z(n480) );
  NAND U718 ( .A(n482), .B(n483), .Z(z3[119]) );
  NANDN U719 ( .A(N262), .B(z2[119]), .Z(n483) );
  NANDN U720 ( .A(n3), .B(N383), .Z(n482) );
  NAND U721 ( .A(n484), .B(n485), .Z(z3[118]) );
  NANDN U722 ( .A(N262), .B(z2[118]), .Z(n485) );
  NANDN U723 ( .A(n3), .B(N382), .Z(n484) );
  NAND U724 ( .A(n486), .B(n487), .Z(z3[117]) );
  NANDN U725 ( .A(N262), .B(z2[117]), .Z(n487) );
  NANDN U726 ( .A(n3), .B(N381), .Z(n486) );
  NAND U727 ( .A(n488), .B(n489), .Z(z3[116]) );
  NANDN U728 ( .A(N262), .B(z2[116]), .Z(n489) );
  NANDN U729 ( .A(n3), .B(N380), .Z(n488) );
  NAND U730 ( .A(n490), .B(n491), .Z(z3[115]) );
  NANDN U731 ( .A(N262), .B(z2[115]), .Z(n491) );
  NANDN U732 ( .A(n3), .B(N379), .Z(n490) );
  NAND U733 ( .A(n492), .B(n493), .Z(z3[114]) );
  NANDN U734 ( .A(N262), .B(z2[114]), .Z(n493) );
  NANDN U735 ( .A(n3), .B(N378), .Z(n492) );
  NAND U736 ( .A(n494), .B(n495), .Z(z3[113]) );
  NANDN U737 ( .A(N262), .B(z2[113]), .Z(n495) );
  NANDN U738 ( .A(n3), .B(N377), .Z(n494) );
  NAND U739 ( .A(n496), .B(n497), .Z(z3[112]) );
  NANDN U740 ( .A(N262), .B(z2[112]), .Z(n497) );
  NANDN U741 ( .A(n3), .B(N376), .Z(n496) );
  NAND U742 ( .A(n498), .B(n499), .Z(z3[111]) );
  NANDN U743 ( .A(N262), .B(z2[111]), .Z(n499) );
  NANDN U744 ( .A(n3), .B(N375), .Z(n498) );
  NAND U745 ( .A(n500), .B(n501), .Z(z3[110]) );
  NANDN U746 ( .A(N262), .B(z2[110]), .Z(n501) );
  NANDN U747 ( .A(n3), .B(N374), .Z(n500) );
  NAND U748 ( .A(n502), .B(n503), .Z(z3[10]) );
  NANDN U749 ( .A(N262), .B(z2[10]), .Z(n503) );
  NANDN U750 ( .A(n3), .B(N274), .Z(n502) );
  NAND U751 ( .A(n504), .B(n505), .Z(z3[109]) );
  NANDN U752 ( .A(N262), .B(z2[109]), .Z(n505) );
  NANDN U753 ( .A(n3), .B(N373), .Z(n504) );
  NAND U754 ( .A(n506), .B(n507), .Z(z3[108]) );
  NANDN U755 ( .A(N262), .B(z2[108]), .Z(n507) );
  NANDN U756 ( .A(n3), .B(N372), .Z(n506) );
  NAND U757 ( .A(n508), .B(n509), .Z(z3[107]) );
  NANDN U758 ( .A(N262), .B(z2[107]), .Z(n509) );
  NANDN U759 ( .A(n3), .B(N371), .Z(n508) );
  NAND U760 ( .A(n510), .B(n511), .Z(z3[106]) );
  NANDN U761 ( .A(N262), .B(z2[106]), .Z(n511) );
  NANDN U762 ( .A(n3), .B(N370), .Z(n510) );
  NAND U763 ( .A(n512), .B(n513), .Z(z3[105]) );
  NANDN U764 ( .A(N262), .B(z2[105]), .Z(n513) );
  NANDN U765 ( .A(n3), .B(N369), .Z(n512) );
  NAND U766 ( .A(n514), .B(n515), .Z(z3[104]) );
  NANDN U767 ( .A(N262), .B(z2[104]), .Z(n515) );
  NANDN U768 ( .A(n3), .B(N368), .Z(n514) );
  NAND U769 ( .A(n516), .B(n517), .Z(z3[103]) );
  NANDN U770 ( .A(N262), .B(z2[103]), .Z(n517) );
  NANDN U771 ( .A(n3), .B(N367), .Z(n516) );
  NAND U772 ( .A(n518), .B(n519), .Z(z3[102]) );
  NANDN U773 ( .A(N262), .B(z2[102]), .Z(n519) );
  NANDN U774 ( .A(n3), .B(N366), .Z(n518) );
  NAND U775 ( .A(n520), .B(n521), .Z(z3[101]) );
  NANDN U776 ( .A(N262), .B(z2[101]), .Z(n521) );
  NANDN U777 ( .A(n3), .B(N365), .Z(n520) );
  NAND U778 ( .A(n522), .B(n523), .Z(z3[100]) );
  NANDN U779 ( .A(N262), .B(z2[100]), .Z(n523) );
  NANDN U780 ( .A(n3), .B(N364), .Z(n522) );
  NAND U781 ( .A(n524), .B(n525), .Z(z3[0]) );
  NANDN U782 ( .A(N262), .B(z2[0]), .Z(n525) );
  NANDN U783 ( .A(n3), .B(N264), .Z(n524) );
  IV U784 ( .A(N262), .Z(n3) );
  NAND U785 ( .A(n526), .B(n527), .Z(z2[9]) );
  NANDN U786 ( .A(xregN_1), .B(zin[8]), .Z(n527) );
  NAND U787 ( .A(N13), .B(xregN_1), .Z(n526) );
  NAND U788 ( .A(n528), .B(n529), .Z(z2[99]) );
  NANDN U789 ( .A(xregN_1), .B(zin[98]), .Z(n529) );
  NAND U790 ( .A(N103), .B(xregN_1), .Z(n528) );
  NAND U791 ( .A(n530), .B(n531), .Z(z2[98]) );
  NANDN U792 ( .A(xregN_1), .B(zin[97]), .Z(n531) );
  NAND U793 ( .A(N102), .B(xregN_1), .Z(n530) );
  NAND U794 ( .A(n532), .B(n533), .Z(z2[97]) );
  NANDN U795 ( .A(xregN_1), .B(zin[96]), .Z(n533) );
  NAND U796 ( .A(N101), .B(xregN_1), .Z(n532) );
  NAND U797 ( .A(n534), .B(n535), .Z(z2[96]) );
  NANDN U798 ( .A(xregN_1), .B(zin[95]), .Z(n535) );
  NAND U799 ( .A(N100), .B(xregN_1), .Z(n534) );
  NAND U800 ( .A(n536), .B(n537), .Z(z2[95]) );
  NANDN U801 ( .A(xregN_1), .B(zin[94]), .Z(n537) );
  NAND U802 ( .A(N99), .B(xregN_1), .Z(n536) );
  NAND U803 ( .A(n538), .B(n539), .Z(z2[94]) );
  NANDN U804 ( .A(xregN_1), .B(zin[93]), .Z(n539) );
  NAND U805 ( .A(N98), .B(xregN_1), .Z(n538) );
  NAND U806 ( .A(n540), .B(n541), .Z(z2[93]) );
  NANDN U807 ( .A(xregN_1), .B(zin[92]), .Z(n541) );
  NAND U808 ( .A(N97), .B(xregN_1), .Z(n540) );
  NAND U809 ( .A(n542), .B(n543), .Z(z2[92]) );
  NANDN U810 ( .A(xregN_1), .B(zin[91]), .Z(n543) );
  NAND U811 ( .A(N96), .B(xregN_1), .Z(n542) );
  NAND U812 ( .A(n544), .B(n545), .Z(z2[91]) );
  NANDN U813 ( .A(xregN_1), .B(zin[90]), .Z(n545) );
  NAND U814 ( .A(N95), .B(xregN_1), .Z(n544) );
  NAND U815 ( .A(n546), .B(n547), .Z(z2[90]) );
  NANDN U816 ( .A(xregN_1), .B(zin[89]), .Z(n547) );
  NAND U817 ( .A(N94), .B(xregN_1), .Z(n546) );
  NAND U818 ( .A(n548), .B(n549), .Z(z2[8]) );
  NANDN U819 ( .A(xregN_1), .B(zin[7]), .Z(n549) );
  NAND U820 ( .A(N12), .B(xregN_1), .Z(n548) );
  NAND U821 ( .A(n550), .B(n551), .Z(z2[89]) );
  NANDN U822 ( .A(xregN_1), .B(zin[88]), .Z(n551) );
  NAND U823 ( .A(N93), .B(xregN_1), .Z(n550) );
  NAND U824 ( .A(n552), .B(n553), .Z(z2[88]) );
  NANDN U825 ( .A(xregN_1), .B(zin[87]), .Z(n553) );
  NAND U826 ( .A(N92), .B(xregN_1), .Z(n552) );
  NAND U827 ( .A(n554), .B(n555), .Z(z2[87]) );
  NANDN U828 ( .A(xregN_1), .B(zin[86]), .Z(n555) );
  NAND U829 ( .A(N91), .B(xregN_1), .Z(n554) );
  NAND U830 ( .A(n556), .B(n557), .Z(z2[86]) );
  NANDN U831 ( .A(xregN_1), .B(zin[85]), .Z(n557) );
  NAND U832 ( .A(N90), .B(xregN_1), .Z(n556) );
  NAND U833 ( .A(n558), .B(n559), .Z(z2[85]) );
  NANDN U834 ( .A(xregN_1), .B(zin[84]), .Z(n559) );
  NAND U835 ( .A(N89), .B(xregN_1), .Z(n558) );
  NAND U836 ( .A(n560), .B(n561), .Z(z2[84]) );
  NANDN U837 ( .A(xregN_1), .B(zin[83]), .Z(n561) );
  NAND U838 ( .A(N88), .B(xregN_1), .Z(n560) );
  NAND U839 ( .A(n562), .B(n563), .Z(z2[83]) );
  NANDN U840 ( .A(xregN_1), .B(zin[82]), .Z(n563) );
  NAND U841 ( .A(N87), .B(xregN_1), .Z(n562) );
  NAND U842 ( .A(n564), .B(n565), .Z(z2[82]) );
  NANDN U843 ( .A(xregN_1), .B(zin[81]), .Z(n565) );
  NAND U844 ( .A(N86), .B(xregN_1), .Z(n564) );
  NAND U845 ( .A(n566), .B(n567), .Z(z2[81]) );
  NANDN U846 ( .A(xregN_1), .B(zin[80]), .Z(n567) );
  NAND U847 ( .A(N85), .B(xregN_1), .Z(n566) );
  NAND U848 ( .A(n568), .B(n569), .Z(z2[80]) );
  NANDN U849 ( .A(xregN_1), .B(zin[79]), .Z(n569) );
  NAND U850 ( .A(N84), .B(xregN_1), .Z(n568) );
  NAND U851 ( .A(n570), .B(n571), .Z(z2[7]) );
  NANDN U852 ( .A(xregN_1), .B(zin[6]), .Z(n571) );
  NAND U853 ( .A(N11), .B(xregN_1), .Z(n570) );
  NAND U854 ( .A(n572), .B(n573), .Z(z2[79]) );
  NANDN U855 ( .A(xregN_1), .B(zin[78]), .Z(n573) );
  NAND U856 ( .A(N83), .B(xregN_1), .Z(n572) );
  NAND U857 ( .A(n574), .B(n575), .Z(z2[78]) );
  NANDN U858 ( .A(xregN_1), .B(zin[77]), .Z(n575) );
  NAND U859 ( .A(N82), .B(xregN_1), .Z(n574) );
  NAND U860 ( .A(n576), .B(n577), .Z(z2[77]) );
  NANDN U861 ( .A(xregN_1), .B(zin[76]), .Z(n577) );
  NAND U862 ( .A(N81), .B(xregN_1), .Z(n576) );
  NAND U863 ( .A(n578), .B(n579), .Z(z2[76]) );
  NANDN U864 ( .A(xregN_1), .B(zin[75]), .Z(n579) );
  NAND U865 ( .A(N80), .B(xregN_1), .Z(n578) );
  NAND U866 ( .A(n580), .B(n581), .Z(z2[75]) );
  NANDN U867 ( .A(xregN_1), .B(zin[74]), .Z(n581) );
  NAND U868 ( .A(N79), .B(xregN_1), .Z(n580) );
  NAND U869 ( .A(n582), .B(n583), .Z(z2[74]) );
  NANDN U870 ( .A(xregN_1), .B(zin[73]), .Z(n583) );
  NAND U871 ( .A(N78), .B(xregN_1), .Z(n582) );
  NAND U872 ( .A(n584), .B(n585), .Z(z2[73]) );
  NANDN U873 ( .A(xregN_1), .B(zin[72]), .Z(n585) );
  NAND U874 ( .A(N77), .B(xregN_1), .Z(n584) );
  NAND U875 ( .A(n586), .B(n587), .Z(z2[72]) );
  NANDN U876 ( .A(xregN_1), .B(zin[71]), .Z(n587) );
  NAND U877 ( .A(N76), .B(xregN_1), .Z(n586) );
  NAND U878 ( .A(n588), .B(n589), .Z(z2[71]) );
  NANDN U879 ( .A(xregN_1), .B(zin[70]), .Z(n589) );
  NAND U880 ( .A(N75), .B(xregN_1), .Z(n588) );
  NAND U881 ( .A(n590), .B(n591), .Z(z2[70]) );
  NANDN U882 ( .A(xregN_1), .B(zin[69]), .Z(n591) );
  NAND U883 ( .A(N74), .B(xregN_1), .Z(n590) );
  NAND U884 ( .A(n592), .B(n593), .Z(z2[6]) );
  NANDN U885 ( .A(xregN_1), .B(zin[5]), .Z(n593) );
  NAND U886 ( .A(N10), .B(xregN_1), .Z(n592) );
  NAND U887 ( .A(n594), .B(n595), .Z(z2[69]) );
  NANDN U888 ( .A(xregN_1), .B(zin[68]), .Z(n595) );
  NAND U889 ( .A(N73), .B(xregN_1), .Z(n594) );
  NAND U890 ( .A(n596), .B(n597), .Z(z2[68]) );
  NANDN U891 ( .A(xregN_1), .B(zin[67]), .Z(n597) );
  NAND U892 ( .A(N72), .B(xregN_1), .Z(n596) );
  NAND U893 ( .A(n598), .B(n599), .Z(z2[67]) );
  NANDN U894 ( .A(xregN_1), .B(zin[66]), .Z(n599) );
  NAND U895 ( .A(N71), .B(xregN_1), .Z(n598) );
  NAND U896 ( .A(n600), .B(n601), .Z(z2[66]) );
  NANDN U897 ( .A(xregN_1), .B(zin[65]), .Z(n601) );
  NAND U898 ( .A(N70), .B(xregN_1), .Z(n600) );
  NAND U899 ( .A(n602), .B(n603), .Z(z2[65]) );
  NANDN U900 ( .A(xregN_1), .B(zin[64]), .Z(n603) );
  NAND U901 ( .A(N69), .B(xregN_1), .Z(n602) );
  NAND U902 ( .A(n604), .B(n605), .Z(z2[64]) );
  NANDN U903 ( .A(xregN_1), .B(zin[63]), .Z(n605) );
  NAND U904 ( .A(N68), .B(xregN_1), .Z(n604) );
  NAND U905 ( .A(n606), .B(n607), .Z(z2[63]) );
  NANDN U906 ( .A(xregN_1), .B(zin[62]), .Z(n607) );
  NAND U907 ( .A(N67), .B(xregN_1), .Z(n606) );
  NAND U908 ( .A(n608), .B(n609), .Z(z2[62]) );
  NANDN U909 ( .A(xregN_1), .B(zin[61]), .Z(n609) );
  NAND U910 ( .A(N66), .B(xregN_1), .Z(n608) );
  NAND U911 ( .A(n610), .B(n611), .Z(z2[61]) );
  NANDN U912 ( .A(xregN_1), .B(zin[60]), .Z(n611) );
  NAND U913 ( .A(N65), .B(xregN_1), .Z(n610) );
  NAND U914 ( .A(n612), .B(n613), .Z(z2[60]) );
  NANDN U915 ( .A(xregN_1), .B(zin[59]), .Z(n613) );
  NAND U916 ( .A(N64), .B(xregN_1), .Z(n612) );
  NAND U917 ( .A(n614), .B(n615), .Z(z2[5]) );
  NANDN U918 ( .A(xregN_1), .B(zin[4]), .Z(n615) );
  NAND U919 ( .A(N9), .B(xregN_1), .Z(n614) );
  NAND U920 ( .A(n616), .B(n617), .Z(z2[59]) );
  NANDN U921 ( .A(xregN_1), .B(zin[58]), .Z(n617) );
  NAND U922 ( .A(N63), .B(xregN_1), .Z(n616) );
  NAND U923 ( .A(n618), .B(n619), .Z(z2[58]) );
  NANDN U924 ( .A(xregN_1), .B(zin[57]), .Z(n619) );
  NAND U925 ( .A(N62), .B(xregN_1), .Z(n618) );
  NAND U926 ( .A(n620), .B(n621), .Z(z2[57]) );
  NANDN U927 ( .A(xregN_1), .B(zin[56]), .Z(n621) );
  NAND U928 ( .A(N61), .B(xregN_1), .Z(n620) );
  NAND U929 ( .A(n622), .B(n623), .Z(z2[56]) );
  NANDN U930 ( .A(xregN_1), .B(zin[55]), .Z(n623) );
  NAND U931 ( .A(N60), .B(xregN_1), .Z(n622) );
  NAND U932 ( .A(n624), .B(n625), .Z(z2[55]) );
  NANDN U933 ( .A(xregN_1), .B(zin[54]), .Z(n625) );
  NAND U934 ( .A(N59), .B(xregN_1), .Z(n624) );
  NAND U935 ( .A(n626), .B(n627), .Z(z2[54]) );
  NANDN U936 ( .A(xregN_1), .B(zin[53]), .Z(n627) );
  NAND U937 ( .A(N58), .B(xregN_1), .Z(n626) );
  NAND U938 ( .A(n628), .B(n629), .Z(z2[53]) );
  NANDN U939 ( .A(xregN_1), .B(zin[52]), .Z(n629) );
  NAND U940 ( .A(N57), .B(xregN_1), .Z(n628) );
  NAND U941 ( .A(n630), .B(n631), .Z(z2[52]) );
  NANDN U942 ( .A(xregN_1), .B(zin[51]), .Z(n631) );
  NAND U943 ( .A(N56), .B(xregN_1), .Z(n630) );
  NAND U944 ( .A(n632), .B(n633), .Z(z2[51]) );
  NANDN U945 ( .A(xregN_1), .B(zin[50]), .Z(n633) );
  NAND U946 ( .A(N55), .B(xregN_1), .Z(n632) );
  NAND U947 ( .A(n634), .B(n635), .Z(z2[50]) );
  NANDN U948 ( .A(xregN_1), .B(zin[49]), .Z(n635) );
  NAND U949 ( .A(N54), .B(xregN_1), .Z(n634) );
  NAND U950 ( .A(n636), .B(n637), .Z(z2[4]) );
  NANDN U951 ( .A(xregN_1), .B(zin[3]), .Z(n637) );
  NAND U952 ( .A(N8), .B(xregN_1), .Z(n636) );
  NAND U953 ( .A(n638), .B(n639), .Z(z2[49]) );
  NANDN U954 ( .A(xregN_1), .B(zin[48]), .Z(n639) );
  NAND U955 ( .A(N53), .B(xregN_1), .Z(n638) );
  NAND U956 ( .A(n640), .B(n641), .Z(z2[48]) );
  NANDN U957 ( .A(xregN_1), .B(zin[47]), .Z(n641) );
  NAND U958 ( .A(N52), .B(xregN_1), .Z(n640) );
  NAND U959 ( .A(n642), .B(n643), .Z(z2[47]) );
  NANDN U960 ( .A(xregN_1), .B(zin[46]), .Z(n643) );
  NAND U961 ( .A(N51), .B(xregN_1), .Z(n642) );
  NAND U962 ( .A(n644), .B(n645), .Z(z2[46]) );
  NANDN U963 ( .A(xregN_1), .B(zin[45]), .Z(n645) );
  NAND U964 ( .A(N50), .B(xregN_1), .Z(n644) );
  NAND U965 ( .A(n646), .B(n647), .Z(z2[45]) );
  NANDN U966 ( .A(xregN_1), .B(zin[44]), .Z(n647) );
  NAND U967 ( .A(N49), .B(xregN_1), .Z(n646) );
  NAND U968 ( .A(n648), .B(n649), .Z(z2[44]) );
  NANDN U969 ( .A(xregN_1), .B(zin[43]), .Z(n649) );
  NAND U970 ( .A(N48), .B(xregN_1), .Z(n648) );
  NAND U971 ( .A(n650), .B(n651), .Z(z2[43]) );
  NANDN U972 ( .A(xregN_1), .B(zin[42]), .Z(n651) );
  NAND U973 ( .A(N47), .B(xregN_1), .Z(n650) );
  NAND U974 ( .A(n652), .B(n653), .Z(z2[42]) );
  NANDN U975 ( .A(xregN_1), .B(zin[41]), .Z(n653) );
  NAND U976 ( .A(N46), .B(xregN_1), .Z(n652) );
  NAND U977 ( .A(n654), .B(n655), .Z(z2[41]) );
  NANDN U978 ( .A(xregN_1), .B(zin[40]), .Z(n655) );
  NAND U979 ( .A(N45), .B(xregN_1), .Z(n654) );
  NAND U980 ( .A(n656), .B(n657), .Z(z2[40]) );
  NANDN U981 ( .A(xregN_1), .B(zin[39]), .Z(n657) );
  NAND U982 ( .A(N44), .B(xregN_1), .Z(n656) );
  NAND U983 ( .A(n658), .B(n659), .Z(z2[3]) );
  NANDN U984 ( .A(xregN_1), .B(zin[2]), .Z(n659) );
  NAND U985 ( .A(N7), .B(xregN_1), .Z(n658) );
  NAND U986 ( .A(n660), .B(n661), .Z(z2[39]) );
  NANDN U987 ( .A(xregN_1), .B(zin[38]), .Z(n661) );
  NAND U988 ( .A(N43), .B(xregN_1), .Z(n660) );
  NAND U989 ( .A(n662), .B(n663), .Z(z2[38]) );
  NANDN U990 ( .A(xregN_1), .B(zin[37]), .Z(n663) );
  NAND U991 ( .A(N42), .B(xregN_1), .Z(n662) );
  NAND U992 ( .A(n664), .B(n665), .Z(z2[37]) );
  NANDN U993 ( .A(xregN_1), .B(zin[36]), .Z(n665) );
  NAND U994 ( .A(N41), .B(xregN_1), .Z(n664) );
  NAND U995 ( .A(n666), .B(n667), .Z(z2[36]) );
  NANDN U996 ( .A(xregN_1), .B(zin[35]), .Z(n667) );
  NAND U997 ( .A(N40), .B(xregN_1), .Z(n666) );
  NAND U998 ( .A(n668), .B(n669), .Z(z2[35]) );
  NANDN U999 ( .A(xregN_1), .B(zin[34]), .Z(n669) );
  NAND U1000 ( .A(N39), .B(xregN_1), .Z(n668) );
  NAND U1001 ( .A(n670), .B(n671), .Z(z2[34]) );
  NANDN U1002 ( .A(xregN_1), .B(zin[33]), .Z(n671) );
  NAND U1003 ( .A(N38), .B(xregN_1), .Z(n670) );
  NAND U1004 ( .A(n672), .B(n673), .Z(z2[33]) );
  NANDN U1005 ( .A(xregN_1), .B(zin[32]), .Z(n673) );
  NAND U1006 ( .A(N37), .B(xregN_1), .Z(n672) );
  NAND U1007 ( .A(n674), .B(n675), .Z(z2[32]) );
  NANDN U1008 ( .A(xregN_1), .B(zin[31]), .Z(n675) );
  NAND U1009 ( .A(N36), .B(xregN_1), .Z(n674) );
  NAND U1010 ( .A(n676), .B(n677), .Z(z2[31]) );
  NANDN U1011 ( .A(xregN_1), .B(zin[30]), .Z(n677) );
  NAND U1012 ( .A(N35), .B(xregN_1), .Z(n676) );
  NAND U1013 ( .A(n678), .B(n679), .Z(z2[30]) );
  NANDN U1014 ( .A(xregN_1), .B(zin[29]), .Z(n679) );
  NAND U1015 ( .A(N34), .B(xregN_1), .Z(n678) );
  NAND U1016 ( .A(n680), .B(n681), .Z(z2[2]) );
  NANDN U1017 ( .A(xregN_1), .B(zin[1]), .Z(n681) );
  NAND U1018 ( .A(N6), .B(xregN_1), .Z(n680) );
  NAND U1019 ( .A(n682), .B(n683), .Z(z2[29]) );
  NANDN U1020 ( .A(xregN_1), .B(zin[28]), .Z(n683) );
  NAND U1021 ( .A(N33), .B(xregN_1), .Z(n682) );
  NAND U1022 ( .A(n684), .B(n685), .Z(z2[28]) );
  NANDN U1023 ( .A(xregN_1), .B(zin[27]), .Z(n685) );
  NAND U1024 ( .A(N32), .B(xregN_1), .Z(n684) );
  NAND U1025 ( .A(n686), .B(n687), .Z(z2[27]) );
  NANDN U1026 ( .A(xregN_1), .B(zin[26]), .Z(n687) );
  NAND U1027 ( .A(N31), .B(xregN_1), .Z(n686) );
  NAND U1028 ( .A(n688), .B(n689), .Z(z2[26]) );
  NANDN U1029 ( .A(xregN_1), .B(zin[25]), .Z(n689) );
  NAND U1030 ( .A(N30), .B(xregN_1), .Z(n688) );
  NAND U1031 ( .A(n690), .B(n691), .Z(z2[25]) );
  NANDN U1032 ( .A(xregN_1), .B(zin[24]), .Z(n691) );
  NAND U1033 ( .A(N29), .B(xregN_1), .Z(n690) );
  NAND U1034 ( .A(n692), .B(n693), .Z(z2[257]) );
  NANDN U1035 ( .A(xregN_1), .B(zin[256]), .Z(n693) );
  NAND U1036 ( .A(N261), .B(xregN_1), .Z(n692) );
  NAND U1037 ( .A(n694), .B(n695), .Z(z2[256]) );
  NANDN U1038 ( .A(xregN_1), .B(zin[255]), .Z(n695) );
  NAND U1039 ( .A(N260), .B(xregN_1), .Z(n694) );
  NAND U1040 ( .A(n696), .B(n697), .Z(z2[255]) );
  NANDN U1041 ( .A(xregN_1), .B(zin[254]), .Z(n697) );
  NAND U1042 ( .A(N259), .B(xregN_1), .Z(n696) );
  NAND U1043 ( .A(n698), .B(n699), .Z(z2[254]) );
  NANDN U1044 ( .A(xregN_1), .B(zin[253]), .Z(n699) );
  NAND U1045 ( .A(N258), .B(xregN_1), .Z(n698) );
  NAND U1046 ( .A(n700), .B(n701), .Z(z2[253]) );
  NANDN U1047 ( .A(xregN_1), .B(zin[252]), .Z(n701) );
  NAND U1048 ( .A(N257), .B(xregN_1), .Z(n700) );
  NAND U1049 ( .A(n702), .B(n703), .Z(z2[252]) );
  NANDN U1050 ( .A(xregN_1), .B(zin[251]), .Z(n703) );
  NAND U1051 ( .A(N256), .B(xregN_1), .Z(n702) );
  NAND U1052 ( .A(n704), .B(n705), .Z(z2[251]) );
  NANDN U1053 ( .A(xregN_1), .B(zin[250]), .Z(n705) );
  NAND U1054 ( .A(N255), .B(xregN_1), .Z(n704) );
  NAND U1055 ( .A(n706), .B(n707), .Z(z2[250]) );
  NANDN U1056 ( .A(xregN_1), .B(zin[249]), .Z(n707) );
  NAND U1057 ( .A(N254), .B(xregN_1), .Z(n706) );
  NAND U1058 ( .A(n708), .B(n709), .Z(z2[24]) );
  NANDN U1059 ( .A(xregN_1), .B(zin[23]), .Z(n709) );
  NAND U1060 ( .A(N28), .B(xregN_1), .Z(n708) );
  NAND U1061 ( .A(n710), .B(n711), .Z(z2[249]) );
  NANDN U1062 ( .A(xregN_1), .B(zin[248]), .Z(n711) );
  NAND U1063 ( .A(N253), .B(xregN_1), .Z(n710) );
  NAND U1064 ( .A(n712), .B(n713), .Z(z2[248]) );
  NANDN U1065 ( .A(xregN_1), .B(zin[247]), .Z(n713) );
  NAND U1066 ( .A(N252), .B(xregN_1), .Z(n712) );
  NAND U1067 ( .A(n714), .B(n715), .Z(z2[247]) );
  NANDN U1068 ( .A(xregN_1), .B(zin[246]), .Z(n715) );
  NAND U1069 ( .A(N251), .B(xregN_1), .Z(n714) );
  NAND U1070 ( .A(n716), .B(n717), .Z(z2[246]) );
  NANDN U1071 ( .A(xregN_1), .B(zin[245]), .Z(n717) );
  NAND U1072 ( .A(N250), .B(xregN_1), .Z(n716) );
  NAND U1073 ( .A(n718), .B(n719), .Z(z2[245]) );
  NANDN U1074 ( .A(xregN_1), .B(zin[244]), .Z(n719) );
  NAND U1075 ( .A(N249), .B(xregN_1), .Z(n718) );
  NAND U1076 ( .A(n720), .B(n721), .Z(z2[244]) );
  NANDN U1077 ( .A(xregN_1), .B(zin[243]), .Z(n721) );
  NAND U1078 ( .A(N248), .B(xregN_1), .Z(n720) );
  NAND U1079 ( .A(n722), .B(n723), .Z(z2[243]) );
  NANDN U1080 ( .A(xregN_1), .B(zin[242]), .Z(n723) );
  NAND U1081 ( .A(N247), .B(xregN_1), .Z(n722) );
  NAND U1082 ( .A(n724), .B(n725), .Z(z2[242]) );
  NANDN U1083 ( .A(xregN_1), .B(zin[241]), .Z(n725) );
  NAND U1084 ( .A(N246), .B(xregN_1), .Z(n724) );
  NAND U1085 ( .A(n726), .B(n727), .Z(z2[241]) );
  NANDN U1086 ( .A(xregN_1), .B(zin[240]), .Z(n727) );
  NAND U1087 ( .A(N245), .B(xregN_1), .Z(n726) );
  NAND U1088 ( .A(n728), .B(n729), .Z(z2[240]) );
  NANDN U1089 ( .A(xregN_1), .B(zin[239]), .Z(n729) );
  NAND U1090 ( .A(N244), .B(xregN_1), .Z(n728) );
  NAND U1091 ( .A(n730), .B(n731), .Z(z2[23]) );
  NANDN U1092 ( .A(xregN_1), .B(zin[22]), .Z(n731) );
  NAND U1093 ( .A(N27), .B(xregN_1), .Z(n730) );
  NAND U1094 ( .A(n732), .B(n733), .Z(z2[239]) );
  NANDN U1095 ( .A(xregN_1), .B(zin[238]), .Z(n733) );
  NAND U1096 ( .A(N243), .B(xregN_1), .Z(n732) );
  NAND U1097 ( .A(n734), .B(n735), .Z(z2[238]) );
  NANDN U1098 ( .A(xregN_1), .B(zin[237]), .Z(n735) );
  NAND U1099 ( .A(N242), .B(xregN_1), .Z(n734) );
  NAND U1100 ( .A(n736), .B(n737), .Z(z2[237]) );
  NANDN U1101 ( .A(xregN_1), .B(zin[236]), .Z(n737) );
  NAND U1102 ( .A(N241), .B(xregN_1), .Z(n736) );
  NAND U1103 ( .A(n738), .B(n739), .Z(z2[236]) );
  NANDN U1104 ( .A(xregN_1), .B(zin[235]), .Z(n739) );
  NAND U1105 ( .A(N240), .B(xregN_1), .Z(n738) );
  NAND U1106 ( .A(n740), .B(n741), .Z(z2[235]) );
  NANDN U1107 ( .A(xregN_1), .B(zin[234]), .Z(n741) );
  NAND U1108 ( .A(N239), .B(xregN_1), .Z(n740) );
  NAND U1109 ( .A(n742), .B(n743), .Z(z2[234]) );
  NANDN U1110 ( .A(xregN_1), .B(zin[233]), .Z(n743) );
  NAND U1111 ( .A(N238), .B(xregN_1), .Z(n742) );
  NAND U1112 ( .A(n744), .B(n745), .Z(z2[233]) );
  NANDN U1113 ( .A(xregN_1), .B(zin[232]), .Z(n745) );
  NAND U1114 ( .A(N237), .B(xregN_1), .Z(n744) );
  NAND U1115 ( .A(n746), .B(n747), .Z(z2[232]) );
  NANDN U1116 ( .A(xregN_1), .B(zin[231]), .Z(n747) );
  NAND U1117 ( .A(N236), .B(xregN_1), .Z(n746) );
  NAND U1118 ( .A(n748), .B(n749), .Z(z2[231]) );
  NANDN U1119 ( .A(xregN_1), .B(zin[230]), .Z(n749) );
  NAND U1120 ( .A(N235), .B(xregN_1), .Z(n748) );
  NAND U1121 ( .A(n750), .B(n751), .Z(z2[230]) );
  NANDN U1122 ( .A(xregN_1), .B(zin[229]), .Z(n751) );
  NAND U1123 ( .A(N234), .B(xregN_1), .Z(n750) );
  NAND U1124 ( .A(n752), .B(n753), .Z(z2[22]) );
  NANDN U1125 ( .A(xregN_1), .B(zin[21]), .Z(n753) );
  NAND U1126 ( .A(N26), .B(xregN_1), .Z(n752) );
  NAND U1127 ( .A(n754), .B(n755), .Z(z2[229]) );
  NANDN U1128 ( .A(xregN_1), .B(zin[228]), .Z(n755) );
  NAND U1129 ( .A(N233), .B(xregN_1), .Z(n754) );
  NAND U1130 ( .A(n756), .B(n757), .Z(z2[228]) );
  NANDN U1131 ( .A(xregN_1), .B(zin[227]), .Z(n757) );
  NAND U1132 ( .A(N232), .B(xregN_1), .Z(n756) );
  NAND U1133 ( .A(n758), .B(n759), .Z(z2[227]) );
  NANDN U1134 ( .A(xregN_1), .B(zin[226]), .Z(n759) );
  NAND U1135 ( .A(N231), .B(xregN_1), .Z(n758) );
  NAND U1136 ( .A(n760), .B(n761), .Z(z2[226]) );
  NANDN U1137 ( .A(xregN_1), .B(zin[225]), .Z(n761) );
  NAND U1138 ( .A(N230), .B(xregN_1), .Z(n760) );
  NAND U1139 ( .A(n762), .B(n763), .Z(z2[225]) );
  NANDN U1140 ( .A(xregN_1), .B(zin[224]), .Z(n763) );
  NAND U1141 ( .A(N229), .B(xregN_1), .Z(n762) );
  NAND U1142 ( .A(n764), .B(n765), .Z(z2[224]) );
  NANDN U1143 ( .A(xregN_1), .B(zin[223]), .Z(n765) );
  NAND U1144 ( .A(N228), .B(xregN_1), .Z(n764) );
  NAND U1145 ( .A(n766), .B(n767), .Z(z2[223]) );
  NANDN U1146 ( .A(xregN_1), .B(zin[222]), .Z(n767) );
  NAND U1147 ( .A(N227), .B(xregN_1), .Z(n766) );
  NAND U1148 ( .A(n768), .B(n769), .Z(z2[222]) );
  NANDN U1149 ( .A(xregN_1), .B(zin[221]), .Z(n769) );
  NAND U1150 ( .A(N226), .B(xregN_1), .Z(n768) );
  NAND U1151 ( .A(n770), .B(n771), .Z(z2[221]) );
  NANDN U1152 ( .A(xregN_1), .B(zin[220]), .Z(n771) );
  NAND U1153 ( .A(N225), .B(xregN_1), .Z(n770) );
  NAND U1154 ( .A(n772), .B(n773), .Z(z2[220]) );
  NANDN U1155 ( .A(xregN_1), .B(zin[219]), .Z(n773) );
  NAND U1156 ( .A(N224), .B(xregN_1), .Z(n772) );
  NAND U1157 ( .A(n774), .B(n775), .Z(z2[21]) );
  NANDN U1158 ( .A(xregN_1), .B(zin[20]), .Z(n775) );
  NAND U1159 ( .A(N25), .B(xregN_1), .Z(n774) );
  NAND U1160 ( .A(n776), .B(n777), .Z(z2[219]) );
  NANDN U1161 ( .A(xregN_1), .B(zin[218]), .Z(n777) );
  NAND U1162 ( .A(N223), .B(xregN_1), .Z(n776) );
  NAND U1163 ( .A(n778), .B(n779), .Z(z2[218]) );
  NANDN U1164 ( .A(xregN_1), .B(zin[217]), .Z(n779) );
  NAND U1165 ( .A(N222), .B(xregN_1), .Z(n778) );
  NAND U1166 ( .A(n780), .B(n781), .Z(z2[217]) );
  NANDN U1167 ( .A(xregN_1), .B(zin[216]), .Z(n781) );
  NAND U1168 ( .A(N221), .B(xregN_1), .Z(n780) );
  NAND U1169 ( .A(n782), .B(n783), .Z(z2[216]) );
  NANDN U1170 ( .A(xregN_1), .B(zin[215]), .Z(n783) );
  NAND U1171 ( .A(N220), .B(xregN_1), .Z(n782) );
  NAND U1172 ( .A(n784), .B(n785), .Z(z2[215]) );
  NANDN U1173 ( .A(xregN_1), .B(zin[214]), .Z(n785) );
  NAND U1174 ( .A(N219), .B(xregN_1), .Z(n784) );
  NAND U1175 ( .A(n786), .B(n787), .Z(z2[214]) );
  NANDN U1176 ( .A(xregN_1), .B(zin[213]), .Z(n787) );
  NAND U1177 ( .A(N218), .B(xregN_1), .Z(n786) );
  NAND U1178 ( .A(n788), .B(n789), .Z(z2[213]) );
  NANDN U1179 ( .A(xregN_1), .B(zin[212]), .Z(n789) );
  NAND U1180 ( .A(N217), .B(xregN_1), .Z(n788) );
  NAND U1181 ( .A(n790), .B(n791), .Z(z2[212]) );
  NANDN U1182 ( .A(xregN_1), .B(zin[211]), .Z(n791) );
  NAND U1183 ( .A(N216), .B(xregN_1), .Z(n790) );
  NAND U1184 ( .A(n792), .B(n793), .Z(z2[211]) );
  NANDN U1185 ( .A(xregN_1), .B(zin[210]), .Z(n793) );
  NAND U1186 ( .A(N215), .B(xregN_1), .Z(n792) );
  NAND U1187 ( .A(n794), .B(n795), .Z(z2[210]) );
  NANDN U1188 ( .A(xregN_1), .B(zin[209]), .Z(n795) );
  NAND U1189 ( .A(N214), .B(xregN_1), .Z(n794) );
  NAND U1190 ( .A(n796), .B(n797), .Z(z2[20]) );
  NANDN U1191 ( .A(xregN_1), .B(zin[19]), .Z(n797) );
  NAND U1192 ( .A(N24), .B(xregN_1), .Z(n796) );
  NAND U1193 ( .A(n798), .B(n799), .Z(z2[209]) );
  NANDN U1194 ( .A(xregN_1), .B(zin[208]), .Z(n799) );
  NAND U1195 ( .A(N213), .B(xregN_1), .Z(n798) );
  NAND U1196 ( .A(n800), .B(n801), .Z(z2[208]) );
  NANDN U1197 ( .A(xregN_1), .B(zin[207]), .Z(n801) );
  NAND U1198 ( .A(N212), .B(xregN_1), .Z(n800) );
  NAND U1199 ( .A(n802), .B(n803), .Z(z2[207]) );
  NANDN U1200 ( .A(xregN_1), .B(zin[206]), .Z(n803) );
  NAND U1201 ( .A(N211), .B(xregN_1), .Z(n802) );
  NAND U1202 ( .A(n804), .B(n805), .Z(z2[206]) );
  NANDN U1203 ( .A(xregN_1), .B(zin[205]), .Z(n805) );
  NAND U1204 ( .A(N210), .B(xregN_1), .Z(n804) );
  NAND U1205 ( .A(n806), .B(n807), .Z(z2[205]) );
  NANDN U1206 ( .A(xregN_1), .B(zin[204]), .Z(n807) );
  NAND U1207 ( .A(N209), .B(xregN_1), .Z(n806) );
  NAND U1208 ( .A(n808), .B(n809), .Z(z2[204]) );
  NANDN U1209 ( .A(xregN_1), .B(zin[203]), .Z(n809) );
  NAND U1210 ( .A(N208), .B(xregN_1), .Z(n808) );
  NAND U1211 ( .A(n810), .B(n811), .Z(z2[203]) );
  NANDN U1212 ( .A(xregN_1), .B(zin[202]), .Z(n811) );
  NAND U1213 ( .A(N207), .B(xregN_1), .Z(n810) );
  NAND U1214 ( .A(n812), .B(n813), .Z(z2[202]) );
  NANDN U1215 ( .A(xregN_1), .B(zin[201]), .Z(n813) );
  NAND U1216 ( .A(N206), .B(xregN_1), .Z(n812) );
  NAND U1217 ( .A(n814), .B(n815), .Z(z2[201]) );
  NANDN U1218 ( .A(xregN_1), .B(zin[200]), .Z(n815) );
  NAND U1219 ( .A(N205), .B(xregN_1), .Z(n814) );
  NAND U1220 ( .A(n816), .B(n817), .Z(z2[200]) );
  NANDN U1221 ( .A(xregN_1), .B(zin[199]), .Z(n817) );
  NAND U1222 ( .A(N204), .B(xregN_1), .Z(n816) );
  NAND U1223 ( .A(n818), .B(n819), .Z(z2[1]) );
  NANDN U1224 ( .A(xregN_1), .B(zin[0]), .Z(n819) );
  NAND U1225 ( .A(N5), .B(xregN_1), .Z(n818) );
  NAND U1226 ( .A(n820), .B(n821), .Z(z2[19]) );
  NANDN U1227 ( .A(xregN_1), .B(zin[18]), .Z(n821) );
  NAND U1228 ( .A(N23), .B(xregN_1), .Z(n820) );
  NAND U1229 ( .A(n822), .B(n823), .Z(z2[199]) );
  NANDN U1230 ( .A(xregN_1), .B(zin[198]), .Z(n823) );
  NAND U1231 ( .A(N203), .B(xregN_1), .Z(n822) );
  NAND U1232 ( .A(n824), .B(n825), .Z(z2[198]) );
  NANDN U1233 ( .A(xregN_1), .B(zin[197]), .Z(n825) );
  NAND U1234 ( .A(N202), .B(xregN_1), .Z(n824) );
  NAND U1235 ( .A(n826), .B(n827), .Z(z2[197]) );
  NANDN U1236 ( .A(xregN_1), .B(zin[196]), .Z(n827) );
  NAND U1237 ( .A(N201), .B(xregN_1), .Z(n826) );
  NAND U1238 ( .A(n828), .B(n829), .Z(z2[196]) );
  NANDN U1239 ( .A(xregN_1), .B(zin[195]), .Z(n829) );
  NAND U1240 ( .A(N200), .B(xregN_1), .Z(n828) );
  NAND U1241 ( .A(n830), .B(n831), .Z(z2[195]) );
  NANDN U1242 ( .A(xregN_1), .B(zin[194]), .Z(n831) );
  NAND U1243 ( .A(N199), .B(xregN_1), .Z(n830) );
  NAND U1244 ( .A(n832), .B(n833), .Z(z2[194]) );
  NANDN U1245 ( .A(xregN_1), .B(zin[193]), .Z(n833) );
  NAND U1246 ( .A(N198), .B(xregN_1), .Z(n832) );
  NAND U1247 ( .A(n834), .B(n835), .Z(z2[193]) );
  NANDN U1248 ( .A(xregN_1), .B(zin[192]), .Z(n835) );
  NAND U1249 ( .A(N197), .B(xregN_1), .Z(n834) );
  NAND U1250 ( .A(n836), .B(n837), .Z(z2[192]) );
  NANDN U1251 ( .A(xregN_1), .B(zin[191]), .Z(n837) );
  NAND U1252 ( .A(N196), .B(xregN_1), .Z(n836) );
  NAND U1253 ( .A(n838), .B(n839), .Z(z2[191]) );
  NANDN U1254 ( .A(xregN_1), .B(zin[190]), .Z(n839) );
  NAND U1255 ( .A(N195), .B(xregN_1), .Z(n838) );
  NAND U1256 ( .A(n840), .B(n841), .Z(z2[190]) );
  NANDN U1257 ( .A(xregN_1), .B(zin[189]), .Z(n841) );
  NAND U1258 ( .A(N194), .B(xregN_1), .Z(n840) );
  NAND U1259 ( .A(n842), .B(n843), .Z(z2[18]) );
  NANDN U1260 ( .A(xregN_1), .B(zin[17]), .Z(n843) );
  NAND U1261 ( .A(N22), .B(xregN_1), .Z(n842) );
  NAND U1262 ( .A(n844), .B(n845), .Z(z2[189]) );
  NANDN U1263 ( .A(xregN_1), .B(zin[188]), .Z(n845) );
  NAND U1264 ( .A(N193), .B(xregN_1), .Z(n844) );
  NAND U1265 ( .A(n846), .B(n847), .Z(z2[188]) );
  NANDN U1266 ( .A(xregN_1), .B(zin[187]), .Z(n847) );
  NAND U1267 ( .A(N192), .B(xregN_1), .Z(n846) );
  NAND U1268 ( .A(n848), .B(n849), .Z(z2[187]) );
  NANDN U1269 ( .A(xregN_1), .B(zin[186]), .Z(n849) );
  NAND U1270 ( .A(N191), .B(xregN_1), .Z(n848) );
  NAND U1271 ( .A(n850), .B(n851), .Z(z2[186]) );
  NANDN U1272 ( .A(xregN_1), .B(zin[185]), .Z(n851) );
  NAND U1273 ( .A(N190), .B(xregN_1), .Z(n850) );
  NAND U1274 ( .A(n852), .B(n853), .Z(z2[185]) );
  NANDN U1275 ( .A(xregN_1), .B(zin[184]), .Z(n853) );
  NAND U1276 ( .A(N189), .B(xregN_1), .Z(n852) );
  NAND U1277 ( .A(n854), .B(n855), .Z(z2[184]) );
  NANDN U1278 ( .A(xregN_1), .B(zin[183]), .Z(n855) );
  NAND U1279 ( .A(N188), .B(xregN_1), .Z(n854) );
  NAND U1280 ( .A(n856), .B(n857), .Z(z2[183]) );
  NANDN U1281 ( .A(xregN_1), .B(zin[182]), .Z(n857) );
  NAND U1282 ( .A(N187), .B(xregN_1), .Z(n856) );
  NAND U1283 ( .A(n858), .B(n859), .Z(z2[182]) );
  NANDN U1284 ( .A(xregN_1), .B(zin[181]), .Z(n859) );
  NAND U1285 ( .A(N186), .B(xregN_1), .Z(n858) );
  NAND U1286 ( .A(n860), .B(n861), .Z(z2[181]) );
  NANDN U1287 ( .A(xregN_1), .B(zin[180]), .Z(n861) );
  NAND U1288 ( .A(N185), .B(xregN_1), .Z(n860) );
  NAND U1289 ( .A(n862), .B(n863), .Z(z2[180]) );
  NANDN U1290 ( .A(xregN_1), .B(zin[179]), .Z(n863) );
  NAND U1291 ( .A(N184), .B(xregN_1), .Z(n862) );
  NAND U1292 ( .A(n864), .B(n865), .Z(z2[17]) );
  NANDN U1293 ( .A(xregN_1), .B(zin[16]), .Z(n865) );
  NAND U1294 ( .A(N21), .B(xregN_1), .Z(n864) );
  NAND U1295 ( .A(n866), .B(n867), .Z(z2[179]) );
  NANDN U1296 ( .A(xregN_1), .B(zin[178]), .Z(n867) );
  NAND U1297 ( .A(N183), .B(xregN_1), .Z(n866) );
  NAND U1298 ( .A(n868), .B(n869), .Z(z2[178]) );
  NANDN U1299 ( .A(xregN_1), .B(zin[177]), .Z(n869) );
  NAND U1300 ( .A(N182), .B(xregN_1), .Z(n868) );
  NAND U1301 ( .A(n870), .B(n871), .Z(z2[177]) );
  NANDN U1302 ( .A(xregN_1), .B(zin[176]), .Z(n871) );
  NAND U1303 ( .A(N181), .B(xregN_1), .Z(n870) );
  NAND U1304 ( .A(n872), .B(n873), .Z(z2[176]) );
  NANDN U1305 ( .A(xregN_1), .B(zin[175]), .Z(n873) );
  NAND U1306 ( .A(N180), .B(xregN_1), .Z(n872) );
  NAND U1307 ( .A(n874), .B(n875), .Z(z2[175]) );
  NANDN U1308 ( .A(xregN_1), .B(zin[174]), .Z(n875) );
  NAND U1309 ( .A(N179), .B(xregN_1), .Z(n874) );
  NAND U1310 ( .A(n876), .B(n877), .Z(z2[174]) );
  NANDN U1311 ( .A(xregN_1), .B(zin[173]), .Z(n877) );
  NAND U1312 ( .A(N178), .B(xregN_1), .Z(n876) );
  NAND U1313 ( .A(n878), .B(n879), .Z(z2[173]) );
  NANDN U1314 ( .A(xregN_1), .B(zin[172]), .Z(n879) );
  NAND U1315 ( .A(N177), .B(xregN_1), .Z(n878) );
  NAND U1316 ( .A(n880), .B(n881), .Z(z2[172]) );
  NANDN U1317 ( .A(xregN_1), .B(zin[171]), .Z(n881) );
  NAND U1318 ( .A(N176), .B(xregN_1), .Z(n880) );
  NAND U1319 ( .A(n882), .B(n883), .Z(z2[171]) );
  NANDN U1320 ( .A(xregN_1), .B(zin[170]), .Z(n883) );
  NAND U1321 ( .A(N175), .B(xregN_1), .Z(n882) );
  NAND U1322 ( .A(n884), .B(n885), .Z(z2[170]) );
  NANDN U1323 ( .A(xregN_1), .B(zin[169]), .Z(n885) );
  NAND U1324 ( .A(N174), .B(xregN_1), .Z(n884) );
  NAND U1325 ( .A(n886), .B(n887), .Z(z2[16]) );
  NANDN U1326 ( .A(xregN_1), .B(zin[15]), .Z(n887) );
  NAND U1327 ( .A(N20), .B(xregN_1), .Z(n886) );
  NAND U1328 ( .A(n888), .B(n889), .Z(z2[169]) );
  NANDN U1329 ( .A(xregN_1), .B(zin[168]), .Z(n889) );
  NAND U1330 ( .A(N173), .B(xregN_1), .Z(n888) );
  NAND U1331 ( .A(n890), .B(n891), .Z(z2[168]) );
  NANDN U1332 ( .A(xregN_1), .B(zin[167]), .Z(n891) );
  NAND U1333 ( .A(N172), .B(xregN_1), .Z(n890) );
  NAND U1334 ( .A(n892), .B(n893), .Z(z2[167]) );
  NANDN U1335 ( .A(xregN_1), .B(zin[166]), .Z(n893) );
  NAND U1336 ( .A(N171), .B(xregN_1), .Z(n892) );
  NAND U1337 ( .A(n894), .B(n895), .Z(z2[166]) );
  NANDN U1338 ( .A(xregN_1), .B(zin[165]), .Z(n895) );
  NAND U1339 ( .A(N170), .B(xregN_1), .Z(n894) );
  NAND U1340 ( .A(n896), .B(n897), .Z(z2[165]) );
  NANDN U1341 ( .A(xregN_1), .B(zin[164]), .Z(n897) );
  NAND U1342 ( .A(N169), .B(xregN_1), .Z(n896) );
  NAND U1343 ( .A(n898), .B(n899), .Z(z2[164]) );
  NANDN U1344 ( .A(xregN_1), .B(zin[163]), .Z(n899) );
  NAND U1345 ( .A(N168), .B(xregN_1), .Z(n898) );
  NAND U1346 ( .A(n900), .B(n901), .Z(z2[163]) );
  NANDN U1347 ( .A(xregN_1), .B(zin[162]), .Z(n901) );
  NAND U1348 ( .A(N167), .B(xregN_1), .Z(n900) );
  NAND U1349 ( .A(n902), .B(n903), .Z(z2[162]) );
  NANDN U1350 ( .A(xregN_1), .B(zin[161]), .Z(n903) );
  NAND U1351 ( .A(N166), .B(xregN_1), .Z(n902) );
  NAND U1352 ( .A(n904), .B(n905), .Z(z2[161]) );
  NANDN U1353 ( .A(xregN_1), .B(zin[160]), .Z(n905) );
  NAND U1354 ( .A(N165), .B(xregN_1), .Z(n904) );
  NAND U1355 ( .A(n906), .B(n907), .Z(z2[160]) );
  NANDN U1356 ( .A(xregN_1), .B(zin[159]), .Z(n907) );
  NAND U1357 ( .A(N164), .B(xregN_1), .Z(n906) );
  NAND U1358 ( .A(n908), .B(n909), .Z(z2[15]) );
  NANDN U1359 ( .A(xregN_1), .B(zin[14]), .Z(n909) );
  NAND U1360 ( .A(N19), .B(xregN_1), .Z(n908) );
  NAND U1361 ( .A(n910), .B(n911), .Z(z2[159]) );
  NANDN U1362 ( .A(xregN_1), .B(zin[158]), .Z(n911) );
  NAND U1363 ( .A(N163), .B(xregN_1), .Z(n910) );
  NAND U1364 ( .A(n912), .B(n913), .Z(z2[158]) );
  NANDN U1365 ( .A(xregN_1), .B(zin[157]), .Z(n913) );
  NAND U1366 ( .A(N162), .B(xregN_1), .Z(n912) );
  NAND U1367 ( .A(n914), .B(n915), .Z(z2[157]) );
  NANDN U1368 ( .A(xregN_1), .B(zin[156]), .Z(n915) );
  NAND U1369 ( .A(N161), .B(xregN_1), .Z(n914) );
  NAND U1370 ( .A(n916), .B(n917), .Z(z2[156]) );
  NANDN U1371 ( .A(xregN_1), .B(zin[155]), .Z(n917) );
  NAND U1372 ( .A(N160), .B(xregN_1), .Z(n916) );
  NAND U1373 ( .A(n918), .B(n919), .Z(z2[155]) );
  NANDN U1374 ( .A(xregN_1), .B(zin[154]), .Z(n919) );
  NAND U1375 ( .A(N159), .B(xregN_1), .Z(n918) );
  NAND U1376 ( .A(n920), .B(n921), .Z(z2[154]) );
  NANDN U1377 ( .A(xregN_1), .B(zin[153]), .Z(n921) );
  NAND U1378 ( .A(N158), .B(xregN_1), .Z(n920) );
  NAND U1379 ( .A(n922), .B(n923), .Z(z2[153]) );
  NANDN U1380 ( .A(xregN_1), .B(zin[152]), .Z(n923) );
  NAND U1381 ( .A(N157), .B(xregN_1), .Z(n922) );
  NAND U1382 ( .A(n924), .B(n925), .Z(z2[152]) );
  NANDN U1383 ( .A(xregN_1), .B(zin[151]), .Z(n925) );
  NAND U1384 ( .A(N156), .B(xregN_1), .Z(n924) );
  NAND U1385 ( .A(n926), .B(n927), .Z(z2[151]) );
  NANDN U1386 ( .A(xregN_1), .B(zin[150]), .Z(n927) );
  NAND U1387 ( .A(N155), .B(xregN_1), .Z(n926) );
  NAND U1388 ( .A(n928), .B(n929), .Z(z2[150]) );
  NANDN U1389 ( .A(xregN_1), .B(zin[149]), .Z(n929) );
  NAND U1390 ( .A(N154), .B(xregN_1), .Z(n928) );
  NAND U1391 ( .A(n930), .B(n931), .Z(z2[14]) );
  NANDN U1392 ( .A(xregN_1), .B(zin[13]), .Z(n931) );
  NAND U1393 ( .A(N18), .B(xregN_1), .Z(n930) );
  NAND U1394 ( .A(n932), .B(n933), .Z(z2[149]) );
  NANDN U1395 ( .A(xregN_1), .B(zin[148]), .Z(n933) );
  NAND U1396 ( .A(N153), .B(xregN_1), .Z(n932) );
  NAND U1397 ( .A(n934), .B(n935), .Z(z2[148]) );
  NANDN U1398 ( .A(xregN_1), .B(zin[147]), .Z(n935) );
  NAND U1399 ( .A(N152), .B(xregN_1), .Z(n934) );
  NAND U1400 ( .A(n936), .B(n937), .Z(z2[147]) );
  NANDN U1401 ( .A(xregN_1), .B(zin[146]), .Z(n937) );
  NAND U1402 ( .A(N151), .B(xregN_1), .Z(n936) );
  NAND U1403 ( .A(n938), .B(n939), .Z(z2[146]) );
  NANDN U1404 ( .A(xregN_1), .B(zin[145]), .Z(n939) );
  NAND U1405 ( .A(N150), .B(xregN_1), .Z(n938) );
  NAND U1406 ( .A(n940), .B(n941), .Z(z2[145]) );
  NANDN U1407 ( .A(xregN_1), .B(zin[144]), .Z(n941) );
  NAND U1408 ( .A(N149), .B(xregN_1), .Z(n940) );
  NAND U1409 ( .A(n942), .B(n943), .Z(z2[144]) );
  NANDN U1410 ( .A(xregN_1), .B(zin[143]), .Z(n943) );
  NAND U1411 ( .A(N148), .B(xregN_1), .Z(n942) );
  NAND U1412 ( .A(n944), .B(n945), .Z(z2[143]) );
  NANDN U1413 ( .A(xregN_1), .B(zin[142]), .Z(n945) );
  NAND U1414 ( .A(N147), .B(xregN_1), .Z(n944) );
  NAND U1415 ( .A(n946), .B(n947), .Z(z2[142]) );
  NANDN U1416 ( .A(xregN_1), .B(zin[141]), .Z(n947) );
  NAND U1417 ( .A(N146), .B(xregN_1), .Z(n946) );
  NAND U1418 ( .A(n948), .B(n949), .Z(z2[141]) );
  NANDN U1419 ( .A(xregN_1), .B(zin[140]), .Z(n949) );
  NAND U1420 ( .A(N145), .B(xregN_1), .Z(n948) );
  NAND U1421 ( .A(n950), .B(n951), .Z(z2[140]) );
  NANDN U1422 ( .A(xregN_1), .B(zin[139]), .Z(n951) );
  NAND U1423 ( .A(N144), .B(xregN_1), .Z(n950) );
  NAND U1424 ( .A(n952), .B(n953), .Z(z2[13]) );
  NANDN U1425 ( .A(xregN_1), .B(zin[12]), .Z(n953) );
  NAND U1426 ( .A(N17), .B(xregN_1), .Z(n952) );
  NAND U1427 ( .A(n954), .B(n955), .Z(z2[139]) );
  NANDN U1428 ( .A(xregN_1), .B(zin[138]), .Z(n955) );
  NAND U1429 ( .A(N143), .B(xregN_1), .Z(n954) );
  NAND U1430 ( .A(n956), .B(n957), .Z(z2[138]) );
  NANDN U1431 ( .A(xregN_1), .B(zin[137]), .Z(n957) );
  NAND U1432 ( .A(N142), .B(xregN_1), .Z(n956) );
  NAND U1433 ( .A(n958), .B(n959), .Z(z2[137]) );
  NANDN U1434 ( .A(xregN_1), .B(zin[136]), .Z(n959) );
  NAND U1435 ( .A(N141), .B(xregN_1), .Z(n958) );
  NAND U1436 ( .A(n960), .B(n961), .Z(z2[136]) );
  NANDN U1437 ( .A(xregN_1), .B(zin[135]), .Z(n961) );
  NAND U1438 ( .A(N140), .B(xregN_1), .Z(n960) );
  NAND U1439 ( .A(n962), .B(n963), .Z(z2[135]) );
  NANDN U1440 ( .A(xregN_1), .B(zin[134]), .Z(n963) );
  NAND U1441 ( .A(N139), .B(xregN_1), .Z(n962) );
  NAND U1442 ( .A(n964), .B(n965), .Z(z2[134]) );
  NANDN U1443 ( .A(xregN_1), .B(zin[133]), .Z(n965) );
  NAND U1444 ( .A(N138), .B(xregN_1), .Z(n964) );
  NAND U1445 ( .A(n966), .B(n967), .Z(z2[133]) );
  NANDN U1446 ( .A(xregN_1), .B(zin[132]), .Z(n967) );
  NAND U1447 ( .A(N137), .B(xregN_1), .Z(n966) );
  NAND U1448 ( .A(n968), .B(n969), .Z(z2[132]) );
  NANDN U1449 ( .A(xregN_1), .B(zin[131]), .Z(n969) );
  NAND U1450 ( .A(N136), .B(xregN_1), .Z(n968) );
  NAND U1451 ( .A(n970), .B(n971), .Z(z2[131]) );
  NANDN U1452 ( .A(xregN_1), .B(zin[130]), .Z(n971) );
  NAND U1453 ( .A(N135), .B(xregN_1), .Z(n970) );
  NAND U1454 ( .A(n972), .B(n973), .Z(z2[130]) );
  NANDN U1455 ( .A(xregN_1), .B(zin[129]), .Z(n973) );
  NAND U1456 ( .A(N134), .B(xregN_1), .Z(n972) );
  NAND U1457 ( .A(n974), .B(n975), .Z(z2[12]) );
  NANDN U1458 ( .A(xregN_1), .B(zin[11]), .Z(n975) );
  NAND U1459 ( .A(N16), .B(xregN_1), .Z(n974) );
  NAND U1460 ( .A(n976), .B(n977), .Z(z2[129]) );
  NANDN U1461 ( .A(xregN_1), .B(zin[128]), .Z(n977) );
  NAND U1462 ( .A(N133), .B(xregN_1), .Z(n976) );
  NAND U1463 ( .A(n978), .B(n979), .Z(z2[128]) );
  NANDN U1464 ( .A(xregN_1), .B(zin[127]), .Z(n979) );
  NAND U1465 ( .A(N132), .B(xregN_1), .Z(n978) );
  NAND U1466 ( .A(n980), .B(n981), .Z(z2[127]) );
  NANDN U1467 ( .A(xregN_1), .B(zin[126]), .Z(n981) );
  NAND U1468 ( .A(N131), .B(xregN_1), .Z(n980) );
  NAND U1469 ( .A(n982), .B(n983), .Z(z2[126]) );
  NANDN U1470 ( .A(xregN_1), .B(zin[125]), .Z(n983) );
  NAND U1471 ( .A(N130), .B(xregN_1), .Z(n982) );
  NAND U1472 ( .A(n984), .B(n985), .Z(z2[125]) );
  NANDN U1473 ( .A(xregN_1), .B(zin[124]), .Z(n985) );
  NAND U1474 ( .A(N129), .B(xregN_1), .Z(n984) );
  NAND U1475 ( .A(n986), .B(n987), .Z(z2[124]) );
  NANDN U1476 ( .A(xregN_1), .B(zin[123]), .Z(n987) );
  NAND U1477 ( .A(N128), .B(xregN_1), .Z(n986) );
  NAND U1478 ( .A(n988), .B(n989), .Z(z2[123]) );
  NANDN U1479 ( .A(xregN_1), .B(zin[122]), .Z(n989) );
  NAND U1480 ( .A(N127), .B(xregN_1), .Z(n988) );
  NAND U1481 ( .A(n990), .B(n991), .Z(z2[122]) );
  NANDN U1482 ( .A(xregN_1), .B(zin[121]), .Z(n991) );
  NAND U1483 ( .A(N126), .B(xregN_1), .Z(n990) );
  NAND U1484 ( .A(n992), .B(n993), .Z(z2[121]) );
  NANDN U1485 ( .A(xregN_1), .B(zin[120]), .Z(n993) );
  NAND U1486 ( .A(N125), .B(xregN_1), .Z(n992) );
  NAND U1487 ( .A(n994), .B(n995), .Z(z2[120]) );
  NANDN U1488 ( .A(xregN_1), .B(zin[119]), .Z(n995) );
  NAND U1489 ( .A(N124), .B(xregN_1), .Z(n994) );
  NAND U1490 ( .A(n996), .B(n997), .Z(z2[11]) );
  NANDN U1491 ( .A(xregN_1), .B(zin[10]), .Z(n997) );
  NAND U1492 ( .A(N15), .B(xregN_1), .Z(n996) );
  NAND U1493 ( .A(n998), .B(n999), .Z(z2[119]) );
  NANDN U1494 ( .A(xregN_1), .B(zin[118]), .Z(n999) );
  NAND U1495 ( .A(N123), .B(xregN_1), .Z(n998) );
  NAND U1496 ( .A(n1000), .B(n1001), .Z(z2[118]) );
  NANDN U1497 ( .A(xregN_1), .B(zin[117]), .Z(n1001) );
  NAND U1498 ( .A(N122), .B(xregN_1), .Z(n1000) );
  NAND U1499 ( .A(n1002), .B(n1003), .Z(z2[117]) );
  NANDN U1500 ( .A(xregN_1), .B(zin[116]), .Z(n1003) );
  NAND U1501 ( .A(N121), .B(xregN_1), .Z(n1002) );
  NAND U1502 ( .A(n1004), .B(n1005), .Z(z2[116]) );
  NANDN U1503 ( .A(xregN_1), .B(zin[115]), .Z(n1005) );
  NAND U1504 ( .A(N120), .B(xregN_1), .Z(n1004) );
  NAND U1505 ( .A(n1006), .B(n1007), .Z(z2[115]) );
  NANDN U1506 ( .A(xregN_1), .B(zin[114]), .Z(n1007) );
  NAND U1507 ( .A(N119), .B(xregN_1), .Z(n1006) );
  NAND U1508 ( .A(n1008), .B(n1009), .Z(z2[114]) );
  NANDN U1509 ( .A(xregN_1), .B(zin[113]), .Z(n1009) );
  NAND U1510 ( .A(N118), .B(xregN_1), .Z(n1008) );
  NAND U1511 ( .A(n1010), .B(n1011), .Z(z2[113]) );
  NANDN U1512 ( .A(xregN_1), .B(zin[112]), .Z(n1011) );
  NAND U1513 ( .A(N117), .B(xregN_1), .Z(n1010) );
  NAND U1514 ( .A(n1012), .B(n1013), .Z(z2[112]) );
  NANDN U1515 ( .A(xregN_1), .B(zin[111]), .Z(n1013) );
  NAND U1516 ( .A(N116), .B(xregN_1), .Z(n1012) );
  NAND U1517 ( .A(n1014), .B(n1015), .Z(z2[111]) );
  NANDN U1518 ( .A(xregN_1), .B(zin[110]), .Z(n1015) );
  NAND U1519 ( .A(N115), .B(xregN_1), .Z(n1014) );
  NAND U1520 ( .A(n1016), .B(n1017), .Z(z2[110]) );
  NANDN U1521 ( .A(xregN_1), .B(zin[109]), .Z(n1017) );
  NAND U1522 ( .A(N114), .B(xregN_1), .Z(n1016) );
  NAND U1523 ( .A(n1018), .B(n1019), .Z(z2[10]) );
  NANDN U1524 ( .A(xregN_1), .B(zin[9]), .Z(n1019) );
  NAND U1525 ( .A(N14), .B(xregN_1), .Z(n1018) );
  NAND U1526 ( .A(n1020), .B(n1021), .Z(z2[109]) );
  NANDN U1527 ( .A(xregN_1), .B(zin[108]), .Z(n1021) );
  NAND U1528 ( .A(N113), .B(xregN_1), .Z(n1020) );
  NAND U1529 ( .A(n1022), .B(n1023), .Z(z2[108]) );
  NANDN U1530 ( .A(xregN_1), .B(zin[107]), .Z(n1023) );
  NAND U1531 ( .A(N112), .B(xregN_1), .Z(n1022) );
  NAND U1532 ( .A(n1024), .B(n1025), .Z(z2[107]) );
  NANDN U1533 ( .A(xregN_1), .B(zin[106]), .Z(n1025) );
  NAND U1534 ( .A(N111), .B(xregN_1), .Z(n1024) );
  NAND U1535 ( .A(n1026), .B(n1027), .Z(z2[106]) );
  NANDN U1536 ( .A(xregN_1), .B(zin[105]), .Z(n1027) );
  NAND U1537 ( .A(N110), .B(xregN_1), .Z(n1026) );
  NAND U1538 ( .A(n1028), .B(n1029), .Z(z2[105]) );
  NANDN U1539 ( .A(xregN_1), .B(zin[104]), .Z(n1029) );
  NAND U1540 ( .A(N109), .B(xregN_1), .Z(n1028) );
  NAND U1541 ( .A(n1030), .B(n1031), .Z(z2[104]) );
  NANDN U1542 ( .A(xregN_1), .B(zin[103]), .Z(n1031) );
  NAND U1543 ( .A(N108), .B(xregN_1), .Z(n1030) );
  NAND U1544 ( .A(n1032), .B(n1033), .Z(z2[103]) );
  NANDN U1545 ( .A(xregN_1), .B(zin[102]), .Z(n1033) );
  NAND U1546 ( .A(N107), .B(xregN_1), .Z(n1032) );
  NAND U1547 ( .A(n1034), .B(n1035), .Z(z2[102]) );
  NANDN U1548 ( .A(xregN_1), .B(zin[101]), .Z(n1035) );
  NAND U1549 ( .A(N106), .B(xregN_1), .Z(n1034) );
  NAND U1550 ( .A(n1036), .B(n1037), .Z(z2[101]) );
  NANDN U1551 ( .A(xregN_1), .B(zin[100]), .Z(n1037) );
  NAND U1552 ( .A(N105), .B(xregN_1), .Z(n1036) );
  NAND U1553 ( .A(n1038), .B(n1039), .Z(z2[100]) );
  NANDN U1554 ( .A(xregN_1), .B(zin[99]), .Z(n1039) );
  NAND U1555 ( .A(N104), .B(xregN_1), .Z(n1038) );
  AND U1556 ( .A(N4), .B(xregN_1), .Z(z2[0]) );
endmodule


module modmult_step_N256_4_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279;

  IV U1 ( .A(n1278), .Z(n1) );
  IV U2 ( .A(A[1]), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(DIFF[9]) );
  XOR U4 ( .A(B[9]), .B(A[9]), .Z(n4) );
  XNOR U5 ( .A(n5), .B(n6), .Z(DIFF[99]) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(DIFF[98]) );
  XOR U8 ( .A(B[98]), .B(A[98]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(DIFF[97]) );
  XOR U10 ( .A(B[97]), .B(A[97]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(DIFF[96]) );
  XOR U12 ( .A(B[96]), .B(A[96]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(DIFF[95]) );
  XOR U14 ( .A(B[95]), .B(A[95]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(DIFF[94]) );
  XOR U16 ( .A(B[94]), .B(A[94]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(DIFF[93]) );
  XOR U18 ( .A(B[93]), .B(A[93]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(DIFF[92]) );
  XOR U20 ( .A(B[92]), .B(A[92]), .Z(n20) );
  XOR U21 ( .A(n21), .B(n22), .Z(DIFF[91]) );
  XOR U22 ( .A(B[91]), .B(A[91]), .Z(n22) );
  XOR U23 ( .A(n23), .B(n24), .Z(DIFF[90]) );
  XOR U24 ( .A(B[90]), .B(A[90]), .Z(n24) );
  XOR U25 ( .A(n25), .B(n26), .Z(DIFF[8]) );
  XOR U26 ( .A(B[8]), .B(A[8]), .Z(n26) );
  XOR U27 ( .A(n27), .B(n28), .Z(DIFF[89]) );
  XOR U28 ( .A(B[89]), .B(A[89]), .Z(n28) );
  XOR U29 ( .A(n29), .B(n30), .Z(DIFF[88]) );
  XOR U30 ( .A(B[88]), .B(A[88]), .Z(n30) );
  XOR U31 ( .A(n31), .B(n32), .Z(DIFF[87]) );
  XOR U32 ( .A(B[87]), .B(A[87]), .Z(n32) );
  XOR U33 ( .A(n33), .B(n34), .Z(DIFF[86]) );
  XOR U34 ( .A(B[86]), .B(A[86]), .Z(n34) );
  XOR U35 ( .A(n35), .B(n36), .Z(DIFF[85]) );
  XOR U36 ( .A(B[85]), .B(A[85]), .Z(n36) );
  XOR U37 ( .A(n37), .B(n38), .Z(DIFF[84]) );
  XOR U38 ( .A(B[84]), .B(A[84]), .Z(n38) );
  XOR U39 ( .A(n39), .B(n40), .Z(DIFF[83]) );
  XOR U40 ( .A(B[83]), .B(A[83]), .Z(n40) );
  XOR U41 ( .A(n41), .B(n42), .Z(DIFF[82]) );
  XOR U42 ( .A(B[82]), .B(A[82]), .Z(n42) );
  XOR U43 ( .A(n43), .B(n44), .Z(DIFF[81]) );
  XOR U44 ( .A(B[81]), .B(A[81]), .Z(n44) );
  XOR U45 ( .A(n45), .B(n46), .Z(DIFF[80]) );
  XOR U46 ( .A(B[80]), .B(A[80]), .Z(n46) );
  XOR U47 ( .A(n47), .B(n48), .Z(DIFF[7]) );
  XOR U48 ( .A(B[7]), .B(A[7]), .Z(n48) );
  XOR U49 ( .A(n49), .B(n50), .Z(DIFF[79]) );
  XOR U50 ( .A(B[79]), .B(A[79]), .Z(n50) );
  XOR U51 ( .A(n51), .B(n52), .Z(DIFF[78]) );
  XOR U52 ( .A(B[78]), .B(A[78]), .Z(n52) );
  XOR U53 ( .A(n53), .B(n54), .Z(DIFF[77]) );
  XOR U54 ( .A(B[77]), .B(A[77]), .Z(n54) );
  XOR U55 ( .A(n55), .B(n56), .Z(DIFF[76]) );
  XOR U56 ( .A(B[76]), .B(A[76]), .Z(n56) );
  XOR U57 ( .A(n57), .B(n58), .Z(DIFF[75]) );
  XOR U58 ( .A(B[75]), .B(A[75]), .Z(n58) );
  XOR U59 ( .A(n59), .B(n60), .Z(DIFF[74]) );
  XOR U60 ( .A(B[74]), .B(A[74]), .Z(n60) );
  XOR U61 ( .A(n61), .B(n62), .Z(DIFF[73]) );
  XOR U62 ( .A(B[73]), .B(A[73]), .Z(n62) );
  XOR U63 ( .A(n63), .B(n64), .Z(DIFF[72]) );
  XOR U64 ( .A(B[72]), .B(A[72]), .Z(n64) );
  XOR U65 ( .A(n65), .B(n66), .Z(DIFF[71]) );
  XOR U66 ( .A(B[71]), .B(A[71]), .Z(n66) );
  XOR U67 ( .A(n67), .B(n68), .Z(DIFF[70]) );
  XOR U68 ( .A(B[70]), .B(A[70]), .Z(n68) );
  XOR U69 ( .A(n69), .B(n70), .Z(DIFF[6]) );
  XOR U70 ( .A(B[6]), .B(A[6]), .Z(n70) );
  XOR U71 ( .A(n71), .B(n72), .Z(DIFF[69]) );
  XOR U72 ( .A(B[69]), .B(A[69]), .Z(n72) );
  XOR U73 ( .A(n73), .B(n74), .Z(DIFF[68]) );
  XOR U74 ( .A(B[68]), .B(A[68]), .Z(n74) );
  XOR U75 ( .A(n75), .B(n76), .Z(DIFF[67]) );
  XOR U76 ( .A(B[67]), .B(A[67]), .Z(n76) );
  XOR U77 ( .A(n77), .B(n78), .Z(DIFF[66]) );
  XOR U78 ( .A(B[66]), .B(A[66]), .Z(n78) );
  XOR U79 ( .A(n79), .B(n80), .Z(DIFF[65]) );
  XOR U80 ( .A(B[65]), .B(A[65]), .Z(n80) );
  XOR U81 ( .A(n81), .B(n82), .Z(DIFF[64]) );
  XOR U82 ( .A(B[64]), .B(A[64]), .Z(n82) );
  XOR U83 ( .A(n83), .B(n84), .Z(DIFF[63]) );
  XOR U84 ( .A(B[63]), .B(A[63]), .Z(n84) );
  XOR U85 ( .A(n85), .B(n86), .Z(DIFF[62]) );
  XOR U86 ( .A(B[62]), .B(A[62]), .Z(n86) );
  XOR U87 ( .A(n87), .B(n88), .Z(DIFF[61]) );
  XOR U88 ( .A(B[61]), .B(A[61]), .Z(n88) );
  XOR U89 ( .A(n89), .B(n90), .Z(DIFF[60]) );
  XOR U90 ( .A(B[60]), .B(A[60]), .Z(n90) );
  XOR U91 ( .A(n91), .B(n92), .Z(DIFF[5]) );
  XOR U92 ( .A(B[5]), .B(A[5]), .Z(n92) );
  XOR U93 ( .A(n93), .B(n94), .Z(DIFF[59]) );
  XOR U94 ( .A(B[59]), .B(A[59]), .Z(n94) );
  XOR U95 ( .A(n95), .B(n96), .Z(DIFF[58]) );
  XOR U96 ( .A(B[58]), .B(A[58]), .Z(n96) );
  XOR U97 ( .A(n97), .B(n98), .Z(DIFF[57]) );
  XOR U98 ( .A(B[57]), .B(A[57]), .Z(n98) );
  XOR U99 ( .A(n99), .B(n100), .Z(DIFF[56]) );
  XOR U100 ( .A(B[56]), .B(A[56]), .Z(n100) );
  XOR U101 ( .A(n101), .B(n102), .Z(DIFF[55]) );
  XOR U102 ( .A(B[55]), .B(A[55]), .Z(n102) );
  XOR U103 ( .A(n103), .B(n104), .Z(DIFF[54]) );
  XOR U104 ( .A(B[54]), .B(A[54]), .Z(n104) );
  XOR U105 ( .A(n105), .B(n106), .Z(DIFF[53]) );
  XOR U106 ( .A(B[53]), .B(A[53]), .Z(n106) );
  XOR U107 ( .A(n107), .B(n108), .Z(DIFF[52]) );
  XOR U108 ( .A(B[52]), .B(A[52]), .Z(n108) );
  XOR U109 ( .A(n109), .B(n110), .Z(DIFF[51]) );
  XOR U110 ( .A(B[51]), .B(A[51]), .Z(n110) );
  XOR U111 ( .A(n111), .B(n112), .Z(DIFF[50]) );
  XOR U112 ( .A(B[50]), .B(A[50]), .Z(n112) );
  XOR U113 ( .A(n113), .B(n114), .Z(DIFF[4]) );
  XOR U114 ( .A(B[4]), .B(A[4]), .Z(n114) );
  XOR U115 ( .A(n115), .B(n116), .Z(DIFF[49]) );
  XOR U116 ( .A(B[49]), .B(A[49]), .Z(n116) );
  XOR U117 ( .A(n117), .B(n118), .Z(DIFF[48]) );
  XOR U118 ( .A(B[48]), .B(A[48]), .Z(n118) );
  XOR U119 ( .A(n119), .B(n120), .Z(DIFF[47]) );
  XOR U120 ( .A(B[47]), .B(A[47]), .Z(n120) );
  XOR U121 ( .A(n121), .B(n122), .Z(DIFF[46]) );
  XOR U122 ( .A(B[46]), .B(A[46]), .Z(n122) );
  XOR U123 ( .A(n123), .B(n124), .Z(DIFF[45]) );
  XOR U124 ( .A(B[45]), .B(A[45]), .Z(n124) );
  XOR U125 ( .A(n125), .B(n126), .Z(DIFF[44]) );
  XOR U126 ( .A(B[44]), .B(A[44]), .Z(n126) );
  XOR U127 ( .A(n127), .B(n128), .Z(DIFF[43]) );
  XOR U128 ( .A(B[43]), .B(A[43]), .Z(n128) );
  XOR U129 ( .A(n129), .B(n130), .Z(DIFF[42]) );
  XOR U130 ( .A(B[42]), .B(A[42]), .Z(n130) );
  XOR U131 ( .A(n131), .B(n132), .Z(DIFF[41]) );
  XOR U132 ( .A(B[41]), .B(A[41]), .Z(n132) );
  XOR U133 ( .A(n133), .B(n134), .Z(DIFF[40]) );
  XOR U134 ( .A(B[40]), .B(A[40]), .Z(n134) );
  XOR U135 ( .A(n135), .B(n136), .Z(DIFF[3]) );
  XOR U136 ( .A(B[3]), .B(A[3]), .Z(n136) );
  XOR U137 ( .A(n137), .B(n138), .Z(DIFF[39]) );
  XOR U138 ( .A(B[39]), .B(A[39]), .Z(n138) );
  XOR U139 ( .A(n139), .B(n140), .Z(DIFF[38]) );
  XOR U140 ( .A(B[38]), .B(A[38]), .Z(n140) );
  XOR U141 ( .A(n141), .B(n142), .Z(DIFF[37]) );
  XOR U142 ( .A(B[37]), .B(A[37]), .Z(n142) );
  XOR U143 ( .A(n143), .B(n144), .Z(DIFF[36]) );
  XOR U144 ( .A(B[36]), .B(A[36]), .Z(n144) );
  XOR U145 ( .A(n145), .B(n146), .Z(DIFF[35]) );
  XOR U146 ( .A(B[35]), .B(A[35]), .Z(n146) );
  XOR U147 ( .A(n147), .B(n148), .Z(DIFF[34]) );
  XOR U148 ( .A(B[34]), .B(A[34]), .Z(n148) );
  XOR U149 ( .A(n149), .B(n150), .Z(DIFF[33]) );
  XOR U150 ( .A(B[33]), .B(A[33]), .Z(n150) );
  XOR U151 ( .A(n151), .B(n152), .Z(DIFF[32]) );
  XOR U152 ( .A(B[32]), .B(A[32]), .Z(n152) );
  XOR U153 ( .A(n153), .B(n154), .Z(DIFF[31]) );
  XOR U154 ( .A(B[31]), .B(A[31]), .Z(n154) );
  XOR U155 ( .A(n155), .B(n156), .Z(DIFF[30]) );
  XOR U156 ( .A(B[30]), .B(A[30]), .Z(n156) );
  XOR U157 ( .A(n157), .B(n158), .Z(DIFF[2]) );
  XOR U158 ( .A(B[2]), .B(A[2]), .Z(n158) );
  XOR U159 ( .A(n159), .B(n160), .Z(DIFF[29]) );
  XOR U160 ( .A(B[29]), .B(A[29]), .Z(n160) );
  XOR U161 ( .A(n161), .B(n162), .Z(DIFF[28]) );
  XOR U162 ( .A(B[28]), .B(A[28]), .Z(n162) );
  XOR U163 ( .A(n163), .B(n164), .Z(DIFF[27]) );
  XOR U164 ( .A(B[27]), .B(A[27]), .Z(n164) );
  XOR U165 ( .A(n165), .B(n166), .Z(DIFF[26]) );
  XOR U166 ( .A(B[26]), .B(A[26]), .Z(n166) );
  XOR U167 ( .A(n167), .B(n168), .Z(DIFF[25]) );
  XOR U168 ( .A(B[25]), .B(A[25]), .Z(n168) );
  XOR U169 ( .A(A[256]), .B(n169), .Z(DIFF[256]) );
  AND U170 ( .A(n170), .B(n171), .Z(n169) );
  NANDN U171 ( .A(B[255]), .B(n172), .Z(n171) );
  NANDN U172 ( .A(A[255]), .B(n173), .Z(n172) );
  NANDN U173 ( .A(n173), .B(A[255]), .Z(n170) );
  XOR U174 ( .A(n173), .B(n174), .Z(DIFF[255]) );
  XOR U175 ( .A(B[255]), .B(A[255]), .Z(n174) );
  AND U176 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U177 ( .A(B[254]), .B(n177), .Z(n176) );
  NANDN U178 ( .A(A[254]), .B(n178), .Z(n177) );
  NANDN U179 ( .A(n178), .B(A[254]), .Z(n175) );
  XOR U180 ( .A(n178), .B(n179), .Z(DIFF[254]) );
  XOR U181 ( .A(B[254]), .B(A[254]), .Z(n179) );
  AND U182 ( .A(n180), .B(n181), .Z(n178) );
  NANDN U183 ( .A(B[253]), .B(n182), .Z(n181) );
  NANDN U184 ( .A(A[253]), .B(n183), .Z(n182) );
  NANDN U185 ( .A(n183), .B(A[253]), .Z(n180) );
  XOR U186 ( .A(n183), .B(n184), .Z(DIFF[253]) );
  XOR U187 ( .A(B[253]), .B(A[253]), .Z(n184) );
  AND U188 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U189 ( .A(B[252]), .B(n187), .Z(n186) );
  NANDN U190 ( .A(A[252]), .B(n188), .Z(n187) );
  NANDN U191 ( .A(n188), .B(A[252]), .Z(n185) );
  XOR U192 ( .A(n188), .B(n189), .Z(DIFF[252]) );
  XOR U193 ( .A(B[252]), .B(A[252]), .Z(n189) );
  AND U194 ( .A(n190), .B(n191), .Z(n188) );
  NANDN U195 ( .A(B[251]), .B(n192), .Z(n191) );
  NANDN U196 ( .A(A[251]), .B(n193), .Z(n192) );
  NANDN U197 ( .A(n193), .B(A[251]), .Z(n190) );
  XOR U198 ( .A(n193), .B(n194), .Z(DIFF[251]) );
  XOR U199 ( .A(B[251]), .B(A[251]), .Z(n194) );
  AND U200 ( .A(n195), .B(n196), .Z(n193) );
  NANDN U201 ( .A(B[250]), .B(n197), .Z(n196) );
  NANDN U202 ( .A(A[250]), .B(n198), .Z(n197) );
  NANDN U203 ( .A(n198), .B(A[250]), .Z(n195) );
  XOR U204 ( .A(n198), .B(n199), .Z(DIFF[250]) );
  XOR U205 ( .A(B[250]), .B(A[250]), .Z(n199) );
  AND U206 ( .A(n200), .B(n201), .Z(n198) );
  NANDN U207 ( .A(B[249]), .B(n202), .Z(n201) );
  NANDN U208 ( .A(A[249]), .B(n203), .Z(n202) );
  NANDN U209 ( .A(n203), .B(A[249]), .Z(n200) );
  XOR U210 ( .A(n204), .B(n205), .Z(DIFF[24]) );
  XOR U211 ( .A(B[24]), .B(A[24]), .Z(n205) );
  XOR U212 ( .A(n203), .B(n206), .Z(DIFF[249]) );
  XOR U213 ( .A(B[249]), .B(A[249]), .Z(n206) );
  AND U214 ( .A(n207), .B(n208), .Z(n203) );
  NANDN U215 ( .A(B[248]), .B(n209), .Z(n208) );
  NANDN U216 ( .A(A[248]), .B(n210), .Z(n209) );
  NANDN U217 ( .A(n210), .B(A[248]), .Z(n207) );
  XOR U218 ( .A(n210), .B(n211), .Z(DIFF[248]) );
  XOR U219 ( .A(B[248]), .B(A[248]), .Z(n211) );
  AND U220 ( .A(n212), .B(n213), .Z(n210) );
  NANDN U221 ( .A(B[247]), .B(n214), .Z(n213) );
  NANDN U222 ( .A(A[247]), .B(n215), .Z(n214) );
  NANDN U223 ( .A(n215), .B(A[247]), .Z(n212) );
  XOR U224 ( .A(n215), .B(n216), .Z(DIFF[247]) );
  XOR U225 ( .A(B[247]), .B(A[247]), .Z(n216) );
  AND U226 ( .A(n217), .B(n218), .Z(n215) );
  NANDN U227 ( .A(B[246]), .B(n219), .Z(n218) );
  NANDN U228 ( .A(A[246]), .B(n220), .Z(n219) );
  NANDN U229 ( .A(n220), .B(A[246]), .Z(n217) );
  XOR U230 ( .A(n220), .B(n221), .Z(DIFF[246]) );
  XOR U231 ( .A(B[246]), .B(A[246]), .Z(n221) );
  AND U232 ( .A(n222), .B(n223), .Z(n220) );
  NANDN U233 ( .A(B[245]), .B(n224), .Z(n223) );
  NANDN U234 ( .A(A[245]), .B(n225), .Z(n224) );
  NANDN U235 ( .A(n225), .B(A[245]), .Z(n222) );
  XOR U236 ( .A(n225), .B(n226), .Z(DIFF[245]) );
  XOR U237 ( .A(B[245]), .B(A[245]), .Z(n226) );
  AND U238 ( .A(n227), .B(n228), .Z(n225) );
  NANDN U239 ( .A(B[244]), .B(n229), .Z(n228) );
  NANDN U240 ( .A(A[244]), .B(n230), .Z(n229) );
  NANDN U241 ( .A(n230), .B(A[244]), .Z(n227) );
  XOR U242 ( .A(n230), .B(n231), .Z(DIFF[244]) );
  XOR U243 ( .A(B[244]), .B(A[244]), .Z(n231) );
  AND U244 ( .A(n232), .B(n233), .Z(n230) );
  NANDN U245 ( .A(B[243]), .B(n234), .Z(n233) );
  NANDN U246 ( .A(A[243]), .B(n235), .Z(n234) );
  NANDN U247 ( .A(n235), .B(A[243]), .Z(n232) );
  XOR U248 ( .A(n235), .B(n236), .Z(DIFF[243]) );
  XOR U249 ( .A(B[243]), .B(A[243]), .Z(n236) );
  AND U250 ( .A(n237), .B(n238), .Z(n235) );
  NANDN U251 ( .A(B[242]), .B(n239), .Z(n238) );
  NANDN U252 ( .A(A[242]), .B(n240), .Z(n239) );
  NANDN U253 ( .A(n240), .B(A[242]), .Z(n237) );
  XOR U254 ( .A(n240), .B(n241), .Z(DIFF[242]) );
  XOR U255 ( .A(B[242]), .B(A[242]), .Z(n241) );
  AND U256 ( .A(n242), .B(n243), .Z(n240) );
  NANDN U257 ( .A(B[241]), .B(n244), .Z(n243) );
  NANDN U258 ( .A(A[241]), .B(n245), .Z(n244) );
  NANDN U259 ( .A(n245), .B(A[241]), .Z(n242) );
  XOR U260 ( .A(n245), .B(n246), .Z(DIFF[241]) );
  XOR U261 ( .A(B[241]), .B(A[241]), .Z(n246) );
  AND U262 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U263 ( .A(B[240]), .B(n249), .Z(n248) );
  NANDN U264 ( .A(A[240]), .B(n250), .Z(n249) );
  NANDN U265 ( .A(n250), .B(A[240]), .Z(n247) );
  XOR U266 ( .A(n250), .B(n251), .Z(DIFF[240]) );
  XOR U267 ( .A(B[240]), .B(A[240]), .Z(n251) );
  AND U268 ( .A(n252), .B(n253), .Z(n250) );
  NANDN U269 ( .A(B[239]), .B(n254), .Z(n253) );
  NANDN U270 ( .A(A[239]), .B(n255), .Z(n254) );
  NANDN U271 ( .A(n255), .B(A[239]), .Z(n252) );
  XOR U272 ( .A(n256), .B(n257), .Z(DIFF[23]) );
  XOR U273 ( .A(B[23]), .B(A[23]), .Z(n257) );
  XOR U274 ( .A(n255), .B(n258), .Z(DIFF[239]) );
  XOR U275 ( .A(B[239]), .B(A[239]), .Z(n258) );
  AND U276 ( .A(n259), .B(n260), .Z(n255) );
  NANDN U277 ( .A(B[238]), .B(n261), .Z(n260) );
  NANDN U278 ( .A(A[238]), .B(n262), .Z(n261) );
  NANDN U279 ( .A(n262), .B(A[238]), .Z(n259) );
  XOR U280 ( .A(n262), .B(n263), .Z(DIFF[238]) );
  XOR U281 ( .A(B[238]), .B(A[238]), .Z(n263) );
  AND U282 ( .A(n264), .B(n265), .Z(n262) );
  NANDN U283 ( .A(B[237]), .B(n266), .Z(n265) );
  NANDN U284 ( .A(A[237]), .B(n267), .Z(n266) );
  NANDN U285 ( .A(n267), .B(A[237]), .Z(n264) );
  XOR U286 ( .A(n267), .B(n268), .Z(DIFF[237]) );
  XOR U287 ( .A(B[237]), .B(A[237]), .Z(n268) );
  AND U288 ( .A(n269), .B(n270), .Z(n267) );
  NANDN U289 ( .A(B[236]), .B(n271), .Z(n270) );
  NANDN U290 ( .A(A[236]), .B(n272), .Z(n271) );
  NANDN U291 ( .A(n272), .B(A[236]), .Z(n269) );
  XOR U292 ( .A(n272), .B(n273), .Z(DIFF[236]) );
  XOR U293 ( .A(B[236]), .B(A[236]), .Z(n273) );
  AND U294 ( .A(n274), .B(n275), .Z(n272) );
  NANDN U295 ( .A(B[235]), .B(n276), .Z(n275) );
  NANDN U296 ( .A(A[235]), .B(n277), .Z(n276) );
  NANDN U297 ( .A(n277), .B(A[235]), .Z(n274) );
  XOR U298 ( .A(n277), .B(n278), .Z(DIFF[235]) );
  XOR U299 ( .A(B[235]), .B(A[235]), .Z(n278) );
  AND U300 ( .A(n279), .B(n280), .Z(n277) );
  NANDN U301 ( .A(B[234]), .B(n281), .Z(n280) );
  NANDN U302 ( .A(A[234]), .B(n282), .Z(n281) );
  NANDN U303 ( .A(n282), .B(A[234]), .Z(n279) );
  XOR U304 ( .A(n282), .B(n283), .Z(DIFF[234]) );
  XOR U305 ( .A(B[234]), .B(A[234]), .Z(n283) );
  AND U306 ( .A(n284), .B(n285), .Z(n282) );
  NANDN U307 ( .A(B[233]), .B(n286), .Z(n285) );
  NANDN U308 ( .A(A[233]), .B(n287), .Z(n286) );
  NANDN U309 ( .A(n287), .B(A[233]), .Z(n284) );
  XOR U310 ( .A(n287), .B(n288), .Z(DIFF[233]) );
  XOR U311 ( .A(B[233]), .B(A[233]), .Z(n288) );
  AND U312 ( .A(n289), .B(n290), .Z(n287) );
  NANDN U313 ( .A(B[232]), .B(n291), .Z(n290) );
  NANDN U314 ( .A(A[232]), .B(n292), .Z(n291) );
  NANDN U315 ( .A(n292), .B(A[232]), .Z(n289) );
  XOR U316 ( .A(n292), .B(n293), .Z(DIFF[232]) );
  XOR U317 ( .A(B[232]), .B(A[232]), .Z(n293) );
  AND U318 ( .A(n294), .B(n295), .Z(n292) );
  NANDN U319 ( .A(B[231]), .B(n296), .Z(n295) );
  NANDN U320 ( .A(A[231]), .B(n297), .Z(n296) );
  NANDN U321 ( .A(n297), .B(A[231]), .Z(n294) );
  XOR U322 ( .A(n297), .B(n298), .Z(DIFF[231]) );
  XOR U323 ( .A(B[231]), .B(A[231]), .Z(n298) );
  AND U324 ( .A(n299), .B(n300), .Z(n297) );
  NANDN U325 ( .A(B[230]), .B(n301), .Z(n300) );
  NANDN U326 ( .A(A[230]), .B(n302), .Z(n301) );
  NANDN U327 ( .A(n302), .B(A[230]), .Z(n299) );
  XOR U328 ( .A(n302), .B(n303), .Z(DIFF[230]) );
  XOR U329 ( .A(B[230]), .B(A[230]), .Z(n303) );
  AND U330 ( .A(n304), .B(n305), .Z(n302) );
  NANDN U331 ( .A(B[229]), .B(n306), .Z(n305) );
  NANDN U332 ( .A(A[229]), .B(n307), .Z(n306) );
  NANDN U333 ( .A(n307), .B(A[229]), .Z(n304) );
  XOR U334 ( .A(n308), .B(n309), .Z(DIFF[22]) );
  XOR U335 ( .A(B[22]), .B(A[22]), .Z(n309) );
  XOR U336 ( .A(n307), .B(n310), .Z(DIFF[229]) );
  XOR U337 ( .A(B[229]), .B(A[229]), .Z(n310) );
  AND U338 ( .A(n311), .B(n312), .Z(n307) );
  NANDN U339 ( .A(B[228]), .B(n313), .Z(n312) );
  NANDN U340 ( .A(A[228]), .B(n314), .Z(n313) );
  NANDN U341 ( .A(n314), .B(A[228]), .Z(n311) );
  XOR U342 ( .A(n314), .B(n315), .Z(DIFF[228]) );
  XOR U343 ( .A(B[228]), .B(A[228]), .Z(n315) );
  AND U344 ( .A(n316), .B(n317), .Z(n314) );
  NANDN U345 ( .A(B[227]), .B(n318), .Z(n317) );
  NANDN U346 ( .A(A[227]), .B(n319), .Z(n318) );
  NANDN U347 ( .A(n319), .B(A[227]), .Z(n316) );
  XOR U348 ( .A(n319), .B(n320), .Z(DIFF[227]) );
  XOR U349 ( .A(B[227]), .B(A[227]), .Z(n320) );
  AND U350 ( .A(n321), .B(n322), .Z(n319) );
  NANDN U351 ( .A(B[226]), .B(n323), .Z(n322) );
  NANDN U352 ( .A(A[226]), .B(n324), .Z(n323) );
  NANDN U353 ( .A(n324), .B(A[226]), .Z(n321) );
  XOR U354 ( .A(n324), .B(n325), .Z(DIFF[226]) );
  XOR U355 ( .A(B[226]), .B(A[226]), .Z(n325) );
  AND U356 ( .A(n326), .B(n327), .Z(n324) );
  NANDN U357 ( .A(B[225]), .B(n328), .Z(n327) );
  NANDN U358 ( .A(A[225]), .B(n329), .Z(n328) );
  NANDN U359 ( .A(n329), .B(A[225]), .Z(n326) );
  XOR U360 ( .A(n329), .B(n330), .Z(DIFF[225]) );
  XOR U361 ( .A(B[225]), .B(A[225]), .Z(n330) );
  AND U362 ( .A(n331), .B(n332), .Z(n329) );
  NANDN U363 ( .A(B[224]), .B(n333), .Z(n332) );
  NANDN U364 ( .A(A[224]), .B(n334), .Z(n333) );
  NANDN U365 ( .A(n334), .B(A[224]), .Z(n331) );
  XOR U366 ( .A(n334), .B(n335), .Z(DIFF[224]) );
  XOR U367 ( .A(B[224]), .B(A[224]), .Z(n335) );
  AND U368 ( .A(n336), .B(n337), .Z(n334) );
  NANDN U369 ( .A(B[223]), .B(n338), .Z(n337) );
  NANDN U370 ( .A(A[223]), .B(n339), .Z(n338) );
  NANDN U371 ( .A(n339), .B(A[223]), .Z(n336) );
  XOR U372 ( .A(n339), .B(n340), .Z(DIFF[223]) );
  XOR U373 ( .A(B[223]), .B(A[223]), .Z(n340) );
  AND U374 ( .A(n341), .B(n342), .Z(n339) );
  NANDN U375 ( .A(B[222]), .B(n343), .Z(n342) );
  NANDN U376 ( .A(A[222]), .B(n344), .Z(n343) );
  NANDN U377 ( .A(n344), .B(A[222]), .Z(n341) );
  XOR U378 ( .A(n344), .B(n345), .Z(DIFF[222]) );
  XOR U379 ( .A(B[222]), .B(A[222]), .Z(n345) );
  AND U380 ( .A(n346), .B(n347), .Z(n344) );
  NANDN U381 ( .A(B[221]), .B(n348), .Z(n347) );
  NANDN U382 ( .A(A[221]), .B(n349), .Z(n348) );
  NANDN U383 ( .A(n349), .B(A[221]), .Z(n346) );
  XOR U384 ( .A(n349), .B(n350), .Z(DIFF[221]) );
  XOR U385 ( .A(B[221]), .B(A[221]), .Z(n350) );
  AND U386 ( .A(n351), .B(n352), .Z(n349) );
  NANDN U387 ( .A(B[220]), .B(n353), .Z(n352) );
  NANDN U388 ( .A(A[220]), .B(n354), .Z(n353) );
  NANDN U389 ( .A(n354), .B(A[220]), .Z(n351) );
  XOR U390 ( .A(n354), .B(n355), .Z(DIFF[220]) );
  XOR U391 ( .A(B[220]), .B(A[220]), .Z(n355) );
  AND U392 ( .A(n356), .B(n357), .Z(n354) );
  NANDN U393 ( .A(B[219]), .B(n358), .Z(n357) );
  NANDN U394 ( .A(A[219]), .B(n359), .Z(n358) );
  NANDN U395 ( .A(n359), .B(A[219]), .Z(n356) );
  XOR U396 ( .A(n360), .B(n361), .Z(DIFF[21]) );
  XOR U397 ( .A(B[21]), .B(A[21]), .Z(n361) );
  XOR U398 ( .A(n359), .B(n362), .Z(DIFF[219]) );
  XOR U399 ( .A(B[219]), .B(A[219]), .Z(n362) );
  AND U400 ( .A(n363), .B(n364), .Z(n359) );
  NANDN U401 ( .A(B[218]), .B(n365), .Z(n364) );
  NANDN U402 ( .A(A[218]), .B(n366), .Z(n365) );
  NANDN U403 ( .A(n366), .B(A[218]), .Z(n363) );
  XOR U404 ( .A(n366), .B(n367), .Z(DIFF[218]) );
  XOR U405 ( .A(B[218]), .B(A[218]), .Z(n367) );
  AND U406 ( .A(n368), .B(n369), .Z(n366) );
  NANDN U407 ( .A(B[217]), .B(n370), .Z(n369) );
  NANDN U408 ( .A(A[217]), .B(n371), .Z(n370) );
  NANDN U409 ( .A(n371), .B(A[217]), .Z(n368) );
  XOR U410 ( .A(n371), .B(n372), .Z(DIFF[217]) );
  XOR U411 ( .A(B[217]), .B(A[217]), .Z(n372) );
  AND U412 ( .A(n373), .B(n374), .Z(n371) );
  NANDN U413 ( .A(B[216]), .B(n375), .Z(n374) );
  NANDN U414 ( .A(A[216]), .B(n376), .Z(n375) );
  NANDN U415 ( .A(n376), .B(A[216]), .Z(n373) );
  XOR U416 ( .A(n376), .B(n377), .Z(DIFF[216]) );
  XOR U417 ( .A(B[216]), .B(A[216]), .Z(n377) );
  AND U418 ( .A(n378), .B(n379), .Z(n376) );
  NANDN U419 ( .A(B[215]), .B(n380), .Z(n379) );
  NANDN U420 ( .A(A[215]), .B(n381), .Z(n380) );
  NANDN U421 ( .A(n381), .B(A[215]), .Z(n378) );
  XOR U422 ( .A(n381), .B(n382), .Z(DIFF[215]) );
  XOR U423 ( .A(B[215]), .B(A[215]), .Z(n382) );
  AND U424 ( .A(n383), .B(n384), .Z(n381) );
  NANDN U425 ( .A(B[214]), .B(n385), .Z(n384) );
  NANDN U426 ( .A(A[214]), .B(n386), .Z(n385) );
  NANDN U427 ( .A(n386), .B(A[214]), .Z(n383) );
  XOR U428 ( .A(n386), .B(n387), .Z(DIFF[214]) );
  XOR U429 ( .A(B[214]), .B(A[214]), .Z(n387) );
  AND U430 ( .A(n388), .B(n389), .Z(n386) );
  NANDN U431 ( .A(B[213]), .B(n390), .Z(n389) );
  NANDN U432 ( .A(A[213]), .B(n391), .Z(n390) );
  NANDN U433 ( .A(n391), .B(A[213]), .Z(n388) );
  XOR U434 ( .A(n391), .B(n392), .Z(DIFF[213]) );
  XOR U435 ( .A(B[213]), .B(A[213]), .Z(n392) );
  AND U436 ( .A(n393), .B(n394), .Z(n391) );
  NANDN U437 ( .A(B[212]), .B(n395), .Z(n394) );
  NANDN U438 ( .A(A[212]), .B(n396), .Z(n395) );
  NANDN U439 ( .A(n396), .B(A[212]), .Z(n393) );
  XOR U440 ( .A(n396), .B(n397), .Z(DIFF[212]) );
  XOR U441 ( .A(B[212]), .B(A[212]), .Z(n397) );
  AND U442 ( .A(n398), .B(n399), .Z(n396) );
  NANDN U443 ( .A(B[211]), .B(n400), .Z(n399) );
  NANDN U444 ( .A(A[211]), .B(n401), .Z(n400) );
  NANDN U445 ( .A(n401), .B(A[211]), .Z(n398) );
  XOR U446 ( .A(n401), .B(n402), .Z(DIFF[211]) );
  XOR U447 ( .A(B[211]), .B(A[211]), .Z(n402) );
  AND U448 ( .A(n403), .B(n404), .Z(n401) );
  NANDN U449 ( .A(B[210]), .B(n405), .Z(n404) );
  NANDN U450 ( .A(A[210]), .B(n406), .Z(n405) );
  NANDN U451 ( .A(n406), .B(A[210]), .Z(n403) );
  XOR U452 ( .A(n406), .B(n407), .Z(DIFF[210]) );
  XOR U453 ( .A(B[210]), .B(A[210]), .Z(n407) );
  AND U454 ( .A(n408), .B(n409), .Z(n406) );
  NANDN U455 ( .A(B[209]), .B(n410), .Z(n409) );
  NANDN U456 ( .A(A[209]), .B(n411), .Z(n410) );
  NANDN U457 ( .A(n411), .B(A[209]), .Z(n408) );
  XOR U458 ( .A(n412), .B(n413), .Z(DIFF[20]) );
  XOR U459 ( .A(B[20]), .B(A[20]), .Z(n413) );
  XOR U460 ( .A(n411), .B(n414), .Z(DIFF[209]) );
  XOR U461 ( .A(B[209]), .B(A[209]), .Z(n414) );
  AND U462 ( .A(n415), .B(n416), .Z(n411) );
  NANDN U463 ( .A(B[208]), .B(n417), .Z(n416) );
  NANDN U464 ( .A(A[208]), .B(n418), .Z(n417) );
  NANDN U465 ( .A(n418), .B(A[208]), .Z(n415) );
  XOR U466 ( .A(n418), .B(n419), .Z(DIFF[208]) );
  XOR U467 ( .A(B[208]), .B(A[208]), .Z(n419) );
  AND U468 ( .A(n420), .B(n421), .Z(n418) );
  NANDN U469 ( .A(B[207]), .B(n422), .Z(n421) );
  NANDN U470 ( .A(A[207]), .B(n423), .Z(n422) );
  NANDN U471 ( .A(n423), .B(A[207]), .Z(n420) );
  XOR U472 ( .A(n423), .B(n424), .Z(DIFF[207]) );
  XOR U473 ( .A(B[207]), .B(A[207]), .Z(n424) );
  AND U474 ( .A(n425), .B(n426), .Z(n423) );
  NANDN U475 ( .A(B[206]), .B(n427), .Z(n426) );
  NANDN U476 ( .A(A[206]), .B(n428), .Z(n427) );
  NANDN U477 ( .A(n428), .B(A[206]), .Z(n425) );
  XOR U478 ( .A(n428), .B(n429), .Z(DIFF[206]) );
  XOR U479 ( .A(B[206]), .B(A[206]), .Z(n429) );
  AND U480 ( .A(n430), .B(n431), .Z(n428) );
  NANDN U481 ( .A(B[205]), .B(n432), .Z(n431) );
  NANDN U482 ( .A(A[205]), .B(n433), .Z(n432) );
  NANDN U483 ( .A(n433), .B(A[205]), .Z(n430) );
  XOR U484 ( .A(n433), .B(n434), .Z(DIFF[205]) );
  XOR U485 ( .A(B[205]), .B(A[205]), .Z(n434) );
  AND U486 ( .A(n435), .B(n436), .Z(n433) );
  NANDN U487 ( .A(B[204]), .B(n437), .Z(n436) );
  NANDN U488 ( .A(A[204]), .B(n438), .Z(n437) );
  NANDN U489 ( .A(n438), .B(A[204]), .Z(n435) );
  XOR U490 ( .A(n438), .B(n439), .Z(DIFF[204]) );
  XOR U491 ( .A(B[204]), .B(A[204]), .Z(n439) );
  AND U492 ( .A(n440), .B(n441), .Z(n438) );
  NANDN U493 ( .A(B[203]), .B(n442), .Z(n441) );
  NANDN U494 ( .A(A[203]), .B(n443), .Z(n442) );
  NANDN U495 ( .A(n443), .B(A[203]), .Z(n440) );
  XOR U496 ( .A(n443), .B(n444), .Z(DIFF[203]) );
  XOR U497 ( .A(B[203]), .B(A[203]), .Z(n444) );
  AND U498 ( .A(n445), .B(n446), .Z(n443) );
  NANDN U499 ( .A(B[202]), .B(n447), .Z(n446) );
  NANDN U500 ( .A(A[202]), .B(n448), .Z(n447) );
  NANDN U501 ( .A(n448), .B(A[202]), .Z(n445) );
  XOR U502 ( .A(n448), .B(n449), .Z(DIFF[202]) );
  XOR U503 ( .A(B[202]), .B(A[202]), .Z(n449) );
  AND U504 ( .A(n450), .B(n451), .Z(n448) );
  NANDN U505 ( .A(B[201]), .B(n452), .Z(n451) );
  NANDN U506 ( .A(A[201]), .B(n453), .Z(n452) );
  NANDN U507 ( .A(n453), .B(A[201]), .Z(n450) );
  XOR U508 ( .A(n453), .B(n454), .Z(DIFF[201]) );
  XOR U509 ( .A(B[201]), .B(A[201]), .Z(n454) );
  AND U510 ( .A(n455), .B(n456), .Z(n453) );
  NANDN U511 ( .A(B[200]), .B(n457), .Z(n456) );
  NANDN U512 ( .A(A[200]), .B(n458), .Z(n457) );
  NANDN U513 ( .A(n458), .B(A[200]), .Z(n455) );
  XOR U514 ( .A(n458), .B(n459), .Z(DIFF[200]) );
  XOR U515 ( .A(B[200]), .B(A[200]), .Z(n459) );
  AND U516 ( .A(n460), .B(n461), .Z(n458) );
  NANDN U517 ( .A(B[199]), .B(n462), .Z(n461) );
  NANDN U518 ( .A(A[199]), .B(n463), .Z(n462) );
  NANDN U519 ( .A(n463), .B(A[199]), .Z(n460) );
  XOR U520 ( .A(n1), .B(n464), .Z(DIFF[1]) );
  XOR U521 ( .A(B[1]), .B(A[1]), .Z(n464) );
  XOR U522 ( .A(n465), .B(n466), .Z(DIFF[19]) );
  XOR U523 ( .A(B[19]), .B(A[19]), .Z(n466) );
  XOR U524 ( .A(n463), .B(n467), .Z(DIFF[199]) );
  XOR U525 ( .A(B[199]), .B(A[199]), .Z(n467) );
  AND U526 ( .A(n468), .B(n469), .Z(n463) );
  NANDN U527 ( .A(B[198]), .B(n470), .Z(n469) );
  NANDN U528 ( .A(A[198]), .B(n471), .Z(n470) );
  NANDN U529 ( .A(n471), .B(A[198]), .Z(n468) );
  XOR U530 ( .A(n471), .B(n472), .Z(DIFF[198]) );
  XOR U531 ( .A(B[198]), .B(A[198]), .Z(n472) );
  AND U532 ( .A(n473), .B(n474), .Z(n471) );
  NANDN U533 ( .A(B[197]), .B(n475), .Z(n474) );
  NANDN U534 ( .A(A[197]), .B(n476), .Z(n475) );
  NANDN U535 ( .A(n476), .B(A[197]), .Z(n473) );
  XOR U536 ( .A(n476), .B(n477), .Z(DIFF[197]) );
  XOR U537 ( .A(B[197]), .B(A[197]), .Z(n477) );
  AND U538 ( .A(n478), .B(n479), .Z(n476) );
  NANDN U539 ( .A(B[196]), .B(n480), .Z(n479) );
  NANDN U540 ( .A(A[196]), .B(n481), .Z(n480) );
  NANDN U541 ( .A(n481), .B(A[196]), .Z(n478) );
  XOR U542 ( .A(n481), .B(n482), .Z(DIFF[196]) );
  XOR U543 ( .A(B[196]), .B(A[196]), .Z(n482) );
  AND U544 ( .A(n483), .B(n484), .Z(n481) );
  NANDN U545 ( .A(B[195]), .B(n485), .Z(n484) );
  NANDN U546 ( .A(A[195]), .B(n486), .Z(n485) );
  NANDN U547 ( .A(n486), .B(A[195]), .Z(n483) );
  XOR U548 ( .A(n486), .B(n487), .Z(DIFF[195]) );
  XOR U549 ( .A(B[195]), .B(A[195]), .Z(n487) );
  AND U550 ( .A(n488), .B(n489), .Z(n486) );
  NANDN U551 ( .A(B[194]), .B(n490), .Z(n489) );
  NANDN U552 ( .A(A[194]), .B(n491), .Z(n490) );
  NANDN U553 ( .A(n491), .B(A[194]), .Z(n488) );
  XOR U554 ( .A(n491), .B(n492), .Z(DIFF[194]) );
  XOR U555 ( .A(B[194]), .B(A[194]), .Z(n492) );
  AND U556 ( .A(n493), .B(n494), .Z(n491) );
  NANDN U557 ( .A(B[193]), .B(n495), .Z(n494) );
  NANDN U558 ( .A(A[193]), .B(n496), .Z(n495) );
  NANDN U559 ( .A(n496), .B(A[193]), .Z(n493) );
  XOR U560 ( .A(n496), .B(n497), .Z(DIFF[193]) );
  XOR U561 ( .A(B[193]), .B(A[193]), .Z(n497) );
  AND U562 ( .A(n498), .B(n499), .Z(n496) );
  NANDN U563 ( .A(B[192]), .B(n500), .Z(n499) );
  NANDN U564 ( .A(A[192]), .B(n501), .Z(n500) );
  NANDN U565 ( .A(n501), .B(A[192]), .Z(n498) );
  XOR U566 ( .A(n501), .B(n502), .Z(DIFF[192]) );
  XOR U567 ( .A(B[192]), .B(A[192]), .Z(n502) );
  AND U568 ( .A(n503), .B(n504), .Z(n501) );
  NANDN U569 ( .A(B[191]), .B(n505), .Z(n504) );
  NANDN U570 ( .A(A[191]), .B(n506), .Z(n505) );
  NANDN U571 ( .A(n506), .B(A[191]), .Z(n503) );
  XOR U572 ( .A(n506), .B(n507), .Z(DIFF[191]) );
  XOR U573 ( .A(B[191]), .B(A[191]), .Z(n507) );
  AND U574 ( .A(n508), .B(n509), .Z(n506) );
  NANDN U575 ( .A(B[190]), .B(n510), .Z(n509) );
  NANDN U576 ( .A(A[190]), .B(n511), .Z(n510) );
  NANDN U577 ( .A(n511), .B(A[190]), .Z(n508) );
  XOR U578 ( .A(n511), .B(n512), .Z(DIFF[190]) );
  XOR U579 ( .A(B[190]), .B(A[190]), .Z(n512) );
  AND U580 ( .A(n513), .B(n514), .Z(n511) );
  NANDN U581 ( .A(B[189]), .B(n515), .Z(n514) );
  NANDN U582 ( .A(A[189]), .B(n516), .Z(n515) );
  NANDN U583 ( .A(n516), .B(A[189]), .Z(n513) );
  XOR U584 ( .A(n517), .B(n518), .Z(DIFF[18]) );
  XOR U585 ( .A(B[18]), .B(A[18]), .Z(n518) );
  XOR U586 ( .A(n516), .B(n519), .Z(DIFF[189]) );
  XOR U587 ( .A(B[189]), .B(A[189]), .Z(n519) );
  AND U588 ( .A(n520), .B(n521), .Z(n516) );
  NANDN U589 ( .A(B[188]), .B(n522), .Z(n521) );
  NANDN U590 ( .A(A[188]), .B(n523), .Z(n522) );
  NANDN U591 ( .A(n523), .B(A[188]), .Z(n520) );
  XOR U592 ( .A(n523), .B(n524), .Z(DIFF[188]) );
  XOR U593 ( .A(B[188]), .B(A[188]), .Z(n524) );
  AND U594 ( .A(n525), .B(n526), .Z(n523) );
  NANDN U595 ( .A(B[187]), .B(n527), .Z(n526) );
  NANDN U596 ( .A(A[187]), .B(n528), .Z(n527) );
  NANDN U597 ( .A(n528), .B(A[187]), .Z(n525) );
  XOR U598 ( .A(n528), .B(n529), .Z(DIFF[187]) );
  XOR U599 ( .A(B[187]), .B(A[187]), .Z(n529) );
  AND U600 ( .A(n530), .B(n531), .Z(n528) );
  NANDN U601 ( .A(B[186]), .B(n532), .Z(n531) );
  NANDN U602 ( .A(A[186]), .B(n533), .Z(n532) );
  NANDN U603 ( .A(n533), .B(A[186]), .Z(n530) );
  XOR U604 ( .A(n533), .B(n534), .Z(DIFF[186]) );
  XOR U605 ( .A(B[186]), .B(A[186]), .Z(n534) );
  AND U606 ( .A(n535), .B(n536), .Z(n533) );
  NANDN U607 ( .A(B[185]), .B(n537), .Z(n536) );
  NANDN U608 ( .A(A[185]), .B(n538), .Z(n537) );
  NANDN U609 ( .A(n538), .B(A[185]), .Z(n535) );
  XOR U610 ( .A(n538), .B(n539), .Z(DIFF[185]) );
  XOR U611 ( .A(B[185]), .B(A[185]), .Z(n539) );
  AND U612 ( .A(n540), .B(n541), .Z(n538) );
  NANDN U613 ( .A(B[184]), .B(n542), .Z(n541) );
  NANDN U614 ( .A(A[184]), .B(n543), .Z(n542) );
  NANDN U615 ( .A(n543), .B(A[184]), .Z(n540) );
  XOR U616 ( .A(n543), .B(n544), .Z(DIFF[184]) );
  XOR U617 ( .A(B[184]), .B(A[184]), .Z(n544) );
  AND U618 ( .A(n545), .B(n546), .Z(n543) );
  NANDN U619 ( .A(B[183]), .B(n547), .Z(n546) );
  NANDN U620 ( .A(A[183]), .B(n548), .Z(n547) );
  NANDN U621 ( .A(n548), .B(A[183]), .Z(n545) );
  XOR U622 ( .A(n548), .B(n549), .Z(DIFF[183]) );
  XOR U623 ( .A(B[183]), .B(A[183]), .Z(n549) );
  AND U624 ( .A(n550), .B(n551), .Z(n548) );
  NANDN U625 ( .A(B[182]), .B(n552), .Z(n551) );
  NANDN U626 ( .A(A[182]), .B(n553), .Z(n552) );
  NANDN U627 ( .A(n553), .B(A[182]), .Z(n550) );
  XOR U628 ( .A(n553), .B(n554), .Z(DIFF[182]) );
  XOR U629 ( .A(B[182]), .B(A[182]), .Z(n554) );
  AND U630 ( .A(n555), .B(n556), .Z(n553) );
  NANDN U631 ( .A(B[181]), .B(n557), .Z(n556) );
  NANDN U632 ( .A(A[181]), .B(n558), .Z(n557) );
  NANDN U633 ( .A(n558), .B(A[181]), .Z(n555) );
  XOR U634 ( .A(n558), .B(n559), .Z(DIFF[181]) );
  XOR U635 ( .A(B[181]), .B(A[181]), .Z(n559) );
  AND U636 ( .A(n560), .B(n561), .Z(n558) );
  NANDN U637 ( .A(B[180]), .B(n562), .Z(n561) );
  NANDN U638 ( .A(A[180]), .B(n563), .Z(n562) );
  NANDN U639 ( .A(n563), .B(A[180]), .Z(n560) );
  XOR U640 ( .A(n563), .B(n564), .Z(DIFF[180]) );
  XOR U641 ( .A(B[180]), .B(A[180]), .Z(n564) );
  AND U642 ( .A(n565), .B(n566), .Z(n563) );
  NANDN U643 ( .A(B[179]), .B(n567), .Z(n566) );
  NANDN U644 ( .A(A[179]), .B(n568), .Z(n567) );
  NANDN U645 ( .A(n568), .B(A[179]), .Z(n565) );
  XOR U646 ( .A(n569), .B(n570), .Z(DIFF[17]) );
  XOR U647 ( .A(B[17]), .B(A[17]), .Z(n570) );
  XOR U648 ( .A(n568), .B(n571), .Z(DIFF[179]) );
  XOR U649 ( .A(B[179]), .B(A[179]), .Z(n571) );
  AND U650 ( .A(n572), .B(n573), .Z(n568) );
  NANDN U651 ( .A(B[178]), .B(n574), .Z(n573) );
  NANDN U652 ( .A(A[178]), .B(n575), .Z(n574) );
  NANDN U653 ( .A(n575), .B(A[178]), .Z(n572) );
  XOR U654 ( .A(n575), .B(n576), .Z(DIFF[178]) );
  XOR U655 ( .A(B[178]), .B(A[178]), .Z(n576) );
  AND U656 ( .A(n577), .B(n578), .Z(n575) );
  NANDN U657 ( .A(B[177]), .B(n579), .Z(n578) );
  NANDN U658 ( .A(A[177]), .B(n580), .Z(n579) );
  NANDN U659 ( .A(n580), .B(A[177]), .Z(n577) );
  XOR U660 ( .A(n580), .B(n581), .Z(DIFF[177]) );
  XOR U661 ( .A(B[177]), .B(A[177]), .Z(n581) );
  AND U662 ( .A(n582), .B(n583), .Z(n580) );
  NANDN U663 ( .A(B[176]), .B(n584), .Z(n583) );
  NANDN U664 ( .A(A[176]), .B(n585), .Z(n584) );
  NANDN U665 ( .A(n585), .B(A[176]), .Z(n582) );
  XOR U666 ( .A(n585), .B(n586), .Z(DIFF[176]) );
  XOR U667 ( .A(B[176]), .B(A[176]), .Z(n586) );
  AND U668 ( .A(n587), .B(n588), .Z(n585) );
  NANDN U669 ( .A(B[175]), .B(n589), .Z(n588) );
  NANDN U670 ( .A(A[175]), .B(n590), .Z(n589) );
  NANDN U671 ( .A(n590), .B(A[175]), .Z(n587) );
  XOR U672 ( .A(n590), .B(n591), .Z(DIFF[175]) );
  XOR U673 ( .A(B[175]), .B(A[175]), .Z(n591) );
  AND U674 ( .A(n592), .B(n593), .Z(n590) );
  NANDN U675 ( .A(B[174]), .B(n594), .Z(n593) );
  NANDN U676 ( .A(A[174]), .B(n595), .Z(n594) );
  NANDN U677 ( .A(n595), .B(A[174]), .Z(n592) );
  XOR U678 ( .A(n595), .B(n596), .Z(DIFF[174]) );
  XOR U679 ( .A(B[174]), .B(A[174]), .Z(n596) );
  AND U680 ( .A(n597), .B(n598), .Z(n595) );
  NANDN U681 ( .A(B[173]), .B(n599), .Z(n598) );
  NANDN U682 ( .A(A[173]), .B(n600), .Z(n599) );
  NANDN U683 ( .A(n600), .B(A[173]), .Z(n597) );
  XOR U684 ( .A(n600), .B(n601), .Z(DIFF[173]) );
  XOR U685 ( .A(B[173]), .B(A[173]), .Z(n601) );
  AND U686 ( .A(n602), .B(n603), .Z(n600) );
  NANDN U687 ( .A(B[172]), .B(n604), .Z(n603) );
  NANDN U688 ( .A(A[172]), .B(n605), .Z(n604) );
  NANDN U689 ( .A(n605), .B(A[172]), .Z(n602) );
  XOR U690 ( .A(n605), .B(n606), .Z(DIFF[172]) );
  XOR U691 ( .A(B[172]), .B(A[172]), .Z(n606) );
  AND U692 ( .A(n607), .B(n608), .Z(n605) );
  NANDN U693 ( .A(B[171]), .B(n609), .Z(n608) );
  NANDN U694 ( .A(A[171]), .B(n610), .Z(n609) );
  NANDN U695 ( .A(n610), .B(A[171]), .Z(n607) );
  XOR U696 ( .A(n610), .B(n611), .Z(DIFF[171]) );
  XOR U697 ( .A(B[171]), .B(A[171]), .Z(n611) );
  AND U698 ( .A(n612), .B(n613), .Z(n610) );
  NANDN U699 ( .A(B[170]), .B(n614), .Z(n613) );
  NANDN U700 ( .A(A[170]), .B(n615), .Z(n614) );
  NANDN U701 ( .A(n615), .B(A[170]), .Z(n612) );
  XOR U702 ( .A(n615), .B(n616), .Z(DIFF[170]) );
  XOR U703 ( .A(B[170]), .B(A[170]), .Z(n616) );
  AND U704 ( .A(n617), .B(n618), .Z(n615) );
  NANDN U705 ( .A(B[169]), .B(n619), .Z(n618) );
  NANDN U706 ( .A(A[169]), .B(n620), .Z(n619) );
  NANDN U707 ( .A(n620), .B(A[169]), .Z(n617) );
  XOR U708 ( .A(n621), .B(n622), .Z(DIFF[16]) );
  XOR U709 ( .A(B[16]), .B(A[16]), .Z(n622) );
  XOR U710 ( .A(n620), .B(n623), .Z(DIFF[169]) );
  XOR U711 ( .A(B[169]), .B(A[169]), .Z(n623) );
  AND U712 ( .A(n624), .B(n625), .Z(n620) );
  NANDN U713 ( .A(B[168]), .B(n626), .Z(n625) );
  NANDN U714 ( .A(A[168]), .B(n627), .Z(n626) );
  NANDN U715 ( .A(n627), .B(A[168]), .Z(n624) );
  XOR U716 ( .A(n627), .B(n628), .Z(DIFF[168]) );
  XOR U717 ( .A(B[168]), .B(A[168]), .Z(n628) );
  AND U718 ( .A(n629), .B(n630), .Z(n627) );
  NANDN U719 ( .A(B[167]), .B(n631), .Z(n630) );
  NANDN U720 ( .A(A[167]), .B(n632), .Z(n631) );
  NANDN U721 ( .A(n632), .B(A[167]), .Z(n629) );
  XOR U722 ( .A(n632), .B(n633), .Z(DIFF[167]) );
  XOR U723 ( .A(B[167]), .B(A[167]), .Z(n633) );
  AND U724 ( .A(n634), .B(n635), .Z(n632) );
  NANDN U725 ( .A(B[166]), .B(n636), .Z(n635) );
  NANDN U726 ( .A(A[166]), .B(n637), .Z(n636) );
  NANDN U727 ( .A(n637), .B(A[166]), .Z(n634) );
  XOR U728 ( .A(n637), .B(n638), .Z(DIFF[166]) );
  XOR U729 ( .A(B[166]), .B(A[166]), .Z(n638) );
  AND U730 ( .A(n639), .B(n640), .Z(n637) );
  NANDN U731 ( .A(B[165]), .B(n641), .Z(n640) );
  NANDN U732 ( .A(A[165]), .B(n642), .Z(n641) );
  NANDN U733 ( .A(n642), .B(A[165]), .Z(n639) );
  XOR U734 ( .A(n642), .B(n643), .Z(DIFF[165]) );
  XOR U735 ( .A(B[165]), .B(A[165]), .Z(n643) );
  AND U736 ( .A(n644), .B(n645), .Z(n642) );
  NANDN U737 ( .A(B[164]), .B(n646), .Z(n645) );
  NANDN U738 ( .A(A[164]), .B(n647), .Z(n646) );
  NANDN U739 ( .A(n647), .B(A[164]), .Z(n644) );
  XOR U740 ( .A(n647), .B(n648), .Z(DIFF[164]) );
  XOR U741 ( .A(B[164]), .B(A[164]), .Z(n648) );
  AND U742 ( .A(n649), .B(n650), .Z(n647) );
  NANDN U743 ( .A(B[163]), .B(n651), .Z(n650) );
  NANDN U744 ( .A(A[163]), .B(n652), .Z(n651) );
  NANDN U745 ( .A(n652), .B(A[163]), .Z(n649) );
  XOR U746 ( .A(n652), .B(n653), .Z(DIFF[163]) );
  XOR U747 ( .A(B[163]), .B(A[163]), .Z(n653) );
  AND U748 ( .A(n654), .B(n655), .Z(n652) );
  NANDN U749 ( .A(B[162]), .B(n656), .Z(n655) );
  NANDN U750 ( .A(A[162]), .B(n657), .Z(n656) );
  NANDN U751 ( .A(n657), .B(A[162]), .Z(n654) );
  XOR U752 ( .A(n657), .B(n658), .Z(DIFF[162]) );
  XOR U753 ( .A(B[162]), .B(A[162]), .Z(n658) );
  AND U754 ( .A(n659), .B(n660), .Z(n657) );
  NANDN U755 ( .A(B[161]), .B(n661), .Z(n660) );
  NANDN U756 ( .A(A[161]), .B(n662), .Z(n661) );
  NANDN U757 ( .A(n662), .B(A[161]), .Z(n659) );
  XOR U758 ( .A(n662), .B(n663), .Z(DIFF[161]) );
  XOR U759 ( .A(B[161]), .B(A[161]), .Z(n663) );
  AND U760 ( .A(n664), .B(n665), .Z(n662) );
  NANDN U761 ( .A(B[160]), .B(n666), .Z(n665) );
  NANDN U762 ( .A(A[160]), .B(n667), .Z(n666) );
  NANDN U763 ( .A(n667), .B(A[160]), .Z(n664) );
  XOR U764 ( .A(n667), .B(n668), .Z(DIFF[160]) );
  XOR U765 ( .A(B[160]), .B(A[160]), .Z(n668) );
  AND U766 ( .A(n669), .B(n670), .Z(n667) );
  NANDN U767 ( .A(B[159]), .B(n671), .Z(n670) );
  NANDN U768 ( .A(A[159]), .B(n672), .Z(n671) );
  NANDN U769 ( .A(n672), .B(A[159]), .Z(n669) );
  XOR U770 ( .A(n673), .B(n674), .Z(DIFF[15]) );
  XOR U771 ( .A(B[15]), .B(A[15]), .Z(n674) );
  XOR U772 ( .A(n672), .B(n675), .Z(DIFF[159]) );
  XOR U773 ( .A(B[159]), .B(A[159]), .Z(n675) );
  AND U774 ( .A(n676), .B(n677), .Z(n672) );
  NANDN U775 ( .A(B[158]), .B(n678), .Z(n677) );
  NANDN U776 ( .A(A[158]), .B(n679), .Z(n678) );
  NANDN U777 ( .A(n679), .B(A[158]), .Z(n676) );
  XOR U778 ( .A(n679), .B(n680), .Z(DIFF[158]) );
  XOR U779 ( .A(B[158]), .B(A[158]), .Z(n680) );
  AND U780 ( .A(n681), .B(n682), .Z(n679) );
  NANDN U781 ( .A(B[157]), .B(n683), .Z(n682) );
  NANDN U782 ( .A(A[157]), .B(n684), .Z(n683) );
  NANDN U783 ( .A(n684), .B(A[157]), .Z(n681) );
  XOR U784 ( .A(n684), .B(n685), .Z(DIFF[157]) );
  XOR U785 ( .A(B[157]), .B(A[157]), .Z(n685) );
  AND U786 ( .A(n686), .B(n687), .Z(n684) );
  NANDN U787 ( .A(B[156]), .B(n688), .Z(n687) );
  NANDN U788 ( .A(A[156]), .B(n689), .Z(n688) );
  NANDN U789 ( .A(n689), .B(A[156]), .Z(n686) );
  XOR U790 ( .A(n689), .B(n690), .Z(DIFF[156]) );
  XOR U791 ( .A(B[156]), .B(A[156]), .Z(n690) );
  AND U792 ( .A(n691), .B(n692), .Z(n689) );
  NANDN U793 ( .A(B[155]), .B(n693), .Z(n692) );
  NANDN U794 ( .A(A[155]), .B(n694), .Z(n693) );
  NANDN U795 ( .A(n694), .B(A[155]), .Z(n691) );
  XOR U796 ( .A(n694), .B(n695), .Z(DIFF[155]) );
  XOR U797 ( .A(B[155]), .B(A[155]), .Z(n695) );
  AND U798 ( .A(n696), .B(n697), .Z(n694) );
  NANDN U799 ( .A(B[154]), .B(n698), .Z(n697) );
  NANDN U800 ( .A(A[154]), .B(n699), .Z(n698) );
  NANDN U801 ( .A(n699), .B(A[154]), .Z(n696) );
  XOR U802 ( .A(n699), .B(n700), .Z(DIFF[154]) );
  XOR U803 ( .A(B[154]), .B(A[154]), .Z(n700) );
  AND U804 ( .A(n701), .B(n702), .Z(n699) );
  NANDN U805 ( .A(B[153]), .B(n703), .Z(n702) );
  NANDN U806 ( .A(A[153]), .B(n704), .Z(n703) );
  NANDN U807 ( .A(n704), .B(A[153]), .Z(n701) );
  XOR U808 ( .A(n704), .B(n705), .Z(DIFF[153]) );
  XOR U809 ( .A(B[153]), .B(A[153]), .Z(n705) );
  AND U810 ( .A(n706), .B(n707), .Z(n704) );
  NANDN U811 ( .A(B[152]), .B(n708), .Z(n707) );
  NANDN U812 ( .A(A[152]), .B(n709), .Z(n708) );
  NANDN U813 ( .A(n709), .B(A[152]), .Z(n706) );
  XOR U814 ( .A(n709), .B(n710), .Z(DIFF[152]) );
  XOR U815 ( .A(B[152]), .B(A[152]), .Z(n710) );
  AND U816 ( .A(n711), .B(n712), .Z(n709) );
  NANDN U817 ( .A(B[151]), .B(n713), .Z(n712) );
  NANDN U818 ( .A(A[151]), .B(n714), .Z(n713) );
  NANDN U819 ( .A(n714), .B(A[151]), .Z(n711) );
  XOR U820 ( .A(n714), .B(n715), .Z(DIFF[151]) );
  XOR U821 ( .A(B[151]), .B(A[151]), .Z(n715) );
  AND U822 ( .A(n716), .B(n717), .Z(n714) );
  NANDN U823 ( .A(B[150]), .B(n718), .Z(n717) );
  NANDN U824 ( .A(A[150]), .B(n719), .Z(n718) );
  NANDN U825 ( .A(n719), .B(A[150]), .Z(n716) );
  XOR U826 ( .A(n719), .B(n720), .Z(DIFF[150]) );
  XOR U827 ( .A(B[150]), .B(A[150]), .Z(n720) );
  AND U828 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U829 ( .A(B[149]), .B(n723), .Z(n722) );
  NANDN U830 ( .A(A[149]), .B(n724), .Z(n723) );
  NANDN U831 ( .A(n724), .B(A[149]), .Z(n721) );
  XOR U832 ( .A(n725), .B(n726), .Z(DIFF[14]) );
  XOR U833 ( .A(B[14]), .B(A[14]), .Z(n726) );
  XOR U834 ( .A(n724), .B(n727), .Z(DIFF[149]) );
  XOR U835 ( .A(B[149]), .B(A[149]), .Z(n727) );
  AND U836 ( .A(n728), .B(n729), .Z(n724) );
  NANDN U837 ( .A(B[148]), .B(n730), .Z(n729) );
  NANDN U838 ( .A(A[148]), .B(n731), .Z(n730) );
  NANDN U839 ( .A(n731), .B(A[148]), .Z(n728) );
  XOR U840 ( .A(n731), .B(n732), .Z(DIFF[148]) );
  XOR U841 ( .A(B[148]), .B(A[148]), .Z(n732) );
  AND U842 ( .A(n733), .B(n734), .Z(n731) );
  NANDN U843 ( .A(B[147]), .B(n735), .Z(n734) );
  NANDN U844 ( .A(A[147]), .B(n736), .Z(n735) );
  NANDN U845 ( .A(n736), .B(A[147]), .Z(n733) );
  XOR U846 ( .A(n736), .B(n737), .Z(DIFF[147]) );
  XOR U847 ( .A(B[147]), .B(A[147]), .Z(n737) );
  AND U848 ( .A(n738), .B(n739), .Z(n736) );
  NANDN U849 ( .A(B[146]), .B(n740), .Z(n739) );
  NANDN U850 ( .A(A[146]), .B(n741), .Z(n740) );
  NANDN U851 ( .A(n741), .B(A[146]), .Z(n738) );
  XOR U852 ( .A(n741), .B(n742), .Z(DIFF[146]) );
  XOR U853 ( .A(B[146]), .B(A[146]), .Z(n742) );
  AND U854 ( .A(n743), .B(n744), .Z(n741) );
  NANDN U855 ( .A(B[145]), .B(n745), .Z(n744) );
  NANDN U856 ( .A(A[145]), .B(n746), .Z(n745) );
  NANDN U857 ( .A(n746), .B(A[145]), .Z(n743) );
  XOR U858 ( .A(n746), .B(n747), .Z(DIFF[145]) );
  XOR U859 ( .A(B[145]), .B(A[145]), .Z(n747) );
  AND U860 ( .A(n748), .B(n749), .Z(n746) );
  NANDN U861 ( .A(B[144]), .B(n750), .Z(n749) );
  NANDN U862 ( .A(A[144]), .B(n751), .Z(n750) );
  NANDN U863 ( .A(n751), .B(A[144]), .Z(n748) );
  XOR U864 ( .A(n751), .B(n752), .Z(DIFF[144]) );
  XOR U865 ( .A(B[144]), .B(A[144]), .Z(n752) );
  AND U866 ( .A(n753), .B(n754), .Z(n751) );
  NANDN U867 ( .A(B[143]), .B(n755), .Z(n754) );
  NANDN U868 ( .A(A[143]), .B(n756), .Z(n755) );
  NANDN U869 ( .A(n756), .B(A[143]), .Z(n753) );
  XOR U870 ( .A(n756), .B(n757), .Z(DIFF[143]) );
  XOR U871 ( .A(B[143]), .B(A[143]), .Z(n757) );
  AND U872 ( .A(n758), .B(n759), .Z(n756) );
  NANDN U873 ( .A(B[142]), .B(n760), .Z(n759) );
  NANDN U874 ( .A(A[142]), .B(n761), .Z(n760) );
  NANDN U875 ( .A(n761), .B(A[142]), .Z(n758) );
  XOR U876 ( .A(n761), .B(n762), .Z(DIFF[142]) );
  XOR U877 ( .A(B[142]), .B(A[142]), .Z(n762) );
  AND U878 ( .A(n763), .B(n764), .Z(n761) );
  NANDN U879 ( .A(B[141]), .B(n765), .Z(n764) );
  NANDN U880 ( .A(A[141]), .B(n766), .Z(n765) );
  NANDN U881 ( .A(n766), .B(A[141]), .Z(n763) );
  XOR U882 ( .A(n766), .B(n767), .Z(DIFF[141]) );
  XOR U883 ( .A(B[141]), .B(A[141]), .Z(n767) );
  AND U884 ( .A(n768), .B(n769), .Z(n766) );
  NANDN U885 ( .A(B[140]), .B(n770), .Z(n769) );
  NANDN U886 ( .A(A[140]), .B(n771), .Z(n770) );
  NANDN U887 ( .A(n771), .B(A[140]), .Z(n768) );
  XOR U888 ( .A(n771), .B(n772), .Z(DIFF[140]) );
  XOR U889 ( .A(B[140]), .B(A[140]), .Z(n772) );
  AND U890 ( .A(n773), .B(n774), .Z(n771) );
  NANDN U891 ( .A(B[139]), .B(n775), .Z(n774) );
  NANDN U892 ( .A(A[139]), .B(n776), .Z(n775) );
  NANDN U893 ( .A(n776), .B(A[139]), .Z(n773) );
  XOR U894 ( .A(n777), .B(n778), .Z(DIFF[13]) );
  XOR U895 ( .A(B[13]), .B(A[13]), .Z(n778) );
  XOR U896 ( .A(n776), .B(n779), .Z(DIFF[139]) );
  XOR U897 ( .A(B[139]), .B(A[139]), .Z(n779) );
  AND U898 ( .A(n780), .B(n781), .Z(n776) );
  NANDN U899 ( .A(B[138]), .B(n782), .Z(n781) );
  NANDN U900 ( .A(A[138]), .B(n783), .Z(n782) );
  NANDN U901 ( .A(n783), .B(A[138]), .Z(n780) );
  XOR U902 ( .A(n783), .B(n784), .Z(DIFF[138]) );
  XOR U903 ( .A(B[138]), .B(A[138]), .Z(n784) );
  AND U904 ( .A(n785), .B(n786), .Z(n783) );
  NANDN U905 ( .A(B[137]), .B(n787), .Z(n786) );
  NANDN U906 ( .A(A[137]), .B(n788), .Z(n787) );
  NANDN U907 ( .A(n788), .B(A[137]), .Z(n785) );
  XOR U908 ( .A(n788), .B(n789), .Z(DIFF[137]) );
  XOR U909 ( .A(B[137]), .B(A[137]), .Z(n789) );
  AND U910 ( .A(n790), .B(n791), .Z(n788) );
  NANDN U911 ( .A(B[136]), .B(n792), .Z(n791) );
  NANDN U912 ( .A(A[136]), .B(n793), .Z(n792) );
  NANDN U913 ( .A(n793), .B(A[136]), .Z(n790) );
  XOR U914 ( .A(n793), .B(n794), .Z(DIFF[136]) );
  XOR U915 ( .A(B[136]), .B(A[136]), .Z(n794) );
  AND U916 ( .A(n795), .B(n796), .Z(n793) );
  NANDN U917 ( .A(B[135]), .B(n797), .Z(n796) );
  NANDN U918 ( .A(A[135]), .B(n798), .Z(n797) );
  NANDN U919 ( .A(n798), .B(A[135]), .Z(n795) );
  XOR U920 ( .A(n798), .B(n799), .Z(DIFF[135]) );
  XOR U921 ( .A(B[135]), .B(A[135]), .Z(n799) );
  AND U922 ( .A(n800), .B(n801), .Z(n798) );
  NANDN U923 ( .A(B[134]), .B(n802), .Z(n801) );
  NANDN U924 ( .A(A[134]), .B(n803), .Z(n802) );
  NANDN U925 ( .A(n803), .B(A[134]), .Z(n800) );
  XOR U926 ( .A(n803), .B(n804), .Z(DIFF[134]) );
  XOR U927 ( .A(B[134]), .B(A[134]), .Z(n804) );
  AND U928 ( .A(n805), .B(n806), .Z(n803) );
  NANDN U929 ( .A(B[133]), .B(n807), .Z(n806) );
  NANDN U930 ( .A(A[133]), .B(n808), .Z(n807) );
  NANDN U931 ( .A(n808), .B(A[133]), .Z(n805) );
  XOR U932 ( .A(n808), .B(n809), .Z(DIFF[133]) );
  XOR U933 ( .A(B[133]), .B(A[133]), .Z(n809) );
  AND U934 ( .A(n810), .B(n811), .Z(n808) );
  NANDN U935 ( .A(B[132]), .B(n812), .Z(n811) );
  NANDN U936 ( .A(A[132]), .B(n813), .Z(n812) );
  NANDN U937 ( .A(n813), .B(A[132]), .Z(n810) );
  XOR U938 ( .A(n813), .B(n814), .Z(DIFF[132]) );
  XOR U939 ( .A(B[132]), .B(A[132]), .Z(n814) );
  AND U940 ( .A(n815), .B(n816), .Z(n813) );
  NANDN U941 ( .A(B[131]), .B(n817), .Z(n816) );
  NANDN U942 ( .A(A[131]), .B(n818), .Z(n817) );
  NANDN U943 ( .A(n818), .B(A[131]), .Z(n815) );
  XOR U944 ( .A(n818), .B(n819), .Z(DIFF[131]) );
  XOR U945 ( .A(B[131]), .B(A[131]), .Z(n819) );
  AND U946 ( .A(n820), .B(n821), .Z(n818) );
  NANDN U947 ( .A(B[130]), .B(n822), .Z(n821) );
  NANDN U948 ( .A(A[130]), .B(n823), .Z(n822) );
  NANDN U949 ( .A(n823), .B(A[130]), .Z(n820) );
  XOR U950 ( .A(n823), .B(n824), .Z(DIFF[130]) );
  XOR U951 ( .A(B[130]), .B(A[130]), .Z(n824) );
  AND U952 ( .A(n825), .B(n826), .Z(n823) );
  NANDN U953 ( .A(B[129]), .B(n827), .Z(n826) );
  NANDN U954 ( .A(A[129]), .B(n828), .Z(n827) );
  NANDN U955 ( .A(n828), .B(A[129]), .Z(n825) );
  XOR U956 ( .A(n829), .B(n830), .Z(DIFF[12]) );
  XOR U957 ( .A(B[12]), .B(A[12]), .Z(n830) );
  XOR U958 ( .A(n828), .B(n831), .Z(DIFF[129]) );
  XOR U959 ( .A(B[129]), .B(A[129]), .Z(n831) );
  AND U960 ( .A(n832), .B(n833), .Z(n828) );
  NANDN U961 ( .A(B[128]), .B(n834), .Z(n833) );
  NANDN U962 ( .A(A[128]), .B(n835), .Z(n834) );
  NANDN U963 ( .A(n835), .B(A[128]), .Z(n832) );
  XOR U964 ( .A(n835), .B(n836), .Z(DIFF[128]) );
  XOR U965 ( .A(B[128]), .B(A[128]), .Z(n836) );
  AND U966 ( .A(n837), .B(n838), .Z(n835) );
  NANDN U967 ( .A(B[127]), .B(n839), .Z(n838) );
  NANDN U968 ( .A(A[127]), .B(n840), .Z(n839) );
  NANDN U969 ( .A(n840), .B(A[127]), .Z(n837) );
  XOR U970 ( .A(n840), .B(n841), .Z(DIFF[127]) );
  XOR U971 ( .A(B[127]), .B(A[127]), .Z(n841) );
  AND U972 ( .A(n842), .B(n843), .Z(n840) );
  NANDN U973 ( .A(B[126]), .B(n844), .Z(n843) );
  NANDN U974 ( .A(A[126]), .B(n845), .Z(n844) );
  NANDN U975 ( .A(n845), .B(A[126]), .Z(n842) );
  XOR U976 ( .A(n845), .B(n846), .Z(DIFF[126]) );
  XOR U977 ( .A(B[126]), .B(A[126]), .Z(n846) );
  AND U978 ( .A(n847), .B(n848), .Z(n845) );
  NANDN U979 ( .A(B[125]), .B(n849), .Z(n848) );
  NANDN U980 ( .A(A[125]), .B(n850), .Z(n849) );
  NANDN U981 ( .A(n850), .B(A[125]), .Z(n847) );
  XOR U982 ( .A(n850), .B(n851), .Z(DIFF[125]) );
  XOR U983 ( .A(B[125]), .B(A[125]), .Z(n851) );
  AND U984 ( .A(n852), .B(n853), .Z(n850) );
  NANDN U985 ( .A(B[124]), .B(n854), .Z(n853) );
  NANDN U986 ( .A(A[124]), .B(n855), .Z(n854) );
  NANDN U987 ( .A(n855), .B(A[124]), .Z(n852) );
  XOR U988 ( .A(n855), .B(n856), .Z(DIFF[124]) );
  XOR U989 ( .A(B[124]), .B(A[124]), .Z(n856) );
  AND U990 ( .A(n857), .B(n858), .Z(n855) );
  NANDN U991 ( .A(B[123]), .B(n859), .Z(n858) );
  NANDN U992 ( .A(A[123]), .B(n860), .Z(n859) );
  NANDN U993 ( .A(n860), .B(A[123]), .Z(n857) );
  XOR U994 ( .A(n860), .B(n861), .Z(DIFF[123]) );
  XOR U995 ( .A(B[123]), .B(A[123]), .Z(n861) );
  AND U996 ( .A(n862), .B(n863), .Z(n860) );
  NANDN U997 ( .A(B[122]), .B(n864), .Z(n863) );
  NANDN U998 ( .A(A[122]), .B(n865), .Z(n864) );
  NANDN U999 ( .A(n865), .B(A[122]), .Z(n862) );
  XOR U1000 ( .A(n865), .B(n866), .Z(DIFF[122]) );
  XOR U1001 ( .A(B[122]), .B(A[122]), .Z(n866) );
  AND U1002 ( .A(n867), .B(n868), .Z(n865) );
  NANDN U1003 ( .A(B[121]), .B(n869), .Z(n868) );
  NANDN U1004 ( .A(A[121]), .B(n870), .Z(n869) );
  NANDN U1005 ( .A(n870), .B(A[121]), .Z(n867) );
  XOR U1006 ( .A(n870), .B(n871), .Z(DIFF[121]) );
  XOR U1007 ( .A(B[121]), .B(A[121]), .Z(n871) );
  AND U1008 ( .A(n872), .B(n873), .Z(n870) );
  NANDN U1009 ( .A(B[120]), .B(n874), .Z(n873) );
  NANDN U1010 ( .A(A[120]), .B(n875), .Z(n874) );
  NANDN U1011 ( .A(n875), .B(A[120]), .Z(n872) );
  XOR U1012 ( .A(n875), .B(n876), .Z(DIFF[120]) );
  XOR U1013 ( .A(B[120]), .B(A[120]), .Z(n876) );
  AND U1014 ( .A(n877), .B(n878), .Z(n875) );
  NANDN U1015 ( .A(B[119]), .B(n879), .Z(n878) );
  NANDN U1016 ( .A(A[119]), .B(n880), .Z(n879) );
  NANDN U1017 ( .A(n880), .B(A[119]), .Z(n877) );
  XOR U1018 ( .A(n881), .B(n882), .Z(DIFF[11]) );
  XOR U1019 ( .A(B[11]), .B(A[11]), .Z(n882) );
  XOR U1020 ( .A(n880), .B(n883), .Z(DIFF[119]) );
  XOR U1021 ( .A(B[119]), .B(A[119]), .Z(n883) );
  AND U1022 ( .A(n884), .B(n885), .Z(n880) );
  NANDN U1023 ( .A(B[118]), .B(n886), .Z(n885) );
  NANDN U1024 ( .A(A[118]), .B(n887), .Z(n886) );
  NANDN U1025 ( .A(n887), .B(A[118]), .Z(n884) );
  XOR U1026 ( .A(n887), .B(n888), .Z(DIFF[118]) );
  XOR U1027 ( .A(B[118]), .B(A[118]), .Z(n888) );
  AND U1028 ( .A(n889), .B(n890), .Z(n887) );
  NANDN U1029 ( .A(B[117]), .B(n891), .Z(n890) );
  NANDN U1030 ( .A(A[117]), .B(n892), .Z(n891) );
  NANDN U1031 ( .A(n892), .B(A[117]), .Z(n889) );
  XOR U1032 ( .A(n892), .B(n893), .Z(DIFF[117]) );
  XOR U1033 ( .A(B[117]), .B(A[117]), .Z(n893) );
  AND U1034 ( .A(n894), .B(n895), .Z(n892) );
  NANDN U1035 ( .A(B[116]), .B(n896), .Z(n895) );
  NANDN U1036 ( .A(A[116]), .B(n897), .Z(n896) );
  NANDN U1037 ( .A(n897), .B(A[116]), .Z(n894) );
  XOR U1038 ( .A(n897), .B(n898), .Z(DIFF[116]) );
  XOR U1039 ( .A(B[116]), .B(A[116]), .Z(n898) );
  AND U1040 ( .A(n899), .B(n900), .Z(n897) );
  NANDN U1041 ( .A(B[115]), .B(n901), .Z(n900) );
  NANDN U1042 ( .A(A[115]), .B(n902), .Z(n901) );
  NANDN U1043 ( .A(n902), .B(A[115]), .Z(n899) );
  XOR U1044 ( .A(n902), .B(n903), .Z(DIFF[115]) );
  XOR U1045 ( .A(B[115]), .B(A[115]), .Z(n903) );
  AND U1046 ( .A(n904), .B(n905), .Z(n902) );
  NANDN U1047 ( .A(B[114]), .B(n906), .Z(n905) );
  NANDN U1048 ( .A(A[114]), .B(n907), .Z(n906) );
  NANDN U1049 ( .A(n907), .B(A[114]), .Z(n904) );
  XOR U1050 ( .A(n907), .B(n908), .Z(DIFF[114]) );
  XOR U1051 ( .A(B[114]), .B(A[114]), .Z(n908) );
  AND U1052 ( .A(n909), .B(n910), .Z(n907) );
  NANDN U1053 ( .A(B[113]), .B(n911), .Z(n910) );
  NANDN U1054 ( .A(A[113]), .B(n912), .Z(n911) );
  NANDN U1055 ( .A(n912), .B(A[113]), .Z(n909) );
  XOR U1056 ( .A(n912), .B(n913), .Z(DIFF[113]) );
  XOR U1057 ( .A(B[113]), .B(A[113]), .Z(n913) );
  AND U1058 ( .A(n914), .B(n915), .Z(n912) );
  NANDN U1059 ( .A(B[112]), .B(n916), .Z(n915) );
  NANDN U1060 ( .A(A[112]), .B(n917), .Z(n916) );
  NANDN U1061 ( .A(n917), .B(A[112]), .Z(n914) );
  XOR U1062 ( .A(n917), .B(n918), .Z(DIFF[112]) );
  XOR U1063 ( .A(B[112]), .B(A[112]), .Z(n918) );
  AND U1064 ( .A(n919), .B(n920), .Z(n917) );
  NANDN U1065 ( .A(B[111]), .B(n921), .Z(n920) );
  NANDN U1066 ( .A(A[111]), .B(n922), .Z(n921) );
  NANDN U1067 ( .A(n922), .B(A[111]), .Z(n919) );
  XOR U1068 ( .A(n922), .B(n923), .Z(DIFF[111]) );
  XOR U1069 ( .A(B[111]), .B(A[111]), .Z(n923) );
  AND U1070 ( .A(n924), .B(n925), .Z(n922) );
  NANDN U1071 ( .A(B[110]), .B(n926), .Z(n925) );
  NANDN U1072 ( .A(A[110]), .B(n927), .Z(n926) );
  NANDN U1073 ( .A(n927), .B(A[110]), .Z(n924) );
  XOR U1074 ( .A(n927), .B(n928), .Z(DIFF[110]) );
  XOR U1075 ( .A(B[110]), .B(A[110]), .Z(n928) );
  AND U1076 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U1077 ( .A(B[109]), .B(n931), .Z(n930) );
  NANDN U1078 ( .A(A[109]), .B(n932), .Z(n931) );
  NANDN U1079 ( .A(n932), .B(A[109]), .Z(n929) );
  XOR U1080 ( .A(n933), .B(n934), .Z(DIFF[10]) );
  XOR U1081 ( .A(B[10]), .B(A[10]), .Z(n934) );
  XOR U1082 ( .A(n932), .B(n935), .Z(DIFF[109]) );
  XOR U1083 ( .A(B[109]), .B(A[109]), .Z(n935) );
  AND U1084 ( .A(n936), .B(n937), .Z(n932) );
  NANDN U1085 ( .A(B[108]), .B(n938), .Z(n937) );
  NANDN U1086 ( .A(A[108]), .B(n939), .Z(n938) );
  NANDN U1087 ( .A(n939), .B(A[108]), .Z(n936) );
  XOR U1088 ( .A(n939), .B(n940), .Z(DIFF[108]) );
  XOR U1089 ( .A(B[108]), .B(A[108]), .Z(n940) );
  AND U1090 ( .A(n941), .B(n942), .Z(n939) );
  NANDN U1091 ( .A(B[107]), .B(n943), .Z(n942) );
  NANDN U1092 ( .A(A[107]), .B(n944), .Z(n943) );
  NANDN U1093 ( .A(n944), .B(A[107]), .Z(n941) );
  XOR U1094 ( .A(n944), .B(n945), .Z(DIFF[107]) );
  XOR U1095 ( .A(B[107]), .B(A[107]), .Z(n945) );
  AND U1096 ( .A(n946), .B(n947), .Z(n944) );
  NANDN U1097 ( .A(B[106]), .B(n948), .Z(n947) );
  NANDN U1098 ( .A(A[106]), .B(n949), .Z(n948) );
  NANDN U1099 ( .A(n949), .B(A[106]), .Z(n946) );
  XOR U1100 ( .A(n949), .B(n950), .Z(DIFF[106]) );
  XOR U1101 ( .A(B[106]), .B(A[106]), .Z(n950) );
  AND U1102 ( .A(n951), .B(n952), .Z(n949) );
  NANDN U1103 ( .A(B[105]), .B(n953), .Z(n952) );
  NANDN U1104 ( .A(A[105]), .B(n954), .Z(n953) );
  NANDN U1105 ( .A(n954), .B(A[105]), .Z(n951) );
  XOR U1106 ( .A(n954), .B(n955), .Z(DIFF[105]) );
  XOR U1107 ( .A(B[105]), .B(A[105]), .Z(n955) );
  AND U1108 ( .A(n956), .B(n957), .Z(n954) );
  NANDN U1109 ( .A(B[104]), .B(n958), .Z(n957) );
  NANDN U1110 ( .A(A[104]), .B(n959), .Z(n958) );
  NANDN U1111 ( .A(n959), .B(A[104]), .Z(n956) );
  XOR U1112 ( .A(n959), .B(n960), .Z(DIFF[104]) );
  XOR U1113 ( .A(B[104]), .B(A[104]), .Z(n960) );
  AND U1114 ( .A(n961), .B(n962), .Z(n959) );
  NANDN U1115 ( .A(B[103]), .B(n963), .Z(n962) );
  NANDN U1116 ( .A(A[103]), .B(n964), .Z(n963) );
  NANDN U1117 ( .A(n964), .B(A[103]), .Z(n961) );
  XOR U1118 ( .A(n964), .B(n965), .Z(DIFF[103]) );
  XOR U1119 ( .A(B[103]), .B(A[103]), .Z(n965) );
  AND U1120 ( .A(n966), .B(n967), .Z(n964) );
  NANDN U1121 ( .A(B[102]), .B(n968), .Z(n967) );
  NANDN U1122 ( .A(A[102]), .B(n969), .Z(n968) );
  NANDN U1123 ( .A(n969), .B(A[102]), .Z(n966) );
  XOR U1124 ( .A(n969), .B(n970), .Z(DIFF[102]) );
  XOR U1125 ( .A(B[102]), .B(A[102]), .Z(n970) );
  AND U1126 ( .A(n971), .B(n972), .Z(n969) );
  NANDN U1127 ( .A(B[101]), .B(n973), .Z(n972) );
  NANDN U1128 ( .A(A[101]), .B(n974), .Z(n973) );
  NANDN U1129 ( .A(n974), .B(A[101]), .Z(n971) );
  XOR U1130 ( .A(n974), .B(n975), .Z(DIFF[101]) );
  XOR U1131 ( .A(B[101]), .B(A[101]), .Z(n975) );
  AND U1132 ( .A(n976), .B(n977), .Z(n974) );
  NANDN U1133 ( .A(B[100]), .B(n978), .Z(n977) );
  NANDN U1134 ( .A(A[100]), .B(n979), .Z(n978) );
  NANDN U1135 ( .A(n979), .B(A[100]), .Z(n976) );
  XOR U1136 ( .A(n979), .B(n980), .Z(DIFF[100]) );
  XOR U1137 ( .A(B[100]), .B(A[100]), .Z(n980) );
  AND U1138 ( .A(n981), .B(n982), .Z(n979) );
  NANDN U1139 ( .A(B[99]), .B(n983), .Z(n982) );
  OR U1140 ( .A(n5), .B(A[99]), .Z(n983) );
  NAND U1141 ( .A(A[99]), .B(n5), .Z(n981) );
  NAND U1142 ( .A(n984), .B(n985), .Z(n5) );
  NANDN U1143 ( .A(B[98]), .B(n986), .Z(n985) );
  NANDN U1144 ( .A(A[98]), .B(n7), .Z(n986) );
  NANDN U1145 ( .A(n7), .B(A[98]), .Z(n984) );
  AND U1146 ( .A(n987), .B(n988), .Z(n7) );
  NANDN U1147 ( .A(B[97]), .B(n989), .Z(n988) );
  NANDN U1148 ( .A(A[97]), .B(n9), .Z(n989) );
  NANDN U1149 ( .A(n9), .B(A[97]), .Z(n987) );
  AND U1150 ( .A(n990), .B(n991), .Z(n9) );
  NANDN U1151 ( .A(B[96]), .B(n992), .Z(n991) );
  NANDN U1152 ( .A(A[96]), .B(n11), .Z(n992) );
  NANDN U1153 ( .A(n11), .B(A[96]), .Z(n990) );
  AND U1154 ( .A(n993), .B(n994), .Z(n11) );
  NANDN U1155 ( .A(B[95]), .B(n995), .Z(n994) );
  NANDN U1156 ( .A(A[95]), .B(n13), .Z(n995) );
  NANDN U1157 ( .A(n13), .B(A[95]), .Z(n993) );
  AND U1158 ( .A(n996), .B(n997), .Z(n13) );
  NANDN U1159 ( .A(B[94]), .B(n998), .Z(n997) );
  NANDN U1160 ( .A(A[94]), .B(n15), .Z(n998) );
  NANDN U1161 ( .A(n15), .B(A[94]), .Z(n996) );
  AND U1162 ( .A(n999), .B(n1000), .Z(n15) );
  NANDN U1163 ( .A(B[93]), .B(n1001), .Z(n1000) );
  NANDN U1164 ( .A(A[93]), .B(n17), .Z(n1001) );
  NANDN U1165 ( .A(n17), .B(A[93]), .Z(n999) );
  AND U1166 ( .A(n1002), .B(n1003), .Z(n17) );
  NANDN U1167 ( .A(B[92]), .B(n1004), .Z(n1003) );
  NANDN U1168 ( .A(A[92]), .B(n19), .Z(n1004) );
  NANDN U1169 ( .A(n19), .B(A[92]), .Z(n1002) );
  AND U1170 ( .A(n1005), .B(n1006), .Z(n19) );
  NANDN U1171 ( .A(B[91]), .B(n1007), .Z(n1006) );
  NANDN U1172 ( .A(A[91]), .B(n21), .Z(n1007) );
  NANDN U1173 ( .A(n21), .B(A[91]), .Z(n1005) );
  AND U1174 ( .A(n1008), .B(n1009), .Z(n21) );
  NANDN U1175 ( .A(B[90]), .B(n1010), .Z(n1009) );
  NANDN U1176 ( .A(A[90]), .B(n23), .Z(n1010) );
  NANDN U1177 ( .A(n23), .B(A[90]), .Z(n1008) );
  AND U1178 ( .A(n1011), .B(n1012), .Z(n23) );
  NANDN U1179 ( .A(B[89]), .B(n1013), .Z(n1012) );
  NANDN U1180 ( .A(A[89]), .B(n27), .Z(n1013) );
  NANDN U1181 ( .A(n27), .B(A[89]), .Z(n1011) );
  AND U1182 ( .A(n1014), .B(n1015), .Z(n27) );
  NANDN U1183 ( .A(B[88]), .B(n1016), .Z(n1015) );
  NANDN U1184 ( .A(A[88]), .B(n29), .Z(n1016) );
  NANDN U1185 ( .A(n29), .B(A[88]), .Z(n1014) );
  AND U1186 ( .A(n1017), .B(n1018), .Z(n29) );
  NANDN U1187 ( .A(B[87]), .B(n1019), .Z(n1018) );
  NANDN U1188 ( .A(A[87]), .B(n31), .Z(n1019) );
  NANDN U1189 ( .A(n31), .B(A[87]), .Z(n1017) );
  AND U1190 ( .A(n1020), .B(n1021), .Z(n31) );
  NANDN U1191 ( .A(B[86]), .B(n1022), .Z(n1021) );
  NANDN U1192 ( .A(A[86]), .B(n33), .Z(n1022) );
  NANDN U1193 ( .A(n33), .B(A[86]), .Z(n1020) );
  AND U1194 ( .A(n1023), .B(n1024), .Z(n33) );
  NANDN U1195 ( .A(B[85]), .B(n1025), .Z(n1024) );
  NANDN U1196 ( .A(A[85]), .B(n35), .Z(n1025) );
  NANDN U1197 ( .A(n35), .B(A[85]), .Z(n1023) );
  AND U1198 ( .A(n1026), .B(n1027), .Z(n35) );
  NANDN U1199 ( .A(B[84]), .B(n1028), .Z(n1027) );
  NANDN U1200 ( .A(A[84]), .B(n37), .Z(n1028) );
  NANDN U1201 ( .A(n37), .B(A[84]), .Z(n1026) );
  AND U1202 ( .A(n1029), .B(n1030), .Z(n37) );
  NANDN U1203 ( .A(B[83]), .B(n1031), .Z(n1030) );
  NANDN U1204 ( .A(A[83]), .B(n39), .Z(n1031) );
  NANDN U1205 ( .A(n39), .B(A[83]), .Z(n1029) );
  AND U1206 ( .A(n1032), .B(n1033), .Z(n39) );
  NANDN U1207 ( .A(B[82]), .B(n1034), .Z(n1033) );
  NANDN U1208 ( .A(A[82]), .B(n41), .Z(n1034) );
  NANDN U1209 ( .A(n41), .B(A[82]), .Z(n1032) );
  AND U1210 ( .A(n1035), .B(n1036), .Z(n41) );
  NANDN U1211 ( .A(B[81]), .B(n1037), .Z(n1036) );
  NANDN U1212 ( .A(A[81]), .B(n43), .Z(n1037) );
  NANDN U1213 ( .A(n43), .B(A[81]), .Z(n1035) );
  AND U1214 ( .A(n1038), .B(n1039), .Z(n43) );
  NANDN U1215 ( .A(B[80]), .B(n1040), .Z(n1039) );
  NANDN U1216 ( .A(A[80]), .B(n45), .Z(n1040) );
  NANDN U1217 ( .A(n45), .B(A[80]), .Z(n1038) );
  AND U1218 ( .A(n1041), .B(n1042), .Z(n45) );
  NANDN U1219 ( .A(B[79]), .B(n1043), .Z(n1042) );
  NANDN U1220 ( .A(A[79]), .B(n49), .Z(n1043) );
  NANDN U1221 ( .A(n49), .B(A[79]), .Z(n1041) );
  AND U1222 ( .A(n1044), .B(n1045), .Z(n49) );
  NANDN U1223 ( .A(B[78]), .B(n1046), .Z(n1045) );
  NANDN U1224 ( .A(A[78]), .B(n51), .Z(n1046) );
  NANDN U1225 ( .A(n51), .B(A[78]), .Z(n1044) );
  AND U1226 ( .A(n1047), .B(n1048), .Z(n51) );
  NANDN U1227 ( .A(B[77]), .B(n1049), .Z(n1048) );
  NANDN U1228 ( .A(A[77]), .B(n53), .Z(n1049) );
  NANDN U1229 ( .A(n53), .B(A[77]), .Z(n1047) );
  AND U1230 ( .A(n1050), .B(n1051), .Z(n53) );
  NANDN U1231 ( .A(B[76]), .B(n1052), .Z(n1051) );
  NANDN U1232 ( .A(A[76]), .B(n55), .Z(n1052) );
  NANDN U1233 ( .A(n55), .B(A[76]), .Z(n1050) );
  AND U1234 ( .A(n1053), .B(n1054), .Z(n55) );
  NANDN U1235 ( .A(B[75]), .B(n1055), .Z(n1054) );
  NANDN U1236 ( .A(A[75]), .B(n57), .Z(n1055) );
  NANDN U1237 ( .A(n57), .B(A[75]), .Z(n1053) );
  AND U1238 ( .A(n1056), .B(n1057), .Z(n57) );
  NANDN U1239 ( .A(B[74]), .B(n1058), .Z(n1057) );
  NANDN U1240 ( .A(A[74]), .B(n59), .Z(n1058) );
  NANDN U1241 ( .A(n59), .B(A[74]), .Z(n1056) );
  AND U1242 ( .A(n1059), .B(n1060), .Z(n59) );
  NANDN U1243 ( .A(B[73]), .B(n1061), .Z(n1060) );
  NANDN U1244 ( .A(A[73]), .B(n61), .Z(n1061) );
  NANDN U1245 ( .A(n61), .B(A[73]), .Z(n1059) );
  AND U1246 ( .A(n1062), .B(n1063), .Z(n61) );
  NANDN U1247 ( .A(B[72]), .B(n1064), .Z(n1063) );
  NANDN U1248 ( .A(A[72]), .B(n63), .Z(n1064) );
  NANDN U1249 ( .A(n63), .B(A[72]), .Z(n1062) );
  AND U1250 ( .A(n1065), .B(n1066), .Z(n63) );
  NANDN U1251 ( .A(B[71]), .B(n1067), .Z(n1066) );
  NANDN U1252 ( .A(A[71]), .B(n65), .Z(n1067) );
  NANDN U1253 ( .A(n65), .B(A[71]), .Z(n1065) );
  AND U1254 ( .A(n1068), .B(n1069), .Z(n65) );
  NANDN U1255 ( .A(B[70]), .B(n1070), .Z(n1069) );
  NANDN U1256 ( .A(A[70]), .B(n67), .Z(n1070) );
  NANDN U1257 ( .A(n67), .B(A[70]), .Z(n1068) );
  AND U1258 ( .A(n1071), .B(n1072), .Z(n67) );
  NANDN U1259 ( .A(B[69]), .B(n1073), .Z(n1072) );
  NANDN U1260 ( .A(A[69]), .B(n71), .Z(n1073) );
  NANDN U1261 ( .A(n71), .B(A[69]), .Z(n1071) );
  AND U1262 ( .A(n1074), .B(n1075), .Z(n71) );
  NANDN U1263 ( .A(B[68]), .B(n1076), .Z(n1075) );
  NANDN U1264 ( .A(A[68]), .B(n73), .Z(n1076) );
  NANDN U1265 ( .A(n73), .B(A[68]), .Z(n1074) );
  AND U1266 ( .A(n1077), .B(n1078), .Z(n73) );
  NANDN U1267 ( .A(B[67]), .B(n1079), .Z(n1078) );
  NANDN U1268 ( .A(A[67]), .B(n75), .Z(n1079) );
  NANDN U1269 ( .A(n75), .B(A[67]), .Z(n1077) );
  AND U1270 ( .A(n1080), .B(n1081), .Z(n75) );
  NANDN U1271 ( .A(B[66]), .B(n1082), .Z(n1081) );
  NANDN U1272 ( .A(A[66]), .B(n77), .Z(n1082) );
  NANDN U1273 ( .A(n77), .B(A[66]), .Z(n1080) );
  AND U1274 ( .A(n1083), .B(n1084), .Z(n77) );
  NANDN U1275 ( .A(B[65]), .B(n1085), .Z(n1084) );
  NANDN U1276 ( .A(A[65]), .B(n79), .Z(n1085) );
  NANDN U1277 ( .A(n79), .B(A[65]), .Z(n1083) );
  AND U1278 ( .A(n1086), .B(n1087), .Z(n79) );
  NANDN U1279 ( .A(B[64]), .B(n1088), .Z(n1087) );
  NANDN U1280 ( .A(A[64]), .B(n81), .Z(n1088) );
  NANDN U1281 ( .A(n81), .B(A[64]), .Z(n1086) );
  AND U1282 ( .A(n1089), .B(n1090), .Z(n81) );
  NANDN U1283 ( .A(B[63]), .B(n1091), .Z(n1090) );
  NANDN U1284 ( .A(A[63]), .B(n83), .Z(n1091) );
  NANDN U1285 ( .A(n83), .B(A[63]), .Z(n1089) );
  AND U1286 ( .A(n1092), .B(n1093), .Z(n83) );
  NANDN U1287 ( .A(B[62]), .B(n1094), .Z(n1093) );
  NANDN U1288 ( .A(A[62]), .B(n85), .Z(n1094) );
  NANDN U1289 ( .A(n85), .B(A[62]), .Z(n1092) );
  AND U1290 ( .A(n1095), .B(n1096), .Z(n85) );
  NANDN U1291 ( .A(B[61]), .B(n1097), .Z(n1096) );
  NANDN U1292 ( .A(A[61]), .B(n87), .Z(n1097) );
  NANDN U1293 ( .A(n87), .B(A[61]), .Z(n1095) );
  AND U1294 ( .A(n1098), .B(n1099), .Z(n87) );
  NANDN U1295 ( .A(B[60]), .B(n1100), .Z(n1099) );
  NANDN U1296 ( .A(A[60]), .B(n89), .Z(n1100) );
  NANDN U1297 ( .A(n89), .B(A[60]), .Z(n1098) );
  AND U1298 ( .A(n1101), .B(n1102), .Z(n89) );
  NANDN U1299 ( .A(B[59]), .B(n1103), .Z(n1102) );
  NANDN U1300 ( .A(A[59]), .B(n93), .Z(n1103) );
  NANDN U1301 ( .A(n93), .B(A[59]), .Z(n1101) );
  AND U1302 ( .A(n1104), .B(n1105), .Z(n93) );
  NANDN U1303 ( .A(B[58]), .B(n1106), .Z(n1105) );
  NANDN U1304 ( .A(A[58]), .B(n95), .Z(n1106) );
  NANDN U1305 ( .A(n95), .B(A[58]), .Z(n1104) );
  AND U1306 ( .A(n1107), .B(n1108), .Z(n95) );
  NANDN U1307 ( .A(B[57]), .B(n1109), .Z(n1108) );
  NANDN U1308 ( .A(A[57]), .B(n97), .Z(n1109) );
  NANDN U1309 ( .A(n97), .B(A[57]), .Z(n1107) );
  AND U1310 ( .A(n1110), .B(n1111), .Z(n97) );
  NANDN U1311 ( .A(B[56]), .B(n1112), .Z(n1111) );
  NANDN U1312 ( .A(A[56]), .B(n99), .Z(n1112) );
  NANDN U1313 ( .A(n99), .B(A[56]), .Z(n1110) );
  AND U1314 ( .A(n1113), .B(n1114), .Z(n99) );
  NANDN U1315 ( .A(B[55]), .B(n1115), .Z(n1114) );
  NANDN U1316 ( .A(A[55]), .B(n101), .Z(n1115) );
  NANDN U1317 ( .A(n101), .B(A[55]), .Z(n1113) );
  AND U1318 ( .A(n1116), .B(n1117), .Z(n101) );
  NANDN U1319 ( .A(B[54]), .B(n1118), .Z(n1117) );
  NANDN U1320 ( .A(A[54]), .B(n103), .Z(n1118) );
  NANDN U1321 ( .A(n103), .B(A[54]), .Z(n1116) );
  AND U1322 ( .A(n1119), .B(n1120), .Z(n103) );
  NANDN U1323 ( .A(B[53]), .B(n1121), .Z(n1120) );
  NANDN U1324 ( .A(A[53]), .B(n105), .Z(n1121) );
  NANDN U1325 ( .A(n105), .B(A[53]), .Z(n1119) );
  AND U1326 ( .A(n1122), .B(n1123), .Z(n105) );
  NANDN U1327 ( .A(B[52]), .B(n1124), .Z(n1123) );
  NANDN U1328 ( .A(A[52]), .B(n107), .Z(n1124) );
  NANDN U1329 ( .A(n107), .B(A[52]), .Z(n1122) );
  AND U1330 ( .A(n1125), .B(n1126), .Z(n107) );
  NANDN U1331 ( .A(B[51]), .B(n1127), .Z(n1126) );
  NANDN U1332 ( .A(A[51]), .B(n109), .Z(n1127) );
  NANDN U1333 ( .A(n109), .B(A[51]), .Z(n1125) );
  AND U1334 ( .A(n1128), .B(n1129), .Z(n109) );
  NANDN U1335 ( .A(B[50]), .B(n1130), .Z(n1129) );
  NANDN U1336 ( .A(A[50]), .B(n111), .Z(n1130) );
  NANDN U1337 ( .A(n111), .B(A[50]), .Z(n1128) );
  AND U1338 ( .A(n1131), .B(n1132), .Z(n111) );
  NANDN U1339 ( .A(B[49]), .B(n1133), .Z(n1132) );
  NANDN U1340 ( .A(A[49]), .B(n115), .Z(n1133) );
  NANDN U1341 ( .A(n115), .B(A[49]), .Z(n1131) );
  AND U1342 ( .A(n1134), .B(n1135), .Z(n115) );
  NANDN U1343 ( .A(B[48]), .B(n1136), .Z(n1135) );
  NANDN U1344 ( .A(A[48]), .B(n117), .Z(n1136) );
  NANDN U1345 ( .A(n117), .B(A[48]), .Z(n1134) );
  AND U1346 ( .A(n1137), .B(n1138), .Z(n117) );
  NANDN U1347 ( .A(B[47]), .B(n1139), .Z(n1138) );
  NANDN U1348 ( .A(A[47]), .B(n119), .Z(n1139) );
  NANDN U1349 ( .A(n119), .B(A[47]), .Z(n1137) );
  AND U1350 ( .A(n1140), .B(n1141), .Z(n119) );
  NANDN U1351 ( .A(B[46]), .B(n1142), .Z(n1141) );
  NANDN U1352 ( .A(A[46]), .B(n121), .Z(n1142) );
  NANDN U1353 ( .A(n121), .B(A[46]), .Z(n1140) );
  AND U1354 ( .A(n1143), .B(n1144), .Z(n121) );
  NANDN U1355 ( .A(B[45]), .B(n1145), .Z(n1144) );
  NANDN U1356 ( .A(A[45]), .B(n123), .Z(n1145) );
  NANDN U1357 ( .A(n123), .B(A[45]), .Z(n1143) );
  AND U1358 ( .A(n1146), .B(n1147), .Z(n123) );
  NANDN U1359 ( .A(B[44]), .B(n1148), .Z(n1147) );
  NANDN U1360 ( .A(A[44]), .B(n125), .Z(n1148) );
  NANDN U1361 ( .A(n125), .B(A[44]), .Z(n1146) );
  AND U1362 ( .A(n1149), .B(n1150), .Z(n125) );
  NANDN U1363 ( .A(B[43]), .B(n1151), .Z(n1150) );
  NANDN U1364 ( .A(A[43]), .B(n127), .Z(n1151) );
  NANDN U1365 ( .A(n127), .B(A[43]), .Z(n1149) );
  AND U1366 ( .A(n1152), .B(n1153), .Z(n127) );
  NANDN U1367 ( .A(B[42]), .B(n1154), .Z(n1153) );
  NANDN U1368 ( .A(A[42]), .B(n129), .Z(n1154) );
  NANDN U1369 ( .A(n129), .B(A[42]), .Z(n1152) );
  AND U1370 ( .A(n1155), .B(n1156), .Z(n129) );
  NANDN U1371 ( .A(B[41]), .B(n1157), .Z(n1156) );
  NANDN U1372 ( .A(A[41]), .B(n131), .Z(n1157) );
  NANDN U1373 ( .A(n131), .B(A[41]), .Z(n1155) );
  AND U1374 ( .A(n1158), .B(n1159), .Z(n131) );
  NANDN U1375 ( .A(B[40]), .B(n1160), .Z(n1159) );
  NANDN U1376 ( .A(A[40]), .B(n133), .Z(n1160) );
  NANDN U1377 ( .A(n133), .B(A[40]), .Z(n1158) );
  AND U1378 ( .A(n1161), .B(n1162), .Z(n133) );
  NANDN U1379 ( .A(B[39]), .B(n1163), .Z(n1162) );
  NANDN U1380 ( .A(A[39]), .B(n137), .Z(n1163) );
  NANDN U1381 ( .A(n137), .B(A[39]), .Z(n1161) );
  AND U1382 ( .A(n1164), .B(n1165), .Z(n137) );
  NANDN U1383 ( .A(B[38]), .B(n1166), .Z(n1165) );
  NANDN U1384 ( .A(A[38]), .B(n139), .Z(n1166) );
  NANDN U1385 ( .A(n139), .B(A[38]), .Z(n1164) );
  AND U1386 ( .A(n1167), .B(n1168), .Z(n139) );
  NANDN U1387 ( .A(B[37]), .B(n1169), .Z(n1168) );
  NANDN U1388 ( .A(A[37]), .B(n141), .Z(n1169) );
  NANDN U1389 ( .A(n141), .B(A[37]), .Z(n1167) );
  AND U1390 ( .A(n1170), .B(n1171), .Z(n141) );
  NANDN U1391 ( .A(B[36]), .B(n1172), .Z(n1171) );
  NANDN U1392 ( .A(A[36]), .B(n143), .Z(n1172) );
  NANDN U1393 ( .A(n143), .B(A[36]), .Z(n1170) );
  AND U1394 ( .A(n1173), .B(n1174), .Z(n143) );
  NANDN U1395 ( .A(B[35]), .B(n1175), .Z(n1174) );
  NANDN U1396 ( .A(A[35]), .B(n145), .Z(n1175) );
  NANDN U1397 ( .A(n145), .B(A[35]), .Z(n1173) );
  AND U1398 ( .A(n1176), .B(n1177), .Z(n145) );
  NANDN U1399 ( .A(B[34]), .B(n1178), .Z(n1177) );
  NANDN U1400 ( .A(A[34]), .B(n147), .Z(n1178) );
  NANDN U1401 ( .A(n147), .B(A[34]), .Z(n1176) );
  AND U1402 ( .A(n1179), .B(n1180), .Z(n147) );
  NANDN U1403 ( .A(B[33]), .B(n1181), .Z(n1180) );
  NANDN U1404 ( .A(A[33]), .B(n149), .Z(n1181) );
  NANDN U1405 ( .A(n149), .B(A[33]), .Z(n1179) );
  AND U1406 ( .A(n1182), .B(n1183), .Z(n149) );
  NANDN U1407 ( .A(B[32]), .B(n1184), .Z(n1183) );
  NANDN U1408 ( .A(A[32]), .B(n151), .Z(n1184) );
  NANDN U1409 ( .A(n151), .B(A[32]), .Z(n1182) );
  AND U1410 ( .A(n1185), .B(n1186), .Z(n151) );
  NANDN U1411 ( .A(B[31]), .B(n1187), .Z(n1186) );
  NANDN U1412 ( .A(A[31]), .B(n153), .Z(n1187) );
  NANDN U1413 ( .A(n153), .B(A[31]), .Z(n1185) );
  AND U1414 ( .A(n1188), .B(n1189), .Z(n153) );
  NANDN U1415 ( .A(B[30]), .B(n1190), .Z(n1189) );
  NANDN U1416 ( .A(A[30]), .B(n155), .Z(n1190) );
  NANDN U1417 ( .A(n155), .B(A[30]), .Z(n1188) );
  AND U1418 ( .A(n1191), .B(n1192), .Z(n155) );
  NANDN U1419 ( .A(B[29]), .B(n1193), .Z(n1192) );
  NANDN U1420 ( .A(A[29]), .B(n159), .Z(n1193) );
  NANDN U1421 ( .A(n159), .B(A[29]), .Z(n1191) );
  AND U1422 ( .A(n1194), .B(n1195), .Z(n159) );
  NANDN U1423 ( .A(B[28]), .B(n1196), .Z(n1195) );
  NANDN U1424 ( .A(A[28]), .B(n161), .Z(n1196) );
  NANDN U1425 ( .A(n161), .B(A[28]), .Z(n1194) );
  AND U1426 ( .A(n1197), .B(n1198), .Z(n161) );
  NANDN U1427 ( .A(B[27]), .B(n1199), .Z(n1198) );
  NANDN U1428 ( .A(A[27]), .B(n163), .Z(n1199) );
  NANDN U1429 ( .A(n163), .B(A[27]), .Z(n1197) );
  AND U1430 ( .A(n1200), .B(n1201), .Z(n163) );
  NANDN U1431 ( .A(B[26]), .B(n1202), .Z(n1201) );
  NANDN U1432 ( .A(A[26]), .B(n165), .Z(n1202) );
  NANDN U1433 ( .A(n165), .B(A[26]), .Z(n1200) );
  AND U1434 ( .A(n1203), .B(n1204), .Z(n165) );
  NANDN U1435 ( .A(B[25]), .B(n1205), .Z(n1204) );
  NANDN U1436 ( .A(A[25]), .B(n167), .Z(n1205) );
  NANDN U1437 ( .A(n167), .B(A[25]), .Z(n1203) );
  AND U1438 ( .A(n1206), .B(n1207), .Z(n167) );
  NANDN U1439 ( .A(B[24]), .B(n1208), .Z(n1207) );
  NANDN U1440 ( .A(A[24]), .B(n204), .Z(n1208) );
  NANDN U1441 ( .A(n204), .B(A[24]), .Z(n1206) );
  AND U1442 ( .A(n1209), .B(n1210), .Z(n204) );
  NANDN U1443 ( .A(B[23]), .B(n1211), .Z(n1210) );
  NANDN U1444 ( .A(A[23]), .B(n256), .Z(n1211) );
  NANDN U1445 ( .A(n256), .B(A[23]), .Z(n1209) );
  AND U1446 ( .A(n1212), .B(n1213), .Z(n256) );
  NANDN U1447 ( .A(B[22]), .B(n1214), .Z(n1213) );
  NANDN U1448 ( .A(A[22]), .B(n308), .Z(n1214) );
  NANDN U1449 ( .A(n308), .B(A[22]), .Z(n1212) );
  AND U1450 ( .A(n1215), .B(n1216), .Z(n308) );
  NANDN U1451 ( .A(B[21]), .B(n1217), .Z(n1216) );
  NANDN U1452 ( .A(A[21]), .B(n360), .Z(n1217) );
  NANDN U1453 ( .A(n360), .B(A[21]), .Z(n1215) );
  AND U1454 ( .A(n1218), .B(n1219), .Z(n360) );
  NANDN U1455 ( .A(B[20]), .B(n1220), .Z(n1219) );
  NANDN U1456 ( .A(A[20]), .B(n412), .Z(n1220) );
  NANDN U1457 ( .A(n412), .B(A[20]), .Z(n1218) );
  AND U1458 ( .A(n1221), .B(n1222), .Z(n412) );
  NANDN U1459 ( .A(B[19]), .B(n1223), .Z(n1222) );
  NANDN U1460 ( .A(A[19]), .B(n465), .Z(n1223) );
  NANDN U1461 ( .A(n465), .B(A[19]), .Z(n1221) );
  AND U1462 ( .A(n1224), .B(n1225), .Z(n465) );
  NANDN U1463 ( .A(B[18]), .B(n1226), .Z(n1225) );
  NANDN U1464 ( .A(A[18]), .B(n517), .Z(n1226) );
  NANDN U1465 ( .A(n517), .B(A[18]), .Z(n1224) );
  AND U1466 ( .A(n1227), .B(n1228), .Z(n517) );
  NANDN U1467 ( .A(B[17]), .B(n1229), .Z(n1228) );
  NANDN U1468 ( .A(A[17]), .B(n569), .Z(n1229) );
  NANDN U1469 ( .A(n569), .B(A[17]), .Z(n1227) );
  AND U1470 ( .A(n1230), .B(n1231), .Z(n569) );
  NANDN U1471 ( .A(B[16]), .B(n1232), .Z(n1231) );
  NANDN U1472 ( .A(A[16]), .B(n621), .Z(n1232) );
  NANDN U1473 ( .A(n621), .B(A[16]), .Z(n1230) );
  AND U1474 ( .A(n1233), .B(n1234), .Z(n621) );
  NANDN U1475 ( .A(B[15]), .B(n1235), .Z(n1234) );
  NANDN U1476 ( .A(A[15]), .B(n673), .Z(n1235) );
  NANDN U1477 ( .A(n673), .B(A[15]), .Z(n1233) );
  AND U1478 ( .A(n1236), .B(n1237), .Z(n673) );
  NANDN U1479 ( .A(B[14]), .B(n1238), .Z(n1237) );
  NANDN U1480 ( .A(A[14]), .B(n725), .Z(n1238) );
  NANDN U1481 ( .A(n725), .B(A[14]), .Z(n1236) );
  AND U1482 ( .A(n1239), .B(n1240), .Z(n725) );
  NANDN U1483 ( .A(B[13]), .B(n1241), .Z(n1240) );
  NANDN U1484 ( .A(A[13]), .B(n777), .Z(n1241) );
  NANDN U1485 ( .A(n777), .B(A[13]), .Z(n1239) );
  AND U1486 ( .A(n1242), .B(n1243), .Z(n777) );
  NANDN U1487 ( .A(B[12]), .B(n1244), .Z(n1243) );
  NANDN U1488 ( .A(A[12]), .B(n829), .Z(n1244) );
  NANDN U1489 ( .A(n829), .B(A[12]), .Z(n1242) );
  AND U1490 ( .A(n1245), .B(n1246), .Z(n829) );
  NANDN U1491 ( .A(B[11]), .B(n1247), .Z(n1246) );
  NANDN U1492 ( .A(A[11]), .B(n881), .Z(n1247) );
  NANDN U1493 ( .A(n881), .B(A[11]), .Z(n1245) );
  AND U1494 ( .A(n1248), .B(n1249), .Z(n881) );
  NANDN U1495 ( .A(B[10]), .B(n1250), .Z(n1249) );
  NANDN U1496 ( .A(A[10]), .B(n933), .Z(n1250) );
  NANDN U1497 ( .A(n933), .B(A[10]), .Z(n1248) );
  AND U1498 ( .A(n1251), .B(n1252), .Z(n933) );
  NANDN U1499 ( .A(B[9]), .B(n1253), .Z(n1252) );
  OR U1500 ( .A(n3), .B(A[9]), .Z(n1253) );
  NAND U1501 ( .A(A[9]), .B(n3), .Z(n1251) );
  NAND U1502 ( .A(n1254), .B(n1255), .Z(n3) );
  NANDN U1503 ( .A(B[8]), .B(n1256), .Z(n1255) );
  NANDN U1504 ( .A(A[8]), .B(n25), .Z(n1256) );
  NANDN U1505 ( .A(n25), .B(A[8]), .Z(n1254) );
  AND U1506 ( .A(n1257), .B(n1258), .Z(n25) );
  NANDN U1507 ( .A(B[7]), .B(n1259), .Z(n1258) );
  NANDN U1508 ( .A(A[7]), .B(n47), .Z(n1259) );
  NANDN U1509 ( .A(n47), .B(A[7]), .Z(n1257) );
  AND U1510 ( .A(n1260), .B(n1261), .Z(n47) );
  NANDN U1511 ( .A(B[6]), .B(n1262), .Z(n1261) );
  NANDN U1512 ( .A(A[6]), .B(n69), .Z(n1262) );
  NANDN U1513 ( .A(n69), .B(A[6]), .Z(n1260) );
  AND U1514 ( .A(n1263), .B(n1264), .Z(n69) );
  NANDN U1515 ( .A(B[5]), .B(n1265), .Z(n1264) );
  NANDN U1516 ( .A(A[5]), .B(n91), .Z(n1265) );
  NANDN U1517 ( .A(n91), .B(A[5]), .Z(n1263) );
  AND U1518 ( .A(n1266), .B(n1267), .Z(n91) );
  NANDN U1519 ( .A(B[4]), .B(n1268), .Z(n1267) );
  NANDN U1520 ( .A(A[4]), .B(n113), .Z(n1268) );
  NANDN U1521 ( .A(n113), .B(A[4]), .Z(n1266) );
  AND U1522 ( .A(n1269), .B(n1270), .Z(n113) );
  NANDN U1523 ( .A(B[3]), .B(n1271), .Z(n1270) );
  NANDN U1524 ( .A(A[3]), .B(n135), .Z(n1271) );
  NANDN U1525 ( .A(n135), .B(A[3]), .Z(n1269) );
  AND U1526 ( .A(n1272), .B(n1273), .Z(n135) );
  NANDN U1527 ( .A(B[2]), .B(n1274), .Z(n1273) );
  NANDN U1528 ( .A(A[2]), .B(n157), .Z(n1274) );
  NANDN U1529 ( .A(n157), .B(A[2]), .Z(n1272) );
  AND U1530 ( .A(n1275), .B(n1276), .Z(n157) );
  NANDN U1531 ( .A(B[1]), .B(n1277), .Z(n1276) );
  NAND U1532 ( .A(n1), .B(n2), .Z(n1277) );
  NAND U1533 ( .A(A[1]), .B(n1278), .Z(n1275) );
  NAND U1534 ( .A(n1278), .B(n1279), .Z(DIFF[0]) );
  NANDN U1535 ( .A(B[0]), .B(A[0]), .Z(n1279) );
  NANDN U1536 ( .A(A[0]), .B(B[0]), .Z(n1278) );
endmodule


module modmult_step_N256_4_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [255:0] A;
  input [0:0] B;
  output [256:0] PRODUCT;
  input TC;


  AND U2 ( .A(A[255]), .B(B[0]), .Z(PRODUCT[255]) );
  AND U3 ( .A(A[254]), .B(B[0]), .Z(PRODUCT[254]) );
  AND U4 ( .A(A[253]), .B(B[0]), .Z(PRODUCT[253]) );
  AND U5 ( .A(A[252]), .B(B[0]), .Z(PRODUCT[252]) );
  AND U6 ( .A(A[251]), .B(B[0]), .Z(PRODUCT[251]) );
  AND U7 ( .A(A[250]), .B(B[0]), .Z(PRODUCT[250]) );
  AND U8 ( .A(A[249]), .B(B[0]), .Z(PRODUCT[249]) );
  AND U9 ( .A(A[248]), .B(B[0]), .Z(PRODUCT[248]) );
  AND U10 ( .A(A[247]), .B(B[0]), .Z(PRODUCT[247]) );
  AND U11 ( .A(A[246]), .B(B[0]), .Z(PRODUCT[246]) );
  AND U12 ( .A(A[245]), .B(B[0]), .Z(PRODUCT[245]) );
  AND U13 ( .A(A[244]), .B(B[0]), .Z(PRODUCT[244]) );
  AND U14 ( .A(A[243]), .B(B[0]), .Z(PRODUCT[243]) );
  AND U15 ( .A(A[242]), .B(B[0]), .Z(PRODUCT[242]) );
  AND U16 ( .A(A[241]), .B(B[0]), .Z(PRODUCT[241]) );
  AND U17 ( .A(A[240]), .B(B[0]), .Z(PRODUCT[240]) );
  AND U18 ( .A(A[239]), .B(B[0]), .Z(PRODUCT[239]) );
  AND U19 ( .A(A[238]), .B(B[0]), .Z(PRODUCT[238]) );
  AND U20 ( .A(A[237]), .B(B[0]), .Z(PRODUCT[237]) );
  AND U21 ( .A(A[236]), .B(B[0]), .Z(PRODUCT[236]) );
  AND U22 ( .A(A[235]), .B(B[0]), .Z(PRODUCT[235]) );
  AND U23 ( .A(A[234]), .B(B[0]), .Z(PRODUCT[234]) );
  AND U24 ( .A(A[233]), .B(B[0]), .Z(PRODUCT[233]) );
  AND U25 ( .A(A[232]), .B(B[0]), .Z(PRODUCT[232]) );
  AND U26 ( .A(A[231]), .B(B[0]), .Z(PRODUCT[231]) );
  AND U27 ( .A(A[230]), .B(B[0]), .Z(PRODUCT[230]) );
  AND U28 ( .A(A[229]), .B(B[0]), .Z(PRODUCT[229]) );
  AND U29 ( .A(A[228]), .B(B[0]), .Z(PRODUCT[228]) );
  AND U30 ( .A(A[227]), .B(B[0]), .Z(PRODUCT[227]) );
  AND U31 ( .A(A[226]), .B(B[0]), .Z(PRODUCT[226]) );
  AND U32 ( .A(A[225]), .B(B[0]), .Z(PRODUCT[225]) );
  AND U33 ( .A(A[224]), .B(B[0]), .Z(PRODUCT[224]) );
  AND U34 ( .A(A[223]), .B(B[0]), .Z(PRODUCT[223]) );
  AND U35 ( .A(A[222]), .B(B[0]), .Z(PRODUCT[222]) );
  AND U36 ( .A(A[221]), .B(B[0]), .Z(PRODUCT[221]) );
  AND U37 ( .A(A[220]), .B(B[0]), .Z(PRODUCT[220]) );
  AND U38 ( .A(A[219]), .B(B[0]), .Z(PRODUCT[219]) );
  AND U39 ( .A(A[218]), .B(B[0]), .Z(PRODUCT[218]) );
  AND U40 ( .A(A[217]), .B(B[0]), .Z(PRODUCT[217]) );
  AND U41 ( .A(A[216]), .B(B[0]), .Z(PRODUCT[216]) );
  AND U42 ( .A(A[215]), .B(B[0]), .Z(PRODUCT[215]) );
  AND U43 ( .A(A[214]), .B(B[0]), .Z(PRODUCT[214]) );
  AND U44 ( .A(A[213]), .B(B[0]), .Z(PRODUCT[213]) );
  AND U45 ( .A(A[212]), .B(B[0]), .Z(PRODUCT[212]) );
  AND U46 ( .A(A[211]), .B(B[0]), .Z(PRODUCT[211]) );
  AND U47 ( .A(A[210]), .B(B[0]), .Z(PRODUCT[210]) );
  AND U48 ( .A(A[209]), .B(B[0]), .Z(PRODUCT[209]) );
  AND U49 ( .A(A[208]), .B(B[0]), .Z(PRODUCT[208]) );
  AND U50 ( .A(A[207]), .B(B[0]), .Z(PRODUCT[207]) );
  AND U51 ( .A(A[206]), .B(B[0]), .Z(PRODUCT[206]) );
  AND U52 ( .A(A[205]), .B(B[0]), .Z(PRODUCT[205]) );
  AND U53 ( .A(A[204]), .B(B[0]), .Z(PRODUCT[204]) );
  AND U54 ( .A(A[203]), .B(B[0]), .Z(PRODUCT[203]) );
  AND U55 ( .A(A[202]), .B(B[0]), .Z(PRODUCT[202]) );
  AND U56 ( .A(A[201]), .B(B[0]), .Z(PRODUCT[201]) );
  AND U57 ( .A(A[200]), .B(B[0]), .Z(PRODUCT[200]) );
  AND U58 ( .A(A[199]), .B(B[0]), .Z(PRODUCT[199]) );
  AND U59 ( .A(A[198]), .B(B[0]), .Z(PRODUCT[198]) );
  AND U60 ( .A(A[197]), .B(B[0]), .Z(PRODUCT[197]) );
  AND U61 ( .A(A[196]), .B(B[0]), .Z(PRODUCT[196]) );
  AND U62 ( .A(A[195]), .B(B[0]), .Z(PRODUCT[195]) );
  AND U63 ( .A(A[194]), .B(B[0]), .Z(PRODUCT[194]) );
  AND U64 ( .A(A[193]), .B(B[0]), .Z(PRODUCT[193]) );
  AND U65 ( .A(A[192]), .B(B[0]), .Z(PRODUCT[192]) );
  AND U66 ( .A(A[191]), .B(B[0]), .Z(PRODUCT[191]) );
  AND U67 ( .A(A[190]), .B(B[0]), .Z(PRODUCT[190]) );
  AND U68 ( .A(A[189]), .B(B[0]), .Z(PRODUCT[189]) );
  AND U69 ( .A(A[188]), .B(B[0]), .Z(PRODUCT[188]) );
  AND U70 ( .A(A[187]), .B(B[0]), .Z(PRODUCT[187]) );
  AND U71 ( .A(A[186]), .B(B[0]), .Z(PRODUCT[186]) );
  AND U72 ( .A(A[185]), .B(B[0]), .Z(PRODUCT[185]) );
  AND U73 ( .A(A[184]), .B(B[0]), .Z(PRODUCT[184]) );
  AND U74 ( .A(A[183]), .B(B[0]), .Z(PRODUCT[183]) );
  AND U75 ( .A(A[182]), .B(B[0]), .Z(PRODUCT[182]) );
  AND U76 ( .A(A[181]), .B(B[0]), .Z(PRODUCT[181]) );
  AND U77 ( .A(A[180]), .B(B[0]), .Z(PRODUCT[180]) );
  AND U78 ( .A(A[179]), .B(B[0]), .Z(PRODUCT[179]) );
  AND U79 ( .A(A[178]), .B(B[0]), .Z(PRODUCT[178]) );
  AND U80 ( .A(A[177]), .B(B[0]), .Z(PRODUCT[177]) );
  AND U81 ( .A(A[176]), .B(B[0]), .Z(PRODUCT[176]) );
  AND U82 ( .A(A[175]), .B(B[0]), .Z(PRODUCT[175]) );
  AND U83 ( .A(A[174]), .B(B[0]), .Z(PRODUCT[174]) );
  AND U84 ( .A(A[173]), .B(B[0]), .Z(PRODUCT[173]) );
  AND U85 ( .A(A[172]), .B(B[0]), .Z(PRODUCT[172]) );
  AND U86 ( .A(A[171]), .B(B[0]), .Z(PRODUCT[171]) );
  AND U87 ( .A(A[170]), .B(B[0]), .Z(PRODUCT[170]) );
  AND U88 ( .A(A[169]), .B(B[0]), .Z(PRODUCT[169]) );
  AND U89 ( .A(A[168]), .B(B[0]), .Z(PRODUCT[168]) );
  AND U90 ( .A(A[167]), .B(B[0]), .Z(PRODUCT[167]) );
  AND U91 ( .A(A[166]), .B(B[0]), .Z(PRODUCT[166]) );
  AND U92 ( .A(A[165]), .B(B[0]), .Z(PRODUCT[165]) );
  AND U93 ( .A(A[164]), .B(B[0]), .Z(PRODUCT[164]) );
  AND U94 ( .A(A[163]), .B(B[0]), .Z(PRODUCT[163]) );
  AND U95 ( .A(A[162]), .B(B[0]), .Z(PRODUCT[162]) );
  AND U96 ( .A(A[161]), .B(B[0]), .Z(PRODUCT[161]) );
  AND U97 ( .A(A[160]), .B(B[0]), .Z(PRODUCT[160]) );
  AND U98 ( .A(A[159]), .B(B[0]), .Z(PRODUCT[159]) );
  AND U99 ( .A(A[158]), .B(B[0]), .Z(PRODUCT[158]) );
  AND U100 ( .A(A[157]), .B(B[0]), .Z(PRODUCT[157]) );
  AND U101 ( .A(A[156]), .B(B[0]), .Z(PRODUCT[156]) );
  AND U102 ( .A(A[155]), .B(B[0]), .Z(PRODUCT[155]) );
  AND U103 ( .A(A[154]), .B(B[0]), .Z(PRODUCT[154]) );
  AND U104 ( .A(A[153]), .B(B[0]), .Z(PRODUCT[153]) );
  AND U105 ( .A(A[152]), .B(B[0]), .Z(PRODUCT[152]) );
  AND U106 ( .A(A[151]), .B(B[0]), .Z(PRODUCT[151]) );
  AND U107 ( .A(A[150]), .B(B[0]), .Z(PRODUCT[150]) );
  AND U108 ( .A(A[149]), .B(B[0]), .Z(PRODUCT[149]) );
  AND U109 ( .A(A[148]), .B(B[0]), .Z(PRODUCT[148]) );
  AND U110 ( .A(A[147]), .B(B[0]), .Z(PRODUCT[147]) );
  AND U111 ( .A(A[146]), .B(B[0]), .Z(PRODUCT[146]) );
  AND U112 ( .A(A[145]), .B(B[0]), .Z(PRODUCT[145]) );
  AND U113 ( .A(A[144]), .B(B[0]), .Z(PRODUCT[144]) );
  AND U114 ( .A(A[143]), .B(B[0]), .Z(PRODUCT[143]) );
  AND U115 ( .A(A[142]), .B(B[0]), .Z(PRODUCT[142]) );
  AND U116 ( .A(A[141]), .B(B[0]), .Z(PRODUCT[141]) );
  AND U117 ( .A(A[140]), .B(B[0]), .Z(PRODUCT[140]) );
  AND U118 ( .A(A[139]), .B(B[0]), .Z(PRODUCT[139]) );
  AND U119 ( .A(A[138]), .B(B[0]), .Z(PRODUCT[138]) );
  AND U120 ( .A(A[137]), .B(B[0]), .Z(PRODUCT[137]) );
  AND U121 ( .A(A[136]), .B(B[0]), .Z(PRODUCT[136]) );
  AND U122 ( .A(A[135]), .B(B[0]), .Z(PRODUCT[135]) );
  AND U123 ( .A(A[134]), .B(B[0]), .Z(PRODUCT[134]) );
  AND U124 ( .A(A[133]), .B(B[0]), .Z(PRODUCT[133]) );
  AND U125 ( .A(A[132]), .B(B[0]), .Z(PRODUCT[132]) );
  AND U126 ( .A(A[131]), .B(B[0]), .Z(PRODUCT[131]) );
  AND U127 ( .A(A[130]), .B(B[0]), .Z(PRODUCT[130]) );
  AND U128 ( .A(A[129]), .B(B[0]), .Z(PRODUCT[129]) );
  AND U129 ( .A(A[128]), .B(B[0]), .Z(PRODUCT[128]) );
  AND U130 ( .A(A[127]), .B(B[0]), .Z(PRODUCT[127]) );
  AND U131 ( .A(A[126]), .B(B[0]), .Z(PRODUCT[126]) );
  AND U132 ( .A(A[125]), .B(B[0]), .Z(PRODUCT[125]) );
  AND U133 ( .A(A[124]), .B(B[0]), .Z(PRODUCT[124]) );
  AND U134 ( .A(A[123]), .B(B[0]), .Z(PRODUCT[123]) );
  AND U135 ( .A(A[122]), .B(B[0]), .Z(PRODUCT[122]) );
  AND U136 ( .A(A[121]), .B(B[0]), .Z(PRODUCT[121]) );
  AND U137 ( .A(A[120]), .B(B[0]), .Z(PRODUCT[120]) );
  AND U138 ( .A(A[119]), .B(B[0]), .Z(PRODUCT[119]) );
  AND U139 ( .A(A[118]), .B(B[0]), .Z(PRODUCT[118]) );
  AND U140 ( .A(A[117]), .B(B[0]), .Z(PRODUCT[117]) );
  AND U141 ( .A(A[116]), .B(B[0]), .Z(PRODUCT[116]) );
  AND U142 ( .A(A[115]), .B(B[0]), .Z(PRODUCT[115]) );
  AND U143 ( .A(A[114]), .B(B[0]), .Z(PRODUCT[114]) );
  AND U144 ( .A(A[113]), .B(B[0]), .Z(PRODUCT[113]) );
  AND U145 ( .A(A[112]), .B(B[0]), .Z(PRODUCT[112]) );
  AND U146 ( .A(A[111]), .B(B[0]), .Z(PRODUCT[111]) );
  AND U147 ( .A(A[110]), .B(B[0]), .Z(PRODUCT[110]) );
  AND U148 ( .A(A[109]), .B(B[0]), .Z(PRODUCT[109]) );
  AND U149 ( .A(A[108]), .B(B[0]), .Z(PRODUCT[108]) );
  AND U150 ( .A(A[107]), .B(B[0]), .Z(PRODUCT[107]) );
  AND U151 ( .A(A[106]), .B(B[0]), .Z(PRODUCT[106]) );
  AND U152 ( .A(A[105]), .B(B[0]), .Z(PRODUCT[105]) );
  AND U153 ( .A(A[104]), .B(B[0]), .Z(PRODUCT[104]) );
  AND U154 ( .A(A[103]), .B(B[0]), .Z(PRODUCT[103]) );
  AND U155 ( .A(A[102]), .B(B[0]), .Z(PRODUCT[102]) );
  AND U156 ( .A(A[101]), .B(B[0]), .Z(PRODUCT[101]) );
  AND U157 ( .A(A[100]), .B(B[0]), .Z(PRODUCT[100]) );
  AND U158 ( .A(A[99]), .B(B[0]), .Z(PRODUCT[99]) );
  AND U159 ( .A(A[98]), .B(B[0]), .Z(PRODUCT[98]) );
  AND U160 ( .A(A[97]), .B(B[0]), .Z(PRODUCT[97]) );
  AND U161 ( .A(A[96]), .B(B[0]), .Z(PRODUCT[96]) );
  AND U162 ( .A(A[95]), .B(B[0]), .Z(PRODUCT[95]) );
  AND U163 ( .A(A[94]), .B(B[0]), .Z(PRODUCT[94]) );
  AND U164 ( .A(A[93]), .B(B[0]), .Z(PRODUCT[93]) );
  AND U165 ( .A(A[92]), .B(B[0]), .Z(PRODUCT[92]) );
  AND U166 ( .A(A[91]), .B(B[0]), .Z(PRODUCT[91]) );
  AND U167 ( .A(A[90]), .B(B[0]), .Z(PRODUCT[90]) );
  AND U168 ( .A(A[89]), .B(B[0]), .Z(PRODUCT[89]) );
  AND U169 ( .A(A[88]), .B(B[0]), .Z(PRODUCT[88]) );
  AND U170 ( .A(A[87]), .B(B[0]), .Z(PRODUCT[87]) );
  AND U171 ( .A(A[86]), .B(B[0]), .Z(PRODUCT[86]) );
  AND U172 ( .A(A[85]), .B(B[0]), .Z(PRODUCT[85]) );
  AND U173 ( .A(A[84]), .B(B[0]), .Z(PRODUCT[84]) );
  AND U174 ( .A(A[83]), .B(B[0]), .Z(PRODUCT[83]) );
  AND U175 ( .A(A[82]), .B(B[0]), .Z(PRODUCT[82]) );
  AND U176 ( .A(A[81]), .B(B[0]), .Z(PRODUCT[81]) );
  AND U177 ( .A(A[80]), .B(B[0]), .Z(PRODUCT[80]) );
  AND U178 ( .A(A[79]), .B(B[0]), .Z(PRODUCT[79]) );
  AND U179 ( .A(A[78]), .B(B[0]), .Z(PRODUCT[78]) );
  AND U180 ( .A(A[77]), .B(B[0]), .Z(PRODUCT[77]) );
  AND U181 ( .A(A[76]), .B(B[0]), .Z(PRODUCT[76]) );
  AND U182 ( .A(A[75]), .B(B[0]), .Z(PRODUCT[75]) );
  AND U183 ( .A(A[74]), .B(B[0]), .Z(PRODUCT[74]) );
  AND U184 ( .A(A[73]), .B(B[0]), .Z(PRODUCT[73]) );
  AND U185 ( .A(A[72]), .B(B[0]), .Z(PRODUCT[72]) );
  AND U186 ( .A(A[71]), .B(B[0]), .Z(PRODUCT[71]) );
  AND U187 ( .A(A[70]), .B(B[0]), .Z(PRODUCT[70]) );
  AND U188 ( .A(A[69]), .B(B[0]), .Z(PRODUCT[69]) );
  AND U189 ( .A(A[68]), .B(B[0]), .Z(PRODUCT[68]) );
  AND U190 ( .A(A[67]), .B(B[0]), .Z(PRODUCT[67]) );
  AND U191 ( .A(A[66]), .B(B[0]), .Z(PRODUCT[66]) );
  AND U192 ( .A(A[65]), .B(B[0]), .Z(PRODUCT[65]) );
  AND U193 ( .A(A[64]), .B(B[0]), .Z(PRODUCT[64]) );
  AND U194 ( .A(A[63]), .B(B[0]), .Z(PRODUCT[63]) );
  AND U195 ( .A(A[62]), .B(B[0]), .Z(PRODUCT[62]) );
  AND U196 ( .A(A[61]), .B(B[0]), .Z(PRODUCT[61]) );
  AND U197 ( .A(A[60]), .B(B[0]), .Z(PRODUCT[60]) );
  AND U198 ( .A(A[59]), .B(B[0]), .Z(PRODUCT[59]) );
  AND U199 ( .A(A[58]), .B(B[0]), .Z(PRODUCT[58]) );
  AND U200 ( .A(A[57]), .B(B[0]), .Z(PRODUCT[57]) );
  AND U201 ( .A(A[56]), .B(B[0]), .Z(PRODUCT[56]) );
  AND U202 ( .A(A[55]), .B(B[0]), .Z(PRODUCT[55]) );
  AND U203 ( .A(A[54]), .B(B[0]), .Z(PRODUCT[54]) );
  AND U204 ( .A(A[53]), .B(B[0]), .Z(PRODUCT[53]) );
  AND U205 ( .A(A[52]), .B(B[0]), .Z(PRODUCT[52]) );
  AND U206 ( .A(A[51]), .B(B[0]), .Z(PRODUCT[51]) );
  AND U207 ( .A(A[50]), .B(B[0]), .Z(PRODUCT[50]) );
  AND U208 ( .A(A[49]), .B(B[0]), .Z(PRODUCT[49]) );
  AND U209 ( .A(A[48]), .B(B[0]), .Z(PRODUCT[48]) );
  AND U210 ( .A(A[47]), .B(B[0]), .Z(PRODUCT[47]) );
  AND U211 ( .A(A[46]), .B(B[0]), .Z(PRODUCT[46]) );
  AND U212 ( .A(A[45]), .B(B[0]), .Z(PRODUCT[45]) );
  AND U213 ( .A(A[44]), .B(B[0]), .Z(PRODUCT[44]) );
  AND U214 ( .A(A[43]), .B(B[0]), .Z(PRODUCT[43]) );
  AND U215 ( .A(A[42]), .B(B[0]), .Z(PRODUCT[42]) );
  AND U216 ( .A(A[41]), .B(B[0]), .Z(PRODUCT[41]) );
  AND U217 ( .A(A[40]), .B(B[0]), .Z(PRODUCT[40]) );
  AND U218 ( .A(A[39]), .B(B[0]), .Z(PRODUCT[39]) );
  AND U219 ( .A(A[38]), .B(B[0]), .Z(PRODUCT[38]) );
  AND U220 ( .A(A[37]), .B(B[0]), .Z(PRODUCT[37]) );
  AND U221 ( .A(A[36]), .B(B[0]), .Z(PRODUCT[36]) );
  AND U222 ( .A(A[35]), .B(B[0]), .Z(PRODUCT[35]) );
  AND U223 ( .A(A[34]), .B(B[0]), .Z(PRODUCT[34]) );
  AND U224 ( .A(A[33]), .B(B[0]), .Z(PRODUCT[33]) );
  AND U225 ( .A(A[32]), .B(B[0]), .Z(PRODUCT[32]) );
  AND U226 ( .A(A[31]), .B(B[0]), .Z(PRODUCT[31]) );
  AND U227 ( .A(A[30]), .B(B[0]), .Z(PRODUCT[30]) );
  AND U228 ( .A(A[29]), .B(B[0]), .Z(PRODUCT[29]) );
  AND U229 ( .A(A[28]), .B(B[0]), .Z(PRODUCT[28]) );
  AND U230 ( .A(A[27]), .B(B[0]), .Z(PRODUCT[27]) );
  AND U231 ( .A(A[26]), .B(B[0]), .Z(PRODUCT[26]) );
  AND U232 ( .A(A[25]), .B(B[0]), .Z(PRODUCT[25]) );
  AND U233 ( .A(A[24]), .B(B[0]), .Z(PRODUCT[24]) );
  AND U234 ( .A(A[23]), .B(B[0]), .Z(PRODUCT[23]) );
  AND U235 ( .A(A[22]), .B(B[0]), .Z(PRODUCT[22]) );
  AND U236 ( .A(A[21]), .B(B[0]), .Z(PRODUCT[21]) );
  AND U237 ( .A(A[20]), .B(B[0]), .Z(PRODUCT[20]) );
  AND U238 ( .A(A[19]), .B(B[0]), .Z(PRODUCT[19]) );
  AND U239 ( .A(A[18]), .B(B[0]), .Z(PRODUCT[18]) );
  AND U240 ( .A(A[17]), .B(B[0]), .Z(PRODUCT[17]) );
  AND U241 ( .A(A[16]), .B(B[0]), .Z(PRODUCT[16]) );
  AND U242 ( .A(A[15]), .B(B[0]), .Z(PRODUCT[15]) );
  AND U243 ( .A(A[14]), .B(B[0]), .Z(PRODUCT[14]) );
  AND U244 ( .A(A[13]), .B(B[0]), .Z(PRODUCT[13]) );
  AND U245 ( .A(A[12]), .B(B[0]), .Z(PRODUCT[12]) );
  AND U246 ( .A(A[11]), .B(B[0]), .Z(PRODUCT[11]) );
  AND U247 ( .A(A[10]), .B(B[0]), .Z(PRODUCT[10]) );
  AND U248 ( .A(B[0]), .B(A[9]), .Z(PRODUCT[9]) );
  AND U249 ( .A(A[8]), .B(B[0]), .Z(PRODUCT[8]) );
  AND U250 ( .A(A[7]), .B(B[0]), .Z(PRODUCT[7]) );
  AND U251 ( .A(A[6]), .B(B[0]), .Z(PRODUCT[6]) );
  AND U252 ( .A(A[5]), .B(B[0]), .Z(PRODUCT[5]) );
  AND U253 ( .A(A[4]), .B(B[0]), .Z(PRODUCT[4]) );
  AND U254 ( .A(A[3]), .B(B[0]), .Z(PRODUCT[3]) );
  AND U255 ( .A(A[2]), .B(B[0]), .Z(PRODUCT[2]) );
  AND U256 ( .A(A[1]), .B(B[0]), .Z(PRODUCT[1]) );
  AND U257 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
endmodule


module modmult_step_N256_4_DW01_cmp2_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [257:0] A;
  input [257:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;

  NAND U1 ( .A(n1), .B(n2), .Z(LT_LE) );
  NOR U2 ( .A(B[257]), .B(B[256]), .Z(n2) );
  AND U3 ( .A(n3), .B(n4), .Z(n1) );
  NAND U4 ( .A(n5), .B(n6), .Z(n4) );
  NANDN U5 ( .A(B[255]), .B(A[255]), .Z(n6) );
  NAND U6 ( .A(n7), .B(n8), .Z(n5) );
  NANDN U7 ( .A(A[254]), .B(B[254]), .Z(n8) );
  NAND U8 ( .A(n9), .B(n10), .Z(n7) );
  NANDN U9 ( .A(B[254]), .B(A[254]), .Z(n10) );
  AND U10 ( .A(n11), .B(n12), .Z(n9) );
  NAND U11 ( .A(n13), .B(n14), .Z(n12) );
  NANDN U12 ( .A(A[253]), .B(B[253]), .Z(n14) );
  AND U13 ( .A(n15), .B(n16), .Z(n13) );
  NANDN U14 ( .A(A[252]), .B(B[252]), .Z(n16) );
  NAND U15 ( .A(n17), .B(n18), .Z(n15) );
  NANDN U16 ( .A(B[252]), .B(A[252]), .Z(n18) );
  AND U17 ( .A(n19), .B(n20), .Z(n17) );
  NAND U18 ( .A(n21), .B(n22), .Z(n20) );
  NANDN U19 ( .A(A[251]), .B(B[251]), .Z(n22) );
  AND U20 ( .A(n23), .B(n24), .Z(n21) );
  NANDN U21 ( .A(A[250]), .B(B[250]), .Z(n24) );
  NAND U22 ( .A(n25), .B(n26), .Z(n23) );
  NANDN U23 ( .A(B[250]), .B(A[250]), .Z(n26) );
  AND U24 ( .A(n27), .B(n28), .Z(n25) );
  NAND U25 ( .A(n29), .B(n30), .Z(n28) );
  NANDN U26 ( .A(A[249]), .B(B[249]), .Z(n30) );
  AND U27 ( .A(n31), .B(n32), .Z(n29) );
  NANDN U28 ( .A(A[248]), .B(B[248]), .Z(n32) );
  NAND U29 ( .A(n33), .B(n34), .Z(n31) );
  NANDN U30 ( .A(B[248]), .B(A[248]), .Z(n34) );
  AND U31 ( .A(n35), .B(n36), .Z(n33) );
  NAND U32 ( .A(n37), .B(n38), .Z(n36) );
  NANDN U33 ( .A(A[247]), .B(B[247]), .Z(n38) );
  AND U34 ( .A(n39), .B(n40), .Z(n37) );
  NANDN U35 ( .A(A[246]), .B(B[246]), .Z(n40) );
  NAND U36 ( .A(n41), .B(n42), .Z(n39) );
  NANDN U37 ( .A(B[246]), .B(A[246]), .Z(n42) );
  AND U38 ( .A(n43), .B(n44), .Z(n41) );
  NAND U39 ( .A(n45), .B(n46), .Z(n44) );
  NANDN U40 ( .A(A[245]), .B(B[245]), .Z(n46) );
  AND U41 ( .A(n47), .B(n48), .Z(n45) );
  NANDN U42 ( .A(A[244]), .B(B[244]), .Z(n48) );
  NAND U43 ( .A(n49), .B(n50), .Z(n47) );
  NANDN U44 ( .A(B[244]), .B(A[244]), .Z(n50) );
  AND U45 ( .A(n51), .B(n52), .Z(n49) );
  NAND U46 ( .A(n53), .B(n54), .Z(n52) );
  NANDN U47 ( .A(A[243]), .B(B[243]), .Z(n54) );
  AND U48 ( .A(n55), .B(n56), .Z(n53) );
  NANDN U49 ( .A(A[242]), .B(B[242]), .Z(n56) );
  NAND U50 ( .A(n57), .B(n58), .Z(n55) );
  NANDN U51 ( .A(B[242]), .B(A[242]), .Z(n58) );
  AND U52 ( .A(n59), .B(n60), .Z(n57) );
  NAND U53 ( .A(n61), .B(n62), .Z(n60) );
  NANDN U54 ( .A(A[241]), .B(B[241]), .Z(n62) );
  AND U55 ( .A(n63), .B(n64), .Z(n61) );
  NANDN U56 ( .A(A[240]), .B(B[240]), .Z(n64) );
  NAND U57 ( .A(n65), .B(n66), .Z(n63) );
  NANDN U58 ( .A(B[240]), .B(A[240]), .Z(n66) );
  AND U59 ( .A(n67), .B(n68), .Z(n65) );
  NAND U60 ( .A(n69), .B(n70), .Z(n68) );
  NANDN U61 ( .A(A[239]), .B(B[239]), .Z(n70) );
  AND U62 ( .A(n71), .B(n72), .Z(n69) );
  NANDN U63 ( .A(A[238]), .B(B[238]), .Z(n72) );
  NAND U64 ( .A(n73), .B(n74), .Z(n71) );
  NANDN U65 ( .A(B[238]), .B(A[238]), .Z(n74) );
  AND U66 ( .A(n75), .B(n76), .Z(n73) );
  NAND U67 ( .A(n77), .B(n78), .Z(n76) );
  NANDN U68 ( .A(A[237]), .B(B[237]), .Z(n78) );
  AND U69 ( .A(n79), .B(n80), .Z(n77) );
  NANDN U70 ( .A(A[236]), .B(B[236]), .Z(n80) );
  NAND U71 ( .A(n81), .B(n82), .Z(n79) );
  NANDN U72 ( .A(B[236]), .B(A[236]), .Z(n82) );
  AND U73 ( .A(n83), .B(n84), .Z(n81) );
  NAND U74 ( .A(n85), .B(n86), .Z(n84) );
  NANDN U75 ( .A(A[235]), .B(B[235]), .Z(n86) );
  AND U76 ( .A(n87), .B(n88), .Z(n85) );
  NANDN U77 ( .A(A[234]), .B(B[234]), .Z(n88) );
  NAND U78 ( .A(n89), .B(n90), .Z(n87) );
  NANDN U79 ( .A(B[234]), .B(A[234]), .Z(n90) );
  AND U80 ( .A(n91), .B(n92), .Z(n89) );
  NAND U81 ( .A(n93), .B(n94), .Z(n92) );
  NANDN U82 ( .A(A[233]), .B(B[233]), .Z(n94) );
  AND U83 ( .A(n95), .B(n96), .Z(n93) );
  NANDN U84 ( .A(A[232]), .B(B[232]), .Z(n96) );
  NAND U85 ( .A(n97), .B(n98), .Z(n95) );
  NANDN U86 ( .A(B[232]), .B(A[232]), .Z(n98) );
  AND U87 ( .A(n99), .B(n100), .Z(n97) );
  NAND U88 ( .A(n101), .B(n102), .Z(n100) );
  NANDN U89 ( .A(A[231]), .B(B[231]), .Z(n102) );
  AND U90 ( .A(n103), .B(n104), .Z(n101) );
  NANDN U91 ( .A(A[230]), .B(B[230]), .Z(n104) );
  NAND U92 ( .A(n105), .B(n106), .Z(n103) );
  NANDN U93 ( .A(B[230]), .B(A[230]), .Z(n106) );
  AND U94 ( .A(n107), .B(n108), .Z(n105) );
  NAND U95 ( .A(n109), .B(n110), .Z(n108) );
  NANDN U96 ( .A(A[229]), .B(B[229]), .Z(n110) );
  AND U97 ( .A(n111), .B(n112), .Z(n109) );
  NANDN U98 ( .A(A[228]), .B(B[228]), .Z(n112) );
  NAND U99 ( .A(n113), .B(n114), .Z(n111) );
  NANDN U100 ( .A(B[228]), .B(A[228]), .Z(n114) );
  AND U101 ( .A(n115), .B(n116), .Z(n113) );
  NAND U102 ( .A(n117), .B(n118), .Z(n116) );
  NANDN U103 ( .A(A[227]), .B(B[227]), .Z(n118) );
  AND U104 ( .A(n119), .B(n120), .Z(n117) );
  NANDN U105 ( .A(A[226]), .B(B[226]), .Z(n120) );
  NAND U106 ( .A(n121), .B(n122), .Z(n119) );
  NANDN U107 ( .A(B[226]), .B(A[226]), .Z(n122) );
  AND U108 ( .A(n123), .B(n124), .Z(n121) );
  NAND U109 ( .A(n125), .B(n126), .Z(n124) );
  NANDN U110 ( .A(A[225]), .B(B[225]), .Z(n126) );
  AND U111 ( .A(n127), .B(n128), .Z(n125) );
  NANDN U112 ( .A(A[224]), .B(B[224]), .Z(n128) );
  NAND U113 ( .A(n129), .B(n130), .Z(n127) );
  NANDN U114 ( .A(B[224]), .B(A[224]), .Z(n130) );
  AND U115 ( .A(n131), .B(n132), .Z(n129) );
  NAND U116 ( .A(n133), .B(n134), .Z(n132) );
  NANDN U117 ( .A(A[223]), .B(B[223]), .Z(n134) );
  AND U118 ( .A(n135), .B(n136), .Z(n133) );
  NANDN U119 ( .A(A[222]), .B(B[222]), .Z(n136) );
  NAND U120 ( .A(n137), .B(n138), .Z(n135) );
  NANDN U121 ( .A(B[222]), .B(A[222]), .Z(n138) );
  AND U122 ( .A(n139), .B(n140), .Z(n137) );
  NAND U123 ( .A(n141), .B(n142), .Z(n140) );
  NANDN U124 ( .A(A[221]), .B(B[221]), .Z(n142) );
  AND U125 ( .A(n143), .B(n144), .Z(n141) );
  NANDN U126 ( .A(A[220]), .B(B[220]), .Z(n144) );
  NAND U127 ( .A(n145), .B(n146), .Z(n143) );
  NANDN U128 ( .A(B[220]), .B(A[220]), .Z(n146) );
  AND U129 ( .A(n147), .B(n148), .Z(n145) );
  NAND U130 ( .A(n149), .B(n150), .Z(n148) );
  NANDN U131 ( .A(A[219]), .B(B[219]), .Z(n150) );
  AND U132 ( .A(n151), .B(n152), .Z(n149) );
  NANDN U133 ( .A(A[218]), .B(B[218]), .Z(n152) );
  NAND U134 ( .A(n153), .B(n154), .Z(n151) );
  NANDN U135 ( .A(B[218]), .B(A[218]), .Z(n154) );
  AND U136 ( .A(n155), .B(n156), .Z(n153) );
  NAND U137 ( .A(n157), .B(n158), .Z(n156) );
  NANDN U138 ( .A(A[217]), .B(B[217]), .Z(n158) );
  AND U139 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U140 ( .A(A[216]), .B(B[216]), .Z(n160) );
  NAND U141 ( .A(n161), .B(n162), .Z(n159) );
  NANDN U142 ( .A(B[216]), .B(A[216]), .Z(n162) );
  AND U143 ( .A(n163), .B(n164), .Z(n161) );
  NAND U144 ( .A(n165), .B(n166), .Z(n164) );
  NANDN U145 ( .A(A[215]), .B(B[215]), .Z(n166) );
  AND U146 ( .A(n167), .B(n168), .Z(n165) );
  NANDN U147 ( .A(A[214]), .B(B[214]), .Z(n168) );
  NAND U148 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U149 ( .A(B[214]), .B(A[214]), .Z(n170) );
  AND U150 ( .A(n171), .B(n172), .Z(n169) );
  NAND U151 ( .A(n173), .B(n174), .Z(n172) );
  NANDN U152 ( .A(A[213]), .B(B[213]), .Z(n174) );
  AND U153 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U154 ( .A(A[212]), .B(B[212]), .Z(n176) );
  NAND U155 ( .A(n177), .B(n178), .Z(n175) );
  NANDN U156 ( .A(B[212]), .B(A[212]), .Z(n178) );
  AND U157 ( .A(n179), .B(n180), .Z(n177) );
  NAND U158 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U159 ( .A(A[211]), .B(B[211]), .Z(n182) );
  AND U160 ( .A(n183), .B(n184), .Z(n181) );
  NANDN U161 ( .A(A[210]), .B(B[210]), .Z(n184) );
  NAND U162 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U163 ( .A(B[210]), .B(A[210]), .Z(n186) );
  AND U164 ( .A(n187), .B(n188), .Z(n185) );
  NAND U165 ( .A(n189), .B(n190), .Z(n188) );
  NANDN U166 ( .A(A[209]), .B(B[209]), .Z(n190) );
  AND U167 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U168 ( .A(A[208]), .B(B[208]), .Z(n192) );
  NAND U169 ( .A(n193), .B(n194), .Z(n191) );
  NANDN U170 ( .A(B[208]), .B(A[208]), .Z(n194) );
  AND U171 ( .A(n195), .B(n196), .Z(n193) );
  NAND U172 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U173 ( .A(A[207]), .B(B[207]), .Z(n198) );
  AND U174 ( .A(n199), .B(n200), .Z(n197) );
  NANDN U175 ( .A(A[206]), .B(B[206]), .Z(n200) );
  NAND U176 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U177 ( .A(B[206]), .B(A[206]), .Z(n202) );
  AND U178 ( .A(n203), .B(n204), .Z(n201) );
  NAND U179 ( .A(n205), .B(n206), .Z(n204) );
  NANDN U180 ( .A(A[205]), .B(B[205]), .Z(n206) );
  AND U181 ( .A(n207), .B(n208), .Z(n205) );
  NANDN U182 ( .A(A[204]), .B(B[204]), .Z(n208) );
  NAND U183 ( .A(n209), .B(n210), .Z(n207) );
  NANDN U184 ( .A(B[204]), .B(A[204]), .Z(n210) );
  AND U185 ( .A(n211), .B(n212), .Z(n209) );
  NAND U186 ( .A(n213), .B(n214), .Z(n212) );
  NANDN U187 ( .A(A[203]), .B(B[203]), .Z(n214) );
  AND U188 ( .A(n215), .B(n216), .Z(n213) );
  NANDN U189 ( .A(A[202]), .B(B[202]), .Z(n216) );
  NAND U190 ( .A(n217), .B(n218), .Z(n215) );
  NANDN U191 ( .A(B[202]), .B(A[202]), .Z(n218) );
  AND U192 ( .A(n219), .B(n220), .Z(n217) );
  NAND U193 ( .A(n221), .B(n222), .Z(n220) );
  NANDN U194 ( .A(A[201]), .B(B[201]), .Z(n222) );
  AND U195 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U196 ( .A(A[200]), .B(B[200]), .Z(n224) );
  NAND U197 ( .A(n225), .B(n226), .Z(n223) );
  NANDN U198 ( .A(B[200]), .B(A[200]), .Z(n226) );
  AND U199 ( .A(n227), .B(n228), .Z(n225) );
  NAND U200 ( .A(n229), .B(n230), .Z(n228) );
  NANDN U201 ( .A(A[199]), .B(B[199]), .Z(n230) );
  AND U202 ( .A(n231), .B(n232), .Z(n229) );
  NANDN U203 ( .A(A[198]), .B(B[198]), .Z(n232) );
  NAND U204 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U205 ( .A(B[198]), .B(A[198]), .Z(n234) );
  AND U206 ( .A(n235), .B(n236), .Z(n233) );
  NAND U207 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U208 ( .A(A[197]), .B(B[197]), .Z(n238) );
  AND U209 ( .A(n239), .B(n240), .Z(n237) );
  NANDN U210 ( .A(A[196]), .B(B[196]), .Z(n240) );
  NAND U211 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U212 ( .A(B[196]), .B(A[196]), .Z(n242) );
  AND U213 ( .A(n243), .B(n244), .Z(n241) );
  NAND U214 ( .A(n245), .B(n246), .Z(n244) );
  NANDN U215 ( .A(A[195]), .B(B[195]), .Z(n246) );
  AND U216 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U217 ( .A(A[194]), .B(B[194]), .Z(n248) );
  NAND U218 ( .A(n249), .B(n250), .Z(n247) );
  NANDN U219 ( .A(B[194]), .B(A[194]), .Z(n250) );
  AND U220 ( .A(n251), .B(n252), .Z(n249) );
  NAND U221 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U222 ( .A(A[193]), .B(B[193]), .Z(n254) );
  AND U223 ( .A(n255), .B(n256), .Z(n253) );
  NANDN U224 ( .A(A[192]), .B(B[192]), .Z(n256) );
  NAND U225 ( .A(n257), .B(n258), .Z(n255) );
  NANDN U226 ( .A(B[192]), .B(A[192]), .Z(n258) );
  AND U227 ( .A(n259), .B(n260), .Z(n257) );
  NAND U228 ( .A(n261), .B(n262), .Z(n260) );
  NANDN U229 ( .A(A[191]), .B(B[191]), .Z(n262) );
  AND U230 ( .A(n263), .B(n264), .Z(n261) );
  NANDN U231 ( .A(A[190]), .B(B[190]), .Z(n264) );
  NAND U232 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U233 ( .A(B[190]), .B(A[190]), .Z(n266) );
  AND U234 ( .A(n267), .B(n268), .Z(n265) );
  NAND U235 ( .A(n269), .B(n270), .Z(n268) );
  NANDN U236 ( .A(A[189]), .B(B[189]), .Z(n270) );
  AND U237 ( .A(n271), .B(n272), .Z(n269) );
  NANDN U238 ( .A(A[188]), .B(B[188]), .Z(n272) );
  NAND U239 ( .A(n273), .B(n274), .Z(n271) );
  NANDN U240 ( .A(B[188]), .B(A[188]), .Z(n274) );
  AND U241 ( .A(n275), .B(n276), .Z(n273) );
  NAND U242 ( .A(n277), .B(n278), .Z(n276) );
  NANDN U243 ( .A(A[187]), .B(B[187]), .Z(n278) );
  AND U244 ( .A(n279), .B(n280), .Z(n277) );
  NANDN U245 ( .A(A[186]), .B(B[186]), .Z(n280) );
  NAND U246 ( .A(n281), .B(n282), .Z(n279) );
  NANDN U247 ( .A(B[186]), .B(A[186]), .Z(n282) );
  AND U248 ( .A(n283), .B(n284), .Z(n281) );
  NAND U249 ( .A(n285), .B(n286), .Z(n284) );
  NANDN U250 ( .A(A[185]), .B(B[185]), .Z(n286) );
  AND U251 ( .A(n287), .B(n288), .Z(n285) );
  NANDN U252 ( .A(A[184]), .B(B[184]), .Z(n288) );
  NAND U253 ( .A(n289), .B(n290), .Z(n287) );
  NANDN U254 ( .A(B[184]), .B(A[184]), .Z(n290) );
  AND U255 ( .A(n291), .B(n292), .Z(n289) );
  NAND U256 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U257 ( .A(A[183]), .B(B[183]), .Z(n294) );
  AND U258 ( .A(n295), .B(n296), .Z(n293) );
  NANDN U259 ( .A(A[182]), .B(B[182]), .Z(n296) );
  NAND U260 ( .A(n297), .B(n298), .Z(n295) );
  NANDN U261 ( .A(B[182]), .B(A[182]), .Z(n298) );
  AND U262 ( .A(n299), .B(n300), .Z(n297) );
  NAND U263 ( .A(n301), .B(n302), .Z(n300) );
  NANDN U264 ( .A(A[181]), .B(B[181]), .Z(n302) );
  AND U265 ( .A(n303), .B(n304), .Z(n301) );
  NANDN U266 ( .A(A[180]), .B(B[180]), .Z(n304) );
  NAND U267 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U268 ( .A(B[180]), .B(A[180]), .Z(n306) );
  AND U269 ( .A(n307), .B(n308), .Z(n305) );
  NAND U270 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U271 ( .A(A[179]), .B(B[179]), .Z(n310) );
  AND U272 ( .A(n311), .B(n312), .Z(n309) );
  NANDN U273 ( .A(A[178]), .B(B[178]), .Z(n312) );
  NAND U274 ( .A(n313), .B(n314), .Z(n311) );
  NANDN U275 ( .A(B[178]), .B(A[178]), .Z(n314) );
  AND U276 ( .A(n315), .B(n316), .Z(n313) );
  NAND U277 ( .A(n317), .B(n318), .Z(n316) );
  NANDN U278 ( .A(A[177]), .B(B[177]), .Z(n318) );
  AND U279 ( .A(n319), .B(n320), .Z(n317) );
  NANDN U280 ( .A(A[176]), .B(B[176]), .Z(n320) );
  NAND U281 ( .A(n321), .B(n322), .Z(n319) );
  NANDN U282 ( .A(B[176]), .B(A[176]), .Z(n322) );
  AND U283 ( .A(n323), .B(n324), .Z(n321) );
  NAND U284 ( .A(n325), .B(n326), .Z(n324) );
  NANDN U285 ( .A(A[175]), .B(B[175]), .Z(n326) );
  AND U286 ( .A(n327), .B(n328), .Z(n325) );
  NANDN U287 ( .A(A[174]), .B(B[174]), .Z(n328) );
  NAND U288 ( .A(n329), .B(n330), .Z(n327) );
  NANDN U289 ( .A(B[174]), .B(A[174]), .Z(n330) );
  AND U290 ( .A(n331), .B(n332), .Z(n329) );
  NAND U291 ( .A(n333), .B(n334), .Z(n332) );
  NANDN U292 ( .A(A[173]), .B(B[173]), .Z(n334) );
  AND U293 ( .A(n335), .B(n336), .Z(n333) );
  NANDN U294 ( .A(A[172]), .B(B[172]), .Z(n336) );
  NAND U295 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U296 ( .A(B[172]), .B(A[172]), .Z(n338) );
  AND U297 ( .A(n339), .B(n340), .Z(n337) );
  NAND U298 ( .A(n341), .B(n342), .Z(n340) );
  NANDN U299 ( .A(A[171]), .B(B[171]), .Z(n342) );
  AND U300 ( .A(n343), .B(n344), .Z(n341) );
  NANDN U301 ( .A(A[170]), .B(B[170]), .Z(n344) );
  NAND U302 ( .A(n345), .B(n346), .Z(n343) );
  NANDN U303 ( .A(B[170]), .B(A[170]), .Z(n346) );
  AND U304 ( .A(n347), .B(n348), .Z(n345) );
  NAND U305 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U306 ( .A(A[169]), .B(B[169]), .Z(n350) );
  AND U307 ( .A(n351), .B(n352), .Z(n349) );
  NANDN U308 ( .A(A[168]), .B(B[168]), .Z(n352) );
  NAND U309 ( .A(n353), .B(n354), .Z(n351) );
  NANDN U310 ( .A(B[168]), .B(A[168]), .Z(n354) );
  AND U311 ( .A(n355), .B(n356), .Z(n353) );
  NAND U312 ( .A(n357), .B(n358), .Z(n356) );
  NANDN U313 ( .A(A[167]), .B(B[167]), .Z(n358) );
  AND U314 ( .A(n359), .B(n360), .Z(n357) );
  NANDN U315 ( .A(A[166]), .B(B[166]), .Z(n360) );
  NAND U316 ( .A(n361), .B(n362), .Z(n359) );
  NANDN U317 ( .A(B[166]), .B(A[166]), .Z(n362) );
  AND U318 ( .A(n363), .B(n364), .Z(n361) );
  NAND U319 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U320 ( .A(A[165]), .B(B[165]), .Z(n366) );
  AND U321 ( .A(n367), .B(n368), .Z(n365) );
  NANDN U322 ( .A(A[164]), .B(B[164]), .Z(n368) );
  NAND U323 ( .A(n369), .B(n370), .Z(n367) );
  NANDN U324 ( .A(B[164]), .B(A[164]), .Z(n370) );
  AND U325 ( .A(n371), .B(n372), .Z(n369) );
  NAND U326 ( .A(n373), .B(n374), .Z(n372) );
  NANDN U327 ( .A(A[163]), .B(B[163]), .Z(n374) );
  AND U328 ( .A(n375), .B(n376), .Z(n373) );
  NANDN U329 ( .A(A[162]), .B(B[162]), .Z(n376) );
  NAND U330 ( .A(n377), .B(n378), .Z(n375) );
  NANDN U331 ( .A(B[162]), .B(A[162]), .Z(n378) );
  AND U332 ( .A(n379), .B(n380), .Z(n377) );
  NAND U333 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U334 ( .A(A[161]), .B(B[161]), .Z(n382) );
  AND U335 ( .A(n383), .B(n384), .Z(n381) );
  NANDN U336 ( .A(A[160]), .B(B[160]), .Z(n384) );
  NAND U337 ( .A(n385), .B(n386), .Z(n383) );
  NANDN U338 ( .A(B[160]), .B(A[160]), .Z(n386) );
  AND U339 ( .A(n387), .B(n388), .Z(n385) );
  NAND U340 ( .A(n389), .B(n390), .Z(n388) );
  NANDN U341 ( .A(A[159]), .B(B[159]), .Z(n390) );
  AND U342 ( .A(n391), .B(n392), .Z(n389) );
  NANDN U343 ( .A(A[158]), .B(B[158]), .Z(n392) );
  NAND U344 ( .A(n393), .B(n394), .Z(n391) );
  NANDN U345 ( .A(B[158]), .B(A[158]), .Z(n394) );
  AND U346 ( .A(n395), .B(n396), .Z(n393) );
  NAND U347 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U348 ( .A(A[157]), .B(B[157]), .Z(n398) );
  AND U349 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U350 ( .A(A[156]), .B(B[156]), .Z(n400) );
  NAND U351 ( .A(n401), .B(n402), .Z(n399) );
  NANDN U352 ( .A(B[156]), .B(A[156]), .Z(n402) );
  AND U353 ( .A(n403), .B(n404), .Z(n401) );
  NAND U354 ( .A(n405), .B(n406), .Z(n404) );
  NANDN U355 ( .A(A[155]), .B(B[155]), .Z(n406) );
  AND U356 ( .A(n407), .B(n408), .Z(n405) );
  NANDN U357 ( .A(A[154]), .B(B[154]), .Z(n408) );
  NAND U358 ( .A(n409), .B(n410), .Z(n407) );
  NANDN U359 ( .A(B[154]), .B(A[154]), .Z(n410) );
  AND U360 ( .A(n411), .B(n412), .Z(n409) );
  NAND U361 ( .A(n413), .B(n414), .Z(n412) );
  NANDN U362 ( .A(A[153]), .B(B[153]), .Z(n414) );
  AND U363 ( .A(n415), .B(n416), .Z(n413) );
  NANDN U364 ( .A(A[152]), .B(B[152]), .Z(n416) );
  NAND U365 ( .A(n417), .B(n418), .Z(n415) );
  NANDN U366 ( .A(B[152]), .B(A[152]), .Z(n418) );
  AND U367 ( .A(n419), .B(n420), .Z(n417) );
  NAND U368 ( .A(n421), .B(n422), .Z(n420) );
  NANDN U369 ( .A(A[151]), .B(B[151]), .Z(n422) );
  AND U370 ( .A(n423), .B(n424), .Z(n421) );
  NANDN U371 ( .A(A[150]), .B(B[150]), .Z(n424) );
  NAND U372 ( .A(n425), .B(n426), .Z(n423) );
  NANDN U373 ( .A(B[150]), .B(A[150]), .Z(n426) );
  AND U374 ( .A(n427), .B(n428), .Z(n425) );
  NAND U375 ( .A(n429), .B(n430), .Z(n428) );
  NANDN U376 ( .A(A[149]), .B(B[149]), .Z(n430) );
  AND U377 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U378 ( .A(A[148]), .B(B[148]), .Z(n432) );
  NAND U379 ( .A(n433), .B(n434), .Z(n431) );
  NANDN U380 ( .A(B[148]), .B(A[148]), .Z(n434) );
  AND U381 ( .A(n435), .B(n436), .Z(n433) );
  NAND U382 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U383 ( .A(A[147]), .B(B[147]), .Z(n438) );
  AND U384 ( .A(n439), .B(n440), .Z(n437) );
  NANDN U385 ( .A(A[146]), .B(B[146]), .Z(n440) );
  NAND U386 ( .A(n441), .B(n442), .Z(n439) );
  NANDN U387 ( .A(B[146]), .B(A[146]), .Z(n442) );
  AND U388 ( .A(n443), .B(n444), .Z(n441) );
  NAND U389 ( .A(n445), .B(n446), .Z(n444) );
  NANDN U390 ( .A(A[145]), .B(B[145]), .Z(n446) );
  AND U391 ( .A(n447), .B(n448), .Z(n445) );
  NANDN U392 ( .A(A[144]), .B(B[144]), .Z(n448) );
  NAND U393 ( .A(n449), .B(n450), .Z(n447) );
  NANDN U394 ( .A(B[144]), .B(A[144]), .Z(n450) );
  AND U395 ( .A(n451), .B(n452), .Z(n449) );
  NAND U396 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U397 ( .A(A[143]), .B(B[143]), .Z(n454) );
  AND U398 ( .A(n455), .B(n456), .Z(n453) );
  NANDN U399 ( .A(A[142]), .B(B[142]), .Z(n456) );
  NAND U400 ( .A(n457), .B(n458), .Z(n455) );
  NANDN U401 ( .A(B[142]), .B(A[142]), .Z(n458) );
  AND U402 ( .A(n459), .B(n460), .Z(n457) );
  NAND U403 ( .A(n461), .B(n462), .Z(n460) );
  NANDN U404 ( .A(A[141]), .B(B[141]), .Z(n462) );
  AND U405 ( .A(n463), .B(n464), .Z(n461) );
  NANDN U406 ( .A(A[140]), .B(B[140]), .Z(n464) );
  NAND U407 ( .A(n465), .B(n466), .Z(n463) );
  NANDN U408 ( .A(B[140]), .B(A[140]), .Z(n466) );
  AND U409 ( .A(n467), .B(n468), .Z(n465) );
  NAND U410 ( .A(n469), .B(n470), .Z(n468) );
  NANDN U411 ( .A(A[139]), .B(B[139]), .Z(n470) );
  AND U412 ( .A(n471), .B(n472), .Z(n469) );
  NANDN U413 ( .A(A[138]), .B(B[138]), .Z(n472) );
  NAND U414 ( .A(n473), .B(n474), .Z(n471) );
  NANDN U415 ( .A(B[138]), .B(A[138]), .Z(n474) );
  AND U416 ( .A(n475), .B(n476), .Z(n473) );
  NAND U417 ( .A(n477), .B(n478), .Z(n476) );
  NANDN U418 ( .A(A[137]), .B(B[137]), .Z(n478) );
  AND U419 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U420 ( .A(A[136]), .B(B[136]), .Z(n480) );
  NAND U421 ( .A(n481), .B(n482), .Z(n479) );
  NANDN U422 ( .A(B[136]), .B(A[136]), .Z(n482) );
  AND U423 ( .A(n483), .B(n484), .Z(n481) );
  NAND U424 ( .A(n485), .B(n486), .Z(n484) );
  NANDN U425 ( .A(A[135]), .B(B[135]), .Z(n486) );
  AND U426 ( .A(n487), .B(n488), .Z(n485) );
  NANDN U427 ( .A(A[134]), .B(B[134]), .Z(n488) );
  NAND U428 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U429 ( .A(B[134]), .B(A[134]), .Z(n490) );
  AND U430 ( .A(n491), .B(n492), .Z(n489) );
  NAND U431 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U432 ( .A(A[133]), .B(B[133]), .Z(n494) );
  AND U433 ( .A(n495), .B(n496), .Z(n493) );
  NANDN U434 ( .A(A[132]), .B(B[132]), .Z(n496) );
  NAND U435 ( .A(n497), .B(n498), .Z(n495) );
  NANDN U436 ( .A(B[132]), .B(A[132]), .Z(n498) );
  AND U437 ( .A(n499), .B(n500), .Z(n497) );
  NAND U438 ( .A(n501), .B(n502), .Z(n500) );
  NANDN U439 ( .A(A[131]), .B(B[131]), .Z(n502) );
  AND U440 ( .A(n503), .B(n504), .Z(n501) );
  NANDN U441 ( .A(A[130]), .B(B[130]), .Z(n504) );
  NAND U442 ( .A(n505), .B(n506), .Z(n503) );
  NANDN U443 ( .A(B[130]), .B(A[130]), .Z(n506) );
  AND U444 ( .A(n507), .B(n508), .Z(n505) );
  NAND U445 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U446 ( .A(A[129]), .B(B[129]), .Z(n510) );
  AND U447 ( .A(n511), .B(n512), .Z(n509) );
  NANDN U448 ( .A(A[128]), .B(B[128]), .Z(n512) );
  NAND U449 ( .A(n513), .B(n514), .Z(n511) );
  NANDN U450 ( .A(B[128]), .B(A[128]), .Z(n514) );
  AND U451 ( .A(n515), .B(n516), .Z(n513) );
  NAND U452 ( .A(n517), .B(n518), .Z(n516) );
  NANDN U453 ( .A(A[127]), .B(B[127]), .Z(n518) );
  AND U454 ( .A(n519), .B(n520), .Z(n517) );
  NANDN U455 ( .A(A[126]), .B(B[126]), .Z(n520) );
  NAND U456 ( .A(n521), .B(n522), .Z(n519) );
  NANDN U457 ( .A(B[126]), .B(A[126]), .Z(n522) );
  AND U458 ( .A(n523), .B(n524), .Z(n521) );
  NAND U459 ( .A(n525), .B(n526), .Z(n524) );
  NANDN U460 ( .A(A[125]), .B(B[125]), .Z(n526) );
  AND U461 ( .A(n527), .B(n528), .Z(n525) );
  NANDN U462 ( .A(A[124]), .B(B[124]), .Z(n528) );
  NAND U463 ( .A(n529), .B(n530), .Z(n527) );
  NANDN U464 ( .A(B[124]), .B(A[124]), .Z(n530) );
  AND U465 ( .A(n531), .B(n532), .Z(n529) );
  NAND U466 ( .A(n533), .B(n534), .Z(n532) );
  NANDN U467 ( .A(A[123]), .B(B[123]), .Z(n534) );
  AND U468 ( .A(n535), .B(n536), .Z(n533) );
  NANDN U469 ( .A(A[122]), .B(B[122]), .Z(n536) );
  NAND U470 ( .A(n537), .B(n538), .Z(n535) );
  NANDN U471 ( .A(B[122]), .B(A[122]), .Z(n538) );
  AND U472 ( .A(n539), .B(n540), .Z(n537) );
  NAND U473 ( .A(n541), .B(n542), .Z(n540) );
  NANDN U474 ( .A(A[121]), .B(B[121]), .Z(n542) );
  AND U475 ( .A(n543), .B(n544), .Z(n541) );
  NANDN U476 ( .A(A[120]), .B(B[120]), .Z(n544) );
  NAND U477 ( .A(n545), .B(n546), .Z(n543) );
  NANDN U478 ( .A(B[120]), .B(A[120]), .Z(n546) );
  AND U479 ( .A(n547), .B(n548), .Z(n545) );
  NAND U480 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U481 ( .A(A[119]), .B(B[119]), .Z(n550) );
  AND U482 ( .A(n551), .B(n552), .Z(n549) );
  NANDN U483 ( .A(A[118]), .B(B[118]), .Z(n552) );
  NAND U484 ( .A(n553), .B(n554), .Z(n551) );
  NANDN U485 ( .A(B[118]), .B(A[118]), .Z(n554) );
  AND U486 ( .A(n555), .B(n556), .Z(n553) );
  NAND U487 ( .A(n557), .B(n558), .Z(n556) );
  NANDN U488 ( .A(A[117]), .B(B[117]), .Z(n558) );
  AND U489 ( .A(n559), .B(n560), .Z(n557) );
  NANDN U490 ( .A(A[116]), .B(B[116]), .Z(n560) );
  NAND U491 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U492 ( .A(B[116]), .B(A[116]), .Z(n562) );
  AND U493 ( .A(n563), .B(n564), .Z(n561) );
  NAND U494 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U495 ( .A(A[115]), .B(B[115]), .Z(n566) );
  AND U496 ( .A(n567), .B(n568), .Z(n565) );
  NANDN U497 ( .A(A[114]), .B(B[114]), .Z(n568) );
  NAND U498 ( .A(n569), .B(n570), .Z(n567) );
  NANDN U499 ( .A(B[114]), .B(A[114]), .Z(n570) );
  AND U500 ( .A(n571), .B(n572), .Z(n569) );
  NAND U501 ( .A(n573), .B(n574), .Z(n572) );
  NANDN U502 ( .A(A[113]), .B(B[113]), .Z(n574) );
  AND U503 ( .A(n575), .B(n576), .Z(n573) );
  NANDN U504 ( .A(A[112]), .B(B[112]), .Z(n576) );
  NAND U505 ( .A(n577), .B(n578), .Z(n575) );
  NANDN U506 ( .A(B[112]), .B(A[112]), .Z(n578) );
  AND U507 ( .A(n579), .B(n580), .Z(n577) );
  NAND U508 ( .A(n581), .B(n582), .Z(n580) );
  NANDN U509 ( .A(A[111]), .B(B[111]), .Z(n582) );
  AND U510 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U511 ( .A(A[110]), .B(B[110]), .Z(n584) );
  NAND U512 ( .A(n585), .B(n586), .Z(n583) );
  NANDN U513 ( .A(B[110]), .B(A[110]), .Z(n586) );
  AND U514 ( .A(n587), .B(n588), .Z(n585) );
  NAND U515 ( .A(n589), .B(n590), .Z(n588) );
  NANDN U516 ( .A(A[109]), .B(B[109]), .Z(n590) );
  AND U517 ( .A(n591), .B(n592), .Z(n589) );
  NANDN U518 ( .A(A[108]), .B(B[108]), .Z(n592) );
  NAND U519 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U520 ( .A(B[108]), .B(A[108]), .Z(n594) );
  AND U521 ( .A(n595), .B(n596), .Z(n593) );
  NAND U522 ( .A(n597), .B(n598), .Z(n596) );
  NANDN U523 ( .A(A[107]), .B(B[107]), .Z(n598) );
  AND U524 ( .A(n599), .B(n600), .Z(n597) );
  NANDN U525 ( .A(A[106]), .B(B[106]), .Z(n600) );
  NAND U526 ( .A(n601), .B(n602), .Z(n599) );
  NANDN U527 ( .A(B[106]), .B(A[106]), .Z(n602) );
  AND U528 ( .A(n603), .B(n604), .Z(n601) );
  NAND U529 ( .A(n605), .B(n606), .Z(n604) );
  NANDN U530 ( .A(A[105]), .B(B[105]), .Z(n606) );
  AND U531 ( .A(n607), .B(n608), .Z(n605) );
  NANDN U532 ( .A(A[104]), .B(B[104]), .Z(n608) );
  NAND U533 ( .A(n609), .B(n610), .Z(n607) );
  NANDN U534 ( .A(B[104]), .B(A[104]), .Z(n610) );
  AND U535 ( .A(n611), .B(n612), .Z(n609) );
  NAND U536 ( .A(n613), .B(n614), .Z(n612) );
  NANDN U537 ( .A(A[103]), .B(B[103]), .Z(n614) );
  AND U538 ( .A(n615), .B(n616), .Z(n613) );
  NANDN U539 ( .A(A[102]), .B(B[102]), .Z(n616) );
  NAND U540 ( .A(n617), .B(n618), .Z(n615) );
  NANDN U541 ( .A(B[102]), .B(A[102]), .Z(n618) );
  AND U542 ( .A(n619), .B(n620), .Z(n617) );
  NAND U543 ( .A(n621), .B(n622), .Z(n620) );
  NANDN U544 ( .A(A[101]), .B(B[101]), .Z(n622) );
  AND U545 ( .A(n623), .B(n624), .Z(n621) );
  NANDN U546 ( .A(A[100]), .B(B[100]), .Z(n624) );
  NAND U547 ( .A(n625), .B(n626), .Z(n623) );
  NANDN U548 ( .A(B[99]), .B(A[99]), .Z(n626) );
  AND U549 ( .A(n627), .B(n628), .Z(n625) );
  NAND U550 ( .A(n629), .B(n630), .Z(n628) );
  NANDN U551 ( .A(A[99]), .B(B[99]), .Z(n630) );
  AND U552 ( .A(n631), .B(n632), .Z(n629) );
  NANDN U553 ( .A(A[98]), .B(B[98]), .Z(n632) );
  NAND U554 ( .A(n633), .B(n634), .Z(n631) );
  NANDN U555 ( .A(B[98]), .B(A[98]), .Z(n634) );
  AND U556 ( .A(n635), .B(n636), .Z(n633) );
  NAND U557 ( .A(n637), .B(n638), .Z(n636) );
  NANDN U558 ( .A(A[97]), .B(B[97]), .Z(n638) );
  AND U559 ( .A(n639), .B(n640), .Z(n637) );
  NANDN U560 ( .A(A[96]), .B(B[96]), .Z(n640) );
  NAND U561 ( .A(n641), .B(n642), .Z(n639) );
  NANDN U562 ( .A(B[96]), .B(A[96]), .Z(n642) );
  AND U563 ( .A(n643), .B(n644), .Z(n641) );
  NAND U564 ( .A(n645), .B(n646), .Z(n644) );
  NANDN U565 ( .A(A[95]), .B(B[95]), .Z(n646) );
  AND U566 ( .A(n647), .B(n648), .Z(n645) );
  NANDN U567 ( .A(A[94]), .B(B[94]), .Z(n648) );
  NAND U568 ( .A(n649), .B(n650), .Z(n647) );
  NANDN U569 ( .A(B[94]), .B(A[94]), .Z(n650) );
  AND U570 ( .A(n651), .B(n652), .Z(n649) );
  NAND U571 ( .A(n653), .B(n654), .Z(n652) );
  NANDN U572 ( .A(A[93]), .B(B[93]), .Z(n654) );
  AND U573 ( .A(n655), .B(n656), .Z(n653) );
  NANDN U574 ( .A(A[92]), .B(B[92]), .Z(n656) );
  NAND U575 ( .A(n657), .B(n658), .Z(n655) );
  NANDN U576 ( .A(B[92]), .B(A[92]), .Z(n658) );
  AND U577 ( .A(n659), .B(n660), .Z(n657) );
  NAND U578 ( .A(n661), .B(n662), .Z(n660) );
  NANDN U579 ( .A(A[91]), .B(B[91]), .Z(n662) );
  AND U580 ( .A(n663), .B(n664), .Z(n661) );
  NANDN U581 ( .A(A[90]), .B(B[90]), .Z(n664) );
  NAND U582 ( .A(n665), .B(n666), .Z(n663) );
  NANDN U583 ( .A(B[90]), .B(A[90]), .Z(n666) );
  AND U584 ( .A(n667), .B(n668), .Z(n665) );
  NAND U585 ( .A(n669), .B(n670), .Z(n668) );
  NANDN U586 ( .A(A[89]), .B(B[89]), .Z(n670) );
  AND U587 ( .A(n671), .B(n672), .Z(n669) );
  NANDN U588 ( .A(A[88]), .B(B[88]), .Z(n672) );
  NAND U589 ( .A(n673), .B(n674), .Z(n671) );
  NANDN U590 ( .A(B[88]), .B(A[88]), .Z(n674) );
  AND U591 ( .A(n675), .B(n676), .Z(n673) );
  NAND U592 ( .A(n677), .B(n678), .Z(n676) );
  NANDN U593 ( .A(A[87]), .B(B[87]), .Z(n678) );
  AND U594 ( .A(n679), .B(n680), .Z(n677) );
  NANDN U595 ( .A(A[86]), .B(B[86]), .Z(n680) );
  NAND U596 ( .A(n681), .B(n682), .Z(n679) );
  NANDN U597 ( .A(B[86]), .B(A[86]), .Z(n682) );
  AND U598 ( .A(n683), .B(n684), .Z(n681) );
  NAND U599 ( .A(n685), .B(n686), .Z(n684) );
  NANDN U600 ( .A(A[85]), .B(B[85]), .Z(n686) );
  AND U601 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U602 ( .A(A[84]), .B(B[84]), .Z(n688) );
  NAND U603 ( .A(n689), .B(n690), .Z(n687) );
  NANDN U604 ( .A(B[84]), .B(A[84]), .Z(n690) );
  AND U605 ( .A(n691), .B(n692), .Z(n689) );
  NAND U606 ( .A(n693), .B(n694), .Z(n692) );
  NANDN U607 ( .A(A[83]), .B(B[83]), .Z(n694) );
  AND U608 ( .A(n695), .B(n696), .Z(n693) );
  NANDN U609 ( .A(A[82]), .B(B[82]), .Z(n696) );
  NAND U610 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U611 ( .A(B[82]), .B(A[82]), .Z(n698) );
  AND U612 ( .A(n699), .B(n700), .Z(n697) );
  NAND U613 ( .A(n701), .B(n702), .Z(n700) );
  NANDN U614 ( .A(A[81]), .B(B[81]), .Z(n702) );
  AND U615 ( .A(n703), .B(n704), .Z(n701) );
  NANDN U616 ( .A(A[80]), .B(B[80]), .Z(n704) );
  NAND U617 ( .A(n705), .B(n706), .Z(n703) );
  NANDN U618 ( .A(B[80]), .B(A[80]), .Z(n706) );
  AND U619 ( .A(n707), .B(n708), .Z(n705) );
  NAND U620 ( .A(n709), .B(n710), .Z(n708) );
  NANDN U621 ( .A(A[79]), .B(B[79]), .Z(n710) );
  AND U622 ( .A(n711), .B(n712), .Z(n709) );
  NANDN U623 ( .A(A[78]), .B(B[78]), .Z(n712) );
  NAND U624 ( .A(n713), .B(n714), .Z(n711) );
  NANDN U625 ( .A(B[78]), .B(A[78]), .Z(n714) );
  AND U626 ( .A(n715), .B(n716), .Z(n713) );
  NAND U627 ( .A(n717), .B(n718), .Z(n716) );
  NANDN U628 ( .A(A[77]), .B(B[77]), .Z(n718) );
  AND U629 ( .A(n719), .B(n720), .Z(n717) );
  NANDN U630 ( .A(A[76]), .B(B[76]), .Z(n720) );
  NAND U631 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U632 ( .A(B[76]), .B(A[76]), .Z(n722) );
  AND U633 ( .A(n723), .B(n724), .Z(n721) );
  NAND U634 ( .A(n725), .B(n726), .Z(n724) );
  NANDN U635 ( .A(A[75]), .B(B[75]), .Z(n726) );
  AND U636 ( .A(n727), .B(n728), .Z(n725) );
  NANDN U637 ( .A(A[74]), .B(B[74]), .Z(n728) );
  NAND U638 ( .A(n729), .B(n730), .Z(n727) );
  NANDN U639 ( .A(B[74]), .B(A[74]), .Z(n730) );
  AND U640 ( .A(n731), .B(n732), .Z(n729) );
  NAND U641 ( .A(n733), .B(n734), .Z(n732) );
  NANDN U642 ( .A(A[73]), .B(B[73]), .Z(n734) );
  AND U643 ( .A(n735), .B(n736), .Z(n733) );
  NANDN U644 ( .A(A[72]), .B(B[72]), .Z(n736) );
  NAND U645 ( .A(n737), .B(n738), .Z(n735) );
  NANDN U646 ( .A(B[72]), .B(A[72]), .Z(n738) );
  AND U647 ( .A(n739), .B(n740), .Z(n737) );
  NAND U648 ( .A(n741), .B(n742), .Z(n740) );
  NANDN U649 ( .A(A[71]), .B(B[71]), .Z(n742) );
  AND U650 ( .A(n743), .B(n744), .Z(n741) );
  NANDN U651 ( .A(A[70]), .B(B[70]), .Z(n744) );
  NAND U652 ( .A(n745), .B(n746), .Z(n743) );
  NANDN U653 ( .A(B[70]), .B(A[70]), .Z(n746) );
  AND U654 ( .A(n747), .B(n748), .Z(n745) );
  NAND U655 ( .A(n749), .B(n750), .Z(n748) );
  NANDN U656 ( .A(A[69]), .B(B[69]), .Z(n750) );
  AND U657 ( .A(n751), .B(n752), .Z(n749) );
  NANDN U658 ( .A(A[68]), .B(B[68]), .Z(n752) );
  NAND U659 ( .A(n753), .B(n754), .Z(n751) );
  NANDN U660 ( .A(B[68]), .B(A[68]), .Z(n754) );
  AND U661 ( .A(n755), .B(n756), .Z(n753) );
  NAND U662 ( .A(n757), .B(n758), .Z(n756) );
  NANDN U663 ( .A(A[67]), .B(B[67]), .Z(n758) );
  AND U664 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U665 ( .A(A[66]), .B(B[66]), .Z(n760) );
  NAND U666 ( .A(n761), .B(n762), .Z(n759) );
  NANDN U667 ( .A(B[66]), .B(A[66]), .Z(n762) );
  AND U668 ( .A(n763), .B(n764), .Z(n761) );
  NAND U669 ( .A(n765), .B(n766), .Z(n764) );
  NANDN U670 ( .A(A[65]), .B(B[65]), .Z(n766) );
  AND U671 ( .A(n767), .B(n768), .Z(n765) );
  NANDN U672 ( .A(A[64]), .B(B[64]), .Z(n768) );
  NAND U673 ( .A(n769), .B(n770), .Z(n767) );
  NANDN U674 ( .A(B[64]), .B(A[64]), .Z(n770) );
  AND U675 ( .A(n771), .B(n772), .Z(n769) );
  NAND U676 ( .A(n773), .B(n774), .Z(n772) );
  NANDN U677 ( .A(A[63]), .B(B[63]), .Z(n774) );
  AND U678 ( .A(n775), .B(n776), .Z(n773) );
  NANDN U679 ( .A(A[62]), .B(B[62]), .Z(n776) );
  NAND U680 ( .A(n777), .B(n778), .Z(n775) );
  NANDN U681 ( .A(B[62]), .B(A[62]), .Z(n778) );
  AND U682 ( .A(n779), .B(n780), .Z(n777) );
  NAND U683 ( .A(n781), .B(n782), .Z(n780) );
  NANDN U684 ( .A(A[61]), .B(B[61]), .Z(n782) );
  AND U685 ( .A(n783), .B(n784), .Z(n781) );
  NANDN U686 ( .A(A[60]), .B(B[60]), .Z(n784) );
  NAND U687 ( .A(n785), .B(n786), .Z(n783) );
  NANDN U688 ( .A(B[60]), .B(A[60]), .Z(n786) );
  AND U689 ( .A(n787), .B(n788), .Z(n785) );
  NAND U690 ( .A(n789), .B(n790), .Z(n788) );
  NANDN U691 ( .A(A[59]), .B(B[59]), .Z(n790) );
  AND U692 ( .A(n791), .B(n792), .Z(n789) );
  NANDN U693 ( .A(A[58]), .B(B[58]), .Z(n792) );
  NAND U694 ( .A(n793), .B(n794), .Z(n791) );
  NANDN U695 ( .A(B[58]), .B(A[58]), .Z(n794) );
  AND U696 ( .A(n795), .B(n796), .Z(n793) );
  NAND U697 ( .A(n797), .B(n798), .Z(n796) );
  NANDN U698 ( .A(A[57]), .B(B[57]), .Z(n798) );
  AND U699 ( .A(n799), .B(n800), .Z(n797) );
  NANDN U700 ( .A(A[56]), .B(B[56]), .Z(n800) );
  NAND U701 ( .A(n801), .B(n802), .Z(n799) );
  NANDN U702 ( .A(B[56]), .B(A[56]), .Z(n802) );
  AND U703 ( .A(n803), .B(n804), .Z(n801) );
  NAND U704 ( .A(n805), .B(n806), .Z(n804) );
  NANDN U705 ( .A(A[55]), .B(B[55]), .Z(n806) );
  AND U706 ( .A(n807), .B(n808), .Z(n805) );
  NANDN U707 ( .A(A[54]), .B(B[54]), .Z(n808) );
  NAND U708 ( .A(n809), .B(n810), .Z(n807) );
  NANDN U709 ( .A(B[54]), .B(A[54]), .Z(n810) );
  AND U710 ( .A(n811), .B(n812), .Z(n809) );
  NAND U711 ( .A(n813), .B(n814), .Z(n812) );
  NANDN U712 ( .A(A[53]), .B(B[53]), .Z(n814) );
  AND U713 ( .A(n815), .B(n816), .Z(n813) );
  NANDN U714 ( .A(A[52]), .B(B[52]), .Z(n816) );
  NAND U715 ( .A(n817), .B(n818), .Z(n815) );
  NANDN U716 ( .A(B[52]), .B(A[52]), .Z(n818) );
  AND U717 ( .A(n819), .B(n820), .Z(n817) );
  NAND U718 ( .A(n821), .B(n822), .Z(n820) );
  NANDN U719 ( .A(A[51]), .B(B[51]), .Z(n822) );
  AND U720 ( .A(n823), .B(n824), .Z(n821) );
  NANDN U721 ( .A(A[50]), .B(B[50]), .Z(n824) );
  NAND U722 ( .A(n825), .B(n826), .Z(n823) );
  NANDN U723 ( .A(B[50]), .B(A[50]), .Z(n826) );
  AND U724 ( .A(n827), .B(n828), .Z(n825) );
  NAND U725 ( .A(n829), .B(n830), .Z(n828) );
  NANDN U726 ( .A(A[49]), .B(B[49]), .Z(n830) );
  AND U727 ( .A(n831), .B(n832), .Z(n829) );
  NANDN U728 ( .A(A[48]), .B(B[48]), .Z(n832) );
  NAND U729 ( .A(n833), .B(n834), .Z(n831) );
  NANDN U730 ( .A(B[48]), .B(A[48]), .Z(n834) );
  AND U731 ( .A(n835), .B(n836), .Z(n833) );
  NAND U732 ( .A(n837), .B(n838), .Z(n836) );
  NANDN U733 ( .A(A[47]), .B(B[47]), .Z(n838) );
  AND U734 ( .A(n839), .B(n840), .Z(n837) );
  NANDN U735 ( .A(A[46]), .B(B[46]), .Z(n840) );
  NAND U736 ( .A(n841), .B(n842), .Z(n839) );
  NANDN U737 ( .A(B[46]), .B(A[46]), .Z(n842) );
  AND U738 ( .A(n843), .B(n844), .Z(n841) );
  NAND U739 ( .A(n845), .B(n846), .Z(n844) );
  NANDN U740 ( .A(A[45]), .B(B[45]), .Z(n846) );
  AND U741 ( .A(n847), .B(n848), .Z(n845) );
  NANDN U742 ( .A(A[44]), .B(B[44]), .Z(n848) );
  NAND U743 ( .A(n849), .B(n850), .Z(n847) );
  NANDN U744 ( .A(B[44]), .B(A[44]), .Z(n850) );
  AND U745 ( .A(n851), .B(n852), .Z(n849) );
  NAND U746 ( .A(n853), .B(n854), .Z(n852) );
  NANDN U747 ( .A(A[43]), .B(B[43]), .Z(n854) );
  AND U748 ( .A(n855), .B(n856), .Z(n853) );
  NANDN U749 ( .A(A[42]), .B(B[42]), .Z(n856) );
  NAND U750 ( .A(n857), .B(n858), .Z(n855) );
  NANDN U751 ( .A(B[42]), .B(A[42]), .Z(n858) );
  AND U752 ( .A(n859), .B(n860), .Z(n857) );
  NAND U753 ( .A(n861), .B(n862), .Z(n860) );
  NANDN U754 ( .A(A[41]), .B(B[41]), .Z(n862) );
  AND U755 ( .A(n863), .B(n864), .Z(n861) );
  NANDN U756 ( .A(A[40]), .B(B[40]), .Z(n864) );
  NAND U757 ( .A(n865), .B(n866), .Z(n863) );
  NANDN U758 ( .A(B[40]), .B(A[40]), .Z(n866) );
  AND U759 ( .A(n867), .B(n868), .Z(n865) );
  NAND U760 ( .A(n869), .B(n870), .Z(n868) );
  NANDN U761 ( .A(A[39]), .B(B[39]), .Z(n870) );
  AND U762 ( .A(n871), .B(n872), .Z(n869) );
  NANDN U763 ( .A(A[38]), .B(B[38]), .Z(n872) );
  NAND U764 ( .A(n873), .B(n874), .Z(n871) );
  NANDN U765 ( .A(B[38]), .B(A[38]), .Z(n874) );
  AND U766 ( .A(n875), .B(n876), .Z(n873) );
  NAND U767 ( .A(n877), .B(n878), .Z(n876) );
  NANDN U768 ( .A(A[37]), .B(B[37]), .Z(n878) );
  AND U769 ( .A(n879), .B(n880), .Z(n877) );
  NANDN U770 ( .A(A[36]), .B(B[36]), .Z(n880) );
  NAND U771 ( .A(n881), .B(n882), .Z(n879) );
  NANDN U772 ( .A(B[36]), .B(A[36]), .Z(n882) );
  AND U773 ( .A(n883), .B(n884), .Z(n881) );
  NAND U774 ( .A(n885), .B(n886), .Z(n884) );
  NANDN U775 ( .A(A[35]), .B(B[35]), .Z(n886) );
  AND U776 ( .A(n887), .B(n888), .Z(n885) );
  NANDN U777 ( .A(A[34]), .B(B[34]), .Z(n888) );
  NAND U778 ( .A(n889), .B(n890), .Z(n887) );
  NANDN U779 ( .A(B[34]), .B(A[34]), .Z(n890) );
  AND U780 ( .A(n891), .B(n892), .Z(n889) );
  NAND U781 ( .A(n893), .B(n894), .Z(n892) );
  NANDN U782 ( .A(A[33]), .B(B[33]), .Z(n894) );
  AND U783 ( .A(n895), .B(n896), .Z(n893) );
  NANDN U784 ( .A(A[32]), .B(B[32]), .Z(n896) );
  NAND U785 ( .A(n897), .B(n898), .Z(n895) );
  NANDN U786 ( .A(B[32]), .B(A[32]), .Z(n898) );
  AND U787 ( .A(n899), .B(n900), .Z(n897) );
  NAND U788 ( .A(n901), .B(n902), .Z(n900) );
  NANDN U789 ( .A(A[31]), .B(B[31]), .Z(n902) );
  AND U790 ( .A(n903), .B(n904), .Z(n901) );
  NANDN U791 ( .A(A[30]), .B(B[30]), .Z(n904) );
  NAND U792 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U793 ( .A(B[30]), .B(A[30]), .Z(n906) );
  AND U794 ( .A(n907), .B(n908), .Z(n905) );
  NAND U795 ( .A(n909), .B(n910), .Z(n908) );
  NANDN U796 ( .A(A[29]), .B(B[29]), .Z(n910) );
  AND U797 ( .A(n911), .B(n912), .Z(n909) );
  NANDN U798 ( .A(A[28]), .B(B[28]), .Z(n912) );
  NAND U799 ( .A(n913), .B(n914), .Z(n911) );
  NANDN U800 ( .A(B[28]), .B(A[28]), .Z(n914) );
  AND U801 ( .A(n915), .B(n916), .Z(n913) );
  NAND U802 ( .A(n917), .B(n918), .Z(n916) );
  NANDN U803 ( .A(A[27]), .B(B[27]), .Z(n918) );
  AND U804 ( .A(n919), .B(n920), .Z(n917) );
  NANDN U805 ( .A(A[26]), .B(B[26]), .Z(n920) );
  NAND U806 ( .A(n921), .B(n922), .Z(n919) );
  NANDN U807 ( .A(B[26]), .B(A[26]), .Z(n922) );
  AND U808 ( .A(n923), .B(n924), .Z(n921) );
  NAND U809 ( .A(n925), .B(n926), .Z(n924) );
  NANDN U810 ( .A(A[25]), .B(B[25]), .Z(n926) );
  AND U811 ( .A(n927), .B(n928), .Z(n925) );
  NANDN U812 ( .A(A[24]), .B(B[24]), .Z(n928) );
  NAND U813 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U814 ( .A(B[24]), .B(A[24]), .Z(n930) );
  AND U815 ( .A(n931), .B(n932), .Z(n929) );
  NAND U816 ( .A(n933), .B(n934), .Z(n932) );
  NANDN U817 ( .A(A[23]), .B(B[23]), .Z(n934) );
  AND U818 ( .A(n935), .B(n936), .Z(n933) );
  NANDN U819 ( .A(A[22]), .B(B[22]), .Z(n936) );
  NAND U820 ( .A(n937), .B(n938), .Z(n935) );
  NANDN U821 ( .A(B[22]), .B(A[22]), .Z(n938) );
  AND U822 ( .A(n939), .B(n940), .Z(n937) );
  NAND U823 ( .A(n941), .B(n942), .Z(n940) );
  NANDN U824 ( .A(A[21]), .B(B[21]), .Z(n942) );
  AND U825 ( .A(n943), .B(n944), .Z(n941) );
  NANDN U826 ( .A(A[20]), .B(B[20]), .Z(n944) );
  NAND U827 ( .A(n945), .B(n946), .Z(n943) );
  NANDN U828 ( .A(B[20]), .B(A[20]), .Z(n946) );
  AND U829 ( .A(n947), .B(n948), .Z(n945) );
  NAND U830 ( .A(n949), .B(n950), .Z(n948) );
  NANDN U831 ( .A(A[19]), .B(B[19]), .Z(n950) );
  AND U832 ( .A(n951), .B(n952), .Z(n949) );
  NANDN U833 ( .A(A[18]), .B(B[18]), .Z(n952) );
  NAND U834 ( .A(n953), .B(n954), .Z(n951) );
  NANDN U835 ( .A(B[18]), .B(A[18]), .Z(n954) );
  AND U836 ( .A(n955), .B(n956), .Z(n953) );
  NAND U837 ( .A(n957), .B(n958), .Z(n956) );
  NANDN U838 ( .A(A[17]), .B(B[17]), .Z(n958) );
  AND U839 ( .A(n959), .B(n960), .Z(n957) );
  NANDN U840 ( .A(A[16]), .B(B[16]), .Z(n960) );
  NAND U841 ( .A(n961), .B(n962), .Z(n959) );
  NANDN U842 ( .A(B[16]), .B(A[16]), .Z(n962) );
  AND U843 ( .A(n963), .B(n964), .Z(n961) );
  NAND U844 ( .A(n965), .B(n966), .Z(n964) );
  NANDN U845 ( .A(A[15]), .B(B[15]), .Z(n966) );
  AND U846 ( .A(n967), .B(n968), .Z(n965) );
  NANDN U847 ( .A(A[14]), .B(B[14]), .Z(n968) );
  NAND U848 ( .A(n969), .B(n970), .Z(n967) );
  NANDN U849 ( .A(B[14]), .B(A[14]), .Z(n970) );
  AND U850 ( .A(n971), .B(n972), .Z(n969) );
  NAND U851 ( .A(n973), .B(n974), .Z(n972) );
  NANDN U852 ( .A(A[13]), .B(B[13]), .Z(n974) );
  AND U853 ( .A(n975), .B(n976), .Z(n973) );
  NANDN U854 ( .A(A[12]), .B(B[12]), .Z(n976) );
  NAND U855 ( .A(n977), .B(n978), .Z(n975) );
  NANDN U856 ( .A(B[12]), .B(A[12]), .Z(n978) );
  AND U857 ( .A(n979), .B(n980), .Z(n977) );
  NAND U858 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U859 ( .A(A[11]), .B(B[11]), .Z(n982) );
  AND U860 ( .A(n983), .B(n984), .Z(n981) );
  NANDN U861 ( .A(A[10]), .B(B[10]), .Z(n984) );
  NAND U862 ( .A(n985), .B(n986), .Z(n983) );
  NANDN U863 ( .A(B[9]), .B(A[9]), .Z(n986) );
  AND U864 ( .A(n987), .B(n988), .Z(n985) );
  NAND U865 ( .A(n989), .B(n990), .Z(n988) );
  NANDN U866 ( .A(A[9]), .B(B[9]), .Z(n990) );
  AND U867 ( .A(n991), .B(n992), .Z(n989) );
  NANDN U868 ( .A(A[8]), .B(B[8]), .Z(n992) );
  NAND U869 ( .A(n993), .B(n994), .Z(n991) );
  NANDN U870 ( .A(B[8]), .B(A[8]), .Z(n994) );
  AND U871 ( .A(n995), .B(n996), .Z(n993) );
  NAND U872 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U873 ( .A(A[7]), .B(B[7]), .Z(n998) );
  AND U874 ( .A(n999), .B(n1000), .Z(n997) );
  NANDN U875 ( .A(A[6]), .B(B[6]), .Z(n1000) );
  NAND U876 ( .A(n1001), .B(n1002), .Z(n999) );
  NANDN U877 ( .A(B[6]), .B(A[6]), .Z(n1002) );
  AND U878 ( .A(n1003), .B(n1004), .Z(n1001) );
  NAND U879 ( .A(n1005), .B(n1006), .Z(n1004) );
  NANDN U880 ( .A(A[5]), .B(B[5]), .Z(n1006) );
  AND U881 ( .A(n1007), .B(n1008), .Z(n1005) );
  NANDN U882 ( .A(A[4]), .B(B[4]), .Z(n1008) );
  NAND U883 ( .A(n1009), .B(n1010), .Z(n1007) );
  NANDN U884 ( .A(B[4]), .B(A[4]), .Z(n1010) );
  AND U885 ( .A(n1011), .B(n1012), .Z(n1009) );
  NAND U886 ( .A(n1013), .B(n1014), .Z(n1012) );
  NANDN U887 ( .A(A[3]), .B(B[3]), .Z(n1014) );
  AND U888 ( .A(n1015), .B(n1016), .Z(n1013) );
  NANDN U889 ( .A(A[2]), .B(B[2]), .Z(n1016) );
  NAND U890 ( .A(n1017), .B(n1018), .Z(n1015) );
  NANDN U891 ( .A(B[2]), .B(A[2]), .Z(n1018) );
  AND U892 ( .A(n1019), .B(n1020), .Z(n1017) );
  NAND U893 ( .A(n1021), .B(A[0]), .Z(n1020) );
  ANDN U894 ( .B(n1022), .A(B[0]), .Z(n1021) );
  NANDN U895 ( .A(A[1]), .B(B[1]), .Z(n1022) );
  NANDN U896 ( .A(B[1]), .B(A[1]), .Z(n1019) );
  NANDN U897 ( .A(B[3]), .B(A[3]), .Z(n1011) );
  NANDN U898 ( .A(B[5]), .B(A[5]), .Z(n1003) );
  NANDN U899 ( .A(B[7]), .B(A[7]), .Z(n995) );
  NANDN U900 ( .A(B[10]), .B(A[10]), .Z(n987) );
  NANDN U901 ( .A(B[11]), .B(A[11]), .Z(n979) );
  NANDN U902 ( .A(B[13]), .B(A[13]), .Z(n971) );
  NANDN U903 ( .A(B[15]), .B(A[15]), .Z(n963) );
  NANDN U904 ( .A(B[17]), .B(A[17]), .Z(n955) );
  NANDN U905 ( .A(B[19]), .B(A[19]), .Z(n947) );
  NANDN U906 ( .A(B[21]), .B(A[21]), .Z(n939) );
  NANDN U907 ( .A(B[23]), .B(A[23]), .Z(n931) );
  NANDN U908 ( .A(B[25]), .B(A[25]), .Z(n923) );
  NANDN U909 ( .A(B[27]), .B(A[27]), .Z(n915) );
  NANDN U910 ( .A(B[29]), .B(A[29]), .Z(n907) );
  NANDN U911 ( .A(B[31]), .B(A[31]), .Z(n899) );
  NANDN U912 ( .A(B[33]), .B(A[33]), .Z(n891) );
  NANDN U913 ( .A(B[35]), .B(A[35]), .Z(n883) );
  NANDN U914 ( .A(B[37]), .B(A[37]), .Z(n875) );
  NANDN U915 ( .A(B[39]), .B(A[39]), .Z(n867) );
  NANDN U916 ( .A(B[41]), .B(A[41]), .Z(n859) );
  NANDN U917 ( .A(B[43]), .B(A[43]), .Z(n851) );
  NANDN U918 ( .A(B[45]), .B(A[45]), .Z(n843) );
  NANDN U919 ( .A(B[47]), .B(A[47]), .Z(n835) );
  NANDN U920 ( .A(B[49]), .B(A[49]), .Z(n827) );
  NANDN U921 ( .A(B[51]), .B(A[51]), .Z(n819) );
  NANDN U922 ( .A(B[53]), .B(A[53]), .Z(n811) );
  NANDN U923 ( .A(B[55]), .B(A[55]), .Z(n803) );
  NANDN U924 ( .A(B[57]), .B(A[57]), .Z(n795) );
  NANDN U925 ( .A(B[59]), .B(A[59]), .Z(n787) );
  NANDN U926 ( .A(B[61]), .B(A[61]), .Z(n779) );
  NANDN U927 ( .A(B[63]), .B(A[63]), .Z(n771) );
  NANDN U928 ( .A(B[65]), .B(A[65]), .Z(n763) );
  NANDN U929 ( .A(B[67]), .B(A[67]), .Z(n755) );
  NANDN U930 ( .A(B[69]), .B(A[69]), .Z(n747) );
  NANDN U931 ( .A(B[71]), .B(A[71]), .Z(n739) );
  NANDN U932 ( .A(B[73]), .B(A[73]), .Z(n731) );
  NANDN U933 ( .A(B[75]), .B(A[75]), .Z(n723) );
  NANDN U934 ( .A(B[77]), .B(A[77]), .Z(n715) );
  NANDN U935 ( .A(B[79]), .B(A[79]), .Z(n707) );
  NANDN U936 ( .A(B[81]), .B(A[81]), .Z(n699) );
  NANDN U937 ( .A(B[83]), .B(A[83]), .Z(n691) );
  NANDN U938 ( .A(B[85]), .B(A[85]), .Z(n683) );
  NANDN U939 ( .A(B[87]), .B(A[87]), .Z(n675) );
  NANDN U940 ( .A(B[89]), .B(A[89]), .Z(n667) );
  NANDN U941 ( .A(B[91]), .B(A[91]), .Z(n659) );
  NANDN U942 ( .A(B[93]), .B(A[93]), .Z(n651) );
  NANDN U943 ( .A(B[95]), .B(A[95]), .Z(n643) );
  NANDN U944 ( .A(B[97]), .B(A[97]), .Z(n635) );
  NANDN U945 ( .A(B[100]), .B(A[100]), .Z(n627) );
  NANDN U946 ( .A(B[101]), .B(A[101]), .Z(n619) );
  NANDN U947 ( .A(B[103]), .B(A[103]), .Z(n611) );
  NANDN U948 ( .A(B[105]), .B(A[105]), .Z(n603) );
  NANDN U949 ( .A(B[107]), .B(A[107]), .Z(n595) );
  NANDN U950 ( .A(B[109]), .B(A[109]), .Z(n587) );
  NANDN U951 ( .A(B[111]), .B(A[111]), .Z(n579) );
  NANDN U952 ( .A(B[113]), .B(A[113]), .Z(n571) );
  NANDN U953 ( .A(B[115]), .B(A[115]), .Z(n563) );
  NANDN U954 ( .A(B[117]), .B(A[117]), .Z(n555) );
  NANDN U955 ( .A(B[119]), .B(A[119]), .Z(n547) );
  NANDN U956 ( .A(B[121]), .B(A[121]), .Z(n539) );
  NANDN U957 ( .A(B[123]), .B(A[123]), .Z(n531) );
  NANDN U958 ( .A(B[125]), .B(A[125]), .Z(n523) );
  NANDN U959 ( .A(B[127]), .B(A[127]), .Z(n515) );
  NANDN U960 ( .A(B[129]), .B(A[129]), .Z(n507) );
  NANDN U961 ( .A(B[131]), .B(A[131]), .Z(n499) );
  NANDN U962 ( .A(B[133]), .B(A[133]), .Z(n491) );
  NANDN U963 ( .A(B[135]), .B(A[135]), .Z(n483) );
  NANDN U964 ( .A(B[137]), .B(A[137]), .Z(n475) );
  NANDN U965 ( .A(B[139]), .B(A[139]), .Z(n467) );
  NANDN U966 ( .A(B[141]), .B(A[141]), .Z(n459) );
  NANDN U967 ( .A(B[143]), .B(A[143]), .Z(n451) );
  NANDN U968 ( .A(B[145]), .B(A[145]), .Z(n443) );
  NANDN U969 ( .A(B[147]), .B(A[147]), .Z(n435) );
  NANDN U970 ( .A(B[149]), .B(A[149]), .Z(n427) );
  NANDN U971 ( .A(B[151]), .B(A[151]), .Z(n419) );
  NANDN U972 ( .A(B[153]), .B(A[153]), .Z(n411) );
  NANDN U973 ( .A(B[155]), .B(A[155]), .Z(n403) );
  NANDN U974 ( .A(B[157]), .B(A[157]), .Z(n395) );
  NANDN U975 ( .A(B[159]), .B(A[159]), .Z(n387) );
  NANDN U976 ( .A(B[161]), .B(A[161]), .Z(n379) );
  NANDN U977 ( .A(B[163]), .B(A[163]), .Z(n371) );
  NANDN U978 ( .A(B[165]), .B(A[165]), .Z(n363) );
  NANDN U979 ( .A(B[167]), .B(A[167]), .Z(n355) );
  NANDN U980 ( .A(B[169]), .B(A[169]), .Z(n347) );
  NANDN U981 ( .A(B[171]), .B(A[171]), .Z(n339) );
  NANDN U982 ( .A(B[173]), .B(A[173]), .Z(n331) );
  NANDN U983 ( .A(B[175]), .B(A[175]), .Z(n323) );
  NANDN U984 ( .A(B[177]), .B(A[177]), .Z(n315) );
  NANDN U985 ( .A(B[179]), .B(A[179]), .Z(n307) );
  NANDN U986 ( .A(B[181]), .B(A[181]), .Z(n299) );
  NANDN U987 ( .A(B[183]), .B(A[183]), .Z(n291) );
  NANDN U988 ( .A(B[185]), .B(A[185]), .Z(n283) );
  NANDN U989 ( .A(B[187]), .B(A[187]), .Z(n275) );
  NANDN U990 ( .A(B[189]), .B(A[189]), .Z(n267) );
  NANDN U991 ( .A(B[191]), .B(A[191]), .Z(n259) );
  NANDN U992 ( .A(B[193]), .B(A[193]), .Z(n251) );
  NANDN U993 ( .A(B[195]), .B(A[195]), .Z(n243) );
  NANDN U994 ( .A(B[197]), .B(A[197]), .Z(n235) );
  NANDN U995 ( .A(B[199]), .B(A[199]), .Z(n227) );
  NANDN U996 ( .A(B[201]), .B(A[201]), .Z(n219) );
  NANDN U997 ( .A(B[203]), .B(A[203]), .Z(n211) );
  NANDN U998 ( .A(B[205]), .B(A[205]), .Z(n203) );
  NANDN U999 ( .A(B[207]), .B(A[207]), .Z(n195) );
  NANDN U1000 ( .A(B[209]), .B(A[209]), .Z(n187) );
  NANDN U1001 ( .A(B[211]), .B(A[211]), .Z(n179) );
  NANDN U1002 ( .A(B[213]), .B(A[213]), .Z(n171) );
  NANDN U1003 ( .A(B[215]), .B(A[215]), .Z(n163) );
  NANDN U1004 ( .A(B[217]), .B(A[217]), .Z(n155) );
  NANDN U1005 ( .A(B[219]), .B(A[219]), .Z(n147) );
  NANDN U1006 ( .A(B[221]), .B(A[221]), .Z(n139) );
  NANDN U1007 ( .A(B[223]), .B(A[223]), .Z(n131) );
  NANDN U1008 ( .A(B[225]), .B(A[225]), .Z(n123) );
  NANDN U1009 ( .A(B[227]), .B(A[227]), .Z(n115) );
  NANDN U1010 ( .A(B[229]), .B(A[229]), .Z(n107) );
  NANDN U1011 ( .A(B[231]), .B(A[231]), .Z(n99) );
  NANDN U1012 ( .A(B[233]), .B(A[233]), .Z(n91) );
  NANDN U1013 ( .A(B[235]), .B(A[235]), .Z(n83) );
  NANDN U1014 ( .A(B[237]), .B(A[237]), .Z(n75) );
  NANDN U1015 ( .A(B[239]), .B(A[239]), .Z(n67) );
  NANDN U1016 ( .A(B[241]), .B(A[241]), .Z(n59) );
  NANDN U1017 ( .A(B[243]), .B(A[243]), .Z(n51) );
  NANDN U1018 ( .A(B[245]), .B(A[245]), .Z(n43) );
  NANDN U1019 ( .A(B[247]), .B(A[247]), .Z(n35) );
  NANDN U1020 ( .A(B[249]), .B(A[249]), .Z(n27) );
  NANDN U1021 ( .A(B[251]), .B(A[251]), .Z(n19) );
  NANDN U1022 ( .A(B[253]), .B(A[253]), .Z(n11) );
  NANDN U1023 ( .A(A[255]), .B(B[255]), .Z(n3) );
endmodule


module modmult_step_N256_4_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280;

  IV U1 ( .A(A[1]), .Z(n1) );
  IV U2 ( .A(n1279), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(DIFF[9]) );
  XOR U4 ( .A(B[9]), .B(A[9]), .Z(n4) );
  XNOR U5 ( .A(n5), .B(n6), .Z(DIFF[99]) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(DIFF[98]) );
  XOR U8 ( .A(B[98]), .B(A[98]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(DIFF[97]) );
  XOR U10 ( .A(B[97]), .B(A[97]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(DIFF[96]) );
  XOR U12 ( .A(B[96]), .B(A[96]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(DIFF[95]) );
  XOR U14 ( .A(B[95]), .B(A[95]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(DIFF[94]) );
  XOR U16 ( .A(B[94]), .B(A[94]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(DIFF[93]) );
  XOR U18 ( .A(B[93]), .B(A[93]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(DIFF[92]) );
  XOR U20 ( .A(B[92]), .B(A[92]), .Z(n20) );
  XOR U21 ( .A(n21), .B(n22), .Z(DIFF[91]) );
  XOR U22 ( .A(B[91]), .B(A[91]), .Z(n22) );
  XOR U23 ( .A(n23), .B(n24), .Z(DIFF[90]) );
  XOR U24 ( .A(B[90]), .B(A[90]), .Z(n24) );
  XOR U25 ( .A(n25), .B(n26), .Z(DIFF[8]) );
  XOR U26 ( .A(B[8]), .B(A[8]), .Z(n26) );
  XOR U27 ( .A(n27), .B(n28), .Z(DIFF[89]) );
  XOR U28 ( .A(B[89]), .B(A[89]), .Z(n28) );
  XOR U29 ( .A(n29), .B(n30), .Z(DIFF[88]) );
  XOR U30 ( .A(B[88]), .B(A[88]), .Z(n30) );
  XOR U31 ( .A(n31), .B(n32), .Z(DIFF[87]) );
  XOR U32 ( .A(B[87]), .B(A[87]), .Z(n32) );
  XOR U33 ( .A(n33), .B(n34), .Z(DIFF[86]) );
  XOR U34 ( .A(B[86]), .B(A[86]), .Z(n34) );
  XOR U35 ( .A(n35), .B(n36), .Z(DIFF[85]) );
  XOR U36 ( .A(B[85]), .B(A[85]), .Z(n36) );
  XOR U37 ( .A(n37), .B(n38), .Z(DIFF[84]) );
  XOR U38 ( .A(B[84]), .B(A[84]), .Z(n38) );
  XOR U39 ( .A(n39), .B(n40), .Z(DIFF[83]) );
  XOR U40 ( .A(B[83]), .B(A[83]), .Z(n40) );
  XOR U41 ( .A(n41), .B(n42), .Z(DIFF[82]) );
  XOR U42 ( .A(B[82]), .B(A[82]), .Z(n42) );
  XOR U43 ( .A(n43), .B(n44), .Z(DIFF[81]) );
  XOR U44 ( .A(B[81]), .B(A[81]), .Z(n44) );
  XOR U45 ( .A(n45), .B(n46), .Z(DIFF[80]) );
  XOR U46 ( .A(B[80]), .B(A[80]), .Z(n46) );
  XOR U47 ( .A(n47), .B(n48), .Z(DIFF[7]) );
  XOR U48 ( .A(B[7]), .B(A[7]), .Z(n48) );
  XOR U49 ( .A(n49), .B(n50), .Z(DIFF[79]) );
  XOR U50 ( .A(B[79]), .B(A[79]), .Z(n50) );
  XOR U51 ( .A(n51), .B(n52), .Z(DIFF[78]) );
  XOR U52 ( .A(B[78]), .B(A[78]), .Z(n52) );
  XOR U53 ( .A(n53), .B(n54), .Z(DIFF[77]) );
  XOR U54 ( .A(B[77]), .B(A[77]), .Z(n54) );
  XOR U55 ( .A(n55), .B(n56), .Z(DIFF[76]) );
  XOR U56 ( .A(B[76]), .B(A[76]), .Z(n56) );
  XOR U57 ( .A(n57), .B(n58), .Z(DIFF[75]) );
  XOR U58 ( .A(B[75]), .B(A[75]), .Z(n58) );
  XOR U59 ( .A(n59), .B(n60), .Z(DIFF[74]) );
  XOR U60 ( .A(B[74]), .B(A[74]), .Z(n60) );
  XOR U61 ( .A(n61), .B(n62), .Z(DIFF[73]) );
  XOR U62 ( .A(B[73]), .B(A[73]), .Z(n62) );
  XOR U63 ( .A(n63), .B(n64), .Z(DIFF[72]) );
  XOR U64 ( .A(B[72]), .B(A[72]), .Z(n64) );
  XOR U65 ( .A(n65), .B(n66), .Z(DIFF[71]) );
  XOR U66 ( .A(B[71]), .B(A[71]), .Z(n66) );
  XOR U67 ( .A(n67), .B(n68), .Z(DIFF[70]) );
  XOR U68 ( .A(B[70]), .B(A[70]), .Z(n68) );
  XOR U69 ( .A(n69), .B(n70), .Z(DIFF[6]) );
  XOR U70 ( .A(B[6]), .B(A[6]), .Z(n70) );
  XOR U71 ( .A(n71), .B(n72), .Z(DIFF[69]) );
  XOR U72 ( .A(B[69]), .B(A[69]), .Z(n72) );
  XOR U73 ( .A(n73), .B(n74), .Z(DIFF[68]) );
  XOR U74 ( .A(B[68]), .B(A[68]), .Z(n74) );
  XOR U75 ( .A(n75), .B(n76), .Z(DIFF[67]) );
  XOR U76 ( .A(B[67]), .B(A[67]), .Z(n76) );
  XOR U77 ( .A(n77), .B(n78), .Z(DIFF[66]) );
  XOR U78 ( .A(B[66]), .B(A[66]), .Z(n78) );
  XOR U79 ( .A(n79), .B(n80), .Z(DIFF[65]) );
  XOR U80 ( .A(B[65]), .B(A[65]), .Z(n80) );
  XOR U81 ( .A(n81), .B(n82), .Z(DIFF[64]) );
  XOR U82 ( .A(B[64]), .B(A[64]), .Z(n82) );
  XOR U83 ( .A(n83), .B(n84), .Z(DIFF[63]) );
  XOR U84 ( .A(B[63]), .B(A[63]), .Z(n84) );
  XOR U85 ( .A(n85), .B(n86), .Z(DIFF[62]) );
  XOR U86 ( .A(B[62]), .B(A[62]), .Z(n86) );
  XOR U87 ( .A(n87), .B(n88), .Z(DIFF[61]) );
  XOR U88 ( .A(B[61]), .B(A[61]), .Z(n88) );
  XOR U89 ( .A(n89), .B(n90), .Z(DIFF[60]) );
  XOR U90 ( .A(B[60]), .B(A[60]), .Z(n90) );
  XOR U91 ( .A(n91), .B(n92), .Z(DIFF[5]) );
  XOR U92 ( .A(B[5]), .B(A[5]), .Z(n92) );
  XOR U93 ( .A(n93), .B(n94), .Z(DIFF[59]) );
  XOR U94 ( .A(B[59]), .B(A[59]), .Z(n94) );
  XOR U95 ( .A(n95), .B(n96), .Z(DIFF[58]) );
  XOR U96 ( .A(B[58]), .B(A[58]), .Z(n96) );
  XOR U97 ( .A(n97), .B(n98), .Z(DIFF[57]) );
  XOR U98 ( .A(B[57]), .B(A[57]), .Z(n98) );
  XOR U99 ( .A(n99), .B(n100), .Z(DIFF[56]) );
  XOR U100 ( .A(B[56]), .B(A[56]), .Z(n100) );
  XOR U101 ( .A(n101), .B(n102), .Z(DIFF[55]) );
  XOR U102 ( .A(B[55]), .B(A[55]), .Z(n102) );
  XOR U103 ( .A(n103), .B(n104), .Z(DIFF[54]) );
  XOR U104 ( .A(B[54]), .B(A[54]), .Z(n104) );
  XOR U105 ( .A(n105), .B(n106), .Z(DIFF[53]) );
  XOR U106 ( .A(B[53]), .B(A[53]), .Z(n106) );
  XOR U107 ( .A(n107), .B(n108), .Z(DIFF[52]) );
  XOR U108 ( .A(B[52]), .B(A[52]), .Z(n108) );
  XOR U109 ( .A(n109), .B(n110), .Z(DIFF[51]) );
  XOR U110 ( .A(B[51]), .B(A[51]), .Z(n110) );
  XOR U111 ( .A(n111), .B(n112), .Z(DIFF[50]) );
  XOR U112 ( .A(B[50]), .B(A[50]), .Z(n112) );
  XOR U113 ( .A(n113), .B(n114), .Z(DIFF[4]) );
  XOR U114 ( .A(B[4]), .B(A[4]), .Z(n114) );
  XOR U115 ( .A(n115), .B(n116), .Z(DIFF[49]) );
  XOR U116 ( .A(B[49]), .B(A[49]), .Z(n116) );
  XOR U117 ( .A(n117), .B(n118), .Z(DIFF[48]) );
  XOR U118 ( .A(B[48]), .B(A[48]), .Z(n118) );
  XOR U119 ( .A(n119), .B(n120), .Z(DIFF[47]) );
  XOR U120 ( .A(B[47]), .B(A[47]), .Z(n120) );
  XOR U121 ( .A(n121), .B(n122), .Z(DIFF[46]) );
  XOR U122 ( .A(B[46]), .B(A[46]), .Z(n122) );
  XOR U123 ( .A(n123), .B(n124), .Z(DIFF[45]) );
  XOR U124 ( .A(B[45]), .B(A[45]), .Z(n124) );
  XOR U125 ( .A(n125), .B(n126), .Z(DIFF[44]) );
  XOR U126 ( .A(B[44]), .B(A[44]), .Z(n126) );
  XOR U127 ( .A(n127), .B(n128), .Z(DIFF[43]) );
  XOR U128 ( .A(B[43]), .B(A[43]), .Z(n128) );
  XOR U129 ( .A(n129), .B(n130), .Z(DIFF[42]) );
  XOR U130 ( .A(B[42]), .B(A[42]), .Z(n130) );
  XOR U131 ( .A(n131), .B(n132), .Z(DIFF[41]) );
  XOR U132 ( .A(B[41]), .B(A[41]), .Z(n132) );
  XOR U133 ( .A(n133), .B(n134), .Z(DIFF[40]) );
  XOR U134 ( .A(B[40]), .B(A[40]), .Z(n134) );
  XOR U135 ( .A(n135), .B(n136), .Z(DIFF[3]) );
  XOR U136 ( .A(B[3]), .B(A[3]), .Z(n136) );
  XOR U137 ( .A(n137), .B(n138), .Z(DIFF[39]) );
  XOR U138 ( .A(B[39]), .B(A[39]), .Z(n138) );
  XOR U139 ( .A(n139), .B(n140), .Z(DIFF[38]) );
  XOR U140 ( .A(B[38]), .B(A[38]), .Z(n140) );
  XOR U141 ( .A(n141), .B(n142), .Z(DIFF[37]) );
  XOR U142 ( .A(B[37]), .B(A[37]), .Z(n142) );
  XOR U143 ( .A(n143), .B(n144), .Z(DIFF[36]) );
  XOR U144 ( .A(B[36]), .B(A[36]), .Z(n144) );
  XOR U145 ( .A(n145), .B(n146), .Z(DIFF[35]) );
  XOR U146 ( .A(B[35]), .B(A[35]), .Z(n146) );
  XOR U147 ( .A(n147), .B(n148), .Z(DIFF[34]) );
  XOR U148 ( .A(B[34]), .B(A[34]), .Z(n148) );
  XOR U149 ( .A(n149), .B(n150), .Z(DIFF[33]) );
  XOR U150 ( .A(B[33]), .B(A[33]), .Z(n150) );
  XOR U151 ( .A(n151), .B(n152), .Z(DIFF[32]) );
  XOR U152 ( .A(B[32]), .B(A[32]), .Z(n152) );
  XOR U153 ( .A(n153), .B(n154), .Z(DIFF[31]) );
  XOR U154 ( .A(B[31]), .B(A[31]), .Z(n154) );
  XOR U155 ( .A(n155), .B(n156), .Z(DIFF[30]) );
  XOR U156 ( .A(B[30]), .B(A[30]), .Z(n156) );
  XOR U157 ( .A(n157), .B(n158), .Z(DIFF[2]) );
  XOR U158 ( .A(B[2]), .B(A[2]), .Z(n158) );
  XOR U159 ( .A(n159), .B(n160), .Z(DIFF[29]) );
  XOR U160 ( .A(B[29]), .B(A[29]), .Z(n160) );
  XOR U161 ( .A(n161), .B(n162), .Z(DIFF[28]) );
  XOR U162 ( .A(B[28]), .B(A[28]), .Z(n162) );
  XOR U163 ( .A(n163), .B(n164), .Z(DIFF[27]) );
  XOR U164 ( .A(B[27]), .B(A[27]), .Z(n164) );
  XOR U165 ( .A(n165), .B(n166), .Z(DIFF[26]) );
  XOR U166 ( .A(B[26]), .B(A[26]), .Z(n166) );
  XOR U167 ( .A(n167), .B(n168), .Z(DIFF[25]) );
  XOR U168 ( .A(B[25]), .B(A[25]), .Z(n168) );
  XOR U169 ( .A(A[257]), .B(n169), .Z(DIFF[257]) );
  ANDN U170 ( .B(n170), .A(A[256]), .Z(n169) );
  XOR U171 ( .A(A[256]), .B(n170), .Z(DIFF[256]) );
  AND U172 ( .A(n171), .B(n172), .Z(n170) );
  NANDN U173 ( .A(B[255]), .B(n173), .Z(n172) );
  NANDN U174 ( .A(A[255]), .B(n174), .Z(n173) );
  NANDN U175 ( .A(n174), .B(A[255]), .Z(n171) );
  XOR U176 ( .A(n174), .B(n175), .Z(DIFF[255]) );
  XOR U177 ( .A(B[255]), .B(A[255]), .Z(n175) );
  AND U178 ( .A(n176), .B(n177), .Z(n174) );
  NANDN U179 ( .A(B[254]), .B(n178), .Z(n177) );
  NANDN U180 ( .A(A[254]), .B(n179), .Z(n178) );
  NANDN U181 ( .A(n179), .B(A[254]), .Z(n176) );
  XOR U182 ( .A(n179), .B(n180), .Z(DIFF[254]) );
  XOR U183 ( .A(B[254]), .B(A[254]), .Z(n180) );
  AND U184 ( .A(n181), .B(n182), .Z(n179) );
  NANDN U185 ( .A(B[253]), .B(n183), .Z(n182) );
  NANDN U186 ( .A(A[253]), .B(n184), .Z(n183) );
  NANDN U187 ( .A(n184), .B(A[253]), .Z(n181) );
  XOR U188 ( .A(n184), .B(n185), .Z(DIFF[253]) );
  XOR U189 ( .A(B[253]), .B(A[253]), .Z(n185) );
  AND U190 ( .A(n186), .B(n187), .Z(n184) );
  NANDN U191 ( .A(B[252]), .B(n188), .Z(n187) );
  NANDN U192 ( .A(A[252]), .B(n189), .Z(n188) );
  NANDN U193 ( .A(n189), .B(A[252]), .Z(n186) );
  XOR U194 ( .A(n189), .B(n190), .Z(DIFF[252]) );
  XOR U195 ( .A(B[252]), .B(A[252]), .Z(n190) );
  AND U196 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U197 ( .A(B[251]), .B(n193), .Z(n192) );
  NANDN U198 ( .A(A[251]), .B(n194), .Z(n193) );
  NANDN U199 ( .A(n194), .B(A[251]), .Z(n191) );
  XOR U200 ( .A(n194), .B(n195), .Z(DIFF[251]) );
  XOR U201 ( .A(B[251]), .B(A[251]), .Z(n195) );
  AND U202 ( .A(n196), .B(n197), .Z(n194) );
  NANDN U203 ( .A(B[250]), .B(n198), .Z(n197) );
  NANDN U204 ( .A(A[250]), .B(n199), .Z(n198) );
  NANDN U205 ( .A(n199), .B(A[250]), .Z(n196) );
  XOR U206 ( .A(n199), .B(n200), .Z(DIFF[250]) );
  XOR U207 ( .A(B[250]), .B(A[250]), .Z(n200) );
  AND U208 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U209 ( .A(B[249]), .B(n203), .Z(n202) );
  NANDN U210 ( .A(A[249]), .B(n204), .Z(n203) );
  NANDN U211 ( .A(n204), .B(A[249]), .Z(n201) );
  XOR U212 ( .A(n205), .B(n206), .Z(DIFF[24]) );
  XOR U213 ( .A(B[24]), .B(A[24]), .Z(n206) );
  XOR U214 ( .A(n204), .B(n207), .Z(DIFF[249]) );
  XOR U215 ( .A(B[249]), .B(A[249]), .Z(n207) );
  AND U216 ( .A(n208), .B(n209), .Z(n204) );
  NANDN U217 ( .A(B[248]), .B(n210), .Z(n209) );
  NANDN U218 ( .A(A[248]), .B(n211), .Z(n210) );
  NANDN U219 ( .A(n211), .B(A[248]), .Z(n208) );
  XOR U220 ( .A(n211), .B(n212), .Z(DIFF[248]) );
  XOR U221 ( .A(B[248]), .B(A[248]), .Z(n212) );
  AND U222 ( .A(n213), .B(n214), .Z(n211) );
  NANDN U223 ( .A(B[247]), .B(n215), .Z(n214) );
  NANDN U224 ( .A(A[247]), .B(n216), .Z(n215) );
  NANDN U225 ( .A(n216), .B(A[247]), .Z(n213) );
  XOR U226 ( .A(n216), .B(n217), .Z(DIFF[247]) );
  XOR U227 ( .A(B[247]), .B(A[247]), .Z(n217) );
  AND U228 ( .A(n218), .B(n219), .Z(n216) );
  NANDN U229 ( .A(B[246]), .B(n220), .Z(n219) );
  NANDN U230 ( .A(A[246]), .B(n221), .Z(n220) );
  NANDN U231 ( .A(n221), .B(A[246]), .Z(n218) );
  XOR U232 ( .A(n221), .B(n222), .Z(DIFF[246]) );
  XOR U233 ( .A(B[246]), .B(A[246]), .Z(n222) );
  AND U234 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U235 ( .A(B[245]), .B(n225), .Z(n224) );
  NANDN U236 ( .A(A[245]), .B(n226), .Z(n225) );
  NANDN U237 ( .A(n226), .B(A[245]), .Z(n223) );
  XOR U238 ( .A(n226), .B(n227), .Z(DIFF[245]) );
  XOR U239 ( .A(B[245]), .B(A[245]), .Z(n227) );
  AND U240 ( .A(n228), .B(n229), .Z(n226) );
  NANDN U241 ( .A(B[244]), .B(n230), .Z(n229) );
  NANDN U242 ( .A(A[244]), .B(n231), .Z(n230) );
  NANDN U243 ( .A(n231), .B(A[244]), .Z(n228) );
  XOR U244 ( .A(n231), .B(n232), .Z(DIFF[244]) );
  XOR U245 ( .A(B[244]), .B(A[244]), .Z(n232) );
  AND U246 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U247 ( .A(B[243]), .B(n235), .Z(n234) );
  NANDN U248 ( .A(A[243]), .B(n236), .Z(n235) );
  NANDN U249 ( .A(n236), .B(A[243]), .Z(n233) );
  XOR U250 ( .A(n236), .B(n237), .Z(DIFF[243]) );
  XOR U251 ( .A(B[243]), .B(A[243]), .Z(n237) );
  AND U252 ( .A(n238), .B(n239), .Z(n236) );
  NANDN U253 ( .A(B[242]), .B(n240), .Z(n239) );
  NANDN U254 ( .A(A[242]), .B(n241), .Z(n240) );
  NANDN U255 ( .A(n241), .B(A[242]), .Z(n238) );
  XOR U256 ( .A(n241), .B(n242), .Z(DIFF[242]) );
  XOR U257 ( .A(B[242]), .B(A[242]), .Z(n242) );
  AND U258 ( .A(n243), .B(n244), .Z(n241) );
  NANDN U259 ( .A(B[241]), .B(n245), .Z(n244) );
  NANDN U260 ( .A(A[241]), .B(n246), .Z(n245) );
  NANDN U261 ( .A(n246), .B(A[241]), .Z(n243) );
  XOR U262 ( .A(n246), .B(n247), .Z(DIFF[241]) );
  XOR U263 ( .A(B[241]), .B(A[241]), .Z(n247) );
  AND U264 ( .A(n248), .B(n249), .Z(n246) );
  NANDN U265 ( .A(B[240]), .B(n250), .Z(n249) );
  NANDN U266 ( .A(A[240]), .B(n251), .Z(n250) );
  NANDN U267 ( .A(n251), .B(A[240]), .Z(n248) );
  XOR U268 ( .A(n251), .B(n252), .Z(DIFF[240]) );
  XOR U269 ( .A(B[240]), .B(A[240]), .Z(n252) );
  AND U270 ( .A(n253), .B(n254), .Z(n251) );
  NANDN U271 ( .A(B[239]), .B(n255), .Z(n254) );
  NANDN U272 ( .A(A[239]), .B(n256), .Z(n255) );
  NANDN U273 ( .A(n256), .B(A[239]), .Z(n253) );
  XOR U274 ( .A(n257), .B(n258), .Z(DIFF[23]) );
  XOR U275 ( .A(B[23]), .B(A[23]), .Z(n258) );
  XOR U276 ( .A(n256), .B(n259), .Z(DIFF[239]) );
  XOR U277 ( .A(B[239]), .B(A[239]), .Z(n259) );
  AND U278 ( .A(n260), .B(n261), .Z(n256) );
  NANDN U279 ( .A(B[238]), .B(n262), .Z(n261) );
  NANDN U280 ( .A(A[238]), .B(n263), .Z(n262) );
  NANDN U281 ( .A(n263), .B(A[238]), .Z(n260) );
  XOR U282 ( .A(n263), .B(n264), .Z(DIFF[238]) );
  XOR U283 ( .A(B[238]), .B(A[238]), .Z(n264) );
  AND U284 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U285 ( .A(B[237]), .B(n267), .Z(n266) );
  NANDN U286 ( .A(A[237]), .B(n268), .Z(n267) );
  NANDN U287 ( .A(n268), .B(A[237]), .Z(n265) );
  XOR U288 ( .A(n268), .B(n269), .Z(DIFF[237]) );
  XOR U289 ( .A(B[237]), .B(A[237]), .Z(n269) );
  AND U290 ( .A(n270), .B(n271), .Z(n268) );
  NANDN U291 ( .A(B[236]), .B(n272), .Z(n271) );
  NANDN U292 ( .A(A[236]), .B(n273), .Z(n272) );
  NANDN U293 ( .A(n273), .B(A[236]), .Z(n270) );
  XOR U294 ( .A(n273), .B(n274), .Z(DIFF[236]) );
  XOR U295 ( .A(B[236]), .B(A[236]), .Z(n274) );
  AND U296 ( .A(n275), .B(n276), .Z(n273) );
  NANDN U297 ( .A(B[235]), .B(n277), .Z(n276) );
  NANDN U298 ( .A(A[235]), .B(n278), .Z(n277) );
  NANDN U299 ( .A(n278), .B(A[235]), .Z(n275) );
  XOR U300 ( .A(n278), .B(n279), .Z(DIFF[235]) );
  XOR U301 ( .A(B[235]), .B(A[235]), .Z(n279) );
  AND U302 ( .A(n280), .B(n281), .Z(n278) );
  NANDN U303 ( .A(B[234]), .B(n282), .Z(n281) );
  NANDN U304 ( .A(A[234]), .B(n283), .Z(n282) );
  NANDN U305 ( .A(n283), .B(A[234]), .Z(n280) );
  XOR U306 ( .A(n283), .B(n284), .Z(DIFF[234]) );
  XOR U307 ( .A(B[234]), .B(A[234]), .Z(n284) );
  AND U308 ( .A(n285), .B(n286), .Z(n283) );
  NANDN U309 ( .A(B[233]), .B(n287), .Z(n286) );
  NANDN U310 ( .A(A[233]), .B(n288), .Z(n287) );
  NANDN U311 ( .A(n288), .B(A[233]), .Z(n285) );
  XOR U312 ( .A(n288), .B(n289), .Z(DIFF[233]) );
  XOR U313 ( .A(B[233]), .B(A[233]), .Z(n289) );
  AND U314 ( .A(n290), .B(n291), .Z(n288) );
  NANDN U315 ( .A(B[232]), .B(n292), .Z(n291) );
  NANDN U316 ( .A(A[232]), .B(n293), .Z(n292) );
  NANDN U317 ( .A(n293), .B(A[232]), .Z(n290) );
  XOR U318 ( .A(n293), .B(n294), .Z(DIFF[232]) );
  XOR U319 ( .A(B[232]), .B(A[232]), .Z(n294) );
  AND U320 ( .A(n295), .B(n296), .Z(n293) );
  NANDN U321 ( .A(B[231]), .B(n297), .Z(n296) );
  NANDN U322 ( .A(A[231]), .B(n298), .Z(n297) );
  NANDN U323 ( .A(n298), .B(A[231]), .Z(n295) );
  XOR U324 ( .A(n298), .B(n299), .Z(DIFF[231]) );
  XOR U325 ( .A(B[231]), .B(A[231]), .Z(n299) );
  AND U326 ( .A(n300), .B(n301), .Z(n298) );
  NANDN U327 ( .A(B[230]), .B(n302), .Z(n301) );
  NANDN U328 ( .A(A[230]), .B(n303), .Z(n302) );
  NANDN U329 ( .A(n303), .B(A[230]), .Z(n300) );
  XOR U330 ( .A(n303), .B(n304), .Z(DIFF[230]) );
  XOR U331 ( .A(B[230]), .B(A[230]), .Z(n304) );
  AND U332 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U333 ( .A(B[229]), .B(n307), .Z(n306) );
  NANDN U334 ( .A(A[229]), .B(n308), .Z(n307) );
  NANDN U335 ( .A(n308), .B(A[229]), .Z(n305) );
  XOR U336 ( .A(n309), .B(n310), .Z(DIFF[22]) );
  XOR U337 ( .A(B[22]), .B(A[22]), .Z(n310) );
  XOR U338 ( .A(n308), .B(n311), .Z(DIFF[229]) );
  XOR U339 ( .A(B[229]), .B(A[229]), .Z(n311) );
  AND U340 ( .A(n312), .B(n313), .Z(n308) );
  NANDN U341 ( .A(B[228]), .B(n314), .Z(n313) );
  NANDN U342 ( .A(A[228]), .B(n315), .Z(n314) );
  NANDN U343 ( .A(n315), .B(A[228]), .Z(n312) );
  XOR U344 ( .A(n315), .B(n316), .Z(DIFF[228]) );
  XOR U345 ( .A(B[228]), .B(A[228]), .Z(n316) );
  AND U346 ( .A(n317), .B(n318), .Z(n315) );
  NANDN U347 ( .A(B[227]), .B(n319), .Z(n318) );
  NANDN U348 ( .A(A[227]), .B(n320), .Z(n319) );
  NANDN U349 ( .A(n320), .B(A[227]), .Z(n317) );
  XOR U350 ( .A(n320), .B(n321), .Z(DIFF[227]) );
  XOR U351 ( .A(B[227]), .B(A[227]), .Z(n321) );
  AND U352 ( .A(n322), .B(n323), .Z(n320) );
  NANDN U353 ( .A(B[226]), .B(n324), .Z(n323) );
  NANDN U354 ( .A(A[226]), .B(n325), .Z(n324) );
  NANDN U355 ( .A(n325), .B(A[226]), .Z(n322) );
  XOR U356 ( .A(n325), .B(n326), .Z(DIFF[226]) );
  XOR U357 ( .A(B[226]), .B(A[226]), .Z(n326) );
  AND U358 ( .A(n327), .B(n328), .Z(n325) );
  NANDN U359 ( .A(B[225]), .B(n329), .Z(n328) );
  NANDN U360 ( .A(A[225]), .B(n330), .Z(n329) );
  NANDN U361 ( .A(n330), .B(A[225]), .Z(n327) );
  XOR U362 ( .A(n330), .B(n331), .Z(DIFF[225]) );
  XOR U363 ( .A(B[225]), .B(A[225]), .Z(n331) );
  AND U364 ( .A(n332), .B(n333), .Z(n330) );
  NANDN U365 ( .A(B[224]), .B(n334), .Z(n333) );
  NANDN U366 ( .A(A[224]), .B(n335), .Z(n334) );
  NANDN U367 ( .A(n335), .B(A[224]), .Z(n332) );
  XOR U368 ( .A(n335), .B(n336), .Z(DIFF[224]) );
  XOR U369 ( .A(B[224]), .B(A[224]), .Z(n336) );
  AND U370 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U371 ( .A(B[223]), .B(n339), .Z(n338) );
  NANDN U372 ( .A(A[223]), .B(n340), .Z(n339) );
  NANDN U373 ( .A(n340), .B(A[223]), .Z(n337) );
  XOR U374 ( .A(n340), .B(n341), .Z(DIFF[223]) );
  XOR U375 ( .A(B[223]), .B(A[223]), .Z(n341) );
  AND U376 ( .A(n342), .B(n343), .Z(n340) );
  NANDN U377 ( .A(B[222]), .B(n344), .Z(n343) );
  NANDN U378 ( .A(A[222]), .B(n345), .Z(n344) );
  NANDN U379 ( .A(n345), .B(A[222]), .Z(n342) );
  XOR U380 ( .A(n345), .B(n346), .Z(DIFF[222]) );
  XOR U381 ( .A(B[222]), .B(A[222]), .Z(n346) );
  AND U382 ( .A(n347), .B(n348), .Z(n345) );
  NANDN U383 ( .A(B[221]), .B(n349), .Z(n348) );
  NANDN U384 ( .A(A[221]), .B(n350), .Z(n349) );
  NANDN U385 ( .A(n350), .B(A[221]), .Z(n347) );
  XOR U386 ( .A(n350), .B(n351), .Z(DIFF[221]) );
  XOR U387 ( .A(B[221]), .B(A[221]), .Z(n351) );
  AND U388 ( .A(n352), .B(n353), .Z(n350) );
  NANDN U389 ( .A(B[220]), .B(n354), .Z(n353) );
  NANDN U390 ( .A(A[220]), .B(n355), .Z(n354) );
  NANDN U391 ( .A(n355), .B(A[220]), .Z(n352) );
  XOR U392 ( .A(n355), .B(n356), .Z(DIFF[220]) );
  XOR U393 ( .A(B[220]), .B(A[220]), .Z(n356) );
  AND U394 ( .A(n357), .B(n358), .Z(n355) );
  NANDN U395 ( .A(B[219]), .B(n359), .Z(n358) );
  NANDN U396 ( .A(A[219]), .B(n360), .Z(n359) );
  NANDN U397 ( .A(n360), .B(A[219]), .Z(n357) );
  XOR U398 ( .A(n361), .B(n362), .Z(DIFF[21]) );
  XOR U399 ( .A(B[21]), .B(A[21]), .Z(n362) );
  XOR U400 ( .A(n360), .B(n363), .Z(DIFF[219]) );
  XOR U401 ( .A(B[219]), .B(A[219]), .Z(n363) );
  AND U402 ( .A(n364), .B(n365), .Z(n360) );
  NANDN U403 ( .A(B[218]), .B(n366), .Z(n365) );
  NANDN U404 ( .A(A[218]), .B(n367), .Z(n366) );
  NANDN U405 ( .A(n367), .B(A[218]), .Z(n364) );
  XOR U406 ( .A(n367), .B(n368), .Z(DIFF[218]) );
  XOR U407 ( .A(B[218]), .B(A[218]), .Z(n368) );
  AND U408 ( .A(n369), .B(n370), .Z(n367) );
  NANDN U409 ( .A(B[217]), .B(n371), .Z(n370) );
  NANDN U410 ( .A(A[217]), .B(n372), .Z(n371) );
  NANDN U411 ( .A(n372), .B(A[217]), .Z(n369) );
  XOR U412 ( .A(n372), .B(n373), .Z(DIFF[217]) );
  XOR U413 ( .A(B[217]), .B(A[217]), .Z(n373) );
  AND U414 ( .A(n374), .B(n375), .Z(n372) );
  NANDN U415 ( .A(B[216]), .B(n376), .Z(n375) );
  NANDN U416 ( .A(A[216]), .B(n377), .Z(n376) );
  NANDN U417 ( .A(n377), .B(A[216]), .Z(n374) );
  XOR U418 ( .A(n377), .B(n378), .Z(DIFF[216]) );
  XOR U419 ( .A(B[216]), .B(A[216]), .Z(n378) );
  AND U420 ( .A(n379), .B(n380), .Z(n377) );
  NANDN U421 ( .A(B[215]), .B(n381), .Z(n380) );
  NANDN U422 ( .A(A[215]), .B(n382), .Z(n381) );
  NANDN U423 ( .A(n382), .B(A[215]), .Z(n379) );
  XOR U424 ( .A(n382), .B(n383), .Z(DIFF[215]) );
  XOR U425 ( .A(B[215]), .B(A[215]), .Z(n383) );
  AND U426 ( .A(n384), .B(n385), .Z(n382) );
  NANDN U427 ( .A(B[214]), .B(n386), .Z(n385) );
  NANDN U428 ( .A(A[214]), .B(n387), .Z(n386) );
  NANDN U429 ( .A(n387), .B(A[214]), .Z(n384) );
  XOR U430 ( .A(n387), .B(n388), .Z(DIFF[214]) );
  XOR U431 ( .A(B[214]), .B(A[214]), .Z(n388) );
  AND U432 ( .A(n389), .B(n390), .Z(n387) );
  NANDN U433 ( .A(B[213]), .B(n391), .Z(n390) );
  NANDN U434 ( .A(A[213]), .B(n392), .Z(n391) );
  NANDN U435 ( .A(n392), .B(A[213]), .Z(n389) );
  XOR U436 ( .A(n392), .B(n393), .Z(DIFF[213]) );
  XOR U437 ( .A(B[213]), .B(A[213]), .Z(n393) );
  AND U438 ( .A(n394), .B(n395), .Z(n392) );
  NANDN U439 ( .A(B[212]), .B(n396), .Z(n395) );
  NANDN U440 ( .A(A[212]), .B(n397), .Z(n396) );
  NANDN U441 ( .A(n397), .B(A[212]), .Z(n394) );
  XOR U442 ( .A(n397), .B(n398), .Z(DIFF[212]) );
  XOR U443 ( .A(B[212]), .B(A[212]), .Z(n398) );
  AND U444 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U445 ( .A(B[211]), .B(n401), .Z(n400) );
  NANDN U446 ( .A(A[211]), .B(n402), .Z(n401) );
  NANDN U447 ( .A(n402), .B(A[211]), .Z(n399) );
  XOR U448 ( .A(n402), .B(n403), .Z(DIFF[211]) );
  XOR U449 ( .A(B[211]), .B(A[211]), .Z(n403) );
  AND U450 ( .A(n404), .B(n405), .Z(n402) );
  NANDN U451 ( .A(B[210]), .B(n406), .Z(n405) );
  NANDN U452 ( .A(A[210]), .B(n407), .Z(n406) );
  NANDN U453 ( .A(n407), .B(A[210]), .Z(n404) );
  XOR U454 ( .A(n407), .B(n408), .Z(DIFF[210]) );
  XOR U455 ( .A(B[210]), .B(A[210]), .Z(n408) );
  AND U456 ( .A(n409), .B(n410), .Z(n407) );
  NANDN U457 ( .A(B[209]), .B(n411), .Z(n410) );
  NANDN U458 ( .A(A[209]), .B(n412), .Z(n411) );
  NANDN U459 ( .A(n412), .B(A[209]), .Z(n409) );
  XOR U460 ( .A(n413), .B(n414), .Z(DIFF[20]) );
  XOR U461 ( .A(B[20]), .B(A[20]), .Z(n414) );
  XOR U462 ( .A(n412), .B(n415), .Z(DIFF[209]) );
  XOR U463 ( .A(B[209]), .B(A[209]), .Z(n415) );
  AND U464 ( .A(n416), .B(n417), .Z(n412) );
  NANDN U465 ( .A(B[208]), .B(n418), .Z(n417) );
  NANDN U466 ( .A(A[208]), .B(n419), .Z(n418) );
  NANDN U467 ( .A(n419), .B(A[208]), .Z(n416) );
  XOR U468 ( .A(n419), .B(n420), .Z(DIFF[208]) );
  XOR U469 ( .A(B[208]), .B(A[208]), .Z(n420) );
  AND U470 ( .A(n421), .B(n422), .Z(n419) );
  NANDN U471 ( .A(B[207]), .B(n423), .Z(n422) );
  NANDN U472 ( .A(A[207]), .B(n424), .Z(n423) );
  NANDN U473 ( .A(n424), .B(A[207]), .Z(n421) );
  XOR U474 ( .A(n424), .B(n425), .Z(DIFF[207]) );
  XOR U475 ( .A(B[207]), .B(A[207]), .Z(n425) );
  AND U476 ( .A(n426), .B(n427), .Z(n424) );
  NANDN U477 ( .A(B[206]), .B(n428), .Z(n427) );
  NANDN U478 ( .A(A[206]), .B(n429), .Z(n428) );
  NANDN U479 ( .A(n429), .B(A[206]), .Z(n426) );
  XOR U480 ( .A(n429), .B(n430), .Z(DIFF[206]) );
  XOR U481 ( .A(B[206]), .B(A[206]), .Z(n430) );
  AND U482 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U483 ( .A(B[205]), .B(n433), .Z(n432) );
  NANDN U484 ( .A(A[205]), .B(n434), .Z(n433) );
  NANDN U485 ( .A(n434), .B(A[205]), .Z(n431) );
  XOR U486 ( .A(n434), .B(n435), .Z(DIFF[205]) );
  XOR U487 ( .A(B[205]), .B(A[205]), .Z(n435) );
  AND U488 ( .A(n436), .B(n437), .Z(n434) );
  NANDN U489 ( .A(B[204]), .B(n438), .Z(n437) );
  NANDN U490 ( .A(A[204]), .B(n439), .Z(n438) );
  NANDN U491 ( .A(n439), .B(A[204]), .Z(n436) );
  XOR U492 ( .A(n439), .B(n440), .Z(DIFF[204]) );
  XOR U493 ( .A(B[204]), .B(A[204]), .Z(n440) );
  AND U494 ( .A(n441), .B(n442), .Z(n439) );
  NANDN U495 ( .A(B[203]), .B(n443), .Z(n442) );
  NANDN U496 ( .A(A[203]), .B(n444), .Z(n443) );
  NANDN U497 ( .A(n444), .B(A[203]), .Z(n441) );
  XOR U498 ( .A(n444), .B(n445), .Z(DIFF[203]) );
  XOR U499 ( .A(B[203]), .B(A[203]), .Z(n445) );
  AND U500 ( .A(n446), .B(n447), .Z(n444) );
  NANDN U501 ( .A(B[202]), .B(n448), .Z(n447) );
  NANDN U502 ( .A(A[202]), .B(n449), .Z(n448) );
  NANDN U503 ( .A(n449), .B(A[202]), .Z(n446) );
  XOR U504 ( .A(n449), .B(n450), .Z(DIFF[202]) );
  XOR U505 ( .A(B[202]), .B(A[202]), .Z(n450) );
  AND U506 ( .A(n451), .B(n452), .Z(n449) );
  NANDN U507 ( .A(B[201]), .B(n453), .Z(n452) );
  NANDN U508 ( .A(A[201]), .B(n454), .Z(n453) );
  NANDN U509 ( .A(n454), .B(A[201]), .Z(n451) );
  XOR U510 ( .A(n454), .B(n455), .Z(DIFF[201]) );
  XOR U511 ( .A(B[201]), .B(A[201]), .Z(n455) );
  AND U512 ( .A(n456), .B(n457), .Z(n454) );
  NANDN U513 ( .A(B[200]), .B(n458), .Z(n457) );
  NANDN U514 ( .A(A[200]), .B(n459), .Z(n458) );
  NANDN U515 ( .A(n459), .B(A[200]), .Z(n456) );
  XOR U516 ( .A(n459), .B(n460), .Z(DIFF[200]) );
  XOR U517 ( .A(B[200]), .B(A[200]), .Z(n460) );
  AND U518 ( .A(n461), .B(n462), .Z(n459) );
  NANDN U519 ( .A(B[199]), .B(n463), .Z(n462) );
  NANDN U520 ( .A(A[199]), .B(n464), .Z(n463) );
  NANDN U521 ( .A(n464), .B(A[199]), .Z(n461) );
  XOR U522 ( .A(n2), .B(n465), .Z(DIFF[1]) );
  XOR U523 ( .A(B[1]), .B(A[1]), .Z(n465) );
  XOR U524 ( .A(n466), .B(n467), .Z(DIFF[19]) );
  XOR U525 ( .A(B[19]), .B(A[19]), .Z(n467) );
  XOR U526 ( .A(n464), .B(n468), .Z(DIFF[199]) );
  XOR U527 ( .A(B[199]), .B(A[199]), .Z(n468) );
  AND U528 ( .A(n469), .B(n470), .Z(n464) );
  NANDN U529 ( .A(B[198]), .B(n471), .Z(n470) );
  NANDN U530 ( .A(A[198]), .B(n472), .Z(n471) );
  NANDN U531 ( .A(n472), .B(A[198]), .Z(n469) );
  XOR U532 ( .A(n472), .B(n473), .Z(DIFF[198]) );
  XOR U533 ( .A(B[198]), .B(A[198]), .Z(n473) );
  AND U534 ( .A(n474), .B(n475), .Z(n472) );
  NANDN U535 ( .A(B[197]), .B(n476), .Z(n475) );
  NANDN U536 ( .A(A[197]), .B(n477), .Z(n476) );
  NANDN U537 ( .A(n477), .B(A[197]), .Z(n474) );
  XOR U538 ( .A(n477), .B(n478), .Z(DIFF[197]) );
  XOR U539 ( .A(B[197]), .B(A[197]), .Z(n478) );
  AND U540 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U541 ( .A(B[196]), .B(n481), .Z(n480) );
  NANDN U542 ( .A(A[196]), .B(n482), .Z(n481) );
  NANDN U543 ( .A(n482), .B(A[196]), .Z(n479) );
  XOR U544 ( .A(n482), .B(n483), .Z(DIFF[196]) );
  XOR U545 ( .A(B[196]), .B(A[196]), .Z(n483) );
  AND U546 ( .A(n484), .B(n485), .Z(n482) );
  NANDN U547 ( .A(B[195]), .B(n486), .Z(n485) );
  NANDN U548 ( .A(A[195]), .B(n487), .Z(n486) );
  NANDN U549 ( .A(n487), .B(A[195]), .Z(n484) );
  XOR U550 ( .A(n487), .B(n488), .Z(DIFF[195]) );
  XOR U551 ( .A(B[195]), .B(A[195]), .Z(n488) );
  AND U552 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U553 ( .A(B[194]), .B(n491), .Z(n490) );
  NANDN U554 ( .A(A[194]), .B(n492), .Z(n491) );
  NANDN U555 ( .A(n492), .B(A[194]), .Z(n489) );
  XOR U556 ( .A(n492), .B(n493), .Z(DIFF[194]) );
  XOR U557 ( .A(B[194]), .B(A[194]), .Z(n493) );
  AND U558 ( .A(n494), .B(n495), .Z(n492) );
  NANDN U559 ( .A(B[193]), .B(n496), .Z(n495) );
  NANDN U560 ( .A(A[193]), .B(n497), .Z(n496) );
  NANDN U561 ( .A(n497), .B(A[193]), .Z(n494) );
  XOR U562 ( .A(n497), .B(n498), .Z(DIFF[193]) );
  XOR U563 ( .A(B[193]), .B(A[193]), .Z(n498) );
  AND U564 ( .A(n499), .B(n500), .Z(n497) );
  NANDN U565 ( .A(B[192]), .B(n501), .Z(n500) );
  NANDN U566 ( .A(A[192]), .B(n502), .Z(n501) );
  NANDN U567 ( .A(n502), .B(A[192]), .Z(n499) );
  XOR U568 ( .A(n502), .B(n503), .Z(DIFF[192]) );
  XOR U569 ( .A(B[192]), .B(A[192]), .Z(n503) );
  AND U570 ( .A(n504), .B(n505), .Z(n502) );
  NANDN U571 ( .A(B[191]), .B(n506), .Z(n505) );
  NANDN U572 ( .A(A[191]), .B(n507), .Z(n506) );
  NANDN U573 ( .A(n507), .B(A[191]), .Z(n504) );
  XOR U574 ( .A(n507), .B(n508), .Z(DIFF[191]) );
  XOR U575 ( .A(B[191]), .B(A[191]), .Z(n508) );
  AND U576 ( .A(n509), .B(n510), .Z(n507) );
  NANDN U577 ( .A(B[190]), .B(n511), .Z(n510) );
  NANDN U578 ( .A(A[190]), .B(n512), .Z(n511) );
  NANDN U579 ( .A(n512), .B(A[190]), .Z(n509) );
  XOR U580 ( .A(n512), .B(n513), .Z(DIFF[190]) );
  XOR U581 ( .A(B[190]), .B(A[190]), .Z(n513) );
  AND U582 ( .A(n514), .B(n515), .Z(n512) );
  NANDN U583 ( .A(B[189]), .B(n516), .Z(n515) );
  NANDN U584 ( .A(A[189]), .B(n517), .Z(n516) );
  NANDN U585 ( .A(n517), .B(A[189]), .Z(n514) );
  XOR U586 ( .A(n518), .B(n519), .Z(DIFF[18]) );
  XOR U587 ( .A(B[18]), .B(A[18]), .Z(n519) );
  XOR U588 ( .A(n517), .B(n520), .Z(DIFF[189]) );
  XOR U589 ( .A(B[189]), .B(A[189]), .Z(n520) );
  AND U590 ( .A(n521), .B(n522), .Z(n517) );
  NANDN U591 ( .A(B[188]), .B(n523), .Z(n522) );
  NANDN U592 ( .A(A[188]), .B(n524), .Z(n523) );
  NANDN U593 ( .A(n524), .B(A[188]), .Z(n521) );
  XOR U594 ( .A(n524), .B(n525), .Z(DIFF[188]) );
  XOR U595 ( .A(B[188]), .B(A[188]), .Z(n525) );
  AND U596 ( .A(n526), .B(n527), .Z(n524) );
  NANDN U597 ( .A(B[187]), .B(n528), .Z(n527) );
  NANDN U598 ( .A(A[187]), .B(n529), .Z(n528) );
  NANDN U599 ( .A(n529), .B(A[187]), .Z(n526) );
  XOR U600 ( .A(n529), .B(n530), .Z(DIFF[187]) );
  XOR U601 ( .A(B[187]), .B(A[187]), .Z(n530) );
  AND U602 ( .A(n531), .B(n532), .Z(n529) );
  NANDN U603 ( .A(B[186]), .B(n533), .Z(n532) );
  NANDN U604 ( .A(A[186]), .B(n534), .Z(n533) );
  NANDN U605 ( .A(n534), .B(A[186]), .Z(n531) );
  XOR U606 ( .A(n534), .B(n535), .Z(DIFF[186]) );
  XOR U607 ( .A(B[186]), .B(A[186]), .Z(n535) );
  AND U608 ( .A(n536), .B(n537), .Z(n534) );
  NANDN U609 ( .A(B[185]), .B(n538), .Z(n537) );
  NANDN U610 ( .A(A[185]), .B(n539), .Z(n538) );
  NANDN U611 ( .A(n539), .B(A[185]), .Z(n536) );
  XOR U612 ( .A(n539), .B(n540), .Z(DIFF[185]) );
  XOR U613 ( .A(B[185]), .B(A[185]), .Z(n540) );
  AND U614 ( .A(n541), .B(n542), .Z(n539) );
  NANDN U615 ( .A(B[184]), .B(n543), .Z(n542) );
  NANDN U616 ( .A(A[184]), .B(n544), .Z(n543) );
  NANDN U617 ( .A(n544), .B(A[184]), .Z(n541) );
  XOR U618 ( .A(n544), .B(n545), .Z(DIFF[184]) );
  XOR U619 ( .A(B[184]), .B(A[184]), .Z(n545) );
  AND U620 ( .A(n546), .B(n547), .Z(n544) );
  NANDN U621 ( .A(B[183]), .B(n548), .Z(n547) );
  NANDN U622 ( .A(A[183]), .B(n549), .Z(n548) );
  NANDN U623 ( .A(n549), .B(A[183]), .Z(n546) );
  XOR U624 ( .A(n549), .B(n550), .Z(DIFF[183]) );
  XOR U625 ( .A(B[183]), .B(A[183]), .Z(n550) );
  AND U626 ( .A(n551), .B(n552), .Z(n549) );
  NANDN U627 ( .A(B[182]), .B(n553), .Z(n552) );
  NANDN U628 ( .A(A[182]), .B(n554), .Z(n553) );
  NANDN U629 ( .A(n554), .B(A[182]), .Z(n551) );
  XOR U630 ( .A(n554), .B(n555), .Z(DIFF[182]) );
  XOR U631 ( .A(B[182]), .B(A[182]), .Z(n555) );
  AND U632 ( .A(n556), .B(n557), .Z(n554) );
  NANDN U633 ( .A(B[181]), .B(n558), .Z(n557) );
  NANDN U634 ( .A(A[181]), .B(n559), .Z(n558) );
  NANDN U635 ( .A(n559), .B(A[181]), .Z(n556) );
  XOR U636 ( .A(n559), .B(n560), .Z(DIFF[181]) );
  XOR U637 ( .A(B[181]), .B(A[181]), .Z(n560) );
  AND U638 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U639 ( .A(B[180]), .B(n563), .Z(n562) );
  NANDN U640 ( .A(A[180]), .B(n564), .Z(n563) );
  NANDN U641 ( .A(n564), .B(A[180]), .Z(n561) );
  XOR U642 ( .A(n564), .B(n565), .Z(DIFF[180]) );
  XOR U643 ( .A(B[180]), .B(A[180]), .Z(n565) );
  AND U644 ( .A(n566), .B(n567), .Z(n564) );
  NANDN U645 ( .A(B[179]), .B(n568), .Z(n567) );
  NANDN U646 ( .A(A[179]), .B(n569), .Z(n568) );
  NANDN U647 ( .A(n569), .B(A[179]), .Z(n566) );
  XOR U648 ( .A(n570), .B(n571), .Z(DIFF[17]) );
  XOR U649 ( .A(B[17]), .B(A[17]), .Z(n571) );
  XOR U650 ( .A(n569), .B(n572), .Z(DIFF[179]) );
  XOR U651 ( .A(B[179]), .B(A[179]), .Z(n572) );
  AND U652 ( .A(n573), .B(n574), .Z(n569) );
  NANDN U653 ( .A(B[178]), .B(n575), .Z(n574) );
  NANDN U654 ( .A(A[178]), .B(n576), .Z(n575) );
  NANDN U655 ( .A(n576), .B(A[178]), .Z(n573) );
  XOR U656 ( .A(n576), .B(n577), .Z(DIFF[178]) );
  XOR U657 ( .A(B[178]), .B(A[178]), .Z(n577) );
  AND U658 ( .A(n578), .B(n579), .Z(n576) );
  NANDN U659 ( .A(B[177]), .B(n580), .Z(n579) );
  NANDN U660 ( .A(A[177]), .B(n581), .Z(n580) );
  NANDN U661 ( .A(n581), .B(A[177]), .Z(n578) );
  XOR U662 ( .A(n581), .B(n582), .Z(DIFF[177]) );
  XOR U663 ( .A(B[177]), .B(A[177]), .Z(n582) );
  AND U664 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U665 ( .A(B[176]), .B(n585), .Z(n584) );
  NANDN U666 ( .A(A[176]), .B(n586), .Z(n585) );
  NANDN U667 ( .A(n586), .B(A[176]), .Z(n583) );
  XOR U668 ( .A(n586), .B(n587), .Z(DIFF[176]) );
  XOR U669 ( .A(B[176]), .B(A[176]), .Z(n587) );
  AND U670 ( .A(n588), .B(n589), .Z(n586) );
  NANDN U671 ( .A(B[175]), .B(n590), .Z(n589) );
  NANDN U672 ( .A(A[175]), .B(n591), .Z(n590) );
  NANDN U673 ( .A(n591), .B(A[175]), .Z(n588) );
  XOR U674 ( .A(n591), .B(n592), .Z(DIFF[175]) );
  XOR U675 ( .A(B[175]), .B(A[175]), .Z(n592) );
  AND U676 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U677 ( .A(B[174]), .B(n595), .Z(n594) );
  NANDN U678 ( .A(A[174]), .B(n596), .Z(n595) );
  NANDN U679 ( .A(n596), .B(A[174]), .Z(n593) );
  XOR U680 ( .A(n596), .B(n597), .Z(DIFF[174]) );
  XOR U681 ( .A(B[174]), .B(A[174]), .Z(n597) );
  AND U682 ( .A(n598), .B(n599), .Z(n596) );
  NANDN U683 ( .A(B[173]), .B(n600), .Z(n599) );
  NANDN U684 ( .A(A[173]), .B(n601), .Z(n600) );
  NANDN U685 ( .A(n601), .B(A[173]), .Z(n598) );
  XOR U686 ( .A(n601), .B(n602), .Z(DIFF[173]) );
  XOR U687 ( .A(B[173]), .B(A[173]), .Z(n602) );
  AND U688 ( .A(n603), .B(n604), .Z(n601) );
  NANDN U689 ( .A(B[172]), .B(n605), .Z(n604) );
  NANDN U690 ( .A(A[172]), .B(n606), .Z(n605) );
  NANDN U691 ( .A(n606), .B(A[172]), .Z(n603) );
  XOR U692 ( .A(n606), .B(n607), .Z(DIFF[172]) );
  XOR U693 ( .A(B[172]), .B(A[172]), .Z(n607) );
  AND U694 ( .A(n608), .B(n609), .Z(n606) );
  NANDN U695 ( .A(B[171]), .B(n610), .Z(n609) );
  NANDN U696 ( .A(A[171]), .B(n611), .Z(n610) );
  NANDN U697 ( .A(n611), .B(A[171]), .Z(n608) );
  XOR U698 ( .A(n611), .B(n612), .Z(DIFF[171]) );
  XOR U699 ( .A(B[171]), .B(A[171]), .Z(n612) );
  AND U700 ( .A(n613), .B(n614), .Z(n611) );
  NANDN U701 ( .A(B[170]), .B(n615), .Z(n614) );
  NANDN U702 ( .A(A[170]), .B(n616), .Z(n615) );
  NANDN U703 ( .A(n616), .B(A[170]), .Z(n613) );
  XOR U704 ( .A(n616), .B(n617), .Z(DIFF[170]) );
  XOR U705 ( .A(B[170]), .B(A[170]), .Z(n617) );
  AND U706 ( .A(n618), .B(n619), .Z(n616) );
  NANDN U707 ( .A(B[169]), .B(n620), .Z(n619) );
  NANDN U708 ( .A(A[169]), .B(n621), .Z(n620) );
  NANDN U709 ( .A(n621), .B(A[169]), .Z(n618) );
  XOR U710 ( .A(n622), .B(n623), .Z(DIFF[16]) );
  XOR U711 ( .A(B[16]), .B(A[16]), .Z(n623) );
  XOR U712 ( .A(n621), .B(n624), .Z(DIFF[169]) );
  XOR U713 ( .A(B[169]), .B(A[169]), .Z(n624) );
  AND U714 ( .A(n625), .B(n626), .Z(n621) );
  NANDN U715 ( .A(B[168]), .B(n627), .Z(n626) );
  NANDN U716 ( .A(A[168]), .B(n628), .Z(n627) );
  NANDN U717 ( .A(n628), .B(A[168]), .Z(n625) );
  XOR U718 ( .A(n628), .B(n629), .Z(DIFF[168]) );
  XOR U719 ( .A(B[168]), .B(A[168]), .Z(n629) );
  AND U720 ( .A(n630), .B(n631), .Z(n628) );
  NANDN U721 ( .A(B[167]), .B(n632), .Z(n631) );
  NANDN U722 ( .A(A[167]), .B(n633), .Z(n632) );
  NANDN U723 ( .A(n633), .B(A[167]), .Z(n630) );
  XOR U724 ( .A(n633), .B(n634), .Z(DIFF[167]) );
  XOR U725 ( .A(B[167]), .B(A[167]), .Z(n634) );
  AND U726 ( .A(n635), .B(n636), .Z(n633) );
  NANDN U727 ( .A(B[166]), .B(n637), .Z(n636) );
  NANDN U728 ( .A(A[166]), .B(n638), .Z(n637) );
  NANDN U729 ( .A(n638), .B(A[166]), .Z(n635) );
  XOR U730 ( .A(n638), .B(n639), .Z(DIFF[166]) );
  XOR U731 ( .A(B[166]), .B(A[166]), .Z(n639) );
  AND U732 ( .A(n640), .B(n641), .Z(n638) );
  NANDN U733 ( .A(B[165]), .B(n642), .Z(n641) );
  NANDN U734 ( .A(A[165]), .B(n643), .Z(n642) );
  NANDN U735 ( .A(n643), .B(A[165]), .Z(n640) );
  XOR U736 ( .A(n643), .B(n644), .Z(DIFF[165]) );
  XOR U737 ( .A(B[165]), .B(A[165]), .Z(n644) );
  AND U738 ( .A(n645), .B(n646), .Z(n643) );
  NANDN U739 ( .A(B[164]), .B(n647), .Z(n646) );
  NANDN U740 ( .A(A[164]), .B(n648), .Z(n647) );
  NANDN U741 ( .A(n648), .B(A[164]), .Z(n645) );
  XOR U742 ( .A(n648), .B(n649), .Z(DIFF[164]) );
  XOR U743 ( .A(B[164]), .B(A[164]), .Z(n649) );
  AND U744 ( .A(n650), .B(n651), .Z(n648) );
  NANDN U745 ( .A(B[163]), .B(n652), .Z(n651) );
  NANDN U746 ( .A(A[163]), .B(n653), .Z(n652) );
  NANDN U747 ( .A(n653), .B(A[163]), .Z(n650) );
  XOR U748 ( .A(n653), .B(n654), .Z(DIFF[163]) );
  XOR U749 ( .A(B[163]), .B(A[163]), .Z(n654) );
  AND U750 ( .A(n655), .B(n656), .Z(n653) );
  NANDN U751 ( .A(B[162]), .B(n657), .Z(n656) );
  NANDN U752 ( .A(A[162]), .B(n658), .Z(n657) );
  NANDN U753 ( .A(n658), .B(A[162]), .Z(n655) );
  XOR U754 ( .A(n658), .B(n659), .Z(DIFF[162]) );
  XOR U755 ( .A(B[162]), .B(A[162]), .Z(n659) );
  AND U756 ( .A(n660), .B(n661), .Z(n658) );
  NANDN U757 ( .A(B[161]), .B(n662), .Z(n661) );
  NANDN U758 ( .A(A[161]), .B(n663), .Z(n662) );
  NANDN U759 ( .A(n663), .B(A[161]), .Z(n660) );
  XOR U760 ( .A(n663), .B(n664), .Z(DIFF[161]) );
  XOR U761 ( .A(B[161]), .B(A[161]), .Z(n664) );
  AND U762 ( .A(n665), .B(n666), .Z(n663) );
  NANDN U763 ( .A(B[160]), .B(n667), .Z(n666) );
  NANDN U764 ( .A(A[160]), .B(n668), .Z(n667) );
  NANDN U765 ( .A(n668), .B(A[160]), .Z(n665) );
  XOR U766 ( .A(n668), .B(n669), .Z(DIFF[160]) );
  XOR U767 ( .A(B[160]), .B(A[160]), .Z(n669) );
  AND U768 ( .A(n670), .B(n671), .Z(n668) );
  NANDN U769 ( .A(B[159]), .B(n672), .Z(n671) );
  NANDN U770 ( .A(A[159]), .B(n673), .Z(n672) );
  NANDN U771 ( .A(n673), .B(A[159]), .Z(n670) );
  XOR U772 ( .A(n674), .B(n675), .Z(DIFF[15]) );
  XOR U773 ( .A(B[15]), .B(A[15]), .Z(n675) );
  XOR U774 ( .A(n673), .B(n676), .Z(DIFF[159]) );
  XOR U775 ( .A(B[159]), .B(A[159]), .Z(n676) );
  AND U776 ( .A(n677), .B(n678), .Z(n673) );
  NANDN U777 ( .A(B[158]), .B(n679), .Z(n678) );
  NANDN U778 ( .A(A[158]), .B(n680), .Z(n679) );
  NANDN U779 ( .A(n680), .B(A[158]), .Z(n677) );
  XOR U780 ( .A(n680), .B(n681), .Z(DIFF[158]) );
  XOR U781 ( .A(B[158]), .B(A[158]), .Z(n681) );
  AND U782 ( .A(n682), .B(n683), .Z(n680) );
  NANDN U783 ( .A(B[157]), .B(n684), .Z(n683) );
  NANDN U784 ( .A(A[157]), .B(n685), .Z(n684) );
  NANDN U785 ( .A(n685), .B(A[157]), .Z(n682) );
  XOR U786 ( .A(n685), .B(n686), .Z(DIFF[157]) );
  XOR U787 ( .A(B[157]), .B(A[157]), .Z(n686) );
  AND U788 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U789 ( .A(B[156]), .B(n689), .Z(n688) );
  NANDN U790 ( .A(A[156]), .B(n690), .Z(n689) );
  NANDN U791 ( .A(n690), .B(A[156]), .Z(n687) );
  XOR U792 ( .A(n690), .B(n691), .Z(DIFF[156]) );
  XOR U793 ( .A(B[156]), .B(A[156]), .Z(n691) );
  AND U794 ( .A(n692), .B(n693), .Z(n690) );
  NANDN U795 ( .A(B[155]), .B(n694), .Z(n693) );
  NANDN U796 ( .A(A[155]), .B(n695), .Z(n694) );
  NANDN U797 ( .A(n695), .B(A[155]), .Z(n692) );
  XOR U798 ( .A(n695), .B(n696), .Z(DIFF[155]) );
  XOR U799 ( .A(B[155]), .B(A[155]), .Z(n696) );
  AND U800 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U801 ( .A(B[154]), .B(n699), .Z(n698) );
  NANDN U802 ( .A(A[154]), .B(n700), .Z(n699) );
  NANDN U803 ( .A(n700), .B(A[154]), .Z(n697) );
  XOR U804 ( .A(n700), .B(n701), .Z(DIFF[154]) );
  XOR U805 ( .A(B[154]), .B(A[154]), .Z(n701) );
  AND U806 ( .A(n702), .B(n703), .Z(n700) );
  NANDN U807 ( .A(B[153]), .B(n704), .Z(n703) );
  NANDN U808 ( .A(A[153]), .B(n705), .Z(n704) );
  NANDN U809 ( .A(n705), .B(A[153]), .Z(n702) );
  XOR U810 ( .A(n705), .B(n706), .Z(DIFF[153]) );
  XOR U811 ( .A(B[153]), .B(A[153]), .Z(n706) );
  AND U812 ( .A(n707), .B(n708), .Z(n705) );
  NANDN U813 ( .A(B[152]), .B(n709), .Z(n708) );
  NANDN U814 ( .A(A[152]), .B(n710), .Z(n709) );
  NANDN U815 ( .A(n710), .B(A[152]), .Z(n707) );
  XOR U816 ( .A(n710), .B(n711), .Z(DIFF[152]) );
  XOR U817 ( .A(B[152]), .B(A[152]), .Z(n711) );
  AND U818 ( .A(n712), .B(n713), .Z(n710) );
  NANDN U819 ( .A(B[151]), .B(n714), .Z(n713) );
  NANDN U820 ( .A(A[151]), .B(n715), .Z(n714) );
  NANDN U821 ( .A(n715), .B(A[151]), .Z(n712) );
  XOR U822 ( .A(n715), .B(n716), .Z(DIFF[151]) );
  XOR U823 ( .A(B[151]), .B(A[151]), .Z(n716) );
  AND U824 ( .A(n717), .B(n718), .Z(n715) );
  NANDN U825 ( .A(B[150]), .B(n719), .Z(n718) );
  NANDN U826 ( .A(A[150]), .B(n720), .Z(n719) );
  NANDN U827 ( .A(n720), .B(A[150]), .Z(n717) );
  XOR U828 ( .A(n720), .B(n721), .Z(DIFF[150]) );
  XOR U829 ( .A(B[150]), .B(A[150]), .Z(n721) );
  AND U830 ( .A(n722), .B(n723), .Z(n720) );
  NANDN U831 ( .A(B[149]), .B(n724), .Z(n723) );
  NANDN U832 ( .A(A[149]), .B(n725), .Z(n724) );
  NANDN U833 ( .A(n725), .B(A[149]), .Z(n722) );
  XOR U834 ( .A(n726), .B(n727), .Z(DIFF[14]) );
  XOR U835 ( .A(B[14]), .B(A[14]), .Z(n727) );
  XOR U836 ( .A(n725), .B(n728), .Z(DIFF[149]) );
  XOR U837 ( .A(B[149]), .B(A[149]), .Z(n728) );
  AND U838 ( .A(n729), .B(n730), .Z(n725) );
  NANDN U839 ( .A(B[148]), .B(n731), .Z(n730) );
  NANDN U840 ( .A(A[148]), .B(n732), .Z(n731) );
  NANDN U841 ( .A(n732), .B(A[148]), .Z(n729) );
  XOR U842 ( .A(n732), .B(n733), .Z(DIFF[148]) );
  XOR U843 ( .A(B[148]), .B(A[148]), .Z(n733) );
  AND U844 ( .A(n734), .B(n735), .Z(n732) );
  NANDN U845 ( .A(B[147]), .B(n736), .Z(n735) );
  NANDN U846 ( .A(A[147]), .B(n737), .Z(n736) );
  NANDN U847 ( .A(n737), .B(A[147]), .Z(n734) );
  XOR U848 ( .A(n737), .B(n738), .Z(DIFF[147]) );
  XOR U849 ( .A(B[147]), .B(A[147]), .Z(n738) );
  AND U850 ( .A(n739), .B(n740), .Z(n737) );
  NANDN U851 ( .A(B[146]), .B(n741), .Z(n740) );
  NANDN U852 ( .A(A[146]), .B(n742), .Z(n741) );
  NANDN U853 ( .A(n742), .B(A[146]), .Z(n739) );
  XOR U854 ( .A(n742), .B(n743), .Z(DIFF[146]) );
  XOR U855 ( .A(B[146]), .B(A[146]), .Z(n743) );
  AND U856 ( .A(n744), .B(n745), .Z(n742) );
  NANDN U857 ( .A(B[145]), .B(n746), .Z(n745) );
  NANDN U858 ( .A(A[145]), .B(n747), .Z(n746) );
  NANDN U859 ( .A(n747), .B(A[145]), .Z(n744) );
  XOR U860 ( .A(n747), .B(n748), .Z(DIFF[145]) );
  XOR U861 ( .A(B[145]), .B(A[145]), .Z(n748) );
  AND U862 ( .A(n749), .B(n750), .Z(n747) );
  NANDN U863 ( .A(B[144]), .B(n751), .Z(n750) );
  NANDN U864 ( .A(A[144]), .B(n752), .Z(n751) );
  NANDN U865 ( .A(n752), .B(A[144]), .Z(n749) );
  XOR U866 ( .A(n752), .B(n753), .Z(DIFF[144]) );
  XOR U867 ( .A(B[144]), .B(A[144]), .Z(n753) );
  AND U868 ( .A(n754), .B(n755), .Z(n752) );
  NANDN U869 ( .A(B[143]), .B(n756), .Z(n755) );
  NANDN U870 ( .A(A[143]), .B(n757), .Z(n756) );
  NANDN U871 ( .A(n757), .B(A[143]), .Z(n754) );
  XOR U872 ( .A(n757), .B(n758), .Z(DIFF[143]) );
  XOR U873 ( .A(B[143]), .B(A[143]), .Z(n758) );
  AND U874 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U875 ( .A(B[142]), .B(n761), .Z(n760) );
  NANDN U876 ( .A(A[142]), .B(n762), .Z(n761) );
  NANDN U877 ( .A(n762), .B(A[142]), .Z(n759) );
  XOR U878 ( .A(n762), .B(n763), .Z(DIFF[142]) );
  XOR U879 ( .A(B[142]), .B(A[142]), .Z(n763) );
  AND U880 ( .A(n764), .B(n765), .Z(n762) );
  NANDN U881 ( .A(B[141]), .B(n766), .Z(n765) );
  NANDN U882 ( .A(A[141]), .B(n767), .Z(n766) );
  NANDN U883 ( .A(n767), .B(A[141]), .Z(n764) );
  XOR U884 ( .A(n767), .B(n768), .Z(DIFF[141]) );
  XOR U885 ( .A(B[141]), .B(A[141]), .Z(n768) );
  AND U886 ( .A(n769), .B(n770), .Z(n767) );
  NANDN U887 ( .A(B[140]), .B(n771), .Z(n770) );
  NANDN U888 ( .A(A[140]), .B(n772), .Z(n771) );
  NANDN U889 ( .A(n772), .B(A[140]), .Z(n769) );
  XOR U890 ( .A(n772), .B(n773), .Z(DIFF[140]) );
  XOR U891 ( .A(B[140]), .B(A[140]), .Z(n773) );
  AND U892 ( .A(n774), .B(n775), .Z(n772) );
  NANDN U893 ( .A(B[139]), .B(n776), .Z(n775) );
  NANDN U894 ( .A(A[139]), .B(n777), .Z(n776) );
  NANDN U895 ( .A(n777), .B(A[139]), .Z(n774) );
  XOR U896 ( .A(n778), .B(n779), .Z(DIFF[13]) );
  XOR U897 ( .A(B[13]), .B(A[13]), .Z(n779) );
  XOR U898 ( .A(n777), .B(n780), .Z(DIFF[139]) );
  XOR U899 ( .A(B[139]), .B(A[139]), .Z(n780) );
  AND U900 ( .A(n781), .B(n782), .Z(n777) );
  NANDN U901 ( .A(B[138]), .B(n783), .Z(n782) );
  NANDN U902 ( .A(A[138]), .B(n784), .Z(n783) );
  NANDN U903 ( .A(n784), .B(A[138]), .Z(n781) );
  XOR U904 ( .A(n784), .B(n785), .Z(DIFF[138]) );
  XOR U905 ( .A(B[138]), .B(A[138]), .Z(n785) );
  AND U906 ( .A(n786), .B(n787), .Z(n784) );
  NANDN U907 ( .A(B[137]), .B(n788), .Z(n787) );
  NANDN U908 ( .A(A[137]), .B(n789), .Z(n788) );
  NANDN U909 ( .A(n789), .B(A[137]), .Z(n786) );
  XOR U910 ( .A(n789), .B(n790), .Z(DIFF[137]) );
  XOR U911 ( .A(B[137]), .B(A[137]), .Z(n790) );
  AND U912 ( .A(n791), .B(n792), .Z(n789) );
  NANDN U913 ( .A(B[136]), .B(n793), .Z(n792) );
  NANDN U914 ( .A(A[136]), .B(n794), .Z(n793) );
  NANDN U915 ( .A(n794), .B(A[136]), .Z(n791) );
  XOR U916 ( .A(n794), .B(n795), .Z(DIFF[136]) );
  XOR U917 ( .A(B[136]), .B(A[136]), .Z(n795) );
  AND U918 ( .A(n796), .B(n797), .Z(n794) );
  NANDN U919 ( .A(B[135]), .B(n798), .Z(n797) );
  NANDN U920 ( .A(A[135]), .B(n799), .Z(n798) );
  NANDN U921 ( .A(n799), .B(A[135]), .Z(n796) );
  XOR U922 ( .A(n799), .B(n800), .Z(DIFF[135]) );
  XOR U923 ( .A(B[135]), .B(A[135]), .Z(n800) );
  AND U924 ( .A(n801), .B(n802), .Z(n799) );
  NANDN U925 ( .A(B[134]), .B(n803), .Z(n802) );
  NANDN U926 ( .A(A[134]), .B(n804), .Z(n803) );
  NANDN U927 ( .A(n804), .B(A[134]), .Z(n801) );
  XOR U928 ( .A(n804), .B(n805), .Z(DIFF[134]) );
  XOR U929 ( .A(B[134]), .B(A[134]), .Z(n805) );
  AND U930 ( .A(n806), .B(n807), .Z(n804) );
  NANDN U931 ( .A(B[133]), .B(n808), .Z(n807) );
  NANDN U932 ( .A(A[133]), .B(n809), .Z(n808) );
  NANDN U933 ( .A(n809), .B(A[133]), .Z(n806) );
  XOR U934 ( .A(n809), .B(n810), .Z(DIFF[133]) );
  XOR U935 ( .A(B[133]), .B(A[133]), .Z(n810) );
  AND U936 ( .A(n811), .B(n812), .Z(n809) );
  NANDN U937 ( .A(B[132]), .B(n813), .Z(n812) );
  NANDN U938 ( .A(A[132]), .B(n814), .Z(n813) );
  NANDN U939 ( .A(n814), .B(A[132]), .Z(n811) );
  XOR U940 ( .A(n814), .B(n815), .Z(DIFF[132]) );
  XOR U941 ( .A(B[132]), .B(A[132]), .Z(n815) );
  AND U942 ( .A(n816), .B(n817), .Z(n814) );
  NANDN U943 ( .A(B[131]), .B(n818), .Z(n817) );
  NANDN U944 ( .A(A[131]), .B(n819), .Z(n818) );
  NANDN U945 ( .A(n819), .B(A[131]), .Z(n816) );
  XOR U946 ( .A(n819), .B(n820), .Z(DIFF[131]) );
  XOR U947 ( .A(B[131]), .B(A[131]), .Z(n820) );
  AND U948 ( .A(n821), .B(n822), .Z(n819) );
  NANDN U949 ( .A(B[130]), .B(n823), .Z(n822) );
  NANDN U950 ( .A(A[130]), .B(n824), .Z(n823) );
  NANDN U951 ( .A(n824), .B(A[130]), .Z(n821) );
  XOR U952 ( .A(n824), .B(n825), .Z(DIFF[130]) );
  XOR U953 ( .A(B[130]), .B(A[130]), .Z(n825) );
  AND U954 ( .A(n826), .B(n827), .Z(n824) );
  NANDN U955 ( .A(B[129]), .B(n828), .Z(n827) );
  NANDN U956 ( .A(A[129]), .B(n829), .Z(n828) );
  NANDN U957 ( .A(n829), .B(A[129]), .Z(n826) );
  XOR U958 ( .A(n830), .B(n831), .Z(DIFF[12]) );
  XOR U959 ( .A(B[12]), .B(A[12]), .Z(n831) );
  XOR U960 ( .A(n829), .B(n832), .Z(DIFF[129]) );
  XOR U961 ( .A(B[129]), .B(A[129]), .Z(n832) );
  AND U962 ( .A(n833), .B(n834), .Z(n829) );
  NANDN U963 ( .A(B[128]), .B(n835), .Z(n834) );
  NANDN U964 ( .A(A[128]), .B(n836), .Z(n835) );
  NANDN U965 ( .A(n836), .B(A[128]), .Z(n833) );
  XOR U966 ( .A(n836), .B(n837), .Z(DIFF[128]) );
  XOR U967 ( .A(B[128]), .B(A[128]), .Z(n837) );
  AND U968 ( .A(n838), .B(n839), .Z(n836) );
  NANDN U969 ( .A(B[127]), .B(n840), .Z(n839) );
  NANDN U970 ( .A(A[127]), .B(n841), .Z(n840) );
  NANDN U971 ( .A(n841), .B(A[127]), .Z(n838) );
  XOR U972 ( .A(n841), .B(n842), .Z(DIFF[127]) );
  XOR U973 ( .A(B[127]), .B(A[127]), .Z(n842) );
  AND U974 ( .A(n843), .B(n844), .Z(n841) );
  NANDN U975 ( .A(B[126]), .B(n845), .Z(n844) );
  NANDN U976 ( .A(A[126]), .B(n846), .Z(n845) );
  NANDN U977 ( .A(n846), .B(A[126]), .Z(n843) );
  XOR U978 ( .A(n846), .B(n847), .Z(DIFF[126]) );
  XOR U979 ( .A(B[126]), .B(A[126]), .Z(n847) );
  AND U980 ( .A(n848), .B(n849), .Z(n846) );
  NANDN U981 ( .A(B[125]), .B(n850), .Z(n849) );
  NANDN U982 ( .A(A[125]), .B(n851), .Z(n850) );
  NANDN U983 ( .A(n851), .B(A[125]), .Z(n848) );
  XOR U984 ( .A(n851), .B(n852), .Z(DIFF[125]) );
  XOR U985 ( .A(B[125]), .B(A[125]), .Z(n852) );
  AND U986 ( .A(n853), .B(n854), .Z(n851) );
  NANDN U987 ( .A(B[124]), .B(n855), .Z(n854) );
  NANDN U988 ( .A(A[124]), .B(n856), .Z(n855) );
  NANDN U989 ( .A(n856), .B(A[124]), .Z(n853) );
  XOR U990 ( .A(n856), .B(n857), .Z(DIFF[124]) );
  XOR U991 ( .A(B[124]), .B(A[124]), .Z(n857) );
  AND U992 ( .A(n858), .B(n859), .Z(n856) );
  NANDN U993 ( .A(B[123]), .B(n860), .Z(n859) );
  NANDN U994 ( .A(A[123]), .B(n861), .Z(n860) );
  NANDN U995 ( .A(n861), .B(A[123]), .Z(n858) );
  XOR U996 ( .A(n861), .B(n862), .Z(DIFF[123]) );
  XOR U997 ( .A(B[123]), .B(A[123]), .Z(n862) );
  AND U998 ( .A(n863), .B(n864), .Z(n861) );
  NANDN U999 ( .A(B[122]), .B(n865), .Z(n864) );
  NANDN U1000 ( .A(A[122]), .B(n866), .Z(n865) );
  NANDN U1001 ( .A(n866), .B(A[122]), .Z(n863) );
  XOR U1002 ( .A(n866), .B(n867), .Z(DIFF[122]) );
  XOR U1003 ( .A(B[122]), .B(A[122]), .Z(n867) );
  AND U1004 ( .A(n868), .B(n869), .Z(n866) );
  NANDN U1005 ( .A(B[121]), .B(n870), .Z(n869) );
  NANDN U1006 ( .A(A[121]), .B(n871), .Z(n870) );
  NANDN U1007 ( .A(n871), .B(A[121]), .Z(n868) );
  XOR U1008 ( .A(n871), .B(n872), .Z(DIFF[121]) );
  XOR U1009 ( .A(B[121]), .B(A[121]), .Z(n872) );
  AND U1010 ( .A(n873), .B(n874), .Z(n871) );
  NANDN U1011 ( .A(B[120]), .B(n875), .Z(n874) );
  NANDN U1012 ( .A(A[120]), .B(n876), .Z(n875) );
  NANDN U1013 ( .A(n876), .B(A[120]), .Z(n873) );
  XOR U1014 ( .A(n876), .B(n877), .Z(DIFF[120]) );
  XOR U1015 ( .A(B[120]), .B(A[120]), .Z(n877) );
  AND U1016 ( .A(n878), .B(n879), .Z(n876) );
  NANDN U1017 ( .A(B[119]), .B(n880), .Z(n879) );
  NANDN U1018 ( .A(A[119]), .B(n881), .Z(n880) );
  NANDN U1019 ( .A(n881), .B(A[119]), .Z(n878) );
  XOR U1020 ( .A(n882), .B(n883), .Z(DIFF[11]) );
  XOR U1021 ( .A(B[11]), .B(A[11]), .Z(n883) );
  XOR U1022 ( .A(n881), .B(n884), .Z(DIFF[119]) );
  XOR U1023 ( .A(B[119]), .B(A[119]), .Z(n884) );
  AND U1024 ( .A(n885), .B(n886), .Z(n881) );
  NANDN U1025 ( .A(B[118]), .B(n887), .Z(n886) );
  NANDN U1026 ( .A(A[118]), .B(n888), .Z(n887) );
  NANDN U1027 ( .A(n888), .B(A[118]), .Z(n885) );
  XOR U1028 ( .A(n888), .B(n889), .Z(DIFF[118]) );
  XOR U1029 ( .A(B[118]), .B(A[118]), .Z(n889) );
  AND U1030 ( .A(n890), .B(n891), .Z(n888) );
  NANDN U1031 ( .A(B[117]), .B(n892), .Z(n891) );
  NANDN U1032 ( .A(A[117]), .B(n893), .Z(n892) );
  NANDN U1033 ( .A(n893), .B(A[117]), .Z(n890) );
  XOR U1034 ( .A(n893), .B(n894), .Z(DIFF[117]) );
  XOR U1035 ( .A(B[117]), .B(A[117]), .Z(n894) );
  AND U1036 ( .A(n895), .B(n896), .Z(n893) );
  NANDN U1037 ( .A(B[116]), .B(n897), .Z(n896) );
  NANDN U1038 ( .A(A[116]), .B(n898), .Z(n897) );
  NANDN U1039 ( .A(n898), .B(A[116]), .Z(n895) );
  XOR U1040 ( .A(n898), .B(n899), .Z(DIFF[116]) );
  XOR U1041 ( .A(B[116]), .B(A[116]), .Z(n899) );
  AND U1042 ( .A(n900), .B(n901), .Z(n898) );
  NANDN U1043 ( .A(B[115]), .B(n902), .Z(n901) );
  NANDN U1044 ( .A(A[115]), .B(n903), .Z(n902) );
  NANDN U1045 ( .A(n903), .B(A[115]), .Z(n900) );
  XOR U1046 ( .A(n903), .B(n904), .Z(DIFF[115]) );
  XOR U1047 ( .A(B[115]), .B(A[115]), .Z(n904) );
  AND U1048 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U1049 ( .A(B[114]), .B(n907), .Z(n906) );
  NANDN U1050 ( .A(A[114]), .B(n908), .Z(n907) );
  NANDN U1051 ( .A(n908), .B(A[114]), .Z(n905) );
  XOR U1052 ( .A(n908), .B(n909), .Z(DIFF[114]) );
  XOR U1053 ( .A(B[114]), .B(A[114]), .Z(n909) );
  AND U1054 ( .A(n910), .B(n911), .Z(n908) );
  NANDN U1055 ( .A(B[113]), .B(n912), .Z(n911) );
  NANDN U1056 ( .A(A[113]), .B(n913), .Z(n912) );
  NANDN U1057 ( .A(n913), .B(A[113]), .Z(n910) );
  XOR U1058 ( .A(n913), .B(n914), .Z(DIFF[113]) );
  XOR U1059 ( .A(B[113]), .B(A[113]), .Z(n914) );
  AND U1060 ( .A(n915), .B(n916), .Z(n913) );
  NANDN U1061 ( .A(B[112]), .B(n917), .Z(n916) );
  NANDN U1062 ( .A(A[112]), .B(n918), .Z(n917) );
  NANDN U1063 ( .A(n918), .B(A[112]), .Z(n915) );
  XOR U1064 ( .A(n918), .B(n919), .Z(DIFF[112]) );
  XOR U1065 ( .A(B[112]), .B(A[112]), .Z(n919) );
  AND U1066 ( .A(n920), .B(n921), .Z(n918) );
  NANDN U1067 ( .A(B[111]), .B(n922), .Z(n921) );
  NANDN U1068 ( .A(A[111]), .B(n923), .Z(n922) );
  NANDN U1069 ( .A(n923), .B(A[111]), .Z(n920) );
  XOR U1070 ( .A(n923), .B(n924), .Z(DIFF[111]) );
  XOR U1071 ( .A(B[111]), .B(A[111]), .Z(n924) );
  AND U1072 ( .A(n925), .B(n926), .Z(n923) );
  NANDN U1073 ( .A(B[110]), .B(n927), .Z(n926) );
  NANDN U1074 ( .A(A[110]), .B(n928), .Z(n927) );
  NANDN U1075 ( .A(n928), .B(A[110]), .Z(n925) );
  XOR U1076 ( .A(n928), .B(n929), .Z(DIFF[110]) );
  XOR U1077 ( .A(B[110]), .B(A[110]), .Z(n929) );
  AND U1078 ( .A(n930), .B(n931), .Z(n928) );
  NANDN U1079 ( .A(B[109]), .B(n932), .Z(n931) );
  NANDN U1080 ( .A(A[109]), .B(n933), .Z(n932) );
  NANDN U1081 ( .A(n933), .B(A[109]), .Z(n930) );
  XOR U1082 ( .A(n934), .B(n935), .Z(DIFF[10]) );
  XOR U1083 ( .A(B[10]), .B(A[10]), .Z(n935) );
  XOR U1084 ( .A(n933), .B(n936), .Z(DIFF[109]) );
  XOR U1085 ( .A(B[109]), .B(A[109]), .Z(n936) );
  AND U1086 ( .A(n937), .B(n938), .Z(n933) );
  NANDN U1087 ( .A(B[108]), .B(n939), .Z(n938) );
  NANDN U1088 ( .A(A[108]), .B(n940), .Z(n939) );
  NANDN U1089 ( .A(n940), .B(A[108]), .Z(n937) );
  XOR U1090 ( .A(n940), .B(n941), .Z(DIFF[108]) );
  XOR U1091 ( .A(B[108]), .B(A[108]), .Z(n941) );
  AND U1092 ( .A(n942), .B(n943), .Z(n940) );
  NANDN U1093 ( .A(B[107]), .B(n944), .Z(n943) );
  NANDN U1094 ( .A(A[107]), .B(n945), .Z(n944) );
  NANDN U1095 ( .A(n945), .B(A[107]), .Z(n942) );
  XOR U1096 ( .A(n945), .B(n946), .Z(DIFF[107]) );
  XOR U1097 ( .A(B[107]), .B(A[107]), .Z(n946) );
  AND U1098 ( .A(n947), .B(n948), .Z(n945) );
  NANDN U1099 ( .A(B[106]), .B(n949), .Z(n948) );
  NANDN U1100 ( .A(A[106]), .B(n950), .Z(n949) );
  NANDN U1101 ( .A(n950), .B(A[106]), .Z(n947) );
  XOR U1102 ( .A(n950), .B(n951), .Z(DIFF[106]) );
  XOR U1103 ( .A(B[106]), .B(A[106]), .Z(n951) );
  AND U1104 ( .A(n952), .B(n953), .Z(n950) );
  NANDN U1105 ( .A(B[105]), .B(n954), .Z(n953) );
  NANDN U1106 ( .A(A[105]), .B(n955), .Z(n954) );
  NANDN U1107 ( .A(n955), .B(A[105]), .Z(n952) );
  XOR U1108 ( .A(n955), .B(n956), .Z(DIFF[105]) );
  XOR U1109 ( .A(B[105]), .B(A[105]), .Z(n956) );
  AND U1110 ( .A(n957), .B(n958), .Z(n955) );
  NANDN U1111 ( .A(B[104]), .B(n959), .Z(n958) );
  NANDN U1112 ( .A(A[104]), .B(n960), .Z(n959) );
  NANDN U1113 ( .A(n960), .B(A[104]), .Z(n957) );
  XOR U1114 ( .A(n960), .B(n961), .Z(DIFF[104]) );
  XOR U1115 ( .A(B[104]), .B(A[104]), .Z(n961) );
  AND U1116 ( .A(n962), .B(n963), .Z(n960) );
  NANDN U1117 ( .A(B[103]), .B(n964), .Z(n963) );
  NANDN U1118 ( .A(A[103]), .B(n965), .Z(n964) );
  NANDN U1119 ( .A(n965), .B(A[103]), .Z(n962) );
  XOR U1120 ( .A(n965), .B(n966), .Z(DIFF[103]) );
  XOR U1121 ( .A(B[103]), .B(A[103]), .Z(n966) );
  AND U1122 ( .A(n967), .B(n968), .Z(n965) );
  NANDN U1123 ( .A(B[102]), .B(n969), .Z(n968) );
  NANDN U1124 ( .A(A[102]), .B(n970), .Z(n969) );
  NANDN U1125 ( .A(n970), .B(A[102]), .Z(n967) );
  XOR U1126 ( .A(n970), .B(n971), .Z(DIFF[102]) );
  XOR U1127 ( .A(B[102]), .B(A[102]), .Z(n971) );
  AND U1128 ( .A(n972), .B(n973), .Z(n970) );
  NANDN U1129 ( .A(B[101]), .B(n974), .Z(n973) );
  NANDN U1130 ( .A(A[101]), .B(n975), .Z(n974) );
  NANDN U1131 ( .A(n975), .B(A[101]), .Z(n972) );
  XOR U1132 ( .A(n975), .B(n976), .Z(DIFF[101]) );
  XOR U1133 ( .A(B[101]), .B(A[101]), .Z(n976) );
  AND U1134 ( .A(n977), .B(n978), .Z(n975) );
  NANDN U1135 ( .A(B[100]), .B(n979), .Z(n978) );
  NANDN U1136 ( .A(A[100]), .B(n980), .Z(n979) );
  NANDN U1137 ( .A(n980), .B(A[100]), .Z(n977) );
  XOR U1138 ( .A(n980), .B(n981), .Z(DIFF[100]) );
  XOR U1139 ( .A(B[100]), .B(A[100]), .Z(n981) );
  AND U1140 ( .A(n982), .B(n983), .Z(n980) );
  NANDN U1141 ( .A(B[99]), .B(n984), .Z(n983) );
  OR U1142 ( .A(n5), .B(A[99]), .Z(n984) );
  NAND U1143 ( .A(A[99]), .B(n5), .Z(n982) );
  NAND U1144 ( .A(n985), .B(n986), .Z(n5) );
  NANDN U1145 ( .A(B[98]), .B(n987), .Z(n986) );
  NANDN U1146 ( .A(A[98]), .B(n7), .Z(n987) );
  NANDN U1147 ( .A(n7), .B(A[98]), .Z(n985) );
  AND U1148 ( .A(n988), .B(n989), .Z(n7) );
  NANDN U1149 ( .A(B[97]), .B(n990), .Z(n989) );
  NANDN U1150 ( .A(A[97]), .B(n9), .Z(n990) );
  NANDN U1151 ( .A(n9), .B(A[97]), .Z(n988) );
  AND U1152 ( .A(n991), .B(n992), .Z(n9) );
  NANDN U1153 ( .A(B[96]), .B(n993), .Z(n992) );
  NANDN U1154 ( .A(A[96]), .B(n11), .Z(n993) );
  NANDN U1155 ( .A(n11), .B(A[96]), .Z(n991) );
  AND U1156 ( .A(n994), .B(n995), .Z(n11) );
  NANDN U1157 ( .A(B[95]), .B(n996), .Z(n995) );
  NANDN U1158 ( .A(A[95]), .B(n13), .Z(n996) );
  NANDN U1159 ( .A(n13), .B(A[95]), .Z(n994) );
  AND U1160 ( .A(n997), .B(n998), .Z(n13) );
  NANDN U1161 ( .A(B[94]), .B(n999), .Z(n998) );
  NANDN U1162 ( .A(A[94]), .B(n15), .Z(n999) );
  NANDN U1163 ( .A(n15), .B(A[94]), .Z(n997) );
  AND U1164 ( .A(n1000), .B(n1001), .Z(n15) );
  NANDN U1165 ( .A(B[93]), .B(n1002), .Z(n1001) );
  NANDN U1166 ( .A(A[93]), .B(n17), .Z(n1002) );
  NANDN U1167 ( .A(n17), .B(A[93]), .Z(n1000) );
  AND U1168 ( .A(n1003), .B(n1004), .Z(n17) );
  NANDN U1169 ( .A(B[92]), .B(n1005), .Z(n1004) );
  NANDN U1170 ( .A(A[92]), .B(n19), .Z(n1005) );
  NANDN U1171 ( .A(n19), .B(A[92]), .Z(n1003) );
  AND U1172 ( .A(n1006), .B(n1007), .Z(n19) );
  NANDN U1173 ( .A(B[91]), .B(n1008), .Z(n1007) );
  NANDN U1174 ( .A(A[91]), .B(n21), .Z(n1008) );
  NANDN U1175 ( .A(n21), .B(A[91]), .Z(n1006) );
  AND U1176 ( .A(n1009), .B(n1010), .Z(n21) );
  NANDN U1177 ( .A(B[90]), .B(n1011), .Z(n1010) );
  NANDN U1178 ( .A(A[90]), .B(n23), .Z(n1011) );
  NANDN U1179 ( .A(n23), .B(A[90]), .Z(n1009) );
  AND U1180 ( .A(n1012), .B(n1013), .Z(n23) );
  NANDN U1181 ( .A(B[89]), .B(n1014), .Z(n1013) );
  NANDN U1182 ( .A(A[89]), .B(n27), .Z(n1014) );
  NANDN U1183 ( .A(n27), .B(A[89]), .Z(n1012) );
  AND U1184 ( .A(n1015), .B(n1016), .Z(n27) );
  NANDN U1185 ( .A(B[88]), .B(n1017), .Z(n1016) );
  NANDN U1186 ( .A(A[88]), .B(n29), .Z(n1017) );
  NANDN U1187 ( .A(n29), .B(A[88]), .Z(n1015) );
  AND U1188 ( .A(n1018), .B(n1019), .Z(n29) );
  NANDN U1189 ( .A(B[87]), .B(n1020), .Z(n1019) );
  NANDN U1190 ( .A(A[87]), .B(n31), .Z(n1020) );
  NANDN U1191 ( .A(n31), .B(A[87]), .Z(n1018) );
  AND U1192 ( .A(n1021), .B(n1022), .Z(n31) );
  NANDN U1193 ( .A(B[86]), .B(n1023), .Z(n1022) );
  NANDN U1194 ( .A(A[86]), .B(n33), .Z(n1023) );
  NANDN U1195 ( .A(n33), .B(A[86]), .Z(n1021) );
  AND U1196 ( .A(n1024), .B(n1025), .Z(n33) );
  NANDN U1197 ( .A(B[85]), .B(n1026), .Z(n1025) );
  NANDN U1198 ( .A(A[85]), .B(n35), .Z(n1026) );
  NANDN U1199 ( .A(n35), .B(A[85]), .Z(n1024) );
  AND U1200 ( .A(n1027), .B(n1028), .Z(n35) );
  NANDN U1201 ( .A(B[84]), .B(n1029), .Z(n1028) );
  NANDN U1202 ( .A(A[84]), .B(n37), .Z(n1029) );
  NANDN U1203 ( .A(n37), .B(A[84]), .Z(n1027) );
  AND U1204 ( .A(n1030), .B(n1031), .Z(n37) );
  NANDN U1205 ( .A(B[83]), .B(n1032), .Z(n1031) );
  NANDN U1206 ( .A(A[83]), .B(n39), .Z(n1032) );
  NANDN U1207 ( .A(n39), .B(A[83]), .Z(n1030) );
  AND U1208 ( .A(n1033), .B(n1034), .Z(n39) );
  NANDN U1209 ( .A(B[82]), .B(n1035), .Z(n1034) );
  NANDN U1210 ( .A(A[82]), .B(n41), .Z(n1035) );
  NANDN U1211 ( .A(n41), .B(A[82]), .Z(n1033) );
  AND U1212 ( .A(n1036), .B(n1037), .Z(n41) );
  NANDN U1213 ( .A(B[81]), .B(n1038), .Z(n1037) );
  NANDN U1214 ( .A(A[81]), .B(n43), .Z(n1038) );
  NANDN U1215 ( .A(n43), .B(A[81]), .Z(n1036) );
  AND U1216 ( .A(n1039), .B(n1040), .Z(n43) );
  NANDN U1217 ( .A(B[80]), .B(n1041), .Z(n1040) );
  NANDN U1218 ( .A(A[80]), .B(n45), .Z(n1041) );
  NANDN U1219 ( .A(n45), .B(A[80]), .Z(n1039) );
  AND U1220 ( .A(n1042), .B(n1043), .Z(n45) );
  NANDN U1221 ( .A(B[79]), .B(n1044), .Z(n1043) );
  NANDN U1222 ( .A(A[79]), .B(n49), .Z(n1044) );
  NANDN U1223 ( .A(n49), .B(A[79]), .Z(n1042) );
  AND U1224 ( .A(n1045), .B(n1046), .Z(n49) );
  NANDN U1225 ( .A(B[78]), .B(n1047), .Z(n1046) );
  NANDN U1226 ( .A(A[78]), .B(n51), .Z(n1047) );
  NANDN U1227 ( .A(n51), .B(A[78]), .Z(n1045) );
  AND U1228 ( .A(n1048), .B(n1049), .Z(n51) );
  NANDN U1229 ( .A(B[77]), .B(n1050), .Z(n1049) );
  NANDN U1230 ( .A(A[77]), .B(n53), .Z(n1050) );
  NANDN U1231 ( .A(n53), .B(A[77]), .Z(n1048) );
  AND U1232 ( .A(n1051), .B(n1052), .Z(n53) );
  NANDN U1233 ( .A(B[76]), .B(n1053), .Z(n1052) );
  NANDN U1234 ( .A(A[76]), .B(n55), .Z(n1053) );
  NANDN U1235 ( .A(n55), .B(A[76]), .Z(n1051) );
  AND U1236 ( .A(n1054), .B(n1055), .Z(n55) );
  NANDN U1237 ( .A(B[75]), .B(n1056), .Z(n1055) );
  NANDN U1238 ( .A(A[75]), .B(n57), .Z(n1056) );
  NANDN U1239 ( .A(n57), .B(A[75]), .Z(n1054) );
  AND U1240 ( .A(n1057), .B(n1058), .Z(n57) );
  NANDN U1241 ( .A(B[74]), .B(n1059), .Z(n1058) );
  NANDN U1242 ( .A(A[74]), .B(n59), .Z(n1059) );
  NANDN U1243 ( .A(n59), .B(A[74]), .Z(n1057) );
  AND U1244 ( .A(n1060), .B(n1061), .Z(n59) );
  NANDN U1245 ( .A(B[73]), .B(n1062), .Z(n1061) );
  NANDN U1246 ( .A(A[73]), .B(n61), .Z(n1062) );
  NANDN U1247 ( .A(n61), .B(A[73]), .Z(n1060) );
  AND U1248 ( .A(n1063), .B(n1064), .Z(n61) );
  NANDN U1249 ( .A(B[72]), .B(n1065), .Z(n1064) );
  NANDN U1250 ( .A(A[72]), .B(n63), .Z(n1065) );
  NANDN U1251 ( .A(n63), .B(A[72]), .Z(n1063) );
  AND U1252 ( .A(n1066), .B(n1067), .Z(n63) );
  NANDN U1253 ( .A(B[71]), .B(n1068), .Z(n1067) );
  NANDN U1254 ( .A(A[71]), .B(n65), .Z(n1068) );
  NANDN U1255 ( .A(n65), .B(A[71]), .Z(n1066) );
  AND U1256 ( .A(n1069), .B(n1070), .Z(n65) );
  NANDN U1257 ( .A(B[70]), .B(n1071), .Z(n1070) );
  NANDN U1258 ( .A(A[70]), .B(n67), .Z(n1071) );
  NANDN U1259 ( .A(n67), .B(A[70]), .Z(n1069) );
  AND U1260 ( .A(n1072), .B(n1073), .Z(n67) );
  NANDN U1261 ( .A(B[69]), .B(n1074), .Z(n1073) );
  NANDN U1262 ( .A(A[69]), .B(n71), .Z(n1074) );
  NANDN U1263 ( .A(n71), .B(A[69]), .Z(n1072) );
  AND U1264 ( .A(n1075), .B(n1076), .Z(n71) );
  NANDN U1265 ( .A(B[68]), .B(n1077), .Z(n1076) );
  NANDN U1266 ( .A(A[68]), .B(n73), .Z(n1077) );
  NANDN U1267 ( .A(n73), .B(A[68]), .Z(n1075) );
  AND U1268 ( .A(n1078), .B(n1079), .Z(n73) );
  NANDN U1269 ( .A(B[67]), .B(n1080), .Z(n1079) );
  NANDN U1270 ( .A(A[67]), .B(n75), .Z(n1080) );
  NANDN U1271 ( .A(n75), .B(A[67]), .Z(n1078) );
  AND U1272 ( .A(n1081), .B(n1082), .Z(n75) );
  NANDN U1273 ( .A(B[66]), .B(n1083), .Z(n1082) );
  NANDN U1274 ( .A(A[66]), .B(n77), .Z(n1083) );
  NANDN U1275 ( .A(n77), .B(A[66]), .Z(n1081) );
  AND U1276 ( .A(n1084), .B(n1085), .Z(n77) );
  NANDN U1277 ( .A(B[65]), .B(n1086), .Z(n1085) );
  NANDN U1278 ( .A(A[65]), .B(n79), .Z(n1086) );
  NANDN U1279 ( .A(n79), .B(A[65]), .Z(n1084) );
  AND U1280 ( .A(n1087), .B(n1088), .Z(n79) );
  NANDN U1281 ( .A(B[64]), .B(n1089), .Z(n1088) );
  NANDN U1282 ( .A(A[64]), .B(n81), .Z(n1089) );
  NANDN U1283 ( .A(n81), .B(A[64]), .Z(n1087) );
  AND U1284 ( .A(n1090), .B(n1091), .Z(n81) );
  NANDN U1285 ( .A(B[63]), .B(n1092), .Z(n1091) );
  NANDN U1286 ( .A(A[63]), .B(n83), .Z(n1092) );
  NANDN U1287 ( .A(n83), .B(A[63]), .Z(n1090) );
  AND U1288 ( .A(n1093), .B(n1094), .Z(n83) );
  NANDN U1289 ( .A(B[62]), .B(n1095), .Z(n1094) );
  NANDN U1290 ( .A(A[62]), .B(n85), .Z(n1095) );
  NANDN U1291 ( .A(n85), .B(A[62]), .Z(n1093) );
  AND U1292 ( .A(n1096), .B(n1097), .Z(n85) );
  NANDN U1293 ( .A(B[61]), .B(n1098), .Z(n1097) );
  NANDN U1294 ( .A(A[61]), .B(n87), .Z(n1098) );
  NANDN U1295 ( .A(n87), .B(A[61]), .Z(n1096) );
  AND U1296 ( .A(n1099), .B(n1100), .Z(n87) );
  NANDN U1297 ( .A(B[60]), .B(n1101), .Z(n1100) );
  NANDN U1298 ( .A(A[60]), .B(n89), .Z(n1101) );
  NANDN U1299 ( .A(n89), .B(A[60]), .Z(n1099) );
  AND U1300 ( .A(n1102), .B(n1103), .Z(n89) );
  NANDN U1301 ( .A(B[59]), .B(n1104), .Z(n1103) );
  NANDN U1302 ( .A(A[59]), .B(n93), .Z(n1104) );
  NANDN U1303 ( .A(n93), .B(A[59]), .Z(n1102) );
  AND U1304 ( .A(n1105), .B(n1106), .Z(n93) );
  NANDN U1305 ( .A(B[58]), .B(n1107), .Z(n1106) );
  NANDN U1306 ( .A(A[58]), .B(n95), .Z(n1107) );
  NANDN U1307 ( .A(n95), .B(A[58]), .Z(n1105) );
  AND U1308 ( .A(n1108), .B(n1109), .Z(n95) );
  NANDN U1309 ( .A(B[57]), .B(n1110), .Z(n1109) );
  NANDN U1310 ( .A(A[57]), .B(n97), .Z(n1110) );
  NANDN U1311 ( .A(n97), .B(A[57]), .Z(n1108) );
  AND U1312 ( .A(n1111), .B(n1112), .Z(n97) );
  NANDN U1313 ( .A(B[56]), .B(n1113), .Z(n1112) );
  NANDN U1314 ( .A(A[56]), .B(n99), .Z(n1113) );
  NANDN U1315 ( .A(n99), .B(A[56]), .Z(n1111) );
  AND U1316 ( .A(n1114), .B(n1115), .Z(n99) );
  NANDN U1317 ( .A(B[55]), .B(n1116), .Z(n1115) );
  NANDN U1318 ( .A(A[55]), .B(n101), .Z(n1116) );
  NANDN U1319 ( .A(n101), .B(A[55]), .Z(n1114) );
  AND U1320 ( .A(n1117), .B(n1118), .Z(n101) );
  NANDN U1321 ( .A(B[54]), .B(n1119), .Z(n1118) );
  NANDN U1322 ( .A(A[54]), .B(n103), .Z(n1119) );
  NANDN U1323 ( .A(n103), .B(A[54]), .Z(n1117) );
  AND U1324 ( .A(n1120), .B(n1121), .Z(n103) );
  NANDN U1325 ( .A(B[53]), .B(n1122), .Z(n1121) );
  NANDN U1326 ( .A(A[53]), .B(n105), .Z(n1122) );
  NANDN U1327 ( .A(n105), .B(A[53]), .Z(n1120) );
  AND U1328 ( .A(n1123), .B(n1124), .Z(n105) );
  NANDN U1329 ( .A(B[52]), .B(n1125), .Z(n1124) );
  NANDN U1330 ( .A(A[52]), .B(n107), .Z(n1125) );
  NANDN U1331 ( .A(n107), .B(A[52]), .Z(n1123) );
  AND U1332 ( .A(n1126), .B(n1127), .Z(n107) );
  NANDN U1333 ( .A(B[51]), .B(n1128), .Z(n1127) );
  NANDN U1334 ( .A(A[51]), .B(n109), .Z(n1128) );
  NANDN U1335 ( .A(n109), .B(A[51]), .Z(n1126) );
  AND U1336 ( .A(n1129), .B(n1130), .Z(n109) );
  NANDN U1337 ( .A(B[50]), .B(n1131), .Z(n1130) );
  NANDN U1338 ( .A(A[50]), .B(n111), .Z(n1131) );
  NANDN U1339 ( .A(n111), .B(A[50]), .Z(n1129) );
  AND U1340 ( .A(n1132), .B(n1133), .Z(n111) );
  NANDN U1341 ( .A(B[49]), .B(n1134), .Z(n1133) );
  NANDN U1342 ( .A(A[49]), .B(n115), .Z(n1134) );
  NANDN U1343 ( .A(n115), .B(A[49]), .Z(n1132) );
  AND U1344 ( .A(n1135), .B(n1136), .Z(n115) );
  NANDN U1345 ( .A(B[48]), .B(n1137), .Z(n1136) );
  NANDN U1346 ( .A(A[48]), .B(n117), .Z(n1137) );
  NANDN U1347 ( .A(n117), .B(A[48]), .Z(n1135) );
  AND U1348 ( .A(n1138), .B(n1139), .Z(n117) );
  NANDN U1349 ( .A(B[47]), .B(n1140), .Z(n1139) );
  NANDN U1350 ( .A(A[47]), .B(n119), .Z(n1140) );
  NANDN U1351 ( .A(n119), .B(A[47]), .Z(n1138) );
  AND U1352 ( .A(n1141), .B(n1142), .Z(n119) );
  NANDN U1353 ( .A(B[46]), .B(n1143), .Z(n1142) );
  NANDN U1354 ( .A(A[46]), .B(n121), .Z(n1143) );
  NANDN U1355 ( .A(n121), .B(A[46]), .Z(n1141) );
  AND U1356 ( .A(n1144), .B(n1145), .Z(n121) );
  NANDN U1357 ( .A(B[45]), .B(n1146), .Z(n1145) );
  NANDN U1358 ( .A(A[45]), .B(n123), .Z(n1146) );
  NANDN U1359 ( .A(n123), .B(A[45]), .Z(n1144) );
  AND U1360 ( .A(n1147), .B(n1148), .Z(n123) );
  NANDN U1361 ( .A(B[44]), .B(n1149), .Z(n1148) );
  NANDN U1362 ( .A(A[44]), .B(n125), .Z(n1149) );
  NANDN U1363 ( .A(n125), .B(A[44]), .Z(n1147) );
  AND U1364 ( .A(n1150), .B(n1151), .Z(n125) );
  NANDN U1365 ( .A(B[43]), .B(n1152), .Z(n1151) );
  NANDN U1366 ( .A(A[43]), .B(n127), .Z(n1152) );
  NANDN U1367 ( .A(n127), .B(A[43]), .Z(n1150) );
  AND U1368 ( .A(n1153), .B(n1154), .Z(n127) );
  NANDN U1369 ( .A(B[42]), .B(n1155), .Z(n1154) );
  NANDN U1370 ( .A(A[42]), .B(n129), .Z(n1155) );
  NANDN U1371 ( .A(n129), .B(A[42]), .Z(n1153) );
  AND U1372 ( .A(n1156), .B(n1157), .Z(n129) );
  NANDN U1373 ( .A(B[41]), .B(n1158), .Z(n1157) );
  NANDN U1374 ( .A(A[41]), .B(n131), .Z(n1158) );
  NANDN U1375 ( .A(n131), .B(A[41]), .Z(n1156) );
  AND U1376 ( .A(n1159), .B(n1160), .Z(n131) );
  NANDN U1377 ( .A(B[40]), .B(n1161), .Z(n1160) );
  NANDN U1378 ( .A(A[40]), .B(n133), .Z(n1161) );
  NANDN U1379 ( .A(n133), .B(A[40]), .Z(n1159) );
  AND U1380 ( .A(n1162), .B(n1163), .Z(n133) );
  NANDN U1381 ( .A(B[39]), .B(n1164), .Z(n1163) );
  NANDN U1382 ( .A(A[39]), .B(n137), .Z(n1164) );
  NANDN U1383 ( .A(n137), .B(A[39]), .Z(n1162) );
  AND U1384 ( .A(n1165), .B(n1166), .Z(n137) );
  NANDN U1385 ( .A(B[38]), .B(n1167), .Z(n1166) );
  NANDN U1386 ( .A(A[38]), .B(n139), .Z(n1167) );
  NANDN U1387 ( .A(n139), .B(A[38]), .Z(n1165) );
  AND U1388 ( .A(n1168), .B(n1169), .Z(n139) );
  NANDN U1389 ( .A(B[37]), .B(n1170), .Z(n1169) );
  NANDN U1390 ( .A(A[37]), .B(n141), .Z(n1170) );
  NANDN U1391 ( .A(n141), .B(A[37]), .Z(n1168) );
  AND U1392 ( .A(n1171), .B(n1172), .Z(n141) );
  NANDN U1393 ( .A(B[36]), .B(n1173), .Z(n1172) );
  NANDN U1394 ( .A(A[36]), .B(n143), .Z(n1173) );
  NANDN U1395 ( .A(n143), .B(A[36]), .Z(n1171) );
  AND U1396 ( .A(n1174), .B(n1175), .Z(n143) );
  NANDN U1397 ( .A(B[35]), .B(n1176), .Z(n1175) );
  NANDN U1398 ( .A(A[35]), .B(n145), .Z(n1176) );
  NANDN U1399 ( .A(n145), .B(A[35]), .Z(n1174) );
  AND U1400 ( .A(n1177), .B(n1178), .Z(n145) );
  NANDN U1401 ( .A(B[34]), .B(n1179), .Z(n1178) );
  NANDN U1402 ( .A(A[34]), .B(n147), .Z(n1179) );
  NANDN U1403 ( .A(n147), .B(A[34]), .Z(n1177) );
  AND U1404 ( .A(n1180), .B(n1181), .Z(n147) );
  NANDN U1405 ( .A(B[33]), .B(n1182), .Z(n1181) );
  NANDN U1406 ( .A(A[33]), .B(n149), .Z(n1182) );
  NANDN U1407 ( .A(n149), .B(A[33]), .Z(n1180) );
  AND U1408 ( .A(n1183), .B(n1184), .Z(n149) );
  NANDN U1409 ( .A(B[32]), .B(n1185), .Z(n1184) );
  NANDN U1410 ( .A(A[32]), .B(n151), .Z(n1185) );
  NANDN U1411 ( .A(n151), .B(A[32]), .Z(n1183) );
  AND U1412 ( .A(n1186), .B(n1187), .Z(n151) );
  NANDN U1413 ( .A(B[31]), .B(n1188), .Z(n1187) );
  NANDN U1414 ( .A(A[31]), .B(n153), .Z(n1188) );
  NANDN U1415 ( .A(n153), .B(A[31]), .Z(n1186) );
  AND U1416 ( .A(n1189), .B(n1190), .Z(n153) );
  NANDN U1417 ( .A(B[30]), .B(n1191), .Z(n1190) );
  NANDN U1418 ( .A(A[30]), .B(n155), .Z(n1191) );
  NANDN U1419 ( .A(n155), .B(A[30]), .Z(n1189) );
  AND U1420 ( .A(n1192), .B(n1193), .Z(n155) );
  NANDN U1421 ( .A(B[29]), .B(n1194), .Z(n1193) );
  NANDN U1422 ( .A(A[29]), .B(n159), .Z(n1194) );
  NANDN U1423 ( .A(n159), .B(A[29]), .Z(n1192) );
  AND U1424 ( .A(n1195), .B(n1196), .Z(n159) );
  NANDN U1425 ( .A(B[28]), .B(n1197), .Z(n1196) );
  NANDN U1426 ( .A(A[28]), .B(n161), .Z(n1197) );
  NANDN U1427 ( .A(n161), .B(A[28]), .Z(n1195) );
  AND U1428 ( .A(n1198), .B(n1199), .Z(n161) );
  NANDN U1429 ( .A(B[27]), .B(n1200), .Z(n1199) );
  NANDN U1430 ( .A(A[27]), .B(n163), .Z(n1200) );
  NANDN U1431 ( .A(n163), .B(A[27]), .Z(n1198) );
  AND U1432 ( .A(n1201), .B(n1202), .Z(n163) );
  NANDN U1433 ( .A(B[26]), .B(n1203), .Z(n1202) );
  NANDN U1434 ( .A(A[26]), .B(n165), .Z(n1203) );
  NANDN U1435 ( .A(n165), .B(A[26]), .Z(n1201) );
  AND U1436 ( .A(n1204), .B(n1205), .Z(n165) );
  NANDN U1437 ( .A(B[25]), .B(n1206), .Z(n1205) );
  NANDN U1438 ( .A(A[25]), .B(n167), .Z(n1206) );
  NANDN U1439 ( .A(n167), .B(A[25]), .Z(n1204) );
  AND U1440 ( .A(n1207), .B(n1208), .Z(n167) );
  NANDN U1441 ( .A(B[24]), .B(n1209), .Z(n1208) );
  NANDN U1442 ( .A(A[24]), .B(n205), .Z(n1209) );
  NANDN U1443 ( .A(n205), .B(A[24]), .Z(n1207) );
  AND U1444 ( .A(n1210), .B(n1211), .Z(n205) );
  NANDN U1445 ( .A(B[23]), .B(n1212), .Z(n1211) );
  NANDN U1446 ( .A(A[23]), .B(n257), .Z(n1212) );
  NANDN U1447 ( .A(n257), .B(A[23]), .Z(n1210) );
  AND U1448 ( .A(n1213), .B(n1214), .Z(n257) );
  NANDN U1449 ( .A(B[22]), .B(n1215), .Z(n1214) );
  NANDN U1450 ( .A(A[22]), .B(n309), .Z(n1215) );
  NANDN U1451 ( .A(n309), .B(A[22]), .Z(n1213) );
  AND U1452 ( .A(n1216), .B(n1217), .Z(n309) );
  NANDN U1453 ( .A(B[21]), .B(n1218), .Z(n1217) );
  NANDN U1454 ( .A(A[21]), .B(n361), .Z(n1218) );
  NANDN U1455 ( .A(n361), .B(A[21]), .Z(n1216) );
  AND U1456 ( .A(n1219), .B(n1220), .Z(n361) );
  NANDN U1457 ( .A(B[20]), .B(n1221), .Z(n1220) );
  NANDN U1458 ( .A(A[20]), .B(n413), .Z(n1221) );
  NANDN U1459 ( .A(n413), .B(A[20]), .Z(n1219) );
  AND U1460 ( .A(n1222), .B(n1223), .Z(n413) );
  NANDN U1461 ( .A(B[19]), .B(n1224), .Z(n1223) );
  NANDN U1462 ( .A(A[19]), .B(n466), .Z(n1224) );
  NANDN U1463 ( .A(n466), .B(A[19]), .Z(n1222) );
  AND U1464 ( .A(n1225), .B(n1226), .Z(n466) );
  NANDN U1465 ( .A(B[18]), .B(n1227), .Z(n1226) );
  NANDN U1466 ( .A(A[18]), .B(n518), .Z(n1227) );
  NANDN U1467 ( .A(n518), .B(A[18]), .Z(n1225) );
  AND U1468 ( .A(n1228), .B(n1229), .Z(n518) );
  NANDN U1469 ( .A(B[17]), .B(n1230), .Z(n1229) );
  NANDN U1470 ( .A(A[17]), .B(n570), .Z(n1230) );
  NANDN U1471 ( .A(n570), .B(A[17]), .Z(n1228) );
  AND U1472 ( .A(n1231), .B(n1232), .Z(n570) );
  NANDN U1473 ( .A(B[16]), .B(n1233), .Z(n1232) );
  NANDN U1474 ( .A(A[16]), .B(n622), .Z(n1233) );
  NANDN U1475 ( .A(n622), .B(A[16]), .Z(n1231) );
  AND U1476 ( .A(n1234), .B(n1235), .Z(n622) );
  NANDN U1477 ( .A(B[15]), .B(n1236), .Z(n1235) );
  NANDN U1478 ( .A(A[15]), .B(n674), .Z(n1236) );
  NANDN U1479 ( .A(n674), .B(A[15]), .Z(n1234) );
  AND U1480 ( .A(n1237), .B(n1238), .Z(n674) );
  NANDN U1481 ( .A(B[14]), .B(n1239), .Z(n1238) );
  NANDN U1482 ( .A(A[14]), .B(n726), .Z(n1239) );
  NANDN U1483 ( .A(n726), .B(A[14]), .Z(n1237) );
  AND U1484 ( .A(n1240), .B(n1241), .Z(n726) );
  NANDN U1485 ( .A(B[13]), .B(n1242), .Z(n1241) );
  NANDN U1486 ( .A(A[13]), .B(n778), .Z(n1242) );
  NANDN U1487 ( .A(n778), .B(A[13]), .Z(n1240) );
  AND U1488 ( .A(n1243), .B(n1244), .Z(n778) );
  NANDN U1489 ( .A(B[12]), .B(n1245), .Z(n1244) );
  NANDN U1490 ( .A(A[12]), .B(n830), .Z(n1245) );
  NANDN U1491 ( .A(n830), .B(A[12]), .Z(n1243) );
  AND U1492 ( .A(n1246), .B(n1247), .Z(n830) );
  NANDN U1493 ( .A(B[11]), .B(n1248), .Z(n1247) );
  NANDN U1494 ( .A(A[11]), .B(n882), .Z(n1248) );
  NANDN U1495 ( .A(n882), .B(A[11]), .Z(n1246) );
  AND U1496 ( .A(n1249), .B(n1250), .Z(n882) );
  NANDN U1497 ( .A(B[10]), .B(n1251), .Z(n1250) );
  NANDN U1498 ( .A(A[10]), .B(n934), .Z(n1251) );
  NANDN U1499 ( .A(n934), .B(A[10]), .Z(n1249) );
  AND U1500 ( .A(n1252), .B(n1253), .Z(n934) );
  NANDN U1501 ( .A(B[9]), .B(n1254), .Z(n1253) );
  OR U1502 ( .A(n3), .B(A[9]), .Z(n1254) );
  NAND U1503 ( .A(A[9]), .B(n3), .Z(n1252) );
  NAND U1504 ( .A(n1255), .B(n1256), .Z(n3) );
  NANDN U1505 ( .A(B[8]), .B(n1257), .Z(n1256) );
  NANDN U1506 ( .A(A[8]), .B(n25), .Z(n1257) );
  NANDN U1507 ( .A(n25), .B(A[8]), .Z(n1255) );
  AND U1508 ( .A(n1258), .B(n1259), .Z(n25) );
  NANDN U1509 ( .A(B[7]), .B(n1260), .Z(n1259) );
  NANDN U1510 ( .A(A[7]), .B(n47), .Z(n1260) );
  NANDN U1511 ( .A(n47), .B(A[7]), .Z(n1258) );
  AND U1512 ( .A(n1261), .B(n1262), .Z(n47) );
  NANDN U1513 ( .A(B[6]), .B(n1263), .Z(n1262) );
  NANDN U1514 ( .A(A[6]), .B(n69), .Z(n1263) );
  NANDN U1515 ( .A(n69), .B(A[6]), .Z(n1261) );
  AND U1516 ( .A(n1264), .B(n1265), .Z(n69) );
  NANDN U1517 ( .A(B[5]), .B(n1266), .Z(n1265) );
  NANDN U1518 ( .A(A[5]), .B(n91), .Z(n1266) );
  NANDN U1519 ( .A(n91), .B(A[5]), .Z(n1264) );
  AND U1520 ( .A(n1267), .B(n1268), .Z(n91) );
  NANDN U1521 ( .A(B[4]), .B(n1269), .Z(n1268) );
  NANDN U1522 ( .A(A[4]), .B(n113), .Z(n1269) );
  NANDN U1523 ( .A(n113), .B(A[4]), .Z(n1267) );
  AND U1524 ( .A(n1270), .B(n1271), .Z(n113) );
  NANDN U1525 ( .A(B[3]), .B(n1272), .Z(n1271) );
  NANDN U1526 ( .A(A[3]), .B(n135), .Z(n1272) );
  NANDN U1527 ( .A(n135), .B(A[3]), .Z(n1270) );
  AND U1528 ( .A(n1273), .B(n1274), .Z(n135) );
  NANDN U1529 ( .A(B[2]), .B(n1275), .Z(n1274) );
  NANDN U1530 ( .A(A[2]), .B(n157), .Z(n1275) );
  NANDN U1531 ( .A(n157), .B(A[2]), .Z(n1273) );
  AND U1532 ( .A(n1276), .B(n1277), .Z(n157) );
  NANDN U1533 ( .A(B[1]), .B(n1278), .Z(n1277) );
  NAND U1534 ( .A(n2), .B(n1), .Z(n1278) );
  NAND U1535 ( .A(A[1]), .B(n1279), .Z(n1276) );
  NAND U1536 ( .A(n1279), .B(n1280), .Z(DIFF[0]) );
  NANDN U1537 ( .A(B[0]), .B(A[0]), .Z(n1280) );
  NANDN U1538 ( .A(A[0]), .B(B[0]), .Z(n1279) );
endmodule


module modmult_step_N256_4_DW01_cmp2_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [257:0] A;
  input [257:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;

  NAND U1 ( .A(n1), .B(n2), .Z(LT_LE) );
  NOR U2 ( .A(B[257]), .B(B[256]), .Z(n2) );
  AND U3 ( .A(n3), .B(n4), .Z(n1) );
  NAND U4 ( .A(n5), .B(n6), .Z(n4) );
  NANDN U5 ( .A(B[255]), .B(A[255]), .Z(n6) );
  NAND U6 ( .A(n7), .B(n8), .Z(n5) );
  NANDN U7 ( .A(A[254]), .B(B[254]), .Z(n8) );
  NAND U8 ( .A(n9), .B(n10), .Z(n7) );
  NANDN U9 ( .A(B[254]), .B(A[254]), .Z(n10) );
  AND U10 ( .A(n11), .B(n12), .Z(n9) );
  NAND U11 ( .A(n13), .B(n14), .Z(n12) );
  NANDN U12 ( .A(A[253]), .B(B[253]), .Z(n14) );
  AND U13 ( .A(n15), .B(n16), .Z(n13) );
  NANDN U14 ( .A(A[252]), .B(B[252]), .Z(n16) );
  NAND U15 ( .A(n17), .B(n18), .Z(n15) );
  NANDN U16 ( .A(B[252]), .B(A[252]), .Z(n18) );
  AND U17 ( .A(n19), .B(n20), .Z(n17) );
  NAND U18 ( .A(n21), .B(n22), .Z(n20) );
  NANDN U19 ( .A(A[251]), .B(B[251]), .Z(n22) );
  AND U20 ( .A(n23), .B(n24), .Z(n21) );
  NANDN U21 ( .A(A[250]), .B(B[250]), .Z(n24) );
  NAND U22 ( .A(n25), .B(n26), .Z(n23) );
  NANDN U23 ( .A(B[250]), .B(A[250]), .Z(n26) );
  AND U24 ( .A(n27), .B(n28), .Z(n25) );
  NAND U25 ( .A(n29), .B(n30), .Z(n28) );
  NANDN U26 ( .A(A[249]), .B(B[249]), .Z(n30) );
  AND U27 ( .A(n31), .B(n32), .Z(n29) );
  NANDN U28 ( .A(A[248]), .B(B[248]), .Z(n32) );
  NAND U29 ( .A(n33), .B(n34), .Z(n31) );
  NANDN U30 ( .A(B[248]), .B(A[248]), .Z(n34) );
  AND U31 ( .A(n35), .B(n36), .Z(n33) );
  NAND U32 ( .A(n37), .B(n38), .Z(n36) );
  NANDN U33 ( .A(A[247]), .B(B[247]), .Z(n38) );
  AND U34 ( .A(n39), .B(n40), .Z(n37) );
  NANDN U35 ( .A(A[246]), .B(B[246]), .Z(n40) );
  NAND U36 ( .A(n41), .B(n42), .Z(n39) );
  NANDN U37 ( .A(B[246]), .B(A[246]), .Z(n42) );
  AND U38 ( .A(n43), .B(n44), .Z(n41) );
  NAND U39 ( .A(n45), .B(n46), .Z(n44) );
  NANDN U40 ( .A(A[245]), .B(B[245]), .Z(n46) );
  AND U41 ( .A(n47), .B(n48), .Z(n45) );
  NANDN U42 ( .A(A[244]), .B(B[244]), .Z(n48) );
  NAND U43 ( .A(n49), .B(n50), .Z(n47) );
  NANDN U44 ( .A(B[244]), .B(A[244]), .Z(n50) );
  AND U45 ( .A(n51), .B(n52), .Z(n49) );
  NAND U46 ( .A(n53), .B(n54), .Z(n52) );
  NANDN U47 ( .A(A[243]), .B(B[243]), .Z(n54) );
  AND U48 ( .A(n55), .B(n56), .Z(n53) );
  NANDN U49 ( .A(A[242]), .B(B[242]), .Z(n56) );
  NAND U50 ( .A(n57), .B(n58), .Z(n55) );
  NANDN U51 ( .A(B[242]), .B(A[242]), .Z(n58) );
  AND U52 ( .A(n59), .B(n60), .Z(n57) );
  NAND U53 ( .A(n61), .B(n62), .Z(n60) );
  NANDN U54 ( .A(A[241]), .B(B[241]), .Z(n62) );
  AND U55 ( .A(n63), .B(n64), .Z(n61) );
  NANDN U56 ( .A(A[240]), .B(B[240]), .Z(n64) );
  NAND U57 ( .A(n65), .B(n66), .Z(n63) );
  NANDN U58 ( .A(B[240]), .B(A[240]), .Z(n66) );
  AND U59 ( .A(n67), .B(n68), .Z(n65) );
  NAND U60 ( .A(n69), .B(n70), .Z(n68) );
  NANDN U61 ( .A(A[239]), .B(B[239]), .Z(n70) );
  AND U62 ( .A(n71), .B(n72), .Z(n69) );
  NANDN U63 ( .A(A[238]), .B(B[238]), .Z(n72) );
  NAND U64 ( .A(n73), .B(n74), .Z(n71) );
  NANDN U65 ( .A(B[238]), .B(A[238]), .Z(n74) );
  AND U66 ( .A(n75), .B(n76), .Z(n73) );
  NAND U67 ( .A(n77), .B(n78), .Z(n76) );
  NANDN U68 ( .A(A[237]), .B(B[237]), .Z(n78) );
  AND U69 ( .A(n79), .B(n80), .Z(n77) );
  NANDN U70 ( .A(A[236]), .B(B[236]), .Z(n80) );
  NAND U71 ( .A(n81), .B(n82), .Z(n79) );
  NANDN U72 ( .A(B[236]), .B(A[236]), .Z(n82) );
  AND U73 ( .A(n83), .B(n84), .Z(n81) );
  NAND U74 ( .A(n85), .B(n86), .Z(n84) );
  NANDN U75 ( .A(A[235]), .B(B[235]), .Z(n86) );
  AND U76 ( .A(n87), .B(n88), .Z(n85) );
  NANDN U77 ( .A(A[234]), .B(B[234]), .Z(n88) );
  NAND U78 ( .A(n89), .B(n90), .Z(n87) );
  NANDN U79 ( .A(B[234]), .B(A[234]), .Z(n90) );
  AND U80 ( .A(n91), .B(n92), .Z(n89) );
  NAND U81 ( .A(n93), .B(n94), .Z(n92) );
  NANDN U82 ( .A(A[233]), .B(B[233]), .Z(n94) );
  AND U83 ( .A(n95), .B(n96), .Z(n93) );
  NANDN U84 ( .A(A[232]), .B(B[232]), .Z(n96) );
  NAND U85 ( .A(n97), .B(n98), .Z(n95) );
  NANDN U86 ( .A(B[232]), .B(A[232]), .Z(n98) );
  AND U87 ( .A(n99), .B(n100), .Z(n97) );
  NAND U88 ( .A(n101), .B(n102), .Z(n100) );
  NANDN U89 ( .A(A[231]), .B(B[231]), .Z(n102) );
  AND U90 ( .A(n103), .B(n104), .Z(n101) );
  NANDN U91 ( .A(A[230]), .B(B[230]), .Z(n104) );
  NAND U92 ( .A(n105), .B(n106), .Z(n103) );
  NANDN U93 ( .A(B[230]), .B(A[230]), .Z(n106) );
  AND U94 ( .A(n107), .B(n108), .Z(n105) );
  NAND U95 ( .A(n109), .B(n110), .Z(n108) );
  NANDN U96 ( .A(A[229]), .B(B[229]), .Z(n110) );
  AND U97 ( .A(n111), .B(n112), .Z(n109) );
  NANDN U98 ( .A(A[228]), .B(B[228]), .Z(n112) );
  NAND U99 ( .A(n113), .B(n114), .Z(n111) );
  NANDN U100 ( .A(B[228]), .B(A[228]), .Z(n114) );
  AND U101 ( .A(n115), .B(n116), .Z(n113) );
  NAND U102 ( .A(n117), .B(n118), .Z(n116) );
  NANDN U103 ( .A(A[227]), .B(B[227]), .Z(n118) );
  AND U104 ( .A(n119), .B(n120), .Z(n117) );
  NANDN U105 ( .A(A[226]), .B(B[226]), .Z(n120) );
  NAND U106 ( .A(n121), .B(n122), .Z(n119) );
  NANDN U107 ( .A(B[226]), .B(A[226]), .Z(n122) );
  AND U108 ( .A(n123), .B(n124), .Z(n121) );
  NAND U109 ( .A(n125), .B(n126), .Z(n124) );
  NANDN U110 ( .A(A[225]), .B(B[225]), .Z(n126) );
  AND U111 ( .A(n127), .B(n128), .Z(n125) );
  NANDN U112 ( .A(A[224]), .B(B[224]), .Z(n128) );
  NAND U113 ( .A(n129), .B(n130), .Z(n127) );
  NANDN U114 ( .A(B[224]), .B(A[224]), .Z(n130) );
  AND U115 ( .A(n131), .B(n132), .Z(n129) );
  NAND U116 ( .A(n133), .B(n134), .Z(n132) );
  NANDN U117 ( .A(A[223]), .B(B[223]), .Z(n134) );
  AND U118 ( .A(n135), .B(n136), .Z(n133) );
  NANDN U119 ( .A(A[222]), .B(B[222]), .Z(n136) );
  NAND U120 ( .A(n137), .B(n138), .Z(n135) );
  NANDN U121 ( .A(B[222]), .B(A[222]), .Z(n138) );
  AND U122 ( .A(n139), .B(n140), .Z(n137) );
  NAND U123 ( .A(n141), .B(n142), .Z(n140) );
  NANDN U124 ( .A(A[221]), .B(B[221]), .Z(n142) );
  AND U125 ( .A(n143), .B(n144), .Z(n141) );
  NANDN U126 ( .A(A[220]), .B(B[220]), .Z(n144) );
  NAND U127 ( .A(n145), .B(n146), .Z(n143) );
  NANDN U128 ( .A(B[220]), .B(A[220]), .Z(n146) );
  AND U129 ( .A(n147), .B(n148), .Z(n145) );
  NAND U130 ( .A(n149), .B(n150), .Z(n148) );
  NANDN U131 ( .A(A[219]), .B(B[219]), .Z(n150) );
  AND U132 ( .A(n151), .B(n152), .Z(n149) );
  NANDN U133 ( .A(A[218]), .B(B[218]), .Z(n152) );
  NAND U134 ( .A(n153), .B(n154), .Z(n151) );
  NANDN U135 ( .A(B[218]), .B(A[218]), .Z(n154) );
  AND U136 ( .A(n155), .B(n156), .Z(n153) );
  NAND U137 ( .A(n157), .B(n158), .Z(n156) );
  NANDN U138 ( .A(A[217]), .B(B[217]), .Z(n158) );
  AND U139 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U140 ( .A(A[216]), .B(B[216]), .Z(n160) );
  NAND U141 ( .A(n161), .B(n162), .Z(n159) );
  NANDN U142 ( .A(B[216]), .B(A[216]), .Z(n162) );
  AND U143 ( .A(n163), .B(n164), .Z(n161) );
  NAND U144 ( .A(n165), .B(n166), .Z(n164) );
  NANDN U145 ( .A(A[215]), .B(B[215]), .Z(n166) );
  AND U146 ( .A(n167), .B(n168), .Z(n165) );
  NANDN U147 ( .A(A[214]), .B(B[214]), .Z(n168) );
  NAND U148 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U149 ( .A(B[214]), .B(A[214]), .Z(n170) );
  AND U150 ( .A(n171), .B(n172), .Z(n169) );
  NAND U151 ( .A(n173), .B(n174), .Z(n172) );
  NANDN U152 ( .A(A[213]), .B(B[213]), .Z(n174) );
  AND U153 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U154 ( .A(A[212]), .B(B[212]), .Z(n176) );
  NAND U155 ( .A(n177), .B(n178), .Z(n175) );
  NANDN U156 ( .A(B[212]), .B(A[212]), .Z(n178) );
  AND U157 ( .A(n179), .B(n180), .Z(n177) );
  NAND U158 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U159 ( .A(A[211]), .B(B[211]), .Z(n182) );
  AND U160 ( .A(n183), .B(n184), .Z(n181) );
  NANDN U161 ( .A(A[210]), .B(B[210]), .Z(n184) );
  NAND U162 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U163 ( .A(B[210]), .B(A[210]), .Z(n186) );
  AND U164 ( .A(n187), .B(n188), .Z(n185) );
  NAND U165 ( .A(n189), .B(n190), .Z(n188) );
  NANDN U166 ( .A(A[209]), .B(B[209]), .Z(n190) );
  AND U167 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U168 ( .A(A[208]), .B(B[208]), .Z(n192) );
  NAND U169 ( .A(n193), .B(n194), .Z(n191) );
  NANDN U170 ( .A(B[208]), .B(A[208]), .Z(n194) );
  AND U171 ( .A(n195), .B(n196), .Z(n193) );
  NAND U172 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U173 ( .A(A[207]), .B(B[207]), .Z(n198) );
  AND U174 ( .A(n199), .B(n200), .Z(n197) );
  NANDN U175 ( .A(A[206]), .B(B[206]), .Z(n200) );
  NAND U176 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U177 ( .A(B[206]), .B(A[206]), .Z(n202) );
  AND U178 ( .A(n203), .B(n204), .Z(n201) );
  NAND U179 ( .A(n205), .B(n206), .Z(n204) );
  NANDN U180 ( .A(A[205]), .B(B[205]), .Z(n206) );
  AND U181 ( .A(n207), .B(n208), .Z(n205) );
  NANDN U182 ( .A(A[204]), .B(B[204]), .Z(n208) );
  NAND U183 ( .A(n209), .B(n210), .Z(n207) );
  NANDN U184 ( .A(B[204]), .B(A[204]), .Z(n210) );
  AND U185 ( .A(n211), .B(n212), .Z(n209) );
  NAND U186 ( .A(n213), .B(n214), .Z(n212) );
  NANDN U187 ( .A(A[203]), .B(B[203]), .Z(n214) );
  AND U188 ( .A(n215), .B(n216), .Z(n213) );
  NANDN U189 ( .A(A[202]), .B(B[202]), .Z(n216) );
  NAND U190 ( .A(n217), .B(n218), .Z(n215) );
  NANDN U191 ( .A(B[202]), .B(A[202]), .Z(n218) );
  AND U192 ( .A(n219), .B(n220), .Z(n217) );
  NAND U193 ( .A(n221), .B(n222), .Z(n220) );
  NANDN U194 ( .A(A[201]), .B(B[201]), .Z(n222) );
  AND U195 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U196 ( .A(A[200]), .B(B[200]), .Z(n224) );
  NAND U197 ( .A(n225), .B(n226), .Z(n223) );
  NANDN U198 ( .A(B[200]), .B(A[200]), .Z(n226) );
  AND U199 ( .A(n227), .B(n228), .Z(n225) );
  NAND U200 ( .A(n229), .B(n230), .Z(n228) );
  NANDN U201 ( .A(A[199]), .B(B[199]), .Z(n230) );
  AND U202 ( .A(n231), .B(n232), .Z(n229) );
  NANDN U203 ( .A(A[198]), .B(B[198]), .Z(n232) );
  NAND U204 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U205 ( .A(B[198]), .B(A[198]), .Z(n234) );
  AND U206 ( .A(n235), .B(n236), .Z(n233) );
  NAND U207 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U208 ( .A(A[197]), .B(B[197]), .Z(n238) );
  AND U209 ( .A(n239), .B(n240), .Z(n237) );
  NANDN U210 ( .A(A[196]), .B(B[196]), .Z(n240) );
  NAND U211 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U212 ( .A(B[196]), .B(A[196]), .Z(n242) );
  AND U213 ( .A(n243), .B(n244), .Z(n241) );
  NAND U214 ( .A(n245), .B(n246), .Z(n244) );
  NANDN U215 ( .A(A[195]), .B(B[195]), .Z(n246) );
  AND U216 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U217 ( .A(A[194]), .B(B[194]), .Z(n248) );
  NAND U218 ( .A(n249), .B(n250), .Z(n247) );
  NANDN U219 ( .A(B[194]), .B(A[194]), .Z(n250) );
  AND U220 ( .A(n251), .B(n252), .Z(n249) );
  NAND U221 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U222 ( .A(A[193]), .B(B[193]), .Z(n254) );
  AND U223 ( .A(n255), .B(n256), .Z(n253) );
  NANDN U224 ( .A(A[192]), .B(B[192]), .Z(n256) );
  NAND U225 ( .A(n257), .B(n258), .Z(n255) );
  NANDN U226 ( .A(B[192]), .B(A[192]), .Z(n258) );
  AND U227 ( .A(n259), .B(n260), .Z(n257) );
  NAND U228 ( .A(n261), .B(n262), .Z(n260) );
  NANDN U229 ( .A(A[191]), .B(B[191]), .Z(n262) );
  AND U230 ( .A(n263), .B(n264), .Z(n261) );
  NANDN U231 ( .A(A[190]), .B(B[190]), .Z(n264) );
  NAND U232 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U233 ( .A(B[190]), .B(A[190]), .Z(n266) );
  AND U234 ( .A(n267), .B(n268), .Z(n265) );
  NAND U235 ( .A(n269), .B(n270), .Z(n268) );
  NANDN U236 ( .A(A[189]), .B(B[189]), .Z(n270) );
  AND U237 ( .A(n271), .B(n272), .Z(n269) );
  NANDN U238 ( .A(A[188]), .B(B[188]), .Z(n272) );
  NAND U239 ( .A(n273), .B(n274), .Z(n271) );
  NANDN U240 ( .A(B[188]), .B(A[188]), .Z(n274) );
  AND U241 ( .A(n275), .B(n276), .Z(n273) );
  NAND U242 ( .A(n277), .B(n278), .Z(n276) );
  NANDN U243 ( .A(A[187]), .B(B[187]), .Z(n278) );
  AND U244 ( .A(n279), .B(n280), .Z(n277) );
  NANDN U245 ( .A(A[186]), .B(B[186]), .Z(n280) );
  NAND U246 ( .A(n281), .B(n282), .Z(n279) );
  NANDN U247 ( .A(B[186]), .B(A[186]), .Z(n282) );
  AND U248 ( .A(n283), .B(n284), .Z(n281) );
  NAND U249 ( .A(n285), .B(n286), .Z(n284) );
  NANDN U250 ( .A(A[185]), .B(B[185]), .Z(n286) );
  AND U251 ( .A(n287), .B(n288), .Z(n285) );
  NANDN U252 ( .A(A[184]), .B(B[184]), .Z(n288) );
  NAND U253 ( .A(n289), .B(n290), .Z(n287) );
  NANDN U254 ( .A(B[184]), .B(A[184]), .Z(n290) );
  AND U255 ( .A(n291), .B(n292), .Z(n289) );
  NAND U256 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U257 ( .A(A[183]), .B(B[183]), .Z(n294) );
  AND U258 ( .A(n295), .B(n296), .Z(n293) );
  NANDN U259 ( .A(A[182]), .B(B[182]), .Z(n296) );
  NAND U260 ( .A(n297), .B(n298), .Z(n295) );
  NANDN U261 ( .A(B[182]), .B(A[182]), .Z(n298) );
  AND U262 ( .A(n299), .B(n300), .Z(n297) );
  NAND U263 ( .A(n301), .B(n302), .Z(n300) );
  NANDN U264 ( .A(A[181]), .B(B[181]), .Z(n302) );
  AND U265 ( .A(n303), .B(n304), .Z(n301) );
  NANDN U266 ( .A(A[180]), .B(B[180]), .Z(n304) );
  NAND U267 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U268 ( .A(B[180]), .B(A[180]), .Z(n306) );
  AND U269 ( .A(n307), .B(n308), .Z(n305) );
  NAND U270 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U271 ( .A(A[179]), .B(B[179]), .Z(n310) );
  AND U272 ( .A(n311), .B(n312), .Z(n309) );
  NANDN U273 ( .A(A[178]), .B(B[178]), .Z(n312) );
  NAND U274 ( .A(n313), .B(n314), .Z(n311) );
  NANDN U275 ( .A(B[178]), .B(A[178]), .Z(n314) );
  AND U276 ( .A(n315), .B(n316), .Z(n313) );
  NAND U277 ( .A(n317), .B(n318), .Z(n316) );
  NANDN U278 ( .A(A[177]), .B(B[177]), .Z(n318) );
  AND U279 ( .A(n319), .B(n320), .Z(n317) );
  NANDN U280 ( .A(A[176]), .B(B[176]), .Z(n320) );
  NAND U281 ( .A(n321), .B(n322), .Z(n319) );
  NANDN U282 ( .A(B[176]), .B(A[176]), .Z(n322) );
  AND U283 ( .A(n323), .B(n324), .Z(n321) );
  NAND U284 ( .A(n325), .B(n326), .Z(n324) );
  NANDN U285 ( .A(A[175]), .B(B[175]), .Z(n326) );
  AND U286 ( .A(n327), .B(n328), .Z(n325) );
  NANDN U287 ( .A(A[174]), .B(B[174]), .Z(n328) );
  NAND U288 ( .A(n329), .B(n330), .Z(n327) );
  NANDN U289 ( .A(B[174]), .B(A[174]), .Z(n330) );
  AND U290 ( .A(n331), .B(n332), .Z(n329) );
  NAND U291 ( .A(n333), .B(n334), .Z(n332) );
  NANDN U292 ( .A(A[173]), .B(B[173]), .Z(n334) );
  AND U293 ( .A(n335), .B(n336), .Z(n333) );
  NANDN U294 ( .A(A[172]), .B(B[172]), .Z(n336) );
  NAND U295 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U296 ( .A(B[172]), .B(A[172]), .Z(n338) );
  AND U297 ( .A(n339), .B(n340), .Z(n337) );
  NAND U298 ( .A(n341), .B(n342), .Z(n340) );
  NANDN U299 ( .A(A[171]), .B(B[171]), .Z(n342) );
  AND U300 ( .A(n343), .B(n344), .Z(n341) );
  NANDN U301 ( .A(A[170]), .B(B[170]), .Z(n344) );
  NAND U302 ( .A(n345), .B(n346), .Z(n343) );
  NANDN U303 ( .A(B[170]), .B(A[170]), .Z(n346) );
  AND U304 ( .A(n347), .B(n348), .Z(n345) );
  NAND U305 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U306 ( .A(A[169]), .B(B[169]), .Z(n350) );
  AND U307 ( .A(n351), .B(n352), .Z(n349) );
  NANDN U308 ( .A(A[168]), .B(B[168]), .Z(n352) );
  NAND U309 ( .A(n353), .B(n354), .Z(n351) );
  NANDN U310 ( .A(B[168]), .B(A[168]), .Z(n354) );
  AND U311 ( .A(n355), .B(n356), .Z(n353) );
  NAND U312 ( .A(n357), .B(n358), .Z(n356) );
  NANDN U313 ( .A(A[167]), .B(B[167]), .Z(n358) );
  AND U314 ( .A(n359), .B(n360), .Z(n357) );
  NANDN U315 ( .A(A[166]), .B(B[166]), .Z(n360) );
  NAND U316 ( .A(n361), .B(n362), .Z(n359) );
  NANDN U317 ( .A(B[166]), .B(A[166]), .Z(n362) );
  AND U318 ( .A(n363), .B(n364), .Z(n361) );
  NAND U319 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U320 ( .A(A[165]), .B(B[165]), .Z(n366) );
  AND U321 ( .A(n367), .B(n368), .Z(n365) );
  NANDN U322 ( .A(A[164]), .B(B[164]), .Z(n368) );
  NAND U323 ( .A(n369), .B(n370), .Z(n367) );
  NANDN U324 ( .A(B[164]), .B(A[164]), .Z(n370) );
  AND U325 ( .A(n371), .B(n372), .Z(n369) );
  NAND U326 ( .A(n373), .B(n374), .Z(n372) );
  NANDN U327 ( .A(A[163]), .B(B[163]), .Z(n374) );
  AND U328 ( .A(n375), .B(n376), .Z(n373) );
  NANDN U329 ( .A(A[162]), .B(B[162]), .Z(n376) );
  NAND U330 ( .A(n377), .B(n378), .Z(n375) );
  NANDN U331 ( .A(B[162]), .B(A[162]), .Z(n378) );
  AND U332 ( .A(n379), .B(n380), .Z(n377) );
  NAND U333 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U334 ( .A(A[161]), .B(B[161]), .Z(n382) );
  AND U335 ( .A(n383), .B(n384), .Z(n381) );
  NANDN U336 ( .A(A[160]), .B(B[160]), .Z(n384) );
  NAND U337 ( .A(n385), .B(n386), .Z(n383) );
  NANDN U338 ( .A(B[160]), .B(A[160]), .Z(n386) );
  AND U339 ( .A(n387), .B(n388), .Z(n385) );
  NAND U340 ( .A(n389), .B(n390), .Z(n388) );
  NANDN U341 ( .A(A[159]), .B(B[159]), .Z(n390) );
  AND U342 ( .A(n391), .B(n392), .Z(n389) );
  NANDN U343 ( .A(A[158]), .B(B[158]), .Z(n392) );
  NAND U344 ( .A(n393), .B(n394), .Z(n391) );
  NANDN U345 ( .A(B[158]), .B(A[158]), .Z(n394) );
  AND U346 ( .A(n395), .B(n396), .Z(n393) );
  NAND U347 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U348 ( .A(A[157]), .B(B[157]), .Z(n398) );
  AND U349 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U350 ( .A(A[156]), .B(B[156]), .Z(n400) );
  NAND U351 ( .A(n401), .B(n402), .Z(n399) );
  NANDN U352 ( .A(B[156]), .B(A[156]), .Z(n402) );
  AND U353 ( .A(n403), .B(n404), .Z(n401) );
  NAND U354 ( .A(n405), .B(n406), .Z(n404) );
  NANDN U355 ( .A(A[155]), .B(B[155]), .Z(n406) );
  AND U356 ( .A(n407), .B(n408), .Z(n405) );
  NANDN U357 ( .A(A[154]), .B(B[154]), .Z(n408) );
  NAND U358 ( .A(n409), .B(n410), .Z(n407) );
  NANDN U359 ( .A(B[154]), .B(A[154]), .Z(n410) );
  AND U360 ( .A(n411), .B(n412), .Z(n409) );
  NAND U361 ( .A(n413), .B(n414), .Z(n412) );
  NANDN U362 ( .A(A[153]), .B(B[153]), .Z(n414) );
  AND U363 ( .A(n415), .B(n416), .Z(n413) );
  NANDN U364 ( .A(A[152]), .B(B[152]), .Z(n416) );
  NAND U365 ( .A(n417), .B(n418), .Z(n415) );
  NANDN U366 ( .A(B[152]), .B(A[152]), .Z(n418) );
  AND U367 ( .A(n419), .B(n420), .Z(n417) );
  NAND U368 ( .A(n421), .B(n422), .Z(n420) );
  NANDN U369 ( .A(A[151]), .B(B[151]), .Z(n422) );
  AND U370 ( .A(n423), .B(n424), .Z(n421) );
  NANDN U371 ( .A(A[150]), .B(B[150]), .Z(n424) );
  NAND U372 ( .A(n425), .B(n426), .Z(n423) );
  NANDN U373 ( .A(B[150]), .B(A[150]), .Z(n426) );
  AND U374 ( .A(n427), .B(n428), .Z(n425) );
  NAND U375 ( .A(n429), .B(n430), .Z(n428) );
  NANDN U376 ( .A(A[149]), .B(B[149]), .Z(n430) );
  AND U377 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U378 ( .A(A[148]), .B(B[148]), .Z(n432) );
  NAND U379 ( .A(n433), .B(n434), .Z(n431) );
  NANDN U380 ( .A(B[148]), .B(A[148]), .Z(n434) );
  AND U381 ( .A(n435), .B(n436), .Z(n433) );
  NAND U382 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U383 ( .A(A[147]), .B(B[147]), .Z(n438) );
  AND U384 ( .A(n439), .B(n440), .Z(n437) );
  NANDN U385 ( .A(A[146]), .B(B[146]), .Z(n440) );
  NAND U386 ( .A(n441), .B(n442), .Z(n439) );
  NANDN U387 ( .A(B[146]), .B(A[146]), .Z(n442) );
  AND U388 ( .A(n443), .B(n444), .Z(n441) );
  NAND U389 ( .A(n445), .B(n446), .Z(n444) );
  NANDN U390 ( .A(A[145]), .B(B[145]), .Z(n446) );
  AND U391 ( .A(n447), .B(n448), .Z(n445) );
  NANDN U392 ( .A(A[144]), .B(B[144]), .Z(n448) );
  NAND U393 ( .A(n449), .B(n450), .Z(n447) );
  NANDN U394 ( .A(B[144]), .B(A[144]), .Z(n450) );
  AND U395 ( .A(n451), .B(n452), .Z(n449) );
  NAND U396 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U397 ( .A(A[143]), .B(B[143]), .Z(n454) );
  AND U398 ( .A(n455), .B(n456), .Z(n453) );
  NANDN U399 ( .A(A[142]), .B(B[142]), .Z(n456) );
  NAND U400 ( .A(n457), .B(n458), .Z(n455) );
  NANDN U401 ( .A(B[142]), .B(A[142]), .Z(n458) );
  AND U402 ( .A(n459), .B(n460), .Z(n457) );
  NAND U403 ( .A(n461), .B(n462), .Z(n460) );
  NANDN U404 ( .A(A[141]), .B(B[141]), .Z(n462) );
  AND U405 ( .A(n463), .B(n464), .Z(n461) );
  NANDN U406 ( .A(A[140]), .B(B[140]), .Z(n464) );
  NAND U407 ( .A(n465), .B(n466), .Z(n463) );
  NANDN U408 ( .A(B[140]), .B(A[140]), .Z(n466) );
  AND U409 ( .A(n467), .B(n468), .Z(n465) );
  NAND U410 ( .A(n469), .B(n470), .Z(n468) );
  NANDN U411 ( .A(A[139]), .B(B[139]), .Z(n470) );
  AND U412 ( .A(n471), .B(n472), .Z(n469) );
  NANDN U413 ( .A(A[138]), .B(B[138]), .Z(n472) );
  NAND U414 ( .A(n473), .B(n474), .Z(n471) );
  NANDN U415 ( .A(B[138]), .B(A[138]), .Z(n474) );
  AND U416 ( .A(n475), .B(n476), .Z(n473) );
  NAND U417 ( .A(n477), .B(n478), .Z(n476) );
  NANDN U418 ( .A(A[137]), .B(B[137]), .Z(n478) );
  AND U419 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U420 ( .A(A[136]), .B(B[136]), .Z(n480) );
  NAND U421 ( .A(n481), .B(n482), .Z(n479) );
  NANDN U422 ( .A(B[136]), .B(A[136]), .Z(n482) );
  AND U423 ( .A(n483), .B(n484), .Z(n481) );
  NAND U424 ( .A(n485), .B(n486), .Z(n484) );
  NANDN U425 ( .A(A[135]), .B(B[135]), .Z(n486) );
  AND U426 ( .A(n487), .B(n488), .Z(n485) );
  NANDN U427 ( .A(A[134]), .B(B[134]), .Z(n488) );
  NAND U428 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U429 ( .A(B[134]), .B(A[134]), .Z(n490) );
  AND U430 ( .A(n491), .B(n492), .Z(n489) );
  NAND U431 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U432 ( .A(A[133]), .B(B[133]), .Z(n494) );
  AND U433 ( .A(n495), .B(n496), .Z(n493) );
  NANDN U434 ( .A(A[132]), .B(B[132]), .Z(n496) );
  NAND U435 ( .A(n497), .B(n498), .Z(n495) );
  NANDN U436 ( .A(B[132]), .B(A[132]), .Z(n498) );
  AND U437 ( .A(n499), .B(n500), .Z(n497) );
  NAND U438 ( .A(n501), .B(n502), .Z(n500) );
  NANDN U439 ( .A(A[131]), .B(B[131]), .Z(n502) );
  AND U440 ( .A(n503), .B(n504), .Z(n501) );
  NANDN U441 ( .A(A[130]), .B(B[130]), .Z(n504) );
  NAND U442 ( .A(n505), .B(n506), .Z(n503) );
  NANDN U443 ( .A(B[130]), .B(A[130]), .Z(n506) );
  AND U444 ( .A(n507), .B(n508), .Z(n505) );
  NAND U445 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U446 ( .A(A[129]), .B(B[129]), .Z(n510) );
  AND U447 ( .A(n511), .B(n512), .Z(n509) );
  NANDN U448 ( .A(A[128]), .B(B[128]), .Z(n512) );
  NAND U449 ( .A(n513), .B(n514), .Z(n511) );
  NANDN U450 ( .A(B[128]), .B(A[128]), .Z(n514) );
  AND U451 ( .A(n515), .B(n516), .Z(n513) );
  NAND U452 ( .A(n517), .B(n518), .Z(n516) );
  NANDN U453 ( .A(A[127]), .B(B[127]), .Z(n518) );
  AND U454 ( .A(n519), .B(n520), .Z(n517) );
  NANDN U455 ( .A(A[126]), .B(B[126]), .Z(n520) );
  NAND U456 ( .A(n521), .B(n522), .Z(n519) );
  NANDN U457 ( .A(B[126]), .B(A[126]), .Z(n522) );
  AND U458 ( .A(n523), .B(n524), .Z(n521) );
  NAND U459 ( .A(n525), .B(n526), .Z(n524) );
  NANDN U460 ( .A(A[125]), .B(B[125]), .Z(n526) );
  AND U461 ( .A(n527), .B(n528), .Z(n525) );
  NANDN U462 ( .A(A[124]), .B(B[124]), .Z(n528) );
  NAND U463 ( .A(n529), .B(n530), .Z(n527) );
  NANDN U464 ( .A(B[124]), .B(A[124]), .Z(n530) );
  AND U465 ( .A(n531), .B(n532), .Z(n529) );
  NAND U466 ( .A(n533), .B(n534), .Z(n532) );
  NANDN U467 ( .A(A[123]), .B(B[123]), .Z(n534) );
  AND U468 ( .A(n535), .B(n536), .Z(n533) );
  NANDN U469 ( .A(A[122]), .B(B[122]), .Z(n536) );
  NAND U470 ( .A(n537), .B(n538), .Z(n535) );
  NANDN U471 ( .A(B[122]), .B(A[122]), .Z(n538) );
  AND U472 ( .A(n539), .B(n540), .Z(n537) );
  NAND U473 ( .A(n541), .B(n542), .Z(n540) );
  NANDN U474 ( .A(A[121]), .B(B[121]), .Z(n542) );
  AND U475 ( .A(n543), .B(n544), .Z(n541) );
  NANDN U476 ( .A(A[120]), .B(B[120]), .Z(n544) );
  NAND U477 ( .A(n545), .B(n546), .Z(n543) );
  NANDN U478 ( .A(B[120]), .B(A[120]), .Z(n546) );
  AND U479 ( .A(n547), .B(n548), .Z(n545) );
  NAND U480 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U481 ( .A(A[119]), .B(B[119]), .Z(n550) );
  AND U482 ( .A(n551), .B(n552), .Z(n549) );
  NANDN U483 ( .A(A[118]), .B(B[118]), .Z(n552) );
  NAND U484 ( .A(n553), .B(n554), .Z(n551) );
  NANDN U485 ( .A(B[118]), .B(A[118]), .Z(n554) );
  AND U486 ( .A(n555), .B(n556), .Z(n553) );
  NAND U487 ( .A(n557), .B(n558), .Z(n556) );
  NANDN U488 ( .A(A[117]), .B(B[117]), .Z(n558) );
  AND U489 ( .A(n559), .B(n560), .Z(n557) );
  NANDN U490 ( .A(A[116]), .B(B[116]), .Z(n560) );
  NAND U491 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U492 ( .A(B[116]), .B(A[116]), .Z(n562) );
  AND U493 ( .A(n563), .B(n564), .Z(n561) );
  NAND U494 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U495 ( .A(A[115]), .B(B[115]), .Z(n566) );
  AND U496 ( .A(n567), .B(n568), .Z(n565) );
  NANDN U497 ( .A(A[114]), .B(B[114]), .Z(n568) );
  NAND U498 ( .A(n569), .B(n570), .Z(n567) );
  NANDN U499 ( .A(B[114]), .B(A[114]), .Z(n570) );
  AND U500 ( .A(n571), .B(n572), .Z(n569) );
  NAND U501 ( .A(n573), .B(n574), .Z(n572) );
  NANDN U502 ( .A(A[113]), .B(B[113]), .Z(n574) );
  AND U503 ( .A(n575), .B(n576), .Z(n573) );
  NANDN U504 ( .A(A[112]), .B(B[112]), .Z(n576) );
  NAND U505 ( .A(n577), .B(n578), .Z(n575) );
  NANDN U506 ( .A(B[112]), .B(A[112]), .Z(n578) );
  AND U507 ( .A(n579), .B(n580), .Z(n577) );
  NAND U508 ( .A(n581), .B(n582), .Z(n580) );
  NANDN U509 ( .A(A[111]), .B(B[111]), .Z(n582) );
  AND U510 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U511 ( .A(A[110]), .B(B[110]), .Z(n584) );
  NAND U512 ( .A(n585), .B(n586), .Z(n583) );
  NANDN U513 ( .A(B[110]), .B(A[110]), .Z(n586) );
  AND U514 ( .A(n587), .B(n588), .Z(n585) );
  NAND U515 ( .A(n589), .B(n590), .Z(n588) );
  NANDN U516 ( .A(A[109]), .B(B[109]), .Z(n590) );
  AND U517 ( .A(n591), .B(n592), .Z(n589) );
  NANDN U518 ( .A(A[108]), .B(B[108]), .Z(n592) );
  NAND U519 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U520 ( .A(B[108]), .B(A[108]), .Z(n594) );
  AND U521 ( .A(n595), .B(n596), .Z(n593) );
  NAND U522 ( .A(n597), .B(n598), .Z(n596) );
  NANDN U523 ( .A(A[107]), .B(B[107]), .Z(n598) );
  AND U524 ( .A(n599), .B(n600), .Z(n597) );
  NANDN U525 ( .A(A[106]), .B(B[106]), .Z(n600) );
  NAND U526 ( .A(n601), .B(n602), .Z(n599) );
  NANDN U527 ( .A(B[106]), .B(A[106]), .Z(n602) );
  AND U528 ( .A(n603), .B(n604), .Z(n601) );
  NAND U529 ( .A(n605), .B(n606), .Z(n604) );
  NANDN U530 ( .A(A[105]), .B(B[105]), .Z(n606) );
  AND U531 ( .A(n607), .B(n608), .Z(n605) );
  NANDN U532 ( .A(A[104]), .B(B[104]), .Z(n608) );
  NAND U533 ( .A(n609), .B(n610), .Z(n607) );
  NANDN U534 ( .A(B[104]), .B(A[104]), .Z(n610) );
  AND U535 ( .A(n611), .B(n612), .Z(n609) );
  NAND U536 ( .A(n613), .B(n614), .Z(n612) );
  NANDN U537 ( .A(A[103]), .B(B[103]), .Z(n614) );
  AND U538 ( .A(n615), .B(n616), .Z(n613) );
  NANDN U539 ( .A(A[102]), .B(B[102]), .Z(n616) );
  NAND U540 ( .A(n617), .B(n618), .Z(n615) );
  NANDN U541 ( .A(B[102]), .B(A[102]), .Z(n618) );
  AND U542 ( .A(n619), .B(n620), .Z(n617) );
  NAND U543 ( .A(n621), .B(n622), .Z(n620) );
  NANDN U544 ( .A(A[101]), .B(B[101]), .Z(n622) );
  AND U545 ( .A(n623), .B(n624), .Z(n621) );
  NANDN U546 ( .A(A[100]), .B(B[100]), .Z(n624) );
  NAND U547 ( .A(n625), .B(n626), .Z(n623) );
  NANDN U548 ( .A(B[99]), .B(A[99]), .Z(n626) );
  AND U549 ( .A(n627), .B(n628), .Z(n625) );
  NAND U550 ( .A(n629), .B(n630), .Z(n628) );
  NANDN U551 ( .A(A[99]), .B(B[99]), .Z(n630) );
  AND U552 ( .A(n631), .B(n632), .Z(n629) );
  NANDN U553 ( .A(A[98]), .B(B[98]), .Z(n632) );
  NAND U554 ( .A(n633), .B(n634), .Z(n631) );
  NANDN U555 ( .A(B[98]), .B(A[98]), .Z(n634) );
  AND U556 ( .A(n635), .B(n636), .Z(n633) );
  NAND U557 ( .A(n637), .B(n638), .Z(n636) );
  NANDN U558 ( .A(A[97]), .B(B[97]), .Z(n638) );
  AND U559 ( .A(n639), .B(n640), .Z(n637) );
  NANDN U560 ( .A(A[96]), .B(B[96]), .Z(n640) );
  NAND U561 ( .A(n641), .B(n642), .Z(n639) );
  NANDN U562 ( .A(B[96]), .B(A[96]), .Z(n642) );
  AND U563 ( .A(n643), .B(n644), .Z(n641) );
  NAND U564 ( .A(n645), .B(n646), .Z(n644) );
  NANDN U565 ( .A(A[95]), .B(B[95]), .Z(n646) );
  AND U566 ( .A(n647), .B(n648), .Z(n645) );
  NANDN U567 ( .A(A[94]), .B(B[94]), .Z(n648) );
  NAND U568 ( .A(n649), .B(n650), .Z(n647) );
  NANDN U569 ( .A(B[94]), .B(A[94]), .Z(n650) );
  AND U570 ( .A(n651), .B(n652), .Z(n649) );
  NAND U571 ( .A(n653), .B(n654), .Z(n652) );
  NANDN U572 ( .A(A[93]), .B(B[93]), .Z(n654) );
  AND U573 ( .A(n655), .B(n656), .Z(n653) );
  NANDN U574 ( .A(A[92]), .B(B[92]), .Z(n656) );
  NAND U575 ( .A(n657), .B(n658), .Z(n655) );
  NANDN U576 ( .A(B[92]), .B(A[92]), .Z(n658) );
  AND U577 ( .A(n659), .B(n660), .Z(n657) );
  NAND U578 ( .A(n661), .B(n662), .Z(n660) );
  NANDN U579 ( .A(A[91]), .B(B[91]), .Z(n662) );
  AND U580 ( .A(n663), .B(n664), .Z(n661) );
  NANDN U581 ( .A(A[90]), .B(B[90]), .Z(n664) );
  NAND U582 ( .A(n665), .B(n666), .Z(n663) );
  NANDN U583 ( .A(B[90]), .B(A[90]), .Z(n666) );
  AND U584 ( .A(n667), .B(n668), .Z(n665) );
  NAND U585 ( .A(n669), .B(n670), .Z(n668) );
  NANDN U586 ( .A(A[89]), .B(B[89]), .Z(n670) );
  AND U587 ( .A(n671), .B(n672), .Z(n669) );
  NANDN U588 ( .A(A[88]), .B(B[88]), .Z(n672) );
  NAND U589 ( .A(n673), .B(n674), .Z(n671) );
  NANDN U590 ( .A(B[88]), .B(A[88]), .Z(n674) );
  AND U591 ( .A(n675), .B(n676), .Z(n673) );
  NAND U592 ( .A(n677), .B(n678), .Z(n676) );
  NANDN U593 ( .A(A[87]), .B(B[87]), .Z(n678) );
  AND U594 ( .A(n679), .B(n680), .Z(n677) );
  NANDN U595 ( .A(A[86]), .B(B[86]), .Z(n680) );
  NAND U596 ( .A(n681), .B(n682), .Z(n679) );
  NANDN U597 ( .A(B[86]), .B(A[86]), .Z(n682) );
  AND U598 ( .A(n683), .B(n684), .Z(n681) );
  NAND U599 ( .A(n685), .B(n686), .Z(n684) );
  NANDN U600 ( .A(A[85]), .B(B[85]), .Z(n686) );
  AND U601 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U602 ( .A(A[84]), .B(B[84]), .Z(n688) );
  NAND U603 ( .A(n689), .B(n690), .Z(n687) );
  NANDN U604 ( .A(B[84]), .B(A[84]), .Z(n690) );
  AND U605 ( .A(n691), .B(n692), .Z(n689) );
  NAND U606 ( .A(n693), .B(n694), .Z(n692) );
  NANDN U607 ( .A(A[83]), .B(B[83]), .Z(n694) );
  AND U608 ( .A(n695), .B(n696), .Z(n693) );
  NANDN U609 ( .A(A[82]), .B(B[82]), .Z(n696) );
  NAND U610 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U611 ( .A(B[82]), .B(A[82]), .Z(n698) );
  AND U612 ( .A(n699), .B(n700), .Z(n697) );
  NAND U613 ( .A(n701), .B(n702), .Z(n700) );
  NANDN U614 ( .A(A[81]), .B(B[81]), .Z(n702) );
  AND U615 ( .A(n703), .B(n704), .Z(n701) );
  NANDN U616 ( .A(A[80]), .B(B[80]), .Z(n704) );
  NAND U617 ( .A(n705), .B(n706), .Z(n703) );
  NANDN U618 ( .A(B[80]), .B(A[80]), .Z(n706) );
  AND U619 ( .A(n707), .B(n708), .Z(n705) );
  NAND U620 ( .A(n709), .B(n710), .Z(n708) );
  NANDN U621 ( .A(A[79]), .B(B[79]), .Z(n710) );
  AND U622 ( .A(n711), .B(n712), .Z(n709) );
  NANDN U623 ( .A(A[78]), .B(B[78]), .Z(n712) );
  NAND U624 ( .A(n713), .B(n714), .Z(n711) );
  NANDN U625 ( .A(B[78]), .B(A[78]), .Z(n714) );
  AND U626 ( .A(n715), .B(n716), .Z(n713) );
  NAND U627 ( .A(n717), .B(n718), .Z(n716) );
  NANDN U628 ( .A(A[77]), .B(B[77]), .Z(n718) );
  AND U629 ( .A(n719), .B(n720), .Z(n717) );
  NANDN U630 ( .A(A[76]), .B(B[76]), .Z(n720) );
  NAND U631 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U632 ( .A(B[76]), .B(A[76]), .Z(n722) );
  AND U633 ( .A(n723), .B(n724), .Z(n721) );
  NAND U634 ( .A(n725), .B(n726), .Z(n724) );
  NANDN U635 ( .A(A[75]), .B(B[75]), .Z(n726) );
  AND U636 ( .A(n727), .B(n728), .Z(n725) );
  NANDN U637 ( .A(A[74]), .B(B[74]), .Z(n728) );
  NAND U638 ( .A(n729), .B(n730), .Z(n727) );
  NANDN U639 ( .A(B[74]), .B(A[74]), .Z(n730) );
  AND U640 ( .A(n731), .B(n732), .Z(n729) );
  NAND U641 ( .A(n733), .B(n734), .Z(n732) );
  NANDN U642 ( .A(A[73]), .B(B[73]), .Z(n734) );
  AND U643 ( .A(n735), .B(n736), .Z(n733) );
  NANDN U644 ( .A(A[72]), .B(B[72]), .Z(n736) );
  NAND U645 ( .A(n737), .B(n738), .Z(n735) );
  NANDN U646 ( .A(B[72]), .B(A[72]), .Z(n738) );
  AND U647 ( .A(n739), .B(n740), .Z(n737) );
  NAND U648 ( .A(n741), .B(n742), .Z(n740) );
  NANDN U649 ( .A(A[71]), .B(B[71]), .Z(n742) );
  AND U650 ( .A(n743), .B(n744), .Z(n741) );
  NANDN U651 ( .A(A[70]), .B(B[70]), .Z(n744) );
  NAND U652 ( .A(n745), .B(n746), .Z(n743) );
  NANDN U653 ( .A(B[70]), .B(A[70]), .Z(n746) );
  AND U654 ( .A(n747), .B(n748), .Z(n745) );
  NAND U655 ( .A(n749), .B(n750), .Z(n748) );
  NANDN U656 ( .A(A[69]), .B(B[69]), .Z(n750) );
  AND U657 ( .A(n751), .B(n752), .Z(n749) );
  NANDN U658 ( .A(A[68]), .B(B[68]), .Z(n752) );
  NAND U659 ( .A(n753), .B(n754), .Z(n751) );
  NANDN U660 ( .A(B[68]), .B(A[68]), .Z(n754) );
  AND U661 ( .A(n755), .B(n756), .Z(n753) );
  NAND U662 ( .A(n757), .B(n758), .Z(n756) );
  NANDN U663 ( .A(A[67]), .B(B[67]), .Z(n758) );
  AND U664 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U665 ( .A(A[66]), .B(B[66]), .Z(n760) );
  NAND U666 ( .A(n761), .B(n762), .Z(n759) );
  NANDN U667 ( .A(B[66]), .B(A[66]), .Z(n762) );
  AND U668 ( .A(n763), .B(n764), .Z(n761) );
  NAND U669 ( .A(n765), .B(n766), .Z(n764) );
  NANDN U670 ( .A(A[65]), .B(B[65]), .Z(n766) );
  AND U671 ( .A(n767), .B(n768), .Z(n765) );
  NANDN U672 ( .A(A[64]), .B(B[64]), .Z(n768) );
  NAND U673 ( .A(n769), .B(n770), .Z(n767) );
  NANDN U674 ( .A(B[64]), .B(A[64]), .Z(n770) );
  AND U675 ( .A(n771), .B(n772), .Z(n769) );
  NAND U676 ( .A(n773), .B(n774), .Z(n772) );
  NANDN U677 ( .A(A[63]), .B(B[63]), .Z(n774) );
  AND U678 ( .A(n775), .B(n776), .Z(n773) );
  NANDN U679 ( .A(A[62]), .B(B[62]), .Z(n776) );
  NAND U680 ( .A(n777), .B(n778), .Z(n775) );
  NANDN U681 ( .A(B[62]), .B(A[62]), .Z(n778) );
  AND U682 ( .A(n779), .B(n780), .Z(n777) );
  NAND U683 ( .A(n781), .B(n782), .Z(n780) );
  NANDN U684 ( .A(A[61]), .B(B[61]), .Z(n782) );
  AND U685 ( .A(n783), .B(n784), .Z(n781) );
  NANDN U686 ( .A(A[60]), .B(B[60]), .Z(n784) );
  NAND U687 ( .A(n785), .B(n786), .Z(n783) );
  NANDN U688 ( .A(B[60]), .B(A[60]), .Z(n786) );
  AND U689 ( .A(n787), .B(n788), .Z(n785) );
  NAND U690 ( .A(n789), .B(n790), .Z(n788) );
  NANDN U691 ( .A(A[59]), .B(B[59]), .Z(n790) );
  AND U692 ( .A(n791), .B(n792), .Z(n789) );
  NANDN U693 ( .A(A[58]), .B(B[58]), .Z(n792) );
  NAND U694 ( .A(n793), .B(n794), .Z(n791) );
  NANDN U695 ( .A(B[58]), .B(A[58]), .Z(n794) );
  AND U696 ( .A(n795), .B(n796), .Z(n793) );
  NAND U697 ( .A(n797), .B(n798), .Z(n796) );
  NANDN U698 ( .A(A[57]), .B(B[57]), .Z(n798) );
  AND U699 ( .A(n799), .B(n800), .Z(n797) );
  NANDN U700 ( .A(A[56]), .B(B[56]), .Z(n800) );
  NAND U701 ( .A(n801), .B(n802), .Z(n799) );
  NANDN U702 ( .A(B[56]), .B(A[56]), .Z(n802) );
  AND U703 ( .A(n803), .B(n804), .Z(n801) );
  NAND U704 ( .A(n805), .B(n806), .Z(n804) );
  NANDN U705 ( .A(A[55]), .B(B[55]), .Z(n806) );
  AND U706 ( .A(n807), .B(n808), .Z(n805) );
  NANDN U707 ( .A(A[54]), .B(B[54]), .Z(n808) );
  NAND U708 ( .A(n809), .B(n810), .Z(n807) );
  NANDN U709 ( .A(B[54]), .B(A[54]), .Z(n810) );
  AND U710 ( .A(n811), .B(n812), .Z(n809) );
  NAND U711 ( .A(n813), .B(n814), .Z(n812) );
  NANDN U712 ( .A(A[53]), .B(B[53]), .Z(n814) );
  AND U713 ( .A(n815), .B(n816), .Z(n813) );
  NANDN U714 ( .A(A[52]), .B(B[52]), .Z(n816) );
  NAND U715 ( .A(n817), .B(n818), .Z(n815) );
  NANDN U716 ( .A(B[52]), .B(A[52]), .Z(n818) );
  AND U717 ( .A(n819), .B(n820), .Z(n817) );
  NAND U718 ( .A(n821), .B(n822), .Z(n820) );
  NANDN U719 ( .A(A[51]), .B(B[51]), .Z(n822) );
  AND U720 ( .A(n823), .B(n824), .Z(n821) );
  NANDN U721 ( .A(A[50]), .B(B[50]), .Z(n824) );
  NAND U722 ( .A(n825), .B(n826), .Z(n823) );
  NANDN U723 ( .A(B[50]), .B(A[50]), .Z(n826) );
  AND U724 ( .A(n827), .B(n828), .Z(n825) );
  NAND U725 ( .A(n829), .B(n830), .Z(n828) );
  NANDN U726 ( .A(A[49]), .B(B[49]), .Z(n830) );
  AND U727 ( .A(n831), .B(n832), .Z(n829) );
  NANDN U728 ( .A(A[48]), .B(B[48]), .Z(n832) );
  NAND U729 ( .A(n833), .B(n834), .Z(n831) );
  NANDN U730 ( .A(B[48]), .B(A[48]), .Z(n834) );
  AND U731 ( .A(n835), .B(n836), .Z(n833) );
  NAND U732 ( .A(n837), .B(n838), .Z(n836) );
  NANDN U733 ( .A(A[47]), .B(B[47]), .Z(n838) );
  AND U734 ( .A(n839), .B(n840), .Z(n837) );
  NANDN U735 ( .A(A[46]), .B(B[46]), .Z(n840) );
  NAND U736 ( .A(n841), .B(n842), .Z(n839) );
  NANDN U737 ( .A(B[46]), .B(A[46]), .Z(n842) );
  AND U738 ( .A(n843), .B(n844), .Z(n841) );
  NAND U739 ( .A(n845), .B(n846), .Z(n844) );
  NANDN U740 ( .A(A[45]), .B(B[45]), .Z(n846) );
  AND U741 ( .A(n847), .B(n848), .Z(n845) );
  NANDN U742 ( .A(A[44]), .B(B[44]), .Z(n848) );
  NAND U743 ( .A(n849), .B(n850), .Z(n847) );
  NANDN U744 ( .A(B[44]), .B(A[44]), .Z(n850) );
  AND U745 ( .A(n851), .B(n852), .Z(n849) );
  NAND U746 ( .A(n853), .B(n854), .Z(n852) );
  NANDN U747 ( .A(A[43]), .B(B[43]), .Z(n854) );
  AND U748 ( .A(n855), .B(n856), .Z(n853) );
  NANDN U749 ( .A(A[42]), .B(B[42]), .Z(n856) );
  NAND U750 ( .A(n857), .B(n858), .Z(n855) );
  NANDN U751 ( .A(B[42]), .B(A[42]), .Z(n858) );
  AND U752 ( .A(n859), .B(n860), .Z(n857) );
  NAND U753 ( .A(n861), .B(n862), .Z(n860) );
  NANDN U754 ( .A(A[41]), .B(B[41]), .Z(n862) );
  AND U755 ( .A(n863), .B(n864), .Z(n861) );
  NANDN U756 ( .A(A[40]), .B(B[40]), .Z(n864) );
  NAND U757 ( .A(n865), .B(n866), .Z(n863) );
  NANDN U758 ( .A(B[40]), .B(A[40]), .Z(n866) );
  AND U759 ( .A(n867), .B(n868), .Z(n865) );
  NAND U760 ( .A(n869), .B(n870), .Z(n868) );
  NANDN U761 ( .A(A[39]), .B(B[39]), .Z(n870) );
  AND U762 ( .A(n871), .B(n872), .Z(n869) );
  NANDN U763 ( .A(A[38]), .B(B[38]), .Z(n872) );
  NAND U764 ( .A(n873), .B(n874), .Z(n871) );
  NANDN U765 ( .A(B[38]), .B(A[38]), .Z(n874) );
  AND U766 ( .A(n875), .B(n876), .Z(n873) );
  NAND U767 ( .A(n877), .B(n878), .Z(n876) );
  NANDN U768 ( .A(A[37]), .B(B[37]), .Z(n878) );
  AND U769 ( .A(n879), .B(n880), .Z(n877) );
  NANDN U770 ( .A(A[36]), .B(B[36]), .Z(n880) );
  NAND U771 ( .A(n881), .B(n882), .Z(n879) );
  NANDN U772 ( .A(B[36]), .B(A[36]), .Z(n882) );
  AND U773 ( .A(n883), .B(n884), .Z(n881) );
  NAND U774 ( .A(n885), .B(n886), .Z(n884) );
  NANDN U775 ( .A(A[35]), .B(B[35]), .Z(n886) );
  AND U776 ( .A(n887), .B(n888), .Z(n885) );
  NANDN U777 ( .A(A[34]), .B(B[34]), .Z(n888) );
  NAND U778 ( .A(n889), .B(n890), .Z(n887) );
  NANDN U779 ( .A(B[34]), .B(A[34]), .Z(n890) );
  AND U780 ( .A(n891), .B(n892), .Z(n889) );
  NAND U781 ( .A(n893), .B(n894), .Z(n892) );
  NANDN U782 ( .A(A[33]), .B(B[33]), .Z(n894) );
  AND U783 ( .A(n895), .B(n896), .Z(n893) );
  NANDN U784 ( .A(A[32]), .B(B[32]), .Z(n896) );
  NAND U785 ( .A(n897), .B(n898), .Z(n895) );
  NANDN U786 ( .A(B[32]), .B(A[32]), .Z(n898) );
  AND U787 ( .A(n899), .B(n900), .Z(n897) );
  NAND U788 ( .A(n901), .B(n902), .Z(n900) );
  NANDN U789 ( .A(A[31]), .B(B[31]), .Z(n902) );
  AND U790 ( .A(n903), .B(n904), .Z(n901) );
  NANDN U791 ( .A(A[30]), .B(B[30]), .Z(n904) );
  NAND U792 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U793 ( .A(B[30]), .B(A[30]), .Z(n906) );
  AND U794 ( .A(n907), .B(n908), .Z(n905) );
  NAND U795 ( .A(n909), .B(n910), .Z(n908) );
  NANDN U796 ( .A(A[29]), .B(B[29]), .Z(n910) );
  AND U797 ( .A(n911), .B(n912), .Z(n909) );
  NANDN U798 ( .A(A[28]), .B(B[28]), .Z(n912) );
  NAND U799 ( .A(n913), .B(n914), .Z(n911) );
  NANDN U800 ( .A(B[28]), .B(A[28]), .Z(n914) );
  AND U801 ( .A(n915), .B(n916), .Z(n913) );
  NAND U802 ( .A(n917), .B(n918), .Z(n916) );
  NANDN U803 ( .A(A[27]), .B(B[27]), .Z(n918) );
  AND U804 ( .A(n919), .B(n920), .Z(n917) );
  NANDN U805 ( .A(A[26]), .B(B[26]), .Z(n920) );
  NAND U806 ( .A(n921), .B(n922), .Z(n919) );
  NANDN U807 ( .A(B[26]), .B(A[26]), .Z(n922) );
  AND U808 ( .A(n923), .B(n924), .Z(n921) );
  NAND U809 ( .A(n925), .B(n926), .Z(n924) );
  NANDN U810 ( .A(A[25]), .B(B[25]), .Z(n926) );
  AND U811 ( .A(n927), .B(n928), .Z(n925) );
  NANDN U812 ( .A(A[24]), .B(B[24]), .Z(n928) );
  NAND U813 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U814 ( .A(B[24]), .B(A[24]), .Z(n930) );
  AND U815 ( .A(n931), .B(n932), .Z(n929) );
  NAND U816 ( .A(n933), .B(n934), .Z(n932) );
  NANDN U817 ( .A(A[23]), .B(B[23]), .Z(n934) );
  AND U818 ( .A(n935), .B(n936), .Z(n933) );
  NANDN U819 ( .A(A[22]), .B(B[22]), .Z(n936) );
  NAND U820 ( .A(n937), .B(n938), .Z(n935) );
  NANDN U821 ( .A(B[22]), .B(A[22]), .Z(n938) );
  AND U822 ( .A(n939), .B(n940), .Z(n937) );
  NAND U823 ( .A(n941), .B(n942), .Z(n940) );
  NANDN U824 ( .A(A[21]), .B(B[21]), .Z(n942) );
  AND U825 ( .A(n943), .B(n944), .Z(n941) );
  NANDN U826 ( .A(A[20]), .B(B[20]), .Z(n944) );
  NAND U827 ( .A(n945), .B(n946), .Z(n943) );
  NANDN U828 ( .A(B[20]), .B(A[20]), .Z(n946) );
  AND U829 ( .A(n947), .B(n948), .Z(n945) );
  NAND U830 ( .A(n949), .B(n950), .Z(n948) );
  NANDN U831 ( .A(A[19]), .B(B[19]), .Z(n950) );
  AND U832 ( .A(n951), .B(n952), .Z(n949) );
  NANDN U833 ( .A(A[18]), .B(B[18]), .Z(n952) );
  NAND U834 ( .A(n953), .B(n954), .Z(n951) );
  NANDN U835 ( .A(B[18]), .B(A[18]), .Z(n954) );
  AND U836 ( .A(n955), .B(n956), .Z(n953) );
  NAND U837 ( .A(n957), .B(n958), .Z(n956) );
  NANDN U838 ( .A(A[17]), .B(B[17]), .Z(n958) );
  AND U839 ( .A(n959), .B(n960), .Z(n957) );
  NANDN U840 ( .A(A[16]), .B(B[16]), .Z(n960) );
  NAND U841 ( .A(n961), .B(n962), .Z(n959) );
  NANDN U842 ( .A(B[16]), .B(A[16]), .Z(n962) );
  AND U843 ( .A(n963), .B(n964), .Z(n961) );
  NAND U844 ( .A(n965), .B(n966), .Z(n964) );
  NANDN U845 ( .A(A[15]), .B(B[15]), .Z(n966) );
  AND U846 ( .A(n967), .B(n968), .Z(n965) );
  NANDN U847 ( .A(A[14]), .B(B[14]), .Z(n968) );
  NAND U848 ( .A(n969), .B(n970), .Z(n967) );
  NANDN U849 ( .A(B[14]), .B(A[14]), .Z(n970) );
  AND U850 ( .A(n971), .B(n972), .Z(n969) );
  NAND U851 ( .A(n973), .B(n974), .Z(n972) );
  NANDN U852 ( .A(A[13]), .B(B[13]), .Z(n974) );
  AND U853 ( .A(n975), .B(n976), .Z(n973) );
  NANDN U854 ( .A(A[12]), .B(B[12]), .Z(n976) );
  NAND U855 ( .A(n977), .B(n978), .Z(n975) );
  NANDN U856 ( .A(B[12]), .B(A[12]), .Z(n978) );
  AND U857 ( .A(n979), .B(n980), .Z(n977) );
  NAND U858 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U859 ( .A(A[11]), .B(B[11]), .Z(n982) );
  AND U860 ( .A(n983), .B(n984), .Z(n981) );
  NANDN U861 ( .A(A[10]), .B(B[10]), .Z(n984) );
  NAND U862 ( .A(n985), .B(n986), .Z(n983) );
  NANDN U863 ( .A(B[9]), .B(A[9]), .Z(n986) );
  AND U864 ( .A(n987), .B(n988), .Z(n985) );
  NAND U865 ( .A(n989), .B(n990), .Z(n988) );
  NANDN U866 ( .A(A[9]), .B(B[9]), .Z(n990) );
  AND U867 ( .A(n991), .B(n992), .Z(n989) );
  NANDN U868 ( .A(A[8]), .B(B[8]), .Z(n992) );
  NAND U869 ( .A(n993), .B(n994), .Z(n991) );
  NANDN U870 ( .A(B[8]), .B(A[8]), .Z(n994) );
  AND U871 ( .A(n995), .B(n996), .Z(n993) );
  NAND U872 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U873 ( .A(A[7]), .B(B[7]), .Z(n998) );
  AND U874 ( .A(n999), .B(n1000), .Z(n997) );
  NANDN U875 ( .A(A[6]), .B(B[6]), .Z(n1000) );
  NAND U876 ( .A(n1001), .B(n1002), .Z(n999) );
  NANDN U877 ( .A(B[6]), .B(A[6]), .Z(n1002) );
  AND U878 ( .A(n1003), .B(n1004), .Z(n1001) );
  NAND U879 ( .A(n1005), .B(n1006), .Z(n1004) );
  NANDN U880 ( .A(A[5]), .B(B[5]), .Z(n1006) );
  AND U881 ( .A(n1007), .B(n1008), .Z(n1005) );
  NANDN U882 ( .A(A[4]), .B(B[4]), .Z(n1008) );
  NAND U883 ( .A(n1009), .B(n1010), .Z(n1007) );
  NANDN U884 ( .A(B[4]), .B(A[4]), .Z(n1010) );
  AND U885 ( .A(n1011), .B(n1012), .Z(n1009) );
  NAND U886 ( .A(n1013), .B(n1014), .Z(n1012) );
  NANDN U887 ( .A(A[3]), .B(B[3]), .Z(n1014) );
  AND U888 ( .A(n1015), .B(n1016), .Z(n1013) );
  NANDN U889 ( .A(A[2]), .B(B[2]), .Z(n1016) );
  NAND U890 ( .A(n1017), .B(n1018), .Z(n1015) );
  NANDN U891 ( .A(B[2]), .B(A[2]), .Z(n1018) );
  AND U892 ( .A(n1019), .B(n1020), .Z(n1017) );
  NANDN U893 ( .A(B[1]), .B(n1021), .Z(n1020) );
  NANDN U894 ( .A(A[1]), .B(n1022), .Z(n1021) );
  NANDN U895 ( .A(n1022), .B(A[1]), .Z(n1019) );
  ANDN U896 ( .B(B[0]), .A(A[0]), .Z(n1022) );
  NANDN U897 ( .A(B[3]), .B(A[3]), .Z(n1011) );
  NANDN U898 ( .A(B[5]), .B(A[5]), .Z(n1003) );
  NANDN U899 ( .A(B[7]), .B(A[7]), .Z(n995) );
  NANDN U900 ( .A(B[10]), .B(A[10]), .Z(n987) );
  NANDN U901 ( .A(B[11]), .B(A[11]), .Z(n979) );
  NANDN U902 ( .A(B[13]), .B(A[13]), .Z(n971) );
  NANDN U903 ( .A(B[15]), .B(A[15]), .Z(n963) );
  NANDN U904 ( .A(B[17]), .B(A[17]), .Z(n955) );
  NANDN U905 ( .A(B[19]), .B(A[19]), .Z(n947) );
  NANDN U906 ( .A(B[21]), .B(A[21]), .Z(n939) );
  NANDN U907 ( .A(B[23]), .B(A[23]), .Z(n931) );
  NANDN U908 ( .A(B[25]), .B(A[25]), .Z(n923) );
  NANDN U909 ( .A(B[27]), .B(A[27]), .Z(n915) );
  NANDN U910 ( .A(B[29]), .B(A[29]), .Z(n907) );
  NANDN U911 ( .A(B[31]), .B(A[31]), .Z(n899) );
  NANDN U912 ( .A(B[33]), .B(A[33]), .Z(n891) );
  NANDN U913 ( .A(B[35]), .B(A[35]), .Z(n883) );
  NANDN U914 ( .A(B[37]), .B(A[37]), .Z(n875) );
  NANDN U915 ( .A(B[39]), .B(A[39]), .Z(n867) );
  NANDN U916 ( .A(B[41]), .B(A[41]), .Z(n859) );
  NANDN U917 ( .A(B[43]), .B(A[43]), .Z(n851) );
  NANDN U918 ( .A(B[45]), .B(A[45]), .Z(n843) );
  NANDN U919 ( .A(B[47]), .B(A[47]), .Z(n835) );
  NANDN U920 ( .A(B[49]), .B(A[49]), .Z(n827) );
  NANDN U921 ( .A(B[51]), .B(A[51]), .Z(n819) );
  NANDN U922 ( .A(B[53]), .B(A[53]), .Z(n811) );
  NANDN U923 ( .A(B[55]), .B(A[55]), .Z(n803) );
  NANDN U924 ( .A(B[57]), .B(A[57]), .Z(n795) );
  NANDN U925 ( .A(B[59]), .B(A[59]), .Z(n787) );
  NANDN U926 ( .A(B[61]), .B(A[61]), .Z(n779) );
  NANDN U927 ( .A(B[63]), .B(A[63]), .Z(n771) );
  NANDN U928 ( .A(B[65]), .B(A[65]), .Z(n763) );
  NANDN U929 ( .A(B[67]), .B(A[67]), .Z(n755) );
  NANDN U930 ( .A(B[69]), .B(A[69]), .Z(n747) );
  NANDN U931 ( .A(B[71]), .B(A[71]), .Z(n739) );
  NANDN U932 ( .A(B[73]), .B(A[73]), .Z(n731) );
  NANDN U933 ( .A(B[75]), .B(A[75]), .Z(n723) );
  NANDN U934 ( .A(B[77]), .B(A[77]), .Z(n715) );
  NANDN U935 ( .A(B[79]), .B(A[79]), .Z(n707) );
  NANDN U936 ( .A(B[81]), .B(A[81]), .Z(n699) );
  NANDN U937 ( .A(B[83]), .B(A[83]), .Z(n691) );
  NANDN U938 ( .A(B[85]), .B(A[85]), .Z(n683) );
  NANDN U939 ( .A(B[87]), .B(A[87]), .Z(n675) );
  NANDN U940 ( .A(B[89]), .B(A[89]), .Z(n667) );
  NANDN U941 ( .A(B[91]), .B(A[91]), .Z(n659) );
  NANDN U942 ( .A(B[93]), .B(A[93]), .Z(n651) );
  NANDN U943 ( .A(B[95]), .B(A[95]), .Z(n643) );
  NANDN U944 ( .A(B[97]), .B(A[97]), .Z(n635) );
  NANDN U945 ( .A(B[100]), .B(A[100]), .Z(n627) );
  NANDN U946 ( .A(B[101]), .B(A[101]), .Z(n619) );
  NANDN U947 ( .A(B[103]), .B(A[103]), .Z(n611) );
  NANDN U948 ( .A(B[105]), .B(A[105]), .Z(n603) );
  NANDN U949 ( .A(B[107]), .B(A[107]), .Z(n595) );
  NANDN U950 ( .A(B[109]), .B(A[109]), .Z(n587) );
  NANDN U951 ( .A(B[111]), .B(A[111]), .Z(n579) );
  NANDN U952 ( .A(B[113]), .B(A[113]), .Z(n571) );
  NANDN U953 ( .A(B[115]), .B(A[115]), .Z(n563) );
  NANDN U954 ( .A(B[117]), .B(A[117]), .Z(n555) );
  NANDN U955 ( .A(B[119]), .B(A[119]), .Z(n547) );
  NANDN U956 ( .A(B[121]), .B(A[121]), .Z(n539) );
  NANDN U957 ( .A(B[123]), .B(A[123]), .Z(n531) );
  NANDN U958 ( .A(B[125]), .B(A[125]), .Z(n523) );
  NANDN U959 ( .A(B[127]), .B(A[127]), .Z(n515) );
  NANDN U960 ( .A(B[129]), .B(A[129]), .Z(n507) );
  NANDN U961 ( .A(B[131]), .B(A[131]), .Z(n499) );
  NANDN U962 ( .A(B[133]), .B(A[133]), .Z(n491) );
  NANDN U963 ( .A(B[135]), .B(A[135]), .Z(n483) );
  NANDN U964 ( .A(B[137]), .B(A[137]), .Z(n475) );
  NANDN U965 ( .A(B[139]), .B(A[139]), .Z(n467) );
  NANDN U966 ( .A(B[141]), .B(A[141]), .Z(n459) );
  NANDN U967 ( .A(B[143]), .B(A[143]), .Z(n451) );
  NANDN U968 ( .A(B[145]), .B(A[145]), .Z(n443) );
  NANDN U969 ( .A(B[147]), .B(A[147]), .Z(n435) );
  NANDN U970 ( .A(B[149]), .B(A[149]), .Z(n427) );
  NANDN U971 ( .A(B[151]), .B(A[151]), .Z(n419) );
  NANDN U972 ( .A(B[153]), .B(A[153]), .Z(n411) );
  NANDN U973 ( .A(B[155]), .B(A[155]), .Z(n403) );
  NANDN U974 ( .A(B[157]), .B(A[157]), .Z(n395) );
  NANDN U975 ( .A(B[159]), .B(A[159]), .Z(n387) );
  NANDN U976 ( .A(B[161]), .B(A[161]), .Z(n379) );
  NANDN U977 ( .A(B[163]), .B(A[163]), .Z(n371) );
  NANDN U978 ( .A(B[165]), .B(A[165]), .Z(n363) );
  NANDN U979 ( .A(B[167]), .B(A[167]), .Z(n355) );
  NANDN U980 ( .A(B[169]), .B(A[169]), .Z(n347) );
  NANDN U981 ( .A(B[171]), .B(A[171]), .Z(n339) );
  NANDN U982 ( .A(B[173]), .B(A[173]), .Z(n331) );
  NANDN U983 ( .A(B[175]), .B(A[175]), .Z(n323) );
  NANDN U984 ( .A(B[177]), .B(A[177]), .Z(n315) );
  NANDN U985 ( .A(B[179]), .B(A[179]), .Z(n307) );
  NANDN U986 ( .A(B[181]), .B(A[181]), .Z(n299) );
  NANDN U987 ( .A(B[183]), .B(A[183]), .Z(n291) );
  NANDN U988 ( .A(B[185]), .B(A[185]), .Z(n283) );
  NANDN U989 ( .A(B[187]), .B(A[187]), .Z(n275) );
  NANDN U990 ( .A(B[189]), .B(A[189]), .Z(n267) );
  NANDN U991 ( .A(B[191]), .B(A[191]), .Z(n259) );
  NANDN U992 ( .A(B[193]), .B(A[193]), .Z(n251) );
  NANDN U993 ( .A(B[195]), .B(A[195]), .Z(n243) );
  NANDN U994 ( .A(B[197]), .B(A[197]), .Z(n235) );
  NANDN U995 ( .A(B[199]), .B(A[199]), .Z(n227) );
  NANDN U996 ( .A(B[201]), .B(A[201]), .Z(n219) );
  NANDN U997 ( .A(B[203]), .B(A[203]), .Z(n211) );
  NANDN U998 ( .A(B[205]), .B(A[205]), .Z(n203) );
  NANDN U999 ( .A(B[207]), .B(A[207]), .Z(n195) );
  NANDN U1000 ( .A(B[209]), .B(A[209]), .Z(n187) );
  NANDN U1001 ( .A(B[211]), .B(A[211]), .Z(n179) );
  NANDN U1002 ( .A(B[213]), .B(A[213]), .Z(n171) );
  NANDN U1003 ( .A(B[215]), .B(A[215]), .Z(n163) );
  NANDN U1004 ( .A(B[217]), .B(A[217]), .Z(n155) );
  NANDN U1005 ( .A(B[219]), .B(A[219]), .Z(n147) );
  NANDN U1006 ( .A(B[221]), .B(A[221]), .Z(n139) );
  NANDN U1007 ( .A(B[223]), .B(A[223]), .Z(n131) );
  NANDN U1008 ( .A(B[225]), .B(A[225]), .Z(n123) );
  NANDN U1009 ( .A(B[227]), .B(A[227]), .Z(n115) );
  NANDN U1010 ( .A(B[229]), .B(A[229]), .Z(n107) );
  NANDN U1011 ( .A(B[231]), .B(A[231]), .Z(n99) );
  NANDN U1012 ( .A(B[233]), .B(A[233]), .Z(n91) );
  NANDN U1013 ( .A(B[235]), .B(A[235]), .Z(n83) );
  NANDN U1014 ( .A(B[237]), .B(A[237]), .Z(n75) );
  NANDN U1015 ( .A(B[239]), .B(A[239]), .Z(n67) );
  NANDN U1016 ( .A(B[241]), .B(A[241]), .Z(n59) );
  NANDN U1017 ( .A(B[243]), .B(A[243]), .Z(n51) );
  NANDN U1018 ( .A(B[245]), .B(A[245]), .Z(n43) );
  NANDN U1019 ( .A(B[247]), .B(A[247]), .Z(n35) );
  NANDN U1020 ( .A(B[249]), .B(A[249]), .Z(n27) );
  NANDN U1021 ( .A(B[251]), .B(A[251]), .Z(n19) );
  NANDN U1022 ( .A(B[253]), .B(A[253]), .Z(n11) );
  NANDN U1023 ( .A(A[255]), .B(B[255]), .Z(n3) );
endmodule


module modmult_step_N256_4_DW01_add_0 ( A, B, CI, SUM, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] SUM;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272;
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];

  XNOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(SUM[99]) );
  XNOR U4 ( .A(B[99]), .B(A[99]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[98]) );
  XNOR U6 ( .A(B[98]), .B(A[98]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[97]) );
  XNOR U8 ( .A(B[97]), .B(A[97]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[96]) );
  XNOR U10 ( .A(B[96]), .B(A[96]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[95]) );
  XNOR U12 ( .A(B[95]), .B(A[95]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[94]) );
  XNOR U14 ( .A(B[94]), .B(A[94]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[93]) );
  XNOR U16 ( .A(B[93]), .B(A[93]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(SUM[92]) );
  XNOR U18 ( .A(B[92]), .B(A[92]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(SUM[91]) );
  XNOR U20 ( .A(B[91]), .B(A[91]), .Z(n20) );
  XOR U21 ( .A(n21), .B(n22), .Z(SUM[90]) );
  XNOR U22 ( .A(B[90]), .B(A[90]), .Z(n22) );
  XOR U23 ( .A(n23), .B(n24), .Z(SUM[8]) );
  XNOR U24 ( .A(B[8]), .B(A[8]), .Z(n24) );
  XOR U25 ( .A(n25), .B(n26), .Z(SUM[89]) );
  XNOR U26 ( .A(B[89]), .B(A[89]), .Z(n26) );
  XOR U27 ( .A(n27), .B(n28), .Z(SUM[88]) );
  XNOR U28 ( .A(B[88]), .B(A[88]), .Z(n28) );
  XOR U29 ( .A(n29), .B(n30), .Z(SUM[87]) );
  XNOR U30 ( .A(B[87]), .B(A[87]), .Z(n30) );
  XOR U31 ( .A(n31), .B(n32), .Z(SUM[86]) );
  XNOR U32 ( .A(B[86]), .B(A[86]), .Z(n32) );
  XOR U33 ( .A(n33), .B(n34), .Z(SUM[85]) );
  XNOR U34 ( .A(B[85]), .B(A[85]), .Z(n34) );
  XOR U35 ( .A(n35), .B(n36), .Z(SUM[84]) );
  XNOR U36 ( .A(B[84]), .B(A[84]), .Z(n36) );
  XOR U37 ( .A(n37), .B(n38), .Z(SUM[83]) );
  XNOR U38 ( .A(B[83]), .B(A[83]), .Z(n38) );
  XOR U39 ( .A(n39), .B(n40), .Z(SUM[82]) );
  XNOR U40 ( .A(B[82]), .B(A[82]), .Z(n40) );
  XOR U41 ( .A(n41), .B(n42), .Z(SUM[81]) );
  XNOR U42 ( .A(B[81]), .B(A[81]), .Z(n42) );
  XOR U43 ( .A(n43), .B(n44), .Z(SUM[80]) );
  XNOR U44 ( .A(B[80]), .B(A[80]), .Z(n44) );
  XOR U45 ( .A(n45), .B(n46), .Z(SUM[7]) );
  XNOR U46 ( .A(B[7]), .B(A[7]), .Z(n46) );
  XOR U47 ( .A(n47), .B(n48), .Z(SUM[79]) );
  XNOR U48 ( .A(B[79]), .B(A[79]), .Z(n48) );
  XOR U49 ( .A(n49), .B(n50), .Z(SUM[78]) );
  XNOR U50 ( .A(B[78]), .B(A[78]), .Z(n50) );
  XOR U51 ( .A(n51), .B(n52), .Z(SUM[77]) );
  XNOR U52 ( .A(B[77]), .B(A[77]), .Z(n52) );
  XOR U53 ( .A(n53), .B(n54), .Z(SUM[76]) );
  XNOR U54 ( .A(B[76]), .B(A[76]), .Z(n54) );
  XOR U55 ( .A(n55), .B(n56), .Z(SUM[75]) );
  XNOR U56 ( .A(B[75]), .B(A[75]), .Z(n56) );
  XOR U57 ( .A(n57), .B(n58), .Z(SUM[74]) );
  XNOR U58 ( .A(B[74]), .B(A[74]), .Z(n58) );
  XOR U59 ( .A(n59), .B(n60), .Z(SUM[73]) );
  XNOR U60 ( .A(B[73]), .B(A[73]), .Z(n60) );
  XOR U61 ( .A(n61), .B(n62), .Z(SUM[72]) );
  XNOR U62 ( .A(B[72]), .B(A[72]), .Z(n62) );
  XOR U63 ( .A(n63), .B(n64), .Z(SUM[71]) );
  XNOR U64 ( .A(B[71]), .B(A[71]), .Z(n64) );
  XOR U65 ( .A(n65), .B(n66), .Z(SUM[70]) );
  XNOR U66 ( .A(B[70]), .B(A[70]), .Z(n66) );
  XOR U67 ( .A(n67), .B(n68), .Z(SUM[6]) );
  XNOR U68 ( .A(B[6]), .B(A[6]), .Z(n68) );
  XOR U69 ( .A(n69), .B(n70), .Z(SUM[69]) );
  XNOR U70 ( .A(B[69]), .B(A[69]), .Z(n70) );
  XOR U71 ( .A(n71), .B(n72), .Z(SUM[68]) );
  XNOR U72 ( .A(B[68]), .B(A[68]), .Z(n72) );
  XOR U73 ( .A(n73), .B(n74), .Z(SUM[67]) );
  XNOR U74 ( .A(B[67]), .B(A[67]), .Z(n74) );
  XOR U75 ( .A(n75), .B(n76), .Z(SUM[66]) );
  XNOR U76 ( .A(B[66]), .B(A[66]), .Z(n76) );
  XOR U77 ( .A(n77), .B(n78), .Z(SUM[65]) );
  XNOR U78 ( .A(B[65]), .B(A[65]), .Z(n78) );
  XOR U79 ( .A(n79), .B(n80), .Z(SUM[64]) );
  XNOR U80 ( .A(B[64]), .B(A[64]), .Z(n80) );
  XOR U81 ( .A(n81), .B(n82), .Z(SUM[63]) );
  XNOR U82 ( .A(B[63]), .B(A[63]), .Z(n82) );
  XOR U83 ( .A(n83), .B(n84), .Z(SUM[62]) );
  XNOR U84 ( .A(B[62]), .B(A[62]), .Z(n84) );
  XOR U85 ( .A(n85), .B(n86), .Z(SUM[61]) );
  XNOR U86 ( .A(B[61]), .B(A[61]), .Z(n86) );
  XOR U87 ( .A(n87), .B(n88), .Z(SUM[60]) );
  XNOR U88 ( .A(B[60]), .B(A[60]), .Z(n88) );
  XOR U89 ( .A(n89), .B(n90), .Z(SUM[5]) );
  XNOR U90 ( .A(B[5]), .B(A[5]), .Z(n90) );
  XOR U91 ( .A(n91), .B(n92), .Z(SUM[59]) );
  XNOR U92 ( .A(B[59]), .B(A[59]), .Z(n92) );
  XOR U93 ( .A(n93), .B(n94), .Z(SUM[58]) );
  XNOR U94 ( .A(B[58]), .B(A[58]), .Z(n94) );
  XOR U95 ( .A(n95), .B(n96), .Z(SUM[57]) );
  XNOR U96 ( .A(B[57]), .B(A[57]), .Z(n96) );
  XOR U97 ( .A(n97), .B(n98), .Z(SUM[56]) );
  XNOR U98 ( .A(B[56]), .B(A[56]), .Z(n98) );
  XOR U99 ( .A(n99), .B(n100), .Z(SUM[55]) );
  XNOR U100 ( .A(B[55]), .B(A[55]), .Z(n100) );
  XOR U101 ( .A(n101), .B(n102), .Z(SUM[54]) );
  XNOR U102 ( .A(B[54]), .B(A[54]), .Z(n102) );
  XOR U103 ( .A(n103), .B(n104), .Z(SUM[53]) );
  XNOR U104 ( .A(B[53]), .B(A[53]), .Z(n104) );
  XOR U105 ( .A(n105), .B(n106), .Z(SUM[52]) );
  XNOR U106 ( .A(B[52]), .B(A[52]), .Z(n106) );
  XOR U107 ( .A(n107), .B(n108), .Z(SUM[51]) );
  XNOR U108 ( .A(B[51]), .B(A[51]), .Z(n108) );
  XOR U109 ( .A(n109), .B(n110), .Z(SUM[50]) );
  XNOR U110 ( .A(B[50]), .B(A[50]), .Z(n110) );
  XOR U111 ( .A(n111), .B(n112), .Z(SUM[4]) );
  XNOR U112 ( .A(B[4]), .B(A[4]), .Z(n112) );
  XOR U113 ( .A(n113), .B(n114), .Z(SUM[49]) );
  XNOR U114 ( .A(B[49]), .B(A[49]), .Z(n114) );
  XOR U115 ( .A(n115), .B(n116), .Z(SUM[48]) );
  XNOR U116 ( .A(B[48]), .B(A[48]), .Z(n116) );
  XOR U117 ( .A(n117), .B(n118), .Z(SUM[47]) );
  XNOR U118 ( .A(B[47]), .B(A[47]), .Z(n118) );
  XOR U119 ( .A(n119), .B(n120), .Z(SUM[46]) );
  XNOR U120 ( .A(B[46]), .B(A[46]), .Z(n120) );
  XOR U121 ( .A(n121), .B(n122), .Z(SUM[45]) );
  XNOR U122 ( .A(B[45]), .B(A[45]), .Z(n122) );
  XOR U123 ( .A(n123), .B(n124), .Z(SUM[44]) );
  XNOR U124 ( .A(B[44]), .B(A[44]), .Z(n124) );
  XOR U125 ( .A(n125), .B(n126), .Z(SUM[43]) );
  XNOR U126 ( .A(B[43]), .B(A[43]), .Z(n126) );
  XOR U127 ( .A(n127), .B(n128), .Z(SUM[42]) );
  XNOR U128 ( .A(B[42]), .B(A[42]), .Z(n128) );
  XOR U129 ( .A(n129), .B(n130), .Z(SUM[41]) );
  XNOR U130 ( .A(B[41]), .B(A[41]), .Z(n130) );
  XOR U131 ( .A(n131), .B(n132), .Z(SUM[40]) );
  XNOR U132 ( .A(B[40]), .B(A[40]), .Z(n132) );
  XOR U133 ( .A(n133), .B(n134), .Z(SUM[3]) );
  XNOR U134 ( .A(B[3]), .B(A[3]), .Z(n134) );
  XOR U135 ( .A(n135), .B(n136), .Z(SUM[39]) );
  XNOR U136 ( .A(B[39]), .B(A[39]), .Z(n136) );
  XOR U137 ( .A(n137), .B(n138), .Z(SUM[38]) );
  XNOR U138 ( .A(B[38]), .B(A[38]), .Z(n138) );
  XOR U139 ( .A(n139), .B(n140), .Z(SUM[37]) );
  XNOR U140 ( .A(B[37]), .B(A[37]), .Z(n140) );
  XOR U141 ( .A(n141), .B(n142), .Z(SUM[36]) );
  XNOR U142 ( .A(B[36]), .B(A[36]), .Z(n142) );
  XOR U143 ( .A(n143), .B(n144), .Z(SUM[35]) );
  XNOR U144 ( .A(B[35]), .B(A[35]), .Z(n144) );
  XOR U145 ( .A(n145), .B(n146), .Z(SUM[34]) );
  XNOR U146 ( .A(B[34]), .B(A[34]), .Z(n146) );
  XOR U147 ( .A(n147), .B(n148), .Z(SUM[33]) );
  XNOR U148 ( .A(B[33]), .B(A[33]), .Z(n148) );
  XOR U149 ( .A(n149), .B(n150), .Z(SUM[32]) );
  XNOR U150 ( .A(B[32]), .B(A[32]), .Z(n150) );
  XOR U151 ( .A(n151), .B(n152), .Z(SUM[31]) );
  XNOR U152 ( .A(B[31]), .B(A[31]), .Z(n152) );
  XOR U153 ( .A(n153), .B(n154), .Z(SUM[30]) );
  XNOR U154 ( .A(B[30]), .B(A[30]), .Z(n154) );
  XOR U155 ( .A(n155), .B(n156), .Z(SUM[2]) );
  XOR U156 ( .A(B[2]), .B(A[2]), .Z(n156) );
  XOR U157 ( .A(n157), .B(n158), .Z(SUM[29]) );
  XNOR U158 ( .A(B[29]), .B(A[29]), .Z(n158) );
  XOR U159 ( .A(n159), .B(n160), .Z(SUM[28]) );
  XNOR U160 ( .A(B[28]), .B(A[28]), .Z(n160) );
  XOR U161 ( .A(n161), .B(n162), .Z(SUM[27]) );
  XNOR U162 ( .A(B[27]), .B(A[27]), .Z(n162) );
  XOR U163 ( .A(n163), .B(n164), .Z(SUM[26]) );
  XNOR U164 ( .A(B[26]), .B(A[26]), .Z(n164) );
  XOR U165 ( .A(n165), .B(n166), .Z(SUM[25]) );
  XNOR U166 ( .A(B[25]), .B(A[25]), .Z(n166) );
  XOR U167 ( .A(A[257]), .B(n167), .Z(SUM[257]) );
  AND U168 ( .A(A[256]), .B(n168), .Z(n167) );
  XOR U169 ( .A(A[256]), .B(n168), .Z(SUM[256]) );
  NAND U170 ( .A(n169), .B(n170), .Z(n168) );
  NAND U171 ( .A(B[255]), .B(n171), .Z(n170) );
  NANDN U172 ( .A(A[255]), .B(n172), .Z(n171) );
  NANDN U173 ( .A(n172), .B(A[255]), .Z(n169) );
  XOR U174 ( .A(n172), .B(n173), .Z(SUM[255]) );
  XNOR U175 ( .A(B[255]), .B(A[255]), .Z(n173) );
  AND U176 ( .A(n174), .B(n175), .Z(n172) );
  NAND U177 ( .A(B[254]), .B(n176), .Z(n175) );
  NANDN U178 ( .A(A[254]), .B(n177), .Z(n176) );
  NANDN U179 ( .A(n177), .B(A[254]), .Z(n174) );
  XOR U180 ( .A(n177), .B(n178), .Z(SUM[254]) );
  XNOR U181 ( .A(B[254]), .B(A[254]), .Z(n178) );
  AND U182 ( .A(n179), .B(n180), .Z(n177) );
  NAND U183 ( .A(B[253]), .B(n181), .Z(n180) );
  NANDN U184 ( .A(A[253]), .B(n182), .Z(n181) );
  NANDN U185 ( .A(n182), .B(A[253]), .Z(n179) );
  XOR U186 ( .A(n182), .B(n183), .Z(SUM[253]) );
  XNOR U187 ( .A(B[253]), .B(A[253]), .Z(n183) );
  AND U188 ( .A(n184), .B(n185), .Z(n182) );
  NAND U189 ( .A(B[252]), .B(n186), .Z(n185) );
  NANDN U190 ( .A(A[252]), .B(n187), .Z(n186) );
  NANDN U191 ( .A(n187), .B(A[252]), .Z(n184) );
  XOR U192 ( .A(n187), .B(n188), .Z(SUM[252]) );
  XNOR U193 ( .A(B[252]), .B(A[252]), .Z(n188) );
  AND U194 ( .A(n189), .B(n190), .Z(n187) );
  NAND U195 ( .A(B[251]), .B(n191), .Z(n190) );
  NANDN U196 ( .A(A[251]), .B(n192), .Z(n191) );
  NANDN U197 ( .A(n192), .B(A[251]), .Z(n189) );
  XOR U198 ( .A(n192), .B(n193), .Z(SUM[251]) );
  XNOR U199 ( .A(B[251]), .B(A[251]), .Z(n193) );
  AND U200 ( .A(n194), .B(n195), .Z(n192) );
  NAND U201 ( .A(B[250]), .B(n196), .Z(n195) );
  NANDN U202 ( .A(A[250]), .B(n197), .Z(n196) );
  NANDN U203 ( .A(n197), .B(A[250]), .Z(n194) );
  XOR U204 ( .A(n197), .B(n198), .Z(SUM[250]) );
  XNOR U205 ( .A(B[250]), .B(A[250]), .Z(n198) );
  AND U206 ( .A(n199), .B(n200), .Z(n197) );
  NAND U207 ( .A(B[249]), .B(n201), .Z(n200) );
  NANDN U208 ( .A(A[249]), .B(n202), .Z(n201) );
  NANDN U209 ( .A(n202), .B(A[249]), .Z(n199) );
  XOR U210 ( .A(n203), .B(n204), .Z(SUM[24]) );
  XNOR U211 ( .A(B[24]), .B(A[24]), .Z(n204) );
  XOR U212 ( .A(n202), .B(n205), .Z(SUM[249]) );
  XNOR U213 ( .A(B[249]), .B(A[249]), .Z(n205) );
  AND U214 ( .A(n206), .B(n207), .Z(n202) );
  NAND U215 ( .A(B[248]), .B(n208), .Z(n207) );
  NANDN U216 ( .A(A[248]), .B(n209), .Z(n208) );
  NANDN U217 ( .A(n209), .B(A[248]), .Z(n206) );
  XOR U218 ( .A(n209), .B(n210), .Z(SUM[248]) );
  XNOR U219 ( .A(B[248]), .B(A[248]), .Z(n210) );
  AND U220 ( .A(n211), .B(n212), .Z(n209) );
  NAND U221 ( .A(B[247]), .B(n213), .Z(n212) );
  NANDN U222 ( .A(A[247]), .B(n214), .Z(n213) );
  NANDN U223 ( .A(n214), .B(A[247]), .Z(n211) );
  XOR U224 ( .A(n214), .B(n215), .Z(SUM[247]) );
  XNOR U225 ( .A(B[247]), .B(A[247]), .Z(n215) );
  AND U226 ( .A(n216), .B(n217), .Z(n214) );
  NAND U227 ( .A(B[246]), .B(n218), .Z(n217) );
  NANDN U228 ( .A(A[246]), .B(n219), .Z(n218) );
  NANDN U229 ( .A(n219), .B(A[246]), .Z(n216) );
  XOR U230 ( .A(n219), .B(n220), .Z(SUM[246]) );
  XNOR U231 ( .A(B[246]), .B(A[246]), .Z(n220) );
  AND U232 ( .A(n221), .B(n222), .Z(n219) );
  NAND U233 ( .A(B[245]), .B(n223), .Z(n222) );
  NANDN U234 ( .A(A[245]), .B(n224), .Z(n223) );
  NANDN U235 ( .A(n224), .B(A[245]), .Z(n221) );
  XOR U236 ( .A(n224), .B(n225), .Z(SUM[245]) );
  XNOR U237 ( .A(B[245]), .B(A[245]), .Z(n225) );
  AND U238 ( .A(n226), .B(n227), .Z(n224) );
  NAND U239 ( .A(B[244]), .B(n228), .Z(n227) );
  NANDN U240 ( .A(A[244]), .B(n229), .Z(n228) );
  NANDN U241 ( .A(n229), .B(A[244]), .Z(n226) );
  XOR U242 ( .A(n229), .B(n230), .Z(SUM[244]) );
  XNOR U243 ( .A(B[244]), .B(A[244]), .Z(n230) );
  AND U244 ( .A(n231), .B(n232), .Z(n229) );
  NAND U245 ( .A(B[243]), .B(n233), .Z(n232) );
  NANDN U246 ( .A(A[243]), .B(n234), .Z(n233) );
  NANDN U247 ( .A(n234), .B(A[243]), .Z(n231) );
  XOR U248 ( .A(n234), .B(n235), .Z(SUM[243]) );
  XNOR U249 ( .A(B[243]), .B(A[243]), .Z(n235) );
  AND U250 ( .A(n236), .B(n237), .Z(n234) );
  NAND U251 ( .A(B[242]), .B(n238), .Z(n237) );
  NANDN U252 ( .A(A[242]), .B(n239), .Z(n238) );
  NANDN U253 ( .A(n239), .B(A[242]), .Z(n236) );
  XOR U254 ( .A(n239), .B(n240), .Z(SUM[242]) );
  XNOR U255 ( .A(B[242]), .B(A[242]), .Z(n240) );
  AND U256 ( .A(n241), .B(n242), .Z(n239) );
  NAND U257 ( .A(B[241]), .B(n243), .Z(n242) );
  NANDN U258 ( .A(A[241]), .B(n244), .Z(n243) );
  NANDN U259 ( .A(n244), .B(A[241]), .Z(n241) );
  XOR U260 ( .A(n244), .B(n245), .Z(SUM[241]) );
  XNOR U261 ( .A(B[241]), .B(A[241]), .Z(n245) );
  AND U262 ( .A(n246), .B(n247), .Z(n244) );
  NAND U263 ( .A(B[240]), .B(n248), .Z(n247) );
  NANDN U264 ( .A(A[240]), .B(n249), .Z(n248) );
  NANDN U265 ( .A(n249), .B(A[240]), .Z(n246) );
  XOR U266 ( .A(n249), .B(n250), .Z(SUM[240]) );
  XNOR U267 ( .A(B[240]), .B(A[240]), .Z(n250) );
  AND U268 ( .A(n251), .B(n252), .Z(n249) );
  NAND U269 ( .A(B[239]), .B(n253), .Z(n252) );
  NANDN U270 ( .A(A[239]), .B(n254), .Z(n253) );
  NANDN U271 ( .A(n254), .B(A[239]), .Z(n251) );
  XOR U272 ( .A(n255), .B(n256), .Z(SUM[23]) );
  XNOR U273 ( .A(B[23]), .B(A[23]), .Z(n256) );
  XOR U274 ( .A(n254), .B(n257), .Z(SUM[239]) );
  XNOR U275 ( .A(B[239]), .B(A[239]), .Z(n257) );
  AND U276 ( .A(n258), .B(n259), .Z(n254) );
  NAND U277 ( .A(B[238]), .B(n260), .Z(n259) );
  NANDN U278 ( .A(A[238]), .B(n261), .Z(n260) );
  NANDN U279 ( .A(n261), .B(A[238]), .Z(n258) );
  XOR U280 ( .A(n261), .B(n262), .Z(SUM[238]) );
  XNOR U281 ( .A(B[238]), .B(A[238]), .Z(n262) );
  AND U282 ( .A(n263), .B(n264), .Z(n261) );
  NAND U283 ( .A(B[237]), .B(n265), .Z(n264) );
  NANDN U284 ( .A(A[237]), .B(n266), .Z(n265) );
  NANDN U285 ( .A(n266), .B(A[237]), .Z(n263) );
  XOR U286 ( .A(n266), .B(n267), .Z(SUM[237]) );
  XNOR U287 ( .A(B[237]), .B(A[237]), .Z(n267) );
  AND U288 ( .A(n268), .B(n269), .Z(n266) );
  NAND U289 ( .A(B[236]), .B(n270), .Z(n269) );
  NANDN U290 ( .A(A[236]), .B(n271), .Z(n270) );
  NANDN U291 ( .A(n271), .B(A[236]), .Z(n268) );
  XOR U292 ( .A(n271), .B(n272), .Z(SUM[236]) );
  XNOR U293 ( .A(B[236]), .B(A[236]), .Z(n272) );
  AND U294 ( .A(n273), .B(n274), .Z(n271) );
  NAND U295 ( .A(B[235]), .B(n275), .Z(n274) );
  NANDN U296 ( .A(A[235]), .B(n276), .Z(n275) );
  NANDN U297 ( .A(n276), .B(A[235]), .Z(n273) );
  XOR U298 ( .A(n276), .B(n277), .Z(SUM[235]) );
  XNOR U299 ( .A(B[235]), .B(A[235]), .Z(n277) );
  AND U300 ( .A(n278), .B(n279), .Z(n276) );
  NAND U301 ( .A(B[234]), .B(n280), .Z(n279) );
  NANDN U302 ( .A(A[234]), .B(n281), .Z(n280) );
  NANDN U303 ( .A(n281), .B(A[234]), .Z(n278) );
  XOR U304 ( .A(n281), .B(n282), .Z(SUM[234]) );
  XNOR U305 ( .A(B[234]), .B(A[234]), .Z(n282) );
  AND U306 ( .A(n283), .B(n284), .Z(n281) );
  NAND U307 ( .A(B[233]), .B(n285), .Z(n284) );
  NANDN U308 ( .A(A[233]), .B(n286), .Z(n285) );
  NANDN U309 ( .A(n286), .B(A[233]), .Z(n283) );
  XOR U310 ( .A(n286), .B(n287), .Z(SUM[233]) );
  XNOR U311 ( .A(B[233]), .B(A[233]), .Z(n287) );
  AND U312 ( .A(n288), .B(n289), .Z(n286) );
  NAND U313 ( .A(B[232]), .B(n290), .Z(n289) );
  NANDN U314 ( .A(A[232]), .B(n291), .Z(n290) );
  NANDN U315 ( .A(n291), .B(A[232]), .Z(n288) );
  XOR U316 ( .A(n291), .B(n292), .Z(SUM[232]) );
  XNOR U317 ( .A(B[232]), .B(A[232]), .Z(n292) );
  AND U318 ( .A(n293), .B(n294), .Z(n291) );
  NAND U319 ( .A(B[231]), .B(n295), .Z(n294) );
  NANDN U320 ( .A(A[231]), .B(n296), .Z(n295) );
  NANDN U321 ( .A(n296), .B(A[231]), .Z(n293) );
  XOR U322 ( .A(n296), .B(n297), .Z(SUM[231]) );
  XNOR U323 ( .A(B[231]), .B(A[231]), .Z(n297) );
  AND U324 ( .A(n298), .B(n299), .Z(n296) );
  NAND U325 ( .A(B[230]), .B(n300), .Z(n299) );
  NANDN U326 ( .A(A[230]), .B(n301), .Z(n300) );
  NANDN U327 ( .A(n301), .B(A[230]), .Z(n298) );
  XOR U328 ( .A(n301), .B(n302), .Z(SUM[230]) );
  XNOR U329 ( .A(B[230]), .B(A[230]), .Z(n302) );
  AND U330 ( .A(n303), .B(n304), .Z(n301) );
  NAND U331 ( .A(B[229]), .B(n305), .Z(n304) );
  NANDN U332 ( .A(A[229]), .B(n306), .Z(n305) );
  NANDN U333 ( .A(n306), .B(A[229]), .Z(n303) );
  XOR U334 ( .A(n307), .B(n308), .Z(SUM[22]) );
  XNOR U335 ( .A(B[22]), .B(A[22]), .Z(n308) );
  XOR U336 ( .A(n306), .B(n309), .Z(SUM[229]) );
  XNOR U337 ( .A(B[229]), .B(A[229]), .Z(n309) );
  AND U338 ( .A(n310), .B(n311), .Z(n306) );
  NAND U339 ( .A(B[228]), .B(n312), .Z(n311) );
  NANDN U340 ( .A(A[228]), .B(n313), .Z(n312) );
  NANDN U341 ( .A(n313), .B(A[228]), .Z(n310) );
  XOR U342 ( .A(n313), .B(n314), .Z(SUM[228]) );
  XNOR U343 ( .A(B[228]), .B(A[228]), .Z(n314) );
  AND U344 ( .A(n315), .B(n316), .Z(n313) );
  NAND U345 ( .A(B[227]), .B(n317), .Z(n316) );
  NANDN U346 ( .A(A[227]), .B(n318), .Z(n317) );
  NANDN U347 ( .A(n318), .B(A[227]), .Z(n315) );
  XOR U348 ( .A(n318), .B(n319), .Z(SUM[227]) );
  XNOR U349 ( .A(B[227]), .B(A[227]), .Z(n319) );
  AND U350 ( .A(n320), .B(n321), .Z(n318) );
  NAND U351 ( .A(B[226]), .B(n322), .Z(n321) );
  NANDN U352 ( .A(A[226]), .B(n323), .Z(n322) );
  NANDN U353 ( .A(n323), .B(A[226]), .Z(n320) );
  XOR U354 ( .A(n323), .B(n324), .Z(SUM[226]) );
  XNOR U355 ( .A(B[226]), .B(A[226]), .Z(n324) );
  AND U356 ( .A(n325), .B(n326), .Z(n323) );
  NAND U357 ( .A(B[225]), .B(n327), .Z(n326) );
  NANDN U358 ( .A(A[225]), .B(n328), .Z(n327) );
  NANDN U359 ( .A(n328), .B(A[225]), .Z(n325) );
  XOR U360 ( .A(n328), .B(n329), .Z(SUM[225]) );
  XNOR U361 ( .A(B[225]), .B(A[225]), .Z(n329) );
  AND U362 ( .A(n330), .B(n331), .Z(n328) );
  NAND U363 ( .A(B[224]), .B(n332), .Z(n331) );
  NANDN U364 ( .A(A[224]), .B(n333), .Z(n332) );
  NANDN U365 ( .A(n333), .B(A[224]), .Z(n330) );
  XOR U366 ( .A(n333), .B(n334), .Z(SUM[224]) );
  XNOR U367 ( .A(B[224]), .B(A[224]), .Z(n334) );
  AND U368 ( .A(n335), .B(n336), .Z(n333) );
  NAND U369 ( .A(B[223]), .B(n337), .Z(n336) );
  NANDN U370 ( .A(A[223]), .B(n338), .Z(n337) );
  NANDN U371 ( .A(n338), .B(A[223]), .Z(n335) );
  XOR U372 ( .A(n338), .B(n339), .Z(SUM[223]) );
  XNOR U373 ( .A(B[223]), .B(A[223]), .Z(n339) );
  AND U374 ( .A(n340), .B(n341), .Z(n338) );
  NAND U375 ( .A(B[222]), .B(n342), .Z(n341) );
  NANDN U376 ( .A(A[222]), .B(n343), .Z(n342) );
  NANDN U377 ( .A(n343), .B(A[222]), .Z(n340) );
  XOR U378 ( .A(n343), .B(n344), .Z(SUM[222]) );
  XNOR U379 ( .A(B[222]), .B(A[222]), .Z(n344) );
  AND U380 ( .A(n345), .B(n346), .Z(n343) );
  NAND U381 ( .A(B[221]), .B(n347), .Z(n346) );
  NANDN U382 ( .A(A[221]), .B(n348), .Z(n347) );
  NANDN U383 ( .A(n348), .B(A[221]), .Z(n345) );
  XOR U384 ( .A(n348), .B(n349), .Z(SUM[221]) );
  XNOR U385 ( .A(B[221]), .B(A[221]), .Z(n349) );
  AND U386 ( .A(n350), .B(n351), .Z(n348) );
  NAND U387 ( .A(B[220]), .B(n352), .Z(n351) );
  NANDN U388 ( .A(A[220]), .B(n353), .Z(n352) );
  NANDN U389 ( .A(n353), .B(A[220]), .Z(n350) );
  XOR U390 ( .A(n353), .B(n354), .Z(SUM[220]) );
  XNOR U391 ( .A(B[220]), .B(A[220]), .Z(n354) );
  AND U392 ( .A(n355), .B(n356), .Z(n353) );
  NAND U393 ( .A(B[219]), .B(n357), .Z(n356) );
  NANDN U394 ( .A(A[219]), .B(n358), .Z(n357) );
  NANDN U395 ( .A(n358), .B(A[219]), .Z(n355) );
  XOR U396 ( .A(n359), .B(n360), .Z(SUM[21]) );
  XNOR U397 ( .A(B[21]), .B(A[21]), .Z(n360) );
  XOR U398 ( .A(n358), .B(n361), .Z(SUM[219]) );
  XNOR U399 ( .A(B[219]), .B(A[219]), .Z(n361) );
  AND U400 ( .A(n362), .B(n363), .Z(n358) );
  NAND U401 ( .A(B[218]), .B(n364), .Z(n363) );
  NANDN U402 ( .A(A[218]), .B(n365), .Z(n364) );
  NANDN U403 ( .A(n365), .B(A[218]), .Z(n362) );
  XOR U404 ( .A(n365), .B(n366), .Z(SUM[218]) );
  XNOR U405 ( .A(B[218]), .B(A[218]), .Z(n366) );
  AND U406 ( .A(n367), .B(n368), .Z(n365) );
  NAND U407 ( .A(B[217]), .B(n369), .Z(n368) );
  NANDN U408 ( .A(A[217]), .B(n370), .Z(n369) );
  NANDN U409 ( .A(n370), .B(A[217]), .Z(n367) );
  XOR U410 ( .A(n370), .B(n371), .Z(SUM[217]) );
  XNOR U411 ( .A(B[217]), .B(A[217]), .Z(n371) );
  AND U412 ( .A(n372), .B(n373), .Z(n370) );
  NAND U413 ( .A(B[216]), .B(n374), .Z(n373) );
  NANDN U414 ( .A(A[216]), .B(n375), .Z(n374) );
  NANDN U415 ( .A(n375), .B(A[216]), .Z(n372) );
  XOR U416 ( .A(n375), .B(n376), .Z(SUM[216]) );
  XNOR U417 ( .A(B[216]), .B(A[216]), .Z(n376) );
  AND U418 ( .A(n377), .B(n378), .Z(n375) );
  NAND U419 ( .A(B[215]), .B(n379), .Z(n378) );
  NANDN U420 ( .A(A[215]), .B(n380), .Z(n379) );
  NANDN U421 ( .A(n380), .B(A[215]), .Z(n377) );
  XOR U422 ( .A(n380), .B(n381), .Z(SUM[215]) );
  XNOR U423 ( .A(B[215]), .B(A[215]), .Z(n381) );
  AND U424 ( .A(n382), .B(n383), .Z(n380) );
  NAND U425 ( .A(B[214]), .B(n384), .Z(n383) );
  NANDN U426 ( .A(A[214]), .B(n385), .Z(n384) );
  NANDN U427 ( .A(n385), .B(A[214]), .Z(n382) );
  XOR U428 ( .A(n385), .B(n386), .Z(SUM[214]) );
  XNOR U429 ( .A(B[214]), .B(A[214]), .Z(n386) );
  AND U430 ( .A(n387), .B(n388), .Z(n385) );
  NAND U431 ( .A(B[213]), .B(n389), .Z(n388) );
  NANDN U432 ( .A(A[213]), .B(n390), .Z(n389) );
  NANDN U433 ( .A(n390), .B(A[213]), .Z(n387) );
  XOR U434 ( .A(n390), .B(n391), .Z(SUM[213]) );
  XNOR U435 ( .A(B[213]), .B(A[213]), .Z(n391) );
  AND U436 ( .A(n392), .B(n393), .Z(n390) );
  NAND U437 ( .A(B[212]), .B(n394), .Z(n393) );
  NANDN U438 ( .A(A[212]), .B(n395), .Z(n394) );
  NANDN U439 ( .A(n395), .B(A[212]), .Z(n392) );
  XOR U440 ( .A(n395), .B(n396), .Z(SUM[212]) );
  XNOR U441 ( .A(B[212]), .B(A[212]), .Z(n396) );
  AND U442 ( .A(n397), .B(n398), .Z(n395) );
  NAND U443 ( .A(B[211]), .B(n399), .Z(n398) );
  NANDN U444 ( .A(A[211]), .B(n400), .Z(n399) );
  NANDN U445 ( .A(n400), .B(A[211]), .Z(n397) );
  XOR U446 ( .A(n400), .B(n401), .Z(SUM[211]) );
  XNOR U447 ( .A(B[211]), .B(A[211]), .Z(n401) );
  AND U448 ( .A(n402), .B(n403), .Z(n400) );
  NAND U449 ( .A(B[210]), .B(n404), .Z(n403) );
  NANDN U450 ( .A(A[210]), .B(n405), .Z(n404) );
  NANDN U451 ( .A(n405), .B(A[210]), .Z(n402) );
  XOR U452 ( .A(n405), .B(n406), .Z(SUM[210]) );
  XNOR U453 ( .A(B[210]), .B(A[210]), .Z(n406) );
  AND U454 ( .A(n407), .B(n408), .Z(n405) );
  NAND U455 ( .A(B[209]), .B(n409), .Z(n408) );
  NANDN U456 ( .A(A[209]), .B(n410), .Z(n409) );
  NANDN U457 ( .A(n410), .B(A[209]), .Z(n407) );
  XOR U458 ( .A(n411), .B(n412), .Z(SUM[20]) );
  XNOR U459 ( .A(B[20]), .B(A[20]), .Z(n412) );
  XOR U460 ( .A(n410), .B(n413), .Z(SUM[209]) );
  XNOR U461 ( .A(B[209]), .B(A[209]), .Z(n413) );
  AND U462 ( .A(n414), .B(n415), .Z(n410) );
  NAND U463 ( .A(B[208]), .B(n416), .Z(n415) );
  NANDN U464 ( .A(A[208]), .B(n417), .Z(n416) );
  NANDN U465 ( .A(n417), .B(A[208]), .Z(n414) );
  XOR U466 ( .A(n417), .B(n418), .Z(SUM[208]) );
  XNOR U467 ( .A(B[208]), .B(A[208]), .Z(n418) );
  AND U468 ( .A(n419), .B(n420), .Z(n417) );
  NAND U469 ( .A(B[207]), .B(n421), .Z(n420) );
  NANDN U470 ( .A(A[207]), .B(n422), .Z(n421) );
  NANDN U471 ( .A(n422), .B(A[207]), .Z(n419) );
  XOR U472 ( .A(n422), .B(n423), .Z(SUM[207]) );
  XNOR U473 ( .A(B[207]), .B(A[207]), .Z(n423) );
  AND U474 ( .A(n424), .B(n425), .Z(n422) );
  NAND U475 ( .A(B[206]), .B(n426), .Z(n425) );
  NANDN U476 ( .A(A[206]), .B(n427), .Z(n426) );
  NANDN U477 ( .A(n427), .B(A[206]), .Z(n424) );
  XOR U478 ( .A(n427), .B(n428), .Z(SUM[206]) );
  XNOR U479 ( .A(B[206]), .B(A[206]), .Z(n428) );
  AND U480 ( .A(n429), .B(n430), .Z(n427) );
  NAND U481 ( .A(B[205]), .B(n431), .Z(n430) );
  NANDN U482 ( .A(A[205]), .B(n432), .Z(n431) );
  NANDN U483 ( .A(n432), .B(A[205]), .Z(n429) );
  XOR U484 ( .A(n432), .B(n433), .Z(SUM[205]) );
  XNOR U485 ( .A(B[205]), .B(A[205]), .Z(n433) );
  AND U486 ( .A(n434), .B(n435), .Z(n432) );
  NAND U487 ( .A(B[204]), .B(n436), .Z(n435) );
  NANDN U488 ( .A(A[204]), .B(n437), .Z(n436) );
  NANDN U489 ( .A(n437), .B(A[204]), .Z(n434) );
  XOR U490 ( .A(n437), .B(n438), .Z(SUM[204]) );
  XNOR U491 ( .A(B[204]), .B(A[204]), .Z(n438) );
  AND U492 ( .A(n439), .B(n440), .Z(n437) );
  NAND U493 ( .A(B[203]), .B(n441), .Z(n440) );
  NANDN U494 ( .A(A[203]), .B(n442), .Z(n441) );
  NANDN U495 ( .A(n442), .B(A[203]), .Z(n439) );
  XOR U496 ( .A(n442), .B(n443), .Z(SUM[203]) );
  XNOR U497 ( .A(B[203]), .B(A[203]), .Z(n443) );
  AND U498 ( .A(n444), .B(n445), .Z(n442) );
  NAND U499 ( .A(B[202]), .B(n446), .Z(n445) );
  NANDN U500 ( .A(A[202]), .B(n447), .Z(n446) );
  NANDN U501 ( .A(n447), .B(A[202]), .Z(n444) );
  XOR U502 ( .A(n447), .B(n448), .Z(SUM[202]) );
  XNOR U503 ( .A(B[202]), .B(A[202]), .Z(n448) );
  AND U504 ( .A(n449), .B(n450), .Z(n447) );
  NAND U505 ( .A(B[201]), .B(n451), .Z(n450) );
  NANDN U506 ( .A(A[201]), .B(n452), .Z(n451) );
  NANDN U507 ( .A(n452), .B(A[201]), .Z(n449) );
  XOR U508 ( .A(n452), .B(n453), .Z(SUM[201]) );
  XNOR U509 ( .A(B[201]), .B(A[201]), .Z(n453) );
  AND U510 ( .A(n454), .B(n455), .Z(n452) );
  NAND U511 ( .A(B[200]), .B(n456), .Z(n455) );
  NANDN U512 ( .A(A[200]), .B(n457), .Z(n456) );
  NANDN U513 ( .A(n457), .B(A[200]), .Z(n454) );
  XOR U514 ( .A(n457), .B(n458), .Z(SUM[200]) );
  XNOR U515 ( .A(B[200]), .B(A[200]), .Z(n458) );
  AND U516 ( .A(n459), .B(n460), .Z(n457) );
  NAND U517 ( .A(B[199]), .B(n461), .Z(n460) );
  NANDN U518 ( .A(A[199]), .B(n462), .Z(n461) );
  NANDN U519 ( .A(n462), .B(A[199]), .Z(n459) );
  XOR U520 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  XOR U521 ( .A(n463), .B(n464), .Z(SUM[19]) );
  XNOR U522 ( .A(B[19]), .B(A[19]), .Z(n464) );
  XOR U523 ( .A(n462), .B(n465), .Z(SUM[199]) );
  XNOR U524 ( .A(B[199]), .B(A[199]), .Z(n465) );
  AND U525 ( .A(n466), .B(n467), .Z(n462) );
  NAND U526 ( .A(B[198]), .B(n468), .Z(n467) );
  NANDN U527 ( .A(A[198]), .B(n469), .Z(n468) );
  NANDN U528 ( .A(n469), .B(A[198]), .Z(n466) );
  XOR U529 ( .A(n469), .B(n470), .Z(SUM[198]) );
  XNOR U530 ( .A(B[198]), .B(A[198]), .Z(n470) );
  AND U531 ( .A(n471), .B(n472), .Z(n469) );
  NAND U532 ( .A(B[197]), .B(n473), .Z(n472) );
  NANDN U533 ( .A(A[197]), .B(n474), .Z(n473) );
  NANDN U534 ( .A(n474), .B(A[197]), .Z(n471) );
  XOR U535 ( .A(n474), .B(n475), .Z(SUM[197]) );
  XNOR U536 ( .A(B[197]), .B(A[197]), .Z(n475) );
  AND U537 ( .A(n476), .B(n477), .Z(n474) );
  NAND U538 ( .A(B[196]), .B(n478), .Z(n477) );
  NANDN U539 ( .A(A[196]), .B(n479), .Z(n478) );
  NANDN U540 ( .A(n479), .B(A[196]), .Z(n476) );
  XOR U541 ( .A(n479), .B(n480), .Z(SUM[196]) );
  XNOR U542 ( .A(B[196]), .B(A[196]), .Z(n480) );
  AND U543 ( .A(n481), .B(n482), .Z(n479) );
  NAND U544 ( .A(B[195]), .B(n483), .Z(n482) );
  NANDN U545 ( .A(A[195]), .B(n484), .Z(n483) );
  NANDN U546 ( .A(n484), .B(A[195]), .Z(n481) );
  XOR U547 ( .A(n484), .B(n485), .Z(SUM[195]) );
  XNOR U548 ( .A(B[195]), .B(A[195]), .Z(n485) );
  AND U549 ( .A(n486), .B(n487), .Z(n484) );
  NAND U550 ( .A(B[194]), .B(n488), .Z(n487) );
  NANDN U551 ( .A(A[194]), .B(n489), .Z(n488) );
  NANDN U552 ( .A(n489), .B(A[194]), .Z(n486) );
  XOR U553 ( .A(n489), .B(n490), .Z(SUM[194]) );
  XNOR U554 ( .A(B[194]), .B(A[194]), .Z(n490) );
  AND U555 ( .A(n491), .B(n492), .Z(n489) );
  NAND U556 ( .A(B[193]), .B(n493), .Z(n492) );
  NANDN U557 ( .A(A[193]), .B(n494), .Z(n493) );
  NANDN U558 ( .A(n494), .B(A[193]), .Z(n491) );
  XOR U559 ( .A(n494), .B(n495), .Z(SUM[193]) );
  XNOR U560 ( .A(B[193]), .B(A[193]), .Z(n495) );
  AND U561 ( .A(n496), .B(n497), .Z(n494) );
  NAND U562 ( .A(B[192]), .B(n498), .Z(n497) );
  NANDN U563 ( .A(A[192]), .B(n499), .Z(n498) );
  NANDN U564 ( .A(n499), .B(A[192]), .Z(n496) );
  XOR U565 ( .A(n499), .B(n500), .Z(SUM[192]) );
  XNOR U566 ( .A(B[192]), .B(A[192]), .Z(n500) );
  AND U567 ( .A(n501), .B(n502), .Z(n499) );
  NAND U568 ( .A(B[191]), .B(n503), .Z(n502) );
  NANDN U569 ( .A(A[191]), .B(n504), .Z(n503) );
  NANDN U570 ( .A(n504), .B(A[191]), .Z(n501) );
  XOR U571 ( .A(n504), .B(n505), .Z(SUM[191]) );
  XNOR U572 ( .A(B[191]), .B(A[191]), .Z(n505) );
  AND U573 ( .A(n506), .B(n507), .Z(n504) );
  NAND U574 ( .A(B[190]), .B(n508), .Z(n507) );
  NANDN U575 ( .A(A[190]), .B(n509), .Z(n508) );
  NANDN U576 ( .A(n509), .B(A[190]), .Z(n506) );
  XOR U577 ( .A(n509), .B(n510), .Z(SUM[190]) );
  XNOR U578 ( .A(B[190]), .B(A[190]), .Z(n510) );
  AND U579 ( .A(n511), .B(n512), .Z(n509) );
  NAND U580 ( .A(B[189]), .B(n513), .Z(n512) );
  NANDN U581 ( .A(A[189]), .B(n514), .Z(n513) );
  NANDN U582 ( .A(n514), .B(A[189]), .Z(n511) );
  XOR U583 ( .A(n515), .B(n516), .Z(SUM[18]) );
  XNOR U584 ( .A(B[18]), .B(A[18]), .Z(n516) );
  XOR U585 ( .A(n514), .B(n517), .Z(SUM[189]) );
  XNOR U586 ( .A(B[189]), .B(A[189]), .Z(n517) );
  AND U587 ( .A(n518), .B(n519), .Z(n514) );
  NAND U588 ( .A(B[188]), .B(n520), .Z(n519) );
  NANDN U589 ( .A(A[188]), .B(n521), .Z(n520) );
  NANDN U590 ( .A(n521), .B(A[188]), .Z(n518) );
  XOR U591 ( .A(n521), .B(n522), .Z(SUM[188]) );
  XNOR U592 ( .A(B[188]), .B(A[188]), .Z(n522) );
  AND U593 ( .A(n523), .B(n524), .Z(n521) );
  NAND U594 ( .A(B[187]), .B(n525), .Z(n524) );
  NANDN U595 ( .A(A[187]), .B(n526), .Z(n525) );
  NANDN U596 ( .A(n526), .B(A[187]), .Z(n523) );
  XOR U597 ( .A(n526), .B(n527), .Z(SUM[187]) );
  XNOR U598 ( .A(B[187]), .B(A[187]), .Z(n527) );
  AND U599 ( .A(n528), .B(n529), .Z(n526) );
  NAND U600 ( .A(B[186]), .B(n530), .Z(n529) );
  NANDN U601 ( .A(A[186]), .B(n531), .Z(n530) );
  NANDN U602 ( .A(n531), .B(A[186]), .Z(n528) );
  XOR U603 ( .A(n531), .B(n532), .Z(SUM[186]) );
  XNOR U604 ( .A(B[186]), .B(A[186]), .Z(n532) );
  AND U605 ( .A(n533), .B(n534), .Z(n531) );
  NAND U606 ( .A(B[185]), .B(n535), .Z(n534) );
  NANDN U607 ( .A(A[185]), .B(n536), .Z(n535) );
  NANDN U608 ( .A(n536), .B(A[185]), .Z(n533) );
  XOR U609 ( .A(n536), .B(n537), .Z(SUM[185]) );
  XNOR U610 ( .A(B[185]), .B(A[185]), .Z(n537) );
  AND U611 ( .A(n538), .B(n539), .Z(n536) );
  NAND U612 ( .A(B[184]), .B(n540), .Z(n539) );
  NANDN U613 ( .A(A[184]), .B(n541), .Z(n540) );
  NANDN U614 ( .A(n541), .B(A[184]), .Z(n538) );
  XOR U615 ( .A(n541), .B(n542), .Z(SUM[184]) );
  XNOR U616 ( .A(B[184]), .B(A[184]), .Z(n542) );
  AND U617 ( .A(n543), .B(n544), .Z(n541) );
  NAND U618 ( .A(B[183]), .B(n545), .Z(n544) );
  NANDN U619 ( .A(A[183]), .B(n546), .Z(n545) );
  NANDN U620 ( .A(n546), .B(A[183]), .Z(n543) );
  XOR U621 ( .A(n546), .B(n547), .Z(SUM[183]) );
  XNOR U622 ( .A(B[183]), .B(A[183]), .Z(n547) );
  AND U623 ( .A(n548), .B(n549), .Z(n546) );
  NAND U624 ( .A(B[182]), .B(n550), .Z(n549) );
  NANDN U625 ( .A(A[182]), .B(n551), .Z(n550) );
  NANDN U626 ( .A(n551), .B(A[182]), .Z(n548) );
  XOR U627 ( .A(n551), .B(n552), .Z(SUM[182]) );
  XNOR U628 ( .A(B[182]), .B(A[182]), .Z(n552) );
  AND U629 ( .A(n553), .B(n554), .Z(n551) );
  NAND U630 ( .A(B[181]), .B(n555), .Z(n554) );
  NANDN U631 ( .A(A[181]), .B(n556), .Z(n555) );
  NANDN U632 ( .A(n556), .B(A[181]), .Z(n553) );
  XOR U633 ( .A(n556), .B(n557), .Z(SUM[181]) );
  XNOR U634 ( .A(B[181]), .B(A[181]), .Z(n557) );
  AND U635 ( .A(n558), .B(n559), .Z(n556) );
  NAND U636 ( .A(B[180]), .B(n560), .Z(n559) );
  NANDN U637 ( .A(A[180]), .B(n561), .Z(n560) );
  NANDN U638 ( .A(n561), .B(A[180]), .Z(n558) );
  XOR U639 ( .A(n561), .B(n562), .Z(SUM[180]) );
  XNOR U640 ( .A(B[180]), .B(A[180]), .Z(n562) );
  AND U641 ( .A(n563), .B(n564), .Z(n561) );
  NAND U642 ( .A(B[179]), .B(n565), .Z(n564) );
  NANDN U643 ( .A(A[179]), .B(n566), .Z(n565) );
  NANDN U644 ( .A(n566), .B(A[179]), .Z(n563) );
  XOR U645 ( .A(n567), .B(n568), .Z(SUM[17]) );
  XNOR U646 ( .A(B[17]), .B(A[17]), .Z(n568) );
  XOR U647 ( .A(n566), .B(n569), .Z(SUM[179]) );
  XNOR U648 ( .A(B[179]), .B(A[179]), .Z(n569) );
  AND U649 ( .A(n570), .B(n571), .Z(n566) );
  NAND U650 ( .A(B[178]), .B(n572), .Z(n571) );
  NANDN U651 ( .A(A[178]), .B(n573), .Z(n572) );
  NANDN U652 ( .A(n573), .B(A[178]), .Z(n570) );
  XOR U653 ( .A(n573), .B(n574), .Z(SUM[178]) );
  XNOR U654 ( .A(B[178]), .B(A[178]), .Z(n574) );
  AND U655 ( .A(n575), .B(n576), .Z(n573) );
  NAND U656 ( .A(B[177]), .B(n577), .Z(n576) );
  NANDN U657 ( .A(A[177]), .B(n578), .Z(n577) );
  NANDN U658 ( .A(n578), .B(A[177]), .Z(n575) );
  XOR U659 ( .A(n578), .B(n579), .Z(SUM[177]) );
  XNOR U660 ( .A(B[177]), .B(A[177]), .Z(n579) );
  AND U661 ( .A(n580), .B(n581), .Z(n578) );
  NAND U662 ( .A(B[176]), .B(n582), .Z(n581) );
  NANDN U663 ( .A(A[176]), .B(n583), .Z(n582) );
  NANDN U664 ( .A(n583), .B(A[176]), .Z(n580) );
  XOR U665 ( .A(n583), .B(n584), .Z(SUM[176]) );
  XNOR U666 ( .A(B[176]), .B(A[176]), .Z(n584) );
  AND U667 ( .A(n585), .B(n586), .Z(n583) );
  NAND U668 ( .A(B[175]), .B(n587), .Z(n586) );
  NANDN U669 ( .A(A[175]), .B(n588), .Z(n587) );
  NANDN U670 ( .A(n588), .B(A[175]), .Z(n585) );
  XOR U671 ( .A(n588), .B(n589), .Z(SUM[175]) );
  XNOR U672 ( .A(B[175]), .B(A[175]), .Z(n589) );
  AND U673 ( .A(n590), .B(n591), .Z(n588) );
  NAND U674 ( .A(B[174]), .B(n592), .Z(n591) );
  NANDN U675 ( .A(A[174]), .B(n593), .Z(n592) );
  NANDN U676 ( .A(n593), .B(A[174]), .Z(n590) );
  XOR U677 ( .A(n593), .B(n594), .Z(SUM[174]) );
  XNOR U678 ( .A(B[174]), .B(A[174]), .Z(n594) );
  AND U679 ( .A(n595), .B(n596), .Z(n593) );
  NAND U680 ( .A(B[173]), .B(n597), .Z(n596) );
  NANDN U681 ( .A(A[173]), .B(n598), .Z(n597) );
  NANDN U682 ( .A(n598), .B(A[173]), .Z(n595) );
  XOR U683 ( .A(n598), .B(n599), .Z(SUM[173]) );
  XNOR U684 ( .A(B[173]), .B(A[173]), .Z(n599) );
  AND U685 ( .A(n600), .B(n601), .Z(n598) );
  NAND U686 ( .A(B[172]), .B(n602), .Z(n601) );
  NANDN U687 ( .A(A[172]), .B(n603), .Z(n602) );
  NANDN U688 ( .A(n603), .B(A[172]), .Z(n600) );
  XOR U689 ( .A(n603), .B(n604), .Z(SUM[172]) );
  XNOR U690 ( .A(B[172]), .B(A[172]), .Z(n604) );
  AND U691 ( .A(n605), .B(n606), .Z(n603) );
  NAND U692 ( .A(B[171]), .B(n607), .Z(n606) );
  NANDN U693 ( .A(A[171]), .B(n608), .Z(n607) );
  NANDN U694 ( .A(n608), .B(A[171]), .Z(n605) );
  XOR U695 ( .A(n608), .B(n609), .Z(SUM[171]) );
  XNOR U696 ( .A(B[171]), .B(A[171]), .Z(n609) );
  AND U697 ( .A(n610), .B(n611), .Z(n608) );
  NAND U698 ( .A(B[170]), .B(n612), .Z(n611) );
  NANDN U699 ( .A(A[170]), .B(n613), .Z(n612) );
  NANDN U700 ( .A(n613), .B(A[170]), .Z(n610) );
  XOR U701 ( .A(n613), .B(n614), .Z(SUM[170]) );
  XNOR U702 ( .A(B[170]), .B(A[170]), .Z(n614) );
  AND U703 ( .A(n615), .B(n616), .Z(n613) );
  NAND U704 ( .A(B[169]), .B(n617), .Z(n616) );
  NANDN U705 ( .A(A[169]), .B(n618), .Z(n617) );
  NANDN U706 ( .A(n618), .B(A[169]), .Z(n615) );
  XOR U707 ( .A(n619), .B(n620), .Z(SUM[16]) );
  XNOR U708 ( .A(B[16]), .B(A[16]), .Z(n620) );
  XOR U709 ( .A(n618), .B(n621), .Z(SUM[169]) );
  XNOR U710 ( .A(B[169]), .B(A[169]), .Z(n621) );
  AND U711 ( .A(n622), .B(n623), .Z(n618) );
  NAND U712 ( .A(B[168]), .B(n624), .Z(n623) );
  NANDN U713 ( .A(A[168]), .B(n625), .Z(n624) );
  NANDN U714 ( .A(n625), .B(A[168]), .Z(n622) );
  XOR U715 ( .A(n625), .B(n626), .Z(SUM[168]) );
  XNOR U716 ( .A(B[168]), .B(A[168]), .Z(n626) );
  AND U717 ( .A(n627), .B(n628), .Z(n625) );
  NAND U718 ( .A(B[167]), .B(n629), .Z(n628) );
  NANDN U719 ( .A(A[167]), .B(n630), .Z(n629) );
  NANDN U720 ( .A(n630), .B(A[167]), .Z(n627) );
  XOR U721 ( .A(n630), .B(n631), .Z(SUM[167]) );
  XNOR U722 ( .A(B[167]), .B(A[167]), .Z(n631) );
  AND U723 ( .A(n632), .B(n633), .Z(n630) );
  NAND U724 ( .A(B[166]), .B(n634), .Z(n633) );
  NANDN U725 ( .A(A[166]), .B(n635), .Z(n634) );
  NANDN U726 ( .A(n635), .B(A[166]), .Z(n632) );
  XOR U727 ( .A(n635), .B(n636), .Z(SUM[166]) );
  XNOR U728 ( .A(B[166]), .B(A[166]), .Z(n636) );
  AND U729 ( .A(n637), .B(n638), .Z(n635) );
  NAND U730 ( .A(B[165]), .B(n639), .Z(n638) );
  NANDN U731 ( .A(A[165]), .B(n640), .Z(n639) );
  NANDN U732 ( .A(n640), .B(A[165]), .Z(n637) );
  XOR U733 ( .A(n640), .B(n641), .Z(SUM[165]) );
  XNOR U734 ( .A(B[165]), .B(A[165]), .Z(n641) );
  AND U735 ( .A(n642), .B(n643), .Z(n640) );
  NAND U736 ( .A(B[164]), .B(n644), .Z(n643) );
  NANDN U737 ( .A(A[164]), .B(n645), .Z(n644) );
  NANDN U738 ( .A(n645), .B(A[164]), .Z(n642) );
  XOR U739 ( .A(n645), .B(n646), .Z(SUM[164]) );
  XNOR U740 ( .A(B[164]), .B(A[164]), .Z(n646) );
  AND U741 ( .A(n647), .B(n648), .Z(n645) );
  NAND U742 ( .A(B[163]), .B(n649), .Z(n648) );
  NANDN U743 ( .A(A[163]), .B(n650), .Z(n649) );
  NANDN U744 ( .A(n650), .B(A[163]), .Z(n647) );
  XOR U745 ( .A(n650), .B(n651), .Z(SUM[163]) );
  XNOR U746 ( .A(B[163]), .B(A[163]), .Z(n651) );
  AND U747 ( .A(n652), .B(n653), .Z(n650) );
  NAND U748 ( .A(B[162]), .B(n654), .Z(n653) );
  NANDN U749 ( .A(A[162]), .B(n655), .Z(n654) );
  NANDN U750 ( .A(n655), .B(A[162]), .Z(n652) );
  XOR U751 ( .A(n655), .B(n656), .Z(SUM[162]) );
  XNOR U752 ( .A(B[162]), .B(A[162]), .Z(n656) );
  AND U753 ( .A(n657), .B(n658), .Z(n655) );
  NAND U754 ( .A(B[161]), .B(n659), .Z(n658) );
  NANDN U755 ( .A(A[161]), .B(n660), .Z(n659) );
  NANDN U756 ( .A(n660), .B(A[161]), .Z(n657) );
  XOR U757 ( .A(n660), .B(n661), .Z(SUM[161]) );
  XNOR U758 ( .A(B[161]), .B(A[161]), .Z(n661) );
  AND U759 ( .A(n662), .B(n663), .Z(n660) );
  NAND U760 ( .A(B[160]), .B(n664), .Z(n663) );
  NANDN U761 ( .A(A[160]), .B(n665), .Z(n664) );
  NANDN U762 ( .A(n665), .B(A[160]), .Z(n662) );
  XOR U763 ( .A(n665), .B(n666), .Z(SUM[160]) );
  XNOR U764 ( .A(B[160]), .B(A[160]), .Z(n666) );
  AND U765 ( .A(n667), .B(n668), .Z(n665) );
  NAND U766 ( .A(B[159]), .B(n669), .Z(n668) );
  NANDN U767 ( .A(A[159]), .B(n670), .Z(n669) );
  NANDN U768 ( .A(n670), .B(A[159]), .Z(n667) );
  XOR U769 ( .A(n671), .B(n672), .Z(SUM[15]) );
  XNOR U770 ( .A(B[15]), .B(A[15]), .Z(n672) );
  XOR U771 ( .A(n670), .B(n673), .Z(SUM[159]) );
  XNOR U772 ( .A(B[159]), .B(A[159]), .Z(n673) );
  AND U773 ( .A(n674), .B(n675), .Z(n670) );
  NAND U774 ( .A(B[158]), .B(n676), .Z(n675) );
  NANDN U775 ( .A(A[158]), .B(n677), .Z(n676) );
  NANDN U776 ( .A(n677), .B(A[158]), .Z(n674) );
  XOR U777 ( .A(n677), .B(n678), .Z(SUM[158]) );
  XNOR U778 ( .A(B[158]), .B(A[158]), .Z(n678) );
  AND U779 ( .A(n679), .B(n680), .Z(n677) );
  NAND U780 ( .A(B[157]), .B(n681), .Z(n680) );
  NANDN U781 ( .A(A[157]), .B(n682), .Z(n681) );
  NANDN U782 ( .A(n682), .B(A[157]), .Z(n679) );
  XOR U783 ( .A(n682), .B(n683), .Z(SUM[157]) );
  XNOR U784 ( .A(B[157]), .B(A[157]), .Z(n683) );
  AND U785 ( .A(n684), .B(n685), .Z(n682) );
  NAND U786 ( .A(B[156]), .B(n686), .Z(n685) );
  NANDN U787 ( .A(A[156]), .B(n687), .Z(n686) );
  NANDN U788 ( .A(n687), .B(A[156]), .Z(n684) );
  XOR U789 ( .A(n687), .B(n688), .Z(SUM[156]) );
  XNOR U790 ( .A(B[156]), .B(A[156]), .Z(n688) );
  AND U791 ( .A(n689), .B(n690), .Z(n687) );
  NAND U792 ( .A(B[155]), .B(n691), .Z(n690) );
  NANDN U793 ( .A(A[155]), .B(n692), .Z(n691) );
  NANDN U794 ( .A(n692), .B(A[155]), .Z(n689) );
  XOR U795 ( .A(n692), .B(n693), .Z(SUM[155]) );
  XNOR U796 ( .A(B[155]), .B(A[155]), .Z(n693) );
  AND U797 ( .A(n694), .B(n695), .Z(n692) );
  NAND U798 ( .A(B[154]), .B(n696), .Z(n695) );
  NANDN U799 ( .A(A[154]), .B(n697), .Z(n696) );
  NANDN U800 ( .A(n697), .B(A[154]), .Z(n694) );
  XOR U801 ( .A(n697), .B(n698), .Z(SUM[154]) );
  XNOR U802 ( .A(B[154]), .B(A[154]), .Z(n698) );
  AND U803 ( .A(n699), .B(n700), .Z(n697) );
  NAND U804 ( .A(B[153]), .B(n701), .Z(n700) );
  NANDN U805 ( .A(A[153]), .B(n702), .Z(n701) );
  NANDN U806 ( .A(n702), .B(A[153]), .Z(n699) );
  XOR U807 ( .A(n702), .B(n703), .Z(SUM[153]) );
  XNOR U808 ( .A(B[153]), .B(A[153]), .Z(n703) );
  AND U809 ( .A(n704), .B(n705), .Z(n702) );
  NAND U810 ( .A(B[152]), .B(n706), .Z(n705) );
  NANDN U811 ( .A(A[152]), .B(n707), .Z(n706) );
  NANDN U812 ( .A(n707), .B(A[152]), .Z(n704) );
  XOR U813 ( .A(n707), .B(n708), .Z(SUM[152]) );
  XNOR U814 ( .A(B[152]), .B(A[152]), .Z(n708) );
  AND U815 ( .A(n709), .B(n710), .Z(n707) );
  NAND U816 ( .A(B[151]), .B(n711), .Z(n710) );
  NANDN U817 ( .A(A[151]), .B(n712), .Z(n711) );
  NANDN U818 ( .A(n712), .B(A[151]), .Z(n709) );
  XOR U819 ( .A(n712), .B(n713), .Z(SUM[151]) );
  XNOR U820 ( .A(B[151]), .B(A[151]), .Z(n713) );
  AND U821 ( .A(n714), .B(n715), .Z(n712) );
  NAND U822 ( .A(B[150]), .B(n716), .Z(n715) );
  NANDN U823 ( .A(A[150]), .B(n717), .Z(n716) );
  NANDN U824 ( .A(n717), .B(A[150]), .Z(n714) );
  XOR U825 ( .A(n717), .B(n718), .Z(SUM[150]) );
  XNOR U826 ( .A(B[150]), .B(A[150]), .Z(n718) );
  AND U827 ( .A(n719), .B(n720), .Z(n717) );
  NAND U828 ( .A(B[149]), .B(n721), .Z(n720) );
  NANDN U829 ( .A(A[149]), .B(n722), .Z(n721) );
  NANDN U830 ( .A(n722), .B(A[149]), .Z(n719) );
  XOR U831 ( .A(n723), .B(n724), .Z(SUM[14]) );
  XNOR U832 ( .A(B[14]), .B(A[14]), .Z(n724) );
  XOR U833 ( .A(n722), .B(n725), .Z(SUM[149]) );
  XNOR U834 ( .A(B[149]), .B(A[149]), .Z(n725) );
  AND U835 ( .A(n726), .B(n727), .Z(n722) );
  NAND U836 ( .A(B[148]), .B(n728), .Z(n727) );
  NANDN U837 ( .A(A[148]), .B(n729), .Z(n728) );
  NANDN U838 ( .A(n729), .B(A[148]), .Z(n726) );
  XOR U839 ( .A(n729), .B(n730), .Z(SUM[148]) );
  XNOR U840 ( .A(B[148]), .B(A[148]), .Z(n730) );
  AND U841 ( .A(n731), .B(n732), .Z(n729) );
  NAND U842 ( .A(B[147]), .B(n733), .Z(n732) );
  NANDN U843 ( .A(A[147]), .B(n734), .Z(n733) );
  NANDN U844 ( .A(n734), .B(A[147]), .Z(n731) );
  XOR U845 ( .A(n734), .B(n735), .Z(SUM[147]) );
  XNOR U846 ( .A(B[147]), .B(A[147]), .Z(n735) );
  AND U847 ( .A(n736), .B(n737), .Z(n734) );
  NAND U848 ( .A(B[146]), .B(n738), .Z(n737) );
  NANDN U849 ( .A(A[146]), .B(n739), .Z(n738) );
  NANDN U850 ( .A(n739), .B(A[146]), .Z(n736) );
  XOR U851 ( .A(n739), .B(n740), .Z(SUM[146]) );
  XNOR U852 ( .A(B[146]), .B(A[146]), .Z(n740) );
  AND U853 ( .A(n741), .B(n742), .Z(n739) );
  NAND U854 ( .A(B[145]), .B(n743), .Z(n742) );
  NANDN U855 ( .A(A[145]), .B(n744), .Z(n743) );
  NANDN U856 ( .A(n744), .B(A[145]), .Z(n741) );
  XOR U857 ( .A(n744), .B(n745), .Z(SUM[145]) );
  XNOR U858 ( .A(B[145]), .B(A[145]), .Z(n745) );
  AND U859 ( .A(n746), .B(n747), .Z(n744) );
  NAND U860 ( .A(B[144]), .B(n748), .Z(n747) );
  NANDN U861 ( .A(A[144]), .B(n749), .Z(n748) );
  NANDN U862 ( .A(n749), .B(A[144]), .Z(n746) );
  XOR U863 ( .A(n749), .B(n750), .Z(SUM[144]) );
  XNOR U864 ( .A(B[144]), .B(A[144]), .Z(n750) );
  AND U865 ( .A(n751), .B(n752), .Z(n749) );
  NAND U866 ( .A(B[143]), .B(n753), .Z(n752) );
  NANDN U867 ( .A(A[143]), .B(n754), .Z(n753) );
  NANDN U868 ( .A(n754), .B(A[143]), .Z(n751) );
  XOR U869 ( .A(n754), .B(n755), .Z(SUM[143]) );
  XNOR U870 ( .A(B[143]), .B(A[143]), .Z(n755) );
  AND U871 ( .A(n756), .B(n757), .Z(n754) );
  NAND U872 ( .A(B[142]), .B(n758), .Z(n757) );
  NANDN U873 ( .A(A[142]), .B(n759), .Z(n758) );
  NANDN U874 ( .A(n759), .B(A[142]), .Z(n756) );
  XOR U875 ( .A(n759), .B(n760), .Z(SUM[142]) );
  XNOR U876 ( .A(B[142]), .B(A[142]), .Z(n760) );
  AND U877 ( .A(n761), .B(n762), .Z(n759) );
  NAND U878 ( .A(B[141]), .B(n763), .Z(n762) );
  NANDN U879 ( .A(A[141]), .B(n764), .Z(n763) );
  NANDN U880 ( .A(n764), .B(A[141]), .Z(n761) );
  XOR U881 ( .A(n764), .B(n765), .Z(SUM[141]) );
  XNOR U882 ( .A(B[141]), .B(A[141]), .Z(n765) );
  AND U883 ( .A(n766), .B(n767), .Z(n764) );
  NAND U884 ( .A(B[140]), .B(n768), .Z(n767) );
  NANDN U885 ( .A(A[140]), .B(n769), .Z(n768) );
  NANDN U886 ( .A(n769), .B(A[140]), .Z(n766) );
  XOR U887 ( .A(n769), .B(n770), .Z(SUM[140]) );
  XNOR U888 ( .A(B[140]), .B(A[140]), .Z(n770) );
  AND U889 ( .A(n771), .B(n772), .Z(n769) );
  NAND U890 ( .A(B[139]), .B(n773), .Z(n772) );
  NANDN U891 ( .A(A[139]), .B(n774), .Z(n773) );
  NANDN U892 ( .A(n774), .B(A[139]), .Z(n771) );
  XOR U893 ( .A(n775), .B(n776), .Z(SUM[13]) );
  XNOR U894 ( .A(B[13]), .B(A[13]), .Z(n776) );
  XOR U895 ( .A(n774), .B(n777), .Z(SUM[139]) );
  XNOR U896 ( .A(B[139]), .B(A[139]), .Z(n777) );
  AND U897 ( .A(n778), .B(n779), .Z(n774) );
  NAND U898 ( .A(B[138]), .B(n780), .Z(n779) );
  NANDN U899 ( .A(A[138]), .B(n781), .Z(n780) );
  NANDN U900 ( .A(n781), .B(A[138]), .Z(n778) );
  XOR U901 ( .A(n781), .B(n782), .Z(SUM[138]) );
  XNOR U902 ( .A(B[138]), .B(A[138]), .Z(n782) );
  AND U903 ( .A(n783), .B(n784), .Z(n781) );
  NAND U904 ( .A(B[137]), .B(n785), .Z(n784) );
  NANDN U905 ( .A(A[137]), .B(n786), .Z(n785) );
  NANDN U906 ( .A(n786), .B(A[137]), .Z(n783) );
  XOR U907 ( .A(n786), .B(n787), .Z(SUM[137]) );
  XNOR U908 ( .A(B[137]), .B(A[137]), .Z(n787) );
  AND U909 ( .A(n788), .B(n789), .Z(n786) );
  NAND U910 ( .A(B[136]), .B(n790), .Z(n789) );
  NANDN U911 ( .A(A[136]), .B(n791), .Z(n790) );
  NANDN U912 ( .A(n791), .B(A[136]), .Z(n788) );
  XOR U913 ( .A(n791), .B(n792), .Z(SUM[136]) );
  XNOR U914 ( .A(B[136]), .B(A[136]), .Z(n792) );
  AND U915 ( .A(n793), .B(n794), .Z(n791) );
  NAND U916 ( .A(B[135]), .B(n795), .Z(n794) );
  NANDN U917 ( .A(A[135]), .B(n796), .Z(n795) );
  NANDN U918 ( .A(n796), .B(A[135]), .Z(n793) );
  XOR U919 ( .A(n796), .B(n797), .Z(SUM[135]) );
  XNOR U920 ( .A(B[135]), .B(A[135]), .Z(n797) );
  AND U921 ( .A(n798), .B(n799), .Z(n796) );
  NAND U922 ( .A(B[134]), .B(n800), .Z(n799) );
  NANDN U923 ( .A(A[134]), .B(n801), .Z(n800) );
  NANDN U924 ( .A(n801), .B(A[134]), .Z(n798) );
  XOR U925 ( .A(n801), .B(n802), .Z(SUM[134]) );
  XNOR U926 ( .A(B[134]), .B(A[134]), .Z(n802) );
  AND U927 ( .A(n803), .B(n804), .Z(n801) );
  NAND U928 ( .A(B[133]), .B(n805), .Z(n804) );
  NANDN U929 ( .A(A[133]), .B(n806), .Z(n805) );
  NANDN U930 ( .A(n806), .B(A[133]), .Z(n803) );
  XOR U931 ( .A(n806), .B(n807), .Z(SUM[133]) );
  XNOR U932 ( .A(B[133]), .B(A[133]), .Z(n807) );
  AND U933 ( .A(n808), .B(n809), .Z(n806) );
  NAND U934 ( .A(B[132]), .B(n810), .Z(n809) );
  NANDN U935 ( .A(A[132]), .B(n811), .Z(n810) );
  NANDN U936 ( .A(n811), .B(A[132]), .Z(n808) );
  XOR U937 ( .A(n811), .B(n812), .Z(SUM[132]) );
  XNOR U938 ( .A(B[132]), .B(A[132]), .Z(n812) );
  AND U939 ( .A(n813), .B(n814), .Z(n811) );
  NAND U940 ( .A(B[131]), .B(n815), .Z(n814) );
  NANDN U941 ( .A(A[131]), .B(n816), .Z(n815) );
  NANDN U942 ( .A(n816), .B(A[131]), .Z(n813) );
  XOR U943 ( .A(n816), .B(n817), .Z(SUM[131]) );
  XNOR U944 ( .A(B[131]), .B(A[131]), .Z(n817) );
  AND U945 ( .A(n818), .B(n819), .Z(n816) );
  NAND U946 ( .A(B[130]), .B(n820), .Z(n819) );
  NANDN U947 ( .A(A[130]), .B(n821), .Z(n820) );
  NANDN U948 ( .A(n821), .B(A[130]), .Z(n818) );
  XOR U949 ( .A(n821), .B(n822), .Z(SUM[130]) );
  XNOR U950 ( .A(B[130]), .B(A[130]), .Z(n822) );
  AND U951 ( .A(n823), .B(n824), .Z(n821) );
  NAND U952 ( .A(B[129]), .B(n825), .Z(n824) );
  NANDN U953 ( .A(A[129]), .B(n826), .Z(n825) );
  NANDN U954 ( .A(n826), .B(A[129]), .Z(n823) );
  XOR U955 ( .A(n827), .B(n828), .Z(SUM[12]) );
  XNOR U956 ( .A(B[12]), .B(A[12]), .Z(n828) );
  XOR U957 ( .A(n826), .B(n829), .Z(SUM[129]) );
  XNOR U958 ( .A(B[129]), .B(A[129]), .Z(n829) );
  AND U959 ( .A(n830), .B(n831), .Z(n826) );
  NAND U960 ( .A(B[128]), .B(n832), .Z(n831) );
  NANDN U961 ( .A(A[128]), .B(n833), .Z(n832) );
  NANDN U962 ( .A(n833), .B(A[128]), .Z(n830) );
  XOR U963 ( .A(n833), .B(n834), .Z(SUM[128]) );
  XNOR U964 ( .A(B[128]), .B(A[128]), .Z(n834) );
  AND U965 ( .A(n835), .B(n836), .Z(n833) );
  NAND U966 ( .A(B[127]), .B(n837), .Z(n836) );
  NANDN U967 ( .A(A[127]), .B(n838), .Z(n837) );
  NANDN U968 ( .A(n838), .B(A[127]), .Z(n835) );
  XOR U969 ( .A(n838), .B(n839), .Z(SUM[127]) );
  XNOR U970 ( .A(B[127]), .B(A[127]), .Z(n839) );
  AND U971 ( .A(n840), .B(n841), .Z(n838) );
  NAND U972 ( .A(B[126]), .B(n842), .Z(n841) );
  NANDN U973 ( .A(A[126]), .B(n843), .Z(n842) );
  NANDN U974 ( .A(n843), .B(A[126]), .Z(n840) );
  XOR U975 ( .A(n843), .B(n844), .Z(SUM[126]) );
  XNOR U976 ( .A(B[126]), .B(A[126]), .Z(n844) );
  AND U977 ( .A(n845), .B(n846), .Z(n843) );
  NAND U978 ( .A(B[125]), .B(n847), .Z(n846) );
  NANDN U979 ( .A(A[125]), .B(n848), .Z(n847) );
  NANDN U980 ( .A(n848), .B(A[125]), .Z(n845) );
  XOR U981 ( .A(n848), .B(n849), .Z(SUM[125]) );
  XNOR U982 ( .A(B[125]), .B(A[125]), .Z(n849) );
  AND U983 ( .A(n850), .B(n851), .Z(n848) );
  NAND U984 ( .A(B[124]), .B(n852), .Z(n851) );
  NANDN U985 ( .A(A[124]), .B(n853), .Z(n852) );
  NANDN U986 ( .A(n853), .B(A[124]), .Z(n850) );
  XOR U987 ( .A(n853), .B(n854), .Z(SUM[124]) );
  XNOR U988 ( .A(B[124]), .B(A[124]), .Z(n854) );
  AND U989 ( .A(n855), .B(n856), .Z(n853) );
  NAND U990 ( .A(B[123]), .B(n857), .Z(n856) );
  NANDN U991 ( .A(A[123]), .B(n858), .Z(n857) );
  NANDN U992 ( .A(n858), .B(A[123]), .Z(n855) );
  XOR U993 ( .A(n858), .B(n859), .Z(SUM[123]) );
  XNOR U994 ( .A(B[123]), .B(A[123]), .Z(n859) );
  AND U995 ( .A(n860), .B(n861), .Z(n858) );
  NAND U996 ( .A(B[122]), .B(n862), .Z(n861) );
  NANDN U997 ( .A(A[122]), .B(n863), .Z(n862) );
  NANDN U998 ( .A(n863), .B(A[122]), .Z(n860) );
  XOR U999 ( .A(n863), .B(n864), .Z(SUM[122]) );
  XNOR U1000 ( .A(B[122]), .B(A[122]), .Z(n864) );
  AND U1001 ( .A(n865), .B(n866), .Z(n863) );
  NAND U1002 ( .A(B[121]), .B(n867), .Z(n866) );
  NANDN U1003 ( .A(A[121]), .B(n868), .Z(n867) );
  NANDN U1004 ( .A(n868), .B(A[121]), .Z(n865) );
  XOR U1005 ( .A(n868), .B(n869), .Z(SUM[121]) );
  XNOR U1006 ( .A(B[121]), .B(A[121]), .Z(n869) );
  AND U1007 ( .A(n870), .B(n871), .Z(n868) );
  NAND U1008 ( .A(B[120]), .B(n872), .Z(n871) );
  NANDN U1009 ( .A(A[120]), .B(n873), .Z(n872) );
  NANDN U1010 ( .A(n873), .B(A[120]), .Z(n870) );
  XOR U1011 ( .A(n873), .B(n874), .Z(SUM[120]) );
  XNOR U1012 ( .A(B[120]), .B(A[120]), .Z(n874) );
  AND U1013 ( .A(n875), .B(n876), .Z(n873) );
  NAND U1014 ( .A(B[119]), .B(n877), .Z(n876) );
  NANDN U1015 ( .A(A[119]), .B(n878), .Z(n877) );
  NANDN U1016 ( .A(n878), .B(A[119]), .Z(n875) );
  XOR U1017 ( .A(n879), .B(n880), .Z(SUM[11]) );
  XNOR U1018 ( .A(B[11]), .B(A[11]), .Z(n880) );
  XOR U1019 ( .A(n878), .B(n881), .Z(SUM[119]) );
  XNOR U1020 ( .A(B[119]), .B(A[119]), .Z(n881) );
  AND U1021 ( .A(n882), .B(n883), .Z(n878) );
  NAND U1022 ( .A(B[118]), .B(n884), .Z(n883) );
  NANDN U1023 ( .A(A[118]), .B(n885), .Z(n884) );
  NANDN U1024 ( .A(n885), .B(A[118]), .Z(n882) );
  XOR U1025 ( .A(n885), .B(n886), .Z(SUM[118]) );
  XNOR U1026 ( .A(B[118]), .B(A[118]), .Z(n886) );
  AND U1027 ( .A(n887), .B(n888), .Z(n885) );
  NAND U1028 ( .A(B[117]), .B(n889), .Z(n888) );
  NANDN U1029 ( .A(A[117]), .B(n890), .Z(n889) );
  NANDN U1030 ( .A(n890), .B(A[117]), .Z(n887) );
  XOR U1031 ( .A(n890), .B(n891), .Z(SUM[117]) );
  XNOR U1032 ( .A(B[117]), .B(A[117]), .Z(n891) );
  AND U1033 ( .A(n892), .B(n893), .Z(n890) );
  NAND U1034 ( .A(B[116]), .B(n894), .Z(n893) );
  NANDN U1035 ( .A(A[116]), .B(n895), .Z(n894) );
  NANDN U1036 ( .A(n895), .B(A[116]), .Z(n892) );
  XOR U1037 ( .A(n895), .B(n896), .Z(SUM[116]) );
  XNOR U1038 ( .A(B[116]), .B(A[116]), .Z(n896) );
  AND U1039 ( .A(n897), .B(n898), .Z(n895) );
  NAND U1040 ( .A(B[115]), .B(n899), .Z(n898) );
  NANDN U1041 ( .A(A[115]), .B(n900), .Z(n899) );
  NANDN U1042 ( .A(n900), .B(A[115]), .Z(n897) );
  XOR U1043 ( .A(n900), .B(n901), .Z(SUM[115]) );
  XNOR U1044 ( .A(B[115]), .B(A[115]), .Z(n901) );
  AND U1045 ( .A(n902), .B(n903), .Z(n900) );
  NAND U1046 ( .A(B[114]), .B(n904), .Z(n903) );
  NANDN U1047 ( .A(A[114]), .B(n905), .Z(n904) );
  NANDN U1048 ( .A(n905), .B(A[114]), .Z(n902) );
  XOR U1049 ( .A(n905), .B(n906), .Z(SUM[114]) );
  XNOR U1050 ( .A(B[114]), .B(A[114]), .Z(n906) );
  AND U1051 ( .A(n907), .B(n908), .Z(n905) );
  NAND U1052 ( .A(B[113]), .B(n909), .Z(n908) );
  NANDN U1053 ( .A(A[113]), .B(n910), .Z(n909) );
  NANDN U1054 ( .A(n910), .B(A[113]), .Z(n907) );
  XOR U1055 ( .A(n910), .B(n911), .Z(SUM[113]) );
  XNOR U1056 ( .A(B[113]), .B(A[113]), .Z(n911) );
  AND U1057 ( .A(n912), .B(n913), .Z(n910) );
  NAND U1058 ( .A(B[112]), .B(n914), .Z(n913) );
  NANDN U1059 ( .A(A[112]), .B(n915), .Z(n914) );
  NANDN U1060 ( .A(n915), .B(A[112]), .Z(n912) );
  XOR U1061 ( .A(n915), .B(n916), .Z(SUM[112]) );
  XNOR U1062 ( .A(B[112]), .B(A[112]), .Z(n916) );
  AND U1063 ( .A(n917), .B(n918), .Z(n915) );
  NAND U1064 ( .A(B[111]), .B(n919), .Z(n918) );
  NANDN U1065 ( .A(A[111]), .B(n920), .Z(n919) );
  NANDN U1066 ( .A(n920), .B(A[111]), .Z(n917) );
  XOR U1067 ( .A(n920), .B(n921), .Z(SUM[111]) );
  XNOR U1068 ( .A(B[111]), .B(A[111]), .Z(n921) );
  AND U1069 ( .A(n922), .B(n923), .Z(n920) );
  NAND U1070 ( .A(B[110]), .B(n924), .Z(n923) );
  NANDN U1071 ( .A(A[110]), .B(n925), .Z(n924) );
  NANDN U1072 ( .A(n925), .B(A[110]), .Z(n922) );
  XOR U1073 ( .A(n925), .B(n926), .Z(SUM[110]) );
  XNOR U1074 ( .A(B[110]), .B(A[110]), .Z(n926) );
  AND U1075 ( .A(n927), .B(n928), .Z(n925) );
  NAND U1076 ( .A(B[109]), .B(n929), .Z(n928) );
  NANDN U1077 ( .A(A[109]), .B(n930), .Z(n929) );
  NANDN U1078 ( .A(n930), .B(A[109]), .Z(n927) );
  XOR U1079 ( .A(n931), .B(n932), .Z(SUM[10]) );
  XNOR U1080 ( .A(B[10]), .B(A[10]), .Z(n932) );
  XOR U1081 ( .A(n930), .B(n933), .Z(SUM[109]) );
  XNOR U1082 ( .A(B[109]), .B(A[109]), .Z(n933) );
  AND U1083 ( .A(n934), .B(n935), .Z(n930) );
  NAND U1084 ( .A(B[108]), .B(n936), .Z(n935) );
  NANDN U1085 ( .A(A[108]), .B(n937), .Z(n936) );
  NANDN U1086 ( .A(n937), .B(A[108]), .Z(n934) );
  XOR U1087 ( .A(n937), .B(n938), .Z(SUM[108]) );
  XNOR U1088 ( .A(B[108]), .B(A[108]), .Z(n938) );
  AND U1089 ( .A(n939), .B(n940), .Z(n937) );
  NAND U1090 ( .A(B[107]), .B(n941), .Z(n940) );
  NANDN U1091 ( .A(A[107]), .B(n942), .Z(n941) );
  NANDN U1092 ( .A(n942), .B(A[107]), .Z(n939) );
  XOR U1093 ( .A(n942), .B(n943), .Z(SUM[107]) );
  XNOR U1094 ( .A(B[107]), .B(A[107]), .Z(n943) );
  AND U1095 ( .A(n944), .B(n945), .Z(n942) );
  NAND U1096 ( .A(B[106]), .B(n946), .Z(n945) );
  NANDN U1097 ( .A(A[106]), .B(n947), .Z(n946) );
  NANDN U1098 ( .A(n947), .B(A[106]), .Z(n944) );
  XOR U1099 ( .A(n947), .B(n948), .Z(SUM[106]) );
  XNOR U1100 ( .A(B[106]), .B(A[106]), .Z(n948) );
  AND U1101 ( .A(n949), .B(n950), .Z(n947) );
  NAND U1102 ( .A(B[105]), .B(n951), .Z(n950) );
  NANDN U1103 ( .A(A[105]), .B(n952), .Z(n951) );
  NANDN U1104 ( .A(n952), .B(A[105]), .Z(n949) );
  XOR U1105 ( .A(n952), .B(n953), .Z(SUM[105]) );
  XNOR U1106 ( .A(B[105]), .B(A[105]), .Z(n953) );
  AND U1107 ( .A(n954), .B(n955), .Z(n952) );
  NAND U1108 ( .A(B[104]), .B(n956), .Z(n955) );
  NANDN U1109 ( .A(A[104]), .B(n957), .Z(n956) );
  NANDN U1110 ( .A(n957), .B(A[104]), .Z(n954) );
  XOR U1111 ( .A(n957), .B(n958), .Z(SUM[104]) );
  XNOR U1112 ( .A(B[104]), .B(A[104]), .Z(n958) );
  AND U1113 ( .A(n959), .B(n960), .Z(n957) );
  NAND U1114 ( .A(B[103]), .B(n961), .Z(n960) );
  NANDN U1115 ( .A(A[103]), .B(n962), .Z(n961) );
  NANDN U1116 ( .A(n962), .B(A[103]), .Z(n959) );
  XOR U1117 ( .A(n962), .B(n963), .Z(SUM[103]) );
  XNOR U1118 ( .A(B[103]), .B(A[103]), .Z(n963) );
  AND U1119 ( .A(n964), .B(n965), .Z(n962) );
  NAND U1120 ( .A(B[102]), .B(n966), .Z(n965) );
  NANDN U1121 ( .A(A[102]), .B(n967), .Z(n966) );
  NANDN U1122 ( .A(n967), .B(A[102]), .Z(n964) );
  XOR U1123 ( .A(n967), .B(n968), .Z(SUM[102]) );
  XNOR U1124 ( .A(B[102]), .B(A[102]), .Z(n968) );
  AND U1125 ( .A(n969), .B(n970), .Z(n967) );
  NAND U1126 ( .A(B[101]), .B(n971), .Z(n970) );
  NANDN U1127 ( .A(A[101]), .B(n972), .Z(n971) );
  NANDN U1128 ( .A(n972), .B(A[101]), .Z(n969) );
  XOR U1129 ( .A(n972), .B(n973), .Z(SUM[101]) );
  XNOR U1130 ( .A(B[101]), .B(A[101]), .Z(n973) );
  AND U1131 ( .A(n974), .B(n975), .Z(n972) );
  NAND U1132 ( .A(B[100]), .B(n976), .Z(n975) );
  NANDN U1133 ( .A(A[100]), .B(n977), .Z(n976) );
  NANDN U1134 ( .A(n977), .B(A[100]), .Z(n974) );
  XOR U1135 ( .A(n977), .B(n978), .Z(SUM[100]) );
  XNOR U1136 ( .A(B[100]), .B(A[100]), .Z(n978) );
  AND U1137 ( .A(n979), .B(n980), .Z(n977) );
  NAND U1138 ( .A(B[99]), .B(n981), .Z(n980) );
  OR U1139 ( .A(n3), .B(A[99]), .Z(n981) );
  NAND U1140 ( .A(A[99]), .B(n3), .Z(n979) );
  NAND U1141 ( .A(n982), .B(n983), .Z(n3) );
  NAND U1142 ( .A(B[98]), .B(n984), .Z(n983) );
  NANDN U1143 ( .A(A[98]), .B(n5), .Z(n984) );
  NANDN U1144 ( .A(n5), .B(A[98]), .Z(n982) );
  AND U1145 ( .A(n985), .B(n986), .Z(n5) );
  NAND U1146 ( .A(B[97]), .B(n987), .Z(n986) );
  NANDN U1147 ( .A(A[97]), .B(n7), .Z(n987) );
  NANDN U1148 ( .A(n7), .B(A[97]), .Z(n985) );
  AND U1149 ( .A(n988), .B(n989), .Z(n7) );
  NAND U1150 ( .A(B[96]), .B(n990), .Z(n989) );
  NANDN U1151 ( .A(A[96]), .B(n9), .Z(n990) );
  NANDN U1152 ( .A(n9), .B(A[96]), .Z(n988) );
  AND U1153 ( .A(n991), .B(n992), .Z(n9) );
  NAND U1154 ( .A(B[95]), .B(n993), .Z(n992) );
  NANDN U1155 ( .A(A[95]), .B(n11), .Z(n993) );
  NANDN U1156 ( .A(n11), .B(A[95]), .Z(n991) );
  AND U1157 ( .A(n994), .B(n995), .Z(n11) );
  NAND U1158 ( .A(B[94]), .B(n996), .Z(n995) );
  NANDN U1159 ( .A(A[94]), .B(n13), .Z(n996) );
  NANDN U1160 ( .A(n13), .B(A[94]), .Z(n994) );
  AND U1161 ( .A(n997), .B(n998), .Z(n13) );
  NAND U1162 ( .A(B[93]), .B(n999), .Z(n998) );
  NANDN U1163 ( .A(A[93]), .B(n15), .Z(n999) );
  NANDN U1164 ( .A(n15), .B(A[93]), .Z(n997) );
  AND U1165 ( .A(n1000), .B(n1001), .Z(n15) );
  NAND U1166 ( .A(B[92]), .B(n1002), .Z(n1001) );
  NANDN U1167 ( .A(A[92]), .B(n17), .Z(n1002) );
  NANDN U1168 ( .A(n17), .B(A[92]), .Z(n1000) );
  AND U1169 ( .A(n1003), .B(n1004), .Z(n17) );
  NAND U1170 ( .A(B[91]), .B(n1005), .Z(n1004) );
  NANDN U1171 ( .A(A[91]), .B(n19), .Z(n1005) );
  NANDN U1172 ( .A(n19), .B(A[91]), .Z(n1003) );
  AND U1173 ( .A(n1006), .B(n1007), .Z(n19) );
  NAND U1174 ( .A(B[90]), .B(n1008), .Z(n1007) );
  NANDN U1175 ( .A(A[90]), .B(n21), .Z(n1008) );
  NANDN U1176 ( .A(n21), .B(A[90]), .Z(n1006) );
  AND U1177 ( .A(n1009), .B(n1010), .Z(n21) );
  NAND U1178 ( .A(B[89]), .B(n1011), .Z(n1010) );
  NANDN U1179 ( .A(A[89]), .B(n25), .Z(n1011) );
  NANDN U1180 ( .A(n25), .B(A[89]), .Z(n1009) );
  AND U1181 ( .A(n1012), .B(n1013), .Z(n25) );
  NAND U1182 ( .A(B[88]), .B(n1014), .Z(n1013) );
  NANDN U1183 ( .A(A[88]), .B(n27), .Z(n1014) );
  NANDN U1184 ( .A(n27), .B(A[88]), .Z(n1012) );
  AND U1185 ( .A(n1015), .B(n1016), .Z(n27) );
  NAND U1186 ( .A(B[87]), .B(n1017), .Z(n1016) );
  NANDN U1187 ( .A(A[87]), .B(n29), .Z(n1017) );
  NANDN U1188 ( .A(n29), .B(A[87]), .Z(n1015) );
  AND U1189 ( .A(n1018), .B(n1019), .Z(n29) );
  NAND U1190 ( .A(B[86]), .B(n1020), .Z(n1019) );
  NANDN U1191 ( .A(A[86]), .B(n31), .Z(n1020) );
  NANDN U1192 ( .A(n31), .B(A[86]), .Z(n1018) );
  AND U1193 ( .A(n1021), .B(n1022), .Z(n31) );
  NAND U1194 ( .A(B[85]), .B(n1023), .Z(n1022) );
  NANDN U1195 ( .A(A[85]), .B(n33), .Z(n1023) );
  NANDN U1196 ( .A(n33), .B(A[85]), .Z(n1021) );
  AND U1197 ( .A(n1024), .B(n1025), .Z(n33) );
  NAND U1198 ( .A(B[84]), .B(n1026), .Z(n1025) );
  NANDN U1199 ( .A(A[84]), .B(n35), .Z(n1026) );
  NANDN U1200 ( .A(n35), .B(A[84]), .Z(n1024) );
  AND U1201 ( .A(n1027), .B(n1028), .Z(n35) );
  NAND U1202 ( .A(B[83]), .B(n1029), .Z(n1028) );
  NANDN U1203 ( .A(A[83]), .B(n37), .Z(n1029) );
  NANDN U1204 ( .A(n37), .B(A[83]), .Z(n1027) );
  AND U1205 ( .A(n1030), .B(n1031), .Z(n37) );
  NAND U1206 ( .A(B[82]), .B(n1032), .Z(n1031) );
  NANDN U1207 ( .A(A[82]), .B(n39), .Z(n1032) );
  NANDN U1208 ( .A(n39), .B(A[82]), .Z(n1030) );
  AND U1209 ( .A(n1033), .B(n1034), .Z(n39) );
  NAND U1210 ( .A(B[81]), .B(n1035), .Z(n1034) );
  NANDN U1211 ( .A(A[81]), .B(n41), .Z(n1035) );
  NANDN U1212 ( .A(n41), .B(A[81]), .Z(n1033) );
  AND U1213 ( .A(n1036), .B(n1037), .Z(n41) );
  NAND U1214 ( .A(B[80]), .B(n1038), .Z(n1037) );
  NANDN U1215 ( .A(A[80]), .B(n43), .Z(n1038) );
  NANDN U1216 ( .A(n43), .B(A[80]), .Z(n1036) );
  AND U1217 ( .A(n1039), .B(n1040), .Z(n43) );
  NAND U1218 ( .A(B[79]), .B(n1041), .Z(n1040) );
  NANDN U1219 ( .A(A[79]), .B(n47), .Z(n1041) );
  NANDN U1220 ( .A(n47), .B(A[79]), .Z(n1039) );
  AND U1221 ( .A(n1042), .B(n1043), .Z(n47) );
  NAND U1222 ( .A(B[78]), .B(n1044), .Z(n1043) );
  NANDN U1223 ( .A(A[78]), .B(n49), .Z(n1044) );
  NANDN U1224 ( .A(n49), .B(A[78]), .Z(n1042) );
  AND U1225 ( .A(n1045), .B(n1046), .Z(n49) );
  NAND U1226 ( .A(B[77]), .B(n1047), .Z(n1046) );
  NANDN U1227 ( .A(A[77]), .B(n51), .Z(n1047) );
  NANDN U1228 ( .A(n51), .B(A[77]), .Z(n1045) );
  AND U1229 ( .A(n1048), .B(n1049), .Z(n51) );
  NAND U1230 ( .A(B[76]), .B(n1050), .Z(n1049) );
  NANDN U1231 ( .A(A[76]), .B(n53), .Z(n1050) );
  NANDN U1232 ( .A(n53), .B(A[76]), .Z(n1048) );
  AND U1233 ( .A(n1051), .B(n1052), .Z(n53) );
  NAND U1234 ( .A(B[75]), .B(n1053), .Z(n1052) );
  NANDN U1235 ( .A(A[75]), .B(n55), .Z(n1053) );
  NANDN U1236 ( .A(n55), .B(A[75]), .Z(n1051) );
  AND U1237 ( .A(n1054), .B(n1055), .Z(n55) );
  NAND U1238 ( .A(B[74]), .B(n1056), .Z(n1055) );
  NANDN U1239 ( .A(A[74]), .B(n57), .Z(n1056) );
  NANDN U1240 ( .A(n57), .B(A[74]), .Z(n1054) );
  AND U1241 ( .A(n1057), .B(n1058), .Z(n57) );
  NAND U1242 ( .A(B[73]), .B(n1059), .Z(n1058) );
  NANDN U1243 ( .A(A[73]), .B(n59), .Z(n1059) );
  NANDN U1244 ( .A(n59), .B(A[73]), .Z(n1057) );
  AND U1245 ( .A(n1060), .B(n1061), .Z(n59) );
  NAND U1246 ( .A(B[72]), .B(n1062), .Z(n1061) );
  NANDN U1247 ( .A(A[72]), .B(n61), .Z(n1062) );
  NANDN U1248 ( .A(n61), .B(A[72]), .Z(n1060) );
  AND U1249 ( .A(n1063), .B(n1064), .Z(n61) );
  NAND U1250 ( .A(B[71]), .B(n1065), .Z(n1064) );
  NANDN U1251 ( .A(A[71]), .B(n63), .Z(n1065) );
  NANDN U1252 ( .A(n63), .B(A[71]), .Z(n1063) );
  AND U1253 ( .A(n1066), .B(n1067), .Z(n63) );
  NAND U1254 ( .A(B[70]), .B(n1068), .Z(n1067) );
  NANDN U1255 ( .A(A[70]), .B(n65), .Z(n1068) );
  NANDN U1256 ( .A(n65), .B(A[70]), .Z(n1066) );
  AND U1257 ( .A(n1069), .B(n1070), .Z(n65) );
  NAND U1258 ( .A(B[69]), .B(n1071), .Z(n1070) );
  NANDN U1259 ( .A(A[69]), .B(n69), .Z(n1071) );
  NANDN U1260 ( .A(n69), .B(A[69]), .Z(n1069) );
  AND U1261 ( .A(n1072), .B(n1073), .Z(n69) );
  NAND U1262 ( .A(B[68]), .B(n1074), .Z(n1073) );
  NANDN U1263 ( .A(A[68]), .B(n71), .Z(n1074) );
  NANDN U1264 ( .A(n71), .B(A[68]), .Z(n1072) );
  AND U1265 ( .A(n1075), .B(n1076), .Z(n71) );
  NAND U1266 ( .A(B[67]), .B(n1077), .Z(n1076) );
  NANDN U1267 ( .A(A[67]), .B(n73), .Z(n1077) );
  NANDN U1268 ( .A(n73), .B(A[67]), .Z(n1075) );
  AND U1269 ( .A(n1078), .B(n1079), .Z(n73) );
  NAND U1270 ( .A(B[66]), .B(n1080), .Z(n1079) );
  NANDN U1271 ( .A(A[66]), .B(n75), .Z(n1080) );
  NANDN U1272 ( .A(n75), .B(A[66]), .Z(n1078) );
  AND U1273 ( .A(n1081), .B(n1082), .Z(n75) );
  NAND U1274 ( .A(B[65]), .B(n1083), .Z(n1082) );
  NANDN U1275 ( .A(A[65]), .B(n77), .Z(n1083) );
  NANDN U1276 ( .A(n77), .B(A[65]), .Z(n1081) );
  AND U1277 ( .A(n1084), .B(n1085), .Z(n77) );
  NAND U1278 ( .A(B[64]), .B(n1086), .Z(n1085) );
  NANDN U1279 ( .A(A[64]), .B(n79), .Z(n1086) );
  NANDN U1280 ( .A(n79), .B(A[64]), .Z(n1084) );
  AND U1281 ( .A(n1087), .B(n1088), .Z(n79) );
  NAND U1282 ( .A(B[63]), .B(n1089), .Z(n1088) );
  NANDN U1283 ( .A(A[63]), .B(n81), .Z(n1089) );
  NANDN U1284 ( .A(n81), .B(A[63]), .Z(n1087) );
  AND U1285 ( .A(n1090), .B(n1091), .Z(n81) );
  NAND U1286 ( .A(B[62]), .B(n1092), .Z(n1091) );
  NANDN U1287 ( .A(A[62]), .B(n83), .Z(n1092) );
  NANDN U1288 ( .A(n83), .B(A[62]), .Z(n1090) );
  AND U1289 ( .A(n1093), .B(n1094), .Z(n83) );
  NAND U1290 ( .A(B[61]), .B(n1095), .Z(n1094) );
  NANDN U1291 ( .A(A[61]), .B(n85), .Z(n1095) );
  NANDN U1292 ( .A(n85), .B(A[61]), .Z(n1093) );
  AND U1293 ( .A(n1096), .B(n1097), .Z(n85) );
  NAND U1294 ( .A(B[60]), .B(n1098), .Z(n1097) );
  NANDN U1295 ( .A(A[60]), .B(n87), .Z(n1098) );
  NANDN U1296 ( .A(n87), .B(A[60]), .Z(n1096) );
  AND U1297 ( .A(n1099), .B(n1100), .Z(n87) );
  NAND U1298 ( .A(B[59]), .B(n1101), .Z(n1100) );
  NANDN U1299 ( .A(A[59]), .B(n91), .Z(n1101) );
  NANDN U1300 ( .A(n91), .B(A[59]), .Z(n1099) );
  AND U1301 ( .A(n1102), .B(n1103), .Z(n91) );
  NAND U1302 ( .A(B[58]), .B(n1104), .Z(n1103) );
  NANDN U1303 ( .A(A[58]), .B(n93), .Z(n1104) );
  NANDN U1304 ( .A(n93), .B(A[58]), .Z(n1102) );
  AND U1305 ( .A(n1105), .B(n1106), .Z(n93) );
  NAND U1306 ( .A(B[57]), .B(n1107), .Z(n1106) );
  NANDN U1307 ( .A(A[57]), .B(n95), .Z(n1107) );
  NANDN U1308 ( .A(n95), .B(A[57]), .Z(n1105) );
  AND U1309 ( .A(n1108), .B(n1109), .Z(n95) );
  NAND U1310 ( .A(B[56]), .B(n1110), .Z(n1109) );
  NANDN U1311 ( .A(A[56]), .B(n97), .Z(n1110) );
  NANDN U1312 ( .A(n97), .B(A[56]), .Z(n1108) );
  AND U1313 ( .A(n1111), .B(n1112), .Z(n97) );
  NAND U1314 ( .A(B[55]), .B(n1113), .Z(n1112) );
  NANDN U1315 ( .A(A[55]), .B(n99), .Z(n1113) );
  NANDN U1316 ( .A(n99), .B(A[55]), .Z(n1111) );
  AND U1317 ( .A(n1114), .B(n1115), .Z(n99) );
  NAND U1318 ( .A(B[54]), .B(n1116), .Z(n1115) );
  NANDN U1319 ( .A(A[54]), .B(n101), .Z(n1116) );
  NANDN U1320 ( .A(n101), .B(A[54]), .Z(n1114) );
  AND U1321 ( .A(n1117), .B(n1118), .Z(n101) );
  NAND U1322 ( .A(B[53]), .B(n1119), .Z(n1118) );
  NANDN U1323 ( .A(A[53]), .B(n103), .Z(n1119) );
  NANDN U1324 ( .A(n103), .B(A[53]), .Z(n1117) );
  AND U1325 ( .A(n1120), .B(n1121), .Z(n103) );
  NAND U1326 ( .A(B[52]), .B(n1122), .Z(n1121) );
  NANDN U1327 ( .A(A[52]), .B(n105), .Z(n1122) );
  NANDN U1328 ( .A(n105), .B(A[52]), .Z(n1120) );
  AND U1329 ( .A(n1123), .B(n1124), .Z(n105) );
  NAND U1330 ( .A(B[51]), .B(n1125), .Z(n1124) );
  NANDN U1331 ( .A(A[51]), .B(n107), .Z(n1125) );
  NANDN U1332 ( .A(n107), .B(A[51]), .Z(n1123) );
  AND U1333 ( .A(n1126), .B(n1127), .Z(n107) );
  NAND U1334 ( .A(B[50]), .B(n1128), .Z(n1127) );
  NANDN U1335 ( .A(A[50]), .B(n109), .Z(n1128) );
  NANDN U1336 ( .A(n109), .B(A[50]), .Z(n1126) );
  AND U1337 ( .A(n1129), .B(n1130), .Z(n109) );
  NAND U1338 ( .A(B[49]), .B(n1131), .Z(n1130) );
  NANDN U1339 ( .A(A[49]), .B(n113), .Z(n1131) );
  NANDN U1340 ( .A(n113), .B(A[49]), .Z(n1129) );
  AND U1341 ( .A(n1132), .B(n1133), .Z(n113) );
  NAND U1342 ( .A(B[48]), .B(n1134), .Z(n1133) );
  NANDN U1343 ( .A(A[48]), .B(n115), .Z(n1134) );
  NANDN U1344 ( .A(n115), .B(A[48]), .Z(n1132) );
  AND U1345 ( .A(n1135), .B(n1136), .Z(n115) );
  NAND U1346 ( .A(B[47]), .B(n1137), .Z(n1136) );
  NANDN U1347 ( .A(A[47]), .B(n117), .Z(n1137) );
  NANDN U1348 ( .A(n117), .B(A[47]), .Z(n1135) );
  AND U1349 ( .A(n1138), .B(n1139), .Z(n117) );
  NAND U1350 ( .A(B[46]), .B(n1140), .Z(n1139) );
  NANDN U1351 ( .A(A[46]), .B(n119), .Z(n1140) );
  NANDN U1352 ( .A(n119), .B(A[46]), .Z(n1138) );
  AND U1353 ( .A(n1141), .B(n1142), .Z(n119) );
  NAND U1354 ( .A(B[45]), .B(n1143), .Z(n1142) );
  NANDN U1355 ( .A(A[45]), .B(n121), .Z(n1143) );
  NANDN U1356 ( .A(n121), .B(A[45]), .Z(n1141) );
  AND U1357 ( .A(n1144), .B(n1145), .Z(n121) );
  NAND U1358 ( .A(B[44]), .B(n1146), .Z(n1145) );
  NANDN U1359 ( .A(A[44]), .B(n123), .Z(n1146) );
  NANDN U1360 ( .A(n123), .B(A[44]), .Z(n1144) );
  AND U1361 ( .A(n1147), .B(n1148), .Z(n123) );
  NAND U1362 ( .A(B[43]), .B(n1149), .Z(n1148) );
  NANDN U1363 ( .A(A[43]), .B(n125), .Z(n1149) );
  NANDN U1364 ( .A(n125), .B(A[43]), .Z(n1147) );
  AND U1365 ( .A(n1150), .B(n1151), .Z(n125) );
  NAND U1366 ( .A(B[42]), .B(n1152), .Z(n1151) );
  NANDN U1367 ( .A(A[42]), .B(n127), .Z(n1152) );
  NANDN U1368 ( .A(n127), .B(A[42]), .Z(n1150) );
  AND U1369 ( .A(n1153), .B(n1154), .Z(n127) );
  NAND U1370 ( .A(B[41]), .B(n1155), .Z(n1154) );
  NANDN U1371 ( .A(A[41]), .B(n129), .Z(n1155) );
  NANDN U1372 ( .A(n129), .B(A[41]), .Z(n1153) );
  AND U1373 ( .A(n1156), .B(n1157), .Z(n129) );
  NAND U1374 ( .A(B[40]), .B(n1158), .Z(n1157) );
  NANDN U1375 ( .A(A[40]), .B(n131), .Z(n1158) );
  NANDN U1376 ( .A(n131), .B(A[40]), .Z(n1156) );
  AND U1377 ( .A(n1159), .B(n1160), .Z(n131) );
  NAND U1378 ( .A(B[39]), .B(n1161), .Z(n1160) );
  NANDN U1379 ( .A(A[39]), .B(n135), .Z(n1161) );
  NANDN U1380 ( .A(n135), .B(A[39]), .Z(n1159) );
  AND U1381 ( .A(n1162), .B(n1163), .Z(n135) );
  NAND U1382 ( .A(B[38]), .B(n1164), .Z(n1163) );
  NANDN U1383 ( .A(A[38]), .B(n137), .Z(n1164) );
  NANDN U1384 ( .A(n137), .B(A[38]), .Z(n1162) );
  AND U1385 ( .A(n1165), .B(n1166), .Z(n137) );
  NAND U1386 ( .A(B[37]), .B(n1167), .Z(n1166) );
  NANDN U1387 ( .A(A[37]), .B(n139), .Z(n1167) );
  NANDN U1388 ( .A(n139), .B(A[37]), .Z(n1165) );
  AND U1389 ( .A(n1168), .B(n1169), .Z(n139) );
  NAND U1390 ( .A(B[36]), .B(n1170), .Z(n1169) );
  NANDN U1391 ( .A(A[36]), .B(n141), .Z(n1170) );
  NANDN U1392 ( .A(n141), .B(A[36]), .Z(n1168) );
  AND U1393 ( .A(n1171), .B(n1172), .Z(n141) );
  NAND U1394 ( .A(B[35]), .B(n1173), .Z(n1172) );
  NANDN U1395 ( .A(A[35]), .B(n143), .Z(n1173) );
  NANDN U1396 ( .A(n143), .B(A[35]), .Z(n1171) );
  AND U1397 ( .A(n1174), .B(n1175), .Z(n143) );
  NAND U1398 ( .A(B[34]), .B(n1176), .Z(n1175) );
  NANDN U1399 ( .A(A[34]), .B(n145), .Z(n1176) );
  NANDN U1400 ( .A(n145), .B(A[34]), .Z(n1174) );
  AND U1401 ( .A(n1177), .B(n1178), .Z(n145) );
  NAND U1402 ( .A(B[33]), .B(n1179), .Z(n1178) );
  NANDN U1403 ( .A(A[33]), .B(n147), .Z(n1179) );
  NANDN U1404 ( .A(n147), .B(A[33]), .Z(n1177) );
  AND U1405 ( .A(n1180), .B(n1181), .Z(n147) );
  NAND U1406 ( .A(B[32]), .B(n1182), .Z(n1181) );
  NANDN U1407 ( .A(A[32]), .B(n149), .Z(n1182) );
  NANDN U1408 ( .A(n149), .B(A[32]), .Z(n1180) );
  AND U1409 ( .A(n1183), .B(n1184), .Z(n149) );
  NAND U1410 ( .A(B[31]), .B(n1185), .Z(n1184) );
  NANDN U1411 ( .A(A[31]), .B(n151), .Z(n1185) );
  NANDN U1412 ( .A(n151), .B(A[31]), .Z(n1183) );
  AND U1413 ( .A(n1186), .B(n1187), .Z(n151) );
  NAND U1414 ( .A(B[30]), .B(n1188), .Z(n1187) );
  NANDN U1415 ( .A(A[30]), .B(n153), .Z(n1188) );
  NANDN U1416 ( .A(n153), .B(A[30]), .Z(n1186) );
  AND U1417 ( .A(n1189), .B(n1190), .Z(n153) );
  NAND U1418 ( .A(B[29]), .B(n1191), .Z(n1190) );
  NANDN U1419 ( .A(A[29]), .B(n157), .Z(n1191) );
  NANDN U1420 ( .A(n157), .B(A[29]), .Z(n1189) );
  AND U1421 ( .A(n1192), .B(n1193), .Z(n157) );
  NAND U1422 ( .A(B[28]), .B(n1194), .Z(n1193) );
  NANDN U1423 ( .A(A[28]), .B(n159), .Z(n1194) );
  NANDN U1424 ( .A(n159), .B(A[28]), .Z(n1192) );
  AND U1425 ( .A(n1195), .B(n1196), .Z(n159) );
  NAND U1426 ( .A(B[27]), .B(n1197), .Z(n1196) );
  NANDN U1427 ( .A(A[27]), .B(n161), .Z(n1197) );
  NANDN U1428 ( .A(n161), .B(A[27]), .Z(n1195) );
  AND U1429 ( .A(n1198), .B(n1199), .Z(n161) );
  NAND U1430 ( .A(B[26]), .B(n1200), .Z(n1199) );
  NANDN U1431 ( .A(A[26]), .B(n163), .Z(n1200) );
  NANDN U1432 ( .A(n163), .B(A[26]), .Z(n1198) );
  AND U1433 ( .A(n1201), .B(n1202), .Z(n163) );
  NAND U1434 ( .A(B[25]), .B(n1203), .Z(n1202) );
  NANDN U1435 ( .A(A[25]), .B(n165), .Z(n1203) );
  NANDN U1436 ( .A(n165), .B(A[25]), .Z(n1201) );
  AND U1437 ( .A(n1204), .B(n1205), .Z(n165) );
  NAND U1438 ( .A(B[24]), .B(n1206), .Z(n1205) );
  NANDN U1439 ( .A(A[24]), .B(n203), .Z(n1206) );
  NANDN U1440 ( .A(n203), .B(A[24]), .Z(n1204) );
  AND U1441 ( .A(n1207), .B(n1208), .Z(n203) );
  NAND U1442 ( .A(B[23]), .B(n1209), .Z(n1208) );
  NANDN U1443 ( .A(A[23]), .B(n255), .Z(n1209) );
  NANDN U1444 ( .A(n255), .B(A[23]), .Z(n1207) );
  AND U1445 ( .A(n1210), .B(n1211), .Z(n255) );
  NAND U1446 ( .A(B[22]), .B(n1212), .Z(n1211) );
  NANDN U1447 ( .A(A[22]), .B(n307), .Z(n1212) );
  NANDN U1448 ( .A(n307), .B(A[22]), .Z(n1210) );
  AND U1449 ( .A(n1213), .B(n1214), .Z(n307) );
  NAND U1450 ( .A(B[21]), .B(n1215), .Z(n1214) );
  NANDN U1451 ( .A(A[21]), .B(n359), .Z(n1215) );
  NANDN U1452 ( .A(n359), .B(A[21]), .Z(n1213) );
  AND U1453 ( .A(n1216), .B(n1217), .Z(n359) );
  NAND U1454 ( .A(B[20]), .B(n1218), .Z(n1217) );
  NANDN U1455 ( .A(A[20]), .B(n411), .Z(n1218) );
  NANDN U1456 ( .A(n411), .B(A[20]), .Z(n1216) );
  AND U1457 ( .A(n1219), .B(n1220), .Z(n411) );
  NAND U1458 ( .A(B[19]), .B(n1221), .Z(n1220) );
  NANDN U1459 ( .A(A[19]), .B(n463), .Z(n1221) );
  NANDN U1460 ( .A(n463), .B(A[19]), .Z(n1219) );
  AND U1461 ( .A(n1222), .B(n1223), .Z(n463) );
  NAND U1462 ( .A(B[18]), .B(n1224), .Z(n1223) );
  NANDN U1463 ( .A(A[18]), .B(n515), .Z(n1224) );
  NANDN U1464 ( .A(n515), .B(A[18]), .Z(n1222) );
  AND U1465 ( .A(n1225), .B(n1226), .Z(n515) );
  NAND U1466 ( .A(B[17]), .B(n1227), .Z(n1226) );
  NANDN U1467 ( .A(A[17]), .B(n567), .Z(n1227) );
  NANDN U1468 ( .A(n567), .B(A[17]), .Z(n1225) );
  AND U1469 ( .A(n1228), .B(n1229), .Z(n567) );
  NAND U1470 ( .A(B[16]), .B(n1230), .Z(n1229) );
  NANDN U1471 ( .A(A[16]), .B(n619), .Z(n1230) );
  NANDN U1472 ( .A(n619), .B(A[16]), .Z(n1228) );
  AND U1473 ( .A(n1231), .B(n1232), .Z(n619) );
  NAND U1474 ( .A(B[15]), .B(n1233), .Z(n1232) );
  NANDN U1475 ( .A(A[15]), .B(n671), .Z(n1233) );
  NANDN U1476 ( .A(n671), .B(A[15]), .Z(n1231) );
  AND U1477 ( .A(n1234), .B(n1235), .Z(n671) );
  NAND U1478 ( .A(B[14]), .B(n1236), .Z(n1235) );
  NANDN U1479 ( .A(A[14]), .B(n723), .Z(n1236) );
  NANDN U1480 ( .A(n723), .B(A[14]), .Z(n1234) );
  AND U1481 ( .A(n1237), .B(n1238), .Z(n723) );
  NAND U1482 ( .A(B[13]), .B(n1239), .Z(n1238) );
  NANDN U1483 ( .A(A[13]), .B(n775), .Z(n1239) );
  NANDN U1484 ( .A(n775), .B(A[13]), .Z(n1237) );
  AND U1485 ( .A(n1240), .B(n1241), .Z(n775) );
  NAND U1486 ( .A(B[12]), .B(n1242), .Z(n1241) );
  NANDN U1487 ( .A(A[12]), .B(n827), .Z(n1242) );
  NANDN U1488 ( .A(n827), .B(A[12]), .Z(n1240) );
  AND U1489 ( .A(n1243), .B(n1244), .Z(n827) );
  NAND U1490 ( .A(B[11]), .B(n1245), .Z(n1244) );
  NANDN U1491 ( .A(A[11]), .B(n879), .Z(n1245) );
  NANDN U1492 ( .A(n879), .B(A[11]), .Z(n1243) );
  AND U1493 ( .A(n1246), .B(n1247), .Z(n879) );
  NAND U1494 ( .A(B[10]), .B(n1248), .Z(n1247) );
  NANDN U1495 ( .A(A[10]), .B(n931), .Z(n1248) );
  NANDN U1496 ( .A(n931), .B(A[10]), .Z(n1246) );
  AND U1497 ( .A(n1249), .B(n1250), .Z(n931) );
  NAND U1498 ( .A(B[9]), .B(n1251), .Z(n1250) );
  OR U1499 ( .A(n1), .B(A[9]), .Z(n1251) );
  NAND U1500 ( .A(A[9]), .B(n1), .Z(n1249) );
  NAND U1501 ( .A(n1252), .B(n1253), .Z(n1) );
  NAND U1502 ( .A(B[8]), .B(n1254), .Z(n1253) );
  NANDN U1503 ( .A(A[8]), .B(n23), .Z(n1254) );
  NANDN U1504 ( .A(n23), .B(A[8]), .Z(n1252) );
  AND U1505 ( .A(n1255), .B(n1256), .Z(n23) );
  NAND U1506 ( .A(B[7]), .B(n1257), .Z(n1256) );
  NANDN U1507 ( .A(A[7]), .B(n45), .Z(n1257) );
  NANDN U1508 ( .A(n45), .B(A[7]), .Z(n1255) );
  AND U1509 ( .A(n1258), .B(n1259), .Z(n45) );
  NAND U1510 ( .A(B[6]), .B(n1260), .Z(n1259) );
  NANDN U1511 ( .A(A[6]), .B(n67), .Z(n1260) );
  NANDN U1512 ( .A(n67), .B(A[6]), .Z(n1258) );
  AND U1513 ( .A(n1261), .B(n1262), .Z(n67) );
  NAND U1514 ( .A(B[5]), .B(n1263), .Z(n1262) );
  NANDN U1515 ( .A(A[5]), .B(n89), .Z(n1263) );
  NANDN U1516 ( .A(n89), .B(A[5]), .Z(n1261) );
  AND U1517 ( .A(n1264), .B(n1265), .Z(n89) );
  NAND U1518 ( .A(B[4]), .B(n1266), .Z(n1265) );
  NANDN U1519 ( .A(A[4]), .B(n111), .Z(n1266) );
  NANDN U1520 ( .A(n111), .B(A[4]), .Z(n1264) );
  AND U1521 ( .A(n1267), .B(n1268), .Z(n111) );
  NAND U1522 ( .A(B[3]), .B(n1269), .Z(n1268) );
  NANDN U1523 ( .A(A[3]), .B(n133), .Z(n1269) );
  NANDN U1524 ( .A(n133), .B(A[3]), .Z(n1267) );
  AND U1525 ( .A(n1270), .B(n1271), .Z(n133) );
  NAND U1526 ( .A(B[2]), .B(n1272), .Z(n1271) );
  OR U1527 ( .A(n155), .B(A[2]), .Z(n1272) );
  NAND U1528 ( .A(A[2]), .B(n155), .Z(n1270) );
  AND U1529 ( .A(B[1]), .B(A[1]), .Z(n155) );
endmodule


module modmult_step_N256_4 ( xregN_1, y, n, zin, zout );
  input [255:0] y;
  input [255:0] n;
  input [257:0] zin;
  output [257:0] zout;
  input xregN_1;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123,
         N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200,
         N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211,
         N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222,
         N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233,
         N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244,
         N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255,
         N256, N257, N258, N259, N260, N261, N262, N264, N265, N266, N267,
         N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278,
         N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289,
         N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300,
         N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311,
         N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322,
         N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333,
         N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344,
         N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366,
         N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377,
         N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410,
         N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421,
         N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432,
         N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443,
         N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454,
         N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465,
         N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476,
         N477, N478, N479, N480, N481, N482, N483, N484, N485, N486, N487,
         N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, N498,
         N499, N500, N501, N502, N503, N504, N505, N506, N507, N508, N509,
         N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, N520,
         N521, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771,
         N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760,
         N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749,
         N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738,
         N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727,
         N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716,
         N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705,
         N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694,
         N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683,
         N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672,
         N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661,
         N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650,
         N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639,
         N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628,
         N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617,
         N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606,
         N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595,
         N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584,
         N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573,
         N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562,
         N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551,
         N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540,
         N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529,
         N528, N527, N526, N525, N522, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039;
  wire   [257:0] z2;
  wire   [257:0] z3;
  wire   SYNOPSYS_UNCONNECTED__0;

  modmult_step_N256_4_DW01_sub_0 sub_129_aco ( .A(z3), .B({1'b0, 1'b0, N780, 
        N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, 
        N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, 
        N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, 
        N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, 
        N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, 
        N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, 
        N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, 
        N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, 
        N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, 
        N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, 
        N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, 
        N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, 
        N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, 
        N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, 
        N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, 
        N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, 
        N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, 
        N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, 
        N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, 
        N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, 
        N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, 
        N527, N526, N525}), .CI(1'b0), .DIFF(zout) );
  modmult_step_N256_4_DW02_mult_0 mult_sub_129_aco ( .A(n), .B(N522), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__0, N780, N779, N778, N777, N776, N775, N774, 
        N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, 
        N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, 
        N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, 
        N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, 
        N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, 
        N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, 
        N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, 
        N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, 
        N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, 
        N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, 
        N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, 
        N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, 
        N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, 
        N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, 
        N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, 
        N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, 
        N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, 
        N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, 
        N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, 
        N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, 
        N533, N532, N531, N530, N529, N528, N527, N526, N525}) );
  modmult_step_N256_4_DW01_cmp2_0 gte_128 ( .A({1'b0, 1'b0, n}), .B(z3), .LEQ(
        1'b1), .TC(1'b0), .LT_LE(N522) );
  modmult_step_N256_4_DW01_sub_1 sub_124 ( .A(z2), .B({1'b0, 1'b0, n}), .CI(
        1'b0), .DIFF({N521, N520, N519, N518, N517, N516, N515, N514, N513, 
        N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, 
        N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, 
        N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, 
        N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, 
        N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, 
        N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, 
        N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, 
        N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, 
        N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, 
        N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, 
        N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, 
        N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, 
        N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, 
        N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, 
        N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, 
        N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, 
        N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, 
        N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, 
        N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, 
        N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, 
        N272, N271, N270, N269, N268, N267, N266, N265, N264}) );
  modmult_step_N256_4_DW01_cmp2_1 gt_123 ( .A({1'b0, 1'b0, n}), .B(z2), .LEQ(
        1'b0), .TC(1'b0), .LT_LE(N262) );
  modmult_step_N256_4_DW01_add_0 add_119 ( .A({zin[256:0], 1'b0}), .B({1'b0, 
        1'b0, y}), .CI(1'b0), .SUM({N261, N260, N259, N258, N257, N256, N255, 
        N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, 
        N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, 
        N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, 
        N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, 
        N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, 
        N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, 
        N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, 
        N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, 
        N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, 
        N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, 
        N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, 
        N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, 
        N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, 
        N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, 
        N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4}) );
  NAND U5 ( .A(n1), .B(n2), .Z(z3[9]) );
  NANDN U6 ( .A(N262), .B(z2[9]), .Z(n2) );
  NANDN U7 ( .A(n3), .B(N273), .Z(n1) );
  NAND U8 ( .A(n4), .B(n5), .Z(z3[99]) );
  NANDN U9 ( .A(N262), .B(z2[99]), .Z(n5) );
  NANDN U10 ( .A(n3), .B(N363), .Z(n4) );
  NAND U11 ( .A(n6), .B(n7), .Z(z3[98]) );
  NANDN U17 ( .A(N262), .B(z2[98]), .Z(n7) );
  NANDN U18 ( .A(n3), .B(N362), .Z(n6) );
  NAND U19 ( .A(n8), .B(n9), .Z(z3[97]) );
  NANDN U20 ( .A(N262), .B(z2[97]), .Z(n9) );
  NANDN U21 ( .A(n3), .B(N361), .Z(n8) );
  NAND U22 ( .A(n10), .B(n11), .Z(z3[96]) );
  NANDN U23 ( .A(N262), .B(z2[96]), .Z(n11) );
  NANDN U24 ( .A(n3), .B(N360), .Z(n10) );
  NAND U25 ( .A(n12), .B(n13), .Z(z3[95]) );
  NANDN U26 ( .A(N262), .B(z2[95]), .Z(n13) );
  NANDN U27 ( .A(n3), .B(N359), .Z(n12) );
  NAND U28 ( .A(n14), .B(n23), .Z(z3[94]) );
  NANDN U29 ( .A(N262), .B(z2[94]), .Z(n23) );
  NANDN U30 ( .A(n3), .B(N358), .Z(n14) );
  NAND U31 ( .A(n24), .B(n25), .Z(z3[93]) );
  NANDN U32 ( .A(N262), .B(z2[93]), .Z(n25) );
  NANDN U33 ( .A(n3), .B(N357), .Z(n24) );
  NAND U34 ( .A(n26), .B(n27), .Z(z3[92]) );
  NANDN U35 ( .A(N262), .B(z2[92]), .Z(n27) );
  NANDN U36 ( .A(n3), .B(N356), .Z(n26) );
  NAND U37 ( .A(n28), .B(n29), .Z(z3[91]) );
  NANDN U38 ( .A(N262), .B(z2[91]), .Z(n29) );
  NANDN U39 ( .A(n3), .B(N355), .Z(n28) );
  NAND U40 ( .A(n30), .B(n31), .Z(z3[90]) );
  NANDN U41 ( .A(N262), .B(z2[90]), .Z(n31) );
  NANDN U42 ( .A(n3), .B(N354), .Z(n30) );
  NAND U43 ( .A(n32), .B(n33), .Z(z3[8]) );
  NANDN U44 ( .A(N262), .B(z2[8]), .Z(n33) );
  NANDN U45 ( .A(n3), .B(N272), .Z(n32) );
  NAND U46 ( .A(n34), .B(n35), .Z(z3[89]) );
  NANDN U47 ( .A(N262), .B(z2[89]), .Z(n35) );
  NANDN U48 ( .A(n3), .B(N353), .Z(n34) );
  NAND U49 ( .A(n36), .B(n37), .Z(z3[88]) );
  NANDN U50 ( .A(N262), .B(z2[88]), .Z(n37) );
  NANDN U51 ( .A(n3), .B(N352), .Z(n36) );
  NAND U52 ( .A(n38), .B(n39), .Z(z3[87]) );
  NANDN U53 ( .A(N262), .B(z2[87]), .Z(n39) );
  NANDN U54 ( .A(n3), .B(N351), .Z(n38) );
  NAND U55 ( .A(n40), .B(n41), .Z(z3[86]) );
  NANDN U56 ( .A(N262), .B(z2[86]), .Z(n41) );
  NANDN U57 ( .A(n3), .B(N350), .Z(n40) );
  NAND U58 ( .A(n42), .B(n43), .Z(z3[85]) );
  NANDN U59 ( .A(N262), .B(z2[85]), .Z(n43) );
  NANDN U60 ( .A(n3), .B(N349), .Z(n42) );
  NAND U61 ( .A(n44), .B(n45), .Z(z3[84]) );
  NANDN U62 ( .A(N262), .B(z2[84]), .Z(n45) );
  NANDN U63 ( .A(n3), .B(N348), .Z(n44) );
  NAND U64 ( .A(n46), .B(n47), .Z(z3[83]) );
  NANDN U65 ( .A(N262), .B(z2[83]), .Z(n47) );
  NANDN U66 ( .A(n3), .B(N347), .Z(n46) );
  NAND U67 ( .A(n48), .B(n49), .Z(z3[82]) );
  NANDN U68 ( .A(N262), .B(z2[82]), .Z(n49) );
  NANDN U69 ( .A(n3), .B(N346), .Z(n48) );
  NAND U70 ( .A(n50), .B(n51), .Z(z3[81]) );
  NANDN U71 ( .A(N262), .B(z2[81]), .Z(n51) );
  NANDN U72 ( .A(n3), .B(N345), .Z(n50) );
  NAND U73 ( .A(n52), .B(n53), .Z(z3[80]) );
  NANDN U74 ( .A(N262), .B(z2[80]), .Z(n53) );
  NANDN U75 ( .A(n3), .B(N344), .Z(n52) );
  NAND U76 ( .A(n54), .B(n55), .Z(z3[7]) );
  NANDN U77 ( .A(N262), .B(z2[7]), .Z(n55) );
  NANDN U78 ( .A(n3), .B(N271), .Z(n54) );
  NAND U79 ( .A(n56), .B(n57), .Z(z3[79]) );
  NANDN U80 ( .A(N262), .B(z2[79]), .Z(n57) );
  NANDN U81 ( .A(n3), .B(N343), .Z(n56) );
  NAND U82 ( .A(n58), .B(n59), .Z(z3[78]) );
  NANDN U83 ( .A(N262), .B(z2[78]), .Z(n59) );
  NANDN U84 ( .A(n3), .B(N342), .Z(n58) );
  NAND U85 ( .A(n60), .B(n61), .Z(z3[77]) );
  NANDN U86 ( .A(N262), .B(z2[77]), .Z(n61) );
  NANDN U87 ( .A(n3), .B(N341), .Z(n60) );
  NAND U88 ( .A(n62), .B(n63), .Z(z3[76]) );
  NANDN U89 ( .A(N262), .B(z2[76]), .Z(n63) );
  NANDN U90 ( .A(n3), .B(N340), .Z(n62) );
  NAND U91 ( .A(n64), .B(n65), .Z(z3[75]) );
  NANDN U92 ( .A(N262), .B(z2[75]), .Z(n65) );
  NANDN U93 ( .A(n3), .B(N339), .Z(n64) );
  NAND U94 ( .A(n66), .B(n67), .Z(z3[74]) );
  NANDN U95 ( .A(N262), .B(z2[74]), .Z(n67) );
  NANDN U96 ( .A(n3), .B(N338), .Z(n66) );
  NAND U97 ( .A(n68), .B(n69), .Z(z3[73]) );
  NANDN U98 ( .A(N262), .B(z2[73]), .Z(n69) );
  NANDN U99 ( .A(n3), .B(N337), .Z(n68) );
  NAND U100 ( .A(n70), .B(n71), .Z(z3[72]) );
  NANDN U101 ( .A(N262), .B(z2[72]), .Z(n71) );
  NANDN U102 ( .A(n3), .B(N336), .Z(n70) );
  NAND U103 ( .A(n72), .B(n73), .Z(z3[71]) );
  NANDN U104 ( .A(N262), .B(z2[71]), .Z(n73) );
  NANDN U105 ( .A(n3), .B(N335), .Z(n72) );
  NAND U106 ( .A(n74), .B(n75), .Z(z3[70]) );
  NANDN U107 ( .A(N262), .B(z2[70]), .Z(n75) );
  NANDN U108 ( .A(n3), .B(N334), .Z(n74) );
  NAND U109 ( .A(n76), .B(n77), .Z(z3[6]) );
  NANDN U110 ( .A(N262), .B(z2[6]), .Z(n77) );
  NANDN U111 ( .A(n3), .B(N270), .Z(n76) );
  NAND U112 ( .A(n78), .B(n79), .Z(z3[69]) );
  NANDN U113 ( .A(N262), .B(z2[69]), .Z(n79) );
  NANDN U114 ( .A(n3), .B(N333), .Z(n78) );
  NAND U115 ( .A(n80), .B(n81), .Z(z3[68]) );
  NANDN U116 ( .A(N262), .B(z2[68]), .Z(n81) );
  NANDN U117 ( .A(n3), .B(N332), .Z(n80) );
  NAND U118 ( .A(n82), .B(n83), .Z(z3[67]) );
  NANDN U119 ( .A(N262), .B(z2[67]), .Z(n83) );
  NANDN U120 ( .A(n3), .B(N331), .Z(n82) );
  NAND U121 ( .A(n84), .B(n85), .Z(z3[66]) );
  NANDN U122 ( .A(N262), .B(z2[66]), .Z(n85) );
  NANDN U123 ( .A(n3), .B(N330), .Z(n84) );
  NAND U124 ( .A(n86), .B(n87), .Z(z3[65]) );
  NANDN U125 ( .A(N262), .B(z2[65]), .Z(n87) );
  NANDN U126 ( .A(n3), .B(N329), .Z(n86) );
  NAND U127 ( .A(n88), .B(n89), .Z(z3[64]) );
  NANDN U128 ( .A(N262), .B(z2[64]), .Z(n89) );
  NANDN U129 ( .A(n3), .B(N328), .Z(n88) );
  NAND U130 ( .A(n90), .B(n91), .Z(z3[63]) );
  NANDN U131 ( .A(N262), .B(z2[63]), .Z(n91) );
  NANDN U132 ( .A(n3), .B(N327), .Z(n90) );
  NAND U133 ( .A(n92), .B(n93), .Z(z3[62]) );
  NANDN U134 ( .A(N262), .B(z2[62]), .Z(n93) );
  NANDN U135 ( .A(n3), .B(N326), .Z(n92) );
  NAND U136 ( .A(n94), .B(n95), .Z(z3[61]) );
  NANDN U137 ( .A(N262), .B(z2[61]), .Z(n95) );
  NANDN U138 ( .A(n3), .B(N325), .Z(n94) );
  NAND U139 ( .A(n96), .B(n97), .Z(z3[60]) );
  NANDN U140 ( .A(N262), .B(z2[60]), .Z(n97) );
  NANDN U141 ( .A(n3), .B(N324), .Z(n96) );
  NAND U142 ( .A(n98), .B(n99), .Z(z3[5]) );
  NANDN U143 ( .A(N262), .B(z2[5]), .Z(n99) );
  NANDN U144 ( .A(n3), .B(N269), .Z(n98) );
  NAND U145 ( .A(n100), .B(n101), .Z(z3[59]) );
  NANDN U146 ( .A(N262), .B(z2[59]), .Z(n101) );
  NANDN U147 ( .A(n3), .B(N323), .Z(n100) );
  NAND U148 ( .A(n102), .B(n103), .Z(z3[58]) );
  NANDN U149 ( .A(N262), .B(z2[58]), .Z(n103) );
  NANDN U150 ( .A(n3), .B(N322), .Z(n102) );
  NAND U151 ( .A(n104), .B(n105), .Z(z3[57]) );
  NANDN U152 ( .A(N262), .B(z2[57]), .Z(n105) );
  NANDN U153 ( .A(n3), .B(N321), .Z(n104) );
  NAND U154 ( .A(n106), .B(n107), .Z(z3[56]) );
  NANDN U155 ( .A(N262), .B(z2[56]), .Z(n107) );
  NANDN U156 ( .A(n3), .B(N320), .Z(n106) );
  NAND U157 ( .A(n108), .B(n109), .Z(z3[55]) );
  NANDN U158 ( .A(N262), .B(z2[55]), .Z(n109) );
  NANDN U159 ( .A(n3), .B(N319), .Z(n108) );
  NAND U160 ( .A(n110), .B(n111), .Z(z3[54]) );
  NANDN U161 ( .A(N262), .B(z2[54]), .Z(n111) );
  NANDN U162 ( .A(n3), .B(N318), .Z(n110) );
  NAND U163 ( .A(n112), .B(n113), .Z(z3[53]) );
  NANDN U164 ( .A(N262), .B(z2[53]), .Z(n113) );
  NANDN U165 ( .A(n3), .B(N317), .Z(n112) );
  NAND U166 ( .A(n114), .B(n115), .Z(z3[52]) );
  NANDN U167 ( .A(N262), .B(z2[52]), .Z(n115) );
  NANDN U168 ( .A(n3), .B(N316), .Z(n114) );
  NAND U169 ( .A(n116), .B(n117), .Z(z3[51]) );
  NANDN U170 ( .A(N262), .B(z2[51]), .Z(n117) );
  NANDN U171 ( .A(n3), .B(N315), .Z(n116) );
  NAND U172 ( .A(n118), .B(n119), .Z(z3[50]) );
  NANDN U173 ( .A(N262), .B(z2[50]), .Z(n119) );
  NANDN U174 ( .A(n3), .B(N314), .Z(n118) );
  NAND U175 ( .A(n120), .B(n121), .Z(z3[4]) );
  NANDN U176 ( .A(N262), .B(z2[4]), .Z(n121) );
  NANDN U177 ( .A(n3), .B(N268), .Z(n120) );
  NAND U178 ( .A(n122), .B(n123), .Z(z3[49]) );
  NANDN U179 ( .A(N262), .B(z2[49]), .Z(n123) );
  NANDN U180 ( .A(n3), .B(N313), .Z(n122) );
  NAND U181 ( .A(n124), .B(n125), .Z(z3[48]) );
  NANDN U182 ( .A(N262), .B(z2[48]), .Z(n125) );
  NANDN U183 ( .A(n3), .B(N312), .Z(n124) );
  NAND U184 ( .A(n126), .B(n127), .Z(z3[47]) );
  NANDN U185 ( .A(N262), .B(z2[47]), .Z(n127) );
  NANDN U186 ( .A(n3), .B(N311), .Z(n126) );
  NAND U187 ( .A(n128), .B(n129), .Z(z3[46]) );
  NANDN U188 ( .A(N262), .B(z2[46]), .Z(n129) );
  NANDN U189 ( .A(n3), .B(N310), .Z(n128) );
  NAND U190 ( .A(n130), .B(n131), .Z(z3[45]) );
  NANDN U191 ( .A(N262), .B(z2[45]), .Z(n131) );
  NANDN U192 ( .A(n3), .B(N309), .Z(n130) );
  NAND U193 ( .A(n132), .B(n133), .Z(z3[44]) );
  NANDN U194 ( .A(N262), .B(z2[44]), .Z(n133) );
  NANDN U195 ( .A(n3), .B(N308), .Z(n132) );
  NAND U196 ( .A(n134), .B(n135), .Z(z3[43]) );
  NANDN U197 ( .A(N262), .B(z2[43]), .Z(n135) );
  NANDN U198 ( .A(n3), .B(N307), .Z(n134) );
  NAND U199 ( .A(n136), .B(n137), .Z(z3[42]) );
  NANDN U200 ( .A(N262), .B(z2[42]), .Z(n137) );
  NANDN U201 ( .A(n3), .B(N306), .Z(n136) );
  NAND U202 ( .A(n138), .B(n139), .Z(z3[41]) );
  NANDN U203 ( .A(N262), .B(z2[41]), .Z(n139) );
  NANDN U204 ( .A(n3), .B(N305), .Z(n138) );
  NAND U205 ( .A(n140), .B(n141), .Z(z3[40]) );
  NANDN U206 ( .A(N262), .B(z2[40]), .Z(n141) );
  NANDN U207 ( .A(n3), .B(N304), .Z(n140) );
  NAND U208 ( .A(n142), .B(n143), .Z(z3[3]) );
  NANDN U209 ( .A(N262), .B(z2[3]), .Z(n143) );
  NANDN U210 ( .A(n3), .B(N267), .Z(n142) );
  NAND U211 ( .A(n144), .B(n145), .Z(z3[39]) );
  NANDN U212 ( .A(N262), .B(z2[39]), .Z(n145) );
  NANDN U213 ( .A(n3), .B(N303), .Z(n144) );
  NAND U214 ( .A(n146), .B(n147), .Z(z3[38]) );
  NANDN U215 ( .A(N262), .B(z2[38]), .Z(n147) );
  NANDN U216 ( .A(n3), .B(N302), .Z(n146) );
  NAND U217 ( .A(n148), .B(n149), .Z(z3[37]) );
  NANDN U218 ( .A(N262), .B(z2[37]), .Z(n149) );
  NANDN U219 ( .A(n3), .B(N301), .Z(n148) );
  NAND U220 ( .A(n150), .B(n151), .Z(z3[36]) );
  NANDN U221 ( .A(N262), .B(z2[36]), .Z(n151) );
  NANDN U222 ( .A(n3), .B(N300), .Z(n150) );
  NAND U223 ( .A(n152), .B(n153), .Z(z3[35]) );
  NANDN U224 ( .A(N262), .B(z2[35]), .Z(n153) );
  NANDN U225 ( .A(n3), .B(N299), .Z(n152) );
  NAND U226 ( .A(n154), .B(n155), .Z(z3[34]) );
  NANDN U227 ( .A(N262), .B(z2[34]), .Z(n155) );
  NANDN U228 ( .A(n3), .B(N298), .Z(n154) );
  NAND U229 ( .A(n156), .B(n157), .Z(z3[33]) );
  NANDN U230 ( .A(N262), .B(z2[33]), .Z(n157) );
  NANDN U231 ( .A(n3), .B(N297), .Z(n156) );
  NAND U232 ( .A(n158), .B(n159), .Z(z3[32]) );
  NANDN U233 ( .A(N262), .B(z2[32]), .Z(n159) );
  NANDN U234 ( .A(n3), .B(N296), .Z(n158) );
  NAND U235 ( .A(n160), .B(n161), .Z(z3[31]) );
  NANDN U236 ( .A(N262), .B(z2[31]), .Z(n161) );
  NANDN U237 ( .A(n3), .B(N295), .Z(n160) );
  NAND U238 ( .A(n162), .B(n163), .Z(z3[30]) );
  NANDN U239 ( .A(N262), .B(z2[30]), .Z(n163) );
  NANDN U240 ( .A(n3), .B(N294), .Z(n162) );
  NAND U241 ( .A(n164), .B(n165), .Z(z3[2]) );
  NANDN U242 ( .A(N262), .B(z2[2]), .Z(n165) );
  NANDN U243 ( .A(n3), .B(N266), .Z(n164) );
  NAND U244 ( .A(n166), .B(n167), .Z(z3[29]) );
  NANDN U245 ( .A(N262), .B(z2[29]), .Z(n167) );
  NANDN U246 ( .A(n3), .B(N293), .Z(n166) );
  NAND U247 ( .A(n168), .B(n169), .Z(z3[28]) );
  NANDN U248 ( .A(N262), .B(z2[28]), .Z(n169) );
  NANDN U249 ( .A(n3), .B(N292), .Z(n168) );
  NAND U250 ( .A(n170), .B(n171), .Z(z3[27]) );
  NANDN U251 ( .A(N262), .B(z2[27]), .Z(n171) );
  NANDN U252 ( .A(n3), .B(N291), .Z(n170) );
  NAND U253 ( .A(n172), .B(n173), .Z(z3[26]) );
  NANDN U254 ( .A(N262), .B(z2[26]), .Z(n173) );
  NANDN U255 ( .A(n3), .B(N290), .Z(n172) );
  NAND U256 ( .A(n174), .B(n175), .Z(z3[25]) );
  NANDN U257 ( .A(N262), .B(z2[25]), .Z(n175) );
  NANDN U258 ( .A(n3), .B(N289), .Z(n174) );
  NAND U259 ( .A(n176), .B(n177), .Z(z3[257]) );
  NANDN U260 ( .A(N262), .B(z2[257]), .Z(n177) );
  NANDN U261 ( .A(n3), .B(N521), .Z(n176) );
  NAND U262 ( .A(n178), .B(n179), .Z(z3[256]) );
  NANDN U263 ( .A(N262), .B(z2[256]), .Z(n179) );
  NANDN U264 ( .A(n3), .B(N520), .Z(n178) );
  NAND U265 ( .A(n180), .B(n181), .Z(z3[255]) );
  NANDN U266 ( .A(N262), .B(z2[255]), .Z(n181) );
  NANDN U267 ( .A(n3), .B(N519), .Z(n180) );
  NAND U268 ( .A(n182), .B(n183), .Z(z3[254]) );
  NANDN U269 ( .A(N262), .B(z2[254]), .Z(n183) );
  NANDN U270 ( .A(n3), .B(N518), .Z(n182) );
  NAND U271 ( .A(n184), .B(n185), .Z(z3[253]) );
  NANDN U272 ( .A(N262), .B(z2[253]), .Z(n185) );
  NANDN U273 ( .A(n3), .B(N517), .Z(n184) );
  NAND U274 ( .A(n186), .B(n187), .Z(z3[252]) );
  NANDN U275 ( .A(N262), .B(z2[252]), .Z(n187) );
  NANDN U276 ( .A(n3), .B(N516), .Z(n186) );
  NAND U277 ( .A(n188), .B(n189), .Z(z3[251]) );
  NANDN U278 ( .A(N262), .B(z2[251]), .Z(n189) );
  NANDN U279 ( .A(n3), .B(N515), .Z(n188) );
  NAND U280 ( .A(n190), .B(n191), .Z(z3[250]) );
  NANDN U281 ( .A(N262), .B(z2[250]), .Z(n191) );
  NANDN U282 ( .A(n3), .B(N514), .Z(n190) );
  NAND U283 ( .A(n192), .B(n193), .Z(z3[24]) );
  NANDN U284 ( .A(N262), .B(z2[24]), .Z(n193) );
  NANDN U285 ( .A(n3), .B(N288), .Z(n192) );
  NAND U286 ( .A(n194), .B(n195), .Z(z3[249]) );
  NANDN U287 ( .A(N262), .B(z2[249]), .Z(n195) );
  NANDN U288 ( .A(n3), .B(N513), .Z(n194) );
  NAND U289 ( .A(n196), .B(n197), .Z(z3[248]) );
  NANDN U290 ( .A(N262), .B(z2[248]), .Z(n197) );
  NANDN U291 ( .A(n3), .B(N512), .Z(n196) );
  NAND U292 ( .A(n198), .B(n199), .Z(z3[247]) );
  NANDN U293 ( .A(N262), .B(z2[247]), .Z(n199) );
  NANDN U294 ( .A(n3), .B(N511), .Z(n198) );
  NAND U295 ( .A(n200), .B(n201), .Z(z3[246]) );
  NANDN U296 ( .A(N262), .B(z2[246]), .Z(n201) );
  NANDN U297 ( .A(n3), .B(N510), .Z(n200) );
  NAND U298 ( .A(n202), .B(n203), .Z(z3[245]) );
  NANDN U299 ( .A(N262), .B(z2[245]), .Z(n203) );
  NANDN U300 ( .A(n3), .B(N509), .Z(n202) );
  NAND U301 ( .A(n204), .B(n205), .Z(z3[244]) );
  NANDN U302 ( .A(N262), .B(z2[244]), .Z(n205) );
  NANDN U303 ( .A(n3), .B(N508), .Z(n204) );
  NAND U304 ( .A(n206), .B(n207), .Z(z3[243]) );
  NANDN U305 ( .A(N262), .B(z2[243]), .Z(n207) );
  NANDN U306 ( .A(n3), .B(N507), .Z(n206) );
  NAND U307 ( .A(n208), .B(n209), .Z(z3[242]) );
  NANDN U308 ( .A(N262), .B(z2[242]), .Z(n209) );
  NANDN U309 ( .A(n3), .B(N506), .Z(n208) );
  NAND U310 ( .A(n210), .B(n211), .Z(z3[241]) );
  NANDN U311 ( .A(N262), .B(z2[241]), .Z(n211) );
  NANDN U312 ( .A(n3), .B(N505), .Z(n210) );
  NAND U313 ( .A(n212), .B(n213), .Z(z3[240]) );
  NANDN U314 ( .A(N262), .B(z2[240]), .Z(n213) );
  NANDN U315 ( .A(n3), .B(N504), .Z(n212) );
  NAND U316 ( .A(n214), .B(n215), .Z(z3[23]) );
  NANDN U317 ( .A(N262), .B(z2[23]), .Z(n215) );
  NANDN U318 ( .A(n3), .B(N287), .Z(n214) );
  NAND U319 ( .A(n216), .B(n217), .Z(z3[239]) );
  NANDN U320 ( .A(N262), .B(z2[239]), .Z(n217) );
  NANDN U321 ( .A(n3), .B(N503), .Z(n216) );
  NAND U322 ( .A(n218), .B(n219), .Z(z3[238]) );
  NANDN U323 ( .A(N262), .B(z2[238]), .Z(n219) );
  NANDN U324 ( .A(n3), .B(N502), .Z(n218) );
  NAND U325 ( .A(n220), .B(n221), .Z(z3[237]) );
  NANDN U326 ( .A(N262), .B(z2[237]), .Z(n221) );
  NANDN U327 ( .A(n3), .B(N501), .Z(n220) );
  NAND U328 ( .A(n222), .B(n223), .Z(z3[236]) );
  NANDN U329 ( .A(N262), .B(z2[236]), .Z(n223) );
  NANDN U330 ( .A(n3), .B(N500), .Z(n222) );
  NAND U331 ( .A(n224), .B(n225), .Z(z3[235]) );
  NANDN U332 ( .A(N262), .B(z2[235]), .Z(n225) );
  NANDN U333 ( .A(n3), .B(N499), .Z(n224) );
  NAND U334 ( .A(n226), .B(n227), .Z(z3[234]) );
  NANDN U335 ( .A(N262), .B(z2[234]), .Z(n227) );
  NANDN U336 ( .A(n3), .B(N498), .Z(n226) );
  NAND U337 ( .A(n228), .B(n229), .Z(z3[233]) );
  NANDN U338 ( .A(N262), .B(z2[233]), .Z(n229) );
  NANDN U339 ( .A(n3), .B(N497), .Z(n228) );
  NAND U340 ( .A(n230), .B(n231), .Z(z3[232]) );
  NANDN U341 ( .A(N262), .B(z2[232]), .Z(n231) );
  NANDN U342 ( .A(n3), .B(N496), .Z(n230) );
  NAND U343 ( .A(n232), .B(n233), .Z(z3[231]) );
  NANDN U344 ( .A(N262), .B(z2[231]), .Z(n233) );
  NANDN U345 ( .A(n3), .B(N495), .Z(n232) );
  NAND U346 ( .A(n234), .B(n235), .Z(z3[230]) );
  NANDN U347 ( .A(N262), .B(z2[230]), .Z(n235) );
  NANDN U348 ( .A(n3), .B(N494), .Z(n234) );
  NAND U349 ( .A(n236), .B(n237), .Z(z3[22]) );
  NANDN U350 ( .A(N262), .B(z2[22]), .Z(n237) );
  NANDN U351 ( .A(n3), .B(N286), .Z(n236) );
  NAND U352 ( .A(n238), .B(n239), .Z(z3[229]) );
  NANDN U353 ( .A(N262), .B(z2[229]), .Z(n239) );
  NANDN U354 ( .A(n3), .B(N493), .Z(n238) );
  NAND U355 ( .A(n240), .B(n241), .Z(z3[228]) );
  NANDN U356 ( .A(N262), .B(z2[228]), .Z(n241) );
  NANDN U357 ( .A(n3), .B(N492), .Z(n240) );
  NAND U358 ( .A(n242), .B(n243), .Z(z3[227]) );
  NANDN U359 ( .A(N262), .B(z2[227]), .Z(n243) );
  NANDN U360 ( .A(n3), .B(N491), .Z(n242) );
  NAND U361 ( .A(n244), .B(n245), .Z(z3[226]) );
  NANDN U362 ( .A(N262), .B(z2[226]), .Z(n245) );
  NANDN U363 ( .A(n3), .B(N490), .Z(n244) );
  NAND U364 ( .A(n246), .B(n247), .Z(z3[225]) );
  NANDN U365 ( .A(N262), .B(z2[225]), .Z(n247) );
  NANDN U366 ( .A(n3), .B(N489), .Z(n246) );
  NAND U367 ( .A(n248), .B(n249), .Z(z3[224]) );
  NANDN U368 ( .A(N262), .B(z2[224]), .Z(n249) );
  NANDN U369 ( .A(n3), .B(N488), .Z(n248) );
  NAND U370 ( .A(n250), .B(n251), .Z(z3[223]) );
  NANDN U371 ( .A(N262), .B(z2[223]), .Z(n251) );
  NANDN U372 ( .A(n3), .B(N487), .Z(n250) );
  NAND U373 ( .A(n252), .B(n253), .Z(z3[222]) );
  NANDN U374 ( .A(N262), .B(z2[222]), .Z(n253) );
  NANDN U375 ( .A(n3), .B(N486), .Z(n252) );
  NAND U376 ( .A(n254), .B(n255), .Z(z3[221]) );
  NANDN U377 ( .A(N262), .B(z2[221]), .Z(n255) );
  NANDN U378 ( .A(n3), .B(N485), .Z(n254) );
  NAND U379 ( .A(n256), .B(n257), .Z(z3[220]) );
  NANDN U380 ( .A(N262), .B(z2[220]), .Z(n257) );
  NANDN U381 ( .A(n3), .B(N484), .Z(n256) );
  NAND U382 ( .A(n258), .B(n259), .Z(z3[21]) );
  NANDN U383 ( .A(N262), .B(z2[21]), .Z(n259) );
  NANDN U384 ( .A(n3), .B(N285), .Z(n258) );
  NAND U385 ( .A(n260), .B(n261), .Z(z3[219]) );
  NANDN U386 ( .A(N262), .B(z2[219]), .Z(n261) );
  NANDN U387 ( .A(n3), .B(N483), .Z(n260) );
  NAND U388 ( .A(n262), .B(n263), .Z(z3[218]) );
  NANDN U389 ( .A(N262), .B(z2[218]), .Z(n263) );
  NANDN U390 ( .A(n3), .B(N482), .Z(n262) );
  NAND U391 ( .A(n264), .B(n265), .Z(z3[217]) );
  NANDN U392 ( .A(N262), .B(z2[217]), .Z(n265) );
  NANDN U393 ( .A(n3), .B(N481), .Z(n264) );
  NAND U394 ( .A(n266), .B(n267), .Z(z3[216]) );
  NANDN U395 ( .A(N262), .B(z2[216]), .Z(n267) );
  NANDN U396 ( .A(n3), .B(N480), .Z(n266) );
  NAND U397 ( .A(n268), .B(n269), .Z(z3[215]) );
  NANDN U398 ( .A(N262), .B(z2[215]), .Z(n269) );
  NANDN U399 ( .A(n3), .B(N479), .Z(n268) );
  NAND U400 ( .A(n270), .B(n271), .Z(z3[214]) );
  NANDN U401 ( .A(N262), .B(z2[214]), .Z(n271) );
  NANDN U402 ( .A(n3), .B(N478), .Z(n270) );
  NAND U403 ( .A(n272), .B(n273), .Z(z3[213]) );
  NANDN U404 ( .A(N262), .B(z2[213]), .Z(n273) );
  NANDN U405 ( .A(n3), .B(N477), .Z(n272) );
  NAND U406 ( .A(n274), .B(n275), .Z(z3[212]) );
  NANDN U407 ( .A(N262), .B(z2[212]), .Z(n275) );
  NANDN U408 ( .A(n3), .B(N476), .Z(n274) );
  NAND U409 ( .A(n276), .B(n277), .Z(z3[211]) );
  NANDN U410 ( .A(N262), .B(z2[211]), .Z(n277) );
  NANDN U411 ( .A(n3), .B(N475), .Z(n276) );
  NAND U412 ( .A(n278), .B(n279), .Z(z3[210]) );
  NANDN U413 ( .A(N262), .B(z2[210]), .Z(n279) );
  NANDN U414 ( .A(n3), .B(N474), .Z(n278) );
  NAND U415 ( .A(n280), .B(n281), .Z(z3[20]) );
  NANDN U416 ( .A(N262), .B(z2[20]), .Z(n281) );
  NANDN U417 ( .A(n3), .B(N284), .Z(n280) );
  NAND U418 ( .A(n282), .B(n283), .Z(z3[209]) );
  NANDN U419 ( .A(N262), .B(z2[209]), .Z(n283) );
  NANDN U420 ( .A(n3), .B(N473), .Z(n282) );
  NAND U421 ( .A(n284), .B(n285), .Z(z3[208]) );
  NANDN U422 ( .A(N262), .B(z2[208]), .Z(n285) );
  NANDN U423 ( .A(n3), .B(N472), .Z(n284) );
  NAND U424 ( .A(n286), .B(n287), .Z(z3[207]) );
  NANDN U425 ( .A(N262), .B(z2[207]), .Z(n287) );
  NANDN U426 ( .A(n3), .B(N471), .Z(n286) );
  NAND U427 ( .A(n288), .B(n289), .Z(z3[206]) );
  NANDN U428 ( .A(N262), .B(z2[206]), .Z(n289) );
  NANDN U429 ( .A(n3), .B(N470), .Z(n288) );
  NAND U430 ( .A(n290), .B(n291), .Z(z3[205]) );
  NANDN U431 ( .A(N262), .B(z2[205]), .Z(n291) );
  NANDN U432 ( .A(n3), .B(N469), .Z(n290) );
  NAND U433 ( .A(n292), .B(n293), .Z(z3[204]) );
  NANDN U434 ( .A(N262), .B(z2[204]), .Z(n293) );
  NANDN U435 ( .A(n3), .B(N468), .Z(n292) );
  NAND U436 ( .A(n294), .B(n295), .Z(z3[203]) );
  NANDN U437 ( .A(N262), .B(z2[203]), .Z(n295) );
  NANDN U438 ( .A(n3), .B(N467), .Z(n294) );
  NAND U439 ( .A(n296), .B(n297), .Z(z3[202]) );
  NANDN U440 ( .A(N262), .B(z2[202]), .Z(n297) );
  NANDN U441 ( .A(n3), .B(N466), .Z(n296) );
  NAND U442 ( .A(n298), .B(n299), .Z(z3[201]) );
  NANDN U443 ( .A(N262), .B(z2[201]), .Z(n299) );
  NANDN U444 ( .A(n3), .B(N465), .Z(n298) );
  NAND U445 ( .A(n300), .B(n301), .Z(z3[200]) );
  NANDN U446 ( .A(N262), .B(z2[200]), .Z(n301) );
  NANDN U447 ( .A(n3), .B(N464), .Z(n300) );
  NAND U448 ( .A(n302), .B(n303), .Z(z3[1]) );
  NANDN U449 ( .A(N262), .B(z2[1]), .Z(n303) );
  NANDN U450 ( .A(n3), .B(N265), .Z(n302) );
  NAND U451 ( .A(n304), .B(n305), .Z(z3[19]) );
  NANDN U452 ( .A(N262), .B(z2[19]), .Z(n305) );
  NANDN U453 ( .A(n3), .B(N283), .Z(n304) );
  NAND U454 ( .A(n306), .B(n307), .Z(z3[199]) );
  NANDN U455 ( .A(N262), .B(z2[199]), .Z(n307) );
  NANDN U456 ( .A(n3), .B(N463), .Z(n306) );
  NAND U457 ( .A(n308), .B(n309), .Z(z3[198]) );
  NANDN U458 ( .A(N262), .B(z2[198]), .Z(n309) );
  NANDN U459 ( .A(n3), .B(N462), .Z(n308) );
  NAND U460 ( .A(n310), .B(n311), .Z(z3[197]) );
  NANDN U461 ( .A(N262), .B(z2[197]), .Z(n311) );
  NANDN U462 ( .A(n3), .B(N461), .Z(n310) );
  NAND U463 ( .A(n312), .B(n313), .Z(z3[196]) );
  NANDN U464 ( .A(N262), .B(z2[196]), .Z(n313) );
  NANDN U465 ( .A(n3), .B(N460), .Z(n312) );
  NAND U466 ( .A(n314), .B(n315), .Z(z3[195]) );
  NANDN U467 ( .A(N262), .B(z2[195]), .Z(n315) );
  NANDN U468 ( .A(n3), .B(N459), .Z(n314) );
  NAND U469 ( .A(n316), .B(n317), .Z(z3[194]) );
  NANDN U470 ( .A(N262), .B(z2[194]), .Z(n317) );
  NANDN U471 ( .A(n3), .B(N458), .Z(n316) );
  NAND U472 ( .A(n318), .B(n319), .Z(z3[193]) );
  NANDN U473 ( .A(N262), .B(z2[193]), .Z(n319) );
  NANDN U474 ( .A(n3), .B(N457), .Z(n318) );
  NAND U475 ( .A(n320), .B(n321), .Z(z3[192]) );
  NANDN U476 ( .A(N262), .B(z2[192]), .Z(n321) );
  NANDN U477 ( .A(n3), .B(N456), .Z(n320) );
  NAND U478 ( .A(n322), .B(n323), .Z(z3[191]) );
  NANDN U479 ( .A(N262), .B(z2[191]), .Z(n323) );
  NANDN U480 ( .A(n3), .B(N455), .Z(n322) );
  NAND U481 ( .A(n324), .B(n325), .Z(z3[190]) );
  NANDN U482 ( .A(N262), .B(z2[190]), .Z(n325) );
  NANDN U483 ( .A(n3), .B(N454), .Z(n324) );
  NAND U484 ( .A(n326), .B(n327), .Z(z3[18]) );
  NANDN U485 ( .A(N262), .B(z2[18]), .Z(n327) );
  NANDN U486 ( .A(n3), .B(N282), .Z(n326) );
  NAND U487 ( .A(n328), .B(n329), .Z(z3[189]) );
  NANDN U488 ( .A(N262), .B(z2[189]), .Z(n329) );
  NANDN U489 ( .A(n3), .B(N453), .Z(n328) );
  NAND U490 ( .A(n330), .B(n331), .Z(z3[188]) );
  NANDN U491 ( .A(N262), .B(z2[188]), .Z(n331) );
  NANDN U492 ( .A(n3), .B(N452), .Z(n330) );
  NAND U493 ( .A(n332), .B(n333), .Z(z3[187]) );
  NANDN U494 ( .A(N262), .B(z2[187]), .Z(n333) );
  NANDN U495 ( .A(n3), .B(N451), .Z(n332) );
  NAND U496 ( .A(n334), .B(n335), .Z(z3[186]) );
  NANDN U497 ( .A(N262), .B(z2[186]), .Z(n335) );
  NANDN U498 ( .A(n3), .B(N450), .Z(n334) );
  NAND U499 ( .A(n336), .B(n337), .Z(z3[185]) );
  NANDN U500 ( .A(N262), .B(z2[185]), .Z(n337) );
  NANDN U501 ( .A(n3), .B(N449), .Z(n336) );
  NAND U502 ( .A(n338), .B(n339), .Z(z3[184]) );
  NANDN U503 ( .A(N262), .B(z2[184]), .Z(n339) );
  NANDN U504 ( .A(n3), .B(N448), .Z(n338) );
  NAND U505 ( .A(n340), .B(n341), .Z(z3[183]) );
  NANDN U506 ( .A(N262), .B(z2[183]), .Z(n341) );
  NANDN U507 ( .A(n3), .B(N447), .Z(n340) );
  NAND U508 ( .A(n342), .B(n343), .Z(z3[182]) );
  NANDN U509 ( .A(N262), .B(z2[182]), .Z(n343) );
  NANDN U510 ( .A(n3), .B(N446), .Z(n342) );
  NAND U511 ( .A(n344), .B(n345), .Z(z3[181]) );
  NANDN U512 ( .A(N262), .B(z2[181]), .Z(n345) );
  NANDN U513 ( .A(n3), .B(N445), .Z(n344) );
  NAND U514 ( .A(n346), .B(n347), .Z(z3[180]) );
  NANDN U515 ( .A(N262), .B(z2[180]), .Z(n347) );
  NANDN U516 ( .A(n3), .B(N444), .Z(n346) );
  NAND U517 ( .A(n348), .B(n349), .Z(z3[17]) );
  NANDN U518 ( .A(N262), .B(z2[17]), .Z(n349) );
  NANDN U519 ( .A(n3), .B(N281), .Z(n348) );
  NAND U520 ( .A(n350), .B(n351), .Z(z3[179]) );
  NANDN U521 ( .A(N262), .B(z2[179]), .Z(n351) );
  NANDN U522 ( .A(n3), .B(N443), .Z(n350) );
  NAND U523 ( .A(n352), .B(n353), .Z(z3[178]) );
  NANDN U524 ( .A(N262), .B(z2[178]), .Z(n353) );
  NANDN U525 ( .A(n3), .B(N442), .Z(n352) );
  NAND U526 ( .A(n354), .B(n355), .Z(z3[177]) );
  NANDN U527 ( .A(N262), .B(z2[177]), .Z(n355) );
  NANDN U528 ( .A(n3), .B(N441), .Z(n354) );
  NAND U529 ( .A(n356), .B(n357), .Z(z3[176]) );
  NANDN U530 ( .A(N262), .B(z2[176]), .Z(n357) );
  NANDN U531 ( .A(n3), .B(N440), .Z(n356) );
  NAND U532 ( .A(n358), .B(n359), .Z(z3[175]) );
  NANDN U533 ( .A(N262), .B(z2[175]), .Z(n359) );
  NANDN U534 ( .A(n3), .B(N439), .Z(n358) );
  NAND U535 ( .A(n360), .B(n361), .Z(z3[174]) );
  NANDN U536 ( .A(N262), .B(z2[174]), .Z(n361) );
  NANDN U537 ( .A(n3), .B(N438), .Z(n360) );
  NAND U538 ( .A(n362), .B(n363), .Z(z3[173]) );
  NANDN U539 ( .A(N262), .B(z2[173]), .Z(n363) );
  NANDN U540 ( .A(n3), .B(N437), .Z(n362) );
  NAND U541 ( .A(n364), .B(n365), .Z(z3[172]) );
  NANDN U542 ( .A(N262), .B(z2[172]), .Z(n365) );
  NANDN U543 ( .A(n3), .B(N436), .Z(n364) );
  NAND U544 ( .A(n366), .B(n367), .Z(z3[171]) );
  NANDN U545 ( .A(N262), .B(z2[171]), .Z(n367) );
  NANDN U546 ( .A(n3), .B(N435), .Z(n366) );
  NAND U547 ( .A(n368), .B(n369), .Z(z3[170]) );
  NANDN U548 ( .A(N262), .B(z2[170]), .Z(n369) );
  NANDN U549 ( .A(n3), .B(N434), .Z(n368) );
  NAND U550 ( .A(n370), .B(n371), .Z(z3[16]) );
  NANDN U551 ( .A(N262), .B(z2[16]), .Z(n371) );
  NANDN U552 ( .A(n3), .B(N280), .Z(n370) );
  NAND U553 ( .A(n372), .B(n373), .Z(z3[169]) );
  NANDN U554 ( .A(N262), .B(z2[169]), .Z(n373) );
  NANDN U555 ( .A(n3), .B(N433), .Z(n372) );
  NAND U556 ( .A(n374), .B(n375), .Z(z3[168]) );
  NANDN U557 ( .A(N262), .B(z2[168]), .Z(n375) );
  NANDN U558 ( .A(n3), .B(N432), .Z(n374) );
  NAND U559 ( .A(n376), .B(n377), .Z(z3[167]) );
  NANDN U560 ( .A(N262), .B(z2[167]), .Z(n377) );
  NANDN U561 ( .A(n3), .B(N431), .Z(n376) );
  NAND U562 ( .A(n378), .B(n379), .Z(z3[166]) );
  NANDN U563 ( .A(N262), .B(z2[166]), .Z(n379) );
  NANDN U564 ( .A(n3), .B(N430), .Z(n378) );
  NAND U565 ( .A(n380), .B(n381), .Z(z3[165]) );
  NANDN U566 ( .A(N262), .B(z2[165]), .Z(n381) );
  NANDN U567 ( .A(n3), .B(N429), .Z(n380) );
  NAND U568 ( .A(n382), .B(n383), .Z(z3[164]) );
  NANDN U569 ( .A(N262), .B(z2[164]), .Z(n383) );
  NANDN U570 ( .A(n3), .B(N428), .Z(n382) );
  NAND U571 ( .A(n384), .B(n385), .Z(z3[163]) );
  NANDN U572 ( .A(N262), .B(z2[163]), .Z(n385) );
  NANDN U573 ( .A(n3), .B(N427), .Z(n384) );
  NAND U574 ( .A(n386), .B(n387), .Z(z3[162]) );
  NANDN U575 ( .A(N262), .B(z2[162]), .Z(n387) );
  NANDN U576 ( .A(n3), .B(N426), .Z(n386) );
  NAND U577 ( .A(n388), .B(n389), .Z(z3[161]) );
  NANDN U578 ( .A(N262), .B(z2[161]), .Z(n389) );
  NANDN U579 ( .A(n3), .B(N425), .Z(n388) );
  NAND U580 ( .A(n390), .B(n391), .Z(z3[160]) );
  NANDN U581 ( .A(N262), .B(z2[160]), .Z(n391) );
  NANDN U582 ( .A(n3), .B(N424), .Z(n390) );
  NAND U583 ( .A(n392), .B(n393), .Z(z3[15]) );
  NANDN U584 ( .A(N262), .B(z2[15]), .Z(n393) );
  NANDN U585 ( .A(n3), .B(N279), .Z(n392) );
  NAND U586 ( .A(n394), .B(n395), .Z(z3[159]) );
  NANDN U587 ( .A(N262), .B(z2[159]), .Z(n395) );
  NANDN U588 ( .A(n3), .B(N423), .Z(n394) );
  NAND U589 ( .A(n396), .B(n397), .Z(z3[158]) );
  NANDN U590 ( .A(N262), .B(z2[158]), .Z(n397) );
  NANDN U591 ( .A(n3), .B(N422), .Z(n396) );
  NAND U592 ( .A(n398), .B(n399), .Z(z3[157]) );
  NANDN U593 ( .A(N262), .B(z2[157]), .Z(n399) );
  NANDN U594 ( .A(n3), .B(N421), .Z(n398) );
  NAND U595 ( .A(n400), .B(n401), .Z(z3[156]) );
  NANDN U596 ( .A(N262), .B(z2[156]), .Z(n401) );
  NANDN U597 ( .A(n3), .B(N420), .Z(n400) );
  NAND U598 ( .A(n402), .B(n403), .Z(z3[155]) );
  NANDN U599 ( .A(N262), .B(z2[155]), .Z(n403) );
  NANDN U600 ( .A(n3), .B(N419), .Z(n402) );
  NAND U601 ( .A(n404), .B(n405), .Z(z3[154]) );
  NANDN U602 ( .A(N262), .B(z2[154]), .Z(n405) );
  NANDN U603 ( .A(n3), .B(N418), .Z(n404) );
  NAND U604 ( .A(n406), .B(n407), .Z(z3[153]) );
  NANDN U605 ( .A(N262), .B(z2[153]), .Z(n407) );
  NANDN U606 ( .A(n3), .B(N417), .Z(n406) );
  NAND U607 ( .A(n408), .B(n409), .Z(z3[152]) );
  NANDN U608 ( .A(N262), .B(z2[152]), .Z(n409) );
  NANDN U609 ( .A(n3), .B(N416), .Z(n408) );
  NAND U610 ( .A(n410), .B(n411), .Z(z3[151]) );
  NANDN U611 ( .A(N262), .B(z2[151]), .Z(n411) );
  NANDN U612 ( .A(n3), .B(N415), .Z(n410) );
  NAND U613 ( .A(n412), .B(n413), .Z(z3[150]) );
  NANDN U614 ( .A(N262), .B(z2[150]), .Z(n413) );
  NANDN U615 ( .A(n3), .B(N414), .Z(n412) );
  NAND U616 ( .A(n414), .B(n415), .Z(z3[14]) );
  NANDN U617 ( .A(N262), .B(z2[14]), .Z(n415) );
  NANDN U618 ( .A(n3), .B(N278), .Z(n414) );
  NAND U619 ( .A(n416), .B(n417), .Z(z3[149]) );
  NANDN U620 ( .A(N262), .B(z2[149]), .Z(n417) );
  NANDN U621 ( .A(n3), .B(N413), .Z(n416) );
  NAND U622 ( .A(n418), .B(n419), .Z(z3[148]) );
  NANDN U623 ( .A(N262), .B(z2[148]), .Z(n419) );
  NANDN U624 ( .A(n3), .B(N412), .Z(n418) );
  NAND U625 ( .A(n420), .B(n421), .Z(z3[147]) );
  NANDN U626 ( .A(N262), .B(z2[147]), .Z(n421) );
  NANDN U627 ( .A(n3), .B(N411), .Z(n420) );
  NAND U628 ( .A(n422), .B(n423), .Z(z3[146]) );
  NANDN U629 ( .A(N262), .B(z2[146]), .Z(n423) );
  NANDN U630 ( .A(n3), .B(N410), .Z(n422) );
  NAND U631 ( .A(n424), .B(n425), .Z(z3[145]) );
  NANDN U632 ( .A(N262), .B(z2[145]), .Z(n425) );
  NANDN U633 ( .A(n3), .B(N409), .Z(n424) );
  NAND U634 ( .A(n426), .B(n427), .Z(z3[144]) );
  NANDN U635 ( .A(N262), .B(z2[144]), .Z(n427) );
  NANDN U636 ( .A(n3), .B(N408), .Z(n426) );
  NAND U637 ( .A(n428), .B(n429), .Z(z3[143]) );
  NANDN U638 ( .A(N262), .B(z2[143]), .Z(n429) );
  NANDN U639 ( .A(n3), .B(N407), .Z(n428) );
  NAND U640 ( .A(n430), .B(n431), .Z(z3[142]) );
  NANDN U641 ( .A(N262), .B(z2[142]), .Z(n431) );
  NANDN U642 ( .A(n3), .B(N406), .Z(n430) );
  NAND U643 ( .A(n432), .B(n433), .Z(z3[141]) );
  NANDN U644 ( .A(N262), .B(z2[141]), .Z(n433) );
  NANDN U645 ( .A(n3), .B(N405), .Z(n432) );
  NAND U646 ( .A(n434), .B(n435), .Z(z3[140]) );
  NANDN U647 ( .A(N262), .B(z2[140]), .Z(n435) );
  NANDN U648 ( .A(n3), .B(N404), .Z(n434) );
  NAND U649 ( .A(n436), .B(n437), .Z(z3[13]) );
  NANDN U650 ( .A(N262), .B(z2[13]), .Z(n437) );
  NANDN U651 ( .A(n3), .B(N277), .Z(n436) );
  NAND U652 ( .A(n438), .B(n439), .Z(z3[139]) );
  NANDN U653 ( .A(N262), .B(z2[139]), .Z(n439) );
  NANDN U654 ( .A(n3), .B(N403), .Z(n438) );
  NAND U655 ( .A(n440), .B(n441), .Z(z3[138]) );
  NANDN U656 ( .A(N262), .B(z2[138]), .Z(n441) );
  NANDN U657 ( .A(n3), .B(N402), .Z(n440) );
  NAND U658 ( .A(n442), .B(n443), .Z(z3[137]) );
  NANDN U659 ( .A(N262), .B(z2[137]), .Z(n443) );
  NANDN U660 ( .A(n3), .B(N401), .Z(n442) );
  NAND U661 ( .A(n444), .B(n445), .Z(z3[136]) );
  NANDN U662 ( .A(N262), .B(z2[136]), .Z(n445) );
  NANDN U663 ( .A(n3), .B(N400), .Z(n444) );
  NAND U664 ( .A(n446), .B(n447), .Z(z3[135]) );
  NANDN U665 ( .A(N262), .B(z2[135]), .Z(n447) );
  NANDN U666 ( .A(n3), .B(N399), .Z(n446) );
  NAND U667 ( .A(n448), .B(n449), .Z(z3[134]) );
  NANDN U668 ( .A(N262), .B(z2[134]), .Z(n449) );
  NANDN U669 ( .A(n3), .B(N398), .Z(n448) );
  NAND U670 ( .A(n450), .B(n451), .Z(z3[133]) );
  NANDN U671 ( .A(N262), .B(z2[133]), .Z(n451) );
  NANDN U672 ( .A(n3), .B(N397), .Z(n450) );
  NAND U673 ( .A(n452), .B(n453), .Z(z3[132]) );
  NANDN U674 ( .A(N262), .B(z2[132]), .Z(n453) );
  NANDN U675 ( .A(n3), .B(N396), .Z(n452) );
  NAND U676 ( .A(n454), .B(n455), .Z(z3[131]) );
  NANDN U677 ( .A(N262), .B(z2[131]), .Z(n455) );
  NANDN U678 ( .A(n3), .B(N395), .Z(n454) );
  NAND U679 ( .A(n456), .B(n457), .Z(z3[130]) );
  NANDN U680 ( .A(N262), .B(z2[130]), .Z(n457) );
  NANDN U681 ( .A(n3), .B(N394), .Z(n456) );
  NAND U682 ( .A(n458), .B(n459), .Z(z3[12]) );
  NANDN U683 ( .A(N262), .B(z2[12]), .Z(n459) );
  NANDN U684 ( .A(n3), .B(N276), .Z(n458) );
  NAND U685 ( .A(n460), .B(n461), .Z(z3[129]) );
  NANDN U686 ( .A(N262), .B(z2[129]), .Z(n461) );
  NANDN U687 ( .A(n3), .B(N393), .Z(n460) );
  NAND U688 ( .A(n462), .B(n463), .Z(z3[128]) );
  NANDN U689 ( .A(N262), .B(z2[128]), .Z(n463) );
  NANDN U690 ( .A(n3), .B(N392), .Z(n462) );
  NAND U691 ( .A(n464), .B(n465), .Z(z3[127]) );
  NANDN U692 ( .A(N262), .B(z2[127]), .Z(n465) );
  NANDN U693 ( .A(n3), .B(N391), .Z(n464) );
  NAND U694 ( .A(n466), .B(n467), .Z(z3[126]) );
  NANDN U695 ( .A(N262), .B(z2[126]), .Z(n467) );
  NANDN U696 ( .A(n3), .B(N390), .Z(n466) );
  NAND U697 ( .A(n468), .B(n469), .Z(z3[125]) );
  NANDN U698 ( .A(N262), .B(z2[125]), .Z(n469) );
  NANDN U699 ( .A(n3), .B(N389), .Z(n468) );
  NAND U700 ( .A(n470), .B(n471), .Z(z3[124]) );
  NANDN U701 ( .A(N262), .B(z2[124]), .Z(n471) );
  NANDN U702 ( .A(n3), .B(N388), .Z(n470) );
  NAND U703 ( .A(n472), .B(n473), .Z(z3[123]) );
  NANDN U704 ( .A(N262), .B(z2[123]), .Z(n473) );
  NANDN U705 ( .A(n3), .B(N387), .Z(n472) );
  NAND U706 ( .A(n474), .B(n475), .Z(z3[122]) );
  NANDN U707 ( .A(N262), .B(z2[122]), .Z(n475) );
  NANDN U708 ( .A(n3), .B(N386), .Z(n474) );
  NAND U709 ( .A(n476), .B(n477), .Z(z3[121]) );
  NANDN U710 ( .A(N262), .B(z2[121]), .Z(n477) );
  NANDN U711 ( .A(n3), .B(N385), .Z(n476) );
  NAND U712 ( .A(n478), .B(n479), .Z(z3[120]) );
  NANDN U713 ( .A(N262), .B(z2[120]), .Z(n479) );
  NANDN U714 ( .A(n3), .B(N384), .Z(n478) );
  NAND U715 ( .A(n480), .B(n481), .Z(z3[11]) );
  NANDN U716 ( .A(N262), .B(z2[11]), .Z(n481) );
  NANDN U717 ( .A(n3), .B(N275), .Z(n480) );
  NAND U718 ( .A(n482), .B(n483), .Z(z3[119]) );
  NANDN U719 ( .A(N262), .B(z2[119]), .Z(n483) );
  NANDN U720 ( .A(n3), .B(N383), .Z(n482) );
  NAND U721 ( .A(n484), .B(n485), .Z(z3[118]) );
  NANDN U722 ( .A(N262), .B(z2[118]), .Z(n485) );
  NANDN U723 ( .A(n3), .B(N382), .Z(n484) );
  NAND U724 ( .A(n486), .B(n487), .Z(z3[117]) );
  NANDN U725 ( .A(N262), .B(z2[117]), .Z(n487) );
  NANDN U726 ( .A(n3), .B(N381), .Z(n486) );
  NAND U727 ( .A(n488), .B(n489), .Z(z3[116]) );
  NANDN U728 ( .A(N262), .B(z2[116]), .Z(n489) );
  NANDN U729 ( .A(n3), .B(N380), .Z(n488) );
  NAND U730 ( .A(n490), .B(n491), .Z(z3[115]) );
  NANDN U731 ( .A(N262), .B(z2[115]), .Z(n491) );
  NANDN U732 ( .A(n3), .B(N379), .Z(n490) );
  NAND U733 ( .A(n492), .B(n493), .Z(z3[114]) );
  NANDN U734 ( .A(N262), .B(z2[114]), .Z(n493) );
  NANDN U735 ( .A(n3), .B(N378), .Z(n492) );
  NAND U736 ( .A(n494), .B(n495), .Z(z3[113]) );
  NANDN U737 ( .A(N262), .B(z2[113]), .Z(n495) );
  NANDN U738 ( .A(n3), .B(N377), .Z(n494) );
  NAND U739 ( .A(n496), .B(n497), .Z(z3[112]) );
  NANDN U740 ( .A(N262), .B(z2[112]), .Z(n497) );
  NANDN U741 ( .A(n3), .B(N376), .Z(n496) );
  NAND U742 ( .A(n498), .B(n499), .Z(z3[111]) );
  NANDN U743 ( .A(N262), .B(z2[111]), .Z(n499) );
  NANDN U744 ( .A(n3), .B(N375), .Z(n498) );
  NAND U745 ( .A(n500), .B(n501), .Z(z3[110]) );
  NANDN U746 ( .A(N262), .B(z2[110]), .Z(n501) );
  NANDN U747 ( .A(n3), .B(N374), .Z(n500) );
  NAND U748 ( .A(n502), .B(n503), .Z(z3[10]) );
  NANDN U749 ( .A(N262), .B(z2[10]), .Z(n503) );
  NANDN U750 ( .A(n3), .B(N274), .Z(n502) );
  NAND U751 ( .A(n504), .B(n505), .Z(z3[109]) );
  NANDN U752 ( .A(N262), .B(z2[109]), .Z(n505) );
  NANDN U753 ( .A(n3), .B(N373), .Z(n504) );
  NAND U754 ( .A(n506), .B(n507), .Z(z3[108]) );
  NANDN U755 ( .A(N262), .B(z2[108]), .Z(n507) );
  NANDN U756 ( .A(n3), .B(N372), .Z(n506) );
  NAND U757 ( .A(n508), .B(n509), .Z(z3[107]) );
  NANDN U758 ( .A(N262), .B(z2[107]), .Z(n509) );
  NANDN U759 ( .A(n3), .B(N371), .Z(n508) );
  NAND U760 ( .A(n510), .B(n511), .Z(z3[106]) );
  NANDN U761 ( .A(N262), .B(z2[106]), .Z(n511) );
  NANDN U762 ( .A(n3), .B(N370), .Z(n510) );
  NAND U763 ( .A(n512), .B(n513), .Z(z3[105]) );
  NANDN U764 ( .A(N262), .B(z2[105]), .Z(n513) );
  NANDN U765 ( .A(n3), .B(N369), .Z(n512) );
  NAND U766 ( .A(n514), .B(n515), .Z(z3[104]) );
  NANDN U767 ( .A(N262), .B(z2[104]), .Z(n515) );
  NANDN U768 ( .A(n3), .B(N368), .Z(n514) );
  NAND U769 ( .A(n516), .B(n517), .Z(z3[103]) );
  NANDN U770 ( .A(N262), .B(z2[103]), .Z(n517) );
  NANDN U771 ( .A(n3), .B(N367), .Z(n516) );
  NAND U772 ( .A(n518), .B(n519), .Z(z3[102]) );
  NANDN U773 ( .A(N262), .B(z2[102]), .Z(n519) );
  NANDN U774 ( .A(n3), .B(N366), .Z(n518) );
  NAND U775 ( .A(n520), .B(n521), .Z(z3[101]) );
  NANDN U776 ( .A(N262), .B(z2[101]), .Z(n521) );
  NANDN U777 ( .A(n3), .B(N365), .Z(n520) );
  NAND U778 ( .A(n522), .B(n523), .Z(z3[100]) );
  NANDN U779 ( .A(N262), .B(z2[100]), .Z(n523) );
  NANDN U780 ( .A(n3), .B(N364), .Z(n522) );
  NAND U781 ( .A(n524), .B(n525), .Z(z3[0]) );
  NANDN U782 ( .A(N262), .B(z2[0]), .Z(n525) );
  NANDN U783 ( .A(n3), .B(N264), .Z(n524) );
  IV U784 ( .A(N262), .Z(n3) );
  NAND U785 ( .A(n526), .B(n527), .Z(z2[9]) );
  NANDN U786 ( .A(xregN_1), .B(zin[8]), .Z(n527) );
  NAND U787 ( .A(N13), .B(xregN_1), .Z(n526) );
  NAND U788 ( .A(n528), .B(n529), .Z(z2[99]) );
  NANDN U789 ( .A(xregN_1), .B(zin[98]), .Z(n529) );
  NAND U790 ( .A(N103), .B(xregN_1), .Z(n528) );
  NAND U791 ( .A(n530), .B(n531), .Z(z2[98]) );
  NANDN U792 ( .A(xregN_1), .B(zin[97]), .Z(n531) );
  NAND U793 ( .A(N102), .B(xregN_1), .Z(n530) );
  NAND U794 ( .A(n532), .B(n533), .Z(z2[97]) );
  NANDN U795 ( .A(xregN_1), .B(zin[96]), .Z(n533) );
  NAND U796 ( .A(N101), .B(xregN_1), .Z(n532) );
  NAND U797 ( .A(n534), .B(n535), .Z(z2[96]) );
  NANDN U798 ( .A(xregN_1), .B(zin[95]), .Z(n535) );
  NAND U799 ( .A(N100), .B(xregN_1), .Z(n534) );
  NAND U800 ( .A(n536), .B(n537), .Z(z2[95]) );
  NANDN U801 ( .A(xregN_1), .B(zin[94]), .Z(n537) );
  NAND U802 ( .A(N99), .B(xregN_1), .Z(n536) );
  NAND U803 ( .A(n538), .B(n539), .Z(z2[94]) );
  NANDN U804 ( .A(xregN_1), .B(zin[93]), .Z(n539) );
  NAND U805 ( .A(N98), .B(xregN_1), .Z(n538) );
  NAND U806 ( .A(n540), .B(n541), .Z(z2[93]) );
  NANDN U807 ( .A(xregN_1), .B(zin[92]), .Z(n541) );
  NAND U808 ( .A(N97), .B(xregN_1), .Z(n540) );
  NAND U809 ( .A(n542), .B(n543), .Z(z2[92]) );
  NANDN U810 ( .A(xregN_1), .B(zin[91]), .Z(n543) );
  NAND U811 ( .A(N96), .B(xregN_1), .Z(n542) );
  NAND U812 ( .A(n544), .B(n545), .Z(z2[91]) );
  NANDN U813 ( .A(xregN_1), .B(zin[90]), .Z(n545) );
  NAND U814 ( .A(N95), .B(xregN_1), .Z(n544) );
  NAND U815 ( .A(n546), .B(n547), .Z(z2[90]) );
  NANDN U816 ( .A(xregN_1), .B(zin[89]), .Z(n547) );
  NAND U817 ( .A(N94), .B(xregN_1), .Z(n546) );
  NAND U818 ( .A(n548), .B(n549), .Z(z2[8]) );
  NANDN U819 ( .A(xregN_1), .B(zin[7]), .Z(n549) );
  NAND U820 ( .A(N12), .B(xregN_1), .Z(n548) );
  NAND U821 ( .A(n550), .B(n551), .Z(z2[89]) );
  NANDN U822 ( .A(xregN_1), .B(zin[88]), .Z(n551) );
  NAND U823 ( .A(N93), .B(xregN_1), .Z(n550) );
  NAND U824 ( .A(n552), .B(n553), .Z(z2[88]) );
  NANDN U825 ( .A(xregN_1), .B(zin[87]), .Z(n553) );
  NAND U826 ( .A(N92), .B(xregN_1), .Z(n552) );
  NAND U827 ( .A(n554), .B(n555), .Z(z2[87]) );
  NANDN U828 ( .A(xregN_1), .B(zin[86]), .Z(n555) );
  NAND U829 ( .A(N91), .B(xregN_1), .Z(n554) );
  NAND U830 ( .A(n556), .B(n557), .Z(z2[86]) );
  NANDN U831 ( .A(xregN_1), .B(zin[85]), .Z(n557) );
  NAND U832 ( .A(N90), .B(xregN_1), .Z(n556) );
  NAND U833 ( .A(n558), .B(n559), .Z(z2[85]) );
  NANDN U834 ( .A(xregN_1), .B(zin[84]), .Z(n559) );
  NAND U835 ( .A(N89), .B(xregN_1), .Z(n558) );
  NAND U836 ( .A(n560), .B(n561), .Z(z2[84]) );
  NANDN U837 ( .A(xregN_1), .B(zin[83]), .Z(n561) );
  NAND U838 ( .A(N88), .B(xregN_1), .Z(n560) );
  NAND U839 ( .A(n562), .B(n563), .Z(z2[83]) );
  NANDN U840 ( .A(xregN_1), .B(zin[82]), .Z(n563) );
  NAND U841 ( .A(N87), .B(xregN_1), .Z(n562) );
  NAND U842 ( .A(n564), .B(n565), .Z(z2[82]) );
  NANDN U843 ( .A(xregN_1), .B(zin[81]), .Z(n565) );
  NAND U844 ( .A(N86), .B(xregN_1), .Z(n564) );
  NAND U845 ( .A(n566), .B(n567), .Z(z2[81]) );
  NANDN U846 ( .A(xregN_1), .B(zin[80]), .Z(n567) );
  NAND U847 ( .A(N85), .B(xregN_1), .Z(n566) );
  NAND U848 ( .A(n568), .B(n569), .Z(z2[80]) );
  NANDN U849 ( .A(xregN_1), .B(zin[79]), .Z(n569) );
  NAND U850 ( .A(N84), .B(xregN_1), .Z(n568) );
  NAND U851 ( .A(n570), .B(n571), .Z(z2[7]) );
  NANDN U852 ( .A(xregN_1), .B(zin[6]), .Z(n571) );
  NAND U853 ( .A(N11), .B(xregN_1), .Z(n570) );
  NAND U854 ( .A(n572), .B(n573), .Z(z2[79]) );
  NANDN U855 ( .A(xregN_1), .B(zin[78]), .Z(n573) );
  NAND U856 ( .A(N83), .B(xregN_1), .Z(n572) );
  NAND U857 ( .A(n574), .B(n575), .Z(z2[78]) );
  NANDN U858 ( .A(xregN_1), .B(zin[77]), .Z(n575) );
  NAND U859 ( .A(N82), .B(xregN_1), .Z(n574) );
  NAND U860 ( .A(n576), .B(n577), .Z(z2[77]) );
  NANDN U861 ( .A(xregN_1), .B(zin[76]), .Z(n577) );
  NAND U862 ( .A(N81), .B(xregN_1), .Z(n576) );
  NAND U863 ( .A(n578), .B(n579), .Z(z2[76]) );
  NANDN U864 ( .A(xregN_1), .B(zin[75]), .Z(n579) );
  NAND U865 ( .A(N80), .B(xregN_1), .Z(n578) );
  NAND U866 ( .A(n580), .B(n581), .Z(z2[75]) );
  NANDN U867 ( .A(xregN_1), .B(zin[74]), .Z(n581) );
  NAND U868 ( .A(N79), .B(xregN_1), .Z(n580) );
  NAND U869 ( .A(n582), .B(n583), .Z(z2[74]) );
  NANDN U870 ( .A(xregN_1), .B(zin[73]), .Z(n583) );
  NAND U871 ( .A(N78), .B(xregN_1), .Z(n582) );
  NAND U872 ( .A(n584), .B(n585), .Z(z2[73]) );
  NANDN U873 ( .A(xregN_1), .B(zin[72]), .Z(n585) );
  NAND U874 ( .A(N77), .B(xregN_1), .Z(n584) );
  NAND U875 ( .A(n586), .B(n587), .Z(z2[72]) );
  NANDN U876 ( .A(xregN_1), .B(zin[71]), .Z(n587) );
  NAND U877 ( .A(N76), .B(xregN_1), .Z(n586) );
  NAND U878 ( .A(n588), .B(n589), .Z(z2[71]) );
  NANDN U879 ( .A(xregN_1), .B(zin[70]), .Z(n589) );
  NAND U880 ( .A(N75), .B(xregN_1), .Z(n588) );
  NAND U881 ( .A(n590), .B(n591), .Z(z2[70]) );
  NANDN U882 ( .A(xregN_1), .B(zin[69]), .Z(n591) );
  NAND U883 ( .A(N74), .B(xregN_1), .Z(n590) );
  NAND U884 ( .A(n592), .B(n593), .Z(z2[6]) );
  NANDN U885 ( .A(xregN_1), .B(zin[5]), .Z(n593) );
  NAND U886 ( .A(N10), .B(xregN_1), .Z(n592) );
  NAND U887 ( .A(n594), .B(n595), .Z(z2[69]) );
  NANDN U888 ( .A(xregN_1), .B(zin[68]), .Z(n595) );
  NAND U889 ( .A(N73), .B(xregN_1), .Z(n594) );
  NAND U890 ( .A(n596), .B(n597), .Z(z2[68]) );
  NANDN U891 ( .A(xregN_1), .B(zin[67]), .Z(n597) );
  NAND U892 ( .A(N72), .B(xregN_1), .Z(n596) );
  NAND U893 ( .A(n598), .B(n599), .Z(z2[67]) );
  NANDN U894 ( .A(xregN_1), .B(zin[66]), .Z(n599) );
  NAND U895 ( .A(N71), .B(xregN_1), .Z(n598) );
  NAND U896 ( .A(n600), .B(n601), .Z(z2[66]) );
  NANDN U897 ( .A(xregN_1), .B(zin[65]), .Z(n601) );
  NAND U898 ( .A(N70), .B(xregN_1), .Z(n600) );
  NAND U899 ( .A(n602), .B(n603), .Z(z2[65]) );
  NANDN U900 ( .A(xregN_1), .B(zin[64]), .Z(n603) );
  NAND U901 ( .A(N69), .B(xregN_1), .Z(n602) );
  NAND U902 ( .A(n604), .B(n605), .Z(z2[64]) );
  NANDN U903 ( .A(xregN_1), .B(zin[63]), .Z(n605) );
  NAND U904 ( .A(N68), .B(xregN_1), .Z(n604) );
  NAND U905 ( .A(n606), .B(n607), .Z(z2[63]) );
  NANDN U906 ( .A(xregN_1), .B(zin[62]), .Z(n607) );
  NAND U907 ( .A(N67), .B(xregN_1), .Z(n606) );
  NAND U908 ( .A(n608), .B(n609), .Z(z2[62]) );
  NANDN U909 ( .A(xregN_1), .B(zin[61]), .Z(n609) );
  NAND U910 ( .A(N66), .B(xregN_1), .Z(n608) );
  NAND U911 ( .A(n610), .B(n611), .Z(z2[61]) );
  NANDN U912 ( .A(xregN_1), .B(zin[60]), .Z(n611) );
  NAND U913 ( .A(N65), .B(xregN_1), .Z(n610) );
  NAND U914 ( .A(n612), .B(n613), .Z(z2[60]) );
  NANDN U915 ( .A(xregN_1), .B(zin[59]), .Z(n613) );
  NAND U916 ( .A(N64), .B(xregN_1), .Z(n612) );
  NAND U917 ( .A(n614), .B(n615), .Z(z2[5]) );
  NANDN U918 ( .A(xregN_1), .B(zin[4]), .Z(n615) );
  NAND U919 ( .A(N9), .B(xregN_1), .Z(n614) );
  NAND U920 ( .A(n616), .B(n617), .Z(z2[59]) );
  NANDN U921 ( .A(xregN_1), .B(zin[58]), .Z(n617) );
  NAND U922 ( .A(N63), .B(xregN_1), .Z(n616) );
  NAND U923 ( .A(n618), .B(n619), .Z(z2[58]) );
  NANDN U924 ( .A(xregN_1), .B(zin[57]), .Z(n619) );
  NAND U925 ( .A(N62), .B(xregN_1), .Z(n618) );
  NAND U926 ( .A(n620), .B(n621), .Z(z2[57]) );
  NANDN U927 ( .A(xregN_1), .B(zin[56]), .Z(n621) );
  NAND U928 ( .A(N61), .B(xregN_1), .Z(n620) );
  NAND U929 ( .A(n622), .B(n623), .Z(z2[56]) );
  NANDN U930 ( .A(xregN_1), .B(zin[55]), .Z(n623) );
  NAND U931 ( .A(N60), .B(xregN_1), .Z(n622) );
  NAND U932 ( .A(n624), .B(n625), .Z(z2[55]) );
  NANDN U933 ( .A(xregN_1), .B(zin[54]), .Z(n625) );
  NAND U934 ( .A(N59), .B(xregN_1), .Z(n624) );
  NAND U935 ( .A(n626), .B(n627), .Z(z2[54]) );
  NANDN U936 ( .A(xregN_1), .B(zin[53]), .Z(n627) );
  NAND U937 ( .A(N58), .B(xregN_1), .Z(n626) );
  NAND U938 ( .A(n628), .B(n629), .Z(z2[53]) );
  NANDN U939 ( .A(xregN_1), .B(zin[52]), .Z(n629) );
  NAND U940 ( .A(N57), .B(xregN_1), .Z(n628) );
  NAND U941 ( .A(n630), .B(n631), .Z(z2[52]) );
  NANDN U942 ( .A(xregN_1), .B(zin[51]), .Z(n631) );
  NAND U943 ( .A(N56), .B(xregN_1), .Z(n630) );
  NAND U944 ( .A(n632), .B(n633), .Z(z2[51]) );
  NANDN U945 ( .A(xregN_1), .B(zin[50]), .Z(n633) );
  NAND U946 ( .A(N55), .B(xregN_1), .Z(n632) );
  NAND U947 ( .A(n634), .B(n635), .Z(z2[50]) );
  NANDN U948 ( .A(xregN_1), .B(zin[49]), .Z(n635) );
  NAND U949 ( .A(N54), .B(xregN_1), .Z(n634) );
  NAND U950 ( .A(n636), .B(n637), .Z(z2[4]) );
  NANDN U951 ( .A(xregN_1), .B(zin[3]), .Z(n637) );
  NAND U952 ( .A(N8), .B(xregN_1), .Z(n636) );
  NAND U953 ( .A(n638), .B(n639), .Z(z2[49]) );
  NANDN U954 ( .A(xregN_1), .B(zin[48]), .Z(n639) );
  NAND U955 ( .A(N53), .B(xregN_1), .Z(n638) );
  NAND U956 ( .A(n640), .B(n641), .Z(z2[48]) );
  NANDN U957 ( .A(xregN_1), .B(zin[47]), .Z(n641) );
  NAND U958 ( .A(N52), .B(xregN_1), .Z(n640) );
  NAND U959 ( .A(n642), .B(n643), .Z(z2[47]) );
  NANDN U960 ( .A(xregN_1), .B(zin[46]), .Z(n643) );
  NAND U961 ( .A(N51), .B(xregN_1), .Z(n642) );
  NAND U962 ( .A(n644), .B(n645), .Z(z2[46]) );
  NANDN U963 ( .A(xregN_1), .B(zin[45]), .Z(n645) );
  NAND U964 ( .A(N50), .B(xregN_1), .Z(n644) );
  NAND U965 ( .A(n646), .B(n647), .Z(z2[45]) );
  NANDN U966 ( .A(xregN_1), .B(zin[44]), .Z(n647) );
  NAND U967 ( .A(N49), .B(xregN_1), .Z(n646) );
  NAND U968 ( .A(n648), .B(n649), .Z(z2[44]) );
  NANDN U969 ( .A(xregN_1), .B(zin[43]), .Z(n649) );
  NAND U970 ( .A(N48), .B(xregN_1), .Z(n648) );
  NAND U971 ( .A(n650), .B(n651), .Z(z2[43]) );
  NANDN U972 ( .A(xregN_1), .B(zin[42]), .Z(n651) );
  NAND U973 ( .A(N47), .B(xregN_1), .Z(n650) );
  NAND U974 ( .A(n652), .B(n653), .Z(z2[42]) );
  NANDN U975 ( .A(xregN_1), .B(zin[41]), .Z(n653) );
  NAND U976 ( .A(N46), .B(xregN_1), .Z(n652) );
  NAND U977 ( .A(n654), .B(n655), .Z(z2[41]) );
  NANDN U978 ( .A(xregN_1), .B(zin[40]), .Z(n655) );
  NAND U979 ( .A(N45), .B(xregN_1), .Z(n654) );
  NAND U980 ( .A(n656), .B(n657), .Z(z2[40]) );
  NANDN U981 ( .A(xregN_1), .B(zin[39]), .Z(n657) );
  NAND U982 ( .A(N44), .B(xregN_1), .Z(n656) );
  NAND U983 ( .A(n658), .B(n659), .Z(z2[3]) );
  NANDN U984 ( .A(xregN_1), .B(zin[2]), .Z(n659) );
  NAND U985 ( .A(N7), .B(xregN_1), .Z(n658) );
  NAND U986 ( .A(n660), .B(n661), .Z(z2[39]) );
  NANDN U987 ( .A(xregN_1), .B(zin[38]), .Z(n661) );
  NAND U988 ( .A(N43), .B(xregN_1), .Z(n660) );
  NAND U989 ( .A(n662), .B(n663), .Z(z2[38]) );
  NANDN U990 ( .A(xregN_1), .B(zin[37]), .Z(n663) );
  NAND U991 ( .A(N42), .B(xregN_1), .Z(n662) );
  NAND U992 ( .A(n664), .B(n665), .Z(z2[37]) );
  NANDN U993 ( .A(xregN_1), .B(zin[36]), .Z(n665) );
  NAND U994 ( .A(N41), .B(xregN_1), .Z(n664) );
  NAND U995 ( .A(n666), .B(n667), .Z(z2[36]) );
  NANDN U996 ( .A(xregN_1), .B(zin[35]), .Z(n667) );
  NAND U997 ( .A(N40), .B(xregN_1), .Z(n666) );
  NAND U998 ( .A(n668), .B(n669), .Z(z2[35]) );
  NANDN U999 ( .A(xregN_1), .B(zin[34]), .Z(n669) );
  NAND U1000 ( .A(N39), .B(xregN_1), .Z(n668) );
  NAND U1001 ( .A(n670), .B(n671), .Z(z2[34]) );
  NANDN U1002 ( .A(xregN_1), .B(zin[33]), .Z(n671) );
  NAND U1003 ( .A(N38), .B(xregN_1), .Z(n670) );
  NAND U1004 ( .A(n672), .B(n673), .Z(z2[33]) );
  NANDN U1005 ( .A(xregN_1), .B(zin[32]), .Z(n673) );
  NAND U1006 ( .A(N37), .B(xregN_1), .Z(n672) );
  NAND U1007 ( .A(n674), .B(n675), .Z(z2[32]) );
  NANDN U1008 ( .A(xregN_1), .B(zin[31]), .Z(n675) );
  NAND U1009 ( .A(N36), .B(xregN_1), .Z(n674) );
  NAND U1010 ( .A(n676), .B(n677), .Z(z2[31]) );
  NANDN U1011 ( .A(xregN_1), .B(zin[30]), .Z(n677) );
  NAND U1012 ( .A(N35), .B(xregN_1), .Z(n676) );
  NAND U1013 ( .A(n678), .B(n679), .Z(z2[30]) );
  NANDN U1014 ( .A(xregN_1), .B(zin[29]), .Z(n679) );
  NAND U1015 ( .A(N34), .B(xregN_1), .Z(n678) );
  NAND U1016 ( .A(n680), .B(n681), .Z(z2[2]) );
  NANDN U1017 ( .A(xregN_1), .B(zin[1]), .Z(n681) );
  NAND U1018 ( .A(N6), .B(xregN_1), .Z(n680) );
  NAND U1019 ( .A(n682), .B(n683), .Z(z2[29]) );
  NANDN U1020 ( .A(xregN_1), .B(zin[28]), .Z(n683) );
  NAND U1021 ( .A(N33), .B(xregN_1), .Z(n682) );
  NAND U1022 ( .A(n684), .B(n685), .Z(z2[28]) );
  NANDN U1023 ( .A(xregN_1), .B(zin[27]), .Z(n685) );
  NAND U1024 ( .A(N32), .B(xregN_1), .Z(n684) );
  NAND U1025 ( .A(n686), .B(n687), .Z(z2[27]) );
  NANDN U1026 ( .A(xregN_1), .B(zin[26]), .Z(n687) );
  NAND U1027 ( .A(N31), .B(xregN_1), .Z(n686) );
  NAND U1028 ( .A(n688), .B(n689), .Z(z2[26]) );
  NANDN U1029 ( .A(xregN_1), .B(zin[25]), .Z(n689) );
  NAND U1030 ( .A(N30), .B(xregN_1), .Z(n688) );
  NAND U1031 ( .A(n690), .B(n691), .Z(z2[25]) );
  NANDN U1032 ( .A(xregN_1), .B(zin[24]), .Z(n691) );
  NAND U1033 ( .A(N29), .B(xregN_1), .Z(n690) );
  NAND U1034 ( .A(n692), .B(n693), .Z(z2[257]) );
  NANDN U1035 ( .A(xregN_1), .B(zin[256]), .Z(n693) );
  NAND U1036 ( .A(N261), .B(xregN_1), .Z(n692) );
  NAND U1037 ( .A(n694), .B(n695), .Z(z2[256]) );
  NANDN U1038 ( .A(xregN_1), .B(zin[255]), .Z(n695) );
  NAND U1039 ( .A(N260), .B(xregN_1), .Z(n694) );
  NAND U1040 ( .A(n696), .B(n697), .Z(z2[255]) );
  NANDN U1041 ( .A(xregN_1), .B(zin[254]), .Z(n697) );
  NAND U1042 ( .A(N259), .B(xregN_1), .Z(n696) );
  NAND U1043 ( .A(n698), .B(n699), .Z(z2[254]) );
  NANDN U1044 ( .A(xregN_1), .B(zin[253]), .Z(n699) );
  NAND U1045 ( .A(N258), .B(xregN_1), .Z(n698) );
  NAND U1046 ( .A(n700), .B(n701), .Z(z2[253]) );
  NANDN U1047 ( .A(xregN_1), .B(zin[252]), .Z(n701) );
  NAND U1048 ( .A(N257), .B(xregN_1), .Z(n700) );
  NAND U1049 ( .A(n702), .B(n703), .Z(z2[252]) );
  NANDN U1050 ( .A(xregN_1), .B(zin[251]), .Z(n703) );
  NAND U1051 ( .A(N256), .B(xregN_1), .Z(n702) );
  NAND U1052 ( .A(n704), .B(n705), .Z(z2[251]) );
  NANDN U1053 ( .A(xregN_1), .B(zin[250]), .Z(n705) );
  NAND U1054 ( .A(N255), .B(xregN_1), .Z(n704) );
  NAND U1055 ( .A(n706), .B(n707), .Z(z2[250]) );
  NANDN U1056 ( .A(xregN_1), .B(zin[249]), .Z(n707) );
  NAND U1057 ( .A(N254), .B(xregN_1), .Z(n706) );
  NAND U1058 ( .A(n708), .B(n709), .Z(z2[24]) );
  NANDN U1059 ( .A(xregN_1), .B(zin[23]), .Z(n709) );
  NAND U1060 ( .A(N28), .B(xregN_1), .Z(n708) );
  NAND U1061 ( .A(n710), .B(n711), .Z(z2[249]) );
  NANDN U1062 ( .A(xregN_1), .B(zin[248]), .Z(n711) );
  NAND U1063 ( .A(N253), .B(xregN_1), .Z(n710) );
  NAND U1064 ( .A(n712), .B(n713), .Z(z2[248]) );
  NANDN U1065 ( .A(xregN_1), .B(zin[247]), .Z(n713) );
  NAND U1066 ( .A(N252), .B(xregN_1), .Z(n712) );
  NAND U1067 ( .A(n714), .B(n715), .Z(z2[247]) );
  NANDN U1068 ( .A(xregN_1), .B(zin[246]), .Z(n715) );
  NAND U1069 ( .A(N251), .B(xregN_1), .Z(n714) );
  NAND U1070 ( .A(n716), .B(n717), .Z(z2[246]) );
  NANDN U1071 ( .A(xregN_1), .B(zin[245]), .Z(n717) );
  NAND U1072 ( .A(N250), .B(xregN_1), .Z(n716) );
  NAND U1073 ( .A(n718), .B(n719), .Z(z2[245]) );
  NANDN U1074 ( .A(xregN_1), .B(zin[244]), .Z(n719) );
  NAND U1075 ( .A(N249), .B(xregN_1), .Z(n718) );
  NAND U1076 ( .A(n720), .B(n721), .Z(z2[244]) );
  NANDN U1077 ( .A(xregN_1), .B(zin[243]), .Z(n721) );
  NAND U1078 ( .A(N248), .B(xregN_1), .Z(n720) );
  NAND U1079 ( .A(n722), .B(n723), .Z(z2[243]) );
  NANDN U1080 ( .A(xregN_1), .B(zin[242]), .Z(n723) );
  NAND U1081 ( .A(N247), .B(xregN_1), .Z(n722) );
  NAND U1082 ( .A(n724), .B(n725), .Z(z2[242]) );
  NANDN U1083 ( .A(xregN_1), .B(zin[241]), .Z(n725) );
  NAND U1084 ( .A(N246), .B(xregN_1), .Z(n724) );
  NAND U1085 ( .A(n726), .B(n727), .Z(z2[241]) );
  NANDN U1086 ( .A(xregN_1), .B(zin[240]), .Z(n727) );
  NAND U1087 ( .A(N245), .B(xregN_1), .Z(n726) );
  NAND U1088 ( .A(n728), .B(n729), .Z(z2[240]) );
  NANDN U1089 ( .A(xregN_1), .B(zin[239]), .Z(n729) );
  NAND U1090 ( .A(N244), .B(xregN_1), .Z(n728) );
  NAND U1091 ( .A(n730), .B(n731), .Z(z2[23]) );
  NANDN U1092 ( .A(xregN_1), .B(zin[22]), .Z(n731) );
  NAND U1093 ( .A(N27), .B(xregN_1), .Z(n730) );
  NAND U1094 ( .A(n732), .B(n733), .Z(z2[239]) );
  NANDN U1095 ( .A(xregN_1), .B(zin[238]), .Z(n733) );
  NAND U1096 ( .A(N243), .B(xregN_1), .Z(n732) );
  NAND U1097 ( .A(n734), .B(n735), .Z(z2[238]) );
  NANDN U1098 ( .A(xregN_1), .B(zin[237]), .Z(n735) );
  NAND U1099 ( .A(N242), .B(xregN_1), .Z(n734) );
  NAND U1100 ( .A(n736), .B(n737), .Z(z2[237]) );
  NANDN U1101 ( .A(xregN_1), .B(zin[236]), .Z(n737) );
  NAND U1102 ( .A(N241), .B(xregN_1), .Z(n736) );
  NAND U1103 ( .A(n738), .B(n739), .Z(z2[236]) );
  NANDN U1104 ( .A(xregN_1), .B(zin[235]), .Z(n739) );
  NAND U1105 ( .A(N240), .B(xregN_1), .Z(n738) );
  NAND U1106 ( .A(n740), .B(n741), .Z(z2[235]) );
  NANDN U1107 ( .A(xregN_1), .B(zin[234]), .Z(n741) );
  NAND U1108 ( .A(N239), .B(xregN_1), .Z(n740) );
  NAND U1109 ( .A(n742), .B(n743), .Z(z2[234]) );
  NANDN U1110 ( .A(xregN_1), .B(zin[233]), .Z(n743) );
  NAND U1111 ( .A(N238), .B(xregN_1), .Z(n742) );
  NAND U1112 ( .A(n744), .B(n745), .Z(z2[233]) );
  NANDN U1113 ( .A(xregN_1), .B(zin[232]), .Z(n745) );
  NAND U1114 ( .A(N237), .B(xregN_1), .Z(n744) );
  NAND U1115 ( .A(n746), .B(n747), .Z(z2[232]) );
  NANDN U1116 ( .A(xregN_1), .B(zin[231]), .Z(n747) );
  NAND U1117 ( .A(N236), .B(xregN_1), .Z(n746) );
  NAND U1118 ( .A(n748), .B(n749), .Z(z2[231]) );
  NANDN U1119 ( .A(xregN_1), .B(zin[230]), .Z(n749) );
  NAND U1120 ( .A(N235), .B(xregN_1), .Z(n748) );
  NAND U1121 ( .A(n750), .B(n751), .Z(z2[230]) );
  NANDN U1122 ( .A(xregN_1), .B(zin[229]), .Z(n751) );
  NAND U1123 ( .A(N234), .B(xregN_1), .Z(n750) );
  NAND U1124 ( .A(n752), .B(n753), .Z(z2[22]) );
  NANDN U1125 ( .A(xregN_1), .B(zin[21]), .Z(n753) );
  NAND U1126 ( .A(N26), .B(xregN_1), .Z(n752) );
  NAND U1127 ( .A(n754), .B(n755), .Z(z2[229]) );
  NANDN U1128 ( .A(xregN_1), .B(zin[228]), .Z(n755) );
  NAND U1129 ( .A(N233), .B(xregN_1), .Z(n754) );
  NAND U1130 ( .A(n756), .B(n757), .Z(z2[228]) );
  NANDN U1131 ( .A(xregN_1), .B(zin[227]), .Z(n757) );
  NAND U1132 ( .A(N232), .B(xregN_1), .Z(n756) );
  NAND U1133 ( .A(n758), .B(n759), .Z(z2[227]) );
  NANDN U1134 ( .A(xregN_1), .B(zin[226]), .Z(n759) );
  NAND U1135 ( .A(N231), .B(xregN_1), .Z(n758) );
  NAND U1136 ( .A(n760), .B(n761), .Z(z2[226]) );
  NANDN U1137 ( .A(xregN_1), .B(zin[225]), .Z(n761) );
  NAND U1138 ( .A(N230), .B(xregN_1), .Z(n760) );
  NAND U1139 ( .A(n762), .B(n763), .Z(z2[225]) );
  NANDN U1140 ( .A(xregN_1), .B(zin[224]), .Z(n763) );
  NAND U1141 ( .A(N229), .B(xregN_1), .Z(n762) );
  NAND U1142 ( .A(n764), .B(n765), .Z(z2[224]) );
  NANDN U1143 ( .A(xregN_1), .B(zin[223]), .Z(n765) );
  NAND U1144 ( .A(N228), .B(xregN_1), .Z(n764) );
  NAND U1145 ( .A(n766), .B(n767), .Z(z2[223]) );
  NANDN U1146 ( .A(xregN_1), .B(zin[222]), .Z(n767) );
  NAND U1147 ( .A(N227), .B(xregN_1), .Z(n766) );
  NAND U1148 ( .A(n768), .B(n769), .Z(z2[222]) );
  NANDN U1149 ( .A(xregN_1), .B(zin[221]), .Z(n769) );
  NAND U1150 ( .A(N226), .B(xregN_1), .Z(n768) );
  NAND U1151 ( .A(n770), .B(n771), .Z(z2[221]) );
  NANDN U1152 ( .A(xregN_1), .B(zin[220]), .Z(n771) );
  NAND U1153 ( .A(N225), .B(xregN_1), .Z(n770) );
  NAND U1154 ( .A(n772), .B(n773), .Z(z2[220]) );
  NANDN U1155 ( .A(xregN_1), .B(zin[219]), .Z(n773) );
  NAND U1156 ( .A(N224), .B(xregN_1), .Z(n772) );
  NAND U1157 ( .A(n774), .B(n775), .Z(z2[21]) );
  NANDN U1158 ( .A(xregN_1), .B(zin[20]), .Z(n775) );
  NAND U1159 ( .A(N25), .B(xregN_1), .Z(n774) );
  NAND U1160 ( .A(n776), .B(n777), .Z(z2[219]) );
  NANDN U1161 ( .A(xregN_1), .B(zin[218]), .Z(n777) );
  NAND U1162 ( .A(N223), .B(xregN_1), .Z(n776) );
  NAND U1163 ( .A(n778), .B(n779), .Z(z2[218]) );
  NANDN U1164 ( .A(xregN_1), .B(zin[217]), .Z(n779) );
  NAND U1165 ( .A(N222), .B(xregN_1), .Z(n778) );
  NAND U1166 ( .A(n780), .B(n781), .Z(z2[217]) );
  NANDN U1167 ( .A(xregN_1), .B(zin[216]), .Z(n781) );
  NAND U1168 ( .A(N221), .B(xregN_1), .Z(n780) );
  NAND U1169 ( .A(n782), .B(n783), .Z(z2[216]) );
  NANDN U1170 ( .A(xregN_1), .B(zin[215]), .Z(n783) );
  NAND U1171 ( .A(N220), .B(xregN_1), .Z(n782) );
  NAND U1172 ( .A(n784), .B(n785), .Z(z2[215]) );
  NANDN U1173 ( .A(xregN_1), .B(zin[214]), .Z(n785) );
  NAND U1174 ( .A(N219), .B(xregN_1), .Z(n784) );
  NAND U1175 ( .A(n786), .B(n787), .Z(z2[214]) );
  NANDN U1176 ( .A(xregN_1), .B(zin[213]), .Z(n787) );
  NAND U1177 ( .A(N218), .B(xregN_1), .Z(n786) );
  NAND U1178 ( .A(n788), .B(n789), .Z(z2[213]) );
  NANDN U1179 ( .A(xregN_1), .B(zin[212]), .Z(n789) );
  NAND U1180 ( .A(N217), .B(xregN_1), .Z(n788) );
  NAND U1181 ( .A(n790), .B(n791), .Z(z2[212]) );
  NANDN U1182 ( .A(xregN_1), .B(zin[211]), .Z(n791) );
  NAND U1183 ( .A(N216), .B(xregN_1), .Z(n790) );
  NAND U1184 ( .A(n792), .B(n793), .Z(z2[211]) );
  NANDN U1185 ( .A(xregN_1), .B(zin[210]), .Z(n793) );
  NAND U1186 ( .A(N215), .B(xregN_1), .Z(n792) );
  NAND U1187 ( .A(n794), .B(n795), .Z(z2[210]) );
  NANDN U1188 ( .A(xregN_1), .B(zin[209]), .Z(n795) );
  NAND U1189 ( .A(N214), .B(xregN_1), .Z(n794) );
  NAND U1190 ( .A(n796), .B(n797), .Z(z2[20]) );
  NANDN U1191 ( .A(xregN_1), .B(zin[19]), .Z(n797) );
  NAND U1192 ( .A(N24), .B(xregN_1), .Z(n796) );
  NAND U1193 ( .A(n798), .B(n799), .Z(z2[209]) );
  NANDN U1194 ( .A(xregN_1), .B(zin[208]), .Z(n799) );
  NAND U1195 ( .A(N213), .B(xregN_1), .Z(n798) );
  NAND U1196 ( .A(n800), .B(n801), .Z(z2[208]) );
  NANDN U1197 ( .A(xregN_1), .B(zin[207]), .Z(n801) );
  NAND U1198 ( .A(N212), .B(xregN_1), .Z(n800) );
  NAND U1199 ( .A(n802), .B(n803), .Z(z2[207]) );
  NANDN U1200 ( .A(xregN_1), .B(zin[206]), .Z(n803) );
  NAND U1201 ( .A(N211), .B(xregN_1), .Z(n802) );
  NAND U1202 ( .A(n804), .B(n805), .Z(z2[206]) );
  NANDN U1203 ( .A(xregN_1), .B(zin[205]), .Z(n805) );
  NAND U1204 ( .A(N210), .B(xregN_1), .Z(n804) );
  NAND U1205 ( .A(n806), .B(n807), .Z(z2[205]) );
  NANDN U1206 ( .A(xregN_1), .B(zin[204]), .Z(n807) );
  NAND U1207 ( .A(N209), .B(xregN_1), .Z(n806) );
  NAND U1208 ( .A(n808), .B(n809), .Z(z2[204]) );
  NANDN U1209 ( .A(xregN_1), .B(zin[203]), .Z(n809) );
  NAND U1210 ( .A(N208), .B(xregN_1), .Z(n808) );
  NAND U1211 ( .A(n810), .B(n811), .Z(z2[203]) );
  NANDN U1212 ( .A(xregN_1), .B(zin[202]), .Z(n811) );
  NAND U1213 ( .A(N207), .B(xregN_1), .Z(n810) );
  NAND U1214 ( .A(n812), .B(n813), .Z(z2[202]) );
  NANDN U1215 ( .A(xregN_1), .B(zin[201]), .Z(n813) );
  NAND U1216 ( .A(N206), .B(xregN_1), .Z(n812) );
  NAND U1217 ( .A(n814), .B(n815), .Z(z2[201]) );
  NANDN U1218 ( .A(xregN_1), .B(zin[200]), .Z(n815) );
  NAND U1219 ( .A(N205), .B(xregN_1), .Z(n814) );
  NAND U1220 ( .A(n816), .B(n817), .Z(z2[200]) );
  NANDN U1221 ( .A(xregN_1), .B(zin[199]), .Z(n817) );
  NAND U1222 ( .A(N204), .B(xregN_1), .Z(n816) );
  NAND U1223 ( .A(n818), .B(n819), .Z(z2[1]) );
  NANDN U1224 ( .A(xregN_1), .B(zin[0]), .Z(n819) );
  NAND U1225 ( .A(N5), .B(xregN_1), .Z(n818) );
  NAND U1226 ( .A(n820), .B(n821), .Z(z2[19]) );
  NANDN U1227 ( .A(xregN_1), .B(zin[18]), .Z(n821) );
  NAND U1228 ( .A(N23), .B(xregN_1), .Z(n820) );
  NAND U1229 ( .A(n822), .B(n823), .Z(z2[199]) );
  NANDN U1230 ( .A(xregN_1), .B(zin[198]), .Z(n823) );
  NAND U1231 ( .A(N203), .B(xregN_1), .Z(n822) );
  NAND U1232 ( .A(n824), .B(n825), .Z(z2[198]) );
  NANDN U1233 ( .A(xregN_1), .B(zin[197]), .Z(n825) );
  NAND U1234 ( .A(N202), .B(xregN_1), .Z(n824) );
  NAND U1235 ( .A(n826), .B(n827), .Z(z2[197]) );
  NANDN U1236 ( .A(xregN_1), .B(zin[196]), .Z(n827) );
  NAND U1237 ( .A(N201), .B(xregN_1), .Z(n826) );
  NAND U1238 ( .A(n828), .B(n829), .Z(z2[196]) );
  NANDN U1239 ( .A(xregN_1), .B(zin[195]), .Z(n829) );
  NAND U1240 ( .A(N200), .B(xregN_1), .Z(n828) );
  NAND U1241 ( .A(n830), .B(n831), .Z(z2[195]) );
  NANDN U1242 ( .A(xregN_1), .B(zin[194]), .Z(n831) );
  NAND U1243 ( .A(N199), .B(xregN_1), .Z(n830) );
  NAND U1244 ( .A(n832), .B(n833), .Z(z2[194]) );
  NANDN U1245 ( .A(xregN_1), .B(zin[193]), .Z(n833) );
  NAND U1246 ( .A(N198), .B(xregN_1), .Z(n832) );
  NAND U1247 ( .A(n834), .B(n835), .Z(z2[193]) );
  NANDN U1248 ( .A(xregN_1), .B(zin[192]), .Z(n835) );
  NAND U1249 ( .A(N197), .B(xregN_1), .Z(n834) );
  NAND U1250 ( .A(n836), .B(n837), .Z(z2[192]) );
  NANDN U1251 ( .A(xregN_1), .B(zin[191]), .Z(n837) );
  NAND U1252 ( .A(N196), .B(xregN_1), .Z(n836) );
  NAND U1253 ( .A(n838), .B(n839), .Z(z2[191]) );
  NANDN U1254 ( .A(xregN_1), .B(zin[190]), .Z(n839) );
  NAND U1255 ( .A(N195), .B(xregN_1), .Z(n838) );
  NAND U1256 ( .A(n840), .B(n841), .Z(z2[190]) );
  NANDN U1257 ( .A(xregN_1), .B(zin[189]), .Z(n841) );
  NAND U1258 ( .A(N194), .B(xregN_1), .Z(n840) );
  NAND U1259 ( .A(n842), .B(n843), .Z(z2[18]) );
  NANDN U1260 ( .A(xregN_1), .B(zin[17]), .Z(n843) );
  NAND U1261 ( .A(N22), .B(xregN_1), .Z(n842) );
  NAND U1262 ( .A(n844), .B(n845), .Z(z2[189]) );
  NANDN U1263 ( .A(xregN_1), .B(zin[188]), .Z(n845) );
  NAND U1264 ( .A(N193), .B(xregN_1), .Z(n844) );
  NAND U1265 ( .A(n846), .B(n847), .Z(z2[188]) );
  NANDN U1266 ( .A(xregN_1), .B(zin[187]), .Z(n847) );
  NAND U1267 ( .A(N192), .B(xregN_1), .Z(n846) );
  NAND U1268 ( .A(n848), .B(n849), .Z(z2[187]) );
  NANDN U1269 ( .A(xregN_1), .B(zin[186]), .Z(n849) );
  NAND U1270 ( .A(N191), .B(xregN_1), .Z(n848) );
  NAND U1271 ( .A(n850), .B(n851), .Z(z2[186]) );
  NANDN U1272 ( .A(xregN_1), .B(zin[185]), .Z(n851) );
  NAND U1273 ( .A(N190), .B(xregN_1), .Z(n850) );
  NAND U1274 ( .A(n852), .B(n853), .Z(z2[185]) );
  NANDN U1275 ( .A(xregN_1), .B(zin[184]), .Z(n853) );
  NAND U1276 ( .A(N189), .B(xregN_1), .Z(n852) );
  NAND U1277 ( .A(n854), .B(n855), .Z(z2[184]) );
  NANDN U1278 ( .A(xregN_1), .B(zin[183]), .Z(n855) );
  NAND U1279 ( .A(N188), .B(xregN_1), .Z(n854) );
  NAND U1280 ( .A(n856), .B(n857), .Z(z2[183]) );
  NANDN U1281 ( .A(xregN_1), .B(zin[182]), .Z(n857) );
  NAND U1282 ( .A(N187), .B(xregN_1), .Z(n856) );
  NAND U1283 ( .A(n858), .B(n859), .Z(z2[182]) );
  NANDN U1284 ( .A(xregN_1), .B(zin[181]), .Z(n859) );
  NAND U1285 ( .A(N186), .B(xregN_1), .Z(n858) );
  NAND U1286 ( .A(n860), .B(n861), .Z(z2[181]) );
  NANDN U1287 ( .A(xregN_1), .B(zin[180]), .Z(n861) );
  NAND U1288 ( .A(N185), .B(xregN_1), .Z(n860) );
  NAND U1289 ( .A(n862), .B(n863), .Z(z2[180]) );
  NANDN U1290 ( .A(xregN_1), .B(zin[179]), .Z(n863) );
  NAND U1291 ( .A(N184), .B(xregN_1), .Z(n862) );
  NAND U1292 ( .A(n864), .B(n865), .Z(z2[17]) );
  NANDN U1293 ( .A(xregN_1), .B(zin[16]), .Z(n865) );
  NAND U1294 ( .A(N21), .B(xregN_1), .Z(n864) );
  NAND U1295 ( .A(n866), .B(n867), .Z(z2[179]) );
  NANDN U1296 ( .A(xregN_1), .B(zin[178]), .Z(n867) );
  NAND U1297 ( .A(N183), .B(xregN_1), .Z(n866) );
  NAND U1298 ( .A(n868), .B(n869), .Z(z2[178]) );
  NANDN U1299 ( .A(xregN_1), .B(zin[177]), .Z(n869) );
  NAND U1300 ( .A(N182), .B(xregN_1), .Z(n868) );
  NAND U1301 ( .A(n870), .B(n871), .Z(z2[177]) );
  NANDN U1302 ( .A(xregN_1), .B(zin[176]), .Z(n871) );
  NAND U1303 ( .A(N181), .B(xregN_1), .Z(n870) );
  NAND U1304 ( .A(n872), .B(n873), .Z(z2[176]) );
  NANDN U1305 ( .A(xregN_1), .B(zin[175]), .Z(n873) );
  NAND U1306 ( .A(N180), .B(xregN_1), .Z(n872) );
  NAND U1307 ( .A(n874), .B(n875), .Z(z2[175]) );
  NANDN U1308 ( .A(xregN_1), .B(zin[174]), .Z(n875) );
  NAND U1309 ( .A(N179), .B(xregN_1), .Z(n874) );
  NAND U1310 ( .A(n876), .B(n877), .Z(z2[174]) );
  NANDN U1311 ( .A(xregN_1), .B(zin[173]), .Z(n877) );
  NAND U1312 ( .A(N178), .B(xregN_1), .Z(n876) );
  NAND U1313 ( .A(n878), .B(n879), .Z(z2[173]) );
  NANDN U1314 ( .A(xregN_1), .B(zin[172]), .Z(n879) );
  NAND U1315 ( .A(N177), .B(xregN_1), .Z(n878) );
  NAND U1316 ( .A(n880), .B(n881), .Z(z2[172]) );
  NANDN U1317 ( .A(xregN_1), .B(zin[171]), .Z(n881) );
  NAND U1318 ( .A(N176), .B(xregN_1), .Z(n880) );
  NAND U1319 ( .A(n882), .B(n883), .Z(z2[171]) );
  NANDN U1320 ( .A(xregN_1), .B(zin[170]), .Z(n883) );
  NAND U1321 ( .A(N175), .B(xregN_1), .Z(n882) );
  NAND U1322 ( .A(n884), .B(n885), .Z(z2[170]) );
  NANDN U1323 ( .A(xregN_1), .B(zin[169]), .Z(n885) );
  NAND U1324 ( .A(N174), .B(xregN_1), .Z(n884) );
  NAND U1325 ( .A(n886), .B(n887), .Z(z2[16]) );
  NANDN U1326 ( .A(xregN_1), .B(zin[15]), .Z(n887) );
  NAND U1327 ( .A(N20), .B(xregN_1), .Z(n886) );
  NAND U1328 ( .A(n888), .B(n889), .Z(z2[169]) );
  NANDN U1329 ( .A(xregN_1), .B(zin[168]), .Z(n889) );
  NAND U1330 ( .A(N173), .B(xregN_1), .Z(n888) );
  NAND U1331 ( .A(n890), .B(n891), .Z(z2[168]) );
  NANDN U1332 ( .A(xregN_1), .B(zin[167]), .Z(n891) );
  NAND U1333 ( .A(N172), .B(xregN_1), .Z(n890) );
  NAND U1334 ( .A(n892), .B(n893), .Z(z2[167]) );
  NANDN U1335 ( .A(xregN_1), .B(zin[166]), .Z(n893) );
  NAND U1336 ( .A(N171), .B(xregN_1), .Z(n892) );
  NAND U1337 ( .A(n894), .B(n895), .Z(z2[166]) );
  NANDN U1338 ( .A(xregN_1), .B(zin[165]), .Z(n895) );
  NAND U1339 ( .A(N170), .B(xregN_1), .Z(n894) );
  NAND U1340 ( .A(n896), .B(n897), .Z(z2[165]) );
  NANDN U1341 ( .A(xregN_1), .B(zin[164]), .Z(n897) );
  NAND U1342 ( .A(N169), .B(xregN_1), .Z(n896) );
  NAND U1343 ( .A(n898), .B(n899), .Z(z2[164]) );
  NANDN U1344 ( .A(xregN_1), .B(zin[163]), .Z(n899) );
  NAND U1345 ( .A(N168), .B(xregN_1), .Z(n898) );
  NAND U1346 ( .A(n900), .B(n901), .Z(z2[163]) );
  NANDN U1347 ( .A(xregN_1), .B(zin[162]), .Z(n901) );
  NAND U1348 ( .A(N167), .B(xregN_1), .Z(n900) );
  NAND U1349 ( .A(n902), .B(n903), .Z(z2[162]) );
  NANDN U1350 ( .A(xregN_1), .B(zin[161]), .Z(n903) );
  NAND U1351 ( .A(N166), .B(xregN_1), .Z(n902) );
  NAND U1352 ( .A(n904), .B(n905), .Z(z2[161]) );
  NANDN U1353 ( .A(xregN_1), .B(zin[160]), .Z(n905) );
  NAND U1354 ( .A(N165), .B(xregN_1), .Z(n904) );
  NAND U1355 ( .A(n906), .B(n907), .Z(z2[160]) );
  NANDN U1356 ( .A(xregN_1), .B(zin[159]), .Z(n907) );
  NAND U1357 ( .A(N164), .B(xregN_1), .Z(n906) );
  NAND U1358 ( .A(n908), .B(n909), .Z(z2[15]) );
  NANDN U1359 ( .A(xregN_1), .B(zin[14]), .Z(n909) );
  NAND U1360 ( .A(N19), .B(xregN_1), .Z(n908) );
  NAND U1361 ( .A(n910), .B(n911), .Z(z2[159]) );
  NANDN U1362 ( .A(xregN_1), .B(zin[158]), .Z(n911) );
  NAND U1363 ( .A(N163), .B(xregN_1), .Z(n910) );
  NAND U1364 ( .A(n912), .B(n913), .Z(z2[158]) );
  NANDN U1365 ( .A(xregN_1), .B(zin[157]), .Z(n913) );
  NAND U1366 ( .A(N162), .B(xregN_1), .Z(n912) );
  NAND U1367 ( .A(n914), .B(n915), .Z(z2[157]) );
  NANDN U1368 ( .A(xregN_1), .B(zin[156]), .Z(n915) );
  NAND U1369 ( .A(N161), .B(xregN_1), .Z(n914) );
  NAND U1370 ( .A(n916), .B(n917), .Z(z2[156]) );
  NANDN U1371 ( .A(xregN_1), .B(zin[155]), .Z(n917) );
  NAND U1372 ( .A(N160), .B(xregN_1), .Z(n916) );
  NAND U1373 ( .A(n918), .B(n919), .Z(z2[155]) );
  NANDN U1374 ( .A(xregN_1), .B(zin[154]), .Z(n919) );
  NAND U1375 ( .A(N159), .B(xregN_1), .Z(n918) );
  NAND U1376 ( .A(n920), .B(n921), .Z(z2[154]) );
  NANDN U1377 ( .A(xregN_1), .B(zin[153]), .Z(n921) );
  NAND U1378 ( .A(N158), .B(xregN_1), .Z(n920) );
  NAND U1379 ( .A(n922), .B(n923), .Z(z2[153]) );
  NANDN U1380 ( .A(xregN_1), .B(zin[152]), .Z(n923) );
  NAND U1381 ( .A(N157), .B(xregN_1), .Z(n922) );
  NAND U1382 ( .A(n924), .B(n925), .Z(z2[152]) );
  NANDN U1383 ( .A(xregN_1), .B(zin[151]), .Z(n925) );
  NAND U1384 ( .A(N156), .B(xregN_1), .Z(n924) );
  NAND U1385 ( .A(n926), .B(n927), .Z(z2[151]) );
  NANDN U1386 ( .A(xregN_1), .B(zin[150]), .Z(n927) );
  NAND U1387 ( .A(N155), .B(xregN_1), .Z(n926) );
  NAND U1388 ( .A(n928), .B(n929), .Z(z2[150]) );
  NANDN U1389 ( .A(xregN_1), .B(zin[149]), .Z(n929) );
  NAND U1390 ( .A(N154), .B(xregN_1), .Z(n928) );
  NAND U1391 ( .A(n930), .B(n931), .Z(z2[14]) );
  NANDN U1392 ( .A(xregN_1), .B(zin[13]), .Z(n931) );
  NAND U1393 ( .A(N18), .B(xregN_1), .Z(n930) );
  NAND U1394 ( .A(n932), .B(n933), .Z(z2[149]) );
  NANDN U1395 ( .A(xregN_1), .B(zin[148]), .Z(n933) );
  NAND U1396 ( .A(N153), .B(xregN_1), .Z(n932) );
  NAND U1397 ( .A(n934), .B(n935), .Z(z2[148]) );
  NANDN U1398 ( .A(xregN_1), .B(zin[147]), .Z(n935) );
  NAND U1399 ( .A(N152), .B(xregN_1), .Z(n934) );
  NAND U1400 ( .A(n936), .B(n937), .Z(z2[147]) );
  NANDN U1401 ( .A(xregN_1), .B(zin[146]), .Z(n937) );
  NAND U1402 ( .A(N151), .B(xregN_1), .Z(n936) );
  NAND U1403 ( .A(n938), .B(n939), .Z(z2[146]) );
  NANDN U1404 ( .A(xregN_1), .B(zin[145]), .Z(n939) );
  NAND U1405 ( .A(N150), .B(xregN_1), .Z(n938) );
  NAND U1406 ( .A(n940), .B(n941), .Z(z2[145]) );
  NANDN U1407 ( .A(xregN_1), .B(zin[144]), .Z(n941) );
  NAND U1408 ( .A(N149), .B(xregN_1), .Z(n940) );
  NAND U1409 ( .A(n942), .B(n943), .Z(z2[144]) );
  NANDN U1410 ( .A(xregN_1), .B(zin[143]), .Z(n943) );
  NAND U1411 ( .A(N148), .B(xregN_1), .Z(n942) );
  NAND U1412 ( .A(n944), .B(n945), .Z(z2[143]) );
  NANDN U1413 ( .A(xregN_1), .B(zin[142]), .Z(n945) );
  NAND U1414 ( .A(N147), .B(xregN_1), .Z(n944) );
  NAND U1415 ( .A(n946), .B(n947), .Z(z2[142]) );
  NANDN U1416 ( .A(xregN_1), .B(zin[141]), .Z(n947) );
  NAND U1417 ( .A(N146), .B(xregN_1), .Z(n946) );
  NAND U1418 ( .A(n948), .B(n949), .Z(z2[141]) );
  NANDN U1419 ( .A(xregN_1), .B(zin[140]), .Z(n949) );
  NAND U1420 ( .A(N145), .B(xregN_1), .Z(n948) );
  NAND U1421 ( .A(n950), .B(n951), .Z(z2[140]) );
  NANDN U1422 ( .A(xregN_1), .B(zin[139]), .Z(n951) );
  NAND U1423 ( .A(N144), .B(xregN_1), .Z(n950) );
  NAND U1424 ( .A(n952), .B(n953), .Z(z2[13]) );
  NANDN U1425 ( .A(xregN_1), .B(zin[12]), .Z(n953) );
  NAND U1426 ( .A(N17), .B(xregN_1), .Z(n952) );
  NAND U1427 ( .A(n954), .B(n955), .Z(z2[139]) );
  NANDN U1428 ( .A(xregN_1), .B(zin[138]), .Z(n955) );
  NAND U1429 ( .A(N143), .B(xregN_1), .Z(n954) );
  NAND U1430 ( .A(n956), .B(n957), .Z(z2[138]) );
  NANDN U1431 ( .A(xregN_1), .B(zin[137]), .Z(n957) );
  NAND U1432 ( .A(N142), .B(xregN_1), .Z(n956) );
  NAND U1433 ( .A(n958), .B(n959), .Z(z2[137]) );
  NANDN U1434 ( .A(xregN_1), .B(zin[136]), .Z(n959) );
  NAND U1435 ( .A(N141), .B(xregN_1), .Z(n958) );
  NAND U1436 ( .A(n960), .B(n961), .Z(z2[136]) );
  NANDN U1437 ( .A(xregN_1), .B(zin[135]), .Z(n961) );
  NAND U1438 ( .A(N140), .B(xregN_1), .Z(n960) );
  NAND U1439 ( .A(n962), .B(n963), .Z(z2[135]) );
  NANDN U1440 ( .A(xregN_1), .B(zin[134]), .Z(n963) );
  NAND U1441 ( .A(N139), .B(xregN_1), .Z(n962) );
  NAND U1442 ( .A(n964), .B(n965), .Z(z2[134]) );
  NANDN U1443 ( .A(xregN_1), .B(zin[133]), .Z(n965) );
  NAND U1444 ( .A(N138), .B(xregN_1), .Z(n964) );
  NAND U1445 ( .A(n966), .B(n967), .Z(z2[133]) );
  NANDN U1446 ( .A(xregN_1), .B(zin[132]), .Z(n967) );
  NAND U1447 ( .A(N137), .B(xregN_1), .Z(n966) );
  NAND U1448 ( .A(n968), .B(n969), .Z(z2[132]) );
  NANDN U1449 ( .A(xregN_1), .B(zin[131]), .Z(n969) );
  NAND U1450 ( .A(N136), .B(xregN_1), .Z(n968) );
  NAND U1451 ( .A(n970), .B(n971), .Z(z2[131]) );
  NANDN U1452 ( .A(xregN_1), .B(zin[130]), .Z(n971) );
  NAND U1453 ( .A(N135), .B(xregN_1), .Z(n970) );
  NAND U1454 ( .A(n972), .B(n973), .Z(z2[130]) );
  NANDN U1455 ( .A(xregN_1), .B(zin[129]), .Z(n973) );
  NAND U1456 ( .A(N134), .B(xregN_1), .Z(n972) );
  NAND U1457 ( .A(n974), .B(n975), .Z(z2[12]) );
  NANDN U1458 ( .A(xregN_1), .B(zin[11]), .Z(n975) );
  NAND U1459 ( .A(N16), .B(xregN_1), .Z(n974) );
  NAND U1460 ( .A(n976), .B(n977), .Z(z2[129]) );
  NANDN U1461 ( .A(xregN_1), .B(zin[128]), .Z(n977) );
  NAND U1462 ( .A(N133), .B(xregN_1), .Z(n976) );
  NAND U1463 ( .A(n978), .B(n979), .Z(z2[128]) );
  NANDN U1464 ( .A(xregN_1), .B(zin[127]), .Z(n979) );
  NAND U1465 ( .A(N132), .B(xregN_1), .Z(n978) );
  NAND U1466 ( .A(n980), .B(n981), .Z(z2[127]) );
  NANDN U1467 ( .A(xregN_1), .B(zin[126]), .Z(n981) );
  NAND U1468 ( .A(N131), .B(xregN_1), .Z(n980) );
  NAND U1469 ( .A(n982), .B(n983), .Z(z2[126]) );
  NANDN U1470 ( .A(xregN_1), .B(zin[125]), .Z(n983) );
  NAND U1471 ( .A(N130), .B(xregN_1), .Z(n982) );
  NAND U1472 ( .A(n984), .B(n985), .Z(z2[125]) );
  NANDN U1473 ( .A(xregN_1), .B(zin[124]), .Z(n985) );
  NAND U1474 ( .A(N129), .B(xregN_1), .Z(n984) );
  NAND U1475 ( .A(n986), .B(n987), .Z(z2[124]) );
  NANDN U1476 ( .A(xregN_1), .B(zin[123]), .Z(n987) );
  NAND U1477 ( .A(N128), .B(xregN_1), .Z(n986) );
  NAND U1478 ( .A(n988), .B(n989), .Z(z2[123]) );
  NANDN U1479 ( .A(xregN_1), .B(zin[122]), .Z(n989) );
  NAND U1480 ( .A(N127), .B(xregN_1), .Z(n988) );
  NAND U1481 ( .A(n990), .B(n991), .Z(z2[122]) );
  NANDN U1482 ( .A(xregN_1), .B(zin[121]), .Z(n991) );
  NAND U1483 ( .A(N126), .B(xregN_1), .Z(n990) );
  NAND U1484 ( .A(n992), .B(n993), .Z(z2[121]) );
  NANDN U1485 ( .A(xregN_1), .B(zin[120]), .Z(n993) );
  NAND U1486 ( .A(N125), .B(xregN_1), .Z(n992) );
  NAND U1487 ( .A(n994), .B(n995), .Z(z2[120]) );
  NANDN U1488 ( .A(xregN_1), .B(zin[119]), .Z(n995) );
  NAND U1489 ( .A(N124), .B(xregN_1), .Z(n994) );
  NAND U1490 ( .A(n996), .B(n997), .Z(z2[11]) );
  NANDN U1491 ( .A(xregN_1), .B(zin[10]), .Z(n997) );
  NAND U1492 ( .A(N15), .B(xregN_1), .Z(n996) );
  NAND U1493 ( .A(n998), .B(n999), .Z(z2[119]) );
  NANDN U1494 ( .A(xregN_1), .B(zin[118]), .Z(n999) );
  NAND U1495 ( .A(N123), .B(xregN_1), .Z(n998) );
  NAND U1496 ( .A(n1000), .B(n1001), .Z(z2[118]) );
  NANDN U1497 ( .A(xregN_1), .B(zin[117]), .Z(n1001) );
  NAND U1498 ( .A(N122), .B(xregN_1), .Z(n1000) );
  NAND U1499 ( .A(n1002), .B(n1003), .Z(z2[117]) );
  NANDN U1500 ( .A(xregN_1), .B(zin[116]), .Z(n1003) );
  NAND U1501 ( .A(N121), .B(xregN_1), .Z(n1002) );
  NAND U1502 ( .A(n1004), .B(n1005), .Z(z2[116]) );
  NANDN U1503 ( .A(xregN_1), .B(zin[115]), .Z(n1005) );
  NAND U1504 ( .A(N120), .B(xregN_1), .Z(n1004) );
  NAND U1505 ( .A(n1006), .B(n1007), .Z(z2[115]) );
  NANDN U1506 ( .A(xregN_1), .B(zin[114]), .Z(n1007) );
  NAND U1507 ( .A(N119), .B(xregN_1), .Z(n1006) );
  NAND U1508 ( .A(n1008), .B(n1009), .Z(z2[114]) );
  NANDN U1509 ( .A(xregN_1), .B(zin[113]), .Z(n1009) );
  NAND U1510 ( .A(N118), .B(xregN_1), .Z(n1008) );
  NAND U1511 ( .A(n1010), .B(n1011), .Z(z2[113]) );
  NANDN U1512 ( .A(xregN_1), .B(zin[112]), .Z(n1011) );
  NAND U1513 ( .A(N117), .B(xregN_1), .Z(n1010) );
  NAND U1514 ( .A(n1012), .B(n1013), .Z(z2[112]) );
  NANDN U1515 ( .A(xregN_1), .B(zin[111]), .Z(n1013) );
  NAND U1516 ( .A(N116), .B(xregN_1), .Z(n1012) );
  NAND U1517 ( .A(n1014), .B(n1015), .Z(z2[111]) );
  NANDN U1518 ( .A(xregN_1), .B(zin[110]), .Z(n1015) );
  NAND U1519 ( .A(N115), .B(xregN_1), .Z(n1014) );
  NAND U1520 ( .A(n1016), .B(n1017), .Z(z2[110]) );
  NANDN U1521 ( .A(xregN_1), .B(zin[109]), .Z(n1017) );
  NAND U1522 ( .A(N114), .B(xregN_1), .Z(n1016) );
  NAND U1523 ( .A(n1018), .B(n1019), .Z(z2[10]) );
  NANDN U1524 ( .A(xregN_1), .B(zin[9]), .Z(n1019) );
  NAND U1525 ( .A(N14), .B(xregN_1), .Z(n1018) );
  NAND U1526 ( .A(n1020), .B(n1021), .Z(z2[109]) );
  NANDN U1527 ( .A(xregN_1), .B(zin[108]), .Z(n1021) );
  NAND U1528 ( .A(N113), .B(xregN_1), .Z(n1020) );
  NAND U1529 ( .A(n1022), .B(n1023), .Z(z2[108]) );
  NANDN U1530 ( .A(xregN_1), .B(zin[107]), .Z(n1023) );
  NAND U1531 ( .A(N112), .B(xregN_1), .Z(n1022) );
  NAND U1532 ( .A(n1024), .B(n1025), .Z(z2[107]) );
  NANDN U1533 ( .A(xregN_1), .B(zin[106]), .Z(n1025) );
  NAND U1534 ( .A(N111), .B(xregN_1), .Z(n1024) );
  NAND U1535 ( .A(n1026), .B(n1027), .Z(z2[106]) );
  NANDN U1536 ( .A(xregN_1), .B(zin[105]), .Z(n1027) );
  NAND U1537 ( .A(N110), .B(xregN_1), .Z(n1026) );
  NAND U1538 ( .A(n1028), .B(n1029), .Z(z2[105]) );
  NANDN U1539 ( .A(xregN_1), .B(zin[104]), .Z(n1029) );
  NAND U1540 ( .A(N109), .B(xregN_1), .Z(n1028) );
  NAND U1541 ( .A(n1030), .B(n1031), .Z(z2[104]) );
  NANDN U1542 ( .A(xregN_1), .B(zin[103]), .Z(n1031) );
  NAND U1543 ( .A(N108), .B(xregN_1), .Z(n1030) );
  NAND U1544 ( .A(n1032), .B(n1033), .Z(z2[103]) );
  NANDN U1545 ( .A(xregN_1), .B(zin[102]), .Z(n1033) );
  NAND U1546 ( .A(N107), .B(xregN_1), .Z(n1032) );
  NAND U1547 ( .A(n1034), .B(n1035), .Z(z2[102]) );
  NANDN U1548 ( .A(xregN_1), .B(zin[101]), .Z(n1035) );
  NAND U1549 ( .A(N106), .B(xregN_1), .Z(n1034) );
  NAND U1550 ( .A(n1036), .B(n1037), .Z(z2[101]) );
  NANDN U1551 ( .A(xregN_1), .B(zin[100]), .Z(n1037) );
  NAND U1552 ( .A(N105), .B(xregN_1), .Z(n1036) );
  NAND U1553 ( .A(n1038), .B(n1039), .Z(z2[100]) );
  NANDN U1554 ( .A(xregN_1), .B(zin[99]), .Z(n1039) );
  NAND U1555 ( .A(N104), .B(xregN_1), .Z(n1038) );
  AND U1556 ( .A(N4), .B(xregN_1), .Z(z2[0]) );
endmodule


module modmult_step_N256_3_DW01_sub_0 ( A, B, CI, DIFF, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280;

  IV U1 ( .A(n1279), .Z(n1) );
  IV U2 ( .A(A[1]), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(DIFF[9]) );
  XOR U4 ( .A(B[9]), .B(A[9]), .Z(n4) );
  XNOR U5 ( .A(n5), .B(n6), .Z(DIFF[99]) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(DIFF[98]) );
  XOR U8 ( .A(B[98]), .B(A[98]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(DIFF[97]) );
  XOR U10 ( .A(B[97]), .B(A[97]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(DIFF[96]) );
  XOR U12 ( .A(B[96]), .B(A[96]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(DIFF[95]) );
  XOR U14 ( .A(B[95]), .B(A[95]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(DIFF[94]) );
  XOR U16 ( .A(B[94]), .B(A[94]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(DIFF[93]) );
  XOR U18 ( .A(B[93]), .B(A[93]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(DIFF[92]) );
  XOR U20 ( .A(B[92]), .B(A[92]), .Z(n20) );
  XOR U21 ( .A(n21), .B(n22), .Z(DIFF[91]) );
  XOR U22 ( .A(B[91]), .B(A[91]), .Z(n22) );
  XOR U23 ( .A(n23), .B(n24), .Z(DIFF[90]) );
  XOR U24 ( .A(B[90]), .B(A[90]), .Z(n24) );
  XOR U25 ( .A(n25), .B(n26), .Z(DIFF[8]) );
  XOR U26 ( .A(B[8]), .B(A[8]), .Z(n26) );
  XOR U27 ( .A(n27), .B(n28), .Z(DIFF[89]) );
  XOR U28 ( .A(B[89]), .B(A[89]), .Z(n28) );
  XOR U29 ( .A(n29), .B(n30), .Z(DIFF[88]) );
  XOR U30 ( .A(B[88]), .B(A[88]), .Z(n30) );
  XOR U31 ( .A(n31), .B(n32), .Z(DIFF[87]) );
  XOR U32 ( .A(B[87]), .B(A[87]), .Z(n32) );
  XOR U33 ( .A(n33), .B(n34), .Z(DIFF[86]) );
  XOR U34 ( .A(B[86]), .B(A[86]), .Z(n34) );
  XOR U35 ( .A(n35), .B(n36), .Z(DIFF[85]) );
  XOR U36 ( .A(B[85]), .B(A[85]), .Z(n36) );
  XOR U37 ( .A(n37), .B(n38), .Z(DIFF[84]) );
  XOR U38 ( .A(B[84]), .B(A[84]), .Z(n38) );
  XOR U39 ( .A(n39), .B(n40), .Z(DIFF[83]) );
  XOR U40 ( .A(B[83]), .B(A[83]), .Z(n40) );
  XOR U41 ( .A(n41), .B(n42), .Z(DIFF[82]) );
  XOR U42 ( .A(B[82]), .B(A[82]), .Z(n42) );
  XOR U43 ( .A(n43), .B(n44), .Z(DIFF[81]) );
  XOR U44 ( .A(B[81]), .B(A[81]), .Z(n44) );
  XOR U45 ( .A(n45), .B(n46), .Z(DIFF[80]) );
  XOR U46 ( .A(B[80]), .B(A[80]), .Z(n46) );
  XOR U47 ( .A(n47), .B(n48), .Z(DIFF[7]) );
  XOR U48 ( .A(B[7]), .B(A[7]), .Z(n48) );
  XOR U49 ( .A(n49), .B(n50), .Z(DIFF[79]) );
  XOR U50 ( .A(B[79]), .B(A[79]), .Z(n50) );
  XOR U51 ( .A(n51), .B(n52), .Z(DIFF[78]) );
  XOR U52 ( .A(B[78]), .B(A[78]), .Z(n52) );
  XOR U53 ( .A(n53), .B(n54), .Z(DIFF[77]) );
  XOR U54 ( .A(B[77]), .B(A[77]), .Z(n54) );
  XOR U55 ( .A(n55), .B(n56), .Z(DIFF[76]) );
  XOR U56 ( .A(B[76]), .B(A[76]), .Z(n56) );
  XOR U57 ( .A(n57), .B(n58), .Z(DIFF[75]) );
  XOR U58 ( .A(B[75]), .B(A[75]), .Z(n58) );
  XOR U59 ( .A(n59), .B(n60), .Z(DIFF[74]) );
  XOR U60 ( .A(B[74]), .B(A[74]), .Z(n60) );
  XOR U61 ( .A(n61), .B(n62), .Z(DIFF[73]) );
  XOR U62 ( .A(B[73]), .B(A[73]), .Z(n62) );
  XOR U63 ( .A(n63), .B(n64), .Z(DIFF[72]) );
  XOR U64 ( .A(B[72]), .B(A[72]), .Z(n64) );
  XOR U65 ( .A(n65), .B(n66), .Z(DIFF[71]) );
  XOR U66 ( .A(B[71]), .B(A[71]), .Z(n66) );
  XOR U67 ( .A(n67), .B(n68), .Z(DIFF[70]) );
  XOR U68 ( .A(B[70]), .B(A[70]), .Z(n68) );
  XOR U69 ( .A(n69), .B(n70), .Z(DIFF[6]) );
  XOR U70 ( .A(B[6]), .B(A[6]), .Z(n70) );
  XOR U71 ( .A(n71), .B(n72), .Z(DIFF[69]) );
  XOR U72 ( .A(B[69]), .B(A[69]), .Z(n72) );
  XOR U73 ( .A(n73), .B(n74), .Z(DIFF[68]) );
  XOR U74 ( .A(B[68]), .B(A[68]), .Z(n74) );
  XOR U75 ( .A(n75), .B(n76), .Z(DIFF[67]) );
  XOR U76 ( .A(B[67]), .B(A[67]), .Z(n76) );
  XOR U77 ( .A(n77), .B(n78), .Z(DIFF[66]) );
  XOR U78 ( .A(B[66]), .B(A[66]), .Z(n78) );
  XOR U79 ( .A(n79), .B(n80), .Z(DIFF[65]) );
  XOR U80 ( .A(B[65]), .B(A[65]), .Z(n80) );
  XOR U81 ( .A(n81), .B(n82), .Z(DIFF[64]) );
  XOR U82 ( .A(B[64]), .B(A[64]), .Z(n82) );
  XOR U83 ( .A(n83), .B(n84), .Z(DIFF[63]) );
  XOR U84 ( .A(B[63]), .B(A[63]), .Z(n84) );
  XOR U85 ( .A(n85), .B(n86), .Z(DIFF[62]) );
  XOR U86 ( .A(B[62]), .B(A[62]), .Z(n86) );
  XOR U87 ( .A(n87), .B(n88), .Z(DIFF[61]) );
  XOR U88 ( .A(B[61]), .B(A[61]), .Z(n88) );
  XOR U89 ( .A(n89), .B(n90), .Z(DIFF[60]) );
  XOR U90 ( .A(B[60]), .B(A[60]), .Z(n90) );
  XOR U91 ( .A(n91), .B(n92), .Z(DIFF[5]) );
  XOR U92 ( .A(B[5]), .B(A[5]), .Z(n92) );
  XOR U93 ( .A(n93), .B(n94), .Z(DIFF[59]) );
  XOR U94 ( .A(B[59]), .B(A[59]), .Z(n94) );
  XOR U95 ( .A(n95), .B(n96), .Z(DIFF[58]) );
  XOR U96 ( .A(B[58]), .B(A[58]), .Z(n96) );
  XOR U97 ( .A(n97), .B(n98), .Z(DIFF[57]) );
  XOR U98 ( .A(B[57]), .B(A[57]), .Z(n98) );
  XOR U99 ( .A(n99), .B(n100), .Z(DIFF[56]) );
  XOR U100 ( .A(B[56]), .B(A[56]), .Z(n100) );
  XOR U101 ( .A(n101), .B(n102), .Z(DIFF[55]) );
  XOR U102 ( .A(B[55]), .B(A[55]), .Z(n102) );
  XOR U103 ( .A(n103), .B(n104), .Z(DIFF[54]) );
  XOR U104 ( .A(B[54]), .B(A[54]), .Z(n104) );
  XOR U105 ( .A(n105), .B(n106), .Z(DIFF[53]) );
  XOR U106 ( .A(B[53]), .B(A[53]), .Z(n106) );
  XOR U107 ( .A(n107), .B(n108), .Z(DIFF[52]) );
  XOR U108 ( .A(B[52]), .B(A[52]), .Z(n108) );
  XOR U109 ( .A(n109), .B(n110), .Z(DIFF[51]) );
  XOR U110 ( .A(B[51]), .B(A[51]), .Z(n110) );
  XOR U111 ( .A(n111), .B(n112), .Z(DIFF[50]) );
  XOR U112 ( .A(B[50]), .B(A[50]), .Z(n112) );
  XOR U113 ( .A(n113), .B(n114), .Z(DIFF[4]) );
  XOR U114 ( .A(B[4]), .B(A[4]), .Z(n114) );
  XOR U115 ( .A(n115), .B(n116), .Z(DIFF[49]) );
  XOR U116 ( .A(B[49]), .B(A[49]), .Z(n116) );
  XOR U117 ( .A(n117), .B(n118), .Z(DIFF[48]) );
  XOR U118 ( .A(B[48]), .B(A[48]), .Z(n118) );
  XOR U119 ( .A(n119), .B(n120), .Z(DIFF[47]) );
  XOR U120 ( .A(B[47]), .B(A[47]), .Z(n120) );
  XOR U121 ( .A(n121), .B(n122), .Z(DIFF[46]) );
  XOR U122 ( .A(B[46]), .B(A[46]), .Z(n122) );
  XOR U123 ( .A(n123), .B(n124), .Z(DIFF[45]) );
  XOR U124 ( .A(B[45]), .B(A[45]), .Z(n124) );
  XOR U125 ( .A(n125), .B(n126), .Z(DIFF[44]) );
  XOR U126 ( .A(B[44]), .B(A[44]), .Z(n126) );
  XOR U127 ( .A(n127), .B(n128), .Z(DIFF[43]) );
  XOR U128 ( .A(B[43]), .B(A[43]), .Z(n128) );
  XOR U129 ( .A(n129), .B(n130), .Z(DIFF[42]) );
  XOR U130 ( .A(B[42]), .B(A[42]), .Z(n130) );
  XOR U131 ( .A(n131), .B(n132), .Z(DIFF[41]) );
  XOR U132 ( .A(B[41]), .B(A[41]), .Z(n132) );
  XOR U133 ( .A(n133), .B(n134), .Z(DIFF[40]) );
  XOR U134 ( .A(B[40]), .B(A[40]), .Z(n134) );
  XOR U135 ( .A(n135), .B(n136), .Z(DIFF[3]) );
  XOR U136 ( .A(B[3]), .B(A[3]), .Z(n136) );
  XOR U137 ( .A(n137), .B(n138), .Z(DIFF[39]) );
  XOR U138 ( .A(B[39]), .B(A[39]), .Z(n138) );
  XOR U139 ( .A(n139), .B(n140), .Z(DIFF[38]) );
  XOR U140 ( .A(B[38]), .B(A[38]), .Z(n140) );
  XOR U141 ( .A(n141), .B(n142), .Z(DIFF[37]) );
  XOR U142 ( .A(B[37]), .B(A[37]), .Z(n142) );
  XOR U143 ( .A(n143), .B(n144), .Z(DIFF[36]) );
  XOR U144 ( .A(B[36]), .B(A[36]), .Z(n144) );
  XOR U145 ( .A(n145), .B(n146), .Z(DIFF[35]) );
  XOR U146 ( .A(B[35]), .B(A[35]), .Z(n146) );
  XOR U147 ( .A(n147), .B(n148), .Z(DIFF[34]) );
  XOR U148 ( .A(B[34]), .B(A[34]), .Z(n148) );
  XOR U149 ( .A(n149), .B(n150), .Z(DIFF[33]) );
  XOR U150 ( .A(B[33]), .B(A[33]), .Z(n150) );
  XOR U151 ( .A(n151), .B(n152), .Z(DIFF[32]) );
  XOR U152 ( .A(B[32]), .B(A[32]), .Z(n152) );
  XOR U153 ( .A(n153), .B(n154), .Z(DIFF[31]) );
  XOR U154 ( .A(B[31]), .B(A[31]), .Z(n154) );
  XOR U155 ( .A(n155), .B(n156), .Z(DIFF[30]) );
  XOR U156 ( .A(B[30]), .B(A[30]), .Z(n156) );
  XOR U157 ( .A(n157), .B(n158), .Z(DIFF[2]) );
  XOR U158 ( .A(B[2]), .B(A[2]), .Z(n158) );
  XOR U159 ( .A(n159), .B(n160), .Z(DIFF[29]) );
  XOR U160 ( .A(B[29]), .B(A[29]), .Z(n160) );
  XOR U161 ( .A(n161), .B(n162), .Z(DIFF[28]) );
  XOR U162 ( .A(B[28]), .B(A[28]), .Z(n162) );
  XOR U163 ( .A(n163), .B(n164), .Z(DIFF[27]) );
  XOR U164 ( .A(B[27]), .B(A[27]), .Z(n164) );
  XOR U165 ( .A(n165), .B(n166), .Z(DIFF[26]) );
  XOR U166 ( .A(B[26]), .B(A[26]), .Z(n166) );
  XOR U167 ( .A(n167), .B(n168), .Z(DIFF[25]) );
  XOR U168 ( .A(B[25]), .B(A[25]), .Z(n168) );
  XOR U169 ( .A(A[257]), .B(n169), .Z(DIFF[257]) );
  ANDN U170 ( .B(n170), .A(A[256]), .Z(n169) );
  XOR U171 ( .A(A[256]), .B(n170), .Z(DIFF[256]) );
  AND U172 ( .A(n171), .B(n172), .Z(n170) );
  NANDN U173 ( .A(B[255]), .B(n173), .Z(n172) );
  NANDN U174 ( .A(A[255]), .B(n174), .Z(n173) );
  NANDN U175 ( .A(n174), .B(A[255]), .Z(n171) );
  XOR U176 ( .A(n174), .B(n175), .Z(DIFF[255]) );
  XOR U177 ( .A(B[255]), .B(A[255]), .Z(n175) );
  AND U178 ( .A(n176), .B(n177), .Z(n174) );
  NANDN U179 ( .A(B[254]), .B(n178), .Z(n177) );
  NANDN U180 ( .A(A[254]), .B(n179), .Z(n178) );
  NANDN U181 ( .A(n179), .B(A[254]), .Z(n176) );
  XOR U182 ( .A(n179), .B(n180), .Z(DIFF[254]) );
  XOR U183 ( .A(B[254]), .B(A[254]), .Z(n180) );
  AND U184 ( .A(n181), .B(n182), .Z(n179) );
  NANDN U185 ( .A(B[253]), .B(n183), .Z(n182) );
  NANDN U186 ( .A(A[253]), .B(n184), .Z(n183) );
  NANDN U187 ( .A(n184), .B(A[253]), .Z(n181) );
  XOR U188 ( .A(n184), .B(n185), .Z(DIFF[253]) );
  XOR U189 ( .A(B[253]), .B(A[253]), .Z(n185) );
  AND U190 ( .A(n186), .B(n187), .Z(n184) );
  NANDN U191 ( .A(B[252]), .B(n188), .Z(n187) );
  NANDN U192 ( .A(A[252]), .B(n189), .Z(n188) );
  NANDN U193 ( .A(n189), .B(A[252]), .Z(n186) );
  XOR U194 ( .A(n189), .B(n190), .Z(DIFF[252]) );
  XOR U195 ( .A(B[252]), .B(A[252]), .Z(n190) );
  AND U196 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U197 ( .A(B[251]), .B(n193), .Z(n192) );
  NANDN U198 ( .A(A[251]), .B(n194), .Z(n193) );
  NANDN U199 ( .A(n194), .B(A[251]), .Z(n191) );
  XOR U200 ( .A(n194), .B(n195), .Z(DIFF[251]) );
  XOR U201 ( .A(B[251]), .B(A[251]), .Z(n195) );
  AND U202 ( .A(n196), .B(n197), .Z(n194) );
  NANDN U203 ( .A(B[250]), .B(n198), .Z(n197) );
  NANDN U204 ( .A(A[250]), .B(n199), .Z(n198) );
  NANDN U205 ( .A(n199), .B(A[250]), .Z(n196) );
  XOR U206 ( .A(n199), .B(n200), .Z(DIFF[250]) );
  XOR U207 ( .A(B[250]), .B(A[250]), .Z(n200) );
  AND U208 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U209 ( .A(B[249]), .B(n203), .Z(n202) );
  NANDN U210 ( .A(A[249]), .B(n204), .Z(n203) );
  NANDN U211 ( .A(n204), .B(A[249]), .Z(n201) );
  XOR U212 ( .A(n205), .B(n206), .Z(DIFF[24]) );
  XOR U213 ( .A(B[24]), .B(A[24]), .Z(n206) );
  XOR U214 ( .A(n204), .B(n207), .Z(DIFF[249]) );
  XOR U215 ( .A(B[249]), .B(A[249]), .Z(n207) );
  AND U216 ( .A(n208), .B(n209), .Z(n204) );
  NANDN U217 ( .A(B[248]), .B(n210), .Z(n209) );
  NANDN U218 ( .A(A[248]), .B(n211), .Z(n210) );
  NANDN U219 ( .A(n211), .B(A[248]), .Z(n208) );
  XOR U220 ( .A(n211), .B(n212), .Z(DIFF[248]) );
  XOR U221 ( .A(B[248]), .B(A[248]), .Z(n212) );
  AND U222 ( .A(n213), .B(n214), .Z(n211) );
  NANDN U223 ( .A(B[247]), .B(n215), .Z(n214) );
  NANDN U224 ( .A(A[247]), .B(n216), .Z(n215) );
  NANDN U225 ( .A(n216), .B(A[247]), .Z(n213) );
  XOR U226 ( .A(n216), .B(n217), .Z(DIFF[247]) );
  XOR U227 ( .A(B[247]), .B(A[247]), .Z(n217) );
  AND U228 ( .A(n218), .B(n219), .Z(n216) );
  NANDN U229 ( .A(B[246]), .B(n220), .Z(n219) );
  NANDN U230 ( .A(A[246]), .B(n221), .Z(n220) );
  NANDN U231 ( .A(n221), .B(A[246]), .Z(n218) );
  XOR U232 ( .A(n221), .B(n222), .Z(DIFF[246]) );
  XOR U233 ( .A(B[246]), .B(A[246]), .Z(n222) );
  AND U234 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U235 ( .A(B[245]), .B(n225), .Z(n224) );
  NANDN U236 ( .A(A[245]), .B(n226), .Z(n225) );
  NANDN U237 ( .A(n226), .B(A[245]), .Z(n223) );
  XOR U238 ( .A(n226), .B(n227), .Z(DIFF[245]) );
  XOR U239 ( .A(B[245]), .B(A[245]), .Z(n227) );
  AND U240 ( .A(n228), .B(n229), .Z(n226) );
  NANDN U241 ( .A(B[244]), .B(n230), .Z(n229) );
  NANDN U242 ( .A(A[244]), .B(n231), .Z(n230) );
  NANDN U243 ( .A(n231), .B(A[244]), .Z(n228) );
  XOR U244 ( .A(n231), .B(n232), .Z(DIFF[244]) );
  XOR U245 ( .A(B[244]), .B(A[244]), .Z(n232) );
  AND U246 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U247 ( .A(B[243]), .B(n235), .Z(n234) );
  NANDN U248 ( .A(A[243]), .B(n236), .Z(n235) );
  NANDN U249 ( .A(n236), .B(A[243]), .Z(n233) );
  XOR U250 ( .A(n236), .B(n237), .Z(DIFF[243]) );
  XOR U251 ( .A(B[243]), .B(A[243]), .Z(n237) );
  AND U252 ( .A(n238), .B(n239), .Z(n236) );
  NANDN U253 ( .A(B[242]), .B(n240), .Z(n239) );
  NANDN U254 ( .A(A[242]), .B(n241), .Z(n240) );
  NANDN U255 ( .A(n241), .B(A[242]), .Z(n238) );
  XOR U256 ( .A(n241), .B(n242), .Z(DIFF[242]) );
  XOR U257 ( .A(B[242]), .B(A[242]), .Z(n242) );
  AND U258 ( .A(n243), .B(n244), .Z(n241) );
  NANDN U259 ( .A(B[241]), .B(n245), .Z(n244) );
  NANDN U260 ( .A(A[241]), .B(n246), .Z(n245) );
  NANDN U261 ( .A(n246), .B(A[241]), .Z(n243) );
  XOR U262 ( .A(n246), .B(n247), .Z(DIFF[241]) );
  XOR U263 ( .A(B[241]), .B(A[241]), .Z(n247) );
  AND U264 ( .A(n248), .B(n249), .Z(n246) );
  NANDN U265 ( .A(B[240]), .B(n250), .Z(n249) );
  NANDN U266 ( .A(A[240]), .B(n251), .Z(n250) );
  NANDN U267 ( .A(n251), .B(A[240]), .Z(n248) );
  XOR U268 ( .A(n251), .B(n252), .Z(DIFF[240]) );
  XOR U269 ( .A(B[240]), .B(A[240]), .Z(n252) );
  AND U270 ( .A(n253), .B(n254), .Z(n251) );
  NANDN U271 ( .A(B[239]), .B(n255), .Z(n254) );
  NANDN U272 ( .A(A[239]), .B(n256), .Z(n255) );
  NANDN U273 ( .A(n256), .B(A[239]), .Z(n253) );
  XOR U274 ( .A(n257), .B(n258), .Z(DIFF[23]) );
  XOR U275 ( .A(B[23]), .B(A[23]), .Z(n258) );
  XOR U276 ( .A(n256), .B(n259), .Z(DIFF[239]) );
  XOR U277 ( .A(B[239]), .B(A[239]), .Z(n259) );
  AND U278 ( .A(n260), .B(n261), .Z(n256) );
  NANDN U279 ( .A(B[238]), .B(n262), .Z(n261) );
  NANDN U280 ( .A(A[238]), .B(n263), .Z(n262) );
  NANDN U281 ( .A(n263), .B(A[238]), .Z(n260) );
  XOR U282 ( .A(n263), .B(n264), .Z(DIFF[238]) );
  XOR U283 ( .A(B[238]), .B(A[238]), .Z(n264) );
  AND U284 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U285 ( .A(B[237]), .B(n267), .Z(n266) );
  NANDN U286 ( .A(A[237]), .B(n268), .Z(n267) );
  NANDN U287 ( .A(n268), .B(A[237]), .Z(n265) );
  XOR U288 ( .A(n268), .B(n269), .Z(DIFF[237]) );
  XOR U289 ( .A(B[237]), .B(A[237]), .Z(n269) );
  AND U290 ( .A(n270), .B(n271), .Z(n268) );
  NANDN U291 ( .A(B[236]), .B(n272), .Z(n271) );
  NANDN U292 ( .A(A[236]), .B(n273), .Z(n272) );
  NANDN U293 ( .A(n273), .B(A[236]), .Z(n270) );
  XOR U294 ( .A(n273), .B(n274), .Z(DIFF[236]) );
  XOR U295 ( .A(B[236]), .B(A[236]), .Z(n274) );
  AND U296 ( .A(n275), .B(n276), .Z(n273) );
  NANDN U297 ( .A(B[235]), .B(n277), .Z(n276) );
  NANDN U298 ( .A(A[235]), .B(n278), .Z(n277) );
  NANDN U299 ( .A(n278), .B(A[235]), .Z(n275) );
  XOR U300 ( .A(n278), .B(n279), .Z(DIFF[235]) );
  XOR U301 ( .A(B[235]), .B(A[235]), .Z(n279) );
  AND U302 ( .A(n280), .B(n281), .Z(n278) );
  NANDN U303 ( .A(B[234]), .B(n282), .Z(n281) );
  NANDN U304 ( .A(A[234]), .B(n283), .Z(n282) );
  NANDN U305 ( .A(n283), .B(A[234]), .Z(n280) );
  XOR U306 ( .A(n283), .B(n284), .Z(DIFF[234]) );
  XOR U307 ( .A(B[234]), .B(A[234]), .Z(n284) );
  AND U308 ( .A(n285), .B(n286), .Z(n283) );
  NANDN U309 ( .A(B[233]), .B(n287), .Z(n286) );
  NANDN U310 ( .A(A[233]), .B(n288), .Z(n287) );
  NANDN U311 ( .A(n288), .B(A[233]), .Z(n285) );
  XOR U312 ( .A(n288), .B(n289), .Z(DIFF[233]) );
  XOR U313 ( .A(B[233]), .B(A[233]), .Z(n289) );
  AND U314 ( .A(n290), .B(n291), .Z(n288) );
  NANDN U315 ( .A(B[232]), .B(n292), .Z(n291) );
  NANDN U316 ( .A(A[232]), .B(n293), .Z(n292) );
  NANDN U317 ( .A(n293), .B(A[232]), .Z(n290) );
  XOR U318 ( .A(n293), .B(n294), .Z(DIFF[232]) );
  XOR U319 ( .A(B[232]), .B(A[232]), .Z(n294) );
  AND U320 ( .A(n295), .B(n296), .Z(n293) );
  NANDN U321 ( .A(B[231]), .B(n297), .Z(n296) );
  NANDN U322 ( .A(A[231]), .B(n298), .Z(n297) );
  NANDN U323 ( .A(n298), .B(A[231]), .Z(n295) );
  XOR U324 ( .A(n298), .B(n299), .Z(DIFF[231]) );
  XOR U325 ( .A(B[231]), .B(A[231]), .Z(n299) );
  AND U326 ( .A(n300), .B(n301), .Z(n298) );
  NANDN U327 ( .A(B[230]), .B(n302), .Z(n301) );
  NANDN U328 ( .A(A[230]), .B(n303), .Z(n302) );
  NANDN U329 ( .A(n303), .B(A[230]), .Z(n300) );
  XOR U330 ( .A(n303), .B(n304), .Z(DIFF[230]) );
  XOR U331 ( .A(B[230]), .B(A[230]), .Z(n304) );
  AND U332 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U333 ( .A(B[229]), .B(n307), .Z(n306) );
  NANDN U334 ( .A(A[229]), .B(n308), .Z(n307) );
  NANDN U335 ( .A(n308), .B(A[229]), .Z(n305) );
  XOR U336 ( .A(n309), .B(n310), .Z(DIFF[22]) );
  XOR U337 ( .A(B[22]), .B(A[22]), .Z(n310) );
  XOR U338 ( .A(n308), .B(n311), .Z(DIFF[229]) );
  XOR U339 ( .A(B[229]), .B(A[229]), .Z(n311) );
  AND U340 ( .A(n312), .B(n313), .Z(n308) );
  NANDN U341 ( .A(B[228]), .B(n314), .Z(n313) );
  NANDN U342 ( .A(A[228]), .B(n315), .Z(n314) );
  NANDN U343 ( .A(n315), .B(A[228]), .Z(n312) );
  XOR U344 ( .A(n315), .B(n316), .Z(DIFF[228]) );
  XOR U345 ( .A(B[228]), .B(A[228]), .Z(n316) );
  AND U346 ( .A(n317), .B(n318), .Z(n315) );
  NANDN U347 ( .A(B[227]), .B(n319), .Z(n318) );
  NANDN U348 ( .A(A[227]), .B(n320), .Z(n319) );
  NANDN U349 ( .A(n320), .B(A[227]), .Z(n317) );
  XOR U350 ( .A(n320), .B(n321), .Z(DIFF[227]) );
  XOR U351 ( .A(B[227]), .B(A[227]), .Z(n321) );
  AND U352 ( .A(n322), .B(n323), .Z(n320) );
  NANDN U353 ( .A(B[226]), .B(n324), .Z(n323) );
  NANDN U354 ( .A(A[226]), .B(n325), .Z(n324) );
  NANDN U355 ( .A(n325), .B(A[226]), .Z(n322) );
  XOR U356 ( .A(n325), .B(n326), .Z(DIFF[226]) );
  XOR U357 ( .A(B[226]), .B(A[226]), .Z(n326) );
  AND U358 ( .A(n327), .B(n328), .Z(n325) );
  NANDN U359 ( .A(B[225]), .B(n329), .Z(n328) );
  NANDN U360 ( .A(A[225]), .B(n330), .Z(n329) );
  NANDN U361 ( .A(n330), .B(A[225]), .Z(n327) );
  XOR U362 ( .A(n330), .B(n331), .Z(DIFF[225]) );
  XOR U363 ( .A(B[225]), .B(A[225]), .Z(n331) );
  AND U364 ( .A(n332), .B(n333), .Z(n330) );
  NANDN U365 ( .A(B[224]), .B(n334), .Z(n333) );
  NANDN U366 ( .A(A[224]), .B(n335), .Z(n334) );
  NANDN U367 ( .A(n335), .B(A[224]), .Z(n332) );
  XOR U368 ( .A(n335), .B(n336), .Z(DIFF[224]) );
  XOR U369 ( .A(B[224]), .B(A[224]), .Z(n336) );
  AND U370 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U371 ( .A(B[223]), .B(n339), .Z(n338) );
  NANDN U372 ( .A(A[223]), .B(n340), .Z(n339) );
  NANDN U373 ( .A(n340), .B(A[223]), .Z(n337) );
  XOR U374 ( .A(n340), .B(n341), .Z(DIFF[223]) );
  XOR U375 ( .A(B[223]), .B(A[223]), .Z(n341) );
  AND U376 ( .A(n342), .B(n343), .Z(n340) );
  NANDN U377 ( .A(B[222]), .B(n344), .Z(n343) );
  NANDN U378 ( .A(A[222]), .B(n345), .Z(n344) );
  NANDN U379 ( .A(n345), .B(A[222]), .Z(n342) );
  XOR U380 ( .A(n345), .B(n346), .Z(DIFF[222]) );
  XOR U381 ( .A(B[222]), .B(A[222]), .Z(n346) );
  AND U382 ( .A(n347), .B(n348), .Z(n345) );
  NANDN U383 ( .A(B[221]), .B(n349), .Z(n348) );
  NANDN U384 ( .A(A[221]), .B(n350), .Z(n349) );
  NANDN U385 ( .A(n350), .B(A[221]), .Z(n347) );
  XOR U386 ( .A(n350), .B(n351), .Z(DIFF[221]) );
  XOR U387 ( .A(B[221]), .B(A[221]), .Z(n351) );
  AND U388 ( .A(n352), .B(n353), .Z(n350) );
  NANDN U389 ( .A(B[220]), .B(n354), .Z(n353) );
  NANDN U390 ( .A(A[220]), .B(n355), .Z(n354) );
  NANDN U391 ( .A(n355), .B(A[220]), .Z(n352) );
  XOR U392 ( .A(n355), .B(n356), .Z(DIFF[220]) );
  XOR U393 ( .A(B[220]), .B(A[220]), .Z(n356) );
  AND U394 ( .A(n357), .B(n358), .Z(n355) );
  NANDN U395 ( .A(B[219]), .B(n359), .Z(n358) );
  NANDN U396 ( .A(A[219]), .B(n360), .Z(n359) );
  NANDN U397 ( .A(n360), .B(A[219]), .Z(n357) );
  XOR U398 ( .A(n361), .B(n362), .Z(DIFF[21]) );
  XOR U399 ( .A(B[21]), .B(A[21]), .Z(n362) );
  XOR U400 ( .A(n360), .B(n363), .Z(DIFF[219]) );
  XOR U401 ( .A(B[219]), .B(A[219]), .Z(n363) );
  AND U402 ( .A(n364), .B(n365), .Z(n360) );
  NANDN U403 ( .A(B[218]), .B(n366), .Z(n365) );
  NANDN U404 ( .A(A[218]), .B(n367), .Z(n366) );
  NANDN U405 ( .A(n367), .B(A[218]), .Z(n364) );
  XOR U406 ( .A(n367), .B(n368), .Z(DIFF[218]) );
  XOR U407 ( .A(B[218]), .B(A[218]), .Z(n368) );
  AND U408 ( .A(n369), .B(n370), .Z(n367) );
  NANDN U409 ( .A(B[217]), .B(n371), .Z(n370) );
  NANDN U410 ( .A(A[217]), .B(n372), .Z(n371) );
  NANDN U411 ( .A(n372), .B(A[217]), .Z(n369) );
  XOR U412 ( .A(n372), .B(n373), .Z(DIFF[217]) );
  XOR U413 ( .A(B[217]), .B(A[217]), .Z(n373) );
  AND U414 ( .A(n374), .B(n375), .Z(n372) );
  NANDN U415 ( .A(B[216]), .B(n376), .Z(n375) );
  NANDN U416 ( .A(A[216]), .B(n377), .Z(n376) );
  NANDN U417 ( .A(n377), .B(A[216]), .Z(n374) );
  XOR U418 ( .A(n377), .B(n378), .Z(DIFF[216]) );
  XOR U419 ( .A(B[216]), .B(A[216]), .Z(n378) );
  AND U420 ( .A(n379), .B(n380), .Z(n377) );
  NANDN U421 ( .A(B[215]), .B(n381), .Z(n380) );
  NANDN U422 ( .A(A[215]), .B(n382), .Z(n381) );
  NANDN U423 ( .A(n382), .B(A[215]), .Z(n379) );
  XOR U424 ( .A(n382), .B(n383), .Z(DIFF[215]) );
  XOR U425 ( .A(B[215]), .B(A[215]), .Z(n383) );
  AND U426 ( .A(n384), .B(n385), .Z(n382) );
  NANDN U427 ( .A(B[214]), .B(n386), .Z(n385) );
  NANDN U428 ( .A(A[214]), .B(n387), .Z(n386) );
  NANDN U429 ( .A(n387), .B(A[214]), .Z(n384) );
  XOR U430 ( .A(n387), .B(n388), .Z(DIFF[214]) );
  XOR U431 ( .A(B[214]), .B(A[214]), .Z(n388) );
  AND U432 ( .A(n389), .B(n390), .Z(n387) );
  NANDN U433 ( .A(B[213]), .B(n391), .Z(n390) );
  NANDN U434 ( .A(A[213]), .B(n392), .Z(n391) );
  NANDN U435 ( .A(n392), .B(A[213]), .Z(n389) );
  XOR U436 ( .A(n392), .B(n393), .Z(DIFF[213]) );
  XOR U437 ( .A(B[213]), .B(A[213]), .Z(n393) );
  AND U438 ( .A(n394), .B(n395), .Z(n392) );
  NANDN U439 ( .A(B[212]), .B(n396), .Z(n395) );
  NANDN U440 ( .A(A[212]), .B(n397), .Z(n396) );
  NANDN U441 ( .A(n397), .B(A[212]), .Z(n394) );
  XOR U442 ( .A(n397), .B(n398), .Z(DIFF[212]) );
  XOR U443 ( .A(B[212]), .B(A[212]), .Z(n398) );
  AND U444 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U445 ( .A(B[211]), .B(n401), .Z(n400) );
  NANDN U446 ( .A(A[211]), .B(n402), .Z(n401) );
  NANDN U447 ( .A(n402), .B(A[211]), .Z(n399) );
  XOR U448 ( .A(n402), .B(n403), .Z(DIFF[211]) );
  XOR U449 ( .A(B[211]), .B(A[211]), .Z(n403) );
  AND U450 ( .A(n404), .B(n405), .Z(n402) );
  NANDN U451 ( .A(B[210]), .B(n406), .Z(n405) );
  NANDN U452 ( .A(A[210]), .B(n407), .Z(n406) );
  NANDN U453 ( .A(n407), .B(A[210]), .Z(n404) );
  XOR U454 ( .A(n407), .B(n408), .Z(DIFF[210]) );
  XOR U455 ( .A(B[210]), .B(A[210]), .Z(n408) );
  AND U456 ( .A(n409), .B(n410), .Z(n407) );
  NANDN U457 ( .A(B[209]), .B(n411), .Z(n410) );
  NANDN U458 ( .A(A[209]), .B(n412), .Z(n411) );
  NANDN U459 ( .A(n412), .B(A[209]), .Z(n409) );
  XOR U460 ( .A(n413), .B(n414), .Z(DIFF[20]) );
  XOR U461 ( .A(B[20]), .B(A[20]), .Z(n414) );
  XOR U462 ( .A(n412), .B(n415), .Z(DIFF[209]) );
  XOR U463 ( .A(B[209]), .B(A[209]), .Z(n415) );
  AND U464 ( .A(n416), .B(n417), .Z(n412) );
  NANDN U465 ( .A(B[208]), .B(n418), .Z(n417) );
  NANDN U466 ( .A(A[208]), .B(n419), .Z(n418) );
  NANDN U467 ( .A(n419), .B(A[208]), .Z(n416) );
  XOR U468 ( .A(n419), .B(n420), .Z(DIFF[208]) );
  XOR U469 ( .A(B[208]), .B(A[208]), .Z(n420) );
  AND U470 ( .A(n421), .B(n422), .Z(n419) );
  NANDN U471 ( .A(B[207]), .B(n423), .Z(n422) );
  NANDN U472 ( .A(A[207]), .B(n424), .Z(n423) );
  NANDN U473 ( .A(n424), .B(A[207]), .Z(n421) );
  XOR U474 ( .A(n424), .B(n425), .Z(DIFF[207]) );
  XOR U475 ( .A(B[207]), .B(A[207]), .Z(n425) );
  AND U476 ( .A(n426), .B(n427), .Z(n424) );
  NANDN U477 ( .A(B[206]), .B(n428), .Z(n427) );
  NANDN U478 ( .A(A[206]), .B(n429), .Z(n428) );
  NANDN U479 ( .A(n429), .B(A[206]), .Z(n426) );
  XOR U480 ( .A(n429), .B(n430), .Z(DIFF[206]) );
  XOR U481 ( .A(B[206]), .B(A[206]), .Z(n430) );
  AND U482 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U483 ( .A(B[205]), .B(n433), .Z(n432) );
  NANDN U484 ( .A(A[205]), .B(n434), .Z(n433) );
  NANDN U485 ( .A(n434), .B(A[205]), .Z(n431) );
  XOR U486 ( .A(n434), .B(n435), .Z(DIFF[205]) );
  XOR U487 ( .A(B[205]), .B(A[205]), .Z(n435) );
  AND U488 ( .A(n436), .B(n437), .Z(n434) );
  NANDN U489 ( .A(B[204]), .B(n438), .Z(n437) );
  NANDN U490 ( .A(A[204]), .B(n439), .Z(n438) );
  NANDN U491 ( .A(n439), .B(A[204]), .Z(n436) );
  XOR U492 ( .A(n439), .B(n440), .Z(DIFF[204]) );
  XOR U493 ( .A(B[204]), .B(A[204]), .Z(n440) );
  AND U494 ( .A(n441), .B(n442), .Z(n439) );
  NANDN U495 ( .A(B[203]), .B(n443), .Z(n442) );
  NANDN U496 ( .A(A[203]), .B(n444), .Z(n443) );
  NANDN U497 ( .A(n444), .B(A[203]), .Z(n441) );
  XOR U498 ( .A(n444), .B(n445), .Z(DIFF[203]) );
  XOR U499 ( .A(B[203]), .B(A[203]), .Z(n445) );
  AND U500 ( .A(n446), .B(n447), .Z(n444) );
  NANDN U501 ( .A(B[202]), .B(n448), .Z(n447) );
  NANDN U502 ( .A(A[202]), .B(n449), .Z(n448) );
  NANDN U503 ( .A(n449), .B(A[202]), .Z(n446) );
  XOR U504 ( .A(n449), .B(n450), .Z(DIFF[202]) );
  XOR U505 ( .A(B[202]), .B(A[202]), .Z(n450) );
  AND U506 ( .A(n451), .B(n452), .Z(n449) );
  NANDN U507 ( .A(B[201]), .B(n453), .Z(n452) );
  NANDN U508 ( .A(A[201]), .B(n454), .Z(n453) );
  NANDN U509 ( .A(n454), .B(A[201]), .Z(n451) );
  XOR U510 ( .A(n454), .B(n455), .Z(DIFF[201]) );
  XOR U511 ( .A(B[201]), .B(A[201]), .Z(n455) );
  AND U512 ( .A(n456), .B(n457), .Z(n454) );
  NANDN U513 ( .A(B[200]), .B(n458), .Z(n457) );
  NANDN U514 ( .A(A[200]), .B(n459), .Z(n458) );
  NANDN U515 ( .A(n459), .B(A[200]), .Z(n456) );
  XOR U516 ( .A(n459), .B(n460), .Z(DIFF[200]) );
  XOR U517 ( .A(B[200]), .B(A[200]), .Z(n460) );
  AND U518 ( .A(n461), .B(n462), .Z(n459) );
  NANDN U519 ( .A(B[199]), .B(n463), .Z(n462) );
  NANDN U520 ( .A(A[199]), .B(n464), .Z(n463) );
  NANDN U521 ( .A(n464), .B(A[199]), .Z(n461) );
  XOR U522 ( .A(n1), .B(n465), .Z(DIFF[1]) );
  XOR U523 ( .A(B[1]), .B(A[1]), .Z(n465) );
  XOR U524 ( .A(n466), .B(n467), .Z(DIFF[19]) );
  XOR U525 ( .A(B[19]), .B(A[19]), .Z(n467) );
  XOR U526 ( .A(n464), .B(n468), .Z(DIFF[199]) );
  XOR U527 ( .A(B[199]), .B(A[199]), .Z(n468) );
  AND U528 ( .A(n469), .B(n470), .Z(n464) );
  NANDN U529 ( .A(B[198]), .B(n471), .Z(n470) );
  NANDN U530 ( .A(A[198]), .B(n472), .Z(n471) );
  NANDN U531 ( .A(n472), .B(A[198]), .Z(n469) );
  XOR U532 ( .A(n472), .B(n473), .Z(DIFF[198]) );
  XOR U533 ( .A(B[198]), .B(A[198]), .Z(n473) );
  AND U534 ( .A(n474), .B(n475), .Z(n472) );
  NANDN U535 ( .A(B[197]), .B(n476), .Z(n475) );
  NANDN U536 ( .A(A[197]), .B(n477), .Z(n476) );
  NANDN U537 ( .A(n477), .B(A[197]), .Z(n474) );
  XOR U538 ( .A(n477), .B(n478), .Z(DIFF[197]) );
  XOR U539 ( .A(B[197]), .B(A[197]), .Z(n478) );
  AND U540 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U541 ( .A(B[196]), .B(n481), .Z(n480) );
  NANDN U542 ( .A(A[196]), .B(n482), .Z(n481) );
  NANDN U543 ( .A(n482), .B(A[196]), .Z(n479) );
  XOR U544 ( .A(n482), .B(n483), .Z(DIFF[196]) );
  XOR U545 ( .A(B[196]), .B(A[196]), .Z(n483) );
  AND U546 ( .A(n484), .B(n485), .Z(n482) );
  NANDN U547 ( .A(B[195]), .B(n486), .Z(n485) );
  NANDN U548 ( .A(A[195]), .B(n487), .Z(n486) );
  NANDN U549 ( .A(n487), .B(A[195]), .Z(n484) );
  XOR U550 ( .A(n487), .B(n488), .Z(DIFF[195]) );
  XOR U551 ( .A(B[195]), .B(A[195]), .Z(n488) );
  AND U552 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U553 ( .A(B[194]), .B(n491), .Z(n490) );
  NANDN U554 ( .A(A[194]), .B(n492), .Z(n491) );
  NANDN U555 ( .A(n492), .B(A[194]), .Z(n489) );
  XOR U556 ( .A(n492), .B(n493), .Z(DIFF[194]) );
  XOR U557 ( .A(B[194]), .B(A[194]), .Z(n493) );
  AND U558 ( .A(n494), .B(n495), .Z(n492) );
  NANDN U559 ( .A(B[193]), .B(n496), .Z(n495) );
  NANDN U560 ( .A(A[193]), .B(n497), .Z(n496) );
  NANDN U561 ( .A(n497), .B(A[193]), .Z(n494) );
  XOR U562 ( .A(n497), .B(n498), .Z(DIFF[193]) );
  XOR U563 ( .A(B[193]), .B(A[193]), .Z(n498) );
  AND U564 ( .A(n499), .B(n500), .Z(n497) );
  NANDN U565 ( .A(B[192]), .B(n501), .Z(n500) );
  NANDN U566 ( .A(A[192]), .B(n502), .Z(n501) );
  NANDN U567 ( .A(n502), .B(A[192]), .Z(n499) );
  XOR U568 ( .A(n502), .B(n503), .Z(DIFF[192]) );
  XOR U569 ( .A(B[192]), .B(A[192]), .Z(n503) );
  AND U570 ( .A(n504), .B(n505), .Z(n502) );
  NANDN U571 ( .A(B[191]), .B(n506), .Z(n505) );
  NANDN U572 ( .A(A[191]), .B(n507), .Z(n506) );
  NANDN U573 ( .A(n507), .B(A[191]), .Z(n504) );
  XOR U574 ( .A(n507), .B(n508), .Z(DIFF[191]) );
  XOR U575 ( .A(B[191]), .B(A[191]), .Z(n508) );
  AND U576 ( .A(n509), .B(n510), .Z(n507) );
  NANDN U577 ( .A(B[190]), .B(n511), .Z(n510) );
  NANDN U578 ( .A(A[190]), .B(n512), .Z(n511) );
  NANDN U579 ( .A(n512), .B(A[190]), .Z(n509) );
  XOR U580 ( .A(n512), .B(n513), .Z(DIFF[190]) );
  XOR U581 ( .A(B[190]), .B(A[190]), .Z(n513) );
  AND U582 ( .A(n514), .B(n515), .Z(n512) );
  NANDN U583 ( .A(B[189]), .B(n516), .Z(n515) );
  NANDN U584 ( .A(A[189]), .B(n517), .Z(n516) );
  NANDN U585 ( .A(n517), .B(A[189]), .Z(n514) );
  XOR U586 ( .A(n518), .B(n519), .Z(DIFF[18]) );
  XOR U587 ( .A(B[18]), .B(A[18]), .Z(n519) );
  XOR U588 ( .A(n517), .B(n520), .Z(DIFF[189]) );
  XOR U589 ( .A(B[189]), .B(A[189]), .Z(n520) );
  AND U590 ( .A(n521), .B(n522), .Z(n517) );
  NANDN U591 ( .A(B[188]), .B(n523), .Z(n522) );
  NANDN U592 ( .A(A[188]), .B(n524), .Z(n523) );
  NANDN U593 ( .A(n524), .B(A[188]), .Z(n521) );
  XOR U594 ( .A(n524), .B(n525), .Z(DIFF[188]) );
  XOR U595 ( .A(B[188]), .B(A[188]), .Z(n525) );
  AND U596 ( .A(n526), .B(n527), .Z(n524) );
  NANDN U597 ( .A(B[187]), .B(n528), .Z(n527) );
  NANDN U598 ( .A(A[187]), .B(n529), .Z(n528) );
  NANDN U599 ( .A(n529), .B(A[187]), .Z(n526) );
  XOR U600 ( .A(n529), .B(n530), .Z(DIFF[187]) );
  XOR U601 ( .A(B[187]), .B(A[187]), .Z(n530) );
  AND U602 ( .A(n531), .B(n532), .Z(n529) );
  NANDN U603 ( .A(B[186]), .B(n533), .Z(n532) );
  NANDN U604 ( .A(A[186]), .B(n534), .Z(n533) );
  NANDN U605 ( .A(n534), .B(A[186]), .Z(n531) );
  XOR U606 ( .A(n534), .B(n535), .Z(DIFF[186]) );
  XOR U607 ( .A(B[186]), .B(A[186]), .Z(n535) );
  AND U608 ( .A(n536), .B(n537), .Z(n534) );
  NANDN U609 ( .A(B[185]), .B(n538), .Z(n537) );
  NANDN U610 ( .A(A[185]), .B(n539), .Z(n538) );
  NANDN U611 ( .A(n539), .B(A[185]), .Z(n536) );
  XOR U612 ( .A(n539), .B(n540), .Z(DIFF[185]) );
  XOR U613 ( .A(B[185]), .B(A[185]), .Z(n540) );
  AND U614 ( .A(n541), .B(n542), .Z(n539) );
  NANDN U615 ( .A(B[184]), .B(n543), .Z(n542) );
  NANDN U616 ( .A(A[184]), .B(n544), .Z(n543) );
  NANDN U617 ( .A(n544), .B(A[184]), .Z(n541) );
  XOR U618 ( .A(n544), .B(n545), .Z(DIFF[184]) );
  XOR U619 ( .A(B[184]), .B(A[184]), .Z(n545) );
  AND U620 ( .A(n546), .B(n547), .Z(n544) );
  NANDN U621 ( .A(B[183]), .B(n548), .Z(n547) );
  NANDN U622 ( .A(A[183]), .B(n549), .Z(n548) );
  NANDN U623 ( .A(n549), .B(A[183]), .Z(n546) );
  XOR U624 ( .A(n549), .B(n550), .Z(DIFF[183]) );
  XOR U625 ( .A(B[183]), .B(A[183]), .Z(n550) );
  AND U626 ( .A(n551), .B(n552), .Z(n549) );
  NANDN U627 ( .A(B[182]), .B(n553), .Z(n552) );
  NANDN U628 ( .A(A[182]), .B(n554), .Z(n553) );
  NANDN U629 ( .A(n554), .B(A[182]), .Z(n551) );
  XOR U630 ( .A(n554), .B(n555), .Z(DIFF[182]) );
  XOR U631 ( .A(B[182]), .B(A[182]), .Z(n555) );
  AND U632 ( .A(n556), .B(n557), .Z(n554) );
  NANDN U633 ( .A(B[181]), .B(n558), .Z(n557) );
  NANDN U634 ( .A(A[181]), .B(n559), .Z(n558) );
  NANDN U635 ( .A(n559), .B(A[181]), .Z(n556) );
  XOR U636 ( .A(n559), .B(n560), .Z(DIFF[181]) );
  XOR U637 ( .A(B[181]), .B(A[181]), .Z(n560) );
  AND U638 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U639 ( .A(B[180]), .B(n563), .Z(n562) );
  NANDN U640 ( .A(A[180]), .B(n564), .Z(n563) );
  NANDN U641 ( .A(n564), .B(A[180]), .Z(n561) );
  XOR U642 ( .A(n564), .B(n565), .Z(DIFF[180]) );
  XOR U643 ( .A(B[180]), .B(A[180]), .Z(n565) );
  AND U644 ( .A(n566), .B(n567), .Z(n564) );
  NANDN U645 ( .A(B[179]), .B(n568), .Z(n567) );
  NANDN U646 ( .A(A[179]), .B(n569), .Z(n568) );
  NANDN U647 ( .A(n569), .B(A[179]), .Z(n566) );
  XOR U648 ( .A(n570), .B(n571), .Z(DIFF[17]) );
  XOR U649 ( .A(B[17]), .B(A[17]), .Z(n571) );
  XOR U650 ( .A(n569), .B(n572), .Z(DIFF[179]) );
  XOR U651 ( .A(B[179]), .B(A[179]), .Z(n572) );
  AND U652 ( .A(n573), .B(n574), .Z(n569) );
  NANDN U653 ( .A(B[178]), .B(n575), .Z(n574) );
  NANDN U654 ( .A(A[178]), .B(n576), .Z(n575) );
  NANDN U655 ( .A(n576), .B(A[178]), .Z(n573) );
  XOR U656 ( .A(n576), .B(n577), .Z(DIFF[178]) );
  XOR U657 ( .A(B[178]), .B(A[178]), .Z(n577) );
  AND U658 ( .A(n578), .B(n579), .Z(n576) );
  NANDN U659 ( .A(B[177]), .B(n580), .Z(n579) );
  NANDN U660 ( .A(A[177]), .B(n581), .Z(n580) );
  NANDN U661 ( .A(n581), .B(A[177]), .Z(n578) );
  XOR U662 ( .A(n581), .B(n582), .Z(DIFF[177]) );
  XOR U663 ( .A(B[177]), .B(A[177]), .Z(n582) );
  AND U664 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U665 ( .A(B[176]), .B(n585), .Z(n584) );
  NANDN U666 ( .A(A[176]), .B(n586), .Z(n585) );
  NANDN U667 ( .A(n586), .B(A[176]), .Z(n583) );
  XOR U668 ( .A(n586), .B(n587), .Z(DIFF[176]) );
  XOR U669 ( .A(B[176]), .B(A[176]), .Z(n587) );
  AND U670 ( .A(n588), .B(n589), .Z(n586) );
  NANDN U671 ( .A(B[175]), .B(n590), .Z(n589) );
  NANDN U672 ( .A(A[175]), .B(n591), .Z(n590) );
  NANDN U673 ( .A(n591), .B(A[175]), .Z(n588) );
  XOR U674 ( .A(n591), .B(n592), .Z(DIFF[175]) );
  XOR U675 ( .A(B[175]), .B(A[175]), .Z(n592) );
  AND U676 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U677 ( .A(B[174]), .B(n595), .Z(n594) );
  NANDN U678 ( .A(A[174]), .B(n596), .Z(n595) );
  NANDN U679 ( .A(n596), .B(A[174]), .Z(n593) );
  XOR U680 ( .A(n596), .B(n597), .Z(DIFF[174]) );
  XOR U681 ( .A(B[174]), .B(A[174]), .Z(n597) );
  AND U682 ( .A(n598), .B(n599), .Z(n596) );
  NANDN U683 ( .A(B[173]), .B(n600), .Z(n599) );
  NANDN U684 ( .A(A[173]), .B(n601), .Z(n600) );
  NANDN U685 ( .A(n601), .B(A[173]), .Z(n598) );
  XOR U686 ( .A(n601), .B(n602), .Z(DIFF[173]) );
  XOR U687 ( .A(B[173]), .B(A[173]), .Z(n602) );
  AND U688 ( .A(n603), .B(n604), .Z(n601) );
  NANDN U689 ( .A(B[172]), .B(n605), .Z(n604) );
  NANDN U690 ( .A(A[172]), .B(n606), .Z(n605) );
  NANDN U691 ( .A(n606), .B(A[172]), .Z(n603) );
  XOR U692 ( .A(n606), .B(n607), .Z(DIFF[172]) );
  XOR U693 ( .A(B[172]), .B(A[172]), .Z(n607) );
  AND U694 ( .A(n608), .B(n609), .Z(n606) );
  NANDN U695 ( .A(B[171]), .B(n610), .Z(n609) );
  NANDN U696 ( .A(A[171]), .B(n611), .Z(n610) );
  NANDN U697 ( .A(n611), .B(A[171]), .Z(n608) );
  XOR U698 ( .A(n611), .B(n612), .Z(DIFF[171]) );
  XOR U699 ( .A(B[171]), .B(A[171]), .Z(n612) );
  AND U700 ( .A(n613), .B(n614), .Z(n611) );
  NANDN U701 ( .A(B[170]), .B(n615), .Z(n614) );
  NANDN U702 ( .A(A[170]), .B(n616), .Z(n615) );
  NANDN U703 ( .A(n616), .B(A[170]), .Z(n613) );
  XOR U704 ( .A(n616), .B(n617), .Z(DIFF[170]) );
  XOR U705 ( .A(B[170]), .B(A[170]), .Z(n617) );
  AND U706 ( .A(n618), .B(n619), .Z(n616) );
  NANDN U707 ( .A(B[169]), .B(n620), .Z(n619) );
  NANDN U708 ( .A(A[169]), .B(n621), .Z(n620) );
  NANDN U709 ( .A(n621), .B(A[169]), .Z(n618) );
  XOR U710 ( .A(n622), .B(n623), .Z(DIFF[16]) );
  XOR U711 ( .A(B[16]), .B(A[16]), .Z(n623) );
  XOR U712 ( .A(n621), .B(n624), .Z(DIFF[169]) );
  XOR U713 ( .A(B[169]), .B(A[169]), .Z(n624) );
  AND U714 ( .A(n625), .B(n626), .Z(n621) );
  NANDN U715 ( .A(B[168]), .B(n627), .Z(n626) );
  NANDN U716 ( .A(A[168]), .B(n628), .Z(n627) );
  NANDN U717 ( .A(n628), .B(A[168]), .Z(n625) );
  XOR U718 ( .A(n628), .B(n629), .Z(DIFF[168]) );
  XOR U719 ( .A(B[168]), .B(A[168]), .Z(n629) );
  AND U720 ( .A(n630), .B(n631), .Z(n628) );
  NANDN U721 ( .A(B[167]), .B(n632), .Z(n631) );
  NANDN U722 ( .A(A[167]), .B(n633), .Z(n632) );
  NANDN U723 ( .A(n633), .B(A[167]), .Z(n630) );
  XOR U724 ( .A(n633), .B(n634), .Z(DIFF[167]) );
  XOR U725 ( .A(B[167]), .B(A[167]), .Z(n634) );
  AND U726 ( .A(n635), .B(n636), .Z(n633) );
  NANDN U727 ( .A(B[166]), .B(n637), .Z(n636) );
  NANDN U728 ( .A(A[166]), .B(n638), .Z(n637) );
  NANDN U729 ( .A(n638), .B(A[166]), .Z(n635) );
  XOR U730 ( .A(n638), .B(n639), .Z(DIFF[166]) );
  XOR U731 ( .A(B[166]), .B(A[166]), .Z(n639) );
  AND U732 ( .A(n640), .B(n641), .Z(n638) );
  NANDN U733 ( .A(B[165]), .B(n642), .Z(n641) );
  NANDN U734 ( .A(A[165]), .B(n643), .Z(n642) );
  NANDN U735 ( .A(n643), .B(A[165]), .Z(n640) );
  XOR U736 ( .A(n643), .B(n644), .Z(DIFF[165]) );
  XOR U737 ( .A(B[165]), .B(A[165]), .Z(n644) );
  AND U738 ( .A(n645), .B(n646), .Z(n643) );
  NANDN U739 ( .A(B[164]), .B(n647), .Z(n646) );
  NANDN U740 ( .A(A[164]), .B(n648), .Z(n647) );
  NANDN U741 ( .A(n648), .B(A[164]), .Z(n645) );
  XOR U742 ( .A(n648), .B(n649), .Z(DIFF[164]) );
  XOR U743 ( .A(B[164]), .B(A[164]), .Z(n649) );
  AND U744 ( .A(n650), .B(n651), .Z(n648) );
  NANDN U745 ( .A(B[163]), .B(n652), .Z(n651) );
  NANDN U746 ( .A(A[163]), .B(n653), .Z(n652) );
  NANDN U747 ( .A(n653), .B(A[163]), .Z(n650) );
  XOR U748 ( .A(n653), .B(n654), .Z(DIFF[163]) );
  XOR U749 ( .A(B[163]), .B(A[163]), .Z(n654) );
  AND U750 ( .A(n655), .B(n656), .Z(n653) );
  NANDN U751 ( .A(B[162]), .B(n657), .Z(n656) );
  NANDN U752 ( .A(A[162]), .B(n658), .Z(n657) );
  NANDN U753 ( .A(n658), .B(A[162]), .Z(n655) );
  XOR U754 ( .A(n658), .B(n659), .Z(DIFF[162]) );
  XOR U755 ( .A(B[162]), .B(A[162]), .Z(n659) );
  AND U756 ( .A(n660), .B(n661), .Z(n658) );
  NANDN U757 ( .A(B[161]), .B(n662), .Z(n661) );
  NANDN U758 ( .A(A[161]), .B(n663), .Z(n662) );
  NANDN U759 ( .A(n663), .B(A[161]), .Z(n660) );
  XOR U760 ( .A(n663), .B(n664), .Z(DIFF[161]) );
  XOR U761 ( .A(B[161]), .B(A[161]), .Z(n664) );
  AND U762 ( .A(n665), .B(n666), .Z(n663) );
  NANDN U763 ( .A(B[160]), .B(n667), .Z(n666) );
  NANDN U764 ( .A(A[160]), .B(n668), .Z(n667) );
  NANDN U765 ( .A(n668), .B(A[160]), .Z(n665) );
  XOR U766 ( .A(n668), .B(n669), .Z(DIFF[160]) );
  XOR U767 ( .A(B[160]), .B(A[160]), .Z(n669) );
  AND U768 ( .A(n670), .B(n671), .Z(n668) );
  NANDN U769 ( .A(B[159]), .B(n672), .Z(n671) );
  NANDN U770 ( .A(A[159]), .B(n673), .Z(n672) );
  NANDN U771 ( .A(n673), .B(A[159]), .Z(n670) );
  XOR U772 ( .A(n674), .B(n675), .Z(DIFF[15]) );
  XOR U773 ( .A(B[15]), .B(A[15]), .Z(n675) );
  XOR U774 ( .A(n673), .B(n676), .Z(DIFF[159]) );
  XOR U775 ( .A(B[159]), .B(A[159]), .Z(n676) );
  AND U776 ( .A(n677), .B(n678), .Z(n673) );
  NANDN U777 ( .A(B[158]), .B(n679), .Z(n678) );
  NANDN U778 ( .A(A[158]), .B(n680), .Z(n679) );
  NANDN U779 ( .A(n680), .B(A[158]), .Z(n677) );
  XOR U780 ( .A(n680), .B(n681), .Z(DIFF[158]) );
  XOR U781 ( .A(B[158]), .B(A[158]), .Z(n681) );
  AND U782 ( .A(n682), .B(n683), .Z(n680) );
  NANDN U783 ( .A(B[157]), .B(n684), .Z(n683) );
  NANDN U784 ( .A(A[157]), .B(n685), .Z(n684) );
  NANDN U785 ( .A(n685), .B(A[157]), .Z(n682) );
  XOR U786 ( .A(n685), .B(n686), .Z(DIFF[157]) );
  XOR U787 ( .A(B[157]), .B(A[157]), .Z(n686) );
  AND U788 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U789 ( .A(B[156]), .B(n689), .Z(n688) );
  NANDN U790 ( .A(A[156]), .B(n690), .Z(n689) );
  NANDN U791 ( .A(n690), .B(A[156]), .Z(n687) );
  XOR U792 ( .A(n690), .B(n691), .Z(DIFF[156]) );
  XOR U793 ( .A(B[156]), .B(A[156]), .Z(n691) );
  AND U794 ( .A(n692), .B(n693), .Z(n690) );
  NANDN U795 ( .A(B[155]), .B(n694), .Z(n693) );
  NANDN U796 ( .A(A[155]), .B(n695), .Z(n694) );
  NANDN U797 ( .A(n695), .B(A[155]), .Z(n692) );
  XOR U798 ( .A(n695), .B(n696), .Z(DIFF[155]) );
  XOR U799 ( .A(B[155]), .B(A[155]), .Z(n696) );
  AND U800 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U801 ( .A(B[154]), .B(n699), .Z(n698) );
  NANDN U802 ( .A(A[154]), .B(n700), .Z(n699) );
  NANDN U803 ( .A(n700), .B(A[154]), .Z(n697) );
  XOR U804 ( .A(n700), .B(n701), .Z(DIFF[154]) );
  XOR U805 ( .A(B[154]), .B(A[154]), .Z(n701) );
  AND U806 ( .A(n702), .B(n703), .Z(n700) );
  NANDN U807 ( .A(B[153]), .B(n704), .Z(n703) );
  NANDN U808 ( .A(A[153]), .B(n705), .Z(n704) );
  NANDN U809 ( .A(n705), .B(A[153]), .Z(n702) );
  XOR U810 ( .A(n705), .B(n706), .Z(DIFF[153]) );
  XOR U811 ( .A(B[153]), .B(A[153]), .Z(n706) );
  AND U812 ( .A(n707), .B(n708), .Z(n705) );
  NANDN U813 ( .A(B[152]), .B(n709), .Z(n708) );
  NANDN U814 ( .A(A[152]), .B(n710), .Z(n709) );
  NANDN U815 ( .A(n710), .B(A[152]), .Z(n707) );
  XOR U816 ( .A(n710), .B(n711), .Z(DIFF[152]) );
  XOR U817 ( .A(B[152]), .B(A[152]), .Z(n711) );
  AND U818 ( .A(n712), .B(n713), .Z(n710) );
  NANDN U819 ( .A(B[151]), .B(n714), .Z(n713) );
  NANDN U820 ( .A(A[151]), .B(n715), .Z(n714) );
  NANDN U821 ( .A(n715), .B(A[151]), .Z(n712) );
  XOR U822 ( .A(n715), .B(n716), .Z(DIFF[151]) );
  XOR U823 ( .A(B[151]), .B(A[151]), .Z(n716) );
  AND U824 ( .A(n717), .B(n718), .Z(n715) );
  NANDN U825 ( .A(B[150]), .B(n719), .Z(n718) );
  NANDN U826 ( .A(A[150]), .B(n720), .Z(n719) );
  NANDN U827 ( .A(n720), .B(A[150]), .Z(n717) );
  XOR U828 ( .A(n720), .B(n721), .Z(DIFF[150]) );
  XOR U829 ( .A(B[150]), .B(A[150]), .Z(n721) );
  AND U830 ( .A(n722), .B(n723), .Z(n720) );
  NANDN U831 ( .A(B[149]), .B(n724), .Z(n723) );
  NANDN U832 ( .A(A[149]), .B(n725), .Z(n724) );
  NANDN U833 ( .A(n725), .B(A[149]), .Z(n722) );
  XOR U834 ( .A(n726), .B(n727), .Z(DIFF[14]) );
  XOR U835 ( .A(B[14]), .B(A[14]), .Z(n727) );
  XOR U836 ( .A(n725), .B(n728), .Z(DIFF[149]) );
  XOR U837 ( .A(B[149]), .B(A[149]), .Z(n728) );
  AND U838 ( .A(n729), .B(n730), .Z(n725) );
  NANDN U839 ( .A(B[148]), .B(n731), .Z(n730) );
  NANDN U840 ( .A(A[148]), .B(n732), .Z(n731) );
  NANDN U841 ( .A(n732), .B(A[148]), .Z(n729) );
  XOR U842 ( .A(n732), .B(n733), .Z(DIFF[148]) );
  XOR U843 ( .A(B[148]), .B(A[148]), .Z(n733) );
  AND U844 ( .A(n734), .B(n735), .Z(n732) );
  NANDN U845 ( .A(B[147]), .B(n736), .Z(n735) );
  NANDN U846 ( .A(A[147]), .B(n737), .Z(n736) );
  NANDN U847 ( .A(n737), .B(A[147]), .Z(n734) );
  XOR U848 ( .A(n737), .B(n738), .Z(DIFF[147]) );
  XOR U849 ( .A(B[147]), .B(A[147]), .Z(n738) );
  AND U850 ( .A(n739), .B(n740), .Z(n737) );
  NANDN U851 ( .A(B[146]), .B(n741), .Z(n740) );
  NANDN U852 ( .A(A[146]), .B(n742), .Z(n741) );
  NANDN U853 ( .A(n742), .B(A[146]), .Z(n739) );
  XOR U854 ( .A(n742), .B(n743), .Z(DIFF[146]) );
  XOR U855 ( .A(B[146]), .B(A[146]), .Z(n743) );
  AND U856 ( .A(n744), .B(n745), .Z(n742) );
  NANDN U857 ( .A(B[145]), .B(n746), .Z(n745) );
  NANDN U858 ( .A(A[145]), .B(n747), .Z(n746) );
  NANDN U859 ( .A(n747), .B(A[145]), .Z(n744) );
  XOR U860 ( .A(n747), .B(n748), .Z(DIFF[145]) );
  XOR U861 ( .A(B[145]), .B(A[145]), .Z(n748) );
  AND U862 ( .A(n749), .B(n750), .Z(n747) );
  NANDN U863 ( .A(B[144]), .B(n751), .Z(n750) );
  NANDN U864 ( .A(A[144]), .B(n752), .Z(n751) );
  NANDN U865 ( .A(n752), .B(A[144]), .Z(n749) );
  XOR U866 ( .A(n752), .B(n753), .Z(DIFF[144]) );
  XOR U867 ( .A(B[144]), .B(A[144]), .Z(n753) );
  AND U868 ( .A(n754), .B(n755), .Z(n752) );
  NANDN U869 ( .A(B[143]), .B(n756), .Z(n755) );
  NANDN U870 ( .A(A[143]), .B(n757), .Z(n756) );
  NANDN U871 ( .A(n757), .B(A[143]), .Z(n754) );
  XOR U872 ( .A(n757), .B(n758), .Z(DIFF[143]) );
  XOR U873 ( .A(B[143]), .B(A[143]), .Z(n758) );
  AND U874 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U875 ( .A(B[142]), .B(n761), .Z(n760) );
  NANDN U876 ( .A(A[142]), .B(n762), .Z(n761) );
  NANDN U877 ( .A(n762), .B(A[142]), .Z(n759) );
  XOR U878 ( .A(n762), .B(n763), .Z(DIFF[142]) );
  XOR U879 ( .A(B[142]), .B(A[142]), .Z(n763) );
  AND U880 ( .A(n764), .B(n765), .Z(n762) );
  NANDN U881 ( .A(B[141]), .B(n766), .Z(n765) );
  NANDN U882 ( .A(A[141]), .B(n767), .Z(n766) );
  NANDN U883 ( .A(n767), .B(A[141]), .Z(n764) );
  XOR U884 ( .A(n767), .B(n768), .Z(DIFF[141]) );
  XOR U885 ( .A(B[141]), .B(A[141]), .Z(n768) );
  AND U886 ( .A(n769), .B(n770), .Z(n767) );
  NANDN U887 ( .A(B[140]), .B(n771), .Z(n770) );
  NANDN U888 ( .A(A[140]), .B(n772), .Z(n771) );
  NANDN U889 ( .A(n772), .B(A[140]), .Z(n769) );
  XOR U890 ( .A(n772), .B(n773), .Z(DIFF[140]) );
  XOR U891 ( .A(B[140]), .B(A[140]), .Z(n773) );
  AND U892 ( .A(n774), .B(n775), .Z(n772) );
  NANDN U893 ( .A(B[139]), .B(n776), .Z(n775) );
  NANDN U894 ( .A(A[139]), .B(n777), .Z(n776) );
  NANDN U895 ( .A(n777), .B(A[139]), .Z(n774) );
  XOR U896 ( .A(n778), .B(n779), .Z(DIFF[13]) );
  XOR U897 ( .A(B[13]), .B(A[13]), .Z(n779) );
  XOR U898 ( .A(n777), .B(n780), .Z(DIFF[139]) );
  XOR U899 ( .A(B[139]), .B(A[139]), .Z(n780) );
  AND U900 ( .A(n781), .B(n782), .Z(n777) );
  NANDN U901 ( .A(B[138]), .B(n783), .Z(n782) );
  NANDN U902 ( .A(A[138]), .B(n784), .Z(n783) );
  NANDN U903 ( .A(n784), .B(A[138]), .Z(n781) );
  XOR U904 ( .A(n784), .B(n785), .Z(DIFF[138]) );
  XOR U905 ( .A(B[138]), .B(A[138]), .Z(n785) );
  AND U906 ( .A(n786), .B(n787), .Z(n784) );
  NANDN U907 ( .A(B[137]), .B(n788), .Z(n787) );
  NANDN U908 ( .A(A[137]), .B(n789), .Z(n788) );
  NANDN U909 ( .A(n789), .B(A[137]), .Z(n786) );
  XOR U910 ( .A(n789), .B(n790), .Z(DIFF[137]) );
  XOR U911 ( .A(B[137]), .B(A[137]), .Z(n790) );
  AND U912 ( .A(n791), .B(n792), .Z(n789) );
  NANDN U913 ( .A(B[136]), .B(n793), .Z(n792) );
  NANDN U914 ( .A(A[136]), .B(n794), .Z(n793) );
  NANDN U915 ( .A(n794), .B(A[136]), .Z(n791) );
  XOR U916 ( .A(n794), .B(n795), .Z(DIFF[136]) );
  XOR U917 ( .A(B[136]), .B(A[136]), .Z(n795) );
  AND U918 ( .A(n796), .B(n797), .Z(n794) );
  NANDN U919 ( .A(B[135]), .B(n798), .Z(n797) );
  NANDN U920 ( .A(A[135]), .B(n799), .Z(n798) );
  NANDN U921 ( .A(n799), .B(A[135]), .Z(n796) );
  XOR U922 ( .A(n799), .B(n800), .Z(DIFF[135]) );
  XOR U923 ( .A(B[135]), .B(A[135]), .Z(n800) );
  AND U924 ( .A(n801), .B(n802), .Z(n799) );
  NANDN U925 ( .A(B[134]), .B(n803), .Z(n802) );
  NANDN U926 ( .A(A[134]), .B(n804), .Z(n803) );
  NANDN U927 ( .A(n804), .B(A[134]), .Z(n801) );
  XOR U928 ( .A(n804), .B(n805), .Z(DIFF[134]) );
  XOR U929 ( .A(B[134]), .B(A[134]), .Z(n805) );
  AND U930 ( .A(n806), .B(n807), .Z(n804) );
  NANDN U931 ( .A(B[133]), .B(n808), .Z(n807) );
  NANDN U932 ( .A(A[133]), .B(n809), .Z(n808) );
  NANDN U933 ( .A(n809), .B(A[133]), .Z(n806) );
  XOR U934 ( .A(n809), .B(n810), .Z(DIFF[133]) );
  XOR U935 ( .A(B[133]), .B(A[133]), .Z(n810) );
  AND U936 ( .A(n811), .B(n812), .Z(n809) );
  NANDN U937 ( .A(B[132]), .B(n813), .Z(n812) );
  NANDN U938 ( .A(A[132]), .B(n814), .Z(n813) );
  NANDN U939 ( .A(n814), .B(A[132]), .Z(n811) );
  XOR U940 ( .A(n814), .B(n815), .Z(DIFF[132]) );
  XOR U941 ( .A(B[132]), .B(A[132]), .Z(n815) );
  AND U942 ( .A(n816), .B(n817), .Z(n814) );
  NANDN U943 ( .A(B[131]), .B(n818), .Z(n817) );
  NANDN U944 ( .A(A[131]), .B(n819), .Z(n818) );
  NANDN U945 ( .A(n819), .B(A[131]), .Z(n816) );
  XOR U946 ( .A(n819), .B(n820), .Z(DIFF[131]) );
  XOR U947 ( .A(B[131]), .B(A[131]), .Z(n820) );
  AND U948 ( .A(n821), .B(n822), .Z(n819) );
  NANDN U949 ( .A(B[130]), .B(n823), .Z(n822) );
  NANDN U950 ( .A(A[130]), .B(n824), .Z(n823) );
  NANDN U951 ( .A(n824), .B(A[130]), .Z(n821) );
  XOR U952 ( .A(n824), .B(n825), .Z(DIFF[130]) );
  XOR U953 ( .A(B[130]), .B(A[130]), .Z(n825) );
  AND U954 ( .A(n826), .B(n827), .Z(n824) );
  NANDN U955 ( .A(B[129]), .B(n828), .Z(n827) );
  NANDN U956 ( .A(A[129]), .B(n829), .Z(n828) );
  NANDN U957 ( .A(n829), .B(A[129]), .Z(n826) );
  XOR U958 ( .A(n830), .B(n831), .Z(DIFF[12]) );
  XOR U959 ( .A(B[12]), .B(A[12]), .Z(n831) );
  XOR U960 ( .A(n829), .B(n832), .Z(DIFF[129]) );
  XOR U961 ( .A(B[129]), .B(A[129]), .Z(n832) );
  AND U962 ( .A(n833), .B(n834), .Z(n829) );
  NANDN U963 ( .A(B[128]), .B(n835), .Z(n834) );
  NANDN U964 ( .A(A[128]), .B(n836), .Z(n835) );
  NANDN U965 ( .A(n836), .B(A[128]), .Z(n833) );
  XOR U966 ( .A(n836), .B(n837), .Z(DIFF[128]) );
  XOR U967 ( .A(B[128]), .B(A[128]), .Z(n837) );
  AND U968 ( .A(n838), .B(n839), .Z(n836) );
  NANDN U969 ( .A(B[127]), .B(n840), .Z(n839) );
  NANDN U970 ( .A(A[127]), .B(n841), .Z(n840) );
  NANDN U971 ( .A(n841), .B(A[127]), .Z(n838) );
  XOR U972 ( .A(n841), .B(n842), .Z(DIFF[127]) );
  XOR U973 ( .A(B[127]), .B(A[127]), .Z(n842) );
  AND U974 ( .A(n843), .B(n844), .Z(n841) );
  NANDN U975 ( .A(B[126]), .B(n845), .Z(n844) );
  NANDN U976 ( .A(A[126]), .B(n846), .Z(n845) );
  NANDN U977 ( .A(n846), .B(A[126]), .Z(n843) );
  XOR U978 ( .A(n846), .B(n847), .Z(DIFF[126]) );
  XOR U979 ( .A(B[126]), .B(A[126]), .Z(n847) );
  AND U980 ( .A(n848), .B(n849), .Z(n846) );
  NANDN U981 ( .A(B[125]), .B(n850), .Z(n849) );
  NANDN U982 ( .A(A[125]), .B(n851), .Z(n850) );
  NANDN U983 ( .A(n851), .B(A[125]), .Z(n848) );
  XOR U984 ( .A(n851), .B(n852), .Z(DIFF[125]) );
  XOR U985 ( .A(B[125]), .B(A[125]), .Z(n852) );
  AND U986 ( .A(n853), .B(n854), .Z(n851) );
  NANDN U987 ( .A(B[124]), .B(n855), .Z(n854) );
  NANDN U988 ( .A(A[124]), .B(n856), .Z(n855) );
  NANDN U989 ( .A(n856), .B(A[124]), .Z(n853) );
  XOR U990 ( .A(n856), .B(n857), .Z(DIFF[124]) );
  XOR U991 ( .A(B[124]), .B(A[124]), .Z(n857) );
  AND U992 ( .A(n858), .B(n859), .Z(n856) );
  NANDN U993 ( .A(B[123]), .B(n860), .Z(n859) );
  NANDN U994 ( .A(A[123]), .B(n861), .Z(n860) );
  NANDN U995 ( .A(n861), .B(A[123]), .Z(n858) );
  XOR U996 ( .A(n861), .B(n862), .Z(DIFF[123]) );
  XOR U997 ( .A(B[123]), .B(A[123]), .Z(n862) );
  AND U998 ( .A(n863), .B(n864), .Z(n861) );
  NANDN U999 ( .A(B[122]), .B(n865), .Z(n864) );
  NANDN U1000 ( .A(A[122]), .B(n866), .Z(n865) );
  NANDN U1001 ( .A(n866), .B(A[122]), .Z(n863) );
  XOR U1002 ( .A(n866), .B(n867), .Z(DIFF[122]) );
  XOR U1003 ( .A(B[122]), .B(A[122]), .Z(n867) );
  AND U1004 ( .A(n868), .B(n869), .Z(n866) );
  NANDN U1005 ( .A(B[121]), .B(n870), .Z(n869) );
  NANDN U1006 ( .A(A[121]), .B(n871), .Z(n870) );
  NANDN U1007 ( .A(n871), .B(A[121]), .Z(n868) );
  XOR U1008 ( .A(n871), .B(n872), .Z(DIFF[121]) );
  XOR U1009 ( .A(B[121]), .B(A[121]), .Z(n872) );
  AND U1010 ( .A(n873), .B(n874), .Z(n871) );
  NANDN U1011 ( .A(B[120]), .B(n875), .Z(n874) );
  NANDN U1012 ( .A(A[120]), .B(n876), .Z(n875) );
  NANDN U1013 ( .A(n876), .B(A[120]), .Z(n873) );
  XOR U1014 ( .A(n876), .B(n877), .Z(DIFF[120]) );
  XOR U1015 ( .A(B[120]), .B(A[120]), .Z(n877) );
  AND U1016 ( .A(n878), .B(n879), .Z(n876) );
  NANDN U1017 ( .A(B[119]), .B(n880), .Z(n879) );
  NANDN U1018 ( .A(A[119]), .B(n881), .Z(n880) );
  NANDN U1019 ( .A(n881), .B(A[119]), .Z(n878) );
  XOR U1020 ( .A(n882), .B(n883), .Z(DIFF[11]) );
  XOR U1021 ( .A(B[11]), .B(A[11]), .Z(n883) );
  XOR U1022 ( .A(n881), .B(n884), .Z(DIFF[119]) );
  XOR U1023 ( .A(B[119]), .B(A[119]), .Z(n884) );
  AND U1024 ( .A(n885), .B(n886), .Z(n881) );
  NANDN U1025 ( .A(B[118]), .B(n887), .Z(n886) );
  NANDN U1026 ( .A(A[118]), .B(n888), .Z(n887) );
  NANDN U1027 ( .A(n888), .B(A[118]), .Z(n885) );
  XOR U1028 ( .A(n888), .B(n889), .Z(DIFF[118]) );
  XOR U1029 ( .A(B[118]), .B(A[118]), .Z(n889) );
  AND U1030 ( .A(n890), .B(n891), .Z(n888) );
  NANDN U1031 ( .A(B[117]), .B(n892), .Z(n891) );
  NANDN U1032 ( .A(A[117]), .B(n893), .Z(n892) );
  NANDN U1033 ( .A(n893), .B(A[117]), .Z(n890) );
  XOR U1034 ( .A(n893), .B(n894), .Z(DIFF[117]) );
  XOR U1035 ( .A(B[117]), .B(A[117]), .Z(n894) );
  AND U1036 ( .A(n895), .B(n896), .Z(n893) );
  NANDN U1037 ( .A(B[116]), .B(n897), .Z(n896) );
  NANDN U1038 ( .A(A[116]), .B(n898), .Z(n897) );
  NANDN U1039 ( .A(n898), .B(A[116]), .Z(n895) );
  XOR U1040 ( .A(n898), .B(n899), .Z(DIFF[116]) );
  XOR U1041 ( .A(B[116]), .B(A[116]), .Z(n899) );
  AND U1042 ( .A(n900), .B(n901), .Z(n898) );
  NANDN U1043 ( .A(B[115]), .B(n902), .Z(n901) );
  NANDN U1044 ( .A(A[115]), .B(n903), .Z(n902) );
  NANDN U1045 ( .A(n903), .B(A[115]), .Z(n900) );
  XOR U1046 ( .A(n903), .B(n904), .Z(DIFF[115]) );
  XOR U1047 ( .A(B[115]), .B(A[115]), .Z(n904) );
  AND U1048 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U1049 ( .A(B[114]), .B(n907), .Z(n906) );
  NANDN U1050 ( .A(A[114]), .B(n908), .Z(n907) );
  NANDN U1051 ( .A(n908), .B(A[114]), .Z(n905) );
  XOR U1052 ( .A(n908), .B(n909), .Z(DIFF[114]) );
  XOR U1053 ( .A(B[114]), .B(A[114]), .Z(n909) );
  AND U1054 ( .A(n910), .B(n911), .Z(n908) );
  NANDN U1055 ( .A(B[113]), .B(n912), .Z(n911) );
  NANDN U1056 ( .A(A[113]), .B(n913), .Z(n912) );
  NANDN U1057 ( .A(n913), .B(A[113]), .Z(n910) );
  XOR U1058 ( .A(n913), .B(n914), .Z(DIFF[113]) );
  XOR U1059 ( .A(B[113]), .B(A[113]), .Z(n914) );
  AND U1060 ( .A(n915), .B(n916), .Z(n913) );
  NANDN U1061 ( .A(B[112]), .B(n917), .Z(n916) );
  NANDN U1062 ( .A(A[112]), .B(n918), .Z(n917) );
  NANDN U1063 ( .A(n918), .B(A[112]), .Z(n915) );
  XOR U1064 ( .A(n918), .B(n919), .Z(DIFF[112]) );
  XOR U1065 ( .A(B[112]), .B(A[112]), .Z(n919) );
  AND U1066 ( .A(n920), .B(n921), .Z(n918) );
  NANDN U1067 ( .A(B[111]), .B(n922), .Z(n921) );
  NANDN U1068 ( .A(A[111]), .B(n923), .Z(n922) );
  NANDN U1069 ( .A(n923), .B(A[111]), .Z(n920) );
  XOR U1070 ( .A(n923), .B(n924), .Z(DIFF[111]) );
  XOR U1071 ( .A(B[111]), .B(A[111]), .Z(n924) );
  AND U1072 ( .A(n925), .B(n926), .Z(n923) );
  NANDN U1073 ( .A(B[110]), .B(n927), .Z(n926) );
  NANDN U1074 ( .A(A[110]), .B(n928), .Z(n927) );
  NANDN U1075 ( .A(n928), .B(A[110]), .Z(n925) );
  XOR U1076 ( .A(n928), .B(n929), .Z(DIFF[110]) );
  XOR U1077 ( .A(B[110]), .B(A[110]), .Z(n929) );
  AND U1078 ( .A(n930), .B(n931), .Z(n928) );
  NANDN U1079 ( .A(B[109]), .B(n932), .Z(n931) );
  NANDN U1080 ( .A(A[109]), .B(n933), .Z(n932) );
  NANDN U1081 ( .A(n933), .B(A[109]), .Z(n930) );
  XOR U1082 ( .A(n934), .B(n935), .Z(DIFF[10]) );
  XOR U1083 ( .A(B[10]), .B(A[10]), .Z(n935) );
  XOR U1084 ( .A(n933), .B(n936), .Z(DIFF[109]) );
  XOR U1085 ( .A(B[109]), .B(A[109]), .Z(n936) );
  AND U1086 ( .A(n937), .B(n938), .Z(n933) );
  NANDN U1087 ( .A(B[108]), .B(n939), .Z(n938) );
  NANDN U1088 ( .A(A[108]), .B(n940), .Z(n939) );
  NANDN U1089 ( .A(n940), .B(A[108]), .Z(n937) );
  XOR U1090 ( .A(n940), .B(n941), .Z(DIFF[108]) );
  XOR U1091 ( .A(B[108]), .B(A[108]), .Z(n941) );
  AND U1092 ( .A(n942), .B(n943), .Z(n940) );
  NANDN U1093 ( .A(B[107]), .B(n944), .Z(n943) );
  NANDN U1094 ( .A(A[107]), .B(n945), .Z(n944) );
  NANDN U1095 ( .A(n945), .B(A[107]), .Z(n942) );
  XOR U1096 ( .A(n945), .B(n946), .Z(DIFF[107]) );
  XOR U1097 ( .A(B[107]), .B(A[107]), .Z(n946) );
  AND U1098 ( .A(n947), .B(n948), .Z(n945) );
  NANDN U1099 ( .A(B[106]), .B(n949), .Z(n948) );
  NANDN U1100 ( .A(A[106]), .B(n950), .Z(n949) );
  NANDN U1101 ( .A(n950), .B(A[106]), .Z(n947) );
  XOR U1102 ( .A(n950), .B(n951), .Z(DIFF[106]) );
  XOR U1103 ( .A(B[106]), .B(A[106]), .Z(n951) );
  AND U1104 ( .A(n952), .B(n953), .Z(n950) );
  NANDN U1105 ( .A(B[105]), .B(n954), .Z(n953) );
  NANDN U1106 ( .A(A[105]), .B(n955), .Z(n954) );
  NANDN U1107 ( .A(n955), .B(A[105]), .Z(n952) );
  XOR U1108 ( .A(n955), .B(n956), .Z(DIFF[105]) );
  XOR U1109 ( .A(B[105]), .B(A[105]), .Z(n956) );
  AND U1110 ( .A(n957), .B(n958), .Z(n955) );
  NANDN U1111 ( .A(B[104]), .B(n959), .Z(n958) );
  NANDN U1112 ( .A(A[104]), .B(n960), .Z(n959) );
  NANDN U1113 ( .A(n960), .B(A[104]), .Z(n957) );
  XOR U1114 ( .A(n960), .B(n961), .Z(DIFF[104]) );
  XOR U1115 ( .A(B[104]), .B(A[104]), .Z(n961) );
  AND U1116 ( .A(n962), .B(n963), .Z(n960) );
  NANDN U1117 ( .A(B[103]), .B(n964), .Z(n963) );
  NANDN U1118 ( .A(A[103]), .B(n965), .Z(n964) );
  NANDN U1119 ( .A(n965), .B(A[103]), .Z(n962) );
  XOR U1120 ( .A(n965), .B(n966), .Z(DIFF[103]) );
  XOR U1121 ( .A(B[103]), .B(A[103]), .Z(n966) );
  AND U1122 ( .A(n967), .B(n968), .Z(n965) );
  NANDN U1123 ( .A(B[102]), .B(n969), .Z(n968) );
  NANDN U1124 ( .A(A[102]), .B(n970), .Z(n969) );
  NANDN U1125 ( .A(n970), .B(A[102]), .Z(n967) );
  XOR U1126 ( .A(n970), .B(n971), .Z(DIFF[102]) );
  XOR U1127 ( .A(B[102]), .B(A[102]), .Z(n971) );
  AND U1128 ( .A(n972), .B(n973), .Z(n970) );
  NANDN U1129 ( .A(B[101]), .B(n974), .Z(n973) );
  NANDN U1130 ( .A(A[101]), .B(n975), .Z(n974) );
  NANDN U1131 ( .A(n975), .B(A[101]), .Z(n972) );
  XOR U1132 ( .A(n975), .B(n976), .Z(DIFF[101]) );
  XOR U1133 ( .A(B[101]), .B(A[101]), .Z(n976) );
  AND U1134 ( .A(n977), .B(n978), .Z(n975) );
  NANDN U1135 ( .A(B[100]), .B(n979), .Z(n978) );
  NANDN U1136 ( .A(A[100]), .B(n980), .Z(n979) );
  NANDN U1137 ( .A(n980), .B(A[100]), .Z(n977) );
  XOR U1138 ( .A(n980), .B(n981), .Z(DIFF[100]) );
  XOR U1139 ( .A(B[100]), .B(A[100]), .Z(n981) );
  AND U1140 ( .A(n982), .B(n983), .Z(n980) );
  NANDN U1141 ( .A(B[99]), .B(n984), .Z(n983) );
  OR U1142 ( .A(n5), .B(A[99]), .Z(n984) );
  NAND U1143 ( .A(A[99]), .B(n5), .Z(n982) );
  NAND U1144 ( .A(n985), .B(n986), .Z(n5) );
  NANDN U1145 ( .A(B[98]), .B(n987), .Z(n986) );
  NANDN U1146 ( .A(A[98]), .B(n7), .Z(n987) );
  NANDN U1147 ( .A(n7), .B(A[98]), .Z(n985) );
  AND U1148 ( .A(n988), .B(n989), .Z(n7) );
  NANDN U1149 ( .A(B[97]), .B(n990), .Z(n989) );
  NANDN U1150 ( .A(A[97]), .B(n9), .Z(n990) );
  NANDN U1151 ( .A(n9), .B(A[97]), .Z(n988) );
  AND U1152 ( .A(n991), .B(n992), .Z(n9) );
  NANDN U1153 ( .A(B[96]), .B(n993), .Z(n992) );
  NANDN U1154 ( .A(A[96]), .B(n11), .Z(n993) );
  NANDN U1155 ( .A(n11), .B(A[96]), .Z(n991) );
  AND U1156 ( .A(n994), .B(n995), .Z(n11) );
  NANDN U1157 ( .A(B[95]), .B(n996), .Z(n995) );
  NANDN U1158 ( .A(A[95]), .B(n13), .Z(n996) );
  NANDN U1159 ( .A(n13), .B(A[95]), .Z(n994) );
  AND U1160 ( .A(n997), .B(n998), .Z(n13) );
  NANDN U1161 ( .A(B[94]), .B(n999), .Z(n998) );
  NANDN U1162 ( .A(A[94]), .B(n15), .Z(n999) );
  NANDN U1163 ( .A(n15), .B(A[94]), .Z(n997) );
  AND U1164 ( .A(n1000), .B(n1001), .Z(n15) );
  NANDN U1165 ( .A(B[93]), .B(n1002), .Z(n1001) );
  NANDN U1166 ( .A(A[93]), .B(n17), .Z(n1002) );
  NANDN U1167 ( .A(n17), .B(A[93]), .Z(n1000) );
  AND U1168 ( .A(n1003), .B(n1004), .Z(n17) );
  NANDN U1169 ( .A(B[92]), .B(n1005), .Z(n1004) );
  NANDN U1170 ( .A(A[92]), .B(n19), .Z(n1005) );
  NANDN U1171 ( .A(n19), .B(A[92]), .Z(n1003) );
  AND U1172 ( .A(n1006), .B(n1007), .Z(n19) );
  NANDN U1173 ( .A(B[91]), .B(n1008), .Z(n1007) );
  NANDN U1174 ( .A(A[91]), .B(n21), .Z(n1008) );
  NANDN U1175 ( .A(n21), .B(A[91]), .Z(n1006) );
  AND U1176 ( .A(n1009), .B(n1010), .Z(n21) );
  NANDN U1177 ( .A(B[90]), .B(n1011), .Z(n1010) );
  NANDN U1178 ( .A(A[90]), .B(n23), .Z(n1011) );
  NANDN U1179 ( .A(n23), .B(A[90]), .Z(n1009) );
  AND U1180 ( .A(n1012), .B(n1013), .Z(n23) );
  NANDN U1181 ( .A(B[89]), .B(n1014), .Z(n1013) );
  NANDN U1182 ( .A(A[89]), .B(n27), .Z(n1014) );
  NANDN U1183 ( .A(n27), .B(A[89]), .Z(n1012) );
  AND U1184 ( .A(n1015), .B(n1016), .Z(n27) );
  NANDN U1185 ( .A(B[88]), .B(n1017), .Z(n1016) );
  NANDN U1186 ( .A(A[88]), .B(n29), .Z(n1017) );
  NANDN U1187 ( .A(n29), .B(A[88]), .Z(n1015) );
  AND U1188 ( .A(n1018), .B(n1019), .Z(n29) );
  NANDN U1189 ( .A(B[87]), .B(n1020), .Z(n1019) );
  NANDN U1190 ( .A(A[87]), .B(n31), .Z(n1020) );
  NANDN U1191 ( .A(n31), .B(A[87]), .Z(n1018) );
  AND U1192 ( .A(n1021), .B(n1022), .Z(n31) );
  NANDN U1193 ( .A(B[86]), .B(n1023), .Z(n1022) );
  NANDN U1194 ( .A(A[86]), .B(n33), .Z(n1023) );
  NANDN U1195 ( .A(n33), .B(A[86]), .Z(n1021) );
  AND U1196 ( .A(n1024), .B(n1025), .Z(n33) );
  NANDN U1197 ( .A(B[85]), .B(n1026), .Z(n1025) );
  NANDN U1198 ( .A(A[85]), .B(n35), .Z(n1026) );
  NANDN U1199 ( .A(n35), .B(A[85]), .Z(n1024) );
  AND U1200 ( .A(n1027), .B(n1028), .Z(n35) );
  NANDN U1201 ( .A(B[84]), .B(n1029), .Z(n1028) );
  NANDN U1202 ( .A(A[84]), .B(n37), .Z(n1029) );
  NANDN U1203 ( .A(n37), .B(A[84]), .Z(n1027) );
  AND U1204 ( .A(n1030), .B(n1031), .Z(n37) );
  NANDN U1205 ( .A(B[83]), .B(n1032), .Z(n1031) );
  NANDN U1206 ( .A(A[83]), .B(n39), .Z(n1032) );
  NANDN U1207 ( .A(n39), .B(A[83]), .Z(n1030) );
  AND U1208 ( .A(n1033), .B(n1034), .Z(n39) );
  NANDN U1209 ( .A(B[82]), .B(n1035), .Z(n1034) );
  NANDN U1210 ( .A(A[82]), .B(n41), .Z(n1035) );
  NANDN U1211 ( .A(n41), .B(A[82]), .Z(n1033) );
  AND U1212 ( .A(n1036), .B(n1037), .Z(n41) );
  NANDN U1213 ( .A(B[81]), .B(n1038), .Z(n1037) );
  NANDN U1214 ( .A(A[81]), .B(n43), .Z(n1038) );
  NANDN U1215 ( .A(n43), .B(A[81]), .Z(n1036) );
  AND U1216 ( .A(n1039), .B(n1040), .Z(n43) );
  NANDN U1217 ( .A(B[80]), .B(n1041), .Z(n1040) );
  NANDN U1218 ( .A(A[80]), .B(n45), .Z(n1041) );
  NANDN U1219 ( .A(n45), .B(A[80]), .Z(n1039) );
  AND U1220 ( .A(n1042), .B(n1043), .Z(n45) );
  NANDN U1221 ( .A(B[79]), .B(n1044), .Z(n1043) );
  NANDN U1222 ( .A(A[79]), .B(n49), .Z(n1044) );
  NANDN U1223 ( .A(n49), .B(A[79]), .Z(n1042) );
  AND U1224 ( .A(n1045), .B(n1046), .Z(n49) );
  NANDN U1225 ( .A(B[78]), .B(n1047), .Z(n1046) );
  NANDN U1226 ( .A(A[78]), .B(n51), .Z(n1047) );
  NANDN U1227 ( .A(n51), .B(A[78]), .Z(n1045) );
  AND U1228 ( .A(n1048), .B(n1049), .Z(n51) );
  NANDN U1229 ( .A(B[77]), .B(n1050), .Z(n1049) );
  NANDN U1230 ( .A(A[77]), .B(n53), .Z(n1050) );
  NANDN U1231 ( .A(n53), .B(A[77]), .Z(n1048) );
  AND U1232 ( .A(n1051), .B(n1052), .Z(n53) );
  NANDN U1233 ( .A(B[76]), .B(n1053), .Z(n1052) );
  NANDN U1234 ( .A(A[76]), .B(n55), .Z(n1053) );
  NANDN U1235 ( .A(n55), .B(A[76]), .Z(n1051) );
  AND U1236 ( .A(n1054), .B(n1055), .Z(n55) );
  NANDN U1237 ( .A(B[75]), .B(n1056), .Z(n1055) );
  NANDN U1238 ( .A(A[75]), .B(n57), .Z(n1056) );
  NANDN U1239 ( .A(n57), .B(A[75]), .Z(n1054) );
  AND U1240 ( .A(n1057), .B(n1058), .Z(n57) );
  NANDN U1241 ( .A(B[74]), .B(n1059), .Z(n1058) );
  NANDN U1242 ( .A(A[74]), .B(n59), .Z(n1059) );
  NANDN U1243 ( .A(n59), .B(A[74]), .Z(n1057) );
  AND U1244 ( .A(n1060), .B(n1061), .Z(n59) );
  NANDN U1245 ( .A(B[73]), .B(n1062), .Z(n1061) );
  NANDN U1246 ( .A(A[73]), .B(n61), .Z(n1062) );
  NANDN U1247 ( .A(n61), .B(A[73]), .Z(n1060) );
  AND U1248 ( .A(n1063), .B(n1064), .Z(n61) );
  NANDN U1249 ( .A(B[72]), .B(n1065), .Z(n1064) );
  NANDN U1250 ( .A(A[72]), .B(n63), .Z(n1065) );
  NANDN U1251 ( .A(n63), .B(A[72]), .Z(n1063) );
  AND U1252 ( .A(n1066), .B(n1067), .Z(n63) );
  NANDN U1253 ( .A(B[71]), .B(n1068), .Z(n1067) );
  NANDN U1254 ( .A(A[71]), .B(n65), .Z(n1068) );
  NANDN U1255 ( .A(n65), .B(A[71]), .Z(n1066) );
  AND U1256 ( .A(n1069), .B(n1070), .Z(n65) );
  NANDN U1257 ( .A(B[70]), .B(n1071), .Z(n1070) );
  NANDN U1258 ( .A(A[70]), .B(n67), .Z(n1071) );
  NANDN U1259 ( .A(n67), .B(A[70]), .Z(n1069) );
  AND U1260 ( .A(n1072), .B(n1073), .Z(n67) );
  NANDN U1261 ( .A(B[69]), .B(n1074), .Z(n1073) );
  NANDN U1262 ( .A(A[69]), .B(n71), .Z(n1074) );
  NANDN U1263 ( .A(n71), .B(A[69]), .Z(n1072) );
  AND U1264 ( .A(n1075), .B(n1076), .Z(n71) );
  NANDN U1265 ( .A(B[68]), .B(n1077), .Z(n1076) );
  NANDN U1266 ( .A(A[68]), .B(n73), .Z(n1077) );
  NANDN U1267 ( .A(n73), .B(A[68]), .Z(n1075) );
  AND U1268 ( .A(n1078), .B(n1079), .Z(n73) );
  NANDN U1269 ( .A(B[67]), .B(n1080), .Z(n1079) );
  NANDN U1270 ( .A(A[67]), .B(n75), .Z(n1080) );
  NANDN U1271 ( .A(n75), .B(A[67]), .Z(n1078) );
  AND U1272 ( .A(n1081), .B(n1082), .Z(n75) );
  NANDN U1273 ( .A(B[66]), .B(n1083), .Z(n1082) );
  NANDN U1274 ( .A(A[66]), .B(n77), .Z(n1083) );
  NANDN U1275 ( .A(n77), .B(A[66]), .Z(n1081) );
  AND U1276 ( .A(n1084), .B(n1085), .Z(n77) );
  NANDN U1277 ( .A(B[65]), .B(n1086), .Z(n1085) );
  NANDN U1278 ( .A(A[65]), .B(n79), .Z(n1086) );
  NANDN U1279 ( .A(n79), .B(A[65]), .Z(n1084) );
  AND U1280 ( .A(n1087), .B(n1088), .Z(n79) );
  NANDN U1281 ( .A(B[64]), .B(n1089), .Z(n1088) );
  NANDN U1282 ( .A(A[64]), .B(n81), .Z(n1089) );
  NANDN U1283 ( .A(n81), .B(A[64]), .Z(n1087) );
  AND U1284 ( .A(n1090), .B(n1091), .Z(n81) );
  NANDN U1285 ( .A(B[63]), .B(n1092), .Z(n1091) );
  NANDN U1286 ( .A(A[63]), .B(n83), .Z(n1092) );
  NANDN U1287 ( .A(n83), .B(A[63]), .Z(n1090) );
  AND U1288 ( .A(n1093), .B(n1094), .Z(n83) );
  NANDN U1289 ( .A(B[62]), .B(n1095), .Z(n1094) );
  NANDN U1290 ( .A(A[62]), .B(n85), .Z(n1095) );
  NANDN U1291 ( .A(n85), .B(A[62]), .Z(n1093) );
  AND U1292 ( .A(n1096), .B(n1097), .Z(n85) );
  NANDN U1293 ( .A(B[61]), .B(n1098), .Z(n1097) );
  NANDN U1294 ( .A(A[61]), .B(n87), .Z(n1098) );
  NANDN U1295 ( .A(n87), .B(A[61]), .Z(n1096) );
  AND U1296 ( .A(n1099), .B(n1100), .Z(n87) );
  NANDN U1297 ( .A(B[60]), .B(n1101), .Z(n1100) );
  NANDN U1298 ( .A(A[60]), .B(n89), .Z(n1101) );
  NANDN U1299 ( .A(n89), .B(A[60]), .Z(n1099) );
  AND U1300 ( .A(n1102), .B(n1103), .Z(n89) );
  NANDN U1301 ( .A(B[59]), .B(n1104), .Z(n1103) );
  NANDN U1302 ( .A(A[59]), .B(n93), .Z(n1104) );
  NANDN U1303 ( .A(n93), .B(A[59]), .Z(n1102) );
  AND U1304 ( .A(n1105), .B(n1106), .Z(n93) );
  NANDN U1305 ( .A(B[58]), .B(n1107), .Z(n1106) );
  NANDN U1306 ( .A(A[58]), .B(n95), .Z(n1107) );
  NANDN U1307 ( .A(n95), .B(A[58]), .Z(n1105) );
  AND U1308 ( .A(n1108), .B(n1109), .Z(n95) );
  NANDN U1309 ( .A(B[57]), .B(n1110), .Z(n1109) );
  NANDN U1310 ( .A(A[57]), .B(n97), .Z(n1110) );
  NANDN U1311 ( .A(n97), .B(A[57]), .Z(n1108) );
  AND U1312 ( .A(n1111), .B(n1112), .Z(n97) );
  NANDN U1313 ( .A(B[56]), .B(n1113), .Z(n1112) );
  NANDN U1314 ( .A(A[56]), .B(n99), .Z(n1113) );
  NANDN U1315 ( .A(n99), .B(A[56]), .Z(n1111) );
  AND U1316 ( .A(n1114), .B(n1115), .Z(n99) );
  NANDN U1317 ( .A(B[55]), .B(n1116), .Z(n1115) );
  NANDN U1318 ( .A(A[55]), .B(n101), .Z(n1116) );
  NANDN U1319 ( .A(n101), .B(A[55]), .Z(n1114) );
  AND U1320 ( .A(n1117), .B(n1118), .Z(n101) );
  NANDN U1321 ( .A(B[54]), .B(n1119), .Z(n1118) );
  NANDN U1322 ( .A(A[54]), .B(n103), .Z(n1119) );
  NANDN U1323 ( .A(n103), .B(A[54]), .Z(n1117) );
  AND U1324 ( .A(n1120), .B(n1121), .Z(n103) );
  NANDN U1325 ( .A(B[53]), .B(n1122), .Z(n1121) );
  NANDN U1326 ( .A(A[53]), .B(n105), .Z(n1122) );
  NANDN U1327 ( .A(n105), .B(A[53]), .Z(n1120) );
  AND U1328 ( .A(n1123), .B(n1124), .Z(n105) );
  NANDN U1329 ( .A(B[52]), .B(n1125), .Z(n1124) );
  NANDN U1330 ( .A(A[52]), .B(n107), .Z(n1125) );
  NANDN U1331 ( .A(n107), .B(A[52]), .Z(n1123) );
  AND U1332 ( .A(n1126), .B(n1127), .Z(n107) );
  NANDN U1333 ( .A(B[51]), .B(n1128), .Z(n1127) );
  NANDN U1334 ( .A(A[51]), .B(n109), .Z(n1128) );
  NANDN U1335 ( .A(n109), .B(A[51]), .Z(n1126) );
  AND U1336 ( .A(n1129), .B(n1130), .Z(n109) );
  NANDN U1337 ( .A(B[50]), .B(n1131), .Z(n1130) );
  NANDN U1338 ( .A(A[50]), .B(n111), .Z(n1131) );
  NANDN U1339 ( .A(n111), .B(A[50]), .Z(n1129) );
  AND U1340 ( .A(n1132), .B(n1133), .Z(n111) );
  NANDN U1341 ( .A(B[49]), .B(n1134), .Z(n1133) );
  NANDN U1342 ( .A(A[49]), .B(n115), .Z(n1134) );
  NANDN U1343 ( .A(n115), .B(A[49]), .Z(n1132) );
  AND U1344 ( .A(n1135), .B(n1136), .Z(n115) );
  NANDN U1345 ( .A(B[48]), .B(n1137), .Z(n1136) );
  NANDN U1346 ( .A(A[48]), .B(n117), .Z(n1137) );
  NANDN U1347 ( .A(n117), .B(A[48]), .Z(n1135) );
  AND U1348 ( .A(n1138), .B(n1139), .Z(n117) );
  NANDN U1349 ( .A(B[47]), .B(n1140), .Z(n1139) );
  NANDN U1350 ( .A(A[47]), .B(n119), .Z(n1140) );
  NANDN U1351 ( .A(n119), .B(A[47]), .Z(n1138) );
  AND U1352 ( .A(n1141), .B(n1142), .Z(n119) );
  NANDN U1353 ( .A(B[46]), .B(n1143), .Z(n1142) );
  NANDN U1354 ( .A(A[46]), .B(n121), .Z(n1143) );
  NANDN U1355 ( .A(n121), .B(A[46]), .Z(n1141) );
  AND U1356 ( .A(n1144), .B(n1145), .Z(n121) );
  NANDN U1357 ( .A(B[45]), .B(n1146), .Z(n1145) );
  NANDN U1358 ( .A(A[45]), .B(n123), .Z(n1146) );
  NANDN U1359 ( .A(n123), .B(A[45]), .Z(n1144) );
  AND U1360 ( .A(n1147), .B(n1148), .Z(n123) );
  NANDN U1361 ( .A(B[44]), .B(n1149), .Z(n1148) );
  NANDN U1362 ( .A(A[44]), .B(n125), .Z(n1149) );
  NANDN U1363 ( .A(n125), .B(A[44]), .Z(n1147) );
  AND U1364 ( .A(n1150), .B(n1151), .Z(n125) );
  NANDN U1365 ( .A(B[43]), .B(n1152), .Z(n1151) );
  NANDN U1366 ( .A(A[43]), .B(n127), .Z(n1152) );
  NANDN U1367 ( .A(n127), .B(A[43]), .Z(n1150) );
  AND U1368 ( .A(n1153), .B(n1154), .Z(n127) );
  NANDN U1369 ( .A(B[42]), .B(n1155), .Z(n1154) );
  NANDN U1370 ( .A(A[42]), .B(n129), .Z(n1155) );
  NANDN U1371 ( .A(n129), .B(A[42]), .Z(n1153) );
  AND U1372 ( .A(n1156), .B(n1157), .Z(n129) );
  NANDN U1373 ( .A(B[41]), .B(n1158), .Z(n1157) );
  NANDN U1374 ( .A(A[41]), .B(n131), .Z(n1158) );
  NANDN U1375 ( .A(n131), .B(A[41]), .Z(n1156) );
  AND U1376 ( .A(n1159), .B(n1160), .Z(n131) );
  NANDN U1377 ( .A(B[40]), .B(n1161), .Z(n1160) );
  NANDN U1378 ( .A(A[40]), .B(n133), .Z(n1161) );
  NANDN U1379 ( .A(n133), .B(A[40]), .Z(n1159) );
  AND U1380 ( .A(n1162), .B(n1163), .Z(n133) );
  NANDN U1381 ( .A(B[39]), .B(n1164), .Z(n1163) );
  NANDN U1382 ( .A(A[39]), .B(n137), .Z(n1164) );
  NANDN U1383 ( .A(n137), .B(A[39]), .Z(n1162) );
  AND U1384 ( .A(n1165), .B(n1166), .Z(n137) );
  NANDN U1385 ( .A(B[38]), .B(n1167), .Z(n1166) );
  NANDN U1386 ( .A(A[38]), .B(n139), .Z(n1167) );
  NANDN U1387 ( .A(n139), .B(A[38]), .Z(n1165) );
  AND U1388 ( .A(n1168), .B(n1169), .Z(n139) );
  NANDN U1389 ( .A(B[37]), .B(n1170), .Z(n1169) );
  NANDN U1390 ( .A(A[37]), .B(n141), .Z(n1170) );
  NANDN U1391 ( .A(n141), .B(A[37]), .Z(n1168) );
  AND U1392 ( .A(n1171), .B(n1172), .Z(n141) );
  NANDN U1393 ( .A(B[36]), .B(n1173), .Z(n1172) );
  NANDN U1394 ( .A(A[36]), .B(n143), .Z(n1173) );
  NANDN U1395 ( .A(n143), .B(A[36]), .Z(n1171) );
  AND U1396 ( .A(n1174), .B(n1175), .Z(n143) );
  NANDN U1397 ( .A(B[35]), .B(n1176), .Z(n1175) );
  NANDN U1398 ( .A(A[35]), .B(n145), .Z(n1176) );
  NANDN U1399 ( .A(n145), .B(A[35]), .Z(n1174) );
  AND U1400 ( .A(n1177), .B(n1178), .Z(n145) );
  NANDN U1401 ( .A(B[34]), .B(n1179), .Z(n1178) );
  NANDN U1402 ( .A(A[34]), .B(n147), .Z(n1179) );
  NANDN U1403 ( .A(n147), .B(A[34]), .Z(n1177) );
  AND U1404 ( .A(n1180), .B(n1181), .Z(n147) );
  NANDN U1405 ( .A(B[33]), .B(n1182), .Z(n1181) );
  NANDN U1406 ( .A(A[33]), .B(n149), .Z(n1182) );
  NANDN U1407 ( .A(n149), .B(A[33]), .Z(n1180) );
  AND U1408 ( .A(n1183), .B(n1184), .Z(n149) );
  NANDN U1409 ( .A(B[32]), .B(n1185), .Z(n1184) );
  NANDN U1410 ( .A(A[32]), .B(n151), .Z(n1185) );
  NANDN U1411 ( .A(n151), .B(A[32]), .Z(n1183) );
  AND U1412 ( .A(n1186), .B(n1187), .Z(n151) );
  NANDN U1413 ( .A(B[31]), .B(n1188), .Z(n1187) );
  NANDN U1414 ( .A(A[31]), .B(n153), .Z(n1188) );
  NANDN U1415 ( .A(n153), .B(A[31]), .Z(n1186) );
  AND U1416 ( .A(n1189), .B(n1190), .Z(n153) );
  NANDN U1417 ( .A(B[30]), .B(n1191), .Z(n1190) );
  NANDN U1418 ( .A(A[30]), .B(n155), .Z(n1191) );
  NANDN U1419 ( .A(n155), .B(A[30]), .Z(n1189) );
  AND U1420 ( .A(n1192), .B(n1193), .Z(n155) );
  NANDN U1421 ( .A(B[29]), .B(n1194), .Z(n1193) );
  NANDN U1422 ( .A(A[29]), .B(n159), .Z(n1194) );
  NANDN U1423 ( .A(n159), .B(A[29]), .Z(n1192) );
  AND U1424 ( .A(n1195), .B(n1196), .Z(n159) );
  NANDN U1425 ( .A(B[28]), .B(n1197), .Z(n1196) );
  NANDN U1426 ( .A(A[28]), .B(n161), .Z(n1197) );
  NANDN U1427 ( .A(n161), .B(A[28]), .Z(n1195) );
  AND U1428 ( .A(n1198), .B(n1199), .Z(n161) );
  NANDN U1429 ( .A(B[27]), .B(n1200), .Z(n1199) );
  NANDN U1430 ( .A(A[27]), .B(n163), .Z(n1200) );
  NANDN U1431 ( .A(n163), .B(A[27]), .Z(n1198) );
  AND U1432 ( .A(n1201), .B(n1202), .Z(n163) );
  NANDN U1433 ( .A(B[26]), .B(n1203), .Z(n1202) );
  NANDN U1434 ( .A(A[26]), .B(n165), .Z(n1203) );
  NANDN U1435 ( .A(n165), .B(A[26]), .Z(n1201) );
  AND U1436 ( .A(n1204), .B(n1205), .Z(n165) );
  NANDN U1437 ( .A(B[25]), .B(n1206), .Z(n1205) );
  NANDN U1438 ( .A(A[25]), .B(n167), .Z(n1206) );
  NANDN U1439 ( .A(n167), .B(A[25]), .Z(n1204) );
  AND U1440 ( .A(n1207), .B(n1208), .Z(n167) );
  NANDN U1441 ( .A(B[24]), .B(n1209), .Z(n1208) );
  NANDN U1442 ( .A(A[24]), .B(n205), .Z(n1209) );
  NANDN U1443 ( .A(n205), .B(A[24]), .Z(n1207) );
  AND U1444 ( .A(n1210), .B(n1211), .Z(n205) );
  NANDN U1445 ( .A(B[23]), .B(n1212), .Z(n1211) );
  NANDN U1446 ( .A(A[23]), .B(n257), .Z(n1212) );
  NANDN U1447 ( .A(n257), .B(A[23]), .Z(n1210) );
  AND U1448 ( .A(n1213), .B(n1214), .Z(n257) );
  NANDN U1449 ( .A(B[22]), .B(n1215), .Z(n1214) );
  NANDN U1450 ( .A(A[22]), .B(n309), .Z(n1215) );
  NANDN U1451 ( .A(n309), .B(A[22]), .Z(n1213) );
  AND U1452 ( .A(n1216), .B(n1217), .Z(n309) );
  NANDN U1453 ( .A(B[21]), .B(n1218), .Z(n1217) );
  NANDN U1454 ( .A(A[21]), .B(n361), .Z(n1218) );
  NANDN U1455 ( .A(n361), .B(A[21]), .Z(n1216) );
  AND U1456 ( .A(n1219), .B(n1220), .Z(n361) );
  NANDN U1457 ( .A(B[20]), .B(n1221), .Z(n1220) );
  NANDN U1458 ( .A(A[20]), .B(n413), .Z(n1221) );
  NANDN U1459 ( .A(n413), .B(A[20]), .Z(n1219) );
  AND U1460 ( .A(n1222), .B(n1223), .Z(n413) );
  NANDN U1461 ( .A(B[19]), .B(n1224), .Z(n1223) );
  NANDN U1462 ( .A(A[19]), .B(n466), .Z(n1224) );
  NANDN U1463 ( .A(n466), .B(A[19]), .Z(n1222) );
  AND U1464 ( .A(n1225), .B(n1226), .Z(n466) );
  NANDN U1465 ( .A(B[18]), .B(n1227), .Z(n1226) );
  NANDN U1466 ( .A(A[18]), .B(n518), .Z(n1227) );
  NANDN U1467 ( .A(n518), .B(A[18]), .Z(n1225) );
  AND U1468 ( .A(n1228), .B(n1229), .Z(n518) );
  NANDN U1469 ( .A(B[17]), .B(n1230), .Z(n1229) );
  NANDN U1470 ( .A(A[17]), .B(n570), .Z(n1230) );
  NANDN U1471 ( .A(n570), .B(A[17]), .Z(n1228) );
  AND U1472 ( .A(n1231), .B(n1232), .Z(n570) );
  NANDN U1473 ( .A(B[16]), .B(n1233), .Z(n1232) );
  NANDN U1474 ( .A(A[16]), .B(n622), .Z(n1233) );
  NANDN U1475 ( .A(n622), .B(A[16]), .Z(n1231) );
  AND U1476 ( .A(n1234), .B(n1235), .Z(n622) );
  NANDN U1477 ( .A(B[15]), .B(n1236), .Z(n1235) );
  NANDN U1478 ( .A(A[15]), .B(n674), .Z(n1236) );
  NANDN U1479 ( .A(n674), .B(A[15]), .Z(n1234) );
  AND U1480 ( .A(n1237), .B(n1238), .Z(n674) );
  NANDN U1481 ( .A(B[14]), .B(n1239), .Z(n1238) );
  NANDN U1482 ( .A(A[14]), .B(n726), .Z(n1239) );
  NANDN U1483 ( .A(n726), .B(A[14]), .Z(n1237) );
  AND U1484 ( .A(n1240), .B(n1241), .Z(n726) );
  NANDN U1485 ( .A(B[13]), .B(n1242), .Z(n1241) );
  NANDN U1486 ( .A(A[13]), .B(n778), .Z(n1242) );
  NANDN U1487 ( .A(n778), .B(A[13]), .Z(n1240) );
  AND U1488 ( .A(n1243), .B(n1244), .Z(n778) );
  NANDN U1489 ( .A(B[12]), .B(n1245), .Z(n1244) );
  NANDN U1490 ( .A(A[12]), .B(n830), .Z(n1245) );
  NANDN U1491 ( .A(n830), .B(A[12]), .Z(n1243) );
  AND U1492 ( .A(n1246), .B(n1247), .Z(n830) );
  NANDN U1493 ( .A(B[11]), .B(n1248), .Z(n1247) );
  NANDN U1494 ( .A(A[11]), .B(n882), .Z(n1248) );
  NANDN U1495 ( .A(n882), .B(A[11]), .Z(n1246) );
  AND U1496 ( .A(n1249), .B(n1250), .Z(n882) );
  NANDN U1497 ( .A(B[10]), .B(n1251), .Z(n1250) );
  NANDN U1498 ( .A(A[10]), .B(n934), .Z(n1251) );
  NANDN U1499 ( .A(n934), .B(A[10]), .Z(n1249) );
  AND U1500 ( .A(n1252), .B(n1253), .Z(n934) );
  NANDN U1501 ( .A(B[9]), .B(n1254), .Z(n1253) );
  OR U1502 ( .A(n3), .B(A[9]), .Z(n1254) );
  NAND U1503 ( .A(A[9]), .B(n3), .Z(n1252) );
  NAND U1504 ( .A(n1255), .B(n1256), .Z(n3) );
  NANDN U1505 ( .A(B[8]), .B(n1257), .Z(n1256) );
  NANDN U1506 ( .A(A[8]), .B(n25), .Z(n1257) );
  NANDN U1507 ( .A(n25), .B(A[8]), .Z(n1255) );
  AND U1508 ( .A(n1258), .B(n1259), .Z(n25) );
  NANDN U1509 ( .A(B[7]), .B(n1260), .Z(n1259) );
  NANDN U1510 ( .A(A[7]), .B(n47), .Z(n1260) );
  NANDN U1511 ( .A(n47), .B(A[7]), .Z(n1258) );
  AND U1512 ( .A(n1261), .B(n1262), .Z(n47) );
  NANDN U1513 ( .A(B[6]), .B(n1263), .Z(n1262) );
  NANDN U1514 ( .A(A[6]), .B(n69), .Z(n1263) );
  NANDN U1515 ( .A(n69), .B(A[6]), .Z(n1261) );
  AND U1516 ( .A(n1264), .B(n1265), .Z(n69) );
  NANDN U1517 ( .A(B[5]), .B(n1266), .Z(n1265) );
  NANDN U1518 ( .A(A[5]), .B(n91), .Z(n1266) );
  NANDN U1519 ( .A(n91), .B(A[5]), .Z(n1264) );
  AND U1520 ( .A(n1267), .B(n1268), .Z(n91) );
  NANDN U1521 ( .A(B[4]), .B(n1269), .Z(n1268) );
  NANDN U1522 ( .A(A[4]), .B(n113), .Z(n1269) );
  NANDN U1523 ( .A(n113), .B(A[4]), .Z(n1267) );
  AND U1524 ( .A(n1270), .B(n1271), .Z(n113) );
  NANDN U1525 ( .A(B[3]), .B(n1272), .Z(n1271) );
  NANDN U1526 ( .A(A[3]), .B(n135), .Z(n1272) );
  NANDN U1527 ( .A(n135), .B(A[3]), .Z(n1270) );
  AND U1528 ( .A(n1273), .B(n1274), .Z(n135) );
  NANDN U1529 ( .A(B[2]), .B(n1275), .Z(n1274) );
  NANDN U1530 ( .A(A[2]), .B(n157), .Z(n1275) );
  NANDN U1531 ( .A(n157), .B(A[2]), .Z(n1273) );
  AND U1532 ( .A(n1276), .B(n1277), .Z(n157) );
  NANDN U1533 ( .A(B[1]), .B(n1278), .Z(n1277) );
  NAND U1534 ( .A(n1), .B(n2), .Z(n1278) );
  NAND U1535 ( .A(A[1]), .B(n1279), .Z(n1276) );
  NAND U1536 ( .A(n1279), .B(n1280), .Z(DIFF[0]) );
  NANDN U1537 ( .A(B[0]), .B(A[0]), .Z(n1280) );
  NANDN U1538 ( .A(A[0]), .B(B[0]), .Z(n1279) );
endmodule


module modmult_step_N256_3_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [255:0] A;
  input [0:0] B;
  output [256:0] PRODUCT;
  input TC;


  AND U2 ( .A(A[255]), .B(B[0]), .Z(PRODUCT[255]) );
  AND U3 ( .A(A[254]), .B(B[0]), .Z(PRODUCT[254]) );
  AND U4 ( .A(A[253]), .B(B[0]), .Z(PRODUCT[253]) );
  AND U5 ( .A(A[252]), .B(B[0]), .Z(PRODUCT[252]) );
  AND U6 ( .A(A[251]), .B(B[0]), .Z(PRODUCT[251]) );
  AND U7 ( .A(A[250]), .B(B[0]), .Z(PRODUCT[250]) );
  AND U8 ( .A(A[249]), .B(B[0]), .Z(PRODUCT[249]) );
  AND U9 ( .A(A[248]), .B(B[0]), .Z(PRODUCT[248]) );
  AND U10 ( .A(A[247]), .B(B[0]), .Z(PRODUCT[247]) );
  AND U11 ( .A(A[246]), .B(B[0]), .Z(PRODUCT[246]) );
  AND U12 ( .A(A[245]), .B(B[0]), .Z(PRODUCT[245]) );
  AND U13 ( .A(A[244]), .B(B[0]), .Z(PRODUCT[244]) );
  AND U14 ( .A(A[243]), .B(B[0]), .Z(PRODUCT[243]) );
  AND U15 ( .A(A[242]), .B(B[0]), .Z(PRODUCT[242]) );
  AND U16 ( .A(A[241]), .B(B[0]), .Z(PRODUCT[241]) );
  AND U17 ( .A(A[240]), .B(B[0]), .Z(PRODUCT[240]) );
  AND U18 ( .A(A[239]), .B(B[0]), .Z(PRODUCT[239]) );
  AND U19 ( .A(A[238]), .B(B[0]), .Z(PRODUCT[238]) );
  AND U20 ( .A(A[237]), .B(B[0]), .Z(PRODUCT[237]) );
  AND U21 ( .A(A[236]), .B(B[0]), .Z(PRODUCT[236]) );
  AND U22 ( .A(A[235]), .B(B[0]), .Z(PRODUCT[235]) );
  AND U23 ( .A(A[234]), .B(B[0]), .Z(PRODUCT[234]) );
  AND U24 ( .A(A[233]), .B(B[0]), .Z(PRODUCT[233]) );
  AND U25 ( .A(A[232]), .B(B[0]), .Z(PRODUCT[232]) );
  AND U26 ( .A(A[231]), .B(B[0]), .Z(PRODUCT[231]) );
  AND U27 ( .A(A[230]), .B(B[0]), .Z(PRODUCT[230]) );
  AND U28 ( .A(A[229]), .B(B[0]), .Z(PRODUCT[229]) );
  AND U29 ( .A(A[228]), .B(B[0]), .Z(PRODUCT[228]) );
  AND U30 ( .A(A[227]), .B(B[0]), .Z(PRODUCT[227]) );
  AND U31 ( .A(A[226]), .B(B[0]), .Z(PRODUCT[226]) );
  AND U32 ( .A(A[225]), .B(B[0]), .Z(PRODUCT[225]) );
  AND U33 ( .A(A[224]), .B(B[0]), .Z(PRODUCT[224]) );
  AND U34 ( .A(A[223]), .B(B[0]), .Z(PRODUCT[223]) );
  AND U35 ( .A(A[222]), .B(B[0]), .Z(PRODUCT[222]) );
  AND U36 ( .A(A[221]), .B(B[0]), .Z(PRODUCT[221]) );
  AND U37 ( .A(A[220]), .B(B[0]), .Z(PRODUCT[220]) );
  AND U38 ( .A(A[219]), .B(B[0]), .Z(PRODUCT[219]) );
  AND U39 ( .A(A[218]), .B(B[0]), .Z(PRODUCT[218]) );
  AND U40 ( .A(A[217]), .B(B[0]), .Z(PRODUCT[217]) );
  AND U41 ( .A(A[216]), .B(B[0]), .Z(PRODUCT[216]) );
  AND U42 ( .A(A[215]), .B(B[0]), .Z(PRODUCT[215]) );
  AND U43 ( .A(A[214]), .B(B[0]), .Z(PRODUCT[214]) );
  AND U44 ( .A(A[213]), .B(B[0]), .Z(PRODUCT[213]) );
  AND U45 ( .A(A[212]), .B(B[0]), .Z(PRODUCT[212]) );
  AND U46 ( .A(A[211]), .B(B[0]), .Z(PRODUCT[211]) );
  AND U47 ( .A(A[210]), .B(B[0]), .Z(PRODUCT[210]) );
  AND U48 ( .A(A[209]), .B(B[0]), .Z(PRODUCT[209]) );
  AND U49 ( .A(A[208]), .B(B[0]), .Z(PRODUCT[208]) );
  AND U50 ( .A(A[207]), .B(B[0]), .Z(PRODUCT[207]) );
  AND U51 ( .A(A[206]), .B(B[0]), .Z(PRODUCT[206]) );
  AND U52 ( .A(A[205]), .B(B[0]), .Z(PRODUCT[205]) );
  AND U53 ( .A(A[204]), .B(B[0]), .Z(PRODUCT[204]) );
  AND U54 ( .A(A[203]), .B(B[0]), .Z(PRODUCT[203]) );
  AND U55 ( .A(A[202]), .B(B[0]), .Z(PRODUCT[202]) );
  AND U56 ( .A(A[201]), .B(B[0]), .Z(PRODUCT[201]) );
  AND U57 ( .A(A[200]), .B(B[0]), .Z(PRODUCT[200]) );
  AND U58 ( .A(A[199]), .B(B[0]), .Z(PRODUCT[199]) );
  AND U59 ( .A(A[198]), .B(B[0]), .Z(PRODUCT[198]) );
  AND U60 ( .A(A[197]), .B(B[0]), .Z(PRODUCT[197]) );
  AND U61 ( .A(A[196]), .B(B[0]), .Z(PRODUCT[196]) );
  AND U62 ( .A(A[195]), .B(B[0]), .Z(PRODUCT[195]) );
  AND U63 ( .A(A[194]), .B(B[0]), .Z(PRODUCT[194]) );
  AND U64 ( .A(A[193]), .B(B[0]), .Z(PRODUCT[193]) );
  AND U65 ( .A(A[192]), .B(B[0]), .Z(PRODUCT[192]) );
  AND U66 ( .A(A[191]), .B(B[0]), .Z(PRODUCT[191]) );
  AND U67 ( .A(A[190]), .B(B[0]), .Z(PRODUCT[190]) );
  AND U68 ( .A(A[189]), .B(B[0]), .Z(PRODUCT[189]) );
  AND U69 ( .A(A[188]), .B(B[0]), .Z(PRODUCT[188]) );
  AND U70 ( .A(A[187]), .B(B[0]), .Z(PRODUCT[187]) );
  AND U71 ( .A(A[186]), .B(B[0]), .Z(PRODUCT[186]) );
  AND U72 ( .A(A[185]), .B(B[0]), .Z(PRODUCT[185]) );
  AND U73 ( .A(A[184]), .B(B[0]), .Z(PRODUCT[184]) );
  AND U74 ( .A(A[183]), .B(B[0]), .Z(PRODUCT[183]) );
  AND U75 ( .A(A[182]), .B(B[0]), .Z(PRODUCT[182]) );
  AND U76 ( .A(A[181]), .B(B[0]), .Z(PRODUCT[181]) );
  AND U77 ( .A(A[180]), .B(B[0]), .Z(PRODUCT[180]) );
  AND U78 ( .A(A[179]), .B(B[0]), .Z(PRODUCT[179]) );
  AND U79 ( .A(A[178]), .B(B[0]), .Z(PRODUCT[178]) );
  AND U80 ( .A(A[177]), .B(B[0]), .Z(PRODUCT[177]) );
  AND U81 ( .A(A[176]), .B(B[0]), .Z(PRODUCT[176]) );
  AND U82 ( .A(A[175]), .B(B[0]), .Z(PRODUCT[175]) );
  AND U83 ( .A(A[174]), .B(B[0]), .Z(PRODUCT[174]) );
  AND U84 ( .A(A[173]), .B(B[0]), .Z(PRODUCT[173]) );
  AND U85 ( .A(A[172]), .B(B[0]), .Z(PRODUCT[172]) );
  AND U86 ( .A(A[171]), .B(B[0]), .Z(PRODUCT[171]) );
  AND U87 ( .A(A[170]), .B(B[0]), .Z(PRODUCT[170]) );
  AND U88 ( .A(A[169]), .B(B[0]), .Z(PRODUCT[169]) );
  AND U89 ( .A(A[168]), .B(B[0]), .Z(PRODUCT[168]) );
  AND U90 ( .A(A[167]), .B(B[0]), .Z(PRODUCT[167]) );
  AND U91 ( .A(A[166]), .B(B[0]), .Z(PRODUCT[166]) );
  AND U92 ( .A(A[165]), .B(B[0]), .Z(PRODUCT[165]) );
  AND U93 ( .A(A[164]), .B(B[0]), .Z(PRODUCT[164]) );
  AND U94 ( .A(A[163]), .B(B[0]), .Z(PRODUCT[163]) );
  AND U95 ( .A(A[162]), .B(B[0]), .Z(PRODUCT[162]) );
  AND U96 ( .A(A[161]), .B(B[0]), .Z(PRODUCT[161]) );
  AND U97 ( .A(A[160]), .B(B[0]), .Z(PRODUCT[160]) );
  AND U98 ( .A(A[159]), .B(B[0]), .Z(PRODUCT[159]) );
  AND U99 ( .A(A[158]), .B(B[0]), .Z(PRODUCT[158]) );
  AND U100 ( .A(A[157]), .B(B[0]), .Z(PRODUCT[157]) );
  AND U101 ( .A(A[156]), .B(B[0]), .Z(PRODUCT[156]) );
  AND U102 ( .A(A[155]), .B(B[0]), .Z(PRODUCT[155]) );
  AND U103 ( .A(A[154]), .B(B[0]), .Z(PRODUCT[154]) );
  AND U104 ( .A(A[153]), .B(B[0]), .Z(PRODUCT[153]) );
  AND U105 ( .A(A[152]), .B(B[0]), .Z(PRODUCT[152]) );
  AND U106 ( .A(A[151]), .B(B[0]), .Z(PRODUCT[151]) );
  AND U107 ( .A(A[150]), .B(B[0]), .Z(PRODUCT[150]) );
  AND U108 ( .A(A[149]), .B(B[0]), .Z(PRODUCT[149]) );
  AND U109 ( .A(A[148]), .B(B[0]), .Z(PRODUCT[148]) );
  AND U110 ( .A(A[147]), .B(B[0]), .Z(PRODUCT[147]) );
  AND U111 ( .A(A[146]), .B(B[0]), .Z(PRODUCT[146]) );
  AND U112 ( .A(A[145]), .B(B[0]), .Z(PRODUCT[145]) );
  AND U113 ( .A(A[144]), .B(B[0]), .Z(PRODUCT[144]) );
  AND U114 ( .A(A[143]), .B(B[0]), .Z(PRODUCT[143]) );
  AND U115 ( .A(A[142]), .B(B[0]), .Z(PRODUCT[142]) );
  AND U116 ( .A(A[141]), .B(B[0]), .Z(PRODUCT[141]) );
  AND U117 ( .A(A[140]), .B(B[0]), .Z(PRODUCT[140]) );
  AND U118 ( .A(A[139]), .B(B[0]), .Z(PRODUCT[139]) );
  AND U119 ( .A(A[138]), .B(B[0]), .Z(PRODUCT[138]) );
  AND U120 ( .A(A[137]), .B(B[0]), .Z(PRODUCT[137]) );
  AND U121 ( .A(A[136]), .B(B[0]), .Z(PRODUCT[136]) );
  AND U122 ( .A(A[135]), .B(B[0]), .Z(PRODUCT[135]) );
  AND U123 ( .A(A[134]), .B(B[0]), .Z(PRODUCT[134]) );
  AND U124 ( .A(A[133]), .B(B[0]), .Z(PRODUCT[133]) );
  AND U125 ( .A(A[132]), .B(B[0]), .Z(PRODUCT[132]) );
  AND U126 ( .A(A[131]), .B(B[0]), .Z(PRODUCT[131]) );
  AND U127 ( .A(A[130]), .B(B[0]), .Z(PRODUCT[130]) );
  AND U128 ( .A(A[129]), .B(B[0]), .Z(PRODUCT[129]) );
  AND U129 ( .A(A[128]), .B(B[0]), .Z(PRODUCT[128]) );
  AND U130 ( .A(A[127]), .B(B[0]), .Z(PRODUCT[127]) );
  AND U131 ( .A(A[126]), .B(B[0]), .Z(PRODUCT[126]) );
  AND U132 ( .A(A[125]), .B(B[0]), .Z(PRODUCT[125]) );
  AND U133 ( .A(A[124]), .B(B[0]), .Z(PRODUCT[124]) );
  AND U134 ( .A(A[123]), .B(B[0]), .Z(PRODUCT[123]) );
  AND U135 ( .A(A[122]), .B(B[0]), .Z(PRODUCT[122]) );
  AND U136 ( .A(A[121]), .B(B[0]), .Z(PRODUCT[121]) );
  AND U137 ( .A(A[120]), .B(B[0]), .Z(PRODUCT[120]) );
  AND U138 ( .A(A[119]), .B(B[0]), .Z(PRODUCT[119]) );
  AND U139 ( .A(A[118]), .B(B[0]), .Z(PRODUCT[118]) );
  AND U140 ( .A(A[117]), .B(B[0]), .Z(PRODUCT[117]) );
  AND U141 ( .A(A[116]), .B(B[0]), .Z(PRODUCT[116]) );
  AND U142 ( .A(A[115]), .B(B[0]), .Z(PRODUCT[115]) );
  AND U143 ( .A(A[114]), .B(B[0]), .Z(PRODUCT[114]) );
  AND U144 ( .A(A[113]), .B(B[0]), .Z(PRODUCT[113]) );
  AND U145 ( .A(A[112]), .B(B[0]), .Z(PRODUCT[112]) );
  AND U146 ( .A(A[111]), .B(B[0]), .Z(PRODUCT[111]) );
  AND U147 ( .A(A[110]), .B(B[0]), .Z(PRODUCT[110]) );
  AND U148 ( .A(A[109]), .B(B[0]), .Z(PRODUCT[109]) );
  AND U149 ( .A(A[108]), .B(B[0]), .Z(PRODUCT[108]) );
  AND U150 ( .A(A[107]), .B(B[0]), .Z(PRODUCT[107]) );
  AND U151 ( .A(A[106]), .B(B[0]), .Z(PRODUCT[106]) );
  AND U152 ( .A(A[105]), .B(B[0]), .Z(PRODUCT[105]) );
  AND U153 ( .A(A[104]), .B(B[0]), .Z(PRODUCT[104]) );
  AND U154 ( .A(A[103]), .B(B[0]), .Z(PRODUCT[103]) );
  AND U155 ( .A(A[102]), .B(B[0]), .Z(PRODUCT[102]) );
  AND U156 ( .A(A[101]), .B(B[0]), .Z(PRODUCT[101]) );
  AND U157 ( .A(A[100]), .B(B[0]), .Z(PRODUCT[100]) );
  AND U158 ( .A(A[99]), .B(B[0]), .Z(PRODUCT[99]) );
  AND U159 ( .A(A[98]), .B(B[0]), .Z(PRODUCT[98]) );
  AND U160 ( .A(A[97]), .B(B[0]), .Z(PRODUCT[97]) );
  AND U161 ( .A(A[96]), .B(B[0]), .Z(PRODUCT[96]) );
  AND U162 ( .A(A[95]), .B(B[0]), .Z(PRODUCT[95]) );
  AND U163 ( .A(A[94]), .B(B[0]), .Z(PRODUCT[94]) );
  AND U164 ( .A(A[93]), .B(B[0]), .Z(PRODUCT[93]) );
  AND U165 ( .A(A[92]), .B(B[0]), .Z(PRODUCT[92]) );
  AND U166 ( .A(A[91]), .B(B[0]), .Z(PRODUCT[91]) );
  AND U167 ( .A(A[90]), .B(B[0]), .Z(PRODUCT[90]) );
  AND U168 ( .A(A[89]), .B(B[0]), .Z(PRODUCT[89]) );
  AND U169 ( .A(A[88]), .B(B[0]), .Z(PRODUCT[88]) );
  AND U170 ( .A(A[87]), .B(B[0]), .Z(PRODUCT[87]) );
  AND U171 ( .A(A[86]), .B(B[0]), .Z(PRODUCT[86]) );
  AND U172 ( .A(A[85]), .B(B[0]), .Z(PRODUCT[85]) );
  AND U173 ( .A(A[84]), .B(B[0]), .Z(PRODUCT[84]) );
  AND U174 ( .A(A[83]), .B(B[0]), .Z(PRODUCT[83]) );
  AND U175 ( .A(A[82]), .B(B[0]), .Z(PRODUCT[82]) );
  AND U176 ( .A(A[81]), .B(B[0]), .Z(PRODUCT[81]) );
  AND U177 ( .A(A[80]), .B(B[0]), .Z(PRODUCT[80]) );
  AND U178 ( .A(A[79]), .B(B[0]), .Z(PRODUCT[79]) );
  AND U179 ( .A(A[78]), .B(B[0]), .Z(PRODUCT[78]) );
  AND U180 ( .A(A[77]), .B(B[0]), .Z(PRODUCT[77]) );
  AND U181 ( .A(A[76]), .B(B[0]), .Z(PRODUCT[76]) );
  AND U182 ( .A(A[75]), .B(B[0]), .Z(PRODUCT[75]) );
  AND U183 ( .A(A[74]), .B(B[0]), .Z(PRODUCT[74]) );
  AND U184 ( .A(A[73]), .B(B[0]), .Z(PRODUCT[73]) );
  AND U185 ( .A(A[72]), .B(B[0]), .Z(PRODUCT[72]) );
  AND U186 ( .A(A[71]), .B(B[0]), .Z(PRODUCT[71]) );
  AND U187 ( .A(A[70]), .B(B[0]), .Z(PRODUCT[70]) );
  AND U188 ( .A(A[69]), .B(B[0]), .Z(PRODUCT[69]) );
  AND U189 ( .A(A[68]), .B(B[0]), .Z(PRODUCT[68]) );
  AND U190 ( .A(A[67]), .B(B[0]), .Z(PRODUCT[67]) );
  AND U191 ( .A(A[66]), .B(B[0]), .Z(PRODUCT[66]) );
  AND U192 ( .A(A[65]), .B(B[0]), .Z(PRODUCT[65]) );
  AND U193 ( .A(A[64]), .B(B[0]), .Z(PRODUCT[64]) );
  AND U194 ( .A(A[63]), .B(B[0]), .Z(PRODUCT[63]) );
  AND U195 ( .A(A[62]), .B(B[0]), .Z(PRODUCT[62]) );
  AND U196 ( .A(A[61]), .B(B[0]), .Z(PRODUCT[61]) );
  AND U197 ( .A(A[60]), .B(B[0]), .Z(PRODUCT[60]) );
  AND U198 ( .A(A[59]), .B(B[0]), .Z(PRODUCT[59]) );
  AND U199 ( .A(A[58]), .B(B[0]), .Z(PRODUCT[58]) );
  AND U200 ( .A(A[57]), .B(B[0]), .Z(PRODUCT[57]) );
  AND U201 ( .A(A[56]), .B(B[0]), .Z(PRODUCT[56]) );
  AND U202 ( .A(A[55]), .B(B[0]), .Z(PRODUCT[55]) );
  AND U203 ( .A(A[54]), .B(B[0]), .Z(PRODUCT[54]) );
  AND U204 ( .A(A[53]), .B(B[0]), .Z(PRODUCT[53]) );
  AND U205 ( .A(A[52]), .B(B[0]), .Z(PRODUCT[52]) );
  AND U206 ( .A(A[51]), .B(B[0]), .Z(PRODUCT[51]) );
  AND U207 ( .A(A[50]), .B(B[0]), .Z(PRODUCT[50]) );
  AND U208 ( .A(A[49]), .B(B[0]), .Z(PRODUCT[49]) );
  AND U209 ( .A(A[48]), .B(B[0]), .Z(PRODUCT[48]) );
  AND U210 ( .A(A[47]), .B(B[0]), .Z(PRODUCT[47]) );
  AND U211 ( .A(A[46]), .B(B[0]), .Z(PRODUCT[46]) );
  AND U212 ( .A(A[45]), .B(B[0]), .Z(PRODUCT[45]) );
  AND U213 ( .A(A[44]), .B(B[0]), .Z(PRODUCT[44]) );
  AND U214 ( .A(A[43]), .B(B[0]), .Z(PRODUCT[43]) );
  AND U215 ( .A(A[42]), .B(B[0]), .Z(PRODUCT[42]) );
  AND U216 ( .A(A[41]), .B(B[0]), .Z(PRODUCT[41]) );
  AND U217 ( .A(A[40]), .B(B[0]), .Z(PRODUCT[40]) );
  AND U218 ( .A(A[39]), .B(B[0]), .Z(PRODUCT[39]) );
  AND U219 ( .A(A[38]), .B(B[0]), .Z(PRODUCT[38]) );
  AND U220 ( .A(A[37]), .B(B[0]), .Z(PRODUCT[37]) );
  AND U221 ( .A(A[36]), .B(B[0]), .Z(PRODUCT[36]) );
  AND U222 ( .A(A[35]), .B(B[0]), .Z(PRODUCT[35]) );
  AND U223 ( .A(A[34]), .B(B[0]), .Z(PRODUCT[34]) );
  AND U224 ( .A(A[33]), .B(B[0]), .Z(PRODUCT[33]) );
  AND U225 ( .A(A[32]), .B(B[0]), .Z(PRODUCT[32]) );
  AND U226 ( .A(A[31]), .B(B[0]), .Z(PRODUCT[31]) );
  AND U227 ( .A(A[30]), .B(B[0]), .Z(PRODUCT[30]) );
  AND U228 ( .A(A[29]), .B(B[0]), .Z(PRODUCT[29]) );
  AND U229 ( .A(A[28]), .B(B[0]), .Z(PRODUCT[28]) );
  AND U230 ( .A(A[27]), .B(B[0]), .Z(PRODUCT[27]) );
  AND U231 ( .A(A[26]), .B(B[0]), .Z(PRODUCT[26]) );
  AND U232 ( .A(A[25]), .B(B[0]), .Z(PRODUCT[25]) );
  AND U233 ( .A(A[24]), .B(B[0]), .Z(PRODUCT[24]) );
  AND U234 ( .A(A[23]), .B(B[0]), .Z(PRODUCT[23]) );
  AND U235 ( .A(A[22]), .B(B[0]), .Z(PRODUCT[22]) );
  AND U236 ( .A(A[21]), .B(B[0]), .Z(PRODUCT[21]) );
  AND U237 ( .A(A[20]), .B(B[0]), .Z(PRODUCT[20]) );
  AND U238 ( .A(A[19]), .B(B[0]), .Z(PRODUCT[19]) );
  AND U239 ( .A(A[18]), .B(B[0]), .Z(PRODUCT[18]) );
  AND U240 ( .A(A[17]), .B(B[0]), .Z(PRODUCT[17]) );
  AND U241 ( .A(A[16]), .B(B[0]), .Z(PRODUCT[16]) );
  AND U242 ( .A(A[15]), .B(B[0]), .Z(PRODUCT[15]) );
  AND U243 ( .A(A[14]), .B(B[0]), .Z(PRODUCT[14]) );
  AND U244 ( .A(A[13]), .B(B[0]), .Z(PRODUCT[13]) );
  AND U245 ( .A(A[12]), .B(B[0]), .Z(PRODUCT[12]) );
  AND U246 ( .A(A[11]), .B(B[0]), .Z(PRODUCT[11]) );
  AND U247 ( .A(A[10]), .B(B[0]), .Z(PRODUCT[10]) );
  AND U248 ( .A(B[0]), .B(A[9]), .Z(PRODUCT[9]) );
  AND U249 ( .A(A[8]), .B(B[0]), .Z(PRODUCT[8]) );
  AND U250 ( .A(A[7]), .B(B[0]), .Z(PRODUCT[7]) );
  AND U251 ( .A(A[6]), .B(B[0]), .Z(PRODUCT[6]) );
  AND U252 ( .A(A[5]), .B(B[0]), .Z(PRODUCT[5]) );
  AND U253 ( .A(A[4]), .B(B[0]), .Z(PRODUCT[4]) );
  AND U254 ( .A(A[3]), .B(B[0]), .Z(PRODUCT[3]) );
  AND U255 ( .A(A[2]), .B(B[0]), .Z(PRODUCT[2]) );
  AND U256 ( .A(A[1]), .B(B[0]), .Z(PRODUCT[1]) );
  AND U257 ( .A(A[0]), .B(B[0]), .Z(PRODUCT[0]) );
endmodule


module modmult_step_N256_3_DW01_cmp2_0 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [257:0] A;
  input [257:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;

  NAND U1 ( .A(n1), .B(n2), .Z(LT_LE) );
  NOR U2 ( .A(B[257]), .B(B[256]), .Z(n2) );
  AND U3 ( .A(n3), .B(n4), .Z(n1) );
  NAND U4 ( .A(n5), .B(n6), .Z(n4) );
  NANDN U5 ( .A(B[255]), .B(A[255]), .Z(n6) );
  NAND U6 ( .A(n7), .B(n8), .Z(n5) );
  NANDN U7 ( .A(A[254]), .B(B[254]), .Z(n8) );
  NAND U8 ( .A(n9), .B(n10), .Z(n7) );
  NANDN U9 ( .A(B[254]), .B(A[254]), .Z(n10) );
  AND U10 ( .A(n11), .B(n12), .Z(n9) );
  NAND U11 ( .A(n13), .B(n14), .Z(n12) );
  NANDN U12 ( .A(A[253]), .B(B[253]), .Z(n14) );
  AND U13 ( .A(n15), .B(n16), .Z(n13) );
  NANDN U14 ( .A(A[252]), .B(B[252]), .Z(n16) );
  NAND U15 ( .A(n17), .B(n18), .Z(n15) );
  NANDN U16 ( .A(B[252]), .B(A[252]), .Z(n18) );
  AND U17 ( .A(n19), .B(n20), .Z(n17) );
  NAND U18 ( .A(n21), .B(n22), .Z(n20) );
  NANDN U19 ( .A(A[251]), .B(B[251]), .Z(n22) );
  AND U20 ( .A(n23), .B(n24), .Z(n21) );
  NANDN U21 ( .A(A[250]), .B(B[250]), .Z(n24) );
  NAND U22 ( .A(n25), .B(n26), .Z(n23) );
  NANDN U23 ( .A(B[250]), .B(A[250]), .Z(n26) );
  AND U24 ( .A(n27), .B(n28), .Z(n25) );
  NAND U25 ( .A(n29), .B(n30), .Z(n28) );
  NANDN U26 ( .A(A[249]), .B(B[249]), .Z(n30) );
  AND U27 ( .A(n31), .B(n32), .Z(n29) );
  NANDN U28 ( .A(A[248]), .B(B[248]), .Z(n32) );
  NAND U29 ( .A(n33), .B(n34), .Z(n31) );
  NANDN U30 ( .A(B[248]), .B(A[248]), .Z(n34) );
  AND U31 ( .A(n35), .B(n36), .Z(n33) );
  NAND U32 ( .A(n37), .B(n38), .Z(n36) );
  NANDN U33 ( .A(A[247]), .B(B[247]), .Z(n38) );
  AND U34 ( .A(n39), .B(n40), .Z(n37) );
  NANDN U35 ( .A(A[246]), .B(B[246]), .Z(n40) );
  NAND U36 ( .A(n41), .B(n42), .Z(n39) );
  NANDN U37 ( .A(B[246]), .B(A[246]), .Z(n42) );
  AND U38 ( .A(n43), .B(n44), .Z(n41) );
  NAND U39 ( .A(n45), .B(n46), .Z(n44) );
  NANDN U40 ( .A(A[245]), .B(B[245]), .Z(n46) );
  AND U41 ( .A(n47), .B(n48), .Z(n45) );
  NANDN U42 ( .A(A[244]), .B(B[244]), .Z(n48) );
  NAND U43 ( .A(n49), .B(n50), .Z(n47) );
  NANDN U44 ( .A(B[244]), .B(A[244]), .Z(n50) );
  AND U45 ( .A(n51), .B(n52), .Z(n49) );
  NAND U46 ( .A(n53), .B(n54), .Z(n52) );
  NANDN U47 ( .A(A[243]), .B(B[243]), .Z(n54) );
  AND U48 ( .A(n55), .B(n56), .Z(n53) );
  NANDN U49 ( .A(A[242]), .B(B[242]), .Z(n56) );
  NAND U50 ( .A(n57), .B(n58), .Z(n55) );
  NANDN U51 ( .A(B[242]), .B(A[242]), .Z(n58) );
  AND U52 ( .A(n59), .B(n60), .Z(n57) );
  NAND U53 ( .A(n61), .B(n62), .Z(n60) );
  NANDN U54 ( .A(A[241]), .B(B[241]), .Z(n62) );
  AND U55 ( .A(n63), .B(n64), .Z(n61) );
  NANDN U56 ( .A(A[240]), .B(B[240]), .Z(n64) );
  NAND U57 ( .A(n65), .B(n66), .Z(n63) );
  NANDN U58 ( .A(B[240]), .B(A[240]), .Z(n66) );
  AND U59 ( .A(n67), .B(n68), .Z(n65) );
  NAND U60 ( .A(n69), .B(n70), .Z(n68) );
  NANDN U61 ( .A(A[239]), .B(B[239]), .Z(n70) );
  AND U62 ( .A(n71), .B(n72), .Z(n69) );
  NANDN U63 ( .A(A[238]), .B(B[238]), .Z(n72) );
  NAND U64 ( .A(n73), .B(n74), .Z(n71) );
  NANDN U65 ( .A(B[238]), .B(A[238]), .Z(n74) );
  AND U66 ( .A(n75), .B(n76), .Z(n73) );
  NAND U67 ( .A(n77), .B(n78), .Z(n76) );
  NANDN U68 ( .A(A[237]), .B(B[237]), .Z(n78) );
  AND U69 ( .A(n79), .B(n80), .Z(n77) );
  NANDN U70 ( .A(A[236]), .B(B[236]), .Z(n80) );
  NAND U71 ( .A(n81), .B(n82), .Z(n79) );
  NANDN U72 ( .A(B[236]), .B(A[236]), .Z(n82) );
  AND U73 ( .A(n83), .B(n84), .Z(n81) );
  NAND U74 ( .A(n85), .B(n86), .Z(n84) );
  NANDN U75 ( .A(A[235]), .B(B[235]), .Z(n86) );
  AND U76 ( .A(n87), .B(n88), .Z(n85) );
  NANDN U77 ( .A(A[234]), .B(B[234]), .Z(n88) );
  NAND U78 ( .A(n89), .B(n90), .Z(n87) );
  NANDN U79 ( .A(B[234]), .B(A[234]), .Z(n90) );
  AND U80 ( .A(n91), .B(n92), .Z(n89) );
  NAND U81 ( .A(n93), .B(n94), .Z(n92) );
  NANDN U82 ( .A(A[233]), .B(B[233]), .Z(n94) );
  AND U83 ( .A(n95), .B(n96), .Z(n93) );
  NANDN U84 ( .A(A[232]), .B(B[232]), .Z(n96) );
  NAND U85 ( .A(n97), .B(n98), .Z(n95) );
  NANDN U86 ( .A(B[232]), .B(A[232]), .Z(n98) );
  AND U87 ( .A(n99), .B(n100), .Z(n97) );
  NAND U88 ( .A(n101), .B(n102), .Z(n100) );
  NANDN U89 ( .A(A[231]), .B(B[231]), .Z(n102) );
  AND U90 ( .A(n103), .B(n104), .Z(n101) );
  NANDN U91 ( .A(A[230]), .B(B[230]), .Z(n104) );
  NAND U92 ( .A(n105), .B(n106), .Z(n103) );
  NANDN U93 ( .A(B[230]), .B(A[230]), .Z(n106) );
  AND U94 ( .A(n107), .B(n108), .Z(n105) );
  NAND U95 ( .A(n109), .B(n110), .Z(n108) );
  NANDN U96 ( .A(A[229]), .B(B[229]), .Z(n110) );
  AND U97 ( .A(n111), .B(n112), .Z(n109) );
  NANDN U98 ( .A(A[228]), .B(B[228]), .Z(n112) );
  NAND U99 ( .A(n113), .B(n114), .Z(n111) );
  NANDN U100 ( .A(B[228]), .B(A[228]), .Z(n114) );
  AND U101 ( .A(n115), .B(n116), .Z(n113) );
  NAND U102 ( .A(n117), .B(n118), .Z(n116) );
  NANDN U103 ( .A(A[227]), .B(B[227]), .Z(n118) );
  AND U104 ( .A(n119), .B(n120), .Z(n117) );
  NANDN U105 ( .A(A[226]), .B(B[226]), .Z(n120) );
  NAND U106 ( .A(n121), .B(n122), .Z(n119) );
  NANDN U107 ( .A(B[226]), .B(A[226]), .Z(n122) );
  AND U108 ( .A(n123), .B(n124), .Z(n121) );
  NAND U109 ( .A(n125), .B(n126), .Z(n124) );
  NANDN U110 ( .A(A[225]), .B(B[225]), .Z(n126) );
  AND U111 ( .A(n127), .B(n128), .Z(n125) );
  NANDN U112 ( .A(A[224]), .B(B[224]), .Z(n128) );
  NAND U113 ( .A(n129), .B(n130), .Z(n127) );
  NANDN U114 ( .A(B[224]), .B(A[224]), .Z(n130) );
  AND U115 ( .A(n131), .B(n132), .Z(n129) );
  NAND U116 ( .A(n133), .B(n134), .Z(n132) );
  NANDN U117 ( .A(A[223]), .B(B[223]), .Z(n134) );
  AND U118 ( .A(n135), .B(n136), .Z(n133) );
  NANDN U119 ( .A(A[222]), .B(B[222]), .Z(n136) );
  NAND U120 ( .A(n137), .B(n138), .Z(n135) );
  NANDN U121 ( .A(B[222]), .B(A[222]), .Z(n138) );
  AND U122 ( .A(n139), .B(n140), .Z(n137) );
  NAND U123 ( .A(n141), .B(n142), .Z(n140) );
  NANDN U124 ( .A(A[221]), .B(B[221]), .Z(n142) );
  AND U125 ( .A(n143), .B(n144), .Z(n141) );
  NANDN U126 ( .A(A[220]), .B(B[220]), .Z(n144) );
  NAND U127 ( .A(n145), .B(n146), .Z(n143) );
  NANDN U128 ( .A(B[220]), .B(A[220]), .Z(n146) );
  AND U129 ( .A(n147), .B(n148), .Z(n145) );
  NAND U130 ( .A(n149), .B(n150), .Z(n148) );
  NANDN U131 ( .A(A[219]), .B(B[219]), .Z(n150) );
  AND U132 ( .A(n151), .B(n152), .Z(n149) );
  NANDN U133 ( .A(A[218]), .B(B[218]), .Z(n152) );
  NAND U134 ( .A(n153), .B(n154), .Z(n151) );
  NANDN U135 ( .A(B[218]), .B(A[218]), .Z(n154) );
  AND U136 ( .A(n155), .B(n156), .Z(n153) );
  NAND U137 ( .A(n157), .B(n158), .Z(n156) );
  NANDN U138 ( .A(A[217]), .B(B[217]), .Z(n158) );
  AND U139 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U140 ( .A(A[216]), .B(B[216]), .Z(n160) );
  NAND U141 ( .A(n161), .B(n162), .Z(n159) );
  NANDN U142 ( .A(B[216]), .B(A[216]), .Z(n162) );
  AND U143 ( .A(n163), .B(n164), .Z(n161) );
  NAND U144 ( .A(n165), .B(n166), .Z(n164) );
  NANDN U145 ( .A(A[215]), .B(B[215]), .Z(n166) );
  AND U146 ( .A(n167), .B(n168), .Z(n165) );
  NANDN U147 ( .A(A[214]), .B(B[214]), .Z(n168) );
  NAND U148 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U149 ( .A(B[214]), .B(A[214]), .Z(n170) );
  AND U150 ( .A(n171), .B(n172), .Z(n169) );
  NAND U151 ( .A(n173), .B(n174), .Z(n172) );
  NANDN U152 ( .A(A[213]), .B(B[213]), .Z(n174) );
  AND U153 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U154 ( .A(A[212]), .B(B[212]), .Z(n176) );
  NAND U155 ( .A(n177), .B(n178), .Z(n175) );
  NANDN U156 ( .A(B[212]), .B(A[212]), .Z(n178) );
  AND U157 ( .A(n179), .B(n180), .Z(n177) );
  NAND U158 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U159 ( .A(A[211]), .B(B[211]), .Z(n182) );
  AND U160 ( .A(n183), .B(n184), .Z(n181) );
  NANDN U161 ( .A(A[210]), .B(B[210]), .Z(n184) );
  NAND U162 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U163 ( .A(B[210]), .B(A[210]), .Z(n186) );
  AND U164 ( .A(n187), .B(n188), .Z(n185) );
  NAND U165 ( .A(n189), .B(n190), .Z(n188) );
  NANDN U166 ( .A(A[209]), .B(B[209]), .Z(n190) );
  AND U167 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U168 ( .A(A[208]), .B(B[208]), .Z(n192) );
  NAND U169 ( .A(n193), .B(n194), .Z(n191) );
  NANDN U170 ( .A(B[208]), .B(A[208]), .Z(n194) );
  AND U171 ( .A(n195), .B(n196), .Z(n193) );
  NAND U172 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U173 ( .A(A[207]), .B(B[207]), .Z(n198) );
  AND U174 ( .A(n199), .B(n200), .Z(n197) );
  NANDN U175 ( .A(A[206]), .B(B[206]), .Z(n200) );
  NAND U176 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U177 ( .A(B[206]), .B(A[206]), .Z(n202) );
  AND U178 ( .A(n203), .B(n204), .Z(n201) );
  NAND U179 ( .A(n205), .B(n206), .Z(n204) );
  NANDN U180 ( .A(A[205]), .B(B[205]), .Z(n206) );
  AND U181 ( .A(n207), .B(n208), .Z(n205) );
  NANDN U182 ( .A(A[204]), .B(B[204]), .Z(n208) );
  NAND U183 ( .A(n209), .B(n210), .Z(n207) );
  NANDN U184 ( .A(B[204]), .B(A[204]), .Z(n210) );
  AND U185 ( .A(n211), .B(n212), .Z(n209) );
  NAND U186 ( .A(n213), .B(n214), .Z(n212) );
  NANDN U187 ( .A(A[203]), .B(B[203]), .Z(n214) );
  AND U188 ( .A(n215), .B(n216), .Z(n213) );
  NANDN U189 ( .A(A[202]), .B(B[202]), .Z(n216) );
  NAND U190 ( .A(n217), .B(n218), .Z(n215) );
  NANDN U191 ( .A(B[202]), .B(A[202]), .Z(n218) );
  AND U192 ( .A(n219), .B(n220), .Z(n217) );
  NAND U193 ( .A(n221), .B(n222), .Z(n220) );
  NANDN U194 ( .A(A[201]), .B(B[201]), .Z(n222) );
  AND U195 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U196 ( .A(A[200]), .B(B[200]), .Z(n224) );
  NAND U197 ( .A(n225), .B(n226), .Z(n223) );
  NANDN U198 ( .A(B[200]), .B(A[200]), .Z(n226) );
  AND U199 ( .A(n227), .B(n228), .Z(n225) );
  NAND U200 ( .A(n229), .B(n230), .Z(n228) );
  NANDN U201 ( .A(A[199]), .B(B[199]), .Z(n230) );
  AND U202 ( .A(n231), .B(n232), .Z(n229) );
  NANDN U203 ( .A(A[198]), .B(B[198]), .Z(n232) );
  NAND U204 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U205 ( .A(B[198]), .B(A[198]), .Z(n234) );
  AND U206 ( .A(n235), .B(n236), .Z(n233) );
  NAND U207 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U208 ( .A(A[197]), .B(B[197]), .Z(n238) );
  AND U209 ( .A(n239), .B(n240), .Z(n237) );
  NANDN U210 ( .A(A[196]), .B(B[196]), .Z(n240) );
  NAND U211 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U212 ( .A(B[196]), .B(A[196]), .Z(n242) );
  AND U213 ( .A(n243), .B(n244), .Z(n241) );
  NAND U214 ( .A(n245), .B(n246), .Z(n244) );
  NANDN U215 ( .A(A[195]), .B(B[195]), .Z(n246) );
  AND U216 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U217 ( .A(A[194]), .B(B[194]), .Z(n248) );
  NAND U218 ( .A(n249), .B(n250), .Z(n247) );
  NANDN U219 ( .A(B[194]), .B(A[194]), .Z(n250) );
  AND U220 ( .A(n251), .B(n252), .Z(n249) );
  NAND U221 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U222 ( .A(A[193]), .B(B[193]), .Z(n254) );
  AND U223 ( .A(n255), .B(n256), .Z(n253) );
  NANDN U224 ( .A(A[192]), .B(B[192]), .Z(n256) );
  NAND U225 ( .A(n257), .B(n258), .Z(n255) );
  NANDN U226 ( .A(B[192]), .B(A[192]), .Z(n258) );
  AND U227 ( .A(n259), .B(n260), .Z(n257) );
  NAND U228 ( .A(n261), .B(n262), .Z(n260) );
  NANDN U229 ( .A(A[191]), .B(B[191]), .Z(n262) );
  AND U230 ( .A(n263), .B(n264), .Z(n261) );
  NANDN U231 ( .A(A[190]), .B(B[190]), .Z(n264) );
  NAND U232 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U233 ( .A(B[190]), .B(A[190]), .Z(n266) );
  AND U234 ( .A(n267), .B(n268), .Z(n265) );
  NAND U235 ( .A(n269), .B(n270), .Z(n268) );
  NANDN U236 ( .A(A[189]), .B(B[189]), .Z(n270) );
  AND U237 ( .A(n271), .B(n272), .Z(n269) );
  NANDN U238 ( .A(A[188]), .B(B[188]), .Z(n272) );
  NAND U239 ( .A(n273), .B(n274), .Z(n271) );
  NANDN U240 ( .A(B[188]), .B(A[188]), .Z(n274) );
  AND U241 ( .A(n275), .B(n276), .Z(n273) );
  NAND U242 ( .A(n277), .B(n278), .Z(n276) );
  NANDN U243 ( .A(A[187]), .B(B[187]), .Z(n278) );
  AND U244 ( .A(n279), .B(n280), .Z(n277) );
  NANDN U245 ( .A(A[186]), .B(B[186]), .Z(n280) );
  NAND U246 ( .A(n281), .B(n282), .Z(n279) );
  NANDN U247 ( .A(B[186]), .B(A[186]), .Z(n282) );
  AND U248 ( .A(n283), .B(n284), .Z(n281) );
  NAND U249 ( .A(n285), .B(n286), .Z(n284) );
  NANDN U250 ( .A(A[185]), .B(B[185]), .Z(n286) );
  AND U251 ( .A(n287), .B(n288), .Z(n285) );
  NANDN U252 ( .A(A[184]), .B(B[184]), .Z(n288) );
  NAND U253 ( .A(n289), .B(n290), .Z(n287) );
  NANDN U254 ( .A(B[184]), .B(A[184]), .Z(n290) );
  AND U255 ( .A(n291), .B(n292), .Z(n289) );
  NAND U256 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U257 ( .A(A[183]), .B(B[183]), .Z(n294) );
  AND U258 ( .A(n295), .B(n296), .Z(n293) );
  NANDN U259 ( .A(A[182]), .B(B[182]), .Z(n296) );
  NAND U260 ( .A(n297), .B(n298), .Z(n295) );
  NANDN U261 ( .A(B[182]), .B(A[182]), .Z(n298) );
  AND U262 ( .A(n299), .B(n300), .Z(n297) );
  NAND U263 ( .A(n301), .B(n302), .Z(n300) );
  NANDN U264 ( .A(A[181]), .B(B[181]), .Z(n302) );
  AND U265 ( .A(n303), .B(n304), .Z(n301) );
  NANDN U266 ( .A(A[180]), .B(B[180]), .Z(n304) );
  NAND U267 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U268 ( .A(B[180]), .B(A[180]), .Z(n306) );
  AND U269 ( .A(n307), .B(n308), .Z(n305) );
  NAND U270 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U271 ( .A(A[179]), .B(B[179]), .Z(n310) );
  AND U272 ( .A(n311), .B(n312), .Z(n309) );
  NANDN U273 ( .A(A[178]), .B(B[178]), .Z(n312) );
  NAND U274 ( .A(n313), .B(n314), .Z(n311) );
  NANDN U275 ( .A(B[178]), .B(A[178]), .Z(n314) );
  AND U276 ( .A(n315), .B(n316), .Z(n313) );
  NAND U277 ( .A(n317), .B(n318), .Z(n316) );
  NANDN U278 ( .A(A[177]), .B(B[177]), .Z(n318) );
  AND U279 ( .A(n319), .B(n320), .Z(n317) );
  NANDN U280 ( .A(A[176]), .B(B[176]), .Z(n320) );
  NAND U281 ( .A(n321), .B(n322), .Z(n319) );
  NANDN U282 ( .A(B[176]), .B(A[176]), .Z(n322) );
  AND U283 ( .A(n323), .B(n324), .Z(n321) );
  NAND U284 ( .A(n325), .B(n326), .Z(n324) );
  NANDN U285 ( .A(A[175]), .B(B[175]), .Z(n326) );
  AND U286 ( .A(n327), .B(n328), .Z(n325) );
  NANDN U287 ( .A(A[174]), .B(B[174]), .Z(n328) );
  NAND U288 ( .A(n329), .B(n330), .Z(n327) );
  NANDN U289 ( .A(B[174]), .B(A[174]), .Z(n330) );
  AND U290 ( .A(n331), .B(n332), .Z(n329) );
  NAND U291 ( .A(n333), .B(n334), .Z(n332) );
  NANDN U292 ( .A(A[173]), .B(B[173]), .Z(n334) );
  AND U293 ( .A(n335), .B(n336), .Z(n333) );
  NANDN U294 ( .A(A[172]), .B(B[172]), .Z(n336) );
  NAND U295 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U296 ( .A(B[172]), .B(A[172]), .Z(n338) );
  AND U297 ( .A(n339), .B(n340), .Z(n337) );
  NAND U298 ( .A(n341), .B(n342), .Z(n340) );
  NANDN U299 ( .A(A[171]), .B(B[171]), .Z(n342) );
  AND U300 ( .A(n343), .B(n344), .Z(n341) );
  NANDN U301 ( .A(A[170]), .B(B[170]), .Z(n344) );
  NAND U302 ( .A(n345), .B(n346), .Z(n343) );
  NANDN U303 ( .A(B[170]), .B(A[170]), .Z(n346) );
  AND U304 ( .A(n347), .B(n348), .Z(n345) );
  NAND U305 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U306 ( .A(A[169]), .B(B[169]), .Z(n350) );
  AND U307 ( .A(n351), .B(n352), .Z(n349) );
  NANDN U308 ( .A(A[168]), .B(B[168]), .Z(n352) );
  NAND U309 ( .A(n353), .B(n354), .Z(n351) );
  NANDN U310 ( .A(B[168]), .B(A[168]), .Z(n354) );
  AND U311 ( .A(n355), .B(n356), .Z(n353) );
  NAND U312 ( .A(n357), .B(n358), .Z(n356) );
  NANDN U313 ( .A(A[167]), .B(B[167]), .Z(n358) );
  AND U314 ( .A(n359), .B(n360), .Z(n357) );
  NANDN U315 ( .A(A[166]), .B(B[166]), .Z(n360) );
  NAND U316 ( .A(n361), .B(n362), .Z(n359) );
  NANDN U317 ( .A(B[166]), .B(A[166]), .Z(n362) );
  AND U318 ( .A(n363), .B(n364), .Z(n361) );
  NAND U319 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U320 ( .A(A[165]), .B(B[165]), .Z(n366) );
  AND U321 ( .A(n367), .B(n368), .Z(n365) );
  NANDN U322 ( .A(A[164]), .B(B[164]), .Z(n368) );
  NAND U323 ( .A(n369), .B(n370), .Z(n367) );
  NANDN U324 ( .A(B[164]), .B(A[164]), .Z(n370) );
  AND U325 ( .A(n371), .B(n372), .Z(n369) );
  NAND U326 ( .A(n373), .B(n374), .Z(n372) );
  NANDN U327 ( .A(A[163]), .B(B[163]), .Z(n374) );
  AND U328 ( .A(n375), .B(n376), .Z(n373) );
  NANDN U329 ( .A(A[162]), .B(B[162]), .Z(n376) );
  NAND U330 ( .A(n377), .B(n378), .Z(n375) );
  NANDN U331 ( .A(B[162]), .B(A[162]), .Z(n378) );
  AND U332 ( .A(n379), .B(n380), .Z(n377) );
  NAND U333 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U334 ( .A(A[161]), .B(B[161]), .Z(n382) );
  AND U335 ( .A(n383), .B(n384), .Z(n381) );
  NANDN U336 ( .A(A[160]), .B(B[160]), .Z(n384) );
  NAND U337 ( .A(n385), .B(n386), .Z(n383) );
  NANDN U338 ( .A(B[160]), .B(A[160]), .Z(n386) );
  AND U339 ( .A(n387), .B(n388), .Z(n385) );
  NAND U340 ( .A(n389), .B(n390), .Z(n388) );
  NANDN U341 ( .A(A[159]), .B(B[159]), .Z(n390) );
  AND U342 ( .A(n391), .B(n392), .Z(n389) );
  NANDN U343 ( .A(A[158]), .B(B[158]), .Z(n392) );
  NAND U344 ( .A(n393), .B(n394), .Z(n391) );
  NANDN U345 ( .A(B[158]), .B(A[158]), .Z(n394) );
  AND U346 ( .A(n395), .B(n396), .Z(n393) );
  NAND U347 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U348 ( .A(A[157]), .B(B[157]), .Z(n398) );
  AND U349 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U350 ( .A(A[156]), .B(B[156]), .Z(n400) );
  NAND U351 ( .A(n401), .B(n402), .Z(n399) );
  NANDN U352 ( .A(B[156]), .B(A[156]), .Z(n402) );
  AND U353 ( .A(n403), .B(n404), .Z(n401) );
  NAND U354 ( .A(n405), .B(n406), .Z(n404) );
  NANDN U355 ( .A(A[155]), .B(B[155]), .Z(n406) );
  AND U356 ( .A(n407), .B(n408), .Z(n405) );
  NANDN U357 ( .A(A[154]), .B(B[154]), .Z(n408) );
  NAND U358 ( .A(n409), .B(n410), .Z(n407) );
  NANDN U359 ( .A(B[154]), .B(A[154]), .Z(n410) );
  AND U360 ( .A(n411), .B(n412), .Z(n409) );
  NAND U361 ( .A(n413), .B(n414), .Z(n412) );
  NANDN U362 ( .A(A[153]), .B(B[153]), .Z(n414) );
  AND U363 ( .A(n415), .B(n416), .Z(n413) );
  NANDN U364 ( .A(A[152]), .B(B[152]), .Z(n416) );
  NAND U365 ( .A(n417), .B(n418), .Z(n415) );
  NANDN U366 ( .A(B[152]), .B(A[152]), .Z(n418) );
  AND U367 ( .A(n419), .B(n420), .Z(n417) );
  NAND U368 ( .A(n421), .B(n422), .Z(n420) );
  NANDN U369 ( .A(A[151]), .B(B[151]), .Z(n422) );
  AND U370 ( .A(n423), .B(n424), .Z(n421) );
  NANDN U371 ( .A(A[150]), .B(B[150]), .Z(n424) );
  NAND U372 ( .A(n425), .B(n426), .Z(n423) );
  NANDN U373 ( .A(B[150]), .B(A[150]), .Z(n426) );
  AND U374 ( .A(n427), .B(n428), .Z(n425) );
  NAND U375 ( .A(n429), .B(n430), .Z(n428) );
  NANDN U376 ( .A(A[149]), .B(B[149]), .Z(n430) );
  AND U377 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U378 ( .A(A[148]), .B(B[148]), .Z(n432) );
  NAND U379 ( .A(n433), .B(n434), .Z(n431) );
  NANDN U380 ( .A(B[148]), .B(A[148]), .Z(n434) );
  AND U381 ( .A(n435), .B(n436), .Z(n433) );
  NAND U382 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U383 ( .A(A[147]), .B(B[147]), .Z(n438) );
  AND U384 ( .A(n439), .B(n440), .Z(n437) );
  NANDN U385 ( .A(A[146]), .B(B[146]), .Z(n440) );
  NAND U386 ( .A(n441), .B(n442), .Z(n439) );
  NANDN U387 ( .A(B[146]), .B(A[146]), .Z(n442) );
  AND U388 ( .A(n443), .B(n444), .Z(n441) );
  NAND U389 ( .A(n445), .B(n446), .Z(n444) );
  NANDN U390 ( .A(A[145]), .B(B[145]), .Z(n446) );
  AND U391 ( .A(n447), .B(n448), .Z(n445) );
  NANDN U392 ( .A(A[144]), .B(B[144]), .Z(n448) );
  NAND U393 ( .A(n449), .B(n450), .Z(n447) );
  NANDN U394 ( .A(B[144]), .B(A[144]), .Z(n450) );
  AND U395 ( .A(n451), .B(n452), .Z(n449) );
  NAND U396 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U397 ( .A(A[143]), .B(B[143]), .Z(n454) );
  AND U398 ( .A(n455), .B(n456), .Z(n453) );
  NANDN U399 ( .A(A[142]), .B(B[142]), .Z(n456) );
  NAND U400 ( .A(n457), .B(n458), .Z(n455) );
  NANDN U401 ( .A(B[142]), .B(A[142]), .Z(n458) );
  AND U402 ( .A(n459), .B(n460), .Z(n457) );
  NAND U403 ( .A(n461), .B(n462), .Z(n460) );
  NANDN U404 ( .A(A[141]), .B(B[141]), .Z(n462) );
  AND U405 ( .A(n463), .B(n464), .Z(n461) );
  NANDN U406 ( .A(A[140]), .B(B[140]), .Z(n464) );
  NAND U407 ( .A(n465), .B(n466), .Z(n463) );
  NANDN U408 ( .A(B[140]), .B(A[140]), .Z(n466) );
  AND U409 ( .A(n467), .B(n468), .Z(n465) );
  NAND U410 ( .A(n469), .B(n470), .Z(n468) );
  NANDN U411 ( .A(A[139]), .B(B[139]), .Z(n470) );
  AND U412 ( .A(n471), .B(n472), .Z(n469) );
  NANDN U413 ( .A(A[138]), .B(B[138]), .Z(n472) );
  NAND U414 ( .A(n473), .B(n474), .Z(n471) );
  NANDN U415 ( .A(B[138]), .B(A[138]), .Z(n474) );
  AND U416 ( .A(n475), .B(n476), .Z(n473) );
  NAND U417 ( .A(n477), .B(n478), .Z(n476) );
  NANDN U418 ( .A(A[137]), .B(B[137]), .Z(n478) );
  AND U419 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U420 ( .A(A[136]), .B(B[136]), .Z(n480) );
  NAND U421 ( .A(n481), .B(n482), .Z(n479) );
  NANDN U422 ( .A(B[136]), .B(A[136]), .Z(n482) );
  AND U423 ( .A(n483), .B(n484), .Z(n481) );
  NAND U424 ( .A(n485), .B(n486), .Z(n484) );
  NANDN U425 ( .A(A[135]), .B(B[135]), .Z(n486) );
  AND U426 ( .A(n487), .B(n488), .Z(n485) );
  NANDN U427 ( .A(A[134]), .B(B[134]), .Z(n488) );
  NAND U428 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U429 ( .A(B[134]), .B(A[134]), .Z(n490) );
  AND U430 ( .A(n491), .B(n492), .Z(n489) );
  NAND U431 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U432 ( .A(A[133]), .B(B[133]), .Z(n494) );
  AND U433 ( .A(n495), .B(n496), .Z(n493) );
  NANDN U434 ( .A(A[132]), .B(B[132]), .Z(n496) );
  NAND U435 ( .A(n497), .B(n498), .Z(n495) );
  NANDN U436 ( .A(B[132]), .B(A[132]), .Z(n498) );
  AND U437 ( .A(n499), .B(n500), .Z(n497) );
  NAND U438 ( .A(n501), .B(n502), .Z(n500) );
  NANDN U439 ( .A(A[131]), .B(B[131]), .Z(n502) );
  AND U440 ( .A(n503), .B(n504), .Z(n501) );
  NANDN U441 ( .A(A[130]), .B(B[130]), .Z(n504) );
  NAND U442 ( .A(n505), .B(n506), .Z(n503) );
  NANDN U443 ( .A(B[130]), .B(A[130]), .Z(n506) );
  AND U444 ( .A(n507), .B(n508), .Z(n505) );
  NAND U445 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U446 ( .A(A[129]), .B(B[129]), .Z(n510) );
  AND U447 ( .A(n511), .B(n512), .Z(n509) );
  NANDN U448 ( .A(A[128]), .B(B[128]), .Z(n512) );
  NAND U449 ( .A(n513), .B(n514), .Z(n511) );
  NANDN U450 ( .A(B[128]), .B(A[128]), .Z(n514) );
  AND U451 ( .A(n515), .B(n516), .Z(n513) );
  NAND U452 ( .A(n517), .B(n518), .Z(n516) );
  NANDN U453 ( .A(A[127]), .B(B[127]), .Z(n518) );
  AND U454 ( .A(n519), .B(n520), .Z(n517) );
  NANDN U455 ( .A(A[126]), .B(B[126]), .Z(n520) );
  NAND U456 ( .A(n521), .B(n522), .Z(n519) );
  NANDN U457 ( .A(B[126]), .B(A[126]), .Z(n522) );
  AND U458 ( .A(n523), .B(n524), .Z(n521) );
  NAND U459 ( .A(n525), .B(n526), .Z(n524) );
  NANDN U460 ( .A(A[125]), .B(B[125]), .Z(n526) );
  AND U461 ( .A(n527), .B(n528), .Z(n525) );
  NANDN U462 ( .A(A[124]), .B(B[124]), .Z(n528) );
  NAND U463 ( .A(n529), .B(n530), .Z(n527) );
  NANDN U464 ( .A(B[124]), .B(A[124]), .Z(n530) );
  AND U465 ( .A(n531), .B(n532), .Z(n529) );
  NAND U466 ( .A(n533), .B(n534), .Z(n532) );
  NANDN U467 ( .A(A[123]), .B(B[123]), .Z(n534) );
  AND U468 ( .A(n535), .B(n536), .Z(n533) );
  NANDN U469 ( .A(A[122]), .B(B[122]), .Z(n536) );
  NAND U470 ( .A(n537), .B(n538), .Z(n535) );
  NANDN U471 ( .A(B[122]), .B(A[122]), .Z(n538) );
  AND U472 ( .A(n539), .B(n540), .Z(n537) );
  NAND U473 ( .A(n541), .B(n542), .Z(n540) );
  NANDN U474 ( .A(A[121]), .B(B[121]), .Z(n542) );
  AND U475 ( .A(n543), .B(n544), .Z(n541) );
  NANDN U476 ( .A(A[120]), .B(B[120]), .Z(n544) );
  NAND U477 ( .A(n545), .B(n546), .Z(n543) );
  NANDN U478 ( .A(B[120]), .B(A[120]), .Z(n546) );
  AND U479 ( .A(n547), .B(n548), .Z(n545) );
  NAND U480 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U481 ( .A(A[119]), .B(B[119]), .Z(n550) );
  AND U482 ( .A(n551), .B(n552), .Z(n549) );
  NANDN U483 ( .A(A[118]), .B(B[118]), .Z(n552) );
  NAND U484 ( .A(n553), .B(n554), .Z(n551) );
  NANDN U485 ( .A(B[118]), .B(A[118]), .Z(n554) );
  AND U486 ( .A(n555), .B(n556), .Z(n553) );
  NAND U487 ( .A(n557), .B(n558), .Z(n556) );
  NANDN U488 ( .A(A[117]), .B(B[117]), .Z(n558) );
  AND U489 ( .A(n559), .B(n560), .Z(n557) );
  NANDN U490 ( .A(A[116]), .B(B[116]), .Z(n560) );
  NAND U491 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U492 ( .A(B[116]), .B(A[116]), .Z(n562) );
  AND U493 ( .A(n563), .B(n564), .Z(n561) );
  NAND U494 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U495 ( .A(A[115]), .B(B[115]), .Z(n566) );
  AND U496 ( .A(n567), .B(n568), .Z(n565) );
  NANDN U497 ( .A(A[114]), .B(B[114]), .Z(n568) );
  NAND U498 ( .A(n569), .B(n570), .Z(n567) );
  NANDN U499 ( .A(B[114]), .B(A[114]), .Z(n570) );
  AND U500 ( .A(n571), .B(n572), .Z(n569) );
  NAND U501 ( .A(n573), .B(n574), .Z(n572) );
  NANDN U502 ( .A(A[113]), .B(B[113]), .Z(n574) );
  AND U503 ( .A(n575), .B(n576), .Z(n573) );
  NANDN U504 ( .A(A[112]), .B(B[112]), .Z(n576) );
  NAND U505 ( .A(n577), .B(n578), .Z(n575) );
  NANDN U506 ( .A(B[112]), .B(A[112]), .Z(n578) );
  AND U507 ( .A(n579), .B(n580), .Z(n577) );
  NAND U508 ( .A(n581), .B(n582), .Z(n580) );
  NANDN U509 ( .A(A[111]), .B(B[111]), .Z(n582) );
  AND U510 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U511 ( .A(A[110]), .B(B[110]), .Z(n584) );
  NAND U512 ( .A(n585), .B(n586), .Z(n583) );
  NANDN U513 ( .A(B[110]), .B(A[110]), .Z(n586) );
  AND U514 ( .A(n587), .B(n588), .Z(n585) );
  NAND U515 ( .A(n589), .B(n590), .Z(n588) );
  NANDN U516 ( .A(A[109]), .B(B[109]), .Z(n590) );
  AND U517 ( .A(n591), .B(n592), .Z(n589) );
  NANDN U518 ( .A(A[108]), .B(B[108]), .Z(n592) );
  NAND U519 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U520 ( .A(B[108]), .B(A[108]), .Z(n594) );
  AND U521 ( .A(n595), .B(n596), .Z(n593) );
  NAND U522 ( .A(n597), .B(n598), .Z(n596) );
  NANDN U523 ( .A(A[107]), .B(B[107]), .Z(n598) );
  AND U524 ( .A(n599), .B(n600), .Z(n597) );
  NANDN U525 ( .A(A[106]), .B(B[106]), .Z(n600) );
  NAND U526 ( .A(n601), .B(n602), .Z(n599) );
  NANDN U527 ( .A(B[106]), .B(A[106]), .Z(n602) );
  AND U528 ( .A(n603), .B(n604), .Z(n601) );
  NAND U529 ( .A(n605), .B(n606), .Z(n604) );
  NANDN U530 ( .A(A[105]), .B(B[105]), .Z(n606) );
  AND U531 ( .A(n607), .B(n608), .Z(n605) );
  NANDN U532 ( .A(A[104]), .B(B[104]), .Z(n608) );
  NAND U533 ( .A(n609), .B(n610), .Z(n607) );
  NANDN U534 ( .A(B[104]), .B(A[104]), .Z(n610) );
  AND U535 ( .A(n611), .B(n612), .Z(n609) );
  NAND U536 ( .A(n613), .B(n614), .Z(n612) );
  NANDN U537 ( .A(A[103]), .B(B[103]), .Z(n614) );
  AND U538 ( .A(n615), .B(n616), .Z(n613) );
  NANDN U539 ( .A(A[102]), .B(B[102]), .Z(n616) );
  NAND U540 ( .A(n617), .B(n618), .Z(n615) );
  NANDN U541 ( .A(B[102]), .B(A[102]), .Z(n618) );
  AND U542 ( .A(n619), .B(n620), .Z(n617) );
  NAND U543 ( .A(n621), .B(n622), .Z(n620) );
  NANDN U544 ( .A(A[101]), .B(B[101]), .Z(n622) );
  AND U545 ( .A(n623), .B(n624), .Z(n621) );
  NANDN U546 ( .A(A[100]), .B(B[100]), .Z(n624) );
  NAND U547 ( .A(n625), .B(n626), .Z(n623) );
  NANDN U548 ( .A(B[99]), .B(A[99]), .Z(n626) );
  AND U549 ( .A(n627), .B(n628), .Z(n625) );
  NAND U550 ( .A(n629), .B(n630), .Z(n628) );
  NANDN U551 ( .A(A[99]), .B(B[99]), .Z(n630) );
  AND U552 ( .A(n631), .B(n632), .Z(n629) );
  NANDN U553 ( .A(A[98]), .B(B[98]), .Z(n632) );
  NAND U554 ( .A(n633), .B(n634), .Z(n631) );
  NANDN U555 ( .A(B[98]), .B(A[98]), .Z(n634) );
  AND U556 ( .A(n635), .B(n636), .Z(n633) );
  NAND U557 ( .A(n637), .B(n638), .Z(n636) );
  NANDN U558 ( .A(A[97]), .B(B[97]), .Z(n638) );
  AND U559 ( .A(n639), .B(n640), .Z(n637) );
  NANDN U560 ( .A(A[96]), .B(B[96]), .Z(n640) );
  NAND U561 ( .A(n641), .B(n642), .Z(n639) );
  NANDN U562 ( .A(B[96]), .B(A[96]), .Z(n642) );
  AND U563 ( .A(n643), .B(n644), .Z(n641) );
  NAND U564 ( .A(n645), .B(n646), .Z(n644) );
  NANDN U565 ( .A(A[95]), .B(B[95]), .Z(n646) );
  AND U566 ( .A(n647), .B(n648), .Z(n645) );
  NANDN U567 ( .A(A[94]), .B(B[94]), .Z(n648) );
  NAND U568 ( .A(n649), .B(n650), .Z(n647) );
  NANDN U569 ( .A(B[94]), .B(A[94]), .Z(n650) );
  AND U570 ( .A(n651), .B(n652), .Z(n649) );
  NAND U571 ( .A(n653), .B(n654), .Z(n652) );
  NANDN U572 ( .A(A[93]), .B(B[93]), .Z(n654) );
  AND U573 ( .A(n655), .B(n656), .Z(n653) );
  NANDN U574 ( .A(A[92]), .B(B[92]), .Z(n656) );
  NAND U575 ( .A(n657), .B(n658), .Z(n655) );
  NANDN U576 ( .A(B[92]), .B(A[92]), .Z(n658) );
  AND U577 ( .A(n659), .B(n660), .Z(n657) );
  NAND U578 ( .A(n661), .B(n662), .Z(n660) );
  NANDN U579 ( .A(A[91]), .B(B[91]), .Z(n662) );
  AND U580 ( .A(n663), .B(n664), .Z(n661) );
  NANDN U581 ( .A(A[90]), .B(B[90]), .Z(n664) );
  NAND U582 ( .A(n665), .B(n666), .Z(n663) );
  NANDN U583 ( .A(B[90]), .B(A[90]), .Z(n666) );
  AND U584 ( .A(n667), .B(n668), .Z(n665) );
  NAND U585 ( .A(n669), .B(n670), .Z(n668) );
  NANDN U586 ( .A(A[89]), .B(B[89]), .Z(n670) );
  AND U587 ( .A(n671), .B(n672), .Z(n669) );
  NANDN U588 ( .A(A[88]), .B(B[88]), .Z(n672) );
  NAND U589 ( .A(n673), .B(n674), .Z(n671) );
  NANDN U590 ( .A(B[88]), .B(A[88]), .Z(n674) );
  AND U591 ( .A(n675), .B(n676), .Z(n673) );
  NAND U592 ( .A(n677), .B(n678), .Z(n676) );
  NANDN U593 ( .A(A[87]), .B(B[87]), .Z(n678) );
  AND U594 ( .A(n679), .B(n680), .Z(n677) );
  NANDN U595 ( .A(A[86]), .B(B[86]), .Z(n680) );
  NAND U596 ( .A(n681), .B(n682), .Z(n679) );
  NANDN U597 ( .A(B[86]), .B(A[86]), .Z(n682) );
  AND U598 ( .A(n683), .B(n684), .Z(n681) );
  NAND U599 ( .A(n685), .B(n686), .Z(n684) );
  NANDN U600 ( .A(A[85]), .B(B[85]), .Z(n686) );
  AND U601 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U602 ( .A(A[84]), .B(B[84]), .Z(n688) );
  NAND U603 ( .A(n689), .B(n690), .Z(n687) );
  NANDN U604 ( .A(B[84]), .B(A[84]), .Z(n690) );
  AND U605 ( .A(n691), .B(n692), .Z(n689) );
  NAND U606 ( .A(n693), .B(n694), .Z(n692) );
  NANDN U607 ( .A(A[83]), .B(B[83]), .Z(n694) );
  AND U608 ( .A(n695), .B(n696), .Z(n693) );
  NANDN U609 ( .A(A[82]), .B(B[82]), .Z(n696) );
  NAND U610 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U611 ( .A(B[82]), .B(A[82]), .Z(n698) );
  AND U612 ( .A(n699), .B(n700), .Z(n697) );
  NAND U613 ( .A(n701), .B(n702), .Z(n700) );
  NANDN U614 ( .A(A[81]), .B(B[81]), .Z(n702) );
  AND U615 ( .A(n703), .B(n704), .Z(n701) );
  NANDN U616 ( .A(A[80]), .B(B[80]), .Z(n704) );
  NAND U617 ( .A(n705), .B(n706), .Z(n703) );
  NANDN U618 ( .A(B[80]), .B(A[80]), .Z(n706) );
  AND U619 ( .A(n707), .B(n708), .Z(n705) );
  NAND U620 ( .A(n709), .B(n710), .Z(n708) );
  NANDN U621 ( .A(A[79]), .B(B[79]), .Z(n710) );
  AND U622 ( .A(n711), .B(n712), .Z(n709) );
  NANDN U623 ( .A(A[78]), .B(B[78]), .Z(n712) );
  NAND U624 ( .A(n713), .B(n714), .Z(n711) );
  NANDN U625 ( .A(B[78]), .B(A[78]), .Z(n714) );
  AND U626 ( .A(n715), .B(n716), .Z(n713) );
  NAND U627 ( .A(n717), .B(n718), .Z(n716) );
  NANDN U628 ( .A(A[77]), .B(B[77]), .Z(n718) );
  AND U629 ( .A(n719), .B(n720), .Z(n717) );
  NANDN U630 ( .A(A[76]), .B(B[76]), .Z(n720) );
  NAND U631 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U632 ( .A(B[76]), .B(A[76]), .Z(n722) );
  AND U633 ( .A(n723), .B(n724), .Z(n721) );
  NAND U634 ( .A(n725), .B(n726), .Z(n724) );
  NANDN U635 ( .A(A[75]), .B(B[75]), .Z(n726) );
  AND U636 ( .A(n727), .B(n728), .Z(n725) );
  NANDN U637 ( .A(A[74]), .B(B[74]), .Z(n728) );
  NAND U638 ( .A(n729), .B(n730), .Z(n727) );
  NANDN U639 ( .A(B[74]), .B(A[74]), .Z(n730) );
  AND U640 ( .A(n731), .B(n732), .Z(n729) );
  NAND U641 ( .A(n733), .B(n734), .Z(n732) );
  NANDN U642 ( .A(A[73]), .B(B[73]), .Z(n734) );
  AND U643 ( .A(n735), .B(n736), .Z(n733) );
  NANDN U644 ( .A(A[72]), .B(B[72]), .Z(n736) );
  NAND U645 ( .A(n737), .B(n738), .Z(n735) );
  NANDN U646 ( .A(B[72]), .B(A[72]), .Z(n738) );
  AND U647 ( .A(n739), .B(n740), .Z(n737) );
  NAND U648 ( .A(n741), .B(n742), .Z(n740) );
  NANDN U649 ( .A(A[71]), .B(B[71]), .Z(n742) );
  AND U650 ( .A(n743), .B(n744), .Z(n741) );
  NANDN U651 ( .A(A[70]), .B(B[70]), .Z(n744) );
  NAND U652 ( .A(n745), .B(n746), .Z(n743) );
  NANDN U653 ( .A(B[70]), .B(A[70]), .Z(n746) );
  AND U654 ( .A(n747), .B(n748), .Z(n745) );
  NAND U655 ( .A(n749), .B(n750), .Z(n748) );
  NANDN U656 ( .A(A[69]), .B(B[69]), .Z(n750) );
  AND U657 ( .A(n751), .B(n752), .Z(n749) );
  NANDN U658 ( .A(A[68]), .B(B[68]), .Z(n752) );
  NAND U659 ( .A(n753), .B(n754), .Z(n751) );
  NANDN U660 ( .A(B[68]), .B(A[68]), .Z(n754) );
  AND U661 ( .A(n755), .B(n756), .Z(n753) );
  NAND U662 ( .A(n757), .B(n758), .Z(n756) );
  NANDN U663 ( .A(A[67]), .B(B[67]), .Z(n758) );
  AND U664 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U665 ( .A(A[66]), .B(B[66]), .Z(n760) );
  NAND U666 ( .A(n761), .B(n762), .Z(n759) );
  NANDN U667 ( .A(B[66]), .B(A[66]), .Z(n762) );
  AND U668 ( .A(n763), .B(n764), .Z(n761) );
  NAND U669 ( .A(n765), .B(n766), .Z(n764) );
  NANDN U670 ( .A(A[65]), .B(B[65]), .Z(n766) );
  AND U671 ( .A(n767), .B(n768), .Z(n765) );
  NANDN U672 ( .A(A[64]), .B(B[64]), .Z(n768) );
  NAND U673 ( .A(n769), .B(n770), .Z(n767) );
  NANDN U674 ( .A(B[64]), .B(A[64]), .Z(n770) );
  AND U675 ( .A(n771), .B(n772), .Z(n769) );
  NAND U676 ( .A(n773), .B(n774), .Z(n772) );
  NANDN U677 ( .A(A[63]), .B(B[63]), .Z(n774) );
  AND U678 ( .A(n775), .B(n776), .Z(n773) );
  NANDN U679 ( .A(A[62]), .B(B[62]), .Z(n776) );
  NAND U680 ( .A(n777), .B(n778), .Z(n775) );
  NANDN U681 ( .A(B[62]), .B(A[62]), .Z(n778) );
  AND U682 ( .A(n779), .B(n780), .Z(n777) );
  NAND U683 ( .A(n781), .B(n782), .Z(n780) );
  NANDN U684 ( .A(A[61]), .B(B[61]), .Z(n782) );
  AND U685 ( .A(n783), .B(n784), .Z(n781) );
  NANDN U686 ( .A(A[60]), .B(B[60]), .Z(n784) );
  NAND U687 ( .A(n785), .B(n786), .Z(n783) );
  NANDN U688 ( .A(B[60]), .B(A[60]), .Z(n786) );
  AND U689 ( .A(n787), .B(n788), .Z(n785) );
  NAND U690 ( .A(n789), .B(n790), .Z(n788) );
  NANDN U691 ( .A(A[59]), .B(B[59]), .Z(n790) );
  AND U692 ( .A(n791), .B(n792), .Z(n789) );
  NANDN U693 ( .A(A[58]), .B(B[58]), .Z(n792) );
  NAND U694 ( .A(n793), .B(n794), .Z(n791) );
  NANDN U695 ( .A(B[58]), .B(A[58]), .Z(n794) );
  AND U696 ( .A(n795), .B(n796), .Z(n793) );
  NAND U697 ( .A(n797), .B(n798), .Z(n796) );
  NANDN U698 ( .A(A[57]), .B(B[57]), .Z(n798) );
  AND U699 ( .A(n799), .B(n800), .Z(n797) );
  NANDN U700 ( .A(A[56]), .B(B[56]), .Z(n800) );
  NAND U701 ( .A(n801), .B(n802), .Z(n799) );
  NANDN U702 ( .A(B[56]), .B(A[56]), .Z(n802) );
  AND U703 ( .A(n803), .B(n804), .Z(n801) );
  NAND U704 ( .A(n805), .B(n806), .Z(n804) );
  NANDN U705 ( .A(A[55]), .B(B[55]), .Z(n806) );
  AND U706 ( .A(n807), .B(n808), .Z(n805) );
  NANDN U707 ( .A(A[54]), .B(B[54]), .Z(n808) );
  NAND U708 ( .A(n809), .B(n810), .Z(n807) );
  NANDN U709 ( .A(B[54]), .B(A[54]), .Z(n810) );
  AND U710 ( .A(n811), .B(n812), .Z(n809) );
  NAND U711 ( .A(n813), .B(n814), .Z(n812) );
  NANDN U712 ( .A(A[53]), .B(B[53]), .Z(n814) );
  AND U713 ( .A(n815), .B(n816), .Z(n813) );
  NANDN U714 ( .A(A[52]), .B(B[52]), .Z(n816) );
  NAND U715 ( .A(n817), .B(n818), .Z(n815) );
  NANDN U716 ( .A(B[52]), .B(A[52]), .Z(n818) );
  AND U717 ( .A(n819), .B(n820), .Z(n817) );
  NAND U718 ( .A(n821), .B(n822), .Z(n820) );
  NANDN U719 ( .A(A[51]), .B(B[51]), .Z(n822) );
  AND U720 ( .A(n823), .B(n824), .Z(n821) );
  NANDN U721 ( .A(A[50]), .B(B[50]), .Z(n824) );
  NAND U722 ( .A(n825), .B(n826), .Z(n823) );
  NANDN U723 ( .A(B[50]), .B(A[50]), .Z(n826) );
  AND U724 ( .A(n827), .B(n828), .Z(n825) );
  NAND U725 ( .A(n829), .B(n830), .Z(n828) );
  NANDN U726 ( .A(A[49]), .B(B[49]), .Z(n830) );
  AND U727 ( .A(n831), .B(n832), .Z(n829) );
  NANDN U728 ( .A(A[48]), .B(B[48]), .Z(n832) );
  NAND U729 ( .A(n833), .B(n834), .Z(n831) );
  NANDN U730 ( .A(B[48]), .B(A[48]), .Z(n834) );
  AND U731 ( .A(n835), .B(n836), .Z(n833) );
  NAND U732 ( .A(n837), .B(n838), .Z(n836) );
  NANDN U733 ( .A(A[47]), .B(B[47]), .Z(n838) );
  AND U734 ( .A(n839), .B(n840), .Z(n837) );
  NANDN U735 ( .A(A[46]), .B(B[46]), .Z(n840) );
  NAND U736 ( .A(n841), .B(n842), .Z(n839) );
  NANDN U737 ( .A(B[46]), .B(A[46]), .Z(n842) );
  AND U738 ( .A(n843), .B(n844), .Z(n841) );
  NAND U739 ( .A(n845), .B(n846), .Z(n844) );
  NANDN U740 ( .A(A[45]), .B(B[45]), .Z(n846) );
  AND U741 ( .A(n847), .B(n848), .Z(n845) );
  NANDN U742 ( .A(A[44]), .B(B[44]), .Z(n848) );
  NAND U743 ( .A(n849), .B(n850), .Z(n847) );
  NANDN U744 ( .A(B[44]), .B(A[44]), .Z(n850) );
  AND U745 ( .A(n851), .B(n852), .Z(n849) );
  NAND U746 ( .A(n853), .B(n854), .Z(n852) );
  NANDN U747 ( .A(A[43]), .B(B[43]), .Z(n854) );
  AND U748 ( .A(n855), .B(n856), .Z(n853) );
  NANDN U749 ( .A(A[42]), .B(B[42]), .Z(n856) );
  NAND U750 ( .A(n857), .B(n858), .Z(n855) );
  NANDN U751 ( .A(B[42]), .B(A[42]), .Z(n858) );
  AND U752 ( .A(n859), .B(n860), .Z(n857) );
  NAND U753 ( .A(n861), .B(n862), .Z(n860) );
  NANDN U754 ( .A(A[41]), .B(B[41]), .Z(n862) );
  AND U755 ( .A(n863), .B(n864), .Z(n861) );
  NANDN U756 ( .A(A[40]), .B(B[40]), .Z(n864) );
  NAND U757 ( .A(n865), .B(n866), .Z(n863) );
  NANDN U758 ( .A(B[40]), .B(A[40]), .Z(n866) );
  AND U759 ( .A(n867), .B(n868), .Z(n865) );
  NAND U760 ( .A(n869), .B(n870), .Z(n868) );
  NANDN U761 ( .A(A[39]), .B(B[39]), .Z(n870) );
  AND U762 ( .A(n871), .B(n872), .Z(n869) );
  NANDN U763 ( .A(A[38]), .B(B[38]), .Z(n872) );
  NAND U764 ( .A(n873), .B(n874), .Z(n871) );
  NANDN U765 ( .A(B[38]), .B(A[38]), .Z(n874) );
  AND U766 ( .A(n875), .B(n876), .Z(n873) );
  NAND U767 ( .A(n877), .B(n878), .Z(n876) );
  NANDN U768 ( .A(A[37]), .B(B[37]), .Z(n878) );
  AND U769 ( .A(n879), .B(n880), .Z(n877) );
  NANDN U770 ( .A(A[36]), .B(B[36]), .Z(n880) );
  NAND U771 ( .A(n881), .B(n882), .Z(n879) );
  NANDN U772 ( .A(B[36]), .B(A[36]), .Z(n882) );
  AND U773 ( .A(n883), .B(n884), .Z(n881) );
  NAND U774 ( .A(n885), .B(n886), .Z(n884) );
  NANDN U775 ( .A(A[35]), .B(B[35]), .Z(n886) );
  AND U776 ( .A(n887), .B(n888), .Z(n885) );
  NANDN U777 ( .A(A[34]), .B(B[34]), .Z(n888) );
  NAND U778 ( .A(n889), .B(n890), .Z(n887) );
  NANDN U779 ( .A(B[34]), .B(A[34]), .Z(n890) );
  AND U780 ( .A(n891), .B(n892), .Z(n889) );
  NAND U781 ( .A(n893), .B(n894), .Z(n892) );
  NANDN U782 ( .A(A[33]), .B(B[33]), .Z(n894) );
  AND U783 ( .A(n895), .B(n896), .Z(n893) );
  NANDN U784 ( .A(A[32]), .B(B[32]), .Z(n896) );
  NAND U785 ( .A(n897), .B(n898), .Z(n895) );
  NANDN U786 ( .A(B[32]), .B(A[32]), .Z(n898) );
  AND U787 ( .A(n899), .B(n900), .Z(n897) );
  NAND U788 ( .A(n901), .B(n902), .Z(n900) );
  NANDN U789 ( .A(A[31]), .B(B[31]), .Z(n902) );
  AND U790 ( .A(n903), .B(n904), .Z(n901) );
  NANDN U791 ( .A(A[30]), .B(B[30]), .Z(n904) );
  NAND U792 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U793 ( .A(B[30]), .B(A[30]), .Z(n906) );
  AND U794 ( .A(n907), .B(n908), .Z(n905) );
  NAND U795 ( .A(n909), .B(n910), .Z(n908) );
  NANDN U796 ( .A(A[29]), .B(B[29]), .Z(n910) );
  AND U797 ( .A(n911), .B(n912), .Z(n909) );
  NANDN U798 ( .A(A[28]), .B(B[28]), .Z(n912) );
  NAND U799 ( .A(n913), .B(n914), .Z(n911) );
  NANDN U800 ( .A(B[28]), .B(A[28]), .Z(n914) );
  AND U801 ( .A(n915), .B(n916), .Z(n913) );
  NAND U802 ( .A(n917), .B(n918), .Z(n916) );
  NANDN U803 ( .A(A[27]), .B(B[27]), .Z(n918) );
  AND U804 ( .A(n919), .B(n920), .Z(n917) );
  NANDN U805 ( .A(A[26]), .B(B[26]), .Z(n920) );
  NAND U806 ( .A(n921), .B(n922), .Z(n919) );
  NANDN U807 ( .A(B[26]), .B(A[26]), .Z(n922) );
  AND U808 ( .A(n923), .B(n924), .Z(n921) );
  NAND U809 ( .A(n925), .B(n926), .Z(n924) );
  NANDN U810 ( .A(A[25]), .B(B[25]), .Z(n926) );
  AND U811 ( .A(n927), .B(n928), .Z(n925) );
  NANDN U812 ( .A(A[24]), .B(B[24]), .Z(n928) );
  NAND U813 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U814 ( .A(B[24]), .B(A[24]), .Z(n930) );
  AND U815 ( .A(n931), .B(n932), .Z(n929) );
  NAND U816 ( .A(n933), .B(n934), .Z(n932) );
  NANDN U817 ( .A(A[23]), .B(B[23]), .Z(n934) );
  AND U818 ( .A(n935), .B(n936), .Z(n933) );
  NANDN U819 ( .A(A[22]), .B(B[22]), .Z(n936) );
  NAND U820 ( .A(n937), .B(n938), .Z(n935) );
  NANDN U821 ( .A(B[22]), .B(A[22]), .Z(n938) );
  AND U822 ( .A(n939), .B(n940), .Z(n937) );
  NAND U823 ( .A(n941), .B(n942), .Z(n940) );
  NANDN U824 ( .A(A[21]), .B(B[21]), .Z(n942) );
  AND U825 ( .A(n943), .B(n944), .Z(n941) );
  NANDN U826 ( .A(A[20]), .B(B[20]), .Z(n944) );
  NAND U827 ( .A(n945), .B(n946), .Z(n943) );
  NANDN U828 ( .A(B[20]), .B(A[20]), .Z(n946) );
  AND U829 ( .A(n947), .B(n948), .Z(n945) );
  NAND U830 ( .A(n949), .B(n950), .Z(n948) );
  NANDN U831 ( .A(A[19]), .B(B[19]), .Z(n950) );
  AND U832 ( .A(n951), .B(n952), .Z(n949) );
  NANDN U833 ( .A(A[18]), .B(B[18]), .Z(n952) );
  NAND U834 ( .A(n953), .B(n954), .Z(n951) );
  NANDN U835 ( .A(B[18]), .B(A[18]), .Z(n954) );
  AND U836 ( .A(n955), .B(n956), .Z(n953) );
  NAND U837 ( .A(n957), .B(n958), .Z(n956) );
  NANDN U838 ( .A(A[17]), .B(B[17]), .Z(n958) );
  AND U839 ( .A(n959), .B(n960), .Z(n957) );
  NANDN U840 ( .A(A[16]), .B(B[16]), .Z(n960) );
  NAND U841 ( .A(n961), .B(n962), .Z(n959) );
  NANDN U842 ( .A(B[16]), .B(A[16]), .Z(n962) );
  AND U843 ( .A(n963), .B(n964), .Z(n961) );
  NAND U844 ( .A(n965), .B(n966), .Z(n964) );
  NANDN U845 ( .A(A[15]), .B(B[15]), .Z(n966) );
  AND U846 ( .A(n967), .B(n968), .Z(n965) );
  NANDN U847 ( .A(A[14]), .B(B[14]), .Z(n968) );
  NAND U848 ( .A(n969), .B(n970), .Z(n967) );
  NANDN U849 ( .A(B[14]), .B(A[14]), .Z(n970) );
  AND U850 ( .A(n971), .B(n972), .Z(n969) );
  NAND U851 ( .A(n973), .B(n974), .Z(n972) );
  NANDN U852 ( .A(A[13]), .B(B[13]), .Z(n974) );
  AND U853 ( .A(n975), .B(n976), .Z(n973) );
  NANDN U854 ( .A(A[12]), .B(B[12]), .Z(n976) );
  NAND U855 ( .A(n977), .B(n978), .Z(n975) );
  NANDN U856 ( .A(B[12]), .B(A[12]), .Z(n978) );
  AND U857 ( .A(n979), .B(n980), .Z(n977) );
  NAND U858 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U859 ( .A(A[11]), .B(B[11]), .Z(n982) );
  AND U860 ( .A(n983), .B(n984), .Z(n981) );
  NANDN U861 ( .A(A[10]), .B(B[10]), .Z(n984) );
  NAND U862 ( .A(n985), .B(n986), .Z(n983) );
  NANDN U863 ( .A(B[9]), .B(A[9]), .Z(n986) );
  AND U864 ( .A(n987), .B(n988), .Z(n985) );
  NAND U865 ( .A(n989), .B(n990), .Z(n988) );
  NANDN U866 ( .A(A[9]), .B(B[9]), .Z(n990) );
  AND U867 ( .A(n991), .B(n992), .Z(n989) );
  NANDN U868 ( .A(A[8]), .B(B[8]), .Z(n992) );
  NAND U869 ( .A(n993), .B(n994), .Z(n991) );
  NANDN U870 ( .A(B[8]), .B(A[8]), .Z(n994) );
  AND U871 ( .A(n995), .B(n996), .Z(n993) );
  NAND U872 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U873 ( .A(A[7]), .B(B[7]), .Z(n998) );
  AND U874 ( .A(n999), .B(n1000), .Z(n997) );
  NANDN U875 ( .A(A[6]), .B(B[6]), .Z(n1000) );
  NAND U876 ( .A(n1001), .B(n1002), .Z(n999) );
  NANDN U877 ( .A(B[6]), .B(A[6]), .Z(n1002) );
  AND U878 ( .A(n1003), .B(n1004), .Z(n1001) );
  NAND U879 ( .A(n1005), .B(n1006), .Z(n1004) );
  NANDN U880 ( .A(A[5]), .B(B[5]), .Z(n1006) );
  AND U881 ( .A(n1007), .B(n1008), .Z(n1005) );
  NANDN U882 ( .A(A[4]), .B(B[4]), .Z(n1008) );
  NAND U883 ( .A(n1009), .B(n1010), .Z(n1007) );
  NANDN U884 ( .A(B[4]), .B(A[4]), .Z(n1010) );
  AND U885 ( .A(n1011), .B(n1012), .Z(n1009) );
  NAND U886 ( .A(n1013), .B(n1014), .Z(n1012) );
  NANDN U887 ( .A(A[3]), .B(B[3]), .Z(n1014) );
  AND U888 ( .A(n1015), .B(n1016), .Z(n1013) );
  NANDN U889 ( .A(A[2]), .B(B[2]), .Z(n1016) );
  NAND U890 ( .A(n1017), .B(n1018), .Z(n1015) );
  NANDN U891 ( .A(B[2]), .B(A[2]), .Z(n1018) );
  AND U892 ( .A(n1019), .B(n1020), .Z(n1017) );
  NAND U893 ( .A(n1021), .B(A[0]), .Z(n1020) );
  ANDN U894 ( .B(n1022), .A(B[0]), .Z(n1021) );
  NANDN U895 ( .A(A[1]), .B(B[1]), .Z(n1022) );
  NANDN U896 ( .A(B[1]), .B(A[1]), .Z(n1019) );
  NANDN U897 ( .A(B[3]), .B(A[3]), .Z(n1011) );
  NANDN U898 ( .A(B[5]), .B(A[5]), .Z(n1003) );
  NANDN U899 ( .A(B[7]), .B(A[7]), .Z(n995) );
  NANDN U900 ( .A(B[10]), .B(A[10]), .Z(n987) );
  NANDN U901 ( .A(B[11]), .B(A[11]), .Z(n979) );
  NANDN U902 ( .A(B[13]), .B(A[13]), .Z(n971) );
  NANDN U903 ( .A(B[15]), .B(A[15]), .Z(n963) );
  NANDN U904 ( .A(B[17]), .B(A[17]), .Z(n955) );
  NANDN U905 ( .A(B[19]), .B(A[19]), .Z(n947) );
  NANDN U906 ( .A(B[21]), .B(A[21]), .Z(n939) );
  NANDN U907 ( .A(B[23]), .B(A[23]), .Z(n931) );
  NANDN U908 ( .A(B[25]), .B(A[25]), .Z(n923) );
  NANDN U909 ( .A(B[27]), .B(A[27]), .Z(n915) );
  NANDN U910 ( .A(B[29]), .B(A[29]), .Z(n907) );
  NANDN U911 ( .A(B[31]), .B(A[31]), .Z(n899) );
  NANDN U912 ( .A(B[33]), .B(A[33]), .Z(n891) );
  NANDN U913 ( .A(B[35]), .B(A[35]), .Z(n883) );
  NANDN U914 ( .A(B[37]), .B(A[37]), .Z(n875) );
  NANDN U915 ( .A(B[39]), .B(A[39]), .Z(n867) );
  NANDN U916 ( .A(B[41]), .B(A[41]), .Z(n859) );
  NANDN U917 ( .A(B[43]), .B(A[43]), .Z(n851) );
  NANDN U918 ( .A(B[45]), .B(A[45]), .Z(n843) );
  NANDN U919 ( .A(B[47]), .B(A[47]), .Z(n835) );
  NANDN U920 ( .A(B[49]), .B(A[49]), .Z(n827) );
  NANDN U921 ( .A(B[51]), .B(A[51]), .Z(n819) );
  NANDN U922 ( .A(B[53]), .B(A[53]), .Z(n811) );
  NANDN U923 ( .A(B[55]), .B(A[55]), .Z(n803) );
  NANDN U924 ( .A(B[57]), .B(A[57]), .Z(n795) );
  NANDN U925 ( .A(B[59]), .B(A[59]), .Z(n787) );
  NANDN U926 ( .A(B[61]), .B(A[61]), .Z(n779) );
  NANDN U927 ( .A(B[63]), .B(A[63]), .Z(n771) );
  NANDN U928 ( .A(B[65]), .B(A[65]), .Z(n763) );
  NANDN U929 ( .A(B[67]), .B(A[67]), .Z(n755) );
  NANDN U930 ( .A(B[69]), .B(A[69]), .Z(n747) );
  NANDN U931 ( .A(B[71]), .B(A[71]), .Z(n739) );
  NANDN U932 ( .A(B[73]), .B(A[73]), .Z(n731) );
  NANDN U933 ( .A(B[75]), .B(A[75]), .Z(n723) );
  NANDN U934 ( .A(B[77]), .B(A[77]), .Z(n715) );
  NANDN U935 ( .A(B[79]), .B(A[79]), .Z(n707) );
  NANDN U936 ( .A(B[81]), .B(A[81]), .Z(n699) );
  NANDN U937 ( .A(B[83]), .B(A[83]), .Z(n691) );
  NANDN U938 ( .A(B[85]), .B(A[85]), .Z(n683) );
  NANDN U939 ( .A(B[87]), .B(A[87]), .Z(n675) );
  NANDN U940 ( .A(B[89]), .B(A[89]), .Z(n667) );
  NANDN U941 ( .A(B[91]), .B(A[91]), .Z(n659) );
  NANDN U942 ( .A(B[93]), .B(A[93]), .Z(n651) );
  NANDN U943 ( .A(B[95]), .B(A[95]), .Z(n643) );
  NANDN U944 ( .A(B[97]), .B(A[97]), .Z(n635) );
  NANDN U945 ( .A(B[100]), .B(A[100]), .Z(n627) );
  NANDN U946 ( .A(B[101]), .B(A[101]), .Z(n619) );
  NANDN U947 ( .A(B[103]), .B(A[103]), .Z(n611) );
  NANDN U948 ( .A(B[105]), .B(A[105]), .Z(n603) );
  NANDN U949 ( .A(B[107]), .B(A[107]), .Z(n595) );
  NANDN U950 ( .A(B[109]), .B(A[109]), .Z(n587) );
  NANDN U951 ( .A(B[111]), .B(A[111]), .Z(n579) );
  NANDN U952 ( .A(B[113]), .B(A[113]), .Z(n571) );
  NANDN U953 ( .A(B[115]), .B(A[115]), .Z(n563) );
  NANDN U954 ( .A(B[117]), .B(A[117]), .Z(n555) );
  NANDN U955 ( .A(B[119]), .B(A[119]), .Z(n547) );
  NANDN U956 ( .A(B[121]), .B(A[121]), .Z(n539) );
  NANDN U957 ( .A(B[123]), .B(A[123]), .Z(n531) );
  NANDN U958 ( .A(B[125]), .B(A[125]), .Z(n523) );
  NANDN U959 ( .A(B[127]), .B(A[127]), .Z(n515) );
  NANDN U960 ( .A(B[129]), .B(A[129]), .Z(n507) );
  NANDN U961 ( .A(B[131]), .B(A[131]), .Z(n499) );
  NANDN U962 ( .A(B[133]), .B(A[133]), .Z(n491) );
  NANDN U963 ( .A(B[135]), .B(A[135]), .Z(n483) );
  NANDN U964 ( .A(B[137]), .B(A[137]), .Z(n475) );
  NANDN U965 ( .A(B[139]), .B(A[139]), .Z(n467) );
  NANDN U966 ( .A(B[141]), .B(A[141]), .Z(n459) );
  NANDN U967 ( .A(B[143]), .B(A[143]), .Z(n451) );
  NANDN U968 ( .A(B[145]), .B(A[145]), .Z(n443) );
  NANDN U969 ( .A(B[147]), .B(A[147]), .Z(n435) );
  NANDN U970 ( .A(B[149]), .B(A[149]), .Z(n427) );
  NANDN U971 ( .A(B[151]), .B(A[151]), .Z(n419) );
  NANDN U972 ( .A(B[153]), .B(A[153]), .Z(n411) );
  NANDN U973 ( .A(B[155]), .B(A[155]), .Z(n403) );
  NANDN U974 ( .A(B[157]), .B(A[157]), .Z(n395) );
  NANDN U975 ( .A(B[159]), .B(A[159]), .Z(n387) );
  NANDN U976 ( .A(B[161]), .B(A[161]), .Z(n379) );
  NANDN U977 ( .A(B[163]), .B(A[163]), .Z(n371) );
  NANDN U978 ( .A(B[165]), .B(A[165]), .Z(n363) );
  NANDN U979 ( .A(B[167]), .B(A[167]), .Z(n355) );
  NANDN U980 ( .A(B[169]), .B(A[169]), .Z(n347) );
  NANDN U981 ( .A(B[171]), .B(A[171]), .Z(n339) );
  NANDN U982 ( .A(B[173]), .B(A[173]), .Z(n331) );
  NANDN U983 ( .A(B[175]), .B(A[175]), .Z(n323) );
  NANDN U984 ( .A(B[177]), .B(A[177]), .Z(n315) );
  NANDN U985 ( .A(B[179]), .B(A[179]), .Z(n307) );
  NANDN U986 ( .A(B[181]), .B(A[181]), .Z(n299) );
  NANDN U987 ( .A(B[183]), .B(A[183]), .Z(n291) );
  NANDN U988 ( .A(B[185]), .B(A[185]), .Z(n283) );
  NANDN U989 ( .A(B[187]), .B(A[187]), .Z(n275) );
  NANDN U990 ( .A(B[189]), .B(A[189]), .Z(n267) );
  NANDN U991 ( .A(B[191]), .B(A[191]), .Z(n259) );
  NANDN U992 ( .A(B[193]), .B(A[193]), .Z(n251) );
  NANDN U993 ( .A(B[195]), .B(A[195]), .Z(n243) );
  NANDN U994 ( .A(B[197]), .B(A[197]), .Z(n235) );
  NANDN U995 ( .A(B[199]), .B(A[199]), .Z(n227) );
  NANDN U996 ( .A(B[201]), .B(A[201]), .Z(n219) );
  NANDN U997 ( .A(B[203]), .B(A[203]), .Z(n211) );
  NANDN U998 ( .A(B[205]), .B(A[205]), .Z(n203) );
  NANDN U999 ( .A(B[207]), .B(A[207]), .Z(n195) );
  NANDN U1000 ( .A(B[209]), .B(A[209]), .Z(n187) );
  NANDN U1001 ( .A(B[211]), .B(A[211]), .Z(n179) );
  NANDN U1002 ( .A(B[213]), .B(A[213]), .Z(n171) );
  NANDN U1003 ( .A(B[215]), .B(A[215]), .Z(n163) );
  NANDN U1004 ( .A(B[217]), .B(A[217]), .Z(n155) );
  NANDN U1005 ( .A(B[219]), .B(A[219]), .Z(n147) );
  NANDN U1006 ( .A(B[221]), .B(A[221]), .Z(n139) );
  NANDN U1007 ( .A(B[223]), .B(A[223]), .Z(n131) );
  NANDN U1008 ( .A(B[225]), .B(A[225]), .Z(n123) );
  NANDN U1009 ( .A(B[227]), .B(A[227]), .Z(n115) );
  NANDN U1010 ( .A(B[229]), .B(A[229]), .Z(n107) );
  NANDN U1011 ( .A(B[231]), .B(A[231]), .Z(n99) );
  NANDN U1012 ( .A(B[233]), .B(A[233]), .Z(n91) );
  NANDN U1013 ( .A(B[235]), .B(A[235]), .Z(n83) );
  NANDN U1014 ( .A(B[237]), .B(A[237]), .Z(n75) );
  NANDN U1015 ( .A(B[239]), .B(A[239]), .Z(n67) );
  NANDN U1016 ( .A(B[241]), .B(A[241]), .Z(n59) );
  NANDN U1017 ( .A(B[243]), .B(A[243]), .Z(n51) );
  NANDN U1018 ( .A(B[245]), .B(A[245]), .Z(n43) );
  NANDN U1019 ( .A(B[247]), .B(A[247]), .Z(n35) );
  NANDN U1020 ( .A(B[249]), .B(A[249]), .Z(n27) );
  NANDN U1021 ( .A(B[251]), .B(A[251]), .Z(n19) );
  NANDN U1022 ( .A(B[253]), .B(A[253]), .Z(n11) );
  NANDN U1023 ( .A(A[255]), .B(B[255]), .Z(n3) );
endmodule


module modmult_step_N256_3_DW01_sub_1 ( A, B, CI, DIFF, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] DIFF;
  input CI;
  output CO;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280;

  IV U1 ( .A(A[1]), .Z(n1) );
  IV U2 ( .A(n1279), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(DIFF[9]) );
  XOR U4 ( .A(B[9]), .B(A[9]), .Z(n4) );
  XNOR U5 ( .A(n5), .B(n6), .Z(DIFF[99]) );
  XOR U6 ( .A(B[99]), .B(A[99]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(DIFF[98]) );
  XOR U8 ( .A(B[98]), .B(A[98]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(DIFF[97]) );
  XOR U10 ( .A(B[97]), .B(A[97]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(DIFF[96]) );
  XOR U12 ( .A(B[96]), .B(A[96]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(DIFF[95]) );
  XOR U14 ( .A(B[95]), .B(A[95]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(DIFF[94]) );
  XOR U16 ( .A(B[94]), .B(A[94]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(DIFF[93]) );
  XOR U18 ( .A(B[93]), .B(A[93]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(DIFF[92]) );
  XOR U20 ( .A(B[92]), .B(A[92]), .Z(n20) );
  XOR U21 ( .A(n21), .B(n22), .Z(DIFF[91]) );
  XOR U22 ( .A(B[91]), .B(A[91]), .Z(n22) );
  XOR U23 ( .A(n23), .B(n24), .Z(DIFF[90]) );
  XOR U24 ( .A(B[90]), .B(A[90]), .Z(n24) );
  XOR U25 ( .A(n25), .B(n26), .Z(DIFF[8]) );
  XOR U26 ( .A(B[8]), .B(A[8]), .Z(n26) );
  XOR U27 ( .A(n27), .B(n28), .Z(DIFF[89]) );
  XOR U28 ( .A(B[89]), .B(A[89]), .Z(n28) );
  XOR U29 ( .A(n29), .B(n30), .Z(DIFF[88]) );
  XOR U30 ( .A(B[88]), .B(A[88]), .Z(n30) );
  XOR U31 ( .A(n31), .B(n32), .Z(DIFF[87]) );
  XOR U32 ( .A(B[87]), .B(A[87]), .Z(n32) );
  XOR U33 ( .A(n33), .B(n34), .Z(DIFF[86]) );
  XOR U34 ( .A(B[86]), .B(A[86]), .Z(n34) );
  XOR U35 ( .A(n35), .B(n36), .Z(DIFF[85]) );
  XOR U36 ( .A(B[85]), .B(A[85]), .Z(n36) );
  XOR U37 ( .A(n37), .B(n38), .Z(DIFF[84]) );
  XOR U38 ( .A(B[84]), .B(A[84]), .Z(n38) );
  XOR U39 ( .A(n39), .B(n40), .Z(DIFF[83]) );
  XOR U40 ( .A(B[83]), .B(A[83]), .Z(n40) );
  XOR U41 ( .A(n41), .B(n42), .Z(DIFF[82]) );
  XOR U42 ( .A(B[82]), .B(A[82]), .Z(n42) );
  XOR U43 ( .A(n43), .B(n44), .Z(DIFF[81]) );
  XOR U44 ( .A(B[81]), .B(A[81]), .Z(n44) );
  XOR U45 ( .A(n45), .B(n46), .Z(DIFF[80]) );
  XOR U46 ( .A(B[80]), .B(A[80]), .Z(n46) );
  XOR U47 ( .A(n47), .B(n48), .Z(DIFF[7]) );
  XOR U48 ( .A(B[7]), .B(A[7]), .Z(n48) );
  XOR U49 ( .A(n49), .B(n50), .Z(DIFF[79]) );
  XOR U50 ( .A(B[79]), .B(A[79]), .Z(n50) );
  XOR U51 ( .A(n51), .B(n52), .Z(DIFF[78]) );
  XOR U52 ( .A(B[78]), .B(A[78]), .Z(n52) );
  XOR U53 ( .A(n53), .B(n54), .Z(DIFF[77]) );
  XOR U54 ( .A(B[77]), .B(A[77]), .Z(n54) );
  XOR U55 ( .A(n55), .B(n56), .Z(DIFF[76]) );
  XOR U56 ( .A(B[76]), .B(A[76]), .Z(n56) );
  XOR U57 ( .A(n57), .B(n58), .Z(DIFF[75]) );
  XOR U58 ( .A(B[75]), .B(A[75]), .Z(n58) );
  XOR U59 ( .A(n59), .B(n60), .Z(DIFF[74]) );
  XOR U60 ( .A(B[74]), .B(A[74]), .Z(n60) );
  XOR U61 ( .A(n61), .B(n62), .Z(DIFF[73]) );
  XOR U62 ( .A(B[73]), .B(A[73]), .Z(n62) );
  XOR U63 ( .A(n63), .B(n64), .Z(DIFF[72]) );
  XOR U64 ( .A(B[72]), .B(A[72]), .Z(n64) );
  XOR U65 ( .A(n65), .B(n66), .Z(DIFF[71]) );
  XOR U66 ( .A(B[71]), .B(A[71]), .Z(n66) );
  XOR U67 ( .A(n67), .B(n68), .Z(DIFF[70]) );
  XOR U68 ( .A(B[70]), .B(A[70]), .Z(n68) );
  XOR U69 ( .A(n69), .B(n70), .Z(DIFF[6]) );
  XOR U70 ( .A(B[6]), .B(A[6]), .Z(n70) );
  XOR U71 ( .A(n71), .B(n72), .Z(DIFF[69]) );
  XOR U72 ( .A(B[69]), .B(A[69]), .Z(n72) );
  XOR U73 ( .A(n73), .B(n74), .Z(DIFF[68]) );
  XOR U74 ( .A(B[68]), .B(A[68]), .Z(n74) );
  XOR U75 ( .A(n75), .B(n76), .Z(DIFF[67]) );
  XOR U76 ( .A(B[67]), .B(A[67]), .Z(n76) );
  XOR U77 ( .A(n77), .B(n78), .Z(DIFF[66]) );
  XOR U78 ( .A(B[66]), .B(A[66]), .Z(n78) );
  XOR U79 ( .A(n79), .B(n80), .Z(DIFF[65]) );
  XOR U80 ( .A(B[65]), .B(A[65]), .Z(n80) );
  XOR U81 ( .A(n81), .B(n82), .Z(DIFF[64]) );
  XOR U82 ( .A(B[64]), .B(A[64]), .Z(n82) );
  XOR U83 ( .A(n83), .B(n84), .Z(DIFF[63]) );
  XOR U84 ( .A(B[63]), .B(A[63]), .Z(n84) );
  XOR U85 ( .A(n85), .B(n86), .Z(DIFF[62]) );
  XOR U86 ( .A(B[62]), .B(A[62]), .Z(n86) );
  XOR U87 ( .A(n87), .B(n88), .Z(DIFF[61]) );
  XOR U88 ( .A(B[61]), .B(A[61]), .Z(n88) );
  XOR U89 ( .A(n89), .B(n90), .Z(DIFF[60]) );
  XOR U90 ( .A(B[60]), .B(A[60]), .Z(n90) );
  XOR U91 ( .A(n91), .B(n92), .Z(DIFF[5]) );
  XOR U92 ( .A(B[5]), .B(A[5]), .Z(n92) );
  XOR U93 ( .A(n93), .B(n94), .Z(DIFF[59]) );
  XOR U94 ( .A(B[59]), .B(A[59]), .Z(n94) );
  XOR U95 ( .A(n95), .B(n96), .Z(DIFF[58]) );
  XOR U96 ( .A(B[58]), .B(A[58]), .Z(n96) );
  XOR U97 ( .A(n97), .B(n98), .Z(DIFF[57]) );
  XOR U98 ( .A(B[57]), .B(A[57]), .Z(n98) );
  XOR U99 ( .A(n99), .B(n100), .Z(DIFF[56]) );
  XOR U100 ( .A(B[56]), .B(A[56]), .Z(n100) );
  XOR U101 ( .A(n101), .B(n102), .Z(DIFF[55]) );
  XOR U102 ( .A(B[55]), .B(A[55]), .Z(n102) );
  XOR U103 ( .A(n103), .B(n104), .Z(DIFF[54]) );
  XOR U104 ( .A(B[54]), .B(A[54]), .Z(n104) );
  XOR U105 ( .A(n105), .B(n106), .Z(DIFF[53]) );
  XOR U106 ( .A(B[53]), .B(A[53]), .Z(n106) );
  XOR U107 ( .A(n107), .B(n108), .Z(DIFF[52]) );
  XOR U108 ( .A(B[52]), .B(A[52]), .Z(n108) );
  XOR U109 ( .A(n109), .B(n110), .Z(DIFF[51]) );
  XOR U110 ( .A(B[51]), .B(A[51]), .Z(n110) );
  XOR U111 ( .A(n111), .B(n112), .Z(DIFF[50]) );
  XOR U112 ( .A(B[50]), .B(A[50]), .Z(n112) );
  XOR U113 ( .A(n113), .B(n114), .Z(DIFF[4]) );
  XOR U114 ( .A(B[4]), .B(A[4]), .Z(n114) );
  XOR U115 ( .A(n115), .B(n116), .Z(DIFF[49]) );
  XOR U116 ( .A(B[49]), .B(A[49]), .Z(n116) );
  XOR U117 ( .A(n117), .B(n118), .Z(DIFF[48]) );
  XOR U118 ( .A(B[48]), .B(A[48]), .Z(n118) );
  XOR U119 ( .A(n119), .B(n120), .Z(DIFF[47]) );
  XOR U120 ( .A(B[47]), .B(A[47]), .Z(n120) );
  XOR U121 ( .A(n121), .B(n122), .Z(DIFF[46]) );
  XOR U122 ( .A(B[46]), .B(A[46]), .Z(n122) );
  XOR U123 ( .A(n123), .B(n124), .Z(DIFF[45]) );
  XOR U124 ( .A(B[45]), .B(A[45]), .Z(n124) );
  XOR U125 ( .A(n125), .B(n126), .Z(DIFF[44]) );
  XOR U126 ( .A(B[44]), .B(A[44]), .Z(n126) );
  XOR U127 ( .A(n127), .B(n128), .Z(DIFF[43]) );
  XOR U128 ( .A(B[43]), .B(A[43]), .Z(n128) );
  XOR U129 ( .A(n129), .B(n130), .Z(DIFF[42]) );
  XOR U130 ( .A(B[42]), .B(A[42]), .Z(n130) );
  XOR U131 ( .A(n131), .B(n132), .Z(DIFF[41]) );
  XOR U132 ( .A(B[41]), .B(A[41]), .Z(n132) );
  XOR U133 ( .A(n133), .B(n134), .Z(DIFF[40]) );
  XOR U134 ( .A(B[40]), .B(A[40]), .Z(n134) );
  XOR U135 ( .A(n135), .B(n136), .Z(DIFF[3]) );
  XOR U136 ( .A(B[3]), .B(A[3]), .Z(n136) );
  XOR U137 ( .A(n137), .B(n138), .Z(DIFF[39]) );
  XOR U138 ( .A(B[39]), .B(A[39]), .Z(n138) );
  XOR U139 ( .A(n139), .B(n140), .Z(DIFF[38]) );
  XOR U140 ( .A(B[38]), .B(A[38]), .Z(n140) );
  XOR U141 ( .A(n141), .B(n142), .Z(DIFF[37]) );
  XOR U142 ( .A(B[37]), .B(A[37]), .Z(n142) );
  XOR U143 ( .A(n143), .B(n144), .Z(DIFF[36]) );
  XOR U144 ( .A(B[36]), .B(A[36]), .Z(n144) );
  XOR U145 ( .A(n145), .B(n146), .Z(DIFF[35]) );
  XOR U146 ( .A(B[35]), .B(A[35]), .Z(n146) );
  XOR U147 ( .A(n147), .B(n148), .Z(DIFF[34]) );
  XOR U148 ( .A(B[34]), .B(A[34]), .Z(n148) );
  XOR U149 ( .A(n149), .B(n150), .Z(DIFF[33]) );
  XOR U150 ( .A(B[33]), .B(A[33]), .Z(n150) );
  XOR U151 ( .A(n151), .B(n152), .Z(DIFF[32]) );
  XOR U152 ( .A(B[32]), .B(A[32]), .Z(n152) );
  XOR U153 ( .A(n153), .B(n154), .Z(DIFF[31]) );
  XOR U154 ( .A(B[31]), .B(A[31]), .Z(n154) );
  XOR U155 ( .A(n155), .B(n156), .Z(DIFF[30]) );
  XOR U156 ( .A(B[30]), .B(A[30]), .Z(n156) );
  XOR U157 ( .A(n157), .B(n158), .Z(DIFF[2]) );
  XOR U158 ( .A(B[2]), .B(A[2]), .Z(n158) );
  XOR U159 ( .A(n159), .B(n160), .Z(DIFF[29]) );
  XOR U160 ( .A(B[29]), .B(A[29]), .Z(n160) );
  XOR U161 ( .A(n161), .B(n162), .Z(DIFF[28]) );
  XOR U162 ( .A(B[28]), .B(A[28]), .Z(n162) );
  XOR U163 ( .A(n163), .B(n164), .Z(DIFF[27]) );
  XOR U164 ( .A(B[27]), .B(A[27]), .Z(n164) );
  XOR U165 ( .A(n165), .B(n166), .Z(DIFF[26]) );
  XOR U166 ( .A(B[26]), .B(A[26]), .Z(n166) );
  XOR U167 ( .A(n167), .B(n168), .Z(DIFF[25]) );
  XOR U168 ( .A(B[25]), .B(A[25]), .Z(n168) );
  XOR U169 ( .A(A[257]), .B(n169), .Z(DIFF[257]) );
  ANDN U170 ( .B(n170), .A(A[256]), .Z(n169) );
  XOR U171 ( .A(A[256]), .B(n170), .Z(DIFF[256]) );
  AND U172 ( .A(n171), .B(n172), .Z(n170) );
  NANDN U173 ( .A(B[255]), .B(n173), .Z(n172) );
  NANDN U174 ( .A(A[255]), .B(n174), .Z(n173) );
  NANDN U175 ( .A(n174), .B(A[255]), .Z(n171) );
  XOR U176 ( .A(n174), .B(n175), .Z(DIFF[255]) );
  XOR U177 ( .A(B[255]), .B(A[255]), .Z(n175) );
  AND U178 ( .A(n176), .B(n177), .Z(n174) );
  NANDN U179 ( .A(B[254]), .B(n178), .Z(n177) );
  NANDN U180 ( .A(A[254]), .B(n179), .Z(n178) );
  NANDN U181 ( .A(n179), .B(A[254]), .Z(n176) );
  XOR U182 ( .A(n179), .B(n180), .Z(DIFF[254]) );
  XOR U183 ( .A(B[254]), .B(A[254]), .Z(n180) );
  AND U184 ( .A(n181), .B(n182), .Z(n179) );
  NANDN U185 ( .A(B[253]), .B(n183), .Z(n182) );
  NANDN U186 ( .A(A[253]), .B(n184), .Z(n183) );
  NANDN U187 ( .A(n184), .B(A[253]), .Z(n181) );
  XOR U188 ( .A(n184), .B(n185), .Z(DIFF[253]) );
  XOR U189 ( .A(B[253]), .B(A[253]), .Z(n185) );
  AND U190 ( .A(n186), .B(n187), .Z(n184) );
  NANDN U191 ( .A(B[252]), .B(n188), .Z(n187) );
  NANDN U192 ( .A(A[252]), .B(n189), .Z(n188) );
  NANDN U193 ( .A(n189), .B(A[252]), .Z(n186) );
  XOR U194 ( .A(n189), .B(n190), .Z(DIFF[252]) );
  XOR U195 ( .A(B[252]), .B(A[252]), .Z(n190) );
  AND U196 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U197 ( .A(B[251]), .B(n193), .Z(n192) );
  NANDN U198 ( .A(A[251]), .B(n194), .Z(n193) );
  NANDN U199 ( .A(n194), .B(A[251]), .Z(n191) );
  XOR U200 ( .A(n194), .B(n195), .Z(DIFF[251]) );
  XOR U201 ( .A(B[251]), .B(A[251]), .Z(n195) );
  AND U202 ( .A(n196), .B(n197), .Z(n194) );
  NANDN U203 ( .A(B[250]), .B(n198), .Z(n197) );
  NANDN U204 ( .A(A[250]), .B(n199), .Z(n198) );
  NANDN U205 ( .A(n199), .B(A[250]), .Z(n196) );
  XOR U206 ( .A(n199), .B(n200), .Z(DIFF[250]) );
  XOR U207 ( .A(B[250]), .B(A[250]), .Z(n200) );
  AND U208 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U209 ( .A(B[249]), .B(n203), .Z(n202) );
  NANDN U210 ( .A(A[249]), .B(n204), .Z(n203) );
  NANDN U211 ( .A(n204), .B(A[249]), .Z(n201) );
  XOR U212 ( .A(n205), .B(n206), .Z(DIFF[24]) );
  XOR U213 ( .A(B[24]), .B(A[24]), .Z(n206) );
  XOR U214 ( .A(n204), .B(n207), .Z(DIFF[249]) );
  XOR U215 ( .A(B[249]), .B(A[249]), .Z(n207) );
  AND U216 ( .A(n208), .B(n209), .Z(n204) );
  NANDN U217 ( .A(B[248]), .B(n210), .Z(n209) );
  NANDN U218 ( .A(A[248]), .B(n211), .Z(n210) );
  NANDN U219 ( .A(n211), .B(A[248]), .Z(n208) );
  XOR U220 ( .A(n211), .B(n212), .Z(DIFF[248]) );
  XOR U221 ( .A(B[248]), .B(A[248]), .Z(n212) );
  AND U222 ( .A(n213), .B(n214), .Z(n211) );
  NANDN U223 ( .A(B[247]), .B(n215), .Z(n214) );
  NANDN U224 ( .A(A[247]), .B(n216), .Z(n215) );
  NANDN U225 ( .A(n216), .B(A[247]), .Z(n213) );
  XOR U226 ( .A(n216), .B(n217), .Z(DIFF[247]) );
  XOR U227 ( .A(B[247]), .B(A[247]), .Z(n217) );
  AND U228 ( .A(n218), .B(n219), .Z(n216) );
  NANDN U229 ( .A(B[246]), .B(n220), .Z(n219) );
  NANDN U230 ( .A(A[246]), .B(n221), .Z(n220) );
  NANDN U231 ( .A(n221), .B(A[246]), .Z(n218) );
  XOR U232 ( .A(n221), .B(n222), .Z(DIFF[246]) );
  XOR U233 ( .A(B[246]), .B(A[246]), .Z(n222) );
  AND U234 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U235 ( .A(B[245]), .B(n225), .Z(n224) );
  NANDN U236 ( .A(A[245]), .B(n226), .Z(n225) );
  NANDN U237 ( .A(n226), .B(A[245]), .Z(n223) );
  XOR U238 ( .A(n226), .B(n227), .Z(DIFF[245]) );
  XOR U239 ( .A(B[245]), .B(A[245]), .Z(n227) );
  AND U240 ( .A(n228), .B(n229), .Z(n226) );
  NANDN U241 ( .A(B[244]), .B(n230), .Z(n229) );
  NANDN U242 ( .A(A[244]), .B(n231), .Z(n230) );
  NANDN U243 ( .A(n231), .B(A[244]), .Z(n228) );
  XOR U244 ( .A(n231), .B(n232), .Z(DIFF[244]) );
  XOR U245 ( .A(B[244]), .B(A[244]), .Z(n232) );
  AND U246 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U247 ( .A(B[243]), .B(n235), .Z(n234) );
  NANDN U248 ( .A(A[243]), .B(n236), .Z(n235) );
  NANDN U249 ( .A(n236), .B(A[243]), .Z(n233) );
  XOR U250 ( .A(n236), .B(n237), .Z(DIFF[243]) );
  XOR U251 ( .A(B[243]), .B(A[243]), .Z(n237) );
  AND U252 ( .A(n238), .B(n239), .Z(n236) );
  NANDN U253 ( .A(B[242]), .B(n240), .Z(n239) );
  NANDN U254 ( .A(A[242]), .B(n241), .Z(n240) );
  NANDN U255 ( .A(n241), .B(A[242]), .Z(n238) );
  XOR U256 ( .A(n241), .B(n242), .Z(DIFF[242]) );
  XOR U257 ( .A(B[242]), .B(A[242]), .Z(n242) );
  AND U258 ( .A(n243), .B(n244), .Z(n241) );
  NANDN U259 ( .A(B[241]), .B(n245), .Z(n244) );
  NANDN U260 ( .A(A[241]), .B(n246), .Z(n245) );
  NANDN U261 ( .A(n246), .B(A[241]), .Z(n243) );
  XOR U262 ( .A(n246), .B(n247), .Z(DIFF[241]) );
  XOR U263 ( .A(B[241]), .B(A[241]), .Z(n247) );
  AND U264 ( .A(n248), .B(n249), .Z(n246) );
  NANDN U265 ( .A(B[240]), .B(n250), .Z(n249) );
  NANDN U266 ( .A(A[240]), .B(n251), .Z(n250) );
  NANDN U267 ( .A(n251), .B(A[240]), .Z(n248) );
  XOR U268 ( .A(n251), .B(n252), .Z(DIFF[240]) );
  XOR U269 ( .A(B[240]), .B(A[240]), .Z(n252) );
  AND U270 ( .A(n253), .B(n254), .Z(n251) );
  NANDN U271 ( .A(B[239]), .B(n255), .Z(n254) );
  NANDN U272 ( .A(A[239]), .B(n256), .Z(n255) );
  NANDN U273 ( .A(n256), .B(A[239]), .Z(n253) );
  XOR U274 ( .A(n257), .B(n258), .Z(DIFF[23]) );
  XOR U275 ( .A(B[23]), .B(A[23]), .Z(n258) );
  XOR U276 ( .A(n256), .B(n259), .Z(DIFF[239]) );
  XOR U277 ( .A(B[239]), .B(A[239]), .Z(n259) );
  AND U278 ( .A(n260), .B(n261), .Z(n256) );
  NANDN U279 ( .A(B[238]), .B(n262), .Z(n261) );
  NANDN U280 ( .A(A[238]), .B(n263), .Z(n262) );
  NANDN U281 ( .A(n263), .B(A[238]), .Z(n260) );
  XOR U282 ( .A(n263), .B(n264), .Z(DIFF[238]) );
  XOR U283 ( .A(B[238]), .B(A[238]), .Z(n264) );
  AND U284 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U285 ( .A(B[237]), .B(n267), .Z(n266) );
  NANDN U286 ( .A(A[237]), .B(n268), .Z(n267) );
  NANDN U287 ( .A(n268), .B(A[237]), .Z(n265) );
  XOR U288 ( .A(n268), .B(n269), .Z(DIFF[237]) );
  XOR U289 ( .A(B[237]), .B(A[237]), .Z(n269) );
  AND U290 ( .A(n270), .B(n271), .Z(n268) );
  NANDN U291 ( .A(B[236]), .B(n272), .Z(n271) );
  NANDN U292 ( .A(A[236]), .B(n273), .Z(n272) );
  NANDN U293 ( .A(n273), .B(A[236]), .Z(n270) );
  XOR U294 ( .A(n273), .B(n274), .Z(DIFF[236]) );
  XOR U295 ( .A(B[236]), .B(A[236]), .Z(n274) );
  AND U296 ( .A(n275), .B(n276), .Z(n273) );
  NANDN U297 ( .A(B[235]), .B(n277), .Z(n276) );
  NANDN U298 ( .A(A[235]), .B(n278), .Z(n277) );
  NANDN U299 ( .A(n278), .B(A[235]), .Z(n275) );
  XOR U300 ( .A(n278), .B(n279), .Z(DIFF[235]) );
  XOR U301 ( .A(B[235]), .B(A[235]), .Z(n279) );
  AND U302 ( .A(n280), .B(n281), .Z(n278) );
  NANDN U303 ( .A(B[234]), .B(n282), .Z(n281) );
  NANDN U304 ( .A(A[234]), .B(n283), .Z(n282) );
  NANDN U305 ( .A(n283), .B(A[234]), .Z(n280) );
  XOR U306 ( .A(n283), .B(n284), .Z(DIFF[234]) );
  XOR U307 ( .A(B[234]), .B(A[234]), .Z(n284) );
  AND U308 ( .A(n285), .B(n286), .Z(n283) );
  NANDN U309 ( .A(B[233]), .B(n287), .Z(n286) );
  NANDN U310 ( .A(A[233]), .B(n288), .Z(n287) );
  NANDN U311 ( .A(n288), .B(A[233]), .Z(n285) );
  XOR U312 ( .A(n288), .B(n289), .Z(DIFF[233]) );
  XOR U313 ( .A(B[233]), .B(A[233]), .Z(n289) );
  AND U314 ( .A(n290), .B(n291), .Z(n288) );
  NANDN U315 ( .A(B[232]), .B(n292), .Z(n291) );
  NANDN U316 ( .A(A[232]), .B(n293), .Z(n292) );
  NANDN U317 ( .A(n293), .B(A[232]), .Z(n290) );
  XOR U318 ( .A(n293), .B(n294), .Z(DIFF[232]) );
  XOR U319 ( .A(B[232]), .B(A[232]), .Z(n294) );
  AND U320 ( .A(n295), .B(n296), .Z(n293) );
  NANDN U321 ( .A(B[231]), .B(n297), .Z(n296) );
  NANDN U322 ( .A(A[231]), .B(n298), .Z(n297) );
  NANDN U323 ( .A(n298), .B(A[231]), .Z(n295) );
  XOR U324 ( .A(n298), .B(n299), .Z(DIFF[231]) );
  XOR U325 ( .A(B[231]), .B(A[231]), .Z(n299) );
  AND U326 ( .A(n300), .B(n301), .Z(n298) );
  NANDN U327 ( .A(B[230]), .B(n302), .Z(n301) );
  NANDN U328 ( .A(A[230]), .B(n303), .Z(n302) );
  NANDN U329 ( .A(n303), .B(A[230]), .Z(n300) );
  XOR U330 ( .A(n303), .B(n304), .Z(DIFF[230]) );
  XOR U331 ( .A(B[230]), .B(A[230]), .Z(n304) );
  AND U332 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U333 ( .A(B[229]), .B(n307), .Z(n306) );
  NANDN U334 ( .A(A[229]), .B(n308), .Z(n307) );
  NANDN U335 ( .A(n308), .B(A[229]), .Z(n305) );
  XOR U336 ( .A(n309), .B(n310), .Z(DIFF[22]) );
  XOR U337 ( .A(B[22]), .B(A[22]), .Z(n310) );
  XOR U338 ( .A(n308), .B(n311), .Z(DIFF[229]) );
  XOR U339 ( .A(B[229]), .B(A[229]), .Z(n311) );
  AND U340 ( .A(n312), .B(n313), .Z(n308) );
  NANDN U341 ( .A(B[228]), .B(n314), .Z(n313) );
  NANDN U342 ( .A(A[228]), .B(n315), .Z(n314) );
  NANDN U343 ( .A(n315), .B(A[228]), .Z(n312) );
  XOR U344 ( .A(n315), .B(n316), .Z(DIFF[228]) );
  XOR U345 ( .A(B[228]), .B(A[228]), .Z(n316) );
  AND U346 ( .A(n317), .B(n318), .Z(n315) );
  NANDN U347 ( .A(B[227]), .B(n319), .Z(n318) );
  NANDN U348 ( .A(A[227]), .B(n320), .Z(n319) );
  NANDN U349 ( .A(n320), .B(A[227]), .Z(n317) );
  XOR U350 ( .A(n320), .B(n321), .Z(DIFF[227]) );
  XOR U351 ( .A(B[227]), .B(A[227]), .Z(n321) );
  AND U352 ( .A(n322), .B(n323), .Z(n320) );
  NANDN U353 ( .A(B[226]), .B(n324), .Z(n323) );
  NANDN U354 ( .A(A[226]), .B(n325), .Z(n324) );
  NANDN U355 ( .A(n325), .B(A[226]), .Z(n322) );
  XOR U356 ( .A(n325), .B(n326), .Z(DIFF[226]) );
  XOR U357 ( .A(B[226]), .B(A[226]), .Z(n326) );
  AND U358 ( .A(n327), .B(n328), .Z(n325) );
  NANDN U359 ( .A(B[225]), .B(n329), .Z(n328) );
  NANDN U360 ( .A(A[225]), .B(n330), .Z(n329) );
  NANDN U361 ( .A(n330), .B(A[225]), .Z(n327) );
  XOR U362 ( .A(n330), .B(n331), .Z(DIFF[225]) );
  XOR U363 ( .A(B[225]), .B(A[225]), .Z(n331) );
  AND U364 ( .A(n332), .B(n333), .Z(n330) );
  NANDN U365 ( .A(B[224]), .B(n334), .Z(n333) );
  NANDN U366 ( .A(A[224]), .B(n335), .Z(n334) );
  NANDN U367 ( .A(n335), .B(A[224]), .Z(n332) );
  XOR U368 ( .A(n335), .B(n336), .Z(DIFF[224]) );
  XOR U369 ( .A(B[224]), .B(A[224]), .Z(n336) );
  AND U370 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U371 ( .A(B[223]), .B(n339), .Z(n338) );
  NANDN U372 ( .A(A[223]), .B(n340), .Z(n339) );
  NANDN U373 ( .A(n340), .B(A[223]), .Z(n337) );
  XOR U374 ( .A(n340), .B(n341), .Z(DIFF[223]) );
  XOR U375 ( .A(B[223]), .B(A[223]), .Z(n341) );
  AND U376 ( .A(n342), .B(n343), .Z(n340) );
  NANDN U377 ( .A(B[222]), .B(n344), .Z(n343) );
  NANDN U378 ( .A(A[222]), .B(n345), .Z(n344) );
  NANDN U379 ( .A(n345), .B(A[222]), .Z(n342) );
  XOR U380 ( .A(n345), .B(n346), .Z(DIFF[222]) );
  XOR U381 ( .A(B[222]), .B(A[222]), .Z(n346) );
  AND U382 ( .A(n347), .B(n348), .Z(n345) );
  NANDN U383 ( .A(B[221]), .B(n349), .Z(n348) );
  NANDN U384 ( .A(A[221]), .B(n350), .Z(n349) );
  NANDN U385 ( .A(n350), .B(A[221]), .Z(n347) );
  XOR U386 ( .A(n350), .B(n351), .Z(DIFF[221]) );
  XOR U387 ( .A(B[221]), .B(A[221]), .Z(n351) );
  AND U388 ( .A(n352), .B(n353), .Z(n350) );
  NANDN U389 ( .A(B[220]), .B(n354), .Z(n353) );
  NANDN U390 ( .A(A[220]), .B(n355), .Z(n354) );
  NANDN U391 ( .A(n355), .B(A[220]), .Z(n352) );
  XOR U392 ( .A(n355), .B(n356), .Z(DIFF[220]) );
  XOR U393 ( .A(B[220]), .B(A[220]), .Z(n356) );
  AND U394 ( .A(n357), .B(n358), .Z(n355) );
  NANDN U395 ( .A(B[219]), .B(n359), .Z(n358) );
  NANDN U396 ( .A(A[219]), .B(n360), .Z(n359) );
  NANDN U397 ( .A(n360), .B(A[219]), .Z(n357) );
  XOR U398 ( .A(n361), .B(n362), .Z(DIFF[21]) );
  XOR U399 ( .A(B[21]), .B(A[21]), .Z(n362) );
  XOR U400 ( .A(n360), .B(n363), .Z(DIFF[219]) );
  XOR U401 ( .A(B[219]), .B(A[219]), .Z(n363) );
  AND U402 ( .A(n364), .B(n365), .Z(n360) );
  NANDN U403 ( .A(B[218]), .B(n366), .Z(n365) );
  NANDN U404 ( .A(A[218]), .B(n367), .Z(n366) );
  NANDN U405 ( .A(n367), .B(A[218]), .Z(n364) );
  XOR U406 ( .A(n367), .B(n368), .Z(DIFF[218]) );
  XOR U407 ( .A(B[218]), .B(A[218]), .Z(n368) );
  AND U408 ( .A(n369), .B(n370), .Z(n367) );
  NANDN U409 ( .A(B[217]), .B(n371), .Z(n370) );
  NANDN U410 ( .A(A[217]), .B(n372), .Z(n371) );
  NANDN U411 ( .A(n372), .B(A[217]), .Z(n369) );
  XOR U412 ( .A(n372), .B(n373), .Z(DIFF[217]) );
  XOR U413 ( .A(B[217]), .B(A[217]), .Z(n373) );
  AND U414 ( .A(n374), .B(n375), .Z(n372) );
  NANDN U415 ( .A(B[216]), .B(n376), .Z(n375) );
  NANDN U416 ( .A(A[216]), .B(n377), .Z(n376) );
  NANDN U417 ( .A(n377), .B(A[216]), .Z(n374) );
  XOR U418 ( .A(n377), .B(n378), .Z(DIFF[216]) );
  XOR U419 ( .A(B[216]), .B(A[216]), .Z(n378) );
  AND U420 ( .A(n379), .B(n380), .Z(n377) );
  NANDN U421 ( .A(B[215]), .B(n381), .Z(n380) );
  NANDN U422 ( .A(A[215]), .B(n382), .Z(n381) );
  NANDN U423 ( .A(n382), .B(A[215]), .Z(n379) );
  XOR U424 ( .A(n382), .B(n383), .Z(DIFF[215]) );
  XOR U425 ( .A(B[215]), .B(A[215]), .Z(n383) );
  AND U426 ( .A(n384), .B(n385), .Z(n382) );
  NANDN U427 ( .A(B[214]), .B(n386), .Z(n385) );
  NANDN U428 ( .A(A[214]), .B(n387), .Z(n386) );
  NANDN U429 ( .A(n387), .B(A[214]), .Z(n384) );
  XOR U430 ( .A(n387), .B(n388), .Z(DIFF[214]) );
  XOR U431 ( .A(B[214]), .B(A[214]), .Z(n388) );
  AND U432 ( .A(n389), .B(n390), .Z(n387) );
  NANDN U433 ( .A(B[213]), .B(n391), .Z(n390) );
  NANDN U434 ( .A(A[213]), .B(n392), .Z(n391) );
  NANDN U435 ( .A(n392), .B(A[213]), .Z(n389) );
  XOR U436 ( .A(n392), .B(n393), .Z(DIFF[213]) );
  XOR U437 ( .A(B[213]), .B(A[213]), .Z(n393) );
  AND U438 ( .A(n394), .B(n395), .Z(n392) );
  NANDN U439 ( .A(B[212]), .B(n396), .Z(n395) );
  NANDN U440 ( .A(A[212]), .B(n397), .Z(n396) );
  NANDN U441 ( .A(n397), .B(A[212]), .Z(n394) );
  XOR U442 ( .A(n397), .B(n398), .Z(DIFF[212]) );
  XOR U443 ( .A(B[212]), .B(A[212]), .Z(n398) );
  AND U444 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U445 ( .A(B[211]), .B(n401), .Z(n400) );
  NANDN U446 ( .A(A[211]), .B(n402), .Z(n401) );
  NANDN U447 ( .A(n402), .B(A[211]), .Z(n399) );
  XOR U448 ( .A(n402), .B(n403), .Z(DIFF[211]) );
  XOR U449 ( .A(B[211]), .B(A[211]), .Z(n403) );
  AND U450 ( .A(n404), .B(n405), .Z(n402) );
  NANDN U451 ( .A(B[210]), .B(n406), .Z(n405) );
  NANDN U452 ( .A(A[210]), .B(n407), .Z(n406) );
  NANDN U453 ( .A(n407), .B(A[210]), .Z(n404) );
  XOR U454 ( .A(n407), .B(n408), .Z(DIFF[210]) );
  XOR U455 ( .A(B[210]), .B(A[210]), .Z(n408) );
  AND U456 ( .A(n409), .B(n410), .Z(n407) );
  NANDN U457 ( .A(B[209]), .B(n411), .Z(n410) );
  NANDN U458 ( .A(A[209]), .B(n412), .Z(n411) );
  NANDN U459 ( .A(n412), .B(A[209]), .Z(n409) );
  XOR U460 ( .A(n413), .B(n414), .Z(DIFF[20]) );
  XOR U461 ( .A(B[20]), .B(A[20]), .Z(n414) );
  XOR U462 ( .A(n412), .B(n415), .Z(DIFF[209]) );
  XOR U463 ( .A(B[209]), .B(A[209]), .Z(n415) );
  AND U464 ( .A(n416), .B(n417), .Z(n412) );
  NANDN U465 ( .A(B[208]), .B(n418), .Z(n417) );
  NANDN U466 ( .A(A[208]), .B(n419), .Z(n418) );
  NANDN U467 ( .A(n419), .B(A[208]), .Z(n416) );
  XOR U468 ( .A(n419), .B(n420), .Z(DIFF[208]) );
  XOR U469 ( .A(B[208]), .B(A[208]), .Z(n420) );
  AND U470 ( .A(n421), .B(n422), .Z(n419) );
  NANDN U471 ( .A(B[207]), .B(n423), .Z(n422) );
  NANDN U472 ( .A(A[207]), .B(n424), .Z(n423) );
  NANDN U473 ( .A(n424), .B(A[207]), .Z(n421) );
  XOR U474 ( .A(n424), .B(n425), .Z(DIFF[207]) );
  XOR U475 ( .A(B[207]), .B(A[207]), .Z(n425) );
  AND U476 ( .A(n426), .B(n427), .Z(n424) );
  NANDN U477 ( .A(B[206]), .B(n428), .Z(n427) );
  NANDN U478 ( .A(A[206]), .B(n429), .Z(n428) );
  NANDN U479 ( .A(n429), .B(A[206]), .Z(n426) );
  XOR U480 ( .A(n429), .B(n430), .Z(DIFF[206]) );
  XOR U481 ( .A(B[206]), .B(A[206]), .Z(n430) );
  AND U482 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U483 ( .A(B[205]), .B(n433), .Z(n432) );
  NANDN U484 ( .A(A[205]), .B(n434), .Z(n433) );
  NANDN U485 ( .A(n434), .B(A[205]), .Z(n431) );
  XOR U486 ( .A(n434), .B(n435), .Z(DIFF[205]) );
  XOR U487 ( .A(B[205]), .B(A[205]), .Z(n435) );
  AND U488 ( .A(n436), .B(n437), .Z(n434) );
  NANDN U489 ( .A(B[204]), .B(n438), .Z(n437) );
  NANDN U490 ( .A(A[204]), .B(n439), .Z(n438) );
  NANDN U491 ( .A(n439), .B(A[204]), .Z(n436) );
  XOR U492 ( .A(n439), .B(n440), .Z(DIFF[204]) );
  XOR U493 ( .A(B[204]), .B(A[204]), .Z(n440) );
  AND U494 ( .A(n441), .B(n442), .Z(n439) );
  NANDN U495 ( .A(B[203]), .B(n443), .Z(n442) );
  NANDN U496 ( .A(A[203]), .B(n444), .Z(n443) );
  NANDN U497 ( .A(n444), .B(A[203]), .Z(n441) );
  XOR U498 ( .A(n444), .B(n445), .Z(DIFF[203]) );
  XOR U499 ( .A(B[203]), .B(A[203]), .Z(n445) );
  AND U500 ( .A(n446), .B(n447), .Z(n444) );
  NANDN U501 ( .A(B[202]), .B(n448), .Z(n447) );
  NANDN U502 ( .A(A[202]), .B(n449), .Z(n448) );
  NANDN U503 ( .A(n449), .B(A[202]), .Z(n446) );
  XOR U504 ( .A(n449), .B(n450), .Z(DIFF[202]) );
  XOR U505 ( .A(B[202]), .B(A[202]), .Z(n450) );
  AND U506 ( .A(n451), .B(n452), .Z(n449) );
  NANDN U507 ( .A(B[201]), .B(n453), .Z(n452) );
  NANDN U508 ( .A(A[201]), .B(n454), .Z(n453) );
  NANDN U509 ( .A(n454), .B(A[201]), .Z(n451) );
  XOR U510 ( .A(n454), .B(n455), .Z(DIFF[201]) );
  XOR U511 ( .A(B[201]), .B(A[201]), .Z(n455) );
  AND U512 ( .A(n456), .B(n457), .Z(n454) );
  NANDN U513 ( .A(B[200]), .B(n458), .Z(n457) );
  NANDN U514 ( .A(A[200]), .B(n459), .Z(n458) );
  NANDN U515 ( .A(n459), .B(A[200]), .Z(n456) );
  XOR U516 ( .A(n459), .B(n460), .Z(DIFF[200]) );
  XOR U517 ( .A(B[200]), .B(A[200]), .Z(n460) );
  AND U518 ( .A(n461), .B(n462), .Z(n459) );
  NANDN U519 ( .A(B[199]), .B(n463), .Z(n462) );
  NANDN U520 ( .A(A[199]), .B(n464), .Z(n463) );
  NANDN U521 ( .A(n464), .B(A[199]), .Z(n461) );
  XOR U522 ( .A(n2), .B(n465), .Z(DIFF[1]) );
  XOR U523 ( .A(B[1]), .B(A[1]), .Z(n465) );
  XOR U524 ( .A(n466), .B(n467), .Z(DIFF[19]) );
  XOR U525 ( .A(B[19]), .B(A[19]), .Z(n467) );
  XOR U526 ( .A(n464), .B(n468), .Z(DIFF[199]) );
  XOR U527 ( .A(B[199]), .B(A[199]), .Z(n468) );
  AND U528 ( .A(n469), .B(n470), .Z(n464) );
  NANDN U529 ( .A(B[198]), .B(n471), .Z(n470) );
  NANDN U530 ( .A(A[198]), .B(n472), .Z(n471) );
  NANDN U531 ( .A(n472), .B(A[198]), .Z(n469) );
  XOR U532 ( .A(n472), .B(n473), .Z(DIFF[198]) );
  XOR U533 ( .A(B[198]), .B(A[198]), .Z(n473) );
  AND U534 ( .A(n474), .B(n475), .Z(n472) );
  NANDN U535 ( .A(B[197]), .B(n476), .Z(n475) );
  NANDN U536 ( .A(A[197]), .B(n477), .Z(n476) );
  NANDN U537 ( .A(n477), .B(A[197]), .Z(n474) );
  XOR U538 ( .A(n477), .B(n478), .Z(DIFF[197]) );
  XOR U539 ( .A(B[197]), .B(A[197]), .Z(n478) );
  AND U540 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U541 ( .A(B[196]), .B(n481), .Z(n480) );
  NANDN U542 ( .A(A[196]), .B(n482), .Z(n481) );
  NANDN U543 ( .A(n482), .B(A[196]), .Z(n479) );
  XOR U544 ( .A(n482), .B(n483), .Z(DIFF[196]) );
  XOR U545 ( .A(B[196]), .B(A[196]), .Z(n483) );
  AND U546 ( .A(n484), .B(n485), .Z(n482) );
  NANDN U547 ( .A(B[195]), .B(n486), .Z(n485) );
  NANDN U548 ( .A(A[195]), .B(n487), .Z(n486) );
  NANDN U549 ( .A(n487), .B(A[195]), .Z(n484) );
  XOR U550 ( .A(n487), .B(n488), .Z(DIFF[195]) );
  XOR U551 ( .A(B[195]), .B(A[195]), .Z(n488) );
  AND U552 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U553 ( .A(B[194]), .B(n491), .Z(n490) );
  NANDN U554 ( .A(A[194]), .B(n492), .Z(n491) );
  NANDN U555 ( .A(n492), .B(A[194]), .Z(n489) );
  XOR U556 ( .A(n492), .B(n493), .Z(DIFF[194]) );
  XOR U557 ( .A(B[194]), .B(A[194]), .Z(n493) );
  AND U558 ( .A(n494), .B(n495), .Z(n492) );
  NANDN U559 ( .A(B[193]), .B(n496), .Z(n495) );
  NANDN U560 ( .A(A[193]), .B(n497), .Z(n496) );
  NANDN U561 ( .A(n497), .B(A[193]), .Z(n494) );
  XOR U562 ( .A(n497), .B(n498), .Z(DIFF[193]) );
  XOR U563 ( .A(B[193]), .B(A[193]), .Z(n498) );
  AND U564 ( .A(n499), .B(n500), .Z(n497) );
  NANDN U565 ( .A(B[192]), .B(n501), .Z(n500) );
  NANDN U566 ( .A(A[192]), .B(n502), .Z(n501) );
  NANDN U567 ( .A(n502), .B(A[192]), .Z(n499) );
  XOR U568 ( .A(n502), .B(n503), .Z(DIFF[192]) );
  XOR U569 ( .A(B[192]), .B(A[192]), .Z(n503) );
  AND U570 ( .A(n504), .B(n505), .Z(n502) );
  NANDN U571 ( .A(B[191]), .B(n506), .Z(n505) );
  NANDN U572 ( .A(A[191]), .B(n507), .Z(n506) );
  NANDN U573 ( .A(n507), .B(A[191]), .Z(n504) );
  XOR U574 ( .A(n507), .B(n508), .Z(DIFF[191]) );
  XOR U575 ( .A(B[191]), .B(A[191]), .Z(n508) );
  AND U576 ( .A(n509), .B(n510), .Z(n507) );
  NANDN U577 ( .A(B[190]), .B(n511), .Z(n510) );
  NANDN U578 ( .A(A[190]), .B(n512), .Z(n511) );
  NANDN U579 ( .A(n512), .B(A[190]), .Z(n509) );
  XOR U580 ( .A(n512), .B(n513), .Z(DIFF[190]) );
  XOR U581 ( .A(B[190]), .B(A[190]), .Z(n513) );
  AND U582 ( .A(n514), .B(n515), .Z(n512) );
  NANDN U583 ( .A(B[189]), .B(n516), .Z(n515) );
  NANDN U584 ( .A(A[189]), .B(n517), .Z(n516) );
  NANDN U585 ( .A(n517), .B(A[189]), .Z(n514) );
  XOR U586 ( .A(n518), .B(n519), .Z(DIFF[18]) );
  XOR U587 ( .A(B[18]), .B(A[18]), .Z(n519) );
  XOR U588 ( .A(n517), .B(n520), .Z(DIFF[189]) );
  XOR U589 ( .A(B[189]), .B(A[189]), .Z(n520) );
  AND U590 ( .A(n521), .B(n522), .Z(n517) );
  NANDN U591 ( .A(B[188]), .B(n523), .Z(n522) );
  NANDN U592 ( .A(A[188]), .B(n524), .Z(n523) );
  NANDN U593 ( .A(n524), .B(A[188]), .Z(n521) );
  XOR U594 ( .A(n524), .B(n525), .Z(DIFF[188]) );
  XOR U595 ( .A(B[188]), .B(A[188]), .Z(n525) );
  AND U596 ( .A(n526), .B(n527), .Z(n524) );
  NANDN U597 ( .A(B[187]), .B(n528), .Z(n527) );
  NANDN U598 ( .A(A[187]), .B(n529), .Z(n528) );
  NANDN U599 ( .A(n529), .B(A[187]), .Z(n526) );
  XOR U600 ( .A(n529), .B(n530), .Z(DIFF[187]) );
  XOR U601 ( .A(B[187]), .B(A[187]), .Z(n530) );
  AND U602 ( .A(n531), .B(n532), .Z(n529) );
  NANDN U603 ( .A(B[186]), .B(n533), .Z(n532) );
  NANDN U604 ( .A(A[186]), .B(n534), .Z(n533) );
  NANDN U605 ( .A(n534), .B(A[186]), .Z(n531) );
  XOR U606 ( .A(n534), .B(n535), .Z(DIFF[186]) );
  XOR U607 ( .A(B[186]), .B(A[186]), .Z(n535) );
  AND U608 ( .A(n536), .B(n537), .Z(n534) );
  NANDN U609 ( .A(B[185]), .B(n538), .Z(n537) );
  NANDN U610 ( .A(A[185]), .B(n539), .Z(n538) );
  NANDN U611 ( .A(n539), .B(A[185]), .Z(n536) );
  XOR U612 ( .A(n539), .B(n540), .Z(DIFF[185]) );
  XOR U613 ( .A(B[185]), .B(A[185]), .Z(n540) );
  AND U614 ( .A(n541), .B(n542), .Z(n539) );
  NANDN U615 ( .A(B[184]), .B(n543), .Z(n542) );
  NANDN U616 ( .A(A[184]), .B(n544), .Z(n543) );
  NANDN U617 ( .A(n544), .B(A[184]), .Z(n541) );
  XOR U618 ( .A(n544), .B(n545), .Z(DIFF[184]) );
  XOR U619 ( .A(B[184]), .B(A[184]), .Z(n545) );
  AND U620 ( .A(n546), .B(n547), .Z(n544) );
  NANDN U621 ( .A(B[183]), .B(n548), .Z(n547) );
  NANDN U622 ( .A(A[183]), .B(n549), .Z(n548) );
  NANDN U623 ( .A(n549), .B(A[183]), .Z(n546) );
  XOR U624 ( .A(n549), .B(n550), .Z(DIFF[183]) );
  XOR U625 ( .A(B[183]), .B(A[183]), .Z(n550) );
  AND U626 ( .A(n551), .B(n552), .Z(n549) );
  NANDN U627 ( .A(B[182]), .B(n553), .Z(n552) );
  NANDN U628 ( .A(A[182]), .B(n554), .Z(n553) );
  NANDN U629 ( .A(n554), .B(A[182]), .Z(n551) );
  XOR U630 ( .A(n554), .B(n555), .Z(DIFF[182]) );
  XOR U631 ( .A(B[182]), .B(A[182]), .Z(n555) );
  AND U632 ( .A(n556), .B(n557), .Z(n554) );
  NANDN U633 ( .A(B[181]), .B(n558), .Z(n557) );
  NANDN U634 ( .A(A[181]), .B(n559), .Z(n558) );
  NANDN U635 ( .A(n559), .B(A[181]), .Z(n556) );
  XOR U636 ( .A(n559), .B(n560), .Z(DIFF[181]) );
  XOR U637 ( .A(B[181]), .B(A[181]), .Z(n560) );
  AND U638 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U639 ( .A(B[180]), .B(n563), .Z(n562) );
  NANDN U640 ( .A(A[180]), .B(n564), .Z(n563) );
  NANDN U641 ( .A(n564), .B(A[180]), .Z(n561) );
  XOR U642 ( .A(n564), .B(n565), .Z(DIFF[180]) );
  XOR U643 ( .A(B[180]), .B(A[180]), .Z(n565) );
  AND U644 ( .A(n566), .B(n567), .Z(n564) );
  NANDN U645 ( .A(B[179]), .B(n568), .Z(n567) );
  NANDN U646 ( .A(A[179]), .B(n569), .Z(n568) );
  NANDN U647 ( .A(n569), .B(A[179]), .Z(n566) );
  XOR U648 ( .A(n570), .B(n571), .Z(DIFF[17]) );
  XOR U649 ( .A(B[17]), .B(A[17]), .Z(n571) );
  XOR U650 ( .A(n569), .B(n572), .Z(DIFF[179]) );
  XOR U651 ( .A(B[179]), .B(A[179]), .Z(n572) );
  AND U652 ( .A(n573), .B(n574), .Z(n569) );
  NANDN U653 ( .A(B[178]), .B(n575), .Z(n574) );
  NANDN U654 ( .A(A[178]), .B(n576), .Z(n575) );
  NANDN U655 ( .A(n576), .B(A[178]), .Z(n573) );
  XOR U656 ( .A(n576), .B(n577), .Z(DIFF[178]) );
  XOR U657 ( .A(B[178]), .B(A[178]), .Z(n577) );
  AND U658 ( .A(n578), .B(n579), .Z(n576) );
  NANDN U659 ( .A(B[177]), .B(n580), .Z(n579) );
  NANDN U660 ( .A(A[177]), .B(n581), .Z(n580) );
  NANDN U661 ( .A(n581), .B(A[177]), .Z(n578) );
  XOR U662 ( .A(n581), .B(n582), .Z(DIFF[177]) );
  XOR U663 ( .A(B[177]), .B(A[177]), .Z(n582) );
  AND U664 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U665 ( .A(B[176]), .B(n585), .Z(n584) );
  NANDN U666 ( .A(A[176]), .B(n586), .Z(n585) );
  NANDN U667 ( .A(n586), .B(A[176]), .Z(n583) );
  XOR U668 ( .A(n586), .B(n587), .Z(DIFF[176]) );
  XOR U669 ( .A(B[176]), .B(A[176]), .Z(n587) );
  AND U670 ( .A(n588), .B(n589), .Z(n586) );
  NANDN U671 ( .A(B[175]), .B(n590), .Z(n589) );
  NANDN U672 ( .A(A[175]), .B(n591), .Z(n590) );
  NANDN U673 ( .A(n591), .B(A[175]), .Z(n588) );
  XOR U674 ( .A(n591), .B(n592), .Z(DIFF[175]) );
  XOR U675 ( .A(B[175]), .B(A[175]), .Z(n592) );
  AND U676 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U677 ( .A(B[174]), .B(n595), .Z(n594) );
  NANDN U678 ( .A(A[174]), .B(n596), .Z(n595) );
  NANDN U679 ( .A(n596), .B(A[174]), .Z(n593) );
  XOR U680 ( .A(n596), .B(n597), .Z(DIFF[174]) );
  XOR U681 ( .A(B[174]), .B(A[174]), .Z(n597) );
  AND U682 ( .A(n598), .B(n599), .Z(n596) );
  NANDN U683 ( .A(B[173]), .B(n600), .Z(n599) );
  NANDN U684 ( .A(A[173]), .B(n601), .Z(n600) );
  NANDN U685 ( .A(n601), .B(A[173]), .Z(n598) );
  XOR U686 ( .A(n601), .B(n602), .Z(DIFF[173]) );
  XOR U687 ( .A(B[173]), .B(A[173]), .Z(n602) );
  AND U688 ( .A(n603), .B(n604), .Z(n601) );
  NANDN U689 ( .A(B[172]), .B(n605), .Z(n604) );
  NANDN U690 ( .A(A[172]), .B(n606), .Z(n605) );
  NANDN U691 ( .A(n606), .B(A[172]), .Z(n603) );
  XOR U692 ( .A(n606), .B(n607), .Z(DIFF[172]) );
  XOR U693 ( .A(B[172]), .B(A[172]), .Z(n607) );
  AND U694 ( .A(n608), .B(n609), .Z(n606) );
  NANDN U695 ( .A(B[171]), .B(n610), .Z(n609) );
  NANDN U696 ( .A(A[171]), .B(n611), .Z(n610) );
  NANDN U697 ( .A(n611), .B(A[171]), .Z(n608) );
  XOR U698 ( .A(n611), .B(n612), .Z(DIFF[171]) );
  XOR U699 ( .A(B[171]), .B(A[171]), .Z(n612) );
  AND U700 ( .A(n613), .B(n614), .Z(n611) );
  NANDN U701 ( .A(B[170]), .B(n615), .Z(n614) );
  NANDN U702 ( .A(A[170]), .B(n616), .Z(n615) );
  NANDN U703 ( .A(n616), .B(A[170]), .Z(n613) );
  XOR U704 ( .A(n616), .B(n617), .Z(DIFF[170]) );
  XOR U705 ( .A(B[170]), .B(A[170]), .Z(n617) );
  AND U706 ( .A(n618), .B(n619), .Z(n616) );
  NANDN U707 ( .A(B[169]), .B(n620), .Z(n619) );
  NANDN U708 ( .A(A[169]), .B(n621), .Z(n620) );
  NANDN U709 ( .A(n621), .B(A[169]), .Z(n618) );
  XOR U710 ( .A(n622), .B(n623), .Z(DIFF[16]) );
  XOR U711 ( .A(B[16]), .B(A[16]), .Z(n623) );
  XOR U712 ( .A(n621), .B(n624), .Z(DIFF[169]) );
  XOR U713 ( .A(B[169]), .B(A[169]), .Z(n624) );
  AND U714 ( .A(n625), .B(n626), .Z(n621) );
  NANDN U715 ( .A(B[168]), .B(n627), .Z(n626) );
  NANDN U716 ( .A(A[168]), .B(n628), .Z(n627) );
  NANDN U717 ( .A(n628), .B(A[168]), .Z(n625) );
  XOR U718 ( .A(n628), .B(n629), .Z(DIFF[168]) );
  XOR U719 ( .A(B[168]), .B(A[168]), .Z(n629) );
  AND U720 ( .A(n630), .B(n631), .Z(n628) );
  NANDN U721 ( .A(B[167]), .B(n632), .Z(n631) );
  NANDN U722 ( .A(A[167]), .B(n633), .Z(n632) );
  NANDN U723 ( .A(n633), .B(A[167]), .Z(n630) );
  XOR U724 ( .A(n633), .B(n634), .Z(DIFF[167]) );
  XOR U725 ( .A(B[167]), .B(A[167]), .Z(n634) );
  AND U726 ( .A(n635), .B(n636), .Z(n633) );
  NANDN U727 ( .A(B[166]), .B(n637), .Z(n636) );
  NANDN U728 ( .A(A[166]), .B(n638), .Z(n637) );
  NANDN U729 ( .A(n638), .B(A[166]), .Z(n635) );
  XOR U730 ( .A(n638), .B(n639), .Z(DIFF[166]) );
  XOR U731 ( .A(B[166]), .B(A[166]), .Z(n639) );
  AND U732 ( .A(n640), .B(n641), .Z(n638) );
  NANDN U733 ( .A(B[165]), .B(n642), .Z(n641) );
  NANDN U734 ( .A(A[165]), .B(n643), .Z(n642) );
  NANDN U735 ( .A(n643), .B(A[165]), .Z(n640) );
  XOR U736 ( .A(n643), .B(n644), .Z(DIFF[165]) );
  XOR U737 ( .A(B[165]), .B(A[165]), .Z(n644) );
  AND U738 ( .A(n645), .B(n646), .Z(n643) );
  NANDN U739 ( .A(B[164]), .B(n647), .Z(n646) );
  NANDN U740 ( .A(A[164]), .B(n648), .Z(n647) );
  NANDN U741 ( .A(n648), .B(A[164]), .Z(n645) );
  XOR U742 ( .A(n648), .B(n649), .Z(DIFF[164]) );
  XOR U743 ( .A(B[164]), .B(A[164]), .Z(n649) );
  AND U744 ( .A(n650), .B(n651), .Z(n648) );
  NANDN U745 ( .A(B[163]), .B(n652), .Z(n651) );
  NANDN U746 ( .A(A[163]), .B(n653), .Z(n652) );
  NANDN U747 ( .A(n653), .B(A[163]), .Z(n650) );
  XOR U748 ( .A(n653), .B(n654), .Z(DIFF[163]) );
  XOR U749 ( .A(B[163]), .B(A[163]), .Z(n654) );
  AND U750 ( .A(n655), .B(n656), .Z(n653) );
  NANDN U751 ( .A(B[162]), .B(n657), .Z(n656) );
  NANDN U752 ( .A(A[162]), .B(n658), .Z(n657) );
  NANDN U753 ( .A(n658), .B(A[162]), .Z(n655) );
  XOR U754 ( .A(n658), .B(n659), .Z(DIFF[162]) );
  XOR U755 ( .A(B[162]), .B(A[162]), .Z(n659) );
  AND U756 ( .A(n660), .B(n661), .Z(n658) );
  NANDN U757 ( .A(B[161]), .B(n662), .Z(n661) );
  NANDN U758 ( .A(A[161]), .B(n663), .Z(n662) );
  NANDN U759 ( .A(n663), .B(A[161]), .Z(n660) );
  XOR U760 ( .A(n663), .B(n664), .Z(DIFF[161]) );
  XOR U761 ( .A(B[161]), .B(A[161]), .Z(n664) );
  AND U762 ( .A(n665), .B(n666), .Z(n663) );
  NANDN U763 ( .A(B[160]), .B(n667), .Z(n666) );
  NANDN U764 ( .A(A[160]), .B(n668), .Z(n667) );
  NANDN U765 ( .A(n668), .B(A[160]), .Z(n665) );
  XOR U766 ( .A(n668), .B(n669), .Z(DIFF[160]) );
  XOR U767 ( .A(B[160]), .B(A[160]), .Z(n669) );
  AND U768 ( .A(n670), .B(n671), .Z(n668) );
  NANDN U769 ( .A(B[159]), .B(n672), .Z(n671) );
  NANDN U770 ( .A(A[159]), .B(n673), .Z(n672) );
  NANDN U771 ( .A(n673), .B(A[159]), .Z(n670) );
  XOR U772 ( .A(n674), .B(n675), .Z(DIFF[15]) );
  XOR U773 ( .A(B[15]), .B(A[15]), .Z(n675) );
  XOR U774 ( .A(n673), .B(n676), .Z(DIFF[159]) );
  XOR U775 ( .A(B[159]), .B(A[159]), .Z(n676) );
  AND U776 ( .A(n677), .B(n678), .Z(n673) );
  NANDN U777 ( .A(B[158]), .B(n679), .Z(n678) );
  NANDN U778 ( .A(A[158]), .B(n680), .Z(n679) );
  NANDN U779 ( .A(n680), .B(A[158]), .Z(n677) );
  XOR U780 ( .A(n680), .B(n681), .Z(DIFF[158]) );
  XOR U781 ( .A(B[158]), .B(A[158]), .Z(n681) );
  AND U782 ( .A(n682), .B(n683), .Z(n680) );
  NANDN U783 ( .A(B[157]), .B(n684), .Z(n683) );
  NANDN U784 ( .A(A[157]), .B(n685), .Z(n684) );
  NANDN U785 ( .A(n685), .B(A[157]), .Z(n682) );
  XOR U786 ( .A(n685), .B(n686), .Z(DIFF[157]) );
  XOR U787 ( .A(B[157]), .B(A[157]), .Z(n686) );
  AND U788 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U789 ( .A(B[156]), .B(n689), .Z(n688) );
  NANDN U790 ( .A(A[156]), .B(n690), .Z(n689) );
  NANDN U791 ( .A(n690), .B(A[156]), .Z(n687) );
  XOR U792 ( .A(n690), .B(n691), .Z(DIFF[156]) );
  XOR U793 ( .A(B[156]), .B(A[156]), .Z(n691) );
  AND U794 ( .A(n692), .B(n693), .Z(n690) );
  NANDN U795 ( .A(B[155]), .B(n694), .Z(n693) );
  NANDN U796 ( .A(A[155]), .B(n695), .Z(n694) );
  NANDN U797 ( .A(n695), .B(A[155]), .Z(n692) );
  XOR U798 ( .A(n695), .B(n696), .Z(DIFF[155]) );
  XOR U799 ( .A(B[155]), .B(A[155]), .Z(n696) );
  AND U800 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U801 ( .A(B[154]), .B(n699), .Z(n698) );
  NANDN U802 ( .A(A[154]), .B(n700), .Z(n699) );
  NANDN U803 ( .A(n700), .B(A[154]), .Z(n697) );
  XOR U804 ( .A(n700), .B(n701), .Z(DIFF[154]) );
  XOR U805 ( .A(B[154]), .B(A[154]), .Z(n701) );
  AND U806 ( .A(n702), .B(n703), .Z(n700) );
  NANDN U807 ( .A(B[153]), .B(n704), .Z(n703) );
  NANDN U808 ( .A(A[153]), .B(n705), .Z(n704) );
  NANDN U809 ( .A(n705), .B(A[153]), .Z(n702) );
  XOR U810 ( .A(n705), .B(n706), .Z(DIFF[153]) );
  XOR U811 ( .A(B[153]), .B(A[153]), .Z(n706) );
  AND U812 ( .A(n707), .B(n708), .Z(n705) );
  NANDN U813 ( .A(B[152]), .B(n709), .Z(n708) );
  NANDN U814 ( .A(A[152]), .B(n710), .Z(n709) );
  NANDN U815 ( .A(n710), .B(A[152]), .Z(n707) );
  XOR U816 ( .A(n710), .B(n711), .Z(DIFF[152]) );
  XOR U817 ( .A(B[152]), .B(A[152]), .Z(n711) );
  AND U818 ( .A(n712), .B(n713), .Z(n710) );
  NANDN U819 ( .A(B[151]), .B(n714), .Z(n713) );
  NANDN U820 ( .A(A[151]), .B(n715), .Z(n714) );
  NANDN U821 ( .A(n715), .B(A[151]), .Z(n712) );
  XOR U822 ( .A(n715), .B(n716), .Z(DIFF[151]) );
  XOR U823 ( .A(B[151]), .B(A[151]), .Z(n716) );
  AND U824 ( .A(n717), .B(n718), .Z(n715) );
  NANDN U825 ( .A(B[150]), .B(n719), .Z(n718) );
  NANDN U826 ( .A(A[150]), .B(n720), .Z(n719) );
  NANDN U827 ( .A(n720), .B(A[150]), .Z(n717) );
  XOR U828 ( .A(n720), .B(n721), .Z(DIFF[150]) );
  XOR U829 ( .A(B[150]), .B(A[150]), .Z(n721) );
  AND U830 ( .A(n722), .B(n723), .Z(n720) );
  NANDN U831 ( .A(B[149]), .B(n724), .Z(n723) );
  NANDN U832 ( .A(A[149]), .B(n725), .Z(n724) );
  NANDN U833 ( .A(n725), .B(A[149]), .Z(n722) );
  XOR U834 ( .A(n726), .B(n727), .Z(DIFF[14]) );
  XOR U835 ( .A(B[14]), .B(A[14]), .Z(n727) );
  XOR U836 ( .A(n725), .B(n728), .Z(DIFF[149]) );
  XOR U837 ( .A(B[149]), .B(A[149]), .Z(n728) );
  AND U838 ( .A(n729), .B(n730), .Z(n725) );
  NANDN U839 ( .A(B[148]), .B(n731), .Z(n730) );
  NANDN U840 ( .A(A[148]), .B(n732), .Z(n731) );
  NANDN U841 ( .A(n732), .B(A[148]), .Z(n729) );
  XOR U842 ( .A(n732), .B(n733), .Z(DIFF[148]) );
  XOR U843 ( .A(B[148]), .B(A[148]), .Z(n733) );
  AND U844 ( .A(n734), .B(n735), .Z(n732) );
  NANDN U845 ( .A(B[147]), .B(n736), .Z(n735) );
  NANDN U846 ( .A(A[147]), .B(n737), .Z(n736) );
  NANDN U847 ( .A(n737), .B(A[147]), .Z(n734) );
  XOR U848 ( .A(n737), .B(n738), .Z(DIFF[147]) );
  XOR U849 ( .A(B[147]), .B(A[147]), .Z(n738) );
  AND U850 ( .A(n739), .B(n740), .Z(n737) );
  NANDN U851 ( .A(B[146]), .B(n741), .Z(n740) );
  NANDN U852 ( .A(A[146]), .B(n742), .Z(n741) );
  NANDN U853 ( .A(n742), .B(A[146]), .Z(n739) );
  XOR U854 ( .A(n742), .B(n743), .Z(DIFF[146]) );
  XOR U855 ( .A(B[146]), .B(A[146]), .Z(n743) );
  AND U856 ( .A(n744), .B(n745), .Z(n742) );
  NANDN U857 ( .A(B[145]), .B(n746), .Z(n745) );
  NANDN U858 ( .A(A[145]), .B(n747), .Z(n746) );
  NANDN U859 ( .A(n747), .B(A[145]), .Z(n744) );
  XOR U860 ( .A(n747), .B(n748), .Z(DIFF[145]) );
  XOR U861 ( .A(B[145]), .B(A[145]), .Z(n748) );
  AND U862 ( .A(n749), .B(n750), .Z(n747) );
  NANDN U863 ( .A(B[144]), .B(n751), .Z(n750) );
  NANDN U864 ( .A(A[144]), .B(n752), .Z(n751) );
  NANDN U865 ( .A(n752), .B(A[144]), .Z(n749) );
  XOR U866 ( .A(n752), .B(n753), .Z(DIFF[144]) );
  XOR U867 ( .A(B[144]), .B(A[144]), .Z(n753) );
  AND U868 ( .A(n754), .B(n755), .Z(n752) );
  NANDN U869 ( .A(B[143]), .B(n756), .Z(n755) );
  NANDN U870 ( .A(A[143]), .B(n757), .Z(n756) );
  NANDN U871 ( .A(n757), .B(A[143]), .Z(n754) );
  XOR U872 ( .A(n757), .B(n758), .Z(DIFF[143]) );
  XOR U873 ( .A(B[143]), .B(A[143]), .Z(n758) );
  AND U874 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U875 ( .A(B[142]), .B(n761), .Z(n760) );
  NANDN U876 ( .A(A[142]), .B(n762), .Z(n761) );
  NANDN U877 ( .A(n762), .B(A[142]), .Z(n759) );
  XOR U878 ( .A(n762), .B(n763), .Z(DIFF[142]) );
  XOR U879 ( .A(B[142]), .B(A[142]), .Z(n763) );
  AND U880 ( .A(n764), .B(n765), .Z(n762) );
  NANDN U881 ( .A(B[141]), .B(n766), .Z(n765) );
  NANDN U882 ( .A(A[141]), .B(n767), .Z(n766) );
  NANDN U883 ( .A(n767), .B(A[141]), .Z(n764) );
  XOR U884 ( .A(n767), .B(n768), .Z(DIFF[141]) );
  XOR U885 ( .A(B[141]), .B(A[141]), .Z(n768) );
  AND U886 ( .A(n769), .B(n770), .Z(n767) );
  NANDN U887 ( .A(B[140]), .B(n771), .Z(n770) );
  NANDN U888 ( .A(A[140]), .B(n772), .Z(n771) );
  NANDN U889 ( .A(n772), .B(A[140]), .Z(n769) );
  XOR U890 ( .A(n772), .B(n773), .Z(DIFF[140]) );
  XOR U891 ( .A(B[140]), .B(A[140]), .Z(n773) );
  AND U892 ( .A(n774), .B(n775), .Z(n772) );
  NANDN U893 ( .A(B[139]), .B(n776), .Z(n775) );
  NANDN U894 ( .A(A[139]), .B(n777), .Z(n776) );
  NANDN U895 ( .A(n777), .B(A[139]), .Z(n774) );
  XOR U896 ( .A(n778), .B(n779), .Z(DIFF[13]) );
  XOR U897 ( .A(B[13]), .B(A[13]), .Z(n779) );
  XOR U898 ( .A(n777), .B(n780), .Z(DIFF[139]) );
  XOR U899 ( .A(B[139]), .B(A[139]), .Z(n780) );
  AND U900 ( .A(n781), .B(n782), .Z(n777) );
  NANDN U901 ( .A(B[138]), .B(n783), .Z(n782) );
  NANDN U902 ( .A(A[138]), .B(n784), .Z(n783) );
  NANDN U903 ( .A(n784), .B(A[138]), .Z(n781) );
  XOR U904 ( .A(n784), .B(n785), .Z(DIFF[138]) );
  XOR U905 ( .A(B[138]), .B(A[138]), .Z(n785) );
  AND U906 ( .A(n786), .B(n787), .Z(n784) );
  NANDN U907 ( .A(B[137]), .B(n788), .Z(n787) );
  NANDN U908 ( .A(A[137]), .B(n789), .Z(n788) );
  NANDN U909 ( .A(n789), .B(A[137]), .Z(n786) );
  XOR U910 ( .A(n789), .B(n790), .Z(DIFF[137]) );
  XOR U911 ( .A(B[137]), .B(A[137]), .Z(n790) );
  AND U912 ( .A(n791), .B(n792), .Z(n789) );
  NANDN U913 ( .A(B[136]), .B(n793), .Z(n792) );
  NANDN U914 ( .A(A[136]), .B(n794), .Z(n793) );
  NANDN U915 ( .A(n794), .B(A[136]), .Z(n791) );
  XOR U916 ( .A(n794), .B(n795), .Z(DIFF[136]) );
  XOR U917 ( .A(B[136]), .B(A[136]), .Z(n795) );
  AND U918 ( .A(n796), .B(n797), .Z(n794) );
  NANDN U919 ( .A(B[135]), .B(n798), .Z(n797) );
  NANDN U920 ( .A(A[135]), .B(n799), .Z(n798) );
  NANDN U921 ( .A(n799), .B(A[135]), .Z(n796) );
  XOR U922 ( .A(n799), .B(n800), .Z(DIFF[135]) );
  XOR U923 ( .A(B[135]), .B(A[135]), .Z(n800) );
  AND U924 ( .A(n801), .B(n802), .Z(n799) );
  NANDN U925 ( .A(B[134]), .B(n803), .Z(n802) );
  NANDN U926 ( .A(A[134]), .B(n804), .Z(n803) );
  NANDN U927 ( .A(n804), .B(A[134]), .Z(n801) );
  XOR U928 ( .A(n804), .B(n805), .Z(DIFF[134]) );
  XOR U929 ( .A(B[134]), .B(A[134]), .Z(n805) );
  AND U930 ( .A(n806), .B(n807), .Z(n804) );
  NANDN U931 ( .A(B[133]), .B(n808), .Z(n807) );
  NANDN U932 ( .A(A[133]), .B(n809), .Z(n808) );
  NANDN U933 ( .A(n809), .B(A[133]), .Z(n806) );
  XOR U934 ( .A(n809), .B(n810), .Z(DIFF[133]) );
  XOR U935 ( .A(B[133]), .B(A[133]), .Z(n810) );
  AND U936 ( .A(n811), .B(n812), .Z(n809) );
  NANDN U937 ( .A(B[132]), .B(n813), .Z(n812) );
  NANDN U938 ( .A(A[132]), .B(n814), .Z(n813) );
  NANDN U939 ( .A(n814), .B(A[132]), .Z(n811) );
  XOR U940 ( .A(n814), .B(n815), .Z(DIFF[132]) );
  XOR U941 ( .A(B[132]), .B(A[132]), .Z(n815) );
  AND U942 ( .A(n816), .B(n817), .Z(n814) );
  NANDN U943 ( .A(B[131]), .B(n818), .Z(n817) );
  NANDN U944 ( .A(A[131]), .B(n819), .Z(n818) );
  NANDN U945 ( .A(n819), .B(A[131]), .Z(n816) );
  XOR U946 ( .A(n819), .B(n820), .Z(DIFF[131]) );
  XOR U947 ( .A(B[131]), .B(A[131]), .Z(n820) );
  AND U948 ( .A(n821), .B(n822), .Z(n819) );
  NANDN U949 ( .A(B[130]), .B(n823), .Z(n822) );
  NANDN U950 ( .A(A[130]), .B(n824), .Z(n823) );
  NANDN U951 ( .A(n824), .B(A[130]), .Z(n821) );
  XOR U952 ( .A(n824), .B(n825), .Z(DIFF[130]) );
  XOR U953 ( .A(B[130]), .B(A[130]), .Z(n825) );
  AND U954 ( .A(n826), .B(n827), .Z(n824) );
  NANDN U955 ( .A(B[129]), .B(n828), .Z(n827) );
  NANDN U956 ( .A(A[129]), .B(n829), .Z(n828) );
  NANDN U957 ( .A(n829), .B(A[129]), .Z(n826) );
  XOR U958 ( .A(n830), .B(n831), .Z(DIFF[12]) );
  XOR U959 ( .A(B[12]), .B(A[12]), .Z(n831) );
  XOR U960 ( .A(n829), .B(n832), .Z(DIFF[129]) );
  XOR U961 ( .A(B[129]), .B(A[129]), .Z(n832) );
  AND U962 ( .A(n833), .B(n834), .Z(n829) );
  NANDN U963 ( .A(B[128]), .B(n835), .Z(n834) );
  NANDN U964 ( .A(A[128]), .B(n836), .Z(n835) );
  NANDN U965 ( .A(n836), .B(A[128]), .Z(n833) );
  XOR U966 ( .A(n836), .B(n837), .Z(DIFF[128]) );
  XOR U967 ( .A(B[128]), .B(A[128]), .Z(n837) );
  AND U968 ( .A(n838), .B(n839), .Z(n836) );
  NANDN U969 ( .A(B[127]), .B(n840), .Z(n839) );
  NANDN U970 ( .A(A[127]), .B(n841), .Z(n840) );
  NANDN U971 ( .A(n841), .B(A[127]), .Z(n838) );
  XOR U972 ( .A(n841), .B(n842), .Z(DIFF[127]) );
  XOR U973 ( .A(B[127]), .B(A[127]), .Z(n842) );
  AND U974 ( .A(n843), .B(n844), .Z(n841) );
  NANDN U975 ( .A(B[126]), .B(n845), .Z(n844) );
  NANDN U976 ( .A(A[126]), .B(n846), .Z(n845) );
  NANDN U977 ( .A(n846), .B(A[126]), .Z(n843) );
  XOR U978 ( .A(n846), .B(n847), .Z(DIFF[126]) );
  XOR U979 ( .A(B[126]), .B(A[126]), .Z(n847) );
  AND U980 ( .A(n848), .B(n849), .Z(n846) );
  NANDN U981 ( .A(B[125]), .B(n850), .Z(n849) );
  NANDN U982 ( .A(A[125]), .B(n851), .Z(n850) );
  NANDN U983 ( .A(n851), .B(A[125]), .Z(n848) );
  XOR U984 ( .A(n851), .B(n852), .Z(DIFF[125]) );
  XOR U985 ( .A(B[125]), .B(A[125]), .Z(n852) );
  AND U986 ( .A(n853), .B(n854), .Z(n851) );
  NANDN U987 ( .A(B[124]), .B(n855), .Z(n854) );
  NANDN U988 ( .A(A[124]), .B(n856), .Z(n855) );
  NANDN U989 ( .A(n856), .B(A[124]), .Z(n853) );
  XOR U990 ( .A(n856), .B(n857), .Z(DIFF[124]) );
  XOR U991 ( .A(B[124]), .B(A[124]), .Z(n857) );
  AND U992 ( .A(n858), .B(n859), .Z(n856) );
  NANDN U993 ( .A(B[123]), .B(n860), .Z(n859) );
  NANDN U994 ( .A(A[123]), .B(n861), .Z(n860) );
  NANDN U995 ( .A(n861), .B(A[123]), .Z(n858) );
  XOR U996 ( .A(n861), .B(n862), .Z(DIFF[123]) );
  XOR U997 ( .A(B[123]), .B(A[123]), .Z(n862) );
  AND U998 ( .A(n863), .B(n864), .Z(n861) );
  NANDN U999 ( .A(B[122]), .B(n865), .Z(n864) );
  NANDN U1000 ( .A(A[122]), .B(n866), .Z(n865) );
  NANDN U1001 ( .A(n866), .B(A[122]), .Z(n863) );
  XOR U1002 ( .A(n866), .B(n867), .Z(DIFF[122]) );
  XOR U1003 ( .A(B[122]), .B(A[122]), .Z(n867) );
  AND U1004 ( .A(n868), .B(n869), .Z(n866) );
  NANDN U1005 ( .A(B[121]), .B(n870), .Z(n869) );
  NANDN U1006 ( .A(A[121]), .B(n871), .Z(n870) );
  NANDN U1007 ( .A(n871), .B(A[121]), .Z(n868) );
  XOR U1008 ( .A(n871), .B(n872), .Z(DIFF[121]) );
  XOR U1009 ( .A(B[121]), .B(A[121]), .Z(n872) );
  AND U1010 ( .A(n873), .B(n874), .Z(n871) );
  NANDN U1011 ( .A(B[120]), .B(n875), .Z(n874) );
  NANDN U1012 ( .A(A[120]), .B(n876), .Z(n875) );
  NANDN U1013 ( .A(n876), .B(A[120]), .Z(n873) );
  XOR U1014 ( .A(n876), .B(n877), .Z(DIFF[120]) );
  XOR U1015 ( .A(B[120]), .B(A[120]), .Z(n877) );
  AND U1016 ( .A(n878), .B(n879), .Z(n876) );
  NANDN U1017 ( .A(B[119]), .B(n880), .Z(n879) );
  NANDN U1018 ( .A(A[119]), .B(n881), .Z(n880) );
  NANDN U1019 ( .A(n881), .B(A[119]), .Z(n878) );
  XOR U1020 ( .A(n882), .B(n883), .Z(DIFF[11]) );
  XOR U1021 ( .A(B[11]), .B(A[11]), .Z(n883) );
  XOR U1022 ( .A(n881), .B(n884), .Z(DIFF[119]) );
  XOR U1023 ( .A(B[119]), .B(A[119]), .Z(n884) );
  AND U1024 ( .A(n885), .B(n886), .Z(n881) );
  NANDN U1025 ( .A(B[118]), .B(n887), .Z(n886) );
  NANDN U1026 ( .A(A[118]), .B(n888), .Z(n887) );
  NANDN U1027 ( .A(n888), .B(A[118]), .Z(n885) );
  XOR U1028 ( .A(n888), .B(n889), .Z(DIFF[118]) );
  XOR U1029 ( .A(B[118]), .B(A[118]), .Z(n889) );
  AND U1030 ( .A(n890), .B(n891), .Z(n888) );
  NANDN U1031 ( .A(B[117]), .B(n892), .Z(n891) );
  NANDN U1032 ( .A(A[117]), .B(n893), .Z(n892) );
  NANDN U1033 ( .A(n893), .B(A[117]), .Z(n890) );
  XOR U1034 ( .A(n893), .B(n894), .Z(DIFF[117]) );
  XOR U1035 ( .A(B[117]), .B(A[117]), .Z(n894) );
  AND U1036 ( .A(n895), .B(n896), .Z(n893) );
  NANDN U1037 ( .A(B[116]), .B(n897), .Z(n896) );
  NANDN U1038 ( .A(A[116]), .B(n898), .Z(n897) );
  NANDN U1039 ( .A(n898), .B(A[116]), .Z(n895) );
  XOR U1040 ( .A(n898), .B(n899), .Z(DIFF[116]) );
  XOR U1041 ( .A(B[116]), .B(A[116]), .Z(n899) );
  AND U1042 ( .A(n900), .B(n901), .Z(n898) );
  NANDN U1043 ( .A(B[115]), .B(n902), .Z(n901) );
  NANDN U1044 ( .A(A[115]), .B(n903), .Z(n902) );
  NANDN U1045 ( .A(n903), .B(A[115]), .Z(n900) );
  XOR U1046 ( .A(n903), .B(n904), .Z(DIFF[115]) );
  XOR U1047 ( .A(B[115]), .B(A[115]), .Z(n904) );
  AND U1048 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U1049 ( .A(B[114]), .B(n907), .Z(n906) );
  NANDN U1050 ( .A(A[114]), .B(n908), .Z(n907) );
  NANDN U1051 ( .A(n908), .B(A[114]), .Z(n905) );
  XOR U1052 ( .A(n908), .B(n909), .Z(DIFF[114]) );
  XOR U1053 ( .A(B[114]), .B(A[114]), .Z(n909) );
  AND U1054 ( .A(n910), .B(n911), .Z(n908) );
  NANDN U1055 ( .A(B[113]), .B(n912), .Z(n911) );
  NANDN U1056 ( .A(A[113]), .B(n913), .Z(n912) );
  NANDN U1057 ( .A(n913), .B(A[113]), .Z(n910) );
  XOR U1058 ( .A(n913), .B(n914), .Z(DIFF[113]) );
  XOR U1059 ( .A(B[113]), .B(A[113]), .Z(n914) );
  AND U1060 ( .A(n915), .B(n916), .Z(n913) );
  NANDN U1061 ( .A(B[112]), .B(n917), .Z(n916) );
  NANDN U1062 ( .A(A[112]), .B(n918), .Z(n917) );
  NANDN U1063 ( .A(n918), .B(A[112]), .Z(n915) );
  XOR U1064 ( .A(n918), .B(n919), .Z(DIFF[112]) );
  XOR U1065 ( .A(B[112]), .B(A[112]), .Z(n919) );
  AND U1066 ( .A(n920), .B(n921), .Z(n918) );
  NANDN U1067 ( .A(B[111]), .B(n922), .Z(n921) );
  NANDN U1068 ( .A(A[111]), .B(n923), .Z(n922) );
  NANDN U1069 ( .A(n923), .B(A[111]), .Z(n920) );
  XOR U1070 ( .A(n923), .B(n924), .Z(DIFF[111]) );
  XOR U1071 ( .A(B[111]), .B(A[111]), .Z(n924) );
  AND U1072 ( .A(n925), .B(n926), .Z(n923) );
  NANDN U1073 ( .A(B[110]), .B(n927), .Z(n926) );
  NANDN U1074 ( .A(A[110]), .B(n928), .Z(n927) );
  NANDN U1075 ( .A(n928), .B(A[110]), .Z(n925) );
  XOR U1076 ( .A(n928), .B(n929), .Z(DIFF[110]) );
  XOR U1077 ( .A(B[110]), .B(A[110]), .Z(n929) );
  AND U1078 ( .A(n930), .B(n931), .Z(n928) );
  NANDN U1079 ( .A(B[109]), .B(n932), .Z(n931) );
  NANDN U1080 ( .A(A[109]), .B(n933), .Z(n932) );
  NANDN U1081 ( .A(n933), .B(A[109]), .Z(n930) );
  XOR U1082 ( .A(n934), .B(n935), .Z(DIFF[10]) );
  XOR U1083 ( .A(B[10]), .B(A[10]), .Z(n935) );
  XOR U1084 ( .A(n933), .B(n936), .Z(DIFF[109]) );
  XOR U1085 ( .A(B[109]), .B(A[109]), .Z(n936) );
  AND U1086 ( .A(n937), .B(n938), .Z(n933) );
  NANDN U1087 ( .A(B[108]), .B(n939), .Z(n938) );
  NANDN U1088 ( .A(A[108]), .B(n940), .Z(n939) );
  NANDN U1089 ( .A(n940), .B(A[108]), .Z(n937) );
  XOR U1090 ( .A(n940), .B(n941), .Z(DIFF[108]) );
  XOR U1091 ( .A(B[108]), .B(A[108]), .Z(n941) );
  AND U1092 ( .A(n942), .B(n943), .Z(n940) );
  NANDN U1093 ( .A(B[107]), .B(n944), .Z(n943) );
  NANDN U1094 ( .A(A[107]), .B(n945), .Z(n944) );
  NANDN U1095 ( .A(n945), .B(A[107]), .Z(n942) );
  XOR U1096 ( .A(n945), .B(n946), .Z(DIFF[107]) );
  XOR U1097 ( .A(B[107]), .B(A[107]), .Z(n946) );
  AND U1098 ( .A(n947), .B(n948), .Z(n945) );
  NANDN U1099 ( .A(B[106]), .B(n949), .Z(n948) );
  NANDN U1100 ( .A(A[106]), .B(n950), .Z(n949) );
  NANDN U1101 ( .A(n950), .B(A[106]), .Z(n947) );
  XOR U1102 ( .A(n950), .B(n951), .Z(DIFF[106]) );
  XOR U1103 ( .A(B[106]), .B(A[106]), .Z(n951) );
  AND U1104 ( .A(n952), .B(n953), .Z(n950) );
  NANDN U1105 ( .A(B[105]), .B(n954), .Z(n953) );
  NANDN U1106 ( .A(A[105]), .B(n955), .Z(n954) );
  NANDN U1107 ( .A(n955), .B(A[105]), .Z(n952) );
  XOR U1108 ( .A(n955), .B(n956), .Z(DIFF[105]) );
  XOR U1109 ( .A(B[105]), .B(A[105]), .Z(n956) );
  AND U1110 ( .A(n957), .B(n958), .Z(n955) );
  NANDN U1111 ( .A(B[104]), .B(n959), .Z(n958) );
  NANDN U1112 ( .A(A[104]), .B(n960), .Z(n959) );
  NANDN U1113 ( .A(n960), .B(A[104]), .Z(n957) );
  XOR U1114 ( .A(n960), .B(n961), .Z(DIFF[104]) );
  XOR U1115 ( .A(B[104]), .B(A[104]), .Z(n961) );
  AND U1116 ( .A(n962), .B(n963), .Z(n960) );
  NANDN U1117 ( .A(B[103]), .B(n964), .Z(n963) );
  NANDN U1118 ( .A(A[103]), .B(n965), .Z(n964) );
  NANDN U1119 ( .A(n965), .B(A[103]), .Z(n962) );
  XOR U1120 ( .A(n965), .B(n966), .Z(DIFF[103]) );
  XOR U1121 ( .A(B[103]), .B(A[103]), .Z(n966) );
  AND U1122 ( .A(n967), .B(n968), .Z(n965) );
  NANDN U1123 ( .A(B[102]), .B(n969), .Z(n968) );
  NANDN U1124 ( .A(A[102]), .B(n970), .Z(n969) );
  NANDN U1125 ( .A(n970), .B(A[102]), .Z(n967) );
  XOR U1126 ( .A(n970), .B(n971), .Z(DIFF[102]) );
  XOR U1127 ( .A(B[102]), .B(A[102]), .Z(n971) );
  AND U1128 ( .A(n972), .B(n973), .Z(n970) );
  NANDN U1129 ( .A(B[101]), .B(n974), .Z(n973) );
  NANDN U1130 ( .A(A[101]), .B(n975), .Z(n974) );
  NANDN U1131 ( .A(n975), .B(A[101]), .Z(n972) );
  XOR U1132 ( .A(n975), .B(n976), .Z(DIFF[101]) );
  XOR U1133 ( .A(B[101]), .B(A[101]), .Z(n976) );
  AND U1134 ( .A(n977), .B(n978), .Z(n975) );
  NANDN U1135 ( .A(B[100]), .B(n979), .Z(n978) );
  NANDN U1136 ( .A(A[100]), .B(n980), .Z(n979) );
  NANDN U1137 ( .A(n980), .B(A[100]), .Z(n977) );
  XOR U1138 ( .A(n980), .B(n981), .Z(DIFF[100]) );
  XOR U1139 ( .A(B[100]), .B(A[100]), .Z(n981) );
  AND U1140 ( .A(n982), .B(n983), .Z(n980) );
  NANDN U1141 ( .A(B[99]), .B(n984), .Z(n983) );
  OR U1142 ( .A(n5), .B(A[99]), .Z(n984) );
  NAND U1143 ( .A(A[99]), .B(n5), .Z(n982) );
  NAND U1144 ( .A(n985), .B(n986), .Z(n5) );
  NANDN U1145 ( .A(B[98]), .B(n987), .Z(n986) );
  NANDN U1146 ( .A(A[98]), .B(n7), .Z(n987) );
  NANDN U1147 ( .A(n7), .B(A[98]), .Z(n985) );
  AND U1148 ( .A(n988), .B(n989), .Z(n7) );
  NANDN U1149 ( .A(B[97]), .B(n990), .Z(n989) );
  NANDN U1150 ( .A(A[97]), .B(n9), .Z(n990) );
  NANDN U1151 ( .A(n9), .B(A[97]), .Z(n988) );
  AND U1152 ( .A(n991), .B(n992), .Z(n9) );
  NANDN U1153 ( .A(B[96]), .B(n993), .Z(n992) );
  NANDN U1154 ( .A(A[96]), .B(n11), .Z(n993) );
  NANDN U1155 ( .A(n11), .B(A[96]), .Z(n991) );
  AND U1156 ( .A(n994), .B(n995), .Z(n11) );
  NANDN U1157 ( .A(B[95]), .B(n996), .Z(n995) );
  NANDN U1158 ( .A(A[95]), .B(n13), .Z(n996) );
  NANDN U1159 ( .A(n13), .B(A[95]), .Z(n994) );
  AND U1160 ( .A(n997), .B(n998), .Z(n13) );
  NANDN U1161 ( .A(B[94]), .B(n999), .Z(n998) );
  NANDN U1162 ( .A(A[94]), .B(n15), .Z(n999) );
  NANDN U1163 ( .A(n15), .B(A[94]), .Z(n997) );
  AND U1164 ( .A(n1000), .B(n1001), .Z(n15) );
  NANDN U1165 ( .A(B[93]), .B(n1002), .Z(n1001) );
  NANDN U1166 ( .A(A[93]), .B(n17), .Z(n1002) );
  NANDN U1167 ( .A(n17), .B(A[93]), .Z(n1000) );
  AND U1168 ( .A(n1003), .B(n1004), .Z(n17) );
  NANDN U1169 ( .A(B[92]), .B(n1005), .Z(n1004) );
  NANDN U1170 ( .A(A[92]), .B(n19), .Z(n1005) );
  NANDN U1171 ( .A(n19), .B(A[92]), .Z(n1003) );
  AND U1172 ( .A(n1006), .B(n1007), .Z(n19) );
  NANDN U1173 ( .A(B[91]), .B(n1008), .Z(n1007) );
  NANDN U1174 ( .A(A[91]), .B(n21), .Z(n1008) );
  NANDN U1175 ( .A(n21), .B(A[91]), .Z(n1006) );
  AND U1176 ( .A(n1009), .B(n1010), .Z(n21) );
  NANDN U1177 ( .A(B[90]), .B(n1011), .Z(n1010) );
  NANDN U1178 ( .A(A[90]), .B(n23), .Z(n1011) );
  NANDN U1179 ( .A(n23), .B(A[90]), .Z(n1009) );
  AND U1180 ( .A(n1012), .B(n1013), .Z(n23) );
  NANDN U1181 ( .A(B[89]), .B(n1014), .Z(n1013) );
  NANDN U1182 ( .A(A[89]), .B(n27), .Z(n1014) );
  NANDN U1183 ( .A(n27), .B(A[89]), .Z(n1012) );
  AND U1184 ( .A(n1015), .B(n1016), .Z(n27) );
  NANDN U1185 ( .A(B[88]), .B(n1017), .Z(n1016) );
  NANDN U1186 ( .A(A[88]), .B(n29), .Z(n1017) );
  NANDN U1187 ( .A(n29), .B(A[88]), .Z(n1015) );
  AND U1188 ( .A(n1018), .B(n1019), .Z(n29) );
  NANDN U1189 ( .A(B[87]), .B(n1020), .Z(n1019) );
  NANDN U1190 ( .A(A[87]), .B(n31), .Z(n1020) );
  NANDN U1191 ( .A(n31), .B(A[87]), .Z(n1018) );
  AND U1192 ( .A(n1021), .B(n1022), .Z(n31) );
  NANDN U1193 ( .A(B[86]), .B(n1023), .Z(n1022) );
  NANDN U1194 ( .A(A[86]), .B(n33), .Z(n1023) );
  NANDN U1195 ( .A(n33), .B(A[86]), .Z(n1021) );
  AND U1196 ( .A(n1024), .B(n1025), .Z(n33) );
  NANDN U1197 ( .A(B[85]), .B(n1026), .Z(n1025) );
  NANDN U1198 ( .A(A[85]), .B(n35), .Z(n1026) );
  NANDN U1199 ( .A(n35), .B(A[85]), .Z(n1024) );
  AND U1200 ( .A(n1027), .B(n1028), .Z(n35) );
  NANDN U1201 ( .A(B[84]), .B(n1029), .Z(n1028) );
  NANDN U1202 ( .A(A[84]), .B(n37), .Z(n1029) );
  NANDN U1203 ( .A(n37), .B(A[84]), .Z(n1027) );
  AND U1204 ( .A(n1030), .B(n1031), .Z(n37) );
  NANDN U1205 ( .A(B[83]), .B(n1032), .Z(n1031) );
  NANDN U1206 ( .A(A[83]), .B(n39), .Z(n1032) );
  NANDN U1207 ( .A(n39), .B(A[83]), .Z(n1030) );
  AND U1208 ( .A(n1033), .B(n1034), .Z(n39) );
  NANDN U1209 ( .A(B[82]), .B(n1035), .Z(n1034) );
  NANDN U1210 ( .A(A[82]), .B(n41), .Z(n1035) );
  NANDN U1211 ( .A(n41), .B(A[82]), .Z(n1033) );
  AND U1212 ( .A(n1036), .B(n1037), .Z(n41) );
  NANDN U1213 ( .A(B[81]), .B(n1038), .Z(n1037) );
  NANDN U1214 ( .A(A[81]), .B(n43), .Z(n1038) );
  NANDN U1215 ( .A(n43), .B(A[81]), .Z(n1036) );
  AND U1216 ( .A(n1039), .B(n1040), .Z(n43) );
  NANDN U1217 ( .A(B[80]), .B(n1041), .Z(n1040) );
  NANDN U1218 ( .A(A[80]), .B(n45), .Z(n1041) );
  NANDN U1219 ( .A(n45), .B(A[80]), .Z(n1039) );
  AND U1220 ( .A(n1042), .B(n1043), .Z(n45) );
  NANDN U1221 ( .A(B[79]), .B(n1044), .Z(n1043) );
  NANDN U1222 ( .A(A[79]), .B(n49), .Z(n1044) );
  NANDN U1223 ( .A(n49), .B(A[79]), .Z(n1042) );
  AND U1224 ( .A(n1045), .B(n1046), .Z(n49) );
  NANDN U1225 ( .A(B[78]), .B(n1047), .Z(n1046) );
  NANDN U1226 ( .A(A[78]), .B(n51), .Z(n1047) );
  NANDN U1227 ( .A(n51), .B(A[78]), .Z(n1045) );
  AND U1228 ( .A(n1048), .B(n1049), .Z(n51) );
  NANDN U1229 ( .A(B[77]), .B(n1050), .Z(n1049) );
  NANDN U1230 ( .A(A[77]), .B(n53), .Z(n1050) );
  NANDN U1231 ( .A(n53), .B(A[77]), .Z(n1048) );
  AND U1232 ( .A(n1051), .B(n1052), .Z(n53) );
  NANDN U1233 ( .A(B[76]), .B(n1053), .Z(n1052) );
  NANDN U1234 ( .A(A[76]), .B(n55), .Z(n1053) );
  NANDN U1235 ( .A(n55), .B(A[76]), .Z(n1051) );
  AND U1236 ( .A(n1054), .B(n1055), .Z(n55) );
  NANDN U1237 ( .A(B[75]), .B(n1056), .Z(n1055) );
  NANDN U1238 ( .A(A[75]), .B(n57), .Z(n1056) );
  NANDN U1239 ( .A(n57), .B(A[75]), .Z(n1054) );
  AND U1240 ( .A(n1057), .B(n1058), .Z(n57) );
  NANDN U1241 ( .A(B[74]), .B(n1059), .Z(n1058) );
  NANDN U1242 ( .A(A[74]), .B(n59), .Z(n1059) );
  NANDN U1243 ( .A(n59), .B(A[74]), .Z(n1057) );
  AND U1244 ( .A(n1060), .B(n1061), .Z(n59) );
  NANDN U1245 ( .A(B[73]), .B(n1062), .Z(n1061) );
  NANDN U1246 ( .A(A[73]), .B(n61), .Z(n1062) );
  NANDN U1247 ( .A(n61), .B(A[73]), .Z(n1060) );
  AND U1248 ( .A(n1063), .B(n1064), .Z(n61) );
  NANDN U1249 ( .A(B[72]), .B(n1065), .Z(n1064) );
  NANDN U1250 ( .A(A[72]), .B(n63), .Z(n1065) );
  NANDN U1251 ( .A(n63), .B(A[72]), .Z(n1063) );
  AND U1252 ( .A(n1066), .B(n1067), .Z(n63) );
  NANDN U1253 ( .A(B[71]), .B(n1068), .Z(n1067) );
  NANDN U1254 ( .A(A[71]), .B(n65), .Z(n1068) );
  NANDN U1255 ( .A(n65), .B(A[71]), .Z(n1066) );
  AND U1256 ( .A(n1069), .B(n1070), .Z(n65) );
  NANDN U1257 ( .A(B[70]), .B(n1071), .Z(n1070) );
  NANDN U1258 ( .A(A[70]), .B(n67), .Z(n1071) );
  NANDN U1259 ( .A(n67), .B(A[70]), .Z(n1069) );
  AND U1260 ( .A(n1072), .B(n1073), .Z(n67) );
  NANDN U1261 ( .A(B[69]), .B(n1074), .Z(n1073) );
  NANDN U1262 ( .A(A[69]), .B(n71), .Z(n1074) );
  NANDN U1263 ( .A(n71), .B(A[69]), .Z(n1072) );
  AND U1264 ( .A(n1075), .B(n1076), .Z(n71) );
  NANDN U1265 ( .A(B[68]), .B(n1077), .Z(n1076) );
  NANDN U1266 ( .A(A[68]), .B(n73), .Z(n1077) );
  NANDN U1267 ( .A(n73), .B(A[68]), .Z(n1075) );
  AND U1268 ( .A(n1078), .B(n1079), .Z(n73) );
  NANDN U1269 ( .A(B[67]), .B(n1080), .Z(n1079) );
  NANDN U1270 ( .A(A[67]), .B(n75), .Z(n1080) );
  NANDN U1271 ( .A(n75), .B(A[67]), .Z(n1078) );
  AND U1272 ( .A(n1081), .B(n1082), .Z(n75) );
  NANDN U1273 ( .A(B[66]), .B(n1083), .Z(n1082) );
  NANDN U1274 ( .A(A[66]), .B(n77), .Z(n1083) );
  NANDN U1275 ( .A(n77), .B(A[66]), .Z(n1081) );
  AND U1276 ( .A(n1084), .B(n1085), .Z(n77) );
  NANDN U1277 ( .A(B[65]), .B(n1086), .Z(n1085) );
  NANDN U1278 ( .A(A[65]), .B(n79), .Z(n1086) );
  NANDN U1279 ( .A(n79), .B(A[65]), .Z(n1084) );
  AND U1280 ( .A(n1087), .B(n1088), .Z(n79) );
  NANDN U1281 ( .A(B[64]), .B(n1089), .Z(n1088) );
  NANDN U1282 ( .A(A[64]), .B(n81), .Z(n1089) );
  NANDN U1283 ( .A(n81), .B(A[64]), .Z(n1087) );
  AND U1284 ( .A(n1090), .B(n1091), .Z(n81) );
  NANDN U1285 ( .A(B[63]), .B(n1092), .Z(n1091) );
  NANDN U1286 ( .A(A[63]), .B(n83), .Z(n1092) );
  NANDN U1287 ( .A(n83), .B(A[63]), .Z(n1090) );
  AND U1288 ( .A(n1093), .B(n1094), .Z(n83) );
  NANDN U1289 ( .A(B[62]), .B(n1095), .Z(n1094) );
  NANDN U1290 ( .A(A[62]), .B(n85), .Z(n1095) );
  NANDN U1291 ( .A(n85), .B(A[62]), .Z(n1093) );
  AND U1292 ( .A(n1096), .B(n1097), .Z(n85) );
  NANDN U1293 ( .A(B[61]), .B(n1098), .Z(n1097) );
  NANDN U1294 ( .A(A[61]), .B(n87), .Z(n1098) );
  NANDN U1295 ( .A(n87), .B(A[61]), .Z(n1096) );
  AND U1296 ( .A(n1099), .B(n1100), .Z(n87) );
  NANDN U1297 ( .A(B[60]), .B(n1101), .Z(n1100) );
  NANDN U1298 ( .A(A[60]), .B(n89), .Z(n1101) );
  NANDN U1299 ( .A(n89), .B(A[60]), .Z(n1099) );
  AND U1300 ( .A(n1102), .B(n1103), .Z(n89) );
  NANDN U1301 ( .A(B[59]), .B(n1104), .Z(n1103) );
  NANDN U1302 ( .A(A[59]), .B(n93), .Z(n1104) );
  NANDN U1303 ( .A(n93), .B(A[59]), .Z(n1102) );
  AND U1304 ( .A(n1105), .B(n1106), .Z(n93) );
  NANDN U1305 ( .A(B[58]), .B(n1107), .Z(n1106) );
  NANDN U1306 ( .A(A[58]), .B(n95), .Z(n1107) );
  NANDN U1307 ( .A(n95), .B(A[58]), .Z(n1105) );
  AND U1308 ( .A(n1108), .B(n1109), .Z(n95) );
  NANDN U1309 ( .A(B[57]), .B(n1110), .Z(n1109) );
  NANDN U1310 ( .A(A[57]), .B(n97), .Z(n1110) );
  NANDN U1311 ( .A(n97), .B(A[57]), .Z(n1108) );
  AND U1312 ( .A(n1111), .B(n1112), .Z(n97) );
  NANDN U1313 ( .A(B[56]), .B(n1113), .Z(n1112) );
  NANDN U1314 ( .A(A[56]), .B(n99), .Z(n1113) );
  NANDN U1315 ( .A(n99), .B(A[56]), .Z(n1111) );
  AND U1316 ( .A(n1114), .B(n1115), .Z(n99) );
  NANDN U1317 ( .A(B[55]), .B(n1116), .Z(n1115) );
  NANDN U1318 ( .A(A[55]), .B(n101), .Z(n1116) );
  NANDN U1319 ( .A(n101), .B(A[55]), .Z(n1114) );
  AND U1320 ( .A(n1117), .B(n1118), .Z(n101) );
  NANDN U1321 ( .A(B[54]), .B(n1119), .Z(n1118) );
  NANDN U1322 ( .A(A[54]), .B(n103), .Z(n1119) );
  NANDN U1323 ( .A(n103), .B(A[54]), .Z(n1117) );
  AND U1324 ( .A(n1120), .B(n1121), .Z(n103) );
  NANDN U1325 ( .A(B[53]), .B(n1122), .Z(n1121) );
  NANDN U1326 ( .A(A[53]), .B(n105), .Z(n1122) );
  NANDN U1327 ( .A(n105), .B(A[53]), .Z(n1120) );
  AND U1328 ( .A(n1123), .B(n1124), .Z(n105) );
  NANDN U1329 ( .A(B[52]), .B(n1125), .Z(n1124) );
  NANDN U1330 ( .A(A[52]), .B(n107), .Z(n1125) );
  NANDN U1331 ( .A(n107), .B(A[52]), .Z(n1123) );
  AND U1332 ( .A(n1126), .B(n1127), .Z(n107) );
  NANDN U1333 ( .A(B[51]), .B(n1128), .Z(n1127) );
  NANDN U1334 ( .A(A[51]), .B(n109), .Z(n1128) );
  NANDN U1335 ( .A(n109), .B(A[51]), .Z(n1126) );
  AND U1336 ( .A(n1129), .B(n1130), .Z(n109) );
  NANDN U1337 ( .A(B[50]), .B(n1131), .Z(n1130) );
  NANDN U1338 ( .A(A[50]), .B(n111), .Z(n1131) );
  NANDN U1339 ( .A(n111), .B(A[50]), .Z(n1129) );
  AND U1340 ( .A(n1132), .B(n1133), .Z(n111) );
  NANDN U1341 ( .A(B[49]), .B(n1134), .Z(n1133) );
  NANDN U1342 ( .A(A[49]), .B(n115), .Z(n1134) );
  NANDN U1343 ( .A(n115), .B(A[49]), .Z(n1132) );
  AND U1344 ( .A(n1135), .B(n1136), .Z(n115) );
  NANDN U1345 ( .A(B[48]), .B(n1137), .Z(n1136) );
  NANDN U1346 ( .A(A[48]), .B(n117), .Z(n1137) );
  NANDN U1347 ( .A(n117), .B(A[48]), .Z(n1135) );
  AND U1348 ( .A(n1138), .B(n1139), .Z(n117) );
  NANDN U1349 ( .A(B[47]), .B(n1140), .Z(n1139) );
  NANDN U1350 ( .A(A[47]), .B(n119), .Z(n1140) );
  NANDN U1351 ( .A(n119), .B(A[47]), .Z(n1138) );
  AND U1352 ( .A(n1141), .B(n1142), .Z(n119) );
  NANDN U1353 ( .A(B[46]), .B(n1143), .Z(n1142) );
  NANDN U1354 ( .A(A[46]), .B(n121), .Z(n1143) );
  NANDN U1355 ( .A(n121), .B(A[46]), .Z(n1141) );
  AND U1356 ( .A(n1144), .B(n1145), .Z(n121) );
  NANDN U1357 ( .A(B[45]), .B(n1146), .Z(n1145) );
  NANDN U1358 ( .A(A[45]), .B(n123), .Z(n1146) );
  NANDN U1359 ( .A(n123), .B(A[45]), .Z(n1144) );
  AND U1360 ( .A(n1147), .B(n1148), .Z(n123) );
  NANDN U1361 ( .A(B[44]), .B(n1149), .Z(n1148) );
  NANDN U1362 ( .A(A[44]), .B(n125), .Z(n1149) );
  NANDN U1363 ( .A(n125), .B(A[44]), .Z(n1147) );
  AND U1364 ( .A(n1150), .B(n1151), .Z(n125) );
  NANDN U1365 ( .A(B[43]), .B(n1152), .Z(n1151) );
  NANDN U1366 ( .A(A[43]), .B(n127), .Z(n1152) );
  NANDN U1367 ( .A(n127), .B(A[43]), .Z(n1150) );
  AND U1368 ( .A(n1153), .B(n1154), .Z(n127) );
  NANDN U1369 ( .A(B[42]), .B(n1155), .Z(n1154) );
  NANDN U1370 ( .A(A[42]), .B(n129), .Z(n1155) );
  NANDN U1371 ( .A(n129), .B(A[42]), .Z(n1153) );
  AND U1372 ( .A(n1156), .B(n1157), .Z(n129) );
  NANDN U1373 ( .A(B[41]), .B(n1158), .Z(n1157) );
  NANDN U1374 ( .A(A[41]), .B(n131), .Z(n1158) );
  NANDN U1375 ( .A(n131), .B(A[41]), .Z(n1156) );
  AND U1376 ( .A(n1159), .B(n1160), .Z(n131) );
  NANDN U1377 ( .A(B[40]), .B(n1161), .Z(n1160) );
  NANDN U1378 ( .A(A[40]), .B(n133), .Z(n1161) );
  NANDN U1379 ( .A(n133), .B(A[40]), .Z(n1159) );
  AND U1380 ( .A(n1162), .B(n1163), .Z(n133) );
  NANDN U1381 ( .A(B[39]), .B(n1164), .Z(n1163) );
  NANDN U1382 ( .A(A[39]), .B(n137), .Z(n1164) );
  NANDN U1383 ( .A(n137), .B(A[39]), .Z(n1162) );
  AND U1384 ( .A(n1165), .B(n1166), .Z(n137) );
  NANDN U1385 ( .A(B[38]), .B(n1167), .Z(n1166) );
  NANDN U1386 ( .A(A[38]), .B(n139), .Z(n1167) );
  NANDN U1387 ( .A(n139), .B(A[38]), .Z(n1165) );
  AND U1388 ( .A(n1168), .B(n1169), .Z(n139) );
  NANDN U1389 ( .A(B[37]), .B(n1170), .Z(n1169) );
  NANDN U1390 ( .A(A[37]), .B(n141), .Z(n1170) );
  NANDN U1391 ( .A(n141), .B(A[37]), .Z(n1168) );
  AND U1392 ( .A(n1171), .B(n1172), .Z(n141) );
  NANDN U1393 ( .A(B[36]), .B(n1173), .Z(n1172) );
  NANDN U1394 ( .A(A[36]), .B(n143), .Z(n1173) );
  NANDN U1395 ( .A(n143), .B(A[36]), .Z(n1171) );
  AND U1396 ( .A(n1174), .B(n1175), .Z(n143) );
  NANDN U1397 ( .A(B[35]), .B(n1176), .Z(n1175) );
  NANDN U1398 ( .A(A[35]), .B(n145), .Z(n1176) );
  NANDN U1399 ( .A(n145), .B(A[35]), .Z(n1174) );
  AND U1400 ( .A(n1177), .B(n1178), .Z(n145) );
  NANDN U1401 ( .A(B[34]), .B(n1179), .Z(n1178) );
  NANDN U1402 ( .A(A[34]), .B(n147), .Z(n1179) );
  NANDN U1403 ( .A(n147), .B(A[34]), .Z(n1177) );
  AND U1404 ( .A(n1180), .B(n1181), .Z(n147) );
  NANDN U1405 ( .A(B[33]), .B(n1182), .Z(n1181) );
  NANDN U1406 ( .A(A[33]), .B(n149), .Z(n1182) );
  NANDN U1407 ( .A(n149), .B(A[33]), .Z(n1180) );
  AND U1408 ( .A(n1183), .B(n1184), .Z(n149) );
  NANDN U1409 ( .A(B[32]), .B(n1185), .Z(n1184) );
  NANDN U1410 ( .A(A[32]), .B(n151), .Z(n1185) );
  NANDN U1411 ( .A(n151), .B(A[32]), .Z(n1183) );
  AND U1412 ( .A(n1186), .B(n1187), .Z(n151) );
  NANDN U1413 ( .A(B[31]), .B(n1188), .Z(n1187) );
  NANDN U1414 ( .A(A[31]), .B(n153), .Z(n1188) );
  NANDN U1415 ( .A(n153), .B(A[31]), .Z(n1186) );
  AND U1416 ( .A(n1189), .B(n1190), .Z(n153) );
  NANDN U1417 ( .A(B[30]), .B(n1191), .Z(n1190) );
  NANDN U1418 ( .A(A[30]), .B(n155), .Z(n1191) );
  NANDN U1419 ( .A(n155), .B(A[30]), .Z(n1189) );
  AND U1420 ( .A(n1192), .B(n1193), .Z(n155) );
  NANDN U1421 ( .A(B[29]), .B(n1194), .Z(n1193) );
  NANDN U1422 ( .A(A[29]), .B(n159), .Z(n1194) );
  NANDN U1423 ( .A(n159), .B(A[29]), .Z(n1192) );
  AND U1424 ( .A(n1195), .B(n1196), .Z(n159) );
  NANDN U1425 ( .A(B[28]), .B(n1197), .Z(n1196) );
  NANDN U1426 ( .A(A[28]), .B(n161), .Z(n1197) );
  NANDN U1427 ( .A(n161), .B(A[28]), .Z(n1195) );
  AND U1428 ( .A(n1198), .B(n1199), .Z(n161) );
  NANDN U1429 ( .A(B[27]), .B(n1200), .Z(n1199) );
  NANDN U1430 ( .A(A[27]), .B(n163), .Z(n1200) );
  NANDN U1431 ( .A(n163), .B(A[27]), .Z(n1198) );
  AND U1432 ( .A(n1201), .B(n1202), .Z(n163) );
  NANDN U1433 ( .A(B[26]), .B(n1203), .Z(n1202) );
  NANDN U1434 ( .A(A[26]), .B(n165), .Z(n1203) );
  NANDN U1435 ( .A(n165), .B(A[26]), .Z(n1201) );
  AND U1436 ( .A(n1204), .B(n1205), .Z(n165) );
  NANDN U1437 ( .A(B[25]), .B(n1206), .Z(n1205) );
  NANDN U1438 ( .A(A[25]), .B(n167), .Z(n1206) );
  NANDN U1439 ( .A(n167), .B(A[25]), .Z(n1204) );
  AND U1440 ( .A(n1207), .B(n1208), .Z(n167) );
  NANDN U1441 ( .A(B[24]), .B(n1209), .Z(n1208) );
  NANDN U1442 ( .A(A[24]), .B(n205), .Z(n1209) );
  NANDN U1443 ( .A(n205), .B(A[24]), .Z(n1207) );
  AND U1444 ( .A(n1210), .B(n1211), .Z(n205) );
  NANDN U1445 ( .A(B[23]), .B(n1212), .Z(n1211) );
  NANDN U1446 ( .A(A[23]), .B(n257), .Z(n1212) );
  NANDN U1447 ( .A(n257), .B(A[23]), .Z(n1210) );
  AND U1448 ( .A(n1213), .B(n1214), .Z(n257) );
  NANDN U1449 ( .A(B[22]), .B(n1215), .Z(n1214) );
  NANDN U1450 ( .A(A[22]), .B(n309), .Z(n1215) );
  NANDN U1451 ( .A(n309), .B(A[22]), .Z(n1213) );
  AND U1452 ( .A(n1216), .B(n1217), .Z(n309) );
  NANDN U1453 ( .A(B[21]), .B(n1218), .Z(n1217) );
  NANDN U1454 ( .A(A[21]), .B(n361), .Z(n1218) );
  NANDN U1455 ( .A(n361), .B(A[21]), .Z(n1216) );
  AND U1456 ( .A(n1219), .B(n1220), .Z(n361) );
  NANDN U1457 ( .A(B[20]), .B(n1221), .Z(n1220) );
  NANDN U1458 ( .A(A[20]), .B(n413), .Z(n1221) );
  NANDN U1459 ( .A(n413), .B(A[20]), .Z(n1219) );
  AND U1460 ( .A(n1222), .B(n1223), .Z(n413) );
  NANDN U1461 ( .A(B[19]), .B(n1224), .Z(n1223) );
  NANDN U1462 ( .A(A[19]), .B(n466), .Z(n1224) );
  NANDN U1463 ( .A(n466), .B(A[19]), .Z(n1222) );
  AND U1464 ( .A(n1225), .B(n1226), .Z(n466) );
  NANDN U1465 ( .A(B[18]), .B(n1227), .Z(n1226) );
  NANDN U1466 ( .A(A[18]), .B(n518), .Z(n1227) );
  NANDN U1467 ( .A(n518), .B(A[18]), .Z(n1225) );
  AND U1468 ( .A(n1228), .B(n1229), .Z(n518) );
  NANDN U1469 ( .A(B[17]), .B(n1230), .Z(n1229) );
  NANDN U1470 ( .A(A[17]), .B(n570), .Z(n1230) );
  NANDN U1471 ( .A(n570), .B(A[17]), .Z(n1228) );
  AND U1472 ( .A(n1231), .B(n1232), .Z(n570) );
  NANDN U1473 ( .A(B[16]), .B(n1233), .Z(n1232) );
  NANDN U1474 ( .A(A[16]), .B(n622), .Z(n1233) );
  NANDN U1475 ( .A(n622), .B(A[16]), .Z(n1231) );
  AND U1476 ( .A(n1234), .B(n1235), .Z(n622) );
  NANDN U1477 ( .A(B[15]), .B(n1236), .Z(n1235) );
  NANDN U1478 ( .A(A[15]), .B(n674), .Z(n1236) );
  NANDN U1479 ( .A(n674), .B(A[15]), .Z(n1234) );
  AND U1480 ( .A(n1237), .B(n1238), .Z(n674) );
  NANDN U1481 ( .A(B[14]), .B(n1239), .Z(n1238) );
  NANDN U1482 ( .A(A[14]), .B(n726), .Z(n1239) );
  NANDN U1483 ( .A(n726), .B(A[14]), .Z(n1237) );
  AND U1484 ( .A(n1240), .B(n1241), .Z(n726) );
  NANDN U1485 ( .A(B[13]), .B(n1242), .Z(n1241) );
  NANDN U1486 ( .A(A[13]), .B(n778), .Z(n1242) );
  NANDN U1487 ( .A(n778), .B(A[13]), .Z(n1240) );
  AND U1488 ( .A(n1243), .B(n1244), .Z(n778) );
  NANDN U1489 ( .A(B[12]), .B(n1245), .Z(n1244) );
  NANDN U1490 ( .A(A[12]), .B(n830), .Z(n1245) );
  NANDN U1491 ( .A(n830), .B(A[12]), .Z(n1243) );
  AND U1492 ( .A(n1246), .B(n1247), .Z(n830) );
  NANDN U1493 ( .A(B[11]), .B(n1248), .Z(n1247) );
  NANDN U1494 ( .A(A[11]), .B(n882), .Z(n1248) );
  NANDN U1495 ( .A(n882), .B(A[11]), .Z(n1246) );
  AND U1496 ( .A(n1249), .B(n1250), .Z(n882) );
  NANDN U1497 ( .A(B[10]), .B(n1251), .Z(n1250) );
  NANDN U1498 ( .A(A[10]), .B(n934), .Z(n1251) );
  NANDN U1499 ( .A(n934), .B(A[10]), .Z(n1249) );
  AND U1500 ( .A(n1252), .B(n1253), .Z(n934) );
  NANDN U1501 ( .A(B[9]), .B(n1254), .Z(n1253) );
  OR U1502 ( .A(n3), .B(A[9]), .Z(n1254) );
  NAND U1503 ( .A(A[9]), .B(n3), .Z(n1252) );
  NAND U1504 ( .A(n1255), .B(n1256), .Z(n3) );
  NANDN U1505 ( .A(B[8]), .B(n1257), .Z(n1256) );
  NANDN U1506 ( .A(A[8]), .B(n25), .Z(n1257) );
  NANDN U1507 ( .A(n25), .B(A[8]), .Z(n1255) );
  AND U1508 ( .A(n1258), .B(n1259), .Z(n25) );
  NANDN U1509 ( .A(B[7]), .B(n1260), .Z(n1259) );
  NANDN U1510 ( .A(A[7]), .B(n47), .Z(n1260) );
  NANDN U1511 ( .A(n47), .B(A[7]), .Z(n1258) );
  AND U1512 ( .A(n1261), .B(n1262), .Z(n47) );
  NANDN U1513 ( .A(B[6]), .B(n1263), .Z(n1262) );
  NANDN U1514 ( .A(A[6]), .B(n69), .Z(n1263) );
  NANDN U1515 ( .A(n69), .B(A[6]), .Z(n1261) );
  AND U1516 ( .A(n1264), .B(n1265), .Z(n69) );
  NANDN U1517 ( .A(B[5]), .B(n1266), .Z(n1265) );
  NANDN U1518 ( .A(A[5]), .B(n91), .Z(n1266) );
  NANDN U1519 ( .A(n91), .B(A[5]), .Z(n1264) );
  AND U1520 ( .A(n1267), .B(n1268), .Z(n91) );
  NANDN U1521 ( .A(B[4]), .B(n1269), .Z(n1268) );
  NANDN U1522 ( .A(A[4]), .B(n113), .Z(n1269) );
  NANDN U1523 ( .A(n113), .B(A[4]), .Z(n1267) );
  AND U1524 ( .A(n1270), .B(n1271), .Z(n113) );
  NANDN U1525 ( .A(B[3]), .B(n1272), .Z(n1271) );
  NANDN U1526 ( .A(A[3]), .B(n135), .Z(n1272) );
  NANDN U1527 ( .A(n135), .B(A[3]), .Z(n1270) );
  AND U1528 ( .A(n1273), .B(n1274), .Z(n135) );
  NANDN U1529 ( .A(B[2]), .B(n1275), .Z(n1274) );
  NANDN U1530 ( .A(A[2]), .B(n157), .Z(n1275) );
  NANDN U1531 ( .A(n157), .B(A[2]), .Z(n1273) );
  AND U1532 ( .A(n1276), .B(n1277), .Z(n157) );
  NANDN U1533 ( .A(B[1]), .B(n1278), .Z(n1277) );
  NAND U1534 ( .A(n2), .B(n1), .Z(n1278) );
  NAND U1535 ( .A(A[1]), .B(n1279), .Z(n1276) );
  NAND U1536 ( .A(n1279), .B(n1280), .Z(DIFF[0]) );
  NANDN U1537 ( .A(B[0]), .B(A[0]), .Z(n1280) );
  NANDN U1538 ( .A(A[0]), .B(B[0]), .Z(n1279) );
endmodule


module modmult_step_N256_3_DW01_cmp2_1 ( A, B, LEQ, TC, LT_LE, GE_GT );
  input [257:0] A;
  input [257:0] B;
  input LEQ, TC;
  output LT_LE, GE_GT;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022;

  NAND U1 ( .A(n1), .B(n2), .Z(LT_LE) );
  NOR U2 ( .A(B[257]), .B(B[256]), .Z(n2) );
  AND U3 ( .A(n3), .B(n4), .Z(n1) );
  NAND U4 ( .A(n5), .B(n6), .Z(n4) );
  NANDN U5 ( .A(B[255]), .B(A[255]), .Z(n6) );
  NAND U6 ( .A(n7), .B(n8), .Z(n5) );
  NANDN U7 ( .A(A[254]), .B(B[254]), .Z(n8) );
  NAND U8 ( .A(n9), .B(n10), .Z(n7) );
  NANDN U9 ( .A(B[254]), .B(A[254]), .Z(n10) );
  AND U10 ( .A(n11), .B(n12), .Z(n9) );
  NAND U11 ( .A(n13), .B(n14), .Z(n12) );
  NANDN U12 ( .A(A[253]), .B(B[253]), .Z(n14) );
  AND U13 ( .A(n15), .B(n16), .Z(n13) );
  NANDN U14 ( .A(A[252]), .B(B[252]), .Z(n16) );
  NAND U15 ( .A(n17), .B(n18), .Z(n15) );
  NANDN U16 ( .A(B[252]), .B(A[252]), .Z(n18) );
  AND U17 ( .A(n19), .B(n20), .Z(n17) );
  NAND U18 ( .A(n21), .B(n22), .Z(n20) );
  NANDN U19 ( .A(A[251]), .B(B[251]), .Z(n22) );
  AND U20 ( .A(n23), .B(n24), .Z(n21) );
  NANDN U21 ( .A(A[250]), .B(B[250]), .Z(n24) );
  NAND U22 ( .A(n25), .B(n26), .Z(n23) );
  NANDN U23 ( .A(B[250]), .B(A[250]), .Z(n26) );
  AND U24 ( .A(n27), .B(n28), .Z(n25) );
  NAND U25 ( .A(n29), .B(n30), .Z(n28) );
  NANDN U26 ( .A(A[249]), .B(B[249]), .Z(n30) );
  AND U27 ( .A(n31), .B(n32), .Z(n29) );
  NANDN U28 ( .A(A[248]), .B(B[248]), .Z(n32) );
  NAND U29 ( .A(n33), .B(n34), .Z(n31) );
  NANDN U30 ( .A(B[248]), .B(A[248]), .Z(n34) );
  AND U31 ( .A(n35), .B(n36), .Z(n33) );
  NAND U32 ( .A(n37), .B(n38), .Z(n36) );
  NANDN U33 ( .A(A[247]), .B(B[247]), .Z(n38) );
  AND U34 ( .A(n39), .B(n40), .Z(n37) );
  NANDN U35 ( .A(A[246]), .B(B[246]), .Z(n40) );
  NAND U36 ( .A(n41), .B(n42), .Z(n39) );
  NANDN U37 ( .A(B[246]), .B(A[246]), .Z(n42) );
  AND U38 ( .A(n43), .B(n44), .Z(n41) );
  NAND U39 ( .A(n45), .B(n46), .Z(n44) );
  NANDN U40 ( .A(A[245]), .B(B[245]), .Z(n46) );
  AND U41 ( .A(n47), .B(n48), .Z(n45) );
  NANDN U42 ( .A(A[244]), .B(B[244]), .Z(n48) );
  NAND U43 ( .A(n49), .B(n50), .Z(n47) );
  NANDN U44 ( .A(B[244]), .B(A[244]), .Z(n50) );
  AND U45 ( .A(n51), .B(n52), .Z(n49) );
  NAND U46 ( .A(n53), .B(n54), .Z(n52) );
  NANDN U47 ( .A(A[243]), .B(B[243]), .Z(n54) );
  AND U48 ( .A(n55), .B(n56), .Z(n53) );
  NANDN U49 ( .A(A[242]), .B(B[242]), .Z(n56) );
  NAND U50 ( .A(n57), .B(n58), .Z(n55) );
  NANDN U51 ( .A(B[242]), .B(A[242]), .Z(n58) );
  AND U52 ( .A(n59), .B(n60), .Z(n57) );
  NAND U53 ( .A(n61), .B(n62), .Z(n60) );
  NANDN U54 ( .A(A[241]), .B(B[241]), .Z(n62) );
  AND U55 ( .A(n63), .B(n64), .Z(n61) );
  NANDN U56 ( .A(A[240]), .B(B[240]), .Z(n64) );
  NAND U57 ( .A(n65), .B(n66), .Z(n63) );
  NANDN U58 ( .A(B[240]), .B(A[240]), .Z(n66) );
  AND U59 ( .A(n67), .B(n68), .Z(n65) );
  NAND U60 ( .A(n69), .B(n70), .Z(n68) );
  NANDN U61 ( .A(A[239]), .B(B[239]), .Z(n70) );
  AND U62 ( .A(n71), .B(n72), .Z(n69) );
  NANDN U63 ( .A(A[238]), .B(B[238]), .Z(n72) );
  NAND U64 ( .A(n73), .B(n74), .Z(n71) );
  NANDN U65 ( .A(B[238]), .B(A[238]), .Z(n74) );
  AND U66 ( .A(n75), .B(n76), .Z(n73) );
  NAND U67 ( .A(n77), .B(n78), .Z(n76) );
  NANDN U68 ( .A(A[237]), .B(B[237]), .Z(n78) );
  AND U69 ( .A(n79), .B(n80), .Z(n77) );
  NANDN U70 ( .A(A[236]), .B(B[236]), .Z(n80) );
  NAND U71 ( .A(n81), .B(n82), .Z(n79) );
  NANDN U72 ( .A(B[236]), .B(A[236]), .Z(n82) );
  AND U73 ( .A(n83), .B(n84), .Z(n81) );
  NAND U74 ( .A(n85), .B(n86), .Z(n84) );
  NANDN U75 ( .A(A[235]), .B(B[235]), .Z(n86) );
  AND U76 ( .A(n87), .B(n88), .Z(n85) );
  NANDN U77 ( .A(A[234]), .B(B[234]), .Z(n88) );
  NAND U78 ( .A(n89), .B(n90), .Z(n87) );
  NANDN U79 ( .A(B[234]), .B(A[234]), .Z(n90) );
  AND U80 ( .A(n91), .B(n92), .Z(n89) );
  NAND U81 ( .A(n93), .B(n94), .Z(n92) );
  NANDN U82 ( .A(A[233]), .B(B[233]), .Z(n94) );
  AND U83 ( .A(n95), .B(n96), .Z(n93) );
  NANDN U84 ( .A(A[232]), .B(B[232]), .Z(n96) );
  NAND U85 ( .A(n97), .B(n98), .Z(n95) );
  NANDN U86 ( .A(B[232]), .B(A[232]), .Z(n98) );
  AND U87 ( .A(n99), .B(n100), .Z(n97) );
  NAND U88 ( .A(n101), .B(n102), .Z(n100) );
  NANDN U89 ( .A(A[231]), .B(B[231]), .Z(n102) );
  AND U90 ( .A(n103), .B(n104), .Z(n101) );
  NANDN U91 ( .A(A[230]), .B(B[230]), .Z(n104) );
  NAND U92 ( .A(n105), .B(n106), .Z(n103) );
  NANDN U93 ( .A(B[230]), .B(A[230]), .Z(n106) );
  AND U94 ( .A(n107), .B(n108), .Z(n105) );
  NAND U95 ( .A(n109), .B(n110), .Z(n108) );
  NANDN U96 ( .A(A[229]), .B(B[229]), .Z(n110) );
  AND U97 ( .A(n111), .B(n112), .Z(n109) );
  NANDN U98 ( .A(A[228]), .B(B[228]), .Z(n112) );
  NAND U99 ( .A(n113), .B(n114), .Z(n111) );
  NANDN U100 ( .A(B[228]), .B(A[228]), .Z(n114) );
  AND U101 ( .A(n115), .B(n116), .Z(n113) );
  NAND U102 ( .A(n117), .B(n118), .Z(n116) );
  NANDN U103 ( .A(A[227]), .B(B[227]), .Z(n118) );
  AND U104 ( .A(n119), .B(n120), .Z(n117) );
  NANDN U105 ( .A(A[226]), .B(B[226]), .Z(n120) );
  NAND U106 ( .A(n121), .B(n122), .Z(n119) );
  NANDN U107 ( .A(B[226]), .B(A[226]), .Z(n122) );
  AND U108 ( .A(n123), .B(n124), .Z(n121) );
  NAND U109 ( .A(n125), .B(n126), .Z(n124) );
  NANDN U110 ( .A(A[225]), .B(B[225]), .Z(n126) );
  AND U111 ( .A(n127), .B(n128), .Z(n125) );
  NANDN U112 ( .A(A[224]), .B(B[224]), .Z(n128) );
  NAND U113 ( .A(n129), .B(n130), .Z(n127) );
  NANDN U114 ( .A(B[224]), .B(A[224]), .Z(n130) );
  AND U115 ( .A(n131), .B(n132), .Z(n129) );
  NAND U116 ( .A(n133), .B(n134), .Z(n132) );
  NANDN U117 ( .A(A[223]), .B(B[223]), .Z(n134) );
  AND U118 ( .A(n135), .B(n136), .Z(n133) );
  NANDN U119 ( .A(A[222]), .B(B[222]), .Z(n136) );
  NAND U120 ( .A(n137), .B(n138), .Z(n135) );
  NANDN U121 ( .A(B[222]), .B(A[222]), .Z(n138) );
  AND U122 ( .A(n139), .B(n140), .Z(n137) );
  NAND U123 ( .A(n141), .B(n142), .Z(n140) );
  NANDN U124 ( .A(A[221]), .B(B[221]), .Z(n142) );
  AND U125 ( .A(n143), .B(n144), .Z(n141) );
  NANDN U126 ( .A(A[220]), .B(B[220]), .Z(n144) );
  NAND U127 ( .A(n145), .B(n146), .Z(n143) );
  NANDN U128 ( .A(B[220]), .B(A[220]), .Z(n146) );
  AND U129 ( .A(n147), .B(n148), .Z(n145) );
  NAND U130 ( .A(n149), .B(n150), .Z(n148) );
  NANDN U131 ( .A(A[219]), .B(B[219]), .Z(n150) );
  AND U132 ( .A(n151), .B(n152), .Z(n149) );
  NANDN U133 ( .A(A[218]), .B(B[218]), .Z(n152) );
  NAND U134 ( .A(n153), .B(n154), .Z(n151) );
  NANDN U135 ( .A(B[218]), .B(A[218]), .Z(n154) );
  AND U136 ( .A(n155), .B(n156), .Z(n153) );
  NAND U137 ( .A(n157), .B(n158), .Z(n156) );
  NANDN U138 ( .A(A[217]), .B(B[217]), .Z(n158) );
  AND U139 ( .A(n159), .B(n160), .Z(n157) );
  NANDN U140 ( .A(A[216]), .B(B[216]), .Z(n160) );
  NAND U141 ( .A(n161), .B(n162), .Z(n159) );
  NANDN U142 ( .A(B[216]), .B(A[216]), .Z(n162) );
  AND U143 ( .A(n163), .B(n164), .Z(n161) );
  NAND U144 ( .A(n165), .B(n166), .Z(n164) );
  NANDN U145 ( .A(A[215]), .B(B[215]), .Z(n166) );
  AND U146 ( .A(n167), .B(n168), .Z(n165) );
  NANDN U147 ( .A(A[214]), .B(B[214]), .Z(n168) );
  NAND U148 ( .A(n169), .B(n170), .Z(n167) );
  NANDN U149 ( .A(B[214]), .B(A[214]), .Z(n170) );
  AND U150 ( .A(n171), .B(n172), .Z(n169) );
  NAND U151 ( .A(n173), .B(n174), .Z(n172) );
  NANDN U152 ( .A(A[213]), .B(B[213]), .Z(n174) );
  AND U153 ( .A(n175), .B(n176), .Z(n173) );
  NANDN U154 ( .A(A[212]), .B(B[212]), .Z(n176) );
  NAND U155 ( .A(n177), .B(n178), .Z(n175) );
  NANDN U156 ( .A(B[212]), .B(A[212]), .Z(n178) );
  AND U157 ( .A(n179), .B(n180), .Z(n177) );
  NAND U158 ( .A(n181), .B(n182), .Z(n180) );
  NANDN U159 ( .A(A[211]), .B(B[211]), .Z(n182) );
  AND U160 ( .A(n183), .B(n184), .Z(n181) );
  NANDN U161 ( .A(A[210]), .B(B[210]), .Z(n184) );
  NAND U162 ( .A(n185), .B(n186), .Z(n183) );
  NANDN U163 ( .A(B[210]), .B(A[210]), .Z(n186) );
  AND U164 ( .A(n187), .B(n188), .Z(n185) );
  NAND U165 ( .A(n189), .B(n190), .Z(n188) );
  NANDN U166 ( .A(A[209]), .B(B[209]), .Z(n190) );
  AND U167 ( .A(n191), .B(n192), .Z(n189) );
  NANDN U168 ( .A(A[208]), .B(B[208]), .Z(n192) );
  NAND U169 ( .A(n193), .B(n194), .Z(n191) );
  NANDN U170 ( .A(B[208]), .B(A[208]), .Z(n194) );
  AND U171 ( .A(n195), .B(n196), .Z(n193) );
  NAND U172 ( .A(n197), .B(n198), .Z(n196) );
  NANDN U173 ( .A(A[207]), .B(B[207]), .Z(n198) );
  AND U174 ( .A(n199), .B(n200), .Z(n197) );
  NANDN U175 ( .A(A[206]), .B(B[206]), .Z(n200) );
  NAND U176 ( .A(n201), .B(n202), .Z(n199) );
  NANDN U177 ( .A(B[206]), .B(A[206]), .Z(n202) );
  AND U178 ( .A(n203), .B(n204), .Z(n201) );
  NAND U179 ( .A(n205), .B(n206), .Z(n204) );
  NANDN U180 ( .A(A[205]), .B(B[205]), .Z(n206) );
  AND U181 ( .A(n207), .B(n208), .Z(n205) );
  NANDN U182 ( .A(A[204]), .B(B[204]), .Z(n208) );
  NAND U183 ( .A(n209), .B(n210), .Z(n207) );
  NANDN U184 ( .A(B[204]), .B(A[204]), .Z(n210) );
  AND U185 ( .A(n211), .B(n212), .Z(n209) );
  NAND U186 ( .A(n213), .B(n214), .Z(n212) );
  NANDN U187 ( .A(A[203]), .B(B[203]), .Z(n214) );
  AND U188 ( .A(n215), .B(n216), .Z(n213) );
  NANDN U189 ( .A(A[202]), .B(B[202]), .Z(n216) );
  NAND U190 ( .A(n217), .B(n218), .Z(n215) );
  NANDN U191 ( .A(B[202]), .B(A[202]), .Z(n218) );
  AND U192 ( .A(n219), .B(n220), .Z(n217) );
  NAND U193 ( .A(n221), .B(n222), .Z(n220) );
  NANDN U194 ( .A(A[201]), .B(B[201]), .Z(n222) );
  AND U195 ( .A(n223), .B(n224), .Z(n221) );
  NANDN U196 ( .A(A[200]), .B(B[200]), .Z(n224) );
  NAND U197 ( .A(n225), .B(n226), .Z(n223) );
  NANDN U198 ( .A(B[200]), .B(A[200]), .Z(n226) );
  AND U199 ( .A(n227), .B(n228), .Z(n225) );
  NAND U200 ( .A(n229), .B(n230), .Z(n228) );
  NANDN U201 ( .A(A[199]), .B(B[199]), .Z(n230) );
  AND U202 ( .A(n231), .B(n232), .Z(n229) );
  NANDN U203 ( .A(A[198]), .B(B[198]), .Z(n232) );
  NAND U204 ( .A(n233), .B(n234), .Z(n231) );
  NANDN U205 ( .A(B[198]), .B(A[198]), .Z(n234) );
  AND U206 ( .A(n235), .B(n236), .Z(n233) );
  NAND U207 ( .A(n237), .B(n238), .Z(n236) );
  NANDN U208 ( .A(A[197]), .B(B[197]), .Z(n238) );
  AND U209 ( .A(n239), .B(n240), .Z(n237) );
  NANDN U210 ( .A(A[196]), .B(B[196]), .Z(n240) );
  NAND U211 ( .A(n241), .B(n242), .Z(n239) );
  NANDN U212 ( .A(B[196]), .B(A[196]), .Z(n242) );
  AND U213 ( .A(n243), .B(n244), .Z(n241) );
  NAND U214 ( .A(n245), .B(n246), .Z(n244) );
  NANDN U215 ( .A(A[195]), .B(B[195]), .Z(n246) );
  AND U216 ( .A(n247), .B(n248), .Z(n245) );
  NANDN U217 ( .A(A[194]), .B(B[194]), .Z(n248) );
  NAND U218 ( .A(n249), .B(n250), .Z(n247) );
  NANDN U219 ( .A(B[194]), .B(A[194]), .Z(n250) );
  AND U220 ( .A(n251), .B(n252), .Z(n249) );
  NAND U221 ( .A(n253), .B(n254), .Z(n252) );
  NANDN U222 ( .A(A[193]), .B(B[193]), .Z(n254) );
  AND U223 ( .A(n255), .B(n256), .Z(n253) );
  NANDN U224 ( .A(A[192]), .B(B[192]), .Z(n256) );
  NAND U225 ( .A(n257), .B(n258), .Z(n255) );
  NANDN U226 ( .A(B[192]), .B(A[192]), .Z(n258) );
  AND U227 ( .A(n259), .B(n260), .Z(n257) );
  NAND U228 ( .A(n261), .B(n262), .Z(n260) );
  NANDN U229 ( .A(A[191]), .B(B[191]), .Z(n262) );
  AND U230 ( .A(n263), .B(n264), .Z(n261) );
  NANDN U231 ( .A(A[190]), .B(B[190]), .Z(n264) );
  NAND U232 ( .A(n265), .B(n266), .Z(n263) );
  NANDN U233 ( .A(B[190]), .B(A[190]), .Z(n266) );
  AND U234 ( .A(n267), .B(n268), .Z(n265) );
  NAND U235 ( .A(n269), .B(n270), .Z(n268) );
  NANDN U236 ( .A(A[189]), .B(B[189]), .Z(n270) );
  AND U237 ( .A(n271), .B(n272), .Z(n269) );
  NANDN U238 ( .A(A[188]), .B(B[188]), .Z(n272) );
  NAND U239 ( .A(n273), .B(n274), .Z(n271) );
  NANDN U240 ( .A(B[188]), .B(A[188]), .Z(n274) );
  AND U241 ( .A(n275), .B(n276), .Z(n273) );
  NAND U242 ( .A(n277), .B(n278), .Z(n276) );
  NANDN U243 ( .A(A[187]), .B(B[187]), .Z(n278) );
  AND U244 ( .A(n279), .B(n280), .Z(n277) );
  NANDN U245 ( .A(A[186]), .B(B[186]), .Z(n280) );
  NAND U246 ( .A(n281), .B(n282), .Z(n279) );
  NANDN U247 ( .A(B[186]), .B(A[186]), .Z(n282) );
  AND U248 ( .A(n283), .B(n284), .Z(n281) );
  NAND U249 ( .A(n285), .B(n286), .Z(n284) );
  NANDN U250 ( .A(A[185]), .B(B[185]), .Z(n286) );
  AND U251 ( .A(n287), .B(n288), .Z(n285) );
  NANDN U252 ( .A(A[184]), .B(B[184]), .Z(n288) );
  NAND U253 ( .A(n289), .B(n290), .Z(n287) );
  NANDN U254 ( .A(B[184]), .B(A[184]), .Z(n290) );
  AND U255 ( .A(n291), .B(n292), .Z(n289) );
  NAND U256 ( .A(n293), .B(n294), .Z(n292) );
  NANDN U257 ( .A(A[183]), .B(B[183]), .Z(n294) );
  AND U258 ( .A(n295), .B(n296), .Z(n293) );
  NANDN U259 ( .A(A[182]), .B(B[182]), .Z(n296) );
  NAND U260 ( .A(n297), .B(n298), .Z(n295) );
  NANDN U261 ( .A(B[182]), .B(A[182]), .Z(n298) );
  AND U262 ( .A(n299), .B(n300), .Z(n297) );
  NAND U263 ( .A(n301), .B(n302), .Z(n300) );
  NANDN U264 ( .A(A[181]), .B(B[181]), .Z(n302) );
  AND U265 ( .A(n303), .B(n304), .Z(n301) );
  NANDN U266 ( .A(A[180]), .B(B[180]), .Z(n304) );
  NAND U267 ( .A(n305), .B(n306), .Z(n303) );
  NANDN U268 ( .A(B[180]), .B(A[180]), .Z(n306) );
  AND U269 ( .A(n307), .B(n308), .Z(n305) );
  NAND U270 ( .A(n309), .B(n310), .Z(n308) );
  NANDN U271 ( .A(A[179]), .B(B[179]), .Z(n310) );
  AND U272 ( .A(n311), .B(n312), .Z(n309) );
  NANDN U273 ( .A(A[178]), .B(B[178]), .Z(n312) );
  NAND U274 ( .A(n313), .B(n314), .Z(n311) );
  NANDN U275 ( .A(B[178]), .B(A[178]), .Z(n314) );
  AND U276 ( .A(n315), .B(n316), .Z(n313) );
  NAND U277 ( .A(n317), .B(n318), .Z(n316) );
  NANDN U278 ( .A(A[177]), .B(B[177]), .Z(n318) );
  AND U279 ( .A(n319), .B(n320), .Z(n317) );
  NANDN U280 ( .A(A[176]), .B(B[176]), .Z(n320) );
  NAND U281 ( .A(n321), .B(n322), .Z(n319) );
  NANDN U282 ( .A(B[176]), .B(A[176]), .Z(n322) );
  AND U283 ( .A(n323), .B(n324), .Z(n321) );
  NAND U284 ( .A(n325), .B(n326), .Z(n324) );
  NANDN U285 ( .A(A[175]), .B(B[175]), .Z(n326) );
  AND U286 ( .A(n327), .B(n328), .Z(n325) );
  NANDN U287 ( .A(A[174]), .B(B[174]), .Z(n328) );
  NAND U288 ( .A(n329), .B(n330), .Z(n327) );
  NANDN U289 ( .A(B[174]), .B(A[174]), .Z(n330) );
  AND U290 ( .A(n331), .B(n332), .Z(n329) );
  NAND U291 ( .A(n333), .B(n334), .Z(n332) );
  NANDN U292 ( .A(A[173]), .B(B[173]), .Z(n334) );
  AND U293 ( .A(n335), .B(n336), .Z(n333) );
  NANDN U294 ( .A(A[172]), .B(B[172]), .Z(n336) );
  NAND U295 ( .A(n337), .B(n338), .Z(n335) );
  NANDN U296 ( .A(B[172]), .B(A[172]), .Z(n338) );
  AND U297 ( .A(n339), .B(n340), .Z(n337) );
  NAND U298 ( .A(n341), .B(n342), .Z(n340) );
  NANDN U299 ( .A(A[171]), .B(B[171]), .Z(n342) );
  AND U300 ( .A(n343), .B(n344), .Z(n341) );
  NANDN U301 ( .A(A[170]), .B(B[170]), .Z(n344) );
  NAND U302 ( .A(n345), .B(n346), .Z(n343) );
  NANDN U303 ( .A(B[170]), .B(A[170]), .Z(n346) );
  AND U304 ( .A(n347), .B(n348), .Z(n345) );
  NAND U305 ( .A(n349), .B(n350), .Z(n348) );
  NANDN U306 ( .A(A[169]), .B(B[169]), .Z(n350) );
  AND U307 ( .A(n351), .B(n352), .Z(n349) );
  NANDN U308 ( .A(A[168]), .B(B[168]), .Z(n352) );
  NAND U309 ( .A(n353), .B(n354), .Z(n351) );
  NANDN U310 ( .A(B[168]), .B(A[168]), .Z(n354) );
  AND U311 ( .A(n355), .B(n356), .Z(n353) );
  NAND U312 ( .A(n357), .B(n358), .Z(n356) );
  NANDN U313 ( .A(A[167]), .B(B[167]), .Z(n358) );
  AND U314 ( .A(n359), .B(n360), .Z(n357) );
  NANDN U315 ( .A(A[166]), .B(B[166]), .Z(n360) );
  NAND U316 ( .A(n361), .B(n362), .Z(n359) );
  NANDN U317 ( .A(B[166]), .B(A[166]), .Z(n362) );
  AND U318 ( .A(n363), .B(n364), .Z(n361) );
  NAND U319 ( .A(n365), .B(n366), .Z(n364) );
  NANDN U320 ( .A(A[165]), .B(B[165]), .Z(n366) );
  AND U321 ( .A(n367), .B(n368), .Z(n365) );
  NANDN U322 ( .A(A[164]), .B(B[164]), .Z(n368) );
  NAND U323 ( .A(n369), .B(n370), .Z(n367) );
  NANDN U324 ( .A(B[164]), .B(A[164]), .Z(n370) );
  AND U325 ( .A(n371), .B(n372), .Z(n369) );
  NAND U326 ( .A(n373), .B(n374), .Z(n372) );
  NANDN U327 ( .A(A[163]), .B(B[163]), .Z(n374) );
  AND U328 ( .A(n375), .B(n376), .Z(n373) );
  NANDN U329 ( .A(A[162]), .B(B[162]), .Z(n376) );
  NAND U330 ( .A(n377), .B(n378), .Z(n375) );
  NANDN U331 ( .A(B[162]), .B(A[162]), .Z(n378) );
  AND U332 ( .A(n379), .B(n380), .Z(n377) );
  NAND U333 ( .A(n381), .B(n382), .Z(n380) );
  NANDN U334 ( .A(A[161]), .B(B[161]), .Z(n382) );
  AND U335 ( .A(n383), .B(n384), .Z(n381) );
  NANDN U336 ( .A(A[160]), .B(B[160]), .Z(n384) );
  NAND U337 ( .A(n385), .B(n386), .Z(n383) );
  NANDN U338 ( .A(B[160]), .B(A[160]), .Z(n386) );
  AND U339 ( .A(n387), .B(n388), .Z(n385) );
  NAND U340 ( .A(n389), .B(n390), .Z(n388) );
  NANDN U341 ( .A(A[159]), .B(B[159]), .Z(n390) );
  AND U342 ( .A(n391), .B(n392), .Z(n389) );
  NANDN U343 ( .A(A[158]), .B(B[158]), .Z(n392) );
  NAND U344 ( .A(n393), .B(n394), .Z(n391) );
  NANDN U345 ( .A(B[158]), .B(A[158]), .Z(n394) );
  AND U346 ( .A(n395), .B(n396), .Z(n393) );
  NAND U347 ( .A(n397), .B(n398), .Z(n396) );
  NANDN U348 ( .A(A[157]), .B(B[157]), .Z(n398) );
  AND U349 ( .A(n399), .B(n400), .Z(n397) );
  NANDN U350 ( .A(A[156]), .B(B[156]), .Z(n400) );
  NAND U351 ( .A(n401), .B(n402), .Z(n399) );
  NANDN U352 ( .A(B[156]), .B(A[156]), .Z(n402) );
  AND U353 ( .A(n403), .B(n404), .Z(n401) );
  NAND U354 ( .A(n405), .B(n406), .Z(n404) );
  NANDN U355 ( .A(A[155]), .B(B[155]), .Z(n406) );
  AND U356 ( .A(n407), .B(n408), .Z(n405) );
  NANDN U357 ( .A(A[154]), .B(B[154]), .Z(n408) );
  NAND U358 ( .A(n409), .B(n410), .Z(n407) );
  NANDN U359 ( .A(B[154]), .B(A[154]), .Z(n410) );
  AND U360 ( .A(n411), .B(n412), .Z(n409) );
  NAND U361 ( .A(n413), .B(n414), .Z(n412) );
  NANDN U362 ( .A(A[153]), .B(B[153]), .Z(n414) );
  AND U363 ( .A(n415), .B(n416), .Z(n413) );
  NANDN U364 ( .A(A[152]), .B(B[152]), .Z(n416) );
  NAND U365 ( .A(n417), .B(n418), .Z(n415) );
  NANDN U366 ( .A(B[152]), .B(A[152]), .Z(n418) );
  AND U367 ( .A(n419), .B(n420), .Z(n417) );
  NAND U368 ( .A(n421), .B(n422), .Z(n420) );
  NANDN U369 ( .A(A[151]), .B(B[151]), .Z(n422) );
  AND U370 ( .A(n423), .B(n424), .Z(n421) );
  NANDN U371 ( .A(A[150]), .B(B[150]), .Z(n424) );
  NAND U372 ( .A(n425), .B(n426), .Z(n423) );
  NANDN U373 ( .A(B[150]), .B(A[150]), .Z(n426) );
  AND U374 ( .A(n427), .B(n428), .Z(n425) );
  NAND U375 ( .A(n429), .B(n430), .Z(n428) );
  NANDN U376 ( .A(A[149]), .B(B[149]), .Z(n430) );
  AND U377 ( .A(n431), .B(n432), .Z(n429) );
  NANDN U378 ( .A(A[148]), .B(B[148]), .Z(n432) );
  NAND U379 ( .A(n433), .B(n434), .Z(n431) );
  NANDN U380 ( .A(B[148]), .B(A[148]), .Z(n434) );
  AND U381 ( .A(n435), .B(n436), .Z(n433) );
  NAND U382 ( .A(n437), .B(n438), .Z(n436) );
  NANDN U383 ( .A(A[147]), .B(B[147]), .Z(n438) );
  AND U384 ( .A(n439), .B(n440), .Z(n437) );
  NANDN U385 ( .A(A[146]), .B(B[146]), .Z(n440) );
  NAND U386 ( .A(n441), .B(n442), .Z(n439) );
  NANDN U387 ( .A(B[146]), .B(A[146]), .Z(n442) );
  AND U388 ( .A(n443), .B(n444), .Z(n441) );
  NAND U389 ( .A(n445), .B(n446), .Z(n444) );
  NANDN U390 ( .A(A[145]), .B(B[145]), .Z(n446) );
  AND U391 ( .A(n447), .B(n448), .Z(n445) );
  NANDN U392 ( .A(A[144]), .B(B[144]), .Z(n448) );
  NAND U393 ( .A(n449), .B(n450), .Z(n447) );
  NANDN U394 ( .A(B[144]), .B(A[144]), .Z(n450) );
  AND U395 ( .A(n451), .B(n452), .Z(n449) );
  NAND U396 ( .A(n453), .B(n454), .Z(n452) );
  NANDN U397 ( .A(A[143]), .B(B[143]), .Z(n454) );
  AND U398 ( .A(n455), .B(n456), .Z(n453) );
  NANDN U399 ( .A(A[142]), .B(B[142]), .Z(n456) );
  NAND U400 ( .A(n457), .B(n458), .Z(n455) );
  NANDN U401 ( .A(B[142]), .B(A[142]), .Z(n458) );
  AND U402 ( .A(n459), .B(n460), .Z(n457) );
  NAND U403 ( .A(n461), .B(n462), .Z(n460) );
  NANDN U404 ( .A(A[141]), .B(B[141]), .Z(n462) );
  AND U405 ( .A(n463), .B(n464), .Z(n461) );
  NANDN U406 ( .A(A[140]), .B(B[140]), .Z(n464) );
  NAND U407 ( .A(n465), .B(n466), .Z(n463) );
  NANDN U408 ( .A(B[140]), .B(A[140]), .Z(n466) );
  AND U409 ( .A(n467), .B(n468), .Z(n465) );
  NAND U410 ( .A(n469), .B(n470), .Z(n468) );
  NANDN U411 ( .A(A[139]), .B(B[139]), .Z(n470) );
  AND U412 ( .A(n471), .B(n472), .Z(n469) );
  NANDN U413 ( .A(A[138]), .B(B[138]), .Z(n472) );
  NAND U414 ( .A(n473), .B(n474), .Z(n471) );
  NANDN U415 ( .A(B[138]), .B(A[138]), .Z(n474) );
  AND U416 ( .A(n475), .B(n476), .Z(n473) );
  NAND U417 ( .A(n477), .B(n478), .Z(n476) );
  NANDN U418 ( .A(A[137]), .B(B[137]), .Z(n478) );
  AND U419 ( .A(n479), .B(n480), .Z(n477) );
  NANDN U420 ( .A(A[136]), .B(B[136]), .Z(n480) );
  NAND U421 ( .A(n481), .B(n482), .Z(n479) );
  NANDN U422 ( .A(B[136]), .B(A[136]), .Z(n482) );
  AND U423 ( .A(n483), .B(n484), .Z(n481) );
  NAND U424 ( .A(n485), .B(n486), .Z(n484) );
  NANDN U425 ( .A(A[135]), .B(B[135]), .Z(n486) );
  AND U426 ( .A(n487), .B(n488), .Z(n485) );
  NANDN U427 ( .A(A[134]), .B(B[134]), .Z(n488) );
  NAND U428 ( .A(n489), .B(n490), .Z(n487) );
  NANDN U429 ( .A(B[134]), .B(A[134]), .Z(n490) );
  AND U430 ( .A(n491), .B(n492), .Z(n489) );
  NAND U431 ( .A(n493), .B(n494), .Z(n492) );
  NANDN U432 ( .A(A[133]), .B(B[133]), .Z(n494) );
  AND U433 ( .A(n495), .B(n496), .Z(n493) );
  NANDN U434 ( .A(A[132]), .B(B[132]), .Z(n496) );
  NAND U435 ( .A(n497), .B(n498), .Z(n495) );
  NANDN U436 ( .A(B[132]), .B(A[132]), .Z(n498) );
  AND U437 ( .A(n499), .B(n500), .Z(n497) );
  NAND U438 ( .A(n501), .B(n502), .Z(n500) );
  NANDN U439 ( .A(A[131]), .B(B[131]), .Z(n502) );
  AND U440 ( .A(n503), .B(n504), .Z(n501) );
  NANDN U441 ( .A(A[130]), .B(B[130]), .Z(n504) );
  NAND U442 ( .A(n505), .B(n506), .Z(n503) );
  NANDN U443 ( .A(B[130]), .B(A[130]), .Z(n506) );
  AND U444 ( .A(n507), .B(n508), .Z(n505) );
  NAND U445 ( .A(n509), .B(n510), .Z(n508) );
  NANDN U446 ( .A(A[129]), .B(B[129]), .Z(n510) );
  AND U447 ( .A(n511), .B(n512), .Z(n509) );
  NANDN U448 ( .A(A[128]), .B(B[128]), .Z(n512) );
  NAND U449 ( .A(n513), .B(n514), .Z(n511) );
  NANDN U450 ( .A(B[128]), .B(A[128]), .Z(n514) );
  AND U451 ( .A(n515), .B(n516), .Z(n513) );
  NAND U452 ( .A(n517), .B(n518), .Z(n516) );
  NANDN U453 ( .A(A[127]), .B(B[127]), .Z(n518) );
  AND U454 ( .A(n519), .B(n520), .Z(n517) );
  NANDN U455 ( .A(A[126]), .B(B[126]), .Z(n520) );
  NAND U456 ( .A(n521), .B(n522), .Z(n519) );
  NANDN U457 ( .A(B[126]), .B(A[126]), .Z(n522) );
  AND U458 ( .A(n523), .B(n524), .Z(n521) );
  NAND U459 ( .A(n525), .B(n526), .Z(n524) );
  NANDN U460 ( .A(A[125]), .B(B[125]), .Z(n526) );
  AND U461 ( .A(n527), .B(n528), .Z(n525) );
  NANDN U462 ( .A(A[124]), .B(B[124]), .Z(n528) );
  NAND U463 ( .A(n529), .B(n530), .Z(n527) );
  NANDN U464 ( .A(B[124]), .B(A[124]), .Z(n530) );
  AND U465 ( .A(n531), .B(n532), .Z(n529) );
  NAND U466 ( .A(n533), .B(n534), .Z(n532) );
  NANDN U467 ( .A(A[123]), .B(B[123]), .Z(n534) );
  AND U468 ( .A(n535), .B(n536), .Z(n533) );
  NANDN U469 ( .A(A[122]), .B(B[122]), .Z(n536) );
  NAND U470 ( .A(n537), .B(n538), .Z(n535) );
  NANDN U471 ( .A(B[122]), .B(A[122]), .Z(n538) );
  AND U472 ( .A(n539), .B(n540), .Z(n537) );
  NAND U473 ( .A(n541), .B(n542), .Z(n540) );
  NANDN U474 ( .A(A[121]), .B(B[121]), .Z(n542) );
  AND U475 ( .A(n543), .B(n544), .Z(n541) );
  NANDN U476 ( .A(A[120]), .B(B[120]), .Z(n544) );
  NAND U477 ( .A(n545), .B(n546), .Z(n543) );
  NANDN U478 ( .A(B[120]), .B(A[120]), .Z(n546) );
  AND U479 ( .A(n547), .B(n548), .Z(n545) );
  NAND U480 ( .A(n549), .B(n550), .Z(n548) );
  NANDN U481 ( .A(A[119]), .B(B[119]), .Z(n550) );
  AND U482 ( .A(n551), .B(n552), .Z(n549) );
  NANDN U483 ( .A(A[118]), .B(B[118]), .Z(n552) );
  NAND U484 ( .A(n553), .B(n554), .Z(n551) );
  NANDN U485 ( .A(B[118]), .B(A[118]), .Z(n554) );
  AND U486 ( .A(n555), .B(n556), .Z(n553) );
  NAND U487 ( .A(n557), .B(n558), .Z(n556) );
  NANDN U488 ( .A(A[117]), .B(B[117]), .Z(n558) );
  AND U489 ( .A(n559), .B(n560), .Z(n557) );
  NANDN U490 ( .A(A[116]), .B(B[116]), .Z(n560) );
  NAND U491 ( .A(n561), .B(n562), .Z(n559) );
  NANDN U492 ( .A(B[116]), .B(A[116]), .Z(n562) );
  AND U493 ( .A(n563), .B(n564), .Z(n561) );
  NAND U494 ( .A(n565), .B(n566), .Z(n564) );
  NANDN U495 ( .A(A[115]), .B(B[115]), .Z(n566) );
  AND U496 ( .A(n567), .B(n568), .Z(n565) );
  NANDN U497 ( .A(A[114]), .B(B[114]), .Z(n568) );
  NAND U498 ( .A(n569), .B(n570), .Z(n567) );
  NANDN U499 ( .A(B[114]), .B(A[114]), .Z(n570) );
  AND U500 ( .A(n571), .B(n572), .Z(n569) );
  NAND U501 ( .A(n573), .B(n574), .Z(n572) );
  NANDN U502 ( .A(A[113]), .B(B[113]), .Z(n574) );
  AND U503 ( .A(n575), .B(n576), .Z(n573) );
  NANDN U504 ( .A(A[112]), .B(B[112]), .Z(n576) );
  NAND U505 ( .A(n577), .B(n578), .Z(n575) );
  NANDN U506 ( .A(B[112]), .B(A[112]), .Z(n578) );
  AND U507 ( .A(n579), .B(n580), .Z(n577) );
  NAND U508 ( .A(n581), .B(n582), .Z(n580) );
  NANDN U509 ( .A(A[111]), .B(B[111]), .Z(n582) );
  AND U510 ( .A(n583), .B(n584), .Z(n581) );
  NANDN U511 ( .A(A[110]), .B(B[110]), .Z(n584) );
  NAND U512 ( .A(n585), .B(n586), .Z(n583) );
  NANDN U513 ( .A(B[110]), .B(A[110]), .Z(n586) );
  AND U514 ( .A(n587), .B(n588), .Z(n585) );
  NAND U515 ( .A(n589), .B(n590), .Z(n588) );
  NANDN U516 ( .A(A[109]), .B(B[109]), .Z(n590) );
  AND U517 ( .A(n591), .B(n592), .Z(n589) );
  NANDN U518 ( .A(A[108]), .B(B[108]), .Z(n592) );
  NAND U519 ( .A(n593), .B(n594), .Z(n591) );
  NANDN U520 ( .A(B[108]), .B(A[108]), .Z(n594) );
  AND U521 ( .A(n595), .B(n596), .Z(n593) );
  NAND U522 ( .A(n597), .B(n598), .Z(n596) );
  NANDN U523 ( .A(A[107]), .B(B[107]), .Z(n598) );
  AND U524 ( .A(n599), .B(n600), .Z(n597) );
  NANDN U525 ( .A(A[106]), .B(B[106]), .Z(n600) );
  NAND U526 ( .A(n601), .B(n602), .Z(n599) );
  NANDN U527 ( .A(B[106]), .B(A[106]), .Z(n602) );
  AND U528 ( .A(n603), .B(n604), .Z(n601) );
  NAND U529 ( .A(n605), .B(n606), .Z(n604) );
  NANDN U530 ( .A(A[105]), .B(B[105]), .Z(n606) );
  AND U531 ( .A(n607), .B(n608), .Z(n605) );
  NANDN U532 ( .A(A[104]), .B(B[104]), .Z(n608) );
  NAND U533 ( .A(n609), .B(n610), .Z(n607) );
  NANDN U534 ( .A(B[104]), .B(A[104]), .Z(n610) );
  AND U535 ( .A(n611), .B(n612), .Z(n609) );
  NAND U536 ( .A(n613), .B(n614), .Z(n612) );
  NANDN U537 ( .A(A[103]), .B(B[103]), .Z(n614) );
  AND U538 ( .A(n615), .B(n616), .Z(n613) );
  NANDN U539 ( .A(A[102]), .B(B[102]), .Z(n616) );
  NAND U540 ( .A(n617), .B(n618), .Z(n615) );
  NANDN U541 ( .A(B[102]), .B(A[102]), .Z(n618) );
  AND U542 ( .A(n619), .B(n620), .Z(n617) );
  NAND U543 ( .A(n621), .B(n622), .Z(n620) );
  NANDN U544 ( .A(A[101]), .B(B[101]), .Z(n622) );
  AND U545 ( .A(n623), .B(n624), .Z(n621) );
  NANDN U546 ( .A(A[100]), .B(B[100]), .Z(n624) );
  NAND U547 ( .A(n625), .B(n626), .Z(n623) );
  NANDN U548 ( .A(B[99]), .B(A[99]), .Z(n626) );
  AND U549 ( .A(n627), .B(n628), .Z(n625) );
  NAND U550 ( .A(n629), .B(n630), .Z(n628) );
  NANDN U551 ( .A(A[99]), .B(B[99]), .Z(n630) );
  AND U552 ( .A(n631), .B(n632), .Z(n629) );
  NANDN U553 ( .A(A[98]), .B(B[98]), .Z(n632) );
  NAND U554 ( .A(n633), .B(n634), .Z(n631) );
  NANDN U555 ( .A(B[98]), .B(A[98]), .Z(n634) );
  AND U556 ( .A(n635), .B(n636), .Z(n633) );
  NAND U557 ( .A(n637), .B(n638), .Z(n636) );
  NANDN U558 ( .A(A[97]), .B(B[97]), .Z(n638) );
  AND U559 ( .A(n639), .B(n640), .Z(n637) );
  NANDN U560 ( .A(A[96]), .B(B[96]), .Z(n640) );
  NAND U561 ( .A(n641), .B(n642), .Z(n639) );
  NANDN U562 ( .A(B[96]), .B(A[96]), .Z(n642) );
  AND U563 ( .A(n643), .B(n644), .Z(n641) );
  NAND U564 ( .A(n645), .B(n646), .Z(n644) );
  NANDN U565 ( .A(A[95]), .B(B[95]), .Z(n646) );
  AND U566 ( .A(n647), .B(n648), .Z(n645) );
  NANDN U567 ( .A(A[94]), .B(B[94]), .Z(n648) );
  NAND U568 ( .A(n649), .B(n650), .Z(n647) );
  NANDN U569 ( .A(B[94]), .B(A[94]), .Z(n650) );
  AND U570 ( .A(n651), .B(n652), .Z(n649) );
  NAND U571 ( .A(n653), .B(n654), .Z(n652) );
  NANDN U572 ( .A(A[93]), .B(B[93]), .Z(n654) );
  AND U573 ( .A(n655), .B(n656), .Z(n653) );
  NANDN U574 ( .A(A[92]), .B(B[92]), .Z(n656) );
  NAND U575 ( .A(n657), .B(n658), .Z(n655) );
  NANDN U576 ( .A(B[92]), .B(A[92]), .Z(n658) );
  AND U577 ( .A(n659), .B(n660), .Z(n657) );
  NAND U578 ( .A(n661), .B(n662), .Z(n660) );
  NANDN U579 ( .A(A[91]), .B(B[91]), .Z(n662) );
  AND U580 ( .A(n663), .B(n664), .Z(n661) );
  NANDN U581 ( .A(A[90]), .B(B[90]), .Z(n664) );
  NAND U582 ( .A(n665), .B(n666), .Z(n663) );
  NANDN U583 ( .A(B[90]), .B(A[90]), .Z(n666) );
  AND U584 ( .A(n667), .B(n668), .Z(n665) );
  NAND U585 ( .A(n669), .B(n670), .Z(n668) );
  NANDN U586 ( .A(A[89]), .B(B[89]), .Z(n670) );
  AND U587 ( .A(n671), .B(n672), .Z(n669) );
  NANDN U588 ( .A(A[88]), .B(B[88]), .Z(n672) );
  NAND U589 ( .A(n673), .B(n674), .Z(n671) );
  NANDN U590 ( .A(B[88]), .B(A[88]), .Z(n674) );
  AND U591 ( .A(n675), .B(n676), .Z(n673) );
  NAND U592 ( .A(n677), .B(n678), .Z(n676) );
  NANDN U593 ( .A(A[87]), .B(B[87]), .Z(n678) );
  AND U594 ( .A(n679), .B(n680), .Z(n677) );
  NANDN U595 ( .A(A[86]), .B(B[86]), .Z(n680) );
  NAND U596 ( .A(n681), .B(n682), .Z(n679) );
  NANDN U597 ( .A(B[86]), .B(A[86]), .Z(n682) );
  AND U598 ( .A(n683), .B(n684), .Z(n681) );
  NAND U599 ( .A(n685), .B(n686), .Z(n684) );
  NANDN U600 ( .A(A[85]), .B(B[85]), .Z(n686) );
  AND U601 ( .A(n687), .B(n688), .Z(n685) );
  NANDN U602 ( .A(A[84]), .B(B[84]), .Z(n688) );
  NAND U603 ( .A(n689), .B(n690), .Z(n687) );
  NANDN U604 ( .A(B[84]), .B(A[84]), .Z(n690) );
  AND U605 ( .A(n691), .B(n692), .Z(n689) );
  NAND U606 ( .A(n693), .B(n694), .Z(n692) );
  NANDN U607 ( .A(A[83]), .B(B[83]), .Z(n694) );
  AND U608 ( .A(n695), .B(n696), .Z(n693) );
  NANDN U609 ( .A(A[82]), .B(B[82]), .Z(n696) );
  NAND U610 ( .A(n697), .B(n698), .Z(n695) );
  NANDN U611 ( .A(B[82]), .B(A[82]), .Z(n698) );
  AND U612 ( .A(n699), .B(n700), .Z(n697) );
  NAND U613 ( .A(n701), .B(n702), .Z(n700) );
  NANDN U614 ( .A(A[81]), .B(B[81]), .Z(n702) );
  AND U615 ( .A(n703), .B(n704), .Z(n701) );
  NANDN U616 ( .A(A[80]), .B(B[80]), .Z(n704) );
  NAND U617 ( .A(n705), .B(n706), .Z(n703) );
  NANDN U618 ( .A(B[80]), .B(A[80]), .Z(n706) );
  AND U619 ( .A(n707), .B(n708), .Z(n705) );
  NAND U620 ( .A(n709), .B(n710), .Z(n708) );
  NANDN U621 ( .A(A[79]), .B(B[79]), .Z(n710) );
  AND U622 ( .A(n711), .B(n712), .Z(n709) );
  NANDN U623 ( .A(A[78]), .B(B[78]), .Z(n712) );
  NAND U624 ( .A(n713), .B(n714), .Z(n711) );
  NANDN U625 ( .A(B[78]), .B(A[78]), .Z(n714) );
  AND U626 ( .A(n715), .B(n716), .Z(n713) );
  NAND U627 ( .A(n717), .B(n718), .Z(n716) );
  NANDN U628 ( .A(A[77]), .B(B[77]), .Z(n718) );
  AND U629 ( .A(n719), .B(n720), .Z(n717) );
  NANDN U630 ( .A(A[76]), .B(B[76]), .Z(n720) );
  NAND U631 ( .A(n721), .B(n722), .Z(n719) );
  NANDN U632 ( .A(B[76]), .B(A[76]), .Z(n722) );
  AND U633 ( .A(n723), .B(n724), .Z(n721) );
  NAND U634 ( .A(n725), .B(n726), .Z(n724) );
  NANDN U635 ( .A(A[75]), .B(B[75]), .Z(n726) );
  AND U636 ( .A(n727), .B(n728), .Z(n725) );
  NANDN U637 ( .A(A[74]), .B(B[74]), .Z(n728) );
  NAND U638 ( .A(n729), .B(n730), .Z(n727) );
  NANDN U639 ( .A(B[74]), .B(A[74]), .Z(n730) );
  AND U640 ( .A(n731), .B(n732), .Z(n729) );
  NAND U641 ( .A(n733), .B(n734), .Z(n732) );
  NANDN U642 ( .A(A[73]), .B(B[73]), .Z(n734) );
  AND U643 ( .A(n735), .B(n736), .Z(n733) );
  NANDN U644 ( .A(A[72]), .B(B[72]), .Z(n736) );
  NAND U645 ( .A(n737), .B(n738), .Z(n735) );
  NANDN U646 ( .A(B[72]), .B(A[72]), .Z(n738) );
  AND U647 ( .A(n739), .B(n740), .Z(n737) );
  NAND U648 ( .A(n741), .B(n742), .Z(n740) );
  NANDN U649 ( .A(A[71]), .B(B[71]), .Z(n742) );
  AND U650 ( .A(n743), .B(n744), .Z(n741) );
  NANDN U651 ( .A(A[70]), .B(B[70]), .Z(n744) );
  NAND U652 ( .A(n745), .B(n746), .Z(n743) );
  NANDN U653 ( .A(B[70]), .B(A[70]), .Z(n746) );
  AND U654 ( .A(n747), .B(n748), .Z(n745) );
  NAND U655 ( .A(n749), .B(n750), .Z(n748) );
  NANDN U656 ( .A(A[69]), .B(B[69]), .Z(n750) );
  AND U657 ( .A(n751), .B(n752), .Z(n749) );
  NANDN U658 ( .A(A[68]), .B(B[68]), .Z(n752) );
  NAND U659 ( .A(n753), .B(n754), .Z(n751) );
  NANDN U660 ( .A(B[68]), .B(A[68]), .Z(n754) );
  AND U661 ( .A(n755), .B(n756), .Z(n753) );
  NAND U662 ( .A(n757), .B(n758), .Z(n756) );
  NANDN U663 ( .A(A[67]), .B(B[67]), .Z(n758) );
  AND U664 ( .A(n759), .B(n760), .Z(n757) );
  NANDN U665 ( .A(A[66]), .B(B[66]), .Z(n760) );
  NAND U666 ( .A(n761), .B(n762), .Z(n759) );
  NANDN U667 ( .A(B[66]), .B(A[66]), .Z(n762) );
  AND U668 ( .A(n763), .B(n764), .Z(n761) );
  NAND U669 ( .A(n765), .B(n766), .Z(n764) );
  NANDN U670 ( .A(A[65]), .B(B[65]), .Z(n766) );
  AND U671 ( .A(n767), .B(n768), .Z(n765) );
  NANDN U672 ( .A(A[64]), .B(B[64]), .Z(n768) );
  NAND U673 ( .A(n769), .B(n770), .Z(n767) );
  NANDN U674 ( .A(B[64]), .B(A[64]), .Z(n770) );
  AND U675 ( .A(n771), .B(n772), .Z(n769) );
  NAND U676 ( .A(n773), .B(n774), .Z(n772) );
  NANDN U677 ( .A(A[63]), .B(B[63]), .Z(n774) );
  AND U678 ( .A(n775), .B(n776), .Z(n773) );
  NANDN U679 ( .A(A[62]), .B(B[62]), .Z(n776) );
  NAND U680 ( .A(n777), .B(n778), .Z(n775) );
  NANDN U681 ( .A(B[62]), .B(A[62]), .Z(n778) );
  AND U682 ( .A(n779), .B(n780), .Z(n777) );
  NAND U683 ( .A(n781), .B(n782), .Z(n780) );
  NANDN U684 ( .A(A[61]), .B(B[61]), .Z(n782) );
  AND U685 ( .A(n783), .B(n784), .Z(n781) );
  NANDN U686 ( .A(A[60]), .B(B[60]), .Z(n784) );
  NAND U687 ( .A(n785), .B(n786), .Z(n783) );
  NANDN U688 ( .A(B[60]), .B(A[60]), .Z(n786) );
  AND U689 ( .A(n787), .B(n788), .Z(n785) );
  NAND U690 ( .A(n789), .B(n790), .Z(n788) );
  NANDN U691 ( .A(A[59]), .B(B[59]), .Z(n790) );
  AND U692 ( .A(n791), .B(n792), .Z(n789) );
  NANDN U693 ( .A(A[58]), .B(B[58]), .Z(n792) );
  NAND U694 ( .A(n793), .B(n794), .Z(n791) );
  NANDN U695 ( .A(B[58]), .B(A[58]), .Z(n794) );
  AND U696 ( .A(n795), .B(n796), .Z(n793) );
  NAND U697 ( .A(n797), .B(n798), .Z(n796) );
  NANDN U698 ( .A(A[57]), .B(B[57]), .Z(n798) );
  AND U699 ( .A(n799), .B(n800), .Z(n797) );
  NANDN U700 ( .A(A[56]), .B(B[56]), .Z(n800) );
  NAND U701 ( .A(n801), .B(n802), .Z(n799) );
  NANDN U702 ( .A(B[56]), .B(A[56]), .Z(n802) );
  AND U703 ( .A(n803), .B(n804), .Z(n801) );
  NAND U704 ( .A(n805), .B(n806), .Z(n804) );
  NANDN U705 ( .A(A[55]), .B(B[55]), .Z(n806) );
  AND U706 ( .A(n807), .B(n808), .Z(n805) );
  NANDN U707 ( .A(A[54]), .B(B[54]), .Z(n808) );
  NAND U708 ( .A(n809), .B(n810), .Z(n807) );
  NANDN U709 ( .A(B[54]), .B(A[54]), .Z(n810) );
  AND U710 ( .A(n811), .B(n812), .Z(n809) );
  NAND U711 ( .A(n813), .B(n814), .Z(n812) );
  NANDN U712 ( .A(A[53]), .B(B[53]), .Z(n814) );
  AND U713 ( .A(n815), .B(n816), .Z(n813) );
  NANDN U714 ( .A(A[52]), .B(B[52]), .Z(n816) );
  NAND U715 ( .A(n817), .B(n818), .Z(n815) );
  NANDN U716 ( .A(B[52]), .B(A[52]), .Z(n818) );
  AND U717 ( .A(n819), .B(n820), .Z(n817) );
  NAND U718 ( .A(n821), .B(n822), .Z(n820) );
  NANDN U719 ( .A(A[51]), .B(B[51]), .Z(n822) );
  AND U720 ( .A(n823), .B(n824), .Z(n821) );
  NANDN U721 ( .A(A[50]), .B(B[50]), .Z(n824) );
  NAND U722 ( .A(n825), .B(n826), .Z(n823) );
  NANDN U723 ( .A(B[50]), .B(A[50]), .Z(n826) );
  AND U724 ( .A(n827), .B(n828), .Z(n825) );
  NAND U725 ( .A(n829), .B(n830), .Z(n828) );
  NANDN U726 ( .A(A[49]), .B(B[49]), .Z(n830) );
  AND U727 ( .A(n831), .B(n832), .Z(n829) );
  NANDN U728 ( .A(A[48]), .B(B[48]), .Z(n832) );
  NAND U729 ( .A(n833), .B(n834), .Z(n831) );
  NANDN U730 ( .A(B[48]), .B(A[48]), .Z(n834) );
  AND U731 ( .A(n835), .B(n836), .Z(n833) );
  NAND U732 ( .A(n837), .B(n838), .Z(n836) );
  NANDN U733 ( .A(A[47]), .B(B[47]), .Z(n838) );
  AND U734 ( .A(n839), .B(n840), .Z(n837) );
  NANDN U735 ( .A(A[46]), .B(B[46]), .Z(n840) );
  NAND U736 ( .A(n841), .B(n842), .Z(n839) );
  NANDN U737 ( .A(B[46]), .B(A[46]), .Z(n842) );
  AND U738 ( .A(n843), .B(n844), .Z(n841) );
  NAND U739 ( .A(n845), .B(n846), .Z(n844) );
  NANDN U740 ( .A(A[45]), .B(B[45]), .Z(n846) );
  AND U741 ( .A(n847), .B(n848), .Z(n845) );
  NANDN U742 ( .A(A[44]), .B(B[44]), .Z(n848) );
  NAND U743 ( .A(n849), .B(n850), .Z(n847) );
  NANDN U744 ( .A(B[44]), .B(A[44]), .Z(n850) );
  AND U745 ( .A(n851), .B(n852), .Z(n849) );
  NAND U746 ( .A(n853), .B(n854), .Z(n852) );
  NANDN U747 ( .A(A[43]), .B(B[43]), .Z(n854) );
  AND U748 ( .A(n855), .B(n856), .Z(n853) );
  NANDN U749 ( .A(A[42]), .B(B[42]), .Z(n856) );
  NAND U750 ( .A(n857), .B(n858), .Z(n855) );
  NANDN U751 ( .A(B[42]), .B(A[42]), .Z(n858) );
  AND U752 ( .A(n859), .B(n860), .Z(n857) );
  NAND U753 ( .A(n861), .B(n862), .Z(n860) );
  NANDN U754 ( .A(A[41]), .B(B[41]), .Z(n862) );
  AND U755 ( .A(n863), .B(n864), .Z(n861) );
  NANDN U756 ( .A(A[40]), .B(B[40]), .Z(n864) );
  NAND U757 ( .A(n865), .B(n866), .Z(n863) );
  NANDN U758 ( .A(B[40]), .B(A[40]), .Z(n866) );
  AND U759 ( .A(n867), .B(n868), .Z(n865) );
  NAND U760 ( .A(n869), .B(n870), .Z(n868) );
  NANDN U761 ( .A(A[39]), .B(B[39]), .Z(n870) );
  AND U762 ( .A(n871), .B(n872), .Z(n869) );
  NANDN U763 ( .A(A[38]), .B(B[38]), .Z(n872) );
  NAND U764 ( .A(n873), .B(n874), .Z(n871) );
  NANDN U765 ( .A(B[38]), .B(A[38]), .Z(n874) );
  AND U766 ( .A(n875), .B(n876), .Z(n873) );
  NAND U767 ( .A(n877), .B(n878), .Z(n876) );
  NANDN U768 ( .A(A[37]), .B(B[37]), .Z(n878) );
  AND U769 ( .A(n879), .B(n880), .Z(n877) );
  NANDN U770 ( .A(A[36]), .B(B[36]), .Z(n880) );
  NAND U771 ( .A(n881), .B(n882), .Z(n879) );
  NANDN U772 ( .A(B[36]), .B(A[36]), .Z(n882) );
  AND U773 ( .A(n883), .B(n884), .Z(n881) );
  NAND U774 ( .A(n885), .B(n886), .Z(n884) );
  NANDN U775 ( .A(A[35]), .B(B[35]), .Z(n886) );
  AND U776 ( .A(n887), .B(n888), .Z(n885) );
  NANDN U777 ( .A(A[34]), .B(B[34]), .Z(n888) );
  NAND U778 ( .A(n889), .B(n890), .Z(n887) );
  NANDN U779 ( .A(B[34]), .B(A[34]), .Z(n890) );
  AND U780 ( .A(n891), .B(n892), .Z(n889) );
  NAND U781 ( .A(n893), .B(n894), .Z(n892) );
  NANDN U782 ( .A(A[33]), .B(B[33]), .Z(n894) );
  AND U783 ( .A(n895), .B(n896), .Z(n893) );
  NANDN U784 ( .A(A[32]), .B(B[32]), .Z(n896) );
  NAND U785 ( .A(n897), .B(n898), .Z(n895) );
  NANDN U786 ( .A(B[32]), .B(A[32]), .Z(n898) );
  AND U787 ( .A(n899), .B(n900), .Z(n897) );
  NAND U788 ( .A(n901), .B(n902), .Z(n900) );
  NANDN U789 ( .A(A[31]), .B(B[31]), .Z(n902) );
  AND U790 ( .A(n903), .B(n904), .Z(n901) );
  NANDN U791 ( .A(A[30]), .B(B[30]), .Z(n904) );
  NAND U792 ( .A(n905), .B(n906), .Z(n903) );
  NANDN U793 ( .A(B[30]), .B(A[30]), .Z(n906) );
  AND U794 ( .A(n907), .B(n908), .Z(n905) );
  NAND U795 ( .A(n909), .B(n910), .Z(n908) );
  NANDN U796 ( .A(A[29]), .B(B[29]), .Z(n910) );
  AND U797 ( .A(n911), .B(n912), .Z(n909) );
  NANDN U798 ( .A(A[28]), .B(B[28]), .Z(n912) );
  NAND U799 ( .A(n913), .B(n914), .Z(n911) );
  NANDN U800 ( .A(B[28]), .B(A[28]), .Z(n914) );
  AND U801 ( .A(n915), .B(n916), .Z(n913) );
  NAND U802 ( .A(n917), .B(n918), .Z(n916) );
  NANDN U803 ( .A(A[27]), .B(B[27]), .Z(n918) );
  AND U804 ( .A(n919), .B(n920), .Z(n917) );
  NANDN U805 ( .A(A[26]), .B(B[26]), .Z(n920) );
  NAND U806 ( .A(n921), .B(n922), .Z(n919) );
  NANDN U807 ( .A(B[26]), .B(A[26]), .Z(n922) );
  AND U808 ( .A(n923), .B(n924), .Z(n921) );
  NAND U809 ( .A(n925), .B(n926), .Z(n924) );
  NANDN U810 ( .A(A[25]), .B(B[25]), .Z(n926) );
  AND U811 ( .A(n927), .B(n928), .Z(n925) );
  NANDN U812 ( .A(A[24]), .B(B[24]), .Z(n928) );
  NAND U813 ( .A(n929), .B(n930), .Z(n927) );
  NANDN U814 ( .A(B[24]), .B(A[24]), .Z(n930) );
  AND U815 ( .A(n931), .B(n932), .Z(n929) );
  NAND U816 ( .A(n933), .B(n934), .Z(n932) );
  NANDN U817 ( .A(A[23]), .B(B[23]), .Z(n934) );
  AND U818 ( .A(n935), .B(n936), .Z(n933) );
  NANDN U819 ( .A(A[22]), .B(B[22]), .Z(n936) );
  NAND U820 ( .A(n937), .B(n938), .Z(n935) );
  NANDN U821 ( .A(B[22]), .B(A[22]), .Z(n938) );
  AND U822 ( .A(n939), .B(n940), .Z(n937) );
  NAND U823 ( .A(n941), .B(n942), .Z(n940) );
  NANDN U824 ( .A(A[21]), .B(B[21]), .Z(n942) );
  AND U825 ( .A(n943), .B(n944), .Z(n941) );
  NANDN U826 ( .A(A[20]), .B(B[20]), .Z(n944) );
  NAND U827 ( .A(n945), .B(n946), .Z(n943) );
  NANDN U828 ( .A(B[20]), .B(A[20]), .Z(n946) );
  AND U829 ( .A(n947), .B(n948), .Z(n945) );
  NAND U830 ( .A(n949), .B(n950), .Z(n948) );
  NANDN U831 ( .A(A[19]), .B(B[19]), .Z(n950) );
  AND U832 ( .A(n951), .B(n952), .Z(n949) );
  NANDN U833 ( .A(A[18]), .B(B[18]), .Z(n952) );
  NAND U834 ( .A(n953), .B(n954), .Z(n951) );
  NANDN U835 ( .A(B[18]), .B(A[18]), .Z(n954) );
  AND U836 ( .A(n955), .B(n956), .Z(n953) );
  NAND U837 ( .A(n957), .B(n958), .Z(n956) );
  NANDN U838 ( .A(A[17]), .B(B[17]), .Z(n958) );
  AND U839 ( .A(n959), .B(n960), .Z(n957) );
  NANDN U840 ( .A(A[16]), .B(B[16]), .Z(n960) );
  NAND U841 ( .A(n961), .B(n962), .Z(n959) );
  NANDN U842 ( .A(B[16]), .B(A[16]), .Z(n962) );
  AND U843 ( .A(n963), .B(n964), .Z(n961) );
  NAND U844 ( .A(n965), .B(n966), .Z(n964) );
  NANDN U845 ( .A(A[15]), .B(B[15]), .Z(n966) );
  AND U846 ( .A(n967), .B(n968), .Z(n965) );
  NANDN U847 ( .A(A[14]), .B(B[14]), .Z(n968) );
  NAND U848 ( .A(n969), .B(n970), .Z(n967) );
  NANDN U849 ( .A(B[14]), .B(A[14]), .Z(n970) );
  AND U850 ( .A(n971), .B(n972), .Z(n969) );
  NAND U851 ( .A(n973), .B(n974), .Z(n972) );
  NANDN U852 ( .A(A[13]), .B(B[13]), .Z(n974) );
  AND U853 ( .A(n975), .B(n976), .Z(n973) );
  NANDN U854 ( .A(A[12]), .B(B[12]), .Z(n976) );
  NAND U855 ( .A(n977), .B(n978), .Z(n975) );
  NANDN U856 ( .A(B[12]), .B(A[12]), .Z(n978) );
  AND U857 ( .A(n979), .B(n980), .Z(n977) );
  NAND U858 ( .A(n981), .B(n982), .Z(n980) );
  NANDN U859 ( .A(A[11]), .B(B[11]), .Z(n982) );
  AND U860 ( .A(n983), .B(n984), .Z(n981) );
  NANDN U861 ( .A(A[10]), .B(B[10]), .Z(n984) );
  NAND U862 ( .A(n985), .B(n986), .Z(n983) );
  NANDN U863 ( .A(B[9]), .B(A[9]), .Z(n986) );
  AND U864 ( .A(n987), .B(n988), .Z(n985) );
  NAND U865 ( .A(n989), .B(n990), .Z(n988) );
  NANDN U866 ( .A(A[9]), .B(B[9]), .Z(n990) );
  AND U867 ( .A(n991), .B(n992), .Z(n989) );
  NANDN U868 ( .A(A[8]), .B(B[8]), .Z(n992) );
  NAND U869 ( .A(n993), .B(n994), .Z(n991) );
  NANDN U870 ( .A(B[8]), .B(A[8]), .Z(n994) );
  AND U871 ( .A(n995), .B(n996), .Z(n993) );
  NAND U872 ( .A(n997), .B(n998), .Z(n996) );
  NANDN U873 ( .A(A[7]), .B(B[7]), .Z(n998) );
  AND U874 ( .A(n999), .B(n1000), .Z(n997) );
  NANDN U875 ( .A(A[6]), .B(B[6]), .Z(n1000) );
  NAND U876 ( .A(n1001), .B(n1002), .Z(n999) );
  NANDN U877 ( .A(B[6]), .B(A[6]), .Z(n1002) );
  AND U878 ( .A(n1003), .B(n1004), .Z(n1001) );
  NAND U879 ( .A(n1005), .B(n1006), .Z(n1004) );
  NANDN U880 ( .A(A[5]), .B(B[5]), .Z(n1006) );
  AND U881 ( .A(n1007), .B(n1008), .Z(n1005) );
  NANDN U882 ( .A(A[4]), .B(B[4]), .Z(n1008) );
  NAND U883 ( .A(n1009), .B(n1010), .Z(n1007) );
  NANDN U884 ( .A(B[4]), .B(A[4]), .Z(n1010) );
  AND U885 ( .A(n1011), .B(n1012), .Z(n1009) );
  NAND U886 ( .A(n1013), .B(n1014), .Z(n1012) );
  NANDN U887 ( .A(A[3]), .B(B[3]), .Z(n1014) );
  AND U888 ( .A(n1015), .B(n1016), .Z(n1013) );
  NANDN U889 ( .A(A[2]), .B(B[2]), .Z(n1016) );
  NAND U890 ( .A(n1017), .B(n1018), .Z(n1015) );
  NANDN U891 ( .A(B[2]), .B(A[2]), .Z(n1018) );
  AND U892 ( .A(n1019), .B(n1020), .Z(n1017) );
  NANDN U893 ( .A(B[1]), .B(n1021), .Z(n1020) );
  NANDN U894 ( .A(A[1]), .B(n1022), .Z(n1021) );
  NANDN U895 ( .A(n1022), .B(A[1]), .Z(n1019) );
  ANDN U896 ( .B(B[0]), .A(A[0]), .Z(n1022) );
  NANDN U897 ( .A(B[3]), .B(A[3]), .Z(n1011) );
  NANDN U898 ( .A(B[5]), .B(A[5]), .Z(n1003) );
  NANDN U899 ( .A(B[7]), .B(A[7]), .Z(n995) );
  NANDN U900 ( .A(B[10]), .B(A[10]), .Z(n987) );
  NANDN U901 ( .A(B[11]), .B(A[11]), .Z(n979) );
  NANDN U902 ( .A(B[13]), .B(A[13]), .Z(n971) );
  NANDN U903 ( .A(B[15]), .B(A[15]), .Z(n963) );
  NANDN U904 ( .A(B[17]), .B(A[17]), .Z(n955) );
  NANDN U905 ( .A(B[19]), .B(A[19]), .Z(n947) );
  NANDN U906 ( .A(B[21]), .B(A[21]), .Z(n939) );
  NANDN U907 ( .A(B[23]), .B(A[23]), .Z(n931) );
  NANDN U908 ( .A(B[25]), .B(A[25]), .Z(n923) );
  NANDN U909 ( .A(B[27]), .B(A[27]), .Z(n915) );
  NANDN U910 ( .A(B[29]), .B(A[29]), .Z(n907) );
  NANDN U911 ( .A(B[31]), .B(A[31]), .Z(n899) );
  NANDN U912 ( .A(B[33]), .B(A[33]), .Z(n891) );
  NANDN U913 ( .A(B[35]), .B(A[35]), .Z(n883) );
  NANDN U914 ( .A(B[37]), .B(A[37]), .Z(n875) );
  NANDN U915 ( .A(B[39]), .B(A[39]), .Z(n867) );
  NANDN U916 ( .A(B[41]), .B(A[41]), .Z(n859) );
  NANDN U917 ( .A(B[43]), .B(A[43]), .Z(n851) );
  NANDN U918 ( .A(B[45]), .B(A[45]), .Z(n843) );
  NANDN U919 ( .A(B[47]), .B(A[47]), .Z(n835) );
  NANDN U920 ( .A(B[49]), .B(A[49]), .Z(n827) );
  NANDN U921 ( .A(B[51]), .B(A[51]), .Z(n819) );
  NANDN U922 ( .A(B[53]), .B(A[53]), .Z(n811) );
  NANDN U923 ( .A(B[55]), .B(A[55]), .Z(n803) );
  NANDN U924 ( .A(B[57]), .B(A[57]), .Z(n795) );
  NANDN U925 ( .A(B[59]), .B(A[59]), .Z(n787) );
  NANDN U926 ( .A(B[61]), .B(A[61]), .Z(n779) );
  NANDN U927 ( .A(B[63]), .B(A[63]), .Z(n771) );
  NANDN U928 ( .A(B[65]), .B(A[65]), .Z(n763) );
  NANDN U929 ( .A(B[67]), .B(A[67]), .Z(n755) );
  NANDN U930 ( .A(B[69]), .B(A[69]), .Z(n747) );
  NANDN U931 ( .A(B[71]), .B(A[71]), .Z(n739) );
  NANDN U932 ( .A(B[73]), .B(A[73]), .Z(n731) );
  NANDN U933 ( .A(B[75]), .B(A[75]), .Z(n723) );
  NANDN U934 ( .A(B[77]), .B(A[77]), .Z(n715) );
  NANDN U935 ( .A(B[79]), .B(A[79]), .Z(n707) );
  NANDN U936 ( .A(B[81]), .B(A[81]), .Z(n699) );
  NANDN U937 ( .A(B[83]), .B(A[83]), .Z(n691) );
  NANDN U938 ( .A(B[85]), .B(A[85]), .Z(n683) );
  NANDN U939 ( .A(B[87]), .B(A[87]), .Z(n675) );
  NANDN U940 ( .A(B[89]), .B(A[89]), .Z(n667) );
  NANDN U941 ( .A(B[91]), .B(A[91]), .Z(n659) );
  NANDN U942 ( .A(B[93]), .B(A[93]), .Z(n651) );
  NANDN U943 ( .A(B[95]), .B(A[95]), .Z(n643) );
  NANDN U944 ( .A(B[97]), .B(A[97]), .Z(n635) );
  NANDN U945 ( .A(B[100]), .B(A[100]), .Z(n627) );
  NANDN U946 ( .A(B[101]), .B(A[101]), .Z(n619) );
  NANDN U947 ( .A(B[103]), .B(A[103]), .Z(n611) );
  NANDN U948 ( .A(B[105]), .B(A[105]), .Z(n603) );
  NANDN U949 ( .A(B[107]), .B(A[107]), .Z(n595) );
  NANDN U950 ( .A(B[109]), .B(A[109]), .Z(n587) );
  NANDN U951 ( .A(B[111]), .B(A[111]), .Z(n579) );
  NANDN U952 ( .A(B[113]), .B(A[113]), .Z(n571) );
  NANDN U953 ( .A(B[115]), .B(A[115]), .Z(n563) );
  NANDN U954 ( .A(B[117]), .B(A[117]), .Z(n555) );
  NANDN U955 ( .A(B[119]), .B(A[119]), .Z(n547) );
  NANDN U956 ( .A(B[121]), .B(A[121]), .Z(n539) );
  NANDN U957 ( .A(B[123]), .B(A[123]), .Z(n531) );
  NANDN U958 ( .A(B[125]), .B(A[125]), .Z(n523) );
  NANDN U959 ( .A(B[127]), .B(A[127]), .Z(n515) );
  NANDN U960 ( .A(B[129]), .B(A[129]), .Z(n507) );
  NANDN U961 ( .A(B[131]), .B(A[131]), .Z(n499) );
  NANDN U962 ( .A(B[133]), .B(A[133]), .Z(n491) );
  NANDN U963 ( .A(B[135]), .B(A[135]), .Z(n483) );
  NANDN U964 ( .A(B[137]), .B(A[137]), .Z(n475) );
  NANDN U965 ( .A(B[139]), .B(A[139]), .Z(n467) );
  NANDN U966 ( .A(B[141]), .B(A[141]), .Z(n459) );
  NANDN U967 ( .A(B[143]), .B(A[143]), .Z(n451) );
  NANDN U968 ( .A(B[145]), .B(A[145]), .Z(n443) );
  NANDN U969 ( .A(B[147]), .B(A[147]), .Z(n435) );
  NANDN U970 ( .A(B[149]), .B(A[149]), .Z(n427) );
  NANDN U971 ( .A(B[151]), .B(A[151]), .Z(n419) );
  NANDN U972 ( .A(B[153]), .B(A[153]), .Z(n411) );
  NANDN U973 ( .A(B[155]), .B(A[155]), .Z(n403) );
  NANDN U974 ( .A(B[157]), .B(A[157]), .Z(n395) );
  NANDN U975 ( .A(B[159]), .B(A[159]), .Z(n387) );
  NANDN U976 ( .A(B[161]), .B(A[161]), .Z(n379) );
  NANDN U977 ( .A(B[163]), .B(A[163]), .Z(n371) );
  NANDN U978 ( .A(B[165]), .B(A[165]), .Z(n363) );
  NANDN U979 ( .A(B[167]), .B(A[167]), .Z(n355) );
  NANDN U980 ( .A(B[169]), .B(A[169]), .Z(n347) );
  NANDN U981 ( .A(B[171]), .B(A[171]), .Z(n339) );
  NANDN U982 ( .A(B[173]), .B(A[173]), .Z(n331) );
  NANDN U983 ( .A(B[175]), .B(A[175]), .Z(n323) );
  NANDN U984 ( .A(B[177]), .B(A[177]), .Z(n315) );
  NANDN U985 ( .A(B[179]), .B(A[179]), .Z(n307) );
  NANDN U986 ( .A(B[181]), .B(A[181]), .Z(n299) );
  NANDN U987 ( .A(B[183]), .B(A[183]), .Z(n291) );
  NANDN U988 ( .A(B[185]), .B(A[185]), .Z(n283) );
  NANDN U989 ( .A(B[187]), .B(A[187]), .Z(n275) );
  NANDN U990 ( .A(B[189]), .B(A[189]), .Z(n267) );
  NANDN U991 ( .A(B[191]), .B(A[191]), .Z(n259) );
  NANDN U992 ( .A(B[193]), .B(A[193]), .Z(n251) );
  NANDN U993 ( .A(B[195]), .B(A[195]), .Z(n243) );
  NANDN U994 ( .A(B[197]), .B(A[197]), .Z(n235) );
  NANDN U995 ( .A(B[199]), .B(A[199]), .Z(n227) );
  NANDN U996 ( .A(B[201]), .B(A[201]), .Z(n219) );
  NANDN U997 ( .A(B[203]), .B(A[203]), .Z(n211) );
  NANDN U998 ( .A(B[205]), .B(A[205]), .Z(n203) );
  NANDN U999 ( .A(B[207]), .B(A[207]), .Z(n195) );
  NANDN U1000 ( .A(B[209]), .B(A[209]), .Z(n187) );
  NANDN U1001 ( .A(B[211]), .B(A[211]), .Z(n179) );
  NANDN U1002 ( .A(B[213]), .B(A[213]), .Z(n171) );
  NANDN U1003 ( .A(B[215]), .B(A[215]), .Z(n163) );
  NANDN U1004 ( .A(B[217]), .B(A[217]), .Z(n155) );
  NANDN U1005 ( .A(B[219]), .B(A[219]), .Z(n147) );
  NANDN U1006 ( .A(B[221]), .B(A[221]), .Z(n139) );
  NANDN U1007 ( .A(B[223]), .B(A[223]), .Z(n131) );
  NANDN U1008 ( .A(B[225]), .B(A[225]), .Z(n123) );
  NANDN U1009 ( .A(B[227]), .B(A[227]), .Z(n115) );
  NANDN U1010 ( .A(B[229]), .B(A[229]), .Z(n107) );
  NANDN U1011 ( .A(B[231]), .B(A[231]), .Z(n99) );
  NANDN U1012 ( .A(B[233]), .B(A[233]), .Z(n91) );
  NANDN U1013 ( .A(B[235]), .B(A[235]), .Z(n83) );
  NANDN U1014 ( .A(B[237]), .B(A[237]), .Z(n75) );
  NANDN U1015 ( .A(B[239]), .B(A[239]), .Z(n67) );
  NANDN U1016 ( .A(B[241]), .B(A[241]), .Z(n59) );
  NANDN U1017 ( .A(B[243]), .B(A[243]), .Z(n51) );
  NANDN U1018 ( .A(B[245]), .B(A[245]), .Z(n43) );
  NANDN U1019 ( .A(B[247]), .B(A[247]), .Z(n35) );
  NANDN U1020 ( .A(B[249]), .B(A[249]), .Z(n27) );
  NANDN U1021 ( .A(B[251]), .B(A[251]), .Z(n19) );
  NANDN U1022 ( .A(B[253]), .B(A[253]), .Z(n11) );
  NANDN U1023 ( .A(A[255]), .B(B[255]), .Z(n3) );
endmodule


module modmult_step_N256_3_DW01_add_0 ( A, B, CI, SUM, CO );
  input [257:0] A;
  input [257:0] B;
  output [257:0] SUM;
  input CI;
  output CO;
  wire   \B[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56,
         n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210, n211, n212, n213, n214, n215, n216, n217, n218, n219, n220,
         n221, n222, n223, n224, n225, n226, n227, n228, n229, n230, n231,
         n232, n233, n234, n235, n236, n237, n238, n239, n240, n241, n242,
         n243, n244, n245, n246, n247, n248, n249, n250, n251, n252, n253,
         n254, n255, n256, n257, n258, n259, n260, n261, n262, n263, n264,
         n265, n266, n267, n268, n269, n270, n271, n272, n273, n274, n275,
         n276, n277, n278, n279, n280, n281, n282, n283, n284, n285, n286,
         n287, n288, n289, n290, n291, n292, n293, n294, n295, n296, n297,
         n298, n299, n300, n301, n302, n303, n304, n305, n306, n307, n308,
         n309, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n327, n328, n329, n330,
         n331, n332, n333, n334, n335, n336, n337, n338, n339, n340, n341,
         n342, n343, n344, n345, n346, n347, n348, n349, n350, n351, n352,
         n353, n354, n355, n356, n357, n358, n359, n360, n361, n362, n363,
         n364, n365, n366, n367, n368, n369, n370, n371, n372, n373, n374,
         n375, n376, n377, n378, n379, n380, n381, n382, n383, n384, n385,
         n386, n387, n388, n389, n390, n391, n392, n393, n394, n395, n396,
         n397, n398, n399, n400, n401, n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161,
         n1162, n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171,
         n1172, n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181,
         n1182, n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191,
         n1192, n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201,
         n1202, n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211,
         n1212, n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221,
         n1222, n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231,
         n1232, n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241,
         n1242, n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251,
         n1252, n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261,
         n1262, n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271,
         n1272;
  assign SUM[0] = \B[0] ;
  assign \B[0]  = B[0];

  XNOR U1 ( .A(n1), .B(n2), .Z(SUM[9]) );
  XNOR U2 ( .A(B[9]), .B(A[9]), .Z(n2) );
  XNOR U3 ( .A(n3), .B(n4), .Z(SUM[99]) );
  XNOR U4 ( .A(B[99]), .B(A[99]), .Z(n4) );
  XOR U5 ( .A(n5), .B(n6), .Z(SUM[98]) );
  XNOR U6 ( .A(B[98]), .B(A[98]), .Z(n6) );
  XOR U7 ( .A(n7), .B(n8), .Z(SUM[97]) );
  XNOR U8 ( .A(B[97]), .B(A[97]), .Z(n8) );
  XOR U9 ( .A(n9), .B(n10), .Z(SUM[96]) );
  XNOR U10 ( .A(B[96]), .B(A[96]), .Z(n10) );
  XOR U11 ( .A(n11), .B(n12), .Z(SUM[95]) );
  XNOR U12 ( .A(B[95]), .B(A[95]), .Z(n12) );
  XOR U13 ( .A(n13), .B(n14), .Z(SUM[94]) );
  XNOR U14 ( .A(B[94]), .B(A[94]), .Z(n14) );
  XOR U15 ( .A(n15), .B(n16), .Z(SUM[93]) );
  XNOR U16 ( .A(B[93]), .B(A[93]), .Z(n16) );
  XOR U17 ( .A(n17), .B(n18), .Z(SUM[92]) );
  XNOR U18 ( .A(B[92]), .B(A[92]), .Z(n18) );
  XOR U19 ( .A(n19), .B(n20), .Z(SUM[91]) );
  XNOR U20 ( .A(B[91]), .B(A[91]), .Z(n20) );
  XOR U21 ( .A(n21), .B(n22), .Z(SUM[90]) );
  XNOR U22 ( .A(B[90]), .B(A[90]), .Z(n22) );
  XOR U23 ( .A(n23), .B(n24), .Z(SUM[8]) );
  XNOR U24 ( .A(B[8]), .B(A[8]), .Z(n24) );
  XOR U25 ( .A(n25), .B(n26), .Z(SUM[89]) );
  XNOR U26 ( .A(B[89]), .B(A[89]), .Z(n26) );
  XOR U27 ( .A(n27), .B(n28), .Z(SUM[88]) );
  XNOR U28 ( .A(B[88]), .B(A[88]), .Z(n28) );
  XOR U29 ( .A(n29), .B(n30), .Z(SUM[87]) );
  XNOR U30 ( .A(B[87]), .B(A[87]), .Z(n30) );
  XOR U31 ( .A(n31), .B(n32), .Z(SUM[86]) );
  XNOR U32 ( .A(B[86]), .B(A[86]), .Z(n32) );
  XOR U33 ( .A(n33), .B(n34), .Z(SUM[85]) );
  XNOR U34 ( .A(B[85]), .B(A[85]), .Z(n34) );
  XOR U35 ( .A(n35), .B(n36), .Z(SUM[84]) );
  XNOR U36 ( .A(B[84]), .B(A[84]), .Z(n36) );
  XOR U37 ( .A(n37), .B(n38), .Z(SUM[83]) );
  XNOR U38 ( .A(B[83]), .B(A[83]), .Z(n38) );
  XOR U39 ( .A(n39), .B(n40), .Z(SUM[82]) );
  XNOR U40 ( .A(B[82]), .B(A[82]), .Z(n40) );
  XOR U41 ( .A(n41), .B(n42), .Z(SUM[81]) );
  XNOR U42 ( .A(B[81]), .B(A[81]), .Z(n42) );
  XOR U43 ( .A(n43), .B(n44), .Z(SUM[80]) );
  XNOR U44 ( .A(B[80]), .B(A[80]), .Z(n44) );
  XOR U45 ( .A(n45), .B(n46), .Z(SUM[7]) );
  XNOR U46 ( .A(B[7]), .B(A[7]), .Z(n46) );
  XOR U47 ( .A(n47), .B(n48), .Z(SUM[79]) );
  XNOR U48 ( .A(B[79]), .B(A[79]), .Z(n48) );
  XOR U49 ( .A(n49), .B(n50), .Z(SUM[78]) );
  XNOR U50 ( .A(B[78]), .B(A[78]), .Z(n50) );
  XOR U51 ( .A(n51), .B(n52), .Z(SUM[77]) );
  XNOR U52 ( .A(B[77]), .B(A[77]), .Z(n52) );
  XOR U53 ( .A(n53), .B(n54), .Z(SUM[76]) );
  XNOR U54 ( .A(B[76]), .B(A[76]), .Z(n54) );
  XOR U55 ( .A(n55), .B(n56), .Z(SUM[75]) );
  XNOR U56 ( .A(B[75]), .B(A[75]), .Z(n56) );
  XOR U57 ( .A(n57), .B(n58), .Z(SUM[74]) );
  XNOR U58 ( .A(B[74]), .B(A[74]), .Z(n58) );
  XOR U59 ( .A(n59), .B(n60), .Z(SUM[73]) );
  XNOR U60 ( .A(B[73]), .B(A[73]), .Z(n60) );
  XOR U61 ( .A(n61), .B(n62), .Z(SUM[72]) );
  XNOR U62 ( .A(B[72]), .B(A[72]), .Z(n62) );
  XOR U63 ( .A(n63), .B(n64), .Z(SUM[71]) );
  XNOR U64 ( .A(B[71]), .B(A[71]), .Z(n64) );
  XOR U65 ( .A(n65), .B(n66), .Z(SUM[70]) );
  XNOR U66 ( .A(B[70]), .B(A[70]), .Z(n66) );
  XOR U67 ( .A(n67), .B(n68), .Z(SUM[6]) );
  XNOR U68 ( .A(B[6]), .B(A[6]), .Z(n68) );
  XOR U69 ( .A(n69), .B(n70), .Z(SUM[69]) );
  XNOR U70 ( .A(B[69]), .B(A[69]), .Z(n70) );
  XOR U71 ( .A(n71), .B(n72), .Z(SUM[68]) );
  XNOR U72 ( .A(B[68]), .B(A[68]), .Z(n72) );
  XOR U73 ( .A(n73), .B(n74), .Z(SUM[67]) );
  XNOR U74 ( .A(B[67]), .B(A[67]), .Z(n74) );
  XOR U75 ( .A(n75), .B(n76), .Z(SUM[66]) );
  XNOR U76 ( .A(B[66]), .B(A[66]), .Z(n76) );
  XOR U77 ( .A(n77), .B(n78), .Z(SUM[65]) );
  XNOR U78 ( .A(B[65]), .B(A[65]), .Z(n78) );
  XOR U79 ( .A(n79), .B(n80), .Z(SUM[64]) );
  XNOR U80 ( .A(B[64]), .B(A[64]), .Z(n80) );
  XOR U81 ( .A(n81), .B(n82), .Z(SUM[63]) );
  XNOR U82 ( .A(B[63]), .B(A[63]), .Z(n82) );
  XOR U83 ( .A(n83), .B(n84), .Z(SUM[62]) );
  XNOR U84 ( .A(B[62]), .B(A[62]), .Z(n84) );
  XOR U85 ( .A(n85), .B(n86), .Z(SUM[61]) );
  XNOR U86 ( .A(B[61]), .B(A[61]), .Z(n86) );
  XOR U87 ( .A(n87), .B(n88), .Z(SUM[60]) );
  XNOR U88 ( .A(B[60]), .B(A[60]), .Z(n88) );
  XOR U89 ( .A(n89), .B(n90), .Z(SUM[5]) );
  XNOR U90 ( .A(B[5]), .B(A[5]), .Z(n90) );
  XOR U91 ( .A(n91), .B(n92), .Z(SUM[59]) );
  XNOR U92 ( .A(B[59]), .B(A[59]), .Z(n92) );
  XOR U93 ( .A(n93), .B(n94), .Z(SUM[58]) );
  XNOR U94 ( .A(B[58]), .B(A[58]), .Z(n94) );
  XOR U95 ( .A(n95), .B(n96), .Z(SUM[57]) );
  XNOR U96 ( .A(B[57]), .B(A[57]), .Z(n96) );
  XOR U97 ( .A(n97), .B(n98), .Z(SUM[56]) );
  XNOR U98 ( .A(B[56]), .B(A[56]), .Z(n98) );
  XOR U99 ( .A(n99), .B(n100), .Z(SUM[55]) );
  XNOR U100 ( .A(B[55]), .B(A[55]), .Z(n100) );
  XOR U101 ( .A(n101), .B(n102), .Z(SUM[54]) );
  XNOR U102 ( .A(B[54]), .B(A[54]), .Z(n102) );
  XOR U103 ( .A(n103), .B(n104), .Z(SUM[53]) );
  XNOR U104 ( .A(B[53]), .B(A[53]), .Z(n104) );
  XOR U105 ( .A(n105), .B(n106), .Z(SUM[52]) );
  XNOR U106 ( .A(B[52]), .B(A[52]), .Z(n106) );
  XOR U107 ( .A(n107), .B(n108), .Z(SUM[51]) );
  XNOR U108 ( .A(B[51]), .B(A[51]), .Z(n108) );
  XOR U109 ( .A(n109), .B(n110), .Z(SUM[50]) );
  XNOR U110 ( .A(B[50]), .B(A[50]), .Z(n110) );
  XOR U111 ( .A(n111), .B(n112), .Z(SUM[4]) );
  XNOR U112 ( .A(B[4]), .B(A[4]), .Z(n112) );
  XOR U113 ( .A(n113), .B(n114), .Z(SUM[49]) );
  XNOR U114 ( .A(B[49]), .B(A[49]), .Z(n114) );
  XOR U115 ( .A(n115), .B(n116), .Z(SUM[48]) );
  XNOR U116 ( .A(B[48]), .B(A[48]), .Z(n116) );
  XOR U117 ( .A(n117), .B(n118), .Z(SUM[47]) );
  XNOR U118 ( .A(B[47]), .B(A[47]), .Z(n118) );
  XOR U119 ( .A(n119), .B(n120), .Z(SUM[46]) );
  XNOR U120 ( .A(B[46]), .B(A[46]), .Z(n120) );
  XOR U121 ( .A(n121), .B(n122), .Z(SUM[45]) );
  XNOR U122 ( .A(B[45]), .B(A[45]), .Z(n122) );
  XOR U123 ( .A(n123), .B(n124), .Z(SUM[44]) );
  XNOR U124 ( .A(B[44]), .B(A[44]), .Z(n124) );
  XOR U125 ( .A(n125), .B(n126), .Z(SUM[43]) );
  XNOR U126 ( .A(B[43]), .B(A[43]), .Z(n126) );
  XOR U127 ( .A(n127), .B(n128), .Z(SUM[42]) );
  XNOR U128 ( .A(B[42]), .B(A[42]), .Z(n128) );
  XOR U129 ( .A(n129), .B(n130), .Z(SUM[41]) );
  XNOR U130 ( .A(B[41]), .B(A[41]), .Z(n130) );
  XOR U131 ( .A(n131), .B(n132), .Z(SUM[40]) );
  XNOR U132 ( .A(B[40]), .B(A[40]), .Z(n132) );
  XOR U133 ( .A(n133), .B(n134), .Z(SUM[3]) );
  XNOR U134 ( .A(B[3]), .B(A[3]), .Z(n134) );
  XOR U135 ( .A(n135), .B(n136), .Z(SUM[39]) );
  XNOR U136 ( .A(B[39]), .B(A[39]), .Z(n136) );
  XOR U137 ( .A(n137), .B(n138), .Z(SUM[38]) );
  XNOR U138 ( .A(B[38]), .B(A[38]), .Z(n138) );
  XOR U139 ( .A(n139), .B(n140), .Z(SUM[37]) );
  XNOR U140 ( .A(B[37]), .B(A[37]), .Z(n140) );
  XOR U141 ( .A(n141), .B(n142), .Z(SUM[36]) );
  XNOR U142 ( .A(B[36]), .B(A[36]), .Z(n142) );
  XOR U143 ( .A(n143), .B(n144), .Z(SUM[35]) );
  XNOR U144 ( .A(B[35]), .B(A[35]), .Z(n144) );
  XOR U145 ( .A(n145), .B(n146), .Z(SUM[34]) );
  XNOR U146 ( .A(B[34]), .B(A[34]), .Z(n146) );
  XOR U147 ( .A(n147), .B(n148), .Z(SUM[33]) );
  XNOR U148 ( .A(B[33]), .B(A[33]), .Z(n148) );
  XOR U149 ( .A(n149), .B(n150), .Z(SUM[32]) );
  XNOR U150 ( .A(B[32]), .B(A[32]), .Z(n150) );
  XOR U151 ( .A(n151), .B(n152), .Z(SUM[31]) );
  XNOR U152 ( .A(B[31]), .B(A[31]), .Z(n152) );
  XOR U153 ( .A(n153), .B(n154), .Z(SUM[30]) );
  XNOR U154 ( .A(B[30]), .B(A[30]), .Z(n154) );
  XOR U155 ( .A(n155), .B(n156), .Z(SUM[2]) );
  XOR U156 ( .A(B[2]), .B(A[2]), .Z(n156) );
  XOR U157 ( .A(n157), .B(n158), .Z(SUM[29]) );
  XNOR U158 ( .A(B[29]), .B(A[29]), .Z(n158) );
  XOR U159 ( .A(n159), .B(n160), .Z(SUM[28]) );
  XNOR U160 ( .A(B[28]), .B(A[28]), .Z(n160) );
  XOR U161 ( .A(n161), .B(n162), .Z(SUM[27]) );
  XNOR U162 ( .A(B[27]), .B(A[27]), .Z(n162) );
  XOR U163 ( .A(n163), .B(n164), .Z(SUM[26]) );
  XNOR U164 ( .A(B[26]), .B(A[26]), .Z(n164) );
  XOR U165 ( .A(n165), .B(n166), .Z(SUM[25]) );
  XNOR U166 ( .A(B[25]), .B(A[25]), .Z(n166) );
  XOR U167 ( .A(A[257]), .B(n167), .Z(SUM[257]) );
  AND U168 ( .A(A[256]), .B(n168), .Z(n167) );
  XOR U169 ( .A(A[256]), .B(n168), .Z(SUM[256]) );
  NAND U170 ( .A(n169), .B(n170), .Z(n168) );
  NAND U171 ( .A(B[255]), .B(n171), .Z(n170) );
  NANDN U172 ( .A(A[255]), .B(n172), .Z(n171) );
  NANDN U173 ( .A(n172), .B(A[255]), .Z(n169) );
  XOR U174 ( .A(n172), .B(n173), .Z(SUM[255]) );
  XNOR U175 ( .A(B[255]), .B(A[255]), .Z(n173) );
  AND U176 ( .A(n174), .B(n175), .Z(n172) );
  NAND U177 ( .A(B[254]), .B(n176), .Z(n175) );
  NANDN U178 ( .A(A[254]), .B(n177), .Z(n176) );
  NANDN U179 ( .A(n177), .B(A[254]), .Z(n174) );
  XOR U180 ( .A(n177), .B(n178), .Z(SUM[254]) );
  XNOR U181 ( .A(B[254]), .B(A[254]), .Z(n178) );
  AND U182 ( .A(n179), .B(n180), .Z(n177) );
  NAND U183 ( .A(B[253]), .B(n181), .Z(n180) );
  NANDN U184 ( .A(A[253]), .B(n182), .Z(n181) );
  NANDN U185 ( .A(n182), .B(A[253]), .Z(n179) );
  XOR U186 ( .A(n182), .B(n183), .Z(SUM[253]) );
  XNOR U187 ( .A(B[253]), .B(A[253]), .Z(n183) );
  AND U188 ( .A(n184), .B(n185), .Z(n182) );
  NAND U189 ( .A(B[252]), .B(n186), .Z(n185) );
  NANDN U190 ( .A(A[252]), .B(n187), .Z(n186) );
  NANDN U191 ( .A(n187), .B(A[252]), .Z(n184) );
  XOR U192 ( .A(n187), .B(n188), .Z(SUM[252]) );
  XNOR U193 ( .A(B[252]), .B(A[252]), .Z(n188) );
  AND U194 ( .A(n189), .B(n190), .Z(n187) );
  NAND U195 ( .A(B[251]), .B(n191), .Z(n190) );
  NANDN U196 ( .A(A[251]), .B(n192), .Z(n191) );
  NANDN U197 ( .A(n192), .B(A[251]), .Z(n189) );
  XOR U198 ( .A(n192), .B(n193), .Z(SUM[251]) );
  XNOR U199 ( .A(B[251]), .B(A[251]), .Z(n193) );
  AND U200 ( .A(n194), .B(n195), .Z(n192) );
  NAND U201 ( .A(B[250]), .B(n196), .Z(n195) );
  NANDN U202 ( .A(A[250]), .B(n197), .Z(n196) );
  NANDN U203 ( .A(n197), .B(A[250]), .Z(n194) );
  XOR U204 ( .A(n197), .B(n198), .Z(SUM[250]) );
  XNOR U205 ( .A(B[250]), .B(A[250]), .Z(n198) );
  AND U206 ( .A(n199), .B(n200), .Z(n197) );
  NAND U207 ( .A(B[249]), .B(n201), .Z(n200) );
  NANDN U208 ( .A(A[249]), .B(n202), .Z(n201) );
  NANDN U209 ( .A(n202), .B(A[249]), .Z(n199) );
  XOR U210 ( .A(n203), .B(n204), .Z(SUM[24]) );
  XNOR U211 ( .A(B[24]), .B(A[24]), .Z(n204) );
  XOR U212 ( .A(n202), .B(n205), .Z(SUM[249]) );
  XNOR U213 ( .A(B[249]), .B(A[249]), .Z(n205) );
  AND U214 ( .A(n206), .B(n207), .Z(n202) );
  NAND U215 ( .A(B[248]), .B(n208), .Z(n207) );
  NANDN U216 ( .A(A[248]), .B(n209), .Z(n208) );
  NANDN U217 ( .A(n209), .B(A[248]), .Z(n206) );
  XOR U218 ( .A(n209), .B(n210), .Z(SUM[248]) );
  XNOR U219 ( .A(B[248]), .B(A[248]), .Z(n210) );
  AND U220 ( .A(n211), .B(n212), .Z(n209) );
  NAND U221 ( .A(B[247]), .B(n213), .Z(n212) );
  NANDN U222 ( .A(A[247]), .B(n214), .Z(n213) );
  NANDN U223 ( .A(n214), .B(A[247]), .Z(n211) );
  XOR U224 ( .A(n214), .B(n215), .Z(SUM[247]) );
  XNOR U225 ( .A(B[247]), .B(A[247]), .Z(n215) );
  AND U226 ( .A(n216), .B(n217), .Z(n214) );
  NAND U227 ( .A(B[246]), .B(n218), .Z(n217) );
  NANDN U228 ( .A(A[246]), .B(n219), .Z(n218) );
  NANDN U229 ( .A(n219), .B(A[246]), .Z(n216) );
  XOR U230 ( .A(n219), .B(n220), .Z(SUM[246]) );
  XNOR U231 ( .A(B[246]), .B(A[246]), .Z(n220) );
  AND U232 ( .A(n221), .B(n222), .Z(n219) );
  NAND U233 ( .A(B[245]), .B(n223), .Z(n222) );
  NANDN U234 ( .A(A[245]), .B(n224), .Z(n223) );
  NANDN U235 ( .A(n224), .B(A[245]), .Z(n221) );
  XOR U236 ( .A(n224), .B(n225), .Z(SUM[245]) );
  XNOR U237 ( .A(B[245]), .B(A[245]), .Z(n225) );
  AND U238 ( .A(n226), .B(n227), .Z(n224) );
  NAND U239 ( .A(B[244]), .B(n228), .Z(n227) );
  NANDN U240 ( .A(A[244]), .B(n229), .Z(n228) );
  NANDN U241 ( .A(n229), .B(A[244]), .Z(n226) );
  XOR U242 ( .A(n229), .B(n230), .Z(SUM[244]) );
  XNOR U243 ( .A(B[244]), .B(A[244]), .Z(n230) );
  AND U244 ( .A(n231), .B(n232), .Z(n229) );
  NAND U245 ( .A(B[243]), .B(n233), .Z(n232) );
  NANDN U246 ( .A(A[243]), .B(n234), .Z(n233) );
  NANDN U247 ( .A(n234), .B(A[243]), .Z(n231) );
  XOR U248 ( .A(n234), .B(n235), .Z(SUM[243]) );
  XNOR U249 ( .A(B[243]), .B(A[243]), .Z(n235) );
  AND U250 ( .A(n236), .B(n237), .Z(n234) );
  NAND U251 ( .A(B[242]), .B(n238), .Z(n237) );
  NANDN U252 ( .A(A[242]), .B(n239), .Z(n238) );
  NANDN U253 ( .A(n239), .B(A[242]), .Z(n236) );
  XOR U254 ( .A(n239), .B(n240), .Z(SUM[242]) );
  XNOR U255 ( .A(B[242]), .B(A[242]), .Z(n240) );
  AND U256 ( .A(n241), .B(n242), .Z(n239) );
  NAND U257 ( .A(B[241]), .B(n243), .Z(n242) );
  NANDN U258 ( .A(A[241]), .B(n244), .Z(n243) );
  NANDN U259 ( .A(n244), .B(A[241]), .Z(n241) );
  XOR U260 ( .A(n244), .B(n245), .Z(SUM[241]) );
  XNOR U261 ( .A(B[241]), .B(A[241]), .Z(n245) );
  AND U262 ( .A(n246), .B(n247), .Z(n244) );
  NAND U263 ( .A(B[240]), .B(n248), .Z(n247) );
  NANDN U264 ( .A(A[240]), .B(n249), .Z(n248) );
  NANDN U265 ( .A(n249), .B(A[240]), .Z(n246) );
  XOR U266 ( .A(n249), .B(n250), .Z(SUM[240]) );
  XNOR U267 ( .A(B[240]), .B(A[240]), .Z(n250) );
  AND U268 ( .A(n251), .B(n252), .Z(n249) );
  NAND U269 ( .A(B[239]), .B(n253), .Z(n252) );
  NANDN U270 ( .A(A[239]), .B(n254), .Z(n253) );
  NANDN U271 ( .A(n254), .B(A[239]), .Z(n251) );
  XOR U272 ( .A(n255), .B(n256), .Z(SUM[23]) );
  XNOR U273 ( .A(B[23]), .B(A[23]), .Z(n256) );
  XOR U274 ( .A(n254), .B(n257), .Z(SUM[239]) );
  XNOR U275 ( .A(B[239]), .B(A[239]), .Z(n257) );
  AND U276 ( .A(n258), .B(n259), .Z(n254) );
  NAND U277 ( .A(B[238]), .B(n260), .Z(n259) );
  NANDN U278 ( .A(A[238]), .B(n261), .Z(n260) );
  NANDN U279 ( .A(n261), .B(A[238]), .Z(n258) );
  XOR U280 ( .A(n261), .B(n262), .Z(SUM[238]) );
  XNOR U281 ( .A(B[238]), .B(A[238]), .Z(n262) );
  AND U282 ( .A(n263), .B(n264), .Z(n261) );
  NAND U283 ( .A(B[237]), .B(n265), .Z(n264) );
  NANDN U284 ( .A(A[237]), .B(n266), .Z(n265) );
  NANDN U285 ( .A(n266), .B(A[237]), .Z(n263) );
  XOR U286 ( .A(n266), .B(n267), .Z(SUM[237]) );
  XNOR U287 ( .A(B[237]), .B(A[237]), .Z(n267) );
  AND U288 ( .A(n268), .B(n269), .Z(n266) );
  NAND U289 ( .A(B[236]), .B(n270), .Z(n269) );
  NANDN U290 ( .A(A[236]), .B(n271), .Z(n270) );
  NANDN U291 ( .A(n271), .B(A[236]), .Z(n268) );
  XOR U292 ( .A(n271), .B(n272), .Z(SUM[236]) );
  XNOR U293 ( .A(B[236]), .B(A[236]), .Z(n272) );
  AND U294 ( .A(n273), .B(n274), .Z(n271) );
  NAND U295 ( .A(B[235]), .B(n275), .Z(n274) );
  NANDN U296 ( .A(A[235]), .B(n276), .Z(n275) );
  NANDN U297 ( .A(n276), .B(A[235]), .Z(n273) );
  XOR U298 ( .A(n276), .B(n277), .Z(SUM[235]) );
  XNOR U299 ( .A(B[235]), .B(A[235]), .Z(n277) );
  AND U300 ( .A(n278), .B(n279), .Z(n276) );
  NAND U301 ( .A(B[234]), .B(n280), .Z(n279) );
  NANDN U302 ( .A(A[234]), .B(n281), .Z(n280) );
  NANDN U303 ( .A(n281), .B(A[234]), .Z(n278) );
  XOR U304 ( .A(n281), .B(n282), .Z(SUM[234]) );
  XNOR U305 ( .A(B[234]), .B(A[234]), .Z(n282) );
  AND U306 ( .A(n283), .B(n284), .Z(n281) );
  NAND U307 ( .A(B[233]), .B(n285), .Z(n284) );
  NANDN U308 ( .A(A[233]), .B(n286), .Z(n285) );
  NANDN U309 ( .A(n286), .B(A[233]), .Z(n283) );
  XOR U310 ( .A(n286), .B(n287), .Z(SUM[233]) );
  XNOR U311 ( .A(B[233]), .B(A[233]), .Z(n287) );
  AND U312 ( .A(n288), .B(n289), .Z(n286) );
  NAND U313 ( .A(B[232]), .B(n290), .Z(n289) );
  NANDN U314 ( .A(A[232]), .B(n291), .Z(n290) );
  NANDN U315 ( .A(n291), .B(A[232]), .Z(n288) );
  XOR U316 ( .A(n291), .B(n292), .Z(SUM[232]) );
  XNOR U317 ( .A(B[232]), .B(A[232]), .Z(n292) );
  AND U318 ( .A(n293), .B(n294), .Z(n291) );
  NAND U319 ( .A(B[231]), .B(n295), .Z(n294) );
  NANDN U320 ( .A(A[231]), .B(n296), .Z(n295) );
  NANDN U321 ( .A(n296), .B(A[231]), .Z(n293) );
  XOR U322 ( .A(n296), .B(n297), .Z(SUM[231]) );
  XNOR U323 ( .A(B[231]), .B(A[231]), .Z(n297) );
  AND U324 ( .A(n298), .B(n299), .Z(n296) );
  NAND U325 ( .A(B[230]), .B(n300), .Z(n299) );
  NANDN U326 ( .A(A[230]), .B(n301), .Z(n300) );
  NANDN U327 ( .A(n301), .B(A[230]), .Z(n298) );
  XOR U328 ( .A(n301), .B(n302), .Z(SUM[230]) );
  XNOR U329 ( .A(B[230]), .B(A[230]), .Z(n302) );
  AND U330 ( .A(n303), .B(n304), .Z(n301) );
  NAND U331 ( .A(B[229]), .B(n305), .Z(n304) );
  NANDN U332 ( .A(A[229]), .B(n306), .Z(n305) );
  NANDN U333 ( .A(n306), .B(A[229]), .Z(n303) );
  XOR U334 ( .A(n307), .B(n308), .Z(SUM[22]) );
  XNOR U335 ( .A(B[22]), .B(A[22]), .Z(n308) );
  XOR U336 ( .A(n306), .B(n309), .Z(SUM[229]) );
  XNOR U337 ( .A(B[229]), .B(A[229]), .Z(n309) );
  AND U338 ( .A(n310), .B(n311), .Z(n306) );
  NAND U339 ( .A(B[228]), .B(n312), .Z(n311) );
  NANDN U340 ( .A(A[228]), .B(n313), .Z(n312) );
  NANDN U341 ( .A(n313), .B(A[228]), .Z(n310) );
  XOR U342 ( .A(n313), .B(n314), .Z(SUM[228]) );
  XNOR U343 ( .A(B[228]), .B(A[228]), .Z(n314) );
  AND U344 ( .A(n315), .B(n316), .Z(n313) );
  NAND U345 ( .A(B[227]), .B(n317), .Z(n316) );
  NANDN U346 ( .A(A[227]), .B(n318), .Z(n317) );
  NANDN U347 ( .A(n318), .B(A[227]), .Z(n315) );
  XOR U348 ( .A(n318), .B(n319), .Z(SUM[227]) );
  XNOR U349 ( .A(B[227]), .B(A[227]), .Z(n319) );
  AND U350 ( .A(n320), .B(n321), .Z(n318) );
  NAND U351 ( .A(B[226]), .B(n322), .Z(n321) );
  NANDN U352 ( .A(A[226]), .B(n323), .Z(n322) );
  NANDN U353 ( .A(n323), .B(A[226]), .Z(n320) );
  XOR U354 ( .A(n323), .B(n324), .Z(SUM[226]) );
  XNOR U355 ( .A(B[226]), .B(A[226]), .Z(n324) );
  AND U356 ( .A(n325), .B(n326), .Z(n323) );
  NAND U357 ( .A(B[225]), .B(n327), .Z(n326) );
  NANDN U358 ( .A(A[225]), .B(n328), .Z(n327) );
  NANDN U359 ( .A(n328), .B(A[225]), .Z(n325) );
  XOR U360 ( .A(n328), .B(n329), .Z(SUM[225]) );
  XNOR U361 ( .A(B[225]), .B(A[225]), .Z(n329) );
  AND U362 ( .A(n330), .B(n331), .Z(n328) );
  NAND U363 ( .A(B[224]), .B(n332), .Z(n331) );
  NANDN U364 ( .A(A[224]), .B(n333), .Z(n332) );
  NANDN U365 ( .A(n333), .B(A[224]), .Z(n330) );
  XOR U366 ( .A(n333), .B(n334), .Z(SUM[224]) );
  XNOR U367 ( .A(B[224]), .B(A[224]), .Z(n334) );
  AND U368 ( .A(n335), .B(n336), .Z(n333) );
  NAND U369 ( .A(B[223]), .B(n337), .Z(n336) );
  NANDN U370 ( .A(A[223]), .B(n338), .Z(n337) );
  NANDN U371 ( .A(n338), .B(A[223]), .Z(n335) );
  XOR U372 ( .A(n338), .B(n339), .Z(SUM[223]) );
  XNOR U373 ( .A(B[223]), .B(A[223]), .Z(n339) );
  AND U374 ( .A(n340), .B(n341), .Z(n338) );
  NAND U375 ( .A(B[222]), .B(n342), .Z(n341) );
  NANDN U376 ( .A(A[222]), .B(n343), .Z(n342) );
  NANDN U377 ( .A(n343), .B(A[222]), .Z(n340) );
  XOR U378 ( .A(n343), .B(n344), .Z(SUM[222]) );
  XNOR U379 ( .A(B[222]), .B(A[222]), .Z(n344) );
  AND U380 ( .A(n345), .B(n346), .Z(n343) );
  NAND U381 ( .A(B[221]), .B(n347), .Z(n346) );
  NANDN U382 ( .A(A[221]), .B(n348), .Z(n347) );
  NANDN U383 ( .A(n348), .B(A[221]), .Z(n345) );
  XOR U384 ( .A(n348), .B(n349), .Z(SUM[221]) );
  XNOR U385 ( .A(B[221]), .B(A[221]), .Z(n349) );
  AND U386 ( .A(n350), .B(n351), .Z(n348) );
  NAND U387 ( .A(B[220]), .B(n352), .Z(n351) );
  NANDN U388 ( .A(A[220]), .B(n353), .Z(n352) );
  NANDN U389 ( .A(n353), .B(A[220]), .Z(n350) );
  XOR U390 ( .A(n353), .B(n354), .Z(SUM[220]) );
  XNOR U391 ( .A(B[220]), .B(A[220]), .Z(n354) );
  AND U392 ( .A(n355), .B(n356), .Z(n353) );
  NAND U393 ( .A(B[219]), .B(n357), .Z(n356) );
  NANDN U394 ( .A(A[219]), .B(n358), .Z(n357) );
  NANDN U395 ( .A(n358), .B(A[219]), .Z(n355) );
  XOR U396 ( .A(n359), .B(n360), .Z(SUM[21]) );
  XNOR U397 ( .A(B[21]), .B(A[21]), .Z(n360) );
  XOR U398 ( .A(n358), .B(n361), .Z(SUM[219]) );
  XNOR U399 ( .A(B[219]), .B(A[219]), .Z(n361) );
  AND U400 ( .A(n362), .B(n363), .Z(n358) );
  NAND U401 ( .A(B[218]), .B(n364), .Z(n363) );
  NANDN U402 ( .A(A[218]), .B(n365), .Z(n364) );
  NANDN U403 ( .A(n365), .B(A[218]), .Z(n362) );
  XOR U404 ( .A(n365), .B(n366), .Z(SUM[218]) );
  XNOR U405 ( .A(B[218]), .B(A[218]), .Z(n366) );
  AND U406 ( .A(n367), .B(n368), .Z(n365) );
  NAND U407 ( .A(B[217]), .B(n369), .Z(n368) );
  NANDN U408 ( .A(A[217]), .B(n370), .Z(n369) );
  NANDN U409 ( .A(n370), .B(A[217]), .Z(n367) );
  XOR U410 ( .A(n370), .B(n371), .Z(SUM[217]) );
  XNOR U411 ( .A(B[217]), .B(A[217]), .Z(n371) );
  AND U412 ( .A(n372), .B(n373), .Z(n370) );
  NAND U413 ( .A(B[216]), .B(n374), .Z(n373) );
  NANDN U414 ( .A(A[216]), .B(n375), .Z(n374) );
  NANDN U415 ( .A(n375), .B(A[216]), .Z(n372) );
  XOR U416 ( .A(n375), .B(n376), .Z(SUM[216]) );
  XNOR U417 ( .A(B[216]), .B(A[216]), .Z(n376) );
  AND U418 ( .A(n377), .B(n378), .Z(n375) );
  NAND U419 ( .A(B[215]), .B(n379), .Z(n378) );
  NANDN U420 ( .A(A[215]), .B(n380), .Z(n379) );
  NANDN U421 ( .A(n380), .B(A[215]), .Z(n377) );
  XOR U422 ( .A(n380), .B(n381), .Z(SUM[215]) );
  XNOR U423 ( .A(B[215]), .B(A[215]), .Z(n381) );
  AND U424 ( .A(n382), .B(n383), .Z(n380) );
  NAND U425 ( .A(B[214]), .B(n384), .Z(n383) );
  NANDN U426 ( .A(A[214]), .B(n385), .Z(n384) );
  NANDN U427 ( .A(n385), .B(A[214]), .Z(n382) );
  XOR U428 ( .A(n385), .B(n386), .Z(SUM[214]) );
  XNOR U429 ( .A(B[214]), .B(A[214]), .Z(n386) );
  AND U430 ( .A(n387), .B(n388), .Z(n385) );
  NAND U431 ( .A(B[213]), .B(n389), .Z(n388) );
  NANDN U432 ( .A(A[213]), .B(n390), .Z(n389) );
  NANDN U433 ( .A(n390), .B(A[213]), .Z(n387) );
  XOR U434 ( .A(n390), .B(n391), .Z(SUM[213]) );
  XNOR U435 ( .A(B[213]), .B(A[213]), .Z(n391) );
  AND U436 ( .A(n392), .B(n393), .Z(n390) );
  NAND U437 ( .A(B[212]), .B(n394), .Z(n393) );
  NANDN U438 ( .A(A[212]), .B(n395), .Z(n394) );
  NANDN U439 ( .A(n395), .B(A[212]), .Z(n392) );
  XOR U440 ( .A(n395), .B(n396), .Z(SUM[212]) );
  XNOR U441 ( .A(B[212]), .B(A[212]), .Z(n396) );
  AND U442 ( .A(n397), .B(n398), .Z(n395) );
  NAND U443 ( .A(B[211]), .B(n399), .Z(n398) );
  NANDN U444 ( .A(A[211]), .B(n400), .Z(n399) );
  NANDN U445 ( .A(n400), .B(A[211]), .Z(n397) );
  XOR U446 ( .A(n400), .B(n401), .Z(SUM[211]) );
  XNOR U447 ( .A(B[211]), .B(A[211]), .Z(n401) );
  AND U448 ( .A(n402), .B(n403), .Z(n400) );
  NAND U449 ( .A(B[210]), .B(n404), .Z(n403) );
  NANDN U450 ( .A(A[210]), .B(n405), .Z(n404) );
  NANDN U451 ( .A(n405), .B(A[210]), .Z(n402) );
  XOR U452 ( .A(n405), .B(n406), .Z(SUM[210]) );
  XNOR U453 ( .A(B[210]), .B(A[210]), .Z(n406) );
  AND U454 ( .A(n407), .B(n408), .Z(n405) );
  NAND U455 ( .A(B[209]), .B(n409), .Z(n408) );
  NANDN U456 ( .A(A[209]), .B(n410), .Z(n409) );
  NANDN U457 ( .A(n410), .B(A[209]), .Z(n407) );
  XOR U458 ( .A(n411), .B(n412), .Z(SUM[20]) );
  XNOR U459 ( .A(B[20]), .B(A[20]), .Z(n412) );
  XOR U460 ( .A(n410), .B(n413), .Z(SUM[209]) );
  XNOR U461 ( .A(B[209]), .B(A[209]), .Z(n413) );
  AND U462 ( .A(n414), .B(n415), .Z(n410) );
  NAND U463 ( .A(B[208]), .B(n416), .Z(n415) );
  NANDN U464 ( .A(A[208]), .B(n417), .Z(n416) );
  NANDN U465 ( .A(n417), .B(A[208]), .Z(n414) );
  XOR U466 ( .A(n417), .B(n418), .Z(SUM[208]) );
  XNOR U467 ( .A(B[208]), .B(A[208]), .Z(n418) );
  AND U468 ( .A(n419), .B(n420), .Z(n417) );
  NAND U469 ( .A(B[207]), .B(n421), .Z(n420) );
  NANDN U470 ( .A(A[207]), .B(n422), .Z(n421) );
  NANDN U471 ( .A(n422), .B(A[207]), .Z(n419) );
  XOR U472 ( .A(n422), .B(n423), .Z(SUM[207]) );
  XNOR U473 ( .A(B[207]), .B(A[207]), .Z(n423) );
  AND U474 ( .A(n424), .B(n425), .Z(n422) );
  NAND U475 ( .A(B[206]), .B(n426), .Z(n425) );
  NANDN U476 ( .A(A[206]), .B(n427), .Z(n426) );
  NANDN U477 ( .A(n427), .B(A[206]), .Z(n424) );
  XOR U478 ( .A(n427), .B(n428), .Z(SUM[206]) );
  XNOR U479 ( .A(B[206]), .B(A[206]), .Z(n428) );
  AND U480 ( .A(n429), .B(n430), .Z(n427) );
  NAND U481 ( .A(B[205]), .B(n431), .Z(n430) );
  NANDN U482 ( .A(A[205]), .B(n432), .Z(n431) );
  NANDN U483 ( .A(n432), .B(A[205]), .Z(n429) );
  XOR U484 ( .A(n432), .B(n433), .Z(SUM[205]) );
  XNOR U485 ( .A(B[205]), .B(A[205]), .Z(n433) );
  AND U486 ( .A(n434), .B(n435), .Z(n432) );
  NAND U487 ( .A(B[204]), .B(n436), .Z(n435) );
  NANDN U488 ( .A(A[204]), .B(n437), .Z(n436) );
  NANDN U489 ( .A(n437), .B(A[204]), .Z(n434) );
  XOR U490 ( .A(n437), .B(n438), .Z(SUM[204]) );
  XNOR U491 ( .A(B[204]), .B(A[204]), .Z(n438) );
  AND U492 ( .A(n439), .B(n440), .Z(n437) );
  NAND U493 ( .A(B[203]), .B(n441), .Z(n440) );
  NANDN U494 ( .A(A[203]), .B(n442), .Z(n441) );
  NANDN U495 ( .A(n442), .B(A[203]), .Z(n439) );
  XOR U496 ( .A(n442), .B(n443), .Z(SUM[203]) );
  XNOR U497 ( .A(B[203]), .B(A[203]), .Z(n443) );
  AND U498 ( .A(n444), .B(n445), .Z(n442) );
  NAND U499 ( .A(B[202]), .B(n446), .Z(n445) );
  NANDN U500 ( .A(A[202]), .B(n447), .Z(n446) );
  NANDN U501 ( .A(n447), .B(A[202]), .Z(n444) );
  XOR U502 ( .A(n447), .B(n448), .Z(SUM[202]) );
  XNOR U503 ( .A(B[202]), .B(A[202]), .Z(n448) );
  AND U504 ( .A(n449), .B(n450), .Z(n447) );
  NAND U505 ( .A(B[201]), .B(n451), .Z(n450) );
  NANDN U506 ( .A(A[201]), .B(n452), .Z(n451) );
  NANDN U507 ( .A(n452), .B(A[201]), .Z(n449) );
  XOR U508 ( .A(n452), .B(n453), .Z(SUM[201]) );
  XNOR U509 ( .A(B[201]), .B(A[201]), .Z(n453) );
  AND U510 ( .A(n454), .B(n455), .Z(n452) );
  NAND U511 ( .A(B[200]), .B(n456), .Z(n455) );
  NANDN U512 ( .A(A[200]), .B(n457), .Z(n456) );
  NANDN U513 ( .A(n457), .B(A[200]), .Z(n454) );
  XOR U514 ( .A(n457), .B(n458), .Z(SUM[200]) );
  XNOR U515 ( .A(B[200]), .B(A[200]), .Z(n458) );
  AND U516 ( .A(n459), .B(n460), .Z(n457) );
  NAND U517 ( .A(B[199]), .B(n461), .Z(n460) );
  NANDN U518 ( .A(A[199]), .B(n462), .Z(n461) );
  NANDN U519 ( .A(n462), .B(A[199]), .Z(n459) );
  XOR U520 ( .A(B[1]), .B(A[1]), .Z(SUM[1]) );
  XOR U521 ( .A(n463), .B(n464), .Z(SUM[19]) );
  XNOR U522 ( .A(B[19]), .B(A[19]), .Z(n464) );
  XOR U523 ( .A(n462), .B(n465), .Z(SUM[199]) );
  XNOR U524 ( .A(B[199]), .B(A[199]), .Z(n465) );
  AND U525 ( .A(n466), .B(n467), .Z(n462) );
  NAND U526 ( .A(B[198]), .B(n468), .Z(n467) );
  NANDN U527 ( .A(A[198]), .B(n469), .Z(n468) );
  NANDN U528 ( .A(n469), .B(A[198]), .Z(n466) );
  XOR U529 ( .A(n469), .B(n470), .Z(SUM[198]) );
  XNOR U530 ( .A(B[198]), .B(A[198]), .Z(n470) );
  AND U531 ( .A(n471), .B(n472), .Z(n469) );
  NAND U532 ( .A(B[197]), .B(n473), .Z(n472) );
  NANDN U533 ( .A(A[197]), .B(n474), .Z(n473) );
  NANDN U534 ( .A(n474), .B(A[197]), .Z(n471) );
  XOR U535 ( .A(n474), .B(n475), .Z(SUM[197]) );
  XNOR U536 ( .A(B[197]), .B(A[197]), .Z(n475) );
  AND U537 ( .A(n476), .B(n477), .Z(n474) );
  NAND U538 ( .A(B[196]), .B(n478), .Z(n477) );
  NANDN U539 ( .A(A[196]), .B(n479), .Z(n478) );
  NANDN U540 ( .A(n479), .B(A[196]), .Z(n476) );
  XOR U541 ( .A(n479), .B(n480), .Z(SUM[196]) );
  XNOR U542 ( .A(B[196]), .B(A[196]), .Z(n480) );
  AND U543 ( .A(n481), .B(n482), .Z(n479) );
  NAND U544 ( .A(B[195]), .B(n483), .Z(n482) );
  NANDN U545 ( .A(A[195]), .B(n484), .Z(n483) );
  NANDN U546 ( .A(n484), .B(A[195]), .Z(n481) );
  XOR U547 ( .A(n484), .B(n485), .Z(SUM[195]) );
  XNOR U548 ( .A(B[195]), .B(A[195]), .Z(n485) );
  AND U549 ( .A(n486), .B(n487), .Z(n484) );
  NAND U550 ( .A(B[194]), .B(n488), .Z(n487) );
  NANDN U551 ( .A(A[194]), .B(n489), .Z(n488) );
  NANDN U552 ( .A(n489), .B(A[194]), .Z(n486) );
  XOR U553 ( .A(n489), .B(n490), .Z(SUM[194]) );
  XNOR U554 ( .A(B[194]), .B(A[194]), .Z(n490) );
  AND U555 ( .A(n491), .B(n492), .Z(n489) );
  NAND U556 ( .A(B[193]), .B(n493), .Z(n492) );
  NANDN U557 ( .A(A[193]), .B(n494), .Z(n493) );
  NANDN U558 ( .A(n494), .B(A[193]), .Z(n491) );
  XOR U559 ( .A(n494), .B(n495), .Z(SUM[193]) );
  XNOR U560 ( .A(B[193]), .B(A[193]), .Z(n495) );
  AND U561 ( .A(n496), .B(n497), .Z(n494) );
  NAND U562 ( .A(B[192]), .B(n498), .Z(n497) );
  NANDN U563 ( .A(A[192]), .B(n499), .Z(n498) );
  NANDN U564 ( .A(n499), .B(A[192]), .Z(n496) );
  XOR U565 ( .A(n499), .B(n500), .Z(SUM[192]) );
  XNOR U566 ( .A(B[192]), .B(A[192]), .Z(n500) );
  AND U567 ( .A(n501), .B(n502), .Z(n499) );
  NAND U568 ( .A(B[191]), .B(n503), .Z(n502) );
  NANDN U569 ( .A(A[191]), .B(n504), .Z(n503) );
  NANDN U570 ( .A(n504), .B(A[191]), .Z(n501) );
  XOR U571 ( .A(n504), .B(n505), .Z(SUM[191]) );
  XNOR U572 ( .A(B[191]), .B(A[191]), .Z(n505) );
  AND U573 ( .A(n506), .B(n507), .Z(n504) );
  NAND U574 ( .A(B[190]), .B(n508), .Z(n507) );
  NANDN U575 ( .A(A[190]), .B(n509), .Z(n508) );
  NANDN U576 ( .A(n509), .B(A[190]), .Z(n506) );
  XOR U577 ( .A(n509), .B(n510), .Z(SUM[190]) );
  XNOR U578 ( .A(B[190]), .B(A[190]), .Z(n510) );
  AND U579 ( .A(n511), .B(n512), .Z(n509) );
  NAND U580 ( .A(B[189]), .B(n513), .Z(n512) );
  NANDN U581 ( .A(A[189]), .B(n514), .Z(n513) );
  NANDN U582 ( .A(n514), .B(A[189]), .Z(n511) );
  XOR U583 ( .A(n515), .B(n516), .Z(SUM[18]) );
  XNOR U584 ( .A(B[18]), .B(A[18]), .Z(n516) );
  XOR U585 ( .A(n514), .B(n517), .Z(SUM[189]) );
  XNOR U586 ( .A(B[189]), .B(A[189]), .Z(n517) );
  AND U587 ( .A(n518), .B(n519), .Z(n514) );
  NAND U588 ( .A(B[188]), .B(n520), .Z(n519) );
  NANDN U589 ( .A(A[188]), .B(n521), .Z(n520) );
  NANDN U590 ( .A(n521), .B(A[188]), .Z(n518) );
  XOR U591 ( .A(n521), .B(n522), .Z(SUM[188]) );
  XNOR U592 ( .A(B[188]), .B(A[188]), .Z(n522) );
  AND U593 ( .A(n523), .B(n524), .Z(n521) );
  NAND U594 ( .A(B[187]), .B(n525), .Z(n524) );
  NANDN U595 ( .A(A[187]), .B(n526), .Z(n525) );
  NANDN U596 ( .A(n526), .B(A[187]), .Z(n523) );
  XOR U597 ( .A(n526), .B(n527), .Z(SUM[187]) );
  XNOR U598 ( .A(B[187]), .B(A[187]), .Z(n527) );
  AND U599 ( .A(n528), .B(n529), .Z(n526) );
  NAND U600 ( .A(B[186]), .B(n530), .Z(n529) );
  NANDN U601 ( .A(A[186]), .B(n531), .Z(n530) );
  NANDN U602 ( .A(n531), .B(A[186]), .Z(n528) );
  XOR U603 ( .A(n531), .B(n532), .Z(SUM[186]) );
  XNOR U604 ( .A(B[186]), .B(A[186]), .Z(n532) );
  AND U605 ( .A(n533), .B(n534), .Z(n531) );
  NAND U606 ( .A(B[185]), .B(n535), .Z(n534) );
  NANDN U607 ( .A(A[185]), .B(n536), .Z(n535) );
  NANDN U608 ( .A(n536), .B(A[185]), .Z(n533) );
  XOR U609 ( .A(n536), .B(n537), .Z(SUM[185]) );
  XNOR U610 ( .A(B[185]), .B(A[185]), .Z(n537) );
  AND U611 ( .A(n538), .B(n539), .Z(n536) );
  NAND U612 ( .A(B[184]), .B(n540), .Z(n539) );
  NANDN U613 ( .A(A[184]), .B(n541), .Z(n540) );
  NANDN U614 ( .A(n541), .B(A[184]), .Z(n538) );
  XOR U615 ( .A(n541), .B(n542), .Z(SUM[184]) );
  XNOR U616 ( .A(B[184]), .B(A[184]), .Z(n542) );
  AND U617 ( .A(n543), .B(n544), .Z(n541) );
  NAND U618 ( .A(B[183]), .B(n545), .Z(n544) );
  NANDN U619 ( .A(A[183]), .B(n546), .Z(n545) );
  NANDN U620 ( .A(n546), .B(A[183]), .Z(n543) );
  XOR U621 ( .A(n546), .B(n547), .Z(SUM[183]) );
  XNOR U622 ( .A(B[183]), .B(A[183]), .Z(n547) );
  AND U623 ( .A(n548), .B(n549), .Z(n546) );
  NAND U624 ( .A(B[182]), .B(n550), .Z(n549) );
  NANDN U625 ( .A(A[182]), .B(n551), .Z(n550) );
  NANDN U626 ( .A(n551), .B(A[182]), .Z(n548) );
  XOR U627 ( .A(n551), .B(n552), .Z(SUM[182]) );
  XNOR U628 ( .A(B[182]), .B(A[182]), .Z(n552) );
  AND U629 ( .A(n553), .B(n554), .Z(n551) );
  NAND U630 ( .A(B[181]), .B(n555), .Z(n554) );
  NANDN U631 ( .A(A[181]), .B(n556), .Z(n555) );
  NANDN U632 ( .A(n556), .B(A[181]), .Z(n553) );
  XOR U633 ( .A(n556), .B(n557), .Z(SUM[181]) );
  XNOR U634 ( .A(B[181]), .B(A[181]), .Z(n557) );
  AND U635 ( .A(n558), .B(n559), .Z(n556) );
  NAND U636 ( .A(B[180]), .B(n560), .Z(n559) );
  NANDN U637 ( .A(A[180]), .B(n561), .Z(n560) );
  NANDN U638 ( .A(n561), .B(A[180]), .Z(n558) );
  XOR U639 ( .A(n561), .B(n562), .Z(SUM[180]) );
  XNOR U640 ( .A(B[180]), .B(A[180]), .Z(n562) );
  AND U641 ( .A(n563), .B(n564), .Z(n561) );
  NAND U642 ( .A(B[179]), .B(n565), .Z(n564) );
  NANDN U643 ( .A(A[179]), .B(n566), .Z(n565) );
  NANDN U644 ( .A(n566), .B(A[179]), .Z(n563) );
  XOR U645 ( .A(n567), .B(n568), .Z(SUM[17]) );
  XNOR U646 ( .A(B[17]), .B(A[17]), .Z(n568) );
  XOR U647 ( .A(n566), .B(n569), .Z(SUM[179]) );
  XNOR U648 ( .A(B[179]), .B(A[179]), .Z(n569) );
  AND U649 ( .A(n570), .B(n571), .Z(n566) );
  NAND U650 ( .A(B[178]), .B(n572), .Z(n571) );
  NANDN U651 ( .A(A[178]), .B(n573), .Z(n572) );
  NANDN U652 ( .A(n573), .B(A[178]), .Z(n570) );
  XOR U653 ( .A(n573), .B(n574), .Z(SUM[178]) );
  XNOR U654 ( .A(B[178]), .B(A[178]), .Z(n574) );
  AND U655 ( .A(n575), .B(n576), .Z(n573) );
  NAND U656 ( .A(B[177]), .B(n577), .Z(n576) );
  NANDN U657 ( .A(A[177]), .B(n578), .Z(n577) );
  NANDN U658 ( .A(n578), .B(A[177]), .Z(n575) );
  XOR U659 ( .A(n578), .B(n579), .Z(SUM[177]) );
  XNOR U660 ( .A(B[177]), .B(A[177]), .Z(n579) );
  AND U661 ( .A(n580), .B(n581), .Z(n578) );
  NAND U662 ( .A(B[176]), .B(n582), .Z(n581) );
  NANDN U663 ( .A(A[176]), .B(n583), .Z(n582) );
  NANDN U664 ( .A(n583), .B(A[176]), .Z(n580) );
  XOR U665 ( .A(n583), .B(n584), .Z(SUM[176]) );
  XNOR U666 ( .A(B[176]), .B(A[176]), .Z(n584) );
  AND U667 ( .A(n585), .B(n586), .Z(n583) );
  NAND U668 ( .A(B[175]), .B(n587), .Z(n586) );
  NANDN U669 ( .A(A[175]), .B(n588), .Z(n587) );
  NANDN U670 ( .A(n588), .B(A[175]), .Z(n585) );
  XOR U671 ( .A(n588), .B(n589), .Z(SUM[175]) );
  XNOR U672 ( .A(B[175]), .B(A[175]), .Z(n589) );
  AND U673 ( .A(n590), .B(n591), .Z(n588) );
  NAND U674 ( .A(B[174]), .B(n592), .Z(n591) );
  NANDN U675 ( .A(A[174]), .B(n593), .Z(n592) );
  NANDN U676 ( .A(n593), .B(A[174]), .Z(n590) );
  XOR U677 ( .A(n593), .B(n594), .Z(SUM[174]) );
  XNOR U678 ( .A(B[174]), .B(A[174]), .Z(n594) );
  AND U679 ( .A(n595), .B(n596), .Z(n593) );
  NAND U680 ( .A(B[173]), .B(n597), .Z(n596) );
  NANDN U681 ( .A(A[173]), .B(n598), .Z(n597) );
  NANDN U682 ( .A(n598), .B(A[173]), .Z(n595) );
  XOR U683 ( .A(n598), .B(n599), .Z(SUM[173]) );
  XNOR U684 ( .A(B[173]), .B(A[173]), .Z(n599) );
  AND U685 ( .A(n600), .B(n601), .Z(n598) );
  NAND U686 ( .A(B[172]), .B(n602), .Z(n601) );
  NANDN U687 ( .A(A[172]), .B(n603), .Z(n602) );
  NANDN U688 ( .A(n603), .B(A[172]), .Z(n600) );
  XOR U689 ( .A(n603), .B(n604), .Z(SUM[172]) );
  XNOR U690 ( .A(B[172]), .B(A[172]), .Z(n604) );
  AND U691 ( .A(n605), .B(n606), .Z(n603) );
  NAND U692 ( .A(B[171]), .B(n607), .Z(n606) );
  NANDN U693 ( .A(A[171]), .B(n608), .Z(n607) );
  NANDN U694 ( .A(n608), .B(A[171]), .Z(n605) );
  XOR U695 ( .A(n608), .B(n609), .Z(SUM[171]) );
  XNOR U696 ( .A(B[171]), .B(A[171]), .Z(n609) );
  AND U697 ( .A(n610), .B(n611), .Z(n608) );
  NAND U698 ( .A(B[170]), .B(n612), .Z(n611) );
  NANDN U699 ( .A(A[170]), .B(n613), .Z(n612) );
  NANDN U700 ( .A(n613), .B(A[170]), .Z(n610) );
  XOR U701 ( .A(n613), .B(n614), .Z(SUM[170]) );
  XNOR U702 ( .A(B[170]), .B(A[170]), .Z(n614) );
  AND U703 ( .A(n615), .B(n616), .Z(n613) );
  NAND U704 ( .A(B[169]), .B(n617), .Z(n616) );
  NANDN U705 ( .A(A[169]), .B(n618), .Z(n617) );
  NANDN U706 ( .A(n618), .B(A[169]), .Z(n615) );
  XOR U707 ( .A(n619), .B(n620), .Z(SUM[16]) );
  XNOR U708 ( .A(B[16]), .B(A[16]), .Z(n620) );
  XOR U709 ( .A(n618), .B(n621), .Z(SUM[169]) );
  XNOR U710 ( .A(B[169]), .B(A[169]), .Z(n621) );
  AND U711 ( .A(n622), .B(n623), .Z(n618) );
  NAND U712 ( .A(B[168]), .B(n624), .Z(n623) );
  NANDN U713 ( .A(A[168]), .B(n625), .Z(n624) );
  NANDN U714 ( .A(n625), .B(A[168]), .Z(n622) );
  XOR U715 ( .A(n625), .B(n626), .Z(SUM[168]) );
  XNOR U716 ( .A(B[168]), .B(A[168]), .Z(n626) );
  AND U717 ( .A(n627), .B(n628), .Z(n625) );
  NAND U718 ( .A(B[167]), .B(n629), .Z(n628) );
  NANDN U719 ( .A(A[167]), .B(n630), .Z(n629) );
  NANDN U720 ( .A(n630), .B(A[167]), .Z(n627) );
  XOR U721 ( .A(n630), .B(n631), .Z(SUM[167]) );
  XNOR U722 ( .A(B[167]), .B(A[167]), .Z(n631) );
  AND U723 ( .A(n632), .B(n633), .Z(n630) );
  NAND U724 ( .A(B[166]), .B(n634), .Z(n633) );
  NANDN U725 ( .A(A[166]), .B(n635), .Z(n634) );
  NANDN U726 ( .A(n635), .B(A[166]), .Z(n632) );
  XOR U727 ( .A(n635), .B(n636), .Z(SUM[166]) );
  XNOR U728 ( .A(B[166]), .B(A[166]), .Z(n636) );
  AND U729 ( .A(n637), .B(n638), .Z(n635) );
  NAND U730 ( .A(B[165]), .B(n639), .Z(n638) );
  NANDN U731 ( .A(A[165]), .B(n640), .Z(n639) );
  NANDN U732 ( .A(n640), .B(A[165]), .Z(n637) );
  XOR U733 ( .A(n640), .B(n641), .Z(SUM[165]) );
  XNOR U734 ( .A(B[165]), .B(A[165]), .Z(n641) );
  AND U735 ( .A(n642), .B(n643), .Z(n640) );
  NAND U736 ( .A(B[164]), .B(n644), .Z(n643) );
  NANDN U737 ( .A(A[164]), .B(n645), .Z(n644) );
  NANDN U738 ( .A(n645), .B(A[164]), .Z(n642) );
  XOR U739 ( .A(n645), .B(n646), .Z(SUM[164]) );
  XNOR U740 ( .A(B[164]), .B(A[164]), .Z(n646) );
  AND U741 ( .A(n647), .B(n648), .Z(n645) );
  NAND U742 ( .A(B[163]), .B(n649), .Z(n648) );
  NANDN U743 ( .A(A[163]), .B(n650), .Z(n649) );
  NANDN U744 ( .A(n650), .B(A[163]), .Z(n647) );
  XOR U745 ( .A(n650), .B(n651), .Z(SUM[163]) );
  XNOR U746 ( .A(B[163]), .B(A[163]), .Z(n651) );
  AND U747 ( .A(n652), .B(n653), .Z(n650) );
  NAND U748 ( .A(B[162]), .B(n654), .Z(n653) );
  NANDN U749 ( .A(A[162]), .B(n655), .Z(n654) );
  NANDN U750 ( .A(n655), .B(A[162]), .Z(n652) );
  XOR U751 ( .A(n655), .B(n656), .Z(SUM[162]) );
  XNOR U752 ( .A(B[162]), .B(A[162]), .Z(n656) );
  AND U753 ( .A(n657), .B(n658), .Z(n655) );
  NAND U754 ( .A(B[161]), .B(n659), .Z(n658) );
  NANDN U755 ( .A(A[161]), .B(n660), .Z(n659) );
  NANDN U756 ( .A(n660), .B(A[161]), .Z(n657) );
  XOR U757 ( .A(n660), .B(n661), .Z(SUM[161]) );
  XNOR U758 ( .A(B[161]), .B(A[161]), .Z(n661) );
  AND U759 ( .A(n662), .B(n663), .Z(n660) );
  NAND U760 ( .A(B[160]), .B(n664), .Z(n663) );
  NANDN U761 ( .A(A[160]), .B(n665), .Z(n664) );
  NANDN U762 ( .A(n665), .B(A[160]), .Z(n662) );
  XOR U763 ( .A(n665), .B(n666), .Z(SUM[160]) );
  XNOR U764 ( .A(B[160]), .B(A[160]), .Z(n666) );
  AND U765 ( .A(n667), .B(n668), .Z(n665) );
  NAND U766 ( .A(B[159]), .B(n669), .Z(n668) );
  NANDN U767 ( .A(A[159]), .B(n670), .Z(n669) );
  NANDN U768 ( .A(n670), .B(A[159]), .Z(n667) );
  XOR U769 ( .A(n671), .B(n672), .Z(SUM[15]) );
  XNOR U770 ( .A(B[15]), .B(A[15]), .Z(n672) );
  XOR U771 ( .A(n670), .B(n673), .Z(SUM[159]) );
  XNOR U772 ( .A(B[159]), .B(A[159]), .Z(n673) );
  AND U773 ( .A(n674), .B(n675), .Z(n670) );
  NAND U774 ( .A(B[158]), .B(n676), .Z(n675) );
  NANDN U775 ( .A(A[158]), .B(n677), .Z(n676) );
  NANDN U776 ( .A(n677), .B(A[158]), .Z(n674) );
  XOR U777 ( .A(n677), .B(n678), .Z(SUM[158]) );
  XNOR U778 ( .A(B[158]), .B(A[158]), .Z(n678) );
  AND U779 ( .A(n679), .B(n680), .Z(n677) );
  NAND U780 ( .A(B[157]), .B(n681), .Z(n680) );
  NANDN U781 ( .A(A[157]), .B(n682), .Z(n681) );
  NANDN U782 ( .A(n682), .B(A[157]), .Z(n679) );
  XOR U783 ( .A(n682), .B(n683), .Z(SUM[157]) );
  XNOR U784 ( .A(B[157]), .B(A[157]), .Z(n683) );
  AND U785 ( .A(n684), .B(n685), .Z(n682) );
  NAND U786 ( .A(B[156]), .B(n686), .Z(n685) );
  NANDN U787 ( .A(A[156]), .B(n687), .Z(n686) );
  NANDN U788 ( .A(n687), .B(A[156]), .Z(n684) );
  XOR U789 ( .A(n687), .B(n688), .Z(SUM[156]) );
  XNOR U790 ( .A(B[156]), .B(A[156]), .Z(n688) );
  AND U791 ( .A(n689), .B(n690), .Z(n687) );
  NAND U792 ( .A(B[155]), .B(n691), .Z(n690) );
  NANDN U793 ( .A(A[155]), .B(n692), .Z(n691) );
  NANDN U794 ( .A(n692), .B(A[155]), .Z(n689) );
  XOR U795 ( .A(n692), .B(n693), .Z(SUM[155]) );
  XNOR U796 ( .A(B[155]), .B(A[155]), .Z(n693) );
  AND U797 ( .A(n694), .B(n695), .Z(n692) );
  NAND U798 ( .A(B[154]), .B(n696), .Z(n695) );
  NANDN U799 ( .A(A[154]), .B(n697), .Z(n696) );
  NANDN U800 ( .A(n697), .B(A[154]), .Z(n694) );
  XOR U801 ( .A(n697), .B(n698), .Z(SUM[154]) );
  XNOR U802 ( .A(B[154]), .B(A[154]), .Z(n698) );
  AND U803 ( .A(n699), .B(n700), .Z(n697) );
  NAND U804 ( .A(B[153]), .B(n701), .Z(n700) );
  NANDN U805 ( .A(A[153]), .B(n702), .Z(n701) );
  NANDN U806 ( .A(n702), .B(A[153]), .Z(n699) );
  XOR U807 ( .A(n702), .B(n703), .Z(SUM[153]) );
  XNOR U808 ( .A(B[153]), .B(A[153]), .Z(n703) );
  AND U809 ( .A(n704), .B(n705), .Z(n702) );
  NAND U810 ( .A(B[152]), .B(n706), .Z(n705) );
  NANDN U811 ( .A(A[152]), .B(n707), .Z(n706) );
  NANDN U812 ( .A(n707), .B(A[152]), .Z(n704) );
  XOR U813 ( .A(n707), .B(n708), .Z(SUM[152]) );
  XNOR U814 ( .A(B[152]), .B(A[152]), .Z(n708) );
  AND U815 ( .A(n709), .B(n710), .Z(n707) );
  NAND U816 ( .A(B[151]), .B(n711), .Z(n710) );
  NANDN U817 ( .A(A[151]), .B(n712), .Z(n711) );
  NANDN U818 ( .A(n712), .B(A[151]), .Z(n709) );
  XOR U819 ( .A(n712), .B(n713), .Z(SUM[151]) );
  XNOR U820 ( .A(B[151]), .B(A[151]), .Z(n713) );
  AND U821 ( .A(n714), .B(n715), .Z(n712) );
  NAND U822 ( .A(B[150]), .B(n716), .Z(n715) );
  NANDN U823 ( .A(A[150]), .B(n717), .Z(n716) );
  NANDN U824 ( .A(n717), .B(A[150]), .Z(n714) );
  XOR U825 ( .A(n717), .B(n718), .Z(SUM[150]) );
  XNOR U826 ( .A(B[150]), .B(A[150]), .Z(n718) );
  AND U827 ( .A(n719), .B(n720), .Z(n717) );
  NAND U828 ( .A(B[149]), .B(n721), .Z(n720) );
  NANDN U829 ( .A(A[149]), .B(n722), .Z(n721) );
  NANDN U830 ( .A(n722), .B(A[149]), .Z(n719) );
  XOR U831 ( .A(n723), .B(n724), .Z(SUM[14]) );
  XNOR U832 ( .A(B[14]), .B(A[14]), .Z(n724) );
  XOR U833 ( .A(n722), .B(n725), .Z(SUM[149]) );
  XNOR U834 ( .A(B[149]), .B(A[149]), .Z(n725) );
  AND U835 ( .A(n726), .B(n727), .Z(n722) );
  NAND U836 ( .A(B[148]), .B(n728), .Z(n727) );
  NANDN U837 ( .A(A[148]), .B(n729), .Z(n728) );
  NANDN U838 ( .A(n729), .B(A[148]), .Z(n726) );
  XOR U839 ( .A(n729), .B(n730), .Z(SUM[148]) );
  XNOR U840 ( .A(B[148]), .B(A[148]), .Z(n730) );
  AND U841 ( .A(n731), .B(n732), .Z(n729) );
  NAND U842 ( .A(B[147]), .B(n733), .Z(n732) );
  NANDN U843 ( .A(A[147]), .B(n734), .Z(n733) );
  NANDN U844 ( .A(n734), .B(A[147]), .Z(n731) );
  XOR U845 ( .A(n734), .B(n735), .Z(SUM[147]) );
  XNOR U846 ( .A(B[147]), .B(A[147]), .Z(n735) );
  AND U847 ( .A(n736), .B(n737), .Z(n734) );
  NAND U848 ( .A(B[146]), .B(n738), .Z(n737) );
  NANDN U849 ( .A(A[146]), .B(n739), .Z(n738) );
  NANDN U850 ( .A(n739), .B(A[146]), .Z(n736) );
  XOR U851 ( .A(n739), .B(n740), .Z(SUM[146]) );
  XNOR U852 ( .A(B[146]), .B(A[146]), .Z(n740) );
  AND U853 ( .A(n741), .B(n742), .Z(n739) );
  NAND U854 ( .A(B[145]), .B(n743), .Z(n742) );
  NANDN U855 ( .A(A[145]), .B(n744), .Z(n743) );
  NANDN U856 ( .A(n744), .B(A[145]), .Z(n741) );
  XOR U857 ( .A(n744), .B(n745), .Z(SUM[145]) );
  XNOR U858 ( .A(B[145]), .B(A[145]), .Z(n745) );
  AND U859 ( .A(n746), .B(n747), .Z(n744) );
  NAND U860 ( .A(B[144]), .B(n748), .Z(n747) );
  NANDN U861 ( .A(A[144]), .B(n749), .Z(n748) );
  NANDN U862 ( .A(n749), .B(A[144]), .Z(n746) );
  XOR U863 ( .A(n749), .B(n750), .Z(SUM[144]) );
  XNOR U864 ( .A(B[144]), .B(A[144]), .Z(n750) );
  AND U865 ( .A(n751), .B(n752), .Z(n749) );
  NAND U866 ( .A(B[143]), .B(n753), .Z(n752) );
  NANDN U867 ( .A(A[143]), .B(n754), .Z(n753) );
  NANDN U868 ( .A(n754), .B(A[143]), .Z(n751) );
  XOR U869 ( .A(n754), .B(n755), .Z(SUM[143]) );
  XNOR U870 ( .A(B[143]), .B(A[143]), .Z(n755) );
  AND U871 ( .A(n756), .B(n757), .Z(n754) );
  NAND U872 ( .A(B[142]), .B(n758), .Z(n757) );
  NANDN U873 ( .A(A[142]), .B(n759), .Z(n758) );
  NANDN U874 ( .A(n759), .B(A[142]), .Z(n756) );
  XOR U875 ( .A(n759), .B(n760), .Z(SUM[142]) );
  XNOR U876 ( .A(B[142]), .B(A[142]), .Z(n760) );
  AND U877 ( .A(n761), .B(n762), .Z(n759) );
  NAND U878 ( .A(B[141]), .B(n763), .Z(n762) );
  NANDN U879 ( .A(A[141]), .B(n764), .Z(n763) );
  NANDN U880 ( .A(n764), .B(A[141]), .Z(n761) );
  XOR U881 ( .A(n764), .B(n765), .Z(SUM[141]) );
  XNOR U882 ( .A(B[141]), .B(A[141]), .Z(n765) );
  AND U883 ( .A(n766), .B(n767), .Z(n764) );
  NAND U884 ( .A(B[140]), .B(n768), .Z(n767) );
  NANDN U885 ( .A(A[140]), .B(n769), .Z(n768) );
  NANDN U886 ( .A(n769), .B(A[140]), .Z(n766) );
  XOR U887 ( .A(n769), .B(n770), .Z(SUM[140]) );
  XNOR U888 ( .A(B[140]), .B(A[140]), .Z(n770) );
  AND U889 ( .A(n771), .B(n772), .Z(n769) );
  NAND U890 ( .A(B[139]), .B(n773), .Z(n772) );
  NANDN U891 ( .A(A[139]), .B(n774), .Z(n773) );
  NANDN U892 ( .A(n774), .B(A[139]), .Z(n771) );
  XOR U893 ( .A(n775), .B(n776), .Z(SUM[13]) );
  XNOR U894 ( .A(B[13]), .B(A[13]), .Z(n776) );
  XOR U895 ( .A(n774), .B(n777), .Z(SUM[139]) );
  XNOR U896 ( .A(B[139]), .B(A[139]), .Z(n777) );
  AND U897 ( .A(n778), .B(n779), .Z(n774) );
  NAND U898 ( .A(B[138]), .B(n780), .Z(n779) );
  NANDN U899 ( .A(A[138]), .B(n781), .Z(n780) );
  NANDN U900 ( .A(n781), .B(A[138]), .Z(n778) );
  XOR U901 ( .A(n781), .B(n782), .Z(SUM[138]) );
  XNOR U902 ( .A(B[138]), .B(A[138]), .Z(n782) );
  AND U903 ( .A(n783), .B(n784), .Z(n781) );
  NAND U904 ( .A(B[137]), .B(n785), .Z(n784) );
  NANDN U905 ( .A(A[137]), .B(n786), .Z(n785) );
  NANDN U906 ( .A(n786), .B(A[137]), .Z(n783) );
  XOR U907 ( .A(n786), .B(n787), .Z(SUM[137]) );
  XNOR U908 ( .A(B[137]), .B(A[137]), .Z(n787) );
  AND U909 ( .A(n788), .B(n789), .Z(n786) );
  NAND U910 ( .A(B[136]), .B(n790), .Z(n789) );
  NANDN U911 ( .A(A[136]), .B(n791), .Z(n790) );
  NANDN U912 ( .A(n791), .B(A[136]), .Z(n788) );
  XOR U913 ( .A(n791), .B(n792), .Z(SUM[136]) );
  XNOR U914 ( .A(B[136]), .B(A[136]), .Z(n792) );
  AND U915 ( .A(n793), .B(n794), .Z(n791) );
  NAND U916 ( .A(B[135]), .B(n795), .Z(n794) );
  NANDN U917 ( .A(A[135]), .B(n796), .Z(n795) );
  NANDN U918 ( .A(n796), .B(A[135]), .Z(n793) );
  XOR U919 ( .A(n796), .B(n797), .Z(SUM[135]) );
  XNOR U920 ( .A(B[135]), .B(A[135]), .Z(n797) );
  AND U921 ( .A(n798), .B(n799), .Z(n796) );
  NAND U922 ( .A(B[134]), .B(n800), .Z(n799) );
  NANDN U923 ( .A(A[134]), .B(n801), .Z(n800) );
  NANDN U924 ( .A(n801), .B(A[134]), .Z(n798) );
  XOR U925 ( .A(n801), .B(n802), .Z(SUM[134]) );
  XNOR U926 ( .A(B[134]), .B(A[134]), .Z(n802) );
  AND U927 ( .A(n803), .B(n804), .Z(n801) );
  NAND U928 ( .A(B[133]), .B(n805), .Z(n804) );
  NANDN U929 ( .A(A[133]), .B(n806), .Z(n805) );
  NANDN U930 ( .A(n806), .B(A[133]), .Z(n803) );
  XOR U931 ( .A(n806), .B(n807), .Z(SUM[133]) );
  XNOR U932 ( .A(B[133]), .B(A[133]), .Z(n807) );
  AND U933 ( .A(n808), .B(n809), .Z(n806) );
  NAND U934 ( .A(B[132]), .B(n810), .Z(n809) );
  NANDN U935 ( .A(A[132]), .B(n811), .Z(n810) );
  NANDN U936 ( .A(n811), .B(A[132]), .Z(n808) );
  XOR U937 ( .A(n811), .B(n812), .Z(SUM[132]) );
  XNOR U938 ( .A(B[132]), .B(A[132]), .Z(n812) );
  AND U939 ( .A(n813), .B(n814), .Z(n811) );
  NAND U940 ( .A(B[131]), .B(n815), .Z(n814) );
  NANDN U941 ( .A(A[131]), .B(n816), .Z(n815) );
  NANDN U942 ( .A(n816), .B(A[131]), .Z(n813) );
  XOR U943 ( .A(n816), .B(n817), .Z(SUM[131]) );
  XNOR U944 ( .A(B[131]), .B(A[131]), .Z(n817) );
  AND U945 ( .A(n818), .B(n819), .Z(n816) );
  NAND U946 ( .A(B[130]), .B(n820), .Z(n819) );
  NANDN U947 ( .A(A[130]), .B(n821), .Z(n820) );
  NANDN U948 ( .A(n821), .B(A[130]), .Z(n818) );
  XOR U949 ( .A(n821), .B(n822), .Z(SUM[130]) );
  XNOR U950 ( .A(B[130]), .B(A[130]), .Z(n822) );
  AND U951 ( .A(n823), .B(n824), .Z(n821) );
  NAND U952 ( .A(B[129]), .B(n825), .Z(n824) );
  NANDN U953 ( .A(A[129]), .B(n826), .Z(n825) );
  NANDN U954 ( .A(n826), .B(A[129]), .Z(n823) );
  XOR U955 ( .A(n827), .B(n828), .Z(SUM[12]) );
  XNOR U956 ( .A(B[12]), .B(A[12]), .Z(n828) );
  XOR U957 ( .A(n826), .B(n829), .Z(SUM[129]) );
  XNOR U958 ( .A(B[129]), .B(A[129]), .Z(n829) );
  AND U959 ( .A(n830), .B(n831), .Z(n826) );
  NAND U960 ( .A(B[128]), .B(n832), .Z(n831) );
  NANDN U961 ( .A(A[128]), .B(n833), .Z(n832) );
  NANDN U962 ( .A(n833), .B(A[128]), .Z(n830) );
  XOR U963 ( .A(n833), .B(n834), .Z(SUM[128]) );
  XNOR U964 ( .A(B[128]), .B(A[128]), .Z(n834) );
  AND U965 ( .A(n835), .B(n836), .Z(n833) );
  NAND U966 ( .A(B[127]), .B(n837), .Z(n836) );
  NANDN U967 ( .A(A[127]), .B(n838), .Z(n837) );
  NANDN U968 ( .A(n838), .B(A[127]), .Z(n835) );
  XOR U969 ( .A(n838), .B(n839), .Z(SUM[127]) );
  XNOR U970 ( .A(B[127]), .B(A[127]), .Z(n839) );
  AND U971 ( .A(n840), .B(n841), .Z(n838) );
  NAND U972 ( .A(B[126]), .B(n842), .Z(n841) );
  NANDN U973 ( .A(A[126]), .B(n843), .Z(n842) );
  NANDN U974 ( .A(n843), .B(A[126]), .Z(n840) );
  XOR U975 ( .A(n843), .B(n844), .Z(SUM[126]) );
  XNOR U976 ( .A(B[126]), .B(A[126]), .Z(n844) );
  AND U977 ( .A(n845), .B(n846), .Z(n843) );
  NAND U978 ( .A(B[125]), .B(n847), .Z(n846) );
  NANDN U979 ( .A(A[125]), .B(n848), .Z(n847) );
  NANDN U980 ( .A(n848), .B(A[125]), .Z(n845) );
  XOR U981 ( .A(n848), .B(n849), .Z(SUM[125]) );
  XNOR U982 ( .A(B[125]), .B(A[125]), .Z(n849) );
  AND U983 ( .A(n850), .B(n851), .Z(n848) );
  NAND U984 ( .A(B[124]), .B(n852), .Z(n851) );
  NANDN U985 ( .A(A[124]), .B(n853), .Z(n852) );
  NANDN U986 ( .A(n853), .B(A[124]), .Z(n850) );
  XOR U987 ( .A(n853), .B(n854), .Z(SUM[124]) );
  XNOR U988 ( .A(B[124]), .B(A[124]), .Z(n854) );
  AND U989 ( .A(n855), .B(n856), .Z(n853) );
  NAND U990 ( .A(B[123]), .B(n857), .Z(n856) );
  NANDN U991 ( .A(A[123]), .B(n858), .Z(n857) );
  NANDN U992 ( .A(n858), .B(A[123]), .Z(n855) );
  XOR U993 ( .A(n858), .B(n859), .Z(SUM[123]) );
  XNOR U994 ( .A(B[123]), .B(A[123]), .Z(n859) );
  AND U995 ( .A(n860), .B(n861), .Z(n858) );
  NAND U996 ( .A(B[122]), .B(n862), .Z(n861) );
  NANDN U997 ( .A(A[122]), .B(n863), .Z(n862) );
  NANDN U998 ( .A(n863), .B(A[122]), .Z(n860) );
  XOR U999 ( .A(n863), .B(n864), .Z(SUM[122]) );
  XNOR U1000 ( .A(B[122]), .B(A[122]), .Z(n864) );
  AND U1001 ( .A(n865), .B(n866), .Z(n863) );
  NAND U1002 ( .A(B[121]), .B(n867), .Z(n866) );
  NANDN U1003 ( .A(A[121]), .B(n868), .Z(n867) );
  NANDN U1004 ( .A(n868), .B(A[121]), .Z(n865) );
  XOR U1005 ( .A(n868), .B(n869), .Z(SUM[121]) );
  XNOR U1006 ( .A(B[121]), .B(A[121]), .Z(n869) );
  AND U1007 ( .A(n870), .B(n871), .Z(n868) );
  NAND U1008 ( .A(B[120]), .B(n872), .Z(n871) );
  NANDN U1009 ( .A(A[120]), .B(n873), .Z(n872) );
  NANDN U1010 ( .A(n873), .B(A[120]), .Z(n870) );
  XOR U1011 ( .A(n873), .B(n874), .Z(SUM[120]) );
  XNOR U1012 ( .A(B[120]), .B(A[120]), .Z(n874) );
  AND U1013 ( .A(n875), .B(n876), .Z(n873) );
  NAND U1014 ( .A(B[119]), .B(n877), .Z(n876) );
  NANDN U1015 ( .A(A[119]), .B(n878), .Z(n877) );
  NANDN U1016 ( .A(n878), .B(A[119]), .Z(n875) );
  XOR U1017 ( .A(n879), .B(n880), .Z(SUM[11]) );
  XNOR U1018 ( .A(B[11]), .B(A[11]), .Z(n880) );
  XOR U1019 ( .A(n878), .B(n881), .Z(SUM[119]) );
  XNOR U1020 ( .A(B[119]), .B(A[119]), .Z(n881) );
  AND U1021 ( .A(n882), .B(n883), .Z(n878) );
  NAND U1022 ( .A(B[118]), .B(n884), .Z(n883) );
  NANDN U1023 ( .A(A[118]), .B(n885), .Z(n884) );
  NANDN U1024 ( .A(n885), .B(A[118]), .Z(n882) );
  XOR U1025 ( .A(n885), .B(n886), .Z(SUM[118]) );
  XNOR U1026 ( .A(B[118]), .B(A[118]), .Z(n886) );
  AND U1027 ( .A(n887), .B(n888), .Z(n885) );
  NAND U1028 ( .A(B[117]), .B(n889), .Z(n888) );
  NANDN U1029 ( .A(A[117]), .B(n890), .Z(n889) );
  NANDN U1030 ( .A(n890), .B(A[117]), .Z(n887) );
  XOR U1031 ( .A(n890), .B(n891), .Z(SUM[117]) );
  XNOR U1032 ( .A(B[117]), .B(A[117]), .Z(n891) );
  AND U1033 ( .A(n892), .B(n893), .Z(n890) );
  NAND U1034 ( .A(B[116]), .B(n894), .Z(n893) );
  NANDN U1035 ( .A(A[116]), .B(n895), .Z(n894) );
  NANDN U1036 ( .A(n895), .B(A[116]), .Z(n892) );
  XOR U1037 ( .A(n895), .B(n896), .Z(SUM[116]) );
  XNOR U1038 ( .A(B[116]), .B(A[116]), .Z(n896) );
  AND U1039 ( .A(n897), .B(n898), .Z(n895) );
  NAND U1040 ( .A(B[115]), .B(n899), .Z(n898) );
  NANDN U1041 ( .A(A[115]), .B(n900), .Z(n899) );
  NANDN U1042 ( .A(n900), .B(A[115]), .Z(n897) );
  XOR U1043 ( .A(n900), .B(n901), .Z(SUM[115]) );
  XNOR U1044 ( .A(B[115]), .B(A[115]), .Z(n901) );
  AND U1045 ( .A(n902), .B(n903), .Z(n900) );
  NAND U1046 ( .A(B[114]), .B(n904), .Z(n903) );
  NANDN U1047 ( .A(A[114]), .B(n905), .Z(n904) );
  NANDN U1048 ( .A(n905), .B(A[114]), .Z(n902) );
  XOR U1049 ( .A(n905), .B(n906), .Z(SUM[114]) );
  XNOR U1050 ( .A(B[114]), .B(A[114]), .Z(n906) );
  AND U1051 ( .A(n907), .B(n908), .Z(n905) );
  NAND U1052 ( .A(B[113]), .B(n909), .Z(n908) );
  NANDN U1053 ( .A(A[113]), .B(n910), .Z(n909) );
  NANDN U1054 ( .A(n910), .B(A[113]), .Z(n907) );
  XOR U1055 ( .A(n910), .B(n911), .Z(SUM[113]) );
  XNOR U1056 ( .A(B[113]), .B(A[113]), .Z(n911) );
  AND U1057 ( .A(n912), .B(n913), .Z(n910) );
  NAND U1058 ( .A(B[112]), .B(n914), .Z(n913) );
  NANDN U1059 ( .A(A[112]), .B(n915), .Z(n914) );
  NANDN U1060 ( .A(n915), .B(A[112]), .Z(n912) );
  XOR U1061 ( .A(n915), .B(n916), .Z(SUM[112]) );
  XNOR U1062 ( .A(B[112]), .B(A[112]), .Z(n916) );
  AND U1063 ( .A(n917), .B(n918), .Z(n915) );
  NAND U1064 ( .A(B[111]), .B(n919), .Z(n918) );
  NANDN U1065 ( .A(A[111]), .B(n920), .Z(n919) );
  NANDN U1066 ( .A(n920), .B(A[111]), .Z(n917) );
  XOR U1067 ( .A(n920), .B(n921), .Z(SUM[111]) );
  XNOR U1068 ( .A(B[111]), .B(A[111]), .Z(n921) );
  AND U1069 ( .A(n922), .B(n923), .Z(n920) );
  NAND U1070 ( .A(B[110]), .B(n924), .Z(n923) );
  NANDN U1071 ( .A(A[110]), .B(n925), .Z(n924) );
  NANDN U1072 ( .A(n925), .B(A[110]), .Z(n922) );
  XOR U1073 ( .A(n925), .B(n926), .Z(SUM[110]) );
  XNOR U1074 ( .A(B[110]), .B(A[110]), .Z(n926) );
  AND U1075 ( .A(n927), .B(n928), .Z(n925) );
  NAND U1076 ( .A(B[109]), .B(n929), .Z(n928) );
  NANDN U1077 ( .A(A[109]), .B(n930), .Z(n929) );
  NANDN U1078 ( .A(n930), .B(A[109]), .Z(n927) );
  XOR U1079 ( .A(n931), .B(n932), .Z(SUM[10]) );
  XNOR U1080 ( .A(B[10]), .B(A[10]), .Z(n932) );
  XOR U1081 ( .A(n930), .B(n933), .Z(SUM[109]) );
  XNOR U1082 ( .A(B[109]), .B(A[109]), .Z(n933) );
  AND U1083 ( .A(n934), .B(n935), .Z(n930) );
  NAND U1084 ( .A(B[108]), .B(n936), .Z(n935) );
  NANDN U1085 ( .A(A[108]), .B(n937), .Z(n936) );
  NANDN U1086 ( .A(n937), .B(A[108]), .Z(n934) );
  XOR U1087 ( .A(n937), .B(n938), .Z(SUM[108]) );
  XNOR U1088 ( .A(B[108]), .B(A[108]), .Z(n938) );
  AND U1089 ( .A(n939), .B(n940), .Z(n937) );
  NAND U1090 ( .A(B[107]), .B(n941), .Z(n940) );
  NANDN U1091 ( .A(A[107]), .B(n942), .Z(n941) );
  NANDN U1092 ( .A(n942), .B(A[107]), .Z(n939) );
  XOR U1093 ( .A(n942), .B(n943), .Z(SUM[107]) );
  XNOR U1094 ( .A(B[107]), .B(A[107]), .Z(n943) );
  AND U1095 ( .A(n944), .B(n945), .Z(n942) );
  NAND U1096 ( .A(B[106]), .B(n946), .Z(n945) );
  NANDN U1097 ( .A(A[106]), .B(n947), .Z(n946) );
  NANDN U1098 ( .A(n947), .B(A[106]), .Z(n944) );
  XOR U1099 ( .A(n947), .B(n948), .Z(SUM[106]) );
  XNOR U1100 ( .A(B[106]), .B(A[106]), .Z(n948) );
  AND U1101 ( .A(n949), .B(n950), .Z(n947) );
  NAND U1102 ( .A(B[105]), .B(n951), .Z(n950) );
  NANDN U1103 ( .A(A[105]), .B(n952), .Z(n951) );
  NANDN U1104 ( .A(n952), .B(A[105]), .Z(n949) );
  XOR U1105 ( .A(n952), .B(n953), .Z(SUM[105]) );
  XNOR U1106 ( .A(B[105]), .B(A[105]), .Z(n953) );
  AND U1107 ( .A(n954), .B(n955), .Z(n952) );
  NAND U1108 ( .A(B[104]), .B(n956), .Z(n955) );
  NANDN U1109 ( .A(A[104]), .B(n957), .Z(n956) );
  NANDN U1110 ( .A(n957), .B(A[104]), .Z(n954) );
  XOR U1111 ( .A(n957), .B(n958), .Z(SUM[104]) );
  XNOR U1112 ( .A(B[104]), .B(A[104]), .Z(n958) );
  AND U1113 ( .A(n959), .B(n960), .Z(n957) );
  NAND U1114 ( .A(B[103]), .B(n961), .Z(n960) );
  NANDN U1115 ( .A(A[103]), .B(n962), .Z(n961) );
  NANDN U1116 ( .A(n962), .B(A[103]), .Z(n959) );
  XOR U1117 ( .A(n962), .B(n963), .Z(SUM[103]) );
  XNOR U1118 ( .A(B[103]), .B(A[103]), .Z(n963) );
  AND U1119 ( .A(n964), .B(n965), .Z(n962) );
  NAND U1120 ( .A(B[102]), .B(n966), .Z(n965) );
  NANDN U1121 ( .A(A[102]), .B(n967), .Z(n966) );
  NANDN U1122 ( .A(n967), .B(A[102]), .Z(n964) );
  XOR U1123 ( .A(n967), .B(n968), .Z(SUM[102]) );
  XNOR U1124 ( .A(B[102]), .B(A[102]), .Z(n968) );
  AND U1125 ( .A(n969), .B(n970), .Z(n967) );
  NAND U1126 ( .A(B[101]), .B(n971), .Z(n970) );
  NANDN U1127 ( .A(A[101]), .B(n972), .Z(n971) );
  NANDN U1128 ( .A(n972), .B(A[101]), .Z(n969) );
  XOR U1129 ( .A(n972), .B(n973), .Z(SUM[101]) );
  XNOR U1130 ( .A(B[101]), .B(A[101]), .Z(n973) );
  AND U1131 ( .A(n974), .B(n975), .Z(n972) );
  NAND U1132 ( .A(B[100]), .B(n976), .Z(n975) );
  NANDN U1133 ( .A(A[100]), .B(n977), .Z(n976) );
  NANDN U1134 ( .A(n977), .B(A[100]), .Z(n974) );
  XOR U1135 ( .A(n977), .B(n978), .Z(SUM[100]) );
  XNOR U1136 ( .A(B[100]), .B(A[100]), .Z(n978) );
  AND U1137 ( .A(n979), .B(n980), .Z(n977) );
  NAND U1138 ( .A(B[99]), .B(n981), .Z(n980) );
  OR U1139 ( .A(n3), .B(A[99]), .Z(n981) );
  NAND U1140 ( .A(A[99]), .B(n3), .Z(n979) );
  NAND U1141 ( .A(n982), .B(n983), .Z(n3) );
  NAND U1142 ( .A(B[98]), .B(n984), .Z(n983) );
  NANDN U1143 ( .A(A[98]), .B(n5), .Z(n984) );
  NANDN U1144 ( .A(n5), .B(A[98]), .Z(n982) );
  AND U1145 ( .A(n985), .B(n986), .Z(n5) );
  NAND U1146 ( .A(B[97]), .B(n987), .Z(n986) );
  NANDN U1147 ( .A(A[97]), .B(n7), .Z(n987) );
  NANDN U1148 ( .A(n7), .B(A[97]), .Z(n985) );
  AND U1149 ( .A(n988), .B(n989), .Z(n7) );
  NAND U1150 ( .A(B[96]), .B(n990), .Z(n989) );
  NANDN U1151 ( .A(A[96]), .B(n9), .Z(n990) );
  NANDN U1152 ( .A(n9), .B(A[96]), .Z(n988) );
  AND U1153 ( .A(n991), .B(n992), .Z(n9) );
  NAND U1154 ( .A(B[95]), .B(n993), .Z(n992) );
  NANDN U1155 ( .A(A[95]), .B(n11), .Z(n993) );
  NANDN U1156 ( .A(n11), .B(A[95]), .Z(n991) );
  AND U1157 ( .A(n994), .B(n995), .Z(n11) );
  NAND U1158 ( .A(B[94]), .B(n996), .Z(n995) );
  NANDN U1159 ( .A(A[94]), .B(n13), .Z(n996) );
  NANDN U1160 ( .A(n13), .B(A[94]), .Z(n994) );
  AND U1161 ( .A(n997), .B(n998), .Z(n13) );
  NAND U1162 ( .A(B[93]), .B(n999), .Z(n998) );
  NANDN U1163 ( .A(A[93]), .B(n15), .Z(n999) );
  NANDN U1164 ( .A(n15), .B(A[93]), .Z(n997) );
  AND U1165 ( .A(n1000), .B(n1001), .Z(n15) );
  NAND U1166 ( .A(B[92]), .B(n1002), .Z(n1001) );
  NANDN U1167 ( .A(A[92]), .B(n17), .Z(n1002) );
  NANDN U1168 ( .A(n17), .B(A[92]), .Z(n1000) );
  AND U1169 ( .A(n1003), .B(n1004), .Z(n17) );
  NAND U1170 ( .A(B[91]), .B(n1005), .Z(n1004) );
  NANDN U1171 ( .A(A[91]), .B(n19), .Z(n1005) );
  NANDN U1172 ( .A(n19), .B(A[91]), .Z(n1003) );
  AND U1173 ( .A(n1006), .B(n1007), .Z(n19) );
  NAND U1174 ( .A(B[90]), .B(n1008), .Z(n1007) );
  NANDN U1175 ( .A(A[90]), .B(n21), .Z(n1008) );
  NANDN U1176 ( .A(n21), .B(A[90]), .Z(n1006) );
  AND U1177 ( .A(n1009), .B(n1010), .Z(n21) );
  NAND U1178 ( .A(B[89]), .B(n1011), .Z(n1010) );
  NANDN U1179 ( .A(A[89]), .B(n25), .Z(n1011) );
  NANDN U1180 ( .A(n25), .B(A[89]), .Z(n1009) );
  AND U1181 ( .A(n1012), .B(n1013), .Z(n25) );
  NAND U1182 ( .A(B[88]), .B(n1014), .Z(n1013) );
  NANDN U1183 ( .A(A[88]), .B(n27), .Z(n1014) );
  NANDN U1184 ( .A(n27), .B(A[88]), .Z(n1012) );
  AND U1185 ( .A(n1015), .B(n1016), .Z(n27) );
  NAND U1186 ( .A(B[87]), .B(n1017), .Z(n1016) );
  NANDN U1187 ( .A(A[87]), .B(n29), .Z(n1017) );
  NANDN U1188 ( .A(n29), .B(A[87]), .Z(n1015) );
  AND U1189 ( .A(n1018), .B(n1019), .Z(n29) );
  NAND U1190 ( .A(B[86]), .B(n1020), .Z(n1019) );
  NANDN U1191 ( .A(A[86]), .B(n31), .Z(n1020) );
  NANDN U1192 ( .A(n31), .B(A[86]), .Z(n1018) );
  AND U1193 ( .A(n1021), .B(n1022), .Z(n31) );
  NAND U1194 ( .A(B[85]), .B(n1023), .Z(n1022) );
  NANDN U1195 ( .A(A[85]), .B(n33), .Z(n1023) );
  NANDN U1196 ( .A(n33), .B(A[85]), .Z(n1021) );
  AND U1197 ( .A(n1024), .B(n1025), .Z(n33) );
  NAND U1198 ( .A(B[84]), .B(n1026), .Z(n1025) );
  NANDN U1199 ( .A(A[84]), .B(n35), .Z(n1026) );
  NANDN U1200 ( .A(n35), .B(A[84]), .Z(n1024) );
  AND U1201 ( .A(n1027), .B(n1028), .Z(n35) );
  NAND U1202 ( .A(B[83]), .B(n1029), .Z(n1028) );
  NANDN U1203 ( .A(A[83]), .B(n37), .Z(n1029) );
  NANDN U1204 ( .A(n37), .B(A[83]), .Z(n1027) );
  AND U1205 ( .A(n1030), .B(n1031), .Z(n37) );
  NAND U1206 ( .A(B[82]), .B(n1032), .Z(n1031) );
  NANDN U1207 ( .A(A[82]), .B(n39), .Z(n1032) );
  NANDN U1208 ( .A(n39), .B(A[82]), .Z(n1030) );
  AND U1209 ( .A(n1033), .B(n1034), .Z(n39) );
  NAND U1210 ( .A(B[81]), .B(n1035), .Z(n1034) );
  NANDN U1211 ( .A(A[81]), .B(n41), .Z(n1035) );
  NANDN U1212 ( .A(n41), .B(A[81]), .Z(n1033) );
  AND U1213 ( .A(n1036), .B(n1037), .Z(n41) );
  NAND U1214 ( .A(B[80]), .B(n1038), .Z(n1037) );
  NANDN U1215 ( .A(A[80]), .B(n43), .Z(n1038) );
  NANDN U1216 ( .A(n43), .B(A[80]), .Z(n1036) );
  AND U1217 ( .A(n1039), .B(n1040), .Z(n43) );
  NAND U1218 ( .A(B[79]), .B(n1041), .Z(n1040) );
  NANDN U1219 ( .A(A[79]), .B(n47), .Z(n1041) );
  NANDN U1220 ( .A(n47), .B(A[79]), .Z(n1039) );
  AND U1221 ( .A(n1042), .B(n1043), .Z(n47) );
  NAND U1222 ( .A(B[78]), .B(n1044), .Z(n1043) );
  NANDN U1223 ( .A(A[78]), .B(n49), .Z(n1044) );
  NANDN U1224 ( .A(n49), .B(A[78]), .Z(n1042) );
  AND U1225 ( .A(n1045), .B(n1046), .Z(n49) );
  NAND U1226 ( .A(B[77]), .B(n1047), .Z(n1046) );
  NANDN U1227 ( .A(A[77]), .B(n51), .Z(n1047) );
  NANDN U1228 ( .A(n51), .B(A[77]), .Z(n1045) );
  AND U1229 ( .A(n1048), .B(n1049), .Z(n51) );
  NAND U1230 ( .A(B[76]), .B(n1050), .Z(n1049) );
  NANDN U1231 ( .A(A[76]), .B(n53), .Z(n1050) );
  NANDN U1232 ( .A(n53), .B(A[76]), .Z(n1048) );
  AND U1233 ( .A(n1051), .B(n1052), .Z(n53) );
  NAND U1234 ( .A(B[75]), .B(n1053), .Z(n1052) );
  NANDN U1235 ( .A(A[75]), .B(n55), .Z(n1053) );
  NANDN U1236 ( .A(n55), .B(A[75]), .Z(n1051) );
  AND U1237 ( .A(n1054), .B(n1055), .Z(n55) );
  NAND U1238 ( .A(B[74]), .B(n1056), .Z(n1055) );
  NANDN U1239 ( .A(A[74]), .B(n57), .Z(n1056) );
  NANDN U1240 ( .A(n57), .B(A[74]), .Z(n1054) );
  AND U1241 ( .A(n1057), .B(n1058), .Z(n57) );
  NAND U1242 ( .A(B[73]), .B(n1059), .Z(n1058) );
  NANDN U1243 ( .A(A[73]), .B(n59), .Z(n1059) );
  NANDN U1244 ( .A(n59), .B(A[73]), .Z(n1057) );
  AND U1245 ( .A(n1060), .B(n1061), .Z(n59) );
  NAND U1246 ( .A(B[72]), .B(n1062), .Z(n1061) );
  NANDN U1247 ( .A(A[72]), .B(n61), .Z(n1062) );
  NANDN U1248 ( .A(n61), .B(A[72]), .Z(n1060) );
  AND U1249 ( .A(n1063), .B(n1064), .Z(n61) );
  NAND U1250 ( .A(B[71]), .B(n1065), .Z(n1064) );
  NANDN U1251 ( .A(A[71]), .B(n63), .Z(n1065) );
  NANDN U1252 ( .A(n63), .B(A[71]), .Z(n1063) );
  AND U1253 ( .A(n1066), .B(n1067), .Z(n63) );
  NAND U1254 ( .A(B[70]), .B(n1068), .Z(n1067) );
  NANDN U1255 ( .A(A[70]), .B(n65), .Z(n1068) );
  NANDN U1256 ( .A(n65), .B(A[70]), .Z(n1066) );
  AND U1257 ( .A(n1069), .B(n1070), .Z(n65) );
  NAND U1258 ( .A(B[69]), .B(n1071), .Z(n1070) );
  NANDN U1259 ( .A(A[69]), .B(n69), .Z(n1071) );
  NANDN U1260 ( .A(n69), .B(A[69]), .Z(n1069) );
  AND U1261 ( .A(n1072), .B(n1073), .Z(n69) );
  NAND U1262 ( .A(B[68]), .B(n1074), .Z(n1073) );
  NANDN U1263 ( .A(A[68]), .B(n71), .Z(n1074) );
  NANDN U1264 ( .A(n71), .B(A[68]), .Z(n1072) );
  AND U1265 ( .A(n1075), .B(n1076), .Z(n71) );
  NAND U1266 ( .A(B[67]), .B(n1077), .Z(n1076) );
  NANDN U1267 ( .A(A[67]), .B(n73), .Z(n1077) );
  NANDN U1268 ( .A(n73), .B(A[67]), .Z(n1075) );
  AND U1269 ( .A(n1078), .B(n1079), .Z(n73) );
  NAND U1270 ( .A(B[66]), .B(n1080), .Z(n1079) );
  NANDN U1271 ( .A(A[66]), .B(n75), .Z(n1080) );
  NANDN U1272 ( .A(n75), .B(A[66]), .Z(n1078) );
  AND U1273 ( .A(n1081), .B(n1082), .Z(n75) );
  NAND U1274 ( .A(B[65]), .B(n1083), .Z(n1082) );
  NANDN U1275 ( .A(A[65]), .B(n77), .Z(n1083) );
  NANDN U1276 ( .A(n77), .B(A[65]), .Z(n1081) );
  AND U1277 ( .A(n1084), .B(n1085), .Z(n77) );
  NAND U1278 ( .A(B[64]), .B(n1086), .Z(n1085) );
  NANDN U1279 ( .A(A[64]), .B(n79), .Z(n1086) );
  NANDN U1280 ( .A(n79), .B(A[64]), .Z(n1084) );
  AND U1281 ( .A(n1087), .B(n1088), .Z(n79) );
  NAND U1282 ( .A(B[63]), .B(n1089), .Z(n1088) );
  NANDN U1283 ( .A(A[63]), .B(n81), .Z(n1089) );
  NANDN U1284 ( .A(n81), .B(A[63]), .Z(n1087) );
  AND U1285 ( .A(n1090), .B(n1091), .Z(n81) );
  NAND U1286 ( .A(B[62]), .B(n1092), .Z(n1091) );
  NANDN U1287 ( .A(A[62]), .B(n83), .Z(n1092) );
  NANDN U1288 ( .A(n83), .B(A[62]), .Z(n1090) );
  AND U1289 ( .A(n1093), .B(n1094), .Z(n83) );
  NAND U1290 ( .A(B[61]), .B(n1095), .Z(n1094) );
  NANDN U1291 ( .A(A[61]), .B(n85), .Z(n1095) );
  NANDN U1292 ( .A(n85), .B(A[61]), .Z(n1093) );
  AND U1293 ( .A(n1096), .B(n1097), .Z(n85) );
  NAND U1294 ( .A(B[60]), .B(n1098), .Z(n1097) );
  NANDN U1295 ( .A(A[60]), .B(n87), .Z(n1098) );
  NANDN U1296 ( .A(n87), .B(A[60]), .Z(n1096) );
  AND U1297 ( .A(n1099), .B(n1100), .Z(n87) );
  NAND U1298 ( .A(B[59]), .B(n1101), .Z(n1100) );
  NANDN U1299 ( .A(A[59]), .B(n91), .Z(n1101) );
  NANDN U1300 ( .A(n91), .B(A[59]), .Z(n1099) );
  AND U1301 ( .A(n1102), .B(n1103), .Z(n91) );
  NAND U1302 ( .A(B[58]), .B(n1104), .Z(n1103) );
  NANDN U1303 ( .A(A[58]), .B(n93), .Z(n1104) );
  NANDN U1304 ( .A(n93), .B(A[58]), .Z(n1102) );
  AND U1305 ( .A(n1105), .B(n1106), .Z(n93) );
  NAND U1306 ( .A(B[57]), .B(n1107), .Z(n1106) );
  NANDN U1307 ( .A(A[57]), .B(n95), .Z(n1107) );
  NANDN U1308 ( .A(n95), .B(A[57]), .Z(n1105) );
  AND U1309 ( .A(n1108), .B(n1109), .Z(n95) );
  NAND U1310 ( .A(B[56]), .B(n1110), .Z(n1109) );
  NANDN U1311 ( .A(A[56]), .B(n97), .Z(n1110) );
  NANDN U1312 ( .A(n97), .B(A[56]), .Z(n1108) );
  AND U1313 ( .A(n1111), .B(n1112), .Z(n97) );
  NAND U1314 ( .A(B[55]), .B(n1113), .Z(n1112) );
  NANDN U1315 ( .A(A[55]), .B(n99), .Z(n1113) );
  NANDN U1316 ( .A(n99), .B(A[55]), .Z(n1111) );
  AND U1317 ( .A(n1114), .B(n1115), .Z(n99) );
  NAND U1318 ( .A(B[54]), .B(n1116), .Z(n1115) );
  NANDN U1319 ( .A(A[54]), .B(n101), .Z(n1116) );
  NANDN U1320 ( .A(n101), .B(A[54]), .Z(n1114) );
  AND U1321 ( .A(n1117), .B(n1118), .Z(n101) );
  NAND U1322 ( .A(B[53]), .B(n1119), .Z(n1118) );
  NANDN U1323 ( .A(A[53]), .B(n103), .Z(n1119) );
  NANDN U1324 ( .A(n103), .B(A[53]), .Z(n1117) );
  AND U1325 ( .A(n1120), .B(n1121), .Z(n103) );
  NAND U1326 ( .A(B[52]), .B(n1122), .Z(n1121) );
  NANDN U1327 ( .A(A[52]), .B(n105), .Z(n1122) );
  NANDN U1328 ( .A(n105), .B(A[52]), .Z(n1120) );
  AND U1329 ( .A(n1123), .B(n1124), .Z(n105) );
  NAND U1330 ( .A(B[51]), .B(n1125), .Z(n1124) );
  NANDN U1331 ( .A(A[51]), .B(n107), .Z(n1125) );
  NANDN U1332 ( .A(n107), .B(A[51]), .Z(n1123) );
  AND U1333 ( .A(n1126), .B(n1127), .Z(n107) );
  NAND U1334 ( .A(B[50]), .B(n1128), .Z(n1127) );
  NANDN U1335 ( .A(A[50]), .B(n109), .Z(n1128) );
  NANDN U1336 ( .A(n109), .B(A[50]), .Z(n1126) );
  AND U1337 ( .A(n1129), .B(n1130), .Z(n109) );
  NAND U1338 ( .A(B[49]), .B(n1131), .Z(n1130) );
  NANDN U1339 ( .A(A[49]), .B(n113), .Z(n1131) );
  NANDN U1340 ( .A(n113), .B(A[49]), .Z(n1129) );
  AND U1341 ( .A(n1132), .B(n1133), .Z(n113) );
  NAND U1342 ( .A(B[48]), .B(n1134), .Z(n1133) );
  NANDN U1343 ( .A(A[48]), .B(n115), .Z(n1134) );
  NANDN U1344 ( .A(n115), .B(A[48]), .Z(n1132) );
  AND U1345 ( .A(n1135), .B(n1136), .Z(n115) );
  NAND U1346 ( .A(B[47]), .B(n1137), .Z(n1136) );
  NANDN U1347 ( .A(A[47]), .B(n117), .Z(n1137) );
  NANDN U1348 ( .A(n117), .B(A[47]), .Z(n1135) );
  AND U1349 ( .A(n1138), .B(n1139), .Z(n117) );
  NAND U1350 ( .A(B[46]), .B(n1140), .Z(n1139) );
  NANDN U1351 ( .A(A[46]), .B(n119), .Z(n1140) );
  NANDN U1352 ( .A(n119), .B(A[46]), .Z(n1138) );
  AND U1353 ( .A(n1141), .B(n1142), .Z(n119) );
  NAND U1354 ( .A(B[45]), .B(n1143), .Z(n1142) );
  NANDN U1355 ( .A(A[45]), .B(n121), .Z(n1143) );
  NANDN U1356 ( .A(n121), .B(A[45]), .Z(n1141) );
  AND U1357 ( .A(n1144), .B(n1145), .Z(n121) );
  NAND U1358 ( .A(B[44]), .B(n1146), .Z(n1145) );
  NANDN U1359 ( .A(A[44]), .B(n123), .Z(n1146) );
  NANDN U1360 ( .A(n123), .B(A[44]), .Z(n1144) );
  AND U1361 ( .A(n1147), .B(n1148), .Z(n123) );
  NAND U1362 ( .A(B[43]), .B(n1149), .Z(n1148) );
  NANDN U1363 ( .A(A[43]), .B(n125), .Z(n1149) );
  NANDN U1364 ( .A(n125), .B(A[43]), .Z(n1147) );
  AND U1365 ( .A(n1150), .B(n1151), .Z(n125) );
  NAND U1366 ( .A(B[42]), .B(n1152), .Z(n1151) );
  NANDN U1367 ( .A(A[42]), .B(n127), .Z(n1152) );
  NANDN U1368 ( .A(n127), .B(A[42]), .Z(n1150) );
  AND U1369 ( .A(n1153), .B(n1154), .Z(n127) );
  NAND U1370 ( .A(B[41]), .B(n1155), .Z(n1154) );
  NANDN U1371 ( .A(A[41]), .B(n129), .Z(n1155) );
  NANDN U1372 ( .A(n129), .B(A[41]), .Z(n1153) );
  AND U1373 ( .A(n1156), .B(n1157), .Z(n129) );
  NAND U1374 ( .A(B[40]), .B(n1158), .Z(n1157) );
  NANDN U1375 ( .A(A[40]), .B(n131), .Z(n1158) );
  NANDN U1376 ( .A(n131), .B(A[40]), .Z(n1156) );
  AND U1377 ( .A(n1159), .B(n1160), .Z(n131) );
  NAND U1378 ( .A(B[39]), .B(n1161), .Z(n1160) );
  NANDN U1379 ( .A(A[39]), .B(n135), .Z(n1161) );
  NANDN U1380 ( .A(n135), .B(A[39]), .Z(n1159) );
  AND U1381 ( .A(n1162), .B(n1163), .Z(n135) );
  NAND U1382 ( .A(B[38]), .B(n1164), .Z(n1163) );
  NANDN U1383 ( .A(A[38]), .B(n137), .Z(n1164) );
  NANDN U1384 ( .A(n137), .B(A[38]), .Z(n1162) );
  AND U1385 ( .A(n1165), .B(n1166), .Z(n137) );
  NAND U1386 ( .A(B[37]), .B(n1167), .Z(n1166) );
  NANDN U1387 ( .A(A[37]), .B(n139), .Z(n1167) );
  NANDN U1388 ( .A(n139), .B(A[37]), .Z(n1165) );
  AND U1389 ( .A(n1168), .B(n1169), .Z(n139) );
  NAND U1390 ( .A(B[36]), .B(n1170), .Z(n1169) );
  NANDN U1391 ( .A(A[36]), .B(n141), .Z(n1170) );
  NANDN U1392 ( .A(n141), .B(A[36]), .Z(n1168) );
  AND U1393 ( .A(n1171), .B(n1172), .Z(n141) );
  NAND U1394 ( .A(B[35]), .B(n1173), .Z(n1172) );
  NANDN U1395 ( .A(A[35]), .B(n143), .Z(n1173) );
  NANDN U1396 ( .A(n143), .B(A[35]), .Z(n1171) );
  AND U1397 ( .A(n1174), .B(n1175), .Z(n143) );
  NAND U1398 ( .A(B[34]), .B(n1176), .Z(n1175) );
  NANDN U1399 ( .A(A[34]), .B(n145), .Z(n1176) );
  NANDN U1400 ( .A(n145), .B(A[34]), .Z(n1174) );
  AND U1401 ( .A(n1177), .B(n1178), .Z(n145) );
  NAND U1402 ( .A(B[33]), .B(n1179), .Z(n1178) );
  NANDN U1403 ( .A(A[33]), .B(n147), .Z(n1179) );
  NANDN U1404 ( .A(n147), .B(A[33]), .Z(n1177) );
  AND U1405 ( .A(n1180), .B(n1181), .Z(n147) );
  NAND U1406 ( .A(B[32]), .B(n1182), .Z(n1181) );
  NANDN U1407 ( .A(A[32]), .B(n149), .Z(n1182) );
  NANDN U1408 ( .A(n149), .B(A[32]), .Z(n1180) );
  AND U1409 ( .A(n1183), .B(n1184), .Z(n149) );
  NAND U1410 ( .A(B[31]), .B(n1185), .Z(n1184) );
  NANDN U1411 ( .A(A[31]), .B(n151), .Z(n1185) );
  NANDN U1412 ( .A(n151), .B(A[31]), .Z(n1183) );
  AND U1413 ( .A(n1186), .B(n1187), .Z(n151) );
  NAND U1414 ( .A(B[30]), .B(n1188), .Z(n1187) );
  NANDN U1415 ( .A(A[30]), .B(n153), .Z(n1188) );
  NANDN U1416 ( .A(n153), .B(A[30]), .Z(n1186) );
  AND U1417 ( .A(n1189), .B(n1190), .Z(n153) );
  NAND U1418 ( .A(B[29]), .B(n1191), .Z(n1190) );
  NANDN U1419 ( .A(A[29]), .B(n157), .Z(n1191) );
  NANDN U1420 ( .A(n157), .B(A[29]), .Z(n1189) );
  AND U1421 ( .A(n1192), .B(n1193), .Z(n157) );
  NAND U1422 ( .A(B[28]), .B(n1194), .Z(n1193) );
  NANDN U1423 ( .A(A[28]), .B(n159), .Z(n1194) );
  NANDN U1424 ( .A(n159), .B(A[28]), .Z(n1192) );
  AND U1425 ( .A(n1195), .B(n1196), .Z(n159) );
  NAND U1426 ( .A(B[27]), .B(n1197), .Z(n1196) );
  NANDN U1427 ( .A(A[27]), .B(n161), .Z(n1197) );
  NANDN U1428 ( .A(n161), .B(A[27]), .Z(n1195) );
  AND U1429 ( .A(n1198), .B(n1199), .Z(n161) );
  NAND U1430 ( .A(B[26]), .B(n1200), .Z(n1199) );
  NANDN U1431 ( .A(A[26]), .B(n163), .Z(n1200) );
  NANDN U1432 ( .A(n163), .B(A[26]), .Z(n1198) );
  AND U1433 ( .A(n1201), .B(n1202), .Z(n163) );
  NAND U1434 ( .A(B[25]), .B(n1203), .Z(n1202) );
  NANDN U1435 ( .A(A[25]), .B(n165), .Z(n1203) );
  NANDN U1436 ( .A(n165), .B(A[25]), .Z(n1201) );
  AND U1437 ( .A(n1204), .B(n1205), .Z(n165) );
  NAND U1438 ( .A(B[24]), .B(n1206), .Z(n1205) );
  NANDN U1439 ( .A(A[24]), .B(n203), .Z(n1206) );
  NANDN U1440 ( .A(n203), .B(A[24]), .Z(n1204) );
  AND U1441 ( .A(n1207), .B(n1208), .Z(n203) );
  NAND U1442 ( .A(B[23]), .B(n1209), .Z(n1208) );
  NANDN U1443 ( .A(A[23]), .B(n255), .Z(n1209) );
  NANDN U1444 ( .A(n255), .B(A[23]), .Z(n1207) );
  AND U1445 ( .A(n1210), .B(n1211), .Z(n255) );
  NAND U1446 ( .A(B[22]), .B(n1212), .Z(n1211) );
  NANDN U1447 ( .A(A[22]), .B(n307), .Z(n1212) );
  NANDN U1448 ( .A(n307), .B(A[22]), .Z(n1210) );
  AND U1449 ( .A(n1213), .B(n1214), .Z(n307) );
  NAND U1450 ( .A(B[21]), .B(n1215), .Z(n1214) );
  NANDN U1451 ( .A(A[21]), .B(n359), .Z(n1215) );
  NANDN U1452 ( .A(n359), .B(A[21]), .Z(n1213) );
  AND U1453 ( .A(n1216), .B(n1217), .Z(n359) );
  NAND U1454 ( .A(B[20]), .B(n1218), .Z(n1217) );
  NANDN U1455 ( .A(A[20]), .B(n411), .Z(n1218) );
  NANDN U1456 ( .A(n411), .B(A[20]), .Z(n1216) );
  AND U1457 ( .A(n1219), .B(n1220), .Z(n411) );
  NAND U1458 ( .A(B[19]), .B(n1221), .Z(n1220) );
  NANDN U1459 ( .A(A[19]), .B(n463), .Z(n1221) );
  NANDN U1460 ( .A(n463), .B(A[19]), .Z(n1219) );
  AND U1461 ( .A(n1222), .B(n1223), .Z(n463) );
  NAND U1462 ( .A(B[18]), .B(n1224), .Z(n1223) );
  NANDN U1463 ( .A(A[18]), .B(n515), .Z(n1224) );
  NANDN U1464 ( .A(n515), .B(A[18]), .Z(n1222) );
  AND U1465 ( .A(n1225), .B(n1226), .Z(n515) );
  NAND U1466 ( .A(B[17]), .B(n1227), .Z(n1226) );
  NANDN U1467 ( .A(A[17]), .B(n567), .Z(n1227) );
  NANDN U1468 ( .A(n567), .B(A[17]), .Z(n1225) );
  AND U1469 ( .A(n1228), .B(n1229), .Z(n567) );
  NAND U1470 ( .A(B[16]), .B(n1230), .Z(n1229) );
  NANDN U1471 ( .A(A[16]), .B(n619), .Z(n1230) );
  NANDN U1472 ( .A(n619), .B(A[16]), .Z(n1228) );
  AND U1473 ( .A(n1231), .B(n1232), .Z(n619) );
  NAND U1474 ( .A(B[15]), .B(n1233), .Z(n1232) );
  NANDN U1475 ( .A(A[15]), .B(n671), .Z(n1233) );
  NANDN U1476 ( .A(n671), .B(A[15]), .Z(n1231) );
  AND U1477 ( .A(n1234), .B(n1235), .Z(n671) );
  NAND U1478 ( .A(B[14]), .B(n1236), .Z(n1235) );
  NANDN U1479 ( .A(A[14]), .B(n723), .Z(n1236) );
  NANDN U1480 ( .A(n723), .B(A[14]), .Z(n1234) );
  AND U1481 ( .A(n1237), .B(n1238), .Z(n723) );
  NAND U1482 ( .A(B[13]), .B(n1239), .Z(n1238) );
  NANDN U1483 ( .A(A[13]), .B(n775), .Z(n1239) );
  NANDN U1484 ( .A(n775), .B(A[13]), .Z(n1237) );
  AND U1485 ( .A(n1240), .B(n1241), .Z(n775) );
  NAND U1486 ( .A(B[12]), .B(n1242), .Z(n1241) );
  NANDN U1487 ( .A(A[12]), .B(n827), .Z(n1242) );
  NANDN U1488 ( .A(n827), .B(A[12]), .Z(n1240) );
  AND U1489 ( .A(n1243), .B(n1244), .Z(n827) );
  NAND U1490 ( .A(B[11]), .B(n1245), .Z(n1244) );
  NANDN U1491 ( .A(A[11]), .B(n879), .Z(n1245) );
  NANDN U1492 ( .A(n879), .B(A[11]), .Z(n1243) );
  AND U1493 ( .A(n1246), .B(n1247), .Z(n879) );
  NAND U1494 ( .A(B[10]), .B(n1248), .Z(n1247) );
  NANDN U1495 ( .A(A[10]), .B(n931), .Z(n1248) );
  NANDN U1496 ( .A(n931), .B(A[10]), .Z(n1246) );
  AND U1497 ( .A(n1249), .B(n1250), .Z(n931) );
  NAND U1498 ( .A(B[9]), .B(n1251), .Z(n1250) );
  OR U1499 ( .A(n1), .B(A[9]), .Z(n1251) );
  NAND U1500 ( .A(A[9]), .B(n1), .Z(n1249) );
  NAND U1501 ( .A(n1252), .B(n1253), .Z(n1) );
  NAND U1502 ( .A(B[8]), .B(n1254), .Z(n1253) );
  NANDN U1503 ( .A(A[8]), .B(n23), .Z(n1254) );
  NANDN U1504 ( .A(n23), .B(A[8]), .Z(n1252) );
  AND U1505 ( .A(n1255), .B(n1256), .Z(n23) );
  NAND U1506 ( .A(B[7]), .B(n1257), .Z(n1256) );
  NANDN U1507 ( .A(A[7]), .B(n45), .Z(n1257) );
  NANDN U1508 ( .A(n45), .B(A[7]), .Z(n1255) );
  AND U1509 ( .A(n1258), .B(n1259), .Z(n45) );
  NAND U1510 ( .A(B[6]), .B(n1260), .Z(n1259) );
  NANDN U1511 ( .A(A[6]), .B(n67), .Z(n1260) );
  NANDN U1512 ( .A(n67), .B(A[6]), .Z(n1258) );
  AND U1513 ( .A(n1261), .B(n1262), .Z(n67) );
  NAND U1514 ( .A(B[5]), .B(n1263), .Z(n1262) );
  NANDN U1515 ( .A(A[5]), .B(n89), .Z(n1263) );
  NANDN U1516 ( .A(n89), .B(A[5]), .Z(n1261) );
  AND U1517 ( .A(n1264), .B(n1265), .Z(n89) );
  NAND U1518 ( .A(B[4]), .B(n1266), .Z(n1265) );
  NANDN U1519 ( .A(A[4]), .B(n111), .Z(n1266) );
  NANDN U1520 ( .A(n111), .B(A[4]), .Z(n1264) );
  AND U1521 ( .A(n1267), .B(n1268), .Z(n111) );
  NAND U1522 ( .A(B[3]), .B(n1269), .Z(n1268) );
  NANDN U1523 ( .A(A[3]), .B(n133), .Z(n1269) );
  NANDN U1524 ( .A(n133), .B(A[3]), .Z(n1267) );
  AND U1525 ( .A(n1270), .B(n1271), .Z(n133) );
  NAND U1526 ( .A(B[2]), .B(n1272), .Z(n1271) );
  OR U1527 ( .A(n155), .B(A[2]), .Z(n1272) );
  NAND U1528 ( .A(A[2]), .B(n155), .Z(n1270) );
  AND U1529 ( .A(B[1]), .B(A[1]), .Z(n155) );
endmodule


module modmult_step_N256_3 ( xregN_1, y, n, zin, zout );
  input [255:0] y;
  input [255:0] n;
  input [257:0] zin;
  output [257:0] zout;
  input xregN_1;
  wire   N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17, N18,
         N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31, N32,
         N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44, N45, N46,
         N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58, N59, N60,
         N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72, N73, N74,
         N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86, N87, N88,
         N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100, N101,
         N102, N103, N104, N105, N106, N107, N108, N109, N110, N111, N112,
         N113, N114, N115, N116, N117, N118, N119, N120, N121, N122, N123,
         N124, N125, N126, N127, N128, N129, N130, N131, N132, N133, N134,
         N135, N136, N137, N138, N139, N140, N141, N142, N143, N144, N145,
         N146, N147, N148, N149, N150, N151, N152, N153, N154, N155, N156,
         N157, N158, N159, N160, N161, N162, N163, N164, N165, N166, N167,
         N168, N169, N170, N171, N172, N173, N174, N175, N176, N177, N178,
         N179, N180, N181, N182, N183, N184, N185, N186, N187, N188, N189,
         N190, N191, N192, N193, N194, N195, N196, N197, N198, N199, N200,
         N201, N202, N203, N204, N205, N206, N207, N208, N209, N210, N211,
         N212, N213, N214, N215, N216, N217, N218, N219, N220, N221, N222,
         N223, N224, N225, N226, N227, N228, N229, N230, N231, N232, N233,
         N234, N235, N236, N237, N238, N239, N240, N241, N242, N243, N244,
         N245, N246, N247, N248, N249, N250, N251, N252, N253, N254, N255,
         N256, N257, N258, N259, N260, N261, N262, N264, N265, N266, N267,
         N268, N269, N270, N271, N272, N273, N274, N275, N276, N277, N278,
         N279, N280, N281, N282, N283, N284, N285, N286, N287, N288, N289,
         N290, N291, N292, N293, N294, N295, N296, N297, N298, N299, N300,
         N301, N302, N303, N304, N305, N306, N307, N308, N309, N310, N311,
         N312, N313, N314, N315, N316, N317, N318, N319, N320, N321, N322,
         N323, N324, N325, N326, N327, N328, N329, N330, N331, N332, N333,
         N334, N335, N336, N337, N338, N339, N340, N341, N342, N343, N344,
         N345, N346, N347, N348, N349, N350, N351, N352, N353, N354, N355,
         N356, N357, N358, N359, N360, N361, N362, N363, N364, N365, N366,
         N367, N368, N369, N370, N371, N372, N373, N374, N375, N376, N377,
         N378, N379, N380, N381, N382, N383, N384, N385, N386, N387, N388,
         N389, N390, N391, N392, N393, N394, N395, N396, N397, N398, N399,
         N400, N401, N402, N403, N404, N405, N406, N407, N408, N409, N410,
         N411, N412, N413, N414, N415, N416, N417, N418, N419, N420, N421,
         N422, N423, N424, N425, N426, N427, N428, N429, N430, N431, N432,
         N433, N434, N435, N436, N437, N438, N439, N440, N441, N442, N443,
         N444, N445, N446, N447, N448, N449, N450, N451, N452, N453, N454,
         N455, N456, N457, N458, N459, N460, N461, N462, N463, N464, N465,
         N466, N467, N468, N469, N470, N471, N472, N473, N474, N475, N476,
         N477, N478, N479, N480, N481, N482, N483, N484, N485, N486, N487,
         N488, N489, N490, N491, N492, N493, N494, N495, N496, N497, N498,
         N499, N500, N501, N502, N503, N504, N505, N506, N507, N508, N509,
         N510, N511, N512, N513, N514, N515, N516, N517, N518, N519, N520,
         N521, N780, N779, N778, N777, N776, N775, N774, N773, N772, N771,
         N770, N769, N768, N767, N766, N765, N764, N763, N762, N761, N760,
         N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, N749,
         N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738,
         N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727,
         N726, N725, N724, N723, N722, N721, N720, N719, N718, N717, N716,
         N715, N714, N713, N712, N711, N710, N709, N708, N707, N706, N705,
         N704, N703, N702, N701, N700, N699, N698, N697, N696, N695, N694,
         N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, N683,
         N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672,
         N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661,
         N660, N659, N658, N657, N656, N655, N654, N653, N652, N651, N650,
         N649, N648, N647, N646, N645, N644, N643, N642, N641, N640, N639,
         N638, N637, N636, N635, N634, N633, N632, N631, N630, N629, N628,
         N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, N617,
         N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606,
         N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595,
         N594, N593, N592, N591, N590, N589, N588, N587, N586, N585, N584,
         N583, N582, N581, N580, N579, N578, N577, N576, N575, N574, N573,
         N572, N571, N570, N569, N568, N567, N566, N565, N564, N563, N562,
         N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, N551,
         N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540,
         N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529,
         N528, N527, N526, N525, N522, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10,
         n11, n12, n13, n14, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101,
         n102, n103, n104, n105, n106, n107, n108, n109, n110, n111, n112,
         n113, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n138, n139, n140, n141, n142, n143, n144, n145,
         n146, n147, n148, n149, n150, n151, n152, n153, n154, n155, n156,
         n157, n158, n159, n160, n161, n162, n163, n164, n165, n166, n167,
         n168, n169, n170, n171, n172, n173, n174, n175, n176, n177, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n209, n210, n211,
         n212, n213, n214, n215, n216, n217, n218, n219, n220, n221, n222,
         n223, n224, n225, n226, n227, n228, n229, n230, n231, n232, n233,
         n234, n235, n236, n237, n238, n239, n240, n241, n242, n243, n244,
         n245, n246, n247, n248, n249, n250, n251, n252, n253, n254, n255,
         n256, n257, n258, n259, n260, n261, n262, n263, n264, n265, n266,
         n267, n268, n269, n270, n271, n272, n273, n274, n275, n276, n277,
         n278, n279, n280, n281, n282, n283, n284, n285, n286, n287, n288,
         n289, n290, n291, n292, n293, n294, n295, n296, n297, n298, n299,
         n300, n301, n302, n303, n304, n305, n306, n307, n308, n309, n310,
         n311, n312, n313, n314, n315, n316, n317, n318, n319, n320, n321,
         n322, n323, n324, n325, n326, n327, n328, n329, n330, n331, n332,
         n333, n334, n335, n336, n337, n338, n339, n340, n341, n342, n343,
         n344, n345, n346, n347, n348, n349, n350, n351, n352, n353, n354,
         n355, n356, n357, n358, n359, n360, n361, n362, n363, n364, n365,
         n366, n367, n368, n369, n370, n371, n372, n373, n374, n375, n376,
         n377, n378, n379, n380, n381, n382, n383, n384, n385, n386, n387,
         n388, n389, n390, n391, n392, n393, n394, n395, n396, n397, n398,
         n399, n400, n401, n402, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, n425, n426, n427, n428, n429, n430, n431,
         n432, n433, n434, n435, n436, n437, n438, n439, n440, n441, n442,
         n443, n444, n445, n446, n447, n448, n449, n450, n451, n452, n453,
         n454, n455, n456, n457, n458, n459, n460, n461, n462, n463, n464,
         n465, n466, n467, n468, n469, n470, n471, n472, n473, n474, n475,
         n476, n477, n478, n479, n480, n481, n482, n483, n484, n485, n486,
         n487, n488, n489, n490, n491, n492, n493, n494, n495, n496, n497,
         n498, n499, n500, n501, n502, n503, n504, n505, n506, n507, n508,
         n509, n510, n511, n512, n513, n514, n515, n516, n517, n518, n519,
         n520, n521, n522, n523, n524, n525, n526, n527, n528, n529, n530,
         n531, n532, n533, n534, n535, n536, n537, n538, n539, n540, n541,
         n542, n543, n544, n545, n546, n547, n548, n549, n550, n551, n552,
         n553, n554, n555, n556, n557, n558, n559, n560, n561, n562, n563,
         n564, n565, n566, n567, n568, n569, n570, n571, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n582, n583, n584, n585,
         n586, n587, n588, n589, n590, n591, n592, n593, n594, n595, n596,
         n597, n598, n599, n600, n601, n602, n603, n604, n605, n606, n607,
         n608, n609, n610, n611, n612, n613, n614, n615, n616, n617, n618,
         n619, n620, n621, n622, n623, n624, n625, n626, n627, n628, n629,
         n630, n631, n632, n633, n634, n635, n636, n637, n638, n639, n640,
         n641, n642, n643, n644, n645, n646, n647, n648, n649, n650, n651,
         n652, n653, n654, n655, n656, n657, n658, n659, n660, n661, n662,
         n663, n664, n665, n666, n667, n668, n669, n670, n671, n672, n673,
         n674, n675, n676, n677, n678, n679, n680, n681, n682, n683, n684,
         n685, n686, n687, n688, n689, n690, n691, n692, n693, n694, n695,
         n696, n697, n698, n699, n700, n701, n702, n703, n704, n705, n706,
         n707, n708, n709, n710, n711, n712, n713, n714, n715, n716, n717,
         n718, n719, n720, n721, n722, n723, n724, n725, n726, n727, n728,
         n729, n730, n731, n732, n733, n734, n735, n736, n737, n738, n739,
         n740, n741, n742, n743, n744, n745, n746, n747, n748, n749, n750,
         n751, n752, n753, n754, n755, n756, n757, n758, n759, n760, n761,
         n762, n763, n764, n765, n766, n767, n768, n769, n770, n771, n772,
         n773, n774, n775, n776, n777, n778, n779, n780, n781, n782, n783,
         n784, n785, n786, n787, n788, n789, n790, n791, n792, n793, n794,
         n795, n796, n797, n798, n799, n800, n801, n802, n803, n804, n805,
         n806, n807, n808, n809, n810, n811, n812, n813, n814, n815, n816,
         n817, n818, n819, n820, n821, n822, n823, n824, n825, n826, n827,
         n828, n829, n830, n831, n832, n833, n834, n835, n836, n837, n838,
         n839, n840, n841, n842, n843, n844, n845, n846, n847, n848, n849,
         n850, n851, n852, n853, n854, n855, n856, n857, n858, n859, n860,
         n861, n862, n863, n864, n865, n866, n867, n868, n869, n870, n871,
         n872, n873, n874, n875, n876, n877, n878, n879, n880, n881, n882,
         n883, n884, n885, n886, n887, n888, n889, n890, n891, n892, n893,
         n894, n895, n896, n897, n898, n899, n900, n901, n902, n903, n904,
         n905, n906, n907, n908, n909, n910, n911, n912, n913, n914, n915,
         n916, n917, n918, n919, n920, n921, n922, n923, n924, n925, n926,
         n927, n928, n929, n930, n931, n932, n933, n934, n935, n936, n937,
         n938, n939, n940, n941, n942, n943, n944, n945, n946, n947, n948,
         n949, n950, n951, n952, n953, n954, n955, n956, n957, n958, n959,
         n960, n961, n962, n963, n964, n965, n966, n967, n968, n969, n970,
         n971, n972, n973, n974, n975, n976, n977, n978, n979, n980, n981,
         n982, n983, n984, n985, n986, n987, n988, n989, n990, n991, n992,
         n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002, n1003,
         n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013,
         n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023,
         n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033,
         n1034, n1035, n1036, n1037, n1038, n1039;
  wire   [257:0] z2;
  wire   [257:0] z3;
  wire   SYNOPSYS_UNCONNECTED__0;

  modmult_step_N256_3_DW01_sub_0 sub_129_aco ( .A(z3), .B({1'b0, 1'b0, N780, 
        N779, N778, N777, N776, N775, N774, N773, N772, N771, N770, N769, N768, 
        N767, N766, N765, N764, N763, N762, N761, N760, N759, N758, N757, N756, 
        N755, N754, N753, N752, N751, N750, N749, N748, N747, N746, N745, N744, 
        N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, 
        N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, 
        N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, 
        N707, N706, N705, N704, N703, N702, N701, N700, N699, N698, N697, N696, 
        N695, N694, N693, N692, N691, N690, N689, N688, N687, N686, N685, N684, 
        N683, N682, N681, N680, N679, N678, N677, N676, N675, N674, N673, N672, 
        N671, N670, N669, N668, N667, N666, N665, N664, N663, N662, N661, N660, 
        N659, N658, N657, N656, N655, N654, N653, N652, N651, N650, N649, N648, 
        N647, N646, N645, N644, N643, N642, N641, N640, N639, N638, N637, N636, 
        N635, N634, N633, N632, N631, N630, N629, N628, N627, N626, N625, N624, 
        N623, N622, N621, N620, N619, N618, N617, N616, N615, N614, N613, N612, 
        N611, N610, N609, N608, N607, N606, N605, N604, N603, N602, N601, N600, 
        N599, N598, N597, N596, N595, N594, N593, N592, N591, N590, N589, N588, 
        N587, N586, N585, N584, N583, N582, N581, N580, N579, N578, N577, N576, 
        N575, N574, N573, N572, N571, N570, N569, N568, N567, N566, N565, N564, 
        N563, N562, N561, N560, N559, N558, N557, N556, N555, N554, N553, N552, 
        N551, N550, N549, N548, N547, N546, N545, N544, N543, N542, N541, N540, 
        N539, N538, N537, N536, N535, N534, N533, N532, N531, N530, N529, N528, 
        N527, N526, N525}), .CI(1'b0), .DIFF(zout) );
  modmult_step_N256_3_DW02_mult_0 mult_sub_129_aco ( .A(n), .B(N522), .TC(1'b0), .PRODUCT({SYNOPSYS_UNCONNECTED__0, N780, N779, N778, N777, N776, N775, N774, 
        N773, N772, N771, N770, N769, N768, N767, N766, N765, N764, N763, N762, 
        N761, N760, N759, N758, N757, N756, N755, N754, N753, N752, N751, N750, 
        N749, N748, N747, N746, N745, N744, N743, N742, N741, N740, N739, N738, 
        N737, N736, N735, N734, N733, N732, N731, N730, N729, N728, N727, N726, 
        N725, N724, N723, N722, N721, N720, N719, N718, N717, N716, N715, N714, 
        N713, N712, N711, N710, N709, N708, N707, N706, N705, N704, N703, N702, 
        N701, N700, N699, N698, N697, N696, N695, N694, N693, N692, N691, N690, 
        N689, N688, N687, N686, N685, N684, N683, N682, N681, N680, N679, N678, 
        N677, N676, N675, N674, N673, N672, N671, N670, N669, N668, N667, N666, 
        N665, N664, N663, N662, N661, N660, N659, N658, N657, N656, N655, N654, 
        N653, N652, N651, N650, N649, N648, N647, N646, N645, N644, N643, N642, 
        N641, N640, N639, N638, N637, N636, N635, N634, N633, N632, N631, N630, 
        N629, N628, N627, N626, N625, N624, N623, N622, N621, N620, N619, N618, 
        N617, N616, N615, N614, N613, N612, N611, N610, N609, N608, N607, N606, 
        N605, N604, N603, N602, N601, N600, N599, N598, N597, N596, N595, N594, 
        N593, N592, N591, N590, N589, N588, N587, N586, N585, N584, N583, N582, 
        N581, N580, N579, N578, N577, N576, N575, N574, N573, N572, N571, N570, 
        N569, N568, N567, N566, N565, N564, N563, N562, N561, N560, N559, N558, 
        N557, N556, N555, N554, N553, N552, N551, N550, N549, N548, N547, N546, 
        N545, N544, N543, N542, N541, N540, N539, N538, N537, N536, N535, N534, 
        N533, N532, N531, N530, N529, N528, N527, N526, N525}) );
  modmult_step_N256_3_DW01_cmp2_0 gte_128 ( .A({1'b0, 1'b0, n}), .B(z3), .LEQ(
        1'b1), .TC(1'b0), .LT_LE(N522) );
  modmult_step_N256_3_DW01_sub_1 sub_124 ( .A(z2), .B({1'b0, 1'b0, n}), .CI(
        1'b0), .DIFF({N521, N520, N519, N518, N517, N516, N515, N514, N513, 
        N512, N511, N510, N509, N508, N507, N506, N505, N504, N503, N502, N501, 
        N500, N499, N498, N497, N496, N495, N494, N493, N492, N491, N490, N489, 
        N488, N487, N486, N485, N484, N483, N482, N481, N480, N479, N478, N477, 
        N476, N475, N474, N473, N472, N471, N470, N469, N468, N467, N466, N465, 
        N464, N463, N462, N461, N460, N459, N458, N457, N456, N455, N454, N453, 
        N452, N451, N450, N449, N448, N447, N446, N445, N444, N443, N442, N441, 
        N440, N439, N438, N437, N436, N435, N434, N433, N432, N431, N430, N429, 
        N428, N427, N426, N425, N424, N423, N422, N421, N420, N419, N418, N417, 
        N416, N415, N414, N413, N412, N411, N410, N409, N408, N407, N406, N405, 
        N404, N403, N402, N401, N400, N399, N398, N397, N396, N395, N394, N393, 
        N392, N391, N390, N389, N388, N387, N386, N385, N384, N383, N382, N381, 
        N380, N379, N378, N377, N376, N375, N374, N373, N372, N371, N370, N369, 
        N368, N367, N366, N365, N364, N363, N362, N361, N360, N359, N358, N357, 
        N356, N355, N354, N353, N352, N351, N350, N349, N348, N347, N346, N345, 
        N344, N343, N342, N341, N340, N339, N338, N337, N336, N335, N334, N333, 
        N332, N331, N330, N329, N328, N327, N326, N325, N324, N323, N322, N321, 
        N320, N319, N318, N317, N316, N315, N314, N313, N312, N311, N310, N309, 
        N308, N307, N306, N305, N304, N303, N302, N301, N300, N299, N298, N297, 
        N296, N295, N294, N293, N292, N291, N290, N289, N288, N287, N286, N285, 
        N284, N283, N282, N281, N280, N279, N278, N277, N276, N275, N274, N273, 
        N272, N271, N270, N269, N268, N267, N266, N265, N264}) );
  modmult_step_N256_3_DW01_cmp2_1 gt_123 ( .A({1'b0, 1'b0, n}), .B(z2), .LEQ(
        1'b0), .TC(1'b0), .LT_LE(N262) );
  modmult_step_N256_3_DW01_add_0 add_119 ( .A({zin[256:0], 1'b0}), .B({1'b0, 
        1'b0, y}), .CI(1'b0), .SUM({N261, N260, N259, N258, N257, N256, N255, 
        N254, N253, N252, N251, N250, N249, N248, N247, N246, N245, N244, N243, 
        N242, N241, N240, N239, N238, N237, N236, N235, N234, N233, N232, N231, 
        N230, N229, N228, N227, N226, N225, N224, N223, N222, N221, N220, N219, 
        N218, N217, N216, N215, N214, N213, N212, N211, N210, N209, N208, N207, 
        N206, N205, N204, N203, N202, N201, N200, N199, N198, N197, N196, N195, 
        N194, N193, N192, N191, N190, N189, N188, N187, N186, N185, N184, N183, 
        N182, N181, N180, N179, N178, N177, N176, N175, N174, N173, N172, N171, 
        N170, N169, N168, N167, N166, N165, N164, N163, N162, N161, N160, N159, 
        N158, N157, N156, N155, N154, N153, N152, N151, N150, N149, N148, N147, 
        N146, N145, N144, N143, N142, N141, N140, N139, N138, N137, N136, N135, 
        N134, N133, N132, N131, N130, N129, N128, N127, N126, N125, N124, N123, 
        N122, N121, N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, 
        N110, N109, N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, 
        N98, N97, N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, 
        N84, N83, N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, 
        N70, N69, N68, N67, N66, N65, N64, N63, N62, N61, N60, N59, N58, N57, 
        N56, N55, N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, 
        N42, N41, N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, 
        N28, N27, N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, 
        N14, N13, N12, N11, N10, N9, N8, N7, N6, N5, N4}) );
  NAND U5 ( .A(n1), .B(n2), .Z(z3[9]) );
  NANDN U6 ( .A(N262), .B(z2[9]), .Z(n2) );
  NANDN U7 ( .A(n3), .B(N273), .Z(n1) );
  NAND U8 ( .A(n4), .B(n5), .Z(z3[99]) );
  NANDN U9 ( .A(N262), .B(z2[99]), .Z(n5) );
  NANDN U10 ( .A(n3), .B(N363), .Z(n4) );
  NAND U11 ( .A(n6), .B(n7), .Z(z3[98]) );
  NANDN U17 ( .A(N262), .B(z2[98]), .Z(n7) );
  NANDN U18 ( .A(n3), .B(N362), .Z(n6) );
  NAND U19 ( .A(n8), .B(n9), .Z(z3[97]) );
  NANDN U20 ( .A(N262), .B(z2[97]), .Z(n9) );
  NANDN U21 ( .A(n3), .B(N361), .Z(n8) );
  NAND U22 ( .A(n10), .B(n11), .Z(z3[96]) );
  NANDN U23 ( .A(N262), .B(z2[96]), .Z(n11) );
  NANDN U24 ( .A(n3), .B(N360), .Z(n10) );
  NAND U25 ( .A(n12), .B(n13), .Z(z3[95]) );
  NANDN U26 ( .A(N262), .B(z2[95]), .Z(n13) );
  NANDN U27 ( .A(n3), .B(N359), .Z(n12) );
  NAND U28 ( .A(n14), .B(n23), .Z(z3[94]) );
  NANDN U29 ( .A(N262), .B(z2[94]), .Z(n23) );
  NANDN U30 ( .A(n3), .B(N358), .Z(n14) );
  NAND U31 ( .A(n24), .B(n25), .Z(z3[93]) );
  NANDN U32 ( .A(N262), .B(z2[93]), .Z(n25) );
  NANDN U33 ( .A(n3), .B(N357), .Z(n24) );
  NAND U34 ( .A(n26), .B(n27), .Z(z3[92]) );
  NANDN U35 ( .A(N262), .B(z2[92]), .Z(n27) );
  NANDN U36 ( .A(n3), .B(N356), .Z(n26) );
  NAND U37 ( .A(n28), .B(n29), .Z(z3[91]) );
  NANDN U38 ( .A(N262), .B(z2[91]), .Z(n29) );
  NANDN U39 ( .A(n3), .B(N355), .Z(n28) );
  NAND U40 ( .A(n30), .B(n31), .Z(z3[90]) );
  NANDN U41 ( .A(N262), .B(z2[90]), .Z(n31) );
  NANDN U42 ( .A(n3), .B(N354), .Z(n30) );
  NAND U43 ( .A(n32), .B(n33), .Z(z3[8]) );
  NANDN U44 ( .A(N262), .B(z2[8]), .Z(n33) );
  NANDN U45 ( .A(n3), .B(N272), .Z(n32) );
  NAND U46 ( .A(n34), .B(n35), .Z(z3[89]) );
  NANDN U47 ( .A(N262), .B(z2[89]), .Z(n35) );
  NANDN U48 ( .A(n3), .B(N353), .Z(n34) );
  NAND U49 ( .A(n36), .B(n37), .Z(z3[88]) );
  NANDN U50 ( .A(N262), .B(z2[88]), .Z(n37) );
  NANDN U51 ( .A(n3), .B(N352), .Z(n36) );
  NAND U52 ( .A(n38), .B(n39), .Z(z3[87]) );
  NANDN U53 ( .A(N262), .B(z2[87]), .Z(n39) );
  NANDN U54 ( .A(n3), .B(N351), .Z(n38) );
  NAND U55 ( .A(n40), .B(n41), .Z(z3[86]) );
  NANDN U56 ( .A(N262), .B(z2[86]), .Z(n41) );
  NANDN U57 ( .A(n3), .B(N350), .Z(n40) );
  NAND U58 ( .A(n42), .B(n43), .Z(z3[85]) );
  NANDN U59 ( .A(N262), .B(z2[85]), .Z(n43) );
  NANDN U60 ( .A(n3), .B(N349), .Z(n42) );
  NAND U61 ( .A(n44), .B(n45), .Z(z3[84]) );
  NANDN U62 ( .A(N262), .B(z2[84]), .Z(n45) );
  NANDN U63 ( .A(n3), .B(N348), .Z(n44) );
  NAND U64 ( .A(n46), .B(n47), .Z(z3[83]) );
  NANDN U65 ( .A(N262), .B(z2[83]), .Z(n47) );
  NANDN U66 ( .A(n3), .B(N347), .Z(n46) );
  NAND U67 ( .A(n48), .B(n49), .Z(z3[82]) );
  NANDN U68 ( .A(N262), .B(z2[82]), .Z(n49) );
  NANDN U69 ( .A(n3), .B(N346), .Z(n48) );
  NAND U70 ( .A(n50), .B(n51), .Z(z3[81]) );
  NANDN U71 ( .A(N262), .B(z2[81]), .Z(n51) );
  NANDN U72 ( .A(n3), .B(N345), .Z(n50) );
  NAND U73 ( .A(n52), .B(n53), .Z(z3[80]) );
  NANDN U74 ( .A(N262), .B(z2[80]), .Z(n53) );
  NANDN U75 ( .A(n3), .B(N344), .Z(n52) );
  NAND U76 ( .A(n54), .B(n55), .Z(z3[7]) );
  NANDN U77 ( .A(N262), .B(z2[7]), .Z(n55) );
  NANDN U78 ( .A(n3), .B(N271), .Z(n54) );
  NAND U79 ( .A(n56), .B(n57), .Z(z3[79]) );
  NANDN U80 ( .A(N262), .B(z2[79]), .Z(n57) );
  NANDN U81 ( .A(n3), .B(N343), .Z(n56) );
  NAND U82 ( .A(n58), .B(n59), .Z(z3[78]) );
  NANDN U83 ( .A(N262), .B(z2[78]), .Z(n59) );
  NANDN U84 ( .A(n3), .B(N342), .Z(n58) );
  NAND U85 ( .A(n60), .B(n61), .Z(z3[77]) );
  NANDN U86 ( .A(N262), .B(z2[77]), .Z(n61) );
  NANDN U87 ( .A(n3), .B(N341), .Z(n60) );
  NAND U88 ( .A(n62), .B(n63), .Z(z3[76]) );
  NANDN U89 ( .A(N262), .B(z2[76]), .Z(n63) );
  NANDN U90 ( .A(n3), .B(N340), .Z(n62) );
  NAND U91 ( .A(n64), .B(n65), .Z(z3[75]) );
  NANDN U92 ( .A(N262), .B(z2[75]), .Z(n65) );
  NANDN U93 ( .A(n3), .B(N339), .Z(n64) );
  NAND U94 ( .A(n66), .B(n67), .Z(z3[74]) );
  NANDN U95 ( .A(N262), .B(z2[74]), .Z(n67) );
  NANDN U96 ( .A(n3), .B(N338), .Z(n66) );
  NAND U97 ( .A(n68), .B(n69), .Z(z3[73]) );
  NANDN U98 ( .A(N262), .B(z2[73]), .Z(n69) );
  NANDN U99 ( .A(n3), .B(N337), .Z(n68) );
  NAND U100 ( .A(n70), .B(n71), .Z(z3[72]) );
  NANDN U101 ( .A(N262), .B(z2[72]), .Z(n71) );
  NANDN U102 ( .A(n3), .B(N336), .Z(n70) );
  NAND U103 ( .A(n72), .B(n73), .Z(z3[71]) );
  NANDN U104 ( .A(N262), .B(z2[71]), .Z(n73) );
  NANDN U105 ( .A(n3), .B(N335), .Z(n72) );
  NAND U106 ( .A(n74), .B(n75), .Z(z3[70]) );
  NANDN U107 ( .A(N262), .B(z2[70]), .Z(n75) );
  NANDN U108 ( .A(n3), .B(N334), .Z(n74) );
  NAND U109 ( .A(n76), .B(n77), .Z(z3[6]) );
  NANDN U110 ( .A(N262), .B(z2[6]), .Z(n77) );
  NANDN U111 ( .A(n3), .B(N270), .Z(n76) );
  NAND U112 ( .A(n78), .B(n79), .Z(z3[69]) );
  NANDN U113 ( .A(N262), .B(z2[69]), .Z(n79) );
  NANDN U114 ( .A(n3), .B(N333), .Z(n78) );
  NAND U115 ( .A(n80), .B(n81), .Z(z3[68]) );
  NANDN U116 ( .A(N262), .B(z2[68]), .Z(n81) );
  NANDN U117 ( .A(n3), .B(N332), .Z(n80) );
  NAND U118 ( .A(n82), .B(n83), .Z(z3[67]) );
  NANDN U119 ( .A(N262), .B(z2[67]), .Z(n83) );
  NANDN U120 ( .A(n3), .B(N331), .Z(n82) );
  NAND U121 ( .A(n84), .B(n85), .Z(z3[66]) );
  NANDN U122 ( .A(N262), .B(z2[66]), .Z(n85) );
  NANDN U123 ( .A(n3), .B(N330), .Z(n84) );
  NAND U124 ( .A(n86), .B(n87), .Z(z3[65]) );
  NANDN U125 ( .A(N262), .B(z2[65]), .Z(n87) );
  NANDN U126 ( .A(n3), .B(N329), .Z(n86) );
  NAND U127 ( .A(n88), .B(n89), .Z(z3[64]) );
  NANDN U128 ( .A(N262), .B(z2[64]), .Z(n89) );
  NANDN U129 ( .A(n3), .B(N328), .Z(n88) );
  NAND U130 ( .A(n90), .B(n91), .Z(z3[63]) );
  NANDN U131 ( .A(N262), .B(z2[63]), .Z(n91) );
  NANDN U132 ( .A(n3), .B(N327), .Z(n90) );
  NAND U133 ( .A(n92), .B(n93), .Z(z3[62]) );
  NANDN U134 ( .A(N262), .B(z2[62]), .Z(n93) );
  NANDN U135 ( .A(n3), .B(N326), .Z(n92) );
  NAND U136 ( .A(n94), .B(n95), .Z(z3[61]) );
  NANDN U137 ( .A(N262), .B(z2[61]), .Z(n95) );
  NANDN U138 ( .A(n3), .B(N325), .Z(n94) );
  NAND U139 ( .A(n96), .B(n97), .Z(z3[60]) );
  NANDN U140 ( .A(N262), .B(z2[60]), .Z(n97) );
  NANDN U141 ( .A(n3), .B(N324), .Z(n96) );
  NAND U142 ( .A(n98), .B(n99), .Z(z3[5]) );
  NANDN U143 ( .A(N262), .B(z2[5]), .Z(n99) );
  NANDN U144 ( .A(n3), .B(N269), .Z(n98) );
  NAND U145 ( .A(n100), .B(n101), .Z(z3[59]) );
  NANDN U146 ( .A(N262), .B(z2[59]), .Z(n101) );
  NANDN U147 ( .A(n3), .B(N323), .Z(n100) );
  NAND U148 ( .A(n102), .B(n103), .Z(z3[58]) );
  NANDN U149 ( .A(N262), .B(z2[58]), .Z(n103) );
  NANDN U150 ( .A(n3), .B(N322), .Z(n102) );
  NAND U151 ( .A(n104), .B(n105), .Z(z3[57]) );
  NANDN U152 ( .A(N262), .B(z2[57]), .Z(n105) );
  NANDN U153 ( .A(n3), .B(N321), .Z(n104) );
  NAND U154 ( .A(n106), .B(n107), .Z(z3[56]) );
  NANDN U155 ( .A(N262), .B(z2[56]), .Z(n107) );
  NANDN U156 ( .A(n3), .B(N320), .Z(n106) );
  NAND U157 ( .A(n108), .B(n109), .Z(z3[55]) );
  NANDN U158 ( .A(N262), .B(z2[55]), .Z(n109) );
  NANDN U159 ( .A(n3), .B(N319), .Z(n108) );
  NAND U160 ( .A(n110), .B(n111), .Z(z3[54]) );
  NANDN U161 ( .A(N262), .B(z2[54]), .Z(n111) );
  NANDN U162 ( .A(n3), .B(N318), .Z(n110) );
  NAND U163 ( .A(n112), .B(n113), .Z(z3[53]) );
  NANDN U164 ( .A(N262), .B(z2[53]), .Z(n113) );
  NANDN U165 ( .A(n3), .B(N317), .Z(n112) );
  NAND U166 ( .A(n114), .B(n115), .Z(z3[52]) );
  NANDN U167 ( .A(N262), .B(z2[52]), .Z(n115) );
  NANDN U168 ( .A(n3), .B(N316), .Z(n114) );
  NAND U169 ( .A(n116), .B(n117), .Z(z3[51]) );
  NANDN U170 ( .A(N262), .B(z2[51]), .Z(n117) );
  NANDN U171 ( .A(n3), .B(N315), .Z(n116) );
  NAND U172 ( .A(n118), .B(n119), .Z(z3[50]) );
  NANDN U173 ( .A(N262), .B(z2[50]), .Z(n119) );
  NANDN U174 ( .A(n3), .B(N314), .Z(n118) );
  NAND U175 ( .A(n120), .B(n121), .Z(z3[4]) );
  NANDN U176 ( .A(N262), .B(z2[4]), .Z(n121) );
  NANDN U177 ( .A(n3), .B(N268), .Z(n120) );
  NAND U178 ( .A(n122), .B(n123), .Z(z3[49]) );
  NANDN U179 ( .A(N262), .B(z2[49]), .Z(n123) );
  NANDN U180 ( .A(n3), .B(N313), .Z(n122) );
  NAND U181 ( .A(n124), .B(n125), .Z(z3[48]) );
  NANDN U182 ( .A(N262), .B(z2[48]), .Z(n125) );
  NANDN U183 ( .A(n3), .B(N312), .Z(n124) );
  NAND U184 ( .A(n126), .B(n127), .Z(z3[47]) );
  NANDN U185 ( .A(N262), .B(z2[47]), .Z(n127) );
  NANDN U186 ( .A(n3), .B(N311), .Z(n126) );
  NAND U187 ( .A(n128), .B(n129), .Z(z3[46]) );
  NANDN U188 ( .A(N262), .B(z2[46]), .Z(n129) );
  NANDN U189 ( .A(n3), .B(N310), .Z(n128) );
  NAND U190 ( .A(n130), .B(n131), .Z(z3[45]) );
  NANDN U191 ( .A(N262), .B(z2[45]), .Z(n131) );
  NANDN U192 ( .A(n3), .B(N309), .Z(n130) );
  NAND U193 ( .A(n132), .B(n133), .Z(z3[44]) );
  NANDN U194 ( .A(N262), .B(z2[44]), .Z(n133) );
  NANDN U195 ( .A(n3), .B(N308), .Z(n132) );
  NAND U196 ( .A(n134), .B(n135), .Z(z3[43]) );
  NANDN U197 ( .A(N262), .B(z2[43]), .Z(n135) );
  NANDN U198 ( .A(n3), .B(N307), .Z(n134) );
  NAND U199 ( .A(n136), .B(n137), .Z(z3[42]) );
  NANDN U200 ( .A(N262), .B(z2[42]), .Z(n137) );
  NANDN U201 ( .A(n3), .B(N306), .Z(n136) );
  NAND U202 ( .A(n138), .B(n139), .Z(z3[41]) );
  NANDN U203 ( .A(N262), .B(z2[41]), .Z(n139) );
  NANDN U204 ( .A(n3), .B(N305), .Z(n138) );
  NAND U205 ( .A(n140), .B(n141), .Z(z3[40]) );
  NANDN U206 ( .A(N262), .B(z2[40]), .Z(n141) );
  NANDN U207 ( .A(n3), .B(N304), .Z(n140) );
  NAND U208 ( .A(n142), .B(n143), .Z(z3[3]) );
  NANDN U209 ( .A(N262), .B(z2[3]), .Z(n143) );
  NANDN U210 ( .A(n3), .B(N267), .Z(n142) );
  NAND U211 ( .A(n144), .B(n145), .Z(z3[39]) );
  NANDN U212 ( .A(N262), .B(z2[39]), .Z(n145) );
  NANDN U213 ( .A(n3), .B(N303), .Z(n144) );
  NAND U214 ( .A(n146), .B(n147), .Z(z3[38]) );
  NANDN U215 ( .A(N262), .B(z2[38]), .Z(n147) );
  NANDN U216 ( .A(n3), .B(N302), .Z(n146) );
  NAND U217 ( .A(n148), .B(n149), .Z(z3[37]) );
  NANDN U218 ( .A(N262), .B(z2[37]), .Z(n149) );
  NANDN U219 ( .A(n3), .B(N301), .Z(n148) );
  NAND U220 ( .A(n150), .B(n151), .Z(z3[36]) );
  NANDN U221 ( .A(N262), .B(z2[36]), .Z(n151) );
  NANDN U222 ( .A(n3), .B(N300), .Z(n150) );
  NAND U223 ( .A(n152), .B(n153), .Z(z3[35]) );
  NANDN U224 ( .A(N262), .B(z2[35]), .Z(n153) );
  NANDN U225 ( .A(n3), .B(N299), .Z(n152) );
  NAND U226 ( .A(n154), .B(n155), .Z(z3[34]) );
  NANDN U227 ( .A(N262), .B(z2[34]), .Z(n155) );
  NANDN U228 ( .A(n3), .B(N298), .Z(n154) );
  NAND U229 ( .A(n156), .B(n157), .Z(z3[33]) );
  NANDN U230 ( .A(N262), .B(z2[33]), .Z(n157) );
  NANDN U231 ( .A(n3), .B(N297), .Z(n156) );
  NAND U232 ( .A(n158), .B(n159), .Z(z3[32]) );
  NANDN U233 ( .A(N262), .B(z2[32]), .Z(n159) );
  NANDN U234 ( .A(n3), .B(N296), .Z(n158) );
  NAND U235 ( .A(n160), .B(n161), .Z(z3[31]) );
  NANDN U236 ( .A(N262), .B(z2[31]), .Z(n161) );
  NANDN U237 ( .A(n3), .B(N295), .Z(n160) );
  NAND U238 ( .A(n162), .B(n163), .Z(z3[30]) );
  NANDN U239 ( .A(N262), .B(z2[30]), .Z(n163) );
  NANDN U240 ( .A(n3), .B(N294), .Z(n162) );
  NAND U241 ( .A(n164), .B(n165), .Z(z3[2]) );
  NANDN U242 ( .A(N262), .B(z2[2]), .Z(n165) );
  NANDN U243 ( .A(n3), .B(N266), .Z(n164) );
  NAND U244 ( .A(n166), .B(n167), .Z(z3[29]) );
  NANDN U245 ( .A(N262), .B(z2[29]), .Z(n167) );
  NANDN U246 ( .A(n3), .B(N293), .Z(n166) );
  NAND U247 ( .A(n168), .B(n169), .Z(z3[28]) );
  NANDN U248 ( .A(N262), .B(z2[28]), .Z(n169) );
  NANDN U249 ( .A(n3), .B(N292), .Z(n168) );
  NAND U250 ( .A(n170), .B(n171), .Z(z3[27]) );
  NANDN U251 ( .A(N262), .B(z2[27]), .Z(n171) );
  NANDN U252 ( .A(n3), .B(N291), .Z(n170) );
  NAND U253 ( .A(n172), .B(n173), .Z(z3[26]) );
  NANDN U254 ( .A(N262), .B(z2[26]), .Z(n173) );
  NANDN U255 ( .A(n3), .B(N290), .Z(n172) );
  NAND U256 ( .A(n174), .B(n175), .Z(z3[25]) );
  NANDN U257 ( .A(N262), .B(z2[25]), .Z(n175) );
  NANDN U258 ( .A(n3), .B(N289), .Z(n174) );
  NAND U259 ( .A(n176), .B(n177), .Z(z3[257]) );
  NANDN U260 ( .A(N262), .B(z2[257]), .Z(n177) );
  NANDN U261 ( .A(n3), .B(N521), .Z(n176) );
  NAND U262 ( .A(n178), .B(n179), .Z(z3[256]) );
  NANDN U263 ( .A(N262), .B(z2[256]), .Z(n179) );
  NANDN U264 ( .A(n3), .B(N520), .Z(n178) );
  NAND U265 ( .A(n180), .B(n181), .Z(z3[255]) );
  NANDN U266 ( .A(N262), .B(z2[255]), .Z(n181) );
  NANDN U267 ( .A(n3), .B(N519), .Z(n180) );
  NAND U268 ( .A(n182), .B(n183), .Z(z3[254]) );
  NANDN U269 ( .A(N262), .B(z2[254]), .Z(n183) );
  NANDN U270 ( .A(n3), .B(N518), .Z(n182) );
  NAND U271 ( .A(n184), .B(n185), .Z(z3[253]) );
  NANDN U272 ( .A(N262), .B(z2[253]), .Z(n185) );
  NANDN U273 ( .A(n3), .B(N517), .Z(n184) );
  NAND U274 ( .A(n186), .B(n187), .Z(z3[252]) );
  NANDN U275 ( .A(N262), .B(z2[252]), .Z(n187) );
  NANDN U276 ( .A(n3), .B(N516), .Z(n186) );
  NAND U277 ( .A(n188), .B(n189), .Z(z3[251]) );
  NANDN U278 ( .A(N262), .B(z2[251]), .Z(n189) );
  NANDN U279 ( .A(n3), .B(N515), .Z(n188) );
  NAND U280 ( .A(n190), .B(n191), .Z(z3[250]) );
  NANDN U281 ( .A(N262), .B(z2[250]), .Z(n191) );
  NANDN U282 ( .A(n3), .B(N514), .Z(n190) );
  NAND U283 ( .A(n192), .B(n193), .Z(z3[24]) );
  NANDN U284 ( .A(N262), .B(z2[24]), .Z(n193) );
  NANDN U285 ( .A(n3), .B(N288), .Z(n192) );
  NAND U286 ( .A(n194), .B(n195), .Z(z3[249]) );
  NANDN U287 ( .A(N262), .B(z2[249]), .Z(n195) );
  NANDN U288 ( .A(n3), .B(N513), .Z(n194) );
  NAND U289 ( .A(n196), .B(n197), .Z(z3[248]) );
  NANDN U290 ( .A(N262), .B(z2[248]), .Z(n197) );
  NANDN U291 ( .A(n3), .B(N512), .Z(n196) );
  NAND U292 ( .A(n198), .B(n199), .Z(z3[247]) );
  NANDN U293 ( .A(N262), .B(z2[247]), .Z(n199) );
  NANDN U294 ( .A(n3), .B(N511), .Z(n198) );
  NAND U295 ( .A(n200), .B(n201), .Z(z3[246]) );
  NANDN U296 ( .A(N262), .B(z2[246]), .Z(n201) );
  NANDN U297 ( .A(n3), .B(N510), .Z(n200) );
  NAND U298 ( .A(n202), .B(n203), .Z(z3[245]) );
  NANDN U299 ( .A(N262), .B(z2[245]), .Z(n203) );
  NANDN U300 ( .A(n3), .B(N509), .Z(n202) );
  NAND U301 ( .A(n204), .B(n205), .Z(z3[244]) );
  NANDN U302 ( .A(N262), .B(z2[244]), .Z(n205) );
  NANDN U303 ( .A(n3), .B(N508), .Z(n204) );
  NAND U304 ( .A(n206), .B(n207), .Z(z3[243]) );
  NANDN U305 ( .A(N262), .B(z2[243]), .Z(n207) );
  NANDN U306 ( .A(n3), .B(N507), .Z(n206) );
  NAND U307 ( .A(n208), .B(n209), .Z(z3[242]) );
  NANDN U308 ( .A(N262), .B(z2[242]), .Z(n209) );
  NANDN U309 ( .A(n3), .B(N506), .Z(n208) );
  NAND U310 ( .A(n210), .B(n211), .Z(z3[241]) );
  NANDN U311 ( .A(N262), .B(z2[241]), .Z(n211) );
  NANDN U312 ( .A(n3), .B(N505), .Z(n210) );
  NAND U313 ( .A(n212), .B(n213), .Z(z3[240]) );
  NANDN U314 ( .A(N262), .B(z2[240]), .Z(n213) );
  NANDN U315 ( .A(n3), .B(N504), .Z(n212) );
  NAND U316 ( .A(n214), .B(n215), .Z(z3[23]) );
  NANDN U317 ( .A(N262), .B(z2[23]), .Z(n215) );
  NANDN U318 ( .A(n3), .B(N287), .Z(n214) );
  NAND U319 ( .A(n216), .B(n217), .Z(z3[239]) );
  NANDN U320 ( .A(N262), .B(z2[239]), .Z(n217) );
  NANDN U321 ( .A(n3), .B(N503), .Z(n216) );
  NAND U322 ( .A(n218), .B(n219), .Z(z3[238]) );
  NANDN U323 ( .A(N262), .B(z2[238]), .Z(n219) );
  NANDN U324 ( .A(n3), .B(N502), .Z(n218) );
  NAND U325 ( .A(n220), .B(n221), .Z(z3[237]) );
  NANDN U326 ( .A(N262), .B(z2[237]), .Z(n221) );
  NANDN U327 ( .A(n3), .B(N501), .Z(n220) );
  NAND U328 ( .A(n222), .B(n223), .Z(z3[236]) );
  NANDN U329 ( .A(N262), .B(z2[236]), .Z(n223) );
  NANDN U330 ( .A(n3), .B(N500), .Z(n222) );
  NAND U331 ( .A(n224), .B(n225), .Z(z3[235]) );
  NANDN U332 ( .A(N262), .B(z2[235]), .Z(n225) );
  NANDN U333 ( .A(n3), .B(N499), .Z(n224) );
  NAND U334 ( .A(n226), .B(n227), .Z(z3[234]) );
  NANDN U335 ( .A(N262), .B(z2[234]), .Z(n227) );
  NANDN U336 ( .A(n3), .B(N498), .Z(n226) );
  NAND U337 ( .A(n228), .B(n229), .Z(z3[233]) );
  NANDN U338 ( .A(N262), .B(z2[233]), .Z(n229) );
  NANDN U339 ( .A(n3), .B(N497), .Z(n228) );
  NAND U340 ( .A(n230), .B(n231), .Z(z3[232]) );
  NANDN U341 ( .A(N262), .B(z2[232]), .Z(n231) );
  NANDN U342 ( .A(n3), .B(N496), .Z(n230) );
  NAND U343 ( .A(n232), .B(n233), .Z(z3[231]) );
  NANDN U344 ( .A(N262), .B(z2[231]), .Z(n233) );
  NANDN U345 ( .A(n3), .B(N495), .Z(n232) );
  NAND U346 ( .A(n234), .B(n235), .Z(z3[230]) );
  NANDN U347 ( .A(N262), .B(z2[230]), .Z(n235) );
  NANDN U348 ( .A(n3), .B(N494), .Z(n234) );
  NAND U349 ( .A(n236), .B(n237), .Z(z3[22]) );
  NANDN U350 ( .A(N262), .B(z2[22]), .Z(n237) );
  NANDN U351 ( .A(n3), .B(N286), .Z(n236) );
  NAND U352 ( .A(n238), .B(n239), .Z(z3[229]) );
  NANDN U353 ( .A(N262), .B(z2[229]), .Z(n239) );
  NANDN U354 ( .A(n3), .B(N493), .Z(n238) );
  NAND U355 ( .A(n240), .B(n241), .Z(z3[228]) );
  NANDN U356 ( .A(N262), .B(z2[228]), .Z(n241) );
  NANDN U357 ( .A(n3), .B(N492), .Z(n240) );
  NAND U358 ( .A(n242), .B(n243), .Z(z3[227]) );
  NANDN U359 ( .A(N262), .B(z2[227]), .Z(n243) );
  NANDN U360 ( .A(n3), .B(N491), .Z(n242) );
  NAND U361 ( .A(n244), .B(n245), .Z(z3[226]) );
  NANDN U362 ( .A(N262), .B(z2[226]), .Z(n245) );
  NANDN U363 ( .A(n3), .B(N490), .Z(n244) );
  NAND U364 ( .A(n246), .B(n247), .Z(z3[225]) );
  NANDN U365 ( .A(N262), .B(z2[225]), .Z(n247) );
  NANDN U366 ( .A(n3), .B(N489), .Z(n246) );
  NAND U367 ( .A(n248), .B(n249), .Z(z3[224]) );
  NANDN U368 ( .A(N262), .B(z2[224]), .Z(n249) );
  NANDN U369 ( .A(n3), .B(N488), .Z(n248) );
  NAND U370 ( .A(n250), .B(n251), .Z(z3[223]) );
  NANDN U371 ( .A(N262), .B(z2[223]), .Z(n251) );
  NANDN U372 ( .A(n3), .B(N487), .Z(n250) );
  NAND U373 ( .A(n252), .B(n253), .Z(z3[222]) );
  NANDN U374 ( .A(N262), .B(z2[222]), .Z(n253) );
  NANDN U375 ( .A(n3), .B(N486), .Z(n252) );
  NAND U376 ( .A(n254), .B(n255), .Z(z3[221]) );
  NANDN U377 ( .A(N262), .B(z2[221]), .Z(n255) );
  NANDN U378 ( .A(n3), .B(N485), .Z(n254) );
  NAND U379 ( .A(n256), .B(n257), .Z(z3[220]) );
  NANDN U380 ( .A(N262), .B(z2[220]), .Z(n257) );
  NANDN U381 ( .A(n3), .B(N484), .Z(n256) );
  NAND U382 ( .A(n258), .B(n259), .Z(z3[21]) );
  NANDN U383 ( .A(N262), .B(z2[21]), .Z(n259) );
  NANDN U384 ( .A(n3), .B(N285), .Z(n258) );
  NAND U385 ( .A(n260), .B(n261), .Z(z3[219]) );
  NANDN U386 ( .A(N262), .B(z2[219]), .Z(n261) );
  NANDN U387 ( .A(n3), .B(N483), .Z(n260) );
  NAND U388 ( .A(n262), .B(n263), .Z(z3[218]) );
  NANDN U389 ( .A(N262), .B(z2[218]), .Z(n263) );
  NANDN U390 ( .A(n3), .B(N482), .Z(n262) );
  NAND U391 ( .A(n264), .B(n265), .Z(z3[217]) );
  NANDN U392 ( .A(N262), .B(z2[217]), .Z(n265) );
  NANDN U393 ( .A(n3), .B(N481), .Z(n264) );
  NAND U394 ( .A(n266), .B(n267), .Z(z3[216]) );
  NANDN U395 ( .A(N262), .B(z2[216]), .Z(n267) );
  NANDN U396 ( .A(n3), .B(N480), .Z(n266) );
  NAND U397 ( .A(n268), .B(n269), .Z(z3[215]) );
  NANDN U398 ( .A(N262), .B(z2[215]), .Z(n269) );
  NANDN U399 ( .A(n3), .B(N479), .Z(n268) );
  NAND U400 ( .A(n270), .B(n271), .Z(z3[214]) );
  NANDN U401 ( .A(N262), .B(z2[214]), .Z(n271) );
  NANDN U402 ( .A(n3), .B(N478), .Z(n270) );
  NAND U403 ( .A(n272), .B(n273), .Z(z3[213]) );
  NANDN U404 ( .A(N262), .B(z2[213]), .Z(n273) );
  NANDN U405 ( .A(n3), .B(N477), .Z(n272) );
  NAND U406 ( .A(n274), .B(n275), .Z(z3[212]) );
  NANDN U407 ( .A(N262), .B(z2[212]), .Z(n275) );
  NANDN U408 ( .A(n3), .B(N476), .Z(n274) );
  NAND U409 ( .A(n276), .B(n277), .Z(z3[211]) );
  NANDN U410 ( .A(N262), .B(z2[211]), .Z(n277) );
  NANDN U411 ( .A(n3), .B(N475), .Z(n276) );
  NAND U412 ( .A(n278), .B(n279), .Z(z3[210]) );
  NANDN U413 ( .A(N262), .B(z2[210]), .Z(n279) );
  NANDN U414 ( .A(n3), .B(N474), .Z(n278) );
  NAND U415 ( .A(n280), .B(n281), .Z(z3[20]) );
  NANDN U416 ( .A(N262), .B(z2[20]), .Z(n281) );
  NANDN U417 ( .A(n3), .B(N284), .Z(n280) );
  NAND U418 ( .A(n282), .B(n283), .Z(z3[209]) );
  NANDN U419 ( .A(N262), .B(z2[209]), .Z(n283) );
  NANDN U420 ( .A(n3), .B(N473), .Z(n282) );
  NAND U421 ( .A(n284), .B(n285), .Z(z3[208]) );
  NANDN U422 ( .A(N262), .B(z2[208]), .Z(n285) );
  NANDN U423 ( .A(n3), .B(N472), .Z(n284) );
  NAND U424 ( .A(n286), .B(n287), .Z(z3[207]) );
  NANDN U425 ( .A(N262), .B(z2[207]), .Z(n287) );
  NANDN U426 ( .A(n3), .B(N471), .Z(n286) );
  NAND U427 ( .A(n288), .B(n289), .Z(z3[206]) );
  NANDN U428 ( .A(N262), .B(z2[206]), .Z(n289) );
  NANDN U429 ( .A(n3), .B(N470), .Z(n288) );
  NAND U430 ( .A(n290), .B(n291), .Z(z3[205]) );
  NANDN U431 ( .A(N262), .B(z2[205]), .Z(n291) );
  NANDN U432 ( .A(n3), .B(N469), .Z(n290) );
  NAND U433 ( .A(n292), .B(n293), .Z(z3[204]) );
  NANDN U434 ( .A(N262), .B(z2[204]), .Z(n293) );
  NANDN U435 ( .A(n3), .B(N468), .Z(n292) );
  NAND U436 ( .A(n294), .B(n295), .Z(z3[203]) );
  NANDN U437 ( .A(N262), .B(z2[203]), .Z(n295) );
  NANDN U438 ( .A(n3), .B(N467), .Z(n294) );
  NAND U439 ( .A(n296), .B(n297), .Z(z3[202]) );
  NANDN U440 ( .A(N262), .B(z2[202]), .Z(n297) );
  NANDN U441 ( .A(n3), .B(N466), .Z(n296) );
  NAND U442 ( .A(n298), .B(n299), .Z(z3[201]) );
  NANDN U443 ( .A(N262), .B(z2[201]), .Z(n299) );
  NANDN U444 ( .A(n3), .B(N465), .Z(n298) );
  NAND U445 ( .A(n300), .B(n301), .Z(z3[200]) );
  NANDN U446 ( .A(N262), .B(z2[200]), .Z(n301) );
  NANDN U447 ( .A(n3), .B(N464), .Z(n300) );
  NAND U448 ( .A(n302), .B(n303), .Z(z3[1]) );
  NANDN U449 ( .A(N262), .B(z2[1]), .Z(n303) );
  NANDN U450 ( .A(n3), .B(N265), .Z(n302) );
  NAND U451 ( .A(n304), .B(n305), .Z(z3[19]) );
  NANDN U452 ( .A(N262), .B(z2[19]), .Z(n305) );
  NANDN U453 ( .A(n3), .B(N283), .Z(n304) );
  NAND U454 ( .A(n306), .B(n307), .Z(z3[199]) );
  NANDN U455 ( .A(N262), .B(z2[199]), .Z(n307) );
  NANDN U456 ( .A(n3), .B(N463), .Z(n306) );
  NAND U457 ( .A(n308), .B(n309), .Z(z3[198]) );
  NANDN U458 ( .A(N262), .B(z2[198]), .Z(n309) );
  NANDN U459 ( .A(n3), .B(N462), .Z(n308) );
  NAND U460 ( .A(n310), .B(n311), .Z(z3[197]) );
  NANDN U461 ( .A(N262), .B(z2[197]), .Z(n311) );
  NANDN U462 ( .A(n3), .B(N461), .Z(n310) );
  NAND U463 ( .A(n312), .B(n313), .Z(z3[196]) );
  NANDN U464 ( .A(N262), .B(z2[196]), .Z(n313) );
  NANDN U465 ( .A(n3), .B(N460), .Z(n312) );
  NAND U466 ( .A(n314), .B(n315), .Z(z3[195]) );
  NANDN U467 ( .A(N262), .B(z2[195]), .Z(n315) );
  NANDN U468 ( .A(n3), .B(N459), .Z(n314) );
  NAND U469 ( .A(n316), .B(n317), .Z(z3[194]) );
  NANDN U470 ( .A(N262), .B(z2[194]), .Z(n317) );
  NANDN U471 ( .A(n3), .B(N458), .Z(n316) );
  NAND U472 ( .A(n318), .B(n319), .Z(z3[193]) );
  NANDN U473 ( .A(N262), .B(z2[193]), .Z(n319) );
  NANDN U474 ( .A(n3), .B(N457), .Z(n318) );
  NAND U475 ( .A(n320), .B(n321), .Z(z3[192]) );
  NANDN U476 ( .A(N262), .B(z2[192]), .Z(n321) );
  NANDN U477 ( .A(n3), .B(N456), .Z(n320) );
  NAND U478 ( .A(n322), .B(n323), .Z(z3[191]) );
  NANDN U479 ( .A(N262), .B(z2[191]), .Z(n323) );
  NANDN U480 ( .A(n3), .B(N455), .Z(n322) );
  NAND U481 ( .A(n324), .B(n325), .Z(z3[190]) );
  NANDN U482 ( .A(N262), .B(z2[190]), .Z(n325) );
  NANDN U483 ( .A(n3), .B(N454), .Z(n324) );
  NAND U484 ( .A(n326), .B(n327), .Z(z3[18]) );
  NANDN U485 ( .A(N262), .B(z2[18]), .Z(n327) );
  NANDN U486 ( .A(n3), .B(N282), .Z(n326) );
  NAND U487 ( .A(n328), .B(n329), .Z(z3[189]) );
  NANDN U488 ( .A(N262), .B(z2[189]), .Z(n329) );
  NANDN U489 ( .A(n3), .B(N453), .Z(n328) );
  NAND U490 ( .A(n330), .B(n331), .Z(z3[188]) );
  NANDN U491 ( .A(N262), .B(z2[188]), .Z(n331) );
  NANDN U492 ( .A(n3), .B(N452), .Z(n330) );
  NAND U493 ( .A(n332), .B(n333), .Z(z3[187]) );
  NANDN U494 ( .A(N262), .B(z2[187]), .Z(n333) );
  NANDN U495 ( .A(n3), .B(N451), .Z(n332) );
  NAND U496 ( .A(n334), .B(n335), .Z(z3[186]) );
  NANDN U497 ( .A(N262), .B(z2[186]), .Z(n335) );
  NANDN U498 ( .A(n3), .B(N450), .Z(n334) );
  NAND U499 ( .A(n336), .B(n337), .Z(z3[185]) );
  NANDN U500 ( .A(N262), .B(z2[185]), .Z(n337) );
  NANDN U501 ( .A(n3), .B(N449), .Z(n336) );
  NAND U502 ( .A(n338), .B(n339), .Z(z3[184]) );
  NANDN U503 ( .A(N262), .B(z2[184]), .Z(n339) );
  NANDN U504 ( .A(n3), .B(N448), .Z(n338) );
  NAND U505 ( .A(n340), .B(n341), .Z(z3[183]) );
  NANDN U506 ( .A(N262), .B(z2[183]), .Z(n341) );
  NANDN U507 ( .A(n3), .B(N447), .Z(n340) );
  NAND U508 ( .A(n342), .B(n343), .Z(z3[182]) );
  NANDN U509 ( .A(N262), .B(z2[182]), .Z(n343) );
  NANDN U510 ( .A(n3), .B(N446), .Z(n342) );
  NAND U511 ( .A(n344), .B(n345), .Z(z3[181]) );
  NANDN U512 ( .A(N262), .B(z2[181]), .Z(n345) );
  NANDN U513 ( .A(n3), .B(N445), .Z(n344) );
  NAND U514 ( .A(n346), .B(n347), .Z(z3[180]) );
  NANDN U515 ( .A(N262), .B(z2[180]), .Z(n347) );
  NANDN U516 ( .A(n3), .B(N444), .Z(n346) );
  NAND U517 ( .A(n348), .B(n349), .Z(z3[17]) );
  NANDN U518 ( .A(N262), .B(z2[17]), .Z(n349) );
  NANDN U519 ( .A(n3), .B(N281), .Z(n348) );
  NAND U520 ( .A(n350), .B(n351), .Z(z3[179]) );
  NANDN U521 ( .A(N262), .B(z2[179]), .Z(n351) );
  NANDN U522 ( .A(n3), .B(N443), .Z(n350) );
  NAND U523 ( .A(n352), .B(n353), .Z(z3[178]) );
  NANDN U524 ( .A(N262), .B(z2[178]), .Z(n353) );
  NANDN U525 ( .A(n3), .B(N442), .Z(n352) );
  NAND U526 ( .A(n354), .B(n355), .Z(z3[177]) );
  NANDN U527 ( .A(N262), .B(z2[177]), .Z(n355) );
  NANDN U528 ( .A(n3), .B(N441), .Z(n354) );
  NAND U529 ( .A(n356), .B(n357), .Z(z3[176]) );
  NANDN U530 ( .A(N262), .B(z2[176]), .Z(n357) );
  NANDN U531 ( .A(n3), .B(N440), .Z(n356) );
  NAND U532 ( .A(n358), .B(n359), .Z(z3[175]) );
  NANDN U533 ( .A(N262), .B(z2[175]), .Z(n359) );
  NANDN U534 ( .A(n3), .B(N439), .Z(n358) );
  NAND U535 ( .A(n360), .B(n361), .Z(z3[174]) );
  NANDN U536 ( .A(N262), .B(z2[174]), .Z(n361) );
  NANDN U537 ( .A(n3), .B(N438), .Z(n360) );
  NAND U538 ( .A(n362), .B(n363), .Z(z3[173]) );
  NANDN U539 ( .A(N262), .B(z2[173]), .Z(n363) );
  NANDN U540 ( .A(n3), .B(N437), .Z(n362) );
  NAND U541 ( .A(n364), .B(n365), .Z(z3[172]) );
  NANDN U542 ( .A(N262), .B(z2[172]), .Z(n365) );
  NANDN U543 ( .A(n3), .B(N436), .Z(n364) );
  NAND U544 ( .A(n366), .B(n367), .Z(z3[171]) );
  NANDN U545 ( .A(N262), .B(z2[171]), .Z(n367) );
  NANDN U546 ( .A(n3), .B(N435), .Z(n366) );
  NAND U547 ( .A(n368), .B(n369), .Z(z3[170]) );
  NANDN U548 ( .A(N262), .B(z2[170]), .Z(n369) );
  NANDN U549 ( .A(n3), .B(N434), .Z(n368) );
  NAND U550 ( .A(n370), .B(n371), .Z(z3[16]) );
  NANDN U551 ( .A(N262), .B(z2[16]), .Z(n371) );
  NANDN U552 ( .A(n3), .B(N280), .Z(n370) );
  NAND U553 ( .A(n372), .B(n373), .Z(z3[169]) );
  NANDN U554 ( .A(N262), .B(z2[169]), .Z(n373) );
  NANDN U555 ( .A(n3), .B(N433), .Z(n372) );
  NAND U556 ( .A(n374), .B(n375), .Z(z3[168]) );
  NANDN U557 ( .A(N262), .B(z2[168]), .Z(n375) );
  NANDN U558 ( .A(n3), .B(N432), .Z(n374) );
  NAND U559 ( .A(n376), .B(n377), .Z(z3[167]) );
  NANDN U560 ( .A(N262), .B(z2[167]), .Z(n377) );
  NANDN U561 ( .A(n3), .B(N431), .Z(n376) );
  NAND U562 ( .A(n378), .B(n379), .Z(z3[166]) );
  NANDN U563 ( .A(N262), .B(z2[166]), .Z(n379) );
  NANDN U564 ( .A(n3), .B(N430), .Z(n378) );
  NAND U565 ( .A(n380), .B(n381), .Z(z3[165]) );
  NANDN U566 ( .A(N262), .B(z2[165]), .Z(n381) );
  NANDN U567 ( .A(n3), .B(N429), .Z(n380) );
  NAND U568 ( .A(n382), .B(n383), .Z(z3[164]) );
  NANDN U569 ( .A(N262), .B(z2[164]), .Z(n383) );
  NANDN U570 ( .A(n3), .B(N428), .Z(n382) );
  NAND U571 ( .A(n384), .B(n385), .Z(z3[163]) );
  NANDN U572 ( .A(N262), .B(z2[163]), .Z(n385) );
  NANDN U573 ( .A(n3), .B(N427), .Z(n384) );
  NAND U574 ( .A(n386), .B(n387), .Z(z3[162]) );
  NANDN U575 ( .A(N262), .B(z2[162]), .Z(n387) );
  NANDN U576 ( .A(n3), .B(N426), .Z(n386) );
  NAND U577 ( .A(n388), .B(n389), .Z(z3[161]) );
  NANDN U578 ( .A(N262), .B(z2[161]), .Z(n389) );
  NANDN U579 ( .A(n3), .B(N425), .Z(n388) );
  NAND U580 ( .A(n390), .B(n391), .Z(z3[160]) );
  NANDN U581 ( .A(N262), .B(z2[160]), .Z(n391) );
  NANDN U582 ( .A(n3), .B(N424), .Z(n390) );
  NAND U583 ( .A(n392), .B(n393), .Z(z3[15]) );
  NANDN U584 ( .A(N262), .B(z2[15]), .Z(n393) );
  NANDN U585 ( .A(n3), .B(N279), .Z(n392) );
  NAND U586 ( .A(n394), .B(n395), .Z(z3[159]) );
  NANDN U587 ( .A(N262), .B(z2[159]), .Z(n395) );
  NANDN U588 ( .A(n3), .B(N423), .Z(n394) );
  NAND U589 ( .A(n396), .B(n397), .Z(z3[158]) );
  NANDN U590 ( .A(N262), .B(z2[158]), .Z(n397) );
  NANDN U591 ( .A(n3), .B(N422), .Z(n396) );
  NAND U592 ( .A(n398), .B(n399), .Z(z3[157]) );
  NANDN U593 ( .A(N262), .B(z2[157]), .Z(n399) );
  NANDN U594 ( .A(n3), .B(N421), .Z(n398) );
  NAND U595 ( .A(n400), .B(n401), .Z(z3[156]) );
  NANDN U596 ( .A(N262), .B(z2[156]), .Z(n401) );
  NANDN U597 ( .A(n3), .B(N420), .Z(n400) );
  NAND U598 ( .A(n402), .B(n403), .Z(z3[155]) );
  NANDN U599 ( .A(N262), .B(z2[155]), .Z(n403) );
  NANDN U600 ( .A(n3), .B(N419), .Z(n402) );
  NAND U601 ( .A(n404), .B(n405), .Z(z3[154]) );
  NANDN U602 ( .A(N262), .B(z2[154]), .Z(n405) );
  NANDN U603 ( .A(n3), .B(N418), .Z(n404) );
  NAND U604 ( .A(n406), .B(n407), .Z(z3[153]) );
  NANDN U605 ( .A(N262), .B(z2[153]), .Z(n407) );
  NANDN U606 ( .A(n3), .B(N417), .Z(n406) );
  NAND U607 ( .A(n408), .B(n409), .Z(z3[152]) );
  NANDN U608 ( .A(N262), .B(z2[152]), .Z(n409) );
  NANDN U609 ( .A(n3), .B(N416), .Z(n408) );
  NAND U610 ( .A(n410), .B(n411), .Z(z3[151]) );
  NANDN U611 ( .A(N262), .B(z2[151]), .Z(n411) );
  NANDN U612 ( .A(n3), .B(N415), .Z(n410) );
  NAND U613 ( .A(n412), .B(n413), .Z(z3[150]) );
  NANDN U614 ( .A(N262), .B(z2[150]), .Z(n413) );
  NANDN U615 ( .A(n3), .B(N414), .Z(n412) );
  NAND U616 ( .A(n414), .B(n415), .Z(z3[14]) );
  NANDN U617 ( .A(N262), .B(z2[14]), .Z(n415) );
  NANDN U618 ( .A(n3), .B(N278), .Z(n414) );
  NAND U619 ( .A(n416), .B(n417), .Z(z3[149]) );
  NANDN U620 ( .A(N262), .B(z2[149]), .Z(n417) );
  NANDN U621 ( .A(n3), .B(N413), .Z(n416) );
  NAND U622 ( .A(n418), .B(n419), .Z(z3[148]) );
  NANDN U623 ( .A(N262), .B(z2[148]), .Z(n419) );
  NANDN U624 ( .A(n3), .B(N412), .Z(n418) );
  NAND U625 ( .A(n420), .B(n421), .Z(z3[147]) );
  NANDN U626 ( .A(N262), .B(z2[147]), .Z(n421) );
  NANDN U627 ( .A(n3), .B(N411), .Z(n420) );
  NAND U628 ( .A(n422), .B(n423), .Z(z3[146]) );
  NANDN U629 ( .A(N262), .B(z2[146]), .Z(n423) );
  NANDN U630 ( .A(n3), .B(N410), .Z(n422) );
  NAND U631 ( .A(n424), .B(n425), .Z(z3[145]) );
  NANDN U632 ( .A(N262), .B(z2[145]), .Z(n425) );
  NANDN U633 ( .A(n3), .B(N409), .Z(n424) );
  NAND U634 ( .A(n426), .B(n427), .Z(z3[144]) );
  NANDN U635 ( .A(N262), .B(z2[144]), .Z(n427) );
  NANDN U636 ( .A(n3), .B(N408), .Z(n426) );
  NAND U637 ( .A(n428), .B(n429), .Z(z3[143]) );
  NANDN U638 ( .A(N262), .B(z2[143]), .Z(n429) );
  NANDN U639 ( .A(n3), .B(N407), .Z(n428) );
  NAND U640 ( .A(n430), .B(n431), .Z(z3[142]) );
  NANDN U641 ( .A(N262), .B(z2[142]), .Z(n431) );
  NANDN U642 ( .A(n3), .B(N406), .Z(n430) );
  NAND U643 ( .A(n432), .B(n433), .Z(z3[141]) );
  NANDN U644 ( .A(N262), .B(z2[141]), .Z(n433) );
  NANDN U645 ( .A(n3), .B(N405), .Z(n432) );
  NAND U646 ( .A(n434), .B(n435), .Z(z3[140]) );
  NANDN U647 ( .A(N262), .B(z2[140]), .Z(n435) );
  NANDN U648 ( .A(n3), .B(N404), .Z(n434) );
  NAND U649 ( .A(n436), .B(n437), .Z(z3[13]) );
  NANDN U650 ( .A(N262), .B(z2[13]), .Z(n437) );
  NANDN U651 ( .A(n3), .B(N277), .Z(n436) );
  NAND U652 ( .A(n438), .B(n439), .Z(z3[139]) );
  NANDN U653 ( .A(N262), .B(z2[139]), .Z(n439) );
  NANDN U654 ( .A(n3), .B(N403), .Z(n438) );
  NAND U655 ( .A(n440), .B(n441), .Z(z3[138]) );
  NANDN U656 ( .A(N262), .B(z2[138]), .Z(n441) );
  NANDN U657 ( .A(n3), .B(N402), .Z(n440) );
  NAND U658 ( .A(n442), .B(n443), .Z(z3[137]) );
  NANDN U659 ( .A(N262), .B(z2[137]), .Z(n443) );
  NANDN U660 ( .A(n3), .B(N401), .Z(n442) );
  NAND U661 ( .A(n444), .B(n445), .Z(z3[136]) );
  NANDN U662 ( .A(N262), .B(z2[136]), .Z(n445) );
  NANDN U663 ( .A(n3), .B(N400), .Z(n444) );
  NAND U664 ( .A(n446), .B(n447), .Z(z3[135]) );
  NANDN U665 ( .A(N262), .B(z2[135]), .Z(n447) );
  NANDN U666 ( .A(n3), .B(N399), .Z(n446) );
  NAND U667 ( .A(n448), .B(n449), .Z(z3[134]) );
  NANDN U668 ( .A(N262), .B(z2[134]), .Z(n449) );
  NANDN U669 ( .A(n3), .B(N398), .Z(n448) );
  NAND U670 ( .A(n450), .B(n451), .Z(z3[133]) );
  NANDN U671 ( .A(N262), .B(z2[133]), .Z(n451) );
  NANDN U672 ( .A(n3), .B(N397), .Z(n450) );
  NAND U673 ( .A(n452), .B(n453), .Z(z3[132]) );
  NANDN U674 ( .A(N262), .B(z2[132]), .Z(n453) );
  NANDN U675 ( .A(n3), .B(N396), .Z(n452) );
  NAND U676 ( .A(n454), .B(n455), .Z(z3[131]) );
  NANDN U677 ( .A(N262), .B(z2[131]), .Z(n455) );
  NANDN U678 ( .A(n3), .B(N395), .Z(n454) );
  NAND U679 ( .A(n456), .B(n457), .Z(z3[130]) );
  NANDN U680 ( .A(N262), .B(z2[130]), .Z(n457) );
  NANDN U681 ( .A(n3), .B(N394), .Z(n456) );
  NAND U682 ( .A(n458), .B(n459), .Z(z3[12]) );
  NANDN U683 ( .A(N262), .B(z2[12]), .Z(n459) );
  NANDN U684 ( .A(n3), .B(N276), .Z(n458) );
  NAND U685 ( .A(n460), .B(n461), .Z(z3[129]) );
  NANDN U686 ( .A(N262), .B(z2[129]), .Z(n461) );
  NANDN U687 ( .A(n3), .B(N393), .Z(n460) );
  NAND U688 ( .A(n462), .B(n463), .Z(z3[128]) );
  NANDN U689 ( .A(N262), .B(z2[128]), .Z(n463) );
  NANDN U690 ( .A(n3), .B(N392), .Z(n462) );
  NAND U691 ( .A(n464), .B(n465), .Z(z3[127]) );
  NANDN U692 ( .A(N262), .B(z2[127]), .Z(n465) );
  NANDN U693 ( .A(n3), .B(N391), .Z(n464) );
  NAND U694 ( .A(n466), .B(n467), .Z(z3[126]) );
  NANDN U695 ( .A(N262), .B(z2[126]), .Z(n467) );
  NANDN U696 ( .A(n3), .B(N390), .Z(n466) );
  NAND U697 ( .A(n468), .B(n469), .Z(z3[125]) );
  NANDN U698 ( .A(N262), .B(z2[125]), .Z(n469) );
  NANDN U699 ( .A(n3), .B(N389), .Z(n468) );
  NAND U700 ( .A(n470), .B(n471), .Z(z3[124]) );
  NANDN U701 ( .A(N262), .B(z2[124]), .Z(n471) );
  NANDN U702 ( .A(n3), .B(N388), .Z(n470) );
  NAND U703 ( .A(n472), .B(n473), .Z(z3[123]) );
  NANDN U704 ( .A(N262), .B(z2[123]), .Z(n473) );
  NANDN U705 ( .A(n3), .B(N387), .Z(n472) );
  NAND U706 ( .A(n474), .B(n475), .Z(z3[122]) );
  NANDN U707 ( .A(N262), .B(z2[122]), .Z(n475) );
  NANDN U708 ( .A(n3), .B(N386), .Z(n474) );
  NAND U709 ( .A(n476), .B(n477), .Z(z3[121]) );
  NANDN U710 ( .A(N262), .B(z2[121]), .Z(n477) );
  NANDN U711 ( .A(n3), .B(N385), .Z(n476) );
  NAND U712 ( .A(n478), .B(n479), .Z(z3[120]) );
  NANDN U713 ( .A(N262), .B(z2[120]), .Z(n479) );
  NANDN U714 ( .A(n3), .B(N384), .Z(n478) );
  NAND U715 ( .A(n480), .B(n481), .Z(z3[11]) );
  NANDN U716 ( .A(N262), .B(z2[11]), .Z(n481) );
  NANDN U717 ( .A(n3), .B(N275), .Z(n480) );
  NAND U718 ( .A(n482), .B(n483), .Z(z3[119]) );
  NANDN U719 ( .A(N262), .B(z2[119]), .Z(n483) );
  NANDN U720 ( .A(n3), .B(N383), .Z(n482) );
  NAND U721 ( .A(n484), .B(n485), .Z(z3[118]) );
  NANDN U722 ( .A(N262), .B(z2[118]), .Z(n485) );
  NANDN U723 ( .A(n3), .B(N382), .Z(n484) );
  NAND U724 ( .A(n486), .B(n487), .Z(z3[117]) );
  NANDN U725 ( .A(N262), .B(z2[117]), .Z(n487) );
  NANDN U726 ( .A(n3), .B(N381), .Z(n486) );
  NAND U727 ( .A(n488), .B(n489), .Z(z3[116]) );
  NANDN U728 ( .A(N262), .B(z2[116]), .Z(n489) );
  NANDN U729 ( .A(n3), .B(N380), .Z(n488) );
  NAND U730 ( .A(n490), .B(n491), .Z(z3[115]) );
  NANDN U731 ( .A(N262), .B(z2[115]), .Z(n491) );
  NANDN U732 ( .A(n3), .B(N379), .Z(n490) );
  NAND U733 ( .A(n492), .B(n493), .Z(z3[114]) );
  NANDN U734 ( .A(N262), .B(z2[114]), .Z(n493) );
  NANDN U735 ( .A(n3), .B(N378), .Z(n492) );
  NAND U736 ( .A(n494), .B(n495), .Z(z3[113]) );
  NANDN U737 ( .A(N262), .B(z2[113]), .Z(n495) );
  NANDN U738 ( .A(n3), .B(N377), .Z(n494) );
  NAND U739 ( .A(n496), .B(n497), .Z(z3[112]) );
  NANDN U740 ( .A(N262), .B(z2[112]), .Z(n497) );
  NANDN U741 ( .A(n3), .B(N376), .Z(n496) );
  NAND U742 ( .A(n498), .B(n499), .Z(z3[111]) );
  NANDN U743 ( .A(N262), .B(z2[111]), .Z(n499) );
  NANDN U744 ( .A(n3), .B(N375), .Z(n498) );
  NAND U745 ( .A(n500), .B(n501), .Z(z3[110]) );
  NANDN U746 ( .A(N262), .B(z2[110]), .Z(n501) );
  NANDN U747 ( .A(n3), .B(N374), .Z(n500) );
  NAND U748 ( .A(n502), .B(n503), .Z(z3[10]) );
  NANDN U749 ( .A(N262), .B(z2[10]), .Z(n503) );
  NANDN U750 ( .A(n3), .B(N274), .Z(n502) );
  NAND U751 ( .A(n504), .B(n505), .Z(z3[109]) );
  NANDN U752 ( .A(N262), .B(z2[109]), .Z(n505) );
  NANDN U753 ( .A(n3), .B(N373), .Z(n504) );
  NAND U754 ( .A(n506), .B(n507), .Z(z3[108]) );
  NANDN U755 ( .A(N262), .B(z2[108]), .Z(n507) );
  NANDN U756 ( .A(n3), .B(N372), .Z(n506) );
  NAND U757 ( .A(n508), .B(n509), .Z(z3[107]) );
  NANDN U758 ( .A(N262), .B(z2[107]), .Z(n509) );
  NANDN U759 ( .A(n3), .B(N371), .Z(n508) );
  NAND U760 ( .A(n510), .B(n511), .Z(z3[106]) );
  NANDN U761 ( .A(N262), .B(z2[106]), .Z(n511) );
  NANDN U762 ( .A(n3), .B(N370), .Z(n510) );
  NAND U763 ( .A(n512), .B(n513), .Z(z3[105]) );
  NANDN U764 ( .A(N262), .B(z2[105]), .Z(n513) );
  NANDN U765 ( .A(n3), .B(N369), .Z(n512) );
  NAND U766 ( .A(n514), .B(n515), .Z(z3[104]) );
  NANDN U767 ( .A(N262), .B(z2[104]), .Z(n515) );
  NANDN U768 ( .A(n3), .B(N368), .Z(n514) );
  NAND U769 ( .A(n516), .B(n517), .Z(z3[103]) );
  NANDN U770 ( .A(N262), .B(z2[103]), .Z(n517) );
  NANDN U771 ( .A(n3), .B(N367), .Z(n516) );
  NAND U772 ( .A(n518), .B(n519), .Z(z3[102]) );
  NANDN U773 ( .A(N262), .B(z2[102]), .Z(n519) );
  NANDN U774 ( .A(n3), .B(N366), .Z(n518) );
  NAND U775 ( .A(n520), .B(n521), .Z(z3[101]) );
  NANDN U776 ( .A(N262), .B(z2[101]), .Z(n521) );
  NANDN U777 ( .A(n3), .B(N365), .Z(n520) );
  NAND U778 ( .A(n522), .B(n523), .Z(z3[100]) );
  NANDN U779 ( .A(N262), .B(z2[100]), .Z(n523) );
  NANDN U780 ( .A(n3), .B(N364), .Z(n522) );
  NAND U781 ( .A(n524), .B(n525), .Z(z3[0]) );
  NANDN U782 ( .A(N262), .B(z2[0]), .Z(n525) );
  NANDN U783 ( .A(n3), .B(N264), .Z(n524) );
  IV U784 ( .A(N262), .Z(n3) );
  NAND U785 ( .A(n526), .B(n527), .Z(z2[9]) );
  NANDN U786 ( .A(xregN_1), .B(zin[8]), .Z(n527) );
  NAND U787 ( .A(N13), .B(xregN_1), .Z(n526) );
  NAND U788 ( .A(n528), .B(n529), .Z(z2[99]) );
  NANDN U789 ( .A(xregN_1), .B(zin[98]), .Z(n529) );
  NAND U790 ( .A(N103), .B(xregN_1), .Z(n528) );
  NAND U791 ( .A(n530), .B(n531), .Z(z2[98]) );
  NANDN U792 ( .A(xregN_1), .B(zin[97]), .Z(n531) );
  NAND U793 ( .A(N102), .B(xregN_1), .Z(n530) );
  NAND U794 ( .A(n532), .B(n533), .Z(z2[97]) );
  NANDN U795 ( .A(xregN_1), .B(zin[96]), .Z(n533) );
  NAND U796 ( .A(N101), .B(xregN_1), .Z(n532) );
  NAND U797 ( .A(n534), .B(n535), .Z(z2[96]) );
  NANDN U798 ( .A(xregN_1), .B(zin[95]), .Z(n535) );
  NAND U799 ( .A(N100), .B(xregN_1), .Z(n534) );
  NAND U800 ( .A(n536), .B(n537), .Z(z2[95]) );
  NANDN U801 ( .A(xregN_1), .B(zin[94]), .Z(n537) );
  NAND U802 ( .A(N99), .B(xregN_1), .Z(n536) );
  NAND U803 ( .A(n538), .B(n539), .Z(z2[94]) );
  NANDN U804 ( .A(xregN_1), .B(zin[93]), .Z(n539) );
  NAND U805 ( .A(N98), .B(xregN_1), .Z(n538) );
  NAND U806 ( .A(n540), .B(n541), .Z(z2[93]) );
  NANDN U807 ( .A(xregN_1), .B(zin[92]), .Z(n541) );
  NAND U808 ( .A(N97), .B(xregN_1), .Z(n540) );
  NAND U809 ( .A(n542), .B(n543), .Z(z2[92]) );
  NANDN U810 ( .A(xregN_1), .B(zin[91]), .Z(n543) );
  NAND U811 ( .A(N96), .B(xregN_1), .Z(n542) );
  NAND U812 ( .A(n544), .B(n545), .Z(z2[91]) );
  NANDN U813 ( .A(xregN_1), .B(zin[90]), .Z(n545) );
  NAND U814 ( .A(N95), .B(xregN_1), .Z(n544) );
  NAND U815 ( .A(n546), .B(n547), .Z(z2[90]) );
  NANDN U816 ( .A(xregN_1), .B(zin[89]), .Z(n547) );
  NAND U817 ( .A(N94), .B(xregN_1), .Z(n546) );
  NAND U818 ( .A(n548), .B(n549), .Z(z2[8]) );
  NANDN U819 ( .A(xregN_1), .B(zin[7]), .Z(n549) );
  NAND U820 ( .A(N12), .B(xregN_1), .Z(n548) );
  NAND U821 ( .A(n550), .B(n551), .Z(z2[89]) );
  NANDN U822 ( .A(xregN_1), .B(zin[88]), .Z(n551) );
  NAND U823 ( .A(N93), .B(xregN_1), .Z(n550) );
  NAND U824 ( .A(n552), .B(n553), .Z(z2[88]) );
  NANDN U825 ( .A(xregN_1), .B(zin[87]), .Z(n553) );
  NAND U826 ( .A(N92), .B(xregN_1), .Z(n552) );
  NAND U827 ( .A(n554), .B(n555), .Z(z2[87]) );
  NANDN U828 ( .A(xregN_1), .B(zin[86]), .Z(n555) );
  NAND U829 ( .A(N91), .B(xregN_1), .Z(n554) );
  NAND U830 ( .A(n556), .B(n557), .Z(z2[86]) );
  NANDN U831 ( .A(xregN_1), .B(zin[85]), .Z(n557) );
  NAND U832 ( .A(N90), .B(xregN_1), .Z(n556) );
  NAND U833 ( .A(n558), .B(n559), .Z(z2[85]) );
  NANDN U834 ( .A(xregN_1), .B(zin[84]), .Z(n559) );
  NAND U835 ( .A(N89), .B(xregN_1), .Z(n558) );
  NAND U836 ( .A(n560), .B(n561), .Z(z2[84]) );
  NANDN U837 ( .A(xregN_1), .B(zin[83]), .Z(n561) );
  NAND U838 ( .A(N88), .B(xregN_1), .Z(n560) );
  NAND U839 ( .A(n562), .B(n563), .Z(z2[83]) );
  NANDN U840 ( .A(xregN_1), .B(zin[82]), .Z(n563) );
  NAND U841 ( .A(N87), .B(xregN_1), .Z(n562) );
  NAND U842 ( .A(n564), .B(n565), .Z(z2[82]) );
  NANDN U843 ( .A(xregN_1), .B(zin[81]), .Z(n565) );
  NAND U844 ( .A(N86), .B(xregN_1), .Z(n564) );
  NAND U845 ( .A(n566), .B(n567), .Z(z2[81]) );
  NANDN U846 ( .A(xregN_1), .B(zin[80]), .Z(n567) );
  NAND U847 ( .A(N85), .B(xregN_1), .Z(n566) );
  NAND U848 ( .A(n568), .B(n569), .Z(z2[80]) );
  NANDN U849 ( .A(xregN_1), .B(zin[79]), .Z(n569) );
  NAND U850 ( .A(N84), .B(xregN_1), .Z(n568) );
  NAND U851 ( .A(n570), .B(n571), .Z(z2[7]) );
  NANDN U852 ( .A(xregN_1), .B(zin[6]), .Z(n571) );
  NAND U853 ( .A(N11), .B(xregN_1), .Z(n570) );
  NAND U854 ( .A(n572), .B(n573), .Z(z2[79]) );
  NANDN U855 ( .A(xregN_1), .B(zin[78]), .Z(n573) );
  NAND U856 ( .A(N83), .B(xregN_1), .Z(n572) );
  NAND U857 ( .A(n574), .B(n575), .Z(z2[78]) );
  NANDN U858 ( .A(xregN_1), .B(zin[77]), .Z(n575) );
  NAND U859 ( .A(N82), .B(xregN_1), .Z(n574) );
  NAND U860 ( .A(n576), .B(n577), .Z(z2[77]) );
  NANDN U861 ( .A(xregN_1), .B(zin[76]), .Z(n577) );
  NAND U862 ( .A(N81), .B(xregN_1), .Z(n576) );
  NAND U863 ( .A(n578), .B(n579), .Z(z2[76]) );
  NANDN U864 ( .A(xregN_1), .B(zin[75]), .Z(n579) );
  NAND U865 ( .A(N80), .B(xregN_1), .Z(n578) );
  NAND U866 ( .A(n580), .B(n581), .Z(z2[75]) );
  NANDN U867 ( .A(xregN_1), .B(zin[74]), .Z(n581) );
  NAND U868 ( .A(N79), .B(xregN_1), .Z(n580) );
  NAND U869 ( .A(n582), .B(n583), .Z(z2[74]) );
  NANDN U870 ( .A(xregN_1), .B(zin[73]), .Z(n583) );
  NAND U871 ( .A(N78), .B(xregN_1), .Z(n582) );
  NAND U872 ( .A(n584), .B(n585), .Z(z2[73]) );
  NANDN U873 ( .A(xregN_1), .B(zin[72]), .Z(n585) );
  NAND U874 ( .A(N77), .B(xregN_1), .Z(n584) );
  NAND U875 ( .A(n586), .B(n587), .Z(z2[72]) );
  NANDN U876 ( .A(xregN_1), .B(zin[71]), .Z(n587) );
  NAND U877 ( .A(N76), .B(xregN_1), .Z(n586) );
  NAND U878 ( .A(n588), .B(n589), .Z(z2[71]) );
  NANDN U879 ( .A(xregN_1), .B(zin[70]), .Z(n589) );
  NAND U880 ( .A(N75), .B(xregN_1), .Z(n588) );
  NAND U881 ( .A(n590), .B(n591), .Z(z2[70]) );
  NANDN U882 ( .A(xregN_1), .B(zin[69]), .Z(n591) );
  NAND U883 ( .A(N74), .B(xregN_1), .Z(n590) );
  NAND U884 ( .A(n592), .B(n593), .Z(z2[6]) );
  NANDN U885 ( .A(xregN_1), .B(zin[5]), .Z(n593) );
  NAND U886 ( .A(N10), .B(xregN_1), .Z(n592) );
  NAND U887 ( .A(n594), .B(n595), .Z(z2[69]) );
  NANDN U888 ( .A(xregN_1), .B(zin[68]), .Z(n595) );
  NAND U889 ( .A(N73), .B(xregN_1), .Z(n594) );
  NAND U890 ( .A(n596), .B(n597), .Z(z2[68]) );
  NANDN U891 ( .A(xregN_1), .B(zin[67]), .Z(n597) );
  NAND U892 ( .A(N72), .B(xregN_1), .Z(n596) );
  NAND U893 ( .A(n598), .B(n599), .Z(z2[67]) );
  NANDN U894 ( .A(xregN_1), .B(zin[66]), .Z(n599) );
  NAND U895 ( .A(N71), .B(xregN_1), .Z(n598) );
  NAND U896 ( .A(n600), .B(n601), .Z(z2[66]) );
  NANDN U897 ( .A(xregN_1), .B(zin[65]), .Z(n601) );
  NAND U898 ( .A(N70), .B(xregN_1), .Z(n600) );
  NAND U899 ( .A(n602), .B(n603), .Z(z2[65]) );
  NANDN U900 ( .A(xregN_1), .B(zin[64]), .Z(n603) );
  NAND U901 ( .A(N69), .B(xregN_1), .Z(n602) );
  NAND U902 ( .A(n604), .B(n605), .Z(z2[64]) );
  NANDN U903 ( .A(xregN_1), .B(zin[63]), .Z(n605) );
  NAND U904 ( .A(N68), .B(xregN_1), .Z(n604) );
  NAND U905 ( .A(n606), .B(n607), .Z(z2[63]) );
  NANDN U906 ( .A(xregN_1), .B(zin[62]), .Z(n607) );
  NAND U907 ( .A(N67), .B(xregN_1), .Z(n606) );
  NAND U908 ( .A(n608), .B(n609), .Z(z2[62]) );
  NANDN U909 ( .A(xregN_1), .B(zin[61]), .Z(n609) );
  NAND U910 ( .A(N66), .B(xregN_1), .Z(n608) );
  NAND U911 ( .A(n610), .B(n611), .Z(z2[61]) );
  NANDN U912 ( .A(xregN_1), .B(zin[60]), .Z(n611) );
  NAND U913 ( .A(N65), .B(xregN_1), .Z(n610) );
  NAND U914 ( .A(n612), .B(n613), .Z(z2[60]) );
  NANDN U915 ( .A(xregN_1), .B(zin[59]), .Z(n613) );
  NAND U916 ( .A(N64), .B(xregN_1), .Z(n612) );
  NAND U917 ( .A(n614), .B(n615), .Z(z2[5]) );
  NANDN U918 ( .A(xregN_1), .B(zin[4]), .Z(n615) );
  NAND U919 ( .A(N9), .B(xregN_1), .Z(n614) );
  NAND U920 ( .A(n616), .B(n617), .Z(z2[59]) );
  NANDN U921 ( .A(xregN_1), .B(zin[58]), .Z(n617) );
  NAND U922 ( .A(N63), .B(xregN_1), .Z(n616) );
  NAND U923 ( .A(n618), .B(n619), .Z(z2[58]) );
  NANDN U924 ( .A(xregN_1), .B(zin[57]), .Z(n619) );
  NAND U925 ( .A(N62), .B(xregN_1), .Z(n618) );
  NAND U926 ( .A(n620), .B(n621), .Z(z2[57]) );
  NANDN U927 ( .A(xregN_1), .B(zin[56]), .Z(n621) );
  NAND U928 ( .A(N61), .B(xregN_1), .Z(n620) );
  NAND U929 ( .A(n622), .B(n623), .Z(z2[56]) );
  NANDN U930 ( .A(xregN_1), .B(zin[55]), .Z(n623) );
  NAND U931 ( .A(N60), .B(xregN_1), .Z(n622) );
  NAND U932 ( .A(n624), .B(n625), .Z(z2[55]) );
  NANDN U933 ( .A(xregN_1), .B(zin[54]), .Z(n625) );
  NAND U934 ( .A(N59), .B(xregN_1), .Z(n624) );
  NAND U935 ( .A(n626), .B(n627), .Z(z2[54]) );
  NANDN U936 ( .A(xregN_1), .B(zin[53]), .Z(n627) );
  NAND U937 ( .A(N58), .B(xregN_1), .Z(n626) );
  NAND U938 ( .A(n628), .B(n629), .Z(z2[53]) );
  NANDN U939 ( .A(xregN_1), .B(zin[52]), .Z(n629) );
  NAND U940 ( .A(N57), .B(xregN_1), .Z(n628) );
  NAND U941 ( .A(n630), .B(n631), .Z(z2[52]) );
  NANDN U942 ( .A(xregN_1), .B(zin[51]), .Z(n631) );
  NAND U943 ( .A(N56), .B(xregN_1), .Z(n630) );
  NAND U944 ( .A(n632), .B(n633), .Z(z2[51]) );
  NANDN U945 ( .A(xregN_1), .B(zin[50]), .Z(n633) );
  NAND U946 ( .A(N55), .B(xregN_1), .Z(n632) );
  NAND U947 ( .A(n634), .B(n635), .Z(z2[50]) );
  NANDN U948 ( .A(xregN_1), .B(zin[49]), .Z(n635) );
  NAND U949 ( .A(N54), .B(xregN_1), .Z(n634) );
  NAND U950 ( .A(n636), .B(n637), .Z(z2[4]) );
  NANDN U951 ( .A(xregN_1), .B(zin[3]), .Z(n637) );
  NAND U952 ( .A(N8), .B(xregN_1), .Z(n636) );
  NAND U953 ( .A(n638), .B(n639), .Z(z2[49]) );
  NANDN U954 ( .A(xregN_1), .B(zin[48]), .Z(n639) );
  NAND U955 ( .A(N53), .B(xregN_1), .Z(n638) );
  NAND U956 ( .A(n640), .B(n641), .Z(z2[48]) );
  NANDN U957 ( .A(xregN_1), .B(zin[47]), .Z(n641) );
  NAND U958 ( .A(N52), .B(xregN_1), .Z(n640) );
  NAND U959 ( .A(n642), .B(n643), .Z(z2[47]) );
  NANDN U960 ( .A(xregN_1), .B(zin[46]), .Z(n643) );
  NAND U961 ( .A(N51), .B(xregN_1), .Z(n642) );
  NAND U962 ( .A(n644), .B(n645), .Z(z2[46]) );
  NANDN U963 ( .A(xregN_1), .B(zin[45]), .Z(n645) );
  NAND U964 ( .A(N50), .B(xregN_1), .Z(n644) );
  NAND U965 ( .A(n646), .B(n647), .Z(z2[45]) );
  NANDN U966 ( .A(xregN_1), .B(zin[44]), .Z(n647) );
  NAND U967 ( .A(N49), .B(xregN_1), .Z(n646) );
  NAND U968 ( .A(n648), .B(n649), .Z(z2[44]) );
  NANDN U969 ( .A(xregN_1), .B(zin[43]), .Z(n649) );
  NAND U970 ( .A(N48), .B(xregN_1), .Z(n648) );
  NAND U971 ( .A(n650), .B(n651), .Z(z2[43]) );
  NANDN U972 ( .A(xregN_1), .B(zin[42]), .Z(n651) );
  NAND U973 ( .A(N47), .B(xregN_1), .Z(n650) );
  NAND U974 ( .A(n652), .B(n653), .Z(z2[42]) );
  NANDN U975 ( .A(xregN_1), .B(zin[41]), .Z(n653) );
  NAND U976 ( .A(N46), .B(xregN_1), .Z(n652) );
  NAND U977 ( .A(n654), .B(n655), .Z(z2[41]) );
  NANDN U978 ( .A(xregN_1), .B(zin[40]), .Z(n655) );
  NAND U979 ( .A(N45), .B(xregN_1), .Z(n654) );
  NAND U980 ( .A(n656), .B(n657), .Z(z2[40]) );
  NANDN U981 ( .A(xregN_1), .B(zin[39]), .Z(n657) );
  NAND U982 ( .A(N44), .B(xregN_1), .Z(n656) );
  NAND U983 ( .A(n658), .B(n659), .Z(z2[3]) );
  NANDN U984 ( .A(xregN_1), .B(zin[2]), .Z(n659) );
  NAND U985 ( .A(N7), .B(xregN_1), .Z(n658) );
  NAND U986 ( .A(n660), .B(n661), .Z(z2[39]) );
  NANDN U987 ( .A(xregN_1), .B(zin[38]), .Z(n661) );
  NAND U988 ( .A(N43), .B(xregN_1), .Z(n660) );
  NAND U989 ( .A(n662), .B(n663), .Z(z2[38]) );
  NANDN U990 ( .A(xregN_1), .B(zin[37]), .Z(n663) );
  NAND U991 ( .A(N42), .B(xregN_1), .Z(n662) );
  NAND U992 ( .A(n664), .B(n665), .Z(z2[37]) );
  NANDN U993 ( .A(xregN_1), .B(zin[36]), .Z(n665) );
  NAND U994 ( .A(N41), .B(xregN_1), .Z(n664) );
  NAND U995 ( .A(n666), .B(n667), .Z(z2[36]) );
  NANDN U996 ( .A(xregN_1), .B(zin[35]), .Z(n667) );
  NAND U997 ( .A(N40), .B(xregN_1), .Z(n666) );
  NAND U998 ( .A(n668), .B(n669), .Z(z2[35]) );
  NANDN U999 ( .A(xregN_1), .B(zin[34]), .Z(n669) );
  NAND U1000 ( .A(N39), .B(xregN_1), .Z(n668) );
  NAND U1001 ( .A(n670), .B(n671), .Z(z2[34]) );
  NANDN U1002 ( .A(xregN_1), .B(zin[33]), .Z(n671) );
  NAND U1003 ( .A(N38), .B(xregN_1), .Z(n670) );
  NAND U1004 ( .A(n672), .B(n673), .Z(z2[33]) );
  NANDN U1005 ( .A(xregN_1), .B(zin[32]), .Z(n673) );
  NAND U1006 ( .A(N37), .B(xregN_1), .Z(n672) );
  NAND U1007 ( .A(n674), .B(n675), .Z(z2[32]) );
  NANDN U1008 ( .A(xregN_1), .B(zin[31]), .Z(n675) );
  NAND U1009 ( .A(N36), .B(xregN_1), .Z(n674) );
  NAND U1010 ( .A(n676), .B(n677), .Z(z2[31]) );
  NANDN U1011 ( .A(xregN_1), .B(zin[30]), .Z(n677) );
  NAND U1012 ( .A(N35), .B(xregN_1), .Z(n676) );
  NAND U1013 ( .A(n678), .B(n679), .Z(z2[30]) );
  NANDN U1014 ( .A(xregN_1), .B(zin[29]), .Z(n679) );
  NAND U1015 ( .A(N34), .B(xregN_1), .Z(n678) );
  NAND U1016 ( .A(n680), .B(n681), .Z(z2[2]) );
  NANDN U1017 ( .A(xregN_1), .B(zin[1]), .Z(n681) );
  NAND U1018 ( .A(N6), .B(xregN_1), .Z(n680) );
  NAND U1019 ( .A(n682), .B(n683), .Z(z2[29]) );
  NANDN U1020 ( .A(xregN_1), .B(zin[28]), .Z(n683) );
  NAND U1021 ( .A(N33), .B(xregN_1), .Z(n682) );
  NAND U1022 ( .A(n684), .B(n685), .Z(z2[28]) );
  NANDN U1023 ( .A(xregN_1), .B(zin[27]), .Z(n685) );
  NAND U1024 ( .A(N32), .B(xregN_1), .Z(n684) );
  NAND U1025 ( .A(n686), .B(n687), .Z(z2[27]) );
  NANDN U1026 ( .A(xregN_1), .B(zin[26]), .Z(n687) );
  NAND U1027 ( .A(N31), .B(xregN_1), .Z(n686) );
  NAND U1028 ( .A(n688), .B(n689), .Z(z2[26]) );
  NANDN U1029 ( .A(xregN_1), .B(zin[25]), .Z(n689) );
  NAND U1030 ( .A(N30), .B(xregN_1), .Z(n688) );
  NAND U1031 ( .A(n690), .B(n691), .Z(z2[25]) );
  NANDN U1032 ( .A(xregN_1), .B(zin[24]), .Z(n691) );
  NAND U1033 ( .A(N29), .B(xregN_1), .Z(n690) );
  NAND U1034 ( .A(n692), .B(n693), .Z(z2[257]) );
  NANDN U1035 ( .A(xregN_1), .B(zin[256]), .Z(n693) );
  NAND U1036 ( .A(N261), .B(xregN_1), .Z(n692) );
  NAND U1037 ( .A(n694), .B(n695), .Z(z2[256]) );
  NANDN U1038 ( .A(xregN_1), .B(zin[255]), .Z(n695) );
  NAND U1039 ( .A(N260), .B(xregN_1), .Z(n694) );
  NAND U1040 ( .A(n696), .B(n697), .Z(z2[255]) );
  NANDN U1041 ( .A(xregN_1), .B(zin[254]), .Z(n697) );
  NAND U1042 ( .A(N259), .B(xregN_1), .Z(n696) );
  NAND U1043 ( .A(n698), .B(n699), .Z(z2[254]) );
  NANDN U1044 ( .A(xregN_1), .B(zin[253]), .Z(n699) );
  NAND U1045 ( .A(N258), .B(xregN_1), .Z(n698) );
  NAND U1046 ( .A(n700), .B(n701), .Z(z2[253]) );
  NANDN U1047 ( .A(xregN_1), .B(zin[252]), .Z(n701) );
  NAND U1048 ( .A(N257), .B(xregN_1), .Z(n700) );
  NAND U1049 ( .A(n702), .B(n703), .Z(z2[252]) );
  NANDN U1050 ( .A(xregN_1), .B(zin[251]), .Z(n703) );
  NAND U1051 ( .A(N256), .B(xregN_1), .Z(n702) );
  NAND U1052 ( .A(n704), .B(n705), .Z(z2[251]) );
  NANDN U1053 ( .A(xregN_1), .B(zin[250]), .Z(n705) );
  NAND U1054 ( .A(N255), .B(xregN_1), .Z(n704) );
  NAND U1055 ( .A(n706), .B(n707), .Z(z2[250]) );
  NANDN U1056 ( .A(xregN_1), .B(zin[249]), .Z(n707) );
  NAND U1057 ( .A(N254), .B(xregN_1), .Z(n706) );
  NAND U1058 ( .A(n708), .B(n709), .Z(z2[24]) );
  NANDN U1059 ( .A(xregN_1), .B(zin[23]), .Z(n709) );
  NAND U1060 ( .A(N28), .B(xregN_1), .Z(n708) );
  NAND U1061 ( .A(n710), .B(n711), .Z(z2[249]) );
  NANDN U1062 ( .A(xregN_1), .B(zin[248]), .Z(n711) );
  NAND U1063 ( .A(N253), .B(xregN_1), .Z(n710) );
  NAND U1064 ( .A(n712), .B(n713), .Z(z2[248]) );
  NANDN U1065 ( .A(xregN_1), .B(zin[247]), .Z(n713) );
  NAND U1066 ( .A(N252), .B(xregN_1), .Z(n712) );
  NAND U1067 ( .A(n714), .B(n715), .Z(z2[247]) );
  NANDN U1068 ( .A(xregN_1), .B(zin[246]), .Z(n715) );
  NAND U1069 ( .A(N251), .B(xregN_1), .Z(n714) );
  NAND U1070 ( .A(n716), .B(n717), .Z(z2[246]) );
  NANDN U1071 ( .A(xregN_1), .B(zin[245]), .Z(n717) );
  NAND U1072 ( .A(N250), .B(xregN_1), .Z(n716) );
  NAND U1073 ( .A(n718), .B(n719), .Z(z2[245]) );
  NANDN U1074 ( .A(xregN_1), .B(zin[244]), .Z(n719) );
  NAND U1075 ( .A(N249), .B(xregN_1), .Z(n718) );
  NAND U1076 ( .A(n720), .B(n721), .Z(z2[244]) );
  NANDN U1077 ( .A(xregN_1), .B(zin[243]), .Z(n721) );
  NAND U1078 ( .A(N248), .B(xregN_1), .Z(n720) );
  NAND U1079 ( .A(n722), .B(n723), .Z(z2[243]) );
  NANDN U1080 ( .A(xregN_1), .B(zin[242]), .Z(n723) );
  NAND U1081 ( .A(N247), .B(xregN_1), .Z(n722) );
  NAND U1082 ( .A(n724), .B(n725), .Z(z2[242]) );
  NANDN U1083 ( .A(xregN_1), .B(zin[241]), .Z(n725) );
  NAND U1084 ( .A(N246), .B(xregN_1), .Z(n724) );
  NAND U1085 ( .A(n726), .B(n727), .Z(z2[241]) );
  NANDN U1086 ( .A(xregN_1), .B(zin[240]), .Z(n727) );
  NAND U1087 ( .A(N245), .B(xregN_1), .Z(n726) );
  NAND U1088 ( .A(n728), .B(n729), .Z(z2[240]) );
  NANDN U1089 ( .A(xregN_1), .B(zin[239]), .Z(n729) );
  NAND U1090 ( .A(N244), .B(xregN_1), .Z(n728) );
  NAND U1091 ( .A(n730), .B(n731), .Z(z2[23]) );
  NANDN U1092 ( .A(xregN_1), .B(zin[22]), .Z(n731) );
  NAND U1093 ( .A(N27), .B(xregN_1), .Z(n730) );
  NAND U1094 ( .A(n732), .B(n733), .Z(z2[239]) );
  NANDN U1095 ( .A(xregN_1), .B(zin[238]), .Z(n733) );
  NAND U1096 ( .A(N243), .B(xregN_1), .Z(n732) );
  NAND U1097 ( .A(n734), .B(n735), .Z(z2[238]) );
  NANDN U1098 ( .A(xregN_1), .B(zin[237]), .Z(n735) );
  NAND U1099 ( .A(N242), .B(xregN_1), .Z(n734) );
  NAND U1100 ( .A(n736), .B(n737), .Z(z2[237]) );
  NANDN U1101 ( .A(xregN_1), .B(zin[236]), .Z(n737) );
  NAND U1102 ( .A(N241), .B(xregN_1), .Z(n736) );
  NAND U1103 ( .A(n738), .B(n739), .Z(z2[236]) );
  NANDN U1104 ( .A(xregN_1), .B(zin[235]), .Z(n739) );
  NAND U1105 ( .A(N240), .B(xregN_1), .Z(n738) );
  NAND U1106 ( .A(n740), .B(n741), .Z(z2[235]) );
  NANDN U1107 ( .A(xregN_1), .B(zin[234]), .Z(n741) );
  NAND U1108 ( .A(N239), .B(xregN_1), .Z(n740) );
  NAND U1109 ( .A(n742), .B(n743), .Z(z2[234]) );
  NANDN U1110 ( .A(xregN_1), .B(zin[233]), .Z(n743) );
  NAND U1111 ( .A(N238), .B(xregN_1), .Z(n742) );
  NAND U1112 ( .A(n744), .B(n745), .Z(z2[233]) );
  NANDN U1113 ( .A(xregN_1), .B(zin[232]), .Z(n745) );
  NAND U1114 ( .A(N237), .B(xregN_1), .Z(n744) );
  NAND U1115 ( .A(n746), .B(n747), .Z(z2[232]) );
  NANDN U1116 ( .A(xregN_1), .B(zin[231]), .Z(n747) );
  NAND U1117 ( .A(N236), .B(xregN_1), .Z(n746) );
  NAND U1118 ( .A(n748), .B(n749), .Z(z2[231]) );
  NANDN U1119 ( .A(xregN_1), .B(zin[230]), .Z(n749) );
  NAND U1120 ( .A(N235), .B(xregN_1), .Z(n748) );
  NAND U1121 ( .A(n750), .B(n751), .Z(z2[230]) );
  NANDN U1122 ( .A(xregN_1), .B(zin[229]), .Z(n751) );
  NAND U1123 ( .A(N234), .B(xregN_1), .Z(n750) );
  NAND U1124 ( .A(n752), .B(n753), .Z(z2[22]) );
  NANDN U1125 ( .A(xregN_1), .B(zin[21]), .Z(n753) );
  NAND U1126 ( .A(N26), .B(xregN_1), .Z(n752) );
  NAND U1127 ( .A(n754), .B(n755), .Z(z2[229]) );
  NANDN U1128 ( .A(xregN_1), .B(zin[228]), .Z(n755) );
  NAND U1129 ( .A(N233), .B(xregN_1), .Z(n754) );
  NAND U1130 ( .A(n756), .B(n757), .Z(z2[228]) );
  NANDN U1131 ( .A(xregN_1), .B(zin[227]), .Z(n757) );
  NAND U1132 ( .A(N232), .B(xregN_1), .Z(n756) );
  NAND U1133 ( .A(n758), .B(n759), .Z(z2[227]) );
  NANDN U1134 ( .A(xregN_1), .B(zin[226]), .Z(n759) );
  NAND U1135 ( .A(N231), .B(xregN_1), .Z(n758) );
  NAND U1136 ( .A(n760), .B(n761), .Z(z2[226]) );
  NANDN U1137 ( .A(xregN_1), .B(zin[225]), .Z(n761) );
  NAND U1138 ( .A(N230), .B(xregN_1), .Z(n760) );
  NAND U1139 ( .A(n762), .B(n763), .Z(z2[225]) );
  NANDN U1140 ( .A(xregN_1), .B(zin[224]), .Z(n763) );
  NAND U1141 ( .A(N229), .B(xregN_1), .Z(n762) );
  NAND U1142 ( .A(n764), .B(n765), .Z(z2[224]) );
  NANDN U1143 ( .A(xregN_1), .B(zin[223]), .Z(n765) );
  NAND U1144 ( .A(N228), .B(xregN_1), .Z(n764) );
  NAND U1145 ( .A(n766), .B(n767), .Z(z2[223]) );
  NANDN U1146 ( .A(xregN_1), .B(zin[222]), .Z(n767) );
  NAND U1147 ( .A(N227), .B(xregN_1), .Z(n766) );
  NAND U1148 ( .A(n768), .B(n769), .Z(z2[222]) );
  NANDN U1149 ( .A(xregN_1), .B(zin[221]), .Z(n769) );
  NAND U1150 ( .A(N226), .B(xregN_1), .Z(n768) );
  NAND U1151 ( .A(n770), .B(n771), .Z(z2[221]) );
  NANDN U1152 ( .A(xregN_1), .B(zin[220]), .Z(n771) );
  NAND U1153 ( .A(N225), .B(xregN_1), .Z(n770) );
  NAND U1154 ( .A(n772), .B(n773), .Z(z2[220]) );
  NANDN U1155 ( .A(xregN_1), .B(zin[219]), .Z(n773) );
  NAND U1156 ( .A(N224), .B(xregN_1), .Z(n772) );
  NAND U1157 ( .A(n774), .B(n775), .Z(z2[21]) );
  NANDN U1158 ( .A(xregN_1), .B(zin[20]), .Z(n775) );
  NAND U1159 ( .A(N25), .B(xregN_1), .Z(n774) );
  NAND U1160 ( .A(n776), .B(n777), .Z(z2[219]) );
  NANDN U1161 ( .A(xregN_1), .B(zin[218]), .Z(n777) );
  NAND U1162 ( .A(N223), .B(xregN_1), .Z(n776) );
  NAND U1163 ( .A(n778), .B(n779), .Z(z2[218]) );
  NANDN U1164 ( .A(xregN_1), .B(zin[217]), .Z(n779) );
  NAND U1165 ( .A(N222), .B(xregN_1), .Z(n778) );
  NAND U1166 ( .A(n780), .B(n781), .Z(z2[217]) );
  NANDN U1167 ( .A(xregN_1), .B(zin[216]), .Z(n781) );
  NAND U1168 ( .A(N221), .B(xregN_1), .Z(n780) );
  NAND U1169 ( .A(n782), .B(n783), .Z(z2[216]) );
  NANDN U1170 ( .A(xregN_1), .B(zin[215]), .Z(n783) );
  NAND U1171 ( .A(N220), .B(xregN_1), .Z(n782) );
  NAND U1172 ( .A(n784), .B(n785), .Z(z2[215]) );
  NANDN U1173 ( .A(xregN_1), .B(zin[214]), .Z(n785) );
  NAND U1174 ( .A(N219), .B(xregN_1), .Z(n784) );
  NAND U1175 ( .A(n786), .B(n787), .Z(z2[214]) );
  NANDN U1176 ( .A(xregN_1), .B(zin[213]), .Z(n787) );
  NAND U1177 ( .A(N218), .B(xregN_1), .Z(n786) );
  NAND U1178 ( .A(n788), .B(n789), .Z(z2[213]) );
  NANDN U1179 ( .A(xregN_1), .B(zin[212]), .Z(n789) );
  NAND U1180 ( .A(N217), .B(xregN_1), .Z(n788) );
  NAND U1181 ( .A(n790), .B(n791), .Z(z2[212]) );
  NANDN U1182 ( .A(xregN_1), .B(zin[211]), .Z(n791) );
  NAND U1183 ( .A(N216), .B(xregN_1), .Z(n790) );
  NAND U1184 ( .A(n792), .B(n793), .Z(z2[211]) );
  NANDN U1185 ( .A(xregN_1), .B(zin[210]), .Z(n793) );
  NAND U1186 ( .A(N215), .B(xregN_1), .Z(n792) );
  NAND U1187 ( .A(n794), .B(n795), .Z(z2[210]) );
  NANDN U1188 ( .A(xregN_1), .B(zin[209]), .Z(n795) );
  NAND U1189 ( .A(N214), .B(xregN_1), .Z(n794) );
  NAND U1190 ( .A(n796), .B(n797), .Z(z2[20]) );
  NANDN U1191 ( .A(xregN_1), .B(zin[19]), .Z(n797) );
  NAND U1192 ( .A(N24), .B(xregN_1), .Z(n796) );
  NAND U1193 ( .A(n798), .B(n799), .Z(z2[209]) );
  NANDN U1194 ( .A(xregN_1), .B(zin[208]), .Z(n799) );
  NAND U1195 ( .A(N213), .B(xregN_1), .Z(n798) );
  NAND U1196 ( .A(n800), .B(n801), .Z(z2[208]) );
  NANDN U1197 ( .A(xregN_1), .B(zin[207]), .Z(n801) );
  NAND U1198 ( .A(N212), .B(xregN_1), .Z(n800) );
  NAND U1199 ( .A(n802), .B(n803), .Z(z2[207]) );
  NANDN U1200 ( .A(xregN_1), .B(zin[206]), .Z(n803) );
  NAND U1201 ( .A(N211), .B(xregN_1), .Z(n802) );
  NAND U1202 ( .A(n804), .B(n805), .Z(z2[206]) );
  NANDN U1203 ( .A(xregN_1), .B(zin[205]), .Z(n805) );
  NAND U1204 ( .A(N210), .B(xregN_1), .Z(n804) );
  NAND U1205 ( .A(n806), .B(n807), .Z(z2[205]) );
  NANDN U1206 ( .A(xregN_1), .B(zin[204]), .Z(n807) );
  NAND U1207 ( .A(N209), .B(xregN_1), .Z(n806) );
  NAND U1208 ( .A(n808), .B(n809), .Z(z2[204]) );
  NANDN U1209 ( .A(xregN_1), .B(zin[203]), .Z(n809) );
  NAND U1210 ( .A(N208), .B(xregN_1), .Z(n808) );
  NAND U1211 ( .A(n810), .B(n811), .Z(z2[203]) );
  NANDN U1212 ( .A(xregN_1), .B(zin[202]), .Z(n811) );
  NAND U1213 ( .A(N207), .B(xregN_1), .Z(n810) );
  NAND U1214 ( .A(n812), .B(n813), .Z(z2[202]) );
  NANDN U1215 ( .A(xregN_1), .B(zin[201]), .Z(n813) );
  NAND U1216 ( .A(N206), .B(xregN_1), .Z(n812) );
  NAND U1217 ( .A(n814), .B(n815), .Z(z2[201]) );
  NANDN U1218 ( .A(xregN_1), .B(zin[200]), .Z(n815) );
  NAND U1219 ( .A(N205), .B(xregN_1), .Z(n814) );
  NAND U1220 ( .A(n816), .B(n817), .Z(z2[200]) );
  NANDN U1221 ( .A(xregN_1), .B(zin[199]), .Z(n817) );
  NAND U1222 ( .A(N204), .B(xregN_1), .Z(n816) );
  NAND U1223 ( .A(n818), .B(n819), .Z(z2[1]) );
  NANDN U1224 ( .A(xregN_1), .B(zin[0]), .Z(n819) );
  NAND U1225 ( .A(N5), .B(xregN_1), .Z(n818) );
  NAND U1226 ( .A(n820), .B(n821), .Z(z2[19]) );
  NANDN U1227 ( .A(xregN_1), .B(zin[18]), .Z(n821) );
  NAND U1228 ( .A(N23), .B(xregN_1), .Z(n820) );
  NAND U1229 ( .A(n822), .B(n823), .Z(z2[199]) );
  NANDN U1230 ( .A(xregN_1), .B(zin[198]), .Z(n823) );
  NAND U1231 ( .A(N203), .B(xregN_1), .Z(n822) );
  NAND U1232 ( .A(n824), .B(n825), .Z(z2[198]) );
  NANDN U1233 ( .A(xregN_1), .B(zin[197]), .Z(n825) );
  NAND U1234 ( .A(N202), .B(xregN_1), .Z(n824) );
  NAND U1235 ( .A(n826), .B(n827), .Z(z2[197]) );
  NANDN U1236 ( .A(xregN_1), .B(zin[196]), .Z(n827) );
  NAND U1237 ( .A(N201), .B(xregN_1), .Z(n826) );
  NAND U1238 ( .A(n828), .B(n829), .Z(z2[196]) );
  NANDN U1239 ( .A(xregN_1), .B(zin[195]), .Z(n829) );
  NAND U1240 ( .A(N200), .B(xregN_1), .Z(n828) );
  NAND U1241 ( .A(n830), .B(n831), .Z(z2[195]) );
  NANDN U1242 ( .A(xregN_1), .B(zin[194]), .Z(n831) );
  NAND U1243 ( .A(N199), .B(xregN_1), .Z(n830) );
  NAND U1244 ( .A(n832), .B(n833), .Z(z2[194]) );
  NANDN U1245 ( .A(xregN_1), .B(zin[193]), .Z(n833) );
  NAND U1246 ( .A(N198), .B(xregN_1), .Z(n832) );
  NAND U1247 ( .A(n834), .B(n835), .Z(z2[193]) );
  NANDN U1248 ( .A(xregN_1), .B(zin[192]), .Z(n835) );
  NAND U1249 ( .A(N197), .B(xregN_1), .Z(n834) );
  NAND U1250 ( .A(n836), .B(n837), .Z(z2[192]) );
  NANDN U1251 ( .A(xregN_1), .B(zin[191]), .Z(n837) );
  NAND U1252 ( .A(N196), .B(xregN_1), .Z(n836) );
  NAND U1253 ( .A(n838), .B(n839), .Z(z2[191]) );
  NANDN U1254 ( .A(xregN_1), .B(zin[190]), .Z(n839) );
  NAND U1255 ( .A(N195), .B(xregN_1), .Z(n838) );
  NAND U1256 ( .A(n840), .B(n841), .Z(z2[190]) );
  NANDN U1257 ( .A(xregN_1), .B(zin[189]), .Z(n841) );
  NAND U1258 ( .A(N194), .B(xregN_1), .Z(n840) );
  NAND U1259 ( .A(n842), .B(n843), .Z(z2[18]) );
  NANDN U1260 ( .A(xregN_1), .B(zin[17]), .Z(n843) );
  NAND U1261 ( .A(N22), .B(xregN_1), .Z(n842) );
  NAND U1262 ( .A(n844), .B(n845), .Z(z2[189]) );
  NANDN U1263 ( .A(xregN_1), .B(zin[188]), .Z(n845) );
  NAND U1264 ( .A(N193), .B(xregN_1), .Z(n844) );
  NAND U1265 ( .A(n846), .B(n847), .Z(z2[188]) );
  NANDN U1266 ( .A(xregN_1), .B(zin[187]), .Z(n847) );
  NAND U1267 ( .A(N192), .B(xregN_1), .Z(n846) );
  NAND U1268 ( .A(n848), .B(n849), .Z(z2[187]) );
  NANDN U1269 ( .A(xregN_1), .B(zin[186]), .Z(n849) );
  NAND U1270 ( .A(N191), .B(xregN_1), .Z(n848) );
  NAND U1271 ( .A(n850), .B(n851), .Z(z2[186]) );
  NANDN U1272 ( .A(xregN_1), .B(zin[185]), .Z(n851) );
  NAND U1273 ( .A(N190), .B(xregN_1), .Z(n850) );
  NAND U1274 ( .A(n852), .B(n853), .Z(z2[185]) );
  NANDN U1275 ( .A(xregN_1), .B(zin[184]), .Z(n853) );
  NAND U1276 ( .A(N189), .B(xregN_1), .Z(n852) );
  NAND U1277 ( .A(n854), .B(n855), .Z(z2[184]) );
  NANDN U1278 ( .A(xregN_1), .B(zin[183]), .Z(n855) );
  NAND U1279 ( .A(N188), .B(xregN_1), .Z(n854) );
  NAND U1280 ( .A(n856), .B(n857), .Z(z2[183]) );
  NANDN U1281 ( .A(xregN_1), .B(zin[182]), .Z(n857) );
  NAND U1282 ( .A(N187), .B(xregN_1), .Z(n856) );
  NAND U1283 ( .A(n858), .B(n859), .Z(z2[182]) );
  NANDN U1284 ( .A(xregN_1), .B(zin[181]), .Z(n859) );
  NAND U1285 ( .A(N186), .B(xregN_1), .Z(n858) );
  NAND U1286 ( .A(n860), .B(n861), .Z(z2[181]) );
  NANDN U1287 ( .A(xregN_1), .B(zin[180]), .Z(n861) );
  NAND U1288 ( .A(N185), .B(xregN_1), .Z(n860) );
  NAND U1289 ( .A(n862), .B(n863), .Z(z2[180]) );
  NANDN U1290 ( .A(xregN_1), .B(zin[179]), .Z(n863) );
  NAND U1291 ( .A(N184), .B(xregN_1), .Z(n862) );
  NAND U1292 ( .A(n864), .B(n865), .Z(z2[17]) );
  NANDN U1293 ( .A(xregN_1), .B(zin[16]), .Z(n865) );
  NAND U1294 ( .A(N21), .B(xregN_1), .Z(n864) );
  NAND U1295 ( .A(n866), .B(n867), .Z(z2[179]) );
  NANDN U1296 ( .A(xregN_1), .B(zin[178]), .Z(n867) );
  NAND U1297 ( .A(N183), .B(xregN_1), .Z(n866) );
  NAND U1298 ( .A(n868), .B(n869), .Z(z2[178]) );
  NANDN U1299 ( .A(xregN_1), .B(zin[177]), .Z(n869) );
  NAND U1300 ( .A(N182), .B(xregN_1), .Z(n868) );
  NAND U1301 ( .A(n870), .B(n871), .Z(z2[177]) );
  NANDN U1302 ( .A(xregN_1), .B(zin[176]), .Z(n871) );
  NAND U1303 ( .A(N181), .B(xregN_1), .Z(n870) );
  NAND U1304 ( .A(n872), .B(n873), .Z(z2[176]) );
  NANDN U1305 ( .A(xregN_1), .B(zin[175]), .Z(n873) );
  NAND U1306 ( .A(N180), .B(xregN_1), .Z(n872) );
  NAND U1307 ( .A(n874), .B(n875), .Z(z2[175]) );
  NANDN U1308 ( .A(xregN_1), .B(zin[174]), .Z(n875) );
  NAND U1309 ( .A(N179), .B(xregN_1), .Z(n874) );
  NAND U1310 ( .A(n876), .B(n877), .Z(z2[174]) );
  NANDN U1311 ( .A(xregN_1), .B(zin[173]), .Z(n877) );
  NAND U1312 ( .A(N178), .B(xregN_1), .Z(n876) );
  NAND U1313 ( .A(n878), .B(n879), .Z(z2[173]) );
  NANDN U1314 ( .A(xregN_1), .B(zin[172]), .Z(n879) );
  NAND U1315 ( .A(N177), .B(xregN_1), .Z(n878) );
  NAND U1316 ( .A(n880), .B(n881), .Z(z2[172]) );
  NANDN U1317 ( .A(xregN_1), .B(zin[171]), .Z(n881) );
  NAND U1318 ( .A(N176), .B(xregN_1), .Z(n880) );
  NAND U1319 ( .A(n882), .B(n883), .Z(z2[171]) );
  NANDN U1320 ( .A(xregN_1), .B(zin[170]), .Z(n883) );
  NAND U1321 ( .A(N175), .B(xregN_1), .Z(n882) );
  NAND U1322 ( .A(n884), .B(n885), .Z(z2[170]) );
  NANDN U1323 ( .A(xregN_1), .B(zin[169]), .Z(n885) );
  NAND U1324 ( .A(N174), .B(xregN_1), .Z(n884) );
  NAND U1325 ( .A(n886), .B(n887), .Z(z2[16]) );
  NANDN U1326 ( .A(xregN_1), .B(zin[15]), .Z(n887) );
  NAND U1327 ( .A(N20), .B(xregN_1), .Z(n886) );
  NAND U1328 ( .A(n888), .B(n889), .Z(z2[169]) );
  NANDN U1329 ( .A(xregN_1), .B(zin[168]), .Z(n889) );
  NAND U1330 ( .A(N173), .B(xregN_1), .Z(n888) );
  NAND U1331 ( .A(n890), .B(n891), .Z(z2[168]) );
  NANDN U1332 ( .A(xregN_1), .B(zin[167]), .Z(n891) );
  NAND U1333 ( .A(N172), .B(xregN_1), .Z(n890) );
  NAND U1334 ( .A(n892), .B(n893), .Z(z2[167]) );
  NANDN U1335 ( .A(xregN_1), .B(zin[166]), .Z(n893) );
  NAND U1336 ( .A(N171), .B(xregN_1), .Z(n892) );
  NAND U1337 ( .A(n894), .B(n895), .Z(z2[166]) );
  NANDN U1338 ( .A(xregN_1), .B(zin[165]), .Z(n895) );
  NAND U1339 ( .A(N170), .B(xregN_1), .Z(n894) );
  NAND U1340 ( .A(n896), .B(n897), .Z(z2[165]) );
  NANDN U1341 ( .A(xregN_1), .B(zin[164]), .Z(n897) );
  NAND U1342 ( .A(N169), .B(xregN_1), .Z(n896) );
  NAND U1343 ( .A(n898), .B(n899), .Z(z2[164]) );
  NANDN U1344 ( .A(xregN_1), .B(zin[163]), .Z(n899) );
  NAND U1345 ( .A(N168), .B(xregN_1), .Z(n898) );
  NAND U1346 ( .A(n900), .B(n901), .Z(z2[163]) );
  NANDN U1347 ( .A(xregN_1), .B(zin[162]), .Z(n901) );
  NAND U1348 ( .A(N167), .B(xregN_1), .Z(n900) );
  NAND U1349 ( .A(n902), .B(n903), .Z(z2[162]) );
  NANDN U1350 ( .A(xregN_1), .B(zin[161]), .Z(n903) );
  NAND U1351 ( .A(N166), .B(xregN_1), .Z(n902) );
  NAND U1352 ( .A(n904), .B(n905), .Z(z2[161]) );
  NANDN U1353 ( .A(xregN_1), .B(zin[160]), .Z(n905) );
  NAND U1354 ( .A(N165), .B(xregN_1), .Z(n904) );
  NAND U1355 ( .A(n906), .B(n907), .Z(z2[160]) );
  NANDN U1356 ( .A(xregN_1), .B(zin[159]), .Z(n907) );
  NAND U1357 ( .A(N164), .B(xregN_1), .Z(n906) );
  NAND U1358 ( .A(n908), .B(n909), .Z(z2[15]) );
  NANDN U1359 ( .A(xregN_1), .B(zin[14]), .Z(n909) );
  NAND U1360 ( .A(N19), .B(xregN_1), .Z(n908) );
  NAND U1361 ( .A(n910), .B(n911), .Z(z2[159]) );
  NANDN U1362 ( .A(xregN_1), .B(zin[158]), .Z(n911) );
  NAND U1363 ( .A(N163), .B(xregN_1), .Z(n910) );
  NAND U1364 ( .A(n912), .B(n913), .Z(z2[158]) );
  NANDN U1365 ( .A(xregN_1), .B(zin[157]), .Z(n913) );
  NAND U1366 ( .A(N162), .B(xregN_1), .Z(n912) );
  NAND U1367 ( .A(n914), .B(n915), .Z(z2[157]) );
  NANDN U1368 ( .A(xregN_1), .B(zin[156]), .Z(n915) );
  NAND U1369 ( .A(N161), .B(xregN_1), .Z(n914) );
  NAND U1370 ( .A(n916), .B(n917), .Z(z2[156]) );
  NANDN U1371 ( .A(xregN_1), .B(zin[155]), .Z(n917) );
  NAND U1372 ( .A(N160), .B(xregN_1), .Z(n916) );
  NAND U1373 ( .A(n918), .B(n919), .Z(z2[155]) );
  NANDN U1374 ( .A(xregN_1), .B(zin[154]), .Z(n919) );
  NAND U1375 ( .A(N159), .B(xregN_1), .Z(n918) );
  NAND U1376 ( .A(n920), .B(n921), .Z(z2[154]) );
  NANDN U1377 ( .A(xregN_1), .B(zin[153]), .Z(n921) );
  NAND U1378 ( .A(N158), .B(xregN_1), .Z(n920) );
  NAND U1379 ( .A(n922), .B(n923), .Z(z2[153]) );
  NANDN U1380 ( .A(xregN_1), .B(zin[152]), .Z(n923) );
  NAND U1381 ( .A(N157), .B(xregN_1), .Z(n922) );
  NAND U1382 ( .A(n924), .B(n925), .Z(z2[152]) );
  NANDN U1383 ( .A(xregN_1), .B(zin[151]), .Z(n925) );
  NAND U1384 ( .A(N156), .B(xregN_1), .Z(n924) );
  NAND U1385 ( .A(n926), .B(n927), .Z(z2[151]) );
  NANDN U1386 ( .A(xregN_1), .B(zin[150]), .Z(n927) );
  NAND U1387 ( .A(N155), .B(xregN_1), .Z(n926) );
  NAND U1388 ( .A(n928), .B(n929), .Z(z2[150]) );
  NANDN U1389 ( .A(xregN_1), .B(zin[149]), .Z(n929) );
  NAND U1390 ( .A(N154), .B(xregN_1), .Z(n928) );
  NAND U1391 ( .A(n930), .B(n931), .Z(z2[14]) );
  NANDN U1392 ( .A(xregN_1), .B(zin[13]), .Z(n931) );
  NAND U1393 ( .A(N18), .B(xregN_1), .Z(n930) );
  NAND U1394 ( .A(n932), .B(n933), .Z(z2[149]) );
  NANDN U1395 ( .A(xregN_1), .B(zin[148]), .Z(n933) );
  NAND U1396 ( .A(N153), .B(xregN_1), .Z(n932) );
  NAND U1397 ( .A(n934), .B(n935), .Z(z2[148]) );
  NANDN U1398 ( .A(xregN_1), .B(zin[147]), .Z(n935) );
  NAND U1399 ( .A(N152), .B(xregN_1), .Z(n934) );
  NAND U1400 ( .A(n936), .B(n937), .Z(z2[147]) );
  NANDN U1401 ( .A(xregN_1), .B(zin[146]), .Z(n937) );
  NAND U1402 ( .A(N151), .B(xregN_1), .Z(n936) );
  NAND U1403 ( .A(n938), .B(n939), .Z(z2[146]) );
  NANDN U1404 ( .A(xregN_1), .B(zin[145]), .Z(n939) );
  NAND U1405 ( .A(N150), .B(xregN_1), .Z(n938) );
  NAND U1406 ( .A(n940), .B(n941), .Z(z2[145]) );
  NANDN U1407 ( .A(xregN_1), .B(zin[144]), .Z(n941) );
  NAND U1408 ( .A(N149), .B(xregN_1), .Z(n940) );
  NAND U1409 ( .A(n942), .B(n943), .Z(z2[144]) );
  NANDN U1410 ( .A(xregN_1), .B(zin[143]), .Z(n943) );
  NAND U1411 ( .A(N148), .B(xregN_1), .Z(n942) );
  NAND U1412 ( .A(n944), .B(n945), .Z(z2[143]) );
  NANDN U1413 ( .A(xregN_1), .B(zin[142]), .Z(n945) );
  NAND U1414 ( .A(N147), .B(xregN_1), .Z(n944) );
  NAND U1415 ( .A(n946), .B(n947), .Z(z2[142]) );
  NANDN U1416 ( .A(xregN_1), .B(zin[141]), .Z(n947) );
  NAND U1417 ( .A(N146), .B(xregN_1), .Z(n946) );
  NAND U1418 ( .A(n948), .B(n949), .Z(z2[141]) );
  NANDN U1419 ( .A(xregN_1), .B(zin[140]), .Z(n949) );
  NAND U1420 ( .A(N145), .B(xregN_1), .Z(n948) );
  NAND U1421 ( .A(n950), .B(n951), .Z(z2[140]) );
  NANDN U1422 ( .A(xregN_1), .B(zin[139]), .Z(n951) );
  NAND U1423 ( .A(N144), .B(xregN_1), .Z(n950) );
  NAND U1424 ( .A(n952), .B(n953), .Z(z2[13]) );
  NANDN U1425 ( .A(xregN_1), .B(zin[12]), .Z(n953) );
  NAND U1426 ( .A(N17), .B(xregN_1), .Z(n952) );
  NAND U1427 ( .A(n954), .B(n955), .Z(z2[139]) );
  NANDN U1428 ( .A(xregN_1), .B(zin[138]), .Z(n955) );
  NAND U1429 ( .A(N143), .B(xregN_1), .Z(n954) );
  NAND U1430 ( .A(n956), .B(n957), .Z(z2[138]) );
  NANDN U1431 ( .A(xregN_1), .B(zin[137]), .Z(n957) );
  NAND U1432 ( .A(N142), .B(xregN_1), .Z(n956) );
  NAND U1433 ( .A(n958), .B(n959), .Z(z2[137]) );
  NANDN U1434 ( .A(xregN_1), .B(zin[136]), .Z(n959) );
  NAND U1435 ( .A(N141), .B(xregN_1), .Z(n958) );
  NAND U1436 ( .A(n960), .B(n961), .Z(z2[136]) );
  NANDN U1437 ( .A(xregN_1), .B(zin[135]), .Z(n961) );
  NAND U1438 ( .A(N140), .B(xregN_1), .Z(n960) );
  NAND U1439 ( .A(n962), .B(n963), .Z(z2[135]) );
  NANDN U1440 ( .A(xregN_1), .B(zin[134]), .Z(n963) );
  NAND U1441 ( .A(N139), .B(xregN_1), .Z(n962) );
  NAND U1442 ( .A(n964), .B(n965), .Z(z2[134]) );
  NANDN U1443 ( .A(xregN_1), .B(zin[133]), .Z(n965) );
  NAND U1444 ( .A(N138), .B(xregN_1), .Z(n964) );
  NAND U1445 ( .A(n966), .B(n967), .Z(z2[133]) );
  NANDN U1446 ( .A(xregN_1), .B(zin[132]), .Z(n967) );
  NAND U1447 ( .A(N137), .B(xregN_1), .Z(n966) );
  NAND U1448 ( .A(n968), .B(n969), .Z(z2[132]) );
  NANDN U1449 ( .A(xregN_1), .B(zin[131]), .Z(n969) );
  NAND U1450 ( .A(N136), .B(xregN_1), .Z(n968) );
  NAND U1451 ( .A(n970), .B(n971), .Z(z2[131]) );
  NANDN U1452 ( .A(xregN_1), .B(zin[130]), .Z(n971) );
  NAND U1453 ( .A(N135), .B(xregN_1), .Z(n970) );
  NAND U1454 ( .A(n972), .B(n973), .Z(z2[130]) );
  NANDN U1455 ( .A(xregN_1), .B(zin[129]), .Z(n973) );
  NAND U1456 ( .A(N134), .B(xregN_1), .Z(n972) );
  NAND U1457 ( .A(n974), .B(n975), .Z(z2[12]) );
  NANDN U1458 ( .A(xregN_1), .B(zin[11]), .Z(n975) );
  NAND U1459 ( .A(N16), .B(xregN_1), .Z(n974) );
  NAND U1460 ( .A(n976), .B(n977), .Z(z2[129]) );
  NANDN U1461 ( .A(xregN_1), .B(zin[128]), .Z(n977) );
  NAND U1462 ( .A(N133), .B(xregN_1), .Z(n976) );
  NAND U1463 ( .A(n978), .B(n979), .Z(z2[128]) );
  NANDN U1464 ( .A(xregN_1), .B(zin[127]), .Z(n979) );
  NAND U1465 ( .A(N132), .B(xregN_1), .Z(n978) );
  NAND U1466 ( .A(n980), .B(n981), .Z(z2[127]) );
  NANDN U1467 ( .A(xregN_1), .B(zin[126]), .Z(n981) );
  NAND U1468 ( .A(N131), .B(xregN_1), .Z(n980) );
  NAND U1469 ( .A(n982), .B(n983), .Z(z2[126]) );
  NANDN U1470 ( .A(xregN_1), .B(zin[125]), .Z(n983) );
  NAND U1471 ( .A(N130), .B(xregN_1), .Z(n982) );
  NAND U1472 ( .A(n984), .B(n985), .Z(z2[125]) );
  NANDN U1473 ( .A(xregN_1), .B(zin[124]), .Z(n985) );
  NAND U1474 ( .A(N129), .B(xregN_1), .Z(n984) );
  NAND U1475 ( .A(n986), .B(n987), .Z(z2[124]) );
  NANDN U1476 ( .A(xregN_1), .B(zin[123]), .Z(n987) );
  NAND U1477 ( .A(N128), .B(xregN_1), .Z(n986) );
  NAND U1478 ( .A(n988), .B(n989), .Z(z2[123]) );
  NANDN U1479 ( .A(xregN_1), .B(zin[122]), .Z(n989) );
  NAND U1480 ( .A(N127), .B(xregN_1), .Z(n988) );
  NAND U1481 ( .A(n990), .B(n991), .Z(z2[122]) );
  NANDN U1482 ( .A(xregN_1), .B(zin[121]), .Z(n991) );
  NAND U1483 ( .A(N126), .B(xregN_1), .Z(n990) );
  NAND U1484 ( .A(n992), .B(n993), .Z(z2[121]) );
  NANDN U1485 ( .A(xregN_1), .B(zin[120]), .Z(n993) );
  NAND U1486 ( .A(N125), .B(xregN_1), .Z(n992) );
  NAND U1487 ( .A(n994), .B(n995), .Z(z2[120]) );
  NANDN U1488 ( .A(xregN_1), .B(zin[119]), .Z(n995) );
  NAND U1489 ( .A(N124), .B(xregN_1), .Z(n994) );
  NAND U1490 ( .A(n996), .B(n997), .Z(z2[11]) );
  NANDN U1491 ( .A(xregN_1), .B(zin[10]), .Z(n997) );
  NAND U1492 ( .A(N15), .B(xregN_1), .Z(n996) );
  NAND U1493 ( .A(n998), .B(n999), .Z(z2[119]) );
  NANDN U1494 ( .A(xregN_1), .B(zin[118]), .Z(n999) );
  NAND U1495 ( .A(N123), .B(xregN_1), .Z(n998) );
  NAND U1496 ( .A(n1000), .B(n1001), .Z(z2[118]) );
  NANDN U1497 ( .A(xregN_1), .B(zin[117]), .Z(n1001) );
  NAND U1498 ( .A(N122), .B(xregN_1), .Z(n1000) );
  NAND U1499 ( .A(n1002), .B(n1003), .Z(z2[117]) );
  NANDN U1500 ( .A(xregN_1), .B(zin[116]), .Z(n1003) );
  NAND U1501 ( .A(N121), .B(xregN_1), .Z(n1002) );
  NAND U1502 ( .A(n1004), .B(n1005), .Z(z2[116]) );
  NANDN U1503 ( .A(xregN_1), .B(zin[115]), .Z(n1005) );
  NAND U1504 ( .A(N120), .B(xregN_1), .Z(n1004) );
  NAND U1505 ( .A(n1006), .B(n1007), .Z(z2[115]) );
  NANDN U1506 ( .A(xregN_1), .B(zin[114]), .Z(n1007) );
  NAND U1507 ( .A(N119), .B(xregN_1), .Z(n1006) );
  NAND U1508 ( .A(n1008), .B(n1009), .Z(z2[114]) );
  NANDN U1509 ( .A(xregN_1), .B(zin[113]), .Z(n1009) );
  NAND U1510 ( .A(N118), .B(xregN_1), .Z(n1008) );
  NAND U1511 ( .A(n1010), .B(n1011), .Z(z2[113]) );
  NANDN U1512 ( .A(xregN_1), .B(zin[112]), .Z(n1011) );
  NAND U1513 ( .A(N117), .B(xregN_1), .Z(n1010) );
  NAND U1514 ( .A(n1012), .B(n1013), .Z(z2[112]) );
  NANDN U1515 ( .A(xregN_1), .B(zin[111]), .Z(n1013) );
  NAND U1516 ( .A(N116), .B(xregN_1), .Z(n1012) );
  NAND U1517 ( .A(n1014), .B(n1015), .Z(z2[111]) );
  NANDN U1518 ( .A(xregN_1), .B(zin[110]), .Z(n1015) );
  NAND U1519 ( .A(N115), .B(xregN_1), .Z(n1014) );
  NAND U1520 ( .A(n1016), .B(n1017), .Z(z2[110]) );
  NANDN U1521 ( .A(xregN_1), .B(zin[109]), .Z(n1017) );
  NAND U1522 ( .A(N114), .B(xregN_1), .Z(n1016) );
  NAND U1523 ( .A(n1018), .B(n1019), .Z(z2[10]) );
  NANDN U1524 ( .A(xregN_1), .B(zin[9]), .Z(n1019) );
  NAND U1525 ( .A(N14), .B(xregN_1), .Z(n1018) );
  NAND U1526 ( .A(n1020), .B(n1021), .Z(z2[109]) );
  NANDN U1527 ( .A(xregN_1), .B(zin[108]), .Z(n1021) );
  NAND U1528 ( .A(N113), .B(xregN_1), .Z(n1020) );
  NAND U1529 ( .A(n1022), .B(n1023), .Z(z2[108]) );
  NANDN U1530 ( .A(xregN_1), .B(zin[107]), .Z(n1023) );
  NAND U1531 ( .A(N112), .B(xregN_1), .Z(n1022) );
  NAND U1532 ( .A(n1024), .B(n1025), .Z(z2[107]) );
  NANDN U1533 ( .A(xregN_1), .B(zin[106]), .Z(n1025) );
  NAND U1534 ( .A(N111), .B(xregN_1), .Z(n1024) );
  NAND U1535 ( .A(n1026), .B(n1027), .Z(z2[106]) );
  NANDN U1536 ( .A(xregN_1), .B(zin[105]), .Z(n1027) );
  NAND U1537 ( .A(N110), .B(xregN_1), .Z(n1026) );
  NAND U1538 ( .A(n1028), .B(n1029), .Z(z2[105]) );
  NANDN U1539 ( .A(xregN_1), .B(zin[104]), .Z(n1029) );
  NAND U1540 ( .A(N109), .B(xregN_1), .Z(n1028) );
  NAND U1541 ( .A(n1030), .B(n1031), .Z(z2[104]) );
  NANDN U1542 ( .A(xregN_1), .B(zin[103]), .Z(n1031) );
  NAND U1543 ( .A(N108), .B(xregN_1), .Z(n1030) );
  NAND U1544 ( .A(n1032), .B(n1033), .Z(z2[103]) );
  NANDN U1545 ( .A(xregN_1), .B(zin[102]), .Z(n1033) );
  NAND U1546 ( .A(N107), .B(xregN_1), .Z(n1032) );
  NAND U1547 ( .A(n1034), .B(n1035), .Z(z2[102]) );
  NANDN U1548 ( .A(xregN_1), .B(zin[101]), .Z(n1035) );
  NAND U1549 ( .A(N106), .B(xregN_1), .Z(n1034) );
  NAND U1550 ( .A(n1036), .B(n1037), .Z(z2[101]) );
  NANDN U1551 ( .A(xregN_1), .B(zin[100]), .Z(n1037) );
  NAND U1552 ( .A(N105), .B(xregN_1), .Z(n1036) );
  NAND U1553 ( .A(n1038), .B(n1039), .Z(z2[100]) );
  NANDN U1554 ( .A(xregN_1), .B(zin[99]), .Z(n1039) );
  NAND U1555 ( .A(N104), .B(xregN_1), .Z(n1038) );
  AND U1556 ( .A(N4), .B(xregN_1), .Z(z2[0]) );
endmodule


module modmult_N256_CC64 ( clk, rst, start, x, y, n, o );
  input [255:0] x;
  input [255:0] y;
  input [255:0] n;
  output [255:0] o;
  input clk, rst, start;
  wire   \zout[3][257] , \zout[3][256] , \zin[3][257] , \zin[3][256] ,
         \zin[3][255] , \zin[3][254] , \zin[3][253] , \zin[3][252] ,
         \zin[3][251] , \zin[3][250] , \zin[3][249] , \zin[3][248] ,
         \zin[3][247] , \zin[3][246] , \zin[3][245] , \zin[3][244] ,
         \zin[3][243] , \zin[3][242] , \zin[3][241] , \zin[3][240] ,
         \zin[3][239] , \zin[3][238] , \zin[3][237] , \zin[3][236] ,
         \zin[3][235] , \zin[3][234] , \zin[3][233] , \zin[3][232] ,
         \zin[3][231] , \zin[3][230] , \zin[3][229] , \zin[3][228] ,
         \zin[3][227] , \zin[3][226] , \zin[3][225] , \zin[3][224] ,
         \zin[3][223] , \zin[3][222] , \zin[3][221] , \zin[3][220] ,
         \zin[3][219] , \zin[3][218] , \zin[3][217] , \zin[3][216] ,
         \zin[3][215] , \zin[3][214] , \zin[3][213] , \zin[3][212] ,
         \zin[3][211] , \zin[3][210] , \zin[3][209] , \zin[3][208] ,
         \zin[3][207] , \zin[3][206] , \zin[3][205] , \zin[3][204] ,
         \zin[3][203] , \zin[3][202] , \zin[3][201] , \zin[3][200] ,
         \zin[3][199] , \zin[3][198] , \zin[3][197] , \zin[3][196] ,
         \zin[3][195] , \zin[3][194] , \zin[3][193] , \zin[3][192] ,
         \zin[3][191] , \zin[3][190] , \zin[3][189] , \zin[3][188] ,
         \zin[3][187] , \zin[3][186] , \zin[3][185] , \zin[3][184] ,
         \zin[3][183] , \zin[3][182] , \zin[3][181] , \zin[3][180] ,
         \zin[3][179] , \zin[3][178] , \zin[3][177] , \zin[3][176] ,
         \zin[3][175] , \zin[3][174] , \zin[3][173] , \zin[3][172] ,
         \zin[3][171] , \zin[3][170] , \zin[3][169] , \zin[3][168] ,
         \zin[3][167] , \zin[3][166] , \zin[3][165] , \zin[3][164] ,
         \zin[3][163] , \zin[3][162] , \zin[3][161] , \zin[3][160] ,
         \zin[3][159] , \zin[3][158] , \zin[3][157] , \zin[3][156] ,
         \zin[3][155] , \zin[3][154] , \zin[3][153] , \zin[3][152] ,
         \zin[3][151] , \zin[3][150] , \zin[3][149] , \zin[3][148] ,
         \zin[3][147] , \zin[3][146] , \zin[3][145] , \zin[3][144] ,
         \zin[3][143] , \zin[3][142] , \zin[3][141] , \zin[3][140] ,
         \zin[3][139] , \zin[3][138] , \zin[3][137] , \zin[3][136] ,
         \zin[3][135] , \zin[3][134] , \zin[3][133] , \zin[3][132] ,
         \zin[3][131] , \zin[3][130] , \zin[3][129] , \zin[3][128] ,
         \zin[3][127] , \zin[3][126] , \zin[3][125] , \zin[3][124] ,
         \zin[3][123] , \zin[3][122] , \zin[3][121] , \zin[3][120] ,
         \zin[3][119] , \zin[3][118] , \zin[3][117] , \zin[3][116] ,
         \zin[3][115] , \zin[3][114] , \zin[3][113] , \zin[3][112] ,
         \zin[3][111] , \zin[3][110] , \zin[3][109] , \zin[3][108] ,
         \zin[3][107] , \zin[3][106] , \zin[3][105] , \zin[3][104] ,
         \zin[3][103] , \zin[3][102] , \zin[3][101] , \zin[3][100] ,
         \zin[3][99] , \zin[3][98] , \zin[3][97] , \zin[3][96] , \zin[3][95] ,
         \zin[3][94] , \zin[3][93] , \zin[3][92] , \zin[3][91] , \zin[3][90] ,
         \zin[3][89] , \zin[3][88] , \zin[3][87] , \zin[3][86] , \zin[3][85] ,
         \zin[3][84] , \zin[3][83] , \zin[3][82] , \zin[3][81] , \zin[3][80] ,
         \zin[3][79] , \zin[3][78] , \zin[3][77] , \zin[3][76] , \zin[3][75] ,
         \zin[3][74] , \zin[3][73] , \zin[3][72] , \zin[3][71] , \zin[3][70] ,
         \zin[3][69] , \zin[3][68] , \zin[3][67] , \zin[3][66] , \zin[3][65] ,
         \zin[3][64] , \zin[3][63] , \zin[3][62] , \zin[3][61] , \zin[3][60] ,
         \zin[3][59] , \zin[3][58] , \zin[3][57] , \zin[3][56] , \zin[3][55] ,
         \zin[3][54] , \zin[3][53] , \zin[3][52] , \zin[3][51] , \zin[3][50] ,
         \zin[3][49] , \zin[3][48] , \zin[3][47] , \zin[3][46] , \zin[3][45] ,
         \zin[3][44] , \zin[3][43] , \zin[3][42] , \zin[3][41] , \zin[3][40] ,
         \zin[3][39] , \zin[3][38] , \zin[3][37] , \zin[3][36] , \zin[3][35] ,
         \zin[3][34] , \zin[3][33] , \zin[3][32] , \zin[3][31] , \zin[3][30] ,
         \zin[3][29] , \zin[3][28] , \zin[3][27] , \zin[3][26] , \zin[3][25] ,
         \zin[3][24] , \zin[3][23] , \zin[3][22] , \zin[3][21] , \zin[3][20] ,
         \zin[3][19] , \zin[3][18] , \zin[3][17] , \zin[3][16] , \zin[3][15] ,
         \zin[3][14] , \zin[3][13] , \zin[3][12] , \zin[3][11] , \zin[3][10] ,
         \zin[3][9] , \zin[3][8] , \zin[3][7] , \zin[3][6] , \zin[3][5] ,
         \zin[3][4] , \zin[3][3] , \zin[3][2] , \zin[3][1] , \zin[3][0] ,
         \zin[2][257] , \zin[2][256] , \zin[2][255] , \zin[2][254] ,
         \zin[2][253] , \zin[2][252] , \zin[2][251] , \zin[2][250] ,
         \zin[2][249] , \zin[2][248] , \zin[2][247] , \zin[2][246] ,
         \zin[2][245] , \zin[2][244] , \zin[2][243] , \zin[2][242] ,
         \zin[2][241] , \zin[2][240] , \zin[2][239] , \zin[2][238] ,
         \zin[2][237] , \zin[2][236] , \zin[2][235] , \zin[2][234] ,
         \zin[2][233] , \zin[2][232] , \zin[2][231] , \zin[2][230] ,
         \zin[2][229] , \zin[2][228] , \zin[2][227] , \zin[2][226] ,
         \zin[2][225] , \zin[2][224] , \zin[2][223] , \zin[2][222] ,
         \zin[2][221] , \zin[2][220] , \zin[2][219] , \zin[2][218] ,
         \zin[2][217] , \zin[2][216] , \zin[2][215] , \zin[2][214] ,
         \zin[2][213] , \zin[2][212] , \zin[2][211] , \zin[2][210] ,
         \zin[2][209] , \zin[2][208] , \zin[2][207] , \zin[2][206] ,
         \zin[2][205] , \zin[2][204] , \zin[2][203] , \zin[2][202] ,
         \zin[2][201] , \zin[2][200] , \zin[2][199] , \zin[2][198] ,
         \zin[2][197] , \zin[2][196] , \zin[2][195] , \zin[2][194] ,
         \zin[2][193] , \zin[2][192] , \zin[2][191] , \zin[2][190] ,
         \zin[2][189] , \zin[2][188] , \zin[2][187] , \zin[2][186] ,
         \zin[2][185] , \zin[2][184] , \zin[2][183] , \zin[2][182] ,
         \zin[2][181] , \zin[2][180] , \zin[2][179] , \zin[2][178] ,
         \zin[2][177] , \zin[2][176] , \zin[2][175] , \zin[2][174] ,
         \zin[2][173] , \zin[2][172] , \zin[2][171] , \zin[2][170] ,
         \zin[2][169] , \zin[2][168] , \zin[2][167] , \zin[2][166] ,
         \zin[2][165] , \zin[2][164] , \zin[2][163] , \zin[2][162] ,
         \zin[2][161] , \zin[2][160] , \zin[2][159] , \zin[2][158] ,
         \zin[2][157] , \zin[2][156] , \zin[2][155] , \zin[2][154] ,
         \zin[2][153] , \zin[2][152] , \zin[2][151] , \zin[2][150] ,
         \zin[2][149] , \zin[2][148] , \zin[2][147] , \zin[2][146] ,
         \zin[2][145] , \zin[2][144] , \zin[2][143] , \zin[2][142] ,
         \zin[2][141] , \zin[2][140] , \zin[2][139] , \zin[2][138] ,
         \zin[2][137] , \zin[2][136] , \zin[2][135] , \zin[2][134] ,
         \zin[2][133] , \zin[2][132] , \zin[2][131] , \zin[2][130] ,
         \zin[2][129] , \zin[2][128] , \zin[2][127] , \zin[2][126] ,
         \zin[2][125] , \zin[2][124] , \zin[2][123] , \zin[2][122] ,
         \zin[2][121] , \zin[2][120] , \zin[2][119] , \zin[2][118] ,
         \zin[2][117] , \zin[2][116] , \zin[2][115] , \zin[2][114] ,
         \zin[2][113] , \zin[2][112] , \zin[2][111] , \zin[2][110] ,
         \zin[2][109] , \zin[2][108] , \zin[2][107] , \zin[2][106] ,
         \zin[2][105] , \zin[2][104] , \zin[2][103] , \zin[2][102] ,
         \zin[2][101] , \zin[2][100] , \zin[2][99] , \zin[2][98] ,
         \zin[2][97] , \zin[2][96] , \zin[2][95] , \zin[2][94] , \zin[2][93] ,
         \zin[2][92] , \zin[2][91] , \zin[2][90] , \zin[2][89] , \zin[2][88] ,
         \zin[2][87] , \zin[2][86] , \zin[2][85] , \zin[2][84] , \zin[2][83] ,
         \zin[2][82] , \zin[2][81] , \zin[2][80] , \zin[2][79] , \zin[2][78] ,
         \zin[2][77] , \zin[2][76] , \zin[2][75] , \zin[2][74] , \zin[2][73] ,
         \zin[2][72] , \zin[2][71] , \zin[2][70] , \zin[2][69] , \zin[2][68] ,
         \zin[2][67] , \zin[2][66] , \zin[2][65] , \zin[2][64] , \zin[2][63] ,
         \zin[2][62] , \zin[2][61] , \zin[2][60] , \zin[2][59] , \zin[2][58] ,
         \zin[2][57] , \zin[2][56] , \zin[2][55] , \zin[2][54] , \zin[2][53] ,
         \zin[2][52] , \zin[2][51] , \zin[2][50] , \zin[2][49] , \zin[2][48] ,
         \zin[2][47] , \zin[2][46] , \zin[2][45] , \zin[2][44] , \zin[2][43] ,
         \zin[2][42] , \zin[2][41] , \zin[2][40] , \zin[2][39] , \zin[2][38] ,
         \zin[2][37] , \zin[2][36] , \zin[2][35] , \zin[2][34] , \zin[2][33] ,
         \zin[2][32] , \zin[2][31] , \zin[2][30] , \zin[2][29] , \zin[2][28] ,
         \zin[2][27] , \zin[2][26] , \zin[2][25] , \zin[2][24] , \zin[2][23] ,
         \zin[2][22] , \zin[2][21] , \zin[2][20] , \zin[2][19] , \zin[2][18] ,
         \zin[2][17] , \zin[2][16] , \zin[2][15] , \zin[2][14] , \zin[2][13] ,
         \zin[2][12] , \zin[2][11] , \zin[2][10] , \zin[2][9] , \zin[2][8] ,
         \zin[2][7] , \zin[2][6] , \zin[2][5] , \zin[2][4] , \zin[2][3] ,
         \zin[2][2] , \zin[2][1] , \zin[2][0] , \zin[1][257] , \zin[1][256] ,
         \zin[1][255] , \zin[1][254] , \zin[1][253] , \zin[1][252] ,
         \zin[1][251] , \zin[1][250] , \zin[1][249] , \zin[1][248] ,
         \zin[1][247] , \zin[1][246] , \zin[1][245] , \zin[1][244] ,
         \zin[1][243] , \zin[1][242] , \zin[1][241] , \zin[1][240] ,
         \zin[1][239] , \zin[1][238] , \zin[1][237] , \zin[1][236] ,
         \zin[1][235] , \zin[1][234] , \zin[1][233] , \zin[1][232] ,
         \zin[1][231] , \zin[1][230] , \zin[1][229] , \zin[1][228] ,
         \zin[1][227] , \zin[1][226] , \zin[1][225] , \zin[1][224] ,
         \zin[1][223] , \zin[1][222] , \zin[1][221] , \zin[1][220] ,
         \zin[1][219] , \zin[1][218] , \zin[1][217] , \zin[1][216] ,
         \zin[1][215] , \zin[1][214] , \zin[1][213] , \zin[1][212] ,
         \zin[1][211] , \zin[1][210] , \zin[1][209] , \zin[1][208] ,
         \zin[1][207] , \zin[1][206] , \zin[1][205] , \zin[1][204] ,
         \zin[1][203] , \zin[1][202] , \zin[1][201] , \zin[1][200] ,
         \zin[1][199] , \zin[1][198] , \zin[1][197] , \zin[1][196] ,
         \zin[1][195] , \zin[1][194] , \zin[1][193] , \zin[1][192] ,
         \zin[1][191] , \zin[1][190] , \zin[1][189] , \zin[1][188] ,
         \zin[1][187] , \zin[1][186] , \zin[1][185] , \zin[1][184] ,
         \zin[1][183] , \zin[1][182] , \zin[1][181] , \zin[1][180] ,
         \zin[1][179] , \zin[1][178] , \zin[1][177] , \zin[1][176] ,
         \zin[1][175] , \zin[1][174] , \zin[1][173] , \zin[1][172] ,
         \zin[1][171] , \zin[1][170] , \zin[1][169] , \zin[1][168] ,
         \zin[1][167] , \zin[1][166] , \zin[1][165] , \zin[1][164] ,
         \zin[1][163] , \zin[1][162] , \zin[1][161] , \zin[1][160] ,
         \zin[1][159] , \zin[1][158] , \zin[1][157] , \zin[1][156] ,
         \zin[1][155] , \zin[1][154] , \zin[1][153] , \zin[1][152] ,
         \zin[1][151] , \zin[1][150] , \zin[1][149] , \zin[1][148] ,
         \zin[1][147] , \zin[1][146] , \zin[1][145] , \zin[1][144] ,
         \zin[1][143] , \zin[1][142] , \zin[1][141] , \zin[1][140] ,
         \zin[1][139] , \zin[1][138] , \zin[1][137] , \zin[1][136] ,
         \zin[1][135] , \zin[1][134] , \zin[1][133] , \zin[1][132] ,
         \zin[1][131] , \zin[1][130] , \zin[1][129] , \zin[1][128] ,
         \zin[1][127] , \zin[1][126] , \zin[1][125] , \zin[1][124] ,
         \zin[1][123] , \zin[1][122] , \zin[1][121] , \zin[1][120] ,
         \zin[1][119] , \zin[1][118] , \zin[1][117] , \zin[1][116] ,
         \zin[1][115] , \zin[1][114] , \zin[1][113] , \zin[1][112] ,
         \zin[1][111] , \zin[1][110] , \zin[1][109] , \zin[1][108] ,
         \zin[1][107] , \zin[1][106] , \zin[1][105] , \zin[1][104] ,
         \zin[1][103] , \zin[1][102] , \zin[1][101] , \zin[1][100] ,
         \zin[1][99] , \zin[1][98] , \zin[1][97] , \zin[1][96] , \zin[1][95] ,
         \zin[1][94] , \zin[1][93] , \zin[1][92] , \zin[1][91] , \zin[1][90] ,
         \zin[1][89] , \zin[1][88] , \zin[1][87] , \zin[1][86] , \zin[1][85] ,
         \zin[1][84] , \zin[1][83] , \zin[1][82] , \zin[1][81] , \zin[1][80] ,
         \zin[1][79] , \zin[1][78] , \zin[1][77] , \zin[1][76] , \zin[1][75] ,
         \zin[1][74] , \zin[1][73] , \zin[1][72] , \zin[1][71] , \zin[1][70] ,
         \zin[1][69] , \zin[1][68] , \zin[1][67] , \zin[1][66] , \zin[1][65] ,
         \zin[1][64] , \zin[1][63] , \zin[1][62] , \zin[1][61] , \zin[1][60] ,
         \zin[1][59] , \zin[1][58] , \zin[1][57] , \zin[1][56] , \zin[1][55] ,
         \zin[1][54] , \zin[1][53] , \zin[1][52] , \zin[1][51] , \zin[1][50] ,
         \zin[1][49] , \zin[1][48] , \zin[1][47] , \zin[1][46] , \zin[1][45] ,
         \zin[1][44] , \zin[1][43] , \zin[1][42] , \zin[1][41] , \zin[1][40] ,
         \zin[1][39] , \zin[1][38] , \zin[1][37] , \zin[1][36] , \zin[1][35] ,
         \zin[1][34] , \zin[1][33] , \zin[1][32] , \zin[1][31] , \zin[1][30] ,
         \zin[1][29] , \zin[1][28] , \zin[1][27] , \zin[1][26] , \zin[1][25] ,
         \zin[1][24] , \zin[1][23] , \zin[1][22] , \zin[1][21] , \zin[1][20] ,
         \zin[1][19] , \zin[1][18] , \zin[1][17] , \zin[1][16] , \zin[1][15] ,
         \zin[1][14] , \zin[1][13] , \zin[1][12] , \zin[1][11] , \zin[1][10] ,
         \zin[1][9] , \zin[1][8] , \zin[1][7] , \zin[1][6] , \zin[1][5] ,
         \zin[1][4] , \zin[1][3] , \zin[1][2] , \zin[1][1] , \zin[1][0] ,
         \zin[0][257] , \zin[0][256] , \zin[0][255] , \zin[0][254] ,
         \zin[0][253] , \zin[0][252] , \zin[0][251] , \zin[0][250] ,
         \zin[0][249] , \zin[0][248] , \zin[0][247] , \zin[0][246] ,
         \zin[0][245] , \zin[0][244] , \zin[0][243] , \zin[0][242] ,
         \zin[0][241] , \zin[0][240] , \zin[0][239] , \zin[0][238] ,
         \zin[0][237] , \zin[0][236] , \zin[0][235] , \zin[0][234] ,
         \zin[0][233] , \zin[0][232] , \zin[0][231] , \zin[0][230] ,
         \zin[0][229] , \zin[0][228] , \zin[0][227] , \zin[0][226] ,
         \zin[0][225] , \zin[0][224] , \zin[0][223] , \zin[0][222] ,
         \zin[0][221] , \zin[0][220] , \zin[0][219] , \zin[0][218] ,
         \zin[0][217] , \zin[0][216] , \zin[0][215] , \zin[0][214] ,
         \zin[0][213] , \zin[0][212] , \zin[0][211] , \zin[0][210] ,
         \zin[0][209] , \zin[0][208] , \zin[0][207] , \zin[0][206] ,
         \zin[0][205] , \zin[0][204] , \zin[0][203] , \zin[0][202] ,
         \zin[0][201] , \zin[0][200] , \zin[0][199] , \zin[0][198] ,
         \zin[0][197] , \zin[0][196] , \zin[0][195] , \zin[0][194] ,
         \zin[0][193] , \zin[0][192] , \zin[0][191] , \zin[0][190] ,
         \zin[0][189] , \zin[0][188] , \zin[0][187] , \zin[0][186] ,
         \zin[0][185] , \zin[0][184] , \zin[0][183] , \zin[0][182] ,
         \zin[0][181] , \zin[0][180] , \zin[0][179] , \zin[0][178] ,
         \zin[0][177] , \zin[0][176] , \zin[0][175] , \zin[0][174] ,
         \zin[0][173] , \zin[0][172] , \zin[0][171] , \zin[0][170] ,
         \zin[0][169] , \zin[0][168] , \zin[0][167] , \zin[0][166] ,
         \zin[0][165] , \zin[0][164] , \zin[0][163] , \zin[0][162] ,
         \zin[0][161] , \zin[0][160] , \zin[0][159] , \zin[0][158] ,
         \zin[0][157] , \zin[0][156] , \zin[0][155] , \zin[0][154] ,
         \zin[0][153] , \zin[0][152] , \zin[0][151] , \zin[0][150] ,
         \zin[0][149] , \zin[0][148] , \zin[0][147] , \zin[0][146] ,
         \zin[0][145] , \zin[0][144] , \zin[0][143] , \zin[0][142] ,
         \zin[0][141] , \zin[0][140] , \zin[0][139] , \zin[0][138] ,
         \zin[0][137] , \zin[0][136] , \zin[0][135] , \zin[0][134] ,
         \zin[0][133] , \zin[0][132] , \zin[0][131] , \zin[0][130] ,
         \zin[0][129] , \zin[0][128] , \zin[0][127] , \zin[0][126] ,
         \zin[0][125] , \zin[0][124] , \zin[0][123] , \zin[0][122] ,
         \zin[0][121] , \zin[0][120] , \zin[0][119] , \zin[0][118] ,
         \zin[0][117] , \zin[0][116] , \zin[0][115] , \zin[0][114] ,
         \zin[0][113] , \zin[0][112] , \zin[0][111] , \zin[0][110] ,
         \zin[0][109] , \zin[0][108] , \zin[0][107] , \zin[0][106] ,
         \zin[0][105] , \zin[0][104] , \zin[0][103] , \zin[0][102] ,
         \zin[0][101] , \zin[0][100] , \zin[0][99] , \zin[0][98] ,
         \zin[0][97] , \zin[0][96] , \zin[0][95] , \zin[0][94] , \zin[0][93] ,
         \zin[0][92] , \zin[0][91] , \zin[0][90] , \zin[0][89] , \zin[0][88] ,
         \zin[0][87] , \zin[0][86] , \zin[0][85] , \zin[0][84] , \zin[0][83] ,
         \zin[0][82] , \zin[0][81] , \zin[0][80] , \zin[0][79] , \zin[0][78] ,
         \zin[0][77] , \zin[0][76] , \zin[0][75] , \zin[0][74] , \zin[0][73] ,
         \zin[0][72] , \zin[0][71] , \zin[0][70] , \zin[0][69] , \zin[0][68] ,
         \zin[0][67] , \zin[0][66] , \zin[0][65] , \zin[0][64] , \zin[0][63] ,
         \zin[0][62] , \zin[0][61] , \zin[0][60] , \zin[0][59] , \zin[0][58] ,
         \zin[0][57] , \zin[0][56] , \zin[0][55] , \zin[0][54] , \zin[0][53] ,
         \zin[0][52] , \zin[0][51] , \zin[0][50] , \zin[0][49] , \zin[0][48] ,
         \zin[0][47] , \zin[0][46] , \zin[0][45] , \zin[0][44] , \zin[0][43] ,
         \zin[0][42] , \zin[0][41] , \zin[0][40] , \zin[0][39] , \zin[0][38] ,
         \zin[0][37] , \zin[0][36] , \zin[0][35] , \zin[0][34] , \zin[0][33] ,
         \zin[0][32] , \zin[0][31] , \zin[0][30] , \zin[0][29] , \zin[0][28] ,
         \zin[0][27] , \zin[0][26] , \zin[0][25] , \zin[0][24] , \zin[0][23] ,
         \zin[0][22] , \zin[0][21] , \zin[0][20] , \zin[0][19] , \zin[0][18] ,
         \zin[0][17] , \zin[0][16] , \zin[0][15] , \zin[0][14] , \zin[0][13] ,
         \zin[0][12] , \zin[0][11] , \zin[0][10] , \zin[0][9] , \zin[0][8] ,
         \zin[0][7] , \zin[0][6] , \zin[0][5] , \zin[0][4] , \zin[0][3] ,
         \zin[0][2] , \zin[0][1] , \zin[0][0] , n1, n2, n3, n4, n5, n6, n7, n8,
         n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22,
         n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35, n36,
         n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50,
         n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204,
         n205, n206, n207, n208, n209, n210, n211, n212, n213, n214, n215,
         n216, n217, n218, n219, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n239, n240, n241, n242, n243, n244, n245, n246, n247, n248,
         n249, n250, n251, n252, n253, n254, n255, n256, n257, n258, n259,
         n260, n261, n262, n263, n264, n265, n266, n267, n268, n269, n270,
         n271, n272, n273, n274, n275, n276, n277, n278, n279, n280, n281,
         n282, n283, n284, n285, n286, n287, n288, n289, n290, n291, n292,
         n293, n294, n295, n296, n297, n298, n299, n300, n301, n302, n303,
         n304, n305, n306, n307, n308, n309, n310, n311, n312, n313, n314,
         n315, n316, n317, n318, n319, n320, n321, n322, n323, n324, n325,
         n326, n327, n328, n329, n330, n331, n332, n333, n334, n335, n336,
         n337, n338, n339, n340, n341, n342, n343, n344, n345, n346, n347,
         n348, n349, n350, n351, n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, n374, n375, n376, n377, n378, n379, n380,
         n381, n382, n383, n384, n385, n386, n387, n388, n389, n390, n391,
         n392, n393, n394, n395, n396, n397, n398, n399, n400, n401, n402,
         n403, n404, n405, n406, n407, n408, n409, n410, n411, n412, n413,
         n414, n415, n416, n417, n418, n419, n420, n421, n422, n423, n424,
         n425, n426, n427, n428, n429, n430, n431, n432, n433, n434, n435,
         n436, n437, n438, n439, n440, n441, n442, n443, n444, n445, n446,
         n447, n448, n449, n450, n451, n452, n453, n454, n455, n456, n457,
         n458, n459, n460, n461, n462, n463, n464, n465, n466, n467, n468,
         n469, n470, n471, n472, n473, n474, n475, n476, n477, n478, n479,
         n480, n481, n482, n483, n484, n485, n486, n487, n488, n489, n490,
         n491, n492, n493, n494, n495, n496, n497, n498, n499, n500, n501,
         n502, n503, n504, n505, n506, n507, n508;
  wire   [257:0] zreg;
  wire   [255:0] xin;
  wire   [255:0] xreg;

  DFF \xreg_reg[7]  ( .D(n505), .CLK(clk), .RST(rst), .Q(xreg[7]) );
  DFF \xreg_reg[11]  ( .D(xin[7]), .CLK(clk), .RST(rst), .Q(xreg[11]) );
  DFF \xreg_reg[15]  ( .D(xin[11]), .CLK(clk), .RST(rst), .Q(xreg[15]) );
  DFF \xreg_reg[19]  ( .D(xin[15]), .CLK(clk), .RST(rst), .Q(xreg[19]) );
  DFF \xreg_reg[23]  ( .D(xin[19]), .CLK(clk), .RST(rst), .Q(xreg[23]) );
  DFF \xreg_reg[27]  ( .D(xin[23]), .CLK(clk), .RST(rst), .Q(xreg[27]) );
  DFF \xreg_reg[31]  ( .D(xin[27]), .CLK(clk), .RST(rst), .Q(xreg[31]) );
  DFF \xreg_reg[35]  ( .D(xin[31]), .CLK(clk), .RST(rst), .Q(xreg[35]) );
  DFF \xreg_reg[39]  ( .D(xin[35]), .CLK(clk), .RST(rst), .Q(xreg[39]) );
  DFF \xreg_reg[43]  ( .D(xin[39]), .CLK(clk), .RST(rst), .Q(xreg[43]) );
  DFF \xreg_reg[47]  ( .D(xin[43]), .CLK(clk), .RST(rst), .Q(xreg[47]) );
  DFF \xreg_reg[51]  ( .D(xin[47]), .CLK(clk), .RST(rst), .Q(xreg[51]) );
  DFF \xreg_reg[55]  ( .D(xin[51]), .CLK(clk), .RST(rst), .Q(xreg[55]) );
  DFF \xreg_reg[59]  ( .D(xin[55]), .CLK(clk), .RST(rst), .Q(xreg[59]) );
  DFF \xreg_reg[63]  ( .D(xin[59]), .CLK(clk), .RST(rst), .Q(xreg[63]) );
  DFF \xreg_reg[67]  ( .D(xin[63]), .CLK(clk), .RST(rst), .Q(xreg[67]) );
  DFF \xreg_reg[71]  ( .D(xin[67]), .CLK(clk), .RST(rst), .Q(xreg[71]) );
  DFF \xreg_reg[75]  ( .D(xin[71]), .CLK(clk), .RST(rst), .Q(xreg[75]) );
  DFF \xreg_reg[79]  ( .D(xin[75]), .CLK(clk), .RST(rst), .Q(xreg[79]) );
  DFF \xreg_reg[83]  ( .D(xin[79]), .CLK(clk), .RST(rst), .Q(xreg[83]) );
  DFF \xreg_reg[87]  ( .D(xin[83]), .CLK(clk), .RST(rst), .Q(xreg[87]) );
  DFF \xreg_reg[91]  ( .D(xin[87]), .CLK(clk), .RST(rst), .Q(xreg[91]) );
  DFF \xreg_reg[95]  ( .D(xin[91]), .CLK(clk), .RST(rst), .Q(xreg[95]) );
  DFF \xreg_reg[99]  ( .D(xin[95]), .CLK(clk), .RST(rst), .Q(xreg[99]) );
  DFF \xreg_reg[103]  ( .D(xin[99]), .CLK(clk), .RST(rst), .Q(xreg[103]) );
  DFF \xreg_reg[107]  ( .D(xin[103]), .CLK(clk), .RST(rst), .Q(xreg[107]) );
  DFF \xreg_reg[111]  ( .D(xin[107]), .CLK(clk), .RST(rst), .Q(xreg[111]) );
  DFF \xreg_reg[115]  ( .D(xin[111]), .CLK(clk), .RST(rst), .Q(xreg[115]) );
  DFF \xreg_reg[119]  ( .D(xin[115]), .CLK(clk), .RST(rst), .Q(xreg[119]) );
  DFF \xreg_reg[123]  ( .D(xin[119]), .CLK(clk), .RST(rst), .Q(xreg[123]) );
  DFF \xreg_reg[127]  ( .D(xin[123]), .CLK(clk), .RST(rst), .Q(xreg[127]) );
  DFF \xreg_reg[131]  ( .D(xin[127]), .CLK(clk), .RST(rst), .Q(xreg[131]) );
  DFF \xreg_reg[135]  ( .D(xin[131]), .CLK(clk), .RST(rst), .Q(xreg[135]) );
  DFF \xreg_reg[139]  ( .D(xin[135]), .CLK(clk), .RST(rst), .Q(xreg[139]) );
  DFF \xreg_reg[143]  ( .D(xin[139]), .CLK(clk), .RST(rst), .Q(xreg[143]) );
  DFF \xreg_reg[147]  ( .D(xin[143]), .CLK(clk), .RST(rst), .Q(xreg[147]) );
  DFF \xreg_reg[151]  ( .D(xin[147]), .CLK(clk), .RST(rst), .Q(xreg[151]) );
  DFF \xreg_reg[155]  ( .D(xin[151]), .CLK(clk), .RST(rst), .Q(xreg[155]) );
  DFF \xreg_reg[159]  ( .D(xin[155]), .CLK(clk), .RST(rst), .Q(xreg[159]) );
  DFF \xreg_reg[163]  ( .D(xin[159]), .CLK(clk), .RST(rst), .Q(xreg[163]) );
  DFF \xreg_reg[167]  ( .D(xin[163]), .CLK(clk), .RST(rst), .Q(xreg[167]) );
  DFF \xreg_reg[171]  ( .D(xin[167]), .CLK(clk), .RST(rst), .Q(xreg[171]) );
  DFF \xreg_reg[175]  ( .D(xin[171]), .CLK(clk), .RST(rst), .Q(xreg[175]) );
  DFF \xreg_reg[179]  ( .D(xin[175]), .CLK(clk), .RST(rst), .Q(xreg[179]) );
  DFF \xreg_reg[183]  ( .D(xin[179]), .CLK(clk), .RST(rst), .Q(xreg[183]) );
  DFF \xreg_reg[187]  ( .D(xin[183]), .CLK(clk), .RST(rst), .Q(xreg[187]) );
  DFF \xreg_reg[191]  ( .D(xin[187]), .CLK(clk), .RST(rst), .Q(xreg[191]) );
  DFF \xreg_reg[195]  ( .D(xin[191]), .CLK(clk), .RST(rst), .Q(xreg[195]) );
  DFF \xreg_reg[199]  ( .D(xin[195]), .CLK(clk), .RST(rst), .Q(xreg[199]) );
  DFF \xreg_reg[203]  ( .D(xin[199]), .CLK(clk), .RST(rst), .Q(xreg[203]) );
  DFF \xreg_reg[207]  ( .D(xin[203]), .CLK(clk), .RST(rst), .Q(xreg[207]) );
  DFF \xreg_reg[211]  ( .D(xin[207]), .CLK(clk), .RST(rst), .Q(xreg[211]) );
  DFF \xreg_reg[215]  ( .D(xin[211]), .CLK(clk), .RST(rst), .Q(xreg[215]) );
  DFF \xreg_reg[219]  ( .D(xin[215]), .CLK(clk), .RST(rst), .Q(xreg[219]) );
  DFF \xreg_reg[223]  ( .D(xin[219]), .CLK(clk), .RST(rst), .Q(xreg[223]) );
  DFF \xreg_reg[227]  ( .D(xin[223]), .CLK(clk), .RST(rst), .Q(xreg[227]) );
  DFF \xreg_reg[231]  ( .D(xin[227]), .CLK(clk), .RST(rst), .Q(xreg[231]) );
  DFF \xreg_reg[235]  ( .D(xin[231]), .CLK(clk), .RST(rst), .Q(xreg[235]) );
  DFF \xreg_reg[239]  ( .D(xin[235]), .CLK(clk), .RST(rst), .Q(xreg[239]) );
  DFF \xreg_reg[243]  ( .D(xin[239]), .CLK(clk), .RST(rst), .Q(xreg[243]) );
  DFF \xreg_reg[247]  ( .D(xin[243]), .CLK(clk), .RST(rst), .Q(xreg[247]) );
  DFF \xreg_reg[251]  ( .D(xin[247]), .CLK(clk), .RST(rst), .Q(xreg[251]) );
  DFF \xreg_reg[255]  ( .D(xin[251]), .CLK(clk), .RST(rst), .Q(xreg[255]) );
  DFF \xreg_reg[6]  ( .D(n506), .CLK(clk), .RST(rst), .Q(xreg[6]) );
  DFF \xreg_reg[10]  ( .D(xin[6]), .CLK(clk), .RST(rst), .Q(xreg[10]) );
  DFF \xreg_reg[14]  ( .D(xin[10]), .CLK(clk), .RST(rst), .Q(xreg[14]) );
  DFF \xreg_reg[18]  ( .D(xin[14]), .CLK(clk), .RST(rst), .Q(xreg[18]) );
  DFF \xreg_reg[22]  ( .D(xin[18]), .CLK(clk), .RST(rst), .Q(xreg[22]) );
  DFF \xreg_reg[26]  ( .D(xin[22]), .CLK(clk), .RST(rst), .Q(xreg[26]) );
  DFF \xreg_reg[30]  ( .D(xin[26]), .CLK(clk), .RST(rst), .Q(xreg[30]) );
  DFF \xreg_reg[34]  ( .D(xin[30]), .CLK(clk), .RST(rst), .Q(xreg[34]) );
  DFF \xreg_reg[38]  ( .D(xin[34]), .CLK(clk), .RST(rst), .Q(xreg[38]) );
  DFF \xreg_reg[42]  ( .D(xin[38]), .CLK(clk), .RST(rst), .Q(xreg[42]) );
  DFF \xreg_reg[46]  ( .D(xin[42]), .CLK(clk), .RST(rst), .Q(xreg[46]) );
  DFF \xreg_reg[50]  ( .D(xin[46]), .CLK(clk), .RST(rst), .Q(xreg[50]) );
  DFF \xreg_reg[54]  ( .D(xin[50]), .CLK(clk), .RST(rst), .Q(xreg[54]) );
  DFF \xreg_reg[58]  ( .D(xin[54]), .CLK(clk), .RST(rst), .Q(xreg[58]) );
  DFF \xreg_reg[62]  ( .D(xin[58]), .CLK(clk), .RST(rst), .Q(xreg[62]) );
  DFF \xreg_reg[66]  ( .D(xin[62]), .CLK(clk), .RST(rst), .Q(xreg[66]) );
  DFF \xreg_reg[70]  ( .D(xin[66]), .CLK(clk), .RST(rst), .Q(xreg[70]) );
  DFF \xreg_reg[74]  ( .D(xin[70]), .CLK(clk), .RST(rst), .Q(xreg[74]) );
  DFF \xreg_reg[78]  ( .D(xin[74]), .CLK(clk), .RST(rst), .Q(xreg[78]) );
  DFF \xreg_reg[82]  ( .D(xin[78]), .CLK(clk), .RST(rst), .Q(xreg[82]) );
  DFF \xreg_reg[86]  ( .D(xin[82]), .CLK(clk), .RST(rst), .Q(xreg[86]) );
  DFF \xreg_reg[90]  ( .D(xin[86]), .CLK(clk), .RST(rst), .Q(xreg[90]) );
  DFF \xreg_reg[94]  ( .D(xin[90]), .CLK(clk), .RST(rst), .Q(xreg[94]) );
  DFF \xreg_reg[98]  ( .D(xin[94]), .CLK(clk), .RST(rst), .Q(xreg[98]) );
  DFF \xreg_reg[102]  ( .D(xin[98]), .CLK(clk), .RST(rst), .Q(xreg[102]) );
  DFF \xreg_reg[106]  ( .D(xin[102]), .CLK(clk), .RST(rst), .Q(xreg[106]) );
  DFF \xreg_reg[110]  ( .D(xin[106]), .CLK(clk), .RST(rst), .Q(xreg[110]) );
  DFF \xreg_reg[114]  ( .D(xin[110]), .CLK(clk), .RST(rst), .Q(xreg[114]) );
  DFF \xreg_reg[118]  ( .D(xin[114]), .CLK(clk), .RST(rst), .Q(xreg[118]) );
  DFF \xreg_reg[122]  ( .D(xin[118]), .CLK(clk), .RST(rst), .Q(xreg[122]) );
  DFF \xreg_reg[126]  ( .D(xin[122]), .CLK(clk), .RST(rst), .Q(xreg[126]) );
  DFF \xreg_reg[130]  ( .D(xin[126]), .CLK(clk), .RST(rst), .Q(xreg[130]) );
  DFF \xreg_reg[134]  ( .D(xin[130]), .CLK(clk), .RST(rst), .Q(xreg[134]) );
  DFF \xreg_reg[138]  ( .D(xin[134]), .CLK(clk), .RST(rst), .Q(xreg[138]) );
  DFF \xreg_reg[142]  ( .D(xin[138]), .CLK(clk), .RST(rst), .Q(xreg[142]) );
  DFF \xreg_reg[146]  ( .D(xin[142]), .CLK(clk), .RST(rst), .Q(xreg[146]) );
  DFF \xreg_reg[150]  ( .D(xin[146]), .CLK(clk), .RST(rst), .Q(xreg[150]) );
  DFF \xreg_reg[154]  ( .D(xin[150]), .CLK(clk), .RST(rst), .Q(xreg[154]) );
  DFF \xreg_reg[158]  ( .D(xin[154]), .CLK(clk), .RST(rst), .Q(xreg[158]) );
  DFF \xreg_reg[162]  ( .D(xin[158]), .CLK(clk), .RST(rst), .Q(xreg[162]) );
  DFF \xreg_reg[166]  ( .D(xin[162]), .CLK(clk), .RST(rst), .Q(xreg[166]) );
  DFF \xreg_reg[170]  ( .D(xin[166]), .CLK(clk), .RST(rst), .Q(xreg[170]) );
  DFF \xreg_reg[174]  ( .D(xin[170]), .CLK(clk), .RST(rst), .Q(xreg[174]) );
  DFF \xreg_reg[178]  ( .D(xin[174]), .CLK(clk), .RST(rst), .Q(xreg[178]) );
  DFF \xreg_reg[182]  ( .D(xin[178]), .CLK(clk), .RST(rst), .Q(xreg[182]) );
  DFF \xreg_reg[186]  ( .D(xin[182]), .CLK(clk), .RST(rst), .Q(xreg[186]) );
  DFF \xreg_reg[190]  ( .D(xin[186]), .CLK(clk), .RST(rst), .Q(xreg[190]) );
  DFF \xreg_reg[194]  ( .D(xin[190]), .CLK(clk), .RST(rst), .Q(xreg[194]) );
  DFF \xreg_reg[198]  ( .D(xin[194]), .CLK(clk), .RST(rst), .Q(xreg[198]) );
  DFF \xreg_reg[202]  ( .D(xin[198]), .CLK(clk), .RST(rst), .Q(xreg[202]) );
  DFF \xreg_reg[206]  ( .D(xin[202]), .CLK(clk), .RST(rst), .Q(xreg[206]) );
  DFF \xreg_reg[210]  ( .D(xin[206]), .CLK(clk), .RST(rst), .Q(xreg[210]) );
  DFF \xreg_reg[214]  ( .D(xin[210]), .CLK(clk), .RST(rst), .Q(xreg[214]) );
  DFF \xreg_reg[218]  ( .D(xin[214]), .CLK(clk), .RST(rst), .Q(xreg[218]) );
  DFF \xreg_reg[222]  ( .D(xin[218]), .CLK(clk), .RST(rst), .Q(xreg[222]) );
  DFF \xreg_reg[226]  ( .D(xin[222]), .CLK(clk), .RST(rst), .Q(xreg[226]) );
  DFF \xreg_reg[230]  ( .D(xin[226]), .CLK(clk), .RST(rst), .Q(xreg[230]) );
  DFF \xreg_reg[234]  ( .D(xin[230]), .CLK(clk), .RST(rst), .Q(xreg[234]) );
  DFF \xreg_reg[238]  ( .D(xin[234]), .CLK(clk), .RST(rst), .Q(xreg[238]) );
  DFF \xreg_reg[242]  ( .D(xin[238]), .CLK(clk), .RST(rst), .Q(xreg[242]) );
  DFF \xreg_reg[246]  ( .D(xin[242]), .CLK(clk), .RST(rst), .Q(xreg[246]) );
  DFF \xreg_reg[250]  ( .D(xin[246]), .CLK(clk), .RST(rst), .Q(xreg[250]) );
  DFF \xreg_reg[254]  ( .D(xin[250]), .CLK(clk), .RST(rst), .Q(xreg[254]) );
  DFF \xreg_reg[5]  ( .D(n507), .CLK(clk), .RST(rst), .Q(xreg[5]) );
  DFF \xreg_reg[9]  ( .D(xin[5]), .CLK(clk), .RST(rst), .Q(xreg[9]) );
  DFF \xreg_reg[13]  ( .D(xin[9]), .CLK(clk), .RST(rst), .Q(xreg[13]) );
  DFF \xreg_reg[17]  ( .D(xin[13]), .CLK(clk), .RST(rst), .Q(xreg[17]) );
  DFF \xreg_reg[21]  ( .D(xin[17]), .CLK(clk), .RST(rst), .Q(xreg[21]) );
  DFF \xreg_reg[25]  ( .D(xin[21]), .CLK(clk), .RST(rst), .Q(xreg[25]) );
  DFF \xreg_reg[29]  ( .D(xin[25]), .CLK(clk), .RST(rst), .Q(xreg[29]) );
  DFF \xreg_reg[33]  ( .D(xin[29]), .CLK(clk), .RST(rst), .Q(xreg[33]) );
  DFF \xreg_reg[37]  ( .D(xin[33]), .CLK(clk), .RST(rst), .Q(xreg[37]) );
  DFF \xreg_reg[41]  ( .D(xin[37]), .CLK(clk), .RST(rst), .Q(xreg[41]) );
  DFF \xreg_reg[45]  ( .D(xin[41]), .CLK(clk), .RST(rst), .Q(xreg[45]) );
  DFF \xreg_reg[49]  ( .D(xin[45]), .CLK(clk), .RST(rst), .Q(xreg[49]) );
  DFF \xreg_reg[53]  ( .D(xin[49]), .CLK(clk), .RST(rst), .Q(xreg[53]) );
  DFF \xreg_reg[57]  ( .D(xin[53]), .CLK(clk), .RST(rst), .Q(xreg[57]) );
  DFF \xreg_reg[61]  ( .D(xin[57]), .CLK(clk), .RST(rst), .Q(xreg[61]) );
  DFF \xreg_reg[65]  ( .D(xin[61]), .CLK(clk), .RST(rst), .Q(xreg[65]) );
  DFF \xreg_reg[69]  ( .D(xin[65]), .CLK(clk), .RST(rst), .Q(xreg[69]) );
  DFF \xreg_reg[73]  ( .D(xin[69]), .CLK(clk), .RST(rst), .Q(xreg[73]) );
  DFF \xreg_reg[77]  ( .D(xin[73]), .CLK(clk), .RST(rst), .Q(xreg[77]) );
  DFF \xreg_reg[81]  ( .D(xin[77]), .CLK(clk), .RST(rst), .Q(xreg[81]) );
  DFF \xreg_reg[85]  ( .D(xin[81]), .CLK(clk), .RST(rst), .Q(xreg[85]) );
  DFF \xreg_reg[89]  ( .D(xin[85]), .CLK(clk), .RST(rst), .Q(xreg[89]) );
  DFF \xreg_reg[93]  ( .D(xin[89]), .CLK(clk), .RST(rst), .Q(xreg[93]) );
  DFF \xreg_reg[97]  ( .D(xin[93]), .CLK(clk), .RST(rst), .Q(xreg[97]) );
  DFF \xreg_reg[101]  ( .D(xin[97]), .CLK(clk), .RST(rst), .Q(xreg[101]) );
  DFF \xreg_reg[105]  ( .D(xin[101]), .CLK(clk), .RST(rst), .Q(xreg[105]) );
  DFF \xreg_reg[109]  ( .D(xin[105]), .CLK(clk), .RST(rst), .Q(xreg[109]) );
  DFF \xreg_reg[113]  ( .D(xin[109]), .CLK(clk), .RST(rst), .Q(xreg[113]) );
  DFF \xreg_reg[117]  ( .D(xin[113]), .CLK(clk), .RST(rst), .Q(xreg[117]) );
  DFF \xreg_reg[121]  ( .D(xin[117]), .CLK(clk), .RST(rst), .Q(xreg[121]) );
  DFF \xreg_reg[125]  ( .D(xin[121]), .CLK(clk), .RST(rst), .Q(xreg[125]) );
  DFF \xreg_reg[129]  ( .D(xin[125]), .CLK(clk), .RST(rst), .Q(xreg[129]) );
  DFF \xreg_reg[133]  ( .D(xin[129]), .CLK(clk), .RST(rst), .Q(xreg[133]) );
  DFF \xreg_reg[137]  ( .D(xin[133]), .CLK(clk), .RST(rst), .Q(xreg[137]) );
  DFF \xreg_reg[141]  ( .D(xin[137]), .CLK(clk), .RST(rst), .Q(xreg[141]) );
  DFF \xreg_reg[145]  ( .D(xin[141]), .CLK(clk), .RST(rst), .Q(xreg[145]) );
  DFF \xreg_reg[149]  ( .D(xin[145]), .CLK(clk), .RST(rst), .Q(xreg[149]) );
  DFF \xreg_reg[153]  ( .D(xin[149]), .CLK(clk), .RST(rst), .Q(xreg[153]) );
  DFF \xreg_reg[157]  ( .D(xin[153]), .CLK(clk), .RST(rst), .Q(xreg[157]) );
  DFF \xreg_reg[161]  ( .D(xin[157]), .CLK(clk), .RST(rst), .Q(xreg[161]) );
  DFF \xreg_reg[165]  ( .D(xin[161]), .CLK(clk), .RST(rst), .Q(xreg[165]) );
  DFF \xreg_reg[169]  ( .D(xin[165]), .CLK(clk), .RST(rst), .Q(xreg[169]) );
  DFF \xreg_reg[173]  ( .D(xin[169]), .CLK(clk), .RST(rst), .Q(xreg[173]) );
  DFF \xreg_reg[177]  ( .D(xin[173]), .CLK(clk), .RST(rst), .Q(xreg[177]) );
  DFF \xreg_reg[181]  ( .D(xin[177]), .CLK(clk), .RST(rst), .Q(xreg[181]) );
  DFF \xreg_reg[185]  ( .D(xin[181]), .CLK(clk), .RST(rst), .Q(xreg[185]) );
  DFF \xreg_reg[189]  ( .D(xin[185]), .CLK(clk), .RST(rst), .Q(xreg[189]) );
  DFF \xreg_reg[193]  ( .D(xin[189]), .CLK(clk), .RST(rst), .Q(xreg[193]) );
  DFF \xreg_reg[197]  ( .D(xin[193]), .CLK(clk), .RST(rst), .Q(xreg[197]) );
  DFF \xreg_reg[201]  ( .D(xin[197]), .CLK(clk), .RST(rst), .Q(xreg[201]) );
  DFF \xreg_reg[205]  ( .D(xin[201]), .CLK(clk), .RST(rst), .Q(xreg[205]) );
  DFF \xreg_reg[209]  ( .D(xin[205]), .CLK(clk), .RST(rst), .Q(xreg[209]) );
  DFF \xreg_reg[213]  ( .D(xin[209]), .CLK(clk), .RST(rst), .Q(xreg[213]) );
  DFF \xreg_reg[217]  ( .D(xin[213]), .CLK(clk), .RST(rst), .Q(xreg[217]) );
  DFF \xreg_reg[221]  ( .D(xin[217]), .CLK(clk), .RST(rst), .Q(xreg[221]) );
  DFF \xreg_reg[225]  ( .D(xin[221]), .CLK(clk), .RST(rst), .Q(xreg[225]) );
  DFF \xreg_reg[229]  ( .D(xin[225]), .CLK(clk), .RST(rst), .Q(xreg[229]) );
  DFF \xreg_reg[233]  ( .D(xin[229]), .CLK(clk), .RST(rst), .Q(xreg[233]) );
  DFF \xreg_reg[237]  ( .D(xin[233]), .CLK(clk), .RST(rst), .Q(xreg[237]) );
  DFF \xreg_reg[241]  ( .D(xin[237]), .CLK(clk), .RST(rst), .Q(xreg[241]) );
  DFF \xreg_reg[245]  ( .D(xin[241]), .CLK(clk), .RST(rst), .Q(xreg[245]) );
  DFF \xreg_reg[249]  ( .D(xin[245]), .CLK(clk), .RST(rst), .Q(xreg[249]) );
  DFF \xreg_reg[253]  ( .D(xin[249]), .CLK(clk), .RST(rst), .Q(xreg[253]) );
  DFF \xreg_reg[4]  ( .D(n508), .CLK(clk), .RST(rst), .Q(xreg[4]) );
  DFF \xreg_reg[8]  ( .D(xin[4]), .CLK(clk), .RST(rst), .Q(xreg[8]) );
  DFF \xreg_reg[12]  ( .D(xin[8]), .CLK(clk), .RST(rst), .Q(xreg[12]) );
  DFF \xreg_reg[16]  ( .D(xin[12]), .CLK(clk), .RST(rst), .Q(xreg[16]) );
  DFF \xreg_reg[20]  ( .D(xin[16]), .CLK(clk), .RST(rst), .Q(xreg[20]) );
  DFF \xreg_reg[24]  ( .D(xin[20]), .CLK(clk), .RST(rst), .Q(xreg[24]) );
  DFF \xreg_reg[28]  ( .D(xin[24]), .CLK(clk), .RST(rst), .Q(xreg[28]) );
  DFF \xreg_reg[32]  ( .D(xin[28]), .CLK(clk), .RST(rst), .Q(xreg[32]) );
  DFF \xreg_reg[36]  ( .D(xin[32]), .CLK(clk), .RST(rst), .Q(xreg[36]) );
  DFF \xreg_reg[40]  ( .D(xin[36]), .CLK(clk), .RST(rst), .Q(xreg[40]) );
  DFF \xreg_reg[44]  ( .D(xin[40]), .CLK(clk), .RST(rst), .Q(xreg[44]) );
  DFF \xreg_reg[48]  ( .D(xin[44]), .CLK(clk), .RST(rst), .Q(xreg[48]) );
  DFF \xreg_reg[52]  ( .D(xin[48]), .CLK(clk), .RST(rst), .Q(xreg[52]) );
  DFF \xreg_reg[56]  ( .D(xin[52]), .CLK(clk), .RST(rst), .Q(xreg[56]) );
  DFF \xreg_reg[60]  ( .D(xin[56]), .CLK(clk), .RST(rst), .Q(xreg[60]) );
  DFF \xreg_reg[64]  ( .D(xin[60]), .CLK(clk), .RST(rst), .Q(xreg[64]) );
  DFF \xreg_reg[68]  ( .D(xin[64]), .CLK(clk), .RST(rst), .Q(xreg[68]) );
  DFF \xreg_reg[72]  ( .D(xin[68]), .CLK(clk), .RST(rst), .Q(xreg[72]) );
  DFF \xreg_reg[76]  ( .D(xin[72]), .CLK(clk), .RST(rst), .Q(xreg[76]) );
  DFF \xreg_reg[80]  ( .D(xin[76]), .CLK(clk), .RST(rst), .Q(xreg[80]) );
  DFF \xreg_reg[84]  ( .D(xin[80]), .CLK(clk), .RST(rst), .Q(xreg[84]) );
  DFF \xreg_reg[88]  ( .D(xin[84]), .CLK(clk), .RST(rst), .Q(xreg[88]) );
  DFF \xreg_reg[92]  ( .D(xin[88]), .CLK(clk), .RST(rst), .Q(xreg[92]) );
  DFF \xreg_reg[96]  ( .D(xin[92]), .CLK(clk), .RST(rst), .Q(xreg[96]) );
  DFF \xreg_reg[100]  ( .D(xin[96]), .CLK(clk), .RST(rst), .Q(xreg[100]) );
  DFF \xreg_reg[104]  ( .D(xin[100]), .CLK(clk), .RST(rst), .Q(xreg[104]) );
  DFF \xreg_reg[108]  ( .D(xin[104]), .CLK(clk), .RST(rst), .Q(xreg[108]) );
  DFF \xreg_reg[112]  ( .D(xin[108]), .CLK(clk), .RST(rst), .Q(xreg[112]) );
  DFF \xreg_reg[116]  ( .D(xin[112]), .CLK(clk), .RST(rst), .Q(xreg[116]) );
  DFF \xreg_reg[120]  ( .D(xin[116]), .CLK(clk), .RST(rst), .Q(xreg[120]) );
  DFF \xreg_reg[124]  ( .D(xin[120]), .CLK(clk), .RST(rst), .Q(xreg[124]) );
  DFF \xreg_reg[128]  ( .D(xin[124]), .CLK(clk), .RST(rst), .Q(xreg[128]) );
  DFF \xreg_reg[132]  ( .D(xin[128]), .CLK(clk), .RST(rst), .Q(xreg[132]) );
  DFF \xreg_reg[136]  ( .D(xin[132]), .CLK(clk), .RST(rst), .Q(xreg[136]) );
  DFF \xreg_reg[140]  ( .D(xin[136]), .CLK(clk), .RST(rst), .Q(xreg[140]) );
  DFF \xreg_reg[144]  ( .D(xin[140]), .CLK(clk), .RST(rst), .Q(xreg[144]) );
  DFF \xreg_reg[148]  ( .D(xin[144]), .CLK(clk), .RST(rst), .Q(xreg[148]) );
  DFF \xreg_reg[152]  ( .D(xin[148]), .CLK(clk), .RST(rst), .Q(xreg[152]) );
  DFF \xreg_reg[156]  ( .D(xin[152]), .CLK(clk), .RST(rst), .Q(xreg[156]) );
  DFF \xreg_reg[160]  ( .D(xin[156]), .CLK(clk), .RST(rst), .Q(xreg[160]) );
  DFF \xreg_reg[164]  ( .D(xin[160]), .CLK(clk), .RST(rst), .Q(xreg[164]) );
  DFF \xreg_reg[168]  ( .D(xin[164]), .CLK(clk), .RST(rst), .Q(xreg[168]) );
  DFF \xreg_reg[172]  ( .D(xin[168]), .CLK(clk), .RST(rst), .Q(xreg[172]) );
  DFF \xreg_reg[176]  ( .D(xin[172]), .CLK(clk), .RST(rst), .Q(xreg[176]) );
  DFF \xreg_reg[180]  ( .D(xin[176]), .CLK(clk), .RST(rst), .Q(xreg[180]) );
  DFF \xreg_reg[184]  ( .D(xin[180]), .CLK(clk), .RST(rst), .Q(xreg[184]) );
  DFF \xreg_reg[188]  ( .D(xin[184]), .CLK(clk), .RST(rst), .Q(xreg[188]) );
  DFF \xreg_reg[192]  ( .D(xin[188]), .CLK(clk), .RST(rst), .Q(xreg[192]) );
  DFF \xreg_reg[196]  ( .D(xin[192]), .CLK(clk), .RST(rst), .Q(xreg[196]) );
  DFF \xreg_reg[200]  ( .D(xin[196]), .CLK(clk), .RST(rst), .Q(xreg[200]) );
  DFF \xreg_reg[204]  ( .D(xin[200]), .CLK(clk), .RST(rst), .Q(xreg[204]) );
  DFF \xreg_reg[208]  ( .D(xin[204]), .CLK(clk), .RST(rst), .Q(xreg[208]) );
  DFF \xreg_reg[212]  ( .D(xin[208]), .CLK(clk), .RST(rst), .Q(xreg[212]) );
  DFF \xreg_reg[216]  ( .D(xin[212]), .CLK(clk), .RST(rst), .Q(xreg[216]) );
  DFF \xreg_reg[220]  ( .D(xin[216]), .CLK(clk), .RST(rst), .Q(xreg[220]) );
  DFF \xreg_reg[224]  ( .D(xin[220]), .CLK(clk), .RST(rst), .Q(xreg[224]) );
  DFF \xreg_reg[228]  ( .D(xin[224]), .CLK(clk), .RST(rst), .Q(xreg[228]) );
  DFF \xreg_reg[232]  ( .D(xin[228]), .CLK(clk), .RST(rst), .Q(xreg[232]) );
  DFF \xreg_reg[236]  ( .D(xin[232]), .CLK(clk), .RST(rst), .Q(xreg[236]) );
  DFF \xreg_reg[240]  ( .D(xin[236]), .CLK(clk), .RST(rst), .Q(xreg[240]) );
  DFF \xreg_reg[244]  ( .D(xin[240]), .CLK(clk), .RST(rst), .Q(xreg[244]) );
  DFF \xreg_reg[248]  ( .D(xin[244]), .CLK(clk), .RST(rst), .Q(xreg[248]) );
  DFF \xreg_reg[252]  ( .D(xin[248]), .CLK(clk), .RST(rst), .Q(xreg[252]) );
  DFF \zreg_reg[0]  ( .D(o[0]), .CLK(clk), .RST(rst), .Q(zreg[0]) );
  DFF \zreg_reg[1]  ( .D(o[1]), .CLK(clk), .RST(rst), .Q(zreg[1]) );
  DFF \zreg_reg[2]  ( .D(o[2]), .CLK(clk), .RST(rst), .Q(zreg[2]) );
  DFF \zreg_reg[3]  ( .D(o[3]), .CLK(clk), .RST(rst), .Q(zreg[3]) );
  DFF \zreg_reg[4]  ( .D(o[4]), .CLK(clk), .RST(rst), .Q(zreg[4]) );
  DFF \zreg_reg[5]  ( .D(o[5]), .CLK(clk), .RST(rst), .Q(zreg[5]) );
  DFF \zreg_reg[6]  ( .D(o[6]), .CLK(clk), .RST(rst), .Q(zreg[6]) );
  DFF \zreg_reg[7]  ( .D(o[7]), .CLK(clk), .RST(rst), .Q(zreg[7]) );
  DFF \zreg_reg[8]  ( .D(o[8]), .CLK(clk), .RST(rst), .Q(zreg[8]) );
  DFF \zreg_reg[9]  ( .D(o[9]), .CLK(clk), .RST(rst), .Q(zreg[9]) );
  DFF \zreg_reg[10]  ( .D(o[10]), .CLK(clk), .RST(rst), .Q(zreg[10]) );
  DFF \zreg_reg[11]  ( .D(o[11]), .CLK(clk), .RST(rst), .Q(zreg[11]) );
  DFF \zreg_reg[12]  ( .D(o[12]), .CLK(clk), .RST(rst), .Q(zreg[12]) );
  DFF \zreg_reg[13]  ( .D(o[13]), .CLK(clk), .RST(rst), .Q(zreg[13]) );
  DFF \zreg_reg[14]  ( .D(o[14]), .CLK(clk), .RST(rst), .Q(zreg[14]) );
  DFF \zreg_reg[15]  ( .D(o[15]), .CLK(clk), .RST(rst), .Q(zreg[15]) );
  DFF \zreg_reg[16]  ( .D(o[16]), .CLK(clk), .RST(rst), .Q(zreg[16]) );
  DFF \zreg_reg[17]  ( .D(o[17]), .CLK(clk), .RST(rst), .Q(zreg[17]) );
  DFF \zreg_reg[18]  ( .D(o[18]), .CLK(clk), .RST(rst), .Q(zreg[18]) );
  DFF \zreg_reg[19]  ( .D(o[19]), .CLK(clk), .RST(rst), .Q(zreg[19]) );
  DFF \zreg_reg[20]  ( .D(o[20]), .CLK(clk), .RST(rst), .Q(zreg[20]) );
  DFF \zreg_reg[21]  ( .D(o[21]), .CLK(clk), .RST(rst), .Q(zreg[21]) );
  DFF \zreg_reg[22]  ( .D(o[22]), .CLK(clk), .RST(rst), .Q(zreg[22]) );
  DFF \zreg_reg[23]  ( .D(o[23]), .CLK(clk), .RST(rst), .Q(zreg[23]) );
  DFF \zreg_reg[24]  ( .D(o[24]), .CLK(clk), .RST(rst), .Q(zreg[24]) );
  DFF \zreg_reg[25]  ( .D(o[25]), .CLK(clk), .RST(rst), .Q(zreg[25]) );
  DFF \zreg_reg[26]  ( .D(o[26]), .CLK(clk), .RST(rst), .Q(zreg[26]) );
  DFF \zreg_reg[27]  ( .D(o[27]), .CLK(clk), .RST(rst), .Q(zreg[27]) );
  DFF \zreg_reg[28]  ( .D(o[28]), .CLK(clk), .RST(rst), .Q(zreg[28]) );
  DFF \zreg_reg[29]  ( .D(o[29]), .CLK(clk), .RST(rst), .Q(zreg[29]) );
  DFF \zreg_reg[30]  ( .D(o[30]), .CLK(clk), .RST(rst), .Q(zreg[30]) );
  DFF \zreg_reg[31]  ( .D(o[31]), .CLK(clk), .RST(rst), .Q(zreg[31]) );
  DFF \zreg_reg[32]  ( .D(o[32]), .CLK(clk), .RST(rst), .Q(zreg[32]) );
  DFF \zreg_reg[33]  ( .D(o[33]), .CLK(clk), .RST(rst), .Q(zreg[33]) );
  DFF \zreg_reg[34]  ( .D(o[34]), .CLK(clk), .RST(rst), .Q(zreg[34]) );
  DFF \zreg_reg[35]  ( .D(o[35]), .CLK(clk), .RST(rst), .Q(zreg[35]) );
  DFF \zreg_reg[36]  ( .D(o[36]), .CLK(clk), .RST(rst), .Q(zreg[36]) );
  DFF \zreg_reg[37]  ( .D(o[37]), .CLK(clk), .RST(rst), .Q(zreg[37]) );
  DFF \zreg_reg[38]  ( .D(o[38]), .CLK(clk), .RST(rst), .Q(zreg[38]) );
  DFF \zreg_reg[39]  ( .D(o[39]), .CLK(clk), .RST(rst), .Q(zreg[39]) );
  DFF \zreg_reg[40]  ( .D(o[40]), .CLK(clk), .RST(rst), .Q(zreg[40]) );
  DFF \zreg_reg[41]  ( .D(o[41]), .CLK(clk), .RST(rst), .Q(zreg[41]) );
  DFF \zreg_reg[42]  ( .D(o[42]), .CLK(clk), .RST(rst), .Q(zreg[42]) );
  DFF \zreg_reg[43]  ( .D(o[43]), .CLK(clk), .RST(rst), .Q(zreg[43]) );
  DFF \zreg_reg[44]  ( .D(o[44]), .CLK(clk), .RST(rst), .Q(zreg[44]) );
  DFF \zreg_reg[45]  ( .D(o[45]), .CLK(clk), .RST(rst), .Q(zreg[45]) );
  DFF \zreg_reg[46]  ( .D(o[46]), .CLK(clk), .RST(rst), .Q(zreg[46]) );
  DFF \zreg_reg[47]  ( .D(o[47]), .CLK(clk), .RST(rst), .Q(zreg[47]) );
  DFF \zreg_reg[48]  ( .D(o[48]), .CLK(clk), .RST(rst), .Q(zreg[48]) );
  DFF \zreg_reg[49]  ( .D(o[49]), .CLK(clk), .RST(rst), .Q(zreg[49]) );
  DFF \zreg_reg[50]  ( .D(o[50]), .CLK(clk), .RST(rst), .Q(zreg[50]) );
  DFF \zreg_reg[51]  ( .D(o[51]), .CLK(clk), .RST(rst), .Q(zreg[51]) );
  DFF \zreg_reg[52]  ( .D(o[52]), .CLK(clk), .RST(rst), .Q(zreg[52]) );
  DFF \zreg_reg[53]  ( .D(o[53]), .CLK(clk), .RST(rst), .Q(zreg[53]) );
  DFF \zreg_reg[54]  ( .D(o[54]), .CLK(clk), .RST(rst), .Q(zreg[54]) );
  DFF \zreg_reg[55]  ( .D(o[55]), .CLK(clk), .RST(rst), .Q(zreg[55]) );
  DFF \zreg_reg[56]  ( .D(o[56]), .CLK(clk), .RST(rst), .Q(zreg[56]) );
  DFF \zreg_reg[57]  ( .D(o[57]), .CLK(clk), .RST(rst), .Q(zreg[57]) );
  DFF \zreg_reg[58]  ( .D(o[58]), .CLK(clk), .RST(rst), .Q(zreg[58]) );
  DFF \zreg_reg[59]  ( .D(o[59]), .CLK(clk), .RST(rst), .Q(zreg[59]) );
  DFF \zreg_reg[60]  ( .D(o[60]), .CLK(clk), .RST(rst), .Q(zreg[60]) );
  DFF \zreg_reg[61]  ( .D(o[61]), .CLK(clk), .RST(rst), .Q(zreg[61]) );
  DFF \zreg_reg[62]  ( .D(o[62]), .CLK(clk), .RST(rst), .Q(zreg[62]) );
  DFF \zreg_reg[63]  ( .D(o[63]), .CLK(clk), .RST(rst), .Q(zreg[63]) );
  DFF \zreg_reg[64]  ( .D(o[64]), .CLK(clk), .RST(rst), .Q(zreg[64]) );
  DFF \zreg_reg[65]  ( .D(o[65]), .CLK(clk), .RST(rst), .Q(zreg[65]) );
  DFF \zreg_reg[66]  ( .D(o[66]), .CLK(clk), .RST(rst), .Q(zreg[66]) );
  DFF \zreg_reg[67]  ( .D(o[67]), .CLK(clk), .RST(rst), .Q(zreg[67]) );
  DFF \zreg_reg[68]  ( .D(o[68]), .CLK(clk), .RST(rst), .Q(zreg[68]) );
  DFF \zreg_reg[69]  ( .D(o[69]), .CLK(clk), .RST(rst), .Q(zreg[69]) );
  DFF \zreg_reg[70]  ( .D(o[70]), .CLK(clk), .RST(rst), .Q(zreg[70]) );
  DFF \zreg_reg[71]  ( .D(o[71]), .CLK(clk), .RST(rst), .Q(zreg[71]) );
  DFF \zreg_reg[72]  ( .D(o[72]), .CLK(clk), .RST(rst), .Q(zreg[72]) );
  DFF \zreg_reg[73]  ( .D(o[73]), .CLK(clk), .RST(rst), .Q(zreg[73]) );
  DFF \zreg_reg[74]  ( .D(o[74]), .CLK(clk), .RST(rst), .Q(zreg[74]) );
  DFF \zreg_reg[75]  ( .D(o[75]), .CLK(clk), .RST(rst), .Q(zreg[75]) );
  DFF \zreg_reg[76]  ( .D(o[76]), .CLK(clk), .RST(rst), .Q(zreg[76]) );
  DFF \zreg_reg[77]  ( .D(o[77]), .CLK(clk), .RST(rst), .Q(zreg[77]) );
  DFF \zreg_reg[78]  ( .D(o[78]), .CLK(clk), .RST(rst), .Q(zreg[78]) );
  DFF \zreg_reg[79]  ( .D(o[79]), .CLK(clk), .RST(rst), .Q(zreg[79]) );
  DFF \zreg_reg[80]  ( .D(o[80]), .CLK(clk), .RST(rst), .Q(zreg[80]) );
  DFF \zreg_reg[81]  ( .D(o[81]), .CLK(clk), .RST(rst), .Q(zreg[81]) );
  DFF \zreg_reg[82]  ( .D(o[82]), .CLK(clk), .RST(rst), .Q(zreg[82]) );
  DFF \zreg_reg[83]  ( .D(o[83]), .CLK(clk), .RST(rst), .Q(zreg[83]) );
  DFF \zreg_reg[84]  ( .D(o[84]), .CLK(clk), .RST(rst), .Q(zreg[84]) );
  DFF \zreg_reg[85]  ( .D(o[85]), .CLK(clk), .RST(rst), .Q(zreg[85]) );
  DFF \zreg_reg[86]  ( .D(o[86]), .CLK(clk), .RST(rst), .Q(zreg[86]) );
  DFF \zreg_reg[87]  ( .D(o[87]), .CLK(clk), .RST(rst), .Q(zreg[87]) );
  DFF \zreg_reg[88]  ( .D(o[88]), .CLK(clk), .RST(rst), .Q(zreg[88]) );
  DFF \zreg_reg[89]  ( .D(o[89]), .CLK(clk), .RST(rst), .Q(zreg[89]) );
  DFF \zreg_reg[90]  ( .D(o[90]), .CLK(clk), .RST(rst), .Q(zreg[90]) );
  DFF \zreg_reg[91]  ( .D(o[91]), .CLK(clk), .RST(rst), .Q(zreg[91]) );
  DFF \zreg_reg[92]  ( .D(o[92]), .CLK(clk), .RST(rst), .Q(zreg[92]) );
  DFF \zreg_reg[93]  ( .D(o[93]), .CLK(clk), .RST(rst), .Q(zreg[93]) );
  DFF \zreg_reg[94]  ( .D(o[94]), .CLK(clk), .RST(rst), .Q(zreg[94]) );
  DFF \zreg_reg[95]  ( .D(o[95]), .CLK(clk), .RST(rst), .Q(zreg[95]) );
  DFF \zreg_reg[96]  ( .D(o[96]), .CLK(clk), .RST(rst), .Q(zreg[96]) );
  DFF \zreg_reg[97]  ( .D(o[97]), .CLK(clk), .RST(rst), .Q(zreg[97]) );
  DFF \zreg_reg[98]  ( .D(o[98]), .CLK(clk), .RST(rst), .Q(zreg[98]) );
  DFF \zreg_reg[99]  ( .D(o[99]), .CLK(clk), .RST(rst), .Q(zreg[99]) );
  DFF \zreg_reg[100]  ( .D(o[100]), .CLK(clk), .RST(rst), .Q(zreg[100]) );
  DFF \zreg_reg[101]  ( .D(o[101]), .CLK(clk), .RST(rst), .Q(zreg[101]) );
  DFF \zreg_reg[102]  ( .D(o[102]), .CLK(clk), .RST(rst), .Q(zreg[102]) );
  DFF \zreg_reg[103]  ( .D(o[103]), .CLK(clk), .RST(rst), .Q(zreg[103]) );
  DFF \zreg_reg[104]  ( .D(o[104]), .CLK(clk), .RST(rst), .Q(zreg[104]) );
  DFF \zreg_reg[105]  ( .D(o[105]), .CLK(clk), .RST(rst), .Q(zreg[105]) );
  DFF \zreg_reg[106]  ( .D(o[106]), .CLK(clk), .RST(rst), .Q(zreg[106]) );
  DFF \zreg_reg[107]  ( .D(o[107]), .CLK(clk), .RST(rst), .Q(zreg[107]) );
  DFF \zreg_reg[108]  ( .D(o[108]), .CLK(clk), .RST(rst), .Q(zreg[108]) );
  DFF \zreg_reg[109]  ( .D(o[109]), .CLK(clk), .RST(rst), .Q(zreg[109]) );
  DFF \zreg_reg[110]  ( .D(o[110]), .CLK(clk), .RST(rst), .Q(zreg[110]) );
  DFF \zreg_reg[111]  ( .D(o[111]), .CLK(clk), .RST(rst), .Q(zreg[111]) );
  DFF \zreg_reg[112]  ( .D(o[112]), .CLK(clk), .RST(rst), .Q(zreg[112]) );
  DFF \zreg_reg[113]  ( .D(o[113]), .CLK(clk), .RST(rst), .Q(zreg[113]) );
  DFF \zreg_reg[114]  ( .D(o[114]), .CLK(clk), .RST(rst), .Q(zreg[114]) );
  DFF \zreg_reg[115]  ( .D(o[115]), .CLK(clk), .RST(rst), .Q(zreg[115]) );
  DFF \zreg_reg[116]  ( .D(o[116]), .CLK(clk), .RST(rst), .Q(zreg[116]) );
  DFF \zreg_reg[117]  ( .D(o[117]), .CLK(clk), .RST(rst), .Q(zreg[117]) );
  DFF \zreg_reg[118]  ( .D(o[118]), .CLK(clk), .RST(rst), .Q(zreg[118]) );
  DFF \zreg_reg[119]  ( .D(o[119]), .CLK(clk), .RST(rst), .Q(zreg[119]) );
  DFF \zreg_reg[120]  ( .D(o[120]), .CLK(clk), .RST(rst), .Q(zreg[120]) );
  DFF \zreg_reg[121]  ( .D(o[121]), .CLK(clk), .RST(rst), .Q(zreg[121]) );
  DFF \zreg_reg[122]  ( .D(o[122]), .CLK(clk), .RST(rst), .Q(zreg[122]) );
  DFF \zreg_reg[123]  ( .D(o[123]), .CLK(clk), .RST(rst), .Q(zreg[123]) );
  DFF \zreg_reg[124]  ( .D(o[124]), .CLK(clk), .RST(rst), .Q(zreg[124]) );
  DFF \zreg_reg[125]  ( .D(o[125]), .CLK(clk), .RST(rst), .Q(zreg[125]) );
  DFF \zreg_reg[126]  ( .D(o[126]), .CLK(clk), .RST(rst), .Q(zreg[126]) );
  DFF \zreg_reg[127]  ( .D(o[127]), .CLK(clk), .RST(rst), .Q(zreg[127]) );
  DFF \zreg_reg[128]  ( .D(o[128]), .CLK(clk), .RST(rst), .Q(zreg[128]) );
  DFF \zreg_reg[129]  ( .D(o[129]), .CLK(clk), .RST(rst), .Q(zreg[129]) );
  DFF \zreg_reg[130]  ( .D(o[130]), .CLK(clk), .RST(rst), .Q(zreg[130]) );
  DFF \zreg_reg[131]  ( .D(o[131]), .CLK(clk), .RST(rst), .Q(zreg[131]) );
  DFF \zreg_reg[132]  ( .D(o[132]), .CLK(clk), .RST(rst), .Q(zreg[132]) );
  DFF \zreg_reg[133]  ( .D(o[133]), .CLK(clk), .RST(rst), .Q(zreg[133]) );
  DFF \zreg_reg[134]  ( .D(o[134]), .CLK(clk), .RST(rst), .Q(zreg[134]) );
  DFF \zreg_reg[135]  ( .D(o[135]), .CLK(clk), .RST(rst), .Q(zreg[135]) );
  DFF \zreg_reg[136]  ( .D(o[136]), .CLK(clk), .RST(rst), .Q(zreg[136]) );
  DFF \zreg_reg[137]  ( .D(o[137]), .CLK(clk), .RST(rst), .Q(zreg[137]) );
  DFF \zreg_reg[138]  ( .D(o[138]), .CLK(clk), .RST(rst), .Q(zreg[138]) );
  DFF \zreg_reg[139]  ( .D(o[139]), .CLK(clk), .RST(rst), .Q(zreg[139]) );
  DFF \zreg_reg[140]  ( .D(o[140]), .CLK(clk), .RST(rst), .Q(zreg[140]) );
  DFF \zreg_reg[141]  ( .D(o[141]), .CLK(clk), .RST(rst), .Q(zreg[141]) );
  DFF \zreg_reg[142]  ( .D(o[142]), .CLK(clk), .RST(rst), .Q(zreg[142]) );
  DFF \zreg_reg[143]  ( .D(o[143]), .CLK(clk), .RST(rst), .Q(zreg[143]) );
  DFF \zreg_reg[144]  ( .D(o[144]), .CLK(clk), .RST(rst), .Q(zreg[144]) );
  DFF \zreg_reg[145]  ( .D(o[145]), .CLK(clk), .RST(rst), .Q(zreg[145]) );
  DFF \zreg_reg[146]  ( .D(o[146]), .CLK(clk), .RST(rst), .Q(zreg[146]) );
  DFF \zreg_reg[147]  ( .D(o[147]), .CLK(clk), .RST(rst), .Q(zreg[147]) );
  DFF \zreg_reg[148]  ( .D(o[148]), .CLK(clk), .RST(rst), .Q(zreg[148]) );
  DFF \zreg_reg[149]  ( .D(o[149]), .CLK(clk), .RST(rst), .Q(zreg[149]) );
  DFF \zreg_reg[150]  ( .D(o[150]), .CLK(clk), .RST(rst), .Q(zreg[150]) );
  DFF \zreg_reg[151]  ( .D(o[151]), .CLK(clk), .RST(rst), .Q(zreg[151]) );
  DFF \zreg_reg[152]  ( .D(o[152]), .CLK(clk), .RST(rst), .Q(zreg[152]) );
  DFF \zreg_reg[153]  ( .D(o[153]), .CLK(clk), .RST(rst), .Q(zreg[153]) );
  DFF \zreg_reg[154]  ( .D(o[154]), .CLK(clk), .RST(rst), .Q(zreg[154]) );
  DFF \zreg_reg[155]  ( .D(o[155]), .CLK(clk), .RST(rst), .Q(zreg[155]) );
  DFF \zreg_reg[156]  ( .D(o[156]), .CLK(clk), .RST(rst), .Q(zreg[156]) );
  DFF \zreg_reg[157]  ( .D(o[157]), .CLK(clk), .RST(rst), .Q(zreg[157]) );
  DFF \zreg_reg[158]  ( .D(o[158]), .CLK(clk), .RST(rst), .Q(zreg[158]) );
  DFF \zreg_reg[159]  ( .D(o[159]), .CLK(clk), .RST(rst), .Q(zreg[159]) );
  DFF \zreg_reg[160]  ( .D(o[160]), .CLK(clk), .RST(rst), .Q(zreg[160]) );
  DFF \zreg_reg[161]  ( .D(o[161]), .CLK(clk), .RST(rst), .Q(zreg[161]) );
  DFF \zreg_reg[162]  ( .D(o[162]), .CLK(clk), .RST(rst), .Q(zreg[162]) );
  DFF \zreg_reg[163]  ( .D(o[163]), .CLK(clk), .RST(rst), .Q(zreg[163]) );
  DFF \zreg_reg[164]  ( .D(o[164]), .CLK(clk), .RST(rst), .Q(zreg[164]) );
  DFF \zreg_reg[165]  ( .D(o[165]), .CLK(clk), .RST(rst), .Q(zreg[165]) );
  DFF \zreg_reg[166]  ( .D(o[166]), .CLK(clk), .RST(rst), .Q(zreg[166]) );
  DFF \zreg_reg[167]  ( .D(o[167]), .CLK(clk), .RST(rst), .Q(zreg[167]) );
  DFF \zreg_reg[168]  ( .D(o[168]), .CLK(clk), .RST(rst), .Q(zreg[168]) );
  DFF \zreg_reg[169]  ( .D(o[169]), .CLK(clk), .RST(rst), .Q(zreg[169]) );
  DFF \zreg_reg[170]  ( .D(o[170]), .CLK(clk), .RST(rst), .Q(zreg[170]) );
  DFF \zreg_reg[171]  ( .D(o[171]), .CLK(clk), .RST(rst), .Q(zreg[171]) );
  DFF \zreg_reg[172]  ( .D(o[172]), .CLK(clk), .RST(rst), .Q(zreg[172]) );
  DFF \zreg_reg[173]  ( .D(o[173]), .CLK(clk), .RST(rst), .Q(zreg[173]) );
  DFF \zreg_reg[174]  ( .D(o[174]), .CLK(clk), .RST(rst), .Q(zreg[174]) );
  DFF \zreg_reg[175]  ( .D(o[175]), .CLK(clk), .RST(rst), .Q(zreg[175]) );
  DFF \zreg_reg[176]  ( .D(o[176]), .CLK(clk), .RST(rst), .Q(zreg[176]) );
  DFF \zreg_reg[177]  ( .D(o[177]), .CLK(clk), .RST(rst), .Q(zreg[177]) );
  DFF \zreg_reg[178]  ( .D(o[178]), .CLK(clk), .RST(rst), .Q(zreg[178]) );
  DFF \zreg_reg[179]  ( .D(o[179]), .CLK(clk), .RST(rst), .Q(zreg[179]) );
  DFF \zreg_reg[180]  ( .D(o[180]), .CLK(clk), .RST(rst), .Q(zreg[180]) );
  DFF \zreg_reg[181]  ( .D(o[181]), .CLK(clk), .RST(rst), .Q(zreg[181]) );
  DFF \zreg_reg[182]  ( .D(o[182]), .CLK(clk), .RST(rst), .Q(zreg[182]) );
  DFF \zreg_reg[183]  ( .D(o[183]), .CLK(clk), .RST(rst), .Q(zreg[183]) );
  DFF \zreg_reg[184]  ( .D(o[184]), .CLK(clk), .RST(rst), .Q(zreg[184]) );
  DFF \zreg_reg[185]  ( .D(o[185]), .CLK(clk), .RST(rst), .Q(zreg[185]) );
  DFF \zreg_reg[186]  ( .D(o[186]), .CLK(clk), .RST(rst), .Q(zreg[186]) );
  DFF \zreg_reg[187]  ( .D(o[187]), .CLK(clk), .RST(rst), .Q(zreg[187]) );
  DFF \zreg_reg[188]  ( .D(o[188]), .CLK(clk), .RST(rst), .Q(zreg[188]) );
  DFF \zreg_reg[189]  ( .D(o[189]), .CLK(clk), .RST(rst), .Q(zreg[189]) );
  DFF \zreg_reg[190]  ( .D(o[190]), .CLK(clk), .RST(rst), .Q(zreg[190]) );
  DFF \zreg_reg[191]  ( .D(o[191]), .CLK(clk), .RST(rst), .Q(zreg[191]) );
  DFF \zreg_reg[192]  ( .D(o[192]), .CLK(clk), .RST(rst), .Q(zreg[192]) );
  DFF \zreg_reg[193]  ( .D(o[193]), .CLK(clk), .RST(rst), .Q(zreg[193]) );
  DFF \zreg_reg[194]  ( .D(o[194]), .CLK(clk), .RST(rst), .Q(zreg[194]) );
  DFF \zreg_reg[195]  ( .D(o[195]), .CLK(clk), .RST(rst), .Q(zreg[195]) );
  DFF \zreg_reg[196]  ( .D(o[196]), .CLK(clk), .RST(rst), .Q(zreg[196]) );
  DFF \zreg_reg[197]  ( .D(o[197]), .CLK(clk), .RST(rst), .Q(zreg[197]) );
  DFF \zreg_reg[198]  ( .D(o[198]), .CLK(clk), .RST(rst), .Q(zreg[198]) );
  DFF \zreg_reg[199]  ( .D(o[199]), .CLK(clk), .RST(rst), .Q(zreg[199]) );
  DFF \zreg_reg[200]  ( .D(o[200]), .CLK(clk), .RST(rst), .Q(zreg[200]) );
  DFF \zreg_reg[201]  ( .D(o[201]), .CLK(clk), .RST(rst), .Q(zreg[201]) );
  DFF \zreg_reg[202]  ( .D(o[202]), .CLK(clk), .RST(rst), .Q(zreg[202]) );
  DFF \zreg_reg[203]  ( .D(o[203]), .CLK(clk), .RST(rst), .Q(zreg[203]) );
  DFF \zreg_reg[204]  ( .D(o[204]), .CLK(clk), .RST(rst), .Q(zreg[204]) );
  DFF \zreg_reg[205]  ( .D(o[205]), .CLK(clk), .RST(rst), .Q(zreg[205]) );
  DFF \zreg_reg[206]  ( .D(o[206]), .CLK(clk), .RST(rst), .Q(zreg[206]) );
  DFF \zreg_reg[207]  ( .D(o[207]), .CLK(clk), .RST(rst), .Q(zreg[207]) );
  DFF \zreg_reg[208]  ( .D(o[208]), .CLK(clk), .RST(rst), .Q(zreg[208]) );
  DFF \zreg_reg[209]  ( .D(o[209]), .CLK(clk), .RST(rst), .Q(zreg[209]) );
  DFF \zreg_reg[210]  ( .D(o[210]), .CLK(clk), .RST(rst), .Q(zreg[210]) );
  DFF \zreg_reg[211]  ( .D(o[211]), .CLK(clk), .RST(rst), .Q(zreg[211]) );
  DFF \zreg_reg[212]  ( .D(o[212]), .CLK(clk), .RST(rst), .Q(zreg[212]) );
  DFF \zreg_reg[213]  ( .D(o[213]), .CLK(clk), .RST(rst), .Q(zreg[213]) );
  DFF \zreg_reg[214]  ( .D(o[214]), .CLK(clk), .RST(rst), .Q(zreg[214]) );
  DFF \zreg_reg[215]  ( .D(o[215]), .CLK(clk), .RST(rst), .Q(zreg[215]) );
  DFF \zreg_reg[216]  ( .D(o[216]), .CLK(clk), .RST(rst), .Q(zreg[216]) );
  DFF \zreg_reg[217]  ( .D(o[217]), .CLK(clk), .RST(rst), .Q(zreg[217]) );
  DFF \zreg_reg[218]  ( .D(o[218]), .CLK(clk), .RST(rst), .Q(zreg[218]) );
  DFF \zreg_reg[219]  ( .D(o[219]), .CLK(clk), .RST(rst), .Q(zreg[219]) );
  DFF \zreg_reg[220]  ( .D(o[220]), .CLK(clk), .RST(rst), .Q(zreg[220]) );
  DFF \zreg_reg[221]  ( .D(o[221]), .CLK(clk), .RST(rst), .Q(zreg[221]) );
  DFF \zreg_reg[222]  ( .D(o[222]), .CLK(clk), .RST(rst), .Q(zreg[222]) );
  DFF \zreg_reg[223]  ( .D(o[223]), .CLK(clk), .RST(rst), .Q(zreg[223]) );
  DFF \zreg_reg[224]  ( .D(o[224]), .CLK(clk), .RST(rst), .Q(zreg[224]) );
  DFF \zreg_reg[225]  ( .D(o[225]), .CLK(clk), .RST(rst), .Q(zreg[225]) );
  DFF \zreg_reg[226]  ( .D(o[226]), .CLK(clk), .RST(rst), .Q(zreg[226]) );
  DFF \zreg_reg[227]  ( .D(o[227]), .CLK(clk), .RST(rst), .Q(zreg[227]) );
  DFF \zreg_reg[228]  ( .D(o[228]), .CLK(clk), .RST(rst), .Q(zreg[228]) );
  DFF \zreg_reg[229]  ( .D(o[229]), .CLK(clk), .RST(rst), .Q(zreg[229]) );
  DFF \zreg_reg[230]  ( .D(o[230]), .CLK(clk), .RST(rst), .Q(zreg[230]) );
  DFF \zreg_reg[231]  ( .D(o[231]), .CLK(clk), .RST(rst), .Q(zreg[231]) );
  DFF \zreg_reg[232]  ( .D(o[232]), .CLK(clk), .RST(rst), .Q(zreg[232]) );
  DFF \zreg_reg[233]  ( .D(o[233]), .CLK(clk), .RST(rst), .Q(zreg[233]) );
  DFF \zreg_reg[234]  ( .D(o[234]), .CLK(clk), .RST(rst), .Q(zreg[234]) );
  DFF \zreg_reg[235]  ( .D(o[235]), .CLK(clk), .RST(rst), .Q(zreg[235]) );
  DFF \zreg_reg[236]  ( .D(o[236]), .CLK(clk), .RST(rst), .Q(zreg[236]) );
  DFF \zreg_reg[237]  ( .D(o[237]), .CLK(clk), .RST(rst), .Q(zreg[237]) );
  DFF \zreg_reg[238]  ( .D(o[238]), .CLK(clk), .RST(rst), .Q(zreg[238]) );
  DFF \zreg_reg[239]  ( .D(o[239]), .CLK(clk), .RST(rst), .Q(zreg[239]) );
  DFF \zreg_reg[240]  ( .D(o[240]), .CLK(clk), .RST(rst), .Q(zreg[240]) );
  DFF \zreg_reg[241]  ( .D(o[241]), .CLK(clk), .RST(rst), .Q(zreg[241]) );
  DFF \zreg_reg[242]  ( .D(o[242]), .CLK(clk), .RST(rst), .Q(zreg[242]) );
  DFF \zreg_reg[243]  ( .D(o[243]), .CLK(clk), .RST(rst), .Q(zreg[243]) );
  DFF \zreg_reg[244]  ( .D(o[244]), .CLK(clk), .RST(rst), .Q(zreg[244]) );
  DFF \zreg_reg[245]  ( .D(o[245]), .CLK(clk), .RST(rst), .Q(zreg[245]) );
  DFF \zreg_reg[246]  ( .D(o[246]), .CLK(clk), .RST(rst), .Q(zreg[246]) );
  DFF \zreg_reg[247]  ( .D(o[247]), .CLK(clk), .RST(rst), .Q(zreg[247]) );
  DFF \zreg_reg[248]  ( .D(o[248]), .CLK(clk), .RST(rst), .Q(zreg[248]) );
  DFF \zreg_reg[249]  ( .D(o[249]), .CLK(clk), .RST(rst), .Q(zreg[249]) );
  DFF \zreg_reg[250]  ( .D(o[250]), .CLK(clk), .RST(rst), .Q(zreg[250]) );
  DFF \zreg_reg[251]  ( .D(o[251]), .CLK(clk), .RST(rst), .Q(zreg[251]) );
  DFF \zreg_reg[252]  ( .D(o[252]), .CLK(clk), .RST(rst), .Q(zreg[252]) );
  DFF \zreg_reg[253]  ( .D(o[253]), .CLK(clk), .RST(rst), .Q(zreg[253]) );
  DFF \zreg_reg[254]  ( .D(o[254]), .CLK(clk), .RST(rst), .Q(zreg[254]) );
  DFF \zreg_reg[255]  ( .D(o[255]), .CLK(clk), .RST(rst), .Q(zreg[255]) );
  DFF \zreg_reg[256]  ( .D(\zout[3][256] ), .CLK(clk), .RST(rst), .Q(zreg[256]) );
  DFF \zreg_reg[257]  ( .D(\zout[3][257] ), .CLK(clk), .RST(rst), .Q(zreg[257]) );
  modmult_step_N256_2 \MODMULT_STEP[0].modmult_step_  ( .xregN_1(xin[255]), 
        .y(y), .n(n), .zin({\zin[0][257] , \zin[0][256] , \zin[0][255] , 
        \zin[0][254] , \zin[0][253] , \zin[0][252] , \zin[0][251] , 
        \zin[0][250] , \zin[0][249] , \zin[0][248] , \zin[0][247] , 
        \zin[0][246] , \zin[0][245] , \zin[0][244] , \zin[0][243] , 
        \zin[0][242] , \zin[0][241] , \zin[0][240] , \zin[0][239] , 
        \zin[0][238] , \zin[0][237] , \zin[0][236] , \zin[0][235] , 
        \zin[0][234] , \zin[0][233] , \zin[0][232] , \zin[0][231] , 
        \zin[0][230] , \zin[0][229] , \zin[0][228] , \zin[0][227] , 
        \zin[0][226] , \zin[0][225] , \zin[0][224] , \zin[0][223] , 
        \zin[0][222] , \zin[0][221] , \zin[0][220] , \zin[0][219] , 
        \zin[0][218] , \zin[0][217] , \zin[0][216] , \zin[0][215] , 
        \zin[0][214] , \zin[0][213] , \zin[0][212] , \zin[0][211] , 
        \zin[0][210] , \zin[0][209] , \zin[0][208] , \zin[0][207] , 
        \zin[0][206] , \zin[0][205] , \zin[0][204] , \zin[0][203] , 
        \zin[0][202] , \zin[0][201] , \zin[0][200] , \zin[0][199] , 
        \zin[0][198] , \zin[0][197] , \zin[0][196] , \zin[0][195] , 
        \zin[0][194] , \zin[0][193] , \zin[0][192] , \zin[0][191] , 
        \zin[0][190] , \zin[0][189] , \zin[0][188] , \zin[0][187] , 
        \zin[0][186] , \zin[0][185] , \zin[0][184] , \zin[0][183] , 
        \zin[0][182] , \zin[0][181] , \zin[0][180] , \zin[0][179] , 
        \zin[0][178] , \zin[0][177] , \zin[0][176] , \zin[0][175] , 
        \zin[0][174] , \zin[0][173] , \zin[0][172] , \zin[0][171] , 
        \zin[0][170] , \zin[0][169] , \zin[0][168] , \zin[0][167] , 
        \zin[0][166] , \zin[0][165] , \zin[0][164] , \zin[0][163] , 
        \zin[0][162] , \zin[0][161] , \zin[0][160] , \zin[0][159] , 
        \zin[0][158] , \zin[0][157] , \zin[0][156] , \zin[0][155] , 
        \zin[0][154] , \zin[0][153] , \zin[0][152] , \zin[0][151] , 
        \zin[0][150] , \zin[0][149] , \zin[0][148] , \zin[0][147] , 
        \zin[0][146] , \zin[0][145] , \zin[0][144] , \zin[0][143] , 
        \zin[0][142] , \zin[0][141] , \zin[0][140] , \zin[0][139] , 
        \zin[0][138] , \zin[0][137] , \zin[0][136] , \zin[0][135] , 
        \zin[0][134] , \zin[0][133] , \zin[0][132] , \zin[0][131] , 
        \zin[0][130] , \zin[0][129] , \zin[0][128] , \zin[0][127] , 
        \zin[0][126] , \zin[0][125] , \zin[0][124] , \zin[0][123] , 
        \zin[0][122] , \zin[0][121] , \zin[0][120] , \zin[0][119] , 
        \zin[0][118] , \zin[0][117] , \zin[0][116] , \zin[0][115] , 
        \zin[0][114] , \zin[0][113] , \zin[0][112] , \zin[0][111] , 
        \zin[0][110] , \zin[0][109] , \zin[0][108] , \zin[0][107] , 
        \zin[0][106] , \zin[0][105] , \zin[0][104] , \zin[0][103] , 
        \zin[0][102] , \zin[0][101] , \zin[0][100] , \zin[0][99] , 
        \zin[0][98] , \zin[0][97] , \zin[0][96] , \zin[0][95] , \zin[0][94] , 
        \zin[0][93] , \zin[0][92] , \zin[0][91] , \zin[0][90] , \zin[0][89] , 
        \zin[0][88] , \zin[0][87] , \zin[0][86] , \zin[0][85] , \zin[0][84] , 
        \zin[0][83] , \zin[0][82] , \zin[0][81] , \zin[0][80] , \zin[0][79] , 
        \zin[0][78] , \zin[0][77] , \zin[0][76] , \zin[0][75] , \zin[0][74] , 
        \zin[0][73] , \zin[0][72] , \zin[0][71] , \zin[0][70] , \zin[0][69] , 
        \zin[0][68] , \zin[0][67] , \zin[0][66] , \zin[0][65] , \zin[0][64] , 
        \zin[0][63] , \zin[0][62] , \zin[0][61] , \zin[0][60] , \zin[0][59] , 
        \zin[0][58] , \zin[0][57] , \zin[0][56] , \zin[0][55] , \zin[0][54] , 
        \zin[0][53] , \zin[0][52] , \zin[0][51] , \zin[0][50] , \zin[0][49] , 
        \zin[0][48] , \zin[0][47] , \zin[0][46] , \zin[0][45] , \zin[0][44] , 
        \zin[0][43] , \zin[0][42] , \zin[0][41] , \zin[0][40] , \zin[0][39] , 
        \zin[0][38] , \zin[0][37] , \zin[0][36] , \zin[0][35] , \zin[0][34] , 
        \zin[0][33] , \zin[0][32] , \zin[0][31] , \zin[0][30] , \zin[0][29] , 
        \zin[0][28] , \zin[0][27] , \zin[0][26] , \zin[0][25] , \zin[0][24] , 
        \zin[0][23] , \zin[0][22] , \zin[0][21] , \zin[0][20] , \zin[0][19] , 
        \zin[0][18] , \zin[0][17] , \zin[0][16] , \zin[0][15] , \zin[0][14] , 
        \zin[0][13] , \zin[0][12] , \zin[0][11] , \zin[0][10] , \zin[0][9] , 
        \zin[0][8] , \zin[0][7] , \zin[0][6] , \zin[0][5] , \zin[0][4] , 
        \zin[0][3] , \zin[0][2] , \zin[0][1] , \zin[0][0] }), .zout({
        \zin[1][257] , \zin[1][256] , \zin[1][255] , \zin[1][254] , 
        \zin[1][253] , \zin[1][252] , \zin[1][251] , \zin[1][250] , 
        \zin[1][249] , \zin[1][248] , \zin[1][247] , \zin[1][246] , 
        \zin[1][245] , \zin[1][244] , \zin[1][243] , \zin[1][242] , 
        \zin[1][241] , \zin[1][240] , \zin[1][239] , \zin[1][238] , 
        \zin[1][237] , \zin[1][236] , \zin[1][235] , \zin[1][234] , 
        \zin[1][233] , \zin[1][232] , \zin[1][231] , \zin[1][230] , 
        \zin[1][229] , \zin[1][228] , \zin[1][227] , \zin[1][226] , 
        \zin[1][225] , \zin[1][224] , \zin[1][223] , \zin[1][222] , 
        \zin[1][221] , \zin[1][220] , \zin[1][219] , \zin[1][218] , 
        \zin[1][217] , \zin[1][216] , \zin[1][215] , \zin[1][214] , 
        \zin[1][213] , \zin[1][212] , \zin[1][211] , \zin[1][210] , 
        \zin[1][209] , \zin[1][208] , \zin[1][207] , \zin[1][206] , 
        \zin[1][205] , \zin[1][204] , \zin[1][203] , \zin[1][202] , 
        \zin[1][201] , \zin[1][200] , \zin[1][199] , \zin[1][198] , 
        \zin[1][197] , \zin[1][196] , \zin[1][195] , \zin[1][194] , 
        \zin[1][193] , \zin[1][192] , \zin[1][191] , \zin[1][190] , 
        \zin[1][189] , \zin[1][188] , \zin[1][187] , \zin[1][186] , 
        \zin[1][185] , \zin[1][184] , \zin[1][183] , \zin[1][182] , 
        \zin[1][181] , \zin[1][180] , \zin[1][179] , \zin[1][178] , 
        \zin[1][177] , \zin[1][176] , \zin[1][175] , \zin[1][174] , 
        \zin[1][173] , \zin[1][172] , \zin[1][171] , \zin[1][170] , 
        \zin[1][169] , \zin[1][168] , \zin[1][167] , \zin[1][166] , 
        \zin[1][165] , \zin[1][164] , \zin[1][163] , \zin[1][162] , 
        \zin[1][161] , \zin[1][160] , \zin[1][159] , \zin[1][158] , 
        \zin[1][157] , \zin[1][156] , \zin[1][155] , \zin[1][154] , 
        \zin[1][153] , \zin[1][152] , \zin[1][151] , \zin[1][150] , 
        \zin[1][149] , \zin[1][148] , \zin[1][147] , \zin[1][146] , 
        \zin[1][145] , \zin[1][144] , \zin[1][143] , \zin[1][142] , 
        \zin[1][141] , \zin[1][140] , \zin[1][139] , \zin[1][138] , 
        \zin[1][137] , \zin[1][136] , \zin[1][135] , \zin[1][134] , 
        \zin[1][133] , \zin[1][132] , \zin[1][131] , \zin[1][130] , 
        \zin[1][129] , \zin[1][128] , \zin[1][127] , \zin[1][126] , 
        \zin[1][125] , \zin[1][124] , \zin[1][123] , \zin[1][122] , 
        \zin[1][121] , \zin[1][120] , \zin[1][119] , \zin[1][118] , 
        \zin[1][117] , \zin[1][116] , \zin[1][115] , \zin[1][114] , 
        \zin[1][113] , \zin[1][112] , \zin[1][111] , \zin[1][110] , 
        \zin[1][109] , \zin[1][108] , \zin[1][107] , \zin[1][106] , 
        \zin[1][105] , \zin[1][104] , \zin[1][103] , \zin[1][102] , 
        \zin[1][101] , \zin[1][100] , \zin[1][99] , \zin[1][98] , \zin[1][97] , 
        \zin[1][96] , \zin[1][95] , \zin[1][94] , \zin[1][93] , \zin[1][92] , 
        \zin[1][91] , \zin[1][90] , \zin[1][89] , \zin[1][88] , \zin[1][87] , 
        \zin[1][86] , \zin[1][85] , \zin[1][84] , \zin[1][83] , \zin[1][82] , 
        \zin[1][81] , \zin[1][80] , \zin[1][79] , \zin[1][78] , \zin[1][77] , 
        \zin[1][76] , \zin[1][75] , \zin[1][74] , \zin[1][73] , \zin[1][72] , 
        \zin[1][71] , \zin[1][70] , \zin[1][69] , \zin[1][68] , \zin[1][67] , 
        \zin[1][66] , \zin[1][65] , \zin[1][64] , \zin[1][63] , \zin[1][62] , 
        \zin[1][61] , \zin[1][60] , \zin[1][59] , \zin[1][58] , \zin[1][57] , 
        \zin[1][56] , \zin[1][55] , \zin[1][54] , \zin[1][53] , \zin[1][52] , 
        \zin[1][51] , \zin[1][50] , \zin[1][49] , \zin[1][48] , \zin[1][47] , 
        \zin[1][46] , \zin[1][45] , \zin[1][44] , \zin[1][43] , \zin[1][42] , 
        \zin[1][41] , \zin[1][40] , \zin[1][39] , \zin[1][38] , \zin[1][37] , 
        \zin[1][36] , \zin[1][35] , \zin[1][34] , \zin[1][33] , \zin[1][32] , 
        \zin[1][31] , \zin[1][30] , \zin[1][29] , \zin[1][28] , \zin[1][27] , 
        \zin[1][26] , \zin[1][25] , \zin[1][24] , \zin[1][23] , \zin[1][22] , 
        \zin[1][21] , \zin[1][20] , \zin[1][19] , \zin[1][18] , \zin[1][17] , 
        \zin[1][16] , \zin[1][15] , \zin[1][14] , \zin[1][13] , \zin[1][12] , 
        \zin[1][11] , \zin[1][10] , \zin[1][9] , \zin[1][8] , \zin[1][7] , 
        \zin[1][6] , \zin[1][5] , \zin[1][4] , \zin[1][3] , \zin[1][2] , 
        \zin[1][1] , \zin[1][0] }) );
  modmult_step_N256_5 \MODMULT_STEP[1].modmult_step_  ( .xregN_1(xin[254]), 
        .y(y), .n(n), .zin({\zin[1][257] , \zin[1][256] , \zin[1][255] , 
        \zin[1][254] , \zin[1][253] , \zin[1][252] , \zin[1][251] , 
        \zin[1][250] , \zin[1][249] , \zin[1][248] , \zin[1][247] , 
        \zin[1][246] , \zin[1][245] , \zin[1][244] , \zin[1][243] , 
        \zin[1][242] , \zin[1][241] , \zin[1][240] , \zin[1][239] , 
        \zin[1][238] , \zin[1][237] , \zin[1][236] , \zin[1][235] , 
        \zin[1][234] , \zin[1][233] , \zin[1][232] , \zin[1][231] , 
        \zin[1][230] , \zin[1][229] , \zin[1][228] , \zin[1][227] , 
        \zin[1][226] , \zin[1][225] , \zin[1][224] , \zin[1][223] , 
        \zin[1][222] , \zin[1][221] , \zin[1][220] , \zin[1][219] , 
        \zin[1][218] , \zin[1][217] , \zin[1][216] , \zin[1][215] , 
        \zin[1][214] , \zin[1][213] , \zin[1][212] , \zin[1][211] , 
        \zin[1][210] , \zin[1][209] , \zin[1][208] , \zin[1][207] , 
        \zin[1][206] , \zin[1][205] , \zin[1][204] , \zin[1][203] , 
        \zin[1][202] , \zin[1][201] , \zin[1][200] , \zin[1][199] , 
        \zin[1][198] , \zin[1][197] , \zin[1][196] , \zin[1][195] , 
        \zin[1][194] , \zin[1][193] , \zin[1][192] , \zin[1][191] , 
        \zin[1][190] , \zin[1][189] , \zin[1][188] , \zin[1][187] , 
        \zin[1][186] , \zin[1][185] , \zin[1][184] , \zin[1][183] , 
        \zin[1][182] , \zin[1][181] , \zin[1][180] , \zin[1][179] , 
        \zin[1][178] , \zin[1][177] , \zin[1][176] , \zin[1][175] , 
        \zin[1][174] , \zin[1][173] , \zin[1][172] , \zin[1][171] , 
        \zin[1][170] , \zin[1][169] , \zin[1][168] , \zin[1][167] , 
        \zin[1][166] , \zin[1][165] , \zin[1][164] , \zin[1][163] , 
        \zin[1][162] , \zin[1][161] , \zin[1][160] , \zin[1][159] , 
        \zin[1][158] , \zin[1][157] , \zin[1][156] , \zin[1][155] , 
        \zin[1][154] , \zin[1][153] , \zin[1][152] , \zin[1][151] , 
        \zin[1][150] , \zin[1][149] , \zin[1][148] , \zin[1][147] , 
        \zin[1][146] , \zin[1][145] , \zin[1][144] , \zin[1][143] , 
        \zin[1][142] , \zin[1][141] , \zin[1][140] , \zin[1][139] , 
        \zin[1][138] , \zin[1][137] , \zin[1][136] , \zin[1][135] , 
        \zin[1][134] , \zin[1][133] , \zin[1][132] , \zin[1][131] , 
        \zin[1][130] , \zin[1][129] , \zin[1][128] , \zin[1][127] , 
        \zin[1][126] , \zin[1][125] , \zin[1][124] , \zin[1][123] , 
        \zin[1][122] , \zin[1][121] , \zin[1][120] , \zin[1][119] , 
        \zin[1][118] , \zin[1][117] , \zin[1][116] , \zin[1][115] , 
        \zin[1][114] , \zin[1][113] , \zin[1][112] , \zin[1][111] , 
        \zin[1][110] , \zin[1][109] , \zin[1][108] , \zin[1][107] , 
        \zin[1][106] , \zin[1][105] , \zin[1][104] , \zin[1][103] , 
        \zin[1][102] , \zin[1][101] , \zin[1][100] , \zin[1][99] , 
        \zin[1][98] , \zin[1][97] , \zin[1][96] , \zin[1][95] , \zin[1][94] , 
        \zin[1][93] , \zin[1][92] , \zin[1][91] , \zin[1][90] , \zin[1][89] , 
        \zin[1][88] , \zin[1][87] , \zin[1][86] , \zin[1][85] , \zin[1][84] , 
        \zin[1][83] , \zin[1][82] , \zin[1][81] , \zin[1][80] , \zin[1][79] , 
        \zin[1][78] , \zin[1][77] , \zin[1][76] , \zin[1][75] , \zin[1][74] , 
        \zin[1][73] , \zin[1][72] , \zin[1][71] , \zin[1][70] , \zin[1][69] , 
        \zin[1][68] , \zin[1][67] , \zin[1][66] , \zin[1][65] , \zin[1][64] , 
        \zin[1][63] , \zin[1][62] , \zin[1][61] , \zin[1][60] , \zin[1][59] , 
        \zin[1][58] , \zin[1][57] , \zin[1][56] , \zin[1][55] , \zin[1][54] , 
        \zin[1][53] , \zin[1][52] , \zin[1][51] , \zin[1][50] , \zin[1][49] , 
        \zin[1][48] , \zin[1][47] , \zin[1][46] , \zin[1][45] , \zin[1][44] , 
        \zin[1][43] , \zin[1][42] , \zin[1][41] , \zin[1][40] , \zin[1][39] , 
        \zin[1][38] , \zin[1][37] , \zin[1][36] , \zin[1][35] , \zin[1][34] , 
        \zin[1][33] , \zin[1][32] , \zin[1][31] , \zin[1][30] , \zin[1][29] , 
        \zin[1][28] , \zin[1][27] , \zin[1][26] , \zin[1][25] , \zin[1][24] , 
        \zin[1][23] , \zin[1][22] , \zin[1][21] , \zin[1][20] , \zin[1][19] , 
        \zin[1][18] , \zin[1][17] , \zin[1][16] , \zin[1][15] , \zin[1][14] , 
        \zin[1][13] , \zin[1][12] , \zin[1][11] , \zin[1][10] , \zin[1][9] , 
        \zin[1][8] , \zin[1][7] , \zin[1][6] , \zin[1][5] , \zin[1][4] , 
        \zin[1][3] , \zin[1][2] , \zin[1][1] , \zin[1][0] }), .zout({
        \zin[2][257] , \zin[2][256] , \zin[2][255] , \zin[2][254] , 
        \zin[2][253] , \zin[2][252] , \zin[2][251] , \zin[2][250] , 
        \zin[2][249] , \zin[2][248] , \zin[2][247] , \zin[2][246] , 
        \zin[2][245] , \zin[2][244] , \zin[2][243] , \zin[2][242] , 
        \zin[2][241] , \zin[2][240] , \zin[2][239] , \zin[2][238] , 
        \zin[2][237] , \zin[2][236] , \zin[2][235] , \zin[2][234] , 
        \zin[2][233] , \zin[2][232] , \zin[2][231] , \zin[2][230] , 
        \zin[2][229] , \zin[2][228] , \zin[2][227] , \zin[2][226] , 
        \zin[2][225] , \zin[2][224] , \zin[2][223] , \zin[2][222] , 
        \zin[2][221] , \zin[2][220] , \zin[2][219] , \zin[2][218] , 
        \zin[2][217] , \zin[2][216] , \zin[2][215] , \zin[2][214] , 
        \zin[2][213] , \zin[2][212] , \zin[2][211] , \zin[2][210] , 
        \zin[2][209] , \zin[2][208] , \zin[2][207] , \zin[2][206] , 
        \zin[2][205] , \zin[2][204] , \zin[2][203] , \zin[2][202] , 
        \zin[2][201] , \zin[2][200] , \zin[2][199] , \zin[2][198] , 
        \zin[2][197] , \zin[2][196] , \zin[2][195] , \zin[2][194] , 
        \zin[2][193] , \zin[2][192] , \zin[2][191] , \zin[2][190] , 
        \zin[2][189] , \zin[2][188] , \zin[2][187] , \zin[2][186] , 
        \zin[2][185] , \zin[2][184] , \zin[2][183] , \zin[2][182] , 
        \zin[2][181] , \zin[2][180] , \zin[2][179] , \zin[2][178] , 
        \zin[2][177] , \zin[2][176] , \zin[2][175] , \zin[2][174] , 
        \zin[2][173] , \zin[2][172] , \zin[2][171] , \zin[2][170] , 
        \zin[2][169] , \zin[2][168] , \zin[2][167] , \zin[2][166] , 
        \zin[2][165] , \zin[2][164] , \zin[2][163] , \zin[2][162] , 
        \zin[2][161] , \zin[2][160] , \zin[2][159] , \zin[2][158] , 
        \zin[2][157] , \zin[2][156] , \zin[2][155] , \zin[2][154] , 
        \zin[2][153] , \zin[2][152] , \zin[2][151] , \zin[2][150] , 
        \zin[2][149] , \zin[2][148] , \zin[2][147] , \zin[2][146] , 
        \zin[2][145] , \zin[2][144] , \zin[2][143] , \zin[2][142] , 
        \zin[2][141] , \zin[2][140] , \zin[2][139] , \zin[2][138] , 
        \zin[2][137] , \zin[2][136] , \zin[2][135] , \zin[2][134] , 
        \zin[2][133] , \zin[2][132] , \zin[2][131] , \zin[2][130] , 
        \zin[2][129] , \zin[2][128] , \zin[2][127] , \zin[2][126] , 
        \zin[2][125] , \zin[2][124] , \zin[2][123] , \zin[2][122] , 
        \zin[2][121] , \zin[2][120] , \zin[2][119] , \zin[2][118] , 
        \zin[2][117] , \zin[2][116] , \zin[2][115] , \zin[2][114] , 
        \zin[2][113] , \zin[2][112] , \zin[2][111] , \zin[2][110] , 
        \zin[2][109] , \zin[2][108] , \zin[2][107] , \zin[2][106] , 
        \zin[2][105] , \zin[2][104] , \zin[2][103] , \zin[2][102] , 
        \zin[2][101] , \zin[2][100] , \zin[2][99] , \zin[2][98] , \zin[2][97] , 
        \zin[2][96] , \zin[2][95] , \zin[2][94] , \zin[2][93] , \zin[2][92] , 
        \zin[2][91] , \zin[2][90] , \zin[2][89] , \zin[2][88] , \zin[2][87] , 
        \zin[2][86] , \zin[2][85] , \zin[2][84] , \zin[2][83] , \zin[2][82] , 
        \zin[2][81] , \zin[2][80] , \zin[2][79] , \zin[2][78] , \zin[2][77] , 
        \zin[2][76] , \zin[2][75] , \zin[2][74] , \zin[2][73] , \zin[2][72] , 
        \zin[2][71] , \zin[2][70] , \zin[2][69] , \zin[2][68] , \zin[2][67] , 
        \zin[2][66] , \zin[2][65] , \zin[2][64] , \zin[2][63] , \zin[2][62] , 
        \zin[2][61] , \zin[2][60] , \zin[2][59] , \zin[2][58] , \zin[2][57] , 
        \zin[2][56] , \zin[2][55] , \zin[2][54] , \zin[2][53] , \zin[2][52] , 
        \zin[2][51] , \zin[2][50] , \zin[2][49] , \zin[2][48] , \zin[2][47] , 
        \zin[2][46] , \zin[2][45] , \zin[2][44] , \zin[2][43] , \zin[2][42] , 
        \zin[2][41] , \zin[2][40] , \zin[2][39] , \zin[2][38] , \zin[2][37] , 
        \zin[2][36] , \zin[2][35] , \zin[2][34] , \zin[2][33] , \zin[2][32] , 
        \zin[2][31] , \zin[2][30] , \zin[2][29] , \zin[2][28] , \zin[2][27] , 
        \zin[2][26] , \zin[2][25] , \zin[2][24] , \zin[2][23] , \zin[2][22] , 
        \zin[2][21] , \zin[2][20] , \zin[2][19] , \zin[2][18] , \zin[2][17] , 
        \zin[2][16] , \zin[2][15] , \zin[2][14] , \zin[2][13] , \zin[2][12] , 
        \zin[2][11] , \zin[2][10] , \zin[2][9] , \zin[2][8] , \zin[2][7] , 
        \zin[2][6] , \zin[2][5] , \zin[2][4] , \zin[2][3] , \zin[2][2] , 
        \zin[2][1] , \zin[2][0] }) );
  modmult_step_N256_4 \MODMULT_STEP[2].modmult_step_  ( .xregN_1(xin[253]), 
        .y(y), .n(n), .zin({\zin[2][257] , \zin[2][256] , \zin[2][255] , 
        \zin[2][254] , \zin[2][253] , \zin[2][252] , \zin[2][251] , 
        \zin[2][250] , \zin[2][249] , \zin[2][248] , \zin[2][247] , 
        \zin[2][246] , \zin[2][245] , \zin[2][244] , \zin[2][243] , 
        \zin[2][242] , \zin[2][241] , \zin[2][240] , \zin[2][239] , 
        \zin[2][238] , \zin[2][237] , \zin[2][236] , \zin[2][235] , 
        \zin[2][234] , \zin[2][233] , \zin[2][232] , \zin[2][231] , 
        \zin[2][230] , \zin[2][229] , \zin[2][228] , \zin[2][227] , 
        \zin[2][226] , \zin[2][225] , \zin[2][224] , \zin[2][223] , 
        \zin[2][222] , \zin[2][221] , \zin[2][220] , \zin[2][219] , 
        \zin[2][218] , \zin[2][217] , \zin[2][216] , \zin[2][215] , 
        \zin[2][214] , \zin[2][213] , \zin[2][212] , \zin[2][211] , 
        \zin[2][210] , \zin[2][209] , \zin[2][208] , \zin[2][207] , 
        \zin[2][206] , \zin[2][205] , \zin[2][204] , \zin[2][203] , 
        \zin[2][202] , \zin[2][201] , \zin[2][200] , \zin[2][199] , 
        \zin[2][198] , \zin[2][197] , \zin[2][196] , \zin[2][195] , 
        \zin[2][194] , \zin[2][193] , \zin[2][192] , \zin[2][191] , 
        \zin[2][190] , \zin[2][189] , \zin[2][188] , \zin[2][187] , 
        \zin[2][186] , \zin[2][185] , \zin[2][184] , \zin[2][183] , 
        \zin[2][182] , \zin[2][181] , \zin[2][180] , \zin[2][179] , 
        \zin[2][178] , \zin[2][177] , \zin[2][176] , \zin[2][175] , 
        \zin[2][174] , \zin[2][173] , \zin[2][172] , \zin[2][171] , 
        \zin[2][170] , \zin[2][169] , \zin[2][168] , \zin[2][167] , 
        \zin[2][166] , \zin[2][165] , \zin[2][164] , \zin[2][163] , 
        \zin[2][162] , \zin[2][161] , \zin[2][160] , \zin[2][159] , 
        \zin[2][158] , \zin[2][157] , \zin[2][156] , \zin[2][155] , 
        \zin[2][154] , \zin[2][153] , \zin[2][152] , \zin[2][151] , 
        \zin[2][150] , \zin[2][149] , \zin[2][148] , \zin[2][147] , 
        \zin[2][146] , \zin[2][145] , \zin[2][144] , \zin[2][143] , 
        \zin[2][142] , \zin[2][141] , \zin[2][140] , \zin[2][139] , 
        \zin[2][138] , \zin[2][137] , \zin[2][136] , \zin[2][135] , 
        \zin[2][134] , \zin[2][133] , \zin[2][132] , \zin[2][131] , 
        \zin[2][130] , \zin[2][129] , \zin[2][128] , \zin[2][127] , 
        \zin[2][126] , \zin[2][125] , \zin[2][124] , \zin[2][123] , 
        \zin[2][122] , \zin[2][121] , \zin[2][120] , \zin[2][119] , 
        \zin[2][118] , \zin[2][117] , \zin[2][116] , \zin[2][115] , 
        \zin[2][114] , \zin[2][113] , \zin[2][112] , \zin[2][111] , 
        \zin[2][110] , \zin[2][109] , \zin[2][108] , \zin[2][107] , 
        \zin[2][106] , \zin[2][105] , \zin[2][104] , \zin[2][103] , 
        \zin[2][102] , \zin[2][101] , \zin[2][100] , \zin[2][99] , 
        \zin[2][98] , \zin[2][97] , \zin[2][96] , \zin[2][95] , \zin[2][94] , 
        \zin[2][93] , \zin[2][92] , \zin[2][91] , \zin[2][90] , \zin[2][89] , 
        \zin[2][88] , \zin[2][87] , \zin[2][86] , \zin[2][85] , \zin[2][84] , 
        \zin[2][83] , \zin[2][82] , \zin[2][81] , \zin[2][80] , \zin[2][79] , 
        \zin[2][78] , \zin[2][77] , \zin[2][76] , \zin[2][75] , \zin[2][74] , 
        \zin[2][73] , \zin[2][72] , \zin[2][71] , \zin[2][70] , \zin[2][69] , 
        \zin[2][68] , \zin[2][67] , \zin[2][66] , \zin[2][65] , \zin[2][64] , 
        \zin[2][63] , \zin[2][62] , \zin[2][61] , \zin[2][60] , \zin[2][59] , 
        \zin[2][58] , \zin[2][57] , \zin[2][56] , \zin[2][55] , \zin[2][54] , 
        \zin[2][53] , \zin[2][52] , \zin[2][51] , \zin[2][50] , \zin[2][49] , 
        \zin[2][48] , \zin[2][47] , \zin[2][46] , \zin[2][45] , \zin[2][44] , 
        \zin[2][43] , \zin[2][42] , \zin[2][41] , \zin[2][40] , \zin[2][39] , 
        \zin[2][38] , \zin[2][37] , \zin[2][36] , \zin[2][35] , \zin[2][34] , 
        \zin[2][33] , \zin[2][32] , \zin[2][31] , \zin[2][30] , \zin[2][29] , 
        \zin[2][28] , \zin[2][27] , \zin[2][26] , \zin[2][25] , \zin[2][24] , 
        \zin[2][23] , \zin[2][22] , \zin[2][21] , \zin[2][20] , \zin[2][19] , 
        \zin[2][18] , \zin[2][17] , \zin[2][16] , \zin[2][15] , \zin[2][14] , 
        \zin[2][13] , \zin[2][12] , \zin[2][11] , \zin[2][10] , \zin[2][9] , 
        \zin[2][8] , \zin[2][7] , \zin[2][6] , \zin[2][5] , \zin[2][4] , 
        \zin[2][3] , \zin[2][2] , \zin[2][1] , \zin[2][0] }), .zout({
        \zin[3][257] , \zin[3][256] , \zin[3][255] , \zin[3][254] , 
        \zin[3][253] , \zin[3][252] , \zin[3][251] , \zin[3][250] , 
        \zin[3][249] , \zin[3][248] , \zin[3][247] , \zin[3][246] , 
        \zin[3][245] , \zin[3][244] , \zin[3][243] , \zin[3][242] , 
        \zin[3][241] , \zin[3][240] , \zin[3][239] , \zin[3][238] , 
        \zin[3][237] , \zin[3][236] , \zin[3][235] , \zin[3][234] , 
        \zin[3][233] , \zin[3][232] , \zin[3][231] , \zin[3][230] , 
        \zin[3][229] , \zin[3][228] , \zin[3][227] , \zin[3][226] , 
        \zin[3][225] , \zin[3][224] , \zin[3][223] , \zin[3][222] , 
        \zin[3][221] , \zin[3][220] , \zin[3][219] , \zin[3][218] , 
        \zin[3][217] , \zin[3][216] , \zin[3][215] , \zin[3][214] , 
        \zin[3][213] , \zin[3][212] , \zin[3][211] , \zin[3][210] , 
        \zin[3][209] , \zin[3][208] , \zin[3][207] , \zin[3][206] , 
        \zin[3][205] , \zin[3][204] , \zin[3][203] , \zin[3][202] , 
        \zin[3][201] , \zin[3][200] , \zin[3][199] , \zin[3][198] , 
        \zin[3][197] , \zin[3][196] , \zin[3][195] , \zin[3][194] , 
        \zin[3][193] , \zin[3][192] , \zin[3][191] , \zin[3][190] , 
        \zin[3][189] , \zin[3][188] , \zin[3][187] , \zin[3][186] , 
        \zin[3][185] , \zin[3][184] , \zin[3][183] , \zin[3][182] , 
        \zin[3][181] , \zin[3][180] , \zin[3][179] , \zin[3][178] , 
        \zin[3][177] , \zin[3][176] , \zin[3][175] , \zin[3][174] , 
        \zin[3][173] , \zin[3][172] , \zin[3][171] , \zin[3][170] , 
        \zin[3][169] , \zin[3][168] , \zin[3][167] , \zin[3][166] , 
        \zin[3][165] , \zin[3][164] , \zin[3][163] , \zin[3][162] , 
        \zin[3][161] , \zin[3][160] , \zin[3][159] , \zin[3][158] , 
        \zin[3][157] , \zin[3][156] , \zin[3][155] , \zin[3][154] , 
        \zin[3][153] , \zin[3][152] , \zin[3][151] , \zin[3][150] , 
        \zin[3][149] , \zin[3][148] , \zin[3][147] , \zin[3][146] , 
        \zin[3][145] , \zin[3][144] , \zin[3][143] , \zin[3][142] , 
        \zin[3][141] , \zin[3][140] , \zin[3][139] , \zin[3][138] , 
        \zin[3][137] , \zin[3][136] , \zin[3][135] , \zin[3][134] , 
        \zin[3][133] , \zin[3][132] , \zin[3][131] , \zin[3][130] , 
        \zin[3][129] , \zin[3][128] , \zin[3][127] , \zin[3][126] , 
        \zin[3][125] , \zin[3][124] , \zin[3][123] , \zin[3][122] , 
        \zin[3][121] , \zin[3][120] , \zin[3][119] , \zin[3][118] , 
        \zin[3][117] , \zin[3][116] , \zin[3][115] , \zin[3][114] , 
        \zin[3][113] , \zin[3][112] , \zin[3][111] , \zin[3][110] , 
        \zin[3][109] , \zin[3][108] , \zin[3][107] , \zin[3][106] , 
        \zin[3][105] , \zin[3][104] , \zin[3][103] , \zin[3][102] , 
        \zin[3][101] , \zin[3][100] , \zin[3][99] , \zin[3][98] , \zin[3][97] , 
        \zin[3][96] , \zin[3][95] , \zin[3][94] , \zin[3][93] , \zin[3][92] , 
        \zin[3][91] , \zin[3][90] , \zin[3][89] , \zin[3][88] , \zin[3][87] , 
        \zin[3][86] , \zin[3][85] , \zin[3][84] , \zin[3][83] , \zin[3][82] , 
        \zin[3][81] , \zin[3][80] , \zin[3][79] , \zin[3][78] , \zin[3][77] , 
        \zin[3][76] , \zin[3][75] , \zin[3][74] , \zin[3][73] , \zin[3][72] , 
        \zin[3][71] , \zin[3][70] , \zin[3][69] , \zin[3][68] , \zin[3][67] , 
        \zin[3][66] , \zin[3][65] , \zin[3][64] , \zin[3][63] , \zin[3][62] , 
        \zin[3][61] , \zin[3][60] , \zin[3][59] , \zin[3][58] , \zin[3][57] , 
        \zin[3][56] , \zin[3][55] , \zin[3][54] , \zin[3][53] , \zin[3][52] , 
        \zin[3][51] , \zin[3][50] , \zin[3][49] , \zin[3][48] , \zin[3][47] , 
        \zin[3][46] , \zin[3][45] , \zin[3][44] , \zin[3][43] , \zin[3][42] , 
        \zin[3][41] , \zin[3][40] , \zin[3][39] , \zin[3][38] , \zin[3][37] , 
        \zin[3][36] , \zin[3][35] , \zin[3][34] , \zin[3][33] , \zin[3][32] , 
        \zin[3][31] , \zin[3][30] , \zin[3][29] , \zin[3][28] , \zin[3][27] , 
        \zin[3][26] , \zin[3][25] , \zin[3][24] , \zin[3][23] , \zin[3][22] , 
        \zin[3][21] , \zin[3][20] , \zin[3][19] , \zin[3][18] , \zin[3][17] , 
        \zin[3][16] , \zin[3][15] , \zin[3][14] , \zin[3][13] , \zin[3][12] , 
        \zin[3][11] , \zin[3][10] , \zin[3][9] , \zin[3][8] , \zin[3][7] , 
        \zin[3][6] , \zin[3][5] , \zin[3][4] , \zin[3][3] , \zin[3][2] , 
        \zin[3][1] , \zin[3][0] }) );
  modmult_step_N256_3 \MODMULT_STEP[3].modmult_step_  ( .xregN_1(xin[252]), 
        .y(y), .n(n), .zin({\zin[3][257] , \zin[3][256] , \zin[3][255] , 
        \zin[3][254] , \zin[3][253] , \zin[3][252] , \zin[3][251] , 
        \zin[3][250] , \zin[3][249] , \zin[3][248] , \zin[3][247] , 
        \zin[3][246] , \zin[3][245] , \zin[3][244] , \zin[3][243] , 
        \zin[3][242] , \zin[3][241] , \zin[3][240] , \zin[3][239] , 
        \zin[3][238] , \zin[3][237] , \zin[3][236] , \zin[3][235] , 
        \zin[3][234] , \zin[3][233] , \zin[3][232] , \zin[3][231] , 
        \zin[3][230] , \zin[3][229] , \zin[3][228] , \zin[3][227] , 
        \zin[3][226] , \zin[3][225] , \zin[3][224] , \zin[3][223] , 
        \zin[3][222] , \zin[3][221] , \zin[3][220] , \zin[3][219] , 
        \zin[3][218] , \zin[3][217] , \zin[3][216] , \zin[3][215] , 
        \zin[3][214] , \zin[3][213] , \zin[3][212] , \zin[3][211] , 
        \zin[3][210] , \zin[3][209] , \zin[3][208] , \zin[3][207] , 
        \zin[3][206] , \zin[3][205] , \zin[3][204] , \zin[3][203] , 
        \zin[3][202] , \zin[3][201] , \zin[3][200] , \zin[3][199] , 
        \zin[3][198] , \zin[3][197] , \zin[3][196] , \zin[3][195] , 
        \zin[3][194] , \zin[3][193] , \zin[3][192] , \zin[3][191] , 
        \zin[3][190] , \zin[3][189] , \zin[3][188] , \zin[3][187] , 
        \zin[3][186] , \zin[3][185] , \zin[3][184] , \zin[3][183] , 
        \zin[3][182] , \zin[3][181] , \zin[3][180] , \zin[3][179] , 
        \zin[3][178] , \zin[3][177] , \zin[3][176] , \zin[3][175] , 
        \zin[3][174] , \zin[3][173] , \zin[3][172] , \zin[3][171] , 
        \zin[3][170] , \zin[3][169] , \zin[3][168] , \zin[3][167] , 
        \zin[3][166] , \zin[3][165] , \zin[3][164] , \zin[3][163] , 
        \zin[3][162] , \zin[3][161] , \zin[3][160] , \zin[3][159] , 
        \zin[3][158] , \zin[3][157] , \zin[3][156] , \zin[3][155] , 
        \zin[3][154] , \zin[3][153] , \zin[3][152] , \zin[3][151] , 
        \zin[3][150] , \zin[3][149] , \zin[3][148] , \zin[3][147] , 
        \zin[3][146] , \zin[3][145] , \zin[3][144] , \zin[3][143] , 
        \zin[3][142] , \zin[3][141] , \zin[3][140] , \zin[3][139] , 
        \zin[3][138] , \zin[3][137] , \zin[3][136] , \zin[3][135] , 
        \zin[3][134] , \zin[3][133] , \zin[3][132] , \zin[3][131] , 
        \zin[3][130] , \zin[3][129] , \zin[3][128] , \zin[3][127] , 
        \zin[3][126] , \zin[3][125] , \zin[3][124] , \zin[3][123] , 
        \zin[3][122] , \zin[3][121] , \zin[3][120] , \zin[3][119] , 
        \zin[3][118] , \zin[3][117] , \zin[3][116] , \zin[3][115] , 
        \zin[3][114] , \zin[3][113] , \zin[3][112] , \zin[3][111] , 
        \zin[3][110] , \zin[3][109] , \zin[3][108] , \zin[3][107] , 
        \zin[3][106] , \zin[3][105] , \zin[3][104] , \zin[3][103] , 
        \zin[3][102] , \zin[3][101] , \zin[3][100] , \zin[3][99] , 
        \zin[3][98] , \zin[3][97] , \zin[3][96] , \zin[3][95] , \zin[3][94] , 
        \zin[3][93] , \zin[3][92] , \zin[3][91] , \zin[3][90] , \zin[3][89] , 
        \zin[3][88] , \zin[3][87] , \zin[3][86] , \zin[3][85] , \zin[3][84] , 
        \zin[3][83] , \zin[3][82] , \zin[3][81] , \zin[3][80] , \zin[3][79] , 
        \zin[3][78] , \zin[3][77] , \zin[3][76] , \zin[3][75] , \zin[3][74] , 
        \zin[3][73] , \zin[3][72] , \zin[3][71] , \zin[3][70] , \zin[3][69] , 
        \zin[3][68] , \zin[3][67] , \zin[3][66] , \zin[3][65] , \zin[3][64] , 
        \zin[3][63] , \zin[3][62] , \zin[3][61] , \zin[3][60] , \zin[3][59] , 
        \zin[3][58] , \zin[3][57] , \zin[3][56] , \zin[3][55] , \zin[3][54] , 
        \zin[3][53] , \zin[3][52] , \zin[3][51] , \zin[3][50] , \zin[3][49] , 
        \zin[3][48] , \zin[3][47] , \zin[3][46] , \zin[3][45] , \zin[3][44] , 
        \zin[3][43] , \zin[3][42] , \zin[3][41] , \zin[3][40] , \zin[3][39] , 
        \zin[3][38] , \zin[3][37] , \zin[3][36] , \zin[3][35] , \zin[3][34] , 
        \zin[3][33] , \zin[3][32] , \zin[3][31] , \zin[3][30] , \zin[3][29] , 
        \zin[3][28] , \zin[3][27] , \zin[3][26] , \zin[3][25] , \zin[3][24] , 
        \zin[3][23] , \zin[3][22] , \zin[3][21] , \zin[3][20] , \zin[3][19] , 
        \zin[3][18] , \zin[3][17] , \zin[3][16] , \zin[3][15] , \zin[3][14] , 
        \zin[3][13] , \zin[3][12] , \zin[3][11] , \zin[3][10] , \zin[3][9] , 
        \zin[3][8] , \zin[3][7] , \zin[3][6] , \zin[3][5] , \zin[3][4] , 
        \zin[3][3] , \zin[3][2] , \zin[3][1] , \zin[3][0] }), .zout({
        \zout[3][257] , \zout[3][256] , o}) );
  ANDN U3 ( .B(zreg[9]), .A(start), .Z(\zin[0][9] ) );
  ANDN U4 ( .B(zreg[99]), .A(start), .Z(\zin[0][99] ) );
  ANDN U5 ( .B(zreg[98]), .A(start), .Z(\zin[0][98] ) );
  ANDN U6 ( .B(zreg[97]), .A(start), .Z(\zin[0][97] ) );
  ANDN U7 ( .B(zreg[96]), .A(start), .Z(\zin[0][96] ) );
  ANDN U8 ( .B(zreg[95]), .A(start), .Z(\zin[0][95] ) );
  ANDN U9 ( .B(zreg[94]), .A(start), .Z(\zin[0][94] ) );
  ANDN U10 ( .B(zreg[93]), .A(start), .Z(\zin[0][93] ) );
  ANDN U11 ( .B(zreg[92]), .A(start), .Z(\zin[0][92] ) );
  ANDN U12 ( .B(zreg[91]), .A(start), .Z(\zin[0][91] ) );
  ANDN U13 ( .B(zreg[90]), .A(start), .Z(\zin[0][90] ) );
  ANDN U14 ( .B(zreg[8]), .A(start), .Z(\zin[0][8] ) );
  ANDN U15 ( .B(zreg[89]), .A(start), .Z(\zin[0][89] ) );
  ANDN U16 ( .B(zreg[88]), .A(start), .Z(\zin[0][88] ) );
  ANDN U17 ( .B(zreg[87]), .A(start), .Z(\zin[0][87] ) );
  ANDN U18 ( .B(zreg[86]), .A(start), .Z(\zin[0][86] ) );
  ANDN U19 ( .B(zreg[85]), .A(start), .Z(\zin[0][85] ) );
  ANDN U20 ( .B(zreg[84]), .A(start), .Z(\zin[0][84] ) );
  ANDN U21 ( .B(zreg[83]), .A(start), .Z(\zin[0][83] ) );
  ANDN U22 ( .B(zreg[82]), .A(start), .Z(\zin[0][82] ) );
  ANDN U23 ( .B(zreg[81]), .A(start), .Z(\zin[0][81] ) );
  ANDN U24 ( .B(zreg[80]), .A(start), .Z(\zin[0][80] ) );
  ANDN U25 ( .B(zreg[7]), .A(start), .Z(\zin[0][7] ) );
  ANDN U26 ( .B(zreg[79]), .A(start), .Z(\zin[0][79] ) );
  ANDN U27 ( .B(zreg[78]), .A(start), .Z(\zin[0][78] ) );
  ANDN U28 ( .B(zreg[77]), .A(start), .Z(\zin[0][77] ) );
  ANDN U29 ( .B(zreg[76]), .A(start), .Z(\zin[0][76] ) );
  ANDN U30 ( .B(zreg[75]), .A(start), .Z(\zin[0][75] ) );
  ANDN U31 ( .B(zreg[74]), .A(start), .Z(\zin[0][74] ) );
  ANDN U32 ( .B(zreg[73]), .A(start), .Z(\zin[0][73] ) );
  ANDN U33 ( .B(zreg[72]), .A(start), .Z(\zin[0][72] ) );
  ANDN U34 ( .B(zreg[71]), .A(start), .Z(\zin[0][71] ) );
  ANDN U35 ( .B(zreg[70]), .A(start), .Z(\zin[0][70] ) );
  ANDN U36 ( .B(zreg[6]), .A(start), .Z(\zin[0][6] ) );
  ANDN U37 ( .B(zreg[69]), .A(start), .Z(\zin[0][69] ) );
  ANDN U38 ( .B(zreg[68]), .A(start), .Z(\zin[0][68] ) );
  ANDN U39 ( .B(zreg[67]), .A(start), .Z(\zin[0][67] ) );
  ANDN U40 ( .B(zreg[66]), .A(start), .Z(\zin[0][66] ) );
  ANDN U41 ( .B(zreg[65]), .A(start), .Z(\zin[0][65] ) );
  ANDN U42 ( .B(zreg[64]), .A(start), .Z(\zin[0][64] ) );
  ANDN U43 ( .B(zreg[63]), .A(start), .Z(\zin[0][63] ) );
  ANDN U44 ( .B(zreg[62]), .A(start), .Z(\zin[0][62] ) );
  ANDN U45 ( .B(zreg[61]), .A(start), .Z(\zin[0][61] ) );
  ANDN U46 ( .B(zreg[60]), .A(start), .Z(\zin[0][60] ) );
  ANDN U47 ( .B(zreg[5]), .A(start), .Z(\zin[0][5] ) );
  ANDN U48 ( .B(zreg[59]), .A(start), .Z(\zin[0][59] ) );
  ANDN U49 ( .B(zreg[58]), .A(start), .Z(\zin[0][58] ) );
  ANDN U50 ( .B(zreg[57]), .A(start), .Z(\zin[0][57] ) );
  ANDN U51 ( .B(zreg[56]), .A(start), .Z(\zin[0][56] ) );
  ANDN U52 ( .B(zreg[55]), .A(start), .Z(\zin[0][55] ) );
  ANDN U53 ( .B(zreg[54]), .A(start), .Z(\zin[0][54] ) );
  ANDN U54 ( .B(zreg[53]), .A(start), .Z(\zin[0][53] ) );
  ANDN U55 ( .B(zreg[52]), .A(start), .Z(\zin[0][52] ) );
  ANDN U56 ( .B(zreg[51]), .A(start), .Z(\zin[0][51] ) );
  ANDN U57 ( .B(zreg[50]), .A(start), .Z(\zin[0][50] ) );
  ANDN U58 ( .B(zreg[4]), .A(start), .Z(\zin[0][4] ) );
  ANDN U59 ( .B(zreg[49]), .A(start), .Z(\zin[0][49] ) );
  ANDN U60 ( .B(zreg[48]), .A(start), .Z(\zin[0][48] ) );
  ANDN U61 ( .B(zreg[47]), .A(start), .Z(\zin[0][47] ) );
  ANDN U62 ( .B(zreg[46]), .A(start), .Z(\zin[0][46] ) );
  ANDN U63 ( .B(zreg[45]), .A(start), .Z(\zin[0][45] ) );
  ANDN U64 ( .B(zreg[44]), .A(start), .Z(\zin[0][44] ) );
  ANDN U65 ( .B(zreg[43]), .A(start), .Z(\zin[0][43] ) );
  ANDN U66 ( .B(zreg[42]), .A(start), .Z(\zin[0][42] ) );
  ANDN U67 ( .B(zreg[41]), .A(start), .Z(\zin[0][41] ) );
  ANDN U68 ( .B(zreg[40]), .A(start), .Z(\zin[0][40] ) );
  ANDN U69 ( .B(zreg[3]), .A(start), .Z(\zin[0][3] ) );
  ANDN U70 ( .B(zreg[39]), .A(start), .Z(\zin[0][39] ) );
  ANDN U71 ( .B(zreg[38]), .A(start), .Z(\zin[0][38] ) );
  ANDN U72 ( .B(zreg[37]), .A(start), .Z(\zin[0][37] ) );
  ANDN U73 ( .B(zreg[36]), .A(start), .Z(\zin[0][36] ) );
  ANDN U74 ( .B(zreg[35]), .A(start), .Z(\zin[0][35] ) );
  ANDN U75 ( .B(zreg[34]), .A(start), .Z(\zin[0][34] ) );
  ANDN U76 ( .B(zreg[33]), .A(start), .Z(\zin[0][33] ) );
  ANDN U77 ( .B(zreg[32]), .A(start), .Z(\zin[0][32] ) );
  ANDN U78 ( .B(zreg[31]), .A(start), .Z(\zin[0][31] ) );
  ANDN U79 ( .B(zreg[30]), .A(start), .Z(\zin[0][30] ) );
  ANDN U80 ( .B(zreg[2]), .A(start), .Z(\zin[0][2] ) );
  ANDN U81 ( .B(zreg[29]), .A(start), .Z(\zin[0][29] ) );
  ANDN U82 ( .B(zreg[28]), .A(start), .Z(\zin[0][28] ) );
  ANDN U83 ( .B(zreg[27]), .A(start), .Z(\zin[0][27] ) );
  ANDN U84 ( .B(zreg[26]), .A(start), .Z(\zin[0][26] ) );
  ANDN U85 ( .B(zreg[25]), .A(start), .Z(\zin[0][25] ) );
  ANDN U86 ( .B(zreg[257]), .A(start), .Z(\zin[0][257] ) );
  ANDN U87 ( .B(zreg[256]), .A(start), .Z(\zin[0][256] ) );
  ANDN U88 ( .B(zreg[255]), .A(start), .Z(\zin[0][255] ) );
  ANDN U89 ( .B(zreg[254]), .A(start), .Z(\zin[0][254] ) );
  ANDN U90 ( .B(zreg[253]), .A(start), .Z(\zin[0][253] ) );
  ANDN U91 ( .B(zreg[252]), .A(start), .Z(\zin[0][252] ) );
  ANDN U92 ( .B(zreg[251]), .A(start), .Z(\zin[0][251] ) );
  ANDN U93 ( .B(zreg[250]), .A(start), .Z(\zin[0][250] ) );
  ANDN U94 ( .B(zreg[24]), .A(start), .Z(\zin[0][24] ) );
  ANDN U95 ( .B(zreg[249]), .A(start), .Z(\zin[0][249] ) );
  ANDN U96 ( .B(zreg[248]), .A(start), .Z(\zin[0][248] ) );
  ANDN U97 ( .B(zreg[247]), .A(start), .Z(\zin[0][247] ) );
  ANDN U98 ( .B(zreg[246]), .A(start), .Z(\zin[0][246] ) );
  ANDN U99 ( .B(zreg[245]), .A(start), .Z(\zin[0][245] ) );
  ANDN U100 ( .B(zreg[244]), .A(start), .Z(\zin[0][244] ) );
  ANDN U101 ( .B(zreg[243]), .A(start), .Z(\zin[0][243] ) );
  ANDN U102 ( .B(zreg[242]), .A(start), .Z(\zin[0][242] ) );
  ANDN U103 ( .B(zreg[241]), .A(start), .Z(\zin[0][241] ) );
  ANDN U104 ( .B(zreg[240]), .A(start), .Z(\zin[0][240] ) );
  ANDN U105 ( .B(zreg[23]), .A(start), .Z(\zin[0][23] ) );
  ANDN U106 ( .B(zreg[239]), .A(start), .Z(\zin[0][239] ) );
  ANDN U107 ( .B(zreg[238]), .A(start), .Z(\zin[0][238] ) );
  ANDN U108 ( .B(zreg[237]), .A(start), .Z(\zin[0][237] ) );
  ANDN U109 ( .B(zreg[236]), .A(start), .Z(\zin[0][236] ) );
  ANDN U110 ( .B(zreg[235]), .A(start), .Z(\zin[0][235] ) );
  ANDN U111 ( .B(zreg[234]), .A(start), .Z(\zin[0][234] ) );
  ANDN U112 ( .B(zreg[233]), .A(start), .Z(\zin[0][233] ) );
  ANDN U113 ( .B(zreg[232]), .A(start), .Z(\zin[0][232] ) );
  ANDN U114 ( .B(zreg[231]), .A(start), .Z(\zin[0][231] ) );
  ANDN U115 ( .B(zreg[230]), .A(start), .Z(\zin[0][230] ) );
  ANDN U116 ( .B(zreg[22]), .A(start), .Z(\zin[0][22] ) );
  ANDN U117 ( .B(zreg[229]), .A(start), .Z(\zin[0][229] ) );
  ANDN U118 ( .B(zreg[228]), .A(start), .Z(\zin[0][228] ) );
  ANDN U119 ( .B(zreg[227]), .A(start), .Z(\zin[0][227] ) );
  ANDN U120 ( .B(zreg[226]), .A(start), .Z(\zin[0][226] ) );
  ANDN U121 ( .B(zreg[225]), .A(start), .Z(\zin[0][225] ) );
  ANDN U122 ( .B(zreg[224]), .A(start), .Z(\zin[0][224] ) );
  ANDN U123 ( .B(zreg[223]), .A(start), .Z(\zin[0][223] ) );
  ANDN U124 ( .B(zreg[222]), .A(start), .Z(\zin[0][222] ) );
  ANDN U125 ( .B(zreg[221]), .A(start), .Z(\zin[0][221] ) );
  ANDN U126 ( .B(zreg[220]), .A(start), .Z(\zin[0][220] ) );
  ANDN U127 ( .B(zreg[21]), .A(start), .Z(\zin[0][21] ) );
  ANDN U128 ( .B(zreg[219]), .A(start), .Z(\zin[0][219] ) );
  ANDN U129 ( .B(zreg[218]), .A(start), .Z(\zin[0][218] ) );
  ANDN U130 ( .B(zreg[217]), .A(start), .Z(\zin[0][217] ) );
  ANDN U131 ( .B(zreg[216]), .A(start), .Z(\zin[0][216] ) );
  ANDN U132 ( .B(zreg[215]), .A(start), .Z(\zin[0][215] ) );
  ANDN U133 ( .B(zreg[214]), .A(start), .Z(\zin[0][214] ) );
  ANDN U134 ( .B(zreg[213]), .A(start), .Z(\zin[0][213] ) );
  ANDN U135 ( .B(zreg[212]), .A(start), .Z(\zin[0][212] ) );
  ANDN U136 ( .B(zreg[211]), .A(start), .Z(\zin[0][211] ) );
  ANDN U137 ( .B(zreg[210]), .A(start), .Z(\zin[0][210] ) );
  ANDN U138 ( .B(zreg[20]), .A(start), .Z(\zin[0][20] ) );
  ANDN U139 ( .B(zreg[209]), .A(start), .Z(\zin[0][209] ) );
  ANDN U140 ( .B(zreg[208]), .A(start), .Z(\zin[0][208] ) );
  ANDN U141 ( .B(zreg[207]), .A(start), .Z(\zin[0][207] ) );
  ANDN U142 ( .B(zreg[206]), .A(start), .Z(\zin[0][206] ) );
  ANDN U143 ( .B(zreg[205]), .A(start), .Z(\zin[0][205] ) );
  ANDN U144 ( .B(zreg[204]), .A(start), .Z(\zin[0][204] ) );
  ANDN U145 ( .B(zreg[203]), .A(start), .Z(\zin[0][203] ) );
  ANDN U146 ( .B(zreg[202]), .A(start), .Z(\zin[0][202] ) );
  ANDN U147 ( .B(zreg[201]), .A(start), .Z(\zin[0][201] ) );
  ANDN U148 ( .B(zreg[200]), .A(start), .Z(\zin[0][200] ) );
  ANDN U149 ( .B(zreg[1]), .A(start), .Z(\zin[0][1] ) );
  ANDN U150 ( .B(zreg[19]), .A(start), .Z(\zin[0][19] ) );
  ANDN U151 ( .B(zreg[199]), .A(start), .Z(\zin[0][199] ) );
  ANDN U152 ( .B(zreg[198]), .A(start), .Z(\zin[0][198] ) );
  ANDN U153 ( .B(zreg[197]), .A(start), .Z(\zin[0][197] ) );
  ANDN U154 ( .B(zreg[196]), .A(start), .Z(\zin[0][196] ) );
  ANDN U155 ( .B(zreg[195]), .A(start), .Z(\zin[0][195] ) );
  ANDN U156 ( .B(zreg[194]), .A(start), .Z(\zin[0][194] ) );
  ANDN U157 ( .B(zreg[193]), .A(start), .Z(\zin[0][193] ) );
  ANDN U158 ( .B(zreg[192]), .A(start), .Z(\zin[0][192] ) );
  ANDN U159 ( .B(zreg[191]), .A(start), .Z(\zin[0][191] ) );
  ANDN U160 ( .B(zreg[190]), .A(start), .Z(\zin[0][190] ) );
  ANDN U161 ( .B(zreg[18]), .A(start), .Z(\zin[0][18] ) );
  ANDN U162 ( .B(zreg[189]), .A(start), .Z(\zin[0][189] ) );
  ANDN U163 ( .B(zreg[188]), .A(start), .Z(\zin[0][188] ) );
  ANDN U164 ( .B(zreg[187]), .A(start), .Z(\zin[0][187] ) );
  ANDN U165 ( .B(zreg[186]), .A(start), .Z(\zin[0][186] ) );
  ANDN U166 ( .B(zreg[185]), .A(start), .Z(\zin[0][185] ) );
  ANDN U167 ( .B(zreg[184]), .A(start), .Z(\zin[0][184] ) );
  ANDN U168 ( .B(zreg[183]), .A(start), .Z(\zin[0][183] ) );
  ANDN U169 ( .B(zreg[182]), .A(start), .Z(\zin[0][182] ) );
  ANDN U170 ( .B(zreg[181]), .A(start), .Z(\zin[0][181] ) );
  ANDN U171 ( .B(zreg[180]), .A(start), .Z(\zin[0][180] ) );
  ANDN U172 ( .B(zreg[17]), .A(start), .Z(\zin[0][17] ) );
  ANDN U173 ( .B(zreg[179]), .A(start), .Z(\zin[0][179] ) );
  ANDN U174 ( .B(zreg[178]), .A(start), .Z(\zin[0][178] ) );
  ANDN U175 ( .B(zreg[177]), .A(start), .Z(\zin[0][177] ) );
  ANDN U176 ( .B(zreg[176]), .A(start), .Z(\zin[0][176] ) );
  ANDN U177 ( .B(zreg[175]), .A(start), .Z(\zin[0][175] ) );
  ANDN U178 ( .B(zreg[174]), .A(start), .Z(\zin[0][174] ) );
  ANDN U179 ( .B(zreg[173]), .A(start), .Z(\zin[0][173] ) );
  ANDN U180 ( .B(zreg[172]), .A(start), .Z(\zin[0][172] ) );
  ANDN U181 ( .B(zreg[171]), .A(start), .Z(\zin[0][171] ) );
  ANDN U182 ( .B(zreg[170]), .A(start), .Z(\zin[0][170] ) );
  ANDN U183 ( .B(zreg[16]), .A(start), .Z(\zin[0][16] ) );
  ANDN U184 ( .B(zreg[169]), .A(start), .Z(\zin[0][169] ) );
  ANDN U185 ( .B(zreg[168]), .A(start), .Z(\zin[0][168] ) );
  ANDN U186 ( .B(zreg[167]), .A(start), .Z(\zin[0][167] ) );
  ANDN U187 ( .B(zreg[166]), .A(start), .Z(\zin[0][166] ) );
  ANDN U188 ( .B(zreg[165]), .A(start), .Z(\zin[0][165] ) );
  ANDN U189 ( .B(zreg[164]), .A(start), .Z(\zin[0][164] ) );
  ANDN U190 ( .B(zreg[163]), .A(start), .Z(\zin[0][163] ) );
  ANDN U191 ( .B(zreg[162]), .A(start), .Z(\zin[0][162] ) );
  ANDN U192 ( .B(zreg[161]), .A(start), .Z(\zin[0][161] ) );
  ANDN U193 ( .B(zreg[160]), .A(start), .Z(\zin[0][160] ) );
  ANDN U194 ( .B(zreg[15]), .A(start), .Z(\zin[0][15] ) );
  ANDN U195 ( .B(zreg[159]), .A(start), .Z(\zin[0][159] ) );
  ANDN U196 ( .B(zreg[158]), .A(start), .Z(\zin[0][158] ) );
  ANDN U197 ( .B(zreg[157]), .A(start), .Z(\zin[0][157] ) );
  ANDN U198 ( .B(zreg[156]), .A(start), .Z(\zin[0][156] ) );
  ANDN U199 ( .B(zreg[155]), .A(start), .Z(\zin[0][155] ) );
  ANDN U200 ( .B(zreg[154]), .A(start), .Z(\zin[0][154] ) );
  ANDN U201 ( .B(zreg[153]), .A(start), .Z(\zin[0][153] ) );
  ANDN U202 ( .B(zreg[152]), .A(start), .Z(\zin[0][152] ) );
  ANDN U203 ( .B(zreg[151]), .A(start), .Z(\zin[0][151] ) );
  ANDN U204 ( .B(zreg[150]), .A(start), .Z(\zin[0][150] ) );
  ANDN U205 ( .B(zreg[14]), .A(start), .Z(\zin[0][14] ) );
  ANDN U206 ( .B(zreg[149]), .A(start), .Z(\zin[0][149] ) );
  ANDN U207 ( .B(zreg[148]), .A(start), .Z(\zin[0][148] ) );
  ANDN U208 ( .B(zreg[147]), .A(start), .Z(\zin[0][147] ) );
  ANDN U209 ( .B(zreg[146]), .A(start), .Z(\zin[0][146] ) );
  ANDN U210 ( .B(zreg[145]), .A(start), .Z(\zin[0][145] ) );
  ANDN U211 ( .B(zreg[144]), .A(start), .Z(\zin[0][144] ) );
  ANDN U212 ( .B(zreg[143]), .A(start), .Z(\zin[0][143] ) );
  ANDN U213 ( .B(zreg[142]), .A(start), .Z(\zin[0][142] ) );
  ANDN U214 ( .B(zreg[141]), .A(start), .Z(\zin[0][141] ) );
  ANDN U215 ( .B(zreg[140]), .A(start), .Z(\zin[0][140] ) );
  ANDN U216 ( .B(zreg[13]), .A(start), .Z(\zin[0][13] ) );
  ANDN U217 ( .B(zreg[139]), .A(start), .Z(\zin[0][139] ) );
  ANDN U218 ( .B(zreg[138]), .A(start), .Z(\zin[0][138] ) );
  ANDN U219 ( .B(zreg[137]), .A(start), .Z(\zin[0][137] ) );
  ANDN U220 ( .B(zreg[136]), .A(start), .Z(\zin[0][136] ) );
  ANDN U221 ( .B(zreg[135]), .A(start), .Z(\zin[0][135] ) );
  ANDN U222 ( .B(zreg[134]), .A(start), .Z(\zin[0][134] ) );
  ANDN U223 ( .B(zreg[133]), .A(start), .Z(\zin[0][133] ) );
  ANDN U224 ( .B(zreg[132]), .A(start), .Z(\zin[0][132] ) );
  ANDN U225 ( .B(zreg[131]), .A(start), .Z(\zin[0][131] ) );
  ANDN U226 ( .B(zreg[130]), .A(start), .Z(\zin[0][130] ) );
  ANDN U227 ( .B(zreg[12]), .A(start), .Z(\zin[0][12] ) );
  ANDN U228 ( .B(zreg[129]), .A(start), .Z(\zin[0][129] ) );
  ANDN U229 ( .B(zreg[128]), .A(start), .Z(\zin[0][128] ) );
  ANDN U230 ( .B(zreg[127]), .A(start), .Z(\zin[0][127] ) );
  ANDN U231 ( .B(zreg[126]), .A(start), .Z(\zin[0][126] ) );
  ANDN U232 ( .B(zreg[125]), .A(start), .Z(\zin[0][125] ) );
  ANDN U233 ( .B(zreg[124]), .A(start), .Z(\zin[0][124] ) );
  ANDN U234 ( .B(zreg[123]), .A(start), .Z(\zin[0][123] ) );
  ANDN U235 ( .B(zreg[122]), .A(start), .Z(\zin[0][122] ) );
  ANDN U236 ( .B(zreg[121]), .A(start), .Z(\zin[0][121] ) );
  ANDN U237 ( .B(zreg[120]), .A(start), .Z(\zin[0][120] ) );
  ANDN U238 ( .B(zreg[11]), .A(start), .Z(\zin[0][11] ) );
  ANDN U239 ( .B(zreg[119]), .A(start), .Z(\zin[0][119] ) );
  ANDN U240 ( .B(zreg[118]), .A(start), .Z(\zin[0][118] ) );
  ANDN U241 ( .B(zreg[117]), .A(start), .Z(\zin[0][117] ) );
  ANDN U242 ( .B(zreg[116]), .A(start), .Z(\zin[0][116] ) );
  ANDN U243 ( .B(zreg[115]), .A(start), .Z(\zin[0][115] ) );
  ANDN U244 ( .B(zreg[114]), .A(start), .Z(\zin[0][114] ) );
  ANDN U245 ( .B(zreg[113]), .A(start), .Z(\zin[0][113] ) );
  ANDN U246 ( .B(zreg[112]), .A(start), .Z(\zin[0][112] ) );
  ANDN U247 ( .B(zreg[111]), .A(start), .Z(\zin[0][111] ) );
  ANDN U248 ( .B(zreg[110]), .A(start), .Z(\zin[0][110] ) );
  ANDN U249 ( .B(zreg[10]), .A(start), .Z(\zin[0][10] ) );
  ANDN U250 ( .B(zreg[109]), .A(start), .Z(\zin[0][109] ) );
  ANDN U251 ( .B(zreg[108]), .A(start), .Z(\zin[0][108] ) );
  ANDN U252 ( .B(zreg[107]), .A(start), .Z(\zin[0][107] ) );
  ANDN U253 ( .B(zreg[106]), .A(start), .Z(\zin[0][106] ) );
  ANDN U254 ( .B(zreg[105]), .A(start), .Z(\zin[0][105] ) );
  ANDN U255 ( .B(zreg[104]), .A(start), .Z(\zin[0][104] ) );
  ANDN U256 ( .B(zreg[103]), .A(start), .Z(\zin[0][103] ) );
  ANDN U257 ( .B(zreg[102]), .A(start), .Z(\zin[0][102] ) );
  ANDN U258 ( .B(zreg[101]), .A(start), .Z(\zin[0][101] ) );
  ANDN U259 ( .B(zreg[100]), .A(start), .Z(\zin[0][100] ) );
  ANDN U260 ( .B(zreg[0]), .A(start), .Z(\zin[0][0] ) );
  NAND U261 ( .A(n1), .B(n2), .Z(xin[9]) );
  NANDN U262 ( .A(start), .B(xreg[9]), .Z(n2) );
  NAND U263 ( .A(x[9]), .B(start), .Z(n1) );
  NAND U264 ( .A(n3), .B(n4), .Z(xin[99]) );
  NANDN U265 ( .A(start), .B(xreg[99]), .Z(n4) );
  NAND U266 ( .A(x[99]), .B(start), .Z(n3) );
  NAND U267 ( .A(n5), .B(n6), .Z(xin[98]) );
  NANDN U268 ( .A(start), .B(xreg[98]), .Z(n6) );
  NAND U269 ( .A(x[98]), .B(start), .Z(n5) );
  NAND U270 ( .A(n7), .B(n8), .Z(xin[97]) );
  NANDN U271 ( .A(start), .B(xreg[97]), .Z(n8) );
  NAND U272 ( .A(x[97]), .B(start), .Z(n7) );
  NAND U273 ( .A(n9), .B(n10), .Z(xin[96]) );
  NANDN U274 ( .A(start), .B(xreg[96]), .Z(n10) );
  NAND U275 ( .A(x[96]), .B(start), .Z(n9) );
  NAND U276 ( .A(n11), .B(n12), .Z(xin[95]) );
  NANDN U277 ( .A(start), .B(xreg[95]), .Z(n12) );
  NAND U278 ( .A(x[95]), .B(start), .Z(n11) );
  NAND U279 ( .A(n13), .B(n14), .Z(xin[94]) );
  NANDN U280 ( .A(start), .B(xreg[94]), .Z(n14) );
  NAND U281 ( .A(x[94]), .B(start), .Z(n13) );
  NAND U282 ( .A(n15), .B(n16), .Z(xin[93]) );
  NANDN U283 ( .A(start), .B(xreg[93]), .Z(n16) );
  NAND U284 ( .A(x[93]), .B(start), .Z(n15) );
  NAND U285 ( .A(n17), .B(n18), .Z(xin[92]) );
  NANDN U286 ( .A(start), .B(xreg[92]), .Z(n18) );
  NAND U287 ( .A(x[92]), .B(start), .Z(n17) );
  NAND U288 ( .A(n19), .B(n20), .Z(xin[91]) );
  NANDN U289 ( .A(start), .B(xreg[91]), .Z(n20) );
  NAND U290 ( .A(x[91]), .B(start), .Z(n19) );
  NAND U291 ( .A(n21), .B(n22), .Z(xin[90]) );
  NANDN U292 ( .A(start), .B(xreg[90]), .Z(n22) );
  NAND U293 ( .A(x[90]), .B(start), .Z(n21) );
  NAND U294 ( .A(n23), .B(n24), .Z(xin[8]) );
  NANDN U295 ( .A(start), .B(xreg[8]), .Z(n24) );
  NAND U296 ( .A(x[8]), .B(start), .Z(n23) );
  NAND U297 ( .A(n25), .B(n26), .Z(xin[89]) );
  NANDN U298 ( .A(start), .B(xreg[89]), .Z(n26) );
  NAND U299 ( .A(x[89]), .B(start), .Z(n25) );
  NAND U300 ( .A(n27), .B(n28), .Z(xin[88]) );
  NANDN U301 ( .A(start), .B(xreg[88]), .Z(n28) );
  NAND U302 ( .A(x[88]), .B(start), .Z(n27) );
  NAND U303 ( .A(n29), .B(n30), .Z(xin[87]) );
  NANDN U304 ( .A(start), .B(xreg[87]), .Z(n30) );
  NAND U305 ( .A(x[87]), .B(start), .Z(n29) );
  NAND U306 ( .A(n31), .B(n32), .Z(xin[86]) );
  NANDN U307 ( .A(start), .B(xreg[86]), .Z(n32) );
  NAND U308 ( .A(x[86]), .B(start), .Z(n31) );
  NAND U309 ( .A(n33), .B(n34), .Z(xin[85]) );
  NANDN U310 ( .A(start), .B(xreg[85]), .Z(n34) );
  NAND U311 ( .A(x[85]), .B(start), .Z(n33) );
  NAND U312 ( .A(n35), .B(n36), .Z(xin[84]) );
  NANDN U313 ( .A(start), .B(xreg[84]), .Z(n36) );
  NAND U314 ( .A(x[84]), .B(start), .Z(n35) );
  NAND U315 ( .A(n37), .B(n38), .Z(xin[83]) );
  NANDN U316 ( .A(start), .B(xreg[83]), .Z(n38) );
  NAND U317 ( .A(x[83]), .B(start), .Z(n37) );
  NAND U318 ( .A(n39), .B(n40), .Z(xin[82]) );
  NANDN U319 ( .A(start), .B(xreg[82]), .Z(n40) );
  NAND U320 ( .A(x[82]), .B(start), .Z(n39) );
  NAND U321 ( .A(n41), .B(n42), .Z(xin[81]) );
  NANDN U322 ( .A(start), .B(xreg[81]), .Z(n42) );
  NAND U323 ( .A(x[81]), .B(start), .Z(n41) );
  NAND U324 ( .A(n43), .B(n44), .Z(xin[80]) );
  NANDN U325 ( .A(start), .B(xreg[80]), .Z(n44) );
  NAND U326 ( .A(x[80]), .B(start), .Z(n43) );
  NAND U327 ( .A(n45), .B(n46), .Z(xin[7]) );
  NANDN U328 ( .A(start), .B(xreg[7]), .Z(n46) );
  NAND U329 ( .A(x[7]), .B(start), .Z(n45) );
  NAND U330 ( .A(n47), .B(n48), .Z(xin[79]) );
  NANDN U331 ( .A(start), .B(xreg[79]), .Z(n48) );
  NAND U332 ( .A(x[79]), .B(start), .Z(n47) );
  NAND U333 ( .A(n49), .B(n50), .Z(xin[78]) );
  NANDN U334 ( .A(start), .B(xreg[78]), .Z(n50) );
  NAND U335 ( .A(x[78]), .B(start), .Z(n49) );
  NAND U336 ( .A(n51), .B(n52), .Z(xin[77]) );
  NANDN U337 ( .A(start), .B(xreg[77]), .Z(n52) );
  NAND U338 ( .A(x[77]), .B(start), .Z(n51) );
  NAND U339 ( .A(n53), .B(n54), .Z(xin[76]) );
  NANDN U340 ( .A(start), .B(xreg[76]), .Z(n54) );
  NAND U341 ( .A(x[76]), .B(start), .Z(n53) );
  NAND U342 ( .A(n55), .B(n56), .Z(xin[75]) );
  NANDN U343 ( .A(start), .B(xreg[75]), .Z(n56) );
  NAND U344 ( .A(x[75]), .B(start), .Z(n55) );
  NAND U345 ( .A(n57), .B(n58), .Z(xin[74]) );
  NANDN U346 ( .A(start), .B(xreg[74]), .Z(n58) );
  NAND U347 ( .A(x[74]), .B(start), .Z(n57) );
  NAND U348 ( .A(n59), .B(n60), .Z(xin[73]) );
  NANDN U349 ( .A(start), .B(xreg[73]), .Z(n60) );
  NAND U350 ( .A(x[73]), .B(start), .Z(n59) );
  NAND U351 ( .A(n61), .B(n62), .Z(xin[72]) );
  NANDN U352 ( .A(start), .B(xreg[72]), .Z(n62) );
  NAND U353 ( .A(x[72]), .B(start), .Z(n61) );
  NAND U354 ( .A(n63), .B(n64), .Z(xin[71]) );
  NANDN U355 ( .A(start), .B(xreg[71]), .Z(n64) );
  NAND U356 ( .A(x[71]), .B(start), .Z(n63) );
  NAND U357 ( .A(n65), .B(n66), .Z(xin[70]) );
  NANDN U358 ( .A(start), .B(xreg[70]), .Z(n66) );
  NAND U359 ( .A(x[70]), .B(start), .Z(n65) );
  NAND U360 ( .A(n67), .B(n68), .Z(xin[6]) );
  NANDN U361 ( .A(start), .B(xreg[6]), .Z(n68) );
  NAND U362 ( .A(x[6]), .B(start), .Z(n67) );
  NAND U363 ( .A(n69), .B(n70), .Z(xin[69]) );
  NANDN U364 ( .A(start), .B(xreg[69]), .Z(n70) );
  NAND U365 ( .A(x[69]), .B(start), .Z(n69) );
  NAND U366 ( .A(n71), .B(n72), .Z(xin[68]) );
  NANDN U367 ( .A(start), .B(xreg[68]), .Z(n72) );
  NAND U368 ( .A(x[68]), .B(start), .Z(n71) );
  NAND U369 ( .A(n73), .B(n74), .Z(xin[67]) );
  NANDN U370 ( .A(start), .B(xreg[67]), .Z(n74) );
  NAND U371 ( .A(x[67]), .B(start), .Z(n73) );
  NAND U372 ( .A(n75), .B(n76), .Z(xin[66]) );
  NANDN U373 ( .A(start), .B(xreg[66]), .Z(n76) );
  NAND U374 ( .A(x[66]), .B(start), .Z(n75) );
  NAND U375 ( .A(n77), .B(n78), .Z(xin[65]) );
  NANDN U376 ( .A(start), .B(xreg[65]), .Z(n78) );
  NAND U377 ( .A(x[65]), .B(start), .Z(n77) );
  NAND U378 ( .A(n79), .B(n80), .Z(xin[64]) );
  NANDN U379 ( .A(start), .B(xreg[64]), .Z(n80) );
  NAND U380 ( .A(x[64]), .B(start), .Z(n79) );
  NAND U381 ( .A(n81), .B(n82), .Z(xin[63]) );
  NANDN U382 ( .A(start), .B(xreg[63]), .Z(n82) );
  NAND U383 ( .A(x[63]), .B(start), .Z(n81) );
  NAND U384 ( .A(n83), .B(n84), .Z(xin[62]) );
  NANDN U385 ( .A(start), .B(xreg[62]), .Z(n84) );
  NAND U386 ( .A(x[62]), .B(start), .Z(n83) );
  NAND U387 ( .A(n85), .B(n86), .Z(xin[61]) );
  NANDN U388 ( .A(start), .B(xreg[61]), .Z(n86) );
  NAND U389 ( .A(x[61]), .B(start), .Z(n85) );
  NAND U390 ( .A(n87), .B(n88), .Z(xin[60]) );
  NANDN U391 ( .A(start), .B(xreg[60]), .Z(n88) );
  NAND U392 ( .A(x[60]), .B(start), .Z(n87) );
  NAND U393 ( .A(n89), .B(n90), .Z(xin[5]) );
  NANDN U394 ( .A(start), .B(xreg[5]), .Z(n90) );
  NAND U395 ( .A(x[5]), .B(start), .Z(n89) );
  NAND U396 ( .A(n91), .B(n92), .Z(xin[59]) );
  NANDN U397 ( .A(start), .B(xreg[59]), .Z(n92) );
  NAND U398 ( .A(x[59]), .B(start), .Z(n91) );
  NAND U399 ( .A(n93), .B(n94), .Z(xin[58]) );
  NANDN U400 ( .A(start), .B(xreg[58]), .Z(n94) );
  NAND U401 ( .A(x[58]), .B(start), .Z(n93) );
  NAND U402 ( .A(n95), .B(n96), .Z(xin[57]) );
  NANDN U403 ( .A(start), .B(xreg[57]), .Z(n96) );
  NAND U404 ( .A(x[57]), .B(start), .Z(n95) );
  NAND U405 ( .A(n97), .B(n98), .Z(xin[56]) );
  NANDN U406 ( .A(start), .B(xreg[56]), .Z(n98) );
  NAND U407 ( .A(x[56]), .B(start), .Z(n97) );
  NAND U408 ( .A(n99), .B(n100), .Z(xin[55]) );
  NANDN U409 ( .A(start), .B(xreg[55]), .Z(n100) );
  NAND U410 ( .A(x[55]), .B(start), .Z(n99) );
  NAND U411 ( .A(n101), .B(n102), .Z(xin[54]) );
  NANDN U412 ( .A(start), .B(xreg[54]), .Z(n102) );
  NAND U413 ( .A(x[54]), .B(start), .Z(n101) );
  NAND U414 ( .A(n103), .B(n104), .Z(xin[53]) );
  NANDN U415 ( .A(start), .B(xreg[53]), .Z(n104) );
  NAND U416 ( .A(x[53]), .B(start), .Z(n103) );
  NAND U417 ( .A(n105), .B(n106), .Z(xin[52]) );
  NANDN U418 ( .A(start), .B(xreg[52]), .Z(n106) );
  NAND U419 ( .A(x[52]), .B(start), .Z(n105) );
  NAND U420 ( .A(n107), .B(n108), .Z(xin[51]) );
  NANDN U421 ( .A(start), .B(xreg[51]), .Z(n108) );
  NAND U422 ( .A(x[51]), .B(start), .Z(n107) );
  NAND U423 ( .A(n109), .B(n110), .Z(xin[50]) );
  NANDN U424 ( .A(start), .B(xreg[50]), .Z(n110) );
  NAND U425 ( .A(x[50]), .B(start), .Z(n109) );
  NAND U426 ( .A(n111), .B(n112), .Z(xin[4]) );
  NANDN U427 ( .A(start), .B(xreg[4]), .Z(n112) );
  NAND U428 ( .A(x[4]), .B(start), .Z(n111) );
  NAND U429 ( .A(n113), .B(n114), .Z(xin[49]) );
  NANDN U430 ( .A(start), .B(xreg[49]), .Z(n114) );
  NAND U431 ( .A(x[49]), .B(start), .Z(n113) );
  NAND U432 ( .A(n115), .B(n116), .Z(xin[48]) );
  NANDN U433 ( .A(start), .B(xreg[48]), .Z(n116) );
  NAND U434 ( .A(x[48]), .B(start), .Z(n115) );
  NAND U435 ( .A(n117), .B(n118), .Z(xin[47]) );
  NANDN U436 ( .A(start), .B(xreg[47]), .Z(n118) );
  NAND U437 ( .A(x[47]), .B(start), .Z(n117) );
  NAND U438 ( .A(n119), .B(n120), .Z(xin[46]) );
  NANDN U439 ( .A(start), .B(xreg[46]), .Z(n120) );
  NAND U440 ( .A(x[46]), .B(start), .Z(n119) );
  NAND U441 ( .A(n121), .B(n122), .Z(xin[45]) );
  NANDN U442 ( .A(start), .B(xreg[45]), .Z(n122) );
  NAND U443 ( .A(x[45]), .B(start), .Z(n121) );
  NAND U444 ( .A(n123), .B(n124), .Z(xin[44]) );
  NANDN U445 ( .A(start), .B(xreg[44]), .Z(n124) );
  NAND U446 ( .A(x[44]), .B(start), .Z(n123) );
  NAND U447 ( .A(n125), .B(n126), .Z(xin[43]) );
  NANDN U448 ( .A(start), .B(xreg[43]), .Z(n126) );
  NAND U449 ( .A(x[43]), .B(start), .Z(n125) );
  NAND U450 ( .A(n127), .B(n128), .Z(xin[42]) );
  NANDN U451 ( .A(start), .B(xreg[42]), .Z(n128) );
  NAND U452 ( .A(x[42]), .B(start), .Z(n127) );
  NAND U453 ( .A(n129), .B(n130), .Z(xin[41]) );
  NANDN U454 ( .A(start), .B(xreg[41]), .Z(n130) );
  NAND U455 ( .A(x[41]), .B(start), .Z(n129) );
  NAND U456 ( .A(n131), .B(n132), .Z(xin[40]) );
  NANDN U457 ( .A(start), .B(xreg[40]), .Z(n132) );
  NAND U458 ( .A(x[40]), .B(start), .Z(n131) );
  NAND U459 ( .A(n133), .B(n134), .Z(xin[39]) );
  NANDN U460 ( .A(start), .B(xreg[39]), .Z(n134) );
  NAND U461 ( .A(x[39]), .B(start), .Z(n133) );
  NAND U462 ( .A(n135), .B(n136), .Z(xin[38]) );
  NANDN U463 ( .A(start), .B(xreg[38]), .Z(n136) );
  NAND U464 ( .A(x[38]), .B(start), .Z(n135) );
  NAND U465 ( .A(n137), .B(n138), .Z(xin[37]) );
  NANDN U466 ( .A(start), .B(xreg[37]), .Z(n138) );
  NAND U467 ( .A(x[37]), .B(start), .Z(n137) );
  NAND U468 ( .A(n139), .B(n140), .Z(xin[36]) );
  NANDN U469 ( .A(start), .B(xreg[36]), .Z(n140) );
  NAND U470 ( .A(x[36]), .B(start), .Z(n139) );
  NAND U471 ( .A(n141), .B(n142), .Z(xin[35]) );
  NANDN U472 ( .A(start), .B(xreg[35]), .Z(n142) );
  NAND U473 ( .A(x[35]), .B(start), .Z(n141) );
  NAND U474 ( .A(n143), .B(n144), .Z(xin[34]) );
  NANDN U475 ( .A(start), .B(xreg[34]), .Z(n144) );
  NAND U476 ( .A(x[34]), .B(start), .Z(n143) );
  NAND U477 ( .A(n145), .B(n146), .Z(xin[33]) );
  NANDN U478 ( .A(start), .B(xreg[33]), .Z(n146) );
  NAND U479 ( .A(x[33]), .B(start), .Z(n145) );
  NAND U480 ( .A(n147), .B(n148), .Z(xin[32]) );
  NANDN U481 ( .A(start), .B(xreg[32]), .Z(n148) );
  NAND U482 ( .A(x[32]), .B(start), .Z(n147) );
  NAND U483 ( .A(n149), .B(n150), .Z(xin[31]) );
  NANDN U484 ( .A(start), .B(xreg[31]), .Z(n150) );
  NAND U485 ( .A(x[31]), .B(start), .Z(n149) );
  NAND U486 ( .A(n151), .B(n152), .Z(xin[30]) );
  NANDN U487 ( .A(start), .B(xreg[30]), .Z(n152) );
  NAND U488 ( .A(x[30]), .B(start), .Z(n151) );
  NAND U489 ( .A(n153), .B(n154), .Z(xin[29]) );
  NANDN U490 ( .A(start), .B(xreg[29]), .Z(n154) );
  NAND U491 ( .A(x[29]), .B(start), .Z(n153) );
  NAND U492 ( .A(n155), .B(n156), .Z(xin[28]) );
  NANDN U493 ( .A(start), .B(xreg[28]), .Z(n156) );
  NAND U494 ( .A(x[28]), .B(start), .Z(n155) );
  NAND U495 ( .A(n157), .B(n158), .Z(xin[27]) );
  NANDN U496 ( .A(start), .B(xreg[27]), .Z(n158) );
  NAND U497 ( .A(x[27]), .B(start), .Z(n157) );
  NAND U498 ( .A(n159), .B(n160), .Z(xin[26]) );
  NANDN U499 ( .A(start), .B(xreg[26]), .Z(n160) );
  NAND U500 ( .A(x[26]), .B(start), .Z(n159) );
  NAND U501 ( .A(n161), .B(n162), .Z(xin[25]) );
  NANDN U502 ( .A(start), .B(xreg[25]), .Z(n162) );
  NAND U503 ( .A(x[25]), .B(start), .Z(n161) );
  NAND U504 ( .A(n163), .B(n164), .Z(xin[255]) );
  NANDN U505 ( .A(start), .B(xreg[255]), .Z(n164) );
  NAND U506 ( .A(x[255]), .B(start), .Z(n163) );
  NAND U507 ( .A(n165), .B(n166), .Z(xin[254]) );
  NANDN U508 ( .A(start), .B(xreg[254]), .Z(n166) );
  NAND U509 ( .A(x[254]), .B(start), .Z(n165) );
  NAND U510 ( .A(n167), .B(n168), .Z(xin[253]) );
  NANDN U511 ( .A(start), .B(xreg[253]), .Z(n168) );
  NAND U512 ( .A(x[253]), .B(start), .Z(n167) );
  NAND U513 ( .A(n169), .B(n170), .Z(xin[252]) );
  NANDN U514 ( .A(start), .B(xreg[252]), .Z(n170) );
  NAND U515 ( .A(x[252]), .B(start), .Z(n169) );
  NAND U516 ( .A(n171), .B(n172), .Z(xin[251]) );
  NANDN U517 ( .A(start), .B(xreg[251]), .Z(n172) );
  NAND U518 ( .A(x[251]), .B(start), .Z(n171) );
  NAND U519 ( .A(n173), .B(n174), .Z(xin[250]) );
  NANDN U520 ( .A(start), .B(xreg[250]), .Z(n174) );
  NAND U521 ( .A(x[250]), .B(start), .Z(n173) );
  NAND U522 ( .A(n175), .B(n176), .Z(xin[24]) );
  NANDN U523 ( .A(start), .B(xreg[24]), .Z(n176) );
  NAND U524 ( .A(x[24]), .B(start), .Z(n175) );
  NAND U525 ( .A(n177), .B(n178), .Z(xin[249]) );
  NANDN U526 ( .A(start), .B(xreg[249]), .Z(n178) );
  NAND U527 ( .A(x[249]), .B(start), .Z(n177) );
  NAND U528 ( .A(n179), .B(n180), .Z(xin[248]) );
  NANDN U529 ( .A(start), .B(xreg[248]), .Z(n180) );
  NAND U530 ( .A(x[248]), .B(start), .Z(n179) );
  NAND U531 ( .A(n181), .B(n182), .Z(xin[247]) );
  NANDN U532 ( .A(start), .B(xreg[247]), .Z(n182) );
  NAND U533 ( .A(x[247]), .B(start), .Z(n181) );
  NAND U534 ( .A(n183), .B(n184), .Z(xin[246]) );
  NANDN U535 ( .A(start), .B(xreg[246]), .Z(n184) );
  NAND U536 ( .A(x[246]), .B(start), .Z(n183) );
  NAND U537 ( .A(n185), .B(n186), .Z(xin[245]) );
  NANDN U538 ( .A(start), .B(xreg[245]), .Z(n186) );
  NAND U539 ( .A(x[245]), .B(start), .Z(n185) );
  NAND U540 ( .A(n187), .B(n188), .Z(xin[244]) );
  NANDN U541 ( .A(start), .B(xreg[244]), .Z(n188) );
  NAND U542 ( .A(x[244]), .B(start), .Z(n187) );
  NAND U543 ( .A(n189), .B(n190), .Z(xin[243]) );
  NANDN U544 ( .A(start), .B(xreg[243]), .Z(n190) );
  NAND U545 ( .A(x[243]), .B(start), .Z(n189) );
  NAND U546 ( .A(n191), .B(n192), .Z(xin[242]) );
  NANDN U547 ( .A(start), .B(xreg[242]), .Z(n192) );
  NAND U548 ( .A(x[242]), .B(start), .Z(n191) );
  NAND U549 ( .A(n193), .B(n194), .Z(xin[241]) );
  NANDN U550 ( .A(start), .B(xreg[241]), .Z(n194) );
  NAND U551 ( .A(x[241]), .B(start), .Z(n193) );
  NAND U552 ( .A(n195), .B(n196), .Z(xin[240]) );
  NANDN U553 ( .A(start), .B(xreg[240]), .Z(n196) );
  NAND U554 ( .A(x[240]), .B(start), .Z(n195) );
  NAND U555 ( .A(n197), .B(n198), .Z(xin[23]) );
  NANDN U556 ( .A(start), .B(xreg[23]), .Z(n198) );
  NAND U557 ( .A(x[23]), .B(start), .Z(n197) );
  NAND U558 ( .A(n199), .B(n200), .Z(xin[239]) );
  NANDN U559 ( .A(start), .B(xreg[239]), .Z(n200) );
  NAND U560 ( .A(x[239]), .B(start), .Z(n199) );
  NAND U561 ( .A(n201), .B(n202), .Z(xin[238]) );
  NANDN U562 ( .A(start), .B(xreg[238]), .Z(n202) );
  NAND U563 ( .A(x[238]), .B(start), .Z(n201) );
  NAND U564 ( .A(n203), .B(n204), .Z(xin[237]) );
  NANDN U565 ( .A(start), .B(xreg[237]), .Z(n204) );
  NAND U566 ( .A(x[237]), .B(start), .Z(n203) );
  NAND U567 ( .A(n205), .B(n206), .Z(xin[236]) );
  NANDN U568 ( .A(start), .B(xreg[236]), .Z(n206) );
  NAND U569 ( .A(x[236]), .B(start), .Z(n205) );
  NAND U570 ( .A(n207), .B(n208), .Z(xin[235]) );
  NANDN U571 ( .A(start), .B(xreg[235]), .Z(n208) );
  NAND U572 ( .A(x[235]), .B(start), .Z(n207) );
  NAND U573 ( .A(n209), .B(n210), .Z(xin[234]) );
  NANDN U574 ( .A(start), .B(xreg[234]), .Z(n210) );
  NAND U575 ( .A(x[234]), .B(start), .Z(n209) );
  NAND U576 ( .A(n211), .B(n212), .Z(xin[233]) );
  NANDN U577 ( .A(start), .B(xreg[233]), .Z(n212) );
  NAND U578 ( .A(x[233]), .B(start), .Z(n211) );
  NAND U579 ( .A(n213), .B(n214), .Z(xin[232]) );
  NANDN U580 ( .A(start), .B(xreg[232]), .Z(n214) );
  NAND U581 ( .A(x[232]), .B(start), .Z(n213) );
  NAND U582 ( .A(n215), .B(n216), .Z(xin[231]) );
  NANDN U583 ( .A(start), .B(xreg[231]), .Z(n216) );
  NAND U584 ( .A(x[231]), .B(start), .Z(n215) );
  NAND U585 ( .A(n217), .B(n218), .Z(xin[230]) );
  NANDN U586 ( .A(start), .B(xreg[230]), .Z(n218) );
  NAND U587 ( .A(x[230]), .B(start), .Z(n217) );
  NAND U588 ( .A(n219), .B(n220), .Z(xin[22]) );
  NANDN U589 ( .A(start), .B(xreg[22]), .Z(n220) );
  NAND U590 ( .A(x[22]), .B(start), .Z(n219) );
  NAND U591 ( .A(n221), .B(n222), .Z(xin[229]) );
  NANDN U592 ( .A(start), .B(xreg[229]), .Z(n222) );
  NAND U593 ( .A(x[229]), .B(start), .Z(n221) );
  NAND U594 ( .A(n223), .B(n224), .Z(xin[228]) );
  NANDN U595 ( .A(start), .B(xreg[228]), .Z(n224) );
  NAND U596 ( .A(x[228]), .B(start), .Z(n223) );
  NAND U597 ( .A(n225), .B(n226), .Z(xin[227]) );
  NANDN U598 ( .A(start), .B(xreg[227]), .Z(n226) );
  NAND U599 ( .A(x[227]), .B(start), .Z(n225) );
  NAND U600 ( .A(n227), .B(n228), .Z(xin[226]) );
  NANDN U601 ( .A(start), .B(xreg[226]), .Z(n228) );
  NAND U602 ( .A(x[226]), .B(start), .Z(n227) );
  NAND U603 ( .A(n229), .B(n230), .Z(xin[225]) );
  NANDN U604 ( .A(start), .B(xreg[225]), .Z(n230) );
  NAND U605 ( .A(x[225]), .B(start), .Z(n229) );
  NAND U606 ( .A(n231), .B(n232), .Z(xin[224]) );
  NANDN U607 ( .A(start), .B(xreg[224]), .Z(n232) );
  NAND U608 ( .A(x[224]), .B(start), .Z(n231) );
  NAND U609 ( .A(n233), .B(n234), .Z(xin[223]) );
  NANDN U610 ( .A(start), .B(xreg[223]), .Z(n234) );
  NAND U611 ( .A(x[223]), .B(start), .Z(n233) );
  NAND U612 ( .A(n235), .B(n236), .Z(xin[222]) );
  NANDN U613 ( .A(start), .B(xreg[222]), .Z(n236) );
  NAND U614 ( .A(x[222]), .B(start), .Z(n235) );
  NAND U615 ( .A(n237), .B(n238), .Z(xin[221]) );
  NANDN U616 ( .A(start), .B(xreg[221]), .Z(n238) );
  NAND U617 ( .A(x[221]), .B(start), .Z(n237) );
  NAND U618 ( .A(n239), .B(n240), .Z(xin[220]) );
  NANDN U619 ( .A(start), .B(xreg[220]), .Z(n240) );
  NAND U620 ( .A(x[220]), .B(start), .Z(n239) );
  NAND U621 ( .A(n241), .B(n242), .Z(xin[21]) );
  NANDN U622 ( .A(start), .B(xreg[21]), .Z(n242) );
  NAND U623 ( .A(x[21]), .B(start), .Z(n241) );
  NAND U624 ( .A(n243), .B(n244), .Z(xin[219]) );
  NANDN U625 ( .A(start), .B(xreg[219]), .Z(n244) );
  NAND U626 ( .A(x[219]), .B(start), .Z(n243) );
  NAND U627 ( .A(n245), .B(n246), .Z(xin[218]) );
  NANDN U628 ( .A(start), .B(xreg[218]), .Z(n246) );
  NAND U629 ( .A(x[218]), .B(start), .Z(n245) );
  NAND U630 ( .A(n247), .B(n248), .Z(xin[217]) );
  NANDN U631 ( .A(start), .B(xreg[217]), .Z(n248) );
  NAND U632 ( .A(x[217]), .B(start), .Z(n247) );
  NAND U633 ( .A(n249), .B(n250), .Z(xin[216]) );
  NANDN U634 ( .A(start), .B(xreg[216]), .Z(n250) );
  NAND U635 ( .A(x[216]), .B(start), .Z(n249) );
  NAND U636 ( .A(n251), .B(n252), .Z(xin[215]) );
  NANDN U637 ( .A(start), .B(xreg[215]), .Z(n252) );
  NAND U638 ( .A(x[215]), .B(start), .Z(n251) );
  NAND U639 ( .A(n253), .B(n254), .Z(xin[214]) );
  NANDN U640 ( .A(start), .B(xreg[214]), .Z(n254) );
  NAND U641 ( .A(x[214]), .B(start), .Z(n253) );
  NAND U642 ( .A(n255), .B(n256), .Z(xin[213]) );
  NANDN U643 ( .A(start), .B(xreg[213]), .Z(n256) );
  NAND U644 ( .A(x[213]), .B(start), .Z(n255) );
  NAND U645 ( .A(n257), .B(n258), .Z(xin[212]) );
  NANDN U646 ( .A(start), .B(xreg[212]), .Z(n258) );
  NAND U647 ( .A(x[212]), .B(start), .Z(n257) );
  NAND U648 ( .A(n259), .B(n260), .Z(xin[211]) );
  NANDN U649 ( .A(start), .B(xreg[211]), .Z(n260) );
  NAND U650 ( .A(x[211]), .B(start), .Z(n259) );
  NAND U651 ( .A(n261), .B(n262), .Z(xin[210]) );
  NANDN U652 ( .A(start), .B(xreg[210]), .Z(n262) );
  NAND U653 ( .A(x[210]), .B(start), .Z(n261) );
  NAND U654 ( .A(n263), .B(n264), .Z(xin[20]) );
  NANDN U655 ( .A(start), .B(xreg[20]), .Z(n264) );
  NAND U656 ( .A(x[20]), .B(start), .Z(n263) );
  NAND U657 ( .A(n265), .B(n266), .Z(xin[209]) );
  NANDN U658 ( .A(start), .B(xreg[209]), .Z(n266) );
  NAND U659 ( .A(x[209]), .B(start), .Z(n265) );
  NAND U660 ( .A(n267), .B(n268), .Z(xin[208]) );
  NANDN U661 ( .A(start), .B(xreg[208]), .Z(n268) );
  NAND U662 ( .A(x[208]), .B(start), .Z(n267) );
  NAND U663 ( .A(n269), .B(n270), .Z(xin[207]) );
  NANDN U664 ( .A(start), .B(xreg[207]), .Z(n270) );
  NAND U665 ( .A(x[207]), .B(start), .Z(n269) );
  NAND U666 ( .A(n271), .B(n272), .Z(xin[206]) );
  NANDN U667 ( .A(start), .B(xreg[206]), .Z(n272) );
  NAND U668 ( .A(x[206]), .B(start), .Z(n271) );
  NAND U669 ( .A(n273), .B(n274), .Z(xin[205]) );
  NANDN U670 ( .A(start), .B(xreg[205]), .Z(n274) );
  NAND U671 ( .A(x[205]), .B(start), .Z(n273) );
  NAND U672 ( .A(n275), .B(n276), .Z(xin[204]) );
  NANDN U673 ( .A(start), .B(xreg[204]), .Z(n276) );
  NAND U674 ( .A(x[204]), .B(start), .Z(n275) );
  NAND U675 ( .A(n277), .B(n278), .Z(xin[203]) );
  NANDN U676 ( .A(start), .B(xreg[203]), .Z(n278) );
  NAND U677 ( .A(x[203]), .B(start), .Z(n277) );
  NAND U678 ( .A(n279), .B(n280), .Z(xin[202]) );
  NANDN U679 ( .A(start), .B(xreg[202]), .Z(n280) );
  NAND U680 ( .A(x[202]), .B(start), .Z(n279) );
  NAND U681 ( .A(n281), .B(n282), .Z(xin[201]) );
  NANDN U682 ( .A(start), .B(xreg[201]), .Z(n282) );
  NAND U683 ( .A(x[201]), .B(start), .Z(n281) );
  NAND U684 ( .A(n283), .B(n284), .Z(xin[200]) );
  NANDN U685 ( .A(start), .B(xreg[200]), .Z(n284) );
  NAND U686 ( .A(x[200]), .B(start), .Z(n283) );
  NAND U687 ( .A(n285), .B(n286), .Z(xin[19]) );
  NANDN U688 ( .A(start), .B(xreg[19]), .Z(n286) );
  NAND U689 ( .A(x[19]), .B(start), .Z(n285) );
  NAND U690 ( .A(n287), .B(n288), .Z(xin[199]) );
  NANDN U691 ( .A(start), .B(xreg[199]), .Z(n288) );
  NAND U692 ( .A(x[199]), .B(start), .Z(n287) );
  NAND U693 ( .A(n289), .B(n290), .Z(xin[198]) );
  NANDN U694 ( .A(start), .B(xreg[198]), .Z(n290) );
  NAND U695 ( .A(x[198]), .B(start), .Z(n289) );
  NAND U696 ( .A(n291), .B(n292), .Z(xin[197]) );
  NANDN U697 ( .A(start), .B(xreg[197]), .Z(n292) );
  NAND U698 ( .A(x[197]), .B(start), .Z(n291) );
  NAND U699 ( .A(n293), .B(n294), .Z(xin[196]) );
  NANDN U700 ( .A(start), .B(xreg[196]), .Z(n294) );
  NAND U701 ( .A(x[196]), .B(start), .Z(n293) );
  NAND U702 ( .A(n295), .B(n296), .Z(xin[195]) );
  NANDN U703 ( .A(start), .B(xreg[195]), .Z(n296) );
  NAND U704 ( .A(x[195]), .B(start), .Z(n295) );
  NAND U705 ( .A(n297), .B(n298), .Z(xin[194]) );
  NANDN U706 ( .A(start), .B(xreg[194]), .Z(n298) );
  NAND U707 ( .A(x[194]), .B(start), .Z(n297) );
  NAND U708 ( .A(n299), .B(n300), .Z(xin[193]) );
  NANDN U709 ( .A(start), .B(xreg[193]), .Z(n300) );
  NAND U710 ( .A(x[193]), .B(start), .Z(n299) );
  NAND U711 ( .A(n301), .B(n302), .Z(xin[192]) );
  NANDN U712 ( .A(start), .B(xreg[192]), .Z(n302) );
  NAND U713 ( .A(x[192]), .B(start), .Z(n301) );
  NAND U714 ( .A(n303), .B(n304), .Z(xin[191]) );
  NANDN U715 ( .A(start), .B(xreg[191]), .Z(n304) );
  NAND U716 ( .A(x[191]), .B(start), .Z(n303) );
  NAND U717 ( .A(n305), .B(n306), .Z(xin[190]) );
  NANDN U718 ( .A(start), .B(xreg[190]), .Z(n306) );
  NAND U719 ( .A(x[190]), .B(start), .Z(n305) );
  NAND U720 ( .A(n307), .B(n308), .Z(xin[18]) );
  NANDN U721 ( .A(start), .B(xreg[18]), .Z(n308) );
  NAND U722 ( .A(x[18]), .B(start), .Z(n307) );
  NAND U723 ( .A(n309), .B(n310), .Z(xin[189]) );
  NANDN U724 ( .A(start), .B(xreg[189]), .Z(n310) );
  NAND U725 ( .A(x[189]), .B(start), .Z(n309) );
  NAND U726 ( .A(n311), .B(n312), .Z(xin[188]) );
  NANDN U727 ( .A(start), .B(xreg[188]), .Z(n312) );
  NAND U728 ( .A(x[188]), .B(start), .Z(n311) );
  NAND U729 ( .A(n313), .B(n314), .Z(xin[187]) );
  NANDN U730 ( .A(start), .B(xreg[187]), .Z(n314) );
  NAND U731 ( .A(x[187]), .B(start), .Z(n313) );
  NAND U732 ( .A(n315), .B(n316), .Z(xin[186]) );
  NANDN U733 ( .A(start), .B(xreg[186]), .Z(n316) );
  NAND U734 ( .A(x[186]), .B(start), .Z(n315) );
  NAND U735 ( .A(n317), .B(n318), .Z(xin[185]) );
  NANDN U736 ( .A(start), .B(xreg[185]), .Z(n318) );
  NAND U737 ( .A(x[185]), .B(start), .Z(n317) );
  NAND U738 ( .A(n319), .B(n320), .Z(xin[184]) );
  NANDN U739 ( .A(start), .B(xreg[184]), .Z(n320) );
  NAND U740 ( .A(x[184]), .B(start), .Z(n319) );
  NAND U741 ( .A(n321), .B(n322), .Z(xin[183]) );
  NANDN U742 ( .A(start), .B(xreg[183]), .Z(n322) );
  NAND U743 ( .A(x[183]), .B(start), .Z(n321) );
  NAND U744 ( .A(n323), .B(n324), .Z(xin[182]) );
  NANDN U745 ( .A(start), .B(xreg[182]), .Z(n324) );
  NAND U746 ( .A(x[182]), .B(start), .Z(n323) );
  NAND U747 ( .A(n325), .B(n326), .Z(xin[181]) );
  NANDN U748 ( .A(start), .B(xreg[181]), .Z(n326) );
  NAND U749 ( .A(x[181]), .B(start), .Z(n325) );
  NAND U750 ( .A(n327), .B(n328), .Z(xin[180]) );
  NANDN U751 ( .A(start), .B(xreg[180]), .Z(n328) );
  NAND U752 ( .A(x[180]), .B(start), .Z(n327) );
  NAND U753 ( .A(n329), .B(n330), .Z(xin[17]) );
  NANDN U754 ( .A(start), .B(xreg[17]), .Z(n330) );
  NAND U755 ( .A(x[17]), .B(start), .Z(n329) );
  NAND U756 ( .A(n331), .B(n332), .Z(xin[179]) );
  NANDN U757 ( .A(start), .B(xreg[179]), .Z(n332) );
  NAND U758 ( .A(x[179]), .B(start), .Z(n331) );
  NAND U759 ( .A(n333), .B(n334), .Z(xin[178]) );
  NANDN U760 ( .A(start), .B(xreg[178]), .Z(n334) );
  NAND U761 ( .A(x[178]), .B(start), .Z(n333) );
  NAND U762 ( .A(n335), .B(n336), .Z(xin[177]) );
  NANDN U763 ( .A(start), .B(xreg[177]), .Z(n336) );
  NAND U764 ( .A(x[177]), .B(start), .Z(n335) );
  NAND U765 ( .A(n337), .B(n338), .Z(xin[176]) );
  NANDN U766 ( .A(start), .B(xreg[176]), .Z(n338) );
  NAND U767 ( .A(x[176]), .B(start), .Z(n337) );
  NAND U768 ( .A(n339), .B(n340), .Z(xin[175]) );
  NANDN U769 ( .A(start), .B(xreg[175]), .Z(n340) );
  NAND U770 ( .A(x[175]), .B(start), .Z(n339) );
  NAND U771 ( .A(n341), .B(n342), .Z(xin[174]) );
  NANDN U772 ( .A(start), .B(xreg[174]), .Z(n342) );
  NAND U773 ( .A(x[174]), .B(start), .Z(n341) );
  NAND U774 ( .A(n343), .B(n344), .Z(xin[173]) );
  NANDN U775 ( .A(start), .B(xreg[173]), .Z(n344) );
  NAND U776 ( .A(x[173]), .B(start), .Z(n343) );
  NAND U777 ( .A(n345), .B(n346), .Z(xin[172]) );
  NANDN U778 ( .A(start), .B(xreg[172]), .Z(n346) );
  NAND U779 ( .A(x[172]), .B(start), .Z(n345) );
  NAND U780 ( .A(n347), .B(n348), .Z(xin[171]) );
  NANDN U781 ( .A(start), .B(xreg[171]), .Z(n348) );
  NAND U782 ( .A(x[171]), .B(start), .Z(n347) );
  NAND U783 ( .A(n349), .B(n350), .Z(xin[170]) );
  NANDN U784 ( .A(start), .B(xreg[170]), .Z(n350) );
  NAND U785 ( .A(x[170]), .B(start), .Z(n349) );
  NAND U786 ( .A(n351), .B(n352), .Z(xin[16]) );
  NANDN U787 ( .A(start), .B(xreg[16]), .Z(n352) );
  NAND U788 ( .A(x[16]), .B(start), .Z(n351) );
  NAND U789 ( .A(n353), .B(n354), .Z(xin[169]) );
  NANDN U790 ( .A(start), .B(xreg[169]), .Z(n354) );
  NAND U791 ( .A(x[169]), .B(start), .Z(n353) );
  NAND U792 ( .A(n355), .B(n356), .Z(xin[168]) );
  NANDN U793 ( .A(start), .B(xreg[168]), .Z(n356) );
  NAND U794 ( .A(x[168]), .B(start), .Z(n355) );
  NAND U795 ( .A(n357), .B(n358), .Z(xin[167]) );
  NANDN U796 ( .A(start), .B(xreg[167]), .Z(n358) );
  NAND U797 ( .A(x[167]), .B(start), .Z(n357) );
  NAND U798 ( .A(n359), .B(n360), .Z(xin[166]) );
  NANDN U799 ( .A(start), .B(xreg[166]), .Z(n360) );
  NAND U800 ( .A(x[166]), .B(start), .Z(n359) );
  NAND U801 ( .A(n361), .B(n362), .Z(xin[165]) );
  NANDN U802 ( .A(start), .B(xreg[165]), .Z(n362) );
  NAND U803 ( .A(x[165]), .B(start), .Z(n361) );
  NAND U804 ( .A(n363), .B(n364), .Z(xin[164]) );
  NANDN U805 ( .A(start), .B(xreg[164]), .Z(n364) );
  NAND U806 ( .A(x[164]), .B(start), .Z(n363) );
  NAND U807 ( .A(n365), .B(n366), .Z(xin[163]) );
  NANDN U808 ( .A(start), .B(xreg[163]), .Z(n366) );
  NAND U809 ( .A(x[163]), .B(start), .Z(n365) );
  NAND U810 ( .A(n367), .B(n368), .Z(xin[162]) );
  NANDN U811 ( .A(start), .B(xreg[162]), .Z(n368) );
  NAND U812 ( .A(x[162]), .B(start), .Z(n367) );
  NAND U813 ( .A(n369), .B(n370), .Z(xin[161]) );
  NANDN U814 ( .A(start), .B(xreg[161]), .Z(n370) );
  NAND U815 ( .A(x[161]), .B(start), .Z(n369) );
  NAND U816 ( .A(n371), .B(n372), .Z(xin[160]) );
  NANDN U817 ( .A(start), .B(xreg[160]), .Z(n372) );
  NAND U818 ( .A(x[160]), .B(start), .Z(n371) );
  NAND U819 ( .A(n373), .B(n374), .Z(xin[15]) );
  NANDN U820 ( .A(start), .B(xreg[15]), .Z(n374) );
  NAND U821 ( .A(x[15]), .B(start), .Z(n373) );
  NAND U822 ( .A(n375), .B(n376), .Z(xin[159]) );
  NANDN U823 ( .A(start), .B(xreg[159]), .Z(n376) );
  NAND U824 ( .A(x[159]), .B(start), .Z(n375) );
  NAND U825 ( .A(n377), .B(n378), .Z(xin[158]) );
  NANDN U826 ( .A(start), .B(xreg[158]), .Z(n378) );
  NAND U827 ( .A(x[158]), .B(start), .Z(n377) );
  NAND U828 ( .A(n379), .B(n380), .Z(xin[157]) );
  NANDN U829 ( .A(start), .B(xreg[157]), .Z(n380) );
  NAND U830 ( .A(x[157]), .B(start), .Z(n379) );
  NAND U831 ( .A(n381), .B(n382), .Z(xin[156]) );
  NANDN U832 ( .A(start), .B(xreg[156]), .Z(n382) );
  NAND U833 ( .A(x[156]), .B(start), .Z(n381) );
  NAND U834 ( .A(n383), .B(n384), .Z(xin[155]) );
  NANDN U835 ( .A(start), .B(xreg[155]), .Z(n384) );
  NAND U836 ( .A(x[155]), .B(start), .Z(n383) );
  NAND U837 ( .A(n385), .B(n386), .Z(xin[154]) );
  NANDN U838 ( .A(start), .B(xreg[154]), .Z(n386) );
  NAND U839 ( .A(x[154]), .B(start), .Z(n385) );
  NAND U840 ( .A(n387), .B(n388), .Z(xin[153]) );
  NANDN U841 ( .A(start), .B(xreg[153]), .Z(n388) );
  NAND U842 ( .A(x[153]), .B(start), .Z(n387) );
  NAND U843 ( .A(n389), .B(n390), .Z(xin[152]) );
  NANDN U844 ( .A(start), .B(xreg[152]), .Z(n390) );
  NAND U845 ( .A(x[152]), .B(start), .Z(n389) );
  NAND U846 ( .A(n391), .B(n392), .Z(xin[151]) );
  NANDN U847 ( .A(start), .B(xreg[151]), .Z(n392) );
  NAND U848 ( .A(x[151]), .B(start), .Z(n391) );
  NAND U849 ( .A(n393), .B(n394), .Z(xin[150]) );
  NANDN U850 ( .A(start), .B(xreg[150]), .Z(n394) );
  NAND U851 ( .A(x[150]), .B(start), .Z(n393) );
  NAND U852 ( .A(n395), .B(n396), .Z(xin[14]) );
  NANDN U853 ( .A(start), .B(xreg[14]), .Z(n396) );
  NAND U854 ( .A(x[14]), .B(start), .Z(n395) );
  NAND U855 ( .A(n397), .B(n398), .Z(xin[149]) );
  NANDN U856 ( .A(start), .B(xreg[149]), .Z(n398) );
  NAND U857 ( .A(x[149]), .B(start), .Z(n397) );
  NAND U858 ( .A(n399), .B(n400), .Z(xin[148]) );
  NANDN U859 ( .A(start), .B(xreg[148]), .Z(n400) );
  NAND U860 ( .A(x[148]), .B(start), .Z(n399) );
  NAND U861 ( .A(n401), .B(n402), .Z(xin[147]) );
  NANDN U862 ( .A(start), .B(xreg[147]), .Z(n402) );
  NAND U863 ( .A(x[147]), .B(start), .Z(n401) );
  NAND U864 ( .A(n403), .B(n404), .Z(xin[146]) );
  NANDN U865 ( .A(start), .B(xreg[146]), .Z(n404) );
  NAND U866 ( .A(x[146]), .B(start), .Z(n403) );
  NAND U867 ( .A(n405), .B(n406), .Z(xin[145]) );
  NANDN U868 ( .A(start), .B(xreg[145]), .Z(n406) );
  NAND U869 ( .A(x[145]), .B(start), .Z(n405) );
  NAND U870 ( .A(n407), .B(n408), .Z(xin[144]) );
  NANDN U871 ( .A(start), .B(xreg[144]), .Z(n408) );
  NAND U872 ( .A(x[144]), .B(start), .Z(n407) );
  NAND U873 ( .A(n409), .B(n410), .Z(xin[143]) );
  NANDN U874 ( .A(start), .B(xreg[143]), .Z(n410) );
  NAND U875 ( .A(x[143]), .B(start), .Z(n409) );
  NAND U876 ( .A(n411), .B(n412), .Z(xin[142]) );
  NANDN U877 ( .A(start), .B(xreg[142]), .Z(n412) );
  NAND U878 ( .A(x[142]), .B(start), .Z(n411) );
  NAND U879 ( .A(n413), .B(n414), .Z(xin[141]) );
  NANDN U880 ( .A(start), .B(xreg[141]), .Z(n414) );
  NAND U881 ( .A(x[141]), .B(start), .Z(n413) );
  NAND U882 ( .A(n415), .B(n416), .Z(xin[140]) );
  NANDN U883 ( .A(start), .B(xreg[140]), .Z(n416) );
  NAND U884 ( .A(x[140]), .B(start), .Z(n415) );
  NAND U885 ( .A(n417), .B(n418), .Z(xin[13]) );
  NANDN U886 ( .A(start), .B(xreg[13]), .Z(n418) );
  NAND U887 ( .A(x[13]), .B(start), .Z(n417) );
  NAND U888 ( .A(n419), .B(n420), .Z(xin[139]) );
  NANDN U889 ( .A(start), .B(xreg[139]), .Z(n420) );
  NAND U890 ( .A(x[139]), .B(start), .Z(n419) );
  NAND U891 ( .A(n421), .B(n422), .Z(xin[138]) );
  NANDN U892 ( .A(start), .B(xreg[138]), .Z(n422) );
  NAND U893 ( .A(x[138]), .B(start), .Z(n421) );
  NAND U894 ( .A(n423), .B(n424), .Z(xin[137]) );
  NANDN U895 ( .A(start), .B(xreg[137]), .Z(n424) );
  NAND U896 ( .A(x[137]), .B(start), .Z(n423) );
  NAND U897 ( .A(n425), .B(n426), .Z(xin[136]) );
  NANDN U898 ( .A(start), .B(xreg[136]), .Z(n426) );
  NAND U899 ( .A(x[136]), .B(start), .Z(n425) );
  NAND U900 ( .A(n427), .B(n428), .Z(xin[135]) );
  NANDN U901 ( .A(start), .B(xreg[135]), .Z(n428) );
  NAND U902 ( .A(x[135]), .B(start), .Z(n427) );
  NAND U903 ( .A(n429), .B(n430), .Z(xin[134]) );
  NANDN U904 ( .A(start), .B(xreg[134]), .Z(n430) );
  NAND U905 ( .A(x[134]), .B(start), .Z(n429) );
  NAND U906 ( .A(n431), .B(n432), .Z(xin[133]) );
  NANDN U907 ( .A(start), .B(xreg[133]), .Z(n432) );
  NAND U908 ( .A(x[133]), .B(start), .Z(n431) );
  NAND U909 ( .A(n433), .B(n434), .Z(xin[132]) );
  NANDN U910 ( .A(start), .B(xreg[132]), .Z(n434) );
  NAND U911 ( .A(x[132]), .B(start), .Z(n433) );
  NAND U912 ( .A(n435), .B(n436), .Z(xin[131]) );
  NANDN U913 ( .A(start), .B(xreg[131]), .Z(n436) );
  NAND U914 ( .A(x[131]), .B(start), .Z(n435) );
  NAND U915 ( .A(n437), .B(n438), .Z(xin[130]) );
  NANDN U916 ( .A(start), .B(xreg[130]), .Z(n438) );
  NAND U917 ( .A(x[130]), .B(start), .Z(n437) );
  NAND U918 ( .A(n439), .B(n440), .Z(xin[12]) );
  NANDN U919 ( .A(start), .B(xreg[12]), .Z(n440) );
  NAND U920 ( .A(x[12]), .B(start), .Z(n439) );
  NAND U921 ( .A(n441), .B(n442), .Z(xin[129]) );
  NANDN U922 ( .A(start), .B(xreg[129]), .Z(n442) );
  NAND U923 ( .A(x[129]), .B(start), .Z(n441) );
  NAND U924 ( .A(n443), .B(n444), .Z(xin[128]) );
  NANDN U925 ( .A(start), .B(xreg[128]), .Z(n444) );
  NAND U926 ( .A(x[128]), .B(start), .Z(n443) );
  NAND U927 ( .A(n445), .B(n446), .Z(xin[127]) );
  NANDN U928 ( .A(start), .B(xreg[127]), .Z(n446) );
  NAND U929 ( .A(x[127]), .B(start), .Z(n445) );
  NAND U930 ( .A(n447), .B(n448), .Z(xin[126]) );
  NANDN U931 ( .A(start), .B(xreg[126]), .Z(n448) );
  NAND U932 ( .A(x[126]), .B(start), .Z(n447) );
  NAND U933 ( .A(n449), .B(n450), .Z(xin[125]) );
  NANDN U934 ( .A(start), .B(xreg[125]), .Z(n450) );
  NAND U935 ( .A(x[125]), .B(start), .Z(n449) );
  NAND U936 ( .A(n451), .B(n452), .Z(xin[124]) );
  NANDN U937 ( .A(start), .B(xreg[124]), .Z(n452) );
  NAND U938 ( .A(x[124]), .B(start), .Z(n451) );
  NAND U939 ( .A(n453), .B(n454), .Z(xin[123]) );
  NANDN U940 ( .A(start), .B(xreg[123]), .Z(n454) );
  NAND U941 ( .A(x[123]), .B(start), .Z(n453) );
  NAND U942 ( .A(n455), .B(n456), .Z(xin[122]) );
  NANDN U943 ( .A(start), .B(xreg[122]), .Z(n456) );
  NAND U944 ( .A(x[122]), .B(start), .Z(n455) );
  NAND U945 ( .A(n457), .B(n458), .Z(xin[121]) );
  NANDN U946 ( .A(start), .B(xreg[121]), .Z(n458) );
  NAND U947 ( .A(x[121]), .B(start), .Z(n457) );
  NAND U948 ( .A(n459), .B(n460), .Z(xin[120]) );
  NANDN U949 ( .A(start), .B(xreg[120]), .Z(n460) );
  NAND U950 ( .A(x[120]), .B(start), .Z(n459) );
  NAND U951 ( .A(n461), .B(n462), .Z(xin[11]) );
  NANDN U952 ( .A(start), .B(xreg[11]), .Z(n462) );
  NAND U953 ( .A(x[11]), .B(start), .Z(n461) );
  NAND U954 ( .A(n463), .B(n464), .Z(xin[119]) );
  NANDN U955 ( .A(start), .B(xreg[119]), .Z(n464) );
  NAND U956 ( .A(x[119]), .B(start), .Z(n463) );
  NAND U957 ( .A(n465), .B(n466), .Z(xin[118]) );
  NANDN U958 ( .A(start), .B(xreg[118]), .Z(n466) );
  NAND U959 ( .A(x[118]), .B(start), .Z(n465) );
  NAND U960 ( .A(n467), .B(n468), .Z(xin[117]) );
  NANDN U961 ( .A(start), .B(xreg[117]), .Z(n468) );
  NAND U962 ( .A(x[117]), .B(start), .Z(n467) );
  NAND U963 ( .A(n469), .B(n470), .Z(xin[116]) );
  NANDN U964 ( .A(start), .B(xreg[116]), .Z(n470) );
  NAND U965 ( .A(x[116]), .B(start), .Z(n469) );
  NAND U966 ( .A(n471), .B(n472), .Z(xin[115]) );
  NANDN U967 ( .A(start), .B(xreg[115]), .Z(n472) );
  NAND U968 ( .A(x[115]), .B(start), .Z(n471) );
  NAND U969 ( .A(n473), .B(n474), .Z(xin[114]) );
  NANDN U970 ( .A(start), .B(xreg[114]), .Z(n474) );
  NAND U971 ( .A(x[114]), .B(start), .Z(n473) );
  NAND U972 ( .A(n475), .B(n476), .Z(xin[113]) );
  NANDN U973 ( .A(start), .B(xreg[113]), .Z(n476) );
  NAND U974 ( .A(x[113]), .B(start), .Z(n475) );
  NAND U975 ( .A(n477), .B(n478), .Z(xin[112]) );
  NANDN U976 ( .A(start), .B(xreg[112]), .Z(n478) );
  NAND U977 ( .A(x[112]), .B(start), .Z(n477) );
  NAND U978 ( .A(n479), .B(n480), .Z(xin[111]) );
  NANDN U979 ( .A(start), .B(xreg[111]), .Z(n480) );
  NAND U980 ( .A(x[111]), .B(start), .Z(n479) );
  NAND U981 ( .A(n481), .B(n482), .Z(xin[110]) );
  NANDN U982 ( .A(start), .B(xreg[110]), .Z(n482) );
  NAND U983 ( .A(x[110]), .B(start), .Z(n481) );
  NAND U984 ( .A(n483), .B(n484), .Z(xin[10]) );
  NANDN U985 ( .A(start), .B(xreg[10]), .Z(n484) );
  NAND U986 ( .A(x[10]), .B(start), .Z(n483) );
  NAND U987 ( .A(n485), .B(n486), .Z(xin[109]) );
  NANDN U988 ( .A(start), .B(xreg[109]), .Z(n486) );
  NAND U989 ( .A(x[109]), .B(start), .Z(n485) );
  NAND U990 ( .A(n487), .B(n488), .Z(xin[108]) );
  NANDN U991 ( .A(start), .B(xreg[108]), .Z(n488) );
  NAND U992 ( .A(x[108]), .B(start), .Z(n487) );
  NAND U993 ( .A(n489), .B(n490), .Z(xin[107]) );
  NANDN U994 ( .A(start), .B(xreg[107]), .Z(n490) );
  NAND U995 ( .A(x[107]), .B(start), .Z(n489) );
  NAND U996 ( .A(n491), .B(n492), .Z(xin[106]) );
  NANDN U997 ( .A(start), .B(xreg[106]), .Z(n492) );
  NAND U998 ( .A(x[106]), .B(start), .Z(n491) );
  NAND U999 ( .A(n493), .B(n494), .Z(xin[105]) );
  NANDN U1000 ( .A(start), .B(xreg[105]), .Z(n494) );
  NAND U1001 ( .A(x[105]), .B(start), .Z(n493) );
  NAND U1002 ( .A(n495), .B(n496), .Z(xin[104]) );
  NANDN U1003 ( .A(start), .B(xreg[104]), .Z(n496) );
  NAND U1004 ( .A(x[104]), .B(start), .Z(n495) );
  NAND U1005 ( .A(n497), .B(n498), .Z(xin[103]) );
  NANDN U1006 ( .A(start), .B(xreg[103]), .Z(n498) );
  NAND U1007 ( .A(x[103]), .B(start), .Z(n497) );
  NAND U1008 ( .A(n499), .B(n500), .Z(xin[102]) );
  NANDN U1009 ( .A(start), .B(xreg[102]), .Z(n500) );
  NAND U1010 ( .A(x[102]), .B(start), .Z(n499) );
  NAND U1011 ( .A(n501), .B(n502), .Z(xin[101]) );
  NANDN U1012 ( .A(start), .B(xreg[101]), .Z(n502) );
  NAND U1013 ( .A(x[101]), .B(start), .Z(n501) );
  NAND U1014 ( .A(n503), .B(n504), .Z(xin[100]) );
  NANDN U1015 ( .A(start), .B(xreg[100]), .Z(n504) );
  NAND U1016 ( .A(x[100]), .B(start), .Z(n503) );
  AND U1017 ( .A(x[3]), .B(start), .Z(n505) );
  AND U1018 ( .A(x[2]), .B(start), .Z(n506) );
  AND U1019 ( .A(x[1]), .B(start), .Z(n507) );
  AND U1020 ( .A(x[0]), .B(start), .Z(n508) );
endmodule


module modexp_2N_NN_N256_CC32768 ( clk, rst, m, e, n, c );
  input [255:0] m;
  input [255:0] e;
  input [255:0] n;
  output [255:0] c;
  input clk, rst;
  wire   init, mul_pow, first_one, n3346, n3347, n3348, n3349, n3350, n3351,
         n3352, n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361,
         n3362, n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371,
         n3372, n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381,
         n3382, n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391,
         n3392, n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401,
         n3402, n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411,
         n3412, n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421,
         n3422, n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431,
         n3432, n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441,
         n3442, n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451,
         n3452, n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461,
         n3462, n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471,
         n3472, n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481,
         n3482, n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491,
         n3492, n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501,
         n3502, n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511,
         n3512, n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521,
         n3522, n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531,
         n3532, n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541,
         n3542, n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551,
         n3552, n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561,
         n3562, n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571,
         n3572, n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581,
         n3582, n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591,
         n3592, n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601,
         n3602, n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611,
         n3612, n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621,
         n3622, n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631,
         n3632, n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641,
         n3642, n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651,
         n3652, n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661,
         n3662, n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671,
         n3672, n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681,
         n3682, n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691,
         n3692, n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701,
         n3702, n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711,
         n3712, n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721,
         n3722, n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731,
         n3732, n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741,
         n3742, n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751,
         n3752, n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761,
         n3762, n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771,
         n3772, n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781,
         n3782, n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791,
         n3792, n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801,
         n3802, n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811,
         n3812, n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821,
         n3822, n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831,
         n3832, n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841,
         n3842, n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851,
         n3852, n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861,
         n3862, n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871,
         n3872, n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881,
         n3882, n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891,
         n3892, n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901,
         n3902, n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911,
         n3912, n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921,
         n3922, n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931,
         n3932, n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941,
         n3942, n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951,
         n3952, n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961,
         n3962, n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971,
         n3972, n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981,
         n3982, n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991,
         n3992, n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001,
         n4002, n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011,
         n4012, n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021,
         n4022, n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031,
         n4032, n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041,
         n4042, n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051,
         n4052, n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061,
         n4062, n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071,
         n4072, n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081,
         n4082, n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091,
         n4092, n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101,
         n4102, n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111,
         n4112, n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121,
         n4122, n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131,
         n4132, n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141,
         n4142, n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151,
         n4152, n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161,
         n4162, n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171,
         n4172, n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181,
         n4182, n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191,
         n4192, n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201,
         n4202, n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211,
         n4212, n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221,
         n4222, n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231,
         n4232, n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241,
         n4242, n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251,
         n4252, n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261,
         n4262, n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271,
         n4272, n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281,
         n4282, n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291,
         n4292, n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301,
         n4302, n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311,
         n4312, n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321,
         n4322, n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331,
         n4332, n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341,
         n4342, n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351,
         n4352, n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361,
         n4362, n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371,
         n4372, n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381,
         n4382, n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391,
         n4392, n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401,
         n4402, n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411,
         n4412, n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421,
         n4422, n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431,
         n4432, n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441,
         n4442, n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451,
         n4452, n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461,
         n4462, n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471,
         n4472, n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481,
         n4482, n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491,
         n4492, n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501,
         n4502, n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511,
         n4512, n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521,
         n4522, n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531,
         n4532, n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541,
         n4542, n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551,
         n4552, n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561,
         n4562, n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571,
         n4572, n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581,
         n4582, n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591,
         n4592, n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601,
         n4602, n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611,
         n4612, n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621,
         n4622, n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631,
         n4632, n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641,
         n4642, n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651,
         n4652, n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661,
         n4662, n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671,
         n4672, n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681,
         n4682, n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691,
         n4692, n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701,
         n4702, n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711,
         n4712, n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721,
         n4722, n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731,
         n4732, n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741,
         n4742, n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751,
         n4752, n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761,
         n4762, n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771,
         n4772, n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781,
         n4782, n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791,
         n4792, n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801,
         n4802, n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811,
         n4812, n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821,
         n4822, n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831,
         n4832, n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841,
         n4842, n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851,
         n4852, n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861,
         n4862, n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871,
         n4872, n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881,
         n4882, n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891,
         n4892, n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901,
         n4902, n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911,
         n4912, n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921,
         n4922, n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931,
         n4932, n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941,
         n4942, n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951,
         n4952, n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961,
         n4962, n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971,
         n4972, n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981,
         n4982, n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991,
         n4992, n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001,
         n5002, n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011,
         n5012, n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021,
         n5022, n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031,
         n5032, n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041,
         n5042, n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051,
         n5052, n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061,
         n5062, n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071,
         n5072, n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081,
         n5082, n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091,
         n5092, n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101,
         n5102, n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111,
         n5112, n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121,
         n5122, n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131,
         n5132, n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141,
         n5142, n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151,
         n5152, n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161,
         n5162, n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171,
         n5172, n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181,
         n5182, n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191,
         n5192, n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201,
         n5202, n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211,
         n5212, n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221,
         n5222, n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231,
         n5232, n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241,
         n5242, n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251,
         n5252, n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261,
         n5262, n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271,
         n5272, n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281,
         n5282, n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291,
         n5292, n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301,
         n5302, n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311,
         n5312, n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321,
         n5322, n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331,
         n5332, n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341,
         n5342, n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351,
         n5352, n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361,
         n5362, n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371,
         n5372, n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381,
         n5382, n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391,
         n5392, n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401,
         n5402, n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411,
         n5412, n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421,
         n5422, n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431,
         n5432, n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441,
         n5442, n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451,
         n5452, n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461,
         n5462, n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471,
         n5472, n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481,
         n5482, n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491,
         n5492, n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501,
         n5502, n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511,
         n5512, n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521,
         n5522, n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531,
         n5532, n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541,
         n5542, n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551,
         n5552, n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561,
         n5562, n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571,
         n5572, n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581,
         n5582, n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591,
         n5592, n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601,
         n5602, n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611,
         n5612, n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621,
         n5622, n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631,
         n5632, n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641,
         n5642, n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651,
         n5652, n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661,
         n5662, n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671,
         n5672, n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681,
         n5682, n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691,
         n5692, n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701,
         n5702, n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711,
         n5712, n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721,
         n5722, n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731,
         n5732, n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741,
         n5742, n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751,
         n5752, n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761,
         n5762, n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771,
         n5772, n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781,
         n5782, n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791,
         n5792, n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801,
         n5802, n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811,
         n5812, n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821,
         n5822, n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831,
         n5832, n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841,
         n5842, n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851,
         n5852, n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861,
         n5862, n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871,
         n5872, n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881,
         n5882, n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891,
         n5892, n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901,
         n5902, n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911,
         n5912, n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921,
         n5922, n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931,
         n5932, n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941,
         n5942, n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951,
         n5952, n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961,
         n5962, n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971,
         n5972, n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981,
         n5982, n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991,
         n5992, n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001,
         n6002, n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011,
         n6012, n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021,
         n6022, n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031,
         n6032, n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041,
         n6042, n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051,
         n6052, n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061,
         n6062, n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071,
         n6072, n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081,
         n6082, n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091,
         n6092, n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101,
         n6102, n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111,
         n6112, n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121,
         n6122, n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131,
         n6132, n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141,
         n6142, n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151,
         n6152, n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161,
         n6162, n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171,
         n6172, n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181,
         n6182, n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191,
         n6192, n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201,
         n6202, n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211,
         n6212, n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221,
         n6222, n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231,
         n6232, n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241,
         n6242, n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251,
         n6252, n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261,
         n6262, n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271,
         n6272, n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281,
         n6282, n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291,
         n6292, n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301,
         n6302, n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311,
         n6312, n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321,
         n6322, n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331,
         n6332, n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341,
         n6342, n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351,
         n6352, n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361,
         n6362, n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371,
         n6372, n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381,
         n6382, n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391,
         n6392, n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401,
         n6402, n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411,
         n6412, n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421,
         n6422, n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431,
         n6432, n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441,
         n6442, n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451,
         n6452, n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461,
         n6462, n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471,
         n6472, n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481,
         n6482, n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491,
         n6492, n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501,
         n6502, n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511,
         n6512, n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521,
         n6522, n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531,
         n6532, n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541,
         n6542, n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551,
         n6552, n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561,
         n6562, n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571,
         n6572, n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581,
         n6582, n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591,
         n6592, n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601,
         n6602, n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611,
         n6612, n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621,
         n6622, n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631,
         n6632, n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641,
         n6642, n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651,
         n6652, n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661,
         n6662, n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671,
         n6672, n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681,
         n6682, n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691,
         n6692, n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701,
         n6702, n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711,
         n6712, n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721,
         n6722, n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731,
         n6732, n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741,
         n6742, n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751,
         n6752, n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761,
         n6762, n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771,
         n6772, n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781,
         n6782, n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791,
         n6792, n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801,
         n6802, n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811,
         n6812, n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821,
         n6822, n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831,
         n6832, n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841,
         n6842, n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851,
         n6852, n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861,
         n6862, n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871,
         n6872, n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881,
         n6882, n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891,
         n6892, n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901,
         n6902, n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911,
         n6912, n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921,
         n6922, n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931,
         n6932, n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941,
         n6942, n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951,
         n6952, n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961,
         n6962, n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971,
         n6972, n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981,
         n6982, n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991,
         n6992, n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001,
         n7002, n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011,
         n7012, n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021,
         n7022, n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031,
         n7032, n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041,
         n7042, n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051,
         n7052, n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061,
         n7062, n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071,
         n7072, n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081,
         n7082, n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091,
         n7092, n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101,
         n7102, n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111,
         n7112, n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121,
         n7122, n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131,
         n7132, n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141,
         n7142, n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151,
         n7152, n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161,
         n7162, n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171,
         n7172, n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181,
         n7182, n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191,
         n7192, n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201,
         n7202, n7203, n7204;
  wire   [63:0] start_in;
  wire   [63:0] start_reg;
  wire   [255:0] ereg;
  wire   [255:0] o;
  wire   [255:0] creg;
  wire   [255:0] x;
  wire   [255:0] y;

  DFF init_reg ( .D(1'b1), .CLK(clk), .RST(rst), .Q(init) );
  DFF \start_reg_reg[0]  ( .D(n7204), .CLK(clk), .RST(rst), .Q(start_reg[0])
         );
  DFF \start_reg_reg[1]  ( .D(start_in[0]), .CLK(clk), .RST(rst), .Q(
        start_reg[1]) );
  DFF \start_reg_reg[2]  ( .D(start_in[1]), .CLK(clk), .RST(rst), .Q(
        start_reg[2]) );
  DFF \start_reg_reg[3]  ( .D(start_in[2]), .CLK(clk), .RST(rst), .Q(
        start_reg[3]) );
  DFF \start_reg_reg[4]  ( .D(start_in[3]), .CLK(clk), .RST(rst), .Q(
        start_reg[4]) );
  DFF \start_reg_reg[5]  ( .D(start_in[4]), .CLK(clk), .RST(rst), .Q(
        start_reg[5]) );
  DFF \start_reg_reg[6]  ( .D(start_in[5]), .CLK(clk), .RST(rst), .Q(
        start_reg[6]) );
  DFF \start_reg_reg[7]  ( .D(start_in[6]), .CLK(clk), .RST(rst), .Q(
        start_reg[7]) );
  DFF \start_reg_reg[8]  ( .D(start_in[7]), .CLK(clk), .RST(rst), .Q(
        start_reg[8]) );
  DFF \start_reg_reg[9]  ( .D(start_in[8]), .CLK(clk), .RST(rst), .Q(
        start_reg[9]) );
  DFF \start_reg_reg[10]  ( .D(start_in[9]), .CLK(clk), .RST(rst), .Q(
        start_reg[10]) );
  DFF \start_reg_reg[11]  ( .D(start_in[10]), .CLK(clk), .RST(rst), .Q(
        start_reg[11]) );
  DFF \start_reg_reg[12]  ( .D(start_in[11]), .CLK(clk), .RST(rst), .Q(
        start_reg[12]) );
  DFF \start_reg_reg[13]  ( .D(start_in[12]), .CLK(clk), .RST(rst), .Q(
        start_reg[13]) );
  DFF \start_reg_reg[14]  ( .D(start_in[13]), .CLK(clk), .RST(rst), .Q(
        start_reg[14]) );
  DFF \start_reg_reg[15]  ( .D(start_in[14]), .CLK(clk), .RST(rst), .Q(
        start_reg[15]) );
  DFF \start_reg_reg[16]  ( .D(start_in[15]), .CLK(clk), .RST(rst), .Q(
        start_reg[16]) );
  DFF \start_reg_reg[17]  ( .D(start_in[16]), .CLK(clk), .RST(rst), .Q(
        start_reg[17]) );
  DFF \start_reg_reg[18]  ( .D(start_in[17]), .CLK(clk), .RST(rst), .Q(
        start_reg[18]) );
  DFF \start_reg_reg[19]  ( .D(start_in[18]), .CLK(clk), .RST(rst), .Q(
        start_reg[19]) );
  DFF \start_reg_reg[20]  ( .D(start_in[19]), .CLK(clk), .RST(rst), .Q(
        start_reg[20]) );
  DFF \start_reg_reg[21]  ( .D(start_in[20]), .CLK(clk), .RST(rst), .Q(
        start_reg[21]) );
  DFF \start_reg_reg[22]  ( .D(start_in[21]), .CLK(clk), .RST(rst), .Q(
        start_reg[22]) );
  DFF \start_reg_reg[23]  ( .D(start_in[22]), .CLK(clk), .RST(rst), .Q(
        start_reg[23]) );
  DFF \start_reg_reg[24]  ( .D(start_in[23]), .CLK(clk), .RST(rst), .Q(
        start_reg[24]) );
  DFF \start_reg_reg[25]  ( .D(start_in[24]), .CLK(clk), .RST(rst), .Q(
        start_reg[25]) );
  DFF \start_reg_reg[26]  ( .D(start_in[25]), .CLK(clk), .RST(rst), .Q(
        start_reg[26]) );
  DFF \start_reg_reg[27]  ( .D(start_in[26]), .CLK(clk), .RST(rst), .Q(
        start_reg[27]) );
  DFF \start_reg_reg[28]  ( .D(start_in[27]), .CLK(clk), .RST(rst), .Q(
        start_reg[28]) );
  DFF \start_reg_reg[29]  ( .D(start_in[28]), .CLK(clk), .RST(rst), .Q(
        start_reg[29]) );
  DFF \start_reg_reg[30]  ( .D(start_in[29]), .CLK(clk), .RST(rst), .Q(
        start_reg[30]) );
  DFF \start_reg_reg[31]  ( .D(start_in[30]), .CLK(clk), .RST(rst), .Q(
        start_reg[31]) );
  DFF \start_reg_reg[32]  ( .D(start_in[31]), .CLK(clk), .RST(rst), .Q(
        start_reg[32]) );
  DFF \start_reg_reg[33]  ( .D(start_in[32]), .CLK(clk), .RST(rst), .Q(
        start_reg[33]) );
  DFF \start_reg_reg[34]  ( .D(start_in[33]), .CLK(clk), .RST(rst), .Q(
        start_reg[34]) );
  DFF \start_reg_reg[35]  ( .D(start_in[34]), .CLK(clk), .RST(rst), .Q(
        start_reg[35]) );
  DFF \start_reg_reg[36]  ( .D(start_in[35]), .CLK(clk), .RST(rst), .Q(
        start_reg[36]) );
  DFF \start_reg_reg[37]  ( .D(start_in[36]), .CLK(clk), .RST(rst), .Q(
        start_reg[37]) );
  DFF \start_reg_reg[38]  ( .D(start_in[37]), .CLK(clk), .RST(rst), .Q(
        start_reg[38]) );
  DFF \start_reg_reg[39]  ( .D(start_in[38]), .CLK(clk), .RST(rst), .Q(
        start_reg[39]) );
  DFF \start_reg_reg[40]  ( .D(start_in[39]), .CLK(clk), .RST(rst), .Q(
        start_reg[40]) );
  DFF \start_reg_reg[41]  ( .D(start_in[40]), .CLK(clk), .RST(rst), .Q(
        start_reg[41]) );
  DFF \start_reg_reg[42]  ( .D(start_in[41]), .CLK(clk), .RST(rst), .Q(
        start_reg[42]) );
  DFF \start_reg_reg[43]  ( .D(start_in[42]), .CLK(clk), .RST(rst), .Q(
        start_reg[43]) );
  DFF \start_reg_reg[44]  ( .D(start_in[43]), .CLK(clk), .RST(rst), .Q(
        start_reg[44]) );
  DFF \start_reg_reg[45]  ( .D(start_in[44]), .CLK(clk), .RST(rst), .Q(
        start_reg[45]) );
  DFF \start_reg_reg[46]  ( .D(start_in[45]), .CLK(clk), .RST(rst), .Q(
        start_reg[46]) );
  DFF \start_reg_reg[47]  ( .D(start_in[46]), .CLK(clk), .RST(rst), .Q(
        start_reg[47]) );
  DFF \start_reg_reg[48]  ( .D(start_in[47]), .CLK(clk), .RST(rst), .Q(
        start_reg[48]) );
  DFF \start_reg_reg[49]  ( .D(start_in[48]), .CLK(clk), .RST(rst), .Q(
        start_reg[49]) );
  DFF \start_reg_reg[50]  ( .D(start_in[49]), .CLK(clk), .RST(rst), .Q(
        start_reg[50]) );
  DFF \start_reg_reg[51]  ( .D(start_in[50]), .CLK(clk), .RST(rst), .Q(
        start_reg[51]) );
  DFF \start_reg_reg[52]  ( .D(start_in[51]), .CLK(clk), .RST(rst), .Q(
        start_reg[52]) );
  DFF \start_reg_reg[53]  ( .D(start_in[52]), .CLK(clk), .RST(rst), .Q(
        start_reg[53]) );
  DFF \start_reg_reg[54]  ( .D(start_in[53]), .CLK(clk), .RST(rst), .Q(
        start_reg[54]) );
  DFF \start_reg_reg[55]  ( .D(start_in[54]), .CLK(clk), .RST(rst), .Q(
        start_reg[55]) );
  DFF \start_reg_reg[56]  ( .D(start_in[55]), .CLK(clk), .RST(rst), .Q(
        start_reg[56]) );
  DFF \start_reg_reg[57]  ( .D(start_in[56]), .CLK(clk), .RST(rst), .Q(
        start_reg[57]) );
  DFF \start_reg_reg[58]  ( .D(start_in[57]), .CLK(clk), .RST(rst), .Q(
        start_reg[58]) );
  DFF \start_reg_reg[59]  ( .D(start_in[58]), .CLK(clk), .RST(rst), .Q(
        start_reg[59]) );
  DFF \start_reg_reg[60]  ( .D(start_in[59]), .CLK(clk), .RST(rst), .Q(
        start_reg[60]) );
  DFF \start_reg_reg[61]  ( .D(start_in[60]), .CLK(clk), .RST(rst), .Q(
        start_reg[61]) );
  DFF \start_reg_reg[62]  ( .D(start_in[61]), .CLK(clk), .RST(rst), .Q(
        start_reg[62]) );
  DFF \start_reg_reg[63]  ( .D(start_in[62]), .CLK(clk), .RST(rst), .Q(
        start_reg[63]) );
  DFF mul_pow_reg ( .D(n3859), .CLK(clk), .RST(rst), .Q(mul_pow) );
  DFF \ereg_reg[0]  ( .D(n3858), .CLK(clk), .RST(rst), .Q(ereg[0]) );
  DFF \ereg_reg[1]  ( .D(n3857), .CLK(clk), .RST(rst), .Q(ereg[1]) );
  DFF \ereg_reg[2]  ( .D(n3856), .CLK(clk), .RST(rst), .Q(ereg[2]) );
  DFF \ereg_reg[3]  ( .D(n3855), .CLK(clk), .RST(rst), .Q(ereg[3]) );
  DFF \ereg_reg[4]  ( .D(n3854), .CLK(clk), .RST(rst), .Q(ereg[4]) );
  DFF \ereg_reg[5]  ( .D(n3853), .CLK(clk), .RST(rst), .Q(ereg[5]) );
  DFF \ereg_reg[6]  ( .D(n3852), .CLK(clk), .RST(rst), .Q(ereg[6]) );
  DFF \ereg_reg[7]  ( .D(n3851), .CLK(clk), .RST(rst), .Q(ereg[7]) );
  DFF \ereg_reg[8]  ( .D(n3850), .CLK(clk), .RST(rst), .Q(ereg[8]) );
  DFF \ereg_reg[9]  ( .D(n3849), .CLK(clk), .RST(rst), .Q(ereg[9]) );
  DFF \ereg_reg[10]  ( .D(n3848), .CLK(clk), .RST(rst), .Q(ereg[10]) );
  DFF \ereg_reg[11]  ( .D(n3847), .CLK(clk), .RST(rst), .Q(ereg[11]) );
  DFF \ereg_reg[12]  ( .D(n3846), .CLK(clk), .RST(rst), .Q(ereg[12]) );
  DFF \ereg_reg[13]  ( .D(n3845), .CLK(clk), .RST(rst), .Q(ereg[13]) );
  DFF \ereg_reg[14]  ( .D(n3844), .CLK(clk), .RST(rst), .Q(ereg[14]) );
  DFF \ereg_reg[15]  ( .D(n3843), .CLK(clk), .RST(rst), .Q(ereg[15]) );
  DFF \ereg_reg[16]  ( .D(n3842), .CLK(clk), .RST(rst), .Q(ereg[16]) );
  DFF \ereg_reg[17]  ( .D(n3841), .CLK(clk), .RST(rst), .Q(ereg[17]) );
  DFF \ereg_reg[18]  ( .D(n3840), .CLK(clk), .RST(rst), .Q(ereg[18]) );
  DFF \ereg_reg[19]  ( .D(n3839), .CLK(clk), .RST(rst), .Q(ereg[19]) );
  DFF \ereg_reg[20]  ( .D(n3838), .CLK(clk), .RST(rst), .Q(ereg[20]) );
  DFF \ereg_reg[21]  ( .D(n3837), .CLK(clk), .RST(rst), .Q(ereg[21]) );
  DFF \ereg_reg[22]  ( .D(n3836), .CLK(clk), .RST(rst), .Q(ereg[22]) );
  DFF \ereg_reg[23]  ( .D(n3835), .CLK(clk), .RST(rst), .Q(ereg[23]) );
  DFF \ereg_reg[24]  ( .D(n3834), .CLK(clk), .RST(rst), .Q(ereg[24]) );
  DFF \ereg_reg[25]  ( .D(n3833), .CLK(clk), .RST(rst), .Q(ereg[25]) );
  DFF \ereg_reg[26]  ( .D(n3832), .CLK(clk), .RST(rst), .Q(ereg[26]) );
  DFF \ereg_reg[27]  ( .D(n3831), .CLK(clk), .RST(rst), .Q(ereg[27]) );
  DFF \ereg_reg[28]  ( .D(n3830), .CLK(clk), .RST(rst), .Q(ereg[28]) );
  DFF \ereg_reg[29]  ( .D(n3829), .CLK(clk), .RST(rst), .Q(ereg[29]) );
  DFF \ereg_reg[30]  ( .D(n3828), .CLK(clk), .RST(rst), .Q(ereg[30]) );
  DFF \ereg_reg[31]  ( .D(n3827), .CLK(clk), .RST(rst), .Q(ereg[31]) );
  DFF \ereg_reg[32]  ( .D(n3826), .CLK(clk), .RST(rst), .Q(ereg[32]) );
  DFF \ereg_reg[33]  ( .D(n3825), .CLK(clk), .RST(rst), .Q(ereg[33]) );
  DFF \ereg_reg[34]  ( .D(n3824), .CLK(clk), .RST(rst), .Q(ereg[34]) );
  DFF \ereg_reg[35]  ( .D(n3823), .CLK(clk), .RST(rst), .Q(ereg[35]) );
  DFF \ereg_reg[36]  ( .D(n3822), .CLK(clk), .RST(rst), .Q(ereg[36]) );
  DFF \ereg_reg[37]  ( .D(n3821), .CLK(clk), .RST(rst), .Q(ereg[37]) );
  DFF \ereg_reg[38]  ( .D(n3820), .CLK(clk), .RST(rst), .Q(ereg[38]) );
  DFF \ereg_reg[39]  ( .D(n3819), .CLK(clk), .RST(rst), .Q(ereg[39]) );
  DFF \ereg_reg[40]  ( .D(n3818), .CLK(clk), .RST(rst), .Q(ereg[40]) );
  DFF \ereg_reg[41]  ( .D(n3817), .CLK(clk), .RST(rst), .Q(ereg[41]) );
  DFF \ereg_reg[42]  ( .D(n3816), .CLK(clk), .RST(rst), .Q(ereg[42]) );
  DFF \ereg_reg[43]  ( .D(n3815), .CLK(clk), .RST(rst), .Q(ereg[43]) );
  DFF \ereg_reg[44]  ( .D(n3814), .CLK(clk), .RST(rst), .Q(ereg[44]) );
  DFF \ereg_reg[45]  ( .D(n3813), .CLK(clk), .RST(rst), .Q(ereg[45]) );
  DFF \ereg_reg[46]  ( .D(n3812), .CLK(clk), .RST(rst), .Q(ereg[46]) );
  DFF \ereg_reg[47]  ( .D(n3811), .CLK(clk), .RST(rst), .Q(ereg[47]) );
  DFF \ereg_reg[48]  ( .D(n3810), .CLK(clk), .RST(rst), .Q(ereg[48]) );
  DFF \ereg_reg[49]  ( .D(n3809), .CLK(clk), .RST(rst), .Q(ereg[49]) );
  DFF \ereg_reg[50]  ( .D(n3808), .CLK(clk), .RST(rst), .Q(ereg[50]) );
  DFF \ereg_reg[51]  ( .D(n3807), .CLK(clk), .RST(rst), .Q(ereg[51]) );
  DFF \ereg_reg[52]  ( .D(n3806), .CLK(clk), .RST(rst), .Q(ereg[52]) );
  DFF \ereg_reg[53]  ( .D(n3805), .CLK(clk), .RST(rst), .Q(ereg[53]) );
  DFF \ereg_reg[54]  ( .D(n3804), .CLK(clk), .RST(rst), .Q(ereg[54]) );
  DFF \ereg_reg[55]  ( .D(n3803), .CLK(clk), .RST(rst), .Q(ereg[55]) );
  DFF \ereg_reg[56]  ( .D(n3802), .CLK(clk), .RST(rst), .Q(ereg[56]) );
  DFF \ereg_reg[57]  ( .D(n3801), .CLK(clk), .RST(rst), .Q(ereg[57]) );
  DFF \ereg_reg[58]  ( .D(n3800), .CLK(clk), .RST(rst), .Q(ereg[58]) );
  DFF \ereg_reg[59]  ( .D(n3799), .CLK(clk), .RST(rst), .Q(ereg[59]) );
  DFF \ereg_reg[60]  ( .D(n3798), .CLK(clk), .RST(rst), .Q(ereg[60]) );
  DFF \ereg_reg[61]  ( .D(n3797), .CLK(clk), .RST(rst), .Q(ereg[61]) );
  DFF \ereg_reg[62]  ( .D(n3796), .CLK(clk), .RST(rst), .Q(ereg[62]) );
  DFF \ereg_reg[63]  ( .D(n3795), .CLK(clk), .RST(rst), .Q(ereg[63]) );
  DFF \ereg_reg[64]  ( .D(n3794), .CLK(clk), .RST(rst), .Q(ereg[64]) );
  DFF \ereg_reg[65]  ( .D(n3793), .CLK(clk), .RST(rst), .Q(ereg[65]) );
  DFF \ereg_reg[66]  ( .D(n3792), .CLK(clk), .RST(rst), .Q(ereg[66]) );
  DFF \ereg_reg[67]  ( .D(n3791), .CLK(clk), .RST(rst), .Q(ereg[67]) );
  DFF \ereg_reg[68]  ( .D(n3790), .CLK(clk), .RST(rst), .Q(ereg[68]) );
  DFF \ereg_reg[69]  ( .D(n3789), .CLK(clk), .RST(rst), .Q(ereg[69]) );
  DFF \ereg_reg[70]  ( .D(n3788), .CLK(clk), .RST(rst), .Q(ereg[70]) );
  DFF \ereg_reg[71]  ( .D(n3787), .CLK(clk), .RST(rst), .Q(ereg[71]) );
  DFF \ereg_reg[72]  ( .D(n3786), .CLK(clk), .RST(rst), .Q(ereg[72]) );
  DFF \ereg_reg[73]  ( .D(n3785), .CLK(clk), .RST(rst), .Q(ereg[73]) );
  DFF \ereg_reg[74]  ( .D(n3784), .CLK(clk), .RST(rst), .Q(ereg[74]) );
  DFF \ereg_reg[75]  ( .D(n3783), .CLK(clk), .RST(rst), .Q(ereg[75]) );
  DFF \ereg_reg[76]  ( .D(n3782), .CLK(clk), .RST(rst), .Q(ereg[76]) );
  DFF \ereg_reg[77]  ( .D(n3781), .CLK(clk), .RST(rst), .Q(ereg[77]) );
  DFF \ereg_reg[78]  ( .D(n3780), .CLK(clk), .RST(rst), .Q(ereg[78]) );
  DFF \ereg_reg[79]  ( .D(n3779), .CLK(clk), .RST(rst), .Q(ereg[79]) );
  DFF \ereg_reg[80]  ( .D(n3778), .CLK(clk), .RST(rst), .Q(ereg[80]) );
  DFF \ereg_reg[81]  ( .D(n3777), .CLK(clk), .RST(rst), .Q(ereg[81]) );
  DFF \ereg_reg[82]  ( .D(n3776), .CLK(clk), .RST(rst), .Q(ereg[82]) );
  DFF \ereg_reg[83]  ( .D(n3775), .CLK(clk), .RST(rst), .Q(ereg[83]) );
  DFF \ereg_reg[84]  ( .D(n3774), .CLK(clk), .RST(rst), .Q(ereg[84]) );
  DFF \ereg_reg[85]  ( .D(n3773), .CLK(clk), .RST(rst), .Q(ereg[85]) );
  DFF \ereg_reg[86]  ( .D(n3772), .CLK(clk), .RST(rst), .Q(ereg[86]) );
  DFF \ereg_reg[87]  ( .D(n3771), .CLK(clk), .RST(rst), .Q(ereg[87]) );
  DFF \ereg_reg[88]  ( .D(n3770), .CLK(clk), .RST(rst), .Q(ereg[88]) );
  DFF \ereg_reg[89]  ( .D(n3769), .CLK(clk), .RST(rst), .Q(ereg[89]) );
  DFF \ereg_reg[90]  ( .D(n3768), .CLK(clk), .RST(rst), .Q(ereg[90]) );
  DFF \ereg_reg[91]  ( .D(n3767), .CLK(clk), .RST(rst), .Q(ereg[91]) );
  DFF \ereg_reg[92]  ( .D(n3766), .CLK(clk), .RST(rst), .Q(ereg[92]) );
  DFF \ereg_reg[93]  ( .D(n3765), .CLK(clk), .RST(rst), .Q(ereg[93]) );
  DFF \ereg_reg[94]  ( .D(n3764), .CLK(clk), .RST(rst), .Q(ereg[94]) );
  DFF \ereg_reg[95]  ( .D(n3763), .CLK(clk), .RST(rst), .Q(ereg[95]) );
  DFF \ereg_reg[96]  ( .D(n3762), .CLK(clk), .RST(rst), .Q(ereg[96]) );
  DFF \ereg_reg[97]  ( .D(n3761), .CLK(clk), .RST(rst), .Q(ereg[97]) );
  DFF \ereg_reg[98]  ( .D(n3760), .CLK(clk), .RST(rst), .Q(ereg[98]) );
  DFF \ereg_reg[99]  ( .D(n3759), .CLK(clk), .RST(rst), .Q(ereg[99]) );
  DFF \ereg_reg[100]  ( .D(n3758), .CLK(clk), .RST(rst), .Q(ereg[100]) );
  DFF \ereg_reg[101]  ( .D(n3757), .CLK(clk), .RST(rst), .Q(ereg[101]) );
  DFF \ereg_reg[102]  ( .D(n3756), .CLK(clk), .RST(rst), .Q(ereg[102]) );
  DFF \ereg_reg[103]  ( .D(n3755), .CLK(clk), .RST(rst), .Q(ereg[103]) );
  DFF \ereg_reg[104]  ( .D(n3754), .CLK(clk), .RST(rst), .Q(ereg[104]) );
  DFF \ereg_reg[105]  ( .D(n3753), .CLK(clk), .RST(rst), .Q(ereg[105]) );
  DFF \ereg_reg[106]  ( .D(n3752), .CLK(clk), .RST(rst), .Q(ereg[106]) );
  DFF \ereg_reg[107]  ( .D(n3751), .CLK(clk), .RST(rst), .Q(ereg[107]) );
  DFF \ereg_reg[108]  ( .D(n3750), .CLK(clk), .RST(rst), .Q(ereg[108]) );
  DFF \ereg_reg[109]  ( .D(n3749), .CLK(clk), .RST(rst), .Q(ereg[109]) );
  DFF \ereg_reg[110]  ( .D(n3748), .CLK(clk), .RST(rst), .Q(ereg[110]) );
  DFF \ereg_reg[111]  ( .D(n3747), .CLK(clk), .RST(rst), .Q(ereg[111]) );
  DFF \ereg_reg[112]  ( .D(n3746), .CLK(clk), .RST(rst), .Q(ereg[112]) );
  DFF \ereg_reg[113]  ( .D(n3745), .CLK(clk), .RST(rst), .Q(ereg[113]) );
  DFF \ereg_reg[114]  ( .D(n3744), .CLK(clk), .RST(rst), .Q(ereg[114]) );
  DFF \ereg_reg[115]  ( .D(n3743), .CLK(clk), .RST(rst), .Q(ereg[115]) );
  DFF \ereg_reg[116]  ( .D(n3742), .CLK(clk), .RST(rst), .Q(ereg[116]) );
  DFF \ereg_reg[117]  ( .D(n3741), .CLK(clk), .RST(rst), .Q(ereg[117]) );
  DFF \ereg_reg[118]  ( .D(n3740), .CLK(clk), .RST(rst), .Q(ereg[118]) );
  DFF \ereg_reg[119]  ( .D(n3739), .CLK(clk), .RST(rst), .Q(ereg[119]) );
  DFF \ereg_reg[120]  ( .D(n3738), .CLK(clk), .RST(rst), .Q(ereg[120]) );
  DFF \ereg_reg[121]  ( .D(n3737), .CLK(clk), .RST(rst), .Q(ereg[121]) );
  DFF \ereg_reg[122]  ( .D(n3736), .CLK(clk), .RST(rst), .Q(ereg[122]) );
  DFF \ereg_reg[123]  ( .D(n3735), .CLK(clk), .RST(rst), .Q(ereg[123]) );
  DFF \ereg_reg[124]  ( .D(n3734), .CLK(clk), .RST(rst), .Q(ereg[124]) );
  DFF \ereg_reg[125]  ( .D(n3733), .CLK(clk), .RST(rst), .Q(ereg[125]) );
  DFF \ereg_reg[126]  ( .D(n3732), .CLK(clk), .RST(rst), .Q(ereg[126]) );
  DFF \ereg_reg[127]  ( .D(n3731), .CLK(clk), .RST(rst), .Q(ereg[127]) );
  DFF \ereg_reg[128]  ( .D(n3730), .CLK(clk), .RST(rst), .Q(ereg[128]) );
  DFF \ereg_reg[129]  ( .D(n3729), .CLK(clk), .RST(rst), .Q(ereg[129]) );
  DFF \ereg_reg[130]  ( .D(n3728), .CLK(clk), .RST(rst), .Q(ereg[130]) );
  DFF \ereg_reg[131]  ( .D(n3727), .CLK(clk), .RST(rst), .Q(ereg[131]) );
  DFF \ereg_reg[132]  ( .D(n3726), .CLK(clk), .RST(rst), .Q(ereg[132]) );
  DFF \ereg_reg[133]  ( .D(n3725), .CLK(clk), .RST(rst), .Q(ereg[133]) );
  DFF \ereg_reg[134]  ( .D(n3724), .CLK(clk), .RST(rst), .Q(ereg[134]) );
  DFF \ereg_reg[135]  ( .D(n3723), .CLK(clk), .RST(rst), .Q(ereg[135]) );
  DFF \ereg_reg[136]  ( .D(n3722), .CLK(clk), .RST(rst), .Q(ereg[136]) );
  DFF \ereg_reg[137]  ( .D(n3721), .CLK(clk), .RST(rst), .Q(ereg[137]) );
  DFF \ereg_reg[138]  ( .D(n3720), .CLK(clk), .RST(rst), .Q(ereg[138]) );
  DFF \ereg_reg[139]  ( .D(n3719), .CLK(clk), .RST(rst), .Q(ereg[139]) );
  DFF \ereg_reg[140]  ( .D(n3718), .CLK(clk), .RST(rst), .Q(ereg[140]) );
  DFF \ereg_reg[141]  ( .D(n3717), .CLK(clk), .RST(rst), .Q(ereg[141]) );
  DFF \ereg_reg[142]  ( .D(n3716), .CLK(clk), .RST(rst), .Q(ereg[142]) );
  DFF \ereg_reg[143]  ( .D(n3715), .CLK(clk), .RST(rst), .Q(ereg[143]) );
  DFF \ereg_reg[144]  ( .D(n3714), .CLK(clk), .RST(rst), .Q(ereg[144]) );
  DFF \ereg_reg[145]  ( .D(n3713), .CLK(clk), .RST(rst), .Q(ereg[145]) );
  DFF \ereg_reg[146]  ( .D(n3712), .CLK(clk), .RST(rst), .Q(ereg[146]) );
  DFF \ereg_reg[147]  ( .D(n3711), .CLK(clk), .RST(rst), .Q(ereg[147]) );
  DFF \ereg_reg[148]  ( .D(n3710), .CLK(clk), .RST(rst), .Q(ereg[148]) );
  DFF \ereg_reg[149]  ( .D(n3709), .CLK(clk), .RST(rst), .Q(ereg[149]) );
  DFF \ereg_reg[150]  ( .D(n3708), .CLK(clk), .RST(rst), .Q(ereg[150]) );
  DFF \ereg_reg[151]  ( .D(n3707), .CLK(clk), .RST(rst), .Q(ereg[151]) );
  DFF \ereg_reg[152]  ( .D(n3706), .CLK(clk), .RST(rst), .Q(ereg[152]) );
  DFF \ereg_reg[153]  ( .D(n3705), .CLK(clk), .RST(rst), .Q(ereg[153]) );
  DFF \ereg_reg[154]  ( .D(n3704), .CLK(clk), .RST(rst), .Q(ereg[154]) );
  DFF \ereg_reg[155]  ( .D(n3703), .CLK(clk), .RST(rst), .Q(ereg[155]) );
  DFF \ereg_reg[156]  ( .D(n3702), .CLK(clk), .RST(rst), .Q(ereg[156]) );
  DFF \ereg_reg[157]  ( .D(n3701), .CLK(clk), .RST(rst), .Q(ereg[157]) );
  DFF \ereg_reg[158]  ( .D(n3700), .CLK(clk), .RST(rst), .Q(ereg[158]) );
  DFF \ereg_reg[159]  ( .D(n3699), .CLK(clk), .RST(rst), .Q(ereg[159]) );
  DFF \ereg_reg[160]  ( .D(n3698), .CLK(clk), .RST(rst), .Q(ereg[160]) );
  DFF \ereg_reg[161]  ( .D(n3697), .CLK(clk), .RST(rst), .Q(ereg[161]) );
  DFF \ereg_reg[162]  ( .D(n3696), .CLK(clk), .RST(rst), .Q(ereg[162]) );
  DFF \ereg_reg[163]  ( .D(n3695), .CLK(clk), .RST(rst), .Q(ereg[163]) );
  DFF \ereg_reg[164]  ( .D(n3694), .CLK(clk), .RST(rst), .Q(ereg[164]) );
  DFF \ereg_reg[165]  ( .D(n3693), .CLK(clk), .RST(rst), .Q(ereg[165]) );
  DFF \ereg_reg[166]  ( .D(n3692), .CLK(clk), .RST(rst), .Q(ereg[166]) );
  DFF \ereg_reg[167]  ( .D(n3691), .CLK(clk), .RST(rst), .Q(ereg[167]) );
  DFF \ereg_reg[168]  ( .D(n3690), .CLK(clk), .RST(rst), .Q(ereg[168]) );
  DFF \ereg_reg[169]  ( .D(n3689), .CLK(clk), .RST(rst), .Q(ereg[169]) );
  DFF \ereg_reg[170]  ( .D(n3688), .CLK(clk), .RST(rst), .Q(ereg[170]) );
  DFF \ereg_reg[171]  ( .D(n3687), .CLK(clk), .RST(rst), .Q(ereg[171]) );
  DFF \ereg_reg[172]  ( .D(n3686), .CLK(clk), .RST(rst), .Q(ereg[172]) );
  DFF \ereg_reg[173]  ( .D(n3685), .CLK(clk), .RST(rst), .Q(ereg[173]) );
  DFF \ereg_reg[174]  ( .D(n3684), .CLK(clk), .RST(rst), .Q(ereg[174]) );
  DFF \ereg_reg[175]  ( .D(n3683), .CLK(clk), .RST(rst), .Q(ereg[175]) );
  DFF \ereg_reg[176]  ( .D(n3682), .CLK(clk), .RST(rst), .Q(ereg[176]) );
  DFF \ereg_reg[177]  ( .D(n3681), .CLK(clk), .RST(rst), .Q(ereg[177]) );
  DFF \ereg_reg[178]  ( .D(n3680), .CLK(clk), .RST(rst), .Q(ereg[178]) );
  DFF \ereg_reg[179]  ( .D(n3679), .CLK(clk), .RST(rst), .Q(ereg[179]) );
  DFF \ereg_reg[180]  ( .D(n3678), .CLK(clk), .RST(rst), .Q(ereg[180]) );
  DFF \ereg_reg[181]  ( .D(n3677), .CLK(clk), .RST(rst), .Q(ereg[181]) );
  DFF \ereg_reg[182]  ( .D(n3676), .CLK(clk), .RST(rst), .Q(ereg[182]) );
  DFF \ereg_reg[183]  ( .D(n3675), .CLK(clk), .RST(rst), .Q(ereg[183]) );
  DFF \ereg_reg[184]  ( .D(n3674), .CLK(clk), .RST(rst), .Q(ereg[184]) );
  DFF \ereg_reg[185]  ( .D(n3673), .CLK(clk), .RST(rst), .Q(ereg[185]) );
  DFF \ereg_reg[186]  ( .D(n3672), .CLK(clk), .RST(rst), .Q(ereg[186]) );
  DFF \ereg_reg[187]  ( .D(n3671), .CLK(clk), .RST(rst), .Q(ereg[187]) );
  DFF \ereg_reg[188]  ( .D(n3670), .CLK(clk), .RST(rst), .Q(ereg[188]) );
  DFF \ereg_reg[189]  ( .D(n3669), .CLK(clk), .RST(rst), .Q(ereg[189]) );
  DFF \ereg_reg[190]  ( .D(n3668), .CLK(clk), .RST(rst), .Q(ereg[190]) );
  DFF \ereg_reg[191]  ( .D(n3667), .CLK(clk), .RST(rst), .Q(ereg[191]) );
  DFF \ereg_reg[192]  ( .D(n3666), .CLK(clk), .RST(rst), .Q(ereg[192]) );
  DFF \ereg_reg[193]  ( .D(n3665), .CLK(clk), .RST(rst), .Q(ereg[193]) );
  DFF \ereg_reg[194]  ( .D(n3664), .CLK(clk), .RST(rst), .Q(ereg[194]) );
  DFF \ereg_reg[195]  ( .D(n3663), .CLK(clk), .RST(rst), .Q(ereg[195]) );
  DFF \ereg_reg[196]  ( .D(n3662), .CLK(clk), .RST(rst), .Q(ereg[196]) );
  DFF \ereg_reg[197]  ( .D(n3661), .CLK(clk), .RST(rst), .Q(ereg[197]) );
  DFF \ereg_reg[198]  ( .D(n3660), .CLK(clk), .RST(rst), .Q(ereg[198]) );
  DFF \ereg_reg[199]  ( .D(n3659), .CLK(clk), .RST(rst), .Q(ereg[199]) );
  DFF \ereg_reg[200]  ( .D(n3658), .CLK(clk), .RST(rst), .Q(ereg[200]) );
  DFF \ereg_reg[201]  ( .D(n3657), .CLK(clk), .RST(rst), .Q(ereg[201]) );
  DFF \ereg_reg[202]  ( .D(n3656), .CLK(clk), .RST(rst), .Q(ereg[202]) );
  DFF \ereg_reg[203]  ( .D(n3655), .CLK(clk), .RST(rst), .Q(ereg[203]) );
  DFF \ereg_reg[204]  ( .D(n3654), .CLK(clk), .RST(rst), .Q(ereg[204]) );
  DFF \ereg_reg[205]  ( .D(n3653), .CLK(clk), .RST(rst), .Q(ereg[205]) );
  DFF \ereg_reg[206]  ( .D(n3652), .CLK(clk), .RST(rst), .Q(ereg[206]) );
  DFF \ereg_reg[207]  ( .D(n3651), .CLK(clk), .RST(rst), .Q(ereg[207]) );
  DFF \ereg_reg[208]  ( .D(n3650), .CLK(clk), .RST(rst), .Q(ereg[208]) );
  DFF \ereg_reg[209]  ( .D(n3649), .CLK(clk), .RST(rst), .Q(ereg[209]) );
  DFF \ereg_reg[210]  ( .D(n3648), .CLK(clk), .RST(rst), .Q(ereg[210]) );
  DFF \ereg_reg[211]  ( .D(n3647), .CLK(clk), .RST(rst), .Q(ereg[211]) );
  DFF \ereg_reg[212]  ( .D(n3646), .CLK(clk), .RST(rst), .Q(ereg[212]) );
  DFF \ereg_reg[213]  ( .D(n3645), .CLK(clk), .RST(rst), .Q(ereg[213]) );
  DFF \ereg_reg[214]  ( .D(n3644), .CLK(clk), .RST(rst), .Q(ereg[214]) );
  DFF \ereg_reg[215]  ( .D(n3643), .CLK(clk), .RST(rst), .Q(ereg[215]) );
  DFF \ereg_reg[216]  ( .D(n3642), .CLK(clk), .RST(rst), .Q(ereg[216]) );
  DFF \ereg_reg[217]  ( .D(n3641), .CLK(clk), .RST(rst), .Q(ereg[217]) );
  DFF \ereg_reg[218]  ( .D(n3640), .CLK(clk), .RST(rst), .Q(ereg[218]) );
  DFF \ereg_reg[219]  ( .D(n3639), .CLK(clk), .RST(rst), .Q(ereg[219]) );
  DFF \ereg_reg[220]  ( .D(n3638), .CLK(clk), .RST(rst), .Q(ereg[220]) );
  DFF \ereg_reg[221]  ( .D(n3637), .CLK(clk), .RST(rst), .Q(ereg[221]) );
  DFF \ereg_reg[222]  ( .D(n3636), .CLK(clk), .RST(rst), .Q(ereg[222]) );
  DFF \ereg_reg[223]  ( .D(n3635), .CLK(clk), .RST(rst), .Q(ereg[223]) );
  DFF \ereg_reg[224]  ( .D(n3634), .CLK(clk), .RST(rst), .Q(ereg[224]) );
  DFF \ereg_reg[225]  ( .D(n3633), .CLK(clk), .RST(rst), .Q(ereg[225]) );
  DFF \ereg_reg[226]  ( .D(n3632), .CLK(clk), .RST(rst), .Q(ereg[226]) );
  DFF \ereg_reg[227]  ( .D(n3631), .CLK(clk), .RST(rst), .Q(ereg[227]) );
  DFF \ereg_reg[228]  ( .D(n3630), .CLK(clk), .RST(rst), .Q(ereg[228]) );
  DFF \ereg_reg[229]  ( .D(n3629), .CLK(clk), .RST(rst), .Q(ereg[229]) );
  DFF \ereg_reg[230]  ( .D(n3628), .CLK(clk), .RST(rst), .Q(ereg[230]) );
  DFF \ereg_reg[231]  ( .D(n3627), .CLK(clk), .RST(rst), .Q(ereg[231]) );
  DFF \ereg_reg[232]  ( .D(n3626), .CLK(clk), .RST(rst), .Q(ereg[232]) );
  DFF \ereg_reg[233]  ( .D(n3625), .CLK(clk), .RST(rst), .Q(ereg[233]) );
  DFF \ereg_reg[234]  ( .D(n3624), .CLK(clk), .RST(rst), .Q(ereg[234]) );
  DFF \ereg_reg[235]  ( .D(n3623), .CLK(clk), .RST(rst), .Q(ereg[235]) );
  DFF \ereg_reg[236]  ( .D(n3622), .CLK(clk), .RST(rst), .Q(ereg[236]) );
  DFF \ereg_reg[237]  ( .D(n3621), .CLK(clk), .RST(rst), .Q(ereg[237]) );
  DFF \ereg_reg[238]  ( .D(n3620), .CLK(clk), .RST(rst), .Q(ereg[238]) );
  DFF \ereg_reg[239]  ( .D(n3619), .CLK(clk), .RST(rst), .Q(ereg[239]) );
  DFF \ereg_reg[240]  ( .D(n3618), .CLK(clk), .RST(rst), .Q(ereg[240]) );
  DFF \ereg_reg[241]  ( .D(n3617), .CLK(clk), .RST(rst), .Q(ereg[241]) );
  DFF \ereg_reg[242]  ( .D(n3616), .CLK(clk), .RST(rst), .Q(ereg[242]) );
  DFF \ereg_reg[243]  ( .D(n3615), .CLK(clk), .RST(rst), .Q(ereg[243]) );
  DFF \ereg_reg[244]  ( .D(n3614), .CLK(clk), .RST(rst), .Q(ereg[244]) );
  DFF \ereg_reg[245]  ( .D(n3613), .CLK(clk), .RST(rst), .Q(ereg[245]) );
  DFF \ereg_reg[246]  ( .D(n3612), .CLK(clk), .RST(rst), .Q(ereg[246]) );
  DFF \ereg_reg[247]  ( .D(n3611), .CLK(clk), .RST(rst), .Q(ereg[247]) );
  DFF \ereg_reg[248]  ( .D(n3610), .CLK(clk), .RST(rst), .Q(ereg[248]) );
  DFF \ereg_reg[249]  ( .D(n3609), .CLK(clk), .RST(rst), .Q(ereg[249]) );
  DFF \ereg_reg[250]  ( .D(n3608), .CLK(clk), .RST(rst), .Q(ereg[250]) );
  DFF \ereg_reg[251]  ( .D(n3607), .CLK(clk), .RST(rst), .Q(ereg[251]) );
  DFF \ereg_reg[252]  ( .D(n3606), .CLK(clk), .RST(rst), .Q(ereg[252]) );
  DFF \ereg_reg[253]  ( .D(n3605), .CLK(clk), .RST(rst), .Q(ereg[253]) );
  DFF \ereg_reg[254]  ( .D(n3604), .CLK(clk), .RST(rst), .Q(ereg[254]) );
  DFF \ereg_reg[255]  ( .D(n3603), .CLK(clk), .RST(rst), .Q(ereg[255]) );
  DFF first_one_reg ( .D(n3346), .CLK(clk), .RST(rst), .Q(first_one) );
  DFF \creg_reg[0]  ( .D(n3601), .CLK(clk), .RST(rst), .Q(creg[0]) );
  DFF \creg_reg[1]  ( .D(n3600), .CLK(clk), .RST(rst), .Q(creg[1]) );
  DFF \creg_reg[2]  ( .D(n3599), .CLK(clk), .RST(rst), .Q(creg[2]) );
  DFF \creg_reg[3]  ( .D(n3598), .CLK(clk), .RST(rst), .Q(creg[3]) );
  DFF \creg_reg[4]  ( .D(n3597), .CLK(clk), .RST(rst), .Q(creg[4]) );
  DFF \creg_reg[5]  ( .D(n3596), .CLK(clk), .RST(rst), .Q(creg[5]) );
  DFF \creg_reg[6]  ( .D(n3595), .CLK(clk), .RST(rst), .Q(creg[6]) );
  DFF \creg_reg[7]  ( .D(n3594), .CLK(clk), .RST(rst), .Q(creg[7]) );
  DFF \creg_reg[8]  ( .D(n3593), .CLK(clk), .RST(rst), .Q(creg[8]) );
  DFF \creg_reg[9]  ( .D(n3592), .CLK(clk), .RST(rst), .Q(creg[9]) );
  DFF \creg_reg[10]  ( .D(n3591), .CLK(clk), .RST(rst), .Q(creg[10]) );
  DFF \creg_reg[11]  ( .D(n3590), .CLK(clk), .RST(rst), .Q(creg[11]) );
  DFF \creg_reg[12]  ( .D(n3589), .CLK(clk), .RST(rst), .Q(creg[12]) );
  DFF \creg_reg[13]  ( .D(n3588), .CLK(clk), .RST(rst), .Q(creg[13]) );
  DFF \creg_reg[14]  ( .D(n3587), .CLK(clk), .RST(rst), .Q(creg[14]) );
  DFF \creg_reg[15]  ( .D(n3586), .CLK(clk), .RST(rst), .Q(creg[15]) );
  DFF \creg_reg[16]  ( .D(n3585), .CLK(clk), .RST(rst), .Q(creg[16]) );
  DFF \creg_reg[17]  ( .D(n3584), .CLK(clk), .RST(rst), .Q(creg[17]) );
  DFF \creg_reg[18]  ( .D(n3583), .CLK(clk), .RST(rst), .Q(creg[18]) );
  DFF \creg_reg[19]  ( .D(n3582), .CLK(clk), .RST(rst), .Q(creg[19]) );
  DFF \creg_reg[20]  ( .D(n3581), .CLK(clk), .RST(rst), .Q(creg[20]) );
  DFF \creg_reg[21]  ( .D(n3580), .CLK(clk), .RST(rst), .Q(creg[21]) );
  DFF \creg_reg[22]  ( .D(n3579), .CLK(clk), .RST(rst), .Q(creg[22]) );
  DFF \creg_reg[23]  ( .D(n3578), .CLK(clk), .RST(rst), .Q(creg[23]) );
  DFF \creg_reg[24]  ( .D(n3577), .CLK(clk), .RST(rst), .Q(creg[24]) );
  DFF \creg_reg[25]  ( .D(n3576), .CLK(clk), .RST(rst), .Q(creg[25]) );
  DFF \creg_reg[26]  ( .D(n3575), .CLK(clk), .RST(rst), .Q(creg[26]) );
  DFF \creg_reg[27]  ( .D(n3574), .CLK(clk), .RST(rst), .Q(creg[27]) );
  DFF \creg_reg[28]  ( .D(n3573), .CLK(clk), .RST(rst), .Q(creg[28]) );
  DFF \creg_reg[29]  ( .D(n3572), .CLK(clk), .RST(rst), .Q(creg[29]) );
  DFF \creg_reg[30]  ( .D(n3571), .CLK(clk), .RST(rst), .Q(creg[30]) );
  DFF \creg_reg[31]  ( .D(n3570), .CLK(clk), .RST(rst), .Q(creg[31]) );
  DFF \creg_reg[32]  ( .D(n3569), .CLK(clk), .RST(rst), .Q(creg[32]) );
  DFF \creg_reg[33]  ( .D(n3568), .CLK(clk), .RST(rst), .Q(creg[33]) );
  DFF \creg_reg[34]  ( .D(n3567), .CLK(clk), .RST(rst), .Q(creg[34]) );
  DFF \creg_reg[35]  ( .D(n3566), .CLK(clk), .RST(rst), .Q(creg[35]) );
  DFF \creg_reg[36]  ( .D(n3565), .CLK(clk), .RST(rst), .Q(creg[36]) );
  DFF \creg_reg[37]  ( .D(n3564), .CLK(clk), .RST(rst), .Q(creg[37]) );
  DFF \creg_reg[38]  ( .D(n3563), .CLK(clk), .RST(rst), .Q(creg[38]) );
  DFF \creg_reg[39]  ( .D(n3562), .CLK(clk), .RST(rst), .Q(creg[39]) );
  DFF \creg_reg[40]  ( .D(n3561), .CLK(clk), .RST(rst), .Q(creg[40]) );
  DFF \creg_reg[41]  ( .D(n3560), .CLK(clk), .RST(rst), .Q(creg[41]) );
  DFF \creg_reg[42]  ( .D(n3559), .CLK(clk), .RST(rst), .Q(creg[42]) );
  DFF \creg_reg[43]  ( .D(n3558), .CLK(clk), .RST(rst), .Q(creg[43]) );
  DFF \creg_reg[44]  ( .D(n3557), .CLK(clk), .RST(rst), .Q(creg[44]) );
  DFF \creg_reg[45]  ( .D(n3556), .CLK(clk), .RST(rst), .Q(creg[45]) );
  DFF \creg_reg[46]  ( .D(n3555), .CLK(clk), .RST(rst), .Q(creg[46]) );
  DFF \creg_reg[47]  ( .D(n3554), .CLK(clk), .RST(rst), .Q(creg[47]) );
  DFF \creg_reg[48]  ( .D(n3553), .CLK(clk), .RST(rst), .Q(creg[48]) );
  DFF \creg_reg[49]  ( .D(n3552), .CLK(clk), .RST(rst), .Q(creg[49]) );
  DFF \creg_reg[50]  ( .D(n3551), .CLK(clk), .RST(rst), .Q(creg[50]) );
  DFF \creg_reg[51]  ( .D(n3550), .CLK(clk), .RST(rst), .Q(creg[51]) );
  DFF \creg_reg[52]  ( .D(n3549), .CLK(clk), .RST(rst), .Q(creg[52]) );
  DFF \creg_reg[53]  ( .D(n3548), .CLK(clk), .RST(rst), .Q(creg[53]) );
  DFF \creg_reg[54]  ( .D(n3547), .CLK(clk), .RST(rst), .Q(creg[54]) );
  DFF \creg_reg[55]  ( .D(n3546), .CLK(clk), .RST(rst), .Q(creg[55]) );
  DFF \creg_reg[56]  ( .D(n3545), .CLK(clk), .RST(rst), .Q(creg[56]) );
  DFF \creg_reg[57]  ( .D(n3544), .CLK(clk), .RST(rst), .Q(creg[57]) );
  DFF \creg_reg[58]  ( .D(n3543), .CLK(clk), .RST(rst), .Q(creg[58]) );
  DFF \creg_reg[59]  ( .D(n3542), .CLK(clk), .RST(rst), .Q(creg[59]) );
  DFF \creg_reg[60]  ( .D(n3541), .CLK(clk), .RST(rst), .Q(creg[60]) );
  DFF \creg_reg[61]  ( .D(n3540), .CLK(clk), .RST(rst), .Q(creg[61]) );
  DFF \creg_reg[62]  ( .D(n3539), .CLK(clk), .RST(rst), .Q(creg[62]) );
  DFF \creg_reg[63]  ( .D(n3538), .CLK(clk), .RST(rst), .Q(creg[63]) );
  DFF \creg_reg[64]  ( .D(n3537), .CLK(clk), .RST(rst), .Q(creg[64]) );
  DFF \creg_reg[65]  ( .D(n3536), .CLK(clk), .RST(rst), .Q(creg[65]) );
  DFF \creg_reg[66]  ( .D(n3535), .CLK(clk), .RST(rst), .Q(creg[66]) );
  DFF \creg_reg[67]  ( .D(n3534), .CLK(clk), .RST(rst), .Q(creg[67]) );
  DFF \creg_reg[68]  ( .D(n3533), .CLK(clk), .RST(rst), .Q(creg[68]) );
  DFF \creg_reg[69]  ( .D(n3532), .CLK(clk), .RST(rst), .Q(creg[69]) );
  DFF \creg_reg[70]  ( .D(n3531), .CLK(clk), .RST(rst), .Q(creg[70]) );
  DFF \creg_reg[71]  ( .D(n3530), .CLK(clk), .RST(rst), .Q(creg[71]) );
  DFF \creg_reg[72]  ( .D(n3529), .CLK(clk), .RST(rst), .Q(creg[72]) );
  DFF \creg_reg[73]  ( .D(n3528), .CLK(clk), .RST(rst), .Q(creg[73]) );
  DFF \creg_reg[74]  ( .D(n3527), .CLK(clk), .RST(rst), .Q(creg[74]) );
  DFF \creg_reg[75]  ( .D(n3526), .CLK(clk), .RST(rst), .Q(creg[75]) );
  DFF \creg_reg[76]  ( .D(n3525), .CLK(clk), .RST(rst), .Q(creg[76]) );
  DFF \creg_reg[77]  ( .D(n3524), .CLK(clk), .RST(rst), .Q(creg[77]) );
  DFF \creg_reg[78]  ( .D(n3523), .CLK(clk), .RST(rst), .Q(creg[78]) );
  DFF \creg_reg[79]  ( .D(n3522), .CLK(clk), .RST(rst), .Q(creg[79]) );
  DFF \creg_reg[80]  ( .D(n3521), .CLK(clk), .RST(rst), .Q(creg[80]) );
  DFF \creg_reg[81]  ( .D(n3520), .CLK(clk), .RST(rst), .Q(creg[81]) );
  DFF \creg_reg[82]  ( .D(n3519), .CLK(clk), .RST(rst), .Q(creg[82]) );
  DFF \creg_reg[83]  ( .D(n3518), .CLK(clk), .RST(rst), .Q(creg[83]) );
  DFF \creg_reg[84]  ( .D(n3517), .CLK(clk), .RST(rst), .Q(creg[84]) );
  DFF \creg_reg[85]  ( .D(n3516), .CLK(clk), .RST(rst), .Q(creg[85]) );
  DFF \creg_reg[86]  ( .D(n3515), .CLK(clk), .RST(rst), .Q(creg[86]) );
  DFF \creg_reg[87]  ( .D(n3514), .CLK(clk), .RST(rst), .Q(creg[87]) );
  DFF \creg_reg[88]  ( .D(n3513), .CLK(clk), .RST(rst), .Q(creg[88]) );
  DFF \creg_reg[89]  ( .D(n3512), .CLK(clk), .RST(rst), .Q(creg[89]) );
  DFF \creg_reg[90]  ( .D(n3511), .CLK(clk), .RST(rst), .Q(creg[90]) );
  DFF \creg_reg[91]  ( .D(n3510), .CLK(clk), .RST(rst), .Q(creg[91]) );
  DFF \creg_reg[92]  ( .D(n3509), .CLK(clk), .RST(rst), .Q(creg[92]) );
  DFF \creg_reg[93]  ( .D(n3508), .CLK(clk), .RST(rst), .Q(creg[93]) );
  DFF \creg_reg[94]  ( .D(n3507), .CLK(clk), .RST(rst), .Q(creg[94]) );
  DFF \creg_reg[95]  ( .D(n3506), .CLK(clk), .RST(rst), .Q(creg[95]) );
  DFF \creg_reg[96]  ( .D(n3505), .CLK(clk), .RST(rst), .Q(creg[96]) );
  DFF \creg_reg[97]  ( .D(n3504), .CLK(clk), .RST(rst), .Q(creg[97]) );
  DFF \creg_reg[98]  ( .D(n3503), .CLK(clk), .RST(rst), .Q(creg[98]) );
  DFF \creg_reg[99]  ( .D(n3502), .CLK(clk), .RST(rst), .Q(creg[99]) );
  DFF \creg_reg[100]  ( .D(n3501), .CLK(clk), .RST(rst), .Q(creg[100]) );
  DFF \creg_reg[101]  ( .D(n3500), .CLK(clk), .RST(rst), .Q(creg[101]) );
  DFF \creg_reg[102]  ( .D(n3499), .CLK(clk), .RST(rst), .Q(creg[102]) );
  DFF \creg_reg[103]  ( .D(n3498), .CLK(clk), .RST(rst), .Q(creg[103]) );
  DFF \creg_reg[104]  ( .D(n3497), .CLK(clk), .RST(rst), .Q(creg[104]) );
  DFF \creg_reg[105]  ( .D(n3496), .CLK(clk), .RST(rst), .Q(creg[105]) );
  DFF \creg_reg[106]  ( .D(n3495), .CLK(clk), .RST(rst), .Q(creg[106]) );
  DFF \creg_reg[107]  ( .D(n3494), .CLK(clk), .RST(rst), .Q(creg[107]) );
  DFF \creg_reg[108]  ( .D(n3493), .CLK(clk), .RST(rst), .Q(creg[108]) );
  DFF \creg_reg[109]  ( .D(n3492), .CLK(clk), .RST(rst), .Q(creg[109]) );
  DFF \creg_reg[110]  ( .D(n3491), .CLK(clk), .RST(rst), .Q(creg[110]) );
  DFF \creg_reg[111]  ( .D(n3490), .CLK(clk), .RST(rst), .Q(creg[111]) );
  DFF \creg_reg[112]  ( .D(n3489), .CLK(clk), .RST(rst), .Q(creg[112]) );
  DFF \creg_reg[113]  ( .D(n3488), .CLK(clk), .RST(rst), .Q(creg[113]) );
  DFF \creg_reg[114]  ( .D(n3487), .CLK(clk), .RST(rst), .Q(creg[114]) );
  DFF \creg_reg[115]  ( .D(n3486), .CLK(clk), .RST(rst), .Q(creg[115]) );
  DFF \creg_reg[116]  ( .D(n3485), .CLK(clk), .RST(rst), .Q(creg[116]) );
  DFF \creg_reg[117]  ( .D(n3484), .CLK(clk), .RST(rst), .Q(creg[117]) );
  DFF \creg_reg[118]  ( .D(n3483), .CLK(clk), .RST(rst), .Q(creg[118]) );
  DFF \creg_reg[119]  ( .D(n3482), .CLK(clk), .RST(rst), .Q(creg[119]) );
  DFF \creg_reg[120]  ( .D(n3481), .CLK(clk), .RST(rst), .Q(creg[120]) );
  DFF \creg_reg[121]  ( .D(n3480), .CLK(clk), .RST(rst), .Q(creg[121]) );
  DFF \creg_reg[122]  ( .D(n3479), .CLK(clk), .RST(rst), .Q(creg[122]) );
  DFF \creg_reg[123]  ( .D(n3478), .CLK(clk), .RST(rst), .Q(creg[123]) );
  DFF \creg_reg[124]  ( .D(n3477), .CLK(clk), .RST(rst), .Q(creg[124]) );
  DFF \creg_reg[125]  ( .D(n3476), .CLK(clk), .RST(rst), .Q(creg[125]) );
  DFF \creg_reg[126]  ( .D(n3475), .CLK(clk), .RST(rst), .Q(creg[126]) );
  DFF \creg_reg[127]  ( .D(n3474), .CLK(clk), .RST(rst), .Q(creg[127]) );
  DFF \creg_reg[128]  ( .D(n3473), .CLK(clk), .RST(rst), .Q(creg[128]) );
  DFF \creg_reg[129]  ( .D(n3472), .CLK(clk), .RST(rst), .Q(creg[129]) );
  DFF \creg_reg[130]  ( .D(n3471), .CLK(clk), .RST(rst), .Q(creg[130]) );
  DFF \creg_reg[131]  ( .D(n3470), .CLK(clk), .RST(rst), .Q(creg[131]) );
  DFF \creg_reg[132]  ( .D(n3469), .CLK(clk), .RST(rst), .Q(creg[132]) );
  DFF \creg_reg[133]  ( .D(n3468), .CLK(clk), .RST(rst), .Q(creg[133]) );
  DFF \creg_reg[134]  ( .D(n3467), .CLK(clk), .RST(rst), .Q(creg[134]) );
  DFF \creg_reg[135]  ( .D(n3466), .CLK(clk), .RST(rst), .Q(creg[135]) );
  DFF \creg_reg[136]  ( .D(n3465), .CLK(clk), .RST(rst), .Q(creg[136]) );
  DFF \creg_reg[137]  ( .D(n3464), .CLK(clk), .RST(rst), .Q(creg[137]) );
  DFF \creg_reg[138]  ( .D(n3463), .CLK(clk), .RST(rst), .Q(creg[138]) );
  DFF \creg_reg[139]  ( .D(n3462), .CLK(clk), .RST(rst), .Q(creg[139]) );
  DFF \creg_reg[140]  ( .D(n3461), .CLK(clk), .RST(rst), .Q(creg[140]) );
  DFF \creg_reg[141]  ( .D(n3460), .CLK(clk), .RST(rst), .Q(creg[141]) );
  DFF \creg_reg[142]  ( .D(n3459), .CLK(clk), .RST(rst), .Q(creg[142]) );
  DFF \creg_reg[143]  ( .D(n3458), .CLK(clk), .RST(rst), .Q(creg[143]) );
  DFF \creg_reg[144]  ( .D(n3457), .CLK(clk), .RST(rst), .Q(creg[144]) );
  DFF \creg_reg[145]  ( .D(n3456), .CLK(clk), .RST(rst), .Q(creg[145]) );
  DFF \creg_reg[146]  ( .D(n3455), .CLK(clk), .RST(rst), .Q(creg[146]) );
  DFF \creg_reg[147]  ( .D(n3454), .CLK(clk), .RST(rst), .Q(creg[147]) );
  DFF \creg_reg[148]  ( .D(n3453), .CLK(clk), .RST(rst), .Q(creg[148]) );
  DFF \creg_reg[149]  ( .D(n3452), .CLK(clk), .RST(rst), .Q(creg[149]) );
  DFF \creg_reg[150]  ( .D(n3451), .CLK(clk), .RST(rst), .Q(creg[150]) );
  DFF \creg_reg[151]  ( .D(n3450), .CLK(clk), .RST(rst), .Q(creg[151]) );
  DFF \creg_reg[152]  ( .D(n3449), .CLK(clk), .RST(rst), .Q(creg[152]) );
  DFF \creg_reg[153]  ( .D(n3448), .CLK(clk), .RST(rst), .Q(creg[153]) );
  DFF \creg_reg[154]  ( .D(n3447), .CLK(clk), .RST(rst), .Q(creg[154]) );
  DFF \creg_reg[155]  ( .D(n3446), .CLK(clk), .RST(rst), .Q(creg[155]) );
  DFF \creg_reg[156]  ( .D(n3445), .CLK(clk), .RST(rst), .Q(creg[156]) );
  DFF \creg_reg[157]  ( .D(n3444), .CLK(clk), .RST(rst), .Q(creg[157]) );
  DFF \creg_reg[158]  ( .D(n3443), .CLK(clk), .RST(rst), .Q(creg[158]) );
  DFF \creg_reg[159]  ( .D(n3442), .CLK(clk), .RST(rst), .Q(creg[159]) );
  DFF \creg_reg[160]  ( .D(n3441), .CLK(clk), .RST(rst), .Q(creg[160]) );
  DFF \creg_reg[161]  ( .D(n3440), .CLK(clk), .RST(rst), .Q(creg[161]) );
  DFF \creg_reg[162]  ( .D(n3439), .CLK(clk), .RST(rst), .Q(creg[162]) );
  DFF \creg_reg[163]  ( .D(n3438), .CLK(clk), .RST(rst), .Q(creg[163]) );
  DFF \creg_reg[164]  ( .D(n3437), .CLK(clk), .RST(rst), .Q(creg[164]) );
  DFF \creg_reg[165]  ( .D(n3436), .CLK(clk), .RST(rst), .Q(creg[165]) );
  DFF \creg_reg[166]  ( .D(n3435), .CLK(clk), .RST(rst), .Q(creg[166]) );
  DFF \creg_reg[167]  ( .D(n3434), .CLK(clk), .RST(rst), .Q(creg[167]) );
  DFF \creg_reg[168]  ( .D(n3433), .CLK(clk), .RST(rst), .Q(creg[168]) );
  DFF \creg_reg[169]  ( .D(n3432), .CLK(clk), .RST(rst), .Q(creg[169]) );
  DFF \creg_reg[170]  ( .D(n3431), .CLK(clk), .RST(rst), .Q(creg[170]) );
  DFF \creg_reg[171]  ( .D(n3430), .CLK(clk), .RST(rst), .Q(creg[171]) );
  DFF \creg_reg[172]  ( .D(n3429), .CLK(clk), .RST(rst), .Q(creg[172]) );
  DFF \creg_reg[173]  ( .D(n3428), .CLK(clk), .RST(rst), .Q(creg[173]) );
  DFF \creg_reg[174]  ( .D(n3427), .CLK(clk), .RST(rst), .Q(creg[174]) );
  DFF \creg_reg[175]  ( .D(n3426), .CLK(clk), .RST(rst), .Q(creg[175]) );
  DFF \creg_reg[176]  ( .D(n3425), .CLK(clk), .RST(rst), .Q(creg[176]) );
  DFF \creg_reg[177]  ( .D(n3424), .CLK(clk), .RST(rst), .Q(creg[177]) );
  DFF \creg_reg[178]  ( .D(n3423), .CLK(clk), .RST(rst), .Q(creg[178]) );
  DFF \creg_reg[179]  ( .D(n3422), .CLK(clk), .RST(rst), .Q(creg[179]) );
  DFF \creg_reg[180]  ( .D(n3421), .CLK(clk), .RST(rst), .Q(creg[180]) );
  DFF \creg_reg[181]  ( .D(n3420), .CLK(clk), .RST(rst), .Q(creg[181]) );
  DFF \creg_reg[182]  ( .D(n3419), .CLK(clk), .RST(rst), .Q(creg[182]) );
  DFF \creg_reg[183]  ( .D(n3418), .CLK(clk), .RST(rst), .Q(creg[183]) );
  DFF \creg_reg[184]  ( .D(n3417), .CLK(clk), .RST(rst), .Q(creg[184]) );
  DFF \creg_reg[185]  ( .D(n3416), .CLK(clk), .RST(rst), .Q(creg[185]) );
  DFF \creg_reg[186]  ( .D(n3415), .CLK(clk), .RST(rst), .Q(creg[186]) );
  DFF \creg_reg[187]  ( .D(n3414), .CLK(clk), .RST(rst), .Q(creg[187]) );
  DFF \creg_reg[188]  ( .D(n3413), .CLK(clk), .RST(rst), .Q(creg[188]) );
  DFF \creg_reg[189]  ( .D(n3412), .CLK(clk), .RST(rst), .Q(creg[189]) );
  DFF \creg_reg[190]  ( .D(n3411), .CLK(clk), .RST(rst), .Q(creg[190]) );
  DFF \creg_reg[191]  ( .D(n3410), .CLK(clk), .RST(rst), .Q(creg[191]) );
  DFF \creg_reg[192]  ( .D(n3409), .CLK(clk), .RST(rst), .Q(creg[192]) );
  DFF \creg_reg[193]  ( .D(n3408), .CLK(clk), .RST(rst), .Q(creg[193]) );
  DFF \creg_reg[194]  ( .D(n3407), .CLK(clk), .RST(rst), .Q(creg[194]) );
  DFF \creg_reg[195]  ( .D(n3406), .CLK(clk), .RST(rst), .Q(creg[195]) );
  DFF \creg_reg[196]  ( .D(n3405), .CLK(clk), .RST(rst), .Q(creg[196]) );
  DFF \creg_reg[197]  ( .D(n3404), .CLK(clk), .RST(rst), .Q(creg[197]) );
  DFF \creg_reg[198]  ( .D(n3403), .CLK(clk), .RST(rst), .Q(creg[198]) );
  DFF \creg_reg[199]  ( .D(n3402), .CLK(clk), .RST(rst), .Q(creg[199]) );
  DFF \creg_reg[200]  ( .D(n3401), .CLK(clk), .RST(rst), .Q(creg[200]) );
  DFF \creg_reg[201]  ( .D(n3400), .CLK(clk), .RST(rst), .Q(creg[201]) );
  DFF \creg_reg[202]  ( .D(n3399), .CLK(clk), .RST(rst), .Q(creg[202]) );
  DFF \creg_reg[203]  ( .D(n3398), .CLK(clk), .RST(rst), .Q(creg[203]) );
  DFF \creg_reg[204]  ( .D(n3397), .CLK(clk), .RST(rst), .Q(creg[204]) );
  DFF \creg_reg[205]  ( .D(n3396), .CLK(clk), .RST(rst), .Q(creg[205]) );
  DFF \creg_reg[206]  ( .D(n3395), .CLK(clk), .RST(rst), .Q(creg[206]) );
  DFF \creg_reg[207]  ( .D(n3394), .CLK(clk), .RST(rst), .Q(creg[207]) );
  DFF \creg_reg[208]  ( .D(n3393), .CLK(clk), .RST(rst), .Q(creg[208]) );
  DFF \creg_reg[209]  ( .D(n3392), .CLK(clk), .RST(rst), .Q(creg[209]) );
  DFF \creg_reg[210]  ( .D(n3391), .CLK(clk), .RST(rst), .Q(creg[210]) );
  DFF \creg_reg[211]  ( .D(n3390), .CLK(clk), .RST(rst), .Q(creg[211]) );
  DFF \creg_reg[212]  ( .D(n3389), .CLK(clk), .RST(rst), .Q(creg[212]) );
  DFF \creg_reg[213]  ( .D(n3388), .CLK(clk), .RST(rst), .Q(creg[213]) );
  DFF \creg_reg[214]  ( .D(n3387), .CLK(clk), .RST(rst), .Q(creg[214]) );
  DFF \creg_reg[215]  ( .D(n3386), .CLK(clk), .RST(rst), .Q(creg[215]) );
  DFF \creg_reg[216]  ( .D(n3385), .CLK(clk), .RST(rst), .Q(creg[216]) );
  DFF \creg_reg[217]  ( .D(n3384), .CLK(clk), .RST(rst), .Q(creg[217]) );
  DFF \creg_reg[218]  ( .D(n3383), .CLK(clk), .RST(rst), .Q(creg[218]) );
  DFF \creg_reg[219]  ( .D(n3382), .CLK(clk), .RST(rst), .Q(creg[219]) );
  DFF \creg_reg[220]  ( .D(n3381), .CLK(clk), .RST(rst), .Q(creg[220]) );
  DFF \creg_reg[221]  ( .D(n3380), .CLK(clk), .RST(rst), .Q(creg[221]) );
  DFF \creg_reg[222]  ( .D(n3379), .CLK(clk), .RST(rst), .Q(creg[222]) );
  DFF \creg_reg[223]  ( .D(n3378), .CLK(clk), .RST(rst), .Q(creg[223]) );
  DFF \creg_reg[224]  ( .D(n3377), .CLK(clk), .RST(rst), .Q(creg[224]) );
  DFF \creg_reg[225]  ( .D(n3376), .CLK(clk), .RST(rst), .Q(creg[225]) );
  DFF \creg_reg[226]  ( .D(n3375), .CLK(clk), .RST(rst), .Q(creg[226]) );
  DFF \creg_reg[227]  ( .D(n3374), .CLK(clk), .RST(rst), .Q(creg[227]) );
  DFF \creg_reg[228]  ( .D(n3373), .CLK(clk), .RST(rst), .Q(creg[228]) );
  DFF \creg_reg[229]  ( .D(n3372), .CLK(clk), .RST(rst), .Q(creg[229]) );
  DFF \creg_reg[230]  ( .D(n3371), .CLK(clk), .RST(rst), .Q(creg[230]) );
  DFF \creg_reg[231]  ( .D(n3370), .CLK(clk), .RST(rst), .Q(creg[231]) );
  DFF \creg_reg[232]  ( .D(n3369), .CLK(clk), .RST(rst), .Q(creg[232]) );
  DFF \creg_reg[233]  ( .D(n3368), .CLK(clk), .RST(rst), .Q(creg[233]) );
  DFF \creg_reg[234]  ( .D(n3367), .CLK(clk), .RST(rst), .Q(creg[234]) );
  DFF \creg_reg[235]  ( .D(n3366), .CLK(clk), .RST(rst), .Q(creg[235]) );
  DFF \creg_reg[236]  ( .D(n3365), .CLK(clk), .RST(rst), .Q(creg[236]) );
  DFF \creg_reg[237]  ( .D(n3364), .CLK(clk), .RST(rst), .Q(creg[237]) );
  DFF \creg_reg[238]  ( .D(n3363), .CLK(clk), .RST(rst), .Q(creg[238]) );
  DFF \creg_reg[239]  ( .D(n3362), .CLK(clk), .RST(rst), .Q(creg[239]) );
  DFF \creg_reg[240]  ( .D(n3361), .CLK(clk), .RST(rst), .Q(creg[240]) );
  DFF \creg_reg[241]  ( .D(n3360), .CLK(clk), .RST(rst), .Q(creg[241]) );
  DFF \creg_reg[242]  ( .D(n3359), .CLK(clk), .RST(rst), .Q(creg[242]) );
  DFF \creg_reg[243]  ( .D(n3358), .CLK(clk), .RST(rst), .Q(creg[243]) );
  DFF \creg_reg[244]  ( .D(n3357), .CLK(clk), .RST(rst), .Q(creg[244]) );
  DFF \creg_reg[245]  ( .D(n3356), .CLK(clk), .RST(rst), .Q(creg[245]) );
  DFF \creg_reg[246]  ( .D(n3355), .CLK(clk), .RST(rst), .Q(creg[246]) );
  DFF \creg_reg[247]  ( .D(n3354), .CLK(clk), .RST(rst), .Q(creg[247]) );
  DFF \creg_reg[248]  ( .D(n3353), .CLK(clk), .RST(rst), .Q(creg[248]) );
  DFF \creg_reg[249]  ( .D(n3352), .CLK(clk), .RST(rst), .Q(creg[249]) );
  DFF \creg_reg[250]  ( .D(n3351), .CLK(clk), .RST(rst), .Q(creg[250]) );
  DFF \creg_reg[251]  ( .D(n3350), .CLK(clk), .RST(rst), .Q(creg[251]) );
  DFF \creg_reg[252]  ( .D(n3349), .CLK(clk), .RST(rst), .Q(creg[252]) );
  DFF \creg_reg[253]  ( .D(n3348), .CLK(clk), .RST(rst), .Q(creg[253]) );
  DFF \creg_reg[254]  ( .D(n3347), .CLK(clk), .RST(rst), .Q(creg[254]) );
  DFF \creg_reg[255]  ( .D(n3602), .CLK(clk), .RST(rst), .Q(creg[255]) );
  modmult_N256_CC64 modmult_1 ( .clk(clk), .rst(rst), .start(start_in[0]), .x(
        x), .y(y), .n(n), .o(o) );
  NAND U4694 ( .A(n3860), .B(n3861), .Z(y[9]) );
  NAND U4695 ( .A(n3862), .B(m[9]), .Z(n3861) );
  NAND U4696 ( .A(n3863), .B(creg[9]), .Z(n3860) );
  NAND U4697 ( .A(n3864), .B(n3865), .Z(y[99]) );
  NAND U4698 ( .A(n3862), .B(m[99]), .Z(n3865) );
  NAND U4699 ( .A(n3863), .B(creg[99]), .Z(n3864) );
  NAND U4700 ( .A(n3866), .B(n3867), .Z(y[98]) );
  NAND U4701 ( .A(n3862), .B(m[98]), .Z(n3867) );
  NAND U4702 ( .A(n3863), .B(creg[98]), .Z(n3866) );
  NAND U4703 ( .A(n3868), .B(n3869), .Z(y[97]) );
  NAND U4704 ( .A(n3862), .B(m[97]), .Z(n3869) );
  NAND U4705 ( .A(n3863), .B(creg[97]), .Z(n3868) );
  NAND U4706 ( .A(n3870), .B(n3871), .Z(y[96]) );
  NAND U4707 ( .A(n3862), .B(m[96]), .Z(n3871) );
  NAND U4708 ( .A(n3863), .B(creg[96]), .Z(n3870) );
  NAND U4709 ( .A(n3872), .B(n3873), .Z(y[95]) );
  NAND U4710 ( .A(n3862), .B(m[95]), .Z(n3873) );
  NAND U4711 ( .A(n3863), .B(creg[95]), .Z(n3872) );
  NAND U4712 ( .A(n3874), .B(n3875), .Z(y[94]) );
  NAND U4713 ( .A(n3862), .B(m[94]), .Z(n3875) );
  NAND U4714 ( .A(n3863), .B(creg[94]), .Z(n3874) );
  NAND U4715 ( .A(n3876), .B(n3877), .Z(y[93]) );
  NAND U4716 ( .A(n3862), .B(m[93]), .Z(n3877) );
  NAND U4717 ( .A(n3863), .B(creg[93]), .Z(n3876) );
  NAND U4718 ( .A(n3878), .B(n3879), .Z(y[92]) );
  NAND U4719 ( .A(n3862), .B(m[92]), .Z(n3879) );
  NAND U4720 ( .A(n3863), .B(creg[92]), .Z(n3878) );
  NAND U4721 ( .A(n3880), .B(n3881), .Z(y[91]) );
  NAND U4722 ( .A(n3862), .B(m[91]), .Z(n3881) );
  NAND U4723 ( .A(n3863), .B(creg[91]), .Z(n3880) );
  NAND U4724 ( .A(n3882), .B(n3883), .Z(y[90]) );
  NAND U4725 ( .A(n3862), .B(m[90]), .Z(n3883) );
  NAND U4726 ( .A(n3863), .B(creg[90]), .Z(n3882) );
  NAND U4727 ( .A(n3884), .B(n3885), .Z(y[8]) );
  NAND U4728 ( .A(n3862), .B(m[8]), .Z(n3885) );
  NAND U4729 ( .A(n3863), .B(creg[8]), .Z(n3884) );
  NAND U4730 ( .A(n3886), .B(n3887), .Z(y[89]) );
  NAND U4731 ( .A(n3862), .B(m[89]), .Z(n3887) );
  NAND U4732 ( .A(n3863), .B(creg[89]), .Z(n3886) );
  NAND U4733 ( .A(n3888), .B(n3889), .Z(y[88]) );
  NAND U4734 ( .A(n3862), .B(m[88]), .Z(n3889) );
  NAND U4735 ( .A(n3863), .B(creg[88]), .Z(n3888) );
  NAND U4736 ( .A(n3890), .B(n3891), .Z(y[87]) );
  NAND U4737 ( .A(n3862), .B(m[87]), .Z(n3891) );
  NAND U4738 ( .A(n3863), .B(creg[87]), .Z(n3890) );
  NAND U4739 ( .A(n3892), .B(n3893), .Z(y[86]) );
  NAND U4740 ( .A(n3862), .B(m[86]), .Z(n3893) );
  NAND U4741 ( .A(n3863), .B(creg[86]), .Z(n3892) );
  NAND U4742 ( .A(n3894), .B(n3895), .Z(y[85]) );
  NAND U4743 ( .A(n3862), .B(m[85]), .Z(n3895) );
  NAND U4744 ( .A(n3863), .B(creg[85]), .Z(n3894) );
  NAND U4745 ( .A(n3896), .B(n3897), .Z(y[84]) );
  NAND U4746 ( .A(n3862), .B(m[84]), .Z(n3897) );
  NAND U4747 ( .A(n3863), .B(creg[84]), .Z(n3896) );
  NAND U4748 ( .A(n3898), .B(n3899), .Z(y[83]) );
  NAND U4749 ( .A(n3862), .B(m[83]), .Z(n3899) );
  NAND U4750 ( .A(n3863), .B(creg[83]), .Z(n3898) );
  NAND U4751 ( .A(n3900), .B(n3901), .Z(y[82]) );
  NAND U4752 ( .A(n3862), .B(m[82]), .Z(n3901) );
  NAND U4753 ( .A(n3863), .B(creg[82]), .Z(n3900) );
  NAND U4754 ( .A(n3902), .B(n3903), .Z(y[81]) );
  NAND U4755 ( .A(n3862), .B(m[81]), .Z(n3903) );
  NAND U4756 ( .A(n3863), .B(creg[81]), .Z(n3902) );
  NAND U4757 ( .A(n3904), .B(n3905), .Z(y[80]) );
  NAND U4758 ( .A(n3862), .B(m[80]), .Z(n3905) );
  NAND U4759 ( .A(n3863), .B(creg[80]), .Z(n3904) );
  NAND U4760 ( .A(n3906), .B(n3907), .Z(y[7]) );
  NAND U4761 ( .A(n3862), .B(m[7]), .Z(n3907) );
  NAND U4762 ( .A(n3863), .B(creg[7]), .Z(n3906) );
  NAND U4763 ( .A(n3908), .B(n3909), .Z(y[79]) );
  NAND U4764 ( .A(n3862), .B(m[79]), .Z(n3909) );
  NAND U4765 ( .A(n3863), .B(creg[79]), .Z(n3908) );
  NAND U4766 ( .A(n3910), .B(n3911), .Z(y[78]) );
  NAND U4767 ( .A(n3862), .B(m[78]), .Z(n3911) );
  NAND U4768 ( .A(n3863), .B(creg[78]), .Z(n3910) );
  NAND U4769 ( .A(n3912), .B(n3913), .Z(y[77]) );
  NAND U4770 ( .A(n3862), .B(m[77]), .Z(n3913) );
  NAND U4771 ( .A(n3863), .B(creg[77]), .Z(n3912) );
  NAND U4772 ( .A(n3914), .B(n3915), .Z(y[76]) );
  NAND U4773 ( .A(n3862), .B(m[76]), .Z(n3915) );
  NAND U4774 ( .A(n3863), .B(creg[76]), .Z(n3914) );
  NAND U4775 ( .A(n3916), .B(n3917), .Z(y[75]) );
  NAND U4776 ( .A(n3862), .B(m[75]), .Z(n3917) );
  NAND U4777 ( .A(n3863), .B(creg[75]), .Z(n3916) );
  NAND U4778 ( .A(n3918), .B(n3919), .Z(y[74]) );
  NAND U4779 ( .A(n3862), .B(m[74]), .Z(n3919) );
  NAND U4780 ( .A(n3863), .B(creg[74]), .Z(n3918) );
  NAND U4781 ( .A(n3920), .B(n3921), .Z(y[73]) );
  NAND U4782 ( .A(n3862), .B(m[73]), .Z(n3921) );
  NAND U4783 ( .A(n3863), .B(creg[73]), .Z(n3920) );
  NAND U4784 ( .A(n3922), .B(n3923), .Z(y[72]) );
  NAND U4785 ( .A(n3862), .B(m[72]), .Z(n3923) );
  NAND U4786 ( .A(n3863), .B(creg[72]), .Z(n3922) );
  NAND U4787 ( .A(n3924), .B(n3925), .Z(y[71]) );
  NAND U4788 ( .A(n3862), .B(m[71]), .Z(n3925) );
  NAND U4789 ( .A(n3863), .B(creg[71]), .Z(n3924) );
  NAND U4790 ( .A(n3926), .B(n3927), .Z(y[70]) );
  NAND U4791 ( .A(n3862), .B(m[70]), .Z(n3927) );
  NAND U4792 ( .A(n3863), .B(creg[70]), .Z(n3926) );
  NAND U4793 ( .A(n3928), .B(n3929), .Z(y[6]) );
  NAND U4794 ( .A(n3862), .B(m[6]), .Z(n3929) );
  NAND U4795 ( .A(n3863), .B(creg[6]), .Z(n3928) );
  NAND U4796 ( .A(n3930), .B(n3931), .Z(y[69]) );
  NAND U4797 ( .A(n3862), .B(m[69]), .Z(n3931) );
  NAND U4798 ( .A(n3863), .B(creg[69]), .Z(n3930) );
  NAND U4799 ( .A(n3932), .B(n3933), .Z(y[68]) );
  NAND U4800 ( .A(n3862), .B(m[68]), .Z(n3933) );
  NAND U4801 ( .A(n3863), .B(creg[68]), .Z(n3932) );
  NAND U4802 ( .A(n3934), .B(n3935), .Z(y[67]) );
  NAND U4803 ( .A(n3862), .B(m[67]), .Z(n3935) );
  NAND U4804 ( .A(n3863), .B(creg[67]), .Z(n3934) );
  NAND U4805 ( .A(n3936), .B(n3937), .Z(y[66]) );
  NAND U4806 ( .A(n3862), .B(m[66]), .Z(n3937) );
  NAND U4807 ( .A(n3863), .B(creg[66]), .Z(n3936) );
  NAND U4808 ( .A(n3938), .B(n3939), .Z(y[65]) );
  NAND U4809 ( .A(n3862), .B(m[65]), .Z(n3939) );
  NAND U4810 ( .A(n3863), .B(creg[65]), .Z(n3938) );
  NAND U4811 ( .A(n3940), .B(n3941), .Z(y[64]) );
  NAND U4812 ( .A(n3862), .B(m[64]), .Z(n3941) );
  NAND U4813 ( .A(n3863), .B(creg[64]), .Z(n3940) );
  NAND U4814 ( .A(n3942), .B(n3943), .Z(y[63]) );
  NAND U4815 ( .A(n3862), .B(m[63]), .Z(n3943) );
  NAND U4816 ( .A(n3863), .B(creg[63]), .Z(n3942) );
  NAND U4817 ( .A(n3944), .B(n3945), .Z(y[62]) );
  NAND U4818 ( .A(n3862), .B(m[62]), .Z(n3945) );
  NAND U4819 ( .A(n3863), .B(creg[62]), .Z(n3944) );
  NAND U4820 ( .A(n3946), .B(n3947), .Z(y[61]) );
  NAND U4821 ( .A(n3862), .B(m[61]), .Z(n3947) );
  NAND U4822 ( .A(n3863), .B(creg[61]), .Z(n3946) );
  NAND U4823 ( .A(n3948), .B(n3949), .Z(y[60]) );
  NAND U4824 ( .A(n3862), .B(m[60]), .Z(n3949) );
  NAND U4825 ( .A(n3863), .B(creg[60]), .Z(n3948) );
  NAND U4826 ( .A(n3950), .B(n3951), .Z(y[5]) );
  NAND U4827 ( .A(n3862), .B(m[5]), .Z(n3951) );
  NAND U4828 ( .A(n3863), .B(creg[5]), .Z(n3950) );
  NAND U4829 ( .A(n3952), .B(n3953), .Z(y[59]) );
  NAND U4830 ( .A(n3862), .B(m[59]), .Z(n3953) );
  NAND U4831 ( .A(n3863), .B(creg[59]), .Z(n3952) );
  NAND U4832 ( .A(n3954), .B(n3955), .Z(y[58]) );
  NAND U4833 ( .A(n3862), .B(m[58]), .Z(n3955) );
  NAND U4834 ( .A(n3863), .B(creg[58]), .Z(n3954) );
  NAND U4835 ( .A(n3956), .B(n3957), .Z(y[57]) );
  NAND U4836 ( .A(n3862), .B(m[57]), .Z(n3957) );
  NAND U4837 ( .A(n3863), .B(creg[57]), .Z(n3956) );
  NAND U4838 ( .A(n3958), .B(n3959), .Z(y[56]) );
  NAND U4839 ( .A(n3862), .B(m[56]), .Z(n3959) );
  NAND U4840 ( .A(n3863), .B(creg[56]), .Z(n3958) );
  NAND U4841 ( .A(n3960), .B(n3961), .Z(y[55]) );
  NAND U4842 ( .A(n3862), .B(m[55]), .Z(n3961) );
  NAND U4843 ( .A(n3863), .B(creg[55]), .Z(n3960) );
  NAND U4844 ( .A(n3962), .B(n3963), .Z(y[54]) );
  NAND U4845 ( .A(n3862), .B(m[54]), .Z(n3963) );
  NAND U4846 ( .A(n3863), .B(creg[54]), .Z(n3962) );
  NAND U4847 ( .A(n3964), .B(n3965), .Z(y[53]) );
  NAND U4848 ( .A(n3862), .B(m[53]), .Z(n3965) );
  NAND U4849 ( .A(n3863), .B(creg[53]), .Z(n3964) );
  NAND U4850 ( .A(n3966), .B(n3967), .Z(y[52]) );
  NAND U4851 ( .A(n3862), .B(m[52]), .Z(n3967) );
  NAND U4852 ( .A(n3863), .B(creg[52]), .Z(n3966) );
  NAND U4853 ( .A(n3968), .B(n3969), .Z(y[51]) );
  NAND U4854 ( .A(n3862), .B(m[51]), .Z(n3969) );
  NAND U4855 ( .A(n3863), .B(creg[51]), .Z(n3968) );
  NAND U4856 ( .A(n3970), .B(n3971), .Z(y[50]) );
  NAND U4857 ( .A(n3862), .B(m[50]), .Z(n3971) );
  NAND U4858 ( .A(n3863), .B(creg[50]), .Z(n3970) );
  NAND U4859 ( .A(n3972), .B(n3973), .Z(y[4]) );
  NAND U4860 ( .A(n3862), .B(m[4]), .Z(n3973) );
  NAND U4861 ( .A(n3863), .B(creg[4]), .Z(n3972) );
  NAND U4862 ( .A(n3974), .B(n3975), .Z(y[49]) );
  NAND U4863 ( .A(n3862), .B(m[49]), .Z(n3975) );
  NAND U4864 ( .A(n3863), .B(creg[49]), .Z(n3974) );
  NAND U4865 ( .A(n3976), .B(n3977), .Z(y[48]) );
  NAND U4866 ( .A(n3862), .B(m[48]), .Z(n3977) );
  NAND U4867 ( .A(n3863), .B(creg[48]), .Z(n3976) );
  NAND U4868 ( .A(n3978), .B(n3979), .Z(y[47]) );
  NAND U4869 ( .A(n3862), .B(m[47]), .Z(n3979) );
  NAND U4870 ( .A(n3863), .B(creg[47]), .Z(n3978) );
  NAND U4871 ( .A(n3980), .B(n3981), .Z(y[46]) );
  NAND U4872 ( .A(n3862), .B(m[46]), .Z(n3981) );
  NAND U4873 ( .A(n3863), .B(creg[46]), .Z(n3980) );
  NAND U4874 ( .A(n3982), .B(n3983), .Z(y[45]) );
  NAND U4875 ( .A(n3862), .B(m[45]), .Z(n3983) );
  NAND U4876 ( .A(n3863), .B(creg[45]), .Z(n3982) );
  NAND U4877 ( .A(n3984), .B(n3985), .Z(y[44]) );
  NAND U4878 ( .A(n3862), .B(m[44]), .Z(n3985) );
  NAND U4879 ( .A(n3863), .B(creg[44]), .Z(n3984) );
  NAND U4880 ( .A(n3986), .B(n3987), .Z(y[43]) );
  NAND U4881 ( .A(n3862), .B(m[43]), .Z(n3987) );
  NAND U4882 ( .A(n3863), .B(creg[43]), .Z(n3986) );
  NAND U4883 ( .A(n3988), .B(n3989), .Z(y[42]) );
  NAND U4884 ( .A(n3862), .B(m[42]), .Z(n3989) );
  NAND U4885 ( .A(n3863), .B(creg[42]), .Z(n3988) );
  NAND U4886 ( .A(n3990), .B(n3991), .Z(y[41]) );
  NAND U4887 ( .A(n3862), .B(m[41]), .Z(n3991) );
  NAND U4888 ( .A(n3863), .B(creg[41]), .Z(n3990) );
  NAND U4889 ( .A(n3992), .B(n3993), .Z(y[40]) );
  NAND U4890 ( .A(n3862), .B(m[40]), .Z(n3993) );
  NAND U4891 ( .A(n3863), .B(creg[40]), .Z(n3992) );
  NAND U4892 ( .A(n3994), .B(n3995), .Z(y[3]) );
  NAND U4893 ( .A(n3862), .B(m[3]), .Z(n3995) );
  NAND U4894 ( .A(n3863), .B(creg[3]), .Z(n3994) );
  NAND U4895 ( .A(n3996), .B(n3997), .Z(y[39]) );
  NAND U4896 ( .A(n3862), .B(m[39]), .Z(n3997) );
  NAND U4897 ( .A(n3863), .B(creg[39]), .Z(n3996) );
  NAND U4898 ( .A(n3998), .B(n3999), .Z(y[38]) );
  NAND U4899 ( .A(n3862), .B(m[38]), .Z(n3999) );
  NAND U4900 ( .A(n3863), .B(creg[38]), .Z(n3998) );
  NAND U4901 ( .A(n4000), .B(n4001), .Z(y[37]) );
  NAND U4902 ( .A(n3862), .B(m[37]), .Z(n4001) );
  NAND U4903 ( .A(n3863), .B(creg[37]), .Z(n4000) );
  NAND U4904 ( .A(n4002), .B(n4003), .Z(y[36]) );
  NAND U4905 ( .A(n3862), .B(m[36]), .Z(n4003) );
  NAND U4906 ( .A(n3863), .B(creg[36]), .Z(n4002) );
  NAND U4907 ( .A(n4004), .B(n4005), .Z(y[35]) );
  NAND U4908 ( .A(n3862), .B(m[35]), .Z(n4005) );
  NAND U4909 ( .A(n3863), .B(creg[35]), .Z(n4004) );
  NAND U4910 ( .A(n4006), .B(n4007), .Z(y[34]) );
  NAND U4911 ( .A(n3862), .B(m[34]), .Z(n4007) );
  NAND U4912 ( .A(n3863), .B(creg[34]), .Z(n4006) );
  NAND U4913 ( .A(n4008), .B(n4009), .Z(y[33]) );
  NAND U4914 ( .A(n3862), .B(m[33]), .Z(n4009) );
  NAND U4915 ( .A(n3863), .B(creg[33]), .Z(n4008) );
  NAND U4916 ( .A(n4010), .B(n4011), .Z(y[32]) );
  NAND U4917 ( .A(n3862), .B(m[32]), .Z(n4011) );
  NAND U4918 ( .A(n3863), .B(creg[32]), .Z(n4010) );
  NAND U4919 ( .A(n4012), .B(n4013), .Z(y[31]) );
  NAND U4920 ( .A(n3862), .B(m[31]), .Z(n4013) );
  NAND U4921 ( .A(n3863), .B(creg[31]), .Z(n4012) );
  NAND U4922 ( .A(n4014), .B(n4015), .Z(y[30]) );
  NAND U4923 ( .A(n3862), .B(m[30]), .Z(n4015) );
  NAND U4924 ( .A(n3863), .B(creg[30]), .Z(n4014) );
  NAND U4925 ( .A(n4016), .B(n4017), .Z(y[2]) );
  NAND U4926 ( .A(n3862), .B(m[2]), .Z(n4017) );
  NAND U4927 ( .A(n3863), .B(creg[2]), .Z(n4016) );
  NAND U4928 ( .A(n4018), .B(n4019), .Z(y[29]) );
  NAND U4929 ( .A(n3862), .B(m[29]), .Z(n4019) );
  NAND U4930 ( .A(n3863), .B(creg[29]), .Z(n4018) );
  NAND U4931 ( .A(n4020), .B(n4021), .Z(y[28]) );
  NAND U4932 ( .A(n3862), .B(m[28]), .Z(n4021) );
  NAND U4933 ( .A(n3863), .B(creg[28]), .Z(n4020) );
  NAND U4934 ( .A(n4022), .B(n4023), .Z(y[27]) );
  NAND U4935 ( .A(n3862), .B(m[27]), .Z(n4023) );
  NAND U4936 ( .A(n3863), .B(creg[27]), .Z(n4022) );
  NAND U4937 ( .A(n4024), .B(n4025), .Z(y[26]) );
  NAND U4938 ( .A(n3862), .B(m[26]), .Z(n4025) );
  NAND U4939 ( .A(n3863), .B(creg[26]), .Z(n4024) );
  NAND U4940 ( .A(n4026), .B(n4027), .Z(y[25]) );
  NAND U4941 ( .A(n3862), .B(m[25]), .Z(n4027) );
  NAND U4942 ( .A(n3863), .B(creg[25]), .Z(n4026) );
  NAND U4943 ( .A(n4028), .B(n4029), .Z(y[255]) );
  NAND U4944 ( .A(n3862), .B(m[255]), .Z(n4029) );
  NAND U4945 ( .A(n3863), .B(creg[255]), .Z(n4028) );
  NAND U4946 ( .A(n4030), .B(n4031), .Z(y[254]) );
  NAND U4947 ( .A(n3862), .B(m[254]), .Z(n4031) );
  NAND U4948 ( .A(n3863), .B(creg[254]), .Z(n4030) );
  NAND U4949 ( .A(n4032), .B(n4033), .Z(y[253]) );
  NAND U4950 ( .A(n3862), .B(m[253]), .Z(n4033) );
  NAND U4951 ( .A(n3863), .B(creg[253]), .Z(n4032) );
  NAND U4952 ( .A(n4034), .B(n4035), .Z(y[252]) );
  NAND U4953 ( .A(n3862), .B(m[252]), .Z(n4035) );
  NAND U4954 ( .A(n3863), .B(creg[252]), .Z(n4034) );
  NAND U4955 ( .A(n4036), .B(n4037), .Z(y[251]) );
  NAND U4956 ( .A(n3862), .B(m[251]), .Z(n4037) );
  NAND U4957 ( .A(n3863), .B(creg[251]), .Z(n4036) );
  NAND U4958 ( .A(n4038), .B(n4039), .Z(y[250]) );
  NAND U4959 ( .A(n3862), .B(m[250]), .Z(n4039) );
  NAND U4960 ( .A(n3863), .B(creg[250]), .Z(n4038) );
  NAND U4961 ( .A(n4040), .B(n4041), .Z(y[24]) );
  NAND U4962 ( .A(n3862), .B(m[24]), .Z(n4041) );
  NAND U4963 ( .A(n3863), .B(creg[24]), .Z(n4040) );
  NAND U4964 ( .A(n4042), .B(n4043), .Z(y[249]) );
  NAND U4965 ( .A(n3862), .B(m[249]), .Z(n4043) );
  NAND U4966 ( .A(n3863), .B(creg[249]), .Z(n4042) );
  NAND U4967 ( .A(n4044), .B(n4045), .Z(y[248]) );
  NAND U4968 ( .A(n3862), .B(m[248]), .Z(n4045) );
  NAND U4969 ( .A(n3863), .B(creg[248]), .Z(n4044) );
  NAND U4970 ( .A(n4046), .B(n4047), .Z(y[247]) );
  NAND U4971 ( .A(n3862), .B(m[247]), .Z(n4047) );
  NAND U4972 ( .A(n3863), .B(creg[247]), .Z(n4046) );
  NAND U4973 ( .A(n4048), .B(n4049), .Z(y[246]) );
  NAND U4974 ( .A(n3862), .B(m[246]), .Z(n4049) );
  NAND U4975 ( .A(n3863), .B(creg[246]), .Z(n4048) );
  NAND U4976 ( .A(n4050), .B(n4051), .Z(y[245]) );
  NAND U4977 ( .A(n3862), .B(m[245]), .Z(n4051) );
  NAND U4978 ( .A(n3863), .B(creg[245]), .Z(n4050) );
  NAND U4979 ( .A(n4052), .B(n4053), .Z(y[244]) );
  NAND U4980 ( .A(n3862), .B(m[244]), .Z(n4053) );
  NAND U4981 ( .A(n3863), .B(creg[244]), .Z(n4052) );
  NAND U4982 ( .A(n4054), .B(n4055), .Z(y[243]) );
  NAND U4983 ( .A(n3862), .B(m[243]), .Z(n4055) );
  NAND U4984 ( .A(n3863), .B(creg[243]), .Z(n4054) );
  NAND U4985 ( .A(n4056), .B(n4057), .Z(y[242]) );
  NAND U4986 ( .A(n3862), .B(m[242]), .Z(n4057) );
  NAND U4987 ( .A(n3863), .B(creg[242]), .Z(n4056) );
  NAND U4988 ( .A(n4058), .B(n4059), .Z(y[241]) );
  NAND U4989 ( .A(n3862), .B(m[241]), .Z(n4059) );
  NAND U4990 ( .A(n3863), .B(creg[241]), .Z(n4058) );
  NAND U4991 ( .A(n4060), .B(n4061), .Z(y[240]) );
  NAND U4992 ( .A(n3862), .B(m[240]), .Z(n4061) );
  NAND U4993 ( .A(n3863), .B(creg[240]), .Z(n4060) );
  NAND U4994 ( .A(n4062), .B(n4063), .Z(y[23]) );
  NAND U4995 ( .A(n3862), .B(m[23]), .Z(n4063) );
  NAND U4996 ( .A(n3863), .B(creg[23]), .Z(n4062) );
  NAND U4997 ( .A(n4064), .B(n4065), .Z(y[239]) );
  NAND U4998 ( .A(n3862), .B(m[239]), .Z(n4065) );
  NAND U4999 ( .A(n3863), .B(creg[239]), .Z(n4064) );
  NAND U5000 ( .A(n4066), .B(n4067), .Z(y[238]) );
  NAND U5001 ( .A(n3862), .B(m[238]), .Z(n4067) );
  NAND U5002 ( .A(n3863), .B(creg[238]), .Z(n4066) );
  NAND U5003 ( .A(n4068), .B(n4069), .Z(y[237]) );
  NAND U5004 ( .A(n3862), .B(m[237]), .Z(n4069) );
  NAND U5005 ( .A(n3863), .B(creg[237]), .Z(n4068) );
  NAND U5006 ( .A(n4070), .B(n4071), .Z(y[236]) );
  NAND U5007 ( .A(n3862), .B(m[236]), .Z(n4071) );
  NAND U5008 ( .A(n3863), .B(creg[236]), .Z(n4070) );
  NAND U5009 ( .A(n4072), .B(n4073), .Z(y[235]) );
  NAND U5010 ( .A(n3862), .B(m[235]), .Z(n4073) );
  NAND U5011 ( .A(n3863), .B(creg[235]), .Z(n4072) );
  NAND U5012 ( .A(n4074), .B(n4075), .Z(y[234]) );
  NAND U5013 ( .A(n3862), .B(m[234]), .Z(n4075) );
  NAND U5014 ( .A(n3863), .B(creg[234]), .Z(n4074) );
  NAND U5015 ( .A(n4076), .B(n4077), .Z(y[233]) );
  NAND U5016 ( .A(n3862), .B(m[233]), .Z(n4077) );
  NAND U5017 ( .A(n3863), .B(creg[233]), .Z(n4076) );
  NAND U5018 ( .A(n4078), .B(n4079), .Z(y[232]) );
  NAND U5019 ( .A(n3862), .B(m[232]), .Z(n4079) );
  NAND U5020 ( .A(n3863), .B(creg[232]), .Z(n4078) );
  NAND U5021 ( .A(n4080), .B(n4081), .Z(y[231]) );
  NAND U5022 ( .A(n3862), .B(m[231]), .Z(n4081) );
  NAND U5023 ( .A(n3863), .B(creg[231]), .Z(n4080) );
  NAND U5024 ( .A(n4082), .B(n4083), .Z(y[230]) );
  NAND U5025 ( .A(n3862), .B(m[230]), .Z(n4083) );
  NAND U5026 ( .A(n3863), .B(creg[230]), .Z(n4082) );
  NAND U5027 ( .A(n4084), .B(n4085), .Z(y[22]) );
  NAND U5028 ( .A(n3862), .B(m[22]), .Z(n4085) );
  NAND U5029 ( .A(n3863), .B(creg[22]), .Z(n4084) );
  NAND U5030 ( .A(n4086), .B(n4087), .Z(y[229]) );
  NAND U5031 ( .A(n3862), .B(m[229]), .Z(n4087) );
  NAND U5032 ( .A(n3863), .B(creg[229]), .Z(n4086) );
  NAND U5033 ( .A(n4088), .B(n4089), .Z(y[228]) );
  NAND U5034 ( .A(n3862), .B(m[228]), .Z(n4089) );
  NAND U5035 ( .A(n3863), .B(creg[228]), .Z(n4088) );
  NAND U5036 ( .A(n4090), .B(n4091), .Z(y[227]) );
  NAND U5037 ( .A(n3862), .B(m[227]), .Z(n4091) );
  NAND U5038 ( .A(n3863), .B(creg[227]), .Z(n4090) );
  NAND U5039 ( .A(n4092), .B(n4093), .Z(y[226]) );
  NAND U5040 ( .A(n3862), .B(m[226]), .Z(n4093) );
  NAND U5041 ( .A(n3863), .B(creg[226]), .Z(n4092) );
  NAND U5042 ( .A(n4094), .B(n4095), .Z(y[225]) );
  NAND U5043 ( .A(n3862), .B(m[225]), .Z(n4095) );
  NAND U5044 ( .A(n3863), .B(creg[225]), .Z(n4094) );
  NAND U5045 ( .A(n4096), .B(n4097), .Z(y[224]) );
  NAND U5046 ( .A(n3862), .B(m[224]), .Z(n4097) );
  NAND U5047 ( .A(n3863), .B(creg[224]), .Z(n4096) );
  NAND U5048 ( .A(n4098), .B(n4099), .Z(y[223]) );
  NAND U5049 ( .A(n3862), .B(m[223]), .Z(n4099) );
  NAND U5050 ( .A(n3863), .B(creg[223]), .Z(n4098) );
  NAND U5051 ( .A(n4100), .B(n4101), .Z(y[222]) );
  NAND U5052 ( .A(n3862), .B(m[222]), .Z(n4101) );
  NAND U5053 ( .A(n3863), .B(creg[222]), .Z(n4100) );
  NAND U5054 ( .A(n4102), .B(n4103), .Z(y[221]) );
  NAND U5055 ( .A(n3862), .B(m[221]), .Z(n4103) );
  NAND U5056 ( .A(n3863), .B(creg[221]), .Z(n4102) );
  NAND U5057 ( .A(n4104), .B(n4105), .Z(y[220]) );
  NAND U5058 ( .A(n3862), .B(m[220]), .Z(n4105) );
  NAND U5059 ( .A(n3863), .B(creg[220]), .Z(n4104) );
  NAND U5060 ( .A(n4106), .B(n4107), .Z(y[21]) );
  NAND U5061 ( .A(n3862), .B(m[21]), .Z(n4107) );
  NAND U5062 ( .A(n3863), .B(creg[21]), .Z(n4106) );
  NAND U5063 ( .A(n4108), .B(n4109), .Z(y[219]) );
  NAND U5064 ( .A(n3862), .B(m[219]), .Z(n4109) );
  NAND U5065 ( .A(n3863), .B(creg[219]), .Z(n4108) );
  NAND U5066 ( .A(n4110), .B(n4111), .Z(y[218]) );
  NAND U5067 ( .A(n3862), .B(m[218]), .Z(n4111) );
  NAND U5068 ( .A(n3863), .B(creg[218]), .Z(n4110) );
  NAND U5069 ( .A(n4112), .B(n4113), .Z(y[217]) );
  NAND U5070 ( .A(n3862), .B(m[217]), .Z(n4113) );
  NAND U5071 ( .A(n3863), .B(creg[217]), .Z(n4112) );
  NAND U5072 ( .A(n4114), .B(n4115), .Z(y[216]) );
  NAND U5073 ( .A(n3862), .B(m[216]), .Z(n4115) );
  NAND U5074 ( .A(n3863), .B(creg[216]), .Z(n4114) );
  NAND U5075 ( .A(n4116), .B(n4117), .Z(y[215]) );
  NAND U5076 ( .A(n3862), .B(m[215]), .Z(n4117) );
  NAND U5077 ( .A(n3863), .B(creg[215]), .Z(n4116) );
  NAND U5078 ( .A(n4118), .B(n4119), .Z(y[214]) );
  NAND U5079 ( .A(n3862), .B(m[214]), .Z(n4119) );
  NAND U5080 ( .A(n3863), .B(creg[214]), .Z(n4118) );
  NAND U5081 ( .A(n4120), .B(n4121), .Z(y[213]) );
  NAND U5082 ( .A(n3862), .B(m[213]), .Z(n4121) );
  NAND U5083 ( .A(n3863), .B(creg[213]), .Z(n4120) );
  NAND U5084 ( .A(n4122), .B(n4123), .Z(y[212]) );
  NAND U5085 ( .A(n3862), .B(m[212]), .Z(n4123) );
  NAND U5086 ( .A(n3863), .B(creg[212]), .Z(n4122) );
  NAND U5087 ( .A(n4124), .B(n4125), .Z(y[211]) );
  NAND U5088 ( .A(n3862), .B(m[211]), .Z(n4125) );
  NAND U5089 ( .A(n3863), .B(creg[211]), .Z(n4124) );
  NAND U5090 ( .A(n4126), .B(n4127), .Z(y[210]) );
  NAND U5091 ( .A(n3862), .B(m[210]), .Z(n4127) );
  NAND U5092 ( .A(n3863), .B(creg[210]), .Z(n4126) );
  NAND U5093 ( .A(n4128), .B(n4129), .Z(y[20]) );
  NAND U5094 ( .A(n3862), .B(m[20]), .Z(n4129) );
  NAND U5095 ( .A(n3863), .B(creg[20]), .Z(n4128) );
  NAND U5096 ( .A(n4130), .B(n4131), .Z(y[209]) );
  NAND U5097 ( .A(n3862), .B(m[209]), .Z(n4131) );
  NAND U5098 ( .A(n3863), .B(creg[209]), .Z(n4130) );
  NAND U5099 ( .A(n4132), .B(n4133), .Z(y[208]) );
  NAND U5100 ( .A(n3862), .B(m[208]), .Z(n4133) );
  NAND U5101 ( .A(n3863), .B(creg[208]), .Z(n4132) );
  NAND U5102 ( .A(n4134), .B(n4135), .Z(y[207]) );
  NAND U5103 ( .A(n3862), .B(m[207]), .Z(n4135) );
  NAND U5104 ( .A(n3863), .B(creg[207]), .Z(n4134) );
  NAND U5105 ( .A(n4136), .B(n4137), .Z(y[206]) );
  NAND U5106 ( .A(n3862), .B(m[206]), .Z(n4137) );
  NAND U5107 ( .A(n3863), .B(creg[206]), .Z(n4136) );
  NAND U5108 ( .A(n4138), .B(n4139), .Z(y[205]) );
  NAND U5109 ( .A(n3862), .B(m[205]), .Z(n4139) );
  NAND U5110 ( .A(n3863), .B(creg[205]), .Z(n4138) );
  NAND U5111 ( .A(n4140), .B(n4141), .Z(y[204]) );
  NAND U5112 ( .A(n3862), .B(m[204]), .Z(n4141) );
  NAND U5113 ( .A(n3863), .B(creg[204]), .Z(n4140) );
  NAND U5114 ( .A(n4142), .B(n4143), .Z(y[203]) );
  NAND U5115 ( .A(n3862), .B(m[203]), .Z(n4143) );
  NAND U5116 ( .A(n3863), .B(creg[203]), .Z(n4142) );
  NAND U5117 ( .A(n4144), .B(n4145), .Z(y[202]) );
  NAND U5118 ( .A(n3862), .B(m[202]), .Z(n4145) );
  NAND U5119 ( .A(n3863), .B(creg[202]), .Z(n4144) );
  NAND U5120 ( .A(n4146), .B(n4147), .Z(y[201]) );
  NAND U5121 ( .A(n3862), .B(m[201]), .Z(n4147) );
  NAND U5122 ( .A(n3863), .B(creg[201]), .Z(n4146) );
  NAND U5123 ( .A(n4148), .B(n4149), .Z(y[200]) );
  NAND U5124 ( .A(n3862), .B(m[200]), .Z(n4149) );
  NAND U5125 ( .A(n3863), .B(creg[200]), .Z(n4148) );
  NAND U5126 ( .A(n4150), .B(n4151), .Z(y[1]) );
  NAND U5127 ( .A(n3862), .B(m[1]), .Z(n4151) );
  NAND U5128 ( .A(n3863), .B(creg[1]), .Z(n4150) );
  NAND U5129 ( .A(n4152), .B(n4153), .Z(y[19]) );
  NAND U5130 ( .A(n3862), .B(m[19]), .Z(n4153) );
  NAND U5131 ( .A(n3863), .B(creg[19]), .Z(n4152) );
  NAND U5132 ( .A(n4154), .B(n4155), .Z(y[199]) );
  NAND U5133 ( .A(n3862), .B(m[199]), .Z(n4155) );
  NAND U5134 ( .A(n3863), .B(creg[199]), .Z(n4154) );
  NAND U5135 ( .A(n4156), .B(n4157), .Z(y[198]) );
  NAND U5136 ( .A(n3862), .B(m[198]), .Z(n4157) );
  NAND U5137 ( .A(n3863), .B(creg[198]), .Z(n4156) );
  NAND U5138 ( .A(n4158), .B(n4159), .Z(y[197]) );
  NAND U5139 ( .A(n3862), .B(m[197]), .Z(n4159) );
  NAND U5140 ( .A(n3863), .B(creg[197]), .Z(n4158) );
  NAND U5141 ( .A(n4160), .B(n4161), .Z(y[196]) );
  NAND U5142 ( .A(n3862), .B(m[196]), .Z(n4161) );
  NAND U5143 ( .A(n3863), .B(creg[196]), .Z(n4160) );
  NAND U5144 ( .A(n4162), .B(n4163), .Z(y[195]) );
  NAND U5145 ( .A(n3862), .B(m[195]), .Z(n4163) );
  NAND U5146 ( .A(n3863), .B(creg[195]), .Z(n4162) );
  NAND U5147 ( .A(n4164), .B(n4165), .Z(y[194]) );
  NAND U5148 ( .A(n3862), .B(m[194]), .Z(n4165) );
  NAND U5149 ( .A(n3863), .B(creg[194]), .Z(n4164) );
  NAND U5150 ( .A(n4166), .B(n4167), .Z(y[193]) );
  NAND U5151 ( .A(n3862), .B(m[193]), .Z(n4167) );
  NAND U5152 ( .A(n3863), .B(creg[193]), .Z(n4166) );
  NAND U5153 ( .A(n4168), .B(n4169), .Z(y[192]) );
  NAND U5154 ( .A(n3862), .B(m[192]), .Z(n4169) );
  NAND U5155 ( .A(n3863), .B(creg[192]), .Z(n4168) );
  NAND U5156 ( .A(n4170), .B(n4171), .Z(y[191]) );
  NAND U5157 ( .A(n3862), .B(m[191]), .Z(n4171) );
  NAND U5158 ( .A(n3863), .B(creg[191]), .Z(n4170) );
  NAND U5159 ( .A(n4172), .B(n4173), .Z(y[190]) );
  NAND U5160 ( .A(n3862), .B(m[190]), .Z(n4173) );
  NAND U5161 ( .A(n3863), .B(creg[190]), .Z(n4172) );
  NAND U5162 ( .A(n4174), .B(n4175), .Z(y[18]) );
  NAND U5163 ( .A(n3862), .B(m[18]), .Z(n4175) );
  NAND U5164 ( .A(n3863), .B(creg[18]), .Z(n4174) );
  NAND U5165 ( .A(n4176), .B(n4177), .Z(y[189]) );
  NAND U5166 ( .A(n3862), .B(m[189]), .Z(n4177) );
  NAND U5167 ( .A(n3863), .B(creg[189]), .Z(n4176) );
  NAND U5168 ( .A(n4178), .B(n4179), .Z(y[188]) );
  NAND U5169 ( .A(n3862), .B(m[188]), .Z(n4179) );
  NAND U5170 ( .A(n3863), .B(creg[188]), .Z(n4178) );
  NAND U5171 ( .A(n4180), .B(n4181), .Z(y[187]) );
  NAND U5172 ( .A(n3862), .B(m[187]), .Z(n4181) );
  NAND U5173 ( .A(n3863), .B(creg[187]), .Z(n4180) );
  NAND U5174 ( .A(n4182), .B(n4183), .Z(y[186]) );
  NAND U5175 ( .A(n3862), .B(m[186]), .Z(n4183) );
  NAND U5176 ( .A(n3863), .B(creg[186]), .Z(n4182) );
  NAND U5177 ( .A(n4184), .B(n4185), .Z(y[185]) );
  NAND U5178 ( .A(n3862), .B(m[185]), .Z(n4185) );
  NAND U5179 ( .A(n3863), .B(creg[185]), .Z(n4184) );
  NAND U5180 ( .A(n4186), .B(n4187), .Z(y[184]) );
  NAND U5181 ( .A(n3862), .B(m[184]), .Z(n4187) );
  NAND U5182 ( .A(n3863), .B(creg[184]), .Z(n4186) );
  NAND U5183 ( .A(n4188), .B(n4189), .Z(y[183]) );
  NAND U5184 ( .A(n3862), .B(m[183]), .Z(n4189) );
  NAND U5185 ( .A(n3863), .B(creg[183]), .Z(n4188) );
  NAND U5186 ( .A(n4190), .B(n4191), .Z(y[182]) );
  NAND U5187 ( .A(n3862), .B(m[182]), .Z(n4191) );
  NAND U5188 ( .A(n3863), .B(creg[182]), .Z(n4190) );
  NAND U5189 ( .A(n4192), .B(n4193), .Z(y[181]) );
  NAND U5190 ( .A(n3862), .B(m[181]), .Z(n4193) );
  NAND U5191 ( .A(n3863), .B(creg[181]), .Z(n4192) );
  NAND U5192 ( .A(n4194), .B(n4195), .Z(y[180]) );
  NAND U5193 ( .A(n3862), .B(m[180]), .Z(n4195) );
  NAND U5194 ( .A(n3863), .B(creg[180]), .Z(n4194) );
  NAND U5195 ( .A(n4196), .B(n4197), .Z(y[17]) );
  NAND U5196 ( .A(n3862), .B(m[17]), .Z(n4197) );
  NAND U5197 ( .A(n3863), .B(creg[17]), .Z(n4196) );
  NAND U5198 ( .A(n4198), .B(n4199), .Z(y[179]) );
  NAND U5199 ( .A(n3862), .B(m[179]), .Z(n4199) );
  NAND U5200 ( .A(n3863), .B(creg[179]), .Z(n4198) );
  NAND U5201 ( .A(n4200), .B(n4201), .Z(y[178]) );
  NAND U5202 ( .A(n3862), .B(m[178]), .Z(n4201) );
  NAND U5203 ( .A(n3863), .B(creg[178]), .Z(n4200) );
  NAND U5204 ( .A(n4202), .B(n4203), .Z(y[177]) );
  NAND U5205 ( .A(n3862), .B(m[177]), .Z(n4203) );
  NAND U5206 ( .A(n3863), .B(creg[177]), .Z(n4202) );
  NAND U5207 ( .A(n4204), .B(n4205), .Z(y[176]) );
  NAND U5208 ( .A(n3862), .B(m[176]), .Z(n4205) );
  NAND U5209 ( .A(n3863), .B(creg[176]), .Z(n4204) );
  NAND U5210 ( .A(n4206), .B(n4207), .Z(y[175]) );
  NAND U5211 ( .A(n3862), .B(m[175]), .Z(n4207) );
  NAND U5212 ( .A(n3863), .B(creg[175]), .Z(n4206) );
  NAND U5213 ( .A(n4208), .B(n4209), .Z(y[174]) );
  NAND U5214 ( .A(n3862), .B(m[174]), .Z(n4209) );
  NAND U5215 ( .A(n3863), .B(creg[174]), .Z(n4208) );
  NAND U5216 ( .A(n4210), .B(n4211), .Z(y[173]) );
  NAND U5217 ( .A(n3862), .B(m[173]), .Z(n4211) );
  NAND U5218 ( .A(n3863), .B(creg[173]), .Z(n4210) );
  NAND U5219 ( .A(n4212), .B(n4213), .Z(y[172]) );
  NAND U5220 ( .A(n3862), .B(m[172]), .Z(n4213) );
  NAND U5221 ( .A(n3863), .B(creg[172]), .Z(n4212) );
  NAND U5222 ( .A(n4214), .B(n4215), .Z(y[171]) );
  NAND U5223 ( .A(n3862), .B(m[171]), .Z(n4215) );
  NAND U5224 ( .A(n3863), .B(creg[171]), .Z(n4214) );
  NAND U5225 ( .A(n4216), .B(n4217), .Z(y[170]) );
  NAND U5226 ( .A(n3862), .B(m[170]), .Z(n4217) );
  NAND U5227 ( .A(n3863), .B(creg[170]), .Z(n4216) );
  NAND U5228 ( .A(n4218), .B(n4219), .Z(y[16]) );
  NAND U5229 ( .A(n3862), .B(m[16]), .Z(n4219) );
  NAND U5230 ( .A(n3863), .B(creg[16]), .Z(n4218) );
  NAND U5231 ( .A(n4220), .B(n4221), .Z(y[169]) );
  NAND U5232 ( .A(n3862), .B(m[169]), .Z(n4221) );
  NAND U5233 ( .A(n3863), .B(creg[169]), .Z(n4220) );
  NAND U5234 ( .A(n4222), .B(n4223), .Z(y[168]) );
  NAND U5235 ( .A(n3862), .B(m[168]), .Z(n4223) );
  NAND U5236 ( .A(n3863), .B(creg[168]), .Z(n4222) );
  NAND U5237 ( .A(n4224), .B(n4225), .Z(y[167]) );
  NAND U5238 ( .A(n3862), .B(m[167]), .Z(n4225) );
  NAND U5239 ( .A(n3863), .B(creg[167]), .Z(n4224) );
  NAND U5240 ( .A(n4226), .B(n4227), .Z(y[166]) );
  NAND U5241 ( .A(n3862), .B(m[166]), .Z(n4227) );
  NAND U5242 ( .A(n3863), .B(creg[166]), .Z(n4226) );
  NAND U5243 ( .A(n4228), .B(n4229), .Z(y[165]) );
  NAND U5244 ( .A(n3862), .B(m[165]), .Z(n4229) );
  NAND U5245 ( .A(n3863), .B(creg[165]), .Z(n4228) );
  NAND U5246 ( .A(n4230), .B(n4231), .Z(y[164]) );
  NAND U5247 ( .A(n3862), .B(m[164]), .Z(n4231) );
  NAND U5248 ( .A(n3863), .B(creg[164]), .Z(n4230) );
  NAND U5249 ( .A(n4232), .B(n4233), .Z(y[163]) );
  NAND U5250 ( .A(n3862), .B(m[163]), .Z(n4233) );
  NAND U5251 ( .A(n3863), .B(creg[163]), .Z(n4232) );
  NAND U5252 ( .A(n4234), .B(n4235), .Z(y[162]) );
  NAND U5253 ( .A(n3862), .B(m[162]), .Z(n4235) );
  NAND U5254 ( .A(n3863), .B(creg[162]), .Z(n4234) );
  NAND U5255 ( .A(n4236), .B(n4237), .Z(y[161]) );
  NAND U5256 ( .A(n3862), .B(m[161]), .Z(n4237) );
  NAND U5257 ( .A(n3863), .B(creg[161]), .Z(n4236) );
  NAND U5258 ( .A(n4238), .B(n4239), .Z(y[160]) );
  NAND U5259 ( .A(n3862), .B(m[160]), .Z(n4239) );
  NAND U5260 ( .A(n3863), .B(creg[160]), .Z(n4238) );
  NAND U5261 ( .A(n4240), .B(n4241), .Z(y[15]) );
  NAND U5262 ( .A(n3862), .B(m[15]), .Z(n4241) );
  NAND U5263 ( .A(n3863), .B(creg[15]), .Z(n4240) );
  NAND U5264 ( .A(n4242), .B(n4243), .Z(y[159]) );
  NAND U5265 ( .A(n3862), .B(m[159]), .Z(n4243) );
  NAND U5266 ( .A(n3863), .B(creg[159]), .Z(n4242) );
  NAND U5267 ( .A(n4244), .B(n4245), .Z(y[158]) );
  NAND U5268 ( .A(n3862), .B(m[158]), .Z(n4245) );
  NAND U5269 ( .A(n3863), .B(creg[158]), .Z(n4244) );
  NAND U5270 ( .A(n4246), .B(n4247), .Z(y[157]) );
  NAND U5271 ( .A(n3862), .B(m[157]), .Z(n4247) );
  NAND U5272 ( .A(n3863), .B(creg[157]), .Z(n4246) );
  NAND U5273 ( .A(n4248), .B(n4249), .Z(y[156]) );
  NAND U5274 ( .A(n3862), .B(m[156]), .Z(n4249) );
  NAND U5275 ( .A(n3863), .B(creg[156]), .Z(n4248) );
  NAND U5276 ( .A(n4250), .B(n4251), .Z(y[155]) );
  NAND U5277 ( .A(n3862), .B(m[155]), .Z(n4251) );
  NAND U5278 ( .A(n3863), .B(creg[155]), .Z(n4250) );
  NAND U5279 ( .A(n4252), .B(n4253), .Z(y[154]) );
  NAND U5280 ( .A(n3862), .B(m[154]), .Z(n4253) );
  NAND U5281 ( .A(n3863), .B(creg[154]), .Z(n4252) );
  NAND U5282 ( .A(n4254), .B(n4255), .Z(y[153]) );
  NAND U5283 ( .A(n3862), .B(m[153]), .Z(n4255) );
  NAND U5284 ( .A(n3863), .B(creg[153]), .Z(n4254) );
  NAND U5285 ( .A(n4256), .B(n4257), .Z(y[152]) );
  NAND U5286 ( .A(n3862), .B(m[152]), .Z(n4257) );
  NAND U5287 ( .A(n3863), .B(creg[152]), .Z(n4256) );
  NAND U5288 ( .A(n4258), .B(n4259), .Z(y[151]) );
  NAND U5289 ( .A(n3862), .B(m[151]), .Z(n4259) );
  NAND U5290 ( .A(n3863), .B(creg[151]), .Z(n4258) );
  NAND U5291 ( .A(n4260), .B(n4261), .Z(y[150]) );
  NAND U5292 ( .A(n3862), .B(m[150]), .Z(n4261) );
  NAND U5293 ( .A(n3863), .B(creg[150]), .Z(n4260) );
  NAND U5294 ( .A(n4262), .B(n4263), .Z(y[14]) );
  NAND U5295 ( .A(n3862), .B(m[14]), .Z(n4263) );
  NAND U5296 ( .A(n3863), .B(creg[14]), .Z(n4262) );
  NAND U5297 ( .A(n4264), .B(n4265), .Z(y[149]) );
  NAND U5298 ( .A(n3862), .B(m[149]), .Z(n4265) );
  NAND U5299 ( .A(n3863), .B(creg[149]), .Z(n4264) );
  NAND U5300 ( .A(n4266), .B(n4267), .Z(y[148]) );
  NAND U5301 ( .A(n3862), .B(m[148]), .Z(n4267) );
  NAND U5302 ( .A(n3863), .B(creg[148]), .Z(n4266) );
  NAND U5303 ( .A(n4268), .B(n4269), .Z(y[147]) );
  NAND U5304 ( .A(n3862), .B(m[147]), .Z(n4269) );
  NAND U5305 ( .A(n3863), .B(creg[147]), .Z(n4268) );
  NAND U5306 ( .A(n4270), .B(n4271), .Z(y[146]) );
  NAND U5307 ( .A(n3862), .B(m[146]), .Z(n4271) );
  NAND U5308 ( .A(n3863), .B(creg[146]), .Z(n4270) );
  NAND U5309 ( .A(n4272), .B(n4273), .Z(y[145]) );
  NAND U5310 ( .A(n3862), .B(m[145]), .Z(n4273) );
  NAND U5311 ( .A(n3863), .B(creg[145]), .Z(n4272) );
  NAND U5312 ( .A(n4274), .B(n4275), .Z(y[144]) );
  NAND U5313 ( .A(n3862), .B(m[144]), .Z(n4275) );
  NAND U5314 ( .A(n3863), .B(creg[144]), .Z(n4274) );
  NAND U5315 ( .A(n4276), .B(n4277), .Z(y[143]) );
  NAND U5316 ( .A(n3862), .B(m[143]), .Z(n4277) );
  NAND U5317 ( .A(n3863), .B(creg[143]), .Z(n4276) );
  NAND U5318 ( .A(n4278), .B(n4279), .Z(y[142]) );
  NAND U5319 ( .A(n3862), .B(m[142]), .Z(n4279) );
  NAND U5320 ( .A(n3863), .B(creg[142]), .Z(n4278) );
  NAND U5321 ( .A(n4280), .B(n4281), .Z(y[141]) );
  NAND U5322 ( .A(n3862), .B(m[141]), .Z(n4281) );
  NAND U5323 ( .A(n3863), .B(creg[141]), .Z(n4280) );
  NAND U5324 ( .A(n4282), .B(n4283), .Z(y[140]) );
  NAND U5325 ( .A(n3862), .B(m[140]), .Z(n4283) );
  NAND U5326 ( .A(n3863), .B(creg[140]), .Z(n4282) );
  NAND U5327 ( .A(n4284), .B(n4285), .Z(y[13]) );
  NAND U5328 ( .A(n3862), .B(m[13]), .Z(n4285) );
  NAND U5329 ( .A(n3863), .B(creg[13]), .Z(n4284) );
  NAND U5330 ( .A(n4286), .B(n4287), .Z(y[139]) );
  NAND U5331 ( .A(n3862), .B(m[139]), .Z(n4287) );
  NAND U5332 ( .A(n3863), .B(creg[139]), .Z(n4286) );
  NAND U5333 ( .A(n4288), .B(n4289), .Z(y[138]) );
  NAND U5334 ( .A(n3862), .B(m[138]), .Z(n4289) );
  NAND U5335 ( .A(n3863), .B(creg[138]), .Z(n4288) );
  NAND U5336 ( .A(n4290), .B(n4291), .Z(y[137]) );
  NAND U5337 ( .A(n3862), .B(m[137]), .Z(n4291) );
  NAND U5338 ( .A(n3863), .B(creg[137]), .Z(n4290) );
  NAND U5339 ( .A(n4292), .B(n4293), .Z(y[136]) );
  NAND U5340 ( .A(n3862), .B(m[136]), .Z(n4293) );
  NAND U5341 ( .A(n3863), .B(creg[136]), .Z(n4292) );
  NAND U5342 ( .A(n4294), .B(n4295), .Z(y[135]) );
  NAND U5343 ( .A(n3862), .B(m[135]), .Z(n4295) );
  NAND U5344 ( .A(n3863), .B(creg[135]), .Z(n4294) );
  NAND U5345 ( .A(n4296), .B(n4297), .Z(y[134]) );
  NAND U5346 ( .A(n3862), .B(m[134]), .Z(n4297) );
  NAND U5347 ( .A(n3863), .B(creg[134]), .Z(n4296) );
  NAND U5348 ( .A(n4298), .B(n4299), .Z(y[133]) );
  NAND U5349 ( .A(n3862), .B(m[133]), .Z(n4299) );
  NAND U5350 ( .A(n3863), .B(creg[133]), .Z(n4298) );
  NAND U5351 ( .A(n4300), .B(n4301), .Z(y[132]) );
  NAND U5352 ( .A(n3862), .B(m[132]), .Z(n4301) );
  NAND U5353 ( .A(n3863), .B(creg[132]), .Z(n4300) );
  NAND U5354 ( .A(n4302), .B(n4303), .Z(y[131]) );
  NAND U5355 ( .A(n3862), .B(m[131]), .Z(n4303) );
  NAND U5356 ( .A(n3863), .B(creg[131]), .Z(n4302) );
  NAND U5357 ( .A(n4304), .B(n4305), .Z(y[130]) );
  NAND U5358 ( .A(n3862), .B(m[130]), .Z(n4305) );
  NAND U5359 ( .A(n3863), .B(creg[130]), .Z(n4304) );
  NAND U5360 ( .A(n4306), .B(n4307), .Z(y[12]) );
  NAND U5361 ( .A(n3862), .B(m[12]), .Z(n4307) );
  NAND U5362 ( .A(n3863), .B(creg[12]), .Z(n4306) );
  NAND U5363 ( .A(n4308), .B(n4309), .Z(y[129]) );
  NAND U5364 ( .A(n3862), .B(m[129]), .Z(n4309) );
  NAND U5365 ( .A(n3863), .B(creg[129]), .Z(n4308) );
  NAND U5366 ( .A(n4310), .B(n4311), .Z(y[128]) );
  NAND U5367 ( .A(n3862), .B(m[128]), .Z(n4311) );
  NAND U5368 ( .A(n3863), .B(creg[128]), .Z(n4310) );
  NAND U5369 ( .A(n4312), .B(n4313), .Z(y[127]) );
  NAND U5370 ( .A(n3862), .B(m[127]), .Z(n4313) );
  NAND U5371 ( .A(n3863), .B(creg[127]), .Z(n4312) );
  NAND U5372 ( .A(n4314), .B(n4315), .Z(y[126]) );
  NAND U5373 ( .A(n3862), .B(m[126]), .Z(n4315) );
  NAND U5374 ( .A(n3863), .B(creg[126]), .Z(n4314) );
  NAND U5375 ( .A(n4316), .B(n4317), .Z(y[125]) );
  NAND U5376 ( .A(n3862), .B(m[125]), .Z(n4317) );
  NAND U5377 ( .A(n3863), .B(creg[125]), .Z(n4316) );
  NAND U5378 ( .A(n4318), .B(n4319), .Z(y[124]) );
  NAND U5379 ( .A(n3862), .B(m[124]), .Z(n4319) );
  NAND U5380 ( .A(n3863), .B(creg[124]), .Z(n4318) );
  NAND U5381 ( .A(n4320), .B(n4321), .Z(y[123]) );
  NAND U5382 ( .A(n3862), .B(m[123]), .Z(n4321) );
  NAND U5383 ( .A(n3863), .B(creg[123]), .Z(n4320) );
  NAND U5384 ( .A(n4322), .B(n4323), .Z(y[122]) );
  NAND U5385 ( .A(n3862), .B(m[122]), .Z(n4323) );
  NAND U5386 ( .A(n3863), .B(creg[122]), .Z(n4322) );
  NAND U5387 ( .A(n4324), .B(n4325), .Z(y[121]) );
  NAND U5388 ( .A(n3862), .B(m[121]), .Z(n4325) );
  NAND U5389 ( .A(n3863), .B(creg[121]), .Z(n4324) );
  NAND U5390 ( .A(n4326), .B(n4327), .Z(y[120]) );
  NAND U5391 ( .A(n3862), .B(m[120]), .Z(n4327) );
  NAND U5392 ( .A(n3863), .B(creg[120]), .Z(n4326) );
  NAND U5393 ( .A(n4328), .B(n4329), .Z(y[11]) );
  NAND U5394 ( .A(n3862), .B(m[11]), .Z(n4329) );
  NAND U5395 ( .A(n3863), .B(creg[11]), .Z(n4328) );
  NAND U5396 ( .A(n4330), .B(n4331), .Z(y[119]) );
  NAND U5397 ( .A(n3862), .B(m[119]), .Z(n4331) );
  NAND U5398 ( .A(n3863), .B(creg[119]), .Z(n4330) );
  NAND U5399 ( .A(n4332), .B(n4333), .Z(y[118]) );
  NAND U5400 ( .A(n3862), .B(m[118]), .Z(n4333) );
  NAND U5401 ( .A(n3863), .B(creg[118]), .Z(n4332) );
  NAND U5402 ( .A(n4334), .B(n4335), .Z(y[117]) );
  NAND U5403 ( .A(n3862), .B(m[117]), .Z(n4335) );
  NAND U5404 ( .A(n3863), .B(creg[117]), .Z(n4334) );
  NAND U5405 ( .A(n4336), .B(n4337), .Z(y[116]) );
  NAND U5406 ( .A(n3862), .B(m[116]), .Z(n4337) );
  NAND U5407 ( .A(n3863), .B(creg[116]), .Z(n4336) );
  NAND U5408 ( .A(n4338), .B(n4339), .Z(y[115]) );
  NAND U5409 ( .A(n3862), .B(m[115]), .Z(n4339) );
  NAND U5410 ( .A(n3863), .B(creg[115]), .Z(n4338) );
  NAND U5411 ( .A(n4340), .B(n4341), .Z(y[114]) );
  NAND U5412 ( .A(n3862), .B(m[114]), .Z(n4341) );
  NAND U5413 ( .A(n3863), .B(creg[114]), .Z(n4340) );
  NAND U5414 ( .A(n4342), .B(n4343), .Z(y[113]) );
  NAND U5415 ( .A(n3862), .B(m[113]), .Z(n4343) );
  NAND U5416 ( .A(n3863), .B(creg[113]), .Z(n4342) );
  NAND U5417 ( .A(n4344), .B(n4345), .Z(y[112]) );
  NAND U5418 ( .A(n3862), .B(m[112]), .Z(n4345) );
  NAND U5419 ( .A(n3863), .B(creg[112]), .Z(n4344) );
  NAND U5420 ( .A(n4346), .B(n4347), .Z(y[111]) );
  NAND U5421 ( .A(n3862), .B(m[111]), .Z(n4347) );
  NAND U5422 ( .A(n3863), .B(creg[111]), .Z(n4346) );
  NAND U5423 ( .A(n4348), .B(n4349), .Z(y[110]) );
  NAND U5424 ( .A(n3862), .B(m[110]), .Z(n4349) );
  NAND U5425 ( .A(n3863), .B(creg[110]), .Z(n4348) );
  NAND U5426 ( .A(n4350), .B(n4351), .Z(y[10]) );
  NAND U5427 ( .A(n3862), .B(m[10]), .Z(n4351) );
  NAND U5428 ( .A(n3863), .B(creg[10]), .Z(n4350) );
  NAND U5429 ( .A(n4352), .B(n4353), .Z(y[109]) );
  NAND U5430 ( .A(n3862), .B(m[109]), .Z(n4353) );
  NAND U5431 ( .A(n3863), .B(creg[109]), .Z(n4352) );
  NAND U5432 ( .A(n4354), .B(n4355), .Z(y[108]) );
  NAND U5433 ( .A(n3862), .B(m[108]), .Z(n4355) );
  NAND U5434 ( .A(n3863), .B(creg[108]), .Z(n4354) );
  NAND U5435 ( .A(n4356), .B(n4357), .Z(y[107]) );
  NAND U5436 ( .A(n3862), .B(m[107]), .Z(n4357) );
  NAND U5437 ( .A(n3863), .B(creg[107]), .Z(n4356) );
  NAND U5438 ( .A(n4358), .B(n4359), .Z(y[106]) );
  NAND U5439 ( .A(n3862), .B(m[106]), .Z(n4359) );
  NAND U5440 ( .A(n3863), .B(creg[106]), .Z(n4358) );
  NAND U5441 ( .A(n4360), .B(n4361), .Z(y[105]) );
  NAND U5442 ( .A(n3862), .B(m[105]), .Z(n4361) );
  NAND U5443 ( .A(n3863), .B(creg[105]), .Z(n4360) );
  NAND U5444 ( .A(n4362), .B(n4363), .Z(y[104]) );
  NAND U5445 ( .A(n3862), .B(m[104]), .Z(n4363) );
  NAND U5446 ( .A(n3863), .B(creg[104]), .Z(n4362) );
  NAND U5447 ( .A(n4364), .B(n4365), .Z(y[103]) );
  NAND U5448 ( .A(n3862), .B(m[103]), .Z(n4365) );
  NAND U5449 ( .A(n3863), .B(creg[103]), .Z(n4364) );
  NAND U5450 ( .A(n4366), .B(n4367), .Z(y[102]) );
  NAND U5451 ( .A(n3862), .B(m[102]), .Z(n4367) );
  NAND U5452 ( .A(n3863), .B(creg[102]), .Z(n4366) );
  NAND U5453 ( .A(n4368), .B(n4369), .Z(y[101]) );
  NAND U5454 ( .A(n3862), .B(m[101]), .Z(n4369) );
  NAND U5455 ( .A(n3863), .B(creg[101]), .Z(n4368) );
  NAND U5456 ( .A(n4370), .B(n4371), .Z(y[100]) );
  NAND U5457 ( .A(n3862), .B(m[100]), .Z(n4371) );
  NAND U5458 ( .A(n3863), .B(creg[100]), .Z(n4370) );
  NAND U5459 ( .A(n4372), .B(n4373), .Z(y[0]) );
  NAND U5460 ( .A(n3862), .B(m[0]), .Z(n4373) );
  NAND U5461 ( .A(n3863), .B(creg[0]), .Z(n4372) );
  NAND U5462 ( .A(n4374), .B(n4375), .Z(x[9]) );
  NAND U5463 ( .A(creg[9]), .B(init), .Z(n4374) );
  NAND U5464 ( .A(n4376), .B(n4377), .Z(x[99]) );
  NAND U5465 ( .A(creg[99]), .B(init), .Z(n4376) );
  NAND U5466 ( .A(n4378), .B(n4379), .Z(x[98]) );
  NAND U5467 ( .A(creg[98]), .B(init), .Z(n4378) );
  NAND U5468 ( .A(n4380), .B(n4381), .Z(x[97]) );
  NAND U5469 ( .A(creg[97]), .B(init), .Z(n4380) );
  NAND U5470 ( .A(n4382), .B(n4383), .Z(x[96]) );
  NAND U5471 ( .A(creg[96]), .B(init), .Z(n4382) );
  NAND U5472 ( .A(n4384), .B(n4385), .Z(x[95]) );
  NAND U5473 ( .A(creg[95]), .B(init), .Z(n4384) );
  NAND U5474 ( .A(n4386), .B(n4387), .Z(x[94]) );
  NAND U5475 ( .A(creg[94]), .B(init), .Z(n4386) );
  NAND U5476 ( .A(n4388), .B(n4389), .Z(x[93]) );
  NAND U5477 ( .A(creg[93]), .B(init), .Z(n4388) );
  NAND U5478 ( .A(n4390), .B(n4391), .Z(x[92]) );
  NAND U5479 ( .A(creg[92]), .B(init), .Z(n4390) );
  NAND U5480 ( .A(n4392), .B(n4393), .Z(x[91]) );
  NAND U5481 ( .A(creg[91]), .B(init), .Z(n4392) );
  NAND U5482 ( .A(n4394), .B(n4395), .Z(x[90]) );
  NAND U5483 ( .A(creg[90]), .B(init), .Z(n4394) );
  NAND U5484 ( .A(n4396), .B(n4397), .Z(x[8]) );
  NAND U5485 ( .A(creg[8]), .B(init), .Z(n4396) );
  NAND U5486 ( .A(n4398), .B(n4399), .Z(x[89]) );
  NAND U5487 ( .A(creg[89]), .B(init), .Z(n4398) );
  NAND U5488 ( .A(n4400), .B(n4401), .Z(x[88]) );
  NAND U5489 ( .A(creg[88]), .B(init), .Z(n4400) );
  NAND U5490 ( .A(n4402), .B(n4403), .Z(x[87]) );
  NAND U5491 ( .A(creg[87]), .B(init), .Z(n4402) );
  NAND U5492 ( .A(n4404), .B(n4405), .Z(x[86]) );
  NAND U5493 ( .A(creg[86]), .B(init), .Z(n4404) );
  NAND U5494 ( .A(n4406), .B(n4407), .Z(x[85]) );
  NAND U5495 ( .A(creg[85]), .B(init), .Z(n4406) );
  NAND U5496 ( .A(n4408), .B(n4409), .Z(x[84]) );
  NAND U5497 ( .A(creg[84]), .B(init), .Z(n4408) );
  NAND U5498 ( .A(n4410), .B(n4411), .Z(x[83]) );
  NAND U5499 ( .A(creg[83]), .B(init), .Z(n4410) );
  NAND U5500 ( .A(n4412), .B(n4413), .Z(x[82]) );
  NAND U5501 ( .A(creg[82]), .B(init), .Z(n4412) );
  NAND U5502 ( .A(n4414), .B(n4415), .Z(x[81]) );
  NAND U5503 ( .A(creg[81]), .B(init), .Z(n4414) );
  NAND U5504 ( .A(n4416), .B(n4417), .Z(x[80]) );
  NAND U5505 ( .A(creg[80]), .B(init), .Z(n4416) );
  NAND U5506 ( .A(n4418), .B(n4419), .Z(x[7]) );
  NAND U5507 ( .A(creg[7]), .B(init), .Z(n4418) );
  NAND U5508 ( .A(n4420), .B(n4421), .Z(x[79]) );
  NAND U5509 ( .A(creg[79]), .B(init), .Z(n4420) );
  NAND U5510 ( .A(n4422), .B(n4423), .Z(x[78]) );
  NAND U5511 ( .A(creg[78]), .B(init), .Z(n4422) );
  NAND U5512 ( .A(n4424), .B(n4425), .Z(x[77]) );
  NAND U5513 ( .A(creg[77]), .B(init), .Z(n4424) );
  NAND U5514 ( .A(n4426), .B(n4427), .Z(x[76]) );
  NAND U5515 ( .A(creg[76]), .B(init), .Z(n4426) );
  NAND U5516 ( .A(n4428), .B(n4429), .Z(x[75]) );
  NAND U5517 ( .A(creg[75]), .B(init), .Z(n4428) );
  NAND U5518 ( .A(n4430), .B(n4431), .Z(x[74]) );
  NAND U5519 ( .A(creg[74]), .B(init), .Z(n4430) );
  NAND U5520 ( .A(n4432), .B(n4433), .Z(x[73]) );
  NAND U5521 ( .A(creg[73]), .B(init), .Z(n4432) );
  NAND U5522 ( .A(n4434), .B(n4435), .Z(x[72]) );
  NAND U5523 ( .A(creg[72]), .B(init), .Z(n4434) );
  NAND U5524 ( .A(n4436), .B(n4437), .Z(x[71]) );
  NAND U5525 ( .A(creg[71]), .B(init), .Z(n4436) );
  NAND U5526 ( .A(n4438), .B(n4439), .Z(x[70]) );
  NAND U5527 ( .A(creg[70]), .B(init), .Z(n4438) );
  NAND U5528 ( .A(n4440), .B(n4441), .Z(x[6]) );
  NAND U5529 ( .A(creg[6]), .B(init), .Z(n4440) );
  NAND U5530 ( .A(n4442), .B(n4443), .Z(x[69]) );
  NAND U5531 ( .A(creg[69]), .B(init), .Z(n4442) );
  NAND U5532 ( .A(n4444), .B(n4445), .Z(x[68]) );
  NAND U5533 ( .A(creg[68]), .B(init), .Z(n4444) );
  NAND U5534 ( .A(n4446), .B(n4447), .Z(x[67]) );
  NAND U5535 ( .A(creg[67]), .B(init), .Z(n4446) );
  NAND U5536 ( .A(n4448), .B(n4449), .Z(x[66]) );
  NAND U5537 ( .A(creg[66]), .B(init), .Z(n4448) );
  NAND U5538 ( .A(n4450), .B(n4451), .Z(x[65]) );
  NAND U5539 ( .A(creg[65]), .B(init), .Z(n4450) );
  NAND U5540 ( .A(n4452), .B(n4453), .Z(x[64]) );
  NAND U5541 ( .A(creg[64]), .B(init), .Z(n4452) );
  NAND U5542 ( .A(n4454), .B(n4455), .Z(x[63]) );
  NAND U5543 ( .A(creg[63]), .B(init), .Z(n4454) );
  NAND U5544 ( .A(n4456), .B(n4457), .Z(x[62]) );
  NAND U5545 ( .A(creg[62]), .B(init), .Z(n4456) );
  NAND U5546 ( .A(n4458), .B(n4459), .Z(x[61]) );
  NAND U5547 ( .A(creg[61]), .B(init), .Z(n4458) );
  NAND U5548 ( .A(n4460), .B(n4461), .Z(x[60]) );
  NAND U5549 ( .A(creg[60]), .B(init), .Z(n4460) );
  NAND U5550 ( .A(n4462), .B(n4463), .Z(x[5]) );
  NAND U5551 ( .A(creg[5]), .B(init), .Z(n4462) );
  NAND U5552 ( .A(n4464), .B(n4465), .Z(x[59]) );
  NAND U5553 ( .A(creg[59]), .B(init), .Z(n4464) );
  NAND U5554 ( .A(n4466), .B(n4467), .Z(x[58]) );
  NAND U5555 ( .A(creg[58]), .B(init), .Z(n4466) );
  NAND U5556 ( .A(n4468), .B(n4469), .Z(x[57]) );
  NAND U5557 ( .A(creg[57]), .B(init), .Z(n4468) );
  NAND U5558 ( .A(n4470), .B(n4471), .Z(x[56]) );
  NAND U5559 ( .A(creg[56]), .B(init), .Z(n4470) );
  NAND U5560 ( .A(n4472), .B(n4473), .Z(x[55]) );
  NAND U5561 ( .A(creg[55]), .B(init), .Z(n4472) );
  NAND U5562 ( .A(n4474), .B(n4475), .Z(x[54]) );
  NAND U5563 ( .A(creg[54]), .B(init), .Z(n4474) );
  NAND U5564 ( .A(n4476), .B(n4477), .Z(x[53]) );
  NAND U5565 ( .A(creg[53]), .B(init), .Z(n4476) );
  NAND U5566 ( .A(n4478), .B(n4479), .Z(x[52]) );
  NAND U5567 ( .A(creg[52]), .B(init), .Z(n4478) );
  NAND U5568 ( .A(n4480), .B(n4481), .Z(x[51]) );
  NAND U5569 ( .A(creg[51]), .B(init), .Z(n4480) );
  NAND U5570 ( .A(n4482), .B(n4483), .Z(x[50]) );
  NAND U5571 ( .A(creg[50]), .B(init), .Z(n4482) );
  NAND U5572 ( .A(n4484), .B(n4485), .Z(x[4]) );
  NAND U5573 ( .A(creg[4]), .B(init), .Z(n4484) );
  NAND U5574 ( .A(n4486), .B(n4487), .Z(x[49]) );
  NAND U5575 ( .A(creg[49]), .B(init), .Z(n4486) );
  NAND U5576 ( .A(n4488), .B(n4489), .Z(x[48]) );
  NAND U5577 ( .A(creg[48]), .B(init), .Z(n4488) );
  NAND U5578 ( .A(n4490), .B(n4491), .Z(x[47]) );
  NAND U5579 ( .A(creg[47]), .B(init), .Z(n4490) );
  NAND U5580 ( .A(n4492), .B(n4493), .Z(x[46]) );
  NAND U5581 ( .A(creg[46]), .B(init), .Z(n4492) );
  NAND U5582 ( .A(n4494), .B(n4495), .Z(x[45]) );
  NAND U5583 ( .A(creg[45]), .B(init), .Z(n4494) );
  NAND U5584 ( .A(n4496), .B(n4497), .Z(x[44]) );
  NAND U5585 ( .A(creg[44]), .B(init), .Z(n4496) );
  NAND U5586 ( .A(n4498), .B(n4499), .Z(x[43]) );
  NAND U5587 ( .A(creg[43]), .B(init), .Z(n4498) );
  NAND U5588 ( .A(n4500), .B(n4501), .Z(x[42]) );
  NAND U5589 ( .A(creg[42]), .B(init), .Z(n4500) );
  NAND U5590 ( .A(n4502), .B(n4503), .Z(x[41]) );
  NAND U5591 ( .A(creg[41]), .B(init), .Z(n4502) );
  NAND U5592 ( .A(n4504), .B(n4505), .Z(x[40]) );
  NAND U5593 ( .A(creg[40]), .B(init), .Z(n4504) );
  NAND U5594 ( .A(n4506), .B(n4507), .Z(x[3]) );
  NAND U5595 ( .A(creg[3]), .B(init), .Z(n4506) );
  NAND U5596 ( .A(n4508), .B(n4509), .Z(x[39]) );
  NAND U5597 ( .A(creg[39]), .B(init), .Z(n4508) );
  NAND U5598 ( .A(n4510), .B(n4511), .Z(x[38]) );
  NAND U5599 ( .A(creg[38]), .B(init), .Z(n4510) );
  NAND U5600 ( .A(n4512), .B(n4513), .Z(x[37]) );
  NAND U5601 ( .A(creg[37]), .B(init), .Z(n4512) );
  NAND U5602 ( .A(n4514), .B(n4515), .Z(x[36]) );
  NAND U5603 ( .A(creg[36]), .B(init), .Z(n4514) );
  NAND U5604 ( .A(n4516), .B(n4517), .Z(x[35]) );
  NAND U5605 ( .A(creg[35]), .B(init), .Z(n4516) );
  NAND U5606 ( .A(n4518), .B(n4519), .Z(x[34]) );
  NAND U5607 ( .A(creg[34]), .B(init), .Z(n4518) );
  NAND U5608 ( .A(n4520), .B(n4521), .Z(x[33]) );
  NAND U5609 ( .A(creg[33]), .B(init), .Z(n4520) );
  NAND U5610 ( .A(n4522), .B(n4523), .Z(x[32]) );
  NAND U5611 ( .A(creg[32]), .B(init), .Z(n4522) );
  NAND U5612 ( .A(n4524), .B(n4525), .Z(x[31]) );
  NAND U5613 ( .A(creg[31]), .B(init), .Z(n4524) );
  NAND U5614 ( .A(n4526), .B(n4527), .Z(x[30]) );
  NAND U5615 ( .A(creg[30]), .B(init), .Z(n4526) );
  NAND U5616 ( .A(n4528), .B(n4529), .Z(x[2]) );
  NAND U5617 ( .A(creg[2]), .B(init), .Z(n4528) );
  NAND U5618 ( .A(n4530), .B(n4531), .Z(x[29]) );
  NAND U5619 ( .A(creg[29]), .B(init), .Z(n4530) );
  NAND U5620 ( .A(n4532), .B(n4533), .Z(x[28]) );
  NAND U5621 ( .A(creg[28]), .B(init), .Z(n4532) );
  NAND U5622 ( .A(n4534), .B(n4535), .Z(x[27]) );
  NAND U5623 ( .A(creg[27]), .B(init), .Z(n4534) );
  NAND U5624 ( .A(n4536), .B(n4537), .Z(x[26]) );
  NAND U5625 ( .A(creg[26]), .B(init), .Z(n4536) );
  NAND U5626 ( .A(n4538), .B(n4539), .Z(x[25]) );
  NAND U5627 ( .A(creg[25]), .B(init), .Z(n4538) );
  NAND U5628 ( .A(n4540), .B(n4541), .Z(x[255]) );
  NAND U5629 ( .A(creg[255]), .B(init), .Z(n4540) );
  NAND U5630 ( .A(n4542), .B(n4543), .Z(x[254]) );
  NAND U5631 ( .A(creg[254]), .B(init), .Z(n4542) );
  NAND U5632 ( .A(n4544), .B(n4545), .Z(x[253]) );
  NAND U5633 ( .A(creg[253]), .B(init), .Z(n4544) );
  NAND U5634 ( .A(n4546), .B(n4547), .Z(x[252]) );
  NAND U5635 ( .A(creg[252]), .B(init), .Z(n4546) );
  NAND U5636 ( .A(n4548), .B(n4549), .Z(x[251]) );
  NAND U5637 ( .A(creg[251]), .B(init), .Z(n4548) );
  NAND U5638 ( .A(n4550), .B(n4551), .Z(x[250]) );
  NAND U5639 ( .A(creg[250]), .B(init), .Z(n4550) );
  NAND U5640 ( .A(n4552), .B(n4553), .Z(x[24]) );
  NAND U5641 ( .A(creg[24]), .B(init), .Z(n4552) );
  NAND U5642 ( .A(n4554), .B(n4555), .Z(x[249]) );
  NAND U5643 ( .A(creg[249]), .B(init), .Z(n4554) );
  NAND U5644 ( .A(n4556), .B(n4557), .Z(x[248]) );
  NAND U5645 ( .A(creg[248]), .B(init), .Z(n4556) );
  NAND U5646 ( .A(n4558), .B(n4559), .Z(x[247]) );
  NAND U5647 ( .A(creg[247]), .B(init), .Z(n4558) );
  NAND U5648 ( .A(n4560), .B(n4561), .Z(x[246]) );
  NAND U5649 ( .A(creg[246]), .B(init), .Z(n4560) );
  NAND U5650 ( .A(n4562), .B(n4563), .Z(x[245]) );
  NAND U5651 ( .A(creg[245]), .B(init), .Z(n4562) );
  NAND U5652 ( .A(n4564), .B(n4565), .Z(x[244]) );
  NAND U5653 ( .A(creg[244]), .B(init), .Z(n4564) );
  NAND U5654 ( .A(n4566), .B(n4567), .Z(x[243]) );
  NAND U5655 ( .A(creg[243]), .B(init), .Z(n4566) );
  NAND U5656 ( .A(n4568), .B(n4569), .Z(x[242]) );
  NAND U5657 ( .A(creg[242]), .B(init), .Z(n4568) );
  NAND U5658 ( .A(n4570), .B(n4571), .Z(x[241]) );
  NAND U5659 ( .A(creg[241]), .B(init), .Z(n4570) );
  NAND U5660 ( .A(n4572), .B(n4573), .Z(x[240]) );
  NAND U5661 ( .A(creg[240]), .B(init), .Z(n4572) );
  NAND U5662 ( .A(n4574), .B(n4575), .Z(x[23]) );
  NAND U5663 ( .A(creg[23]), .B(init), .Z(n4574) );
  NAND U5664 ( .A(n4576), .B(n4577), .Z(x[239]) );
  NAND U5665 ( .A(creg[239]), .B(init), .Z(n4576) );
  NAND U5666 ( .A(n4578), .B(n4579), .Z(x[238]) );
  NAND U5667 ( .A(creg[238]), .B(init), .Z(n4578) );
  NAND U5668 ( .A(n4580), .B(n4581), .Z(x[237]) );
  NAND U5669 ( .A(creg[237]), .B(init), .Z(n4580) );
  NAND U5670 ( .A(n4582), .B(n4583), .Z(x[236]) );
  NAND U5671 ( .A(creg[236]), .B(init), .Z(n4582) );
  NAND U5672 ( .A(n4584), .B(n4585), .Z(x[235]) );
  NAND U5673 ( .A(creg[235]), .B(init), .Z(n4584) );
  NAND U5674 ( .A(n4586), .B(n4587), .Z(x[234]) );
  NAND U5675 ( .A(creg[234]), .B(init), .Z(n4586) );
  NAND U5676 ( .A(n4588), .B(n4589), .Z(x[233]) );
  NAND U5677 ( .A(creg[233]), .B(init), .Z(n4588) );
  NAND U5678 ( .A(n4590), .B(n4591), .Z(x[232]) );
  NAND U5679 ( .A(creg[232]), .B(init), .Z(n4590) );
  NAND U5680 ( .A(n4592), .B(n4593), .Z(x[231]) );
  NAND U5681 ( .A(creg[231]), .B(init), .Z(n4592) );
  NAND U5682 ( .A(n4594), .B(n4595), .Z(x[230]) );
  NAND U5683 ( .A(creg[230]), .B(init), .Z(n4594) );
  NAND U5684 ( .A(n4596), .B(n4597), .Z(x[22]) );
  NAND U5685 ( .A(creg[22]), .B(init), .Z(n4596) );
  NAND U5686 ( .A(n4598), .B(n4599), .Z(x[229]) );
  NAND U5687 ( .A(creg[229]), .B(init), .Z(n4598) );
  NAND U5688 ( .A(n4600), .B(n4601), .Z(x[228]) );
  NAND U5689 ( .A(creg[228]), .B(init), .Z(n4600) );
  NAND U5690 ( .A(n4602), .B(n4603), .Z(x[227]) );
  NAND U5691 ( .A(creg[227]), .B(init), .Z(n4602) );
  NAND U5692 ( .A(n4604), .B(n4605), .Z(x[226]) );
  NAND U5693 ( .A(creg[226]), .B(init), .Z(n4604) );
  NAND U5694 ( .A(n4606), .B(n4607), .Z(x[225]) );
  NAND U5695 ( .A(creg[225]), .B(init), .Z(n4606) );
  NAND U5696 ( .A(n4608), .B(n4609), .Z(x[224]) );
  NAND U5697 ( .A(creg[224]), .B(init), .Z(n4608) );
  NAND U5698 ( .A(n4610), .B(n4611), .Z(x[223]) );
  NAND U5699 ( .A(creg[223]), .B(init), .Z(n4610) );
  NAND U5700 ( .A(n4612), .B(n4613), .Z(x[222]) );
  NAND U5701 ( .A(creg[222]), .B(init), .Z(n4612) );
  NAND U5702 ( .A(n4614), .B(n4615), .Z(x[221]) );
  NAND U5703 ( .A(creg[221]), .B(init), .Z(n4614) );
  NAND U5704 ( .A(n4616), .B(n4617), .Z(x[220]) );
  NAND U5705 ( .A(creg[220]), .B(init), .Z(n4616) );
  NAND U5706 ( .A(n4618), .B(n4619), .Z(x[21]) );
  NAND U5707 ( .A(creg[21]), .B(init), .Z(n4618) );
  NAND U5708 ( .A(n4620), .B(n4621), .Z(x[219]) );
  NAND U5709 ( .A(creg[219]), .B(init), .Z(n4620) );
  NAND U5710 ( .A(n4622), .B(n4623), .Z(x[218]) );
  NAND U5711 ( .A(creg[218]), .B(init), .Z(n4622) );
  NAND U5712 ( .A(n4624), .B(n4625), .Z(x[217]) );
  NAND U5713 ( .A(creg[217]), .B(init), .Z(n4624) );
  NAND U5714 ( .A(n4626), .B(n4627), .Z(x[216]) );
  NAND U5715 ( .A(creg[216]), .B(init), .Z(n4626) );
  NAND U5716 ( .A(n4628), .B(n4629), .Z(x[215]) );
  NAND U5717 ( .A(creg[215]), .B(init), .Z(n4628) );
  NAND U5718 ( .A(n4630), .B(n4631), .Z(x[214]) );
  NAND U5719 ( .A(creg[214]), .B(init), .Z(n4630) );
  NAND U5720 ( .A(n4632), .B(n4633), .Z(x[213]) );
  NAND U5721 ( .A(creg[213]), .B(init), .Z(n4632) );
  NAND U5722 ( .A(n4634), .B(n4635), .Z(x[212]) );
  NAND U5723 ( .A(creg[212]), .B(init), .Z(n4634) );
  NAND U5724 ( .A(n4636), .B(n4637), .Z(x[211]) );
  NAND U5725 ( .A(creg[211]), .B(init), .Z(n4636) );
  NAND U5726 ( .A(n4638), .B(n4639), .Z(x[210]) );
  NAND U5727 ( .A(creg[210]), .B(init), .Z(n4638) );
  NAND U5728 ( .A(n4640), .B(n4641), .Z(x[20]) );
  NAND U5729 ( .A(creg[20]), .B(init), .Z(n4640) );
  NAND U5730 ( .A(n4642), .B(n4643), .Z(x[209]) );
  NAND U5731 ( .A(creg[209]), .B(init), .Z(n4642) );
  NAND U5732 ( .A(n4644), .B(n4645), .Z(x[208]) );
  NAND U5733 ( .A(creg[208]), .B(init), .Z(n4644) );
  NAND U5734 ( .A(n4646), .B(n4647), .Z(x[207]) );
  NAND U5735 ( .A(creg[207]), .B(init), .Z(n4646) );
  NAND U5736 ( .A(n4648), .B(n4649), .Z(x[206]) );
  NAND U5737 ( .A(creg[206]), .B(init), .Z(n4648) );
  NAND U5738 ( .A(n4650), .B(n4651), .Z(x[205]) );
  NAND U5739 ( .A(creg[205]), .B(init), .Z(n4650) );
  NAND U5740 ( .A(n4652), .B(n4653), .Z(x[204]) );
  NAND U5741 ( .A(creg[204]), .B(init), .Z(n4652) );
  NAND U5742 ( .A(n4654), .B(n4655), .Z(x[203]) );
  NAND U5743 ( .A(creg[203]), .B(init), .Z(n4654) );
  NAND U5744 ( .A(n4656), .B(n4657), .Z(x[202]) );
  NAND U5745 ( .A(creg[202]), .B(init), .Z(n4656) );
  NAND U5746 ( .A(n4658), .B(n4659), .Z(x[201]) );
  NAND U5747 ( .A(creg[201]), .B(init), .Z(n4658) );
  NAND U5748 ( .A(n4660), .B(n4661), .Z(x[200]) );
  NAND U5749 ( .A(creg[200]), .B(init), .Z(n4660) );
  NAND U5750 ( .A(n4662), .B(n4663), .Z(x[1]) );
  NAND U5751 ( .A(creg[1]), .B(init), .Z(n4662) );
  NAND U5752 ( .A(n4664), .B(n4665), .Z(x[19]) );
  NAND U5753 ( .A(creg[19]), .B(init), .Z(n4664) );
  NAND U5754 ( .A(n4666), .B(n4667), .Z(x[199]) );
  NAND U5755 ( .A(creg[199]), .B(init), .Z(n4666) );
  NAND U5756 ( .A(n4668), .B(n4669), .Z(x[198]) );
  NAND U5757 ( .A(creg[198]), .B(init), .Z(n4668) );
  NAND U5758 ( .A(n4670), .B(n4671), .Z(x[197]) );
  NAND U5759 ( .A(creg[197]), .B(init), .Z(n4670) );
  NAND U5760 ( .A(n4672), .B(n4673), .Z(x[196]) );
  NAND U5761 ( .A(creg[196]), .B(init), .Z(n4672) );
  NAND U5762 ( .A(n4674), .B(n4675), .Z(x[195]) );
  NAND U5763 ( .A(creg[195]), .B(init), .Z(n4674) );
  NAND U5764 ( .A(n4676), .B(n4677), .Z(x[194]) );
  NAND U5765 ( .A(creg[194]), .B(init), .Z(n4676) );
  NAND U5766 ( .A(n4678), .B(n4679), .Z(x[193]) );
  NAND U5767 ( .A(creg[193]), .B(init), .Z(n4678) );
  NAND U5768 ( .A(n4680), .B(n4681), .Z(x[192]) );
  NAND U5769 ( .A(creg[192]), .B(init), .Z(n4680) );
  NAND U5770 ( .A(n4682), .B(n4683), .Z(x[191]) );
  NAND U5771 ( .A(creg[191]), .B(init), .Z(n4682) );
  NAND U5772 ( .A(n4684), .B(n4685), .Z(x[190]) );
  NAND U5773 ( .A(creg[190]), .B(init), .Z(n4684) );
  NAND U5774 ( .A(n4686), .B(n4687), .Z(x[18]) );
  NAND U5775 ( .A(creg[18]), .B(init), .Z(n4686) );
  NAND U5776 ( .A(n4688), .B(n4689), .Z(x[189]) );
  NAND U5777 ( .A(creg[189]), .B(init), .Z(n4688) );
  NAND U5778 ( .A(n4690), .B(n4691), .Z(x[188]) );
  NAND U5779 ( .A(creg[188]), .B(init), .Z(n4690) );
  NAND U5780 ( .A(n4692), .B(n4693), .Z(x[187]) );
  NAND U5781 ( .A(creg[187]), .B(init), .Z(n4692) );
  NAND U5782 ( .A(n4694), .B(n4695), .Z(x[186]) );
  NAND U5783 ( .A(creg[186]), .B(init), .Z(n4694) );
  NAND U5784 ( .A(n4696), .B(n4697), .Z(x[185]) );
  NAND U5785 ( .A(creg[185]), .B(init), .Z(n4696) );
  NAND U5786 ( .A(n4698), .B(n4699), .Z(x[184]) );
  NAND U5787 ( .A(creg[184]), .B(init), .Z(n4698) );
  NAND U5788 ( .A(n4700), .B(n4701), .Z(x[183]) );
  NAND U5789 ( .A(creg[183]), .B(init), .Z(n4700) );
  NAND U5790 ( .A(n4702), .B(n4703), .Z(x[182]) );
  NAND U5791 ( .A(creg[182]), .B(init), .Z(n4702) );
  NAND U5792 ( .A(n4704), .B(n4705), .Z(x[181]) );
  NAND U5793 ( .A(creg[181]), .B(init), .Z(n4704) );
  NAND U5794 ( .A(n4706), .B(n4707), .Z(x[180]) );
  NAND U5795 ( .A(creg[180]), .B(init), .Z(n4706) );
  NAND U5796 ( .A(n4708), .B(n4709), .Z(x[17]) );
  NAND U5797 ( .A(creg[17]), .B(init), .Z(n4708) );
  NAND U5798 ( .A(n4710), .B(n4711), .Z(x[179]) );
  NAND U5799 ( .A(creg[179]), .B(init), .Z(n4710) );
  NAND U5800 ( .A(n4712), .B(n4713), .Z(x[178]) );
  NAND U5801 ( .A(creg[178]), .B(init), .Z(n4712) );
  NAND U5802 ( .A(n4714), .B(n4715), .Z(x[177]) );
  NAND U5803 ( .A(creg[177]), .B(init), .Z(n4714) );
  NAND U5804 ( .A(n4716), .B(n4717), .Z(x[176]) );
  NAND U5805 ( .A(creg[176]), .B(init), .Z(n4716) );
  NAND U5806 ( .A(n4718), .B(n4719), .Z(x[175]) );
  NAND U5807 ( .A(creg[175]), .B(init), .Z(n4718) );
  NAND U5808 ( .A(n4720), .B(n4721), .Z(x[174]) );
  NAND U5809 ( .A(creg[174]), .B(init), .Z(n4720) );
  NAND U5810 ( .A(n4722), .B(n4723), .Z(x[173]) );
  NAND U5811 ( .A(creg[173]), .B(init), .Z(n4722) );
  NAND U5812 ( .A(n4724), .B(n4725), .Z(x[172]) );
  NAND U5813 ( .A(creg[172]), .B(init), .Z(n4724) );
  NAND U5814 ( .A(n4726), .B(n4727), .Z(x[171]) );
  NAND U5815 ( .A(creg[171]), .B(init), .Z(n4726) );
  NAND U5816 ( .A(n4728), .B(n4729), .Z(x[170]) );
  NAND U5817 ( .A(creg[170]), .B(init), .Z(n4728) );
  NAND U5818 ( .A(n4730), .B(n4731), .Z(x[16]) );
  NAND U5819 ( .A(creg[16]), .B(init), .Z(n4730) );
  NAND U5820 ( .A(n4732), .B(n4733), .Z(x[169]) );
  NAND U5821 ( .A(creg[169]), .B(init), .Z(n4732) );
  NAND U5822 ( .A(n4734), .B(n4735), .Z(x[168]) );
  NAND U5823 ( .A(creg[168]), .B(init), .Z(n4734) );
  NAND U5824 ( .A(n4736), .B(n4737), .Z(x[167]) );
  NAND U5825 ( .A(creg[167]), .B(init), .Z(n4736) );
  NAND U5826 ( .A(n4738), .B(n4739), .Z(x[166]) );
  NAND U5827 ( .A(creg[166]), .B(init), .Z(n4738) );
  NAND U5828 ( .A(n4740), .B(n4741), .Z(x[165]) );
  NAND U5829 ( .A(creg[165]), .B(init), .Z(n4740) );
  NAND U5830 ( .A(n4742), .B(n4743), .Z(x[164]) );
  NAND U5831 ( .A(creg[164]), .B(init), .Z(n4742) );
  NAND U5832 ( .A(n4744), .B(n4745), .Z(x[163]) );
  NAND U5833 ( .A(creg[163]), .B(init), .Z(n4744) );
  NAND U5834 ( .A(n4746), .B(n4747), .Z(x[162]) );
  NAND U5835 ( .A(creg[162]), .B(init), .Z(n4746) );
  NAND U5836 ( .A(n4748), .B(n4749), .Z(x[161]) );
  NAND U5837 ( .A(creg[161]), .B(init), .Z(n4748) );
  NAND U5838 ( .A(n4750), .B(n4751), .Z(x[160]) );
  NAND U5839 ( .A(creg[160]), .B(init), .Z(n4750) );
  NAND U5840 ( .A(n4752), .B(n4753), .Z(x[15]) );
  NAND U5841 ( .A(creg[15]), .B(init), .Z(n4752) );
  NAND U5842 ( .A(n4754), .B(n4755), .Z(x[159]) );
  NAND U5843 ( .A(creg[159]), .B(init), .Z(n4754) );
  NAND U5844 ( .A(n4756), .B(n4757), .Z(x[158]) );
  NAND U5845 ( .A(creg[158]), .B(init), .Z(n4756) );
  NAND U5846 ( .A(n4758), .B(n4759), .Z(x[157]) );
  NAND U5847 ( .A(creg[157]), .B(init), .Z(n4758) );
  NAND U5848 ( .A(n4760), .B(n4761), .Z(x[156]) );
  NAND U5849 ( .A(creg[156]), .B(init), .Z(n4760) );
  NAND U5850 ( .A(n4762), .B(n4763), .Z(x[155]) );
  NAND U5851 ( .A(creg[155]), .B(init), .Z(n4762) );
  NAND U5852 ( .A(n4764), .B(n4765), .Z(x[154]) );
  NAND U5853 ( .A(creg[154]), .B(init), .Z(n4764) );
  NAND U5854 ( .A(n4766), .B(n4767), .Z(x[153]) );
  NAND U5855 ( .A(creg[153]), .B(init), .Z(n4766) );
  NAND U5856 ( .A(n4768), .B(n4769), .Z(x[152]) );
  NAND U5857 ( .A(creg[152]), .B(init), .Z(n4768) );
  NAND U5858 ( .A(n4770), .B(n4771), .Z(x[151]) );
  NAND U5859 ( .A(creg[151]), .B(init), .Z(n4770) );
  NAND U5860 ( .A(n4772), .B(n4773), .Z(x[150]) );
  NAND U5861 ( .A(creg[150]), .B(init), .Z(n4772) );
  NAND U5862 ( .A(n4774), .B(n4775), .Z(x[14]) );
  NAND U5863 ( .A(creg[14]), .B(init), .Z(n4774) );
  NAND U5864 ( .A(n4776), .B(n4777), .Z(x[149]) );
  NAND U5865 ( .A(creg[149]), .B(init), .Z(n4776) );
  NAND U5866 ( .A(n4778), .B(n4779), .Z(x[148]) );
  NAND U5867 ( .A(creg[148]), .B(init), .Z(n4778) );
  NAND U5868 ( .A(n4780), .B(n4781), .Z(x[147]) );
  NAND U5869 ( .A(creg[147]), .B(init), .Z(n4780) );
  NAND U5870 ( .A(n4782), .B(n4783), .Z(x[146]) );
  NAND U5871 ( .A(creg[146]), .B(init), .Z(n4782) );
  NAND U5872 ( .A(n4784), .B(n4785), .Z(x[145]) );
  NAND U5873 ( .A(creg[145]), .B(init), .Z(n4784) );
  NAND U5874 ( .A(n4786), .B(n4787), .Z(x[144]) );
  NAND U5875 ( .A(creg[144]), .B(init), .Z(n4786) );
  NAND U5876 ( .A(n4788), .B(n4789), .Z(x[143]) );
  NAND U5877 ( .A(creg[143]), .B(init), .Z(n4788) );
  NAND U5878 ( .A(n4790), .B(n4791), .Z(x[142]) );
  NAND U5879 ( .A(creg[142]), .B(init), .Z(n4790) );
  NAND U5880 ( .A(n4792), .B(n4793), .Z(x[141]) );
  NAND U5881 ( .A(creg[141]), .B(init), .Z(n4792) );
  NAND U5882 ( .A(n4794), .B(n4795), .Z(x[140]) );
  NAND U5883 ( .A(creg[140]), .B(init), .Z(n4794) );
  NAND U5884 ( .A(n4796), .B(n4797), .Z(x[13]) );
  NAND U5885 ( .A(creg[13]), .B(init), .Z(n4796) );
  NAND U5886 ( .A(n4798), .B(n4799), .Z(x[139]) );
  NAND U5887 ( .A(creg[139]), .B(init), .Z(n4798) );
  NAND U5888 ( .A(n4800), .B(n4801), .Z(x[138]) );
  NAND U5889 ( .A(creg[138]), .B(init), .Z(n4800) );
  NAND U5890 ( .A(n4802), .B(n4803), .Z(x[137]) );
  NAND U5891 ( .A(creg[137]), .B(init), .Z(n4802) );
  NAND U5892 ( .A(n4804), .B(n4805), .Z(x[136]) );
  NAND U5893 ( .A(creg[136]), .B(init), .Z(n4804) );
  NAND U5894 ( .A(n4806), .B(n4807), .Z(x[135]) );
  NAND U5895 ( .A(creg[135]), .B(init), .Z(n4806) );
  NAND U5896 ( .A(n4808), .B(n4809), .Z(x[134]) );
  NAND U5897 ( .A(creg[134]), .B(init), .Z(n4808) );
  NAND U5898 ( .A(n4810), .B(n4811), .Z(x[133]) );
  NAND U5899 ( .A(creg[133]), .B(init), .Z(n4810) );
  NAND U5900 ( .A(n4812), .B(n4813), .Z(x[132]) );
  NAND U5901 ( .A(creg[132]), .B(init), .Z(n4812) );
  NAND U5902 ( .A(n4814), .B(n4815), .Z(x[131]) );
  NAND U5903 ( .A(creg[131]), .B(init), .Z(n4814) );
  NAND U5904 ( .A(n4816), .B(n4817), .Z(x[130]) );
  NAND U5905 ( .A(creg[130]), .B(init), .Z(n4816) );
  NAND U5906 ( .A(n4818), .B(n4819), .Z(x[12]) );
  NAND U5907 ( .A(creg[12]), .B(init), .Z(n4818) );
  NAND U5908 ( .A(n4820), .B(n4821), .Z(x[129]) );
  NAND U5909 ( .A(creg[129]), .B(init), .Z(n4820) );
  NAND U5910 ( .A(n4822), .B(n4823), .Z(x[128]) );
  NAND U5911 ( .A(creg[128]), .B(init), .Z(n4822) );
  NAND U5912 ( .A(n4824), .B(n4825), .Z(x[127]) );
  NAND U5913 ( .A(creg[127]), .B(init), .Z(n4824) );
  NAND U5914 ( .A(n4826), .B(n4827), .Z(x[126]) );
  NAND U5915 ( .A(creg[126]), .B(init), .Z(n4826) );
  NAND U5916 ( .A(n4828), .B(n4829), .Z(x[125]) );
  NAND U5917 ( .A(creg[125]), .B(init), .Z(n4828) );
  NAND U5918 ( .A(n4830), .B(n4831), .Z(x[124]) );
  NAND U5919 ( .A(creg[124]), .B(init), .Z(n4830) );
  NAND U5920 ( .A(n4832), .B(n4833), .Z(x[123]) );
  NAND U5921 ( .A(creg[123]), .B(init), .Z(n4832) );
  NAND U5922 ( .A(n4834), .B(n4835), .Z(x[122]) );
  NAND U5923 ( .A(creg[122]), .B(init), .Z(n4834) );
  NAND U5924 ( .A(n4836), .B(n4837), .Z(x[121]) );
  NAND U5925 ( .A(creg[121]), .B(init), .Z(n4836) );
  NAND U5926 ( .A(n4838), .B(n4839), .Z(x[120]) );
  NAND U5927 ( .A(creg[120]), .B(init), .Z(n4838) );
  NAND U5928 ( .A(n4840), .B(n4841), .Z(x[11]) );
  NAND U5929 ( .A(creg[11]), .B(init), .Z(n4840) );
  NAND U5930 ( .A(n4842), .B(n4843), .Z(x[119]) );
  NAND U5931 ( .A(creg[119]), .B(init), .Z(n4842) );
  NAND U5932 ( .A(n4844), .B(n4845), .Z(x[118]) );
  NAND U5933 ( .A(creg[118]), .B(init), .Z(n4844) );
  NAND U5934 ( .A(n4846), .B(n4847), .Z(x[117]) );
  NAND U5935 ( .A(creg[117]), .B(init), .Z(n4846) );
  NAND U5936 ( .A(n4848), .B(n4849), .Z(x[116]) );
  NAND U5937 ( .A(creg[116]), .B(init), .Z(n4848) );
  NAND U5938 ( .A(n4850), .B(n4851), .Z(x[115]) );
  NAND U5939 ( .A(creg[115]), .B(init), .Z(n4850) );
  NAND U5940 ( .A(n4852), .B(n4853), .Z(x[114]) );
  NAND U5941 ( .A(creg[114]), .B(init), .Z(n4852) );
  NAND U5942 ( .A(n4854), .B(n4855), .Z(x[113]) );
  NAND U5943 ( .A(creg[113]), .B(init), .Z(n4854) );
  NAND U5944 ( .A(n4856), .B(n4857), .Z(x[112]) );
  NAND U5945 ( .A(creg[112]), .B(init), .Z(n4856) );
  NAND U5946 ( .A(n4858), .B(n4859), .Z(x[111]) );
  NAND U5947 ( .A(creg[111]), .B(init), .Z(n4858) );
  NAND U5948 ( .A(n4860), .B(n4861), .Z(x[110]) );
  NAND U5949 ( .A(creg[110]), .B(init), .Z(n4860) );
  NAND U5950 ( .A(n4862), .B(n4863), .Z(x[10]) );
  NAND U5951 ( .A(creg[10]), .B(init), .Z(n4862) );
  NAND U5952 ( .A(n4864), .B(n4865), .Z(x[109]) );
  NAND U5953 ( .A(creg[109]), .B(init), .Z(n4864) );
  NAND U5954 ( .A(n4866), .B(n4867), .Z(x[108]) );
  NAND U5955 ( .A(creg[108]), .B(init), .Z(n4866) );
  NAND U5956 ( .A(n4868), .B(n4869), .Z(x[107]) );
  NAND U5957 ( .A(creg[107]), .B(init), .Z(n4868) );
  NAND U5958 ( .A(n4870), .B(n4871), .Z(x[106]) );
  NAND U5959 ( .A(creg[106]), .B(init), .Z(n4870) );
  NAND U5960 ( .A(n4872), .B(n4873), .Z(x[105]) );
  NAND U5961 ( .A(creg[105]), .B(init), .Z(n4872) );
  NAND U5962 ( .A(n4874), .B(n4875), .Z(x[104]) );
  NAND U5963 ( .A(creg[104]), .B(init), .Z(n4874) );
  NAND U5964 ( .A(n4876), .B(n4877), .Z(x[103]) );
  NAND U5965 ( .A(creg[103]), .B(init), .Z(n4876) );
  NAND U5966 ( .A(n4878), .B(n4879), .Z(x[102]) );
  NAND U5967 ( .A(creg[102]), .B(init), .Z(n4878) );
  NAND U5968 ( .A(n4880), .B(n4881), .Z(x[101]) );
  NAND U5969 ( .A(creg[101]), .B(init), .Z(n4880) );
  NAND U5970 ( .A(n4882), .B(n4883), .Z(x[100]) );
  NAND U5971 ( .A(creg[100]), .B(init), .Z(n4882) );
  NAND U5972 ( .A(n4884), .B(n4885), .Z(x[0]) );
  NAND U5973 ( .A(creg[0]), .B(init), .Z(n4884) );
  AND U5974 ( .A(start_reg[9]), .B(init), .Z(start_in[9]) );
  AND U5975 ( .A(start_reg[8]), .B(init), .Z(start_in[8]) );
  AND U5976 ( .A(start_reg[7]), .B(init), .Z(start_in[7]) );
  AND U5977 ( .A(start_reg[6]), .B(init), .Z(start_in[6]) );
  AND U5978 ( .A(start_reg[62]), .B(init), .Z(start_in[62]) );
  AND U5979 ( .A(start_reg[61]), .B(init), .Z(start_in[61]) );
  AND U5980 ( .A(start_reg[60]), .B(init), .Z(start_in[60]) );
  AND U5981 ( .A(start_reg[5]), .B(init), .Z(start_in[5]) );
  AND U5982 ( .A(start_reg[59]), .B(init), .Z(start_in[59]) );
  AND U5983 ( .A(start_reg[58]), .B(init), .Z(start_in[58]) );
  AND U5984 ( .A(start_reg[57]), .B(init), .Z(start_in[57]) );
  AND U5985 ( .A(start_reg[56]), .B(init), .Z(start_in[56]) );
  AND U5986 ( .A(start_reg[55]), .B(init), .Z(start_in[55]) );
  AND U5987 ( .A(start_reg[54]), .B(init), .Z(start_in[54]) );
  AND U5988 ( .A(start_reg[53]), .B(init), .Z(start_in[53]) );
  AND U5989 ( .A(start_reg[52]), .B(init), .Z(start_in[52]) );
  AND U5990 ( .A(start_reg[51]), .B(init), .Z(start_in[51]) );
  AND U5991 ( .A(start_reg[50]), .B(init), .Z(start_in[50]) );
  AND U5992 ( .A(start_reg[4]), .B(init), .Z(start_in[4]) );
  AND U5993 ( .A(start_reg[49]), .B(init), .Z(start_in[49]) );
  AND U5994 ( .A(start_reg[48]), .B(init), .Z(start_in[48]) );
  AND U5995 ( .A(start_reg[47]), .B(init), .Z(start_in[47]) );
  AND U5996 ( .A(start_reg[46]), .B(init), .Z(start_in[46]) );
  AND U5997 ( .A(start_reg[45]), .B(init), .Z(start_in[45]) );
  AND U5998 ( .A(start_reg[44]), .B(init), .Z(start_in[44]) );
  AND U5999 ( .A(start_reg[43]), .B(init), .Z(start_in[43]) );
  AND U6000 ( .A(start_reg[42]), .B(init), .Z(start_in[42]) );
  AND U6001 ( .A(start_reg[41]), .B(init), .Z(start_in[41]) );
  AND U6002 ( .A(start_reg[40]), .B(init), .Z(start_in[40]) );
  AND U6003 ( .A(start_reg[3]), .B(init), .Z(start_in[3]) );
  AND U6004 ( .A(start_reg[39]), .B(init), .Z(start_in[39]) );
  AND U6005 ( .A(start_reg[38]), .B(init), .Z(start_in[38]) );
  AND U6006 ( .A(start_reg[37]), .B(init), .Z(start_in[37]) );
  AND U6007 ( .A(start_reg[36]), .B(init), .Z(start_in[36]) );
  AND U6008 ( .A(start_reg[35]), .B(init), .Z(start_in[35]) );
  AND U6009 ( .A(start_reg[34]), .B(init), .Z(start_in[34]) );
  AND U6010 ( .A(start_reg[33]), .B(init), .Z(start_in[33]) );
  AND U6011 ( .A(start_reg[32]), .B(init), .Z(start_in[32]) );
  AND U6012 ( .A(start_reg[31]), .B(init), .Z(start_in[31]) );
  AND U6013 ( .A(start_reg[30]), .B(init), .Z(start_in[30]) );
  AND U6014 ( .A(start_reg[2]), .B(init), .Z(start_in[2]) );
  AND U6015 ( .A(start_reg[29]), .B(init), .Z(start_in[29]) );
  AND U6016 ( .A(start_reg[28]), .B(init), .Z(start_in[28]) );
  AND U6017 ( .A(start_reg[27]), .B(init), .Z(start_in[27]) );
  AND U6018 ( .A(start_reg[26]), .B(init), .Z(start_in[26]) );
  AND U6019 ( .A(start_reg[25]), .B(init), .Z(start_in[25]) );
  AND U6020 ( .A(start_reg[24]), .B(init), .Z(start_in[24]) );
  AND U6021 ( .A(start_reg[23]), .B(init), .Z(start_in[23]) );
  AND U6022 ( .A(start_reg[22]), .B(init), .Z(start_in[22]) );
  AND U6023 ( .A(start_reg[21]), .B(init), .Z(start_in[21]) );
  AND U6024 ( .A(start_reg[20]), .B(init), .Z(start_in[20]) );
  AND U6025 ( .A(start_reg[1]), .B(init), .Z(start_in[1]) );
  AND U6026 ( .A(start_reg[19]), .B(init), .Z(start_in[19]) );
  AND U6027 ( .A(start_reg[18]), .B(init), .Z(start_in[18]) );
  AND U6028 ( .A(start_reg[17]), .B(init), .Z(start_in[17]) );
  AND U6029 ( .A(start_reg[16]), .B(init), .Z(start_in[16]) );
  AND U6030 ( .A(start_reg[15]), .B(init), .Z(start_in[15]) );
  AND U6031 ( .A(start_reg[14]), .B(init), .Z(start_in[14]) );
  AND U6032 ( .A(start_reg[13]), .B(init), .Z(start_in[13]) );
  AND U6033 ( .A(start_reg[12]), .B(init), .Z(start_in[12]) );
  AND U6034 ( .A(start_reg[11]), .B(init), .Z(start_in[11]) );
  AND U6035 ( .A(start_reg[10]), .B(init), .Z(start_in[10]) );
  NANDN U6036 ( .A(start_reg[0]), .B(init), .Z(start_in[0]) );
  NAND U6037 ( .A(n4886), .B(n4887), .Z(n3859) );
  NAND U6038 ( .A(n3863), .B(start_reg[63]), .Z(n4887) );
  IV U6039 ( .A(n3862), .Z(n3863) );
  NANDN U6040 ( .A(n7204), .B(mul_pow), .Z(n4886) );
  NAND U6041 ( .A(n4888), .B(n4889), .Z(n3858) );
  NANDN U6042 ( .A(n4890), .B(ereg[0]), .Z(n4889) );
  NANDN U6043 ( .A(init), .B(e[0]), .Z(n4888) );
  NAND U6044 ( .A(n4891), .B(n4892), .Z(n3857) );
  NANDN U6045 ( .A(init), .B(e[1]), .Z(n4892) );
  AND U6046 ( .A(n4893), .B(n4894), .Z(n4891) );
  NAND U6047 ( .A(n4895), .B(ereg[0]), .Z(n4894) );
  NANDN U6048 ( .A(n4890), .B(ereg[1]), .Z(n4893) );
  NAND U6049 ( .A(n4896), .B(n4897), .Z(n3856) );
  NANDN U6050 ( .A(init), .B(e[2]), .Z(n4897) );
  AND U6051 ( .A(n4898), .B(n4899), .Z(n4896) );
  NAND U6052 ( .A(ereg[1]), .B(n4895), .Z(n4899) );
  NANDN U6053 ( .A(n4890), .B(ereg[2]), .Z(n4898) );
  NAND U6054 ( .A(n4900), .B(n4901), .Z(n3855) );
  NANDN U6055 ( .A(init), .B(e[3]), .Z(n4901) );
  AND U6056 ( .A(n4902), .B(n4903), .Z(n4900) );
  NAND U6057 ( .A(ereg[2]), .B(n4895), .Z(n4903) );
  NANDN U6058 ( .A(n4890), .B(ereg[3]), .Z(n4902) );
  NAND U6059 ( .A(n4904), .B(n4905), .Z(n3854) );
  NANDN U6060 ( .A(init), .B(e[4]), .Z(n4905) );
  AND U6061 ( .A(n4906), .B(n4907), .Z(n4904) );
  NAND U6062 ( .A(ereg[3]), .B(n4895), .Z(n4907) );
  NANDN U6063 ( .A(n4890), .B(ereg[4]), .Z(n4906) );
  NAND U6064 ( .A(n4908), .B(n4909), .Z(n3853) );
  NANDN U6065 ( .A(init), .B(e[5]), .Z(n4909) );
  AND U6066 ( .A(n4910), .B(n4911), .Z(n4908) );
  NAND U6067 ( .A(ereg[4]), .B(n4895), .Z(n4911) );
  NANDN U6068 ( .A(n4890), .B(ereg[5]), .Z(n4910) );
  NAND U6069 ( .A(n4912), .B(n4913), .Z(n3852) );
  NANDN U6070 ( .A(init), .B(e[6]), .Z(n4913) );
  AND U6071 ( .A(n4914), .B(n4915), .Z(n4912) );
  NAND U6072 ( .A(ereg[5]), .B(n4895), .Z(n4915) );
  NANDN U6073 ( .A(n4890), .B(ereg[6]), .Z(n4914) );
  NAND U6074 ( .A(n4916), .B(n4917), .Z(n3851) );
  NANDN U6075 ( .A(init), .B(e[7]), .Z(n4917) );
  AND U6076 ( .A(n4918), .B(n4919), .Z(n4916) );
  NAND U6077 ( .A(ereg[6]), .B(n4895), .Z(n4919) );
  NANDN U6078 ( .A(n4890), .B(ereg[7]), .Z(n4918) );
  NAND U6079 ( .A(n4920), .B(n4921), .Z(n3850) );
  NANDN U6080 ( .A(init), .B(e[8]), .Z(n4921) );
  AND U6081 ( .A(n4922), .B(n4923), .Z(n4920) );
  NAND U6082 ( .A(ereg[7]), .B(n4895), .Z(n4923) );
  NANDN U6083 ( .A(n4890), .B(ereg[8]), .Z(n4922) );
  NAND U6084 ( .A(n4924), .B(n4925), .Z(n3849) );
  NANDN U6085 ( .A(init), .B(e[9]), .Z(n4925) );
  AND U6086 ( .A(n4926), .B(n4927), .Z(n4924) );
  NAND U6087 ( .A(ereg[8]), .B(n4895), .Z(n4927) );
  NANDN U6088 ( .A(n4890), .B(ereg[9]), .Z(n4926) );
  NAND U6089 ( .A(n4928), .B(n4929), .Z(n3848) );
  NANDN U6090 ( .A(init), .B(e[10]), .Z(n4929) );
  AND U6091 ( .A(n4930), .B(n4931), .Z(n4928) );
  NAND U6092 ( .A(ereg[9]), .B(n4895), .Z(n4931) );
  NANDN U6093 ( .A(n4890), .B(ereg[10]), .Z(n4930) );
  NAND U6094 ( .A(n4932), .B(n4933), .Z(n3847) );
  NANDN U6095 ( .A(init), .B(e[11]), .Z(n4933) );
  AND U6096 ( .A(n4934), .B(n4935), .Z(n4932) );
  NAND U6097 ( .A(ereg[10]), .B(n4895), .Z(n4935) );
  NANDN U6098 ( .A(n4890), .B(ereg[11]), .Z(n4934) );
  NAND U6099 ( .A(n4936), .B(n4937), .Z(n3846) );
  NANDN U6100 ( .A(init), .B(e[12]), .Z(n4937) );
  AND U6101 ( .A(n4938), .B(n4939), .Z(n4936) );
  NAND U6102 ( .A(ereg[11]), .B(n4895), .Z(n4939) );
  NANDN U6103 ( .A(n4890), .B(ereg[12]), .Z(n4938) );
  NAND U6104 ( .A(n4940), .B(n4941), .Z(n3845) );
  NANDN U6105 ( .A(init), .B(e[13]), .Z(n4941) );
  AND U6106 ( .A(n4942), .B(n4943), .Z(n4940) );
  NAND U6107 ( .A(ereg[12]), .B(n4895), .Z(n4943) );
  NANDN U6108 ( .A(n4890), .B(ereg[13]), .Z(n4942) );
  NAND U6109 ( .A(n4944), .B(n4945), .Z(n3844) );
  NANDN U6110 ( .A(init), .B(e[14]), .Z(n4945) );
  AND U6111 ( .A(n4946), .B(n4947), .Z(n4944) );
  NAND U6112 ( .A(ereg[13]), .B(n4895), .Z(n4947) );
  NANDN U6113 ( .A(n4890), .B(ereg[14]), .Z(n4946) );
  NAND U6114 ( .A(n4948), .B(n4949), .Z(n3843) );
  NANDN U6115 ( .A(init), .B(e[15]), .Z(n4949) );
  AND U6116 ( .A(n4950), .B(n4951), .Z(n4948) );
  NAND U6117 ( .A(ereg[14]), .B(n4895), .Z(n4951) );
  NANDN U6118 ( .A(n4890), .B(ereg[15]), .Z(n4950) );
  NAND U6119 ( .A(n4952), .B(n4953), .Z(n3842) );
  NANDN U6120 ( .A(init), .B(e[16]), .Z(n4953) );
  AND U6121 ( .A(n4954), .B(n4955), .Z(n4952) );
  NAND U6122 ( .A(ereg[15]), .B(n4895), .Z(n4955) );
  NANDN U6123 ( .A(n4890), .B(ereg[16]), .Z(n4954) );
  NAND U6124 ( .A(n4956), .B(n4957), .Z(n3841) );
  NANDN U6125 ( .A(init), .B(e[17]), .Z(n4957) );
  AND U6126 ( .A(n4958), .B(n4959), .Z(n4956) );
  NAND U6127 ( .A(ereg[16]), .B(n4895), .Z(n4959) );
  NANDN U6128 ( .A(n4890), .B(ereg[17]), .Z(n4958) );
  NAND U6129 ( .A(n4960), .B(n4961), .Z(n3840) );
  NANDN U6130 ( .A(init), .B(e[18]), .Z(n4961) );
  AND U6131 ( .A(n4962), .B(n4963), .Z(n4960) );
  NAND U6132 ( .A(ereg[17]), .B(n4895), .Z(n4963) );
  NANDN U6133 ( .A(n4890), .B(ereg[18]), .Z(n4962) );
  NAND U6134 ( .A(n4964), .B(n4965), .Z(n3839) );
  NANDN U6135 ( .A(init), .B(e[19]), .Z(n4965) );
  AND U6136 ( .A(n4966), .B(n4967), .Z(n4964) );
  NAND U6137 ( .A(ereg[18]), .B(n4895), .Z(n4967) );
  NANDN U6138 ( .A(n4890), .B(ereg[19]), .Z(n4966) );
  NAND U6139 ( .A(n4968), .B(n4969), .Z(n3838) );
  NANDN U6140 ( .A(init), .B(e[20]), .Z(n4969) );
  AND U6141 ( .A(n4970), .B(n4971), .Z(n4968) );
  NAND U6142 ( .A(ereg[19]), .B(n4895), .Z(n4971) );
  NANDN U6143 ( .A(n4890), .B(ereg[20]), .Z(n4970) );
  NAND U6144 ( .A(n4972), .B(n4973), .Z(n3837) );
  NANDN U6145 ( .A(init), .B(e[21]), .Z(n4973) );
  AND U6146 ( .A(n4974), .B(n4975), .Z(n4972) );
  NAND U6147 ( .A(ereg[20]), .B(n4895), .Z(n4975) );
  NANDN U6148 ( .A(n4890), .B(ereg[21]), .Z(n4974) );
  NAND U6149 ( .A(n4976), .B(n4977), .Z(n3836) );
  NANDN U6150 ( .A(init), .B(e[22]), .Z(n4977) );
  AND U6151 ( .A(n4978), .B(n4979), .Z(n4976) );
  NAND U6152 ( .A(ereg[21]), .B(n4895), .Z(n4979) );
  NANDN U6153 ( .A(n4890), .B(ereg[22]), .Z(n4978) );
  NAND U6154 ( .A(n4980), .B(n4981), .Z(n3835) );
  NANDN U6155 ( .A(init), .B(e[23]), .Z(n4981) );
  AND U6156 ( .A(n4982), .B(n4983), .Z(n4980) );
  NAND U6157 ( .A(ereg[22]), .B(n4895), .Z(n4983) );
  NANDN U6158 ( .A(n4890), .B(ereg[23]), .Z(n4982) );
  NAND U6159 ( .A(n4984), .B(n4985), .Z(n3834) );
  NANDN U6160 ( .A(init), .B(e[24]), .Z(n4985) );
  AND U6161 ( .A(n4986), .B(n4987), .Z(n4984) );
  NAND U6162 ( .A(ereg[23]), .B(n4895), .Z(n4987) );
  NANDN U6163 ( .A(n4890), .B(ereg[24]), .Z(n4986) );
  NAND U6164 ( .A(n4988), .B(n4989), .Z(n3833) );
  NANDN U6165 ( .A(init), .B(e[25]), .Z(n4989) );
  AND U6166 ( .A(n4990), .B(n4991), .Z(n4988) );
  NAND U6167 ( .A(ereg[24]), .B(n4895), .Z(n4991) );
  NANDN U6168 ( .A(n4890), .B(ereg[25]), .Z(n4990) );
  NAND U6169 ( .A(n4992), .B(n4993), .Z(n3832) );
  NANDN U6170 ( .A(init), .B(e[26]), .Z(n4993) );
  AND U6171 ( .A(n4994), .B(n4995), .Z(n4992) );
  NAND U6172 ( .A(ereg[25]), .B(n4895), .Z(n4995) );
  NANDN U6173 ( .A(n4890), .B(ereg[26]), .Z(n4994) );
  NAND U6174 ( .A(n4996), .B(n4997), .Z(n3831) );
  NANDN U6175 ( .A(init), .B(e[27]), .Z(n4997) );
  AND U6176 ( .A(n4998), .B(n4999), .Z(n4996) );
  NAND U6177 ( .A(ereg[26]), .B(n4895), .Z(n4999) );
  NANDN U6178 ( .A(n4890), .B(ereg[27]), .Z(n4998) );
  NAND U6179 ( .A(n5000), .B(n5001), .Z(n3830) );
  NANDN U6180 ( .A(init), .B(e[28]), .Z(n5001) );
  AND U6181 ( .A(n5002), .B(n5003), .Z(n5000) );
  NAND U6182 ( .A(ereg[27]), .B(n4895), .Z(n5003) );
  NANDN U6183 ( .A(n4890), .B(ereg[28]), .Z(n5002) );
  NAND U6184 ( .A(n5004), .B(n5005), .Z(n3829) );
  NANDN U6185 ( .A(init), .B(e[29]), .Z(n5005) );
  AND U6186 ( .A(n5006), .B(n5007), .Z(n5004) );
  NAND U6187 ( .A(ereg[28]), .B(n4895), .Z(n5007) );
  NANDN U6188 ( .A(n4890), .B(ereg[29]), .Z(n5006) );
  NAND U6189 ( .A(n5008), .B(n5009), .Z(n3828) );
  NANDN U6190 ( .A(init), .B(e[30]), .Z(n5009) );
  AND U6191 ( .A(n5010), .B(n5011), .Z(n5008) );
  NAND U6192 ( .A(ereg[29]), .B(n4895), .Z(n5011) );
  NANDN U6193 ( .A(n4890), .B(ereg[30]), .Z(n5010) );
  NAND U6194 ( .A(n5012), .B(n5013), .Z(n3827) );
  NANDN U6195 ( .A(init), .B(e[31]), .Z(n5013) );
  AND U6196 ( .A(n5014), .B(n5015), .Z(n5012) );
  NAND U6197 ( .A(ereg[30]), .B(n4895), .Z(n5015) );
  NANDN U6198 ( .A(n4890), .B(ereg[31]), .Z(n5014) );
  NAND U6199 ( .A(n5016), .B(n5017), .Z(n3826) );
  NANDN U6200 ( .A(init), .B(e[32]), .Z(n5017) );
  AND U6201 ( .A(n5018), .B(n5019), .Z(n5016) );
  NAND U6202 ( .A(ereg[31]), .B(n4895), .Z(n5019) );
  NANDN U6203 ( .A(n4890), .B(ereg[32]), .Z(n5018) );
  NAND U6204 ( .A(n5020), .B(n5021), .Z(n3825) );
  NANDN U6205 ( .A(init), .B(e[33]), .Z(n5021) );
  AND U6206 ( .A(n5022), .B(n5023), .Z(n5020) );
  NAND U6207 ( .A(ereg[32]), .B(n4895), .Z(n5023) );
  NANDN U6208 ( .A(n4890), .B(ereg[33]), .Z(n5022) );
  NAND U6209 ( .A(n5024), .B(n5025), .Z(n3824) );
  NANDN U6210 ( .A(init), .B(e[34]), .Z(n5025) );
  AND U6211 ( .A(n5026), .B(n5027), .Z(n5024) );
  NAND U6212 ( .A(ereg[33]), .B(n4895), .Z(n5027) );
  NANDN U6213 ( .A(n4890), .B(ereg[34]), .Z(n5026) );
  NAND U6214 ( .A(n5028), .B(n5029), .Z(n3823) );
  NANDN U6215 ( .A(init), .B(e[35]), .Z(n5029) );
  AND U6216 ( .A(n5030), .B(n5031), .Z(n5028) );
  NAND U6217 ( .A(ereg[34]), .B(n4895), .Z(n5031) );
  NANDN U6218 ( .A(n4890), .B(ereg[35]), .Z(n5030) );
  NAND U6219 ( .A(n5032), .B(n5033), .Z(n3822) );
  NANDN U6220 ( .A(init), .B(e[36]), .Z(n5033) );
  AND U6221 ( .A(n5034), .B(n5035), .Z(n5032) );
  NAND U6222 ( .A(ereg[35]), .B(n4895), .Z(n5035) );
  NANDN U6223 ( .A(n4890), .B(ereg[36]), .Z(n5034) );
  NAND U6224 ( .A(n5036), .B(n5037), .Z(n3821) );
  NANDN U6225 ( .A(init), .B(e[37]), .Z(n5037) );
  AND U6226 ( .A(n5038), .B(n5039), .Z(n5036) );
  NAND U6227 ( .A(ereg[36]), .B(n4895), .Z(n5039) );
  NANDN U6228 ( .A(n4890), .B(ereg[37]), .Z(n5038) );
  NAND U6229 ( .A(n5040), .B(n5041), .Z(n3820) );
  NANDN U6230 ( .A(init), .B(e[38]), .Z(n5041) );
  AND U6231 ( .A(n5042), .B(n5043), .Z(n5040) );
  NAND U6232 ( .A(ereg[37]), .B(n4895), .Z(n5043) );
  NANDN U6233 ( .A(n4890), .B(ereg[38]), .Z(n5042) );
  NAND U6234 ( .A(n5044), .B(n5045), .Z(n3819) );
  NANDN U6235 ( .A(init), .B(e[39]), .Z(n5045) );
  AND U6236 ( .A(n5046), .B(n5047), .Z(n5044) );
  NAND U6237 ( .A(ereg[38]), .B(n4895), .Z(n5047) );
  NANDN U6238 ( .A(n4890), .B(ereg[39]), .Z(n5046) );
  NAND U6239 ( .A(n5048), .B(n5049), .Z(n3818) );
  NANDN U6240 ( .A(init), .B(e[40]), .Z(n5049) );
  AND U6241 ( .A(n5050), .B(n5051), .Z(n5048) );
  NAND U6242 ( .A(ereg[39]), .B(n4895), .Z(n5051) );
  NANDN U6243 ( .A(n4890), .B(ereg[40]), .Z(n5050) );
  NAND U6244 ( .A(n5052), .B(n5053), .Z(n3817) );
  NANDN U6245 ( .A(init), .B(e[41]), .Z(n5053) );
  AND U6246 ( .A(n5054), .B(n5055), .Z(n5052) );
  NAND U6247 ( .A(ereg[40]), .B(n4895), .Z(n5055) );
  NANDN U6248 ( .A(n4890), .B(ereg[41]), .Z(n5054) );
  NAND U6249 ( .A(n5056), .B(n5057), .Z(n3816) );
  NANDN U6250 ( .A(init), .B(e[42]), .Z(n5057) );
  AND U6251 ( .A(n5058), .B(n5059), .Z(n5056) );
  NAND U6252 ( .A(ereg[41]), .B(n4895), .Z(n5059) );
  NANDN U6253 ( .A(n4890), .B(ereg[42]), .Z(n5058) );
  NAND U6254 ( .A(n5060), .B(n5061), .Z(n3815) );
  NANDN U6255 ( .A(init), .B(e[43]), .Z(n5061) );
  AND U6256 ( .A(n5062), .B(n5063), .Z(n5060) );
  NAND U6257 ( .A(ereg[42]), .B(n4895), .Z(n5063) );
  NANDN U6258 ( .A(n4890), .B(ereg[43]), .Z(n5062) );
  NAND U6259 ( .A(n5064), .B(n5065), .Z(n3814) );
  NANDN U6260 ( .A(init), .B(e[44]), .Z(n5065) );
  AND U6261 ( .A(n5066), .B(n5067), .Z(n5064) );
  NAND U6262 ( .A(ereg[43]), .B(n4895), .Z(n5067) );
  NANDN U6263 ( .A(n4890), .B(ereg[44]), .Z(n5066) );
  NAND U6264 ( .A(n5068), .B(n5069), .Z(n3813) );
  NANDN U6265 ( .A(init), .B(e[45]), .Z(n5069) );
  AND U6266 ( .A(n5070), .B(n5071), .Z(n5068) );
  NAND U6267 ( .A(ereg[44]), .B(n4895), .Z(n5071) );
  NANDN U6268 ( .A(n4890), .B(ereg[45]), .Z(n5070) );
  NAND U6269 ( .A(n5072), .B(n5073), .Z(n3812) );
  NANDN U6270 ( .A(init), .B(e[46]), .Z(n5073) );
  AND U6271 ( .A(n5074), .B(n5075), .Z(n5072) );
  NAND U6272 ( .A(ereg[45]), .B(n4895), .Z(n5075) );
  NANDN U6273 ( .A(n4890), .B(ereg[46]), .Z(n5074) );
  NAND U6274 ( .A(n5076), .B(n5077), .Z(n3811) );
  NANDN U6275 ( .A(init), .B(e[47]), .Z(n5077) );
  AND U6276 ( .A(n5078), .B(n5079), .Z(n5076) );
  NAND U6277 ( .A(ereg[46]), .B(n4895), .Z(n5079) );
  NANDN U6278 ( .A(n4890), .B(ereg[47]), .Z(n5078) );
  NAND U6279 ( .A(n5080), .B(n5081), .Z(n3810) );
  NANDN U6280 ( .A(init), .B(e[48]), .Z(n5081) );
  AND U6281 ( .A(n5082), .B(n5083), .Z(n5080) );
  NAND U6282 ( .A(ereg[47]), .B(n4895), .Z(n5083) );
  NANDN U6283 ( .A(n4890), .B(ereg[48]), .Z(n5082) );
  NAND U6284 ( .A(n5084), .B(n5085), .Z(n3809) );
  NANDN U6285 ( .A(init), .B(e[49]), .Z(n5085) );
  AND U6286 ( .A(n5086), .B(n5087), .Z(n5084) );
  NAND U6287 ( .A(ereg[48]), .B(n4895), .Z(n5087) );
  NANDN U6288 ( .A(n4890), .B(ereg[49]), .Z(n5086) );
  NAND U6289 ( .A(n5088), .B(n5089), .Z(n3808) );
  NANDN U6290 ( .A(init), .B(e[50]), .Z(n5089) );
  AND U6291 ( .A(n5090), .B(n5091), .Z(n5088) );
  NAND U6292 ( .A(ereg[49]), .B(n4895), .Z(n5091) );
  NANDN U6293 ( .A(n4890), .B(ereg[50]), .Z(n5090) );
  NAND U6294 ( .A(n5092), .B(n5093), .Z(n3807) );
  NANDN U6295 ( .A(init), .B(e[51]), .Z(n5093) );
  AND U6296 ( .A(n5094), .B(n5095), .Z(n5092) );
  NAND U6297 ( .A(ereg[50]), .B(n4895), .Z(n5095) );
  NANDN U6298 ( .A(n4890), .B(ereg[51]), .Z(n5094) );
  NAND U6299 ( .A(n5096), .B(n5097), .Z(n3806) );
  NANDN U6300 ( .A(init), .B(e[52]), .Z(n5097) );
  AND U6301 ( .A(n5098), .B(n5099), .Z(n5096) );
  NAND U6302 ( .A(ereg[51]), .B(n4895), .Z(n5099) );
  NANDN U6303 ( .A(n4890), .B(ereg[52]), .Z(n5098) );
  NAND U6304 ( .A(n5100), .B(n5101), .Z(n3805) );
  NANDN U6305 ( .A(init), .B(e[53]), .Z(n5101) );
  AND U6306 ( .A(n5102), .B(n5103), .Z(n5100) );
  NAND U6307 ( .A(ereg[52]), .B(n4895), .Z(n5103) );
  NANDN U6308 ( .A(n4890), .B(ereg[53]), .Z(n5102) );
  NAND U6309 ( .A(n5104), .B(n5105), .Z(n3804) );
  NANDN U6310 ( .A(init), .B(e[54]), .Z(n5105) );
  AND U6311 ( .A(n5106), .B(n5107), .Z(n5104) );
  NAND U6312 ( .A(ereg[53]), .B(n4895), .Z(n5107) );
  NANDN U6313 ( .A(n4890), .B(ereg[54]), .Z(n5106) );
  NAND U6314 ( .A(n5108), .B(n5109), .Z(n3803) );
  NANDN U6315 ( .A(init), .B(e[55]), .Z(n5109) );
  AND U6316 ( .A(n5110), .B(n5111), .Z(n5108) );
  NAND U6317 ( .A(ereg[54]), .B(n4895), .Z(n5111) );
  NANDN U6318 ( .A(n4890), .B(ereg[55]), .Z(n5110) );
  NAND U6319 ( .A(n5112), .B(n5113), .Z(n3802) );
  NANDN U6320 ( .A(init), .B(e[56]), .Z(n5113) );
  AND U6321 ( .A(n5114), .B(n5115), .Z(n5112) );
  NAND U6322 ( .A(ereg[55]), .B(n4895), .Z(n5115) );
  NANDN U6323 ( .A(n4890), .B(ereg[56]), .Z(n5114) );
  NAND U6324 ( .A(n5116), .B(n5117), .Z(n3801) );
  NANDN U6325 ( .A(init), .B(e[57]), .Z(n5117) );
  AND U6326 ( .A(n5118), .B(n5119), .Z(n5116) );
  NAND U6327 ( .A(ereg[56]), .B(n4895), .Z(n5119) );
  NANDN U6328 ( .A(n4890), .B(ereg[57]), .Z(n5118) );
  NAND U6329 ( .A(n5120), .B(n5121), .Z(n3800) );
  NANDN U6330 ( .A(init), .B(e[58]), .Z(n5121) );
  AND U6331 ( .A(n5122), .B(n5123), .Z(n5120) );
  NAND U6332 ( .A(ereg[57]), .B(n4895), .Z(n5123) );
  NANDN U6333 ( .A(n4890), .B(ereg[58]), .Z(n5122) );
  NAND U6334 ( .A(n5124), .B(n5125), .Z(n3799) );
  NANDN U6335 ( .A(init), .B(e[59]), .Z(n5125) );
  AND U6336 ( .A(n5126), .B(n5127), .Z(n5124) );
  NAND U6337 ( .A(ereg[58]), .B(n4895), .Z(n5127) );
  NANDN U6338 ( .A(n4890), .B(ereg[59]), .Z(n5126) );
  NAND U6339 ( .A(n5128), .B(n5129), .Z(n3798) );
  NANDN U6340 ( .A(init), .B(e[60]), .Z(n5129) );
  AND U6341 ( .A(n5130), .B(n5131), .Z(n5128) );
  NAND U6342 ( .A(ereg[59]), .B(n4895), .Z(n5131) );
  NANDN U6343 ( .A(n4890), .B(ereg[60]), .Z(n5130) );
  NAND U6344 ( .A(n5132), .B(n5133), .Z(n3797) );
  NANDN U6345 ( .A(init), .B(e[61]), .Z(n5133) );
  AND U6346 ( .A(n5134), .B(n5135), .Z(n5132) );
  NAND U6347 ( .A(ereg[60]), .B(n4895), .Z(n5135) );
  NANDN U6348 ( .A(n4890), .B(ereg[61]), .Z(n5134) );
  NAND U6349 ( .A(n5136), .B(n5137), .Z(n3796) );
  NANDN U6350 ( .A(init), .B(e[62]), .Z(n5137) );
  AND U6351 ( .A(n5138), .B(n5139), .Z(n5136) );
  NAND U6352 ( .A(ereg[61]), .B(n4895), .Z(n5139) );
  NANDN U6353 ( .A(n4890), .B(ereg[62]), .Z(n5138) );
  NAND U6354 ( .A(n5140), .B(n5141), .Z(n3795) );
  NANDN U6355 ( .A(init), .B(e[63]), .Z(n5141) );
  AND U6356 ( .A(n5142), .B(n5143), .Z(n5140) );
  NAND U6357 ( .A(ereg[62]), .B(n4895), .Z(n5143) );
  NANDN U6358 ( .A(n4890), .B(ereg[63]), .Z(n5142) );
  NAND U6359 ( .A(n5144), .B(n5145), .Z(n3794) );
  NANDN U6360 ( .A(init), .B(e[64]), .Z(n5145) );
  AND U6361 ( .A(n5146), .B(n5147), .Z(n5144) );
  NAND U6362 ( .A(ereg[63]), .B(n4895), .Z(n5147) );
  NANDN U6363 ( .A(n4890), .B(ereg[64]), .Z(n5146) );
  NAND U6364 ( .A(n5148), .B(n5149), .Z(n3793) );
  NANDN U6365 ( .A(init), .B(e[65]), .Z(n5149) );
  AND U6366 ( .A(n5150), .B(n5151), .Z(n5148) );
  NAND U6367 ( .A(ereg[64]), .B(n4895), .Z(n5151) );
  NANDN U6368 ( .A(n4890), .B(ereg[65]), .Z(n5150) );
  NAND U6369 ( .A(n5152), .B(n5153), .Z(n3792) );
  NANDN U6370 ( .A(init), .B(e[66]), .Z(n5153) );
  AND U6371 ( .A(n5154), .B(n5155), .Z(n5152) );
  NAND U6372 ( .A(ereg[65]), .B(n4895), .Z(n5155) );
  NANDN U6373 ( .A(n4890), .B(ereg[66]), .Z(n5154) );
  NAND U6374 ( .A(n5156), .B(n5157), .Z(n3791) );
  NANDN U6375 ( .A(init), .B(e[67]), .Z(n5157) );
  AND U6376 ( .A(n5158), .B(n5159), .Z(n5156) );
  NAND U6377 ( .A(ereg[66]), .B(n4895), .Z(n5159) );
  NANDN U6378 ( .A(n4890), .B(ereg[67]), .Z(n5158) );
  NAND U6379 ( .A(n5160), .B(n5161), .Z(n3790) );
  NANDN U6380 ( .A(init), .B(e[68]), .Z(n5161) );
  AND U6381 ( .A(n5162), .B(n5163), .Z(n5160) );
  NAND U6382 ( .A(ereg[67]), .B(n4895), .Z(n5163) );
  NANDN U6383 ( .A(n4890), .B(ereg[68]), .Z(n5162) );
  NAND U6384 ( .A(n5164), .B(n5165), .Z(n3789) );
  NANDN U6385 ( .A(init), .B(e[69]), .Z(n5165) );
  AND U6386 ( .A(n5166), .B(n5167), .Z(n5164) );
  NAND U6387 ( .A(ereg[68]), .B(n4895), .Z(n5167) );
  NANDN U6388 ( .A(n4890), .B(ereg[69]), .Z(n5166) );
  NAND U6389 ( .A(n5168), .B(n5169), .Z(n3788) );
  NANDN U6390 ( .A(init), .B(e[70]), .Z(n5169) );
  AND U6391 ( .A(n5170), .B(n5171), .Z(n5168) );
  NAND U6392 ( .A(ereg[69]), .B(n4895), .Z(n5171) );
  NANDN U6393 ( .A(n4890), .B(ereg[70]), .Z(n5170) );
  NAND U6394 ( .A(n5172), .B(n5173), .Z(n3787) );
  NANDN U6395 ( .A(init), .B(e[71]), .Z(n5173) );
  AND U6396 ( .A(n5174), .B(n5175), .Z(n5172) );
  NAND U6397 ( .A(ereg[70]), .B(n4895), .Z(n5175) );
  NANDN U6398 ( .A(n4890), .B(ereg[71]), .Z(n5174) );
  NAND U6399 ( .A(n5176), .B(n5177), .Z(n3786) );
  NANDN U6400 ( .A(init), .B(e[72]), .Z(n5177) );
  AND U6401 ( .A(n5178), .B(n5179), .Z(n5176) );
  NAND U6402 ( .A(ereg[71]), .B(n4895), .Z(n5179) );
  NANDN U6403 ( .A(n4890), .B(ereg[72]), .Z(n5178) );
  NAND U6404 ( .A(n5180), .B(n5181), .Z(n3785) );
  NANDN U6405 ( .A(init), .B(e[73]), .Z(n5181) );
  AND U6406 ( .A(n5182), .B(n5183), .Z(n5180) );
  NAND U6407 ( .A(ereg[72]), .B(n4895), .Z(n5183) );
  NANDN U6408 ( .A(n4890), .B(ereg[73]), .Z(n5182) );
  NAND U6409 ( .A(n5184), .B(n5185), .Z(n3784) );
  NANDN U6410 ( .A(init), .B(e[74]), .Z(n5185) );
  AND U6411 ( .A(n5186), .B(n5187), .Z(n5184) );
  NAND U6412 ( .A(ereg[73]), .B(n4895), .Z(n5187) );
  NANDN U6413 ( .A(n4890), .B(ereg[74]), .Z(n5186) );
  NAND U6414 ( .A(n5188), .B(n5189), .Z(n3783) );
  NANDN U6415 ( .A(init), .B(e[75]), .Z(n5189) );
  AND U6416 ( .A(n5190), .B(n5191), .Z(n5188) );
  NAND U6417 ( .A(ereg[74]), .B(n4895), .Z(n5191) );
  NANDN U6418 ( .A(n4890), .B(ereg[75]), .Z(n5190) );
  NAND U6419 ( .A(n5192), .B(n5193), .Z(n3782) );
  NANDN U6420 ( .A(init), .B(e[76]), .Z(n5193) );
  AND U6421 ( .A(n5194), .B(n5195), .Z(n5192) );
  NAND U6422 ( .A(ereg[75]), .B(n4895), .Z(n5195) );
  NANDN U6423 ( .A(n4890), .B(ereg[76]), .Z(n5194) );
  NAND U6424 ( .A(n5196), .B(n5197), .Z(n3781) );
  NANDN U6425 ( .A(init), .B(e[77]), .Z(n5197) );
  AND U6426 ( .A(n5198), .B(n5199), .Z(n5196) );
  NAND U6427 ( .A(ereg[76]), .B(n4895), .Z(n5199) );
  NANDN U6428 ( .A(n4890), .B(ereg[77]), .Z(n5198) );
  NAND U6429 ( .A(n5200), .B(n5201), .Z(n3780) );
  NANDN U6430 ( .A(init), .B(e[78]), .Z(n5201) );
  AND U6431 ( .A(n5202), .B(n5203), .Z(n5200) );
  NAND U6432 ( .A(ereg[77]), .B(n4895), .Z(n5203) );
  NANDN U6433 ( .A(n4890), .B(ereg[78]), .Z(n5202) );
  NAND U6434 ( .A(n5204), .B(n5205), .Z(n3779) );
  NANDN U6435 ( .A(init), .B(e[79]), .Z(n5205) );
  AND U6436 ( .A(n5206), .B(n5207), .Z(n5204) );
  NAND U6437 ( .A(ereg[78]), .B(n4895), .Z(n5207) );
  NANDN U6438 ( .A(n4890), .B(ereg[79]), .Z(n5206) );
  NAND U6439 ( .A(n5208), .B(n5209), .Z(n3778) );
  NANDN U6440 ( .A(init), .B(e[80]), .Z(n5209) );
  AND U6441 ( .A(n5210), .B(n5211), .Z(n5208) );
  NAND U6442 ( .A(ereg[79]), .B(n4895), .Z(n5211) );
  NANDN U6443 ( .A(n4890), .B(ereg[80]), .Z(n5210) );
  NAND U6444 ( .A(n5212), .B(n5213), .Z(n3777) );
  NANDN U6445 ( .A(init), .B(e[81]), .Z(n5213) );
  AND U6446 ( .A(n5214), .B(n5215), .Z(n5212) );
  NAND U6447 ( .A(ereg[80]), .B(n4895), .Z(n5215) );
  NANDN U6448 ( .A(n4890), .B(ereg[81]), .Z(n5214) );
  NAND U6449 ( .A(n5216), .B(n5217), .Z(n3776) );
  NANDN U6450 ( .A(init), .B(e[82]), .Z(n5217) );
  AND U6451 ( .A(n5218), .B(n5219), .Z(n5216) );
  NAND U6452 ( .A(ereg[81]), .B(n4895), .Z(n5219) );
  NANDN U6453 ( .A(n4890), .B(ereg[82]), .Z(n5218) );
  NAND U6454 ( .A(n5220), .B(n5221), .Z(n3775) );
  NANDN U6455 ( .A(init), .B(e[83]), .Z(n5221) );
  AND U6456 ( .A(n5222), .B(n5223), .Z(n5220) );
  NAND U6457 ( .A(ereg[82]), .B(n4895), .Z(n5223) );
  NANDN U6458 ( .A(n4890), .B(ereg[83]), .Z(n5222) );
  NAND U6459 ( .A(n5224), .B(n5225), .Z(n3774) );
  NANDN U6460 ( .A(init), .B(e[84]), .Z(n5225) );
  AND U6461 ( .A(n5226), .B(n5227), .Z(n5224) );
  NAND U6462 ( .A(ereg[83]), .B(n4895), .Z(n5227) );
  NANDN U6463 ( .A(n4890), .B(ereg[84]), .Z(n5226) );
  NAND U6464 ( .A(n5228), .B(n5229), .Z(n3773) );
  NANDN U6465 ( .A(init), .B(e[85]), .Z(n5229) );
  AND U6466 ( .A(n5230), .B(n5231), .Z(n5228) );
  NAND U6467 ( .A(ereg[84]), .B(n4895), .Z(n5231) );
  NANDN U6468 ( .A(n4890), .B(ereg[85]), .Z(n5230) );
  NAND U6469 ( .A(n5232), .B(n5233), .Z(n3772) );
  NANDN U6470 ( .A(init), .B(e[86]), .Z(n5233) );
  AND U6471 ( .A(n5234), .B(n5235), .Z(n5232) );
  NAND U6472 ( .A(ereg[85]), .B(n4895), .Z(n5235) );
  NANDN U6473 ( .A(n4890), .B(ereg[86]), .Z(n5234) );
  NAND U6474 ( .A(n5236), .B(n5237), .Z(n3771) );
  NANDN U6475 ( .A(init), .B(e[87]), .Z(n5237) );
  AND U6476 ( .A(n5238), .B(n5239), .Z(n5236) );
  NAND U6477 ( .A(ereg[86]), .B(n4895), .Z(n5239) );
  NANDN U6478 ( .A(n4890), .B(ereg[87]), .Z(n5238) );
  NAND U6479 ( .A(n5240), .B(n5241), .Z(n3770) );
  NANDN U6480 ( .A(init), .B(e[88]), .Z(n5241) );
  AND U6481 ( .A(n5242), .B(n5243), .Z(n5240) );
  NAND U6482 ( .A(ereg[87]), .B(n4895), .Z(n5243) );
  NANDN U6483 ( .A(n4890), .B(ereg[88]), .Z(n5242) );
  NAND U6484 ( .A(n5244), .B(n5245), .Z(n3769) );
  NANDN U6485 ( .A(init), .B(e[89]), .Z(n5245) );
  AND U6486 ( .A(n5246), .B(n5247), .Z(n5244) );
  NAND U6487 ( .A(ereg[88]), .B(n4895), .Z(n5247) );
  NANDN U6488 ( .A(n4890), .B(ereg[89]), .Z(n5246) );
  NAND U6489 ( .A(n5248), .B(n5249), .Z(n3768) );
  NANDN U6490 ( .A(init), .B(e[90]), .Z(n5249) );
  AND U6491 ( .A(n5250), .B(n5251), .Z(n5248) );
  NAND U6492 ( .A(ereg[89]), .B(n4895), .Z(n5251) );
  NANDN U6493 ( .A(n4890), .B(ereg[90]), .Z(n5250) );
  NAND U6494 ( .A(n5252), .B(n5253), .Z(n3767) );
  NANDN U6495 ( .A(init), .B(e[91]), .Z(n5253) );
  AND U6496 ( .A(n5254), .B(n5255), .Z(n5252) );
  NAND U6497 ( .A(ereg[90]), .B(n4895), .Z(n5255) );
  NANDN U6498 ( .A(n4890), .B(ereg[91]), .Z(n5254) );
  NAND U6499 ( .A(n5256), .B(n5257), .Z(n3766) );
  NANDN U6500 ( .A(init), .B(e[92]), .Z(n5257) );
  AND U6501 ( .A(n5258), .B(n5259), .Z(n5256) );
  NAND U6502 ( .A(ereg[91]), .B(n4895), .Z(n5259) );
  NANDN U6503 ( .A(n4890), .B(ereg[92]), .Z(n5258) );
  NAND U6504 ( .A(n5260), .B(n5261), .Z(n3765) );
  NANDN U6505 ( .A(init), .B(e[93]), .Z(n5261) );
  AND U6506 ( .A(n5262), .B(n5263), .Z(n5260) );
  NAND U6507 ( .A(ereg[92]), .B(n4895), .Z(n5263) );
  NANDN U6508 ( .A(n4890), .B(ereg[93]), .Z(n5262) );
  NAND U6509 ( .A(n5264), .B(n5265), .Z(n3764) );
  NANDN U6510 ( .A(init), .B(e[94]), .Z(n5265) );
  AND U6511 ( .A(n5266), .B(n5267), .Z(n5264) );
  NAND U6512 ( .A(ereg[93]), .B(n4895), .Z(n5267) );
  NANDN U6513 ( .A(n4890), .B(ereg[94]), .Z(n5266) );
  NAND U6514 ( .A(n5268), .B(n5269), .Z(n3763) );
  NANDN U6515 ( .A(init), .B(e[95]), .Z(n5269) );
  AND U6516 ( .A(n5270), .B(n5271), .Z(n5268) );
  NAND U6517 ( .A(ereg[94]), .B(n4895), .Z(n5271) );
  NANDN U6518 ( .A(n4890), .B(ereg[95]), .Z(n5270) );
  NAND U6519 ( .A(n5272), .B(n5273), .Z(n3762) );
  NANDN U6520 ( .A(init), .B(e[96]), .Z(n5273) );
  AND U6521 ( .A(n5274), .B(n5275), .Z(n5272) );
  NAND U6522 ( .A(ereg[95]), .B(n4895), .Z(n5275) );
  NANDN U6523 ( .A(n4890), .B(ereg[96]), .Z(n5274) );
  NAND U6524 ( .A(n5276), .B(n5277), .Z(n3761) );
  NANDN U6525 ( .A(init), .B(e[97]), .Z(n5277) );
  AND U6526 ( .A(n5278), .B(n5279), .Z(n5276) );
  NAND U6527 ( .A(ereg[96]), .B(n4895), .Z(n5279) );
  NANDN U6528 ( .A(n4890), .B(ereg[97]), .Z(n5278) );
  NAND U6529 ( .A(n5280), .B(n5281), .Z(n3760) );
  NANDN U6530 ( .A(init), .B(e[98]), .Z(n5281) );
  AND U6531 ( .A(n5282), .B(n5283), .Z(n5280) );
  NAND U6532 ( .A(ereg[97]), .B(n4895), .Z(n5283) );
  NANDN U6533 ( .A(n4890), .B(ereg[98]), .Z(n5282) );
  NAND U6534 ( .A(n5284), .B(n5285), .Z(n3759) );
  NANDN U6535 ( .A(init), .B(e[99]), .Z(n5285) );
  AND U6536 ( .A(n5286), .B(n5287), .Z(n5284) );
  NAND U6537 ( .A(ereg[98]), .B(n4895), .Z(n5287) );
  NANDN U6538 ( .A(n4890), .B(ereg[99]), .Z(n5286) );
  NAND U6539 ( .A(n5288), .B(n5289), .Z(n3758) );
  NANDN U6540 ( .A(init), .B(e[100]), .Z(n5289) );
  AND U6541 ( .A(n5290), .B(n5291), .Z(n5288) );
  NAND U6542 ( .A(ereg[99]), .B(n4895), .Z(n5291) );
  NANDN U6543 ( .A(n4890), .B(ereg[100]), .Z(n5290) );
  NAND U6544 ( .A(n5292), .B(n5293), .Z(n3757) );
  NANDN U6545 ( .A(init), .B(e[101]), .Z(n5293) );
  AND U6546 ( .A(n5294), .B(n5295), .Z(n5292) );
  NAND U6547 ( .A(ereg[100]), .B(n4895), .Z(n5295) );
  NANDN U6548 ( .A(n4890), .B(ereg[101]), .Z(n5294) );
  NAND U6549 ( .A(n5296), .B(n5297), .Z(n3756) );
  NANDN U6550 ( .A(init), .B(e[102]), .Z(n5297) );
  AND U6551 ( .A(n5298), .B(n5299), .Z(n5296) );
  NAND U6552 ( .A(ereg[101]), .B(n4895), .Z(n5299) );
  NANDN U6553 ( .A(n4890), .B(ereg[102]), .Z(n5298) );
  NAND U6554 ( .A(n5300), .B(n5301), .Z(n3755) );
  NANDN U6555 ( .A(init), .B(e[103]), .Z(n5301) );
  AND U6556 ( .A(n5302), .B(n5303), .Z(n5300) );
  NAND U6557 ( .A(ereg[102]), .B(n4895), .Z(n5303) );
  NANDN U6558 ( .A(n4890), .B(ereg[103]), .Z(n5302) );
  NAND U6559 ( .A(n5304), .B(n5305), .Z(n3754) );
  NANDN U6560 ( .A(init), .B(e[104]), .Z(n5305) );
  AND U6561 ( .A(n5306), .B(n5307), .Z(n5304) );
  NAND U6562 ( .A(ereg[103]), .B(n4895), .Z(n5307) );
  NANDN U6563 ( .A(n4890), .B(ereg[104]), .Z(n5306) );
  NAND U6564 ( .A(n5308), .B(n5309), .Z(n3753) );
  NANDN U6565 ( .A(init), .B(e[105]), .Z(n5309) );
  AND U6566 ( .A(n5310), .B(n5311), .Z(n5308) );
  NAND U6567 ( .A(ereg[104]), .B(n4895), .Z(n5311) );
  NANDN U6568 ( .A(n4890), .B(ereg[105]), .Z(n5310) );
  NAND U6569 ( .A(n5312), .B(n5313), .Z(n3752) );
  NANDN U6570 ( .A(init), .B(e[106]), .Z(n5313) );
  AND U6571 ( .A(n5314), .B(n5315), .Z(n5312) );
  NAND U6572 ( .A(ereg[105]), .B(n4895), .Z(n5315) );
  NANDN U6573 ( .A(n4890), .B(ereg[106]), .Z(n5314) );
  NAND U6574 ( .A(n5316), .B(n5317), .Z(n3751) );
  NANDN U6575 ( .A(init), .B(e[107]), .Z(n5317) );
  AND U6576 ( .A(n5318), .B(n5319), .Z(n5316) );
  NAND U6577 ( .A(ereg[106]), .B(n4895), .Z(n5319) );
  NANDN U6578 ( .A(n4890), .B(ereg[107]), .Z(n5318) );
  NAND U6579 ( .A(n5320), .B(n5321), .Z(n3750) );
  NANDN U6580 ( .A(init), .B(e[108]), .Z(n5321) );
  AND U6581 ( .A(n5322), .B(n5323), .Z(n5320) );
  NAND U6582 ( .A(ereg[107]), .B(n4895), .Z(n5323) );
  NANDN U6583 ( .A(n4890), .B(ereg[108]), .Z(n5322) );
  NAND U6584 ( .A(n5324), .B(n5325), .Z(n3749) );
  NANDN U6585 ( .A(init), .B(e[109]), .Z(n5325) );
  AND U6586 ( .A(n5326), .B(n5327), .Z(n5324) );
  NAND U6587 ( .A(ereg[108]), .B(n4895), .Z(n5327) );
  NANDN U6588 ( .A(n4890), .B(ereg[109]), .Z(n5326) );
  NAND U6589 ( .A(n5328), .B(n5329), .Z(n3748) );
  NANDN U6590 ( .A(init), .B(e[110]), .Z(n5329) );
  AND U6591 ( .A(n5330), .B(n5331), .Z(n5328) );
  NAND U6592 ( .A(ereg[109]), .B(n4895), .Z(n5331) );
  NANDN U6593 ( .A(n4890), .B(ereg[110]), .Z(n5330) );
  NAND U6594 ( .A(n5332), .B(n5333), .Z(n3747) );
  NANDN U6595 ( .A(init), .B(e[111]), .Z(n5333) );
  AND U6596 ( .A(n5334), .B(n5335), .Z(n5332) );
  NAND U6597 ( .A(ereg[110]), .B(n4895), .Z(n5335) );
  NANDN U6598 ( .A(n4890), .B(ereg[111]), .Z(n5334) );
  NAND U6599 ( .A(n5336), .B(n5337), .Z(n3746) );
  NANDN U6600 ( .A(init), .B(e[112]), .Z(n5337) );
  AND U6601 ( .A(n5338), .B(n5339), .Z(n5336) );
  NAND U6602 ( .A(ereg[111]), .B(n4895), .Z(n5339) );
  NANDN U6603 ( .A(n4890), .B(ereg[112]), .Z(n5338) );
  NAND U6604 ( .A(n5340), .B(n5341), .Z(n3745) );
  NANDN U6605 ( .A(init), .B(e[113]), .Z(n5341) );
  AND U6606 ( .A(n5342), .B(n5343), .Z(n5340) );
  NAND U6607 ( .A(ereg[112]), .B(n4895), .Z(n5343) );
  NANDN U6608 ( .A(n4890), .B(ereg[113]), .Z(n5342) );
  NAND U6609 ( .A(n5344), .B(n5345), .Z(n3744) );
  NANDN U6610 ( .A(init), .B(e[114]), .Z(n5345) );
  AND U6611 ( .A(n5346), .B(n5347), .Z(n5344) );
  NAND U6612 ( .A(ereg[113]), .B(n4895), .Z(n5347) );
  NANDN U6613 ( .A(n4890), .B(ereg[114]), .Z(n5346) );
  NAND U6614 ( .A(n5348), .B(n5349), .Z(n3743) );
  NANDN U6615 ( .A(init), .B(e[115]), .Z(n5349) );
  AND U6616 ( .A(n5350), .B(n5351), .Z(n5348) );
  NAND U6617 ( .A(ereg[114]), .B(n4895), .Z(n5351) );
  NANDN U6618 ( .A(n4890), .B(ereg[115]), .Z(n5350) );
  NAND U6619 ( .A(n5352), .B(n5353), .Z(n3742) );
  NANDN U6620 ( .A(init), .B(e[116]), .Z(n5353) );
  AND U6621 ( .A(n5354), .B(n5355), .Z(n5352) );
  NAND U6622 ( .A(ereg[115]), .B(n4895), .Z(n5355) );
  NANDN U6623 ( .A(n4890), .B(ereg[116]), .Z(n5354) );
  NAND U6624 ( .A(n5356), .B(n5357), .Z(n3741) );
  NANDN U6625 ( .A(init), .B(e[117]), .Z(n5357) );
  AND U6626 ( .A(n5358), .B(n5359), .Z(n5356) );
  NAND U6627 ( .A(ereg[116]), .B(n4895), .Z(n5359) );
  NANDN U6628 ( .A(n4890), .B(ereg[117]), .Z(n5358) );
  NAND U6629 ( .A(n5360), .B(n5361), .Z(n3740) );
  NANDN U6630 ( .A(init), .B(e[118]), .Z(n5361) );
  AND U6631 ( .A(n5362), .B(n5363), .Z(n5360) );
  NAND U6632 ( .A(ereg[117]), .B(n4895), .Z(n5363) );
  NANDN U6633 ( .A(n4890), .B(ereg[118]), .Z(n5362) );
  NAND U6634 ( .A(n5364), .B(n5365), .Z(n3739) );
  NANDN U6635 ( .A(init), .B(e[119]), .Z(n5365) );
  AND U6636 ( .A(n5366), .B(n5367), .Z(n5364) );
  NAND U6637 ( .A(ereg[118]), .B(n4895), .Z(n5367) );
  NANDN U6638 ( .A(n4890), .B(ereg[119]), .Z(n5366) );
  NAND U6639 ( .A(n5368), .B(n5369), .Z(n3738) );
  NANDN U6640 ( .A(init), .B(e[120]), .Z(n5369) );
  AND U6641 ( .A(n5370), .B(n5371), .Z(n5368) );
  NAND U6642 ( .A(ereg[119]), .B(n4895), .Z(n5371) );
  NANDN U6643 ( .A(n4890), .B(ereg[120]), .Z(n5370) );
  NAND U6644 ( .A(n5372), .B(n5373), .Z(n3737) );
  NANDN U6645 ( .A(init), .B(e[121]), .Z(n5373) );
  AND U6646 ( .A(n5374), .B(n5375), .Z(n5372) );
  NAND U6647 ( .A(ereg[120]), .B(n4895), .Z(n5375) );
  NANDN U6648 ( .A(n4890), .B(ereg[121]), .Z(n5374) );
  NAND U6649 ( .A(n5376), .B(n5377), .Z(n3736) );
  NANDN U6650 ( .A(init), .B(e[122]), .Z(n5377) );
  AND U6651 ( .A(n5378), .B(n5379), .Z(n5376) );
  NAND U6652 ( .A(ereg[121]), .B(n4895), .Z(n5379) );
  NANDN U6653 ( .A(n4890), .B(ereg[122]), .Z(n5378) );
  NAND U6654 ( .A(n5380), .B(n5381), .Z(n3735) );
  NANDN U6655 ( .A(init), .B(e[123]), .Z(n5381) );
  AND U6656 ( .A(n5382), .B(n5383), .Z(n5380) );
  NAND U6657 ( .A(ereg[122]), .B(n4895), .Z(n5383) );
  NANDN U6658 ( .A(n4890), .B(ereg[123]), .Z(n5382) );
  NAND U6659 ( .A(n5384), .B(n5385), .Z(n3734) );
  NANDN U6660 ( .A(init), .B(e[124]), .Z(n5385) );
  AND U6661 ( .A(n5386), .B(n5387), .Z(n5384) );
  NAND U6662 ( .A(ereg[123]), .B(n4895), .Z(n5387) );
  NANDN U6663 ( .A(n4890), .B(ereg[124]), .Z(n5386) );
  NAND U6664 ( .A(n5388), .B(n5389), .Z(n3733) );
  NANDN U6665 ( .A(init), .B(e[125]), .Z(n5389) );
  AND U6666 ( .A(n5390), .B(n5391), .Z(n5388) );
  NAND U6667 ( .A(ereg[124]), .B(n4895), .Z(n5391) );
  NANDN U6668 ( .A(n4890), .B(ereg[125]), .Z(n5390) );
  NAND U6669 ( .A(n5392), .B(n5393), .Z(n3732) );
  NANDN U6670 ( .A(init), .B(e[126]), .Z(n5393) );
  AND U6671 ( .A(n5394), .B(n5395), .Z(n5392) );
  NAND U6672 ( .A(ereg[125]), .B(n4895), .Z(n5395) );
  NANDN U6673 ( .A(n4890), .B(ereg[126]), .Z(n5394) );
  NAND U6674 ( .A(n5396), .B(n5397), .Z(n3731) );
  NANDN U6675 ( .A(init), .B(e[127]), .Z(n5397) );
  AND U6676 ( .A(n5398), .B(n5399), .Z(n5396) );
  NAND U6677 ( .A(ereg[126]), .B(n4895), .Z(n5399) );
  NANDN U6678 ( .A(n4890), .B(ereg[127]), .Z(n5398) );
  NAND U6679 ( .A(n5400), .B(n5401), .Z(n3730) );
  NANDN U6680 ( .A(init), .B(e[128]), .Z(n5401) );
  AND U6681 ( .A(n5402), .B(n5403), .Z(n5400) );
  NAND U6682 ( .A(ereg[127]), .B(n4895), .Z(n5403) );
  NANDN U6683 ( .A(n4890), .B(ereg[128]), .Z(n5402) );
  NAND U6684 ( .A(n5404), .B(n5405), .Z(n3729) );
  NANDN U6685 ( .A(init), .B(e[129]), .Z(n5405) );
  AND U6686 ( .A(n5406), .B(n5407), .Z(n5404) );
  NAND U6687 ( .A(ereg[128]), .B(n4895), .Z(n5407) );
  NANDN U6688 ( .A(n4890), .B(ereg[129]), .Z(n5406) );
  NAND U6689 ( .A(n5408), .B(n5409), .Z(n3728) );
  NANDN U6690 ( .A(init), .B(e[130]), .Z(n5409) );
  AND U6691 ( .A(n5410), .B(n5411), .Z(n5408) );
  NAND U6692 ( .A(ereg[129]), .B(n4895), .Z(n5411) );
  NANDN U6693 ( .A(n4890), .B(ereg[130]), .Z(n5410) );
  NAND U6694 ( .A(n5412), .B(n5413), .Z(n3727) );
  NANDN U6695 ( .A(init), .B(e[131]), .Z(n5413) );
  AND U6696 ( .A(n5414), .B(n5415), .Z(n5412) );
  NAND U6697 ( .A(ereg[130]), .B(n4895), .Z(n5415) );
  NANDN U6698 ( .A(n4890), .B(ereg[131]), .Z(n5414) );
  NAND U6699 ( .A(n5416), .B(n5417), .Z(n3726) );
  NANDN U6700 ( .A(init), .B(e[132]), .Z(n5417) );
  AND U6701 ( .A(n5418), .B(n5419), .Z(n5416) );
  NAND U6702 ( .A(ereg[131]), .B(n4895), .Z(n5419) );
  NANDN U6703 ( .A(n4890), .B(ereg[132]), .Z(n5418) );
  NAND U6704 ( .A(n5420), .B(n5421), .Z(n3725) );
  NANDN U6705 ( .A(init), .B(e[133]), .Z(n5421) );
  AND U6706 ( .A(n5422), .B(n5423), .Z(n5420) );
  NAND U6707 ( .A(ereg[132]), .B(n4895), .Z(n5423) );
  NANDN U6708 ( .A(n4890), .B(ereg[133]), .Z(n5422) );
  NAND U6709 ( .A(n5424), .B(n5425), .Z(n3724) );
  NANDN U6710 ( .A(init), .B(e[134]), .Z(n5425) );
  AND U6711 ( .A(n5426), .B(n5427), .Z(n5424) );
  NAND U6712 ( .A(ereg[133]), .B(n4895), .Z(n5427) );
  NANDN U6713 ( .A(n4890), .B(ereg[134]), .Z(n5426) );
  NAND U6714 ( .A(n5428), .B(n5429), .Z(n3723) );
  NANDN U6715 ( .A(init), .B(e[135]), .Z(n5429) );
  AND U6716 ( .A(n5430), .B(n5431), .Z(n5428) );
  NAND U6717 ( .A(ereg[134]), .B(n4895), .Z(n5431) );
  NANDN U6718 ( .A(n4890), .B(ereg[135]), .Z(n5430) );
  NAND U6719 ( .A(n5432), .B(n5433), .Z(n3722) );
  NANDN U6720 ( .A(init), .B(e[136]), .Z(n5433) );
  AND U6721 ( .A(n5434), .B(n5435), .Z(n5432) );
  NAND U6722 ( .A(ereg[135]), .B(n4895), .Z(n5435) );
  NANDN U6723 ( .A(n4890), .B(ereg[136]), .Z(n5434) );
  NAND U6724 ( .A(n5436), .B(n5437), .Z(n3721) );
  NANDN U6725 ( .A(init), .B(e[137]), .Z(n5437) );
  AND U6726 ( .A(n5438), .B(n5439), .Z(n5436) );
  NAND U6727 ( .A(ereg[136]), .B(n4895), .Z(n5439) );
  NANDN U6728 ( .A(n4890), .B(ereg[137]), .Z(n5438) );
  NAND U6729 ( .A(n5440), .B(n5441), .Z(n3720) );
  NANDN U6730 ( .A(init), .B(e[138]), .Z(n5441) );
  AND U6731 ( .A(n5442), .B(n5443), .Z(n5440) );
  NAND U6732 ( .A(ereg[137]), .B(n4895), .Z(n5443) );
  NANDN U6733 ( .A(n4890), .B(ereg[138]), .Z(n5442) );
  NAND U6734 ( .A(n5444), .B(n5445), .Z(n3719) );
  NANDN U6735 ( .A(init), .B(e[139]), .Z(n5445) );
  AND U6736 ( .A(n5446), .B(n5447), .Z(n5444) );
  NAND U6737 ( .A(ereg[138]), .B(n4895), .Z(n5447) );
  NANDN U6738 ( .A(n4890), .B(ereg[139]), .Z(n5446) );
  NAND U6739 ( .A(n5448), .B(n5449), .Z(n3718) );
  NANDN U6740 ( .A(init), .B(e[140]), .Z(n5449) );
  AND U6741 ( .A(n5450), .B(n5451), .Z(n5448) );
  NAND U6742 ( .A(ereg[139]), .B(n4895), .Z(n5451) );
  NANDN U6743 ( .A(n4890), .B(ereg[140]), .Z(n5450) );
  NAND U6744 ( .A(n5452), .B(n5453), .Z(n3717) );
  NANDN U6745 ( .A(init), .B(e[141]), .Z(n5453) );
  AND U6746 ( .A(n5454), .B(n5455), .Z(n5452) );
  NAND U6747 ( .A(ereg[140]), .B(n4895), .Z(n5455) );
  NANDN U6748 ( .A(n4890), .B(ereg[141]), .Z(n5454) );
  NAND U6749 ( .A(n5456), .B(n5457), .Z(n3716) );
  NANDN U6750 ( .A(init), .B(e[142]), .Z(n5457) );
  AND U6751 ( .A(n5458), .B(n5459), .Z(n5456) );
  NAND U6752 ( .A(ereg[141]), .B(n4895), .Z(n5459) );
  NANDN U6753 ( .A(n4890), .B(ereg[142]), .Z(n5458) );
  NAND U6754 ( .A(n5460), .B(n5461), .Z(n3715) );
  NANDN U6755 ( .A(init), .B(e[143]), .Z(n5461) );
  AND U6756 ( .A(n5462), .B(n5463), .Z(n5460) );
  NAND U6757 ( .A(ereg[142]), .B(n4895), .Z(n5463) );
  NANDN U6758 ( .A(n4890), .B(ereg[143]), .Z(n5462) );
  NAND U6759 ( .A(n5464), .B(n5465), .Z(n3714) );
  NANDN U6760 ( .A(init), .B(e[144]), .Z(n5465) );
  AND U6761 ( .A(n5466), .B(n5467), .Z(n5464) );
  NAND U6762 ( .A(ereg[143]), .B(n4895), .Z(n5467) );
  NANDN U6763 ( .A(n4890), .B(ereg[144]), .Z(n5466) );
  NAND U6764 ( .A(n5468), .B(n5469), .Z(n3713) );
  NANDN U6765 ( .A(init), .B(e[145]), .Z(n5469) );
  AND U6766 ( .A(n5470), .B(n5471), .Z(n5468) );
  NAND U6767 ( .A(ereg[144]), .B(n4895), .Z(n5471) );
  NANDN U6768 ( .A(n4890), .B(ereg[145]), .Z(n5470) );
  NAND U6769 ( .A(n5472), .B(n5473), .Z(n3712) );
  NANDN U6770 ( .A(init), .B(e[146]), .Z(n5473) );
  AND U6771 ( .A(n5474), .B(n5475), .Z(n5472) );
  NAND U6772 ( .A(ereg[145]), .B(n4895), .Z(n5475) );
  NANDN U6773 ( .A(n4890), .B(ereg[146]), .Z(n5474) );
  NAND U6774 ( .A(n5476), .B(n5477), .Z(n3711) );
  NANDN U6775 ( .A(init), .B(e[147]), .Z(n5477) );
  AND U6776 ( .A(n5478), .B(n5479), .Z(n5476) );
  NAND U6777 ( .A(ereg[146]), .B(n4895), .Z(n5479) );
  NANDN U6778 ( .A(n4890), .B(ereg[147]), .Z(n5478) );
  NAND U6779 ( .A(n5480), .B(n5481), .Z(n3710) );
  NANDN U6780 ( .A(init), .B(e[148]), .Z(n5481) );
  AND U6781 ( .A(n5482), .B(n5483), .Z(n5480) );
  NAND U6782 ( .A(ereg[147]), .B(n4895), .Z(n5483) );
  NANDN U6783 ( .A(n4890), .B(ereg[148]), .Z(n5482) );
  NAND U6784 ( .A(n5484), .B(n5485), .Z(n3709) );
  NANDN U6785 ( .A(init), .B(e[149]), .Z(n5485) );
  AND U6786 ( .A(n5486), .B(n5487), .Z(n5484) );
  NAND U6787 ( .A(ereg[148]), .B(n4895), .Z(n5487) );
  NANDN U6788 ( .A(n4890), .B(ereg[149]), .Z(n5486) );
  NAND U6789 ( .A(n5488), .B(n5489), .Z(n3708) );
  NANDN U6790 ( .A(init), .B(e[150]), .Z(n5489) );
  AND U6791 ( .A(n5490), .B(n5491), .Z(n5488) );
  NAND U6792 ( .A(ereg[149]), .B(n4895), .Z(n5491) );
  NANDN U6793 ( .A(n4890), .B(ereg[150]), .Z(n5490) );
  NAND U6794 ( .A(n5492), .B(n5493), .Z(n3707) );
  NANDN U6795 ( .A(init), .B(e[151]), .Z(n5493) );
  AND U6796 ( .A(n5494), .B(n5495), .Z(n5492) );
  NAND U6797 ( .A(ereg[150]), .B(n4895), .Z(n5495) );
  NANDN U6798 ( .A(n4890), .B(ereg[151]), .Z(n5494) );
  NAND U6799 ( .A(n5496), .B(n5497), .Z(n3706) );
  NANDN U6800 ( .A(init), .B(e[152]), .Z(n5497) );
  AND U6801 ( .A(n5498), .B(n5499), .Z(n5496) );
  NAND U6802 ( .A(ereg[151]), .B(n4895), .Z(n5499) );
  NANDN U6803 ( .A(n4890), .B(ereg[152]), .Z(n5498) );
  NAND U6804 ( .A(n5500), .B(n5501), .Z(n3705) );
  NANDN U6805 ( .A(init), .B(e[153]), .Z(n5501) );
  AND U6806 ( .A(n5502), .B(n5503), .Z(n5500) );
  NAND U6807 ( .A(ereg[152]), .B(n4895), .Z(n5503) );
  NANDN U6808 ( .A(n4890), .B(ereg[153]), .Z(n5502) );
  NAND U6809 ( .A(n5504), .B(n5505), .Z(n3704) );
  NANDN U6810 ( .A(init), .B(e[154]), .Z(n5505) );
  AND U6811 ( .A(n5506), .B(n5507), .Z(n5504) );
  NAND U6812 ( .A(ereg[153]), .B(n4895), .Z(n5507) );
  NANDN U6813 ( .A(n4890), .B(ereg[154]), .Z(n5506) );
  NAND U6814 ( .A(n5508), .B(n5509), .Z(n3703) );
  NANDN U6815 ( .A(init), .B(e[155]), .Z(n5509) );
  AND U6816 ( .A(n5510), .B(n5511), .Z(n5508) );
  NAND U6817 ( .A(ereg[154]), .B(n4895), .Z(n5511) );
  NANDN U6818 ( .A(n4890), .B(ereg[155]), .Z(n5510) );
  NAND U6819 ( .A(n5512), .B(n5513), .Z(n3702) );
  NANDN U6820 ( .A(init), .B(e[156]), .Z(n5513) );
  AND U6821 ( .A(n5514), .B(n5515), .Z(n5512) );
  NAND U6822 ( .A(ereg[155]), .B(n4895), .Z(n5515) );
  NANDN U6823 ( .A(n4890), .B(ereg[156]), .Z(n5514) );
  NAND U6824 ( .A(n5516), .B(n5517), .Z(n3701) );
  NANDN U6825 ( .A(init), .B(e[157]), .Z(n5517) );
  AND U6826 ( .A(n5518), .B(n5519), .Z(n5516) );
  NAND U6827 ( .A(ereg[156]), .B(n4895), .Z(n5519) );
  NANDN U6828 ( .A(n4890), .B(ereg[157]), .Z(n5518) );
  NAND U6829 ( .A(n5520), .B(n5521), .Z(n3700) );
  NANDN U6830 ( .A(init), .B(e[158]), .Z(n5521) );
  AND U6831 ( .A(n5522), .B(n5523), .Z(n5520) );
  NAND U6832 ( .A(ereg[157]), .B(n4895), .Z(n5523) );
  NANDN U6833 ( .A(n4890), .B(ereg[158]), .Z(n5522) );
  NAND U6834 ( .A(n5524), .B(n5525), .Z(n3699) );
  NANDN U6835 ( .A(init), .B(e[159]), .Z(n5525) );
  AND U6836 ( .A(n5526), .B(n5527), .Z(n5524) );
  NAND U6837 ( .A(ereg[158]), .B(n4895), .Z(n5527) );
  NANDN U6838 ( .A(n4890), .B(ereg[159]), .Z(n5526) );
  NAND U6839 ( .A(n5528), .B(n5529), .Z(n3698) );
  NANDN U6840 ( .A(init), .B(e[160]), .Z(n5529) );
  AND U6841 ( .A(n5530), .B(n5531), .Z(n5528) );
  NAND U6842 ( .A(ereg[159]), .B(n4895), .Z(n5531) );
  NANDN U6843 ( .A(n4890), .B(ereg[160]), .Z(n5530) );
  NAND U6844 ( .A(n5532), .B(n5533), .Z(n3697) );
  NANDN U6845 ( .A(init), .B(e[161]), .Z(n5533) );
  AND U6846 ( .A(n5534), .B(n5535), .Z(n5532) );
  NAND U6847 ( .A(ereg[160]), .B(n4895), .Z(n5535) );
  NANDN U6848 ( .A(n4890), .B(ereg[161]), .Z(n5534) );
  NAND U6849 ( .A(n5536), .B(n5537), .Z(n3696) );
  NANDN U6850 ( .A(init), .B(e[162]), .Z(n5537) );
  AND U6851 ( .A(n5538), .B(n5539), .Z(n5536) );
  NAND U6852 ( .A(ereg[161]), .B(n4895), .Z(n5539) );
  NANDN U6853 ( .A(n4890), .B(ereg[162]), .Z(n5538) );
  NAND U6854 ( .A(n5540), .B(n5541), .Z(n3695) );
  NANDN U6855 ( .A(init), .B(e[163]), .Z(n5541) );
  AND U6856 ( .A(n5542), .B(n5543), .Z(n5540) );
  NAND U6857 ( .A(ereg[162]), .B(n4895), .Z(n5543) );
  NANDN U6858 ( .A(n4890), .B(ereg[163]), .Z(n5542) );
  NAND U6859 ( .A(n5544), .B(n5545), .Z(n3694) );
  NANDN U6860 ( .A(init), .B(e[164]), .Z(n5545) );
  AND U6861 ( .A(n5546), .B(n5547), .Z(n5544) );
  NAND U6862 ( .A(ereg[163]), .B(n4895), .Z(n5547) );
  NANDN U6863 ( .A(n4890), .B(ereg[164]), .Z(n5546) );
  NAND U6864 ( .A(n5548), .B(n5549), .Z(n3693) );
  NANDN U6865 ( .A(init), .B(e[165]), .Z(n5549) );
  AND U6866 ( .A(n5550), .B(n5551), .Z(n5548) );
  NAND U6867 ( .A(ereg[164]), .B(n4895), .Z(n5551) );
  NANDN U6868 ( .A(n4890), .B(ereg[165]), .Z(n5550) );
  NAND U6869 ( .A(n5552), .B(n5553), .Z(n3692) );
  NANDN U6870 ( .A(init), .B(e[166]), .Z(n5553) );
  AND U6871 ( .A(n5554), .B(n5555), .Z(n5552) );
  NAND U6872 ( .A(ereg[165]), .B(n4895), .Z(n5555) );
  NANDN U6873 ( .A(n4890), .B(ereg[166]), .Z(n5554) );
  NAND U6874 ( .A(n5556), .B(n5557), .Z(n3691) );
  NANDN U6875 ( .A(init), .B(e[167]), .Z(n5557) );
  AND U6876 ( .A(n5558), .B(n5559), .Z(n5556) );
  NAND U6877 ( .A(ereg[166]), .B(n4895), .Z(n5559) );
  NANDN U6878 ( .A(n4890), .B(ereg[167]), .Z(n5558) );
  NAND U6879 ( .A(n5560), .B(n5561), .Z(n3690) );
  NANDN U6880 ( .A(init), .B(e[168]), .Z(n5561) );
  AND U6881 ( .A(n5562), .B(n5563), .Z(n5560) );
  NAND U6882 ( .A(ereg[167]), .B(n4895), .Z(n5563) );
  NANDN U6883 ( .A(n4890), .B(ereg[168]), .Z(n5562) );
  NAND U6884 ( .A(n5564), .B(n5565), .Z(n3689) );
  NANDN U6885 ( .A(init), .B(e[169]), .Z(n5565) );
  AND U6886 ( .A(n5566), .B(n5567), .Z(n5564) );
  NAND U6887 ( .A(ereg[168]), .B(n4895), .Z(n5567) );
  NANDN U6888 ( .A(n4890), .B(ereg[169]), .Z(n5566) );
  NAND U6889 ( .A(n5568), .B(n5569), .Z(n3688) );
  NANDN U6890 ( .A(init), .B(e[170]), .Z(n5569) );
  AND U6891 ( .A(n5570), .B(n5571), .Z(n5568) );
  NAND U6892 ( .A(ereg[169]), .B(n4895), .Z(n5571) );
  NANDN U6893 ( .A(n4890), .B(ereg[170]), .Z(n5570) );
  NAND U6894 ( .A(n5572), .B(n5573), .Z(n3687) );
  NANDN U6895 ( .A(init), .B(e[171]), .Z(n5573) );
  AND U6896 ( .A(n5574), .B(n5575), .Z(n5572) );
  NAND U6897 ( .A(ereg[170]), .B(n4895), .Z(n5575) );
  NANDN U6898 ( .A(n4890), .B(ereg[171]), .Z(n5574) );
  NAND U6899 ( .A(n5576), .B(n5577), .Z(n3686) );
  NANDN U6900 ( .A(init), .B(e[172]), .Z(n5577) );
  AND U6901 ( .A(n5578), .B(n5579), .Z(n5576) );
  NAND U6902 ( .A(ereg[171]), .B(n4895), .Z(n5579) );
  NANDN U6903 ( .A(n4890), .B(ereg[172]), .Z(n5578) );
  NAND U6904 ( .A(n5580), .B(n5581), .Z(n3685) );
  NANDN U6905 ( .A(init), .B(e[173]), .Z(n5581) );
  AND U6906 ( .A(n5582), .B(n5583), .Z(n5580) );
  NAND U6907 ( .A(ereg[172]), .B(n4895), .Z(n5583) );
  NANDN U6908 ( .A(n4890), .B(ereg[173]), .Z(n5582) );
  NAND U6909 ( .A(n5584), .B(n5585), .Z(n3684) );
  NANDN U6910 ( .A(init), .B(e[174]), .Z(n5585) );
  AND U6911 ( .A(n5586), .B(n5587), .Z(n5584) );
  NAND U6912 ( .A(ereg[173]), .B(n4895), .Z(n5587) );
  NANDN U6913 ( .A(n4890), .B(ereg[174]), .Z(n5586) );
  NAND U6914 ( .A(n5588), .B(n5589), .Z(n3683) );
  NANDN U6915 ( .A(init), .B(e[175]), .Z(n5589) );
  AND U6916 ( .A(n5590), .B(n5591), .Z(n5588) );
  NAND U6917 ( .A(ereg[174]), .B(n4895), .Z(n5591) );
  NANDN U6918 ( .A(n4890), .B(ereg[175]), .Z(n5590) );
  NAND U6919 ( .A(n5592), .B(n5593), .Z(n3682) );
  NANDN U6920 ( .A(init), .B(e[176]), .Z(n5593) );
  AND U6921 ( .A(n5594), .B(n5595), .Z(n5592) );
  NAND U6922 ( .A(ereg[175]), .B(n4895), .Z(n5595) );
  NANDN U6923 ( .A(n4890), .B(ereg[176]), .Z(n5594) );
  NAND U6924 ( .A(n5596), .B(n5597), .Z(n3681) );
  NANDN U6925 ( .A(init), .B(e[177]), .Z(n5597) );
  AND U6926 ( .A(n5598), .B(n5599), .Z(n5596) );
  NAND U6927 ( .A(ereg[176]), .B(n4895), .Z(n5599) );
  NANDN U6928 ( .A(n4890), .B(ereg[177]), .Z(n5598) );
  NAND U6929 ( .A(n5600), .B(n5601), .Z(n3680) );
  NANDN U6930 ( .A(init), .B(e[178]), .Z(n5601) );
  AND U6931 ( .A(n5602), .B(n5603), .Z(n5600) );
  NAND U6932 ( .A(ereg[177]), .B(n4895), .Z(n5603) );
  NANDN U6933 ( .A(n4890), .B(ereg[178]), .Z(n5602) );
  NAND U6934 ( .A(n5604), .B(n5605), .Z(n3679) );
  NANDN U6935 ( .A(init), .B(e[179]), .Z(n5605) );
  AND U6936 ( .A(n5606), .B(n5607), .Z(n5604) );
  NAND U6937 ( .A(ereg[178]), .B(n4895), .Z(n5607) );
  NANDN U6938 ( .A(n4890), .B(ereg[179]), .Z(n5606) );
  NAND U6939 ( .A(n5608), .B(n5609), .Z(n3678) );
  NANDN U6940 ( .A(init), .B(e[180]), .Z(n5609) );
  AND U6941 ( .A(n5610), .B(n5611), .Z(n5608) );
  NAND U6942 ( .A(ereg[179]), .B(n4895), .Z(n5611) );
  NANDN U6943 ( .A(n4890), .B(ereg[180]), .Z(n5610) );
  NAND U6944 ( .A(n5612), .B(n5613), .Z(n3677) );
  NANDN U6945 ( .A(init), .B(e[181]), .Z(n5613) );
  AND U6946 ( .A(n5614), .B(n5615), .Z(n5612) );
  NAND U6947 ( .A(ereg[180]), .B(n4895), .Z(n5615) );
  NANDN U6948 ( .A(n4890), .B(ereg[181]), .Z(n5614) );
  NAND U6949 ( .A(n5616), .B(n5617), .Z(n3676) );
  NANDN U6950 ( .A(init), .B(e[182]), .Z(n5617) );
  AND U6951 ( .A(n5618), .B(n5619), .Z(n5616) );
  NAND U6952 ( .A(ereg[181]), .B(n4895), .Z(n5619) );
  NANDN U6953 ( .A(n4890), .B(ereg[182]), .Z(n5618) );
  NAND U6954 ( .A(n5620), .B(n5621), .Z(n3675) );
  NANDN U6955 ( .A(init), .B(e[183]), .Z(n5621) );
  AND U6956 ( .A(n5622), .B(n5623), .Z(n5620) );
  NAND U6957 ( .A(ereg[182]), .B(n4895), .Z(n5623) );
  NANDN U6958 ( .A(n4890), .B(ereg[183]), .Z(n5622) );
  NAND U6959 ( .A(n5624), .B(n5625), .Z(n3674) );
  NANDN U6960 ( .A(init), .B(e[184]), .Z(n5625) );
  AND U6961 ( .A(n5626), .B(n5627), .Z(n5624) );
  NAND U6962 ( .A(ereg[183]), .B(n4895), .Z(n5627) );
  NANDN U6963 ( .A(n4890), .B(ereg[184]), .Z(n5626) );
  NAND U6964 ( .A(n5628), .B(n5629), .Z(n3673) );
  NANDN U6965 ( .A(init), .B(e[185]), .Z(n5629) );
  AND U6966 ( .A(n5630), .B(n5631), .Z(n5628) );
  NAND U6967 ( .A(ereg[184]), .B(n4895), .Z(n5631) );
  NANDN U6968 ( .A(n4890), .B(ereg[185]), .Z(n5630) );
  NAND U6969 ( .A(n5632), .B(n5633), .Z(n3672) );
  NANDN U6970 ( .A(init), .B(e[186]), .Z(n5633) );
  AND U6971 ( .A(n5634), .B(n5635), .Z(n5632) );
  NAND U6972 ( .A(ereg[185]), .B(n4895), .Z(n5635) );
  NANDN U6973 ( .A(n4890), .B(ereg[186]), .Z(n5634) );
  NAND U6974 ( .A(n5636), .B(n5637), .Z(n3671) );
  NANDN U6975 ( .A(init), .B(e[187]), .Z(n5637) );
  AND U6976 ( .A(n5638), .B(n5639), .Z(n5636) );
  NAND U6977 ( .A(ereg[186]), .B(n4895), .Z(n5639) );
  NANDN U6978 ( .A(n4890), .B(ereg[187]), .Z(n5638) );
  NAND U6979 ( .A(n5640), .B(n5641), .Z(n3670) );
  NANDN U6980 ( .A(init), .B(e[188]), .Z(n5641) );
  AND U6981 ( .A(n5642), .B(n5643), .Z(n5640) );
  NAND U6982 ( .A(ereg[187]), .B(n4895), .Z(n5643) );
  NANDN U6983 ( .A(n4890), .B(ereg[188]), .Z(n5642) );
  NAND U6984 ( .A(n5644), .B(n5645), .Z(n3669) );
  NANDN U6985 ( .A(init), .B(e[189]), .Z(n5645) );
  AND U6986 ( .A(n5646), .B(n5647), .Z(n5644) );
  NAND U6987 ( .A(ereg[188]), .B(n4895), .Z(n5647) );
  NANDN U6988 ( .A(n4890), .B(ereg[189]), .Z(n5646) );
  NAND U6989 ( .A(n5648), .B(n5649), .Z(n3668) );
  NANDN U6990 ( .A(init), .B(e[190]), .Z(n5649) );
  AND U6991 ( .A(n5650), .B(n5651), .Z(n5648) );
  NAND U6992 ( .A(ereg[189]), .B(n4895), .Z(n5651) );
  NANDN U6993 ( .A(n4890), .B(ereg[190]), .Z(n5650) );
  NAND U6994 ( .A(n5652), .B(n5653), .Z(n3667) );
  NANDN U6995 ( .A(init), .B(e[191]), .Z(n5653) );
  AND U6996 ( .A(n5654), .B(n5655), .Z(n5652) );
  NAND U6997 ( .A(ereg[190]), .B(n4895), .Z(n5655) );
  NANDN U6998 ( .A(n4890), .B(ereg[191]), .Z(n5654) );
  NAND U6999 ( .A(n5656), .B(n5657), .Z(n3666) );
  NANDN U7000 ( .A(init), .B(e[192]), .Z(n5657) );
  AND U7001 ( .A(n5658), .B(n5659), .Z(n5656) );
  NAND U7002 ( .A(ereg[191]), .B(n4895), .Z(n5659) );
  NANDN U7003 ( .A(n4890), .B(ereg[192]), .Z(n5658) );
  NAND U7004 ( .A(n5660), .B(n5661), .Z(n3665) );
  NANDN U7005 ( .A(init), .B(e[193]), .Z(n5661) );
  AND U7006 ( .A(n5662), .B(n5663), .Z(n5660) );
  NAND U7007 ( .A(ereg[192]), .B(n4895), .Z(n5663) );
  NANDN U7008 ( .A(n4890), .B(ereg[193]), .Z(n5662) );
  NAND U7009 ( .A(n5664), .B(n5665), .Z(n3664) );
  NANDN U7010 ( .A(init), .B(e[194]), .Z(n5665) );
  AND U7011 ( .A(n5666), .B(n5667), .Z(n5664) );
  NAND U7012 ( .A(ereg[193]), .B(n4895), .Z(n5667) );
  NANDN U7013 ( .A(n4890), .B(ereg[194]), .Z(n5666) );
  NAND U7014 ( .A(n5668), .B(n5669), .Z(n3663) );
  NANDN U7015 ( .A(init), .B(e[195]), .Z(n5669) );
  AND U7016 ( .A(n5670), .B(n5671), .Z(n5668) );
  NAND U7017 ( .A(ereg[194]), .B(n4895), .Z(n5671) );
  NANDN U7018 ( .A(n4890), .B(ereg[195]), .Z(n5670) );
  NAND U7019 ( .A(n5672), .B(n5673), .Z(n3662) );
  NANDN U7020 ( .A(init), .B(e[196]), .Z(n5673) );
  AND U7021 ( .A(n5674), .B(n5675), .Z(n5672) );
  NAND U7022 ( .A(ereg[195]), .B(n4895), .Z(n5675) );
  NANDN U7023 ( .A(n4890), .B(ereg[196]), .Z(n5674) );
  NAND U7024 ( .A(n5676), .B(n5677), .Z(n3661) );
  NANDN U7025 ( .A(init), .B(e[197]), .Z(n5677) );
  AND U7026 ( .A(n5678), .B(n5679), .Z(n5676) );
  NAND U7027 ( .A(ereg[196]), .B(n4895), .Z(n5679) );
  NANDN U7028 ( .A(n4890), .B(ereg[197]), .Z(n5678) );
  NAND U7029 ( .A(n5680), .B(n5681), .Z(n3660) );
  NANDN U7030 ( .A(init), .B(e[198]), .Z(n5681) );
  AND U7031 ( .A(n5682), .B(n5683), .Z(n5680) );
  NAND U7032 ( .A(ereg[197]), .B(n4895), .Z(n5683) );
  NANDN U7033 ( .A(n4890), .B(ereg[198]), .Z(n5682) );
  NAND U7034 ( .A(n5684), .B(n5685), .Z(n3659) );
  NANDN U7035 ( .A(init), .B(e[199]), .Z(n5685) );
  AND U7036 ( .A(n5686), .B(n5687), .Z(n5684) );
  NAND U7037 ( .A(ereg[198]), .B(n4895), .Z(n5687) );
  NANDN U7038 ( .A(n4890), .B(ereg[199]), .Z(n5686) );
  NAND U7039 ( .A(n5688), .B(n5689), .Z(n3658) );
  NANDN U7040 ( .A(init), .B(e[200]), .Z(n5689) );
  AND U7041 ( .A(n5690), .B(n5691), .Z(n5688) );
  NAND U7042 ( .A(ereg[199]), .B(n4895), .Z(n5691) );
  NANDN U7043 ( .A(n4890), .B(ereg[200]), .Z(n5690) );
  NAND U7044 ( .A(n5692), .B(n5693), .Z(n3657) );
  NANDN U7045 ( .A(init), .B(e[201]), .Z(n5693) );
  AND U7046 ( .A(n5694), .B(n5695), .Z(n5692) );
  NAND U7047 ( .A(ereg[200]), .B(n4895), .Z(n5695) );
  NANDN U7048 ( .A(n4890), .B(ereg[201]), .Z(n5694) );
  NAND U7049 ( .A(n5696), .B(n5697), .Z(n3656) );
  NANDN U7050 ( .A(init), .B(e[202]), .Z(n5697) );
  AND U7051 ( .A(n5698), .B(n5699), .Z(n5696) );
  NAND U7052 ( .A(ereg[201]), .B(n4895), .Z(n5699) );
  NANDN U7053 ( .A(n4890), .B(ereg[202]), .Z(n5698) );
  NAND U7054 ( .A(n5700), .B(n5701), .Z(n3655) );
  NANDN U7055 ( .A(init), .B(e[203]), .Z(n5701) );
  AND U7056 ( .A(n5702), .B(n5703), .Z(n5700) );
  NAND U7057 ( .A(ereg[202]), .B(n4895), .Z(n5703) );
  NANDN U7058 ( .A(n4890), .B(ereg[203]), .Z(n5702) );
  NAND U7059 ( .A(n5704), .B(n5705), .Z(n3654) );
  NANDN U7060 ( .A(init), .B(e[204]), .Z(n5705) );
  AND U7061 ( .A(n5706), .B(n5707), .Z(n5704) );
  NAND U7062 ( .A(ereg[203]), .B(n4895), .Z(n5707) );
  NANDN U7063 ( .A(n4890), .B(ereg[204]), .Z(n5706) );
  NAND U7064 ( .A(n5708), .B(n5709), .Z(n3653) );
  NANDN U7065 ( .A(init), .B(e[205]), .Z(n5709) );
  AND U7066 ( .A(n5710), .B(n5711), .Z(n5708) );
  NAND U7067 ( .A(ereg[204]), .B(n4895), .Z(n5711) );
  NANDN U7068 ( .A(n4890), .B(ereg[205]), .Z(n5710) );
  NAND U7069 ( .A(n5712), .B(n5713), .Z(n3652) );
  NANDN U7070 ( .A(init), .B(e[206]), .Z(n5713) );
  AND U7071 ( .A(n5714), .B(n5715), .Z(n5712) );
  NAND U7072 ( .A(ereg[205]), .B(n4895), .Z(n5715) );
  NANDN U7073 ( .A(n4890), .B(ereg[206]), .Z(n5714) );
  NAND U7074 ( .A(n5716), .B(n5717), .Z(n3651) );
  NANDN U7075 ( .A(init), .B(e[207]), .Z(n5717) );
  AND U7076 ( .A(n5718), .B(n5719), .Z(n5716) );
  NAND U7077 ( .A(ereg[206]), .B(n4895), .Z(n5719) );
  NANDN U7078 ( .A(n4890), .B(ereg[207]), .Z(n5718) );
  NAND U7079 ( .A(n5720), .B(n5721), .Z(n3650) );
  NANDN U7080 ( .A(init), .B(e[208]), .Z(n5721) );
  AND U7081 ( .A(n5722), .B(n5723), .Z(n5720) );
  NAND U7082 ( .A(ereg[207]), .B(n4895), .Z(n5723) );
  NANDN U7083 ( .A(n4890), .B(ereg[208]), .Z(n5722) );
  NAND U7084 ( .A(n5724), .B(n5725), .Z(n3649) );
  NANDN U7085 ( .A(init), .B(e[209]), .Z(n5725) );
  AND U7086 ( .A(n5726), .B(n5727), .Z(n5724) );
  NAND U7087 ( .A(ereg[208]), .B(n4895), .Z(n5727) );
  NANDN U7088 ( .A(n4890), .B(ereg[209]), .Z(n5726) );
  NAND U7089 ( .A(n5728), .B(n5729), .Z(n3648) );
  NANDN U7090 ( .A(init), .B(e[210]), .Z(n5729) );
  AND U7091 ( .A(n5730), .B(n5731), .Z(n5728) );
  NAND U7092 ( .A(ereg[209]), .B(n4895), .Z(n5731) );
  NANDN U7093 ( .A(n4890), .B(ereg[210]), .Z(n5730) );
  NAND U7094 ( .A(n5732), .B(n5733), .Z(n3647) );
  NANDN U7095 ( .A(init), .B(e[211]), .Z(n5733) );
  AND U7096 ( .A(n5734), .B(n5735), .Z(n5732) );
  NAND U7097 ( .A(ereg[210]), .B(n4895), .Z(n5735) );
  NANDN U7098 ( .A(n4890), .B(ereg[211]), .Z(n5734) );
  NAND U7099 ( .A(n5736), .B(n5737), .Z(n3646) );
  NANDN U7100 ( .A(init), .B(e[212]), .Z(n5737) );
  AND U7101 ( .A(n5738), .B(n5739), .Z(n5736) );
  NAND U7102 ( .A(ereg[211]), .B(n4895), .Z(n5739) );
  NANDN U7103 ( .A(n4890), .B(ereg[212]), .Z(n5738) );
  NAND U7104 ( .A(n5740), .B(n5741), .Z(n3645) );
  NANDN U7105 ( .A(init), .B(e[213]), .Z(n5741) );
  AND U7106 ( .A(n5742), .B(n5743), .Z(n5740) );
  NAND U7107 ( .A(ereg[212]), .B(n4895), .Z(n5743) );
  NANDN U7108 ( .A(n4890), .B(ereg[213]), .Z(n5742) );
  NAND U7109 ( .A(n5744), .B(n5745), .Z(n3644) );
  NANDN U7110 ( .A(init), .B(e[214]), .Z(n5745) );
  AND U7111 ( .A(n5746), .B(n5747), .Z(n5744) );
  NAND U7112 ( .A(ereg[213]), .B(n4895), .Z(n5747) );
  NANDN U7113 ( .A(n4890), .B(ereg[214]), .Z(n5746) );
  NAND U7114 ( .A(n5748), .B(n5749), .Z(n3643) );
  NANDN U7115 ( .A(init), .B(e[215]), .Z(n5749) );
  AND U7116 ( .A(n5750), .B(n5751), .Z(n5748) );
  NAND U7117 ( .A(ereg[214]), .B(n4895), .Z(n5751) );
  NANDN U7118 ( .A(n4890), .B(ereg[215]), .Z(n5750) );
  NAND U7119 ( .A(n5752), .B(n5753), .Z(n3642) );
  NANDN U7120 ( .A(init), .B(e[216]), .Z(n5753) );
  AND U7121 ( .A(n5754), .B(n5755), .Z(n5752) );
  NAND U7122 ( .A(ereg[215]), .B(n4895), .Z(n5755) );
  NANDN U7123 ( .A(n4890), .B(ereg[216]), .Z(n5754) );
  NAND U7124 ( .A(n5756), .B(n5757), .Z(n3641) );
  NANDN U7125 ( .A(init), .B(e[217]), .Z(n5757) );
  AND U7126 ( .A(n5758), .B(n5759), .Z(n5756) );
  NAND U7127 ( .A(ereg[216]), .B(n4895), .Z(n5759) );
  NANDN U7128 ( .A(n4890), .B(ereg[217]), .Z(n5758) );
  NAND U7129 ( .A(n5760), .B(n5761), .Z(n3640) );
  NANDN U7130 ( .A(init), .B(e[218]), .Z(n5761) );
  AND U7131 ( .A(n5762), .B(n5763), .Z(n5760) );
  NAND U7132 ( .A(ereg[217]), .B(n4895), .Z(n5763) );
  NANDN U7133 ( .A(n4890), .B(ereg[218]), .Z(n5762) );
  NAND U7134 ( .A(n5764), .B(n5765), .Z(n3639) );
  NANDN U7135 ( .A(init), .B(e[219]), .Z(n5765) );
  AND U7136 ( .A(n5766), .B(n5767), .Z(n5764) );
  NAND U7137 ( .A(ereg[218]), .B(n4895), .Z(n5767) );
  NANDN U7138 ( .A(n4890), .B(ereg[219]), .Z(n5766) );
  NAND U7139 ( .A(n5768), .B(n5769), .Z(n3638) );
  NANDN U7140 ( .A(init), .B(e[220]), .Z(n5769) );
  AND U7141 ( .A(n5770), .B(n5771), .Z(n5768) );
  NAND U7142 ( .A(ereg[219]), .B(n4895), .Z(n5771) );
  NANDN U7143 ( .A(n4890), .B(ereg[220]), .Z(n5770) );
  NAND U7144 ( .A(n5772), .B(n5773), .Z(n3637) );
  NANDN U7145 ( .A(init), .B(e[221]), .Z(n5773) );
  AND U7146 ( .A(n5774), .B(n5775), .Z(n5772) );
  NAND U7147 ( .A(ereg[220]), .B(n4895), .Z(n5775) );
  NANDN U7148 ( .A(n4890), .B(ereg[221]), .Z(n5774) );
  NAND U7149 ( .A(n5776), .B(n5777), .Z(n3636) );
  NANDN U7150 ( .A(init), .B(e[222]), .Z(n5777) );
  AND U7151 ( .A(n5778), .B(n5779), .Z(n5776) );
  NAND U7152 ( .A(ereg[221]), .B(n4895), .Z(n5779) );
  NANDN U7153 ( .A(n4890), .B(ereg[222]), .Z(n5778) );
  NAND U7154 ( .A(n5780), .B(n5781), .Z(n3635) );
  NANDN U7155 ( .A(init), .B(e[223]), .Z(n5781) );
  AND U7156 ( .A(n5782), .B(n5783), .Z(n5780) );
  NAND U7157 ( .A(ereg[222]), .B(n4895), .Z(n5783) );
  NANDN U7158 ( .A(n4890), .B(ereg[223]), .Z(n5782) );
  NAND U7159 ( .A(n5784), .B(n5785), .Z(n3634) );
  NANDN U7160 ( .A(init), .B(e[224]), .Z(n5785) );
  AND U7161 ( .A(n5786), .B(n5787), .Z(n5784) );
  NAND U7162 ( .A(ereg[223]), .B(n4895), .Z(n5787) );
  NANDN U7163 ( .A(n4890), .B(ereg[224]), .Z(n5786) );
  NAND U7164 ( .A(n5788), .B(n5789), .Z(n3633) );
  NANDN U7165 ( .A(init), .B(e[225]), .Z(n5789) );
  AND U7166 ( .A(n5790), .B(n5791), .Z(n5788) );
  NAND U7167 ( .A(ereg[224]), .B(n4895), .Z(n5791) );
  NANDN U7168 ( .A(n4890), .B(ereg[225]), .Z(n5790) );
  NAND U7169 ( .A(n5792), .B(n5793), .Z(n3632) );
  NANDN U7170 ( .A(init), .B(e[226]), .Z(n5793) );
  AND U7171 ( .A(n5794), .B(n5795), .Z(n5792) );
  NAND U7172 ( .A(ereg[225]), .B(n4895), .Z(n5795) );
  NANDN U7173 ( .A(n4890), .B(ereg[226]), .Z(n5794) );
  NAND U7174 ( .A(n5796), .B(n5797), .Z(n3631) );
  NANDN U7175 ( .A(init), .B(e[227]), .Z(n5797) );
  AND U7176 ( .A(n5798), .B(n5799), .Z(n5796) );
  NAND U7177 ( .A(ereg[226]), .B(n4895), .Z(n5799) );
  NANDN U7178 ( .A(n4890), .B(ereg[227]), .Z(n5798) );
  NAND U7179 ( .A(n5800), .B(n5801), .Z(n3630) );
  NANDN U7180 ( .A(init), .B(e[228]), .Z(n5801) );
  AND U7181 ( .A(n5802), .B(n5803), .Z(n5800) );
  NAND U7182 ( .A(ereg[227]), .B(n4895), .Z(n5803) );
  NANDN U7183 ( .A(n4890), .B(ereg[228]), .Z(n5802) );
  NAND U7184 ( .A(n5804), .B(n5805), .Z(n3629) );
  NANDN U7185 ( .A(init), .B(e[229]), .Z(n5805) );
  AND U7186 ( .A(n5806), .B(n5807), .Z(n5804) );
  NAND U7187 ( .A(ereg[228]), .B(n4895), .Z(n5807) );
  NANDN U7188 ( .A(n4890), .B(ereg[229]), .Z(n5806) );
  NAND U7189 ( .A(n5808), .B(n5809), .Z(n3628) );
  NANDN U7190 ( .A(init), .B(e[230]), .Z(n5809) );
  AND U7191 ( .A(n5810), .B(n5811), .Z(n5808) );
  NAND U7192 ( .A(ereg[229]), .B(n4895), .Z(n5811) );
  NANDN U7193 ( .A(n4890), .B(ereg[230]), .Z(n5810) );
  NAND U7194 ( .A(n5812), .B(n5813), .Z(n3627) );
  NANDN U7195 ( .A(init), .B(e[231]), .Z(n5813) );
  AND U7196 ( .A(n5814), .B(n5815), .Z(n5812) );
  NAND U7197 ( .A(ereg[230]), .B(n4895), .Z(n5815) );
  NANDN U7198 ( .A(n4890), .B(ereg[231]), .Z(n5814) );
  NAND U7199 ( .A(n5816), .B(n5817), .Z(n3626) );
  NANDN U7200 ( .A(init), .B(e[232]), .Z(n5817) );
  AND U7201 ( .A(n5818), .B(n5819), .Z(n5816) );
  NAND U7202 ( .A(ereg[231]), .B(n4895), .Z(n5819) );
  NANDN U7203 ( .A(n4890), .B(ereg[232]), .Z(n5818) );
  NAND U7204 ( .A(n5820), .B(n5821), .Z(n3625) );
  NANDN U7205 ( .A(init), .B(e[233]), .Z(n5821) );
  AND U7206 ( .A(n5822), .B(n5823), .Z(n5820) );
  NAND U7207 ( .A(ereg[232]), .B(n4895), .Z(n5823) );
  NANDN U7208 ( .A(n4890), .B(ereg[233]), .Z(n5822) );
  NAND U7209 ( .A(n5824), .B(n5825), .Z(n3624) );
  NANDN U7210 ( .A(init), .B(e[234]), .Z(n5825) );
  AND U7211 ( .A(n5826), .B(n5827), .Z(n5824) );
  NAND U7212 ( .A(ereg[233]), .B(n4895), .Z(n5827) );
  NANDN U7213 ( .A(n4890), .B(ereg[234]), .Z(n5826) );
  NAND U7214 ( .A(n5828), .B(n5829), .Z(n3623) );
  NANDN U7215 ( .A(init), .B(e[235]), .Z(n5829) );
  AND U7216 ( .A(n5830), .B(n5831), .Z(n5828) );
  NAND U7217 ( .A(ereg[234]), .B(n4895), .Z(n5831) );
  NANDN U7218 ( .A(n4890), .B(ereg[235]), .Z(n5830) );
  NAND U7219 ( .A(n5832), .B(n5833), .Z(n3622) );
  NANDN U7220 ( .A(init), .B(e[236]), .Z(n5833) );
  AND U7221 ( .A(n5834), .B(n5835), .Z(n5832) );
  NAND U7222 ( .A(ereg[235]), .B(n4895), .Z(n5835) );
  NANDN U7223 ( .A(n4890), .B(ereg[236]), .Z(n5834) );
  NAND U7224 ( .A(n5836), .B(n5837), .Z(n3621) );
  NANDN U7225 ( .A(init), .B(e[237]), .Z(n5837) );
  AND U7226 ( .A(n5838), .B(n5839), .Z(n5836) );
  NAND U7227 ( .A(ereg[236]), .B(n4895), .Z(n5839) );
  NANDN U7228 ( .A(n4890), .B(ereg[237]), .Z(n5838) );
  NAND U7229 ( .A(n5840), .B(n5841), .Z(n3620) );
  NANDN U7230 ( .A(init), .B(e[238]), .Z(n5841) );
  AND U7231 ( .A(n5842), .B(n5843), .Z(n5840) );
  NAND U7232 ( .A(ereg[237]), .B(n4895), .Z(n5843) );
  NANDN U7233 ( .A(n4890), .B(ereg[238]), .Z(n5842) );
  NAND U7234 ( .A(n5844), .B(n5845), .Z(n3619) );
  NANDN U7235 ( .A(init), .B(e[239]), .Z(n5845) );
  AND U7236 ( .A(n5846), .B(n5847), .Z(n5844) );
  NAND U7237 ( .A(ereg[238]), .B(n4895), .Z(n5847) );
  NANDN U7238 ( .A(n4890), .B(ereg[239]), .Z(n5846) );
  NAND U7239 ( .A(n5848), .B(n5849), .Z(n3618) );
  NANDN U7240 ( .A(init), .B(e[240]), .Z(n5849) );
  AND U7241 ( .A(n5850), .B(n5851), .Z(n5848) );
  NAND U7242 ( .A(ereg[239]), .B(n4895), .Z(n5851) );
  NANDN U7243 ( .A(n4890), .B(ereg[240]), .Z(n5850) );
  NAND U7244 ( .A(n5852), .B(n5853), .Z(n3617) );
  NANDN U7245 ( .A(init), .B(e[241]), .Z(n5853) );
  AND U7246 ( .A(n5854), .B(n5855), .Z(n5852) );
  NAND U7247 ( .A(ereg[240]), .B(n4895), .Z(n5855) );
  NANDN U7248 ( .A(n4890), .B(ereg[241]), .Z(n5854) );
  NAND U7249 ( .A(n5856), .B(n5857), .Z(n3616) );
  NANDN U7250 ( .A(init), .B(e[242]), .Z(n5857) );
  AND U7251 ( .A(n5858), .B(n5859), .Z(n5856) );
  NAND U7252 ( .A(ereg[241]), .B(n4895), .Z(n5859) );
  NANDN U7253 ( .A(n4890), .B(ereg[242]), .Z(n5858) );
  NAND U7254 ( .A(n5860), .B(n5861), .Z(n3615) );
  NANDN U7255 ( .A(init), .B(e[243]), .Z(n5861) );
  AND U7256 ( .A(n5862), .B(n5863), .Z(n5860) );
  NAND U7257 ( .A(ereg[242]), .B(n4895), .Z(n5863) );
  NANDN U7258 ( .A(n4890), .B(ereg[243]), .Z(n5862) );
  NAND U7259 ( .A(n5864), .B(n5865), .Z(n3614) );
  NANDN U7260 ( .A(init), .B(e[244]), .Z(n5865) );
  AND U7261 ( .A(n5866), .B(n5867), .Z(n5864) );
  NAND U7262 ( .A(ereg[243]), .B(n4895), .Z(n5867) );
  NANDN U7263 ( .A(n4890), .B(ereg[244]), .Z(n5866) );
  NAND U7264 ( .A(n5868), .B(n5869), .Z(n3613) );
  NANDN U7265 ( .A(init), .B(e[245]), .Z(n5869) );
  AND U7266 ( .A(n5870), .B(n5871), .Z(n5868) );
  NAND U7267 ( .A(ereg[244]), .B(n4895), .Z(n5871) );
  NANDN U7268 ( .A(n4890), .B(ereg[245]), .Z(n5870) );
  NAND U7269 ( .A(n5872), .B(n5873), .Z(n3612) );
  NANDN U7270 ( .A(init), .B(e[246]), .Z(n5873) );
  AND U7271 ( .A(n5874), .B(n5875), .Z(n5872) );
  NAND U7272 ( .A(ereg[245]), .B(n4895), .Z(n5875) );
  NANDN U7273 ( .A(n4890), .B(ereg[246]), .Z(n5874) );
  NAND U7274 ( .A(n5876), .B(n5877), .Z(n3611) );
  NANDN U7275 ( .A(init), .B(e[247]), .Z(n5877) );
  AND U7276 ( .A(n5878), .B(n5879), .Z(n5876) );
  NAND U7277 ( .A(ereg[246]), .B(n4895), .Z(n5879) );
  NANDN U7278 ( .A(n4890), .B(ereg[247]), .Z(n5878) );
  NAND U7279 ( .A(n5880), .B(n5881), .Z(n3610) );
  NANDN U7280 ( .A(init), .B(e[248]), .Z(n5881) );
  AND U7281 ( .A(n5882), .B(n5883), .Z(n5880) );
  NAND U7282 ( .A(ereg[247]), .B(n4895), .Z(n5883) );
  NANDN U7283 ( .A(n4890), .B(ereg[248]), .Z(n5882) );
  NAND U7284 ( .A(n5884), .B(n5885), .Z(n3609) );
  NANDN U7285 ( .A(init), .B(e[249]), .Z(n5885) );
  AND U7286 ( .A(n5886), .B(n5887), .Z(n5884) );
  NAND U7287 ( .A(ereg[248]), .B(n4895), .Z(n5887) );
  NANDN U7288 ( .A(n4890), .B(ereg[249]), .Z(n5886) );
  NAND U7289 ( .A(n5888), .B(n5889), .Z(n3608) );
  NANDN U7290 ( .A(init), .B(e[250]), .Z(n5889) );
  AND U7291 ( .A(n5890), .B(n5891), .Z(n5888) );
  NAND U7292 ( .A(ereg[249]), .B(n4895), .Z(n5891) );
  NANDN U7293 ( .A(n4890), .B(ereg[250]), .Z(n5890) );
  NAND U7294 ( .A(n5892), .B(n5893), .Z(n3607) );
  NANDN U7295 ( .A(init), .B(e[251]), .Z(n5893) );
  AND U7296 ( .A(n5894), .B(n5895), .Z(n5892) );
  NAND U7297 ( .A(ereg[250]), .B(n4895), .Z(n5895) );
  NANDN U7298 ( .A(n4890), .B(ereg[251]), .Z(n5894) );
  NAND U7299 ( .A(n5896), .B(n5897), .Z(n3606) );
  NANDN U7300 ( .A(init), .B(e[252]), .Z(n5897) );
  AND U7301 ( .A(n5898), .B(n5899), .Z(n5896) );
  NAND U7302 ( .A(ereg[251]), .B(n4895), .Z(n5899) );
  NANDN U7303 ( .A(n4890), .B(ereg[252]), .Z(n5898) );
  NAND U7304 ( .A(n5900), .B(n5901), .Z(n3605) );
  NANDN U7305 ( .A(init), .B(e[253]), .Z(n5901) );
  AND U7306 ( .A(n5902), .B(n5903), .Z(n5900) );
  NAND U7307 ( .A(ereg[252]), .B(n4895), .Z(n5903) );
  NANDN U7308 ( .A(n4890), .B(ereg[253]), .Z(n5902) );
  NAND U7309 ( .A(n5904), .B(n5905), .Z(n3604) );
  NANDN U7310 ( .A(init), .B(e[254]), .Z(n5905) );
  AND U7311 ( .A(n5906), .B(n5907), .Z(n5904) );
  NAND U7312 ( .A(ereg[253]), .B(n4895), .Z(n5907) );
  NANDN U7313 ( .A(n4890), .B(ereg[254]), .Z(n5906) );
  NAND U7314 ( .A(n5908), .B(n5909), .Z(n3603) );
  NANDN U7315 ( .A(init), .B(e[255]), .Z(n5909) );
  AND U7316 ( .A(n5910), .B(n5911), .Z(n5908) );
  NAND U7317 ( .A(ereg[254]), .B(n4895), .Z(n5911) );
  AND U7318 ( .A(n4890), .B(n7204), .Z(n4895) );
  NANDN U7319 ( .A(n4890), .B(ereg[255]), .Z(n5910) );
  AND U7320 ( .A(n5912), .B(n3862), .Z(n4890) );
  NANDN U7321 ( .A(mul_pow), .B(init), .Z(n3862) );
  NANDN U7322 ( .A(start_reg[63]), .B(init), .Z(n5912) );
  NAND U7323 ( .A(n5913), .B(n4541), .Z(n3602) );
  NANDN U7324 ( .A(init), .B(m[255]), .Z(n4541) );
  AND U7325 ( .A(n5914), .B(n5915), .Z(n5913) );
  NAND U7326 ( .A(o[255]), .B(n5916), .Z(n5915) );
  NANDN U7327 ( .A(n5917), .B(creg[255]), .Z(n5914) );
  NAND U7328 ( .A(n5918), .B(n4885), .Z(n3601) );
  NANDN U7329 ( .A(init), .B(m[0]), .Z(n4885) );
  AND U7330 ( .A(n5919), .B(n5920), .Z(n5918) );
  NAND U7331 ( .A(o[0]), .B(n5916), .Z(n5920) );
  NANDN U7332 ( .A(n5917), .B(creg[0]), .Z(n5919) );
  NAND U7333 ( .A(n5921), .B(n4663), .Z(n3600) );
  NANDN U7334 ( .A(init), .B(m[1]), .Z(n4663) );
  AND U7335 ( .A(n5922), .B(n5923), .Z(n5921) );
  NAND U7336 ( .A(o[1]), .B(n5916), .Z(n5923) );
  NANDN U7337 ( .A(n5917), .B(creg[1]), .Z(n5922) );
  NAND U7338 ( .A(n5924), .B(n4529), .Z(n3599) );
  NANDN U7339 ( .A(init), .B(m[2]), .Z(n4529) );
  AND U7340 ( .A(n5925), .B(n5926), .Z(n5924) );
  NAND U7341 ( .A(o[2]), .B(n5916), .Z(n5926) );
  NANDN U7342 ( .A(n5917), .B(creg[2]), .Z(n5925) );
  NAND U7343 ( .A(n5927), .B(n4507), .Z(n3598) );
  NANDN U7344 ( .A(init), .B(m[3]), .Z(n4507) );
  AND U7345 ( .A(n5928), .B(n5929), .Z(n5927) );
  NAND U7346 ( .A(o[3]), .B(n5916), .Z(n5929) );
  NANDN U7347 ( .A(n5917), .B(creg[3]), .Z(n5928) );
  NAND U7348 ( .A(n5930), .B(n4485), .Z(n3597) );
  NANDN U7349 ( .A(init), .B(m[4]), .Z(n4485) );
  AND U7350 ( .A(n5931), .B(n5932), .Z(n5930) );
  NAND U7351 ( .A(o[4]), .B(n5916), .Z(n5932) );
  NANDN U7352 ( .A(n5917), .B(creg[4]), .Z(n5931) );
  NAND U7353 ( .A(n5933), .B(n4463), .Z(n3596) );
  NANDN U7354 ( .A(init), .B(m[5]), .Z(n4463) );
  AND U7355 ( .A(n5934), .B(n5935), .Z(n5933) );
  NAND U7356 ( .A(o[5]), .B(n5916), .Z(n5935) );
  NANDN U7357 ( .A(n5917), .B(creg[5]), .Z(n5934) );
  NAND U7358 ( .A(n5936), .B(n4441), .Z(n3595) );
  NANDN U7359 ( .A(init), .B(m[6]), .Z(n4441) );
  AND U7360 ( .A(n5937), .B(n5938), .Z(n5936) );
  NAND U7361 ( .A(o[6]), .B(n5916), .Z(n5938) );
  NANDN U7362 ( .A(n5917), .B(creg[6]), .Z(n5937) );
  NAND U7363 ( .A(n5939), .B(n4419), .Z(n3594) );
  NANDN U7364 ( .A(init), .B(m[7]), .Z(n4419) );
  AND U7365 ( .A(n5940), .B(n5941), .Z(n5939) );
  NAND U7366 ( .A(o[7]), .B(n5916), .Z(n5941) );
  NANDN U7367 ( .A(n5917), .B(creg[7]), .Z(n5940) );
  NAND U7368 ( .A(n5942), .B(n4397), .Z(n3593) );
  NANDN U7369 ( .A(init), .B(m[8]), .Z(n4397) );
  AND U7370 ( .A(n5943), .B(n5944), .Z(n5942) );
  NAND U7371 ( .A(o[8]), .B(n5916), .Z(n5944) );
  NANDN U7372 ( .A(n5917), .B(creg[8]), .Z(n5943) );
  NAND U7373 ( .A(n5945), .B(n4375), .Z(n3592) );
  NANDN U7374 ( .A(init), .B(m[9]), .Z(n4375) );
  AND U7375 ( .A(n5946), .B(n5947), .Z(n5945) );
  NAND U7376 ( .A(o[9]), .B(n5916), .Z(n5947) );
  NANDN U7377 ( .A(n5917), .B(creg[9]), .Z(n5946) );
  NAND U7378 ( .A(n5948), .B(n4863), .Z(n3591) );
  NANDN U7379 ( .A(init), .B(m[10]), .Z(n4863) );
  AND U7380 ( .A(n5949), .B(n5950), .Z(n5948) );
  NAND U7381 ( .A(o[10]), .B(n5916), .Z(n5950) );
  NANDN U7382 ( .A(n5917), .B(creg[10]), .Z(n5949) );
  NAND U7383 ( .A(n5951), .B(n4841), .Z(n3590) );
  NANDN U7384 ( .A(init), .B(m[11]), .Z(n4841) );
  AND U7385 ( .A(n5952), .B(n5953), .Z(n5951) );
  NAND U7386 ( .A(o[11]), .B(n5916), .Z(n5953) );
  NANDN U7387 ( .A(n5917), .B(creg[11]), .Z(n5952) );
  NAND U7388 ( .A(n5954), .B(n4819), .Z(n3589) );
  NANDN U7389 ( .A(init), .B(m[12]), .Z(n4819) );
  AND U7390 ( .A(n5955), .B(n5956), .Z(n5954) );
  NAND U7391 ( .A(o[12]), .B(n5916), .Z(n5956) );
  NANDN U7392 ( .A(n5917), .B(creg[12]), .Z(n5955) );
  NAND U7393 ( .A(n5957), .B(n4797), .Z(n3588) );
  NANDN U7394 ( .A(init), .B(m[13]), .Z(n4797) );
  AND U7395 ( .A(n5958), .B(n5959), .Z(n5957) );
  NAND U7396 ( .A(o[13]), .B(n5916), .Z(n5959) );
  NANDN U7397 ( .A(n5917), .B(creg[13]), .Z(n5958) );
  NAND U7398 ( .A(n5960), .B(n4775), .Z(n3587) );
  NANDN U7399 ( .A(init), .B(m[14]), .Z(n4775) );
  AND U7400 ( .A(n5961), .B(n5962), .Z(n5960) );
  NAND U7401 ( .A(o[14]), .B(n5916), .Z(n5962) );
  NANDN U7402 ( .A(n5917), .B(creg[14]), .Z(n5961) );
  NAND U7403 ( .A(n5963), .B(n4753), .Z(n3586) );
  NANDN U7404 ( .A(init), .B(m[15]), .Z(n4753) );
  AND U7405 ( .A(n5964), .B(n5965), .Z(n5963) );
  NAND U7406 ( .A(o[15]), .B(n5916), .Z(n5965) );
  NANDN U7407 ( .A(n5917), .B(creg[15]), .Z(n5964) );
  NAND U7408 ( .A(n5966), .B(n4731), .Z(n3585) );
  NANDN U7409 ( .A(init), .B(m[16]), .Z(n4731) );
  AND U7410 ( .A(n5967), .B(n5968), .Z(n5966) );
  NAND U7411 ( .A(o[16]), .B(n5916), .Z(n5968) );
  NANDN U7412 ( .A(n5917), .B(creg[16]), .Z(n5967) );
  NAND U7413 ( .A(n5969), .B(n4709), .Z(n3584) );
  NANDN U7414 ( .A(init), .B(m[17]), .Z(n4709) );
  AND U7415 ( .A(n5970), .B(n5971), .Z(n5969) );
  NAND U7416 ( .A(o[17]), .B(n5916), .Z(n5971) );
  NANDN U7417 ( .A(n5917), .B(creg[17]), .Z(n5970) );
  NAND U7418 ( .A(n5972), .B(n4687), .Z(n3583) );
  NANDN U7419 ( .A(init), .B(m[18]), .Z(n4687) );
  AND U7420 ( .A(n5973), .B(n5974), .Z(n5972) );
  NAND U7421 ( .A(o[18]), .B(n5916), .Z(n5974) );
  NANDN U7422 ( .A(n5917), .B(creg[18]), .Z(n5973) );
  NAND U7423 ( .A(n5975), .B(n4665), .Z(n3582) );
  NANDN U7424 ( .A(init), .B(m[19]), .Z(n4665) );
  AND U7425 ( .A(n5976), .B(n5977), .Z(n5975) );
  NAND U7426 ( .A(o[19]), .B(n5916), .Z(n5977) );
  NANDN U7427 ( .A(n5917), .B(creg[19]), .Z(n5976) );
  NAND U7428 ( .A(n5978), .B(n4641), .Z(n3581) );
  NANDN U7429 ( .A(init), .B(m[20]), .Z(n4641) );
  AND U7430 ( .A(n5979), .B(n5980), .Z(n5978) );
  NAND U7431 ( .A(o[20]), .B(n5916), .Z(n5980) );
  NANDN U7432 ( .A(n5917), .B(creg[20]), .Z(n5979) );
  NAND U7433 ( .A(n5981), .B(n4619), .Z(n3580) );
  NANDN U7434 ( .A(init), .B(m[21]), .Z(n4619) );
  AND U7435 ( .A(n5982), .B(n5983), .Z(n5981) );
  NAND U7436 ( .A(o[21]), .B(n5916), .Z(n5983) );
  NANDN U7437 ( .A(n5917), .B(creg[21]), .Z(n5982) );
  NAND U7438 ( .A(n5984), .B(n4597), .Z(n3579) );
  NANDN U7439 ( .A(init), .B(m[22]), .Z(n4597) );
  AND U7440 ( .A(n5985), .B(n5986), .Z(n5984) );
  NAND U7441 ( .A(o[22]), .B(n5916), .Z(n5986) );
  NANDN U7442 ( .A(n5917), .B(creg[22]), .Z(n5985) );
  NAND U7443 ( .A(n5987), .B(n4575), .Z(n3578) );
  NANDN U7444 ( .A(init), .B(m[23]), .Z(n4575) );
  AND U7445 ( .A(n5988), .B(n5989), .Z(n5987) );
  NAND U7446 ( .A(o[23]), .B(n5916), .Z(n5989) );
  NANDN U7447 ( .A(n5917), .B(creg[23]), .Z(n5988) );
  NAND U7448 ( .A(n5990), .B(n4553), .Z(n3577) );
  NANDN U7449 ( .A(init), .B(m[24]), .Z(n4553) );
  AND U7450 ( .A(n5991), .B(n5992), .Z(n5990) );
  NAND U7451 ( .A(o[24]), .B(n5916), .Z(n5992) );
  NANDN U7452 ( .A(n5917), .B(creg[24]), .Z(n5991) );
  NAND U7453 ( .A(n5993), .B(n4539), .Z(n3576) );
  NANDN U7454 ( .A(init), .B(m[25]), .Z(n4539) );
  AND U7455 ( .A(n5994), .B(n5995), .Z(n5993) );
  NAND U7456 ( .A(o[25]), .B(n5916), .Z(n5995) );
  NANDN U7457 ( .A(n5917), .B(creg[25]), .Z(n5994) );
  NAND U7458 ( .A(n5996), .B(n4537), .Z(n3575) );
  NANDN U7459 ( .A(init), .B(m[26]), .Z(n4537) );
  AND U7460 ( .A(n5997), .B(n5998), .Z(n5996) );
  NAND U7461 ( .A(o[26]), .B(n5916), .Z(n5998) );
  NANDN U7462 ( .A(n5917), .B(creg[26]), .Z(n5997) );
  NAND U7463 ( .A(n5999), .B(n4535), .Z(n3574) );
  NANDN U7464 ( .A(init), .B(m[27]), .Z(n4535) );
  AND U7465 ( .A(n6000), .B(n6001), .Z(n5999) );
  NAND U7466 ( .A(o[27]), .B(n5916), .Z(n6001) );
  NANDN U7467 ( .A(n5917), .B(creg[27]), .Z(n6000) );
  NAND U7468 ( .A(n6002), .B(n4533), .Z(n3573) );
  NANDN U7469 ( .A(init), .B(m[28]), .Z(n4533) );
  AND U7470 ( .A(n6003), .B(n6004), .Z(n6002) );
  NAND U7471 ( .A(o[28]), .B(n5916), .Z(n6004) );
  NANDN U7472 ( .A(n5917), .B(creg[28]), .Z(n6003) );
  NAND U7473 ( .A(n6005), .B(n4531), .Z(n3572) );
  NANDN U7474 ( .A(init), .B(m[29]), .Z(n4531) );
  AND U7475 ( .A(n6006), .B(n6007), .Z(n6005) );
  NAND U7476 ( .A(o[29]), .B(n5916), .Z(n6007) );
  NANDN U7477 ( .A(n5917), .B(creg[29]), .Z(n6006) );
  NAND U7478 ( .A(n6008), .B(n4527), .Z(n3571) );
  NANDN U7479 ( .A(init), .B(m[30]), .Z(n4527) );
  AND U7480 ( .A(n6009), .B(n6010), .Z(n6008) );
  NAND U7481 ( .A(o[30]), .B(n5916), .Z(n6010) );
  NANDN U7482 ( .A(n5917), .B(creg[30]), .Z(n6009) );
  NAND U7483 ( .A(n6011), .B(n4525), .Z(n3570) );
  NANDN U7484 ( .A(init), .B(m[31]), .Z(n4525) );
  AND U7485 ( .A(n6012), .B(n6013), .Z(n6011) );
  NAND U7486 ( .A(o[31]), .B(n5916), .Z(n6013) );
  NANDN U7487 ( .A(n5917), .B(creg[31]), .Z(n6012) );
  NAND U7488 ( .A(n6014), .B(n4523), .Z(n3569) );
  NANDN U7489 ( .A(init), .B(m[32]), .Z(n4523) );
  AND U7490 ( .A(n6015), .B(n6016), .Z(n6014) );
  NAND U7491 ( .A(o[32]), .B(n5916), .Z(n6016) );
  NANDN U7492 ( .A(n5917), .B(creg[32]), .Z(n6015) );
  NAND U7493 ( .A(n6017), .B(n4521), .Z(n3568) );
  NANDN U7494 ( .A(init), .B(m[33]), .Z(n4521) );
  AND U7495 ( .A(n6018), .B(n6019), .Z(n6017) );
  NAND U7496 ( .A(o[33]), .B(n5916), .Z(n6019) );
  NANDN U7497 ( .A(n5917), .B(creg[33]), .Z(n6018) );
  NAND U7498 ( .A(n6020), .B(n4519), .Z(n3567) );
  NANDN U7499 ( .A(init), .B(m[34]), .Z(n4519) );
  AND U7500 ( .A(n6021), .B(n6022), .Z(n6020) );
  NAND U7501 ( .A(o[34]), .B(n5916), .Z(n6022) );
  NANDN U7502 ( .A(n5917), .B(creg[34]), .Z(n6021) );
  NAND U7503 ( .A(n6023), .B(n4517), .Z(n3566) );
  NANDN U7504 ( .A(init), .B(m[35]), .Z(n4517) );
  AND U7505 ( .A(n6024), .B(n6025), .Z(n6023) );
  NAND U7506 ( .A(o[35]), .B(n5916), .Z(n6025) );
  NANDN U7507 ( .A(n5917), .B(creg[35]), .Z(n6024) );
  NAND U7508 ( .A(n6026), .B(n4515), .Z(n3565) );
  NANDN U7509 ( .A(init), .B(m[36]), .Z(n4515) );
  AND U7510 ( .A(n6027), .B(n6028), .Z(n6026) );
  NAND U7511 ( .A(o[36]), .B(n5916), .Z(n6028) );
  NANDN U7512 ( .A(n5917), .B(creg[36]), .Z(n6027) );
  NAND U7513 ( .A(n6029), .B(n4513), .Z(n3564) );
  NANDN U7514 ( .A(init), .B(m[37]), .Z(n4513) );
  AND U7515 ( .A(n6030), .B(n6031), .Z(n6029) );
  NAND U7516 ( .A(o[37]), .B(n5916), .Z(n6031) );
  NANDN U7517 ( .A(n5917), .B(creg[37]), .Z(n6030) );
  NAND U7518 ( .A(n6032), .B(n4511), .Z(n3563) );
  NANDN U7519 ( .A(init), .B(m[38]), .Z(n4511) );
  AND U7520 ( .A(n6033), .B(n6034), .Z(n6032) );
  NAND U7521 ( .A(o[38]), .B(n5916), .Z(n6034) );
  NANDN U7522 ( .A(n5917), .B(creg[38]), .Z(n6033) );
  NAND U7523 ( .A(n6035), .B(n4509), .Z(n3562) );
  NANDN U7524 ( .A(init), .B(m[39]), .Z(n4509) );
  AND U7525 ( .A(n6036), .B(n6037), .Z(n6035) );
  NAND U7526 ( .A(o[39]), .B(n5916), .Z(n6037) );
  NANDN U7527 ( .A(n5917), .B(creg[39]), .Z(n6036) );
  NAND U7528 ( .A(n6038), .B(n4505), .Z(n3561) );
  NANDN U7529 ( .A(init), .B(m[40]), .Z(n4505) );
  AND U7530 ( .A(n6039), .B(n6040), .Z(n6038) );
  NAND U7531 ( .A(o[40]), .B(n5916), .Z(n6040) );
  NANDN U7532 ( .A(n5917), .B(creg[40]), .Z(n6039) );
  NAND U7533 ( .A(n6041), .B(n4503), .Z(n3560) );
  NANDN U7534 ( .A(init), .B(m[41]), .Z(n4503) );
  AND U7535 ( .A(n6042), .B(n6043), .Z(n6041) );
  NAND U7536 ( .A(o[41]), .B(n5916), .Z(n6043) );
  NANDN U7537 ( .A(n5917), .B(creg[41]), .Z(n6042) );
  NAND U7538 ( .A(n6044), .B(n4501), .Z(n3559) );
  NANDN U7539 ( .A(init), .B(m[42]), .Z(n4501) );
  AND U7540 ( .A(n6045), .B(n6046), .Z(n6044) );
  NAND U7541 ( .A(o[42]), .B(n5916), .Z(n6046) );
  NANDN U7542 ( .A(n5917), .B(creg[42]), .Z(n6045) );
  NAND U7543 ( .A(n6047), .B(n4499), .Z(n3558) );
  NANDN U7544 ( .A(init), .B(m[43]), .Z(n4499) );
  AND U7545 ( .A(n6048), .B(n6049), .Z(n6047) );
  NAND U7546 ( .A(o[43]), .B(n5916), .Z(n6049) );
  NANDN U7547 ( .A(n5917), .B(creg[43]), .Z(n6048) );
  NAND U7548 ( .A(n6050), .B(n4497), .Z(n3557) );
  NANDN U7549 ( .A(init), .B(m[44]), .Z(n4497) );
  AND U7550 ( .A(n6051), .B(n6052), .Z(n6050) );
  NAND U7551 ( .A(o[44]), .B(n5916), .Z(n6052) );
  NANDN U7552 ( .A(n5917), .B(creg[44]), .Z(n6051) );
  NAND U7553 ( .A(n6053), .B(n4495), .Z(n3556) );
  NANDN U7554 ( .A(init), .B(m[45]), .Z(n4495) );
  AND U7555 ( .A(n6054), .B(n6055), .Z(n6053) );
  NAND U7556 ( .A(o[45]), .B(n5916), .Z(n6055) );
  NANDN U7557 ( .A(n5917), .B(creg[45]), .Z(n6054) );
  NAND U7558 ( .A(n6056), .B(n4493), .Z(n3555) );
  NANDN U7559 ( .A(init), .B(m[46]), .Z(n4493) );
  AND U7560 ( .A(n6057), .B(n6058), .Z(n6056) );
  NAND U7561 ( .A(o[46]), .B(n5916), .Z(n6058) );
  NANDN U7562 ( .A(n5917), .B(creg[46]), .Z(n6057) );
  NAND U7563 ( .A(n6059), .B(n4491), .Z(n3554) );
  NANDN U7564 ( .A(init), .B(m[47]), .Z(n4491) );
  AND U7565 ( .A(n6060), .B(n6061), .Z(n6059) );
  NAND U7566 ( .A(o[47]), .B(n5916), .Z(n6061) );
  NANDN U7567 ( .A(n5917), .B(creg[47]), .Z(n6060) );
  NAND U7568 ( .A(n6062), .B(n4489), .Z(n3553) );
  NANDN U7569 ( .A(init), .B(m[48]), .Z(n4489) );
  AND U7570 ( .A(n6063), .B(n6064), .Z(n6062) );
  NAND U7571 ( .A(o[48]), .B(n5916), .Z(n6064) );
  NANDN U7572 ( .A(n5917), .B(creg[48]), .Z(n6063) );
  NAND U7573 ( .A(n6065), .B(n4487), .Z(n3552) );
  NANDN U7574 ( .A(init), .B(m[49]), .Z(n4487) );
  AND U7575 ( .A(n6066), .B(n6067), .Z(n6065) );
  NAND U7576 ( .A(o[49]), .B(n5916), .Z(n6067) );
  NANDN U7577 ( .A(n5917), .B(creg[49]), .Z(n6066) );
  NAND U7578 ( .A(n6068), .B(n4483), .Z(n3551) );
  NANDN U7579 ( .A(init), .B(m[50]), .Z(n4483) );
  AND U7580 ( .A(n6069), .B(n6070), .Z(n6068) );
  NAND U7581 ( .A(o[50]), .B(n5916), .Z(n6070) );
  NANDN U7582 ( .A(n5917), .B(creg[50]), .Z(n6069) );
  NAND U7583 ( .A(n6071), .B(n4481), .Z(n3550) );
  NANDN U7584 ( .A(init), .B(m[51]), .Z(n4481) );
  AND U7585 ( .A(n6072), .B(n6073), .Z(n6071) );
  NAND U7586 ( .A(o[51]), .B(n5916), .Z(n6073) );
  NANDN U7587 ( .A(n5917), .B(creg[51]), .Z(n6072) );
  NAND U7588 ( .A(n6074), .B(n4479), .Z(n3549) );
  NANDN U7589 ( .A(init), .B(m[52]), .Z(n4479) );
  AND U7590 ( .A(n6075), .B(n6076), .Z(n6074) );
  NAND U7591 ( .A(o[52]), .B(n5916), .Z(n6076) );
  NANDN U7592 ( .A(n5917), .B(creg[52]), .Z(n6075) );
  NAND U7593 ( .A(n6077), .B(n4477), .Z(n3548) );
  NANDN U7594 ( .A(init), .B(m[53]), .Z(n4477) );
  AND U7595 ( .A(n6078), .B(n6079), .Z(n6077) );
  NAND U7596 ( .A(o[53]), .B(n5916), .Z(n6079) );
  NANDN U7597 ( .A(n5917), .B(creg[53]), .Z(n6078) );
  NAND U7598 ( .A(n6080), .B(n4475), .Z(n3547) );
  NANDN U7599 ( .A(init), .B(m[54]), .Z(n4475) );
  AND U7600 ( .A(n6081), .B(n6082), .Z(n6080) );
  NAND U7601 ( .A(o[54]), .B(n5916), .Z(n6082) );
  NANDN U7602 ( .A(n5917), .B(creg[54]), .Z(n6081) );
  NAND U7603 ( .A(n6083), .B(n4473), .Z(n3546) );
  NANDN U7604 ( .A(init), .B(m[55]), .Z(n4473) );
  AND U7605 ( .A(n6084), .B(n6085), .Z(n6083) );
  NAND U7606 ( .A(o[55]), .B(n5916), .Z(n6085) );
  NANDN U7607 ( .A(n5917), .B(creg[55]), .Z(n6084) );
  NAND U7608 ( .A(n6086), .B(n4471), .Z(n3545) );
  NANDN U7609 ( .A(init), .B(m[56]), .Z(n4471) );
  AND U7610 ( .A(n6087), .B(n6088), .Z(n6086) );
  NAND U7611 ( .A(o[56]), .B(n5916), .Z(n6088) );
  NANDN U7612 ( .A(n5917), .B(creg[56]), .Z(n6087) );
  NAND U7613 ( .A(n6089), .B(n4469), .Z(n3544) );
  NANDN U7614 ( .A(init), .B(m[57]), .Z(n4469) );
  AND U7615 ( .A(n6090), .B(n6091), .Z(n6089) );
  NAND U7616 ( .A(o[57]), .B(n5916), .Z(n6091) );
  NANDN U7617 ( .A(n5917), .B(creg[57]), .Z(n6090) );
  NAND U7618 ( .A(n6092), .B(n4467), .Z(n3543) );
  NANDN U7619 ( .A(init), .B(m[58]), .Z(n4467) );
  AND U7620 ( .A(n6093), .B(n6094), .Z(n6092) );
  NAND U7621 ( .A(o[58]), .B(n5916), .Z(n6094) );
  NANDN U7622 ( .A(n5917), .B(creg[58]), .Z(n6093) );
  NAND U7623 ( .A(n6095), .B(n4465), .Z(n3542) );
  NANDN U7624 ( .A(init), .B(m[59]), .Z(n4465) );
  AND U7625 ( .A(n6096), .B(n6097), .Z(n6095) );
  NAND U7626 ( .A(o[59]), .B(n5916), .Z(n6097) );
  NANDN U7627 ( .A(n5917), .B(creg[59]), .Z(n6096) );
  NAND U7628 ( .A(n6098), .B(n4461), .Z(n3541) );
  NANDN U7629 ( .A(init), .B(m[60]), .Z(n4461) );
  AND U7630 ( .A(n6099), .B(n6100), .Z(n6098) );
  NAND U7631 ( .A(o[60]), .B(n5916), .Z(n6100) );
  NANDN U7632 ( .A(n5917), .B(creg[60]), .Z(n6099) );
  NAND U7633 ( .A(n6101), .B(n4459), .Z(n3540) );
  NANDN U7634 ( .A(init), .B(m[61]), .Z(n4459) );
  AND U7635 ( .A(n6102), .B(n6103), .Z(n6101) );
  NAND U7636 ( .A(o[61]), .B(n5916), .Z(n6103) );
  NANDN U7637 ( .A(n5917), .B(creg[61]), .Z(n6102) );
  NAND U7638 ( .A(n6104), .B(n4457), .Z(n3539) );
  NANDN U7639 ( .A(init), .B(m[62]), .Z(n4457) );
  AND U7640 ( .A(n6105), .B(n6106), .Z(n6104) );
  NAND U7641 ( .A(o[62]), .B(n5916), .Z(n6106) );
  NANDN U7642 ( .A(n5917), .B(creg[62]), .Z(n6105) );
  NAND U7643 ( .A(n6107), .B(n4455), .Z(n3538) );
  NANDN U7644 ( .A(init), .B(m[63]), .Z(n4455) );
  AND U7645 ( .A(n6108), .B(n6109), .Z(n6107) );
  NAND U7646 ( .A(o[63]), .B(n5916), .Z(n6109) );
  NANDN U7647 ( .A(n5917), .B(creg[63]), .Z(n6108) );
  NAND U7648 ( .A(n6110), .B(n4453), .Z(n3537) );
  NANDN U7649 ( .A(init), .B(m[64]), .Z(n4453) );
  AND U7650 ( .A(n6111), .B(n6112), .Z(n6110) );
  NAND U7651 ( .A(o[64]), .B(n5916), .Z(n6112) );
  NANDN U7652 ( .A(n5917), .B(creg[64]), .Z(n6111) );
  NAND U7653 ( .A(n6113), .B(n4451), .Z(n3536) );
  NANDN U7654 ( .A(init), .B(m[65]), .Z(n4451) );
  AND U7655 ( .A(n6114), .B(n6115), .Z(n6113) );
  NAND U7656 ( .A(o[65]), .B(n5916), .Z(n6115) );
  NANDN U7657 ( .A(n5917), .B(creg[65]), .Z(n6114) );
  NAND U7658 ( .A(n6116), .B(n4449), .Z(n3535) );
  NANDN U7659 ( .A(init), .B(m[66]), .Z(n4449) );
  AND U7660 ( .A(n6117), .B(n6118), .Z(n6116) );
  NAND U7661 ( .A(o[66]), .B(n5916), .Z(n6118) );
  NANDN U7662 ( .A(n5917), .B(creg[66]), .Z(n6117) );
  NAND U7663 ( .A(n6119), .B(n4447), .Z(n3534) );
  NANDN U7664 ( .A(init), .B(m[67]), .Z(n4447) );
  AND U7665 ( .A(n6120), .B(n6121), .Z(n6119) );
  NAND U7666 ( .A(o[67]), .B(n5916), .Z(n6121) );
  NANDN U7667 ( .A(n5917), .B(creg[67]), .Z(n6120) );
  NAND U7668 ( .A(n6122), .B(n4445), .Z(n3533) );
  NANDN U7669 ( .A(init), .B(m[68]), .Z(n4445) );
  AND U7670 ( .A(n6123), .B(n6124), .Z(n6122) );
  NAND U7671 ( .A(o[68]), .B(n5916), .Z(n6124) );
  NANDN U7672 ( .A(n5917), .B(creg[68]), .Z(n6123) );
  NAND U7673 ( .A(n6125), .B(n4443), .Z(n3532) );
  NANDN U7674 ( .A(init), .B(m[69]), .Z(n4443) );
  AND U7675 ( .A(n6126), .B(n6127), .Z(n6125) );
  NAND U7676 ( .A(o[69]), .B(n5916), .Z(n6127) );
  NANDN U7677 ( .A(n5917), .B(creg[69]), .Z(n6126) );
  NAND U7678 ( .A(n6128), .B(n4439), .Z(n3531) );
  NANDN U7679 ( .A(init), .B(m[70]), .Z(n4439) );
  AND U7680 ( .A(n6129), .B(n6130), .Z(n6128) );
  NAND U7681 ( .A(o[70]), .B(n5916), .Z(n6130) );
  NANDN U7682 ( .A(n5917), .B(creg[70]), .Z(n6129) );
  NAND U7683 ( .A(n6131), .B(n4437), .Z(n3530) );
  NANDN U7684 ( .A(init), .B(m[71]), .Z(n4437) );
  AND U7685 ( .A(n6132), .B(n6133), .Z(n6131) );
  NAND U7686 ( .A(o[71]), .B(n5916), .Z(n6133) );
  NANDN U7687 ( .A(n5917), .B(creg[71]), .Z(n6132) );
  NAND U7688 ( .A(n6134), .B(n4435), .Z(n3529) );
  NANDN U7689 ( .A(init), .B(m[72]), .Z(n4435) );
  AND U7690 ( .A(n6135), .B(n6136), .Z(n6134) );
  NAND U7691 ( .A(o[72]), .B(n5916), .Z(n6136) );
  NANDN U7692 ( .A(n5917), .B(creg[72]), .Z(n6135) );
  NAND U7693 ( .A(n6137), .B(n4433), .Z(n3528) );
  NANDN U7694 ( .A(init), .B(m[73]), .Z(n4433) );
  AND U7695 ( .A(n6138), .B(n6139), .Z(n6137) );
  NAND U7696 ( .A(o[73]), .B(n5916), .Z(n6139) );
  NANDN U7697 ( .A(n5917), .B(creg[73]), .Z(n6138) );
  NAND U7698 ( .A(n6140), .B(n4431), .Z(n3527) );
  NANDN U7699 ( .A(init), .B(m[74]), .Z(n4431) );
  AND U7700 ( .A(n6141), .B(n6142), .Z(n6140) );
  NAND U7701 ( .A(o[74]), .B(n5916), .Z(n6142) );
  NANDN U7702 ( .A(n5917), .B(creg[74]), .Z(n6141) );
  NAND U7703 ( .A(n6143), .B(n4429), .Z(n3526) );
  NANDN U7704 ( .A(init), .B(m[75]), .Z(n4429) );
  AND U7705 ( .A(n6144), .B(n6145), .Z(n6143) );
  NAND U7706 ( .A(o[75]), .B(n5916), .Z(n6145) );
  NANDN U7707 ( .A(n5917), .B(creg[75]), .Z(n6144) );
  NAND U7708 ( .A(n6146), .B(n4427), .Z(n3525) );
  NANDN U7709 ( .A(init), .B(m[76]), .Z(n4427) );
  AND U7710 ( .A(n6147), .B(n6148), .Z(n6146) );
  NAND U7711 ( .A(o[76]), .B(n5916), .Z(n6148) );
  NANDN U7712 ( .A(n5917), .B(creg[76]), .Z(n6147) );
  NAND U7713 ( .A(n6149), .B(n4425), .Z(n3524) );
  NANDN U7714 ( .A(init), .B(m[77]), .Z(n4425) );
  AND U7715 ( .A(n6150), .B(n6151), .Z(n6149) );
  NAND U7716 ( .A(o[77]), .B(n5916), .Z(n6151) );
  NANDN U7717 ( .A(n5917), .B(creg[77]), .Z(n6150) );
  NAND U7718 ( .A(n6152), .B(n4423), .Z(n3523) );
  NANDN U7719 ( .A(init), .B(m[78]), .Z(n4423) );
  AND U7720 ( .A(n6153), .B(n6154), .Z(n6152) );
  NAND U7721 ( .A(o[78]), .B(n5916), .Z(n6154) );
  NANDN U7722 ( .A(n5917), .B(creg[78]), .Z(n6153) );
  NAND U7723 ( .A(n6155), .B(n4421), .Z(n3522) );
  NANDN U7724 ( .A(init), .B(m[79]), .Z(n4421) );
  AND U7725 ( .A(n6156), .B(n6157), .Z(n6155) );
  NAND U7726 ( .A(o[79]), .B(n5916), .Z(n6157) );
  NANDN U7727 ( .A(n5917), .B(creg[79]), .Z(n6156) );
  NAND U7728 ( .A(n6158), .B(n4417), .Z(n3521) );
  NANDN U7729 ( .A(init), .B(m[80]), .Z(n4417) );
  AND U7730 ( .A(n6159), .B(n6160), .Z(n6158) );
  NAND U7731 ( .A(o[80]), .B(n5916), .Z(n6160) );
  NANDN U7732 ( .A(n5917), .B(creg[80]), .Z(n6159) );
  NAND U7733 ( .A(n6161), .B(n4415), .Z(n3520) );
  NANDN U7734 ( .A(init), .B(m[81]), .Z(n4415) );
  AND U7735 ( .A(n6162), .B(n6163), .Z(n6161) );
  NAND U7736 ( .A(o[81]), .B(n5916), .Z(n6163) );
  NANDN U7737 ( .A(n5917), .B(creg[81]), .Z(n6162) );
  NAND U7738 ( .A(n6164), .B(n4413), .Z(n3519) );
  NANDN U7739 ( .A(init), .B(m[82]), .Z(n4413) );
  AND U7740 ( .A(n6165), .B(n6166), .Z(n6164) );
  NAND U7741 ( .A(o[82]), .B(n5916), .Z(n6166) );
  NANDN U7742 ( .A(n5917), .B(creg[82]), .Z(n6165) );
  NAND U7743 ( .A(n6167), .B(n4411), .Z(n3518) );
  NANDN U7744 ( .A(init), .B(m[83]), .Z(n4411) );
  AND U7745 ( .A(n6168), .B(n6169), .Z(n6167) );
  NAND U7746 ( .A(o[83]), .B(n5916), .Z(n6169) );
  NANDN U7747 ( .A(n5917), .B(creg[83]), .Z(n6168) );
  NAND U7748 ( .A(n6170), .B(n4409), .Z(n3517) );
  NANDN U7749 ( .A(init), .B(m[84]), .Z(n4409) );
  AND U7750 ( .A(n6171), .B(n6172), .Z(n6170) );
  NAND U7751 ( .A(o[84]), .B(n5916), .Z(n6172) );
  NANDN U7752 ( .A(n5917), .B(creg[84]), .Z(n6171) );
  NAND U7753 ( .A(n6173), .B(n4407), .Z(n3516) );
  NANDN U7754 ( .A(init), .B(m[85]), .Z(n4407) );
  AND U7755 ( .A(n6174), .B(n6175), .Z(n6173) );
  NAND U7756 ( .A(o[85]), .B(n5916), .Z(n6175) );
  NANDN U7757 ( .A(n5917), .B(creg[85]), .Z(n6174) );
  NAND U7758 ( .A(n6176), .B(n4405), .Z(n3515) );
  NANDN U7759 ( .A(init), .B(m[86]), .Z(n4405) );
  AND U7760 ( .A(n6177), .B(n6178), .Z(n6176) );
  NAND U7761 ( .A(o[86]), .B(n5916), .Z(n6178) );
  NANDN U7762 ( .A(n5917), .B(creg[86]), .Z(n6177) );
  NAND U7763 ( .A(n6179), .B(n4403), .Z(n3514) );
  NANDN U7764 ( .A(init), .B(m[87]), .Z(n4403) );
  AND U7765 ( .A(n6180), .B(n6181), .Z(n6179) );
  NAND U7766 ( .A(o[87]), .B(n5916), .Z(n6181) );
  NANDN U7767 ( .A(n5917), .B(creg[87]), .Z(n6180) );
  NAND U7768 ( .A(n6182), .B(n4401), .Z(n3513) );
  NANDN U7769 ( .A(init), .B(m[88]), .Z(n4401) );
  AND U7770 ( .A(n6183), .B(n6184), .Z(n6182) );
  NAND U7771 ( .A(o[88]), .B(n5916), .Z(n6184) );
  NANDN U7772 ( .A(n5917), .B(creg[88]), .Z(n6183) );
  NAND U7773 ( .A(n6185), .B(n4399), .Z(n3512) );
  NANDN U7774 ( .A(init), .B(m[89]), .Z(n4399) );
  AND U7775 ( .A(n6186), .B(n6187), .Z(n6185) );
  NAND U7776 ( .A(o[89]), .B(n5916), .Z(n6187) );
  NANDN U7777 ( .A(n5917), .B(creg[89]), .Z(n6186) );
  NAND U7778 ( .A(n6188), .B(n4395), .Z(n3511) );
  NANDN U7779 ( .A(init), .B(m[90]), .Z(n4395) );
  AND U7780 ( .A(n6189), .B(n6190), .Z(n6188) );
  NAND U7781 ( .A(o[90]), .B(n5916), .Z(n6190) );
  NANDN U7782 ( .A(n5917), .B(creg[90]), .Z(n6189) );
  NAND U7783 ( .A(n6191), .B(n4393), .Z(n3510) );
  NANDN U7784 ( .A(init), .B(m[91]), .Z(n4393) );
  AND U7785 ( .A(n6192), .B(n6193), .Z(n6191) );
  NAND U7786 ( .A(o[91]), .B(n5916), .Z(n6193) );
  NANDN U7787 ( .A(n5917), .B(creg[91]), .Z(n6192) );
  NAND U7788 ( .A(n6194), .B(n4391), .Z(n3509) );
  NANDN U7789 ( .A(init), .B(m[92]), .Z(n4391) );
  AND U7790 ( .A(n6195), .B(n6196), .Z(n6194) );
  NAND U7791 ( .A(o[92]), .B(n5916), .Z(n6196) );
  NANDN U7792 ( .A(n5917), .B(creg[92]), .Z(n6195) );
  NAND U7793 ( .A(n6197), .B(n4389), .Z(n3508) );
  NANDN U7794 ( .A(init), .B(m[93]), .Z(n4389) );
  AND U7795 ( .A(n6198), .B(n6199), .Z(n6197) );
  NAND U7796 ( .A(o[93]), .B(n5916), .Z(n6199) );
  NANDN U7797 ( .A(n5917), .B(creg[93]), .Z(n6198) );
  NAND U7798 ( .A(n6200), .B(n4387), .Z(n3507) );
  NANDN U7799 ( .A(init), .B(m[94]), .Z(n4387) );
  AND U7800 ( .A(n6201), .B(n6202), .Z(n6200) );
  NAND U7801 ( .A(o[94]), .B(n5916), .Z(n6202) );
  NANDN U7802 ( .A(n5917), .B(creg[94]), .Z(n6201) );
  NAND U7803 ( .A(n6203), .B(n4385), .Z(n3506) );
  NANDN U7804 ( .A(init), .B(m[95]), .Z(n4385) );
  AND U7805 ( .A(n6204), .B(n6205), .Z(n6203) );
  NAND U7806 ( .A(o[95]), .B(n5916), .Z(n6205) );
  NANDN U7807 ( .A(n5917), .B(creg[95]), .Z(n6204) );
  NAND U7808 ( .A(n6206), .B(n4383), .Z(n3505) );
  NANDN U7809 ( .A(init), .B(m[96]), .Z(n4383) );
  AND U7810 ( .A(n6207), .B(n6208), .Z(n6206) );
  NAND U7811 ( .A(o[96]), .B(n5916), .Z(n6208) );
  NANDN U7812 ( .A(n5917), .B(creg[96]), .Z(n6207) );
  NAND U7813 ( .A(n6209), .B(n4381), .Z(n3504) );
  NANDN U7814 ( .A(init), .B(m[97]), .Z(n4381) );
  AND U7815 ( .A(n6210), .B(n6211), .Z(n6209) );
  NAND U7816 ( .A(o[97]), .B(n5916), .Z(n6211) );
  NANDN U7817 ( .A(n5917), .B(creg[97]), .Z(n6210) );
  NAND U7818 ( .A(n6212), .B(n4379), .Z(n3503) );
  NANDN U7819 ( .A(init), .B(m[98]), .Z(n4379) );
  AND U7820 ( .A(n6213), .B(n6214), .Z(n6212) );
  NAND U7821 ( .A(o[98]), .B(n5916), .Z(n6214) );
  NANDN U7822 ( .A(n5917), .B(creg[98]), .Z(n6213) );
  NAND U7823 ( .A(n6215), .B(n4377), .Z(n3502) );
  NANDN U7824 ( .A(init), .B(m[99]), .Z(n4377) );
  AND U7825 ( .A(n6216), .B(n6217), .Z(n6215) );
  NAND U7826 ( .A(o[99]), .B(n5916), .Z(n6217) );
  NANDN U7827 ( .A(n5917), .B(creg[99]), .Z(n6216) );
  NAND U7828 ( .A(n6218), .B(n4883), .Z(n3501) );
  NANDN U7829 ( .A(init), .B(m[100]), .Z(n4883) );
  AND U7830 ( .A(n6219), .B(n6220), .Z(n6218) );
  NAND U7831 ( .A(o[100]), .B(n5916), .Z(n6220) );
  NANDN U7832 ( .A(n5917), .B(creg[100]), .Z(n6219) );
  NAND U7833 ( .A(n6221), .B(n4881), .Z(n3500) );
  NANDN U7834 ( .A(init), .B(m[101]), .Z(n4881) );
  AND U7835 ( .A(n6222), .B(n6223), .Z(n6221) );
  NAND U7836 ( .A(o[101]), .B(n5916), .Z(n6223) );
  NANDN U7837 ( .A(n5917), .B(creg[101]), .Z(n6222) );
  NAND U7838 ( .A(n6224), .B(n4879), .Z(n3499) );
  NANDN U7839 ( .A(init), .B(m[102]), .Z(n4879) );
  AND U7840 ( .A(n6225), .B(n6226), .Z(n6224) );
  NAND U7841 ( .A(o[102]), .B(n5916), .Z(n6226) );
  NANDN U7842 ( .A(n5917), .B(creg[102]), .Z(n6225) );
  NAND U7843 ( .A(n6227), .B(n4877), .Z(n3498) );
  NANDN U7844 ( .A(init), .B(m[103]), .Z(n4877) );
  AND U7845 ( .A(n6228), .B(n6229), .Z(n6227) );
  NAND U7846 ( .A(o[103]), .B(n5916), .Z(n6229) );
  NANDN U7847 ( .A(n5917), .B(creg[103]), .Z(n6228) );
  NAND U7848 ( .A(n6230), .B(n4875), .Z(n3497) );
  NANDN U7849 ( .A(init), .B(m[104]), .Z(n4875) );
  AND U7850 ( .A(n6231), .B(n6232), .Z(n6230) );
  NAND U7851 ( .A(o[104]), .B(n5916), .Z(n6232) );
  NANDN U7852 ( .A(n5917), .B(creg[104]), .Z(n6231) );
  NAND U7853 ( .A(n6233), .B(n4873), .Z(n3496) );
  NANDN U7854 ( .A(init), .B(m[105]), .Z(n4873) );
  AND U7855 ( .A(n6234), .B(n6235), .Z(n6233) );
  NAND U7856 ( .A(o[105]), .B(n5916), .Z(n6235) );
  NANDN U7857 ( .A(n5917), .B(creg[105]), .Z(n6234) );
  NAND U7858 ( .A(n6236), .B(n4871), .Z(n3495) );
  NANDN U7859 ( .A(init), .B(m[106]), .Z(n4871) );
  AND U7860 ( .A(n6237), .B(n6238), .Z(n6236) );
  NAND U7861 ( .A(o[106]), .B(n5916), .Z(n6238) );
  NANDN U7862 ( .A(n5917), .B(creg[106]), .Z(n6237) );
  NAND U7863 ( .A(n6239), .B(n4869), .Z(n3494) );
  NANDN U7864 ( .A(init), .B(m[107]), .Z(n4869) );
  AND U7865 ( .A(n6240), .B(n6241), .Z(n6239) );
  NAND U7866 ( .A(o[107]), .B(n5916), .Z(n6241) );
  NANDN U7867 ( .A(n5917), .B(creg[107]), .Z(n6240) );
  NAND U7868 ( .A(n6242), .B(n4867), .Z(n3493) );
  NANDN U7869 ( .A(init), .B(m[108]), .Z(n4867) );
  AND U7870 ( .A(n6243), .B(n6244), .Z(n6242) );
  NAND U7871 ( .A(o[108]), .B(n5916), .Z(n6244) );
  NANDN U7872 ( .A(n5917), .B(creg[108]), .Z(n6243) );
  NAND U7873 ( .A(n6245), .B(n4865), .Z(n3492) );
  NANDN U7874 ( .A(init), .B(m[109]), .Z(n4865) );
  AND U7875 ( .A(n6246), .B(n6247), .Z(n6245) );
  NAND U7876 ( .A(o[109]), .B(n5916), .Z(n6247) );
  NANDN U7877 ( .A(n5917), .B(creg[109]), .Z(n6246) );
  NAND U7878 ( .A(n6248), .B(n4861), .Z(n3491) );
  NANDN U7879 ( .A(init), .B(m[110]), .Z(n4861) );
  AND U7880 ( .A(n6249), .B(n6250), .Z(n6248) );
  NAND U7881 ( .A(o[110]), .B(n5916), .Z(n6250) );
  NANDN U7882 ( .A(n5917), .B(creg[110]), .Z(n6249) );
  NAND U7883 ( .A(n6251), .B(n4859), .Z(n3490) );
  NANDN U7884 ( .A(init), .B(m[111]), .Z(n4859) );
  AND U7885 ( .A(n6252), .B(n6253), .Z(n6251) );
  NAND U7886 ( .A(o[111]), .B(n5916), .Z(n6253) );
  NANDN U7887 ( .A(n5917), .B(creg[111]), .Z(n6252) );
  NAND U7888 ( .A(n6254), .B(n4857), .Z(n3489) );
  NANDN U7889 ( .A(init), .B(m[112]), .Z(n4857) );
  AND U7890 ( .A(n6255), .B(n6256), .Z(n6254) );
  NAND U7891 ( .A(o[112]), .B(n5916), .Z(n6256) );
  NANDN U7892 ( .A(n5917), .B(creg[112]), .Z(n6255) );
  NAND U7893 ( .A(n6257), .B(n4855), .Z(n3488) );
  NANDN U7894 ( .A(init), .B(m[113]), .Z(n4855) );
  AND U7895 ( .A(n6258), .B(n6259), .Z(n6257) );
  NAND U7896 ( .A(o[113]), .B(n5916), .Z(n6259) );
  NANDN U7897 ( .A(n5917), .B(creg[113]), .Z(n6258) );
  NAND U7898 ( .A(n6260), .B(n4853), .Z(n3487) );
  NANDN U7899 ( .A(init), .B(m[114]), .Z(n4853) );
  AND U7900 ( .A(n6261), .B(n6262), .Z(n6260) );
  NAND U7901 ( .A(o[114]), .B(n5916), .Z(n6262) );
  NANDN U7902 ( .A(n5917), .B(creg[114]), .Z(n6261) );
  NAND U7903 ( .A(n6263), .B(n4851), .Z(n3486) );
  NANDN U7904 ( .A(init), .B(m[115]), .Z(n4851) );
  AND U7905 ( .A(n6264), .B(n6265), .Z(n6263) );
  NAND U7906 ( .A(o[115]), .B(n5916), .Z(n6265) );
  NANDN U7907 ( .A(n5917), .B(creg[115]), .Z(n6264) );
  NAND U7908 ( .A(n6266), .B(n4849), .Z(n3485) );
  NANDN U7909 ( .A(init), .B(m[116]), .Z(n4849) );
  AND U7910 ( .A(n6267), .B(n6268), .Z(n6266) );
  NAND U7911 ( .A(o[116]), .B(n5916), .Z(n6268) );
  NANDN U7912 ( .A(n5917), .B(creg[116]), .Z(n6267) );
  NAND U7913 ( .A(n6269), .B(n4847), .Z(n3484) );
  NANDN U7914 ( .A(init), .B(m[117]), .Z(n4847) );
  AND U7915 ( .A(n6270), .B(n6271), .Z(n6269) );
  NAND U7916 ( .A(o[117]), .B(n5916), .Z(n6271) );
  NANDN U7917 ( .A(n5917), .B(creg[117]), .Z(n6270) );
  NAND U7918 ( .A(n6272), .B(n4845), .Z(n3483) );
  NANDN U7919 ( .A(init), .B(m[118]), .Z(n4845) );
  AND U7920 ( .A(n6273), .B(n6274), .Z(n6272) );
  NAND U7921 ( .A(o[118]), .B(n5916), .Z(n6274) );
  NANDN U7922 ( .A(n5917), .B(creg[118]), .Z(n6273) );
  NAND U7923 ( .A(n6275), .B(n4843), .Z(n3482) );
  NANDN U7924 ( .A(init), .B(m[119]), .Z(n4843) );
  AND U7925 ( .A(n6276), .B(n6277), .Z(n6275) );
  NAND U7926 ( .A(o[119]), .B(n5916), .Z(n6277) );
  NANDN U7927 ( .A(n5917), .B(creg[119]), .Z(n6276) );
  NAND U7928 ( .A(n6278), .B(n4839), .Z(n3481) );
  NANDN U7929 ( .A(init), .B(m[120]), .Z(n4839) );
  AND U7930 ( .A(n6279), .B(n6280), .Z(n6278) );
  NAND U7931 ( .A(o[120]), .B(n5916), .Z(n6280) );
  NANDN U7932 ( .A(n5917), .B(creg[120]), .Z(n6279) );
  NAND U7933 ( .A(n6281), .B(n4837), .Z(n3480) );
  NANDN U7934 ( .A(init), .B(m[121]), .Z(n4837) );
  AND U7935 ( .A(n6282), .B(n6283), .Z(n6281) );
  NAND U7936 ( .A(o[121]), .B(n5916), .Z(n6283) );
  NANDN U7937 ( .A(n5917), .B(creg[121]), .Z(n6282) );
  NAND U7938 ( .A(n6284), .B(n4835), .Z(n3479) );
  NANDN U7939 ( .A(init), .B(m[122]), .Z(n4835) );
  AND U7940 ( .A(n6285), .B(n6286), .Z(n6284) );
  NAND U7941 ( .A(o[122]), .B(n5916), .Z(n6286) );
  NANDN U7942 ( .A(n5917), .B(creg[122]), .Z(n6285) );
  NAND U7943 ( .A(n6287), .B(n4833), .Z(n3478) );
  NANDN U7944 ( .A(init), .B(m[123]), .Z(n4833) );
  AND U7945 ( .A(n6288), .B(n6289), .Z(n6287) );
  NAND U7946 ( .A(o[123]), .B(n5916), .Z(n6289) );
  NANDN U7947 ( .A(n5917), .B(creg[123]), .Z(n6288) );
  NAND U7948 ( .A(n6290), .B(n4831), .Z(n3477) );
  NANDN U7949 ( .A(init), .B(m[124]), .Z(n4831) );
  AND U7950 ( .A(n6291), .B(n6292), .Z(n6290) );
  NAND U7951 ( .A(o[124]), .B(n5916), .Z(n6292) );
  NANDN U7952 ( .A(n5917), .B(creg[124]), .Z(n6291) );
  NAND U7953 ( .A(n6293), .B(n4829), .Z(n3476) );
  NANDN U7954 ( .A(init), .B(m[125]), .Z(n4829) );
  AND U7955 ( .A(n6294), .B(n6295), .Z(n6293) );
  NAND U7956 ( .A(o[125]), .B(n5916), .Z(n6295) );
  NANDN U7957 ( .A(n5917), .B(creg[125]), .Z(n6294) );
  NAND U7958 ( .A(n6296), .B(n4827), .Z(n3475) );
  NANDN U7959 ( .A(init), .B(m[126]), .Z(n4827) );
  AND U7960 ( .A(n6297), .B(n6298), .Z(n6296) );
  NAND U7961 ( .A(o[126]), .B(n5916), .Z(n6298) );
  NANDN U7962 ( .A(n5917), .B(creg[126]), .Z(n6297) );
  NAND U7963 ( .A(n6299), .B(n4825), .Z(n3474) );
  NANDN U7964 ( .A(init), .B(m[127]), .Z(n4825) );
  AND U7965 ( .A(n6300), .B(n6301), .Z(n6299) );
  NAND U7966 ( .A(o[127]), .B(n5916), .Z(n6301) );
  NANDN U7967 ( .A(n5917), .B(creg[127]), .Z(n6300) );
  NAND U7968 ( .A(n6302), .B(n4823), .Z(n3473) );
  NANDN U7969 ( .A(init), .B(m[128]), .Z(n4823) );
  AND U7970 ( .A(n6303), .B(n6304), .Z(n6302) );
  NAND U7971 ( .A(o[128]), .B(n5916), .Z(n6304) );
  NANDN U7972 ( .A(n5917), .B(creg[128]), .Z(n6303) );
  NAND U7973 ( .A(n6305), .B(n4821), .Z(n3472) );
  NANDN U7974 ( .A(init), .B(m[129]), .Z(n4821) );
  AND U7975 ( .A(n6306), .B(n6307), .Z(n6305) );
  NAND U7976 ( .A(o[129]), .B(n5916), .Z(n6307) );
  NANDN U7977 ( .A(n5917), .B(creg[129]), .Z(n6306) );
  NAND U7978 ( .A(n6308), .B(n4817), .Z(n3471) );
  NANDN U7979 ( .A(init), .B(m[130]), .Z(n4817) );
  AND U7980 ( .A(n6309), .B(n6310), .Z(n6308) );
  NAND U7981 ( .A(o[130]), .B(n5916), .Z(n6310) );
  NANDN U7982 ( .A(n5917), .B(creg[130]), .Z(n6309) );
  NAND U7983 ( .A(n6311), .B(n4815), .Z(n3470) );
  NANDN U7984 ( .A(init), .B(m[131]), .Z(n4815) );
  AND U7985 ( .A(n6312), .B(n6313), .Z(n6311) );
  NAND U7986 ( .A(o[131]), .B(n5916), .Z(n6313) );
  NANDN U7987 ( .A(n5917), .B(creg[131]), .Z(n6312) );
  NAND U7988 ( .A(n6314), .B(n4813), .Z(n3469) );
  NANDN U7989 ( .A(init), .B(m[132]), .Z(n4813) );
  AND U7990 ( .A(n6315), .B(n6316), .Z(n6314) );
  NAND U7991 ( .A(o[132]), .B(n5916), .Z(n6316) );
  NANDN U7992 ( .A(n5917), .B(creg[132]), .Z(n6315) );
  NAND U7993 ( .A(n6317), .B(n4811), .Z(n3468) );
  NANDN U7994 ( .A(init), .B(m[133]), .Z(n4811) );
  AND U7995 ( .A(n6318), .B(n6319), .Z(n6317) );
  NAND U7996 ( .A(o[133]), .B(n5916), .Z(n6319) );
  NANDN U7997 ( .A(n5917), .B(creg[133]), .Z(n6318) );
  NAND U7998 ( .A(n6320), .B(n4809), .Z(n3467) );
  NANDN U7999 ( .A(init), .B(m[134]), .Z(n4809) );
  AND U8000 ( .A(n6321), .B(n6322), .Z(n6320) );
  NAND U8001 ( .A(o[134]), .B(n5916), .Z(n6322) );
  NANDN U8002 ( .A(n5917), .B(creg[134]), .Z(n6321) );
  NAND U8003 ( .A(n6323), .B(n4807), .Z(n3466) );
  NANDN U8004 ( .A(init), .B(m[135]), .Z(n4807) );
  AND U8005 ( .A(n6324), .B(n6325), .Z(n6323) );
  NAND U8006 ( .A(o[135]), .B(n5916), .Z(n6325) );
  NANDN U8007 ( .A(n5917), .B(creg[135]), .Z(n6324) );
  NAND U8008 ( .A(n6326), .B(n4805), .Z(n3465) );
  NANDN U8009 ( .A(init), .B(m[136]), .Z(n4805) );
  AND U8010 ( .A(n6327), .B(n6328), .Z(n6326) );
  NAND U8011 ( .A(o[136]), .B(n5916), .Z(n6328) );
  NANDN U8012 ( .A(n5917), .B(creg[136]), .Z(n6327) );
  NAND U8013 ( .A(n6329), .B(n4803), .Z(n3464) );
  NANDN U8014 ( .A(init), .B(m[137]), .Z(n4803) );
  AND U8015 ( .A(n6330), .B(n6331), .Z(n6329) );
  NAND U8016 ( .A(o[137]), .B(n5916), .Z(n6331) );
  NANDN U8017 ( .A(n5917), .B(creg[137]), .Z(n6330) );
  NAND U8018 ( .A(n6332), .B(n4801), .Z(n3463) );
  NANDN U8019 ( .A(init), .B(m[138]), .Z(n4801) );
  AND U8020 ( .A(n6333), .B(n6334), .Z(n6332) );
  NAND U8021 ( .A(o[138]), .B(n5916), .Z(n6334) );
  NANDN U8022 ( .A(n5917), .B(creg[138]), .Z(n6333) );
  NAND U8023 ( .A(n6335), .B(n4799), .Z(n3462) );
  NANDN U8024 ( .A(init), .B(m[139]), .Z(n4799) );
  AND U8025 ( .A(n6336), .B(n6337), .Z(n6335) );
  NAND U8026 ( .A(o[139]), .B(n5916), .Z(n6337) );
  NANDN U8027 ( .A(n5917), .B(creg[139]), .Z(n6336) );
  NAND U8028 ( .A(n6338), .B(n4795), .Z(n3461) );
  NANDN U8029 ( .A(init), .B(m[140]), .Z(n4795) );
  AND U8030 ( .A(n6339), .B(n6340), .Z(n6338) );
  NAND U8031 ( .A(o[140]), .B(n5916), .Z(n6340) );
  NANDN U8032 ( .A(n5917), .B(creg[140]), .Z(n6339) );
  NAND U8033 ( .A(n6341), .B(n4793), .Z(n3460) );
  NANDN U8034 ( .A(init), .B(m[141]), .Z(n4793) );
  AND U8035 ( .A(n6342), .B(n6343), .Z(n6341) );
  NAND U8036 ( .A(o[141]), .B(n5916), .Z(n6343) );
  NANDN U8037 ( .A(n5917), .B(creg[141]), .Z(n6342) );
  NAND U8038 ( .A(n6344), .B(n4791), .Z(n3459) );
  NANDN U8039 ( .A(init), .B(m[142]), .Z(n4791) );
  AND U8040 ( .A(n6345), .B(n6346), .Z(n6344) );
  NAND U8041 ( .A(o[142]), .B(n5916), .Z(n6346) );
  NANDN U8042 ( .A(n5917), .B(creg[142]), .Z(n6345) );
  NAND U8043 ( .A(n6347), .B(n4789), .Z(n3458) );
  NANDN U8044 ( .A(init), .B(m[143]), .Z(n4789) );
  AND U8045 ( .A(n6348), .B(n6349), .Z(n6347) );
  NAND U8046 ( .A(o[143]), .B(n5916), .Z(n6349) );
  NANDN U8047 ( .A(n5917), .B(creg[143]), .Z(n6348) );
  NAND U8048 ( .A(n6350), .B(n4787), .Z(n3457) );
  NANDN U8049 ( .A(init), .B(m[144]), .Z(n4787) );
  AND U8050 ( .A(n6351), .B(n6352), .Z(n6350) );
  NAND U8051 ( .A(o[144]), .B(n5916), .Z(n6352) );
  NANDN U8052 ( .A(n5917), .B(creg[144]), .Z(n6351) );
  NAND U8053 ( .A(n6353), .B(n4785), .Z(n3456) );
  NANDN U8054 ( .A(init), .B(m[145]), .Z(n4785) );
  AND U8055 ( .A(n6354), .B(n6355), .Z(n6353) );
  NAND U8056 ( .A(o[145]), .B(n5916), .Z(n6355) );
  NANDN U8057 ( .A(n5917), .B(creg[145]), .Z(n6354) );
  NAND U8058 ( .A(n6356), .B(n4783), .Z(n3455) );
  NANDN U8059 ( .A(init), .B(m[146]), .Z(n4783) );
  AND U8060 ( .A(n6357), .B(n6358), .Z(n6356) );
  NAND U8061 ( .A(o[146]), .B(n5916), .Z(n6358) );
  NANDN U8062 ( .A(n5917), .B(creg[146]), .Z(n6357) );
  NAND U8063 ( .A(n6359), .B(n4781), .Z(n3454) );
  NANDN U8064 ( .A(init), .B(m[147]), .Z(n4781) );
  AND U8065 ( .A(n6360), .B(n6361), .Z(n6359) );
  NAND U8066 ( .A(o[147]), .B(n5916), .Z(n6361) );
  NANDN U8067 ( .A(n5917), .B(creg[147]), .Z(n6360) );
  NAND U8068 ( .A(n6362), .B(n4779), .Z(n3453) );
  NANDN U8069 ( .A(init), .B(m[148]), .Z(n4779) );
  AND U8070 ( .A(n6363), .B(n6364), .Z(n6362) );
  NAND U8071 ( .A(o[148]), .B(n5916), .Z(n6364) );
  NANDN U8072 ( .A(n5917), .B(creg[148]), .Z(n6363) );
  NAND U8073 ( .A(n6365), .B(n4777), .Z(n3452) );
  NANDN U8074 ( .A(init), .B(m[149]), .Z(n4777) );
  AND U8075 ( .A(n6366), .B(n6367), .Z(n6365) );
  NAND U8076 ( .A(o[149]), .B(n5916), .Z(n6367) );
  NANDN U8077 ( .A(n5917), .B(creg[149]), .Z(n6366) );
  NAND U8078 ( .A(n6368), .B(n4773), .Z(n3451) );
  NANDN U8079 ( .A(init), .B(m[150]), .Z(n4773) );
  AND U8080 ( .A(n6369), .B(n6370), .Z(n6368) );
  NAND U8081 ( .A(o[150]), .B(n5916), .Z(n6370) );
  NANDN U8082 ( .A(n5917), .B(creg[150]), .Z(n6369) );
  NAND U8083 ( .A(n6371), .B(n4771), .Z(n3450) );
  NANDN U8084 ( .A(init), .B(m[151]), .Z(n4771) );
  AND U8085 ( .A(n6372), .B(n6373), .Z(n6371) );
  NAND U8086 ( .A(o[151]), .B(n5916), .Z(n6373) );
  NANDN U8087 ( .A(n5917), .B(creg[151]), .Z(n6372) );
  NAND U8088 ( .A(n6374), .B(n4769), .Z(n3449) );
  NANDN U8089 ( .A(init), .B(m[152]), .Z(n4769) );
  AND U8090 ( .A(n6375), .B(n6376), .Z(n6374) );
  NAND U8091 ( .A(o[152]), .B(n5916), .Z(n6376) );
  NANDN U8092 ( .A(n5917), .B(creg[152]), .Z(n6375) );
  NAND U8093 ( .A(n6377), .B(n4767), .Z(n3448) );
  NANDN U8094 ( .A(init), .B(m[153]), .Z(n4767) );
  AND U8095 ( .A(n6378), .B(n6379), .Z(n6377) );
  NAND U8096 ( .A(o[153]), .B(n5916), .Z(n6379) );
  NANDN U8097 ( .A(n5917), .B(creg[153]), .Z(n6378) );
  NAND U8098 ( .A(n6380), .B(n4765), .Z(n3447) );
  NANDN U8099 ( .A(init), .B(m[154]), .Z(n4765) );
  AND U8100 ( .A(n6381), .B(n6382), .Z(n6380) );
  NAND U8101 ( .A(o[154]), .B(n5916), .Z(n6382) );
  NANDN U8102 ( .A(n5917), .B(creg[154]), .Z(n6381) );
  NAND U8103 ( .A(n6383), .B(n4763), .Z(n3446) );
  NANDN U8104 ( .A(init), .B(m[155]), .Z(n4763) );
  AND U8105 ( .A(n6384), .B(n6385), .Z(n6383) );
  NAND U8106 ( .A(o[155]), .B(n5916), .Z(n6385) );
  NANDN U8107 ( .A(n5917), .B(creg[155]), .Z(n6384) );
  NAND U8108 ( .A(n6386), .B(n4761), .Z(n3445) );
  NANDN U8109 ( .A(init), .B(m[156]), .Z(n4761) );
  AND U8110 ( .A(n6387), .B(n6388), .Z(n6386) );
  NAND U8111 ( .A(o[156]), .B(n5916), .Z(n6388) );
  NANDN U8112 ( .A(n5917), .B(creg[156]), .Z(n6387) );
  NAND U8113 ( .A(n6389), .B(n4759), .Z(n3444) );
  NANDN U8114 ( .A(init), .B(m[157]), .Z(n4759) );
  AND U8115 ( .A(n6390), .B(n6391), .Z(n6389) );
  NAND U8116 ( .A(o[157]), .B(n5916), .Z(n6391) );
  NANDN U8117 ( .A(n5917), .B(creg[157]), .Z(n6390) );
  NAND U8118 ( .A(n6392), .B(n4757), .Z(n3443) );
  NANDN U8119 ( .A(init), .B(m[158]), .Z(n4757) );
  AND U8120 ( .A(n6393), .B(n6394), .Z(n6392) );
  NAND U8121 ( .A(o[158]), .B(n5916), .Z(n6394) );
  NANDN U8122 ( .A(n5917), .B(creg[158]), .Z(n6393) );
  NAND U8123 ( .A(n6395), .B(n4755), .Z(n3442) );
  NANDN U8124 ( .A(init), .B(m[159]), .Z(n4755) );
  AND U8125 ( .A(n6396), .B(n6397), .Z(n6395) );
  NAND U8126 ( .A(o[159]), .B(n5916), .Z(n6397) );
  NANDN U8127 ( .A(n5917), .B(creg[159]), .Z(n6396) );
  NAND U8128 ( .A(n6398), .B(n4751), .Z(n3441) );
  NANDN U8129 ( .A(init), .B(m[160]), .Z(n4751) );
  AND U8130 ( .A(n6399), .B(n6400), .Z(n6398) );
  NAND U8131 ( .A(o[160]), .B(n5916), .Z(n6400) );
  NANDN U8132 ( .A(n5917), .B(creg[160]), .Z(n6399) );
  NAND U8133 ( .A(n6401), .B(n4749), .Z(n3440) );
  NANDN U8134 ( .A(init), .B(m[161]), .Z(n4749) );
  AND U8135 ( .A(n6402), .B(n6403), .Z(n6401) );
  NAND U8136 ( .A(o[161]), .B(n5916), .Z(n6403) );
  NANDN U8137 ( .A(n5917), .B(creg[161]), .Z(n6402) );
  NAND U8138 ( .A(n6404), .B(n4747), .Z(n3439) );
  NANDN U8139 ( .A(init), .B(m[162]), .Z(n4747) );
  AND U8140 ( .A(n6405), .B(n6406), .Z(n6404) );
  NAND U8141 ( .A(o[162]), .B(n5916), .Z(n6406) );
  NANDN U8142 ( .A(n5917), .B(creg[162]), .Z(n6405) );
  NAND U8143 ( .A(n6407), .B(n4745), .Z(n3438) );
  NANDN U8144 ( .A(init), .B(m[163]), .Z(n4745) );
  AND U8145 ( .A(n6408), .B(n6409), .Z(n6407) );
  NAND U8146 ( .A(o[163]), .B(n5916), .Z(n6409) );
  NANDN U8147 ( .A(n5917), .B(creg[163]), .Z(n6408) );
  NAND U8148 ( .A(n6410), .B(n4743), .Z(n3437) );
  NANDN U8149 ( .A(init), .B(m[164]), .Z(n4743) );
  AND U8150 ( .A(n6411), .B(n6412), .Z(n6410) );
  NAND U8151 ( .A(o[164]), .B(n5916), .Z(n6412) );
  NANDN U8152 ( .A(n5917), .B(creg[164]), .Z(n6411) );
  NAND U8153 ( .A(n6413), .B(n4741), .Z(n3436) );
  NANDN U8154 ( .A(init), .B(m[165]), .Z(n4741) );
  AND U8155 ( .A(n6414), .B(n6415), .Z(n6413) );
  NAND U8156 ( .A(o[165]), .B(n5916), .Z(n6415) );
  NANDN U8157 ( .A(n5917), .B(creg[165]), .Z(n6414) );
  NAND U8158 ( .A(n6416), .B(n4739), .Z(n3435) );
  NANDN U8159 ( .A(init), .B(m[166]), .Z(n4739) );
  AND U8160 ( .A(n6417), .B(n6418), .Z(n6416) );
  NAND U8161 ( .A(o[166]), .B(n5916), .Z(n6418) );
  NANDN U8162 ( .A(n5917), .B(creg[166]), .Z(n6417) );
  NAND U8163 ( .A(n6419), .B(n4737), .Z(n3434) );
  NANDN U8164 ( .A(init), .B(m[167]), .Z(n4737) );
  AND U8165 ( .A(n6420), .B(n6421), .Z(n6419) );
  NAND U8166 ( .A(o[167]), .B(n5916), .Z(n6421) );
  NANDN U8167 ( .A(n5917), .B(creg[167]), .Z(n6420) );
  NAND U8168 ( .A(n6422), .B(n4735), .Z(n3433) );
  NANDN U8169 ( .A(init), .B(m[168]), .Z(n4735) );
  AND U8170 ( .A(n6423), .B(n6424), .Z(n6422) );
  NAND U8171 ( .A(o[168]), .B(n5916), .Z(n6424) );
  NANDN U8172 ( .A(n5917), .B(creg[168]), .Z(n6423) );
  NAND U8173 ( .A(n6425), .B(n4733), .Z(n3432) );
  NANDN U8174 ( .A(init), .B(m[169]), .Z(n4733) );
  AND U8175 ( .A(n6426), .B(n6427), .Z(n6425) );
  NAND U8176 ( .A(o[169]), .B(n5916), .Z(n6427) );
  NANDN U8177 ( .A(n5917), .B(creg[169]), .Z(n6426) );
  NAND U8178 ( .A(n6428), .B(n4729), .Z(n3431) );
  NANDN U8179 ( .A(init), .B(m[170]), .Z(n4729) );
  AND U8180 ( .A(n6429), .B(n6430), .Z(n6428) );
  NAND U8181 ( .A(o[170]), .B(n5916), .Z(n6430) );
  NANDN U8182 ( .A(n5917), .B(creg[170]), .Z(n6429) );
  NAND U8183 ( .A(n6431), .B(n4727), .Z(n3430) );
  NANDN U8184 ( .A(init), .B(m[171]), .Z(n4727) );
  AND U8185 ( .A(n6432), .B(n6433), .Z(n6431) );
  NAND U8186 ( .A(o[171]), .B(n5916), .Z(n6433) );
  NANDN U8187 ( .A(n5917), .B(creg[171]), .Z(n6432) );
  NAND U8188 ( .A(n6434), .B(n4725), .Z(n3429) );
  NANDN U8189 ( .A(init), .B(m[172]), .Z(n4725) );
  AND U8190 ( .A(n6435), .B(n6436), .Z(n6434) );
  NAND U8191 ( .A(o[172]), .B(n5916), .Z(n6436) );
  NANDN U8192 ( .A(n5917), .B(creg[172]), .Z(n6435) );
  NAND U8193 ( .A(n6437), .B(n4723), .Z(n3428) );
  NANDN U8194 ( .A(init), .B(m[173]), .Z(n4723) );
  AND U8195 ( .A(n6438), .B(n6439), .Z(n6437) );
  NAND U8196 ( .A(o[173]), .B(n5916), .Z(n6439) );
  NANDN U8197 ( .A(n5917), .B(creg[173]), .Z(n6438) );
  NAND U8198 ( .A(n6440), .B(n4721), .Z(n3427) );
  NANDN U8199 ( .A(init), .B(m[174]), .Z(n4721) );
  AND U8200 ( .A(n6441), .B(n6442), .Z(n6440) );
  NAND U8201 ( .A(o[174]), .B(n5916), .Z(n6442) );
  NANDN U8202 ( .A(n5917), .B(creg[174]), .Z(n6441) );
  NAND U8203 ( .A(n6443), .B(n4719), .Z(n3426) );
  NANDN U8204 ( .A(init), .B(m[175]), .Z(n4719) );
  AND U8205 ( .A(n6444), .B(n6445), .Z(n6443) );
  NAND U8206 ( .A(o[175]), .B(n5916), .Z(n6445) );
  NANDN U8207 ( .A(n5917), .B(creg[175]), .Z(n6444) );
  NAND U8208 ( .A(n6446), .B(n4717), .Z(n3425) );
  NANDN U8209 ( .A(init), .B(m[176]), .Z(n4717) );
  AND U8210 ( .A(n6447), .B(n6448), .Z(n6446) );
  NAND U8211 ( .A(o[176]), .B(n5916), .Z(n6448) );
  NANDN U8212 ( .A(n5917), .B(creg[176]), .Z(n6447) );
  NAND U8213 ( .A(n6449), .B(n4715), .Z(n3424) );
  NANDN U8214 ( .A(init), .B(m[177]), .Z(n4715) );
  AND U8215 ( .A(n6450), .B(n6451), .Z(n6449) );
  NAND U8216 ( .A(o[177]), .B(n5916), .Z(n6451) );
  NANDN U8217 ( .A(n5917), .B(creg[177]), .Z(n6450) );
  NAND U8218 ( .A(n6452), .B(n4713), .Z(n3423) );
  NANDN U8219 ( .A(init), .B(m[178]), .Z(n4713) );
  AND U8220 ( .A(n6453), .B(n6454), .Z(n6452) );
  NAND U8221 ( .A(o[178]), .B(n5916), .Z(n6454) );
  NANDN U8222 ( .A(n5917), .B(creg[178]), .Z(n6453) );
  NAND U8223 ( .A(n6455), .B(n4711), .Z(n3422) );
  NANDN U8224 ( .A(init), .B(m[179]), .Z(n4711) );
  AND U8225 ( .A(n6456), .B(n6457), .Z(n6455) );
  NAND U8226 ( .A(o[179]), .B(n5916), .Z(n6457) );
  NANDN U8227 ( .A(n5917), .B(creg[179]), .Z(n6456) );
  NAND U8228 ( .A(n6458), .B(n4707), .Z(n3421) );
  NANDN U8229 ( .A(init), .B(m[180]), .Z(n4707) );
  AND U8230 ( .A(n6459), .B(n6460), .Z(n6458) );
  NAND U8231 ( .A(o[180]), .B(n5916), .Z(n6460) );
  NANDN U8232 ( .A(n5917), .B(creg[180]), .Z(n6459) );
  NAND U8233 ( .A(n6461), .B(n4705), .Z(n3420) );
  NANDN U8234 ( .A(init), .B(m[181]), .Z(n4705) );
  AND U8235 ( .A(n6462), .B(n6463), .Z(n6461) );
  NAND U8236 ( .A(o[181]), .B(n5916), .Z(n6463) );
  NANDN U8237 ( .A(n5917), .B(creg[181]), .Z(n6462) );
  NAND U8238 ( .A(n6464), .B(n4703), .Z(n3419) );
  NANDN U8239 ( .A(init), .B(m[182]), .Z(n4703) );
  AND U8240 ( .A(n6465), .B(n6466), .Z(n6464) );
  NAND U8241 ( .A(o[182]), .B(n5916), .Z(n6466) );
  NANDN U8242 ( .A(n5917), .B(creg[182]), .Z(n6465) );
  NAND U8243 ( .A(n6467), .B(n4701), .Z(n3418) );
  NANDN U8244 ( .A(init), .B(m[183]), .Z(n4701) );
  AND U8245 ( .A(n6468), .B(n6469), .Z(n6467) );
  NAND U8246 ( .A(o[183]), .B(n5916), .Z(n6469) );
  NANDN U8247 ( .A(n5917), .B(creg[183]), .Z(n6468) );
  NAND U8248 ( .A(n6470), .B(n4699), .Z(n3417) );
  NANDN U8249 ( .A(init), .B(m[184]), .Z(n4699) );
  AND U8250 ( .A(n6471), .B(n6472), .Z(n6470) );
  NAND U8251 ( .A(o[184]), .B(n5916), .Z(n6472) );
  NANDN U8252 ( .A(n5917), .B(creg[184]), .Z(n6471) );
  NAND U8253 ( .A(n6473), .B(n4697), .Z(n3416) );
  NANDN U8254 ( .A(init), .B(m[185]), .Z(n4697) );
  AND U8255 ( .A(n6474), .B(n6475), .Z(n6473) );
  NAND U8256 ( .A(o[185]), .B(n5916), .Z(n6475) );
  NANDN U8257 ( .A(n5917), .B(creg[185]), .Z(n6474) );
  NAND U8258 ( .A(n6476), .B(n4695), .Z(n3415) );
  NANDN U8259 ( .A(init), .B(m[186]), .Z(n4695) );
  AND U8260 ( .A(n6477), .B(n6478), .Z(n6476) );
  NAND U8261 ( .A(o[186]), .B(n5916), .Z(n6478) );
  NANDN U8262 ( .A(n5917), .B(creg[186]), .Z(n6477) );
  NAND U8263 ( .A(n6479), .B(n4693), .Z(n3414) );
  NANDN U8264 ( .A(init), .B(m[187]), .Z(n4693) );
  AND U8265 ( .A(n6480), .B(n6481), .Z(n6479) );
  NAND U8266 ( .A(o[187]), .B(n5916), .Z(n6481) );
  NANDN U8267 ( .A(n5917), .B(creg[187]), .Z(n6480) );
  NAND U8268 ( .A(n6482), .B(n4691), .Z(n3413) );
  NANDN U8269 ( .A(init), .B(m[188]), .Z(n4691) );
  AND U8270 ( .A(n6483), .B(n6484), .Z(n6482) );
  NAND U8271 ( .A(o[188]), .B(n5916), .Z(n6484) );
  NANDN U8272 ( .A(n5917), .B(creg[188]), .Z(n6483) );
  NAND U8273 ( .A(n6485), .B(n4689), .Z(n3412) );
  NANDN U8274 ( .A(init), .B(m[189]), .Z(n4689) );
  AND U8275 ( .A(n6486), .B(n6487), .Z(n6485) );
  NAND U8276 ( .A(o[189]), .B(n5916), .Z(n6487) );
  NANDN U8277 ( .A(n5917), .B(creg[189]), .Z(n6486) );
  NAND U8278 ( .A(n6488), .B(n4685), .Z(n3411) );
  NANDN U8279 ( .A(init), .B(m[190]), .Z(n4685) );
  AND U8280 ( .A(n6489), .B(n6490), .Z(n6488) );
  NAND U8281 ( .A(o[190]), .B(n5916), .Z(n6490) );
  NANDN U8282 ( .A(n5917), .B(creg[190]), .Z(n6489) );
  NAND U8283 ( .A(n6491), .B(n4683), .Z(n3410) );
  NANDN U8284 ( .A(init), .B(m[191]), .Z(n4683) );
  AND U8285 ( .A(n6492), .B(n6493), .Z(n6491) );
  NAND U8286 ( .A(o[191]), .B(n5916), .Z(n6493) );
  NANDN U8287 ( .A(n5917), .B(creg[191]), .Z(n6492) );
  NAND U8288 ( .A(n6494), .B(n4681), .Z(n3409) );
  NANDN U8289 ( .A(init), .B(m[192]), .Z(n4681) );
  AND U8290 ( .A(n6495), .B(n6496), .Z(n6494) );
  NAND U8291 ( .A(o[192]), .B(n5916), .Z(n6496) );
  NANDN U8292 ( .A(n5917), .B(creg[192]), .Z(n6495) );
  NAND U8293 ( .A(n6497), .B(n4679), .Z(n3408) );
  NANDN U8294 ( .A(init), .B(m[193]), .Z(n4679) );
  AND U8295 ( .A(n6498), .B(n6499), .Z(n6497) );
  NAND U8296 ( .A(o[193]), .B(n5916), .Z(n6499) );
  NANDN U8297 ( .A(n5917), .B(creg[193]), .Z(n6498) );
  NAND U8298 ( .A(n6500), .B(n4677), .Z(n3407) );
  NANDN U8299 ( .A(init), .B(m[194]), .Z(n4677) );
  AND U8300 ( .A(n6501), .B(n6502), .Z(n6500) );
  NAND U8301 ( .A(o[194]), .B(n5916), .Z(n6502) );
  NANDN U8302 ( .A(n5917), .B(creg[194]), .Z(n6501) );
  NAND U8303 ( .A(n6503), .B(n4675), .Z(n3406) );
  NANDN U8304 ( .A(init), .B(m[195]), .Z(n4675) );
  AND U8305 ( .A(n6504), .B(n6505), .Z(n6503) );
  NAND U8306 ( .A(o[195]), .B(n5916), .Z(n6505) );
  NANDN U8307 ( .A(n5917), .B(creg[195]), .Z(n6504) );
  NAND U8308 ( .A(n6506), .B(n4673), .Z(n3405) );
  NANDN U8309 ( .A(init), .B(m[196]), .Z(n4673) );
  AND U8310 ( .A(n6507), .B(n6508), .Z(n6506) );
  NAND U8311 ( .A(o[196]), .B(n5916), .Z(n6508) );
  NANDN U8312 ( .A(n5917), .B(creg[196]), .Z(n6507) );
  NAND U8313 ( .A(n6509), .B(n4671), .Z(n3404) );
  NANDN U8314 ( .A(init), .B(m[197]), .Z(n4671) );
  AND U8315 ( .A(n6510), .B(n6511), .Z(n6509) );
  NAND U8316 ( .A(o[197]), .B(n5916), .Z(n6511) );
  NANDN U8317 ( .A(n5917), .B(creg[197]), .Z(n6510) );
  NAND U8318 ( .A(n6512), .B(n4669), .Z(n3403) );
  NANDN U8319 ( .A(init), .B(m[198]), .Z(n4669) );
  AND U8320 ( .A(n6513), .B(n6514), .Z(n6512) );
  NAND U8321 ( .A(o[198]), .B(n5916), .Z(n6514) );
  NANDN U8322 ( .A(n5917), .B(creg[198]), .Z(n6513) );
  NAND U8323 ( .A(n6515), .B(n4667), .Z(n3402) );
  NANDN U8324 ( .A(init), .B(m[199]), .Z(n4667) );
  AND U8325 ( .A(n6516), .B(n6517), .Z(n6515) );
  NAND U8326 ( .A(o[199]), .B(n5916), .Z(n6517) );
  NANDN U8327 ( .A(n5917), .B(creg[199]), .Z(n6516) );
  NAND U8328 ( .A(n6518), .B(n4661), .Z(n3401) );
  NANDN U8329 ( .A(init), .B(m[200]), .Z(n4661) );
  AND U8330 ( .A(n6519), .B(n6520), .Z(n6518) );
  NAND U8331 ( .A(o[200]), .B(n5916), .Z(n6520) );
  NANDN U8332 ( .A(n5917), .B(creg[200]), .Z(n6519) );
  NAND U8333 ( .A(n6521), .B(n4659), .Z(n3400) );
  NANDN U8334 ( .A(init), .B(m[201]), .Z(n4659) );
  AND U8335 ( .A(n6522), .B(n6523), .Z(n6521) );
  NAND U8336 ( .A(o[201]), .B(n5916), .Z(n6523) );
  NANDN U8337 ( .A(n5917), .B(creg[201]), .Z(n6522) );
  NAND U8338 ( .A(n6524), .B(n4657), .Z(n3399) );
  NANDN U8339 ( .A(init), .B(m[202]), .Z(n4657) );
  AND U8340 ( .A(n6525), .B(n6526), .Z(n6524) );
  NAND U8341 ( .A(o[202]), .B(n5916), .Z(n6526) );
  NANDN U8342 ( .A(n5917), .B(creg[202]), .Z(n6525) );
  NAND U8343 ( .A(n6527), .B(n4655), .Z(n3398) );
  NANDN U8344 ( .A(init), .B(m[203]), .Z(n4655) );
  AND U8345 ( .A(n6528), .B(n6529), .Z(n6527) );
  NAND U8346 ( .A(o[203]), .B(n5916), .Z(n6529) );
  NANDN U8347 ( .A(n5917), .B(creg[203]), .Z(n6528) );
  NAND U8348 ( .A(n6530), .B(n4653), .Z(n3397) );
  NANDN U8349 ( .A(init), .B(m[204]), .Z(n4653) );
  AND U8350 ( .A(n6531), .B(n6532), .Z(n6530) );
  NAND U8351 ( .A(o[204]), .B(n5916), .Z(n6532) );
  NANDN U8352 ( .A(n5917), .B(creg[204]), .Z(n6531) );
  NAND U8353 ( .A(n6533), .B(n4651), .Z(n3396) );
  NANDN U8354 ( .A(init), .B(m[205]), .Z(n4651) );
  AND U8355 ( .A(n6534), .B(n6535), .Z(n6533) );
  NAND U8356 ( .A(o[205]), .B(n5916), .Z(n6535) );
  NANDN U8357 ( .A(n5917), .B(creg[205]), .Z(n6534) );
  NAND U8358 ( .A(n6536), .B(n4649), .Z(n3395) );
  NANDN U8359 ( .A(init), .B(m[206]), .Z(n4649) );
  AND U8360 ( .A(n6537), .B(n6538), .Z(n6536) );
  NAND U8361 ( .A(o[206]), .B(n5916), .Z(n6538) );
  NANDN U8362 ( .A(n5917), .B(creg[206]), .Z(n6537) );
  NAND U8363 ( .A(n6539), .B(n4647), .Z(n3394) );
  NANDN U8364 ( .A(init), .B(m[207]), .Z(n4647) );
  AND U8365 ( .A(n6540), .B(n6541), .Z(n6539) );
  NAND U8366 ( .A(o[207]), .B(n5916), .Z(n6541) );
  NANDN U8367 ( .A(n5917), .B(creg[207]), .Z(n6540) );
  NAND U8368 ( .A(n6542), .B(n4645), .Z(n3393) );
  NANDN U8369 ( .A(init), .B(m[208]), .Z(n4645) );
  AND U8370 ( .A(n6543), .B(n6544), .Z(n6542) );
  NAND U8371 ( .A(o[208]), .B(n5916), .Z(n6544) );
  NANDN U8372 ( .A(n5917), .B(creg[208]), .Z(n6543) );
  NAND U8373 ( .A(n6545), .B(n4643), .Z(n3392) );
  NANDN U8374 ( .A(init), .B(m[209]), .Z(n4643) );
  AND U8375 ( .A(n6546), .B(n6547), .Z(n6545) );
  NAND U8376 ( .A(o[209]), .B(n5916), .Z(n6547) );
  NANDN U8377 ( .A(n5917), .B(creg[209]), .Z(n6546) );
  NAND U8378 ( .A(n6548), .B(n4639), .Z(n3391) );
  NANDN U8379 ( .A(init), .B(m[210]), .Z(n4639) );
  AND U8380 ( .A(n6549), .B(n6550), .Z(n6548) );
  NAND U8381 ( .A(o[210]), .B(n5916), .Z(n6550) );
  NANDN U8382 ( .A(n5917), .B(creg[210]), .Z(n6549) );
  NAND U8383 ( .A(n6551), .B(n4637), .Z(n3390) );
  NANDN U8384 ( .A(init), .B(m[211]), .Z(n4637) );
  AND U8385 ( .A(n6552), .B(n6553), .Z(n6551) );
  NAND U8386 ( .A(o[211]), .B(n5916), .Z(n6553) );
  NANDN U8387 ( .A(n5917), .B(creg[211]), .Z(n6552) );
  NAND U8388 ( .A(n6554), .B(n4635), .Z(n3389) );
  NANDN U8389 ( .A(init), .B(m[212]), .Z(n4635) );
  AND U8390 ( .A(n6555), .B(n6556), .Z(n6554) );
  NAND U8391 ( .A(o[212]), .B(n5916), .Z(n6556) );
  NANDN U8392 ( .A(n5917), .B(creg[212]), .Z(n6555) );
  NAND U8393 ( .A(n6557), .B(n4633), .Z(n3388) );
  NANDN U8394 ( .A(init), .B(m[213]), .Z(n4633) );
  AND U8395 ( .A(n6558), .B(n6559), .Z(n6557) );
  NAND U8396 ( .A(o[213]), .B(n5916), .Z(n6559) );
  NANDN U8397 ( .A(n5917), .B(creg[213]), .Z(n6558) );
  NAND U8398 ( .A(n6560), .B(n4631), .Z(n3387) );
  NANDN U8399 ( .A(init), .B(m[214]), .Z(n4631) );
  AND U8400 ( .A(n6561), .B(n6562), .Z(n6560) );
  NAND U8401 ( .A(o[214]), .B(n5916), .Z(n6562) );
  NANDN U8402 ( .A(n5917), .B(creg[214]), .Z(n6561) );
  NAND U8403 ( .A(n6563), .B(n4629), .Z(n3386) );
  NANDN U8404 ( .A(init), .B(m[215]), .Z(n4629) );
  AND U8405 ( .A(n6564), .B(n6565), .Z(n6563) );
  NAND U8406 ( .A(o[215]), .B(n5916), .Z(n6565) );
  NANDN U8407 ( .A(n5917), .B(creg[215]), .Z(n6564) );
  NAND U8408 ( .A(n6566), .B(n4627), .Z(n3385) );
  NANDN U8409 ( .A(init), .B(m[216]), .Z(n4627) );
  AND U8410 ( .A(n6567), .B(n6568), .Z(n6566) );
  NAND U8411 ( .A(o[216]), .B(n5916), .Z(n6568) );
  NANDN U8412 ( .A(n5917), .B(creg[216]), .Z(n6567) );
  NAND U8413 ( .A(n6569), .B(n4625), .Z(n3384) );
  NANDN U8414 ( .A(init), .B(m[217]), .Z(n4625) );
  AND U8415 ( .A(n6570), .B(n6571), .Z(n6569) );
  NAND U8416 ( .A(o[217]), .B(n5916), .Z(n6571) );
  NANDN U8417 ( .A(n5917), .B(creg[217]), .Z(n6570) );
  NAND U8418 ( .A(n6572), .B(n4623), .Z(n3383) );
  NANDN U8419 ( .A(init), .B(m[218]), .Z(n4623) );
  AND U8420 ( .A(n6573), .B(n6574), .Z(n6572) );
  NAND U8421 ( .A(o[218]), .B(n5916), .Z(n6574) );
  NANDN U8422 ( .A(n5917), .B(creg[218]), .Z(n6573) );
  NAND U8423 ( .A(n6575), .B(n4621), .Z(n3382) );
  NANDN U8424 ( .A(init), .B(m[219]), .Z(n4621) );
  AND U8425 ( .A(n6576), .B(n6577), .Z(n6575) );
  NAND U8426 ( .A(o[219]), .B(n5916), .Z(n6577) );
  NANDN U8427 ( .A(n5917), .B(creg[219]), .Z(n6576) );
  NAND U8428 ( .A(n6578), .B(n4617), .Z(n3381) );
  NANDN U8429 ( .A(init), .B(m[220]), .Z(n4617) );
  AND U8430 ( .A(n6579), .B(n6580), .Z(n6578) );
  NAND U8431 ( .A(o[220]), .B(n5916), .Z(n6580) );
  NANDN U8432 ( .A(n5917), .B(creg[220]), .Z(n6579) );
  NAND U8433 ( .A(n6581), .B(n4615), .Z(n3380) );
  NANDN U8434 ( .A(init), .B(m[221]), .Z(n4615) );
  AND U8435 ( .A(n6582), .B(n6583), .Z(n6581) );
  NAND U8436 ( .A(o[221]), .B(n5916), .Z(n6583) );
  NANDN U8437 ( .A(n5917), .B(creg[221]), .Z(n6582) );
  NAND U8438 ( .A(n6584), .B(n4613), .Z(n3379) );
  NANDN U8439 ( .A(init), .B(m[222]), .Z(n4613) );
  AND U8440 ( .A(n6585), .B(n6586), .Z(n6584) );
  NAND U8441 ( .A(o[222]), .B(n5916), .Z(n6586) );
  NANDN U8442 ( .A(n5917), .B(creg[222]), .Z(n6585) );
  NAND U8443 ( .A(n6587), .B(n4611), .Z(n3378) );
  NANDN U8444 ( .A(init), .B(m[223]), .Z(n4611) );
  AND U8445 ( .A(n6588), .B(n6589), .Z(n6587) );
  NAND U8446 ( .A(o[223]), .B(n5916), .Z(n6589) );
  NANDN U8447 ( .A(n5917), .B(creg[223]), .Z(n6588) );
  NAND U8448 ( .A(n6590), .B(n4609), .Z(n3377) );
  NANDN U8449 ( .A(init), .B(m[224]), .Z(n4609) );
  AND U8450 ( .A(n6591), .B(n6592), .Z(n6590) );
  NAND U8451 ( .A(o[224]), .B(n5916), .Z(n6592) );
  NANDN U8452 ( .A(n5917), .B(creg[224]), .Z(n6591) );
  NAND U8453 ( .A(n6593), .B(n4607), .Z(n3376) );
  NANDN U8454 ( .A(init), .B(m[225]), .Z(n4607) );
  AND U8455 ( .A(n6594), .B(n6595), .Z(n6593) );
  NAND U8456 ( .A(o[225]), .B(n5916), .Z(n6595) );
  NANDN U8457 ( .A(n5917), .B(creg[225]), .Z(n6594) );
  NAND U8458 ( .A(n6596), .B(n4605), .Z(n3375) );
  NANDN U8459 ( .A(init), .B(m[226]), .Z(n4605) );
  AND U8460 ( .A(n6597), .B(n6598), .Z(n6596) );
  NAND U8461 ( .A(o[226]), .B(n5916), .Z(n6598) );
  NANDN U8462 ( .A(n5917), .B(creg[226]), .Z(n6597) );
  NAND U8463 ( .A(n6599), .B(n4603), .Z(n3374) );
  NANDN U8464 ( .A(init), .B(m[227]), .Z(n4603) );
  AND U8465 ( .A(n6600), .B(n6601), .Z(n6599) );
  NAND U8466 ( .A(o[227]), .B(n5916), .Z(n6601) );
  NANDN U8467 ( .A(n5917), .B(creg[227]), .Z(n6600) );
  NAND U8468 ( .A(n6602), .B(n4601), .Z(n3373) );
  NANDN U8469 ( .A(init), .B(m[228]), .Z(n4601) );
  AND U8470 ( .A(n6603), .B(n6604), .Z(n6602) );
  NAND U8471 ( .A(o[228]), .B(n5916), .Z(n6604) );
  NANDN U8472 ( .A(n5917), .B(creg[228]), .Z(n6603) );
  NAND U8473 ( .A(n6605), .B(n4599), .Z(n3372) );
  NANDN U8474 ( .A(init), .B(m[229]), .Z(n4599) );
  AND U8475 ( .A(n6606), .B(n6607), .Z(n6605) );
  NAND U8476 ( .A(o[229]), .B(n5916), .Z(n6607) );
  NANDN U8477 ( .A(n5917), .B(creg[229]), .Z(n6606) );
  NAND U8478 ( .A(n6608), .B(n4595), .Z(n3371) );
  NANDN U8479 ( .A(init), .B(m[230]), .Z(n4595) );
  AND U8480 ( .A(n6609), .B(n6610), .Z(n6608) );
  NAND U8481 ( .A(o[230]), .B(n5916), .Z(n6610) );
  NANDN U8482 ( .A(n5917), .B(creg[230]), .Z(n6609) );
  NAND U8483 ( .A(n6611), .B(n4593), .Z(n3370) );
  NANDN U8484 ( .A(init), .B(m[231]), .Z(n4593) );
  AND U8485 ( .A(n6612), .B(n6613), .Z(n6611) );
  NAND U8486 ( .A(o[231]), .B(n5916), .Z(n6613) );
  NANDN U8487 ( .A(n5917), .B(creg[231]), .Z(n6612) );
  NAND U8488 ( .A(n6614), .B(n4591), .Z(n3369) );
  NANDN U8489 ( .A(init), .B(m[232]), .Z(n4591) );
  AND U8490 ( .A(n6615), .B(n6616), .Z(n6614) );
  NAND U8491 ( .A(o[232]), .B(n5916), .Z(n6616) );
  NANDN U8492 ( .A(n5917), .B(creg[232]), .Z(n6615) );
  NAND U8493 ( .A(n6617), .B(n4589), .Z(n3368) );
  NANDN U8494 ( .A(init), .B(m[233]), .Z(n4589) );
  AND U8495 ( .A(n6618), .B(n6619), .Z(n6617) );
  NAND U8496 ( .A(o[233]), .B(n5916), .Z(n6619) );
  NANDN U8497 ( .A(n5917), .B(creg[233]), .Z(n6618) );
  NAND U8498 ( .A(n6620), .B(n4587), .Z(n3367) );
  NANDN U8499 ( .A(init), .B(m[234]), .Z(n4587) );
  AND U8500 ( .A(n6621), .B(n6622), .Z(n6620) );
  NAND U8501 ( .A(o[234]), .B(n5916), .Z(n6622) );
  NANDN U8502 ( .A(n5917), .B(creg[234]), .Z(n6621) );
  NAND U8503 ( .A(n6623), .B(n4585), .Z(n3366) );
  NANDN U8504 ( .A(init), .B(m[235]), .Z(n4585) );
  AND U8505 ( .A(n6624), .B(n6625), .Z(n6623) );
  NAND U8506 ( .A(o[235]), .B(n5916), .Z(n6625) );
  NANDN U8507 ( .A(n5917), .B(creg[235]), .Z(n6624) );
  NAND U8508 ( .A(n6626), .B(n4583), .Z(n3365) );
  NANDN U8509 ( .A(init), .B(m[236]), .Z(n4583) );
  AND U8510 ( .A(n6627), .B(n6628), .Z(n6626) );
  NAND U8511 ( .A(o[236]), .B(n5916), .Z(n6628) );
  NANDN U8512 ( .A(n5917), .B(creg[236]), .Z(n6627) );
  NAND U8513 ( .A(n6629), .B(n4581), .Z(n3364) );
  NANDN U8514 ( .A(init), .B(m[237]), .Z(n4581) );
  AND U8515 ( .A(n6630), .B(n6631), .Z(n6629) );
  NAND U8516 ( .A(o[237]), .B(n5916), .Z(n6631) );
  NANDN U8517 ( .A(n5917), .B(creg[237]), .Z(n6630) );
  NAND U8518 ( .A(n6632), .B(n4579), .Z(n3363) );
  NANDN U8519 ( .A(init), .B(m[238]), .Z(n4579) );
  AND U8520 ( .A(n6633), .B(n6634), .Z(n6632) );
  NAND U8521 ( .A(o[238]), .B(n5916), .Z(n6634) );
  NANDN U8522 ( .A(n5917), .B(creg[238]), .Z(n6633) );
  NAND U8523 ( .A(n6635), .B(n4577), .Z(n3362) );
  NANDN U8524 ( .A(init), .B(m[239]), .Z(n4577) );
  AND U8525 ( .A(n6636), .B(n6637), .Z(n6635) );
  NAND U8526 ( .A(o[239]), .B(n5916), .Z(n6637) );
  NANDN U8527 ( .A(n5917), .B(creg[239]), .Z(n6636) );
  NAND U8528 ( .A(n6638), .B(n4573), .Z(n3361) );
  NANDN U8529 ( .A(init), .B(m[240]), .Z(n4573) );
  AND U8530 ( .A(n6639), .B(n6640), .Z(n6638) );
  NAND U8531 ( .A(o[240]), .B(n5916), .Z(n6640) );
  NANDN U8532 ( .A(n5917), .B(creg[240]), .Z(n6639) );
  NAND U8533 ( .A(n6641), .B(n4571), .Z(n3360) );
  NANDN U8534 ( .A(init), .B(m[241]), .Z(n4571) );
  AND U8535 ( .A(n6642), .B(n6643), .Z(n6641) );
  NAND U8536 ( .A(o[241]), .B(n5916), .Z(n6643) );
  NANDN U8537 ( .A(n5917), .B(creg[241]), .Z(n6642) );
  NAND U8538 ( .A(n6644), .B(n4569), .Z(n3359) );
  NANDN U8539 ( .A(init), .B(m[242]), .Z(n4569) );
  AND U8540 ( .A(n6645), .B(n6646), .Z(n6644) );
  NAND U8541 ( .A(o[242]), .B(n5916), .Z(n6646) );
  NANDN U8542 ( .A(n5917), .B(creg[242]), .Z(n6645) );
  NAND U8543 ( .A(n6647), .B(n4567), .Z(n3358) );
  NANDN U8544 ( .A(init), .B(m[243]), .Z(n4567) );
  AND U8545 ( .A(n6648), .B(n6649), .Z(n6647) );
  NAND U8546 ( .A(o[243]), .B(n5916), .Z(n6649) );
  NANDN U8547 ( .A(n5917), .B(creg[243]), .Z(n6648) );
  NAND U8548 ( .A(n6650), .B(n4565), .Z(n3357) );
  NANDN U8549 ( .A(init), .B(m[244]), .Z(n4565) );
  AND U8550 ( .A(n6651), .B(n6652), .Z(n6650) );
  NAND U8551 ( .A(o[244]), .B(n5916), .Z(n6652) );
  NANDN U8552 ( .A(n5917), .B(creg[244]), .Z(n6651) );
  NAND U8553 ( .A(n6653), .B(n4563), .Z(n3356) );
  NANDN U8554 ( .A(init), .B(m[245]), .Z(n4563) );
  AND U8555 ( .A(n6654), .B(n6655), .Z(n6653) );
  NAND U8556 ( .A(o[245]), .B(n5916), .Z(n6655) );
  NANDN U8557 ( .A(n5917), .B(creg[245]), .Z(n6654) );
  NAND U8558 ( .A(n6656), .B(n4561), .Z(n3355) );
  NANDN U8559 ( .A(init), .B(m[246]), .Z(n4561) );
  AND U8560 ( .A(n6657), .B(n6658), .Z(n6656) );
  NAND U8561 ( .A(o[246]), .B(n5916), .Z(n6658) );
  NANDN U8562 ( .A(n5917), .B(creg[246]), .Z(n6657) );
  NAND U8563 ( .A(n6659), .B(n4559), .Z(n3354) );
  NANDN U8564 ( .A(init), .B(m[247]), .Z(n4559) );
  AND U8565 ( .A(n6660), .B(n6661), .Z(n6659) );
  NAND U8566 ( .A(o[247]), .B(n5916), .Z(n6661) );
  NANDN U8567 ( .A(n5917), .B(creg[247]), .Z(n6660) );
  NAND U8568 ( .A(n6662), .B(n4557), .Z(n3353) );
  NANDN U8569 ( .A(init), .B(m[248]), .Z(n4557) );
  AND U8570 ( .A(n6663), .B(n6664), .Z(n6662) );
  NAND U8571 ( .A(o[248]), .B(n5916), .Z(n6664) );
  NANDN U8572 ( .A(n5917), .B(creg[248]), .Z(n6663) );
  NAND U8573 ( .A(n6665), .B(n4555), .Z(n3352) );
  NANDN U8574 ( .A(init), .B(m[249]), .Z(n4555) );
  AND U8575 ( .A(n6666), .B(n6667), .Z(n6665) );
  NAND U8576 ( .A(o[249]), .B(n5916), .Z(n6667) );
  NANDN U8577 ( .A(n5917), .B(creg[249]), .Z(n6666) );
  NAND U8578 ( .A(n6668), .B(n4551), .Z(n3351) );
  NANDN U8579 ( .A(init), .B(m[250]), .Z(n4551) );
  AND U8580 ( .A(n6669), .B(n6670), .Z(n6668) );
  NAND U8581 ( .A(o[250]), .B(n5916), .Z(n6670) );
  NANDN U8582 ( .A(n5917), .B(creg[250]), .Z(n6669) );
  NAND U8583 ( .A(n6671), .B(n4549), .Z(n3350) );
  NANDN U8584 ( .A(init), .B(m[251]), .Z(n4549) );
  AND U8585 ( .A(n6672), .B(n6673), .Z(n6671) );
  NAND U8586 ( .A(o[251]), .B(n5916), .Z(n6673) );
  NANDN U8587 ( .A(n5917), .B(creg[251]), .Z(n6672) );
  NAND U8588 ( .A(n6674), .B(n4547), .Z(n3349) );
  NANDN U8589 ( .A(init), .B(m[252]), .Z(n4547) );
  AND U8590 ( .A(n6675), .B(n6676), .Z(n6674) );
  NAND U8591 ( .A(o[252]), .B(n5916), .Z(n6676) );
  NANDN U8592 ( .A(n5917), .B(creg[252]), .Z(n6675) );
  NAND U8593 ( .A(n6677), .B(n4545), .Z(n3348) );
  NANDN U8594 ( .A(init), .B(m[253]), .Z(n4545) );
  AND U8595 ( .A(n6678), .B(n6679), .Z(n6677) );
  NAND U8596 ( .A(o[253]), .B(n5916), .Z(n6679) );
  NANDN U8597 ( .A(n5917), .B(creg[253]), .Z(n6678) );
  NAND U8598 ( .A(n6680), .B(n4543), .Z(n3347) );
  NANDN U8599 ( .A(init), .B(m[254]), .Z(n4543) );
  AND U8600 ( .A(n6681), .B(n6682), .Z(n6680) );
  NAND U8601 ( .A(o[254]), .B(n5916), .Z(n6682) );
  AND U8602 ( .A(n7204), .B(n5917), .Z(n5916) );
  NANDN U8603 ( .A(n5917), .B(creg[254]), .Z(n6681) );
  NAND U8604 ( .A(init), .B(n6683), .Z(n5917) );
  NAND U8605 ( .A(first_one), .B(n6684), .Z(n6683) );
  AND U8606 ( .A(start_reg[63]), .B(n6685), .Z(n6684) );
  NAND U8607 ( .A(n6686), .B(mul_pow), .Z(n6685) );
  NANDN U8608 ( .A(first_one), .B(n6687), .Z(n3346) );
  NAND U8609 ( .A(n6688), .B(ereg[255]), .Z(n6687) );
  AND U8610 ( .A(n7204), .B(mul_pow), .Z(n6688) );
  AND U8611 ( .A(start_reg[63]), .B(init), .Z(n7204) );
  NAND U8612 ( .A(n6689), .B(n6690), .Z(c[9]) );
  NAND U8613 ( .A(n6691), .B(o[9]), .Z(n6690) );
  NAND U8614 ( .A(n6686), .B(creg[9]), .Z(n6689) );
  NAND U8615 ( .A(n6692), .B(n6693), .Z(c[99]) );
  NAND U8616 ( .A(n6691), .B(o[99]), .Z(n6693) );
  NAND U8617 ( .A(n6686), .B(creg[99]), .Z(n6692) );
  NAND U8618 ( .A(n6694), .B(n6695), .Z(c[98]) );
  NAND U8619 ( .A(n6691), .B(o[98]), .Z(n6695) );
  NAND U8620 ( .A(n6686), .B(creg[98]), .Z(n6694) );
  NAND U8621 ( .A(n6696), .B(n6697), .Z(c[97]) );
  NAND U8622 ( .A(n6691), .B(o[97]), .Z(n6697) );
  NAND U8623 ( .A(n6686), .B(creg[97]), .Z(n6696) );
  NAND U8624 ( .A(n6698), .B(n6699), .Z(c[96]) );
  NAND U8625 ( .A(n6691), .B(o[96]), .Z(n6699) );
  NAND U8626 ( .A(n6686), .B(creg[96]), .Z(n6698) );
  NAND U8627 ( .A(n6700), .B(n6701), .Z(c[95]) );
  NAND U8628 ( .A(n6691), .B(o[95]), .Z(n6701) );
  NAND U8629 ( .A(n6686), .B(creg[95]), .Z(n6700) );
  NAND U8630 ( .A(n6702), .B(n6703), .Z(c[94]) );
  NAND U8631 ( .A(n6691), .B(o[94]), .Z(n6703) );
  NAND U8632 ( .A(n6686), .B(creg[94]), .Z(n6702) );
  NAND U8633 ( .A(n6704), .B(n6705), .Z(c[93]) );
  NAND U8634 ( .A(n6691), .B(o[93]), .Z(n6705) );
  NAND U8635 ( .A(n6686), .B(creg[93]), .Z(n6704) );
  NAND U8636 ( .A(n6706), .B(n6707), .Z(c[92]) );
  NAND U8637 ( .A(n6691), .B(o[92]), .Z(n6707) );
  NAND U8638 ( .A(n6686), .B(creg[92]), .Z(n6706) );
  NAND U8639 ( .A(n6708), .B(n6709), .Z(c[91]) );
  NAND U8640 ( .A(n6691), .B(o[91]), .Z(n6709) );
  NAND U8641 ( .A(n6686), .B(creg[91]), .Z(n6708) );
  NAND U8642 ( .A(n6710), .B(n6711), .Z(c[90]) );
  NAND U8643 ( .A(n6691), .B(o[90]), .Z(n6711) );
  NAND U8644 ( .A(n6686), .B(creg[90]), .Z(n6710) );
  NAND U8645 ( .A(n6712), .B(n6713), .Z(c[8]) );
  NAND U8646 ( .A(n6691), .B(o[8]), .Z(n6713) );
  NAND U8647 ( .A(n6686), .B(creg[8]), .Z(n6712) );
  NAND U8648 ( .A(n6714), .B(n6715), .Z(c[89]) );
  NAND U8649 ( .A(n6691), .B(o[89]), .Z(n6715) );
  NAND U8650 ( .A(n6686), .B(creg[89]), .Z(n6714) );
  NAND U8651 ( .A(n6716), .B(n6717), .Z(c[88]) );
  NAND U8652 ( .A(n6691), .B(o[88]), .Z(n6717) );
  NAND U8653 ( .A(n6686), .B(creg[88]), .Z(n6716) );
  NAND U8654 ( .A(n6718), .B(n6719), .Z(c[87]) );
  NAND U8655 ( .A(n6691), .B(o[87]), .Z(n6719) );
  NAND U8656 ( .A(n6686), .B(creg[87]), .Z(n6718) );
  NAND U8657 ( .A(n6720), .B(n6721), .Z(c[86]) );
  NAND U8658 ( .A(n6691), .B(o[86]), .Z(n6721) );
  NAND U8659 ( .A(n6686), .B(creg[86]), .Z(n6720) );
  NAND U8660 ( .A(n6722), .B(n6723), .Z(c[85]) );
  NAND U8661 ( .A(n6691), .B(o[85]), .Z(n6723) );
  NAND U8662 ( .A(n6686), .B(creg[85]), .Z(n6722) );
  NAND U8663 ( .A(n6724), .B(n6725), .Z(c[84]) );
  NAND U8664 ( .A(n6691), .B(o[84]), .Z(n6725) );
  NAND U8665 ( .A(n6686), .B(creg[84]), .Z(n6724) );
  NAND U8666 ( .A(n6726), .B(n6727), .Z(c[83]) );
  NAND U8667 ( .A(n6691), .B(o[83]), .Z(n6727) );
  NAND U8668 ( .A(n6686), .B(creg[83]), .Z(n6726) );
  NAND U8669 ( .A(n6728), .B(n6729), .Z(c[82]) );
  NAND U8670 ( .A(n6691), .B(o[82]), .Z(n6729) );
  NAND U8671 ( .A(n6686), .B(creg[82]), .Z(n6728) );
  NAND U8672 ( .A(n6730), .B(n6731), .Z(c[81]) );
  NAND U8673 ( .A(n6691), .B(o[81]), .Z(n6731) );
  NAND U8674 ( .A(n6686), .B(creg[81]), .Z(n6730) );
  NAND U8675 ( .A(n6732), .B(n6733), .Z(c[80]) );
  NAND U8676 ( .A(n6691), .B(o[80]), .Z(n6733) );
  NAND U8677 ( .A(n6686), .B(creg[80]), .Z(n6732) );
  NAND U8678 ( .A(n6734), .B(n6735), .Z(c[7]) );
  NAND U8679 ( .A(n6691), .B(o[7]), .Z(n6735) );
  NAND U8680 ( .A(n6686), .B(creg[7]), .Z(n6734) );
  NAND U8681 ( .A(n6736), .B(n6737), .Z(c[79]) );
  NAND U8682 ( .A(n6691), .B(o[79]), .Z(n6737) );
  NAND U8683 ( .A(n6686), .B(creg[79]), .Z(n6736) );
  NAND U8684 ( .A(n6738), .B(n6739), .Z(c[78]) );
  NAND U8685 ( .A(n6691), .B(o[78]), .Z(n6739) );
  NAND U8686 ( .A(n6686), .B(creg[78]), .Z(n6738) );
  NAND U8687 ( .A(n6740), .B(n6741), .Z(c[77]) );
  NAND U8688 ( .A(n6691), .B(o[77]), .Z(n6741) );
  NAND U8689 ( .A(n6686), .B(creg[77]), .Z(n6740) );
  NAND U8690 ( .A(n6742), .B(n6743), .Z(c[76]) );
  NAND U8691 ( .A(n6691), .B(o[76]), .Z(n6743) );
  NAND U8692 ( .A(n6686), .B(creg[76]), .Z(n6742) );
  NAND U8693 ( .A(n6744), .B(n6745), .Z(c[75]) );
  NAND U8694 ( .A(n6691), .B(o[75]), .Z(n6745) );
  NAND U8695 ( .A(n6686), .B(creg[75]), .Z(n6744) );
  NAND U8696 ( .A(n6746), .B(n6747), .Z(c[74]) );
  NAND U8697 ( .A(n6691), .B(o[74]), .Z(n6747) );
  NAND U8698 ( .A(n6686), .B(creg[74]), .Z(n6746) );
  NAND U8699 ( .A(n6748), .B(n6749), .Z(c[73]) );
  NAND U8700 ( .A(n6691), .B(o[73]), .Z(n6749) );
  NAND U8701 ( .A(n6686), .B(creg[73]), .Z(n6748) );
  NAND U8702 ( .A(n6750), .B(n6751), .Z(c[72]) );
  NAND U8703 ( .A(n6691), .B(o[72]), .Z(n6751) );
  NAND U8704 ( .A(n6686), .B(creg[72]), .Z(n6750) );
  NAND U8705 ( .A(n6752), .B(n6753), .Z(c[71]) );
  NAND U8706 ( .A(n6691), .B(o[71]), .Z(n6753) );
  NAND U8707 ( .A(n6686), .B(creg[71]), .Z(n6752) );
  NAND U8708 ( .A(n6754), .B(n6755), .Z(c[70]) );
  NAND U8709 ( .A(n6691), .B(o[70]), .Z(n6755) );
  NAND U8710 ( .A(n6686), .B(creg[70]), .Z(n6754) );
  NAND U8711 ( .A(n6756), .B(n6757), .Z(c[6]) );
  NAND U8712 ( .A(n6691), .B(o[6]), .Z(n6757) );
  NAND U8713 ( .A(n6686), .B(creg[6]), .Z(n6756) );
  NAND U8714 ( .A(n6758), .B(n6759), .Z(c[69]) );
  NAND U8715 ( .A(n6691), .B(o[69]), .Z(n6759) );
  NAND U8716 ( .A(n6686), .B(creg[69]), .Z(n6758) );
  NAND U8717 ( .A(n6760), .B(n6761), .Z(c[68]) );
  NAND U8718 ( .A(n6691), .B(o[68]), .Z(n6761) );
  NAND U8719 ( .A(n6686), .B(creg[68]), .Z(n6760) );
  NAND U8720 ( .A(n6762), .B(n6763), .Z(c[67]) );
  NAND U8721 ( .A(n6691), .B(o[67]), .Z(n6763) );
  NAND U8722 ( .A(n6686), .B(creg[67]), .Z(n6762) );
  NAND U8723 ( .A(n6764), .B(n6765), .Z(c[66]) );
  NAND U8724 ( .A(n6691), .B(o[66]), .Z(n6765) );
  NAND U8725 ( .A(n6686), .B(creg[66]), .Z(n6764) );
  NAND U8726 ( .A(n6766), .B(n6767), .Z(c[65]) );
  NAND U8727 ( .A(n6691), .B(o[65]), .Z(n6767) );
  NAND U8728 ( .A(n6686), .B(creg[65]), .Z(n6766) );
  NAND U8729 ( .A(n6768), .B(n6769), .Z(c[64]) );
  NAND U8730 ( .A(n6691), .B(o[64]), .Z(n6769) );
  NAND U8731 ( .A(n6686), .B(creg[64]), .Z(n6768) );
  NAND U8732 ( .A(n6770), .B(n6771), .Z(c[63]) );
  NAND U8733 ( .A(n6691), .B(o[63]), .Z(n6771) );
  NAND U8734 ( .A(n6686), .B(creg[63]), .Z(n6770) );
  NAND U8735 ( .A(n6772), .B(n6773), .Z(c[62]) );
  NAND U8736 ( .A(n6691), .B(o[62]), .Z(n6773) );
  NAND U8737 ( .A(n6686), .B(creg[62]), .Z(n6772) );
  NAND U8738 ( .A(n6774), .B(n6775), .Z(c[61]) );
  NAND U8739 ( .A(n6691), .B(o[61]), .Z(n6775) );
  NAND U8740 ( .A(n6686), .B(creg[61]), .Z(n6774) );
  NAND U8741 ( .A(n6776), .B(n6777), .Z(c[60]) );
  NAND U8742 ( .A(n6691), .B(o[60]), .Z(n6777) );
  NAND U8743 ( .A(n6686), .B(creg[60]), .Z(n6776) );
  NAND U8744 ( .A(n6778), .B(n6779), .Z(c[5]) );
  NAND U8745 ( .A(n6691), .B(o[5]), .Z(n6779) );
  NAND U8746 ( .A(n6686), .B(creg[5]), .Z(n6778) );
  NAND U8747 ( .A(n6780), .B(n6781), .Z(c[59]) );
  NAND U8748 ( .A(n6691), .B(o[59]), .Z(n6781) );
  NAND U8749 ( .A(n6686), .B(creg[59]), .Z(n6780) );
  NAND U8750 ( .A(n6782), .B(n6783), .Z(c[58]) );
  NAND U8751 ( .A(n6691), .B(o[58]), .Z(n6783) );
  NAND U8752 ( .A(n6686), .B(creg[58]), .Z(n6782) );
  NAND U8753 ( .A(n6784), .B(n6785), .Z(c[57]) );
  NAND U8754 ( .A(n6691), .B(o[57]), .Z(n6785) );
  NAND U8755 ( .A(n6686), .B(creg[57]), .Z(n6784) );
  NAND U8756 ( .A(n6786), .B(n6787), .Z(c[56]) );
  NAND U8757 ( .A(n6691), .B(o[56]), .Z(n6787) );
  NAND U8758 ( .A(n6686), .B(creg[56]), .Z(n6786) );
  NAND U8759 ( .A(n6788), .B(n6789), .Z(c[55]) );
  NAND U8760 ( .A(n6691), .B(o[55]), .Z(n6789) );
  NAND U8761 ( .A(n6686), .B(creg[55]), .Z(n6788) );
  NAND U8762 ( .A(n6790), .B(n6791), .Z(c[54]) );
  NAND U8763 ( .A(n6691), .B(o[54]), .Z(n6791) );
  NAND U8764 ( .A(n6686), .B(creg[54]), .Z(n6790) );
  NAND U8765 ( .A(n6792), .B(n6793), .Z(c[53]) );
  NAND U8766 ( .A(n6691), .B(o[53]), .Z(n6793) );
  NAND U8767 ( .A(n6686), .B(creg[53]), .Z(n6792) );
  NAND U8768 ( .A(n6794), .B(n6795), .Z(c[52]) );
  NAND U8769 ( .A(n6691), .B(o[52]), .Z(n6795) );
  NAND U8770 ( .A(n6686), .B(creg[52]), .Z(n6794) );
  NAND U8771 ( .A(n6796), .B(n6797), .Z(c[51]) );
  NAND U8772 ( .A(n6691), .B(o[51]), .Z(n6797) );
  NAND U8773 ( .A(n6686), .B(creg[51]), .Z(n6796) );
  NAND U8774 ( .A(n6798), .B(n6799), .Z(c[50]) );
  NAND U8775 ( .A(n6691), .B(o[50]), .Z(n6799) );
  NAND U8776 ( .A(n6686), .B(creg[50]), .Z(n6798) );
  NAND U8777 ( .A(n6800), .B(n6801), .Z(c[4]) );
  NAND U8778 ( .A(n6691), .B(o[4]), .Z(n6801) );
  NAND U8779 ( .A(n6686), .B(creg[4]), .Z(n6800) );
  NAND U8780 ( .A(n6802), .B(n6803), .Z(c[49]) );
  NAND U8781 ( .A(n6691), .B(o[49]), .Z(n6803) );
  NAND U8782 ( .A(n6686), .B(creg[49]), .Z(n6802) );
  NAND U8783 ( .A(n6804), .B(n6805), .Z(c[48]) );
  NAND U8784 ( .A(n6691), .B(o[48]), .Z(n6805) );
  NAND U8785 ( .A(n6686), .B(creg[48]), .Z(n6804) );
  NAND U8786 ( .A(n6806), .B(n6807), .Z(c[47]) );
  NAND U8787 ( .A(n6691), .B(o[47]), .Z(n6807) );
  NAND U8788 ( .A(n6686), .B(creg[47]), .Z(n6806) );
  NAND U8789 ( .A(n6808), .B(n6809), .Z(c[46]) );
  NAND U8790 ( .A(n6691), .B(o[46]), .Z(n6809) );
  NAND U8791 ( .A(n6686), .B(creg[46]), .Z(n6808) );
  NAND U8792 ( .A(n6810), .B(n6811), .Z(c[45]) );
  NAND U8793 ( .A(n6691), .B(o[45]), .Z(n6811) );
  NAND U8794 ( .A(n6686), .B(creg[45]), .Z(n6810) );
  NAND U8795 ( .A(n6812), .B(n6813), .Z(c[44]) );
  NAND U8796 ( .A(n6691), .B(o[44]), .Z(n6813) );
  NAND U8797 ( .A(n6686), .B(creg[44]), .Z(n6812) );
  NAND U8798 ( .A(n6814), .B(n6815), .Z(c[43]) );
  NAND U8799 ( .A(n6691), .B(o[43]), .Z(n6815) );
  NAND U8800 ( .A(n6686), .B(creg[43]), .Z(n6814) );
  NAND U8801 ( .A(n6816), .B(n6817), .Z(c[42]) );
  NAND U8802 ( .A(n6691), .B(o[42]), .Z(n6817) );
  NAND U8803 ( .A(n6686), .B(creg[42]), .Z(n6816) );
  NAND U8804 ( .A(n6818), .B(n6819), .Z(c[41]) );
  NAND U8805 ( .A(n6691), .B(o[41]), .Z(n6819) );
  NAND U8806 ( .A(n6686), .B(creg[41]), .Z(n6818) );
  NAND U8807 ( .A(n6820), .B(n6821), .Z(c[40]) );
  NAND U8808 ( .A(n6691), .B(o[40]), .Z(n6821) );
  NAND U8809 ( .A(n6686), .B(creg[40]), .Z(n6820) );
  NAND U8810 ( .A(n6822), .B(n6823), .Z(c[3]) );
  NAND U8811 ( .A(n6691), .B(o[3]), .Z(n6823) );
  NAND U8812 ( .A(n6686), .B(creg[3]), .Z(n6822) );
  NAND U8813 ( .A(n6824), .B(n6825), .Z(c[39]) );
  NAND U8814 ( .A(n6691), .B(o[39]), .Z(n6825) );
  NAND U8815 ( .A(n6686), .B(creg[39]), .Z(n6824) );
  NAND U8816 ( .A(n6826), .B(n6827), .Z(c[38]) );
  NAND U8817 ( .A(n6691), .B(o[38]), .Z(n6827) );
  NAND U8818 ( .A(n6686), .B(creg[38]), .Z(n6826) );
  NAND U8819 ( .A(n6828), .B(n6829), .Z(c[37]) );
  NAND U8820 ( .A(n6691), .B(o[37]), .Z(n6829) );
  NAND U8821 ( .A(n6686), .B(creg[37]), .Z(n6828) );
  NAND U8822 ( .A(n6830), .B(n6831), .Z(c[36]) );
  NAND U8823 ( .A(n6691), .B(o[36]), .Z(n6831) );
  NAND U8824 ( .A(n6686), .B(creg[36]), .Z(n6830) );
  NAND U8825 ( .A(n6832), .B(n6833), .Z(c[35]) );
  NAND U8826 ( .A(n6691), .B(o[35]), .Z(n6833) );
  NAND U8827 ( .A(n6686), .B(creg[35]), .Z(n6832) );
  NAND U8828 ( .A(n6834), .B(n6835), .Z(c[34]) );
  NAND U8829 ( .A(n6691), .B(o[34]), .Z(n6835) );
  NAND U8830 ( .A(n6686), .B(creg[34]), .Z(n6834) );
  NAND U8831 ( .A(n6836), .B(n6837), .Z(c[33]) );
  NAND U8832 ( .A(n6691), .B(o[33]), .Z(n6837) );
  NAND U8833 ( .A(n6686), .B(creg[33]), .Z(n6836) );
  NAND U8834 ( .A(n6838), .B(n6839), .Z(c[32]) );
  NAND U8835 ( .A(n6691), .B(o[32]), .Z(n6839) );
  NAND U8836 ( .A(n6686), .B(creg[32]), .Z(n6838) );
  NAND U8837 ( .A(n6840), .B(n6841), .Z(c[31]) );
  NAND U8838 ( .A(n6691), .B(o[31]), .Z(n6841) );
  NAND U8839 ( .A(n6686), .B(creg[31]), .Z(n6840) );
  NAND U8840 ( .A(n6842), .B(n6843), .Z(c[30]) );
  NAND U8841 ( .A(n6691), .B(o[30]), .Z(n6843) );
  NAND U8842 ( .A(n6686), .B(creg[30]), .Z(n6842) );
  NAND U8843 ( .A(n6844), .B(n6845), .Z(c[2]) );
  NAND U8844 ( .A(n6691), .B(o[2]), .Z(n6845) );
  NAND U8845 ( .A(n6686), .B(creg[2]), .Z(n6844) );
  NAND U8846 ( .A(n6846), .B(n6847), .Z(c[29]) );
  NAND U8847 ( .A(n6691), .B(o[29]), .Z(n6847) );
  NAND U8848 ( .A(n6686), .B(creg[29]), .Z(n6846) );
  NAND U8849 ( .A(n6848), .B(n6849), .Z(c[28]) );
  NAND U8850 ( .A(n6691), .B(o[28]), .Z(n6849) );
  NAND U8851 ( .A(n6686), .B(creg[28]), .Z(n6848) );
  NAND U8852 ( .A(n6850), .B(n6851), .Z(c[27]) );
  NAND U8853 ( .A(n6691), .B(o[27]), .Z(n6851) );
  NAND U8854 ( .A(n6686), .B(creg[27]), .Z(n6850) );
  NAND U8855 ( .A(n6852), .B(n6853), .Z(c[26]) );
  NAND U8856 ( .A(n6691), .B(o[26]), .Z(n6853) );
  NAND U8857 ( .A(n6686), .B(creg[26]), .Z(n6852) );
  NAND U8858 ( .A(n6854), .B(n6855), .Z(c[25]) );
  NAND U8859 ( .A(n6691), .B(o[25]), .Z(n6855) );
  NAND U8860 ( .A(n6686), .B(creg[25]), .Z(n6854) );
  NAND U8861 ( .A(n6856), .B(n6857), .Z(c[255]) );
  NAND U8862 ( .A(n6691), .B(o[255]), .Z(n6857) );
  NAND U8863 ( .A(n6686), .B(creg[255]), .Z(n6856) );
  NAND U8864 ( .A(n6858), .B(n6859), .Z(c[254]) );
  NAND U8865 ( .A(n6691), .B(o[254]), .Z(n6859) );
  NAND U8866 ( .A(n6686), .B(creg[254]), .Z(n6858) );
  NAND U8867 ( .A(n6860), .B(n6861), .Z(c[253]) );
  NAND U8868 ( .A(n6691), .B(o[253]), .Z(n6861) );
  NAND U8869 ( .A(n6686), .B(creg[253]), .Z(n6860) );
  NAND U8870 ( .A(n6862), .B(n6863), .Z(c[252]) );
  NAND U8871 ( .A(n6691), .B(o[252]), .Z(n6863) );
  NAND U8872 ( .A(n6686), .B(creg[252]), .Z(n6862) );
  NAND U8873 ( .A(n6864), .B(n6865), .Z(c[251]) );
  NAND U8874 ( .A(n6691), .B(o[251]), .Z(n6865) );
  NAND U8875 ( .A(n6686), .B(creg[251]), .Z(n6864) );
  NAND U8876 ( .A(n6866), .B(n6867), .Z(c[250]) );
  NAND U8877 ( .A(n6691), .B(o[250]), .Z(n6867) );
  NAND U8878 ( .A(n6686), .B(creg[250]), .Z(n6866) );
  NAND U8879 ( .A(n6868), .B(n6869), .Z(c[24]) );
  NAND U8880 ( .A(n6691), .B(o[24]), .Z(n6869) );
  NAND U8881 ( .A(n6686), .B(creg[24]), .Z(n6868) );
  NAND U8882 ( .A(n6870), .B(n6871), .Z(c[249]) );
  NAND U8883 ( .A(n6691), .B(o[249]), .Z(n6871) );
  NAND U8884 ( .A(n6686), .B(creg[249]), .Z(n6870) );
  NAND U8885 ( .A(n6872), .B(n6873), .Z(c[248]) );
  NAND U8886 ( .A(n6691), .B(o[248]), .Z(n6873) );
  NAND U8887 ( .A(n6686), .B(creg[248]), .Z(n6872) );
  NAND U8888 ( .A(n6874), .B(n6875), .Z(c[247]) );
  NAND U8889 ( .A(n6691), .B(o[247]), .Z(n6875) );
  NAND U8890 ( .A(n6686), .B(creg[247]), .Z(n6874) );
  NAND U8891 ( .A(n6876), .B(n6877), .Z(c[246]) );
  NAND U8892 ( .A(n6691), .B(o[246]), .Z(n6877) );
  NAND U8893 ( .A(n6686), .B(creg[246]), .Z(n6876) );
  NAND U8894 ( .A(n6878), .B(n6879), .Z(c[245]) );
  NAND U8895 ( .A(n6691), .B(o[245]), .Z(n6879) );
  NAND U8896 ( .A(n6686), .B(creg[245]), .Z(n6878) );
  NAND U8897 ( .A(n6880), .B(n6881), .Z(c[244]) );
  NAND U8898 ( .A(n6691), .B(o[244]), .Z(n6881) );
  NAND U8899 ( .A(n6686), .B(creg[244]), .Z(n6880) );
  NAND U8900 ( .A(n6882), .B(n6883), .Z(c[243]) );
  NAND U8901 ( .A(n6691), .B(o[243]), .Z(n6883) );
  NAND U8902 ( .A(n6686), .B(creg[243]), .Z(n6882) );
  NAND U8903 ( .A(n6884), .B(n6885), .Z(c[242]) );
  NAND U8904 ( .A(n6691), .B(o[242]), .Z(n6885) );
  NAND U8905 ( .A(n6686), .B(creg[242]), .Z(n6884) );
  NAND U8906 ( .A(n6886), .B(n6887), .Z(c[241]) );
  NAND U8907 ( .A(n6691), .B(o[241]), .Z(n6887) );
  NAND U8908 ( .A(n6686), .B(creg[241]), .Z(n6886) );
  NAND U8909 ( .A(n6888), .B(n6889), .Z(c[240]) );
  NAND U8910 ( .A(n6691), .B(o[240]), .Z(n6889) );
  NAND U8911 ( .A(n6686), .B(creg[240]), .Z(n6888) );
  NAND U8912 ( .A(n6890), .B(n6891), .Z(c[23]) );
  NAND U8913 ( .A(n6691), .B(o[23]), .Z(n6891) );
  NAND U8914 ( .A(n6686), .B(creg[23]), .Z(n6890) );
  NAND U8915 ( .A(n6892), .B(n6893), .Z(c[239]) );
  NAND U8916 ( .A(n6691), .B(o[239]), .Z(n6893) );
  NAND U8917 ( .A(n6686), .B(creg[239]), .Z(n6892) );
  NAND U8918 ( .A(n6894), .B(n6895), .Z(c[238]) );
  NAND U8919 ( .A(n6691), .B(o[238]), .Z(n6895) );
  NAND U8920 ( .A(n6686), .B(creg[238]), .Z(n6894) );
  NAND U8921 ( .A(n6896), .B(n6897), .Z(c[237]) );
  NAND U8922 ( .A(n6691), .B(o[237]), .Z(n6897) );
  NAND U8923 ( .A(n6686), .B(creg[237]), .Z(n6896) );
  NAND U8924 ( .A(n6898), .B(n6899), .Z(c[236]) );
  NAND U8925 ( .A(n6691), .B(o[236]), .Z(n6899) );
  NAND U8926 ( .A(n6686), .B(creg[236]), .Z(n6898) );
  NAND U8927 ( .A(n6900), .B(n6901), .Z(c[235]) );
  NAND U8928 ( .A(n6691), .B(o[235]), .Z(n6901) );
  NAND U8929 ( .A(n6686), .B(creg[235]), .Z(n6900) );
  NAND U8930 ( .A(n6902), .B(n6903), .Z(c[234]) );
  NAND U8931 ( .A(n6691), .B(o[234]), .Z(n6903) );
  NAND U8932 ( .A(n6686), .B(creg[234]), .Z(n6902) );
  NAND U8933 ( .A(n6904), .B(n6905), .Z(c[233]) );
  NAND U8934 ( .A(n6691), .B(o[233]), .Z(n6905) );
  NAND U8935 ( .A(n6686), .B(creg[233]), .Z(n6904) );
  NAND U8936 ( .A(n6906), .B(n6907), .Z(c[232]) );
  NAND U8937 ( .A(n6691), .B(o[232]), .Z(n6907) );
  NAND U8938 ( .A(n6686), .B(creg[232]), .Z(n6906) );
  NAND U8939 ( .A(n6908), .B(n6909), .Z(c[231]) );
  NAND U8940 ( .A(n6691), .B(o[231]), .Z(n6909) );
  NAND U8941 ( .A(n6686), .B(creg[231]), .Z(n6908) );
  NAND U8942 ( .A(n6910), .B(n6911), .Z(c[230]) );
  NAND U8943 ( .A(n6691), .B(o[230]), .Z(n6911) );
  NAND U8944 ( .A(n6686), .B(creg[230]), .Z(n6910) );
  NAND U8945 ( .A(n6912), .B(n6913), .Z(c[22]) );
  NAND U8946 ( .A(n6691), .B(o[22]), .Z(n6913) );
  NAND U8947 ( .A(n6686), .B(creg[22]), .Z(n6912) );
  NAND U8948 ( .A(n6914), .B(n6915), .Z(c[229]) );
  NAND U8949 ( .A(n6691), .B(o[229]), .Z(n6915) );
  NAND U8950 ( .A(n6686), .B(creg[229]), .Z(n6914) );
  NAND U8951 ( .A(n6916), .B(n6917), .Z(c[228]) );
  NAND U8952 ( .A(n6691), .B(o[228]), .Z(n6917) );
  NAND U8953 ( .A(n6686), .B(creg[228]), .Z(n6916) );
  NAND U8954 ( .A(n6918), .B(n6919), .Z(c[227]) );
  NAND U8955 ( .A(n6691), .B(o[227]), .Z(n6919) );
  NAND U8956 ( .A(n6686), .B(creg[227]), .Z(n6918) );
  NAND U8957 ( .A(n6920), .B(n6921), .Z(c[226]) );
  NAND U8958 ( .A(n6691), .B(o[226]), .Z(n6921) );
  NAND U8959 ( .A(n6686), .B(creg[226]), .Z(n6920) );
  NAND U8960 ( .A(n6922), .B(n6923), .Z(c[225]) );
  NAND U8961 ( .A(n6691), .B(o[225]), .Z(n6923) );
  NAND U8962 ( .A(n6686), .B(creg[225]), .Z(n6922) );
  NAND U8963 ( .A(n6924), .B(n6925), .Z(c[224]) );
  NAND U8964 ( .A(n6691), .B(o[224]), .Z(n6925) );
  NAND U8965 ( .A(n6686), .B(creg[224]), .Z(n6924) );
  NAND U8966 ( .A(n6926), .B(n6927), .Z(c[223]) );
  NAND U8967 ( .A(n6691), .B(o[223]), .Z(n6927) );
  NAND U8968 ( .A(n6686), .B(creg[223]), .Z(n6926) );
  NAND U8969 ( .A(n6928), .B(n6929), .Z(c[222]) );
  NAND U8970 ( .A(n6691), .B(o[222]), .Z(n6929) );
  NAND U8971 ( .A(n6686), .B(creg[222]), .Z(n6928) );
  NAND U8972 ( .A(n6930), .B(n6931), .Z(c[221]) );
  NAND U8973 ( .A(n6691), .B(o[221]), .Z(n6931) );
  NAND U8974 ( .A(n6686), .B(creg[221]), .Z(n6930) );
  NAND U8975 ( .A(n6932), .B(n6933), .Z(c[220]) );
  NAND U8976 ( .A(n6691), .B(o[220]), .Z(n6933) );
  NAND U8977 ( .A(n6686), .B(creg[220]), .Z(n6932) );
  NAND U8978 ( .A(n6934), .B(n6935), .Z(c[21]) );
  NAND U8979 ( .A(n6691), .B(o[21]), .Z(n6935) );
  NAND U8980 ( .A(n6686), .B(creg[21]), .Z(n6934) );
  NAND U8981 ( .A(n6936), .B(n6937), .Z(c[219]) );
  NAND U8982 ( .A(n6691), .B(o[219]), .Z(n6937) );
  NAND U8983 ( .A(n6686), .B(creg[219]), .Z(n6936) );
  NAND U8984 ( .A(n6938), .B(n6939), .Z(c[218]) );
  NAND U8985 ( .A(n6691), .B(o[218]), .Z(n6939) );
  NAND U8986 ( .A(n6686), .B(creg[218]), .Z(n6938) );
  NAND U8987 ( .A(n6940), .B(n6941), .Z(c[217]) );
  NAND U8988 ( .A(n6691), .B(o[217]), .Z(n6941) );
  NAND U8989 ( .A(n6686), .B(creg[217]), .Z(n6940) );
  NAND U8990 ( .A(n6942), .B(n6943), .Z(c[216]) );
  NAND U8991 ( .A(n6691), .B(o[216]), .Z(n6943) );
  NAND U8992 ( .A(n6686), .B(creg[216]), .Z(n6942) );
  NAND U8993 ( .A(n6944), .B(n6945), .Z(c[215]) );
  NAND U8994 ( .A(n6691), .B(o[215]), .Z(n6945) );
  NAND U8995 ( .A(n6686), .B(creg[215]), .Z(n6944) );
  NAND U8996 ( .A(n6946), .B(n6947), .Z(c[214]) );
  NAND U8997 ( .A(n6691), .B(o[214]), .Z(n6947) );
  NAND U8998 ( .A(n6686), .B(creg[214]), .Z(n6946) );
  NAND U8999 ( .A(n6948), .B(n6949), .Z(c[213]) );
  NAND U9000 ( .A(n6691), .B(o[213]), .Z(n6949) );
  NAND U9001 ( .A(n6686), .B(creg[213]), .Z(n6948) );
  NAND U9002 ( .A(n6950), .B(n6951), .Z(c[212]) );
  NAND U9003 ( .A(n6691), .B(o[212]), .Z(n6951) );
  NAND U9004 ( .A(n6686), .B(creg[212]), .Z(n6950) );
  NAND U9005 ( .A(n6952), .B(n6953), .Z(c[211]) );
  NAND U9006 ( .A(n6691), .B(o[211]), .Z(n6953) );
  NAND U9007 ( .A(n6686), .B(creg[211]), .Z(n6952) );
  NAND U9008 ( .A(n6954), .B(n6955), .Z(c[210]) );
  NAND U9009 ( .A(n6691), .B(o[210]), .Z(n6955) );
  NAND U9010 ( .A(n6686), .B(creg[210]), .Z(n6954) );
  NAND U9011 ( .A(n6956), .B(n6957), .Z(c[20]) );
  NAND U9012 ( .A(n6691), .B(o[20]), .Z(n6957) );
  NAND U9013 ( .A(n6686), .B(creg[20]), .Z(n6956) );
  NAND U9014 ( .A(n6958), .B(n6959), .Z(c[209]) );
  NAND U9015 ( .A(n6691), .B(o[209]), .Z(n6959) );
  NAND U9016 ( .A(n6686), .B(creg[209]), .Z(n6958) );
  NAND U9017 ( .A(n6960), .B(n6961), .Z(c[208]) );
  NAND U9018 ( .A(n6691), .B(o[208]), .Z(n6961) );
  NAND U9019 ( .A(n6686), .B(creg[208]), .Z(n6960) );
  NAND U9020 ( .A(n6962), .B(n6963), .Z(c[207]) );
  NAND U9021 ( .A(n6691), .B(o[207]), .Z(n6963) );
  NAND U9022 ( .A(n6686), .B(creg[207]), .Z(n6962) );
  NAND U9023 ( .A(n6964), .B(n6965), .Z(c[206]) );
  NAND U9024 ( .A(n6691), .B(o[206]), .Z(n6965) );
  NAND U9025 ( .A(n6686), .B(creg[206]), .Z(n6964) );
  NAND U9026 ( .A(n6966), .B(n6967), .Z(c[205]) );
  NAND U9027 ( .A(n6691), .B(o[205]), .Z(n6967) );
  NAND U9028 ( .A(n6686), .B(creg[205]), .Z(n6966) );
  NAND U9029 ( .A(n6968), .B(n6969), .Z(c[204]) );
  NAND U9030 ( .A(n6691), .B(o[204]), .Z(n6969) );
  NAND U9031 ( .A(n6686), .B(creg[204]), .Z(n6968) );
  NAND U9032 ( .A(n6970), .B(n6971), .Z(c[203]) );
  NAND U9033 ( .A(n6691), .B(o[203]), .Z(n6971) );
  NAND U9034 ( .A(n6686), .B(creg[203]), .Z(n6970) );
  NAND U9035 ( .A(n6972), .B(n6973), .Z(c[202]) );
  NAND U9036 ( .A(n6691), .B(o[202]), .Z(n6973) );
  NAND U9037 ( .A(n6686), .B(creg[202]), .Z(n6972) );
  NAND U9038 ( .A(n6974), .B(n6975), .Z(c[201]) );
  NAND U9039 ( .A(n6691), .B(o[201]), .Z(n6975) );
  NAND U9040 ( .A(n6686), .B(creg[201]), .Z(n6974) );
  NAND U9041 ( .A(n6976), .B(n6977), .Z(c[200]) );
  NAND U9042 ( .A(n6691), .B(o[200]), .Z(n6977) );
  NAND U9043 ( .A(n6686), .B(creg[200]), .Z(n6976) );
  NAND U9044 ( .A(n6978), .B(n6979), .Z(c[1]) );
  NAND U9045 ( .A(n6691), .B(o[1]), .Z(n6979) );
  NAND U9046 ( .A(n6686), .B(creg[1]), .Z(n6978) );
  NAND U9047 ( .A(n6980), .B(n6981), .Z(c[19]) );
  NAND U9048 ( .A(n6691), .B(o[19]), .Z(n6981) );
  NAND U9049 ( .A(n6686), .B(creg[19]), .Z(n6980) );
  NAND U9050 ( .A(n6982), .B(n6983), .Z(c[199]) );
  NAND U9051 ( .A(n6691), .B(o[199]), .Z(n6983) );
  NAND U9052 ( .A(n6686), .B(creg[199]), .Z(n6982) );
  NAND U9053 ( .A(n6984), .B(n6985), .Z(c[198]) );
  NAND U9054 ( .A(n6691), .B(o[198]), .Z(n6985) );
  NAND U9055 ( .A(n6686), .B(creg[198]), .Z(n6984) );
  NAND U9056 ( .A(n6986), .B(n6987), .Z(c[197]) );
  NAND U9057 ( .A(n6691), .B(o[197]), .Z(n6987) );
  NAND U9058 ( .A(n6686), .B(creg[197]), .Z(n6986) );
  NAND U9059 ( .A(n6988), .B(n6989), .Z(c[196]) );
  NAND U9060 ( .A(n6691), .B(o[196]), .Z(n6989) );
  NAND U9061 ( .A(n6686), .B(creg[196]), .Z(n6988) );
  NAND U9062 ( .A(n6990), .B(n6991), .Z(c[195]) );
  NAND U9063 ( .A(n6691), .B(o[195]), .Z(n6991) );
  NAND U9064 ( .A(n6686), .B(creg[195]), .Z(n6990) );
  NAND U9065 ( .A(n6992), .B(n6993), .Z(c[194]) );
  NAND U9066 ( .A(n6691), .B(o[194]), .Z(n6993) );
  NAND U9067 ( .A(n6686), .B(creg[194]), .Z(n6992) );
  NAND U9068 ( .A(n6994), .B(n6995), .Z(c[193]) );
  NAND U9069 ( .A(n6691), .B(o[193]), .Z(n6995) );
  NAND U9070 ( .A(n6686), .B(creg[193]), .Z(n6994) );
  NAND U9071 ( .A(n6996), .B(n6997), .Z(c[192]) );
  NAND U9072 ( .A(n6691), .B(o[192]), .Z(n6997) );
  NAND U9073 ( .A(n6686), .B(creg[192]), .Z(n6996) );
  NAND U9074 ( .A(n6998), .B(n6999), .Z(c[191]) );
  NAND U9075 ( .A(n6691), .B(o[191]), .Z(n6999) );
  NAND U9076 ( .A(n6686), .B(creg[191]), .Z(n6998) );
  NAND U9077 ( .A(n7000), .B(n7001), .Z(c[190]) );
  NAND U9078 ( .A(n6691), .B(o[190]), .Z(n7001) );
  NAND U9079 ( .A(n6686), .B(creg[190]), .Z(n7000) );
  NAND U9080 ( .A(n7002), .B(n7003), .Z(c[18]) );
  NAND U9081 ( .A(n6691), .B(o[18]), .Z(n7003) );
  NAND U9082 ( .A(n6686), .B(creg[18]), .Z(n7002) );
  NAND U9083 ( .A(n7004), .B(n7005), .Z(c[189]) );
  NAND U9084 ( .A(n6691), .B(o[189]), .Z(n7005) );
  NAND U9085 ( .A(n6686), .B(creg[189]), .Z(n7004) );
  NAND U9086 ( .A(n7006), .B(n7007), .Z(c[188]) );
  NAND U9087 ( .A(n6691), .B(o[188]), .Z(n7007) );
  NAND U9088 ( .A(n6686), .B(creg[188]), .Z(n7006) );
  NAND U9089 ( .A(n7008), .B(n7009), .Z(c[187]) );
  NAND U9090 ( .A(n6691), .B(o[187]), .Z(n7009) );
  NAND U9091 ( .A(n6686), .B(creg[187]), .Z(n7008) );
  NAND U9092 ( .A(n7010), .B(n7011), .Z(c[186]) );
  NAND U9093 ( .A(n6691), .B(o[186]), .Z(n7011) );
  NAND U9094 ( .A(n6686), .B(creg[186]), .Z(n7010) );
  NAND U9095 ( .A(n7012), .B(n7013), .Z(c[185]) );
  NAND U9096 ( .A(n6691), .B(o[185]), .Z(n7013) );
  NAND U9097 ( .A(n6686), .B(creg[185]), .Z(n7012) );
  NAND U9098 ( .A(n7014), .B(n7015), .Z(c[184]) );
  NAND U9099 ( .A(n6691), .B(o[184]), .Z(n7015) );
  NAND U9100 ( .A(n6686), .B(creg[184]), .Z(n7014) );
  NAND U9101 ( .A(n7016), .B(n7017), .Z(c[183]) );
  NAND U9102 ( .A(n6691), .B(o[183]), .Z(n7017) );
  NAND U9103 ( .A(n6686), .B(creg[183]), .Z(n7016) );
  NAND U9104 ( .A(n7018), .B(n7019), .Z(c[182]) );
  NAND U9105 ( .A(n6691), .B(o[182]), .Z(n7019) );
  NAND U9106 ( .A(n6686), .B(creg[182]), .Z(n7018) );
  NAND U9107 ( .A(n7020), .B(n7021), .Z(c[181]) );
  NAND U9108 ( .A(n6691), .B(o[181]), .Z(n7021) );
  NAND U9109 ( .A(n6686), .B(creg[181]), .Z(n7020) );
  NAND U9110 ( .A(n7022), .B(n7023), .Z(c[180]) );
  NAND U9111 ( .A(n6691), .B(o[180]), .Z(n7023) );
  NAND U9112 ( .A(n6686), .B(creg[180]), .Z(n7022) );
  NAND U9113 ( .A(n7024), .B(n7025), .Z(c[17]) );
  NAND U9114 ( .A(n6691), .B(o[17]), .Z(n7025) );
  NAND U9115 ( .A(n6686), .B(creg[17]), .Z(n7024) );
  NAND U9116 ( .A(n7026), .B(n7027), .Z(c[179]) );
  NAND U9117 ( .A(n6691), .B(o[179]), .Z(n7027) );
  NAND U9118 ( .A(n6686), .B(creg[179]), .Z(n7026) );
  NAND U9119 ( .A(n7028), .B(n7029), .Z(c[178]) );
  NAND U9120 ( .A(n6691), .B(o[178]), .Z(n7029) );
  NAND U9121 ( .A(n6686), .B(creg[178]), .Z(n7028) );
  NAND U9122 ( .A(n7030), .B(n7031), .Z(c[177]) );
  NAND U9123 ( .A(n6691), .B(o[177]), .Z(n7031) );
  NAND U9124 ( .A(n6686), .B(creg[177]), .Z(n7030) );
  NAND U9125 ( .A(n7032), .B(n7033), .Z(c[176]) );
  NAND U9126 ( .A(n6691), .B(o[176]), .Z(n7033) );
  NAND U9127 ( .A(n6686), .B(creg[176]), .Z(n7032) );
  NAND U9128 ( .A(n7034), .B(n7035), .Z(c[175]) );
  NAND U9129 ( .A(n6691), .B(o[175]), .Z(n7035) );
  NAND U9130 ( .A(n6686), .B(creg[175]), .Z(n7034) );
  NAND U9131 ( .A(n7036), .B(n7037), .Z(c[174]) );
  NAND U9132 ( .A(n6691), .B(o[174]), .Z(n7037) );
  NAND U9133 ( .A(n6686), .B(creg[174]), .Z(n7036) );
  NAND U9134 ( .A(n7038), .B(n7039), .Z(c[173]) );
  NAND U9135 ( .A(n6691), .B(o[173]), .Z(n7039) );
  NAND U9136 ( .A(n6686), .B(creg[173]), .Z(n7038) );
  NAND U9137 ( .A(n7040), .B(n7041), .Z(c[172]) );
  NAND U9138 ( .A(n6691), .B(o[172]), .Z(n7041) );
  NAND U9139 ( .A(n6686), .B(creg[172]), .Z(n7040) );
  NAND U9140 ( .A(n7042), .B(n7043), .Z(c[171]) );
  NAND U9141 ( .A(n6691), .B(o[171]), .Z(n7043) );
  NAND U9142 ( .A(n6686), .B(creg[171]), .Z(n7042) );
  NAND U9143 ( .A(n7044), .B(n7045), .Z(c[170]) );
  NAND U9144 ( .A(n6691), .B(o[170]), .Z(n7045) );
  NAND U9145 ( .A(n6686), .B(creg[170]), .Z(n7044) );
  NAND U9146 ( .A(n7046), .B(n7047), .Z(c[16]) );
  NAND U9147 ( .A(n6691), .B(o[16]), .Z(n7047) );
  NAND U9148 ( .A(n6686), .B(creg[16]), .Z(n7046) );
  NAND U9149 ( .A(n7048), .B(n7049), .Z(c[169]) );
  NAND U9150 ( .A(n6691), .B(o[169]), .Z(n7049) );
  NAND U9151 ( .A(n6686), .B(creg[169]), .Z(n7048) );
  NAND U9152 ( .A(n7050), .B(n7051), .Z(c[168]) );
  NAND U9153 ( .A(n6691), .B(o[168]), .Z(n7051) );
  NAND U9154 ( .A(n6686), .B(creg[168]), .Z(n7050) );
  NAND U9155 ( .A(n7052), .B(n7053), .Z(c[167]) );
  NAND U9156 ( .A(n6691), .B(o[167]), .Z(n7053) );
  NAND U9157 ( .A(n6686), .B(creg[167]), .Z(n7052) );
  NAND U9158 ( .A(n7054), .B(n7055), .Z(c[166]) );
  NAND U9159 ( .A(n6691), .B(o[166]), .Z(n7055) );
  NAND U9160 ( .A(n6686), .B(creg[166]), .Z(n7054) );
  NAND U9161 ( .A(n7056), .B(n7057), .Z(c[165]) );
  NAND U9162 ( .A(n6691), .B(o[165]), .Z(n7057) );
  NAND U9163 ( .A(n6686), .B(creg[165]), .Z(n7056) );
  NAND U9164 ( .A(n7058), .B(n7059), .Z(c[164]) );
  NAND U9165 ( .A(n6691), .B(o[164]), .Z(n7059) );
  NAND U9166 ( .A(n6686), .B(creg[164]), .Z(n7058) );
  NAND U9167 ( .A(n7060), .B(n7061), .Z(c[163]) );
  NAND U9168 ( .A(n6691), .B(o[163]), .Z(n7061) );
  NAND U9169 ( .A(n6686), .B(creg[163]), .Z(n7060) );
  NAND U9170 ( .A(n7062), .B(n7063), .Z(c[162]) );
  NAND U9171 ( .A(n6691), .B(o[162]), .Z(n7063) );
  NAND U9172 ( .A(n6686), .B(creg[162]), .Z(n7062) );
  NAND U9173 ( .A(n7064), .B(n7065), .Z(c[161]) );
  NAND U9174 ( .A(n6691), .B(o[161]), .Z(n7065) );
  NAND U9175 ( .A(n6686), .B(creg[161]), .Z(n7064) );
  NAND U9176 ( .A(n7066), .B(n7067), .Z(c[160]) );
  NAND U9177 ( .A(n6691), .B(o[160]), .Z(n7067) );
  NAND U9178 ( .A(n6686), .B(creg[160]), .Z(n7066) );
  NAND U9179 ( .A(n7068), .B(n7069), .Z(c[15]) );
  NAND U9180 ( .A(n6691), .B(o[15]), .Z(n7069) );
  NAND U9181 ( .A(n6686), .B(creg[15]), .Z(n7068) );
  NAND U9182 ( .A(n7070), .B(n7071), .Z(c[159]) );
  NAND U9183 ( .A(n6691), .B(o[159]), .Z(n7071) );
  NAND U9184 ( .A(n6686), .B(creg[159]), .Z(n7070) );
  NAND U9185 ( .A(n7072), .B(n7073), .Z(c[158]) );
  NAND U9186 ( .A(n6691), .B(o[158]), .Z(n7073) );
  NAND U9187 ( .A(n6686), .B(creg[158]), .Z(n7072) );
  NAND U9188 ( .A(n7074), .B(n7075), .Z(c[157]) );
  NAND U9189 ( .A(n6691), .B(o[157]), .Z(n7075) );
  NAND U9190 ( .A(n6686), .B(creg[157]), .Z(n7074) );
  NAND U9191 ( .A(n7076), .B(n7077), .Z(c[156]) );
  NAND U9192 ( .A(n6691), .B(o[156]), .Z(n7077) );
  NAND U9193 ( .A(n6686), .B(creg[156]), .Z(n7076) );
  NAND U9194 ( .A(n7078), .B(n7079), .Z(c[155]) );
  NAND U9195 ( .A(n6691), .B(o[155]), .Z(n7079) );
  NAND U9196 ( .A(n6686), .B(creg[155]), .Z(n7078) );
  NAND U9197 ( .A(n7080), .B(n7081), .Z(c[154]) );
  NAND U9198 ( .A(n6691), .B(o[154]), .Z(n7081) );
  NAND U9199 ( .A(n6686), .B(creg[154]), .Z(n7080) );
  NAND U9200 ( .A(n7082), .B(n7083), .Z(c[153]) );
  NAND U9201 ( .A(n6691), .B(o[153]), .Z(n7083) );
  NAND U9202 ( .A(n6686), .B(creg[153]), .Z(n7082) );
  NAND U9203 ( .A(n7084), .B(n7085), .Z(c[152]) );
  NAND U9204 ( .A(n6691), .B(o[152]), .Z(n7085) );
  NAND U9205 ( .A(n6686), .B(creg[152]), .Z(n7084) );
  NAND U9206 ( .A(n7086), .B(n7087), .Z(c[151]) );
  NAND U9207 ( .A(n6691), .B(o[151]), .Z(n7087) );
  NAND U9208 ( .A(n6686), .B(creg[151]), .Z(n7086) );
  NAND U9209 ( .A(n7088), .B(n7089), .Z(c[150]) );
  NAND U9210 ( .A(n6691), .B(o[150]), .Z(n7089) );
  NAND U9211 ( .A(n6686), .B(creg[150]), .Z(n7088) );
  NAND U9212 ( .A(n7090), .B(n7091), .Z(c[14]) );
  NAND U9213 ( .A(n6691), .B(o[14]), .Z(n7091) );
  NAND U9214 ( .A(n6686), .B(creg[14]), .Z(n7090) );
  NAND U9215 ( .A(n7092), .B(n7093), .Z(c[149]) );
  NAND U9216 ( .A(n6691), .B(o[149]), .Z(n7093) );
  NAND U9217 ( .A(n6686), .B(creg[149]), .Z(n7092) );
  NAND U9218 ( .A(n7094), .B(n7095), .Z(c[148]) );
  NAND U9219 ( .A(n6691), .B(o[148]), .Z(n7095) );
  NAND U9220 ( .A(n6686), .B(creg[148]), .Z(n7094) );
  NAND U9221 ( .A(n7096), .B(n7097), .Z(c[147]) );
  NAND U9222 ( .A(n6691), .B(o[147]), .Z(n7097) );
  NAND U9223 ( .A(n6686), .B(creg[147]), .Z(n7096) );
  NAND U9224 ( .A(n7098), .B(n7099), .Z(c[146]) );
  NAND U9225 ( .A(n6691), .B(o[146]), .Z(n7099) );
  NAND U9226 ( .A(n6686), .B(creg[146]), .Z(n7098) );
  NAND U9227 ( .A(n7100), .B(n7101), .Z(c[145]) );
  NAND U9228 ( .A(n6691), .B(o[145]), .Z(n7101) );
  NAND U9229 ( .A(n6686), .B(creg[145]), .Z(n7100) );
  NAND U9230 ( .A(n7102), .B(n7103), .Z(c[144]) );
  NAND U9231 ( .A(n6691), .B(o[144]), .Z(n7103) );
  NAND U9232 ( .A(n6686), .B(creg[144]), .Z(n7102) );
  NAND U9233 ( .A(n7104), .B(n7105), .Z(c[143]) );
  NAND U9234 ( .A(n6691), .B(o[143]), .Z(n7105) );
  NAND U9235 ( .A(n6686), .B(creg[143]), .Z(n7104) );
  NAND U9236 ( .A(n7106), .B(n7107), .Z(c[142]) );
  NAND U9237 ( .A(n6691), .B(o[142]), .Z(n7107) );
  NAND U9238 ( .A(n6686), .B(creg[142]), .Z(n7106) );
  NAND U9239 ( .A(n7108), .B(n7109), .Z(c[141]) );
  NAND U9240 ( .A(n6691), .B(o[141]), .Z(n7109) );
  NAND U9241 ( .A(n6686), .B(creg[141]), .Z(n7108) );
  NAND U9242 ( .A(n7110), .B(n7111), .Z(c[140]) );
  NAND U9243 ( .A(n6691), .B(o[140]), .Z(n7111) );
  NAND U9244 ( .A(n6686), .B(creg[140]), .Z(n7110) );
  NAND U9245 ( .A(n7112), .B(n7113), .Z(c[13]) );
  NAND U9246 ( .A(n6691), .B(o[13]), .Z(n7113) );
  NAND U9247 ( .A(n6686), .B(creg[13]), .Z(n7112) );
  NAND U9248 ( .A(n7114), .B(n7115), .Z(c[139]) );
  NAND U9249 ( .A(n6691), .B(o[139]), .Z(n7115) );
  NAND U9250 ( .A(n6686), .B(creg[139]), .Z(n7114) );
  NAND U9251 ( .A(n7116), .B(n7117), .Z(c[138]) );
  NAND U9252 ( .A(n6691), .B(o[138]), .Z(n7117) );
  NAND U9253 ( .A(n6686), .B(creg[138]), .Z(n7116) );
  NAND U9254 ( .A(n7118), .B(n7119), .Z(c[137]) );
  NAND U9255 ( .A(n6691), .B(o[137]), .Z(n7119) );
  NAND U9256 ( .A(n6686), .B(creg[137]), .Z(n7118) );
  NAND U9257 ( .A(n7120), .B(n7121), .Z(c[136]) );
  NAND U9258 ( .A(n6691), .B(o[136]), .Z(n7121) );
  NAND U9259 ( .A(n6686), .B(creg[136]), .Z(n7120) );
  NAND U9260 ( .A(n7122), .B(n7123), .Z(c[135]) );
  NAND U9261 ( .A(n6691), .B(o[135]), .Z(n7123) );
  NAND U9262 ( .A(n6686), .B(creg[135]), .Z(n7122) );
  NAND U9263 ( .A(n7124), .B(n7125), .Z(c[134]) );
  NAND U9264 ( .A(n6691), .B(o[134]), .Z(n7125) );
  NAND U9265 ( .A(n6686), .B(creg[134]), .Z(n7124) );
  NAND U9266 ( .A(n7126), .B(n7127), .Z(c[133]) );
  NAND U9267 ( .A(n6691), .B(o[133]), .Z(n7127) );
  NAND U9268 ( .A(n6686), .B(creg[133]), .Z(n7126) );
  NAND U9269 ( .A(n7128), .B(n7129), .Z(c[132]) );
  NAND U9270 ( .A(n6691), .B(o[132]), .Z(n7129) );
  NAND U9271 ( .A(n6686), .B(creg[132]), .Z(n7128) );
  NAND U9272 ( .A(n7130), .B(n7131), .Z(c[131]) );
  NAND U9273 ( .A(n6691), .B(o[131]), .Z(n7131) );
  NAND U9274 ( .A(n6686), .B(creg[131]), .Z(n7130) );
  NAND U9275 ( .A(n7132), .B(n7133), .Z(c[130]) );
  NAND U9276 ( .A(n6691), .B(o[130]), .Z(n7133) );
  NAND U9277 ( .A(n6686), .B(creg[130]), .Z(n7132) );
  NAND U9278 ( .A(n7134), .B(n7135), .Z(c[12]) );
  NAND U9279 ( .A(n6691), .B(o[12]), .Z(n7135) );
  NAND U9280 ( .A(n6686), .B(creg[12]), .Z(n7134) );
  NAND U9281 ( .A(n7136), .B(n7137), .Z(c[129]) );
  NAND U9282 ( .A(n6691), .B(o[129]), .Z(n7137) );
  NAND U9283 ( .A(n6686), .B(creg[129]), .Z(n7136) );
  NAND U9284 ( .A(n7138), .B(n7139), .Z(c[128]) );
  NAND U9285 ( .A(n6691), .B(o[128]), .Z(n7139) );
  NAND U9286 ( .A(n6686), .B(creg[128]), .Z(n7138) );
  NAND U9287 ( .A(n7140), .B(n7141), .Z(c[127]) );
  NAND U9288 ( .A(n6691), .B(o[127]), .Z(n7141) );
  NAND U9289 ( .A(n6686), .B(creg[127]), .Z(n7140) );
  NAND U9290 ( .A(n7142), .B(n7143), .Z(c[126]) );
  NAND U9291 ( .A(n6691), .B(o[126]), .Z(n7143) );
  NAND U9292 ( .A(n6686), .B(creg[126]), .Z(n7142) );
  NAND U9293 ( .A(n7144), .B(n7145), .Z(c[125]) );
  NAND U9294 ( .A(n6691), .B(o[125]), .Z(n7145) );
  NAND U9295 ( .A(n6686), .B(creg[125]), .Z(n7144) );
  NAND U9296 ( .A(n7146), .B(n7147), .Z(c[124]) );
  NAND U9297 ( .A(n6691), .B(o[124]), .Z(n7147) );
  NAND U9298 ( .A(n6686), .B(creg[124]), .Z(n7146) );
  NAND U9299 ( .A(n7148), .B(n7149), .Z(c[123]) );
  NAND U9300 ( .A(n6691), .B(o[123]), .Z(n7149) );
  NAND U9301 ( .A(n6686), .B(creg[123]), .Z(n7148) );
  NAND U9302 ( .A(n7150), .B(n7151), .Z(c[122]) );
  NAND U9303 ( .A(n6691), .B(o[122]), .Z(n7151) );
  NAND U9304 ( .A(n6686), .B(creg[122]), .Z(n7150) );
  NAND U9305 ( .A(n7152), .B(n7153), .Z(c[121]) );
  NAND U9306 ( .A(n6691), .B(o[121]), .Z(n7153) );
  NAND U9307 ( .A(n6686), .B(creg[121]), .Z(n7152) );
  NAND U9308 ( .A(n7154), .B(n7155), .Z(c[120]) );
  NAND U9309 ( .A(n6691), .B(o[120]), .Z(n7155) );
  NAND U9310 ( .A(n6686), .B(creg[120]), .Z(n7154) );
  NAND U9311 ( .A(n7156), .B(n7157), .Z(c[11]) );
  NAND U9312 ( .A(n6691), .B(o[11]), .Z(n7157) );
  NAND U9313 ( .A(n6686), .B(creg[11]), .Z(n7156) );
  NAND U9314 ( .A(n7158), .B(n7159), .Z(c[119]) );
  NAND U9315 ( .A(n6691), .B(o[119]), .Z(n7159) );
  NAND U9316 ( .A(n6686), .B(creg[119]), .Z(n7158) );
  NAND U9317 ( .A(n7160), .B(n7161), .Z(c[118]) );
  NAND U9318 ( .A(n6691), .B(o[118]), .Z(n7161) );
  NAND U9319 ( .A(n6686), .B(creg[118]), .Z(n7160) );
  NAND U9320 ( .A(n7162), .B(n7163), .Z(c[117]) );
  NAND U9321 ( .A(n6691), .B(o[117]), .Z(n7163) );
  NAND U9322 ( .A(n6686), .B(creg[117]), .Z(n7162) );
  NAND U9323 ( .A(n7164), .B(n7165), .Z(c[116]) );
  NAND U9324 ( .A(n6691), .B(o[116]), .Z(n7165) );
  NAND U9325 ( .A(n6686), .B(creg[116]), .Z(n7164) );
  NAND U9326 ( .A(n7166), .B(n7167), .Z(c[115]) );
  NAND U9327 ( .A(n6691), .B(o[115]), .Z(n7167) );
  NAND U9328 ( .A(n6686), .B(creg[115]), .Z(n7166) );
  NAND U9329 ( .A(n7168), .B(n7169), .Z(c[114]) );
  NAND U9330 ( .A(n6691), .B(o[114]), .Z(n7169) );
  NAND U9331 ( .A(n6686), .B(creg[114]), .Z(n7168) );
  NAND U9332 ( .A(n7170), .B(n7171), .Z(c[113]) );
  NAND U9333 ( .A(n6691), .B(o[113]), .Z(n7171) );
  NAND U9334 ( .A(n6686), .B(creg[113]), .Z(n7170) );
  NAND U9335 ( .A(n7172), .B(n7173), .Z(c[112]) );
  NAND U9336 ( .A(n6691), .B(o[112]), .Z(n7173) );
  NAND U9337 ( .A(n6686), .B(creg[112]), .Z(n7172) );
  NAND U9338 ( .A(n7174), .B(n7175), .Z(c[111]) );
  NAND U9339 ( .A(n6691), .B(o[111]), .Z(n7175) );
  NAND U9340 ( .A(n6686), .B(creg[111]), .Z(n7174) );
  NAND U9341 ( .A(n7176), .B(n7177), .Z(c[110]) );
  NAND U9342 ( .A(n6691), .B(o[110]), .Z(n7177) );
  NAND U9343 ( .A(n6686), .B(creg[110]), .Z(n7176) );
  NAND U9344 ( .A(n7178), .B(n7179), .Z(c[10]) );
  NAND U9345 ( .A(n6691), .B(o[10]), .Z(n7179) );
  NAND U9346 ( .A(n6686), .B(creg[10]), .Z(n7178) );
  NAND U9347 ( .A(n7180), .B(n7181), .Z(c[109]) );
  NAND U9348 ( .A(n6691), .B(o[109]), .Z(n7181) );
  NAND U9349 ( .A(n6686), .B(creg[109]), .Z(n7180) );
  NAND U9350 ( .A(n7182), .B(n7183), .Z(c[108]) );
  NAND U9351 ( .A(n6691), .B(o[108]), .Z(n7183) );
  NAND U9352 ( .A(n6686), .B(creg[108]), .Z(n7182) );
  NAND U9353 ( .A(n7184), .B(n7185), .Z(c[107]) );
  NAND U9354 ( .A(n6691), .B(o[107]), .Z(n7185) );
  NAND U9355 ( .A(n6686), .B(creg[107]), .Z(n7184) );
  NAND U9356 ( .A(n7186), .B(n7187), .Z(c[106]) );
  NAND U9357 ( .A(n6691), .B(o[106]), .Z(n7187) );
  NAND U9358 ( .A(n6686), .B(creg[106]), .Z(n7186) );
  NAND U9359 ( .A(n7188), .B(n7189), .Z(c[105]) );
  NAND U9360 ( .A(n6691), .B(o[105]), .Z(n7189) );
  NAND U9361 ( .A(n6686), .B(creg[105]), .Z(n7188) );
  NAND U9362 ( .A(n7190), .B(n7191), .Z(c[104]) );
  NAND U9363 ( .A(n6691), .B(o[104]), .Z(n7191) );
  NAND U9364 ( .A(n6686), .B(creg[104]), .Z(n7190) );
  NAND U9365 ( .A(n7192), .B(n7193), .Z(c[103]) );
  NAND U9366 ( .A(n6691), .B(o[103]), .Z(n7193) );
  NAND U9367 ( .A(n6686), .B(creg[103]), .Z(n7192) );
  NAND U9368 ( .A(n7194), .B(n7195), .Z(c[102]) );
  NAND U9369 ( .A(n6691), .B(o[102]), .Z(n7195) );
  NAND U9370 ( .A(n6686), .B(creg[102]), .Z(n7194) );
  NAND U9371 ( .A(n7196), .B(n7197), .Z(c[101]) );
  NAND U9372 ( .A(n6691), .B(o[101]), .Z(n7197) );
  NAND U9373 ( .A(n6686), .B(creg[101]), .Z(n7196) );
  NAND U9374 ( .A(n7198), .B(n7199), .Z(c[100]) );
  NAND U9375 ( .A(n6691), .B(o[100]), .Z(n7199) );
  NAND U9376 ( .A(n6686), .B(creg[100]), .Z(n7198) );
  NAND U9377 ( .A(n7200), .B(n7201), .Z(c[0]) );
  NAND U9378 ( .A(n6691), .B(o[0]), .Z(n7201) );
  IV U9379 ( .A(n6686), .Z(n6691) );
  NAND U9380 ( .A(n6686), .B(creg[0]), .Z(n7200) );
  NAND U9381 ( .A(n7202), .B(n7203), .Z(n6686) );
  NANDN U9382 ( .A(ereg[255]), .B(init), .Z(n7203) );
  OR U9383 ( .A(init), .B(e[255]), .Z(n7202) );
endmodule

