
module mult_N128_CC32 ( clk, rst, a, b, c );
  input [127:0] a;
  input [3:0] b;
  output [127:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378;
  wire   [127:4] swire;
  wire   [255:128] sreg;

  DFF \sreg_reg[128]  ( .D(swire[4]), .CLK(clk), .RST(rst), .Q(sreg[128]) );
  DFF \sreg_reg[129]  ( .D(swire[5]), .CLK(clk), .RST(rst), .Q(sreg[129]) );
  DFF \sreg_reg[130]  ( .D(swire[6]), .CLK(clk), .RST(rst), .Q(sreg[130]) );
  DFF \sreg_reg[131]  ( .D(swire[7]), .CLK(clk), .RST(rst), .Q(sreg[131]) );
  DFF \sreg_reg[132]  ( .D(swire[8]), .CLK(clk), .RST(rst), .Q(sreg[132]) );
  DFF \sreg_reg[133]  ( .D(swire[9]), .CLK(clk), .RST(rst), .Q(sreg[133]) );
  DFF \sreg_reg[134]  ( .D(swire[10]), .CLK(clk), .RST(rst), .Q(sreg[134]) );
  DFF \sreg_reg[135]  ( .D(swire[11]), .CLK(clk), .RST(rst), .Q(sreg[135]) );
  DFF \sreg_reg[136]  ( .D(swire[12]), .CLK(clk), .RST(rst), .Q(sreg[136]) );
  DFF \sreg_reg[137]  ( .D(swire[13]), .CLK(clk), .RST(rst), .Q(sreg[137]) );
  DFF \sreg_reg[138]  ( .D(swire[14]), .CLK(clk), .RST(rst), .Q(sreg[138]) );
  DFF \sreg_reg[139]  ( .D(swire[15]), .CLK(clk), .RST(rst), .Q(sreg[139]) );
  DFF \sreg_reg[140]  ( .D(swire[16]), .CLK(clk), .RST(rst), .Q(sreg[140]) );
  DFF \sreg_reg[141]  ( .D(swire[17]), .CLK(clk), .RST(rst), .Q(sreg[141]) );
  DFF \sreg_reg[142]  ( .D(swire[18]), .CLK(clk), .RST(rst), .Q(sreg[142]) );
  DFF \sreg_reg[143]  ( .D(swire[19]), .CLK(clk), .RST(rst), .Q(sreg[143]) );
  DFF \sreg_reg[144]  ( .D(swire[20]), .CLK(clk), .RST(rst), .Q(sreg[144]) );
  DFF \sreg_reg[145]  ( .D(swire[21]), .CLK(clk), .RST(rst), .Q(sreg[145]) );
  DFF \sreg_reg[146]  ( .D(swire[22]), .CLK(clk), .RST(rst), .Q(sreg[146]) );
  DFF \sreg_reg[147]  ( .D(swire[23]), .CLK(clk), .RST(rst), .Q(sreg[147]) );
  DFF \sreg_reg[148]  ( .D(swire[24]), .CLK(clk), .RST(rst), .Q(sreg[148]) );
  DFF \sreg_reg[149]  ( .D(swire[25]), .CLK(clk), .RST(rst), .Q(sreg[149]) );
  DFF \sreg_reg[150]  ( .D(swire[26]), .CLK(clk), .RST(rst), .Q(sreg[150]) );
  DFF \sreg_reg[151]  ( .D(swire[27]), .CLK(clk), .RST(rst), .Q(sreg[151]) );
  DFF \sreg_reg[152]  ( .D(swire[28]), .CLK(clk), .RST(rst), .Q(sreg[152]) );
  DFF \sreg_reg[153]  ( .D(swire[29]), .CLK(clk), .RST(rst), .Q(sreg[153]) );
  DFF \sreg_reg[154]  ( .D(swire[30]), .CLK(clk), .RST(rst), .Q(sreg[154]) );
  DFF \sreg_reg[155]  ( .D(swire[31]), .CLK(clk), .RST(rst), .Q(sreg[155]) );
  DFF \sreg_reg[156]  ( .D(swire[32]), .CLK(clk), .RST(rst), .Q(sreg[156]) );
  DFF \sreg_reg[157]  ( .D(swire[33]), .CLK(clk), .RST(rst), .Q(sreg[157]) );
  DFF \sreg_reg[158]  ( .D(swire[34]), .CLK(clk), .RST(rst), .Q(sreg[158]) );
  DFF \sreg_reg[159]  ( .D(swire[35]), .CLK(clk), .RST(rst), .Q(sreg[159]) );
  DFF \sreg_reg[160]  ( .D(swire[36]), .CLK(clk), .RST(rst), .Q(sreg[160]) );
  DFF \sreg_reg[161]  ( .D(swire[37]), .CLK(clk), .RST(rst), .Q(sreg[161]) );
  DFF \sreg_reg[162]  ( .D(swire[38]), .CLK(clk), .RST(rst), .Q(sreg[162]) );
  DFF \sreg_reg[163]  ( .D(swire[39]), .CLK(clk), .RST(rst), .Q(sreg[163]) );
  DFF \sreg_reg[164]  ( .D(swire[40]), .CLK(clk), .RST(rst), .Q(sreg[164]) );
  DFF \sreg_reg[165]  ( .D(swire[41]), .CLK(clk), .RST(rst), .Q(sreg[165]) );
  DFF \sreg_reg[166]  ( .D(swire[42]), .CLK(clk), .RST(rst), .Q(sreg[166]) );
  DFF \sreg_reg[167]  ( .D(swire[43]), .CLK(clk), .RST(rst), .Q(sreg[167]) );
  DFF \sreg_reg[168]  ( .D(swire[44]), .CLK(clk), .RST(rst), .Q(sreg[168]) );
  DFF \sreg_reg[169]  ( .D(swire[45]), .CLK(clk), .RST(rst), .Q(sreg[169]) );
  DFF \sreg_reg[170]  ( .D(swire[46]), .CLK(clk), .RST(rst), .Q(sreg[170]) );
  DFF \sreg_reg[171]  ( .D(swire[47]), .CLK(clk), .RST(rst), .Q(sreg[171]) );
  DFF \sreg_reg[172]  ( .D(swire[48]), .CLK(clk), .RST(rst), .Q(sreg[172]) );
  DFF \sreg_reg[173]  ( .D(swire[49]), .CLK(clk), .RST(rst), .Q(sreg[173]) );
  DFF \sreg_reg[174]  ( .D(swire[50]), .CLK(clk), .RST(rst), .Q(sreg[174]) );
  DFF \sreg_reg[175]  ( .D(swire[51]), .CLK(clk), .RST(rst), .Q(sreg[175]) );
  DFF \sreg_reg[176]  ( .D(swire[52]), .CLK(clk), .RST(rst), .Q(sreg[176]) );
  DFF \sreg_reg[177]  ( .D(swire[53]), .CLK(clk), .RST(rst), .Q(sreg[177]) );
  DFF \sreg_reg[178]  ( .D(swire[54]), .CLK(clk), .RST(rst), .Q(sreg[178]) );
  DFF \sreg_reg[179]  ( .D(swire[55]), .CLK(clk), .RST(rst), .Q(sreg[179]) );
  DFF \sreg_reg[180]  ( .D(swire[56]), .CLK(clk), .RST(rst), .Q(sreg[180]) );
  DFF \sreg_reg[181]  ( .D(swire[57]), .CLK(clk), .RST(rst), .Q(sreg[181]) );
  DFF \sreg_reg[182]  ( .D(swire[58]), .CLK(clk), .RST(rst), .Q(sreg[182]) );
  DFF \sreg_reg[183]  ( .D(swire[59]), .CLK(clk), .RST(rst), .Q(sreg[183]) );
  DFF \sreg_reg[184]  ( .D(swire[60]), .CLK(clk), .RST(rst), .Q(sreg[184]) );
  DFF \sreg_reg[185]  ( .D(swire[61]), .CLK(clk), .RST(rst), .Q(sreg[185]) );
  DFF \sreg_reg[186]  ( .D(swire[62]), .CLK(clk), .RST(rst), .Q(sreg[186]) );
  DFF \sreg_reg[187]  ( .D(swire[63]), .CLK(clk), .RST(rst), .Q(sreg[187]) );
  DFF \sreg_reg[188]  ( .D(swire[64]), .CLK(clk), .RST(rst), .Q(sreg[188]) );
  DFF \sreg_reg[189]  ( .D(swire[65]), .CLK(clk), .RST(rst), .Q(sreg[189]) );
  DFF \sreg_reg[190]  ( .D(swire[66]), .CLK(clk), .RST(rst), .Q(sreg[190]) );
  DFF \sreg_reg[191]  ( .D(swire[67]), .CLK(clk), .RST(rst), .Q(sreg[191]) );
  DFF \sreg_reg[192]  ( .D(swire[68]), .CLK(clk), .RST(rst), .Q(sreg[192]) );
  DFF \sreg_reg[193]  ( .D(swire[69]), .CLK(clk), .RST(rst), .Q(sreg[193]) );
  DFF \sreg_reg[194]  ( .D(swire[70]), .CLK(clk), .RST(rst), .Q(sreg[194]) );
  DFF \sreg_reg[195]  ( .D(swire[71]), .CLK(clk), .RST(rst), .Q(sreg[195]) );
  DFF \sreg_reg[196]  ( .D(swire[72]), .CLK(clk), .RST(rst), .Q(sreg[196]) );
  DFF \sreg_reg[197]  ( .D(swire[73]), .CLK(clk), .RST(rst), .Q(sreg[197]) );
  DFF \sreg_reg[198]  ( .D(swire[74]), .CLK(clk), .RST(rst), .Q(sreg[198]) );
  DFF \sreg_reg[199]  ( .D(swire[75]), .CLK(clk), .RST(rst), .Q(sreg[199]) );
  DFF \sreg_reg[200]  ( .D(swire[76]), .CLK(clk), .RST(rst), .Q(sreg[200]) );
  DFF \sreg_reg[201]  ( .D(swire[77]), .CLK(clk), .RST(rst), .Q(sreg[201]) );
  DFF \sreg_reg[202]  ( .D(swire[78]), .CLK(clk), .RST(rst), .Q(sreg[202]) );
  DFF \sreg_reg[203]  ( .D(swire[79]), .CLK(clk), .RST(rst), .Q(sreg[203]) );
  DFF \sreg_reg[204]  ( .D(swire[80]), .CLK(clk), .RST(rst), .Q(sreg[204]) );
  DFF \sreg_reg[205]  ( .D(swire[81]), .CLK(clk), .RST(rst), .Q(sreg[205]) );
  DFF \sreg_reg[206]  ( .D(swire[82]), .CLK(clk), .RST(rst), .Q(sreg[206]) );
  DFF \sreg_reg[207]  ( .D(swire[83]), .CLK(clk), .RST(rst), .Q(sreg[207]) );
  DFF \sreg_reg[208]  ( .D(swire[84]), .CLK(clk), .RST(rst), .Q(sreg[208]) );
  DFF \sreg_reg[209]  ( .D(swire[85]), .CLK(clk), .RST(rst), .Q(sreg[209]) );
  DFF \sreg_reg[210]  ( .D(swire[86]), .CLK(clk), .RST(rst), .Q(sreg[210]) );
  DFF \sreg_reg[211]  ( .D(swire[87]), .CLK(clk), .RST(rst), .Q(sreg[211]) );
  DFF \sreg_reg[212]  ( .D(swire[88]), .CLK(clk), .RST(rst), .Q(sreg[212]) );
  DFF \sreg_reg[213]  ( .D(swire[89]), .CLK(clk), .RST(rst), .Q(sreg[213]) );
  DFF \sreg_reg[214]  ( .D(swire[90]), .CLK(clk), .RST(rst), .Q(sreg[214]) );
  DFF \sreg_reg[215]  ( .D(swire[91]), .CLK(clk), .RST(rst), .Q(sreg[215]) );
  DFF \sreg_reg[216]  ( .D(swire[92]), .CLK(clk), .RST(rst), .Q(sreg[216]) );
  DFF \sreg_reg[217]  ( .D(swire[93]), .CLK(clk), .RST(rst), .Q(sreg[217]) );
  DFF \sreg_reg[218]  ( .D(swire[94]), .CLK(clk), .RST(rst), .Q(sreg[218]) );
  DFF \sreg_reg[219]  ( .D(swire[95]), .CLK(clk), .RST(rst), .Q(sreg[219]) );
  DFF \sreg_reg[220]  ( .D(swire[96]), .CLK(clk), .RST(rst), .Q(sreg[220]) );
  DFF \sreg_reg[221]  ( .D(swire[97]), .CLK(clk), .RST(rst), .Q(sreg[221]) );
  DFF \sreg_reg[222]  ( .D(swire[98]), .CLK(clk), .RST(rst), .Q(sreg[222]) );
  DFF \sreg_reg[223]  ( .D(swire[99]), .CLK(clk), .RST(rst), .Q(sreg[223]) );
  DFF \sreg_reg[224]  ( .D(swire[100]), .CLK(clk), .RST(rst), .Q(sreg[224]) );
  DFF \sreg_reg[225]  ( .D(swire[101]), .CLK(clk), .RST(rst), .Q(sreg[225]) );
  DFF \sreg_reg[226]  ( .D(swire[102]), .CLK(clk), .RST(rst), .Q(sreg[226]) );
  DFF \sreg_reg[227]  ( .D(swire[103]), .CLK(clk), .RST(rst), .Q(sreg[227]) );
  DFF \sreg_reg[228]  ( .D(swire[104]), .CLK(clk), .RST(rst), .Q(sreg[228]) );
  DFF \sreg_reg[229]  ( .D(swire[105]), .CLK(clk), .RST(rst), .Q(sreg[229]) );
  DFF \sreg_reg[230]  ( .D(swire[106]), .CLK(clk), .RST(rst), .Q(sreg[230]) );
  DFF \sreg_reg[231]  ( .D(swire[107]), .CLK(clk), .RST(rst), .Q(sreg[231]) );
  DFF \sreg_reg[232]  ( .D(swire[108]), .CLK(clk), .RST(rst), .Q(sreg[232]) );
  DFF \sreg_reg[233]  ( .D(swire[109]), .CLK(clk), .RST(rst), .Q(sreg[233]) );
  DFF \sreg_reg[234]  ( .D(swire[110]), .CLK(clk), .RST(rst), .Q(sreg[234]) );
  DFF \sreg_reg[235]  ( .D(swire[111]), .CLK(clk), .RST(rst), .Q(sreg[235]) );
  DFF \sreg_reg[236]  ( .D(swire[112]), .CLK(clk), .RST(rst), .Q(sreg[236]) );
  DFF \sreg_reg[237]  ( .D(swire[113]), .CLK(clk), .RST(rst), .Q(sreg[237]) );
  DFF \sreg_reg[238]  ( .D(swire[114]), .CLK(clk), .RST(rst), .Q(sreg[238]) );
  DFF \sreg_reg[239]  ( .D(swire[115]), .CLK(clk), .RST(rst), .Q(sreg[239]) );
  DFF \sreg_reg[240]  ( .D(swire[116]), .CLK(clk), .RST(rst), .Q(sreg[240]) );
  DFF \sreg_reg[241]  ( .D(swire[117]), .CLK(clk), .RST(rst), .Q(sreg[241]) );
  DFF \sreg_reg[242]  ( .D(swire[118]), .CLK(clk), .RST(rst), .Q(sreg[242]) );
  DFF \sreg_reg[243]  ( .D(swire[119]), .CLK(clk), .RST(rst), .Q(sreg[243]) );
  DFF \sreg_reg[244]  ( .D(swire[120]), .CLK(clk), .RST(rst), .Q(sreg[244]) );
  DFF \sreg_reg[245]  ( .D(swire[121]), .CLK(clk), .RST(rst), .Q(sreg[245]) );
  DFF \sreg_reg[246]  ( .D(swire[122]), .CLK(clk), .RST(rst), .Q(sreg[246]) );
  DFF \sreg_reg[247]  ( .D(swire[123]), .CLK(clk), .RST(rst), .Q(sreg[247]) );
  DFF \sreg_reg[248]  ( .D(swire[124]), .CLK(clk), .RST(rst), .Q(sreg[248]) );
  DFF \sreg_reg[249]  ( .D(swire[125]), .CLK(clk), .RST(rst), .Q(sreg[249]) );
  DFF \sreg_reg[250]  ( .D(swire[126]), .CLK(clk), .RST(rst), .Q(sreg[250]) );
  DFF \sreg_reg[251]  ( .D(swire[127]), .CLK(clk), .RST(rst), .Q(sreg[251]) );
  DFF \sreg_reg[127]  ( .D(c[127]), .CLK(clk), .RST(rst), .Q(c[123]) );
  DFF \sreg_reg[126]  ( .D(c[126]), .CLK(clk), .RST(rst), .Q(c[122]) );
  DFF \sreg_reg[125]  ( .D(c[125]), .CLK(clk), .RST(rst), .Q(c[121]) );
  DFF \sreg_reg[124]  ( .D(c[124]), .CLK(clk), .RST(rst), .Q(c[120]) );
  DFF \sreg_reg[123]  ( .D(c[123]), .CLK(clk), .RST(rst), .Q(c[119]) );
  DFF \sreg_reg[122]  ( .D(c[122]), .CLK(clk), .RST(rst), .Q(c[118]) );
  DFF \sreg_reg[121]  ( .D(c[121]), .CLK(clk), .RST(rst), .Q(c[117]) );
  DFF \sreg_reg[120]  ( .D(c[120]), .CLK(clk), .RST(rst), .Q(c[116]) );
  DFF \sreg_reg[119]  ( .D(c[119]), .CLK(clk), .RST(rst), .Q(c[115]) );
  DFF \sreg_reg[118]  ( .D(c[118]), .CLK(clk), .RST(rst), .Q(c[114]) );
  DFF \sreg_reg[117]  ( .D(c[117]), .CLK(clk), .RST(rst), .Q(c[113]) );
  DFF \sreg_reg[116]  ( .D(c[116]), .CLK(clk), .RST(rst), .Q(c[112]) );
  DFF \sreg_reg[115]  ( .D(c[115]), .CLK(clk), .RST(rst), .Q(c[111]) );
  DFF \sreg_reg[114]  ( .D(c[114]), .CLK(clk), .RST(rst), .Q(c[110]) );
  DFF \sreg_reg[113]  ( .D(c[113]), .CLK(clk), .RST(rst), .Q(c[109]) );
  DFF \sreg_reg[112]  ( .D(c[112]), .CLK(clk), .RST(rst), .Q(c[108]) );
  DFF \sreg_reg[111]  ( .D(c[111]), .CLK(clk), .RST(rst), .Q(c[107]) );
  DFF \sreg_reg[110]  ( .D(c[110]), .CLK(clk), .RST(rst), .Q(c[106]) );
  DFF \sreg_reg[109]  ( .D(c[109]), .CLK(clk), .RST(rst), .Q(c[105]) );
  DFF \sreg_reg[108]  ( .D(c[108]), .CLK(clk), .RST(rst), .Q(c[104]) );
  DFF \sreg_reg[107]  ( .D(c[107]), .CLK(clk), .RST(rst), .Q(c[103]) );
  DFF \sreg_reg[106]  ( .D(c[106]), .CLK(clk), .RST(rst), .Q(c[102]) );
  DFF \sreg_reg[105]  ( .D(c[105]), .CLK(clk), .RST(rst), .Q(c[101]) );
  DFF \sreg_reg[104]  ( .D(c[104]), .CLK(clk), .RST(rst), .Q(c[100]) );
  DFF \sreg_reg[103]  ( .D(c[103]), .CLK(clk), .RST(rst), .Q(c[99]) );
  DFF \sreg_reg[102]  ( .D(c[102]), .CLK(clk), .RST(rst), .Q(c[98]) );
  DFF \sreg_reg[101]  ( .D(c[101]), .CLK(clk), .RST(rst), .Q(c[97]) );
  DFF \sreg_reg[100]  ( .D(c[100]), .CLK(clk), .RST(rst), .Q(c[96]) );
  DFF \sreg_reg[99]  ( .D(c[99]), .CLK(clk), .RST(rst), .Q(c[95]) );
  DFF \sreg_reg[98]  ( .D(c[98]), .CLK(clk), .RST(rst), .Q(c[94]) );
  DFF \sreg_reg[97]  ( .D(c[97]), .CLK(clk), .RST(rst), .Q(c[93]) );
  DFF \sreg_reg[96]  ( .D(c[96]), .CLK(clk), .RST(rst), .Q(c[92]) );
  DFF \sreg_reg[95]  ( .D(c[95]), .CLK(clk), .RST(rst), .Q(c[91]) );
  DFF \sreg_reg[94]  ( .D(c[94]), .CLK(clk), .RST(rst), .Q(c[90]) );
  DFF \sreg_reg[93]  ( .D(c[93]), .CLK(clk), .RST(rst), .Q(c[89]) );
  DFF \sreg_reg[92]  ( .D(c[92]), .CLK(clk), .RST(rst), .Q(c[88]) );
  DFF \sreg_reg[91]  ( .D(c[91]), .CLK(clk), .RST(rst), .Q(c[87]) );
  DFF \sreg_reg[90]  ( .D(c[90]), .CLK(clk), .RST(rst), .Q(c[86]) );
  DFF \sreg_reg[89]  ( .D(c[89]), .CLK(clk), .RST(rst), .Q(c[85]) );
  DFF \sreg_reg[88]  ( .D(c[88]), .CLK(clk), .RST(rst), .Q(c[84]) );
  DFF \sreg_reg[87]  ( .D(c[87]), .CLK(clk), .RST(rst), .Q(c[83]) );
  DFF \sreg_reg[86]  ( .D(c[86]), .CLK(clk), .RST(rst), .Q(c[82]) );
  DFF \sreg_reg[85]  ( .D(c[85]), .CLK(clk), .RST(rst), .Q(c[81]) );
  DFF \sreg_reg[84]  ( .D(c[84]), .CLK(clk), .RST(rst), .Q(c[80]) );
  DFF \sreg_reg[83]  ( .D(c[83]), .CLK(clk), .RST(rst), .Q(c[79]) );
  DFF \sreg_reg[82]  ( .D(c[82]), .CLK(clk), .RST(rst), .Q(c[78]) );
  DFF \sreg_reg[81]  ( .D(c[81]), .CLK(clk), .RST(rst), .Q(c[77]) );
  DFF \sreg_reg[80]  ( .D(c[80]), .CLK(clk), .RST(rst), .Q(c[76]) );
  DFF \sreg_reg[79]  ( .D(c[79]), .CLK(clk), .RST(rst), .Q(c[75]) );
  DFF \sreg_reg[78]  ( .D(c[78]), .CLK(clk), .RST(rst), .Q(c[74]) );
  DFF \sreg_reg[77]  ( .D(c[77]), .CLK(clk), .RST(rst), .Q(c[73]) );
  DFF \sreg_reg[76]  ( .D(c[76]), .CLK(clk), .RST(rst), .Q(c[72]) );
  DFF \sreg_reg[75]  ( .D(c[75]), .CLK(clk), .RST(rst), .Q(c[71]) );
  DFF \sreg_reg[74]  ( .D(c[74]), .CLK(clk), .RST(rst), .Q(c[70]) );
  DFF \sreg_reg[73]  ( .D(c[73]), .CLK(clk), .RST(rst), .Q(c[69]) );
  DFF \sreg_reg[72]  ( .D(c[72]), .CLK(clk), .RST(rst), .Q(c[68]) );
  DFF \sreg_reg[71]  ( .D(c[71]), .CLK(clk), .RST(rst), .Q(c[67]) );
  DFF \sreg_reg[70]  ( .D(c[70]), .CLK(clk), .RST(rst), .Q(c[66]) );
  DFF \sreg_reg[69]  ( .D(c[69]), .CLK(clk), .RST(rst), .Q(c[65]) );
  DFF \sreg_reg[68]  ( .D(c[68]), .CLK(clk), .RST(rst), .Q(c[64]) );
  DFF \sreg_reg[67]  ( .D(c[67]), .CLK(clk), .RST(rst), .Q(c[63]) );
  DFF \sreg_reg[66]  ( .D(c[66]), .CLK(clk), .RST(rst), .Q(c[62]) );
  DFF \sreg_reg[65]  ( .D(c[65]), .CLK(clk), .RST(rst), .Q(c[61]) );
  DFF \sreg_reg[64]  ( .D(c[64]), .CLK(clk), .RST(rst), .Q(c[60]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[59]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[58]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[57]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[56]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[55]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[54]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[53]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[52]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[51]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[50]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[49]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[48]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[47]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[46]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[45]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[44]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[43]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[42]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[41]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[40]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[39]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[38]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[37]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[36]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[35]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[34]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[33]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[32]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[31]  ( .D(c[31]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[30]  ( .D(c[30]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[29]  ( .D(c[29]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[28]  ( .D(c[28]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[27]  ( .D(c[27]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[26]  ( .D(c[26]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[25]  ( .D(c[25]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[24]  ( .D(c[24]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[23]  ( .D(c[23]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[22]  ( .D(c[22]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[21]  ( .D(c[21]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[20]  ( .D(c[20]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[19]  ( .D(c[19]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[18]  ( .D(c[18]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[17]  ( .D(c[17]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[16]  ( .D(c[16]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[15]  ( .D(c[15]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[14]  ( .D(c[14]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[13]  ( .D(c[13]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[12]  ( .D(c[12]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[11]  ( .D(c[11]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[10]  ( .D(c[10]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[9]  ( .D(c[9]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[8]  ( .D(c[8]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[7]  ( .D(c[7]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[6]  ( .D(c[6]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[5]  ( .D(c[5]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[4]  ( .D(c[4]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XOR U7 ( .A(n1368), .B(n1359), .Z(n1367) );
  NAND U8 ( .A(n211), .B(n210), .Z(n201) );
  XOR U9 ( .A(n1), .B(n2), .Z(swire[9]) );
  XOR U10 ( .A(n3), .B(n4), .Z(swire[99]) );
  XOR U11 ( .A(n5), .B(n6), .Z(swire[98]) );
  XOR U12 ( .A(n7), .B(n8), .Z(swire[97]) );
  XOR U13 ( .A(n9), .B(n10), .Z(swire[96]) );
  XOR U14 ( .A(n11), .B(n12), .Z(swire[95]) );
  XOR U15 ( .A(n13), .B(n14), .Z(swire[94]) );
  XOR U16 ( .A(n15), .B(n16), .Z(swire[93]) );
  XOR U17 ( .A(n17), .B(n18), .Z(swire[92]) );
  XOR U18 ( .A(n19), .B(n20), .Z(swire[91]) );
  XOR U19 ( .A(n21), .B(n22), .Z(swire[90]) );
  XOR U20 ( .A(n23), .B(n24), .Z(swire[8]) );
  XOR U21 ( .A(n25), .B(n26), .Z(swire[89]) );
  XOR U22 ( .A(n27), .B(n28), .Z(swire[88]) );
  XOR U23 ( .A(n29), .B(n30), .Z(swire[87]) );
  XOR U24 ( .A(n31), .B(n32), .Z(swire[86]) );
  XOR U25 ( .A(n33), .B(n34), .Z(swire[85]) );
  XOR U26 ( .A(n35), .B(n36), .Z(swire[84]) );
  XOR U27 ( .A(n37), .B(n38), .Z(swire[83]) );
  XOR U28 ( .A(n39), .B(n40), .Z(swire[82]) );
  XOR U29 ( .A(n41), .B(n42), .Z(swire[81]) );
  XOR U30 ( .A(n43), .B(n44), .Z(swire[80]) );
  XOR U31 ( .A(n45), .B(n46), .Z(swire[7]) );
  XOR U32 ( .A(n47), .B(n48), .Z(swire[79]) );
  XOR U33 ( .A(n49), .B(n50), .Z(swire[78]) );
  XOR U34 ( .A(n51), .B(n52), .Z(swire[77]) );
  XOR U35 ( .A(n53), .B(n54), .Z(swire[76]) );
  XOR U36 ( .A(n55), .B(n56), .Z(swire[75]) );
  XOR U37 ( .A(n57), .B(n58), .Z(swire[74]) );
  XOR U38 ( .A(n59), .B(n60), .Z(swire[73]) );
  XOR U39 ( .A(n61), .B(n62), .Z(swire[72]) );
  XOR U40 ( .A(n63), .B(n64), .Z(swire[71]) );
  XOR U41 ( .A(n65), .B(n66), .Z(swire[70]) );
  XOR U42 ( .A(n67), .B(n68), .Z(swire[6]) );
  XOR U43 ( .A(n69), .B(n70), .Z(swire[69]) );
  XOR U44 ( .A(n71), .B(n72), .Z(swire[68]) );
  XOR U45 ( .A(n73), .B(n74), .Z(swire[67]) );
  XOR U46 ( .A(n75), .B(n76), .Z(swire[66]) );
  XOR U47 ( .A(n77), .B(n78), .Z(swire[65]) );
  XOR U48 ( .A(n79), .B(n80), .Z(swire[64]) );
  XOR U49 ( .A(n81), .B(n82), .Z(swire[63]) );
  XOR U50 ( .A(n83), .B(n84), .Z(swire[62]) );
  XOR U51 ( .A(n85), .B(n86), .Z(swire[61]) );
  XOR U52 ( .A(n87), .B(n88), .Z(swire[60]) );
  XOR U53 ( .A(n89), .B(n90), .Z(swire[5]) );
  XOR U54 ( .A(n91), .B(n92), .Z(swire[59]) );
  XOR U55 ( .A(n93), .B(n94), .Z(swire[58]) );
  XOR U56 ( .A(n95), .B(n96), .Z(swire[57]) );
  XOR U57 ( .A(n97), .B(n98), .Z(swire[56]) );
  XOR U58 ( .A(n99), .B(n100), .Z(swire[55]) );
  XOR U59 ( .A(n101), .B(n102), .Z(swire[54]) );
  XOR U60 ( .A(n103), .B(n104), .Z(swire[53]) );
  XOR U61 ( .A(n105), .B(n106), .Z(swire[52]) );
  XOR U62 ( .A(n107), .B(n108), .Z(swire[51]) );
  XOR U63 ( .A(n109), .B(n110), .Z(swire[50]) );
  XOR U64 ( .A(n111), .B(n112), .Z(swire[4]) );
  XOR U65 ( .A(n113), .B(n114), .Z(swire[49]) );
  XOR U66 ( .A(n115), .B(n116), .Z(swire[48]) );
  XOR U67 ( .A(n117), .B(n118), .Z(swire[47]) );
  XOR U68 ( .A(n119), .B(n120), .Z(swire[46]) );
  XOR U69 ( .A(n121), .B(n122), .Z(swire[45]) );
  XOR U70 ( .A(n123), .B(n124), .Z(swire[44]) );
  XOR U71 ( .A(n125), .B(n126), .Z(swire[43]) );
  XOR U72 ( .A(n127), .B(n128), .Z(swire[42]) );
  XOR U73 ( .A(n129), .B(n130), .Z(swire[41]) );
  XOR U74 ( .A(n131), .B(n132), .Z(swire[40]) );
  XOR U75 ( .A(n133), .B(n134), .Z(swire[39]) );
  XOR U76 ( .A(n135), .B(n136), .Z(swire[38]) );
  XOR U77 ( .A(n137), .B(n138), .Z(swire[37]) );
  XOR U78 ( .A(n139), .B(n140), .Z(swire[36]) );
  XOR U79 ( .A(n141), .B(n142), .Z(swire[35]) );
  XOR U80 ( .A(n143), .B(n144), .Z(swire[34]) );
  XOR U81 ( .A(n145), .B(n146), .Z(swire[33]) );
  XOR U82 ( .A(n147), .B(n148), .Z(swire[32]) );
  XOR U83 ( .A(n149), .B(n150), .Z(swire[31]) );
  XOR U84 ( .A(n151), .B(n152), .Z(swire[30]) );
  XOR U85 ( .A(n153), .B(n154), .Z(swire[29]) );
  XOR U86 ( .A(n155), .B(n156), .Z(swire[28]) );
  XOR U87 ( .A(n157), .B(n158), .Z(swire[27]) );
  XOR U88 ( .A(n159), .B(n160), .Z(swire[26]) );
  XOR U89 ( .A(n161), .B(n162), .Z(swire[25]) );
  XOR U90 ( .A(n163), .B(n164), .Z(swire[24]) );
  XOR U91 ( .A(n165), .B(n166), .Z(swire[23]) );
  XOR U92 ( .A(n167), .B(n168), .Z(swire[22]) );
  XOR U93 ( .A(n169), .B(n170), .Z(swire[21]) );
  XOR U94 ( .A(n171), .B(n172), .Z(swire[20]) );
  XOR U95 ( .A(n173), .B(n174), .Z(swire[19]) );
  XOR U96 ( .A(n175), .B(n176), .Z(swire[18]) );
  XOR U97 ( .A(n177), .B(n178), .Z(swire[17]) );
  XOR U98 ( .A(n179), .B(n180), .Z(swire[16]) );
  XOR U99 ( .A(n181), .B(n182), .Z(swire[15]) );
  XOR U100 ( .A(n183), .B(n184), .Z(swire[14]) );
  XOR U101 ( .A(n185), .B(n186), .Z(swire[13]) );
  XOR U102 ( .A(n187), .B(n188), .Z(swire[12]) );
  XOR U103 ( .A(n189), .B(n190), .Z(swire[127]) );
  XOR U104 ( .A(n191), .B(n192), .Z(n190) );
  AND U105 ( .A(a[127]), .B(b[0]), .Z(n192) );
  AND U106 ( .A(b[1]), .B(a[126]), .Z(n191) );
  XOR U107 ( .A(n193), .B(n194), .Z(n189) );
  AND U108 ( .A(b[2]), .B(a[125]), .Z(n194) );
  AND U109 ( .A(b[3]), .B(a[124]), .Z(n193) );
  XOR U110 ( .A(n195), .B(n196), .Z(swire[126]) );
  XOR U111 ( .A(n197), .B(n198), .Z(n196) );
  AND U112 ( .A(a[126]), .B(b[0]), .Z(n198) );
  AND U113 ( .A(b[1]), .B(a[125]), .Z(n197) );
  XOR U114 ( .A(n199), .B(n200), .Z(n195) );
  AND U115 ( .A(b[2]), .B(a[124]), .Z(n200) );
  AND U116 ( .A(b[3]), .B(a[123]), .Z(n199) );
  XNOR U117 ( .A(n201), .B(n202), .Z(swire[125]) );
  XOR U118 ( .A(n203), .B(n204), .Z(n202) );
  XNOR U119 ( .A(n205), .B(n201), .Z(n204) );
  AND U120 ( .A(a[125]), .B(b[0]), .Z(n205) );
  XOR U121 ( .A(n206), .B(n207), .Z(n203) );
  XOR U122 ( .A(n208), .B(n209), .Z(n207) );
  AND U123 ( .A(a[123]), .B(b[2]), .Z(n209) );
  AND U124 ( .A(a[122]), .B(b[3]), .Z(n208) );
  AND U125 ( .A(a[124]), .B(b[1]), .Z(n206) );
  XNOR U126 ( .A(n210), .B(n211), .Z(swire[124]) );
  XOR U127 ( .A(n212), .B(n213), .Z(n211) );
  XNOR U128 ( .A(n214), .B(n210), .Z(n213) );
  AND U129 ( .A(b[0]), .B(a[124]), .Z(n214) );
  XOR U130 ( .A(n215), .B(n216), .Z(n212) );
  XOR U131 ( .A(n217), .B(n218), .Z(n216) );
  AND U132 ( .A(b[2]), .B(a[122]), .Z(n218) );
  AND U133 ( .A(a[121]), .B(b[3]), .Z(n217) );
  AND U134 ( .A(b[1]), .B(a[123]), .Z(n215) );
  XNOR U135 ( .A(n219), .B(n220), .Z(n210) );
  NOR U136 ( .A(n221), .B(n222), .Z(n219) );
  XOR U137 ( .A(n222), .B(n221), .Z(swire[123]) );
  XOR U138 ( .A(sreg[251]), .B(n220), .Z(n221) );
  XOR U139 ( .A(n223), .B(n224), .Z(n222) );
  XOR U140 ( .A(n225), .B(n220), .Z(n224) );
  XOR U141 ( .A(n226), .B(n227), .Z(n220) );
  NOR U142 ( .A(n228), .B(n229), .Z(n226) );
  AND U143 ( .A(b[0]), .B(a[123]), .Z(n225) );
  XOR U144 ( .A(n230), .B(n231), .Z(n223) );
  XOR U145 ( .A(n232), .B(n233), .Z(n231) );
  AND U146 ( .A(b[2]), .B(a[121]), .Z(n233) );
  AND U147 ( .A(a[120]), .B(b[3]), .Z(n232) );
  AND U148 ( .A(b[1]), .B(a[122]), .Z(n230) );
  XOR U149 ( .A(n229), .B(n228), .Z(swire[122]) );
  XOR U150 ( .A(sreg[250]), .B(n227), .Z(n228) );
  XOR U151 ( .A(n234), .B(n235), .Z(n229) );
  XOR U152 ( .A(n236), .B(n227), .Z(n235) );
  XOR U153 ( .A(n237), .B(n238), .Z(n227) );
  NOR U154 ( .A(n239), .B(n240), .Z(n237) );
  AND U155 ( .A(b[0]), .B(a[122]), .Z(n236) );
  XOR U156 ( .A(n241), .B(n242), .Z(n234) );
  XOR U157 ( .A(n243), .B(n244), .Z(n242) );
  AND U158 ( .A(b[2]), .B(a[120]), .Z(n244) );
  AND U159 ( .A(a[119]), .B(b[3]), .Z(n243) );
  AND U160 ( .A(b[1]), .B(a[121]), .Z(n241) );
  XOR U161 ( .A(n240), .B(n239), .Z(swire[121]) );
  XOR U162 ( .A(sreg[249]), .B(n238), .Z(n239) );
  XOR U163 ( .A(n245), .B(n246), .Z(n240) );
  XOR U164 ( .A(n247), .B(n238), .Z(n246) );
  XOR U165 ( .A(n248), .B(n249), .Z(n238) );
  NOR U166 ( .A(n250), .B(n251), .Z(n248) );
  AND U167 ( .A(b[0]), .B(a[121]), .Z(n247) );
  XOR U168 ( .A(n252), .B(n253), .Z(n245) );
  XOR U169 ( .A(n254), .B(n255), .Z(n253) );
  AND U170 ( .A(b[2]), .B(a[119]), .Z(n255) );
  AND U171 ( .A(a[118]), .B(b[3]), .Z(n254) );
  AND U172 ( .A(b[1]), .B(a[120]), .Z(n252) );
  XOR U173 ( .A(n251), .B(n250), .Z(swire[120]) );
  XOR U174 ( .A(sreg[248]), .B(n249), .Z(n250) );
  XOR U175 ( .A(n256), .B(n257), .Z(n251) );
  XOR U176 ( .A(n258), .B(n249), .Z(n257) );
  XOR U177 ( .A(n259), .B(n260), .Z(n249) );
  NOR U178 ( .A(n261), .B(n262), .Z(n259) );
  AND U179 ( .A(b[0]), .B(a[120]), .Z(n258) );
  XOR U180 ( .A(n263), .B(n264), .Z(n256) );
  XOR U181 ( .A(n265), .B(n266), .Z(n264) );
  AND U182 ( .A(b[2]), .B(a[118]), .Z(n266) );
  AND U183 ( .A(a[117]), .B(b[3]), .Z(n265) );
  AND U184 ( .A(b[1]), .B(a[119]), .Z(n263) );
  XOR U185 ( .A(n267), .B(n268), .Z(swire[11]) );
  XOR U186 ( .A(n262), .B(n261), .Z(swire[119]) );
  XOR U187 ( .A(sreg[247]), .B(n260), .Z(n261) );
  XOR U188 ( .A(n269), .B(n270), .Z(n262) );
  XOR U189 ( .A(n271), .B(n260), .Z(n270) );
  XOR U190 ( .A(n272), .B(n273), .Z(n260) );
  NOR U191 ( .A(n274), .B(n275), .Z(n272) );
  AND U192 ( .A(b[0]), .B(a[119]), .Z(n271) );
  XOR U193 ( .A(n276), .B(n277), .Z(n269) );
  XOR U194 ( .A(n278), .B(n279), .Z(n277) );
  AND U195 ( .A(b[2]), .B(a[117]), .Z(n279) );
  AND U196 ( .A(a[116]), .B(b[3]), .Z(n278) );
  AND U197 ( .A(b[1]), .B(a[118]), .Z(n276) );
  XOR U198 ( .A(n275), .B(n274), .Z(swire[118]) );
  XOR U199 ( .A(sreg[246]), .B(n273), .Z(n274) );
  XOR U200 ( .A(n280), .B(n281), .Z(n275) );
  XOR U201 ( .A(n282), .B(n273), .Z(n281) );
  XOR U202 ( .A(n283), .B(n284), .Z(n273) );
  NOR U203 ( .A(n285), .B(n286), .Z(n283) );
  AND U204 ( .A(b[0]), .B(a[118]), .Z(n282) );
  XOR U205 ( .A(n287), .B(n288), .Z(n280) );
  XOR U206 ( .A(n289), .B(n290), .Z(n288) );
  AND U207 ( .A(b[2]), .B(a[116]), .Z(n290) );
  AND U208 ( .A(a[115]), .B(b[3]), .Z(n289) );
  AND U209 ( .A(b[1]), .B(a[117]), .Z(n287) );
  XOR U210 ( .A(n286), .B(n285), .Z(swire[117]) );
  XOR U211 ( .A(sreg[245]), .B(n284), .Z(n285) );
  XOR U212 ( .A(n291), .B(n292), .Z(n286) );
  XOR U213 ( .A(n293), .B(n284), .Z(n292) );
  XOR U214 ( .A(n294), .B(n295), .Z(n284) );
  NOR U215 ( .A(n296), .B(n297), .Z(n294) );
  AND U216 ( .A(b[0]), .B(a[117]), .Z(n293) );
  XOR U217 ( .A(n298), .B(n299), .Z(n291) );
  XOR U218 ( .A(n300), .B(n301), .Z(n299) );
  AND U219 ( .A(b[2]), .B(a[115]), .Z(n301) );
  AND U220 ( .A(a[114]), .B(b[3]), .Z(n300) );
  AND U221 ( .A(b[1]), .B(a[116]), .Z(n298) );
  XOR U222 ( .A(n297), .B(n296), .Z(swire[116]) );
  XOR U223 ( .A(sreg[244]), .B(n295), .Z(n296) );
  XOR U224 ( .A(n302), .B(n303), .Z(n297) );
  XOR U225 ( .A(n304), .B(n295), .Z(n303) );
  XOR U226 ( .A(n305), .B(n306), .Z(n295) );
  NOR U227 ( .A(n307), .B(n308), .Z(n305) );
  AND U228 ( .A(b[0]), .B(a[116]), .Z(n304) );
  XOR U229 ( .A(n309), .B(n310), .Z(n302) );
  XOR U230 ( .A(n311), .B(n312), .Z(n310) );
  AND U231 ( .A(b[2]), .B(a[114]), .Z(n312) );
  AND U232 ( .A(a[113]), .B(b[3]), .Z(n311) );
  AND U233 ( .A(b[1]), .B(a[115]), .Z(n309) );
  XOR U234 ( .A(n308), .B(n307), .Z(swire[115]) );
  XOR U235 ( .A(sreg[243]), .B(n306), .Z(n307) );
  XOR U236 ( .A(n313), .B(n314), .Z(n308) );
  XOR U237 ( .A(n315), .B(n306), .Z(n314) );
  XOR U238 ( .A(n316), .B(n317), .Z(n306) );
  NOR U239 ( .A(n318), .B(n319), .Z(n316) );
  AND U240 ( .A(b[0]), .B(a[115]), .Z(n315) );
  XOR U241 ( .A(n320), .B(n321), .Z(n313) );
  XOR U242 ( .A(n322), .B(n323), .Z(n321) );
  AND U243 ( .A(b[2]), .B(a[113]), .Z(n323) );
  AND U244 ( .A(a[112]), .B(b[3]), .Z(n322) );
  AND U245 ( .A(b[1]), .B(a[114]), .Z(n320) );
  XOR U246 ( .A(n319), .B(n318), .Z(swire[114]) );
  XOR U247 ( .A(sreg[242]), .B(n317), .Z(n318) );
  XOR U248 ( .A(n324), .B(n325), .Z(n319) );
  XOR U249 ( .A(n326), .B(n317), .Z(n325) );
  XOR U250 ( .A(n327), .B(n328), .Z(n317) );
  NOR U251 ( .A(n329), .B(n330), .Z(n327) );
  AND U252 ( .A(b[0]), .B(a[114]), .Z(n326) );
  XOR U253 ( .A(n331), .B(n332), .Z(n324) );
  XOR U254 ( .A(n333), .B(n334), .Z(n332) );
  AND U255 ( .A(b[2]), .B(a[112]), .Z(n334) );
  AND U256 ( .A(a[111]), .B(b[3]), .Z(n333) );
  AND U257 ( .A(b[1]), .B(a[113]), .Z(n331) );
  XOR U258 ( .A(n330), .B(n329), .Z(swire[113]) );
  XOR U259 ( .A(sreg[241]), .B(n328), .Z(n329) );
  XOR U260 ( .A(n335), .B(n336), .Z(n330) );
  XOR U261 ( .A(n337), .B(n328), .Z(n336) );
  XOR U262 ( .A(n338), .B(n339), .Z(n328) );
  NOR U263 ( .A(n340), .B(n341), .Z(n338) );
  AND U264 ( .A(b[0]), .B(a[113]), .Z(n337) );
  XOR U265 ( .A(n342), .B(n343), .Z(n335) );
  XOR U266 ( .A(n344), .B(n345), .Z(n343) );
  AND U267 ( .A(b[2]), .B(a[111]), .Z(n345) );
  AND U268 ( .A(a[110]), .B(b[3]), .Z(n344) );
  AND U269 ( .A(b[1]), .B(a[112]), .Z(n342) );
  XOR U270 ( .A(n341), .B(n340), .Z(swire[112]) );
  XOR U271 ( .A(sreg[240]), .B(n339), .Z(n340) );
  XOR U272 ( .A(n346), .B(n347), .Z(n341) );
  XOR U273 ( .A(n348), .B(n339), .Z(n347) );
  XOR U274 ( .A(n349), .B(n350), .Z(n339) );
  NOR U275 ( .A(n351), .B(n352), .Z(n349) );
  AND U276 ( .A(b[0]), .B(a[112]), .Z(n348) );
  XOR U277 ( .A(n353), .B(n354), .Z(n346) );
  XOR U278 ( .A(n355), .B(n356), .Z(n354) );
  AND U279 ( .A(b[2]), .B(a[110]), .Z(n356) );
  AND U280 ( .A(a[109]), .B(b[3]), .Z(n355) );
  AND U281 ( .A(b[1]), .B(a[111]), .Z(n353) );
  XOR U282 ( .A(n352), .B(n351), .Z(swire[111]) );
  XOR U283 ( .A(sreg[239]), .B(n350), .Z(n351) );
  XOR U284 ( .A(n357), .B(n358), .Z(n352) );
  XOR U285 ( .A(n359), .B(n350), .Z(n358) );
  XOR U286 ( .A(n360), .B(n361), .Z(n350) );
  NOR U287 ( .A(n362), .B(n363), .Z(n360) );
  AND U288 ( .A(b[0]), .B(a[111]), .Z(n359) );
  XOR U289 ( .A(n364), .B(n365), .Z(n357) );
  XOR U290 ( .A(n366), .B(n367), .Z(n365) );
  AND U291 ( .A(b[2]), .B(a[109]), .Z(n367) );
  AND U292 ( .A(a[108]), .B(b[3]), .Z(n366) );
  AND U293 ( .A(b[1]), .B(a[110]), .Z(n364) );
  XOR U294 ( .A(n363), .B(n362), .Z(swire[110]) );
  XOR U295 ( .A(sreg[238]), .B(n361), .Z(n362) );
  XOR U296 ( .A(n368), .B(n369), .Z(n363) );
  XOR U297 ( .A(n370), .B(n361), .Z(n369) );
  XOR U298 ( .A(n371), .B(n372), .Z(n361) );
  NOR U299 ( .A(n373), .B(n374), .Z(n371) );
  AND U300 ( .A(b[0]), .B(a[110]), .Z(n370) );
  XOR U301 ( .A(n375), .B(n376), .Z(n368) );
  XOR U302 ( .A(n377), .B(n378), .Z(n376) );
  AND U303 ( .A(b[2]), .B(a[108]), .Z(n378) );
  AND U304 ( .A(a[107]), .B(b[3]), .Z(n377) );
  AND U305 ( .A(b[1]), .B(a[109]), .Z(n375) );
  XOR U306 ( .A(n379), .B(n380), .Z(swire[10]) );
  XOR U307 ( .A(n374), .B(n373), .Z(swire[109]) );
  XOR U308 ( .A(sreg[237]), .B(n372), .Z(n373) );
  XOR U309 ( .A(n381), .B(n382), .Z(n374) );
  XOR U310 ( .A(n383), .B(n372), .Z(n382) );
  XOR U311 ( .A(n384), .B(n385), .Z(n372) );
  NOR U312 ( .A(n386), .B(n387), .Z(n384) );
  AND U313 ( .A(b[0]), .B(a[109]), .Z(n383) );
  XOR U314 ( .A(n388), .B(n389), .Z(n381) );
  XOR U315 ( .A(n390), .B(n391), .Z(n389) );
  AND U316 ( .A(b[2]), .B(a[107]), .Z(n391) );
  AND U317 ( .A(a[106]), .B(b[3]), .Z(n390) );
  AND U318 ( .A(b[1]), .B(a[108]), .Z(n388) );
  XOR U319 ( .A(n387), .B(n386), .Z(swire[108]) );
  XOR U320 ( .A(sreg[236]), .B(n385), .Z(n386) );
  XOR U321 ( .A(n392), .B(n393), .Z(n387) );
  XOR U322 ( .A(n394), .B(n385), .Z(n393) );
  XOR U323 ( .A(n395), .B(n396), .Z(n385) );
  NOR U324 ( .A(n397), .B(n398), .Z(n395) );
  AND U325 ( .A(b[0]), .B(a[108]), .Z(n394) );
  XOR U326 ( .A(n399), .B(n400), .Z(n392) );
  XOR U327 ( .A(n401), .B(n402), .Z(n400) );
  AND U328 ( .A(b[2]), .B(a[106]), .Z(n402) );
  AND U329 ( .A(a[105]), .B(b[3]), .Z(n401) );
  AND U330 ( .A(b[1]), .B(a[107]), .Z(n399) );
  XOR U331 ( .A(n398), .B(n397), .Z(swire[107]) );
  XOR U332 ( .A(sreg[235]), .B(n396), .Z(n397) );
  XOR U333 ( .A(n403), .B(n404), .Z(n398) );
  XOR U334 ( .A(n405), .B(n396), .Z(n404) );
  XOR U335 ( .A(n406), .B(n407), .Z(n396) );
  NOR U336 ( .A(n408), .B(n409), .Z(n406) );
  AND U337 ( .A(b[0]), .B(a[107]), .Z(n405) );
  XOR U338 ( .A(n410), .B(n411), .Z(n403) );
  XOR U339 ( .A(n412), .B(n413), .Z(n411) );
  AND U340 ( .A(b[2]), .B(a[105]), .Z(n413) );
  AND U341 ( .A(a[104]), .B(b[3]), .Z(n412) );
  AND U342 ( .A(b[1]), .B(a[106]), .Z(n410) );
  XOR U343 ( .A(n409), .B(n408), .Z(swire[106]) );
  XOR U344 ( .A(sreg[234]), .B(n407), .Z(n408) );
  XOR U345 ( .A(n414), .B(n415), .Z(n409) );
  XOR U346 ( .A(n416), .B(n407), .Z(n415) );
  XOR U347 ( .A(n417), .B(n418), .Z(n407) );
  NOR U348 ( .A(n419), .B(n420), .Z(n417) );
  AND U349 ( .A(b[0]), .B(a[106]), .Z(n416) );
  XOR U350 ( .A(n421), .B(n422), .Z(n414) );
  XOR U351 ( .A(n423), .B(n424), .Z(n422) );
  AND U352 ( .A(b[2]), .B(a[104]), .Z(n424) );
  AND U353 ( .A(a[103]), .B(b[3]), .Z(n423) );
  AND U354 ( .A(b[1]), .B(a[105]), .Z(n421) );
  XOR U355 ( .A(n420), .B(n419), .Z(swire[105]) );
  XOR U356 ( .A(sreg[233]), .B(n418), .Z(n419) );
  XOR U357 ( .A(n425), .B(n426), .Z(n420) );
  XOR U358 ( .A(n427), .B(n418), .Z(n426) );
  XOR U359 ( .A(n428), .B(n429), .Z(n418) );
  NOR U360 ( .A(n430), .B(n431), .Z(n428) );
  AND U361 ( .A(b[0]), .B(a[105]), .Z(n427) );
  XOR U362 ( .A(n432), .B(n433), .Z(n425) );
  XOR U363 ( .A(n434), .B(n435), .Z(n433) );
  AND U364 ( .A(b[2]), .B(a[103]), .Z(n435) );
  AND U365 ( .A(a[102]), .B(b[3]), .Z(n434) );
  AND U366 ( .A(b[1]), .B(a[104]), .Z(n432) );
  XOR U367 ( .A(n431), .B(n430), .Z(swire[104]) );
  XOR U368 ( .A(sreg[232]), .B(n429), .Z(n430) );
  XOR U369 ( .A(n436), .B(n437), .Z(n431) );
  XOR U370 ( .A(n438), .B(n429), .Z(n437) );
  XOR U371 ( .A(n439), .B(n440), .Z(n429) );
  NOR U372 ( .A(n441), .B(n442), .Z(n439) );
  AND U373 ( .A(b[0]), .B(a[104]), .Z(n438) );
  XOR U374 ( .A(n443), .B(n444), .Z(n436) );
  XOR U375 ( .A(n445), .B(n446), .Z(n444) );
  AND U376 ( .A(b[2]), .B(a[102]), .Z(n446) );
  AND U377 ( .A(a[101]), .B(b[3]), .Z(n445) );
  AND U378 ( .A(b[1]), .B(a[103]), .Z(n443) );
  XOR U379 ( .A(n442), .B(n441), .Z(swire[103]) );
  XOR U380 ( .A(sreg[231]), .B(n440), .Z(n441) );
  XOR U381 ( .A(n447), .B(n448), .Z(n442) );
  XOR U382 ( .A(n449), .B(n440), .Z(n448) );
  XOR U383 ( .A(n450), .B(n451), .Z(n440) );
  NOR U384 ( .A(n452), .B(n453), .Z(n450) );
  AND U385 ( .A(b[0]), .B(a[103]), .Z(n449) );
  XOR U386 ( .A(n454), .B(n455), .Z(n447) );
  XOR U387 ( .A(n456), .B(n457), .Z(n455) );
  AND U388 ( .A(b[2]), .B(a[101]), .Z(n457) );
  AND U389 ( .A(a[100]), .B(b[3]), .Z(n456) );
  AND U390 ( .A(b[1]), .B(a[102]), .Z(n454) );
  XOR U391 ( .A(n453), .B(n452), .Z(swire[102]) );
  XOR U392 ( .A(sreg[230]), .B(n451), .Z(n452) );
  XOR U393 ( .A(n458), .B(n459), .Z(n453) );
  XOR U394 ( .A(n460), .B(n451), .Z(n459) );
  XOR U395 ( .A(n461), .B(n462), .Z(n451) );
  NOR U396 ( .A(n463), .B(n464), .Z(n461) );
  AND U397 ( .A(b[0]), .B(a[102]), .Z(n460) );
  XOR U398 ( .A(n465), .B(n466), .Z(n458) );
  XOR U399 ( .A(n467), .B(n468), .Z(n466) );
  AND U400 ( .A(b[2]), .B(a[100]), .Z(n468) );
  AND U401 ( .A(a[99]), .B(b[3]), .Z(n467) );
  AND U402 ( .A(b[1]), .B(a[101]), .Z(n465) );
  XOR U403 ( .A(n464), .B(n463), .Z(swire[101]) );
  XOR U404 ( .A(sreg[229]), .B(n462), .Z(n463) );
  XOR U405 ( .A(n469), .B(n470), .Z(n464) );
  XOR U406 ( .A(n471), .B(n462), .Z(n470) );
  XOR U407 ( .A(n472), .B(n473), .Z(n462) );
  NOR U408 ( .A(n474), .B(n475), .Z(n472) );
  AND U409 ( .A(b[0]), .B(a[101]), .Z(n471) );
  XOR U410 ( .A(n476), .B(n477), .Z(n469) );
  XOR U411 ( .A(n478), .B(n479), .Z(n477) );
  AND U412 ( .A(b[2]), .B(a[99]), .Z(n479) );
  AND U413 ( .A(a[98]), .B(b[3]), .Z(n478) );
  AND U414 ( .A(b[1]), .B(a[100]), .Z(n476) );
  XOR U415 ( .A(n475), .B(n474), .Z(swire[100]) );
  XOR U416 ( .A(sreg[228]), .B(n473), .Z(n474) );
  XOR U417 ( .A(n480), .B(n481), .Z(n475) );
  XOR U418 ( .A(n482), .B(n473), .Z(n481) );
  XOR U419 ( .A(n483), .B(n484), .Z(n473) );
  NOR U420 ( .A(n4), .B(n3), .Z(n483) );
  XOR U421 ( .A(sreg[227]), .B(n484), .Z(n3) );
  XOR U422 ( .A(n485), .B(n486), .Z(n4) );
  XOR U423 ( .A(n487), .B(n484), .Z(n486) );
  XOR U424 ( .A(n488), .B(n489), .Z(n484) );
  NOR U425 ( .A(n6), .B(n5), .Z(n488) );
  XOR U426 ( .A(n490), .B(n491), .Z(n5) );
  XOR U427 ( .A(n492), .B(n489), .Z(n491) );
  AND U428 ( .A(b[0]), .B(a[98]), .Z(n492) );
  XOR U429 ( .A(n493), .B(n494), .Z(n490) );
  XOR U430 ( .A(n495), .B(n496), .Z(n494) );
  AND U431 ( .A(a[95]), .B(b[3]), .Z(n496) );
  AND U432 ( .A(b[1]), .B(a[97]), .Z(n495) );
  AND U433 ( .A(b[2]), .B(a[96]), .Z(n493) );
  XOR U434 ( .A(sreg[226]), .B(n489), .Z(n6) );
  XOR U435 ( .A(n497), .B(n498), .Z(n489) );
  NOR U436 ( .A(n8), .B(n7), .Z(n497) );
  XOR U437 ( .A(n499), .B(n500), .Z(n7) );
  XOR U438 ( .A(n501), .B(n498), .Z(n500) );
  AND U439 ( .A(b[0]), .B(a[97]), .Z(n501) );
  XOR U440 ( .A(n502), .B(n503), .Z(n499) );
  XOR U441 ( .A(n504), .B(n505), .Z(n503) );
  AND U442 ( .A(b[2]), .B(a[95]), .Z(n505) );
  AND U443 ( .A(a[94]), .B(b[3]), .Z(n504) );
  AND U444 ( .A(b[1]), .B(a[96]), .Z(n502) );
  XOR U445 ( .A(sreg[225]), .B(n498), .Z(n8) );
  XOR U446 ( .A(n506), .B(n507), .Z(n498) );
  NOR U447 ( .A(n10), .B(n9), .Z(n506) );
  XOR U448 ( .A(n508), .B(n509), .Z(n9) );
  XOR U449 ( .A(n510), .B(n507), .Z(n509) );
  AND U450 ( .A(b[0]), .B(a[96]), .Z(n510) );
  XOR U451 ( .A(n511), .B(n512), .Z(n508) );
  XOR U452 ( .A(n513), .B(n514), .Z(n512) );
  AND U453 ( .A(a[93]), .B(b[3]), .Z(n514) );
  AND U454 ( .A(b[2]), .B(a[94]), .Z(n513) );
  AND U455 ( .A(b[1]), .B(a[95]), .Z(n511) );
  XOR U456 ( .A(sreg[224]), .B(n507), .Z(n10) );
  XOR U457 ( .A(n515), .B(n516), .Z(n507) );
  NOR U458 ( .A(n12), .B(n11), .Z(n515) );
  XOR U459 ( .A(n517), .B(n518), .Z(n11) );
  XOR U460 ( .A(n519), .B(n516), .Z(n518) );
  AND U461 ( .A(b[0]), .B(a[95]), .Z(n519) );
  XOR U462 ( .A(n520), .B(n521), .Z(n517) );
  XOR U463 ( .A(n522), .B(n523), .Z(n521) );
  AND U464 ( .A(a[92]), .B(b[3]), .Z(n523) );
  AND U465 ( .A(b[1]), .B(a[94]), .Z(n522) );
  AND U466 ( .A(b[2]), .B(a[93]), .Z(n520) );
  XOR U467 ( .A(sreg[223]), .B(n516), .Z(n12) );
  XOR U468 ( .A(n524), .B(n525), .Z(n516) );
  NOR U469 ( .A(n14), .B(n13), .Z(n524) );
  XOR U470 ( .A(n526), .B(n527), .Z(n13) );
  XOR U471 ( .A(n528), .B(n525), .Z(n527) );
  AND U472 ( .A(b[0]), .B(a[94]), .Z(n528) );
  XOR U473 ( .A(n529), .B(n530), .Z(n526) );
  XOR U474 ( .A(n531), .B(n532), .Z(n530) );
  AND U475 ( .A(b[2]), .B(a[92]), .Z(n532) );
  AND U476 ( .A(a[91]), .B(b[3]), .Z(n531) );
  AND U477 ( .A(b[1]), .B(a[93]), .Z(n529) );
  XOR U478 ( .A(sreg[222]), .B(n525), .Z(n14) );
  XOR U479 ( .A(n533), .B(n534), .Z(n525) );
  NOR U480 ( .A(n16), .B(n15), .Z(n533) );
  XOR U481 ( .A(n535), .B(n536), .Z(n15) );
  XOR U482 ( .A(n537), .B(n534), .Z(n536) );
  AND U483 ( .A(b[0]), .B(a[93]), .Z(n537) );
  XOR U484 ( .A(n538), .B(n539), .Z(n535) );
  XOR U485 ( .A(n540), .B(n541), .Z(n539) );
  AND U486 ( .A(a[90]), .B(b[3]), .Z(n541) );
  AND U487 ( .A(b[2]), .B(a[91]), .Z(n540) );
  AND U488 ( .A(b[1]), .B(a[92]), .Z(n538) );
  XOR U489 ( .A(sreg[221]), .B(n534), .Z(n16) );
  XOR U490 ( .A(n542), .B(n543), .Z(n534) );
  NOR U491 ( .A(n18), .B(n17), .Z(n542) );
  XOR U492 ( .A(n544), .B(n545), .Z(n17) );
  XOR U493 ( .A(n546), .B(n543), .Z(n545) );
  AND U494 ( .A(b[0]), .B(a[92]), .Z(n546) );
  XOR U495 ( .A(n547), .B(n548), .Z(n544) );
  XOR U496 ( .A(n549), .B(n550), .Z(n548) );
  AND U497 ( .A(a[89]), .B(b[3]), .Z(n550) );
  AND U498 ( .A(b[1]), .B(a[91]), .Z(n549) );
  AND U499 ( .A(b[2]), .B(a[90]), .Z(n547) );
  XOR U500 ( .A(sreg[220]), .B(n543), .Z(n18) );
  XOR U501 ( .A(n551), .B(n552), .Z(n543) );
  NOR U502 ( .A(n20), .B(n19), .Z(n551) );
  XOR U503 ( .A(n553), .B(n554), .Z(n19) );
  XOR U504 ( .A(n555), .B(n552), .Z(n554) );
  AND U505 ( .A(b[0]), .B(a[91]), .Z(n555) );
  XOR U506 ( .A(n556), .B(n557), .Z(n553) );
  XOR U507 ( .A(n558), .B(n559), .Z(n557) );
  AND U508 ( .A(b[2]), .B(a[89]), .Z(n559) );
  AND U509 ( .A(a[88]), .B(b[3]), .Z(n558) );
  AND U510 ( .A(b[1]), .B(a[90]), .Z(n556) );
  XOR U511 ( .A(sreg[219]), .B(n552), .Z(n20) );
  XOR U512 ( .A(n560), .B(n561), .Z(n552) );
  NOR U513 ( .A(n22), .B(n21), .Z(n560) );
  XOR U514 ( .A(n562), .B(n563), .Z(n21) );
  XOR U515 ( .A(n564), .B(n561), .Z(n563) );
  AND U516 ( .A(b[0]), .B(a[90]), .Z(n564) );
  XOR U517 ( .A(n565), .B(n566), .Z(n562) );
  XOR U518 ( .A(n567), .B(n568), .Z(n566) );
  AND U519 ( .A(a[87]), .B(b[3]), .Z(n568) );
  AND U520 ( .A(b[2]), .B(a[88]), .Z(n567) );
  AND U521 ( .A(b[1]), .B(a[89]), .Z(n565) );
  XOR U522 ( .A(sreg[218]), .B(n561), .Z(n22) );
  XOR U523 ( .A(n569), .B(n570), .Z(n561) );
  NOR U524 ( .A(n26), .B(n25), .Z(n569) );
  XOR U525 ( .A(n571), .B(n572), .Z(n25) );
  XOR U526 ( .A(n573), .B(n570), .Z(n572) );
  AND U527 ( .A(b[0]), .B(a[89]), .Z(n573) );
  XOR U528 ( .A(n574), .B(n575), .Z(n571) );
  XOR U529 ( .A(n576), .B(n577), .Z(n575) );
  AND U530 ( .A(a[86]), .B(b[3]), .Z(n577) );
  AND U531 ( .A(b[1]), .B(a[88]), .Z(n576) );
  AND U532 ( .A(b[2]), .B(a[87]), .Z(n574) );
  XOR U533 ( .A(sreg[217]), .B(n570), .Z(n26) );
  XOR U534 ( .A(n578), .B(n579), .Z(n570) );
  NOR U535 ( .A(n28), .B(n27), .Z(n578) );
  XOR U536 ( .A(n580), .B(n581), .Z(n27) );
  XOR U537 ( .A(n582), .B(n579), .Z(n581) );
  AND U538 ( .A(b[0]), .B(a[88]), .Z(n582) );
  XOR U539 ( .A(n583), .B(n584), .Z(n580) );
  XOR U540 ( .A(n585), .B(n586), .Z(n584) );
  AND U541 ( .A(b[2]), .B(a[86]), .Z(n586) );
  AND U542 ( .A(a[85]), .B(b[3]), .Z(n585) );
  AND U543 ( .A(b[1]), .B(a[87]), .Z(n583) );
  XOR U544 ( .A(sreg[216]), .B(n579), .Z(n28) );
  XOR U545 ( .A(n587), .B(n588), .Z(n579) );
  NOR U546 ( .A(n30), .B(n29), .Z(n587) );
  XOR U547 ( .A(n589), .B(n590), .Z(n29) );
  XOR U548 ( .A(n591), .B(n588), .Z(n590) );
  AND U549 ( .A(b[0]), .B(a[87]), .Z(n591) );
  XOR U550 ( .A(n592), .B(n593), .Z(n589) );
  XOR U551 ( .A(n594), .B(n595), .Z(n593) );
  AND U552 ( .A(a[84]), .B(b[3]), .Z(n595) );
  AND U553 ( .A(b[2]), .B(a[85]), .Z(n594) );
  AND U554 ( .A(b[1]), .B(a[86]), .Z(n592) );
  XOR U555 ( .A(sreg[215]), .B(n588), .Z(n30) );
  XOR U556 ( .A(n596), .B(n597), .Z(n588) );
  NOR U557 ( .A(n32), .B(n31), .Z(n596) );
  XOR U558 ( .A(n598), .B(n599), .Z(n31) );
  XOR U559 ( .A(n600), .B(n597), .Z(n599) );
  AND U560 ( .A(b[0]), .B(a[86]), .Z(n600) );
  XOR U561 ( .A(n601), .B(n602), .Z(n598) );
  XOR U562 ( .A(n603), .B(n604), .Z(n602) );
  AND U563 ( .A(a[83]), .B(b[3]), .Z(n604) );
  AND U564 ( .A(b[1]), .B(a[85]), .Z(n603) );
  AND U565 ( .A(b[2]), .B(a[84]), .Z(n601) );
  XOR U566 ( .A(sreg[214]), .B(n597), .Z(n32) );
  XOR U567 ( .A(n605), .B(n606), .Z(n597) );
  NOR U568 ( .A(n34), .B(n33), .Z(n605) );
  XOR U569 ( .A(n607), .B(n608), .Z(n33) );
  XOR U570 ( .A(n609), .B(n606), .Z(n608) );
  AND U571 ( .A(b[0]), .B(a[85]), .Z(n609) );
  XOR U572 ( .A(n610), .B(n611), .Z(n607) );
  XOR U573 ( .A(n612), .B(n613), .Z(n611) );
  AND U574 ( .A(b[2]), .B(a[83]), .Z(n613) );
  AND U575 ( .A(a[82]), .B(b[3]), .Z(n612) );
  AND U576 ( .A(b[1]), .B(a[84]), .Z(n610) );
  XOR U577 ( .A(sreg[213]), .B(n606), .Z(n34) );
  XOR U578 ( .A(n614), .B(n615), .Z(n606) );
  NOR U579 ( .A(n36), .B(n35), .Z(n614) );
  XOR U580 ( .A(n616), .B(n617), .Z(n35) );
  XOR U581 ( .A(n618), .B(n615), .Z(n617) );
  AND U582 ( .A(b[0]), .B(a[84]), .Z(n618) );
  XOR U583 ( .A(n619), .B(n620), .Z(n616) );
  XOR U584 ( .A(n621), .B(n622), .Z(n620) );
  AND U585 ( .A(a[81]), .B(b[3]), .Z(n622) );
  AND U586 ( .A(b[2]), .B(a[82]), .Z(n621) );
  AND U587 ( .A(b[1]), .B(a[83]), .Z(n619) );
  XOR U588 ( .A(sreg[212]), .B(n615), .Z(n36) );
  XOR U589 ( .A(n623), .B(n624), .Z(n615) );
  NOR U590 ( .A(n38), .B(n37), .Z(n623) );
  XOR U591 ( .A(n625), .B(n626), .Z(n37) );
  XOR U592 ( .A(n627), .B(n624), .Z(n626) );
  AND U593 ( .A(b[0]), .B(a[83]), .Z(n627) );
  XOR U594 ( .A(n628), .B(n629), .Z(n625) );
  XOR U595 ( .A(n630), .B(n631), .Z(n629) );
  AND U596 ( .A(a[80]), .B(b[3]), .Z(n631) );
  AND U597 ( .A(b[1]), .B(a[82]), .Z(n630) );
  AND U598 ( .A(b[2]), .B(a[81]), .Z(n628) );
  XOR U599 ( .A(sreg[211]), .B(n624), .Z(n38) );
  XOR U600 ( .A(n632), .B(n633), .Z(n624) );
  NOR U601 ( .A(n40), .B(n39), .Z(n632) );
  XOR U602 ( .A(n634), .B(n635), .Z(n39) );
  XOR U603 ( .A(n636), .B(n633), .Z(n635) );
  AND U604 ( .A(b[0]), .B(a[82]), .Z(n636) );
  XOR U605 ( .A(n637), .B(n638), .Z(n634) );
  XOR U606 ( .A(n639), .B(n640), .Z(n638) );
  AND U607 ( .A(b[2]), .B(a[80]), .Z(n640) );
  AND U608 ( .A(a[79]), .B(b[3]), .Z(n639) );
  AND U609 ( .A(b[1]), .B(a[81]), .Z(n637) );
  XOR U610 ( .A(sreg[210]), .B(n633), .Z(n40) );
  XOR U611 ( .A(n641), .B(n642), .Z(n633) );
  NOR U612 ( .A(n42), .B(n41), .Z(n641) );
  XOR U613 ( .A(n643), .B(n644), .Z(n41) );
  XOR U614 ( .A(n645), .B(n642), .Z(n644) );
  AND U615 ( .A(b[0]), .B(a[81]), .Z(n645) );
  XOR U616 ( .A(n646), .B(n647), .Z(n643) );
  XOR U617 ( .A(n648), .B(n649), .Z(n647) );
  AND U618 ( .A(a[78]), .B(b[3]), .Z(n649) );
  AND U619 ( .A(b[2]), .B(a[79]), .Z(n648) );
  AND U620 ( .A(b[1]), .B(a[80]), .Z(n646) );
  XOR U621 ( .A(sreg[209]), .B(n642), .Z(n42) );
  XOR U622 ( .A(n650), .B(n651), .Z(n642) );
  NOR U623 ( .A(n44), .B(n43), .Z(n650) );
  XOR U624 ( .A(n652), .B(n653), .Z(n43) );
  XOR U625 ( .A(n654), .B(n651), .Z(n653) );
  AND U626 ( .A(b[0]), .B(a[80]), .Z(n654) );
  XOR U627 ( .A(n655), .B(n656), .Z(n652) );
  XOR U628 ( .A(n657), .B(n658), .Z(n656) );
  AND U629 ( .A(a[77]), .B(b[3]), .Z(n658) );
  AND U630 ( .A(b[1]), .B(a[79]), .Z(n657) );
  AND U631 ( .A(b[2]), .B(a[78]), .Z(n655) );
  XOR U632 ( .A(sreg[208]), .B(n651), .Z(n44) );
  XOR U633 ( .A(n659), .B(n660), .Z(n651) );
  NOR U634 ( .A(n48), .B(n47), .Z(n659) );
  XOR U635 ( .A(n661), .B(n662), .Z(n47) );
  XOR U636 ( .A(n663), .B(n660), .Z(n662) );
  AND U637 ( .A(b[0]), .B(a[79]), .Z(n663) );
  XOR U638 ( .A(n664), .B(n665), .Z(n661) );
  XOR U639 ( .A(n666), .B(n667), .Z(n665) );
  AND U640 ( .A(b[2]), .B(a[77]), .Z(n667) );
  AND U641 ( .A(a[76]), .B(b[3]), .Z(n666) );
  AND U642 ( .A(b[1]), .B(a[78]), .Z(n664) );
  XOR U643 ( .A(sreg[207]), .B(n660), .Z(n48) );
  XOR U644 ( .A(n668), .B(n669), .Z(n660) );
  NOR U645 ( .A(n50), .B(n49), .Z(n668) );
  XOR U646 ( .A(n670), .B(n671), .Z(n49) );
  XOR U647 ( .A(n672), .B(n669), .Z(n671) );
  AND U648 ( .A(b[0]), .B(a[78]), .Z(n672) );
  XOR U649 ( .A(n673), .B(n674), .Z(n670) );
  XOR U650 ( .A(n675), .B(n676), .Z(n674) );
  AND U651 ( .A(a[75]), .B(b[3]), .Z(n676) );
  AND U652 ( .A(b[2]), .B(a[76]), .Z(n675) );
  AND U653 ( .A(b[1]), .B(a[77]), .Z(n673) );
  XOR U654 ( .A(sreg[206]), .B(n669), .Z(n50) );
  XOR U655 ( .A(n677), .B(n678), .Z(n669) );
  NOR U656 ( .A(n52), .B(n51), .Z(n677) );
  XOR U657 ( .A(n679), .B(n680), .Z(n51) );
  XOR U658 ( .A(n681), .B(n678), .Z(n680) );
  AND U659 ( .A(b[0]), .B(a[77]), .Z(n681) );
  XOR U660 ( .A(n682), .B(n683), .Z(n679) );
  XOR U661 ( .A(n684), .B(n685), .Z(n683) );
  AND U662 ( .A(a[74]), .B(b[3]), .Z(n685) );
  AND U663 ( .A(b[1]), .B(a[76]), .Z(n684) );
  AND U664 ( .A(b[2]), .B(a[75]), .Z(n682) );
  XOR U665 ( .A(sreg[205]), .B(n678), .Z(n52) );
  XOR U666 ( .A(n686), .B(n687), .Z(n678) );
  NOR U667 ( .A(n54), .B(n53), .Z(n686) );
  XOR U668 ( .A(n688), .B(n689), .Z(n53) );
  XOR U669 ( .A(n690), .B(n687), .Z(n689) );
  AND U670 ( .A(b[0]), .B(a[76]), .Z(n690) );
  XOR U671 ( .A(n691), .B(n692), .Z(n688) );
  XOR U672 ( .A(n693), .B(n694), .Z(n692) );
  AND U673 ( .A(b[2]), .B(a[74]), .Z(n694) );
  AND U674 ( .A(a[73]), .B(b[3]), .Z(n693) );
  AND U675 ( .A(b[1]), .B(a[75]), .Z(n691) );
  XOR U676 ( .A(sreg[204]), .B(n687), .Z(n54) );
  XOR U677 ( .A(n695), .B(n696), .Z(n687) );
  NOR U678 ( .A(n56), .B(n55), .Z(n695) );
  XOR U679 ( .A(n697), .B(n698), .Z(n55) );
  XOR U680 ( .A(n699), .B(n696), .Z(n698) );
  AND U681 ( .A(b[0]), .B(a[75]), .Z(n699) );
  XOR U682 ( .A(n700), .B(n701), .Z(n697) );
  XOR U683 ( .A(n702), .B(n703), .Z(n701) );
  AND U684 ( .A(a[72]), .B(b[3]), .Z(n703) );
  AND U685 ( .A(b[2]), .B(a[73]), .Z(n702) );
  AND U686 ( .A(b[1]), .B(a[74]), .Z(n700) );
  XOR U687 ( .A(sreg[203]), .B(n696), .Z(n56) );
  XOR U688 ( .A(n704), .B(n705), .Z(n696) );
  NOR U689 ( .A(n58), .B(n57), .Z(n704) );
  XOR U690 ( .A(n706), .B(n707), .Z(n57) );
  XOR U691 ( .A(n708), .B(n705), .Z(n707) );
  AND U692 ( .A(b[0]), .B(a[74]), .Z(n708) );
  XOR U693 ( .A(n709), .B(n710), .Z(n706) );
  XOR U694 ( .A(n711), .B(n712), .Z(n710) );
  AND U695 ( .A(a[71]), .B(b[3]), .Z(n712) );
  AND U696 ( .A(b[1]), .B(a[73]), .Z(n711) );
  AND U697 ( .A(b[2]), .B(a[72]), .Z(n709) );
  XOR U698 ( .A(sreg[202]), .B(n705), .Z(n58) );
  XOR U699 ( .A(n713), .B(n714), .Z(n705) );
  NOR U700 ( .A(n60), .B(n59), .Z(n713) );
  XOR U701 ( .A(n715), .B(n716), .Z(n59) );
  XOR U702 ( .A(n717), .B(n714), .Z(n716) );
  AND U703 ( .A(b[0]), .B(a[73]), .Z(n717) );
  XOR U704 ( .A(n718), .B(n719), .Z(n715) );
  XOR U705 ( .A(n720), .B(n721), .Z(n719) );
  AND U706 ( .A(b[2]), .B(a[71]), .Z(n721) );
  AND U707 ( .A(a[70]), .B(b[3]), .Z(n720) );
  AND U708 ( .A(b[1]), .B(a[72]), .Z(n718) );
  XOR U709 ( .A(sreg[201]), .B(n714), .Z(n60) );
  XOR U710 ( .A(n722), .B(n723), .Z(n714) );
  NOR U711 ( .A(n62), .B(n61), .Z(n722) );
  XOR U712 ( .A(n724), .B(n725), .Z(n61) );
  XOR U713 ( .A(n726), .B(n723), .Z(n725) );
  AND U714 ( .A(b[0]), .B(a[72]), .Z(n726) );
  XOR U715 ( .A(n727), .B(n728), .Z(n724) );
  XOR U716 ( .A(n729), .B(n730), .Z(n728) );
  AND U717 ( .A(a[69]), .B(b[3]), .Z(n730) );
  AND U718 ( .A(b[2]), .B(a[70]), .Z(n729) );
  AND U719 ( .A(b[1]), .B(a[71]), .Z(n727) );
  XOR U720 ( .A(sreg[200]), .B(n723), .Z(n62) );
  XOR U721 ( .A(n731), .B(n732), .Z(n723) );
  NOR U722 ( .A(n64), .B(n63), .Z(n731) );
  XOR U723 ( .A(n733), .B(n734), .Z(n63) );
  XOR U724 ( .A(n735), .B(n732), .Z(n734) );
  AND U725 ( .A(b[0]), .B(a[71]), .Z(n735) );
  XOR U726 ( .A(n736), .B(n737), .Z(n733) );
  XOR U727 ( .A(n738), .B(n739), .Z(n737) );
  AND U728 ( .A(a[68]), .B(b[3]), .Z(n739) );
  AND U729 ( .A(b[1]), .B(a[70]), .Z(n738) );
  AND U730 ( .A(b[2]), .B(a[69]), .Z(n736) );
  XOR U731 ( .A(sreg[199]), .B(n732), .Z(n64) );
  XOR U732 ( .A(n740), .B(n741), .Z(n732) );
  NOR U733 ( .A(n66), .B(n65), .Z(n740) );
  XOR U734 ( .A(n742), .B(n743), .Z(n65) );
  XOR U735 ( .A(n744), .B(n741), .Z(n743) );
  AND U736 ( .A(b[0]), .B(a[70]), .Z(n744) );
  XOR U737 ( .A(n745), .B(n746), .Z(n742) );
  XOR U738 ( .A(n747), .B(n748), .Z(n746) );
  AND U739 ( .A(b[2]), .B(a[68]), .Z(n748) );
  AND U740 ( .A(a[67]), .B(b[3]), .Z(n747) );
  AND U741 ( .A(b[1]), .B(a[69]), .Z(n745) );
  XOR U742 ( .A(sreg[198]), .B(n741), .Z(n66) );
  XOR U743 ( .A(n749), .B(n750), .Z(n741) );
  NOR U744 ( .A(n70), .B(n69), .Z(n749) );
  XOR U745 ( .A(n751), .B(n752), .Z(n69) );
  XOR U746 ( .A(n753), .B(n750), .Z(n752) );
  AND U747 ( .A(b[0]), .B(a[69]), .Z(n753) );
  XOR U748 ( .A(n754), .B(n755), .Z(n751) );
  XOR U749 ( .A(n756), .B(n757), .Z(n755) );
  AND U750 ( .A(a[66]), .B(b[3]), .Z(n757) );
  AND U751 ( .A(b[2]), .B(a[67]), .Z(n756) );
  AND U752 ( .A(b[1]), .B(a[68]), .Z(n754) );
  XOR U753 ( .A(sreg[197]), .B(n750), .Z(n70) );
  XOR U754 ( .A(n758), .B(n759), .Z(n750) );
  NOR U755 ( .A(n72), .B(n71), .Z(n758) );
  XOR U756 ( .A(n760), .B(n761), .Z(n71) );
  XOR U757 ( .A(n762), .B(n759), .Z(n761) );
  AND U758 ( .A(b[0]), .B(a[68]), .Z(n762) );
  XOR U759 ( .A(n763), .B(n764), .Z(n760) );
  XOR U760 ( .A(n765), .B(n766), .Z(n764) );
  AND U761 ( .A(a[65]), .B(b[3]), .Z(n766) );
  AND U762 ( .A(b[1]), .B(a[67]), .Z(n765) );
  AND U763 ( .A(b[2]), .B(a[66]), .Z(n763) );
  XOR U764 ( .A(sreg[196]), .B(n759), .Z(n72) );
  XOR U765 ( .A(n767), .B(n768), .Z(n759) );
  NOR U766 ( .A(n74), .B(n73), .Z(n767) );
  XOR U767 ( .A(n769), .B(n770), .Z(n73) );
  XOR U768 ( .A(n771), .B(n768), .Z(n770) );
  AND U769 ( .A(b[0]), .B(a[67]), .Z(n771) );
  XOR U770 ( .A(n772), .B(n773), .Z(n769) );
  XOR U771 ( .A(n774), .B(n775), .Z(n773) );
  AND U772 ( .A(b[2]), .B(a[65]), .Z(n775) );
  AND U773 ( .A(a[64]), .B(b[3]), .Z(n774) );
  AND U774 ( .A(b[1]), .B(a[66]), .Z(n772) );
  XOR U775 ( .A(sreg[195]), .B(n768), .Z(n74) );
  XOR U776 ( .A(n776), .B(n777), .Z(n768) );
  NOR U777 ( .A(n76), .B(n75), .Z(n776) );
  XOR U778 ( .A(n778), .B(n779), .Z(n75) );
  XOR U779 ( .A(n780), .B(n777), .Z(n779) );
  AND U780 ( .A(b[0]), .B(a[66]), .Z(n780) );
  XOR U781 ( .A(n781), .B(n782), .Z(n778) );
  XOR U782 ( .A(n783), .B(n784), .Z(n782) );
  AND U783 ( .A(a[63]), .B(b[3]), .Z(n784) );
  AND U784 ( .A(b[2]), .B(a[64]), .Z(n783) );
  AND U785 ( .A(b[1]), .B(a[65]), .Z(n781) );
  XOR U786 ( .A(sreg[194]), .B(n777), .Z(n76) );
  XOR U787 ( .A(n785), .B(n786), .Z(n777) );
  NOR U788 ( .A(n78), .B(n77), .Z(n785) );
  XOR U789 ( .A(n787), .B(n788), .Z(n77) );
  XOR U790 ( .A(n789), .B(n786), .Z(n788) );
  AND U791 ( .A(b[0]), .B(a[65]), .Z(n789) );
  XOR U792 ( .A(n790), .B(n791), .Z(n787) );
  XOR U793 ( .A(n792), .B(n793), .Z(n791) );
  AND U794 ( .A(a[62]), .B(b[3]), .Z(n793) );
  AND U795 ( .A(b[1]), .B(a[64]), .Z(n792) );
  AND U796 ( .A(b[2]), .B(a[63]), .Z(n790) );
  XOR U797 ( .A(sreg[193]), .B(n786), .Z(n78) );
  XOR U798 ( .A(n794), .B(n795), .Z(n786) );
  NOR U799 ( .A(n80), .B(n79), .Z(n794) );
  XOR U800 ( .A(n796), .B(n797), .Z(n79) );
  XOR U801 ( .A(n798), .B(n795), .Z(n797) );
  AND U802 ( .A(b[0]), .B(a[64]), .Z(n798) );
  XOR U803 ( .A(n799), .B(n800), .Z(n796) );
  XOR U804 ( .A(n801), .B(n802), .Z(n800) );
  AND U805 ( .A(b[2]), .B(a[62]), .Z(n802) );
  AND U806 ( .A(a[61]), .B(b[3]), .Z(n801) );
  AND U807 ( .A(b[1]), .B(a[63]), .Z(n799) );
  XOR U808 ( .A(sreg[192]), .B(n795), .Z(n80) );
  XOR U809 ( .A(n803), .B(n804), .Z(n795) );
  NOR U810 ( .A(n82), .B(n81), .Z(n803) );
  XOR U811 ( .A(n805), .B(n806), .Z(n81) );
  XOR U812 ( .A(n807), .B(n804), .Z(n806) );
  AND U813 ( .A(b[0]), .B(a[63]), .Z(n807) );
  XOR U814 ( .A(n808), .B(n809), .Z(n805) );
  XOR U815 ( .A(n810), .B(n811), .Z(n809) );
  AND U816 ( .A(a[60]), .B(b[3]), .Z(n811) );
  AND U817 ( .A(b[2]), .B(a[61]), .Z(n810) );
  AND U818 ( .A(b[1]), .B(a[62]), .Z(n808) );
  XOR U819 ( .A(sreg[191]), .B(n804), .Z(n82) );
  XOR U820 ( .A(n812), .B(n813), .Z(n804) );
  NOR U821 ( .A(n84), .B(n83), .Z(n812) );
  XOR U822 ( .A(n814), .B(n815), .Z(n83) );
  XOR U823 ( .A(n816), .B(n813), .Z(n815) );
  AND U824 ( .A(b[0]), .B(a[62]), .Z(n816) );
  XOR U825 ( .A(n817), .B(n818), .Z(n814) );
  XOR U826 ( .A(n819), .B(n820), .Z(n818) );
  AND U827 ( .A(a[59]), .B(b[3]), .Z(n820) );
  AND U828 ( .A(b[1]), .B(a[61]), .Z(n819) );
  AND U829 ( .A(b[2]), .B(a[60]), .Z(n817) );
  XOR U830 ( .A(sreg[190]), .B(n813), .Z(n84) );
  XOR U831 ( .A(n821), .B(n822), .Z(n813) );
  NOR U832 ( .A(n86), .B(n85), .Z(n821) );
  XOR U833 ( .A(n823), .B(n824), .Z(n85) );
  XOR U834 ( .A(n825), .B(n822), .Z(n824) );
  AND U835 ( .A(b[0]), .B(a[61]), .Z(n825) );
  XOR U836 ( .A(n826), .B(n827), .Z(n823) );
  XOR U837 ( .A(n828), .B(n829), .Z(n827) );
  AND U838 ( .A(b[2]), .B(a[59]), .Z(n829) );
  AND U839 ( .A(a[58]), .B(b[3]), .Z(n828) );
  AND U840 ( .A(b[1]), .B(a[60]), .Z(n826) );
  XOR U841 ( .A(sreg[189]), .B(n822), .Z(n86) );
  XOR U842 ( .A(n830), .B(n831), .Z(n822) );
  NOR U843 ( .A(n88), .B(n87), .Z(n830) );
  XOR U844 ( .A(n832), .B(n833), .Z(n87) );
  XOR U845 ( .A(n834), .B(n831), .Z(n833) );
  AND U846 ( .A(b[0]), .B(a[60]), .Z(n834) );
  XOR U847 ( .A(n835), .B(n836), .Z(n832) );
  XOR U848 ( .A(n837), .B(n838), .Z(n836) );
  AND U849 ( .A(a[57]), .B(b[3]), .Z(n838) );
  AND U850 ( .A(b[2]), .B(a[58]), .Z(n837) );
  AND U851 ( .A(b[1]), .B(a[59]), .Z(n835) );
  XOR U852 ( .A(sreg[188]), .B(n831), .Z(n88) );
  XOR U853 ( .A(n839), .B(n840), .Z(n831) );
  NOR U854 ( .A(n92), .B(n91), .Z(n839) );
  XOR U855 ( .A(n841), .B(n842), .Z(n91) );
  XOR U856 ( .A(n843), .B(n840), .Z(n842) );
  AND U857 ( .A(b[0]), .B(a[59]), .Z(n843) );
  XOR U858 ( .A(n844), .B(n845), .Z(n841) );
  XOR U859 ( .A(n846), .B(n847), .Z(n845) );
  AND U860 ( .A(a[56]), .B(b[3]), .Z(n847) );
  AND U861 ( .A(b[1]), .B(a[58]), .Z(n846) );
  AND U862 ( .A(b[2]), .B(a[57]), .Z(n844) );
  XOR U863 ( .A(sreg[187]), .B(n840), .Z(n92) );
  XOR U864 ( .A(n848), .B(n849), .Z(n840) );
  NOR U865 ( .A(n94), .B(n93), .Z(n848) );
  XOR U866 ( .A(n850), .B(n851), .Z(n93) );
  XOR U867 ( .A(n852), .B(n849), .Z(n851) );
  AND U868 ( .A(b[0]), .B(a[58]), .Z(n852) );
  XOR U869 ( .A(n853), .B(n854), .Z(n850) );
  XOR U870 ( .A(n855), .B(n856), .Z(n854) );
  AND U871 ( .A(b[2]), .B(a[56]), .Z(n856) );
  AND U872 ( .A(a[55]), .B(b[3]), .Z(n855) );
  AND U873 ( .A(b[1]), .B(a[57]), .Z(n853) );
  XOR U874 ( .A(sreg[186]), .B(n849), .Z(n94) );
  XOR U875 ( .A(n857), .B(n858), .Z(n849) );
  NOR U876 ( .A(n96), .B(n95), .Z(n857) );
  XOR U877 ( .A(n859), .B(n860), .Z(n95) );
  XOR U878 ( .A(n861), .B(n858), .Z(n860) );
  AND U879 ( .A(b[0]), .B(a[57]), .Z(n861) );
  XOR U880 ( .A(n862), .B(n863), .Z(n859) );
  XOR U881 ( .A(n864), .B(n865), .Z(n863) );
  AND U882 ( .A(a[54]), .B(b[3]), .Z(n865) );
  AND U883 ( .A(b[2]), .B(a[55]), .Z(n864) );
  AND U884 ( .A(b[1]), .B(a[56]), .Z(n862) );
  XOR U885 ( .A(sreg[185]), .B(n858), .Z(n96) );
  XOR U886 ( .A(n866), .B(n867), .Z(n858) );
  NOR U887 ( .A(n98), .B(n97), .Z(n866) );
  XOR U888 ( .A(n868), .B(n869), .Z(n97) );
  XOR U889 ( .A(n870), .B(n867), .Z(n869) );
  AND U890 ( .A(b[0]), .B(a[56]), .Z(n870) );
  XOR U891 ( .A(n871), .B(n872), .Z(n868) );
  XOR U892 ( .A(n873), .B(n874), .Z(n872) );
  AND U893 ( .A(a[53]), .B(b[3]), .Z(n874) );
  AND U894 ( .A(b[1]), .B(a[55]), .Z(n873) );
  AND U895 ( .A(b[2]), .B(a[54]), .Z(n871) );
  XOR U896 ( .A(sreg[184]), .B(n867), .Z(n98) );
  XOR U897 ( .A(n875), .B(n876), .Z(n867) );
  NOR U898 ( .A(n100), .B(n99), .Z(n875) );
  XOR U899 ( .A(n877), .B(n878), .Z(n99) );
  XOR U900 ( .A(n879), .B(n876), .Z(n878) );
  AND U901 ( .A(b[0]), .B(a[55]), .Z(n879) );
  XOR U902 ( .A(n880), .B(n881), .Z(n877) );
  XOR U903 ( .A(n882), .B(n883), .Z(n881) );
  AND U904 ( .A(b[2]), .B(a[53]), .Z(n883) );
  AND U905 ( .A(a[52]), .B(b[3]), .Z(n882) );
  AND U906 ( .A(b[1]), .B(a[54]), .Z(n880) );
  XOR U907 ( .A(sreg[183]), .B(n876), .Z(n100) );
  XOR U908 ( .A(n884), .B(n885), .Z(n876) );
  NOR U909 ( .A(n102), .B(n101), .Z(n884) );
  XOR U910 ( .A(n886), .B(n887), .Z(n101) );
  XOR U911 ( .A(n888), .B(n885), .Z(n887) );
  AND U912 ( .A(b[0]), .B(a[54]), .Z(n888) );
  XOR U913 ( .A(n889), .B(n890), .Z(n886) );
  XOR U914 ( .A(n891), .B(n892), .Z(n890) );
  AND U915 ( .A(a[51]), .B(b[3]), .Z(n892) );
  AND U916 ( .A(b[2]), .B(a[52]), .Z(n891) );
  AND U917 ( .A(b[1]), .B(a[53]), .Z(n889) );
  XOR U918 ( .A(sreg[182]), .B(n885), .Z(n102) );
  XOR U919 ( .A(n893), .B(n894), .Z(n885) );
  NOR U920 ( .A(n104), .B(n103), .Z(n893) );
  XOR U921 ( .A(n895), .B(n896), .Z(n103) );
  XOR U922 ( .A(n897), .B(n894), .Z(n896) );
  AND U923 ( .A(b[0]), .B(a[53]), .Z(n897) );
  XOR U924 ( .A(n898), .B(n899), .Z(n895) );
  XOR U925 ( .A(n900), .B(n901), .Z(n899) );
  AND U926 ( .A(a[50]), .B(b[3]), .Z(n901) );
  AND U927 ( .A(b[1]), .B(a[52]), .Z(n900) );
  AND U928 ( .A(b[2]), .B(a[51]), .Z(n898) );
  XOR U929 ( .A(sreg[181]), .B(n894), .Z(n104) );
  XOR U930 ( .A(n902), .B(n903), .Z(n894) );
  NOR U931 ( .A(n106), .B(n105), .Z(n902) );
  XOR U932 ( .A(n904), .B(n905), .Z(n105) );
  XOR U933 ( .A(n906), .B(n903), .Z(n905) );
  AND U934 ( .A(b[0]), .B(a[52]), .Z(n906) );
  XOR U935 ( .A(n907), .B(n908), .Z(n904) );
  XOR U936 ( .A(n909), .B(n910), .Z(n908) );
  AND U937 ( .A(b[2]), .B(a[50]), .Z(n910) );
  AND U938 ( .A(a[49]), .B(b[3]), .Z(n909) );
  AND U939 ( .A(b[1]), .B(a[51]), .Z(n907) );
  XOR U940 ( .A(sreg[180]), .B(n903), .Z(n106) );
  XOR U941 ( .A(n911), .B(n912), .Z(n903) );
  NOR U942 ( .A(n108), .B(n107), .Z(n911) );
  XOR U943 ( .A(n913), .B(n914), .Z(n107) );
  XOR U944 ( .A(n915), .B(n912), .Z(n914) );
  AND U945 ( .A(b[0]), .B(a[51]), .Z(n915) );
  XOR U946 ( .A(n916), .B(n917), .Z(n913) );
  XOR U947 ( .A(n918), .B(n919), .Z(n917) );
  AND U948 ( .A(a[48]), .B(b[3]), .Z(n919) );
  AND U949 ( .A(b[2]), .B(a[49]), .Z(n918) );
  AND U950 ( .A(b[1]), .B(a[50]), .Z(n916) );
  XOR U951 ( .A(sreg[179]), .B(n912), .Z(n108) );
  XOR U952 ( .A(n920), .B(n921), .Z(n912) );
  NOR U953 ( .A(n110), .B(n109), .Z(n920) );
  XOR U954 ( .A(n922), .B(n923), .Z(n109) );
  XOR U955 ( .A(n924), .B(n921), .Z(n923) );
  AND U956 ( .A(b[0]), .B(a[50]), .Z(n924) );
  XOR U957 ( .A(n925), .B(n926), .Z(n922) );
  XOR U958 ( .A(n927), .B(n928), .Z(n926) );
  AND U959 ( .A(a[47]), .B(b[3]), .Z(n928) );
  AND U960 ( .A(b[1]), .B(a[49]), .Z(n927) );
  AND U961 ( .A(b[2]), .B(a[48]), .Z(n925) );
  XOR U962 ( .A(sreg[178]), .B(n921), .Z(n110) );
  XOR U963 ( .A(n929), .B(n930), .Z(n921) );
  NOR U964 ( .A(n114), .B(n113), .Z(n929) );
  XOR U965 ( .A(n931), .B(n932), .Z(n113) );
  XOR U966 ( .A(n933), .B(n930), .Z(n932) );
  AND U967 ( .A(b[0]), .B(a[49]), .Z(n933) );
  XOR U968 ( .A(n934), .B(n935), .Z(n931) );
  XOR U969 ( .A(n936), .B(n937), .Z(n935) );
  AND U970 ( .A(b[2]), .B(a[47]), .Z(n937) );
  AND U971 ( .A(a[46]), .B(b[3]), .Z(n936) );
  AND U972 ( .A(b[1]), .B(a[48]), .Z(n934) );
  XOR U973 ( .A(sreg[177]), .B(n930), .Z(n114) );
  XOR U974 ( .A(n938), .B(n939), .Z(n930) );
  NOR U975 ( .A(n116), .B(n115), .Z(n938) );
  XOR U976 ( .A(n940), .B(n941), .Z(n115) );
  XOR U977 ( .A(n942), .B(n939), .Z(n941) );
  AND U978 ( .A(b[0]), .B(a[48]), .Z(n942) );
  XOR U979 ( .A(n943), .B(n944), .Z(n940) );
  XOR U980 ( .A(n945), .B(n946), .Z(n944) );
  AND U981 ( .A(a[45]), .B(b[3]), .Z(n946) );
  AND U982 ( .A(b[2]), .B(a[46]), .Z(n945) );
  AND U983 ( .A(b[1]), .B(a[47]), .Z(n943) );
  XOR U984 ( .A(sreg[176]), .B(n939), .Z(n116) );
  XOR U985 ( .A(n947), .B(n948), .Z(n939) );
  NOR U986 ( .A(n118), .B(n117), .Z(n947) );
  XOR U987 ( .A(n949), .B(n950), .Z(n117) );
  XOR U988 ( .A(n951), .B(n948), .Z(n950) );
  AND U989 ( .A(b[0]), .B(a[47]), .Z(n951) );
  XOR U990 ( .A(n952), .B(n953), .Z(n949) );
  XOR U991 ( .A(n954), .B(n955), .Z(n953) );
  AND U992 ( .A(a[44]), .B(b[3]), .Z(n955) );
  AND U993 ( .A(b[1]), .B(a[46]), .Z(n954) );
  AND U994 ( .A(b[2]), .B(a[45]), .Z(n952) );
  XOR U995 ( .A(sreg[175]), .B(n948), .Z(n118) );
  XOR U996 ( .A(n956), .B(n957), .Z(n948) );
  NOR U997 ( .A(n120), .B(n119), .Z(n956) );
  XOR U998 ( .A(n958), .B(n959), .Z(n119) );
  XOR U999 ( .A(n960), .B(n957), .Z(n959) );
  AND U1000 ( .A(b[0]), .B(a[46]), .Z(n960) );
  XOR U1001 ( .A(n961), .B(n962), .Z(n958) );
  XOR U1002 ( .A(n963), .B(n964), .Z(n962) );
  AND U1003 ( .A(b[2]), .B(a[44]), .Z(n964) );
  AND U1004 ( .A(a[43]), .B(b[3]), .Z(n963) );
  AND U1005 ( .A(b[1]), .B(a[45]), .Z(n961) );
  XOR U1006 ( .A(sreg[174]), .B(n957), .Z(n120) );
  XOR U1007 ( .A(n965), .B(n966), .Z(n957) );
  NOR U1008 ( .A(n122), .B(n121), .Z(n965) );
  XOR U1009 ( .A(n967), .B(n968), .Z(n121) );
  XOR U1010 ( .A(n969), .B(n966), .Z(n968) );
  AND U1011 ( .A(b[0]), .B(a[45]), .Z(n969) );
  XOR U1012 ( .A(n970), .B(n971), .Z(n967) );
  XOR U1013 ( .A(n972), .B(n973), .Z(n971) );
  AND U1014 ( .A(a[42]), .B(b[3]), .Z(n973) );
  AND U1015 ( .A(b[2]), .B(a[43]), .Z(n972) );
  AND U1016 ( .A(b[1]), .B(a[44]), .Z(n970) );
  XOR U1017 ( .A(sreg[173]), .B(n966), .Z(n122) );
  XOR U1018 ( .A(n974), .B(n975), .Z(n966) );
  NOR U1019 ( .A(n124), .B(n123), .Z(n974) );
  XOR U1020 ( .A(n976), .B(n977), .Z(n123) );
  XOR U1021 ( .A(n978), .B(n975), .Z(n977) );
  AND U1022 ( .A(b[0]), .B(a[44]), .Z(n978) );
  XOR U1023 ( .A(n979), .B(n980), .Z(n976) );
  XOR U1024 ( .A(n981), .B(n982), .Z(n980) );
  AND U1025 ( .A(a[41]), .B(b[3]), .Z(n982) );
  AND U1026 ( .A(b[1]), .B(a[43]), .Z(n981) );
  AND U1027 ( .A(b[2]), .B(a[42]), .Z(n979) );
  XOR U1028 ( .A(sreg[172]), .B(n975), .Z(n124) );
  XOR U1029 ( .A(n983), .B(n984), .Z(n975) );
  NOR U1030 ( .A(n126), .B(n125), .Z(n983) );
  XOR U1031 ( .A(n985), .B(n986), .Z(n125) );
  XOR U1032 ( .A(n987), .B(n984), .Z(n986) );
  AND U1033 ( .A(b[0]), .B(a[43]), .Z(n987) );
  XOR U1034 ( .A(n988), .B(n989), .Z(n985) );
  XOR U1035 ( .A(n990), .B(n991), .Z(n989) );
  AND U1036 ( .A(b[2]), .B(a[41]), .Z(n991) );
  AND U1037 ( .A(a[40]), .B(b[3]), .Z(n990) );
  AND U1038 ( .A(b[1]), .B(a[42]), .Z(n988) );
  XOR U1039 ( .A(sreg[171]), .B(n984), .Z(n126) );
  XOR U1040 ( .A(n992), .B(n993), .Z(n984) );
  NOR U1041 ( .A(n128), .B(n127), .Z(n992) );
  XOR U1042 ( .A(n994), .B(n995), .Z(n127) );
  XOR U1043 ( .A(n996), .B(n993), .Z(n995) );
  AND U1044 ( .A(b[0]), .B(a[42]), .Z(n996) );
  XOR U1045 ( .A(n997), .B(n998), .Z(n994) );
  XOR U1046 ( .A(n999), .B(n1000), .Z(n998) );
  AND U1047 ( .A(a[39]), .B(b[3]), .Z(n1000) );
  AND U1048 ( .A(b[2]), .B(a[40]), .Z(n999) );
  AND U1049 ( .A(b[1]), .B(a[41]), .Z(n997) );
  XOR U1050 ( .A(sreg[170]), .B(n993), .Z(n128) );
  XOR U1051 ( .A(n1001), .B(n1002), .Z(n993) );
  NOR U1052 ( .A(n130), .B(n129), .Z(n1001) );
  XOR U1053 ( .A(n1003), .B(n1004), .Z(n129) );
  XOR U1054 ( .A(n1005), .B(n1002), .Z(n1004) );
  AND U1055 ( .A(b[0]), .B(a[41]), .Z(n1005) );
  XOR U1056 ( .A(n1006), .B(n1007), .Z(n1003) );
  XOR U1057 ( .A(n1008), .B(n1009), .Z(n1007) );
  AND U1058 ( .A(a[38]), .B(b[3]), .Z(n1009) );
  AND U1059 ( .A(b[1]), .B(a[40]), .Z(n1008) );
  AND U1060 ( .A(b[2]), .B(a[39]), .Z(n1006) );
  XOR U1061 ( .A(sreg[169]), .B(n1002), .Z(n130) );
  XOR U1062 ( .A(n1010), .B(n1011), .Z(n1002) );
  NOR U1063 ( .A(n132), .B(n131), .Z(n1010) );
  XOR U1064 ( .A(n1012), .B(n1013), .Z(n131) );
  XOR U1065 ( .A(n1014), .B(n1011), .Z(n1013) );
  AND U1066 ( .A(b[0]), .B(a[40]), .Z(n1014) );
  XOR U1067 ( .A(n1015), .B(n1016), .Z(n1012) );
  XOR U1068 ( .A(n1017), .B(n1018), .Z(n1016) );
  AND U1069 ( .A(b[2]), .B(a[38]), .Z(n1018) );
  AND U1070 ( .A(a[37]), .B(b[3]), .Z(n1017) );
  AND U1071 ( .A(b[1]), .B(a[39]), .Z(n1015) );
  XOR U1072 ( .A(sreg[168]), .B(n1011), .Z(n132) );
  XOR U1073 ( .A(n1019), .B(n1020), .Z(n1011) );
  NOR U1074 ( .A(n134), .B(n133), .Z(n1019) );
  XOR U1075 ( .A(n1021), .B(n1022), .Z(n133) );
  XOR U1076 ( .A(n1023), .B(n1020), .Z(n1022) );
  AND U1077 ( .A(b[0]), .B(a[39]), .Z(n1023) );
  XOR U1078 ( .A(n1024), .B(n1025), .Z(n1021) );
  XOR U1079 ( .A(n1026), .B(n1027), .Z(n1025) );
  AND U1080 ( .A(a[36]), .B(b[3]), .Z(n1027) );
  AND U1081 ( .A(b[2]), .B(a[37]), .Z(n1026) );
  AND U1082 ( .A(b[1]), .B(a[38]), .Z(n1024) );
  XOR U1083 ( .A(sreg[167]), .B(n1020), .Z(n134) );
  XOR U1084 ( .A(n1028), .B(n1029), .Z(n1020) );
  NOR U1085 ( .A(n136), .B(n135), .Z(n1028) );
  XOR U1086 ( .A(n1030), .B(n1031), .Z(n135) );
  XOR U1087 ( .A(n1032), .B(n1029), .Z(n1031) );
  AND U1088 ( .A(b[0]), .B(a[38]), .Z(n1032) );
  XOR U1089 ( .A(n1033), .B(n1034), .Z(n1030) );
  XOR U1090 ( .A(n1035), .B(n1036), .Z(n1034) );
  AND U1091 ( .A(a[35]), .B(b[3]), .Z(n1036) );
  AND U1092 ( .A(b[1]), .B(a[37]), .Z(n1035) );
  AND U1093 ( .A(b[2]), .B(a[36]), .Z(n1033) );
  XOR U1094 ( .A(sreg[166]), .B(n1029), .Z(n136) );
  XOR U1095 ( .A(n1037), .B(n1038), .Z(n1029) );
  NOR U1096 ( .A(n138), .B(n137), .Z(n1037) );
  XOR U1097 ( .A(n1039), .B(n1040), .Z(n137) );
  XOR U1098 ( .A(n1041), .B(n1038), .Z(n1040) );
  AND U1099 ( .A(b[0]), .B(a[37]), .Z(n1041) );
  XOR U1100 ( .A(n1042), .B(n1043), .Z(n1039) );
  XOR U1101 ( .A(n1044), .B(n1045), .Z(n1043) );
  AND U1102 ( .A(b[2]), .B(a[35]), .Z(n1045) );
  AND U1103 ( .A(a[34]), .B(b[3]), .Z(n1044) );
  AND U1104 ( .A(b[1]), .B(a[36]), .Z(n1042) );
  XOR U1105 ( .A(sreg[165]), .B(n1038), .Z(n138) );
  XOR U1106 ( .A(n1046), .B(n1047), .Z(n1038) );
  NOR U1107 ( .A(n140), .B(n139), .Z(n1046) );
  XOR U1108 ( .A(n1048), .B(n1049), .Z(n139) );
  XOR U1109 ( .A(n1050), .B(n1047), .Z(n1049) );
  AND U1110 ( .A(b[0]), .B(a[36]), .Z(n1050) );
  XOR U1111 ( .A(n1051), .B(n1052), .Z(n1048) );
  XOR U1112 ( .A(n1053), .B(n1054), .Z(n1052) );
  AND U1113 ( .A(a[33]), .B(b[3]), .Z(n1054) );
  AND U1114 ( .A(b[2]), .B(a[34]), .Z(n1053) );
  AND U1115 ( .A(b[1]), .B(a[35]), .Z(n1051) );
  XOR U1116 ( .A(sreg[164]), .B(n1047), .Z(n140) );
  XOR U1117 ( .A(n1055), .B(n1056), .Z(n1047) );
  NOR U1118 ( .A(n142), .B(n141), .Z(n1055) );
  XOR U1119 ( .A(n1057), .B(n1058), .Z(n141) );
  XOR U1120 ( .A(n1059), .B(n1056), .Z(n1058) );
  AND U1121 ( .A(b[0]), .B(a[35]), .Z(n1059) );
  XOR U1122 ( .A(n1060), .B(n1061), .Z(n1057) );
  XOR U1123 ( .A(n1062), .B(n1063), .Z(n1061) );
  AND U1124 ( .A(a[32]), .B(b[3]), .Z(n1063) );
  AND U1125 ( .A(b[1]), .B(a[34]), .Z(n1062) );
  AND U1126 ( .A(b[2]), .B(a[33]), .Z(n1060) );
  XOR U1127 ( .A(sreg[163]), .B(n1056), .Z(n142) );
  XOR U1128 ( .A(n1064), .B(n1065), .Z(n1056) );
  NOR U1129 ( .A(n144), .B(n143), .Z(n1064) );
  XOR U1130 ( .A(n1066), .B(n1067), .Z(n143) );
  XOR U1131 ( .A(n1068), .B(n1065), .Z(n1067) );
  AND U1132 ( .A(b[0]), .B(a[34]), .Z(n1068) );
  XOR U1133 ( .A(n1069), .B(n1070), .Z(n1066) );
  XOR U1134 ( .A(n1071), .B(n1072), .Z(n1070) );
  AND U1135 ( .A(b[2]), .B(a[32]), .Z(n1072) );
  AND U1136 ( .A(a[31]), .B(b[3]), .Z(n1071) );
  AND U1137 ( .A(b[1]), .B(a[33]), .Z(n1069) );
  XOR U1138 ( .A(sreg[162]), .B(n1065), .Z(n144) );
  XOR U1139 ( .A(n1073), .B(n1074), .Z(n1065) );
  NOR U1140 ( .A(n146), .B(n145), .Z(n1073) );
  XOR U1141 ( .A(n1075), .B(n1076), .Z(n145) );
  XOR U1142 ( .A(n1077), .B(n1074), .Z(n1076) );
  AND U1143 ( .A(b[0]), .B(a[33]), .Z(n1077) );
  XOR U1144 ( .A(n1078), .B(n1079), .Z(n1075) );
  XOR U1145 ( .A(n1080), .B(n1081), .Z(n1079) );
  AND U1146 ( .A(a[30]), .B(b[3]), .Z(n1081) );
  AND U1147 ( .A(b[2]), .B(a[31]), .Z(n1080) );
  AND U1148 ( .A(b[1]), .B(a[32]), .Z(n1078) );
  XOR U1149 ( .A(sreg[161]), .B(n1074), .Z(n146) );
  XOR U1150 ( .A(n1082), .B(n1083), .Z(n1074) );
  NOR U1151 ( .A(n148), .B(n147), .Z(n1082) );
  XOR U1152 ( .A(n1084), .B(n1085), .Z(n147) );
  XOR U1153 ( .A(n1086), .B(n1083), .Z(n1085) );
  AND U1154 ( .A(b[0]), .B(a[32]), .Z(n1086) );
  XOR U1155 ( .A(n1087), .B(n1088), .Z(n1084) );
  XOR U1156 ( .A(n1089), .B(n1090), .Z(n1088) );
  AND U1157 ( .A(a[29]), .B(b[3]), .Z(n1090) );
  AND U1158 ( .A(b[1]), .B(a[31]), .Z(n1089) );
  AND U1159 ( .A(b[2]), .B(a[30]), .Z(n1087) );
  XOR U1160 ( .A(sreg[160]), .B(n1083), .Z(n148) );
  XOR U1161 ( .A(n1091), .B(n1092), .Z(n1083) );
  NOR U1162 ( .A(n150), .B(n149), .Z(n1091) );
  XOR U1163 ( .A(n1093), .B(n1094), .Z(n149) );
  XOR U1164 ( .A(n1095), .B(n1092), .Z(n1094) );
  AND U1165 ( .A(b[0]), .B(a[31]), .Z(n1095) );
  XOR U1166 ( .A(n1096), .B(n1097), .Z(n1093) );
  XOR U1167 ( .A(n1098), .B(n1099), .Z(n1097) );
  AND U1168 ( .A(b[2]), .B(a[29]), .Z(n1099) );
  AND U1169 ( .A(a[28]), .B(b[3]), .Z(n1098) );
  AND U1170 ( .A(b[1]), .B(a[30]), .Z(n1096) );
  XOR U1171 ( .A(sreg[159]), .B(n1092), .Z(n150) );
  XOR U1172 ( .A(n1100), .B(n1101), .Z(n1092) );
  NOR U1173 ( .A(n152), .B(n151), .Z(n1100) );
  XOR U1174 ( .A(n1102), .B(n1103), .Z(n151) );
  XOR U1175 ( .A(n1104), .B(n1101), .Z(n1103) );
  AND U1176 ( .A(b[0]), .B(a[30]), .Z(n1104) );
  XOR U1177 ( .A(n1105), .B(n1106), .Z(n1102) );
  XOR U1178 ( .A(n1107), .B(n1108), .Z(n1106) );
  AND U1179 ( .A(a[27]), .B(b[3]), .Z(n1108) );
  AND U1180 ( .A(b[2]), .B(a[28]), .Z(n1107) );
  AND U1181 ( .A(b[1]), .B(a[29]), .Z(n1105) );
  XOR U1182 ( .A(sreg[158]), .B(n1101), .Z(n152) );
  XOR U1183 ( .A(n1109), .B(n1110), .Z(n1101) );
  NOR U1184 ( .A(n154), .B(n153), .Z(n1109) );
  XOR U1185 ( .A(n1111), .B(n1112), .Z(n153) );
  XOR U1186 ( .A(n1113), .B(n1110), .Z(n1112) );
  AND U1187 ( .A(b[0]), .B(a[29]), .Z(n1113) );
  XOR U1188 ( .A(n1114), .B(n1115), .Z(n1111) );
  XOR U1189 ( .A(n1116), .B(n1117), .Z(n1115) );
  AND U1190 ( .A(a[26]), .B(b[3]), .Z(n1117) );
  AND U1191 ( .A(b[1]), .B(a[28]), .Z(n1116) );
  AND U1192 ( .A(b[2]), .B(a[27]), .Z(n1114) );
  XOR U1193 ( .A(sreg[157]), .B(n1110), .Z(n154) );
  XOR U1194 ( .A(n1118), .B(n1119), .Z(n1110) );
  NOR U1195 ( .A(n156), .B(n155), .Z(n1118) );
  XOR U1196 ( .A(n1120), .B(n1121), .Z(n155) );
  XOR U1197 ( .A(n1122), .B(n1119), .Z(n1121) );
  AND U1198 ( .A(b[0]), .B(a[28]), .Z(n1122) );
  XOR U1199 ( .A(n1123), .B(n1124), .Z(n1120) );
  XOR U1200 ( .A(n1125), .B(n1126), .Z(n1124) );
  AND U1201 ( .A(b[2]), .B(a[26]), .Z(n1126) );
  AND U1202 ( .A(a[25]), .B(b[3]), .Z(n1125) );
  AND U1203 ( .A(b[1]), .B(a[27]), .Z(n1123) );
  XOR U1204 ( .A(sreg[156]), .B(n1119), .Z(n156) );
  XOR U1205 ( .A(n1127), .B(n1128), .Z(n1119) );
  NOR U1206 ( .A(n158), .B(n157), .Z(n1127) );
  XOR U1207 ( .A(n1129), .B(n1130), .Z(n157) );
  XOR U1208 ( .A(n1131), .B(n1128), .Z(n1130) );
  AND U1209 ( .A(b[0]), .B(a[27]), .Z(n1131) );
  XOR U1210 ( .A(n1132), .B(n1133), .Z(n1129) );
  XOR U1211 ( .A(n1134), .B(n1135), .Z(n1133) );
  AND U1212 ( .A(a[24]), .B(b[3]), .Z(n1135) );
  AND U1213 ( .A(b[2]), .B(a[25]), .Z(n1134) );
  AND U1214 ( .A(b[1]), .B(a[26]), .Z(n1132) );
  XOR U1215 ( .A(sreg[155]), .B(n1128), .Z(n158) );
  XOR U1216 ( .A(n1136), .B(n1137), .Z(n1128) );
  NOR U1217 ( .A(n160), .B(n159), .Z(n1136) );
  XOR U1218 ( .A(n1138), .B(n1139), .Z(n159) );
  XOR U1219 ( .A(n1140), .B(n1137), .Z(n1139) );
  AND U1220 ( .A(b[0]), .B(a[26]), .Z(n1140) );
  XOR U1221 ( .A(n1141), .B(n1142), .Z(n1138) );
  XOR U1222 ( .A(n1143), .B(n1144), .Z(n1142) );
  AND U1223 ( .A(a[23]), .B(b[3]), .Z(n1144) );
  AND U1224 ( .A(b[1]), .B(a[25]), .Z(n1143) );
  AND U1225 ( .A(b[2]), .B(a[24]), .Z(n1141) );
  XOR U1226 ( .A(sreg[154]), .B(n1137), .Z(n160) );
  XOR U1227 ( .A(n1145), .B(n1146), .Z(n1137) );
  NOR U1228 ( .A(n162), .B(n161), .Z(n1145) );
  XOR U1229 ( .A(n1147), .B(n1148), .Z(n161) );
  XOR U1230 ( .A(n1149), .B(n1146), .Z(n1148) );
  AND U1231 ( .A(b[0]), .B(a[25]), .Z(n1149) );
  XOR U1232 ( .A(n1150), .B(n1151), .Z(n1147) );
  XOR U1233 ( .A(n1152), .B(n1153), .Z(n1151) );
  AND U1234 ( .A(b[2]), .B(a[23]), .Z(n1153) );
  AND U1235 ( .A(a[22]), .B(b[3]), .Z(n1152) );
  AND U1236 ( .A(b[1]), .B(a[24]), .Z(n1150) );
  XOR U1237 ( .A(sreg[153]), .B(n1146), .Z(n162) );
  XOR U1238 ( .A(n1154), .B(n1155), .Z(n1146) );
  NOR U1239 ( .A(n164), .B(n163), .Z(n1154) );
  XOR U1240 ( .A(n1156), .B(n1157), .Z(n163) );
  XOR U1241 ( .A(n1158), .B(n1155), .Z(n1157) );
  AND U1242 ( .A(b[0]), .B(a[24]), .Z(n1158) );
  XOR U1243 ( .A(n1159), .B(n1160), .Z(n1156) );
  XOR U1244 ( .A(n1161), .B(n1162), .Z(n1160) );
  AND U1245 ( .A(a[21]), .B(b[3]), .Z(n1162) );
  AND U1246 ( .A(b[2]), .B(a[22]), .Z(n1161) );
  AND U1247 ( .A(b[1]), .B(a[23]), .Z(n1159) );
  XOR U1248 ( .A(sreg[152]), .B(n1155), .Z(n164) );
  XOR U1249 ( .A(n1163), .B(n1164), .Z(n1155) );
  NOR U1250 ( .A(n166), .B(n165), .Z(n1163) );
  XOR U1251 ( .A(n1165), .B(n1166), .Z(n165) );
  XOR U1252 ( .A(n1167), .B(n1164), .Z(n1166) );
  AND U1253 ( .A(b[0]), .B(a[23]), .Z(n1167) );
  XOR U1254 ( .A(n1168), .B(n1169), .Z(n1165) );
  XOR U1255 ( .A(n1170), .B(n1171), .Z(n1169) );
  AND U1256 ( .A(a[20]), .B(b[3]), .Z(n1171) );
  AND U1257 ( .A(b[1]), .B(a[22]), .Z(n1170) );
  AND U1258 ( .A(b[2]), .B(a[21]), .Z(n1168) );
  XOR U1259 ( .A(sreg[151]), .B(n1164), .Z(n166) );
  XOR U1260 ( .A(n1172), .B(n1173), .Z(n1164) );
  NOR U1261 ( .A(n168), .B(n167), .Z(n1172) );
  XOR U1262 ( .A(n1174), .B(n1175), .Z(n167) );
  XOR U1263 ( .A(n1176), .B(n1173), .Z(n1175) );
  AND U1264 ( .A(b[0]), .B(a[22]), .Z(n1176) );
  XOR U1265 ( .A(n1177), .B(n1178), .Z(n1174) );
  XOR U1266 ( .A(n1179), .B(n1180), .Z(n1178) );
  AND U1267 ( .A(b[2]), .B(a[20]), .Z(n1180) );
  AND U1268 ( .A(a[19]), .B(b[3]), .Z(n1179) );
  AND U1269 ( .A(b[1]), .B(a[21]), .Z(n1177) );
  XOR U1270 ( .A(sreg[150]), .B(n1173), .Z(n168) );
  XOR U1271 ( .A(n1181), .B(n1182), .Z(n1173) );
  NOR U1272 ( .A(n170), .B(n169), .Z(n1181) );
  XOR U1273 ( .A(n1183), .B(n1184), .Z(n169) );
  XOR U1274 ( .A(n1185), .B(n1182), .Z(n1184) );
  AND U1275 ( .A(b[0]), .B(a[21]), .Z(n1185) );
  XOR U1276 ( .A(n1186), .B(n1187), .Z(n1183) );
  XOR U1277 ( .A(n1188), .B(n1189), .Z(n1187) );
  AND U1278 ( .A(a[18]), .B(b[3]), .Z(n1189) );
  AND U1279 ( .A(b[2]), .B(a[19]), .Z(n1188) );
  AND U1280 ( .A(b[1]), .B(a[20]), .Z(n1186) );
  XOR U1281 ( .A(sreg[149]), .B(n1182), .Z(n170) );
  XOR U1282 ( .A(n1190), .B(n1191), .Z(n1182) );
  NOR U1283 ( .A(n172), .B(n171), .Z(n1190) );
  XOR U1284 ( .A(n1192), .B(n1193), .Z(n171) );
  XOR U1285 ( .A(n1194), .B(n1191), .Z(n1193) );
  AND U1286 ( .A(b[0]), .B(a[20]), .Z(n1194) );
  XOR U1287 ( .A(n1195), .B(n1196), .Z(n1192) );
  XOR U1288 ( .A(n1197), .B(n1198), .Z(n1196) );
  AND U1289 ( .A(a[17]), .B(b[3]), .Z(n1198) );
  AND U1290 ( .A(b[1]), .B(a[19]), .Z(n1197) );
  AND U1291 ( .A(b[2]), .B(a[18]), .Z(n1195) );
  XOR U1292 ( .A(sreg[148]), .B(n1191), .Z(n172) );
  XOR U1293 ( .A(n1199), .B(n1200), .Z(n1191) );
  NOR U1294 ( .A(n174), .B(n173), .Z(n1199) );
  XOR U1295 ( .A(n1201), .B(n1202), .Z(n173) );
  XOR U1296 ( .A(n1203), .B(n1200), .Z(n1202) );
  AND U1297 ( .A(b[0]), .B(a[19]), .Z(n1203) );
  XOR U1298 ( .A(n1204), .B(n1205), .Z(n1201) );
  XOR U1299 ( .A(n1206), .B(n1207), .Z(n1205) );
  AND U1300 ( .A(b[2]), .B(a[17]), .Z(n1207) );
  AND U1301 ( .A(a[16]), .B(b[3]), .Z(n1206) );
  AND U1302 ( .A(b[1]), .B(a[18]), .Z(n1204) );
  XOR U1303 ( .A(sreg[147]), .B(n1200), .Z(n174) );
  XOR U1304 ( .A(n1208), .B(n1209), .Z(n1200) );
  NOR U1305 ( .A(n176), .B(n175), .Z(n1208) );
  XOR U1306 ( .A(n1210), .B(n1211), .Z(n175) );
  XOR U1307 ( .A(n1212), .B(n1209), .Z(n1211) );
  AND U1308 ( .A(b[0]), .B(a[18]), .Z(n1212) );
  XOR U1309 ( .A(n1213), .B(n1214), .Z(n1210) );
  XOR U1310 ( .A(n1215), .B(n1216), .Z(n1214) );
  AND U1311 ( .A(a[15]), .B(b[3]), .Z(n1216) );
  AND U1312 ( .A(b[2]), .B(a[16]), .Z(n1215) );
  AND U1313 ( .A(b[1]), .B(a[17]), .Z(n1213) );
  XOR U1314 ( .A(sreg[146]), .B(n1209), .Z(n176) );
  XOR U1315 ( .A(n1217), .B(n1218), .Z(n1209) );
  NOR U1316 ( .A(n178), .B(n177), .Z(n1217) );
  XOR U1317 ( .A(n1219), .B(n1220), .Z(n177) );
  XOR U1318 ( .A(n1221), .B(n1218), .Z(n1220) );
  AND U1319 ( .A(b[0]), .B(a[17]), .Z(n1221) );
  XOR U1320 ( .A(n1222), .B(n1223), .Z(n1219) );
  XOR U1321 ( .A(n1224), .B(n1225), .Z(n1223) );
  AND U1322 ( .A(a[14]), .B(b[3]), .Z(n1225) );
  AND U1323 ( .A(b[1]), .B(a[16]), .Z(n1224) );
  AND U1324 ( .A(b[2]), .B(a[15]), .Z(n1222) );
  XOR U1325 ( .A(sreg[145]), .B(n1218), .Z(n178) );
  XOR U1326 ( .A(n1226), .B(n1227), .Z(n1218) );
  NOR U1327 ( .A(n180), .B(n179), .Z(n1226) );
  XOR U1328 ( .A(n1228), .B(n1229), .Z(n179) );
  XOR U1329 ( .A(n1230), .B(n1227), .Z(n1229) );
  AND U1330 ( .A(b[0]), .B(a[16]), .Z(n1230) );
  XOR U1331 ( .A(n1231), .B(n1232), .Z(n1228) );
  XOR U1332 ( .A(n1233), .B(n1234), .Z(n1232) );
  AND U1333 ( .A(b[2]), .B(a[14]), .Z(n1234) );
  AND U1334 ( .A(a[13]), .B(b[3]), .Z(n1233) );
  AND U1335 ( .A(b[1]), .B(a[15]), .Z(n1231) );
  XOR U1336 ( .A(sreg[144]), .B(n1227), .Z(n180) );
  XOR U1337 ( .A(n1235), .B(n1236), .Z(n1227) );
  NOR U1338 ( .A(n182), .B(n181), .Z(n1235) );
  XOR U1339 ( .A(n1237), .B(n1238), .Z(n181) );
  XOR U1340 ( .A(n1239), .B(n1236), .Z(n1238) );
  AND U1341 ( .A(b[0]), .B(a[15]), .Z(n1239) );
  XOR U1342 ( .A(n1240), .B(n1241), .Z(n1237) );
  XOR U1343 ( .A(n1242), .B(n1243), .Z(n1241) );
  AND U1344 ( .A(a[12]), .B(b[3]), .Z(n1243) );
  AND U1345 ( .A(b[2]), .B(a[13]), .Z(n1242) );
  AND U1346 ( .A(b[1]), .B(a[14]), .Z(n1240) );
  XOR U1347 ( .A(sreg[143]), .B(n1236), .Z(n182) );
  XOR U1348 ( .A(n1244), .B(n1245), .Z(n1236) );
  NOR U1349 ( .A(n184), .B(n183), .Z(n1244) );
  XOR U1350 ( .A(n1246), .B(n1247), .Z(n183) );
  XOR U1351 ( .A(n1248), .B(n1245), .Z(n1247) );
  AND U1352 ( .A(b[0]), .B(a[14]), .Z(n1248) );
  XOR U1353 ( .A(n1249), .B(n1250), .Z(n1246) );
  XOR U1354 ( .A(n1251), .B(n1252), .Z(n1250) );
  AND U1355 ( .A(a[11]), .B(b[3]), .Z(n1252) );
  AND U1356 ( .A(b[1]), .B(a[13]), .Z(n1251) );
  AND U1357 ( .A(b[2]), .B(a[12]), .Z(n1249) );
  XOR U1358 ( .A(sreg[142]), .B(n1245), .Z(n184) );
  XOR U1359 ( .A(n1253), .B(n1254), .Z(n1245) );
  NOR U1360 ( .A(n186), .B(n185), .Z(n1253) );
  XOR U1361 ( .A(n1255), .B(n1256), .Z(n185) );
  XOR U1362 ( .A(n1257), .B(n1254), .Z(n1256) );
  AND U1363 ( .A(b[0]), .B(a[13]), .Z(n1257) );
  XOR U1364 ( .A(n1258), .B(n1259), .Z(n1255) );
  XOR U1365 ( .A(n1260), .B(n1261), .Z(n1259) );
  AND U1366 ( .A(b[2]), .B(a[11]), .Z(n1261) );
  AND U1367 ( .A(a[10]), .B(b[3]), .Z(n1260) );
  AND U1368 ( .A(b[1]), .B(a[12]), .Z(n1258) );
  XOR U1369 ( .A(sreg[141]), .B(n1254), .Z(n186) );
  XOR U1370 ( .A(n1262), .B(n1263), .Z(n1254) );
  NOR U1371 ( .A(n188), .B(n187), .Z(n1262) );
  XOR U1372 ( .A(n1264), .B(n1265), .Z(n187) );
  XOR U1373 ( .A(n1266), .B(n1263), .Z(n1265) );
  AND U1374 ( .A(b[0]), .B(a[12]), .Z(n1266) );
  XOR U1375 ( .A(n1267), .B(n1268), .Z(n1264) );
  XOR U1376 ( .A(n1269), .B(n1270), .Z(n1268) );
  AND U1377 ( .A(a[9]), .B(b[3]), .Z(n1270) );
  AND U1378 ( .A(b[2]), .B(a[10]), .Z(n1269) );
  AND U1379 ( .A(b[1]), .B(a[11]), .Z(n1267) );
  XOR U1380 ( .A(sreg[140]), .B(n1263), .Z(n188) );
  XOR U1381 ( .A(n1271), .B(n1272), .Z(n1263) );
  NOR U1382 ( .A(n268), .B(n267), .Z(n1271) );
  XOR U1383 ( .A(n1273), .B(n1274), .Z(n267) );
  XOR U1384 ( .A(n1275), .B(n1272), .Z(n1274) );
  AND U1385 ( .A(b[0]), .B(a[11]), .Z(n1275) );
  XOR U1386 ( .A(n1276), .B(n1277), .Z(n1273) );
  XOR U1387 ( .A(n1278), .B(n1279), .Z(n1277) );
  AND U1388 ( .A(a[8]), .B(b[3]), .Z(n1279) );
  AND U1389 ( .A(b[1]), .B(a[10]), .Z(n1278) );
  AND U1390 ( .A(b[2]), .B(a[9]), .Z(n1276) );
  XOR U1391 ( .A(sreg[139]), .B(n1272), .Z(n268) );
  XOR U1392 ( .A(n1280), .B(n1281), .Z(n1272) );
  NOR U1393 ( .A(n380), .B(n379), .Z(n1280) );
  XOR U1394 ( .A(n1282), .B(n1283), .Z(n379) );
  XOR U1395 ( .A(n1284), .B(n1281), .Z(n1283) );
  AND U1396 ( .A(b[0]), .B(a[10]), .Z(n1284) );
  XOR U1397 ( .A(n1285), .B(n1286), .Z(n1282) );
  XOR U1398 ( .A(n1287), .B(n1288), .Z(n1286) );
  AND U1399 ( .A(b[2]), .B(a[8]), .Z(n1288) );
  AND U1400 ( .A(a[7]), .B(b[3]), .Z(n1287) );
  AND U1401 ( .A(b[1]), .B(a[9]), .Z(n1285) );
  XOR U1402 ( .A(sreg[138]), .B(n1281), .Z(n380) );
  XOR U1403 ( .A(n1289), .B(n1290), .Z(n1281) );
  NOR U1404 ( .A(n2), .B(n1), .Z(n1289) );
  XOR U1405 ( .A(sreg[137]), .B(n1290), .Z(n1) );
  XOR U1406 ( .A(n1291), .B(n1292), .Z(n2) );
  XOR U1407 ( .A(n1293), .B(n1290), .Z(n1292) );
  XOR U1408 ( .A(n1294), .B(n1295), .Z(n1290) );
  NOR U1409 ( .A(n24), .B(n23), .Z(n1294) );
  XOR U1410 ( .A(n1296), .B(n1297), .Z(n23) );
  XOR U1411 ( .A(n1298), .B(n1295), .Z(n1297) );
  AND U1412 ( .A(b[0]), .B(a[8]), .Z(n1298) );
  XOR U1413 ( .A(n1299), .B(n1300), .Z(n1296) );
  XOR U1414 ( .A(n1301), .B(n1302), .Z(n1300) );
  AND U1415 ( .A(a[5]), .B(b[3]), .Z(n1302) );
  AND U1416 ( .A(a[7]), .B(b[1]), .Z(n1301) );
  AND U1417 ( .A(b[2]), .B(a[6]), .Z(n1299) );
  XOR U1418 ( .A(sreg[136]), .B(n1295), .Z(n24) );
  XOR U1419 ( .A(n1303), .B(n1304), .Z(n1295) );
  NOR U1420 ( .A(n46), .B(n45), .Z(n1303) );
  XOR U1421 ( .A(n1305), .B(n1306), .Z(n45) );
  XOR U1422 ( .A(n1307), .B(n1304), .Z(n1306) );
  AND U1423 ( .A(a[7]), .B(b[0]), .Z(n1307) );
  XOR U1424 ( .A(n1308), .B(n1309), .Z(n1305) );
  XOR U1425 ( .A(n1310), .B(n1311), .Z(n1309) );
  AND U1426 ( .A(a[5]), .B(b[2]), .Z(n1311) );
  AND U1427 ( .A(a[4]), .B(b[3]), .Z(n1310) );
  AND U1428 ( .A(b[1]), .B(a[6]), .Z(n1308) );
  XOR U1429 ( .A(sreg[135]), .B(n1304), .Z(n46) );
  XOR U1430 ( .A(n1312), .B(n1313), .Z(n1304) );
  NOR U1431 ( .A(n68), .B(n67), .Z(n1312) );
  XOR U1432 ( .A(n1314), .B(n1315), .Z(n67) );
  XOR U1433 ( .A(n1316), .B(n1313), .Z(n1315) );
  AND U1434 ( .A(b[0]), .B(a[6]), .Z(n1316) );
  XOR U1435 ( .A(n1317), .B(n1318), .Z(n1314) );
  XOR U1436 ( .A(n1319), .B(n1320), .Z(n1318) );
  AND U1437 ( .A(a[3]), .B(b[3]), .Z(n1320) );
  AND U1438 ( .A(b[2]), .B(a[4]), .Z(n1319) );
  AND U1439 ( .A(a[5]), .B(b[1]), .Z(n1317) );
  XOR U1440 ( .A(sreg[134]), .B(n1313), .Z(n68) );
  XOR U1441 ( .A(n1321), .B(n1322), .Z(n1313) );
  NOR U1442 ( .A(n90), .B(n89), .Z(n1321) );
  XOR U1443 ( .A(n1323), .B(n1324), .Z(n89) );
  XOR U1444 ( .A(n1325), .B(n1322), .Z(n1324) );
  AND U1445 ( .A(b[0]), .B(a[5]), .Z(n1325) );
  XOR U1446 ( .A(n1326), .B(n1327), .Z(n1323) );
  XOR U1447 ( .A(n1328), .B(n1329), .Z(n1327) );
  AND U1448 ( .A(a[2]), .B(b[3]), .Z(n1329) );
  AND U1449 ( .A(a[4]), .B(b[1]), .Z(n1328) );
  AND U1450 ( .A(b[2]), .B(a[3]), .Z(n1326) );
  XOR U1451 ( .A(sreg[133]), .B(n1322), .Z(n90) );
  XOR U1452 ( .A(n1330), .B(n1331), .Z(n1322) );
  NOR U1453 ( .A(n112), .B(n111), .Z(n1330) );
  XOR U1454 ( .A(n1332), .B(n1333), .Z(n111) );
  XOR U1455 ( .A(n1334), .B(n1331), .Z(n1333) );
  AND U1456 ( .A(b[0]), .B(a[4]), .Z(n1334) );
  XOR U1457 ( .A(n1335), .B(n1336), .Z(n1332) );
  XOR U1458 ( .A(n1337), .B(n1338), .Z(n1336) );
  AND U1459 ( .A(b[2]), .B(a[2]), .Z(n1338) );
  AND U1460 ( .A(a[1]), .B(b[3]), .Z(n1337) );
  AND U1461 ( .A(a[3]), .B(b[1]), .Z(n1335) );
  XOR U1462 ( .A(sreg[132]), .B(n1331), .Z(n112) );
  XOR U1463 ( .A(n1339), .B(n1340), .Z(n1331) );
  NOR U1464 ( .A(n1341), .B(n1342), .Z(n1339) );
  AND U1465 ( .A(b[0]), .B(a[9]), .Z(n1293) );
  XOR U1466 ( .A(n1343), .B(n1344), .Z(n1291) );
  XOR U1467 ( .A(n1345), .B(n1346), .Z(n1344) );
  AND U1468 ( .A(a[6]), .B(b[3]), .Z(n1346) );
  AND U1469 ( .A(a[7]), .B(b[2]), .Z(n1345) );
  AND U1470 ( .A(b[1]), .B(a[8]), .Z(n1343) );
  AND U1471 ( .A(b[0]), .B(a[99]), .Z(n487) );
  XOR U1472 ( .A(n1347), .B(n1348), .Z(n485) );
  XOR U1473 ( .A(n1349), .B(n1350), .Z(n1348) );
  AND U1474 ( .A(a[96]), .B(b[3]), .Z(n1350) );
  AND U1475 ( .A(b[2]), .B(a[97]), .Z(n1349) );
  AND U1476 ( .A(b[1]), .B(a[98]), .Z(n1347) );
  AND U1477 ( .A(b[0]), .B(a[100]), .Z(n482) );
  XOR U1478 ( .A(n1351), .B(n1352), .Z(n480) );
  XOR U1479 ( .A(n1353), .B(n1354), .Z(n1352) );
  AND U1480 ( .A(b[2]), .B(a[98]), .Z(n1354) );
  AND U1481 ( .A(a[97]), .B(b[3]), .Z(n1353) );
  AND U1482 ( .A(b[1]), .B(a[99]), .Z(n1351) );
  XOR U1483 ( .A(n1342), .B(n1341), .Z(c[127]) );
  XOR U1484 ( .A(sreg[131]), .B(n1340), .Z(n1341) );
  XOR U1485 ( .A(n1355), .B(n1356), .Z(n1342) );
  XOR U1486 ( .A(n1357), .B(n1340), .Z(n1356) );
  XOR U1487 ( .A(n1358), .B(n1359), .Z(n1340) );
  NOR U1488 ( .A(n1360), .B(n1361), .Z(n1358) );
  AND U1489 ( .A(b[0]), .B(a[3]), .Z(n1357) );
  XOR U1490 ( .A(n1362), .B(n1363), .Z(n1355) );
  XOR U1491 ( .A(n1364), .B(n1365), .Z(n1363) );
  AND U1492 ( .A(b[2]), .B(a[1]), .Z(n1365) );
  AND U1493 ( .A(a[0]), .B(b[3]), .Z(n1364) );
  AND U1494 ( .A(a[2]), .B(b[1]), .Z(n1362) );
  XOR U1495 ( .A(n1361), .B(n1360), .Z(c[126]) );
  XOR U1496 ( .A(sreg[130]), .B(n1359), .Z(n1360) );
  XOR U1497 ( .A(n1366), .B(n1367), .Z(n1361) );
  XOR U1498 ( .A(n1369), .B(n1370), .Z(n1359) );
  NAND U1499 ( .A(n1371), .B(n1372), .Z(n1370) );
  AND U1500 ( .A(b[0]), .B(a[2]), .Z(n1368) );
  XOR U1501 ( .A(n1373), .B(n1374), .Z(n1366) );
  AND U1502 ( .A(a[1]), .B(b[1]), .Z(n1374) );
  AND U1503 ( .A(b[2]), .B(a[0]), .Z(n1373) );
  XOR U1504 ( .A(n1371), .B(n1372), .Z(c[125]) );
  XOR U1505 ( .A(sreg[129]), .B(n1369), .Z(n1372) );
  XNOR U1506 ( .A(n1369), .B(n1375), .Z(n1371) );
  XOR U1507 ( .A(n1376), .B(n1377), .Z(n1375) );
  NAND U1508 ( .A(b[0]), .B(a[1]), .Z(n1377) );
  AND U1509 ( .A(a[0]), .B(b[1]), .Z(n1376) );
  ANDN U1510 ( .B(sreg[128]), .A(n1378), .Z(n1369) );
  XNOR U1511 ( .A(sreg[128]), .B(n1378), .Z(c[124]) );
  NAND U1512 ( .A(a[0]), .B(b[0]), .Z(n1378) );
endmodule

