
module mult_N64_CC2 ( clk, rst, a, b, c );
  input [63:0] a;
  input [31:0] b;
  output [63:0] c;
  input clk, rst;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72,
         n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86,
         n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100,
         n101, n102, n103, n104, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n121, n122,
         n123, n124, n125, n126, n127, n128, n129, n130, n131, n132, n133,
         n134, n135, n136, n137, n138, n139, n140, n141, n142, n143, n144,
         n145, n146, n147, n148, n149, n150, n151, n152, n153, n154, n155,
         n156, n157, n158, n159, n160, n161, n162, n163, n164, n165, n166,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n177,
         n178, n179, n180, n181, n182, n183, n184, n185, n186, n187, n188,
         n189, n190, n191, n192, n193, n194, n195, n196, n197, n198, n199,
         n200, n201, n202, n203, n204, n205, n206, n207, n208, n209, n210,
         n211, n212, n213, n214, n215, n216, n217, n218, n219, n220, n221,
         n222, n223, n224, n225, n226, n227, n228, n229, n230, n231, n232,
         n233, n234, n235, n236, n237, n238, n239, n240, n241, n242, n243,
         n244, n245, n246, n247, n248, n249, n250, n251, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n274, n275, n276,
         n277, n278, n279, n280, n281, n282, n283, n284, n285, n286, n287,
         n288, n289, n290, n291, n292, n293, n294, n295, n296, n297, n298,
         n299, n300, n301, n302, n303, n304, n305, n306, n307, n308, n309,
         n310, n311, n312, n313, n314, n315, n316, n317, n318, n319, n320,
         n321, n322, n323, n324, n325, n326, n327, n328, n329, n330, n331,
         n332, n333, n334, n335, n336, n337, n338, n339, n340, n341, n342,
         n343, n344, n345, n346, n347, n348, n349, n350, n351, n352, n353,
         n354, n355, n356, n357, n358, n359, n360, n361, n362, n363, n364,
         n365, n366, n367, n368, n369, n370, n371, n372, n373, n374, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, n399, n400, n401, n402, n403, n404, n405, n406, n407, n408,
         n409, n410, n411, n412, n413, n414, n415, n416, n417, n418, n419,
         n420, n421, n422, n423, n424, n425, n426, n427, n428, n429, n430,
         n431, n432, n433, n434, n435, n436, n437, n438, n439, n440, n441,
         n442, n443, n444, n445, n446, n447, n448, n449, n450, n451, n452,
         n453, n454, n455, n456, n457, n458, n459, n460, n461, n462, n463,
         n464, n465, n466, n467, n468, n469, n470, n471, n472, n473, n474,
         n475, n476, n477, n478, n479, n480, n481, n482, n483, n484, n485,
         n486, n487, n488, n489, n490, n491, n492, n493, n494, n495, n496,
         n497, n498, n499, n500, n501, n502, n503, n504, n505, n506, n507,
         n508, n509, n510, n511, n512, n513, n514, n515, n516, n517, n518,
         n519, n520, n521, n522, n523, n524, n525, n526, n527, n528, n529,
         n530, n531, n532, n533, n534, n535, n536, n537, n538, n539, n540,
         n541, n542, n543, n544, n545, n546, n547, n548, n549, n550, n551,
         n552, n553, n554, n555, n556, n557, n558, n559, n560, n561, n562,
         n563, n564, n565, n566, n567, n568, n569, n570, n571, n572, n573,
         n574, n575, n576, n577, n578, n579, n580, n581, n582, n583, n584,
         n585, n586, n587, n588, n589, n590, n591, n592, n593, n594, n595,
         n596, n597, n598, n599, n600, n601, n602, n603, n604, n605, n606,
         n607, n608, n609, n610, n611, n612, n613, n614, n615, n616, n617,
         n618, n619, n620, n621, n622, n623, n624, n625, n626, n627, n628,
         n629, n630, n631, n632, n633, n634, n635, n636, n637, n638, n639,
         n640, n641, n642, n643, n644, n645, n646, n647, n648, n649, n650,
         n651, n652, n653, n654, n655, n656, n657, n658, n659, n660, n661,
         n662, n663, n664, n665, n666, n667, n668, n669, n670, n671, n672,
         n673, n674, n675, n676, n677, n678, n679, n680, n681, n682, n683,
         n684, n685, n686, n687, n688, n689, n690, n691, n692, n693, n694,
         n695, n696, n697, n698, n699, n700, n701, n702, n703, n704, n705,
         n706, n707, n708, n709, n710, n711, n712, n713, n714, n715, n716,
         n717, n718, n719, n720, n721, n722, n723, n724, n725, n726, n727,
         n728, n729, n730, n731, n732, n733, n734, n735, n736, n737, n738,
         n739, n740, n741, n742, n743, n744, n745, n746, n747, n748, n749,
         n750, n751, n752, n753, n754, n755, n756, n757, n758, n759, n760,
         n761, n762, n763, n764, n765, n766, n767, n768, n769, n770, n771,
         n772, n773, n774, n775, n776, n777, n778, n779, n780, n781, n782,
         n783, n784, n785, n786, n787, n788, n789, n790, n791, n792, n793,
         n794, n795, n796, n797, n798, n799, n800, n801, n802, n803, n804,
         n805, n806, n807, n808, n809, n810, n811, n812, n813, n814, n815,
         n816, n817, n818, n819, n820, n821, n822, n823, n824, n825, n826,
         n827, n828, n829, n830, n831, n832, n833, n834, n835, n836, n837,
         n838, n839, n840, n841, n842, n843, n844, n845, n846, n847, n848,
         n849, n850, n851, n852, n853, n854, n855, n856, n857, n858, n859,
         n860, n861, n862, n863, n864, n865, n866, n867, n868, n869, n870,
         n871, n872, n873, n874, n875, n876, n877, n878, n879, n880, n881,
         n882, n883, n884, n885, n886, n887, n888, n889, n890, n891, n892,
         n893, n894, n895, n896, n897, n898, n899, n900, n901, n902, n903,
         n904, n905, n906, n907, n908, n909, n910, n911, n912, n913, n914,
         n915, n916, n917, n918, n919, n920, n921, n922, n923, n924, n925,
         n926, n927, n928, n929, n930, n931, n932, n933, n934, n935, n936,
         n937, n938, n939, n940, n941, n942, n943, n944, n945, n946, n947,
         n948, n949, n950, n951, n952, n953, n954, n955, n956, n957, n958,
         n959, n960, n961, n962, n963, n964, n965, n966, n967, n968, n969,
         n970, n971, n972, n973, n974, n975, n976, n977, n978, n979, n980,
         n981, n982, n983, n984, n985, n986, n987, n988, n989, n990, n991,
         n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001, n1002,
         n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011, n1012,
         n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021, n1022,
         n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031, n1032,
         n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041, n1042,
         n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051, n1052,
         n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061, n1062,
         n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071, n1072,
         n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081, n1082,
         n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091, n1092,
         n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101, n1102,
         n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111, n1112,
         n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121, n1122,
         n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131, n1132,
         n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141, n1142,
         n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151, n1152,
         n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160, n1161, n1162,
         n1163, n1164, n1165, n1166, n1167, n1168, n1169, n1170, n1171, n1172,
         n1173, n1174, n1175, n1176, n1177, n1178, n1179, n1180, n1181, n1182,
         n1183, n1184, n1185, n1186, n1187, n1188, n1189, n1190, n1191, n1192,
         n1193, n1194, n1195, n1196, n1197, n1198, n1199, n1200, n1201, n1202,
         n1203, n1204, n1205, n1206, n1207, n1208, n1209, n1210, n1211, n1212,
         n1213, n1214, n1215, n1216, n1217, n1218, n1219, n1220, n1221, n1222,
         n1223, n1224, n1225, n1226, n1227, n1228, n1229, n1230, n1231, n1232,
         n1233, n1234, n1235, n1236, n1237, n1238, n1239, n1240, n1241, n1242,
         n1243, n1244, n1245, n1246, n1247, n1248, n1249, n1250, n1251, n1252,
         n1253, n1254, n1255, n1256, n1257, n1258, n1259, n1260, n1261, n1262,
         n1263, n1264, n1265, n1266, n1267, n1268, n1269, n1270, n1271, n1272,
         n1273, n1274, n1275, n1276, n1277, n1278, n1279, n1280, n1281, n1282,
         n1283, n1284, n1285, n1286, n1287, n1288, n1289, n1290, n1291, n1292,
         n1293, n1294, n1295, n1296, n1297, n1298, n1299, n1300, n1301, n1302,
         n1303, n1304, n1305, n1306, n1307, n1308, n1309, n1310, n1311, n1312,
         n1313, n1314, n1315, n1316, n1317, n1318, n1319, n1320, n1321, n1322,
         n1323, n1324, n1325, n1326, n1327, n1328, n1329, n1330, n1331, n1332,
         n1333, n1334, n1335, n1336, n1337, n1338, n1339, n1340, n1341, n1342,
         n1343, n1344, n1345, n1346, n1347, n1348, n1349, n1350, n1351, n1352,
         n1353, n1354, n1355, n1356, n1357, n1358, n1359, n1360, n1361, n1362,
         n1363, n1364, n1365, n1366, n1367, n1368, n1369, n1370, n1371, n1372,
         n1373, n1374, n1375, n1376, n1377, n1378, n1379, n1380, n1381, n1382,
         n1383, n1384, n1385, n1386, n1387, n1388, n1389, n1390, n1391, n1392,
         n1393, n1394, n1395, n1396, n1397, n1398, n1399, n1400, n1401, n1402,
         n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411, n1412,
         n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421, n1422,
         n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431, n1432,
         n1433, n1434, n1435, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1456, n1457, n1458, n1459, n1460, n1461, n1462,
         n1463, n1464, n1465, n1466, n1467, n1468, n1469, n1470, n1471, n1472,
         n1473, n1474, n1475, n1476, n1477, n1478, n1479, n1480, n1481, n1482,
         n1483, n1484, n1485, n1486, n1487, n1488, n1489, n1490, n1491, n1492,
         n1493, n1494, n1495, n1496, n1497, n1498, n1499, n1500, n1501, n1502,
         n1503, n1504, n1505, n1506, n1507, n1508, n1509, n1510, n1511, n1512,
         n1513, n1514, n1515, n1516, n1517, n1518, n1519, n1520, n1521, n1522,
         n1523, n1524, n1525, n1526, n1527, n1528, n1529, n1530, n1531, n1532,
         n1533, n1534, n1535, n1536, n1537, n1538, n1539, n1540, n1541, n1542,
         n1543, n1544, n1545, n1546, n1547, n1548, n1549, n1550, n1551, n1552,
         n1553, n1554, n1555, n1556, n1557, n1558, n1559, n1560, n1561, n1562,
         n1563, n1564, n1565, n1566, n1567, n1568, n1569, n1570, n1571, n1572,
         n1573, n1574, n1575, n1576, n1577, n1578, n1579, n1580, n1581, n1582,
         n1583, n1584, n1585, n1586, n1587, n1588, n1589, n1590, n1591, n1592,
         n1593, n1594, n1595, n1596, n1597, n1598, n1599, n1600, n1601, n1602,
         n1603, n1604, n1605, n1606, n1607, n1608, n1609, n1610, n1611, n1612,
         n1613, n1614, n1615, n1616, n1617, n1618, n1619, n1620, n1621, n1622,
         n1623, n1624, n1625, n1626, n1627, n1628, n1629, n1630, n1631, n1632,
         n1633, n1634, n1635, n1636, n1637, n1638, n1639, n1640, n1641, n1642,
         n1643, n1644, n1645, n1646, n1647, n1648, n1649, n1650, n1651, n1652,
         n1653, n1654, n1655, n1656, n1657, n1658, n1659, n1660, n1661, n1662,
         n1663, n1664, n1665, n1666, n1667, n1668, n1669, n1670, n1671, n1672,
         n1673, n1674, n1675, n1676, n1677, n1678, n1679, n1680, n1681, n1682,
         n1683, n1684, n1685, n1686, n1687, n1688, n1689, n1690, n1691, n1692,
         n1693, n1694, n1695, n1696, n1697, n1698, n1699, n1700, n1701, n1702,
         n1703, n1704, n1705, n1706, n1707, n1708, n1709, n1710, n1711, n1712,
         n1713, n1714, n1715, n1716, n1717, n1718, n1719, n1720, n1721, n1722,
         n1723, n1724, n1725, n1726, n1727, n1728, n1729, n1730, n1731, n1732,
         n1733, n1734, n1735, n1736, n1737, n1738, n1739, n1740, n1741, n1742,
         n1743, n1744, n1745, n1746, n1747, n1748, n1749, n1750, n1751, n1752,
         n1753, n1754, n1755, n1756, n1757, n1758, n1759, n1760, n1761, n1762,
         n1763, n1764, n1765, n1766, n1767, n1768, n1769, n1770, n1771, n1772,
         n1773, n1774, n1775, n1776, n1777, n1778, n1779, n1780, n1781, n1782,
         n1783, n1784, n1785, n1786, n1787, n1788, n1789, n1790, n1791, n1792,
         n1793, n1794, n1795, n1796, n1797, n1798, n1799, n1800, n1801, n1802,
         n1803, n1804, n1805, n1806, n1807, n1808, n1809, n1810, n1811, n1812,
         n1813, n1814, n1815, n1816, n1817, n1818, n1819, n1820, n1821, n1822,
         n1823, n1824, n1825, n1826, n1827, n1828, n1829, n1830, n1831, n1832,
         n1833, n1834, n1835, n1836, n1837, n1838, n1839, n1840, n1841, n1842,
         n1843, n1844, n1845, n1846, n1847, n1848, n1849, n1850, n1851, n1852,
         n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861, n1862,
         n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871, n1872,
         n1873, n1874, n1875, n1876, n1877, n1878, n1879, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n1989, n1990, n1991, n1992,
         n1993, n1994, n1995, n1996, n1997, n1998, n1999, n2000, n2001, n2002,
         n2003, n2004, n2005, n2006, n2007, n2008, n2009, n2010, n2011, n2012,
         n2013, n2014, n2015, n2016, n2017, n2018, n2019, n2020, n2021, n2022,
         n2023, n2024, n2025, n2026, n2027, n2028, n2029, n2030, n2031, n2032,
         n2033, n2034, n2035, n2036, n2037, n2038, n2039, n2040, n2041, n2042,
         n2043, n2044, n2045, n2046, n2047, n2048, n2049, n2050, n2051, n2052,
         n2053, n2054, n2055, n2056, n2057, n2058, n2059, n2060, n2061, n2062,
         n2063, n2064, n2065, n2066, n2067, n2068, n2069, n2070, n2071, n2072,
         n2073, n2074, n2075, n2076, n2077, n2078, n2079, n2080, n2081, n2082,
         n2083, n2084, n2085, n2086, n2087, n2088, n2089, n2090, n2091, n2092,
         n2093, n2094, n2095, n2096, n2097, n2098, n2099, n2100, n2101, n2102,
         n2103, n2104, n2105, n2106, n2107, n2108, n2109, n2110, n2111, n2112,
         n2113, n2114, n2115, n2116, n2117, n2118, n2119, n2120, n2121, n2122,
         n2123, n2124, n2125, n2126, n2127, n2128, n2129, n2130, n2131, n2132,
         n2133, n2134, n2135, n2136, n2137, n2138, n2139, n2140, n2141, n2142,
         n2143, n2144, n2145, n2146, n2147, n2148, n2149, n2150, n2151, n2152,
         n2153, n2154, n2155, n2156, n2157, n2158, n2159, n2160, n2161, n2162,
         n2163, n2164, n2165, n2166, n2167, n2168, n2169, n2170, n2171, n2172,
         n2173, n2174, n2175, n2176, n2177, n2178, n2179, n2180, n2181, n2182,
         n2183, n2184, n2185, n2186, n2187, n2188, n2189, n2190, n2191, n2192,
         n2193, n2194, n2195, n2196, n2197, n2198, n2199, n2200, n2201, n2202,
         n2203, n2204, n2205, n2206, n2207, n2208, n2209, n2210, n2211, n2212,
         n2213, n2214, n2215, n2216, n2217, n2218, n2219, n2220, n2221, n2222,
         n2223, n2224, n2225, n2226, n2227, n2228, n2229, n2230, n2231, n2232,
         n2233, n2234, n2235, n2236, n2237, n2238, n2239, n2240, n2241, n2242,
         n2243, n2244, n2245, n2246, n2247, n2248, n2249, n2250, n2251, n2252,
         n2253, n2254, n2255, n2256, n2257, n2258, n2259, n2260, n2261, n2262,
         n2263, n2264, n2265, n2266, n2267, n2268, n2269, n2270, n2271, n2272,
         n2273, n2274, n2275, n2276, n2277, n2278, n2279, n2280, n2281, n2282,
         n2283, n2284, n2285, n2286, n2287, n2288, n2289, n2290, n2291, n2292,
         n2293, n2294, n2295, n2296, n2297, n2298, n2299, n2300, n2301, n2302,
         n2303, n2304, n2305, n2306, n2307, n2308, n2309, n2310, n2311, n2312,
         n2313, n2314, n2315, n2316, n2317, n2318, n2319, n2320, n2321, n2322,
         n2323, n2324, n2325, n2326, n2327, n2328, n2329, n2330, n2331, n2332,
         n2333, n2334, n2335, n2336, n2337, n2338, n2339, n2340, n2341, n2342,
         n2343, n2344, n2345, n2346, n2347, n2348, n2349, n2350, n2351, n2352,
         n2353, n2354, n2355, n2356, n2357, n2358, n2359, n2360, n2361, n2362,
         n2363, n2364, n2365, n2366, n2367, n2368, n2369, n2370, n2371, n2372,
         n2373, n2374, n2375, n2376, n2377, n2378, n2379, n2380, n2381, n2382,
         n2383, n2384, n2385, n2386, n2387, n2388, n2389, n2390, n2391, n2392,
         n2393, n2394, n2395, n2396, n2397, n2398, n2399, n2400, n2401, n2402,
         n2403, n2404, n2405, n2406, n2407, n2408, n2409, n2410, n2411, n2412,
         n2413, n2414, n2415, n2416, n2417, n2418, n2419, n2420, n2421, n2422,
         n2423, n2424, n2425, n2426, n2427, n2428, n2429, n2430, n2431, n2432,
         n2433, n2434, n2435, n2436, n2437, n2438, n2439, n2440, n2441, n2442,
         n2443, n2444, n2445, n2446, n2447, n2448, n2449, n2450, n2451, n2452,
         n2453, n2454, n2455, n2456, n2457, n2458, n2459, n2460, n2461, n2462,
         n2463, n2464, n2465, n2466, n2467, n2468, n2469, n2470, n2471, n2472,
         n2473, n2474, n2475, n2476, n2477, n2478, n2479, n2480, n2481, n2482,
         n2483, n2484, n2485, n2486, n2487, n2488, n2489, n2490, n2491, n2492,
         n2493, n2494, n2495, n2496, n2497, n2498, n2499, n2500, n2501, n2502,
         n2503, n2504, n2505, n2506, n2507, n2508, n2509, n2510, n2511, n2512,
         n2513, n2514, n2515, n2516, n2517, n2518, n2519, n2520, n2521, n2522,
         n2523, n2524, n2525, n2526, n2527, n2528, n2529, n2530, n2531, n2532,
         n2533, n2534, n2535, n2536, n2537, n2538, n2539, n2540, n2541, n2542,
         n2543, n2544, n2545, n2546, n2547, n2548, n2549, n2550, n2551, n2552,
         n2553, n2554, n2555, n2556, n2557, n2558, n2559, n2560, n2561, n2562,
         n2563, n2564, n2565, n2566, n2567, n2568, n2569, n2570, n2571, n2572,
         n2573, n2574, n2575, n2576, n2577, n2578, n2579, n2580, n2581, n2582,
         n2583, n2584, n2585, n2586, n2587, n2588, n2589, n2590, n2591, n2592,
         n2593, n2594, n2595, n2596, n2597, n2598, n2599, n2600, n2601, n2602,
         n2603, n2604, n2605, n2606, n2607, n2608, n2609, n2610, n2611, n2612,
         n2613, n2614, n2615, n2616, n2617, n2618, n2619, n2620, n2621, n2622,
         n2623, n2624, n2625, n2626, n2627, n2628, n2629, n2630, n2631, n2632,
         n2633, n2634, n2635, n2636, n2637, n2638, n2639, n2640, n2641, n2642,
         n2643, n2644, n2645, n2646, n2647, n2648, n2649, n2650, n2651, n2652,
         n2653, n2654, n2655, n2656, n2657, n2658, n2659, n2660, n2661, n2662,
         n2663, n2664, n2665, n2666, n2667, n2668, n2669, n2670, n2671, n2672,
         n2673, n2674, n2675, n2676, n2677, n2678, n2679, n2680, n2681, n2682,
         n2683, n2684, n2685, n2686, n2687, n2688, n2689, n2690, n2691, n2692,
         n2693, n2694, n2695, n2696, n2697, n2698, n2699, n2700, n2701, n2702,
         n2703, n2704, n2705, n2706, n2707, n2708, n2709, n2710, n2711, n2712,
         n2713, n2714, n2715, n2716, n2717, n2718, n2719, n2720, n2721, n2722,
         n2723, n2724, n2725, n2726, n2727, n2728, n2729, n2730, n2731, n2732,
         n2733, n2734, n2735, n2736, n2737, n2738, n2739, n2740, n2741, n2742,
         n2743, n2744, n2745, n2746, n2747, n2748, n2749, n2750, n2751, n2752,
         n2753, n2754, n2755, n2756, n2757, n2758, n2759, n2760, n2761, n2762,
         n2763, n2764, n2765, n2766, n2767, n2768, n2769, n2770, n2771, n2772,
         n2773, n2774, n2775, n2776, n2777, n2778, n2779, n2780, n2781, n2782,
         n2783, n2784, n2785, n2786, n2787, n2788, n2789, n2790, n2791, n2792,
         n2793, n2794, n2795, n2796, n2797, n2798, n2799, n2800, n2801, n2802,
         n2803, n2804, n2805, n2806, n2807, n2808, n2809, n2810, n2811, n2812,
         n2813, n2814, n2815, n2816, n2817, n2818, n2819, n2820, n2821, n2822,
         n2823, n2824, n2825, n2826, n2827, n2828, n2829, n2830, n2831, n2832,
         n2833, n2834, n2835, n2836, n2837, n2838, n2839, n2840, n2841, n2842,
         n2843, n2844, n2845, n2846, n2847, n2848, n2849, n2850, n2851, n2852,
         n2853, n2854, n2855, n2856, n2857, n2858, n2859, n2860, n2861, n2862,
         n2863, n2864, n2865, n2866, n2867, n2868, n2869, n2870, n2871, n2872,
         n2873, n2874, n2875, n2876, n2877, n2878, n2879, n2880, n2881, n2882,
         n2883, n2884, n2885, n2886, n2887, n2888, n2889, n2890, n2891, n2892,
         n2893, n2894, n2895, n2896, n2897, n2898, n2899, n2900, n2901, n2902,
         n2903, n2904, n2905, n2906, n2907, n2908, n2909, n2910, n2911, n2912,
         n2913, n2914, n2915, n2916, n2917, n2918, n2919, n2920, n2921, n2922,
         n2923, n2924, n2925, n2926, n2927, n2928, n2929, n2930, n2931, n2932,
         n2933, n2934, n2935, n2936, n2937, n2938, n2939, n2940, n2941, n2942,
         n2943, n2944, n2945, n2946, n2947, n2948, n2949, n2950, n2951, n2952,
         n2953, n2954, n2955, n2956, n2957, n2958, n2959, n2960, n2961, n2962,
         n2963, n2964, n2965, n2966, n2967, n2968, n2969, n2970, n2971, n2972,
         n2973, n2974, n2975, n2976, n2977, n2978, n2979, n2980, n2981, n2982,
         n2983, n2984, n2985, n2986, n2987, n2988, n2989, n2990, n2991, n2992,
         n2993, n2994, n2995, n2996, n2997, n2998, n2999, n3000, n3001, n3002,
         n3003, n3004, n3005, n3006, n3007, n3008, n3009, n3010, n3011, n3012,
         n3013, n3014, n3015, n3016, n3017, n3018, n3019, n3020, n3021, n3022,
         n3023, n3024, n3025, n3026, n3027, n3028, n3029, n3030, n3031, n3032,
         n3033, n3034, n3035, n3036, n3037, n3038, n3039, n3040, n3041, n3042,
         n3043, n3044, n3045, n3046, n3047, n3048, n3049, n3050, n3051, n3052,
         n3053, n3054, n3055, n3056, n3057, n3058, n3059, n3060, n3061, n3062,
         n3063, n3064, n3065, n3066, n3067, n3068, n3069, n3070, n3071, n3072,
         n3073, n3074, n3075, n3076, n3077, n3078, n3079, n3080, n3081, n3082,
         n3083, n3084, n3085, n3086, n3087, n3088, n3089, n3090, n3091, n3092,
         n3093, n3094, n3095, n3096, n3097, n3098, n3099, n3100, n3101, n3102,
         n3103, n3104, n3105, n3106, n3107, n3108, n3109, n3110, n3111, n3112,
         n3113, n3114, n3115, n3116, n3117, n3118, n3119, n3120, n3121, n3122,
         n3123, n3124, n3125, n3126, n3127, n3128, n3129, n3130, n3131, n3132,
         n3133, n3134, n3135, n3136, n3137, n3138, n3139, n3140, n3141, n3142,
         n3143, n3144, n3145, n3146, n3147, n3148, n3149, n3150, n3151, n3152,
         n3153, n3154, n3155, n3156, n3157, n3158, n3159, n3160, n3161, n3162,
         n3163, n3164, n3165, n3166, n3167, n3168, n3169, n3170, n3171, n3172,
         n3173, n3174, n3175, n3176, n3177, n3178, n3179, n3180, n3181, n3182,
         n3183, n3184, n3185, n3186, n3187, n3188, n3189, n3190, n3191, n3192,
         n3193, n3194, n3195, n3196, n3197, n3198, n3199, n3200, n3201, n3202,
         n3203, n3204, n3205, n3206, n3207, n3208, n3209, n3210, n3211, n3212,
         n3213, n3214, n3215, n3216, n3217, n3218, n3219, n3220, n3221, n3222,
         n3223, n3224, n3225, n3226, n3227, n3228, n3229, n3230, n3231, n3232,
         n3233, n3234, n3235, n3236, n3237, n3238, n3239, n3240, n3241, n3242,
         n3243, n3244, n3245, n3246, n3247, n3248, n3249, n3250, n3251, n3252,
         n3253, n3254, n3255, n3256, n3257, n3258, n3259, n3260, n3261, n3262,
         n3263, n3264, n3265, n3266, n3267, n3268, n3269, n3270, n3271, n3272,
         n3273, n3274, n3275, n3276, n3277, n3278, n3279, n3280, n3281, n3282,
         n3283, n3284, n3285, n3286, n3287, n3288, n3289, n3290, n3291, n3292,
         n3293, n3294, n3295, n3296, n3297, n3298, n3299, n3300, n3301, n3302,
         n3303, n3304, n3305, n3306, n3307, n3308, n3309, n3310, n3311, n3312,
         n3313, n3314, n3315, n3316, n3317, n3318, n3319, n3320, n3321, n3322,
         n3323, n3324, n3325, n3326, n3327, n3328, n3329, n3330, n3331, n3332,
         n3333, n3334, n3335, n3336, n3337, n3338, n3339, n3340, n3341, n3342,
         n3343, n3344, n3345, n3346, n3347, n3348, n3349, n3350, n3351, n3352,
         n3353, n3354, n3355, n3356, n3357, n3358, n3359, n3360, n3361, n3362,
         n3363, n3364, n3365, n3366, n3367, n3368, n3369, n3370, n3371, n3372,
         n3373, n3374, n3375, n3376, n3377, n3378, n3379, n3380, n3381, n3382,
         n3383, n3384, n3385, n3386, n3387, n3388, n3389, n3390, n3391, n3392,
         n3393, n3394, n3395, n3396, n3397, n3398, n3399, n3400, n3401, n3402,
         n3403, n3404, n3405, n3406, n3407, n3408, n3409, n3410, n3411, n3412,
         n3413, n3414, n3415, n3416, n3417, n3418, n3419, n3420, n3421, n3422,
         n3423, n3424, n3425, n3426, n3427, n3428, n3429, n3430, n3431, n3432,
         n3433, n3434, n3435, n3436, n3437, n3438, n3439, n3440, n3441, n3442,
         n3443, n3444, n3445, n3446, n3447, n3448, n3449, n3450, n3451, n3452,
         n3453, n3454, n3455, n3456, n3457, n3458, n3459, n3460, n3461, n3462,
         n3463, n3464, n3465, n3466, n3467, n3468, n3469, n3470, n3471, n3472,
         n3473, n3474, n3475, n3476, n3477, n3478, n3479, n3480, n3481, n3482,
         n3483, n3484, n3485, n3486, n3487, n3488, n3489, n3490, n3491, n3492,
         n3493, n3494, n3495, n3496, n3497, n3498, n3499, n3500, n3501, n3502,
         n3503, n3504, n3505, n3506, n3507, n3508, n3509, n3510, n3511, n3512,
         n3513, n3514, n3515, n3516, n3517, n3518, n3519, n3520, n3521, n3522,
         n3523, n3524, n3525, n3526, n3527, n3528, n3529, n3530, n3531, n3532,
         n3533, n3534, n3535, n3536, n3537, n3538, n3539, n3540, n3541, n3542,
         n3543, n3544, n3545, n3546, n3547, n3548, n3549, n3550, n3551, n3552,
         n3553, n3554, n3555, n3556, n3557, n3558, n3559, n3560, n3561, n3562,
         n3563, n3564, n3565, n3566, n3567, n3568, n3569, n3570, n3571, n3572,
         n3573, n3574, n3575, n3576, n3577, n3578, n3579, n3580, n3581, n3582,
         n3583, n3584, n3585, n3586, n3587, n3588, n3589, n3590, n3591, n3592,
         n3593, n3594, n3595, n3596, n3597, n3598, n3599, n3600, n3601, n3602,
         n3603, n3604, n3605, n3606, n3607, n3608, n3609, n3610, n3611, n3612,
         n3613, n3614, n3615, n3616, n3617, n3618, n3619, n3620, n3621, n3622,
         n3623, n3624, n3625, n3626, n3627, n3628, n3629, n3630, n3631, n3632,
         n3633, n3634, n3635, n3636, n3637, n3638, n3639, n3640, n3641, n3642,
         n3643, n3644, n3645, n3646, n3647, n3648, n3649, n3650, n3651, n3652,
         n3653, n3654, n3655, n3656, n3657, n3658, n3659, n3660, n3661, n3662,
         n3663, n3664, n3665, n3666, n3667, n3668, n3669, n3670, n3671, n3672,
         n3673, n3674, n3675, n3676, n3677, n3678, n3679, n3680, n3681, n3682,
         n3683, n3684, n3685, n3686, n3687, n3688, n3689, n3690, n3691, n3692,
         n3693, n3694, n3695, n3696, n3697, n3698, n3699, n3700, n3701, n3702,
         n3703, n3704, n3705, n3706, n3707, n3708, n3709, n3710, n3711, n3712,
         n3713, n3714, n3715, n3716, n3717, n3718, n3719, n3720, n3721, n3722,
         n3723, n3724, n3725, n3726, n3727, n3728, n3729, n3730, n3731, n3732,
         n3733, n3734, n3735, n3736, n3737, n3738, n3739, n3740, n3741, n3742,
         n3743, n3744, n3745, n3746, n3747, n3748, n3749, n3750, n3751, n3752,
         n3753, n3754, n3755, n3756, n3757, n3758, n3759, n3760, n3761, n3762,
         n3763, n3764, n3765, n3766, n3767, n3768, n3769, n3770, n3771, n3772,
         n3773, n3774, n3775, n3776, n3777, n3778, n3779, n3780, n3781, n3782,
         n3783, n3784, n3785, n3786, n3787, n3788, n3789, n3790, n3791, n3792,
         n3793, n3794, n3795, n3796, n3797, n3798, n3799, n3800, n3801, n3802,
         n3803, n3804, n3805, n3806, n3807, n3808, n3809, n3810, n3811, n3812,
         n3813, n3814, n3815, n3816, n3817, n3818, n3819, n3820, n3821, n3822,
         n3823, n3824, n3825, n3826, n3827, n3828, n3829, n3830, n3831, n3832,
         n3833, n3834, n3835, n3836, n3837, n3838, n3839, n3840, n3841, n3842,
         n3843, n3844, n3845, n3846, n3847, n3848, n3849, n3850, n3851, n3852,
         n3853, n3854, n3855, n3856, n3857, n3858, n3859, n3860, n3861, n3862,
         n3863, n3864, n3865, n3866, n3867, n3868, n3869, n3870, n3871, n3872,
         n3873, n3874, n3875, n3876, n3877, n3878, n3879, n3880, n3881, n3882,
         n3883, n3884, n3885, n3886, n3887, n3888, n3889, n3890, n3891, n3892,
         n3893, n3894, n3895, n3896, n3897, n3898, n3899, n3900, n3901, n3902,
         n3903, n3904, n3905, n3906, n3907, n3908, n3909, n3910, n3911, n3912,
         n3913, n3914, n3915, n3916, n3917, n3918, n3919, n3920, n3921, n3922,
         n3923, n3924, n3925, n3926, n3927, n3928, n3929, n3930, n3931, n3932,
         n3933, n3934, n3935, n3936, n3937, n3938, n3939, n3940, n3941, n3942,
         n3943, n3944, n3945, n3946, n3947, n3948, n3949, n3950, n3951, n3952,
         n3953, n3954, n3955, n3956, n3957, n3958, n3959, n3960, n3961, n3962,
         n3963, n3964, n3965, n3966, n3967, n3968, n3969, n3970, n3971, n3972,
         n3973, n3974, n3975, n3976, n3977, n3978, n3979, n3980, n3981, n3982,
         n3983, n3984, n3985, n3986, n3987, n3988, n3989, n3990, n3991, n3992,
         n3993, n3994, n3995, n3996, n3997, n3998, n3999, n4000, n4001, n4002,
         n4003, n4004, n4005, n4006, n4007, n4008, n4009, n4010, n4011, n4012,
         n4013, n4014, n4015, n4016, n4017, n4018, n4019, n4020, n4021, n4022,
         n4023, n4024, n4025, n4026, n4027, n4028, n4029, n4030, n4031, n4032,
         n4033, n4034, n4035, n4036, n4037, n4038, n4039, n4040, n4041, n4042,
         n4043, n4044, n4045, n4046, n4047, n4048, n4049, n4050, n4051, n4052,
         n4053, n4054, n4055, n4056, n4057, n4058, n4059, n4060, n4061, n4062,
         n4063, n4064, n4065, n4066, n4067, n4068, n4069, n4070, n4071, n4072,
         n4073, n4074, n4075, n4076, n4077, n4078, n4079, n4080, n4081, n4082,
         n4083, n4084, n4085, n4086, n4087, n4088, n4089, n4090, n4091, n4092,
         n4093, n4094, n4095, n4096, n4097, n4098, n4099, n4100, n4101, n4102,
         n4103, n4104, n4105, n4106, n4107, n4108, n4109, n4110, n4111, n4112,
         n4113, n4114, n4115, n4116, n4117, n4118, n4119, n4120, n4121, n4122,
         n4123, n4124, n4125, n4126, n4127, n4128, n4129, n4130, n4131, n4132,
         n4133, n4134, n4135, n4136, n4137, n4138, n4139, n4140, n4141, n4142,
         n4143, n4144, n4145, n4146, n4147, n4148, n4149, n4150, n4151, n4152,
         n4153, n4154, n4155, n4156, n4157, n4158, n4159, n4160, n4161, n4162,
         n4163, n4164, n4165, n4166, n4167, n4168, n4169, n4170, n4171, n4172,
         n4173, n4174, n4175, n4176, n4177, n4178, n4179, n4180, n4181, n4182,
         n4183, n4184, n4185, n4186, n4187, n4188, n4189, n4190, n4191, n4192,
         n4193, n4194, n4195, n4196, n4197, n4198, n4199, n4200, n4201, n4202,
         n4203, n4204, n4205, n4206, n4207, n4208, n4209, n4210, n4211, n4212,
         n4213, n4214, n4215, n4216, n4217, n4218, n4219, n4220, n4221, n4222,
         n4223, n4224, n4225, n4226, n4227, n4228, n4229, n4230, n4231, n4232,
         n4233, n4234, n4235, n4236, n4237, n4238, n4239, n4240, n4241, n4242,
         n4243, n4244, n4245, n4246, n4247, n4248, n4249, n4250, n4251, n4252,
         n4253, n4254, n4255, n4256, n4257, n4258, n4259, n4260, n4261, n4262,
         n4263, n4264, n4265, n4266, n4267, n4268, n4269, n4270, n4271, n4272,
         n4273, n4274, n4275, n4276, n4277, n4278, n4279, n4280, n4281, n4282,
         n4283, n4284, n4285, n4286, n4287, n4288, n4289, n4290, n4291, n4292,
         n4293, n4294, n4295, n4296, n4297, n4298, n4299, n4300, n4301, n4302,
         n4303, n4304, n4305, n4306, n4307, n4308, n4309, n4310, n4311, n4312,
         n4313, n4314, n4315, n4316, n4317, n4318, n4319, n4320, n4321, n4322,
         n4323, n4324, n4325, n4326, n4327, n4328, n4329, n4330, n4331, n4332,
         n4333, n4334, n4335, n4336, n4337, n4338, n4339, n4340, n4341, n4342,
         n4343, n4344, n4345, n4346, n4347, n4348, n4349, n4350, n4351, n4352,
         n4353, n4354, n4355, n4356, n4357, n4358, n4359, n4360, n4361, n4362,
         n4363, n4364, n4365, n4366, n4367, n4368, n4369, n4370, n4371, n4372,
         n4373, n4374, n4375, n4376, n4377, n4378, n4379, n4380, n4381, n4382,
         n4383, n4384, n4385, n4386, n4387, n4388, n4389, n4390, n4391, n4392,
         n4393, n4394, n4395, n4396, n4397, n4398, n4399, n4400, n4401, n4402,
         n4403, n4404, n4405, n4406, n4407, n4408, n4409, n4410, n4411, n4412,
         n4413, n4414, n4415, n4416, n4417, n4418, n4419, n4420, n4421, n4422,
         n4423, n4424, n4425, n4426, n4427, n4428, n4429, n4430, n4431, n4432,
         n4433, n4434, n4435, n4436, n4437, n4438, n4439, n4440, n4441, n4442,
         n4443, n4444, n4445, n4446, n4447, n4448, n4449, n4450, n4451, n4452,
         n4453, n4454, n4455, n4456, n4457, n4458, n4459, n4460, n4461, n4462,
         n4463, n4464, n4465, n4466, n4467, n4468, n4469, n4470, n4471, n4472,
         n4473, n4474, n4475, n4476, n4477, n4478, n4479, n4480, n4481, n4482,
         n4483, n4484, n4485, n4486, n4487, n4488, n4489, n4490, n4491, n4492,
         n4493, n4494, n4495, n4496, n4497, n4498, n4499, n4500, n4501, n4502,
         n4503, n4504, n4505, n4506, n4507, n4508, n4509, n4510, n4511, n4512,
         n4513, n4514, n4515, n4516, n4517, n4518, n4519, n4520, n4521, n4522,
         n4523, n4524, n4525, n4526, n4527, n4528, n4529, n4530, n4531, n4532,
         n4533, n4534, n4535, n4536, n4537, n4538, n4539, n4540, n4541, n4542,
         n4543, n4544, n4545, n4546, n4547, n4548, n4549, n4550, n4551, n4552,
         n4553, n4554, n4555, n4556, n4557, n4558, n4559, n4560, n4561, n4562,
         n4563, n4564, n4565, n4566, n4567, n4568, n4569, n4570, n4571, n4572,
         n4573, n4574, n4575, n4576, n4577, n4578, n4579, n4580, n4581, n4582,
         n4583, n4584, n4585, n4586, n4587, n4588, n4589, n4590, n4591, n4592,
         n4593, n4594, n4595, n4596, n4597, n4598, n4599, n4600, n4601, n4602,
         n4603, n4604, n4605, n4606, n4607, n4608, n4609, n4610, n4611, n4612,
         n4613, n4614, n4615, n4616, n4617, n4618, n4619, n4620, n4621, n4622,
         n4623, n4624, n4625, n4626, n4627, n4628, n4629, n4630, n4631, n4632,
         n4633, n4634, n4635, n4636, n4637, n4638, n4639, n4640, n4641, n4642,
         n4643, n4644, n4645, n4646, n4647, n4648, n4649, n4650, n4651, n4652,
         n4653, n4654, n4655, n4656, n4657, n4658, n4659, n4660, n4661, n4662,
         n4663, n4664, n4665, n4666, n4667, n4668, n4669, n4670, n4671, n4672,
         n4673, n4674, n4675, n4676, n4677, n4678, n4679, n4680, n4681, n4682,
         n4683, n4684, n4685, n4686, n4687, n4688, n4689, n4690, n4691, n4692,
         n4693, n4694, n4695, n4696, n4697, n4698, n4699, n4700, n4701, n4702,
         n4703, n4704, n4705, n4706, n4707, n4708, n4709, n4710, n4711, n4712,
         n4713, n4714, n4715, n4716, n4717, n4718, n4719, n4720, n4721, n4722,
         n4723, n4724, n4725, n4726, n4727, n4728, n4729, n4730, n4731, n4732,
         n4733, n4734, n4735, n4736, n4737, n4738, n4739, n4740, n4741, n4742,
         n4743, n4744, n4745, n4746, n4747, n4748, n4749, n4750, n4751, n4752,
         n4753, n4754, n4755, n4756, n4757, n4758, n4759, n4760, n4761, n4762,
         n4763, n4764, n4765, n4766, n4767, n4768, n4769, n4770, n4771, n4772,
         n4773, n4774, n4775, n4776, n4777, n4778, n4779, n4780, n4781, n4782,
         n4783, n4784, n4785, n4786, n4787, n4788, n4789, n4790, n4791, n4792,
         n4793, n4794, n4795, n4796, n4797, n4798, n4799, n4800, n4801, n4802,
         n4803, n4804, n4805, n4806, n4807, n4808, n4809, n4810, n4811, n4812,
         n4813, n4814, n4815, n4816, n4817, n4818, n4819, n4820, n4821, n4822,
         n4823, n4824, n4825, n4826, n4827, n4828, n4829, n4830, n4831, n4832,
         n4833, n4834, n4835, n4836, n4837, n4838, n4839, n4840, n4841, n4842,
         n4843, n4844, n4845, n4846, n4847, n4848, n4849, n4850, n4851, n4852,
         n4853, n4854, n4855, n4856, n4857, n4858, n4859, n4860, n4861, n4862,
         n4863, n4864, n4865, n4866, n4867, n4868, n4869, n4870, n4871, n4872,
         n4873, n4874, n4875, n4876, n4877, n4878, n4879, n4880, n4881, n4882,
         n4883, n4884, n4885, n4886, n4887, n4888, n4889, n4890, n4891, n4892,
         n4893, n4894, n4895, n4896, n4897, n4898, n4899, n4900, n4901, n4902,
         n4903, n4904, n4905, n4906, n4907, n4908, n4909, n4910, n4911, n4912,
         n4913, n4914, n4915, n4916, n4917, n4918, n4919, n4920, n4921, n4922,
         n4923, n4924, n4925, n4926, n4927, n4928, n4929, n4930, n4931, n4932,
         n4933, n4934, n4935, n4936, n4937, n4938, n4939, n4940, n4941, n4942,
         n4943, n4944, n4945, n4946, n4947, n4948, n4949, n4950, n4951, n4952,
         n4953, n4954, n4955, n4956, n4957, n4958, n4959, n4960, n4961, n4962,
         n4963, n4964, n4965, n4966, n4967, n4968, n4969, n4970, n4971, n4972,
         n4973, n4974, n4975, n4976, n4977, n4978, n4979, n4980, n4981, n4982,
         n4983, n4984, n4985, n4986, n4987, n4988, n4989, n4990, n4991, n4992,
         n4993, n4994, n4995, n4996, n4997, n4998, n4999, n5000, n5001, n5002,
         n5003, n5004, n5005, n5006, n5007, n5008, n5009, n5010, n5011, n5012,
         n5013, n5014, n5015, n5016, n5017, n5018, n5019, n5020, n5021, n5022,
         n5023, n5024, n5025, n5026, n5027, n5028, n5029, n5030, n5031, n5032,
         n5033, n5034, n5035, n5036, n5037, n5038, n5039, n5040, n5041, n5042,
         n5043, n5044, n5045, n5046, n5047, n5048, n5049, n5050, n5051, n5052,
         n5053, n5054, n5055, n5056, n5057, n5058, n5059, n5060, n5061, n5062,
         n5063, n5064, n5065, n5066, n5067, n5068, n5069, n5070, n5071, n5072,
         n5073, n5074, n5075, n5076, n5077, n5078, n5079, n5080, n5081, n5082,
         n5083, n5084, n5085, n5086, n5087, n5088, n5089, n5090, n5091, n5092,
         n5093, n5094, n5095, n5096, n5097, n5098, n5099, n5100, n5101, n5102,
         n5103, n5104, n5105, n5106, n5107, n5108, n5109, n5110, n5111, n5112,
         n5113, n5114, n5115, n5116, n5117, n5118, n5119, n5120, n5121, n5122,
         n5123, n5124, n5125, n5126, n5127, n5128, n5129, n5130, n5131, n5132,
         n5133, n5134, n5135, n5136, n5137, n5138, n5139, n5140, n5141, n5142,
         n5143, n5144, n5145, n5146, n5147, n5148, n5149, n5150, n5151, n5152,
         n5153, n5154, n5155, n5156, n5157, n5158, n5159, n5160, n5161, n5162,
         n5163, n5164, n5165, n5166, n5167, n5168, n5169, n5170, n5171, n5172,
         n5173, n5174, n5175, n5176, n5177, n5178, n5179, n5180, n5181, n5182,
         n5183, n5184, n5185, n5186, n5187, n5188, n5189, n5190, n5191, n5192,
         n5193, n5194, n5195, n5196, n5197, n5198, n5199, n5200, n5201, n5202,
         n5203, n5204, n5205, n5206, n5207, n5208, n5209, n5210, n5211, n5212,
         n5213, n5214, n5215, n5216, n5217, n5218, n5219, n5220, n5221, n5222,
         n5223, n5224, n5225, n5226, n5227, n5228, n5229, n5230, n5231, n5232,
         n5233, n5234, n5235, n5236, n5237, n5238, n5239, n5240, n5241, n5242,
         n5243, n5244, n5245, n5246, n5247, n5248, n5249, n5250, n5251, n5252,
         n5253, n5254, n5255, n5256, n5257, n5258, n5259, n5260, n5261, n5262,
         n5263, n5264, n5265, n5266, n5267, n5268, n5269, n5270, n5271, n5272,
         n5273, n5274, n5275, n5276, n5277, n5278, n5279, n5280, n5281, n5282,
         n5283, n5284, n5285, n5286, n5287, n5288, n5289, n5290, n5291, n5292,
         n5293, n5294, n5295, n5296, n5297, n5298, n5299, n5300, n5301, n5302,
         n5303, n5304, n5305, n5306, n5307, n5308, n5309, n5310, n5311, n5312,
         n5313, n5314, n5315, n5316, n5317, n5318, n5319, n5320, n5321, n5322,
         n5323, n5324, n5325, n5326, n5327, n5328, n5329, n5330, n5331, n5332,
         n5333, n5334, n5335, n5336, n5337, n5338, n5339, n5340, n5341, n5342,
         n5343, n5344, n5345, n5346, n5347, n5348, n5349, n5350, n5351, n5352,
         n5353, n5354, n5355, n5356, n5357, n5358, n5359, n5360, n5361, n5362,
         n5363, n5364, n5365, n5366, n5367, n5368, n5369, n5370, n5371, n5372,
         n5373, n5374, n5375, n5376, n5377, n5378, n5379, n5380, n5381, n5382,
         n5383, n5384, n5385, n5386, n5387, n5388, n5389, n5390, n5391, n5392,
         n5393, n5394, n5395, n5396, n5397, n5398, n5399, n5400, n5401, n5402,
         n5403, n5404, n5405, n5406, n5407, n5408, n5409, n5410, n5411, n5412,
         n5413, n5414, n5415, n5416, n5417, n5418, n5419, n5420, n5421, n5422,
         n5423, n5424, n5425, n5426, n5427, n5428, n5429, n5430, n5431, n5432,
         n5433, n5434, n5435, n5436, n5437, n5438, n5439, n5440, n5441, n5442,
         n5443, n5444, n5445, n5446, n5447, n5448, n5449, n5450, n5451, n5452,
         n5453, n5454, n5455, n5456, n5457, n5458, n5459, n5460, n5461, n5462,
         n5463, n5464, n5465, n5466, n5467, n5468, n5469, n5470, n5471, n5472,
         n5473, n5474, n5475, n5476, n5477, n5478, n5479, n5480, n5481, n5482,
         n5483, n5484, n5485, n5486, n5487, n5488, n5489, n5490, n5491, n5492,
         n5493, n5494, n5495, n5496, n5497, n5498, n5499, n5500, n5501, n5502,
         n5503, n5504, n5505, n5506, n5507, n5508, n5509, n5510, n5511, n5512,
         n5513, n5514, n5515, n5516, n5517, n5518, n5519, n5520, n5521, n5522,
         n5523, n5524, n5525, n5526, n5527, n5528, n5529, n5530, n5531, n5532,
         n5533, n5534, n5535, n5536, n5537, n5538, n5539, n5540, n5541, n5542,
         n5543, n5544, n5545, n5546, n5547, n5548, n5549, n5550, n5551, n5552,
         n5553, n5554, n5555, n5556, n5557, n5558, n5559, n5560, n5561, n5562,
         n5563, n5564, n5565, n5566, n5567, n5568, n5569, n5570, n5571, n5572,
         n5573, n5574, n5575, n5576, n5577, n5578, n5579, n5580, n5581, n5582,
         n5583, n5584, n5585, n5586, n5587, n5588, n5589, n5590, n5591, n5592,
         n5593, n5594, n5595, n5596, n5597, n5598, n5599, n5600, n5601, n5602,
         n5603, n5604, n5605, n5606, n5607, n5608, n5609, n5610, n5611, n5612,
         n5613, n5614, n5615, n5616, n5617, n5618, n5619, n5620, n5621, n5622,
         n5623, n5624, n5625, n5626, n5627, n5628, n5629, n5630, n5631, n5632,
         n5633, n5634, n5635, n5636, n5637, n5638, n5639, n5640, n5641, n5642,
         n5643, n5644, n5645, n5646, n5647, n5648, n5649, n5650, n5651, n5652,
         n5653, n5654, n5655, n5656, n5657, n5658, n5659, n5660, n5661, n5662,
         n5663, n5664, n5665, n5666, n5667, n5668, n5669, n5670, n5671, n5672,
         n5673, n5674, n5675, n5676, n5677, n5678, n5679, n5680, n5681, n5682,
         n5683, n5684, n5685, n5686, n5687, n5688, n5689, n5690, n5691, n5692,
         n5693, n5694, n5695, n5696, n5697, n5698, n5699, n5700, n5701, n5702,
         n5703, n5704, n5705, n5706, n5707, n5708, n5709, n5710, n5711, n5712,
         n5713, n5714, n5715, n5716, n5717, n5718, n5719, n5720, n5721, n5722,
         n5723, n5724, n5725, n5726, n5727, n5728, n5729, n5730, n5731, n5732,
         n5733, n5734, n5735, n5736, n5737, n5738, n5739, n5740, n5741, n5742,
         n5743, n5744, n5745, n5746, n5747, n5748, n5749, n5750, n5751, n5752,
         n5753, n5754, n5755, n5756, n5757, n5758, n5759, n5760, n5761, n5762,
         n5763, n5764, n5765, n5766, n5767, n5768, n5769, n5770, n5771, n5772,
         n5773, n5774, n5775, n5776, n5777, n5778, n5779, n5780, n5781, n5782,
         n5783, n5784, n5785, n5786, n5787, n5788, n5789, n5790, n5791, n5792,
         n5793, n5794, n5795, n5796, n5797, n5798, n5799, n5800, n5801, n5802,
         n5803, n5804, n5805, n5806, n5807, n5808, n5809, n5810, n5811, n5812,
         n5813, n5814, n5815, n5816, n5817, n5818, n5819, n5820, n5821, n5822,
         n5823, n5824, n5825, n5826, n5827, n5828, n5829, n5830, n5831, n5832,
         n5833, n5834, n5835, n5836, n5837, n5838, n5839, n5840, n5841, n5842,
         n5843, n5844, n5845, n5846, n5847, n5848, n5849, n5850, n5851, n5852,
         n5853, n5854, n5855, n5856, n5857, n5858, n5859, n5860, n5861, n5862,
         n5863, n5864, n5865, n5866, n5867, n5868, n5869, n5870, n5871, n5872,
         n5873, n5874, n5875, n5876, n5877, n5878, n5879, n5880, n5881, n5882,
         n5883, n5884, n5885, n5886, n5887, n5888, n5889, n5890, n5891, n5892,
         n5893, n5894, n5895, n5896, n5897, n5898, n5899, n5900, n5901, n5902,
         n5903, n5904, n5905, n5906, n5907, n5908, n5909, n5910, n5911, n5912,
         n5913, n5914, n5915, n5916, n5917, n5918, n5919, n5920, n5921, n5922,
         n5923, n5924, n5925, n5926, n5927, n5928, n5929, n5930, n5931, n5932,
         n5933, n5934, n5935, n5936, n5937, n5938, n5939, n5940, n5941, n5942,
         n5943, n5944, n5945, n5946, n5947, n5948, n5949, n5950, n5951, n5952,
         n5953, n5954, n5955, n5956, n5957, n5958, n5959, n5960, n5961, n5962,
         n5963, n5964, n5965, n5966, n5967, n5968, n5969, n5970, n5971, n5972,
         n5973, n5974, n5975, n5976, n5977, n5978, n5979, n5980, n5981, n5982,
         n5983, n5984, n5985, n5986, n5987, n5988, n5989, n5990, n5991, n5992,
         n5993, n5994, n5995, n5996, n5997, n5998, n5999, n6000, n6001, n6002,
         n6003, n6004, n6005, n6006, n6007, n6008, n6009, n6010, n6011, n6012,
         n6013, n6014, n6015, n6016, n6017, n6018, n6019, n6020, n6021, n6022,
         n6023, n6024, n6025, n6026, n6027, n6028, n6029, n6030, n6031, n6032,
         n6033, n6034, n6035, n6036, n6037, n6038, n6039, n6040, n6041, n6042,
         n6043, n6044, n6045, n6046, n6047, n6048, n6049, n6050, n6051, n6052,
         n6053, n6054, n6055, n6056, n6057, n6058, n6059, n6060, n6061, n6062,
         n6063, n6064, n6065, n6066, n6067, n6068, n6069, n6070, n6071, n6072,
         n6073, n6074, n6075, n6076, n6077, n6078, n6079, n6080, n6081, n6082,
         n6083, n6084, n6085, n6086, n6087, n6088, n6089, n6090, n6091, n6092,
         n6093, n6094, n6095, n6096, n6097, n6098, n6099, n6100, n6101, n6102,
         n6103, n6104, n6105, n6106, n6107, n6108, n6109, n6110, n6111, n6112,
         n6113, n6114, n6115, n6116, n6117, n6118, n6119, n6120, n6121, n6122,
         n6123, n6124, n6125, n6126, n6127, n6128, n6129, n6130, n6131, n6132,
         n6133, n6134, n6135, n6136, n6137, n6138, n6139, n6140, n6141, n6142,
         n6143, n6144, n6145, n6146, n6147, n6148, n6149, n6150, n6151, n6152,
         n6153, n6154, n6155, n6156, n6157, n6158, n6159, n6160, n6161, n6162,
         n6163, n6164, n6165, n6166, n6167, n6168, n6169, n6170, n6171, n6172,
         n6173, n6174, n6175, n6176, n6177, n6178, n6179, n6180, n6181, n6182,
         n6183, n6184, n6185, n6186, n6187, n6188, n6189, n6190, n6191, n6192,
         n6193, n6194, n6195, n6196, n6197, n6198, n6199, n6200, n6201, n6202,
         n6203, n6204, n6205, n6206, n6207, n6208, n6209, n6210, n6211, n6212,
         n6213, n6214, n6215, n6216, n6217, n6218, n6219, n6220, n6221, n6222,
         n6223, n6224, n6225, n6226, n6227, n6228, n6229, n6230, n6231, n6232,
         n6233, n6234, n6235, n6236, n6237, n6238, n6239, n6240, n6241, n6242,
         n6243, n6244, n6245, n6246, n6247, n6248, n6249, n6250, n6251, n6252,
         n6253, n6254, n6255, n6256, n6257, n6258, n6259, n6260, n6261, n6262,
         n6263, n6264, n6265, n6266, n6267, n6268, n6269, n6270, n6271, n6272,
         n6273, n6274, n6275, n6276, n6277, n6278, n6279, n6280, n6281, n6282,
         n6283, n6284, n6285, n6286, n6287, n6288, n6289, n6290, n6291, n6292,
         n6293, n6294, n6295, n6296, n6297, n6298, n6299, n6300, n6301, n6302,
         n6303, n6304, n6305, n6306, n6307, n6308, n6309, n6310, n6311, n6312,
         n6313, n6314, n6315, n6316, n6317, n6318, n6319, n6320, n6321, n6322,
         n6323, n6324, n6325, n6326, n6327, n6328, n6329, n6330, n6331, n6332,
         n6333, n6334, n6335, n6336, n6337, n6338, n6339, n6340, n6341, n6342,
         n6343, n6344, n6345, n6346, n6347, n6348, n6349, n6350, n6351, n6352,
         n6353, n6354, n6355, n6356, n6357, n6358, n6359, n6360, n6361, n6362,
         n6363, n6364, n6365, n6366, n6367, n6368, n6369, n6370, n6371, n6372,
         n6373, n6374, n6375, n6376, n6377, n6378, n6379, n6380, n6381, n6382,
         n6383, n6384, n6385, n6386, n6387, n6388, n6389, n6390, n6391, n6392,
         n6393, n6394, n6395, n6396, n6397, n6398, n6399, n6400, n6401, n6402,
         n6403, n6404, n6405, n6406, n6407, n6408, n6409, n6410, n6411, n6412,
         n6413, n6414, n6415, n6416, n6417, n6418, n6419, n6420, n6421, n6422,
         n6423, n6424, n6425, n6426, n6427, n6428, n6429, n6430, n6431, n6432,
         n6433, n6434, n6435, n6436, n6437, n6438, n6439, n6440, n6441, n6442,
         n6443, n6444, n6445, n6446, n6447, n6448, n6449, n6450, n6451, n6452,
         n6453, n6454, n6455, n6456, n6457, n6458, n6459, n6460, n6461, n6462,
         n6463, n6464, n6465, n6466, n6467, n6468, n6469, n6470, n6471, n6472,
         n6473, n6474, n6475, n6476, n6477, n6478, n6479, n6480, n6481, n6482,
         n6483, n6484, n6485, n6486, n6487, n6488, n6489, n6490, n6491, n6492,
         n6493, n6494, n6495, n6496, n6497, n6498, n6499, n6500, n6501, n6502,
         n6503, n6504, n6505, n6506, n6507, n6508, n6509, n6510, n6511, n6512,
         n6513, n6514, n6515, n6516, n6517, n6518, n6519, n6520, n6521, n6522,
         n6523, n6524, n6525, n6526, n6527, n6528, n6529, n6530, n6531, n6532,
         n6533, n6534, n6535, n6536, n6537, n6538, n6539, n6540, n6541, n6542,
         n6543, n6544, n6545, n6546, n6547, n6548, n6549, n6550, n6551, n6552,
         n6553, n6554, n6555, n6556, n6557, n6558, n6559, n6560, n6561, n6562,
         n6563, n6564, n6565, n6566, n6567, n6568, n6569, n6570, n6571, n6572,
         n6573, n6574, n6575, n6576, n6577, n6578, n6579, n6580, n6581, n6582,
         n6583, n6584, n6585, n6586, n6587, n6588, n6589, n6590, n6591, n6592,
         n6593, n6594, n6595, n6596, n6597, n6598, n6599, n6600, n6601, n6602,
         n6603, n6604, n6605, n6606, n6607, n6608, n6609, n6610, n6611, n6612,
         n6613, n6614, n6615, n6616, n6617, n6618, n6619, n6620, n6621, n6622,
         n6623, n6624, n6625, n6626, n6627, n6628, n6629, n6630, n6631, n6632,
         n6633, n6634, n6635, n6636, n6637, n6638, n6639, n6640, n6641, n6642,
         n6643, n6644, n6645, n6646, n6647, n6648, n6649, n6650, n6651, n6652,
         n6653, n6654, n6655, n6656, n6657, n6658, n6659, n6660, n6661, n6662,
         n6663, n6664, n6665, n6666, n6667, n6668, n6669, n6670, n6671, n6672,
         n6673, n6674, n6675, n6676, n6677, n6678, n6679, n6680, n6681, n6682,
         n6683, n6684, n6685, n6686, n6687, n6688, n6689, n6690, n6691, n6692,
         n6693, n6694, n6695, n6696, n6697, n6698, n6699, n6700, n6701, n6702,
         n6703, n6704, n6705, n6706, n6707, n6708, n6709, n6710, n6711, n6712,
         n6713, n6714, n6715, n6716, n6717, n6718, n6719, n6720, n6721, n6722,
         n6723, n6724, n6725, n6726, n6727, n6728, n6729, n6730, n6731, n6732,
         n6733, n6734, n6735, n6736, n6737, n6738, n6739, n6740, n6741, n6742,
         n6743, n6744, n6745, n6746, n6747, n6748, n6749, n6750, n6751, n6752,
         n6753, n6754, n6755, n6756, n6757, n6758, n6759, n6760, n6761, n6762,
         n6763, n6764, n6765, n6766, n6767, n6768, n6769, n6770, n6771, n6772,
         n6773, n6774, n6775, n6776, n6777, n6778, n6779, n6780, n6781, n6782,
         n6783, n6784, n6785, n6786, n6787, n6788, n6789, n6790, n6791, n6792,
         n6793, n6794, n6795, n6796, n6797, n6798, n6799, n6800, n6801, n6802,
         n6803, n6804, n6805, n6806, n6807, n6808, n6809, n6810, n6811, n6812,
         n6813, n6814, n6815, n6816, n6817, n6818, n6819, n6820, n6821, n6822,
         n6823, n6824, n6825, n6826, n6827, n6828, n6829, n6830, n6831, n6832,
         n6833, n6834, n6835, n6836, n6837, n6838, n6839, n6840, n6841, n6842,
         n6843, n6844, n6845, n6846, n6847, n6848, n6849, n6850, n6851, n6852,
         n6853, n6854, n6855, n6856, n6857, n6858, n6859, n6860, n6861, n6862,
         n6863, n6864, n6865, n6866, n6867, n6868, n6869, n6870, n6871, n6872,
         n6873, n6874, n6875, n6876, n6877, n6878, n6879, n6880, n6881, n6882,
         n6883, n6884, n6885, n6886, n6887, n6888, n6889, n6890, n6891, n6892,
         n6893, n6894, n6895, n6896, n6897, n6898, n6899, n6900, n6901, n6902,
         n6903, n6904, n6905, n6906, n6907, n6908, n6909, n6910, n6911, n6912,
         n6913, n6914, n6915, n6916, n6917, n6918, n6919, n6920, n6921, n6922,
         n6923, n6924, n6925, n6926, n6927, n6928, n6929, n6930, n6931, n6932,
         n6933, n6934, n6935, n6936, n6937, n6938, n6939, n6940, n6941, n6942,
         n6943, n6944, n6945, n6946, n6947, n6948, n6949, n6950, n6951, n6952,
         n6953, n6954, n6955, n6956, n6957, n6958, n6959, n6960, n6961, n6962,
         n6963, n6964, n6965, n6966, n6967, n6968, n6969, n6970, n6971, n6972,
         n6973, n6974, n6975, n6976, n6977, n6978, n6979, n6980, n6981, n6982,
         n6983, n6984, n6985, n6986, n6987, n6988, n6989, n6990, n6991, n6992,
         n6993, n6994, n6995, n6996, n6997, n6998, n6999, n7000, n7001, n7002,
         n7003, n7004, n7005, n7006, n7007, n7008, n7009, n7010, n7011, n7012,
         n7013, n7014, n7015, n7016, n7017, n7018, n7019, n7020, n7021, n7022,
         n7023, n7024, n7025, n7026, n7027, n7028, n7029, n7030, n7031, n7032,
         n7033, n7034, n7035, n7036, n7037, n7038, n7039, n7040, n7041, n7042,
         n7043, n7044, n7045, n7046, n7047, n7048, n7049, n7050, n7051, n7052,
         n7053, n7054, n7055, n7056, n7057, n7058, n7059, n7060, n7061, n7062,
         n7063, n7064, n7065, n7066, n7067, n7068, n7069, n7070, n7071, n7072,
         n7073, n7074, n7075, n7076, n7077, n7078, n7079, n7080, n7081, n7082,
         n7083, n7084, n7085, n7086, n7087, n7088, n7089, n7090, n7091, n7092,
         n7093, n7094, n7095, n7096, n7097, n7098, n7099, n7100, n7101, n7102,
         n7103, n7104, n7105, n7106, n7107, n7108, n7109, n7110, n7111, n7112,
         n7113, n7114, n7115, n7116, n7117, n7118, n7119, n7120, n7121, n7122,
         n7123, n7124, n7125, n7126, n7127, n7128, n7129, n7130, n7131, n7132,
         n7133, n7134, n7135, n7136, n7137, n7138, n7139, n7140, n7141, n7142,
         n7143, n7144, n7145, n7146, n7147, n7148, n7149, n7150, n7151, n7152,
         n7153, n7154, n7155, n7156, n7157, n7158, n7159, n7160, n7161, n7162,
         n7163, n7164, n7165, n7166, n7167, n7168, n7169, n7170, n7171, n7172,
         n7173, n7174, n7175, n7176, n7177, n7178, n7179, n7180, n7181, n7182,
         n7183, n7184, n7185, n7186, n7187, n7188, n7189, n7190, n7191, n7192,
         n7193, n7194, n7195, n7196, n7197, n7198, n7199, n7200, n7201, n7202,
         n7203, n7204, n7205, n7206, n7207, n7208, n7209, n7210, n7211, n7212,
         n7213, n7214, n7215, n7216, n7217, n7218, n7219, n7220, n7221, n7222,
         n7223, n7224, n7225, n7226, n7227, n7228, n7229, n7230, n7231, n7232,
         n7233, n7234, n7235, n7236, n7237, n7238, n7239, n7240, n7241, n7242,
         n7243, n7244, n7245, n7246, n7247, n7248, n7249, n7250, n7251, n7252,
         n7253, n7254, n7255, n7256, n7257, n7258, n7259, n7260, n7261, n7262,
         n7263, n7264, n7265, n7266, n7267, n7268, n7269, n7270, n7271, n7272,
         n7273, n7274, n7275, n7276, n7277, n7278, n7279, n7280, n7281, n7282,
         n7283, n7284, n7285, n7286, n7287, n7288, n7289, n7290, n7291, n7292,
         n7293, n7294, n7295, n7296, n7297, n7298, n7299, n7300, n7301, n7302,
         n7303, n7304, n7305, n7306, n7307, n7308, n7309, n7310, n7311, n7312,
         n7313, n7314, n7315, n7316, n7317, n7318, n7319, n7320, n7321, n7322,
         n7323, n7324, n7325, n7326, n7327, n7328, n7329, n7330, n7331, n7332,
         n7333, n7334, n7335, n7336, n7337, n7338, n7339, n7340, n7341, n7342,
         n7343, n7344, n7345, n7346, n7347, n7348, n7349, n7350, n7351, n7352,
         n7353, n7354, n7355, n7356, n7357, n7358, n7359, n7360, n7361, n7362,
         n7363, n7364, n7365, n7366, n7367, n7368, n7369, n7370, n7371, n7372,
         n7373, n7374, n7375, n7376, n7377, n7378, n7379, n7380, n7381, n7382,
         n7383, n7384, n7385, n7386, n7387, n7388, n7389, n7390, n7391, n7392,
         n7393, n7394, n7395, n7396, n7397, n7398, n7399, n7400, n7401, n7402,
         n7403, n7404, n7405, n7406, n7407, n7408, n7409, n7410, n7411, n7412,
         n7413, n7414, n7415, n7416, n7417, n7418, n7419, n7420, n7421, n7422,
         n7423, n7424, n7425, n7426, n7427, n7428, n7429, n7430, n7431, n7432,
         n7433, n7434, n7435, n7436, n7437, n7438, n7439, n7440, n7441, n7442,
         n7443, n7444, n7445, n7446, n7447, n7448, n7449, n7450, n7451, n7452,
         n7453, n7454, n7455, n7456, n7457, n7458, n7459, n7460, n7461, n7462,
         n7463, n7464, n7465, n7466, n7467, n7468, n7469, n7470, n7471, n7472,
         n7473, n7474, n7475, n7476, n7477, n7478, n7479, n7480, n7481, n7482,
         n7483, n7484, n7485, n7486, n7487, n7488, n7489, n7490, n7491, n7492,
         n7493, n7494, n7495, n7496, n7497, n7498, n7499, n7500, n7501, n7502,
         n7503, n7504, n7505, n7506, n7507, n7508, n7509, n7510, n7511, n7512,
         n7513, n7514, n7515, n7516, n7517, n7518, n7519, n7520, n7521, n7522,
         n7523, n7524, n7525, n7526, n7527, n7528, n7529, n7530, n7531, n7532,
         n7533, n7534, n7535, n7536, n7537, n7538, n7539, n7540, n7541, n7542,
         n7543, n7544, n7545, n7546, n7547, n7548, n7549, n7550, n7551, n7552,
         n7553, n7554, n7555, n7556, n7557, n7558, n7559, n7560, n7561, n7562,
         n7563, n7564, n7565, n7566, n7567, n7568, n7569, n7570, n7571, n7572,
         n7573, n7574, n7575, n7576, n7577, n7578, n7579, n7580, n7581, n7582,
         n7583, n7584, n7585, n7586, n7587, n7588, n7589, n7590, n7591, n7592,
         n7593, n7594, n7595, n7596, n7597, n7598, n7599, n7600, n7601, n7602,
         n7603, n7604, n7605, n7606, n7607, n7608, n7609, n7610, n7611, n7612,
         n7613, n7614, n7615, n7616, n7617, n7618, n7619, n7620, n7621, n7622,
         n7623, n7624, n7625, n7626, n7627, n7628, n7629, n7630, n7631, n7632,
         n7633, n7634, n7635, n7636, n7637, n7638, n7639, n7640, n7641, n7642,
         n7643, n7644, n7645, n7646, n7647, n7648, n7649, n7650, n7651, n7652,
         n7653, n7654, n7655, n7656, n7657, n7658, n7659, n7660, n7661, n7662,
         n7663, n7664, n7665, n7666, n7667, n7668, n7669, n7670, n7671, n7672,
         n7673, n7674, n7675, n7676, n7677, n7678, n7679, n7680, n7681, n7682,
         n7683, n7684, n7685, n7686, n7687, n7688, n7689, n7690, n7691, n7692,
         n7693, n7694, n7695, n7696, n7697, n7698, n7699, n7700, n7701, n7702,
         n7703, n7704, n7705, n7706, n7707, n7708, n7709, n7710, n7711, n7712,
         n7713, n7714, n7715, n7716, n7717, n7718, n7719, n7720, n7721, n7722,
         n7723, n7724, n7725, n7726, n7727, n7728, n7729, n7730, n7731, n7732,
         n7733, n7734, n7735, n7736, n7737, n7738, n7739, n7740, n7741, n7742,
         n7743, n7744, n7745, n7746, n7747, n7748, n7749, n7750, n7751, n7752,
         n7753, n7754, n7755, n7756, n7757, n7758, n7759, n7760, n7761, n7762,
         n7763, n7764, n7765, n7766, n7767, n7768, n7769, n7770, n7771, n7772,
         n7773, n7774, n7775, n7776, n7777, n7778, n7779, n7780, n7781, n7782,
         n7783, n7784, n7785, n7786, n7787, n7788, n7789, n7790, n7791, n7792,
         n7793, n7794, n7795, n7796, n7797, n7798, n7799, n7800, n7801, n7802,
         n7803, n7804, n7805, n7806, n7807, n7808, n7809, n7810, n7811, n7812,
         n7813, n7814, n7815, n7816, n7817, n7818, n7819, n7820, n7821, n7822,
         n7823, n7824, n7825, n7826, n7827, n7828, n7829, n7830, n7831, n7832,
         n7833, n7834, n7835, n7836, n7837, n7838, n7839, n7840, n7841, n7842,
         n7843, n7844, n7845, n7846, n7847, n7848, n7849, n7850, n7851, n7852,
         n7853, n7854, n7855, n7856, n7857, n7858, n7859, n7860, n7861, n7862,
         n7863, n7864, n7865, n7866, n7867, n7868, n7869, n7870, n7871, n7872,
         n7873, n7874, n7875, n7876, n7877, n7878, n7879, n7880, n7881, n7882,
         n7883, n7884, n7885, n7886, n7887, n7888, n7889, n7890, n7891, n7892,
         n7893, n7894, n7895, n7896, n7897, n7898, n7899, n7900, n7901, n7902,
         n7903, n7904, n7905, n7906, n7907, n7908, n7909, n7910, n7911, n7912,
         n7913, n7914, n7915, n7916, n7917, n7918, n7919, n7920, n7921, n7922,
         n7923, n7924, n7925, n7926, n7927, n7928, n7929, n7930, n7931, n7932,
         n7933, n7934, n7935, n7936, n7937, n7938, n7939, n7940, n7941, n7942,
         n7943, n7944, n7945, n7946, n7947, n7948, n7949, n7950, n7951, n7952,
         n7953, n7954, n7955, n7956, n7957, n7958, n7959, n7960, n7961, n7962,
         n7963, n7964, n7965, n7966, n7967, n7968, n7969, n7970, n7971, n7972,
         n7973, n7974, n7975, n7976, n7977, n7978, n7979, n7980, n7981, n7982,
         n7983, n7984, n7985, n7986, n7987, n7988, n7989, n7990, n7991, n7992,
         n7993, n7994, n7995, n7996, n7997, n7998, n7999, n8000, n8001, n8002,
         n8003, n8004, n8005, n8006, n8007, n8008, n8009, n8010, n8011, n8012,
         n8013, n8014, n8015, n8016, n8017, n8018, n8019, n8020, n8021, n8022,
         n8023, n8024, n8025, n8026, n8027, n8028, n8029, n8030, n8031, n8032,
         n8033, n8034, n8035, n8036, n8037, n8038, n8039, n8040, n8041, n8042,
         n8043, n8044, n8045, n8046, n8047, n8048, n8049, n8050, n8051, n8052,
         n8053, n8054, n8055, n8056, n8057, n8058, n8059, n8060, n8061, n8062,
         n8063, n8064, n8065, n8066, n8067, n8068, n8069, n8070, n8071, n8072,
         n8073, n8074, n8075, n8076, n8077, n8078, n8079, n8080, n8081, n8082,
         n8083, n8084, n8085, n8086, n8087, n8088, n8089, n8090, n8091, n8092,
         n8093, n8094, n8095, n8096, n8097, n8098, n8099, n8100, n8101, n8102,
         n8103, n8104, n8105, n8106, n8107, n8108, n8109, n8110, n8111, n8112,
         n8113, n8114, n8115, n8116, n8117, n8118, n8119, n8120, n8121, n8122,
         n8123, n8124, n8125, n8126, n8127, n8128, n8129, n8130, n8131, n8132,
         n8133, n8134, n8135, n8136, n8137, n8138, n8139, n8140, n8141, n8142,
         n8143, n8144, n8145, n8146, n8147, n8148, n8149, n8150, n8151, n8152,
         n8153, n8154, n8155, n8156, n8157, n8158, n8159, n8160, n8161, n8162,
         n8163, n8164, n8165, n8166, n8167, n8168, n8169, n8170, n8171, n8172,
         n8173, n8174, n8175, n8176, n8177, n8178, n8179, n8180, n8181, n8182,
         n8183, n8184, n8185, n8186, n8187, n8188, n8189, n8190, n8191, n8192,
         n8193, n8194, n8195, n8196, n8197, n8198, n8199, n8200, n8201, n8202,
         n8203, n8204, n8205, n8206, n8207, n8208, n8209, n8210, n8211, n8212,
         n8213, n8214, n8215, n8216, n8217, n8218, n8219, n8220, n8221, n8222,
         n8223, n8224, n8225, n8226, n8227, n8228, n8229, n8230, n8231, n8232,
         n8233, n8234, n8235, n8236, n8237, n8238, n8239, n8240, n8241, n8242,
         n8243, n8244, n8245, n8246, n8247, n8248, n8249, n8250, n8251, n8252,
         n8253, n8254, n8255, n8256, n8257, n8258, n8259, n8260, n8261, n8262,
         n8263, n8264, n8265, n8266, n8267, n8268, n8269, n8270, n8271, n8272,
         n8273, n8274, n8275, n8276, n8277, n8278, n8279, n8280, n8281, n8282,
         n8283, n8284, n8285, n8286, n8287, n8288, n8289, n8290, n8291, n8292,
         n8293, n8294, n8295, n8296, n8297, n8298, n8299, n8300, n8301, n8302,
         n8303, n8304, n8305, n8306, n8307, n8308, n8309, n8310, n8311, n8312,
         n8313, n8314, n8315, n8316, n8317, n8318, n8319, n8320, n8321, n8322,
         n8323, n8324, n8325, n8326, n8327, n8328, n8329, n8330, n8331, n8332,
         n8333, n8334, n8335, n8336, n8337, n8338, n8339, n8340, n8341, n8342,
         n8343, n8344, n8345, n8346, n8347, n8348, n8349, n8350, n8351, n8352,
         n8353, n8354, n8355, n8356, n8357, n8358, n8359, n8360, n8361, n8362,
         n8363, n8364, n8365, n8366, n8367, n8368, n8369, n8370, n8371, n8372,
         n8373, n8374, n8375, n8376, n8377, n8378, n8379, n8380, n8381, n8382,
         n8383, n8384, n8385, n8386, n8387, n8388, n8389, n8390, n8391, n8392,
         n8393, n8394, n8395, n8396, n8397, n8398, n8399, n8400, n8401, n8402,
         n8403, n8404, n8405, n8406, n8407, n8408, n8409, n8410, n8411, n8412,
         n8413, n8414, n8415, n8416, n8417, n8418, n8419, n8420, n8421, n8422,
         n8423, n8424, n8425, n8426, n8427, n8428, n8429, n8430, n8431, n8432,
         n8433, n8434, n8435, n8436, n8437, n8438, n8439, n8440, n8441, n8442,
         n8443, n8444, n8445, n8446, n8447, n8448, n8449, n8450, n8451, n8452,
         n8453, n8454, n8455, n8456, n8457, n8458, n8459, n8460, n8461, n8462,
         n8463, n8464, n8465, n8466, n8467, n8468, n8469, n8470, n8471, n8472,
         n8473, n8474, n8475, n8476, n8477, n8478, n8479, n8480, n8481, n8482,
         n8483, n8484, n8485, n8486, n8487, n8488, n8489, n8490, n8491, n8492,
         n8493, n8494, n8495, n8496, n8497, n8498, n8499, n8500, n8501, n8502,
         n8503, n8504, n8505, n8506, n8507, n8508, n8509, n8510, n8511, n8512,
         n8513, n8514, n8515, n8516, n8517, n8518, n8519, n8520, n8521, n8522,
         n8523, n8524, n8525, n8526, n8527, n8528, n8529, n8530, n8531, n8532,
         n8533, n8534, n8535, n8536, n8537, n8538, n8539, n8540, n8541, n8542,
         n8543, n8544, n8545, n8546, n8547, n8548, n8549, n8550, n8551, n8552,
         n8553, n8554, n8555, n8556, n8557, n8558, n8559, n8560, n8561, n8562,
         n8563, n8564, n8565, n8566, n8567, n8568, n8569, n8570, n8571, n8572,
         n8573, n8574, n8575, n8576, n8577, n8578, n8579, n8580;
  wire   [63:32] swire;
  wire   [127:64] sreg;

  DFF \sreg_reg[64]  ( .D(swire[32]), .CLK(clk), .RST(rst), .Q(sreg[64]) );
  DFF \sreg_reg[65]  ( .D(swire[33]), .CLK(clk), .RST(rst), .Q(sreg[65]) );
  DFF \sreg_reg[66]  ( .D(swire[34]), .CLK(clk), .RST(rst), .Q(sreg[66]) );
  DFF \sreg_reg[67]  ( .D(swire[35]), .CLK(clk), .RST(rst), .Q(sreg[67]) );
  DFF \sreg_reg[68]  ( .D(swire[36]), .CLK(clk), .RST(rst), .Q(sreg[68]) );
  DFF \sreg_reg[69]  ( .D(swire[37]), .CLK(clk), .RST(rst), .Q(sreg[69]) );
  DFF \sreg_reg[70]  ( .D(swire[38]), .CLK(clk), .RST(rst), .Q(sreg[70]) );
  DFF \sreg_reg[71]  ( .D(swire[39]), .CLK(clk), .RST(rst), .Q(sreg[71]) );
  DFF \sreg_reg[72]  ( .D(swire[40]), .CLK(clk), .RST(rst), .Q(sreg[72]) );
  DFF \sreg_reg[73]  ( .D(swire[41]), .CLK(clk), .RST(rst), .Q(sreg[73]) );
  DFF \sreg_reg[74]  ( .D(swire[42]), .CLK(clk), .RST(rst), .Q(sreg[74]) );
  DFF \sreg_reg[75]  ( .D(swire[43]), .CLK(clk), .RST(rst), .Q(sreg[75]) );
  DFF \sreg_reg[76]  ( .D(swire[44]), .CLK(clk), .RST(rst), .Q(sreg[76]) );
  DFF \sreg_reg[77]  ( .D(swire[45]), .CLK(clk), .RST(rst), .Q(sreg[77]) );
  DFF \sreg_reg[78]  ( .D(swire[46]), .CLK(clk), .RST(rst), .Q(sreg[78]) );
  DFF \sreg_reg[79]  ( .D(swire[47]), .CLK(clk), .RST(rst), .Q(sreg[79]) );
  DFF \sreg_reg[80]  ( .D(swire[48]), .CLK(clk), .RST(rst), .Q(sreg[80]) );
  DFF \sreg_reg[81]  ( .D(swire[49]), .CLK(clk), .RST(rst), .Q(sreg[81]) );
  DFF \sreg_reg[82]  ( .D(swire[50]), .CLK(clk), .RST(rst), .Q(sreg[82]) );
  DFF \sreg_reg[83]  ( .D(swire[51]), .CLK(clk), .RST(rst), .Q(sreg[83]) );
  DFF \sreg_reg[84]  ( .D(swire[52]), .CLK(clk), .RST(rst), .Q(sreg[84]) );
  DFF \sreg_reg[85]  ( .D(swire[53]), .CLK(clk), .RST(rst), .Q(sreg[85]) );
  DFF \sreg_reg[86]  ( .D(swire[54]), .CLK(clk), .RST(rst), .Q(sreg[86]) );
  DFF \sreg_reg[87]  ( .D(swire[55]), .CLK(clk), .RST(rst), .Q(sreg[87]) );
  DFF \sreg_reg[88]  ( .D(swire[56]), .CLK(clk), .RST(rst), .Q(sreg[88]) );
  DFF \sreg_reg[89]  ( .D(swire[57]), .CLK(clk), .RST(rst), .Q(sreg[89]) );
  DFF \sreg_reg[90]  ( .D(swire[58]), .CLK(clk), .RST(rst), .Q(sreg[90]) );
  DFF \sreg_reg[91]  ( .D(swire[59]), .CLK(clk), .RST(rst), .Q(sreg[91]) );
  DFF \sreg_reg[92]  ( .D(swire[60]), .CLK(clk), .RST(rst), .Q(sreg[92]) );
  DFF \sreg_reg[93]  ( .D(swire[61]), .CLK(clk), .RST(rst), .Q(sreg[93]) );
  DFF \sreg_reg[94]  ( .D(swire[62]), .CLK(clk), .RST(rst), .Q(sreg[94]) );
  DFF \sreg_reg[95]  ( .D(swire[63]), .CLK(clk), .RST(rst), .Q(sreg[95]) );
  DFF \sreg_reg[63]  ( .D(c[63]), .CLK(clk), .RST(rst), .Q(c[31]) );
  DFF \sreg_reg[62]  ( .D(c[62]), .CLK(clk), .RST(rst), .Q(c[30]) );
  DFF \sreg_reg[61]  ( .D(c[61]), .CLK(clk), .RST(rst), .Q(c[29]) );
  DFF \sreg_reg[60]  ( .D(c[60]), .CLK(clk), .RST(rst), .Q(c[28]) );
  DFF \sreg_reg[59]  ( .D(c[59]), .CLK(clk), .RST(rst), .Q(c[27]) );
  DFF \sreg_reg[58]  ( .D(c[58]), .CLK(clk), .RST(rst), .Q(c[26]) );
  DFF \sreg_reg[57]  ( .D(c[57]), .CLK(clk), .RST(rst), .Q(c[25]) );
  DFF \sreg_reg[56]  ( .D(c[56]), .CLK(clk), .RST(rst), .Q(c[24]) );
  DFF \sreg_reg[55]  ( .D(c[55]), .CLK(clk), .RST(rst), .Q(c[23]) );
  DFF \sreg_reg[54]  ( .D(c[54]), .CLK(clk), .RST(rst), .Q(c[22]) );
  DFF \sreg_reg[53]  ( .D(c[53]), .CLK(clk), .RST(rst), .Q(c[21]) );
  DFF \sreg_reg[52]  ( .D(c[52]), .CLK(clk), .RST(rst), .Q(c[20]) );
  DFF \sreg_reg[51]  ( .D(c[51]), .CLK(clk), .RST(rst), .Q(c[19]) );
  DFF \sreg_reg[50]  ( .D(c[50]), .CLK(clk), .RST(rst), .Q(c[18]) );
  DFF \sreg_reg[49]  ( .D(c[49]), .CLK(clk), .RST(rst), .Q(c[17]) );
  DFF \sreg_reg[48]  ( .D(c[48]), .CLK(clk), .RST(rst), .Q(c[16]) );
  DFF \sreg_reg[47]  ( .D(c[47]), .CLK(clk), .RST(rst), .Q(c[15]) );
  DFF \sreg_reg[46]  ( .D(c[46]), .CLK(clk), .RST(rst), .Q(c[14]) );
  DFF \sreg_reg[45]  ( .D(c[45]), .CLK(clk), .RST(rst), .Q(c[13]) );
  DFF \sreg_reg[44]  ( .D(c[44]), .CLK(clk), .RST(rst), .Q(c[12]) );
  DFF \sreg_reg[43]  ( .D(c[43]), .CLK(clk), .RST(rst), .Q(c[11]) );
  DFF \sreg_reg[42]  ( .D(c[42]), .CLK(clk), .RST(rst), .Q(c[10]) );
  DFF \sreg_reg[41]  ( .D(c[41]), .CLK(clk), .RST(rst), .Q(c[9]) );
  DFF \sreg_reg[40]  ( .D(c[40]), .CLK(clk), .RST(rst), .Q(c[8]) );
  DFF \sreg_reg[39]  ( .D(c[39]), .CLK(clk), .RST(rst), .Q(c[7]) );
  DFF \sreg_reg[38]  ( .D(c[38]), .CLK(clk), .RST(rst), .Q(c[6]) );
  DFF \sreg_reg[37]  ( .D(c[37]), .CLK(clk), .RST(rst), .Q(c[5]) );
  DFF \sreg_reg[36]  ( .D(c[36]), .CLK(clk), .RST(rst), .Q(c[4]) );
  DFF \sreg_reg[35]  ( .D(c[35]), .CLK(clk), .RST(rst), .Q(c[3]) );
  DFF \sreg_reg[34]  ( .D(c[34]), .CLK(clk), .RST(rst), .Q(c[2]) );
  DFF \sreg_reg[33]  ( .D(c[33]), .CLK(clk), .RST(rst), .Q(c[1]) );
  DFF \sreg_reg[32]  ( .D(c[32]), .CLK(clk), .RST(rst), .Q(c[0]) );
  XOR U35 ( .A(n1566), .B(n1724), .Z(n1570) );
  XOR U36 ( .A(n1394), .B(n1540), .Z(n1398) );
  XOR U37 ( .A(n1596), .B(n1717), .Z(n1600) );
  XOR U38 ( .A(n1616), .B(n1712), .Z(n1620) );
  XOR U39 ( .A(n1071), .B(n1168), .Z(n1075) );
  XOR U40 ( .A(n687), .B(n809), .Z(n691) );
  XOR U41 ( .A(n1268), .B(n1346), .Z(n1272) );
  XOR U42 ( .A(n531), .B(n622), .Z(n535) );
  XOR U43 ( .A(n737), .B(n798), .Z(n741) );
  XOR U44 ( .A(n6241), .B(n6400), .Z(n6245) );
  XOR U45 ( .A(n5903), .B(n6062), .Z(n5907) );
  XOR U46 ( .A(n5539), .B(n5698), .Z(n5543) );
  XOR U47 ( .A(n1929), .B(n2085), .Z(n1933) );
  XOR U48 ( .A(n2290), .B(n2446), .Z(n2294) );
  XOR U49 ( .A(n2651), .B(n2807), .Z(n2655) );
  XOR U50 ( .A(n3012), .B(n3168), .Z(n3016) );
  XOR U51 ( .A(n3373), .B(n3529), .Z(n3377) );
  XOR U52 ( .A(n3734), .B(n3890), .Z(n3738) );
  XOR U53 ( .A(n4095), .B(n4251), .Z(n4099) );
  XOR U54 ( .A(n4456), .B(n4612), .Z(n4460) );
  XOR U55 ( .A(n4817), .B(n4973), .Z(n4821) );
  XOR U56 ( .A(n5178), .B(n5334), .Z(n5182) );
  XOR U57 ( .A(n1379), .B(n1543), .Z(n1383) );
  XOR U58 ( .A(n6570), .B(n6711), .Z(n6574) );
  XOR U59 ( .A(n6256), .B(n6397), .Z(n6260) );
  XOR U60 ( .A(n5918), .B(n6059), .Z(n5922) );
  XOR U61 ( .A(n5554), .B(n5695), .Z(n5558) );
  XOR U62 ( .A(n1944), .B(n2082), .Z(n1948) );
  XOR U63 ( .A(n2305), .B(n2443), .Z(n2309) );
  XOR U64 ( .A(n2666), .B(n2804), .Z(n2670) );
  XOR U65 ( .A(n3027), .B(n3165), .Z(n3031) );
  XOR U66 ( .A(n3388), .B(n3526), .Z(n3392) );
  XOR U67 ( .A(n3749), .B(n3887), .Z(n3753) );
  XOR U68 ( .A(n4110), .B(n4248), .Z(n4114) );
  XOR U69 ( .A(n4471), .B(n4609), .Z(n4475) );
  XOR U70 ( .A(n4832), .B(n4970), .Z(n4836) );
  XOR U71 ( .A(n5193), .B(n5331), .Z(n5197) );
  XOR U72 ( .A(n1208), .B(n1359), .Z(n1212) );
  XOR U73 ( .A(n1591), .B(n1718), .Z(n1595) );
  XOR U74 ( .A(n7141), .B(n7264), .Z(n7145) );
  XOR U75 ( .A(n6875), .B(n6998), .Z(n6879) );
  XOR U76 ( .A(n6585), .B(n6708), .Z(n6589) );
  XOR U77 ( .A(n6271), .B(n6394), .Z(n6275) );
  XOR U78 ( .A(n5933), .B(n6056), .Z(n5937) );
  XOR U79 ( .A(n5569), .B(n5692), .Z(n5573) );
  XOR U80 ( .A(n1959), .B(n2079), .Z(n1963) );
  XOR U81 ( .A(n2320), .B(n2440), .Z(n2324) );
  XOR U82 ( .A(n2681), .B(n2801), .Z(n2685) );
  XOR U83 ( .A(n3042), .B(n3162), .Z(n3046) );
  XOR U84 ( .A(n3403), .B(n3523), .Z(n3407) );
  XOR U85 ( .A(n3764), .B(n3884), .Z(n3768) );
  XOR U86 ( .A(n4125), .B(n4245), .Z(n4129) );
  XOR U87 ( .A(n4486), .B(n4606), .Z(n4490) );
  XOR U88 ( .A(n4847), .B(n4967), .Z(n4851) );
  XOR U89 ( .A(n5208), .B(n5328), .Z(n5212) );
  XOR U90 ( .A(n1223), .B(n1356), .Z(n1227) );
  XOR U91 ( .A(n839), .B(n997), .Z(n843) );
  XOR U92 ( .A(n7398), .B(n7503), .Z(n7402) );
  XOR U93 ( .A(n7156), .B(n7261), .Z(n7160) );
  XOR U94 ( .A(n6890), .B(n6995), .Z(n6894) );
  XOR U95 ( .A(n6600), .B(n6705), .Z(n6604) );
  XOR U96 ( .A(n6286), .B(n6391), .Z(n6290) );
  XOR U97 ( .A(n5948), .B(n6053), .Z(n5952) );
  XOR U98 ( .A(n5584), .B(n5689), .Z(n5588) );
  XOR U99 ( .A(n1248), .B(n1351), .Z(n1252) );
  XOR U100 ( .A(n1974), .B(n2076), .Z(n1978) );
  XOR U101 ( .A(n2335), .B(n2437), .Z(n2339) );
  XOR U102 ( .A(n2696), .B(n2798), .Z(n2700) );
  XOR U103 ( .A(n3057), .B(n3159), .Z(n3061) );
  XOR U104 ( .A(n3418), .B(n3520), .Z(n3422) );
  XOR U105 ( .A(n3779), .B(n3881), .Z(n3783) );
  XOR U106 ( .A(n4140), .B(n4242), .Z(n4144) );
  XOR U107 ( .A(n4501), .B(n4603), .Z(n4505) );
  XOR U108 ( .A(n4862), .B(n4964), .Z(n4866) );
  XOR U109 ( .A(n5223), .B(n5325), .Z(n5227) );
  XOR U110 ( .A(n1424), .B(n1533), .Z(n1428) );
  XOR U111 ( .A(n1046), .B(n1174), .Z(n1050) );
  XOR U112 ( .A(n662), .B(n814), .Z(n666) );
  XOR U113 ( .A(n7825), .B(n7912), .Z(n7829) );
  XOR U114 ( .A(n7631), .B(n7718), .Z(n7635) );
  XOR U115 ( .A(n7413), .B(n7500), .Z(n7417) );
  XOR U116 ( .A(n7171), .B(n7258), .Z(n7175) );
  XOR U117 ( .A(n6905), .B(n6992), .Z(n6909) );
  XOR U118 ( .A(n6615), .B(n6702), .Z(n6619) );
  XOR U119 ( .A(n6301), .B(n6388), .Z(n6305) );
  XOR U120 ( .A(n5963), .B(n6050), .Z(n5967) );
  XOR U121 ( .A(n5599), .B(n5686), .Z(n5603) );
  XOR U122 ( .A(n1076), .B(n1167), .Z(n1080) );
  XOR U123 ( .A(n899), .B(n985), .Z(n903) );
  XOR U124 ( .A(n1626), .B(n1710), .Z(n1630) );
  XOR U125 ( .A(n1989), .B(n2073), .Z(n1993) );
  XOR U126 ( .A(n2350), .B(n2434), .Z(n2354) );
  XOR U127 ( .A(n2711), .B(n2795), .Z(n2715) );
  XOR U128 ( .A(n3072), .B(n3156), .Z(n3076) );
  XOR U129 ( .A(n3433), .B(n3517), .Z(n3437) );
  XOR U130 ( .A(n3794), .B(n3878), .Z(n3798) );
  XOR U131 ( .A(n4155), .B(n4239), .Z(n4159) );
  XOR U132 ( .A(n4516), .B(n4600), .Z(n4520) );
  XOR U133 ( .A(n4877), .B(n4961), .Z(n4881) );
  XOR U134 ( .A(n5238), .B(n5322), .Z(n5242) );
  XOR U135 ( .A(n697), .B(n807), .Z(n701) );
  XOR U136 ( .A(n486), .B(n631), .Z(n490) );
  XOR U137 ( .A(n8010), .B(n8079), .Z(n8014) );
  XOR U138 ( .A(n7840), .B(n7909), .Z(n7844) );
  XOR U139 ( .A(n7646), .B(n7715), .Z(n7650) );
  XOR U140 ( .A(n7428), .B(n7497), .Z(n7432) );
  XOR U141 ( .A(n7186), .B(n7255), .Z(n7190) );
  XOR U142 ( .A(n6920), .B(n6989), .Z(n6924) );
  XOR U143 ( .A(n6630), .B(n6699), .Z(n6634) );
  XOR U144 ( .A(n6316), .B(n6385), .Z(n6320) );
  XOR U145 ( .A(n5978), .B(n6047), .Z(n5982) );
  XOR U146 ( .A(n5614), .B(n5683), .Z(n5618) );
  XOR U147 ( .A(n536), .B(n621), .Z(n540) );
  XOR U148 ( .A(n1278), .B(n1344), .Z(n1282) );
  XOR U149 ( .A(n1641), .B(n1707), .Z(n1645) );
  XOR U150 ( .A(n2004), .B(n2070), .Z(n2008) );
  XOR U151 ( .A(n2365), .B(n2431), .Z(n2369) );
  XOR U152 ( .A(n2726), .B(n2792), .Z(n2730) );
  XOR U153 ( .A(n3087), .B(n3153), .Z(n3091) );
  XOR U154 ( .A(n3448), .B(n3514), .Z(n3452) );
  XOR U155 ( .A(n3809), .B(n3875), .Z(n3813) );
  XOR U156 ( .A(n4170), .B(n4236), .Z(n4174) );
  XOR U157 ( .A(n4531), .B(n4597), .Z(n4535) );
  XOR U158 ( .A(n4892), .B(n4958), .Z(n4896) );
  XOR U159 ( .A(n5253), .B(n5319), .Z(n5257) );
  XOR U160 ( .A(n732), .B(n799), .Z(n736) );
  XOR U161 ( .A(n8293), .B(n8344), .Z(n8297) );
  XOR U162 ( .A(n8171), .B(n8222), .Z(n8175) );
  XOR U163 ( .A(n8025), .B(n8076), .Z(n8029) );
  XOR U164 ( .A(n7855), .B(n7906), .Z(n7859) );
  XOR U165 ( .A(n7661), .B(n7712), .Z(n7665) );
  XOR U166 ( .A(n7443), .B(n7494), .Z(n7447) );
  XOR U167 ( .A(n7201), .B(n7252), .Z(n7205) );
  XOR U168 ( .A(n6935), .B(n6986), .Z(n6939) );
  XOR U169 ( .A(n6645), .B(n6696), .Z(n6649) );
  XOR U170 ( .A(n6331), .B(n6382), .Z(n6335) );
  XOR U171 ( .A(n5993), .B(n6044), .Z(n5997) );
  XOR U172 ( .A(n5629), .B(n5680), .Z(n5633) );
  XOR U173 ( .A(n566), .B(n614), .Z(n570) );
  XOR U174 ( .A(n929), .B(n977), .Z(n933) );
  XOR U175 ( .A(n1293), .B(n1341), .Z(n1297) );
  XOR U176 ( .A(n1656), .B(n1704), .Z(n1660) );
  XOR U177 ( .A(n2019), .B(n2067), .Z(n2023) );
  XOR U178 ( .A(n2380), .B(n2428), .Z(n2384) );
  XOR U179 ( .A(n2741), .B(n2789), .Z(n2745) );
  XOR U180 ( .A(n3102), .B(n3150), .Z(n3106) );
  XOR U181 ( .A(n3463), .B(n3511), .Z(n3467) );
  XOR U182 ( .A(n3824), .B(n3872), .Z(n3828) );
  XOR U183 ( .A(n4185), .B(n4233), .Z(n4189) );
  XOR U184 ( .A(n4546), .B(n4594), .Z(n4550) );
  XOR U185 ( .A(n4907), .B(n4955), .Z(n4911) );
  XOR U186 ( .A(n5268), .B(n5316), .Z(n5272) );
  XOR U187 ( .A(n8406), .B(n8439), .Z(n8410) );
  XOR U188 ( .A(n8308), .B(n8341), .Z(n8312) );
  XOR U189 ( .A(n8186), .B(n8219), .Z(n8190) );
  XOR U190 ( .A(n8040), .B(n8073), .Z(n8044) );
  XOR U191 ( .A(n7870), .B(n7903), .Z(n7874) );
  XOR U192 ( .A(n7676), .B(n7709), .Z(n7680) );
  XOR U193 ( .A(n7458), .B(n7491), .Z(n7462) );
  XOR U194 ( .A(n7216), .B(n7249), .Z(n7220) );
  XOR U195 ( .A(n6950), .B(n6983), .Z(n6954) );
  XOR U196 ( .A(n6660), .B(n6693), .Z(n6664) );
  XOR U197 ( .A(n6346), .B(n6379), .Z(n6350) );
  XOR U198 ( .A(n6008), .B(n6041), .Z(n6012) );
  XOR U199 ( .A(n5644), .B(n5677), .Z(n5648) );
  XOR U200 ( .A(n581), .B(n611), .Z(n585) );
  XOR U201 ( .A(n944), .B(n974), .Z(n948) );
  XOR U202 ( .A(n1308), .B(n1338), .Z(n1312) );
  XOR U203 ( .A(n1671), .B(n1701), .Z(n1675) );
  XOR U204 ( .A(n2034), .B(n2064), .Z(n2038) );
  XOR U205 ( .A(n2395), .B(n2425), .Z(n2399) );
  XOR U206 ( .A(n2756), .B(n2786), .Z(n2760) );
  XOR U207 ( .A(n3117), .B(n3147), .Z(n3121) );
  XOR U208 ( .A(n3478), .B(n3508), .Z(n3482) );
  XOR U209 ( .A(n3839), .B(n3869), .Z(n3843) );
  XOR U210 ( .A(n4200), .B(n4230), .Z(n4204) );
  XOR U211 ( .A(n4561), .B(n4591), .Z(n4565) );
  XOR U212 ( .A(n4922), .B(n4952), .Z(n4926) );
  XOR U213 ( .A(n5283), .B(n5313), .Z(n5287) );
  XOR U214 ( .A(n6075), .B(n6234), .Z(n6079) );
  XOR U215 ( .A(n5722), .B(n5881), .Z(n5726) );
  XOR U216 ( .A(n1748), .B(n1905), .Z(n1752) );
  XOR U217 ( .A(n2109), .B(n2266), .Z(n2113) );
  XOR U218 ( .A(n2470), .B(n2627), .Z(n2474) );
  XOR U219 ( .A(n2831), .B(n2988), .Z(n2835) );
  XOR U220 ( .A(n3192), .B(n3349), .Z(n3196) );
  XOR U221 ( .A(n3553), .B(n3710), .Z(n3557) );
  XOR U222 ( .A(n3914), .B(n4071), .Z(n3918) );
  XOR U223 ( .A(n4275), .B(n4432), .Z(n4279) );
  XOR U224 ( .A(n4636), .B(n4793), .Z(n4640) );
  XOR U225 ( .A(n4997), .B(n5154), .Z(n5001) );
  XOR U226 ( .A(n5358), .B(n5515), .Z(n5362) );
  XOR U227 ( .A(n1384), .B(n1542), .Z(n1388) );
  XOR U228 ( .A(n6718), .B(n6859), .Z(n6722) );
  XOR U229 ( .A(n6416), .B(n6557), .Z(n6420) );
  XOR U230 ( .A(n6090), .B(n6231), .Z(n6094) );
  XOR U231 ( .A(n5737), .B(n5878), .Z(n5741) );
  XOR U232 ( .A(n1763), .B(n1902), .Z(n1767) );
  XOR U233 ( .A(n2124), .B(n2263), .Z(n2128) );
  XOR U234 ( .A(n2485), .B(n2624), .Z(n2489) );
  XOR U235 ( .A(n2846), .B(n2985), .Z(n2850) );
  XOR U236 ( .A(n3207), .B(n3346), .Z(n3211) );
  XOR U237 ( .A(n3568), .B(n3707), .Z(n3572) );
  XOR U238 ( .A(n3929), .B(n4068), .Z(n3933) );
  XOR U239 ( .A(n4290), .B(n4429), .Z(n4294) );
  XOR U240 ( .A(n4651), .B(n4790), .Z(n4655) );
  XOR U241 ( .A(n5012), .B(n5151), .Z(n5016) );
  XOR U242 ( .A(n5373), .B(n5512), .Z(n5377) );
  XOR U243 ( .A(n7011), .B(n7134), .Z(n7015) );
  XOR U244 ( .A(n6733), .B(n6856), .Z(n6737) );
  XOR U245 ( .A(n6431), .B(n6554), .Z(n6435) );
  XOR U246 ( .A(n6105), .B(n6228), .Z(n6109) );
  XOR U247 ( .A(n5752), .B(n5875), .Z(n5756) );
  XOR U248 ( .A(n1021), .B(n1179), .Z(n1025) );
  XOR U249 ( .A(n1778), .B(n1899), .Z(n1782) );
  XOR U250 ( .A(n2139), .B(n2260), .Z(n2143) );
  XOR U251 ( .A(n2500), .B(n2621), .Z(n2504) );
  XOR U252 ( .A(n2861), .B(n2982), .Z(n2865) );
  XOR U253 ( .A(n3222), .B(n3343), .Z(n3226) );
  XOR U254 ( .A(n3583), .B(n3704), .Z(n3587) );
  XOR U255 ( .A(n3944), .B(n4065), .Z(n3948) );
  XOR U256 ( .A(n4305), .B(n4426), .Z(n4309) );
  XOR U257 ( .A(n4666), .B(n4787), .Z(n4670) );
  XOR U258 ( .A(n5027), .B(n5148), .Z(n5031) );
  XOR U259 ( .A(n5388), .B(n5509), .Z(n5392) );
  XOR U260 ( .A(n7510), .B(n7615), .Z(n7514) );
  XOR U261 ( .A(n7280), .B(n7385), .Z(n7284) );
  XOR U262 ( .A(n7026), .B(n7131), .Z(n7030) );
  XOR U263 ( .A(n6748), .B(n6853), .Z(n6752) );
  XOR U264 ( .A(n6446), .B(n6551), .Z(n6450) );
  XOR U265 ( .A(n6120), .B(n6225), .Z(n6124) );
  XOR U266 ( .A(n5767), .B(n5872), .Z(n5771) );
  XOR U267 ( .A(n1228), .B(n1355), .Z(n1232) );
  XOR U268 ( .A(n844), .B(n996), .Z(n848) );
  XOR U269 ( .A(n1793), .B(n1896), .Z(n1797) );
  XOR U270 ( .A(n2154), .B(n2257), .Z(n2158) );
  XOR U271 ( .A(n2515), .B(n2618), .Z(n2519) );
  XOR U272 ( .A(n2876), .B(n2979), .Z(n2880) );
  XOR U273 ( .A(n3237), .B(n3340), .Z(n3241) );
  XOR U274 ( .A(n3598), .B(n3701), .Z(n3602) );
  XOR U275 ( .A(n3959), .B(n4062), .Z(n3963) );
  XOR U276 ( .A(n4320), .B(n4423), .Z(n4324) );
  XOR U277 ( .A(n4681), .B(n4784), .Z(n4685) );
  XOR U278 ( .A(n5042), .B(n5145), .Z(n5046) );
  XOR U279 ( .A(n5403), .B(n5506), .Z(n5407) );
  XOR U280 ( .A(n874), .B(n990), .Z(n878) );
  XOR U281 ( .A(n1429), .B(n1532), .Z(n1433) );
  XOR U282 ( .A(n7731), .B(n7818), .Z(n7735) );
  XOR U283 ( .A(n7525), .B(n7612), .Z(n7529) );
  XOR U284 ( .A(n7295), .B(n7382), .Z(n7299) );
  XOR U285 ( .A(n7041), .B(n7128), .Z(n7045) );
  XOR U286 ( .A(n6763), .B(n6850), .Z(n6767) );
  XOR U287 ( .A(n6461), .B(n6548), .Z(n6465) );
  XOR U288 ( .A(n6135), .B(n6222), .Z(n6139) );
  XOR U289 ( .A(n5782), .B(n5869), .Z(n5786) );
  XOR U290 ( .A(n859), .B(n993), .Z(n863) );
  XOR U291 ( .A(n476), .B(n633), .Z(n480) );
  XOR U292 ( .A(n1444), .B(n1529), .Z(n1448) );
  XOR U293 ( .A(n1808), .B(n1893), .Z(n1812) );
  XOR U294 ( .A(n2169), .B(n2254), .Z(n2173) );
  XOR U295 ( .A(n2530), .B(n2615), .Z(n2534) );
  XOR U296 ( .A(n2891), .B(n2976), .Z(n2895) );
  XOR U297 ( .A(n3252), .B(n3337), .Z(n3256) );
  XOR U298 ( .A(n3613), .B(n3698), .Z(n3617) );
  XOR U299 ( .A(n3974), .B(n4059), .Z(n3978) );
  XOR U300 ( .A(n4335), .B(n4420), .Z(n4339) );
  XOR U301 ( .A(n4696), .B(n4781), .Z(n4700) );
  XOR U302 ( .A(n5057), .B(n5142), .Z(n5061) );
  XOR U303 ( .A(n5418), .B(n5503), .Z(n5422) );
  XOR U304 ( .A(n1081), .B(n1166), .Z(n1085) );
  XOR U305 ( .A(n316), .B(n448), .Z(n320) );
  XOR U306 ( .A(n526), .B(n623), .Z(n530) );
  XOR U307 ( .A(n511), .B(n626), .Z(n515) );
  XOR U308 ( .A(n8086), .B(n8155), .Z(n8090) );
  XOR U309 ( .A(n7928), .B(n7997), .Z(n7932) );
  XOR U310 ( .A(n7746), .B(n7815), .Z(n7750) );
  XOR U311 ( .A(n7540), .B(n7609), .Z(n7544) );
  XOR U312 ( .A(n7310), .B(n7379), .Z(n7314) );
  XOR U313 ( .A(n7056), .B(n7125), .Z(n7060) );
  XOR U314 ( .A(n6778), .B(n6847), .Z(n6782) );
  XOR U315 ( .A(n6476), .B(n6545), .Z(n6480) );
  XOR U316 ( .A(n6150), .B(n6219), .Z(n6154) );
  XOR U317 ( .A(n5797), .B(n5866), .Z(n5801) );
  XOR U318 ( .A(n491), .B(n630), .Z(n495) );
  XOR U319 ( .A(n1096), .B(n1163), .Z(n1100) );
  XOR U320 ( .A(n1459), .B(n1526), .Z(n1463) );
  XOR U321 ( .A(n1823), .B(n1890), .Z(n1827) );
  XOR U322 ( .A(n2184), .B(n2251), .Z(n2188) );
  XOR U323 ( .A(n2545), .B(n2612), .Z(n2549) );
  XOR U324 ( .A(n2906), .B(n2973), .Z(n2910) );
  XOR U325 ( .A(n3267), .B(n3334), .Z(n3271) );
  XOR U326 ( .A(n3628), .B(n3695), .Z(n3632) );
  XOR U327 ( .A(n3989), .B(n4056), .Z(n3993) );
  XOR U328 ( .A(n4350), .B(n4417), .Z(n4354) );
  XOR U329 ( .A(n4711), .B(n4778), .Z(n4715) );
  XOR U330 ( .A(n5072), .B(n5139), .Z(n5076) );
  XOR U331 ( .A(n5433), .B(n5500), .Z(n5437) );
  XOR U332 ( .A(n541), .B(n620), .Z(n545) );
  XOR U333 ( .A(n8235), .B(n8286), .Z(n8239) );
  XOR U334 ( .A(n8101), .B(n8152), .Z(n8105) );
  XOR U335 ( .A(n7943), .B(n7994), .Z(n7947) );
  XOR U336 ( .A(n7761), .B(n7812), .Z(n7765) );
  XOR U337 ( .A(n7555), .B(n7606), .Z(n7559) );
  XOR U338 ( .A(n7325), .B(n7376), .Z(n7329) );
  XOR U339 ( .A(n7071), .B(n7122), .Z(n7075) );
  XOR U340 ( .A(n6793), .B(n6844), .Z(n6797) );
  XOR U341 ( .A(n6491), .B(n6542), .Z(n6495) );
  XOR U342 ( .A(n6165), .B(n6216), .Z(n6169) );
  XOR U343 ( .A(n5812), .B(n5863), .Z(n5816) );
  XOR U344 ( .A(n386), .B(n434), .Z(n390) );
  XOR U345 ( .A(n747), .B(n796), .Z(n751) );
  XOR U346 ( .A(n1111), .B(n1160), .Z(n1115) );
  XOR U347 ( .A(n1474), .B(n1523), .Z(n1478) );
  XOR U348 ( .A(n1838), .B(n1887), .Z(n1842) );
  XOR U349 ( .A(n2199), .B(n2248), .Z(n2203) );
  XOR U350 ( .A(n2560), .B(n2609), .Z(n2564) );
  XOR U351 ( .A(n2921), .B(n2970), .Z(n2925) );
  XOR U352 ( .A(n3282), .B(n3331), .Z(n3286) );
  XOR U353 ( .A(n3643), .B(n3692), .Z(n3647) );
  XOR U354 ( .A(n4004), .B(n4053), .Z(n4008) );
  XOR U355 ( .A(n4365), .B(n4414), .Z(n4369) );
  XOR U356 ( .A(n4726), .B(n4775), .Z(n4730) );
  XOR U357 ( .A(n5087), .B(n5136), .Z(n5091) );
  XOR U358 ( .A(n5448), .B(n5497), .Z(n5452) );
  XOR U359 ( .A(n8446), .B(n8479), .Z(n8450) );
  XOR U360 ( .A(n8360), .B(n8393), .Z(n8364) );
  XOR U361 ( .A(n8250), .B(n8283), .Z(n8254) );
  XOR U362 ( .A(n8116), .B(n8149), .Z(n8120) );
  XOR U363 ( .A(n7958), .B(n7991), .Z(n7962) );
  XOR U364 ( .A(n7776), .B(n7809), .Z(n7780) );
  XOR U365 ( .A(n7570), .B(n7603), .Z(n7574) );
  XOR U366 ( .A(n7340), .B(n7373), .Z(n7344) );
  XOR U367 ( .A(n7086), .B(n7119), .Z(n7090) );
  XOR U368 ( .A(n6808), .B(n6841), .Z(n6812) );
  XOR U369 ( .A(n6506), .B(n6539), .Z(n6510) );
  XOR U370 ( .A(n6180), .B(n6213), .Z(n6184) );
  XOR U371 ( .A(n5827), .B(n5860), .Z(n5831) );
  XOR U372 ( .A(n401), .B(n431), .Z(n405) );
  XOR U373 ( .A(n762), .B(n793), .Z(n766) );
  XOR U374 ( .A(n1126), .B(n1157), .Z(n1130) );
  XOR U375 ( .A(n1489), .B(n1520), .Z(n1493) );
  XOR U376 ( .A(n1853), .B(n1884), .Z(n1857) );
  XOR U377 ( .A(n2214), .B(n2245), .Z(n2218) );
  XOR U378 ( .A(n2575), .B(n2606), .Z(n2579) );
  XOR U379 ( .A(n2936), .B(n2967), .Z(n2940) );
  XOR U380 ( .A(n3297), .B(n3328), .Z(n3301) );
  XOR U381 ( .A(n3658), .B(n3689), .Z(n3662) );
  XOR U382 ( .A(n4019), .B(n4050), .Z(n4023) );
  XOR U383 ( .A(n4380), .B(n4411), .Z(n4384) );
  XOR U384 ( .A(n4741), .B(n4772), .Z(n4745) );
  XOR U385 ( .A(n5102), .B(n5133), .Z(n5106) );
  XOR U386 ( .A(n5463), .B(n5494), .Z(n5467) );
  XOR U387 ( .A(n5893), .B(n6064), .Z(n5897) );
  XOR U388 ( .A(n5528), .B(n5700), .Z(n5533) );
  XOR U389 ( .A(n1555), .B(n1726), .Z(n1560) );
  XOR U390 ( .A(n1918), .B(n2087), .Z(n1923) );
  XOR U391 ( .A(n2279), .B(n2448), .Z(n2284) );
  XOR U392 ( .A(n2640), .B(n2809), .Z(n2645) );
  XOR U393 ( .A(n3001), .B(n3170), .Z(n3006) );
  XOR U394 ( .A(n3362), .B(n3531), .Z(n3367) );
  XOR U395 ( .A(n3723), .B(n3892), .Z(n3728) );
  XOR U396 ( .A(n4084), .B(n4253), .Z(n4089) );
  XOR U397 ( .A(n4445), .B(n4614), .Z(n4450) );
  XOR U398 ( .A(n4806), .B(n4975), .Z(n4811) );
  XOR U399 ( .A(n5167), .B(n5336), .Z(n5172) );
  XOR U400 ( .A(n6246), .B(n6399), .Z(n6250) );
  XOR U401 ( .A(n5908), .B(n6061), .Z(n5912) );
  XOR U402 ( .A(n5544), .B(n5697), .Z(n5548) );
  XOR U403 ( .A(n1571), .B(n1723), .Z(n1575) );
  XOR U404 ( .A(n1934), .B(n2084), .Z(n1938) );
  XOR U405 ( .A(n2295), .B(n2445), .Z(n2299) );
  XOR U406 ( .A(n2656), .B(n2806), .Z(n2660) );
  XOR U407 ( .A(n3017), .B(n3167), .Z(n3021) );
  XOR U408 ( .A(n3378), .B(n3528), .Z(n3382) );
  XOR U409 ( .A(n3739), .B(n3889), .Z(n3743) );
  XOR U410 ( .A(n4100), .B(n4250), .Z(n4104) );
  XOR U411 ( .A(n4461), .B(n4611), .Z(n4465) );
  XOR U412 ( .A(n4822), .B(n4972), .Z(n4826) );
  XOR U413 ( .A(n5183), .B(n5333), .Z(n5187) );
  XOR U414 ( .A(n6865), .B(n7000), .Z(n6869) );
  XOR U415 ( .A(n6575), .B(n6710), .Z(n6579) );
  XOR U416 ( .A(n6261), .B(n6396), .Z(n6265) );
  XOR U417 ( .A(n5923), .B(n6058), .Z(n5927) );
  XOR U418 ( .A(n5559), .B(n5694), .Z(n5563) );
  XOR U419 ( .A(n1203), .B(n1360), .Z(n1207) );
  XOR U420 ( .A(n1586), .B(n1719), .Z(n1590) );
  XOR U421 ( .A(n1949), .B(n2081), .Z(n1953) );
  XOR U422 ( .A(n2310), .B(n2442), .Z(n2314) );
  XOR U423 ( .A(n2671), .B(n2803), .Z(n2675) );
  XOR U424 ( .A(n3032), .B(n3164), .Z(n3036) );
  XOR U425 ( .A(n3393), .B(n3525), .Z(n3397) );
  XOR U426 ( .A(n3754), .B(n3886), .Z(n3758) );
  XOR U427 ( .A(n4115), .B(n4247), .Z(n4119) );
  XOR U428 ( .A(n4476), .B(n4608), .Z(n4480) );
  XOR U429 ( .A(n4837), .B(n4969), .Z(n4841) );
  XOR U430 ( .A(n5198), .B(n5330), .Z(n5202) );
  XOR U431 ( .A(n7146), .B(n7263), .Z(n7150) );
  XOR U432 ( .A(n6880), .B(n6997), .Z(n6884) );
  XOR U433 ( .A(n6590), .B(n6707), .Z(n6594) );
  XOR U434 ( .A(n6276), .B(n6393), .Z(n6280) );
  XOR U435 ( .A(n5938), .B(n6055), .Z(n5942) );
  XOR U436 ( .A(n5574), .B(n5691), .Z(n5578) );
  XOR U437 ( .A(n1409), .B(n1536), .Z(n1413) );
  XOR U438 ( .A(n1026), .B(n1178), .Z(n1030) );
  XOR U439 ( .A(n1964), .B(n2078), .Z(n1968) );
  XOR U440 ( .A(n2325), .B(n2439), .Z(n2329) );
  XOR U441 ( .A(n2686), .B(n2800), .Z(n2690) );
  XOR U442 ( .A(n3047), .B(n3161), .Z(n3051) );
  XOR U443 ( .A(n3408), .B(n3522), .Z(n3412) );
  XOR U444 ( .A(n3769), .B(n3883), .Z(n3773) );
  XOR U445 ( .A(n4130), .B(n4244), .Z(n4134) );
  XOR U446 ( .A(n4491), .B(n4605), .Z(n4495) );
  XOR U447 ( .A(n4852), .B(n4966), .Z(n4856) );
  XOR U448 ( .A(n5213), .B(n5327), .Z(n5217) );
  XOR U449 ( .A(n1611), .B(n1713), .Z(n1615) );
  XOR U450 ( .A(n7621), .B(n7720), .Z(n7625) );
  XOR U451 ( .A(n7403), .B(n7502), .Z(n7407) );
  XOR U452 ( .A(n7161), .B(n7260), .Z(n7165) );
  XOR U453 ( .A(n6895), .B(n6994), .Z(n6899) );
  XOR U454 ( .A(n6605), .B(n6704), .Z(n6609) );
  XOR U455 ( .A(n6291), .B(n6390), .Z(n6295) );
  XOR U456 ( .A(n5953), .B(n6052), .Z(n5957) );
  XOR U457 ( .A(n5589), .B(n5688), .Z(n5593) );
  XOR U458 ( .A(n1041), .B(n1175), .Z(n1045) );
  XOR U459 ( .A(n657), .B(n815), .Z(n661) );
  XOR U460 ( .A(n1979), .B(n2075), .Z(n1983) );
  XOR U461 ( .A(n2340), .B(n2436), .Z(n2344) );
  XOR U462 ( .A(n2701), .B(n2797), .Z(n2705) );
  XOR U463 ( .A(n3062), .B(n3158), .Z(n3066) );
  XOR U464 ( .A(n3423), .B(n3519), .Z(n3427) );
  XOR U465 ( .A(n3784), .B(n3880), .Z(n3788) );
  XOR U466 ( .A(n4145), .B(n4241), .Z(n4149) );
  XOR U467 ( .A(n4506), .B(n4602), .Z(n4510) );
  XOR U468 ( .A(n4867), .B(n4963), .Z(n4871) );
  XOR U469 ( .A(n5228), .B(n5324), .Z(n5232) );
  XOR U470 ( .A(n692), .B(n808), .Z(n696) );
  XOR U471 ( .A(n1243), .B(n1352), .Z(n1247) );
  XOR U472 ( .A(n1263), .B(n1347), .Z(n1267) );
  XOR U473 ( .A(n7830), .B(n7911), .Z(n7834) );
  XOR U474 ( .A(n7636), .B(n7717), .Z(n7640) );
  XOR U475 ( .A(n7418), .B(n7499), .Z(n7422) );
  XOR U476 ( .A(n7176), .B(n7257), .Z(n7180) );
  XOR U477 ( .A(n6910), .B(n6991), .Z(n6914) );
  XOR U478 ( .A(n6620), .B(n6701), .Z(n6624) );
  XOR U479 ( .A(n6306), .B(n6387), .Z(n6310) );
  XOR U480 ( .A(n5968), .B(n6049), .Z(n5972) );
  XOR U481 ( .A(n5604), .B(n5685), .Z(n5608) );
  XOR U482 ( .A(n864), .B(n992), .Z(n868) );
  XOR U483 ( .A(n481), .B(n632), .Z(n485) );
  XOR U484 ( .A(n717), .B(n802), .Z(n721) );
  XOR U485 ( .A(n1631), .B(n1709), .Z(n1635) );
  XOR U486 ( .A(n1994), .B(n2072), .Z(n1998) );
  XOR U487 ( .A(n2355), .B(n2433), .Z(n2359) );
  XOR U488 ( .A(n2716), .B(n2794), .Z(n2720) );
  XOR U489 ( .A(n3077), .B(n3155), .Z(n3081) );
  XOR U490 ( .A(n3438), .B(n3516), .Z(n3442) );
  XOR U491 ( .A(n3799), .B(n3877), .Z(n3803) );
  XOR U492 ( .A(n4160), .B(n4238), .Z(n4164) );
  XOR U493 ( .A(n4521), .B(n4599), .Z(n4525) );
  XOR U494 ( .A(n4882), .B(n4960), .Z(n4886) );
  XOR U495 ( .A(n5243), .B(n5321), .Z(n5247) );
  XOR U496 ( .A(n894), .B(n986), .Z(n898) );
  XOR U497 ( .A(n341), .B(n443), .Z(n345) );
  XOR U498 ( .A(n516), .B(n625), .Z(n520) );
  XOR U499 ( .A(n371), .B(n437), .Z(n375) );
  XOR U500 ( .A(n914), .B(n981), .Z(n918) );
  XOR U501 ( .A(n8161), .B(n8224), .Z(n8165) );
  XOR U502 ( .A(n8015), .B(n8078), .Z(n8019) );
  XOR U503 ( .A(n7845), .B(n7908), .Z(n7849) );
  XOR U504 ( .A(n7651), .B(n7714), .Z(n7655) );
  XOR U505 ( .A(n7433), .B(n7496), .Z(n7437) );
  XOR U506 ( .A(n7191), .B(n7254), .Z(n7195) );
  XOR U507 ( .A(n6925), .B(n6988), .Z(n6929) );
  XOR U508 ( .A(n6635), .B(n6698), .Z(n6639) );
  XOR U509 ( .A(n6321), .B(n6384), .Z(n6325) );
  XOR U510 ( .A(n5983), .B(n6046), .Z(n5987) );
  XOR U511 ( .A(n5619), .B(n5682), .Z(n5623) );
  XOR U512 ( .A(n496), .B(n629), .Z(n500) );
  XOR U513 ( .A(n1283), .B(n1343), .Z(n1287) );
  XOR U514 ( .A(n1646), .B(n1706), .Z(n1650) );
  XOR U515 ( .A(n2009), .B(n2069), .Z(n2013) );
  XOR U516 ( .A(n2370), .B(n2430), .Z(n2374) );
  XOR U517 ( .A(n2731), .B(n2791), .Z(n2735) );
  XOR U518 ( .A(n3092), .B(n3152), .Z(n3096) );
  XOR U519 ( .A(n3453), .B(n3513), .Z(n3457) );
  XOR U520 ( .A(n3814), .B(n3874), .Z(n3818) );
  XOR U521 ( .A(n4175), .B(n4235), .Z(n4179) );
  XOR U522 ( .A(n4536), .B(n4596), .Z(n4540) );
  XOR U523 ( .A(n4897), .B(n4957), .Z(n4901) );
  XOR U524 ( .A(n5258), .B(n5318), .Z(n5262) );
  XOR U525 ( .A(n546), .B(n619), .Z(n550) );
  XOR U526 ( .A(n8298), .B(n8343), .Z(n8302) );
  XOR U527 ( .A(n8176), .B(n8221), .Z(n8180) );
  XOR U528 ( .A(n8030), .B(n8075), .Z(n8034) );
  XOR U529 ( .A(n7860), .B(n7905), .Z(n7864) );
  XOR U530 ( .A(n7666), .B(n7711), .Z(n7670) );
  XOR U531 ( .A(n7448), .B(n7493), .Z(n7452) );
  XOR U532 ( .A(n7206), .B(n7251), .Z(n7210) );
  XOR U533 ( .A(n6940), .B(n6985), .Z(n6944) );
  XOR U534 ( .A(n6650), .B(n6695), .Z(n6654) );
  XOR U535 ( .A(n6336), .B(n6381), .Z(n6340) );
  XOR U536 ( .A(n5998), .B(n6043), .Z(n6002) );
  XOR U537 ( .A(n5634), .B(n5679), .Z(n5638) );
  XOR U538 ( .A(n571), .B(n613), .Z(n575) );
  XOR U539 ( .A(n934), .B(n976), .Z(n938) );
  XOR U540 ( .A(n1298), .B(n1340), .Z(n1302) );
  XOR U541 ( .A(n1661), .B(n1703), .Z(n1665) );
  XOR U542 ( .A(n2024), .B(n2066), .Z(n2028) );
  XOR U543 ( .A(n2385), .B(n2427), .Z(n2389) );
  XOR U544 ( .A(n2746), .B(n2788), .Z(n2750) );
  XOR U545 ( .A(n3107), .B(n3149), .Z(n3111) );
  XOR U546 ( .A(n3468), .B(n3510), .Z(n3472) );
  XOR U547 ( .A(n3829), .B(n3871), .Z(n3833) );
  XOR U548 ( .A(n4190), .B(n4232), .Z(n4194) );
  XOR U549 ( .A(n4551), .B(n4593), .Z(n4555) );
  XOR U550 ( .A(n4912), .B(n4954), .Z(n4916) );
  XOR U551 ( .A(n5273), .B(n5315), .Z(n5277) );
  XOR U552 ( .A(n8485), .B(n8512), .Z(n8489) );
  XOR U553 ( .A(n8411), .B(n8438), .Z(n8415) );
  XOR U554 ( .A(n8313), .B(n8340), .Z(n8317) );
  XOR U555 ( .A(n8191), .B(n8218), .Z(n8195) );
  XOR U556 ( .A(n8045), .B(n8072), .Z(n8049) );
  XOR U557 ( .A(n7875), .B(n7902), .Z(n7879) );
  XOR U558 ( .A(n7681), .B(n7708), .Z(n7685) );
  XOR U559 ( .A(n7463), .B(n7490), .Z(n7467) );
  XOR U560 ( .A(n7221), .B(n7248), .Z(n7225) );
  XOR U561 ( .A(n6955), .B(n6982), .Z(n6959) );
  XOR U562 ( .A(n6665), .B(n6692), .Z(n6669) );
  XOR U563 ( .A(n6351), .B(n6378), .Z(n6355) );
  XOR U564 ( .A(n6013), .B(n6040), .Z(n6017) );
  XOR U565 ( .A(n5649), .B(n5676), .Z(n5653) );
  XOR U566 ( .A(n586), .B(n610), .Z(n590) );
  XOR U567 ( .A(n949), .B(n973), .Z(n953) );
  XOR U568 ( .A(n1313), .B(n1337), .Z(n1317) );
  XOR U569 ( .A(n1676), .B(n1700), .Z(n1680) );
  XOR U570 ( .A(n2039), .B(n2063), .Z(n2043) );
  XOR U571 ( .A(n2400), .B(n2424), .Z(n2404) );
  XOR U572 ( .A(n2761), .B(n2785), .Z(n2765) );
  XOR U573 ( .A(n3122), .B(n3146), .Z(n3126) );
  XOR U574 ( .A(n3483), .B(n3507), .Z(n3487) );
  XOR U575 ( .A(n3844), .B(n3868), .Z(n3848) );
  XOR U576 ( .A(n4205), .B(n4229), .Z(n4209) );
  XOR U577 ( .A(n4566), .B(n4590), .Z(n4570) );
  XOR U578 ( .A(n4927), .B(n4951), .Z(n4931) );
  XOR U579 ( .A(n5288), .B(n5312), .Z(n5292) );
  AND U580 ( .A(n602), .B(n601), .Z(n421) );
  AND U581 ( .A(n1329), .B(n1328), .Z(n1146) );
  AND U582 ( .A(n2055), .B(n2054), .Z(n1873) );
  AND U583 ( .A(n2777), .B(n2776), .Z(n2595) );
  AND U584 ( .A(n3499), .B(n3498), .Z(n3317) );
  AND U585 ( .A(n4221), .B(n4220), .Z(n4039) );
  AND U586 ( .A(n4943), .B(n4942), .Z(n4761) );
  XOR U587 ( .A(n5711), .B(n5883), .Z(n5716) );
  XOR U588 ( .A(n1737), .B(n1907), .Z(n1742) );
  XOR U589 ( .A(n2098), .B(n2268), .Z(n2103) );
  XOR U590 ( .A(n2459), .B(n2629), .Z(n2464) );
  XOR U591 ( .A(n2820), .B(n2990), .Z(n2825) );
  XOR U592 ( .A(n3181), .B(n3351), .Z(n3186) );
  XOR U593 ( .A(n3542), .B(n3712), .Z(n3547) );
  XOR U594 ( .A(n3903), .B(n4073), .Z(n3908) );
  XOR U595 ( .A(n4264), .B(n4434), .Z(n4269) );
  XOR U596 ( .A(n4625), .B(n4795), .Z(n4630) );
  XOR U597 ( .A(n4986), .B(n5156), .Z(n4991) );
  XOR U598 ( .A(n5347), .B(n5517), .Z(n5352) );
  XOR U599 ( .A(n6406), .B(n6559), .Z(n6410) );
  XOR U600 ( .A(n6080), .B(n6233), .Z(n6084) );
  XOR U601 ( .A(n5727), .B(n5880), .Z(n5731) );
  XOR U602 ( .A(n1753), .B(n1904), .Z(n1757) );
  XOR U603 ( .A(n2114), .B(n2265), .Z(n2118) );
  XOR U604 ( .A(n2475), .B(n2626), .Z(n2479) );
  XOR U605 ( .A(n2836), .B(n2987), .Z(n2840) );
  XOR U606 ( .A(n3197), .B(n3348), .Z(n3201) );
  XOR U607 ( .A(n3558), .B(n3709), .Z(n3562) );
  XOR U608 ( .A(n3919), .B(n4070), .Z(n3923) );
  XOR U609 ( .A(n4280), .B(n4431), .Z(n4284) );
  XOR U610 ( .A(n4641), .B(n4792), .Z(n4645) );
  XOR U611 ( .A(n5002), .B(n5153), .Z(n5006) );
  XOR U612 ( .A(n5363), .B(n5514), .Z(n5367) );
  XOR U613 ( .A(n1389), .B(n1541), .Z(n1393) );
  XOR U614 ( .A(n6723), .B(n6858), .Z(n6727) );
  XOR U615 ( .A(n6421), .B(n6556), .Z(n6425) );
  XOR U616 ( .A(n6095), .B(n6230), .Z(n6099) );
  XOR U617 ( .A(n5742), .B(n5877), .Z(n5746) );
  XOR U618 ( .A(n1010), .B(n1181), .Z(n1015) );
  XOR U619 ( .A(n1768), .B(n1901), .Z(n1772) );
  XOR U620 ( .A(n2129), .B(n2262), .Z(n2133) );
  XOR U621 ( .A(n2490), .B(n2623), .Z(n2494) );
  XOR U622 ( .A(n2851), .B(n2984), .Z(n2855) );
  XOR U623 ( .A(n3212), .B(n3345), .Z(n3216) );
  XOR U624 ( .A(n3573), .B(n3706), .Z(n3577) );
  XOR U625 ( .A(n3934), .B(n4067), .Z(n3938) );
  XOR U626 ( .A(n4295), .B(n4428), .Z(n4299) );
  XOR U627 ( .A(n4656), .B(n4789), .Z(n4660) );
  XOR U628 ( .A(n5017), .B(n5150), .Z(n5021) );
  XOR U629 ( .A(n5378), .B(n5511), .Z(n5382) );
  XOR U630 ( .A(n7270), .B(n7387), .Z(n7274) );
  XOR U631 ( .A(n7016), .B(n7133), .Z(n7020) );
  XOR U632 ( .A(n6738), .B(n6855), .Z(n6742) );
  XOR U633 ( .A(n6436), .B(n6553), .Z(n6440) );
  XOR U634 ( .A(n6110), .B(n6227), .Z(n6114) );
  XOR U635 ( .A(n5757), .B(n5874), .Z(n5761) );
  XOR U636 ( .A(n1218), .B(n1357), .Z(n1222) );
  XOR U637 ( .A(n834), .B(n998), .Z(n838) );
  XOR U638 ( .A(n1783), .B(n1898), .Z(n1787) );
  XOR U639 ( .A(n2144), .B(n2259), .Z(n2148) );
  XOR U640 ( .A(n2505), .B(n2620), .Z(n2509) );
  XOR U641 ( .A(n2866), .B(n2981), .Z(n2870) );
  XOR U642 ( .A(n3227), .B(n3342), .Z(n3231) );
  XOR U643 ( .A(n3588), .B(n3703), .Z(n3592) );
  XOR U644 ( .A(n3949), .B(n4064), .Z(n3953) );
  XOR U645 ( .A(n4310), .B(n4425), .Z(n4314) );
  XOR U646 ( .A(n4671), .B(n4786), .Z(n4675) );
  XOR U647 ( .A(n5032), .B(n5147), .Z(n5036) );
  XOR U648 ( .A(n5393), .B(n5508), .Z(n5397) );
  XOR U649 ( .A(n1414), .B(n1535), .Z(n1418) );
  XOR U650 ( .A(n7515), .B(n7614), .Z(n7519) );
  XOR U651 ( .A(n7285), .B(n7384), .Z(n7289) );
  XOR U652 ( .A(n7031), .B(n7130), .Z(n7035) );
  XOR U653 ( .A(n6753), .B(n6852), .Z(n6757) );
  XOR U654 ( .A(n6451), .B(n6550), .Z(n6455) );
  XOR U655 ( .A(n6125), .B(n6224), .Z(n6129) );
  XOR U656 ( .A(n5772), .B(n5871), .Z(n5776) );
  XOR U657 ( .A(n1066), .B(n1169), .Z(n1070) );
  XOR U658 ( .A(n849), .B(n995), .Z(n853) );
  XOR U659 ( .A(n465), .B(n635), .Z(n470) );
  XOR U660 ( .A(n1434), .B(n1531), .Z(n1438) );
  XOR U661 ( .A(n1798), .B(n1895), .Z(n1802) );
  XOR U662 ( .A(n2159), .B(n2256), .Z(n2163) );
  XOR U663 ( .A(n2520), .B(n2617), .Z(n2524) );
  XOR U664 ( .A(n2881), .B(n2978), .Z(n2885) );
  XOR U665 ( .A(n3242), .B(n3339), .Z(n3246) );
  XOR U666 ( .A(n3603), .B(n3700), .Z(n3607) );
  XOR U667 ( .A(n3964), .B(n4061), .Z(n3968) );
  XOR U668 ( .A(n4325), .B(n4422), .Z(n4329) );
  XOR U669 ( .A(n4686), .B(n4783), .Z(n4690) );
  XOR U670 ( .A(n5047), .B(n5144), .Z(n5051) );
  XOR U671 ( .A(n5408), .B(n5505), .Z(n5412) );
  XOR U672 ( .A(n1238), .B(n1353), .Z(n1242) );
  XOR U673 ( .A(n501), .B(n628), .Z(n505) );
  XOR U674 ( .A(n7918), .B(n7999), .Z(n7922) );
  XOR U675 ( .A(n7736), .B(n7817), .Z(n7740) );
  XOR U676 ( .A(n7530), .B(n7611), .Z(n7534) );
  XOR U677 ( .A(n7300), .B(n7381), .Z(n7304) );
  XOR U678 ( .A(n7046), .B(n7127), .Z(n7050) );
  XOR U679 ( .A(n6768), .B(n6849), .Z(n6772) );
  XOR U680 ( .A(n6466), .B(n6547), .Z(n6470) );
  XOR U681 ( .A(n6140), .B(n6221), .Z(n6144) );
  XOR U682 ( .A(n5787), .B(n5868), .Z(n5791) );
  XOR U683 ( .A(n889), .B(n987), .Z(n893) );
  XOR U684 ( .A(n672), .B(n812), .Z(n676) );
  XOR U685 ( .A(n291), .B(n453), .Z(n295) );
  XOR U686 ( .A(n1086), .B(n1165), .Z(n1090) );
  XOR U687 ( .A(n1449), .B(n1528), .Z(n1453) );
  XOR U688 ( .A(n1813), .B(n1892), .Z(n1817) );
  XOR U689 ( .A(n2174), .B(n2253), .Z(n2178) );
  XOR U690 ( .A(n2535), .B(n2614), .Z(n2539) );
  XOR U691 ( .A(n2896), .B(n2975), .Z(n2900) );
  XOR U692 ( .A(n3257), .B(n3336), .Z(n3261) );
  XOR U693 ( .A(n3618), .B(n3697), .Z(n3622) );
  XOR U694 ( .A(n3979), .B(n4058), .Z(n3983) );
  XOR U695 ( .A(n4340), .B(n4419), .Z(n4344) );
  XOR U696 ( .A(n4701), .B(n4780), .Z(n4705) );
  XOR U697 ( .A(n5062), .B(n5141), .Z(n5066) );
  XOR U698 ( .A(n5423), .B(n5502), .Z(n5427) );
  XOR U699 ( .A(n869), .B(n991), .Z(n873) );
  XOR U700 ( .A(n722), .B(n801), .Z(n726) );
  XOR U701 ( .A(n326), .B(n446), .Z(n330) );
  XOR U702 ( .A(n8091), .B(n8154), .Z(n8095) );
  XOR U703 ( .A(n7933), .B(n7996), .Z(n7937) );
  XOR U704 ( .A(n7751), .B(n7814), .Z(n7755) );
  XOR U705 ( .A(n7545), .B(n7608), .Z(n7549) );
  XOR U706 ( .A(n7315), .B(n7378), .Z(n7319) );
  XOR U707 ( .A(n7061), .B(n7124), .Z(n7065) );
  XOR U708 ( .A(n6783), .B(n6846), .Z(n6787) );
  XOR U709 ( .A(n6481), .B(n6544), .Z(n6485) );
  XOR U710 ( .A(n6155), .B(n6218), .Z(n6159) );
  XOR U711 ( .A(n5802), .B(n5865), .Z(n5806) );
  XOR U712 ( .A(n521), .B(n624), .Z(n525) );
  XOR U713 ( .A(n306), .B(n450), .Z(n310) );
  XOR U714 ( .A(n376), .B(n436), .Z(n380) );
  XOR U715 ( .A(n1101), .B(n1162), .Z(n1105) );
  XOR U716 ( .A(n1464), .B(n1525), .Z(n1468) );
  XOR U717 ( .A(n1828), .B(n1889), .Z(n1832) );
  XOR U718 ( .A(n2189), .B(n2250), .Z(n2193) );
  XOR U719 ( .A(n2550), .B(n2611), .Z(n2554) );
  XOR U720 ( .A(n2911), .B(n2972), .Z(n2915) );
  XOR U721 ( .A(n3272), .B(n3333), .Z(n3276) );
  XOR U722 ( .A(n3633), .B(n3694), .Z(n3637) );
  XOR U723 ( .A(n3994), .B(n4055), .Z(n3998) );
  XOR U724 ( .A(n4355), .B(n4416), .Z(n4359) );
  XOR U725 ( .A(n4716), .B(n4777), .Z(n4720) );
  XOR U726 ( .A(n5077), .B(n5138), .Z(n5081) );
  XOR U727 ( .A(n5438), .B(n5499), .Z(n5442) );
  XOR U728 ( .A(n356), .B(n440), .Z(n360) );
  XOR U729 ( .A(n551), .B(n618), .Z(n555) );
  XOR U730 ( .A(n8350), .B(n8395), .Z(n8354) );
  XOR U731 ( .A(n8240), .B(n8285), .Z(n8244) );
  XOR U732 ( .A(n8106), .B(n8151), .Z(n8110) );
  XOR U733 ( .A(n7948), .B(n7993), .Z(n7952) );
  XOR U734 ( .A(n7766), .B(n7811), .Z(n7770) );
  XOR U735 ( .A(n7560), .B(n7605), .Z(n7564) );
  XOR U736 ( .A(n7330), .B(n7375), .Z(n7334) );
  XOR U737 ( .A(n7076), .B(n7121), .Z(n7080) );
  XOR U738 ( .A(n6798), .B(n6843), .Z(n6802) );
  XOR U739 ( .A(n6496), .B(n6541), .Z(n6500) );
  XOR U740 ( .A(n6170), .B(n6215), .Z(n6174) );
  XOR U741 ( .A(n5817), .B(n5862), .Z(n5821) );
  XOR U742 ( .A(n391), .B(n433), .Z(n395) );
  XOR U743 ( .A(n752), .B(n795), .Z(n756) );
  XOR U744 ( .A(n1116), .B(n1159), .Z(n1120) );
  XOR U745 ( .A(n1479), .B(n1522), .Z(n1483) );
  XOR U746 ( .A(n1843), .B(n1886), .Z(n1847) );
  XOR U747 ( .A(n2204), .B(n2247), .Z(n2208) );
  XOR U748 ( .A(n2565), .B(n2608), .Z(n2569) );
  XOR U749 ( .A(n2926), .B(n2969), .Z(n2930) );
  XOR U750 ( .A(n3287), .B(n3330), .Z(n3291) );
  XOR U751 ( .A(n3648), .B(n3691), .Z(n3652) );
  XOR U752 ( .A(n4009), .B(n4052), .Z(n4013) );
  XOR U753 ( .A(n4370), .B(n4413), .Z(n4374) );
  XOR U754 ( .A(n4731), .B(n4774), .Z(n4735) );
  XOR U755 ( .A(n5092), .B(n5135), .Z(n5096) );
  XOR U756 ( .A(n5453), .B(n5496), .Z(n5457) );
  XOR U757 ( .A(n8451), .B(n8478), .Z(n8455) );
  XOR U758 ( .A(n8365), .B(n8392), .Z(n8369) );
  XOR U759 ( .A(n8255), .B(n8282), .Z(n8259) );
  XOR U760 ( .A(n8121), .B(n8148), .Z(n8125) );
  XOR U761 ( .A(n7963), .B(n7990), .Z(n7967) );
  XOR U762 ( .A(n7781), .B(n7808), .Z(n7785) );
  XOR U763 ( .A(n7575), .B(n7602), .Z(n7579) );
  XOR U764 ( .A(n7345), .B(n7372), .Z(n7349) );
  XOR U765 ( .A(n7091), .B(n7118), .Z(n7095) );
  XOR U766 ( .A(n6813), .B(n6840), .Z(n6817) );
  XOR U767 ( .A(n6511), .B(n6538), .Z(n6515) );
  XOR U768 ( .A(n6185), .B(n6212), .Z(n6189) );
  XOR U769 ( .A(n5832), .B(n5859), .Z(n5836) );
  XOR U770 ( .A(n406), .B(n430), .Z(n410) );
  XOR U771 ( .A(n767), .B(n792), .Z(n771) );
  XOR U772 ( .A(n1131), .B(n1156), .Z(n1135) );
  XOR U773 ( .A(n1494), .B(n1519), .Z(n1498) );
  XOR U774 ( .A(n1858), .B(n1883), .Z(n1862) );
  XOR U775 ( .A(n2219), .B(n2244), .Z(n2223) );
  XOR U776 ( .A(n2580), .B(n2605), .Z(n2584) );
  XOR U777 ( .A(n2941), .B(n2966), .Z(n2945) );
  XOR U778 ( .A(n3302), .B(n3327), .Z(n3306) );
  XOR U779 ( .A(n3663), .B(n3688), .Z(n3667) );
  XOR U780 ( .A(n4024), .B(n4049), .Z(n4028) );
  XOR U781 ( .A(n4385), .B(n4410), .Z(n4389) );
  XOR U782 ( .A(n4746), .B(n4771), .Z(n4750) );
  XOR U783 ( .A(n5107), .B(n5132), .Z(n5111) );
  XOR U784 ( .A(n5468), .B(n5493), .Z(n5472) );
  AND U785 ( .A(n783), .B(n782), .Z(n601) );
  AND U786 ( .A(n1510), .B(n1509), .Z(n1328) );
  AND U787 ( .A(n2235), .B(n2234), .Z(n2054) );
  AND U788 ( .A(n2957), .B(n2956), .Z(n2776) );
  AND U789 ( .A(n3679), .B(n3678), .Z(n3498) );
  AND U790 ( .A(n4401), .B(n4400), .Z(n4220) );
  AND U791 ( .A(n5123), .B(n5122), .Z(n4942) );
  XOR U792 ( .A(n5898), .B(n6063), .Z(n5902) );
  XOR U793 ( .A(n5534), .B(n5699), .Z(n5538) );
  XOR U794 ( .A(n1561), .B(n1725), .Z(n1565) );
  XOR U795 ( .A(n1924), .B(n2086), .Z(n1928) );
  XOR U796 ( .A(n2285), .B(n2447), .Z(n2289) );
  XOR U797 ( .A(n2646), .B(n2808), .Z(n2650) );
  XOR U798 ( .A(n3007), .B(n3169), .Z(n3011) );
  XOR U799 ( .A(n3368), .B(n3530), .Z(n3372) );
  XOR U800 ( .A(n3729), .B(n3891), .Z(n3733) );
  XOR U801 ( .A(n4090), .B(n4252), .Z(n4094) );
  XOR U802 ( .A(n4451), .B(n4613), .Z(n4455) );
  XOR U803 ( .A(n4812), .B(n4974), .Z(n4816) );
  XOR U804 ( .A(n5173), .B(n5335), .Z(n5177) );
  XOR U805 ( .A(n6565), .B(n6712), .Z(n6569) );
  XOR U806 ( .A(n6251), .B(n6398), .Z(n6255) );
  XOR U807 ( .A(n5913), .B(n6060), .Z(n5917) );
  XOR U808 ( .A(n5549), .B(n5696), .Z(n5553) );
  XOR U809 ( .A(n1192), .B(n1362), .Z(n1197) );
  XOR U810 ( .A(n1576), .B(n1722), .Z(n1580) );
  XOR U811 ( .A(n1939), .B(n2083), .Z(n1943) );
  XOR U812 ( .A(n2300), .B(n2444), .Z(n2304) );
  XOR U813 ( .A(n2661), .B(n2805), .Z(n2665) );
  XOR U814 ( .A(n3022), .B(n3166), .Z(n3026) );
  XOR U815 ( .A(n3383), .B(n3527), .Z(n3387) );
  XOR U816 ( .A(n3744), .B(n3888), .Z(n3748) );
  XOR U817 ( .A(n4105), .B(n4249), .Z(n4109) );
  XOR U818 ( .A(n4466), .B(n4610), .Z(n4470) );
  XOR U819 ( .A(n4827), .B(n4971), .Z(n4831) );
  XOR U820 ( .A(n5188), .B(n5332), .Z(n5192) );
  XOR U821 ( .A(n6870), .B(n6999), .Z(n6874) );
  XOR U822 ( .A(n6580), .B(n6709), .Z(n6584) );
  XOR U823 ( .A(n6266), .B(n6395), .Z(n6270) );
  XOR U824 ( .A(n5928), .B(n6057), .Z(n5932) );
  XOR U825 ( .A(n5564), .B(n5693), .Z(n5568) );
  XOR U826 ( .A(n1399), .B(n1539), .Z(n1403) );
  XOR U827 ( .A(n1016), .B(n1180), .Z(n1020) );
  XOR U828 ( .A(n1954), .B(n2080), .Z(n1958) );
  XOR U829 ( .A(n2315), .B(n2441), .Z(n2319) );
  XOR U830 ( .A(n2676), .B(n2802), .Z(n2680) );
  XOR U831 ( .A(n3037), .B(n3163), .Z(n3041) );
  XOR U832 ( .A(n3398), .B(n3524), .Z(n3402) );
  XOR U833 ( .A(n3759), .B(n3885), .Z(n3763) );
  XOR U834 ( .A(n4120), .B(n4246), .Z(n4124) );
  XOR U835 ( .A(n4481), .B(n4607), .Z(n4485) );
  XOR U836 ( .A(n4842), .B(n4968), .Z(n4846) );
  XOR U837 ( .A(n5203), .B(n5329), .Z(n5207) );
  XOR U838 ( .A(n1601), .B(n1716), .Z(n1605) );
  XOR U839 ( .A(n7393), .B(n7504), .Z(n7397) );
  XOR U840 ( .A(n7151), .B(n7262), .Z(n7155) );
  XOR U841 ( .A(n6885), .B(n6996), .Z(n6889) );
  XOR U842 ( .A(n6595), .B(n6706), .Z(n6599) );
  XOR U843 ( .A(n6281), .B(n6392), .Z(n6285) );
  XOR U844 ( .A(n5943), .B(n6054), .Z(n5947) );
  XOR U845 ( .A(n5579), .B(n5690), .Z(n5583) );
  XOR U846 ( .A(n1031), .B(n1177), .Z(n1035) );
  XOR U847 ( .A(n646), .B(n817), .Z(n651) );
  XOR U848 ( .A(n1969), .B(n2077), .Z(n1973) );
  XOR U849 ( .A(n2330), .B(n2438), .Z(n2334) );
  XOR U850 ( .A(n2691), .B(n2799), .Z(n2695) );
  XOR U851 ( .A(n3052), .B(n3160), .Z(n3056) );
  XOR U852 ( .A(n3413), .B(n3521), .Z(n3417) );
  XOR U853 ( .A(n3774), .B(n3882), .Z(n3778) );
  XOR U854 ( .A(n4135), .B(n4243), .Z(n4139) );
  XOR U855 ( .A(n4496), .B(n4604), .Z(n4500) );
  XOR U856 ( .A(n4857), .B(n4965), .Z(n4861) );
  XOR U857 ( .A(n5218), .B(n5326), .Z(n5222) );
  XOR U858 ( .A(n1233), .B(n1354), .Z(n1237) );
  XOR U859 ( .A(n1253), .B(n1350), .Z(n1257) );
  XOR U860 ( .A(n7626), .B(n7719), .Z(n7630) );
  XOR U861 ( .A(n7408), .B(n7501), .Z(n7412) );
  XOR U862 ( .A(n7166), .B(n7259), .Z(n7170) );
  XOR U863 ( .A(n6900), .B(n6993), .Z(n6904) );
  XOR U864 ( .A(n6610), .B(n6703), .Z(n6614) );
  XOR U865 ( .A(n6296), .B(n6389), .Z(n6300) );
  XOR U866 ( .A(n5958), .B(n6051), .Z(n5962) );
  XOR U867 ( .A(n5594), .B(n5687), .Z(n5598) );
  XOR U868 ( .A(n854), .B(n994), .Z(n858) );
  XOR U869 ( .A(n471), .B(n634), .Z(n475) );
  XOR U870 ( .A(n1621), .B(n1711), .Z(n1625) );
  XOR U871 ( .A(n1984), .B(n2074), .Z(n1988) );
  XOR U872 ( .A(n2345), .B(n2435), .Z(n2349) );
  XOR U873 ( .A(n2706), .B(n2796), .Z(n2710) );
  XOR U874 ( .A(n3067), .B(n3157), .Z(n3071) );
  XOR U875 ( .A(n3428), .B(n3518), .Z(n3432) );
  XOR U876 ( .A(n3789), .B(n3879), .Z(n3793) );
  XOR U877 ( .A(n4150), .B(n4240), .Z(n4154) );
  XOR U878 ( .A(n4511), .B(n4601), .Z(n4515) );
  XOR U879 ( .A(n4872), .B(n4962), .Z(n4876) );
  XOR U880 ( .A(n5233), .B(n5323), .Z(n5237) );
  XOR U881 ( .A(n884), .B(n988), .Z(n888) );
  XOR U882 ( .A(n506), .B(n627), .Z(n510) );
  XOR U883 ( .A(n1056), .B(n1172), .Z(n1060) );
  XOR U884 ( .A(n8005), .B(n8080), .Z(n8009) );
  XOR U885 ( .A(n7835), .B(n7910), .Z(n7839) );
  XOR U886 ( .A(n7641), .B(n7716), .Z(n7645) );
  XOR U887 ( .A(n7423), .B(n7498), .Z(n7427) );
  XOR U888 ( .A(n7181), .B(n7256), .Z(n7185) );
  XOR U889 ( .A(n6915), .B(n6990), .Z(n6919) );
  XOR U890 ( .A(n6625), .B(n6700), .Z(n6629) );
  XOR U891 ( .A(n6311), .B(n6386), .Z(n6315) );
  XOR U892 ( .A(n5973), .B(n6048), .Z(n5977) );
  XOR U893 ( .A(n5609), .B(n5684), .Z(n5613) );
  XOR U894 ( .A(n677), .B(n811), .Z(n681) );
  XOR U895 ( .A(n296), .B(n452), .Z(n300) );
  XOR U896 ( .A(n909), .B(n982), .Z(n913) );
  XOR U897 ( .A(n1273), .B(n1345), .Z(n1277) );
  XOR U898 ( .A(n1636), .B(n1708), .Z(n1640) );
  XOR U899 ( .A(n1999), .B(n2071), .Z(n2003) );
  XOR U900 ( .A(n2360), .B(n2432), .Z(n2364) );
  XOR U901 ( .A(n2721), .B(n2793), .Z(n2725) );
  XOR U902 ( .A(n3082), .B(n3154), .Z(n3086) );
  XOR U903 ( .A(n3443), .B(n3515), .Z(n3447) );
  XOR U904 ( .A(n3804), .B(n3876), .Z(n3808) );
  XOR U905 ( .A(n4165), .B(n4237), .Z(n4169) );
  XOR U906 ( .A(n4526), .B(n4598), .Z(n4530) );
  XOR U907 ( .A(n4887), .B(n4959), .Z(n4891) );
  XOR U908 ( .A(n5248), .B(n5320), .Z(n5252) );
  XOR U909 ( .A(n707), .B(n805), .Z(n711) );
  XOR U910 ( .A(n346), .B(n442), .Z(n350) );
  XOR U911 ( .A(n331), .B(n445), .Z(n335) );
  XOR U912 ( .A(n8166), .B(n8223), .Z(n8170) );
  XOR U913 ( .A(n8020), .B(n8077), .Z(n8024) );
  XOR U914 ( .A(n7850), .B(n7907), .Z(n7854) );
  XOR U915 ( .A(n7656), .B(n7713), .Z(n7660) );
  XOR U916 ( .A(n7438), .B(n7495), .Z(n7442) );
  XOR U917 ( .A(n7196), .B(n7253), .Z(n7200) );
  XOR U918 ( .A(n6930), .B(n6987), .Z(n6934) );
  XOR U919 ( .A(n6640), .B(n6697), .Z(n6644) );
  XOR U920 ( .A(n6326), .B(n6383), .Z(n6330) );
  XOR U921 ( .A(n5988), .B(n6045), .Z(n5992) );
  XOR U922 ( .A(n5624), .B(n5681), .Z(n5628) );
  XOR U923 ( .A(n311), .B(n449), .Z(n315) );
  XOR U924 ( .A(n561), .B(n615), .Z(n565) );
  XOR U925 ( .A(n924), .B(n978), .Z(n928) );
  XOR U926 ( .A(n1288), .B(n1342), .Z(n1292) );
  XOR U927 ( .A(n1651), .B(n1705), .Z(n1655) );
  XOR U928 ( .A(n2014), .B(n2068), .Z(n2018) );
  XOR U929 ( .A(n2375), .B(n2429), .Z(n2379) );
  XOR U930 ( .A(n2736), .B(n2790), .Z(n2740) );
  XOR U931 ( .A(n3097), .B(n3151), .Z(n3101) );
  XOR U932 ( .A(n3458), .B(n3512), .Z(n3462) );
  XOR U933 ( .A(n3819), .B(n3873), .Z(n3823) );
  XOR U934 ( .A(n4180), .B(n4234), .Z(n4184) );
  XOR U935 ( .A(n4541), .B(n4595), .Z(n4545) );
  XOR U936 ( .A(n4902), .B(n4956), .Z(n4906) );
  XOR U937 ( .A(n5263), .B(n5317), .Z(n5267) );
  XOR U938 ( .A(n361), .B(n439), .Z(n365) );
  XOR U939 ( .A(n8401), .B(n8440), .Z(n8405) );
  XOR U940 ( .A(n8303), .B(n8342), .Z(n8307) );
  XOR U941 ( .A(n8181), .B(n8220), .Z(n8185) );
  XOR U942 ( .A(n8035), .B(n8074), .Z(n8039) );
  XOR U943 ( .A(n7865), .B(n7904), .Z(n7869) );
  XOR U944 ( .A(n7671), .B(n7710), .Z(n7675) );
  XOR U945 ( .A(n7453), .B(n7492), .Z(n7457) );
  XOR U946 ( .A(n7211), .B(n7250), .Z(n7215) );
  XOR U947 ( .A(n6945), .B(n6984), .Z(n6949) );
  XOR U948 ( .A(n6655), .B(n6694), .Z(n6659) );
  XOR U949 ( .A(n6341), .B(n6380), .Z(n6345) );
  XOR U950 ( .A(n6003), .B(n6042), .Z(n6007) );
  XOR U951 ( .A(n5639), .B(n5678), .Z(n5643) );
  XOR U952 ( .A(n576), .B(n612), .Z(n580) );
  XOR U953 ( .A(n939), .B(n975), .Z(n943) );
  XOR U954 ( .A(n1303), .B(n1339), .Z(n1307) );
  XOR U955 ( .A(n1666), .B(n1702), .Z(n1670) );
  XOR U956 ( .A(n2029), .B(n2065), .Z(n2033) );
  XOR U957 ( .A(n2390), .B(n2426), .Z(n2394) );
  XOR U958 ( .A(n2751), .B(n2787), .Z(n2755) );
  XOR U959 ( .A(n3112), .B(n3148), .Z(n3116) );
  XOR U960 ( .A(n3473), .B(n3509), .Z(n3477) );
  XOR U961 ( .A(n3834), .B(n3870), .Z(n3838) );
  XOR U962 ( .A(n4195), .B(n4231), .Z(n4199) );
  XOR U963 ( .A(n4556), .B(n4592), .Z(n4560) );
  XOR U964 ( .A(n4917), .B(n4953), .Z(n4921) );
  XOR U965 ( .A(n5278), .B(n5314), .Z(n5282) );
  XOR U966 ( .A(n8490), .B(n8511), .Z(n8499) );
  XOR U967 ( .A(n8416), .B(n8437), .Z(n8425) );
  XOR U968 ( .A(n8318), .B(n8339), .Z(n8327) );
  XOR U969 ( .A(n8196), .B(n8217), .Z(n8205) );
  XOR U970 ( .A(n8050), .B(n8071), .Z(n8059) );
  XOR U971 ( .A(n7880), .B(n7901), .Z(n7889) );
  XOR U972 ( .A(n7686), .B(n7707), .Z(n7695) );
  XOR U973 ( .A(n7468), .B(n7489), .Z(n7477) );
  XOR U974 ( .A(n7226), .B(n7247), .Z(n7235) );
  XOR U975 ( .A(n6960), .B(n6981), .Z(n6969) );
  XOR U976 ( .A(n6670), .B(n6691), .Z(n6679) );
  XOR U977 ( .A(n6356), .B(n6377), .Z(n6365) );
  XOR U978 ( .A(n6018), .B(n6039), .Z(n6027) );
  XOR U979 ( .A(n5654), .B(n5675), .Z(n5663) );
  XOR U980 ( .A(n591), .B(n609), .Z(n600) );
  XOR U981 ( .A(n954), .B(n972), .Z(n963) );
  XOR U982 ( .A(n1318), .B(n1336), .Z(n1327) );
  XOR U983 ( .A(n1681), .B(n1699), .Z(n1690) );
  XOR U984 ( .A(n2044), .B(n2062), .Z(n2053) );
  XOR U985 ( .A(n2405), .B(n2423), .Z(n2414) );
  XOR U986 ( .A(n2766), .B(n2784), .Z(n2775) );
  XOR U987 ( .A(n3127), .B(n3145), .Z(n3136) );
  XOR U988 ( .A(n3488), .B(n3506), .Z(n3497) );
  XOR U989 ( .A(n3849), .B(n3867), .Z(n3858) );
  XOR U990 ( .A(n4210), .B(n4228), .Z(n4219) );
  XOR U991 ( .A(n4571), .B(n4589), .Z(n4580) );
  XOR U992 ( .A(n4932), .B(n4950), .Z(n4941) );
  XOR U993 ( .A(n5293), .B(n5311), .Z(n5302) );
  AND U994 ( .A(n965), .B(n964), .Z(n782) );
  AND U995 ( .A(n1692), .B(n1691), .Z(n1509) );
  AND U996 ( .A(n2416), .B(n2415), .Z(n2234) );
  AND U997 ( .A(n3138), .B(n3137), .Z(n2956) );
  AND U998 ( .A(n3860), .B(n3859), .Z(n3678) );
  AND U999 ( .A(n4582), .B(n4581), .Z(n4400) );
  AND U1000 ( .A(n5304), .B(n5303), .Z(n5122) );
  XOR U1001 ( .A(n6070), .B(n6235), .Z(n6074) );
  XOR U1002 ( .A(n5717), .B(n5882), .Z(n5721) );
  XOR U1003 ( .A(n1743), .B(n1906), .Z(n1747) );
  XOR U1004 ( .A(n2104), .B(n2267), .Z(n2108) );
  XOR U1005 ( .A(n2465), .B(n2628), .Z(n2469) );
  XOR U1006 ( .A(n2826), .B(n2989), .Z(n2830) );
  XOR U1007 ( .A(n3187), .B(n3350), .Z(n3191) );
  XOR U1008 ( .A(n3548), .B(n3711), .Z(n3552) );
  XOR U1009 ( .A(n3909), .B(n4072), .Z(n3913) );
  XOR U1010 ( .A(n4270), .B(n4433), .Z(n4274) );
  XOR U1011 ( .A(n4631), .B(n4794), .Z(n4635) );
  XOR U1012 ( .A(n4992), .B(n5155), .Z(n4996) );
  XOR U1013 ( .A(n5353), .B(n5516), .Z(n5357) );
  XOR U1014 ( .A(n1373), .B(n1544), .Z(n1378) );
  XOR U1015 ( .A(n6411), .B(n6558), .Z(n6415) );
  XOR U1016 ( .A(n6085), .B(n6232), .Z(n6089) );
  XOR U1017 ( .A(n5732), .B(n5879), .Z(n5736) );
  XOR U1018 ( .A(n1758), .B(n1903), .Z(n1762) );
  XOR U1019 ( .A(n2119), .B(n2264), .Z(n2123) );
  XOR U1020 ( .A(n2480), .B(n2625), .Z(n2484) );
  XOR U1021 ( .A(n2841), .B(n2986), .Z(n2845) );
  XOR U1022 ( .A(n3202), .B(n3347), .Z(n3206) );
  XOR U1023 ( .A(n3563), .B(n3708), .Z(n3567) );
  XOR U1024 ( .A(n3924), .B(n4069), .Z(n3928) );
  XOR U1025 ( .A(n4285), .B(n4430), .Z(n4289) );
  XOR U1026 ( .A(n4646), .B(n4791), .Z(n4650) );
  XOR U1027 ( .A(n5007), .B(n5152), .Z(n5011) );
  XOR U1028 ( .A(n5368), .B(n5513), .Z(n5372) );
  XOR U1029 ( .A(n1198), .B(n1361), .Z(n1202) );
  XOR U1030 ( .A(n7006), .B(n7135), .Z(n7010) );
  XOR U1031 ( .A(n6728), .B(n6857), .Z(n6732) );
  XOR U1032 ( .A(n6426), .B(n6555), .Z(n6430) );
  XOR U1033 ( .A(n6100), .B(n6229), .Z(n6104) );
  XOR U1034 ( .A(n5747), .B(n5876), .Z(n5751) );
  XOR U1035 ( .A(n1773), .B(n1900), .Z(n1777) );
  XOR U1036 ( .A(n2134), .B(n2261), .Z(n2138) );
  XOR U1037 ( .A(n2495), .B(n2622), .Z(n2499) );
  XOR U1038 ( .A(n2856), .B(n2983), .Z(n2860) );
  XOR U1039 ( .A(n3217), .B(n3344), .Z(n3221) );
  XOR U1040 ( .A(n3578), .B(n3705), .Z(n3582) );
  XOR U1041 ( .A(n3939), .B(n4066), .Z(n3943) );
  XOR U1042 ( .A(n4300), .B(n4427), .Z(n4304) );
  XOR U1043 ( .A(n4661), .B(n4788), .Z(n4665) );
  XOR U1044 ( .A(n5022), .B(n5149), .Z(n5026) );
  XOR U1045 ( .A(n5383), .B(n5510), .Z(n5387) );
  XOR U1046 ( .A(n1213), .B(n1358), .Z(n1217) );
  XOR U1047 ( .A(n828), .B(n999), .Z(n833) );
  XOR U1048 ( .A(n7275), .B(n7386), .Z(n7279) );
  XOR U1049 ( .A(n7021), .B(n7132), .Z(n7025) );
  XOR U1050 ( .A(n6743), .B(n6854), .Z(n6747) );
  XOR U1051 ( .A(n6441), .B(n6552), .Z(n6445) );
  XOR U1052 ( .A(n6115), .B(n6226), .Z(n6119) );
  XOR U1053 ( .A(n5762), .B(n5873), .Z(n5766) );
  XOR U1054 ( .A(n1788), .B(n1897), .Z(n1792) );
  XOR U1055 ( .A(n2149), .B(n2258), .Z(n2153) );
  XOR U1056 ( .A(n2510), .B(n2619), .Z(n2514) );
  XOR U1057 ( .A(n2871), .B(n2980), .Z(n2875) );
  XOR U1058 ( .A(n3232), .B(n3341), .Z(n3236) );
  XOR U1059 ( .A(n3593), .B(n3702), .Z(n3597) );
  XOR U1060 ( .A(n3954), .B(n4063), .Z(n3958) );
  XOR U1061 ( .A(n4315), .B(n4424), .Z(n4319) );
  XOR U1062 ( .A(n4676), .B(n4785), .Z(n4680) );
  XOR U1063 ( .A(n5037), .B(n5146), .Z(n5041) );
  XOR U1064 ( .A(n5398), .B(n5507), .Z(n5402) );
  XOR U1065 ( .A(n1419), .B(n1534), .Z(n1423) );
  XOR U1066 ( .A(n1036), .B(n1176), .Z(n1040) );
  XOR U1067 ( .A(n652), .B(n816), .Z(n656) );
  XOR U1068 ( .A(n7726), .B(n7819), .Z(n7730) );
  XOR U1069 ( .A(n7520), .B(n7613), .Z(n7524) );
  XOR U1070 ( .A(n7290), .B(n7383), .Z(n7294) );
  XOR U1071 ( .A(n7036), .B(n7129), .Z(n7040) );
  XOR U1072 ( .A(n6758), .B(n6851), .Z(n6762) );
  XOR U1073 ( .A(n6456), .B(n6549), .Z(n6460) );
  XOR U1074 ( .A(n6130), .B(n6223), .Z(n6134) );
  XOR U1075 ( .A(n5777), .B(n5870), .Z(n5781) );
  XOR U1076 ( .A(n879), .B(n989), .Z(n883) );
  XOR U1077 ( .A(n1439), .B(n1530), .Z(n1443) );
  XOR U1078 ( .A(n1803), .B(n1894), .Z(n1807) );
  XOR U1079 ( .A(n2164), .B(n2255), .Z(n2168) );
  XOR U1080 ( .A(n2525), .B(n2616), .Z(n2529) );
  XOR U1081 ( .A(n2886), .B(n2977), .Z(n2890) );
  XOR U1082 ( .A(n3247), .B(n3338), .Z(n3251) );
  XOR U1083 ( .A(n3608), .B(n3699), .Z(n3612) );
  XOR U1084 ( .A(n3969), .B(n4060), .Z(n3973) );
  XOR U1085 ( .A(n4330), .B(n4421), .Z(n4334) );
  XOR U1086 ( .A(n4691), .B(n4782), .Z(n4695) );
  XOR U1087 ( .A(n5052), .B(n5143), .Z(n5056) );
  XOR U1088 ( .A(n5413), .B(n5504), .Z(n5417) );
  XOR U1089 ( .A(n1051), .B(n1173), .Z(n1055) );
  XOR U1090 ( .A(n667), .B(n813), .Z(n671) );
  XOR U1091 ( .A(n285), .B(n454), .Z(n290) );
  XOR U1092 ( .A(n7923), .B(n7998), .Z(n7927) );
  XOR U1093 ( .A(n7741), .B(n7816), .Z(n7745) );
  XOR U1094 ( .A(n7535), .B(n7610), .Z(n7539) );
  XOR U1095 ( .A(n7305), .B(n7380), .Z(n7309) );
  XOR U1096 ( .A(n7051), .B(n7126), .Z(n7055) );
  XOR U1097 ( .A(n6773), .B(n6848), .Z(n6777) );
  XOR U1098 ( .A(n6471), .B(n6546), .Z(n6475) );
  XOR U1099 ( .A(n6145), .B(n6220), .Z(n6149) );
  XOR U1100 ( .A(n5792), .B(n5867), .Z(n5796) );
  XOR U1101 ( .A(n702), .B(n806), .Z(n706) );
  XOR U1102 ( .A(n321), .B(n447), .Z(n325) );
  XOR U1103 ( .A(n1091), .B(n1164), .Z(n1095) );
  XOR U1104 ( .A(n1454), .B(n1527), .Z(n1458) );
  XOR U1105 ( .A(n1818), .B(n1891), .Z(n1822) );
  XOR U1106 ( .A(n2179), .B(n2252), .Z(n2183) );
  XOR U1107 ( .A(n2540), .B(n2613), .Z(n2544) );
  XOR U1108 ( .A(n2901), .B(n2974), .Z(n2905) );
  XOR U1109 ( .A(n3262), .B(n3335), .Z(n3266) );
  XOR U1110 ( .A(n3623), .B(n3696), .Z(n3627) );
  XOR U1111 ( .A(n3984), .B(n4057), .Z(n3988) );
  XOR U1112 ( .A(n4345), .B(n4418), .Z(n4349) );
  XOR U1113 ( .A(n4706), .B(n4779), .Z(n4710) );
  XOR U1114 ( .A(n5067), .B(n5140), .Z(n5071) );
  XOR U1115 ( .A(n5428), .B(n5501), .Z(n5432) );
  XOR U1116 ( .A(n682), .B(n810), .Z(n686) );
  XOR U1117 ( .A(n301), .B(n451), .Z(n305) );
  XOR U1118 ( .A(n727), .B(n800), .Z(n731) );
  XOR U1119 ( .A(n351), .B(n441), .Z(n355) );
  XOR U1120 ( .A(n8230), .B(n8287), .Z(n8234) );
  XOR U1121 ( .A(n8096), .B(n8153), .Z(n8100) );
  XOR U1122 ( .A(n7938), .B(n7995), .Z(n7942) );
  XOR U1123 ( .A(n7756), .B(n7813), .Z(n7760) );
  XOR U1124 ( .A(n7550), .B(n7607), .Z(n7554) );
  XOR U1125 ( .A(n7320), .B(n7377), .Z(n7324) );
  XOR U1126 ( .A(n7066), .B(n7123), .Z(n7070) );
  XOR U1127 ( .A(n6788), .B(n6845), .Z(n6792) );
  XOR U1128 ( .A(n6486), .B(n6543), .Z(n6490) );
  XOR U1129 ( .A(n6160), .B(n6217), .Z(n6164) );
  XOR U1130 ( .A(n5807), .B(n5864), .Z(n5811) );
  XOR U1131 ( .A(n336), .B(n444), .Z(n340) );
  XOR U1132 ( .A(n381), .B(n435), .Z(n385) );
  XOR U1133 ( .A(n742), .B(n797), .Z(n746) );
  XOR U1134 ( .A(n1106), .B(n1161), .Z(n1110) );
  XOR U1135 ( .A(n1469), .B(n1524), .Z(n1473) );
  XOR U1136 ( .A(n1833), .B(n1888), .Z(n1837) );
  XOR U1137 ( .A(n2194), .B(n2249), .Z(n2198) );
  XOR U1138 ( .A(n2555), .B(n2610), .Z(n2559) );
  XOR U1139 ( .A(n2916), .B(n2971), .Z(n2920) );
  XOR U1140 ( .A(n3277), .B(n3332), .Z(n3281) );
  XOR U1141 ( .A(n3638), .B(n3693), .Z(n3642) );
  XOR U1142 ( .A(n3999), .B(n4054), .Z(n4003) );
  XOR U1143 ( .A(n4360), .B(n4415), .Z(n4364) );
  XOR U1144 ( .A(n4721), .B(n4776), .Z(n4725) );
  XOR U1145 ( .A(n5082), .B(n5137), .Z(n5086) );
  XOR U1146 ( .A(n5443), .B(n5498), .Z(n5447) );
  XOR U1147 ( .A(n114), .B(n258), .Z(n126) );
  XOR U1148 ( .A(n366), .B(n438), .Z(n370) );
  XOR U1149 ( .A(n8355), .B(n8394), .Z(n8359) );
  XOR U1150 ( .A(n8245), .B(n8284), .Z(n8249) );
  XOR U1151 ( .A(n8111), .B(n8150), .Z(n8115) );
  XOR U1152 ( .A(n7953), .B(n7992), .Z(n7957) );
  XOR U1153 ( .A(n7771), .B(n7810), .Z(n7775) );
  XOR U1154 ( .A(n7565), .B(n7604), .Z(n7569) );
  XOR U1155 ( .A(n7335), .B(n7374), .Z(n7339) );
  XOR U1156 ( .A(n7081), .B(n7120), .Z(n7085) );
  XOR U1157 ( .A(n6803), .B(n6842), .Z(n6807) );
  XOR U1158 ( .A(n6501), .B(n6540), .Z(n6505) );
  XOR U1159 ( .A(n6175), .B(n6214), .Z(n6179) );
  XOR U1160 ( .A(n5822), .B(n5861), .Z(n5826) );
  XOR U1161 ( .A(n396), .B(n432), .Z(n400) );
  XOR U1162 ( .A(n757), .B(n794), .Z(n761) );
  XOR U1163 ( .A(n1121), .B(n1158), .Z(n1125) );
  XOR U1164 ( .A(n1484), .B(n1521), .Z(n1488) );
  XOR U1165 ( .A(n1848), .B(n1885), .Z(n1852) );
  XOR U1166 ( .A(n2209), .B(n2246), .Z(n2213) );
  XOR U1167 ( .A(n2570), .B(n2607), .Z(n2574) );
  XOR U1168 ( .A(n2931), .B(n2968), .Z(n2935) );
  XOR U1169 ( .A(n3292), .B(n3329), .Z(n3296) );
  XOR U1170 ( .A(n3653), .B(n3690), .Z(n3657) );
  XOR U1171 ( .A(n4014), .B(n4051), .Z(n4018) );
  XOR U1172 ( .A(n4375), .B(n4412), .Z(n4379) );
  XOR U1173 ( .A(n4736), .B(n4773), .Z(n4740) );
  XOR U1174 ( .A(n5097), .B(n5134), .Z(n5101) );
  XOR U1175 ( .A(n5458), .B(n5495), .Z(n5462) );
  XOR U1176 ( .A(n8518), .B(n8539), .Z(n8527) );
  XOR U1177 ( .A(n8456), .B(n8477), .Z(n8465) );
  XOR U1178 ( .A(n8370), .B(n8391), .Z(n8379) );
  XOR U1179 ( .A(n8260), .B(n8281), .Z(n8269) );
  XOR U1180 ( .A(n8126), .B(n8147), .Z(n8135) );
  XOR U1181 ( .A(n7968), .B(n7989), .Z(n7977) );
  XOR U1182 ( .A(n7786), .B(n7807), .Z(n7795) );
  XOR U1183 ( .A(n7580), .B(n7601), .Z(n7589) );
  XOR U1184 ( .A(n7350), .B(n7371), .Z(n7359) );
  XOR U1185 ( .A(n7096), .B(n7117), .Z(n7105) );
  XOR U1186 ( .A(n6818), .B(n6839), .Z(n6827) );
  XOR U1187 ( .A(n6516), .B(n6537), .Z(n6525) );
  XOR U1188 ( .A(n6190), .B(n6211), .Z(n6199) );
  XOR U1189 ( .A(n5837), .B(n5858), .Z(n5846) );
  XOR U1190 ( .A(n411), .B(n429), .Z(n420) );
  XOR U1191 ( .A(n772), .B(n791), .Z(n781) );
  XOR U1192 ( .A(n1136), .B(n1155), .Z(n1145) );
  XOR U1193 ( .A(n1499), .B(n1518), .Z(n1508) );
  XOR U1194 ( .A(n1863), .B(n1882), .Z(n1872) );
  XOR U1195 ( .A(n2224), .B(n2243), .Z(n2233) );
  XOR U1196 ( .A(n2585), .B(n2604), .Z(n2594) );
  XOR U1197 ( .A(n2946), .B(n2965), .Z(n2955) );
  XOR U1198 ( .A(n3307), .B(n3326), .Z(n3316) );
  XOR U1199 ( .A(n3668), .B(n3687), .Z(n3677) );
  XOR U1200 ( .A(n4029), .B(n4048), .Z(n4038) );
  XOR U1201 ( .A(n4390), .B(n4409), .Z(n4399) );
  XOR U1202 ( .A(n4751), .B(n4770), .Z(n4760) );
  XOR U1203 ( .A(n5112), .B(n5131), .Z(n5121) );
  XOR U1204 ( .A(n5473), .B(n5492), .Z(n5482) );
  AND U1205 ( .A(n1147), .B(n1146), .Z(n964) );
  AND U1206 ( .A(n1874), .B(n1873), .Z(n1691) );
  AND U1207 ( .A(n2596), .B(n2595), .Z(n2415) );
  AND U1208 ( .A(n3318), .B(n3317), .Z(n3137) );
  AND U1209 ( .A(n4040), .B(n4039), .Z(n3859) );
  AND U1210 ( .A(n4762), .B(n4761), .Z(n4581) );
  ANDN U1211 ( .B(n5483), .A(n5485), .Z(n5303) );
  NAND U1212 ( .A(n422), .B(n421), .Z(n175) );
  XOR U1213 ( .A(n1), .B(n2), .Z(swire[63]) );
  XOR U1214 ( .A(n3), .B(n4), .Z(n2) );
  XOR U1215 ( .A(n5), .B(n6), .Z(n4) );
  XOR U1216 ( .A(n7), .B(n8), .Z(n6) );
  XOR U1217 ( .A(n9), .B(n10), .Z(n8) );
  XNOR U1218 ( .A(n11), .B(n12), .Z(n10) );
  AND U1219 ( .A(a[62]), .B(b[1]), .Z(n12) );
  XOR U1220 ( .A(n13), .B(n14), .Z(n9) );
  XOR U1221 ( .A(n15), .B(n16), .Z(n14) );
  XOR U1222 ( .A(n17), .B(n18), .Z(n16) );
  AND U1223 ( .A(a[56]), .B(b[7]), .Z(n18) );
  AND U1224 ( .A(b[8]), .B(a[55]), .Z(n17) );
  XOR U1225 ( .A(n19), .B(n20), .Z(n15) );
  XOR U1226 ( .A(n21), .B(n22), .Z(n20) );
  XOR U1227 ( .A(n23), .B(n24), .Z(n22) );
  XOR U1228 ( .A(n25), .B(n26), .Z(n24) );
  XOR U1229 ( .A(n27), .B(n28), .Z(n26) );
  XOR U1230 ( .A(n29), .B(n30), .Z(n28) );
  AND U1231 ( .A(b[20]), .B(a[43]), .Z(n30) );
  AND U1232 ( .A(a[38]), .B(b[25]), .Z(n29) );
  XOR U1233 ( .A(n31), .B(n32), .Z(n27) );
  AND U1234 ( .A(b[26]), .B(a[37]), .Z(n32) );
  AND U1235 ( .A(a[36]), .B(b[27]), .Z(n31) );
  XOR U1236 ( .A(n33), .B(n34), .Z(n25) );
  XOR U1237 ( .A(n35), .B(n36), .Z(n34) );
  AND U1238 ( .A(b[28]), .B(a[35]), .Z(n36) );
  AND U1239 ( .A(a[34]), .B(b[29]), .Z(n35) );
  XOR U1240 ( .A(n37), .B(n38), .Z(n33) );
  AND U1241 ( .A(b[30]), .B(a[33]), .Z(n38) );
  AND U1242 ( .A(a[32]), .B(b[31]), .Z(n37) );
  AND U1243 ( .A(a[50]), .B(b[13]), .Z(n23) );
  XOR U1244 ( .A(n39), .B(n40), .Z(n21) );
  AND U1245 ( .A(b[14]), .B(a[49]), .Z(n40) );
  AND U1246 ( .A(a[44]), .B(b[19]), .Z(n39) );
  XOR U1247 ( .A(n41), .B(n42), .Z(n19) );
  XOR U1248 ( .A(n43), .B(n44), .Z(n42) );
  AND U1249 ( .A(a[42]), .B(b[21]), .Z(n44) );
  AND U1250 ( .A(b[22]), .B(a[41]), .Z(n43) );
  XOR U1251 ( .A(n45), .B(n46), .Z(n41) );
  AND U1252 ( .A(a[40]), .B(b[23]), .Z(n46) );
  AND U1253 ( .A(b[24]), .B(a[39]), .Z(n45) );
  XOR U1254 ( .A(n47), .B(n48), .Z(n13) );
  XOR U1255 ( .A(n49), .B(n50), .Z(n48) );
  AND U1256 ( .A(a[48]), .B(b[15]), .Z(n50) );
  AND U1257 ( .A(b[16]), .B(a[47]), .Z(n49) );
  XOR U1258 ( .A(n51), .B(n52), .Z(n47) );
  AND U1259 ( .A(a[46]), .B(b[17]), .Z(n52) );
  AND U1260 ( .A(b[18]), .B(a[45]), .Z(n51) );
  XOR U1261 ( .A(n53), .B(n54), .Z(n7) );
  XOR U1262 ( .A(n55), .B(n56), .Z(n54) );
  AND U1263 ( .A(a[54]), .B(b[9]), .Z(n56) );
  AND U1264 ( .A(b[10]), .B(a[53]), .Z(n55) );
  XOR U1265 ( .A(n57), .B(n58), .Z(n53) );
  AND U1266 ( .A(a[52]), .B(b[11]), .Z(n58) );
  AND U1267 ( .A(b[12]), .B(a[51]), .Z(n57) );
  AND U1268 ( .A(a[63]), .B(b[0]), .Z(n5) );
  XNOR U1269 ( .A(n59), .B(n11), .Z(n3) );
  OR U1270 ( .A(n60), .B(n61), .Z(n11) );
  AND U1271 ( .A(a[61]), .B(b[2]), .Z(n59) );
  XOR U1272 ( .A(n62), .B(n63), .Z(n1) );
  XOR U1273 ( .A(n64), .B(n65), .Z(n63) );
  AND U1274 ( .A(a[60]), .B(b[3]), .Z(n65) );
  AND U1275 ( .A(a[59]), .B(b[4]), .Z(n64) );
  XOR U1276 ( .A(n66), .B(n67), .Z(n62) );
  AND U1277 ( .A(a[58]), .B(b[5]), .Z(n67) );
  AND U1278 ( .A(a[57]), .B(b[6]), .Z(n66) );
  XOR U1279 ( .A(n60), .B(n61), .Z(swire[62]) );
  XOR U1280 ( .A(n68), .B(n69), .Z(n61) );
  XNOR U1281 ( .A(n70), .B(n71), .Z(n69) );
  XOR U1282 ( .A(n72), .B(n73), .Z(n71) );
  XOR U1283 ( .A(n74), .B(n75), .Z(n73) );
  XNOR U1284 ( .A(n76), .B(n70), .Z(n75) );
  XOR U1285 ( .A(n77), .B(n78), .Z(n74) );
  XOR U1286 ( .A(n79), .B(n80), .Z(n78) );
  XOR U1287 ( .A(n81), .B(n82), .Z(n80) );
  XOR U1288 ( .A(n83), .B(n84), .Z(n82) );
  AND U1289 ( .A(b[7]), .B(a[55]), .Z(n83) );
  XOR U1290 ( .A(n85), .B(n86), .Z(n81) );
  XOR U1291 ( .A(n87), .B(n88), .Z(n86) );
  XOR U1292 ( .A(n89), .B(n90), .Z(n88) );
  XOR U1293 ( .A(n91), .B(n92), .Z(n90) );
  AND U1294 ( .A(b[13]), .B(a[49]), .Z(n91) );
  XOR U1295 ( .A(n93), .B(n94), .Z(n89) );
  XOR U1296 ( .A(n95), .B(n96), .Z(n94) );
  XOR U1297 ( .A(n97), .B(n98), .Z(n96) );
  XOR U1298 ( .A(n99), .B(n100), .Z(n98) );
  AND U1299 ( .A(b[19]), .B(a[43]), .Z(n99) );
  XOR U1300 ( .A(n101), .B(n102), .Z(n97) );
  AND U1301 ( .A(a[38]), .B(b[24]), .Z(n101) );
  XOR U1302 ( .A(n100), .B(n103), .Z(n95) );
  XOR U1303 ( .A(n102), .B(n104), .Z(n103) );
  XOR U1304 ( .A(n105), .B(n106), .Z(n104) );
  XOR U1305 ( .A(n107), .B(n108), .Z(n106) );
  XOR U1306 ( .A(n109), .B(n110), .Z(n108) );
  XOR U1307 ( .A(n111), .B(n109), .Z(n110) );
  AND U1308 ( .A(b[25]), .B(a[37]), .Z(n111) );
  XOR U1309 ( .A(n112), .B(n113), .Z(n109) );
  NOR U1310 ( .A(n114), .B(n115), .Z(n112) );
  XOR U1311 ( .A(n116), .B(n117), .Z(n107) );
  AND U1312 ( .A(a[36]), .B(b[26]), .Z(n117) );
  AND U1313 ( .A(b[27]), .B(a[35]), .Z(n116) );
  XOR U1314 ( .A(n118), .B(n119), .Z(n105) );
  XOR U1315 ( .A(n120), .B(n121), .Z(n119) );
  AND U1316 ( .A(a[34]), .B(b[28]), .Z(n121) );
  AND U1317 ( .A(b[29]), .B(a[33]), .Z(n120) );
  XOR U1318 ( .A(n122), .B(n123), .Z(n118) );
  AND U1319 ( .A(a[32]), .B(b[30]), .Z(n123) );
  AND U1320 ( .A(b[31]), .B(a[31]), .Z(n122) );
  XOR U1321 ( .A(n124), .B(n125), .Z(n102) );
  AND U1322 ( .A(n126), .B(n127), .Z(n124) );
  XOR U1323 ( .A(n128), .B(n129), .Z(n100) );
  ANDN U1324 ( .B(n130), .A(n131), .Z(n128) );
  XOR U1325 ( .A(n132), .B(n133), .Z(n93) );
  XOR U1326 ( .A(n134), .B(n135), .Z(n133) );
  AND U1327 ( .A(a[42]), .B(b[20]), .Z(n135) );
  AND U1328 ( .A(b[21]), .B(a[41]), .Z(n134) );
  XOR U1329 ( .A(n136), .B(n137), .Z(n132) );
  AND U1330 ( .A(a[40]), .B(b[22]), .Z(n137) );
  AND U1331 ( .A(b[23]), .B(a[39]), .Z(n136) );
  XOR U1332 ( .A(n138), .B(n92), .Z(n87) );
  XOR U1333 ( .A(n139), .B(n140), .Z(n92) );
  ANDN U1334 ( .B(n141), .A(n142), .Z(n139) );
  AND U1335 ( .A(a[48]), .B(b[14]), .Z(n138) );
  XOR U1336 ( .A(n143), .B(n144), .Z(n85) );
  XOR U1337 ( .A(n145), .B(n146), .Z(n144) );
  AND U1338 ( .A(b[15]), .B(a[47]), .Z(n146) );
  AND U1339 ( .A(a[46]), .B(b[16]), .Z(n145) );
  XOR U1340 ( .A(n147), .B(n148), .Z(n143) );
  AND U1341 ( .A(b[17]), .B(a[45]), .Z(n148) );
  AND U1342 ( .A(a[44]), .B(b[18]), .Z(n147) );
  XOR U1343 ( .A(n149), .B(n84), .Z(n79) );
  XOR U1344 ( .A(n150), .B(n151), .Z(n84) );
  ANDN U1345 ( .B(n152), .A(n153), .Z(n150) );
  AND U1346 ( .A(a[54]), .B(b[8]), .Z(n149) );
  XOR U1347 ( .A(n154), .B(n155), .Z(n77) );
  XOR U1348 ( .A(n156), .B(n157), .Z(n155) );
  AND U1349 ( .A(b[9]), .B(a[53]), .Z(n157) );
  AND U1350 ( .A(a[52]), .B(b[10]), .Z(n156) );
  XOR U1351 ( .A(n158), .B(n159), .Z(n154) );
  AND U1352 ( .A(b[11]), .B(a[51]), .Z(n159) );
  AND U1353 ( .A(a[50]), .B(b[12]), .Z(n158) );
  XOR U1354 ( .A(n160), .B(n161), .Z(n72) );
  XOR U1355 ( .A(n162), .B(n163), .Z(n161) );
  AND U1356 ( .A(a[59]), .B(b[3]), .Z(n163) );
  AND U1357 ( .A(a[58]), .B(b[4]), .Z(n162) );
  XOR U1358 ( .A(n164), .B(n165), .Z(n160) );
  AND U1359 ( .A(a[57]), .B(b[5]), .Z(n165) );
  AND U1360 ( .A(b[6]), .B(a[56]), .Z(n164) );
  XOR U1361 ( .A(n166), .B(n167), .Z(n70) );
  OR U1362 ( .A(n168), .B(n169), .Z(n167) );
  XOR U1363 ( .A(n170), .B(n171), .Z(n68) );
  XNOR U1364 ( .A(n172), .B(n76), .Z(n171) );
  NANDN U1365 ( .A(n173), .B(n174), .Z(n76) );
  AND U1366 ( .A(a[60]), .B(b[2]), .Z(n172) );
  AND U1367 ( .A(a[61]), .B(b[1]), .Z(n170) );
  NAND U1368 ( .A(a[62]), .B(b[0]), .Z(n60) );
  XNOR U1369 ( .A(n175), .B(n176), .Z(swire[61]) );
  XOR U1370 ( .A(n174), .B(n177), .Z(n176) );
  XOR U1371 ( .A(n173), .B(n175), .Z(n177) );
  NAND U1372 ( .A(a[61]), .B(b[0]), .Z(n173) );
  XOR U1373 ( .A(n168), .B(n169), .Z(n174) );
  XOR U1374 ( .A(n166), .B(n178), .Z(n169) );
  NAND U1375 ( .A(a[60]), .B(b[1]), .Z(n178) );
  XOR U1376 ( .A(n179), .B(n180), .Z(n168) );
  XOR U1377 ( .A(n166), .B(n181), .Z(n180) );
  XOR U1378 ( .A(n182), .B(n183), .Z(n181) );
  AND U1379 ( .A(a[59]), .B(b[2]), .Z(n182) );
  ANDN U1380 ( .B(n184), .A(n185), .Z(n166) );
  XOR U1381 ( .A(n186), .B(n187), .Z(n179) );
  XNOR U1382 ( .A(n183), .B(n188), .Z(n187) );
  XOR U1383 ( .A(n189), .B(n190), .Z(n188) );
  XOR U1384 ( .A(n191), .B(n192), .Z(n190) );
  XOR U1385 ( .A(n193), .B(n194), .Z(n192) );
  XOR U1386 ( .A(n195), .B(n196), .Z(n194) );
  XOR U1387 ( .A(n152), .B(n197), .Z(n196) );
  XNOR U1388 ( .A(n198), .B(n153), .Z(n197) );
  XOR U1389 ( .A(n199), .B(n200), .Z(n153) );
  XOR U1390 ( .A(n151), .B(n201), .Z(n200) );
  XOR U1391 ( .A(n202), .B(n203), .Z(n201) );
  XOR U1392 ( .A(n204), .B(n205), .Z(n203) );
  XOR U1393 ( .A(n206), .B(n207), .Z(n205) );
  XOR U1394 ( .A(n208), .B(n209), .Z(n207) );
  XOR U1395 ( .A(n210), .B(n211), .Z(n209) );
  XOR U1396 ( .A(n212), .B(n213), .Z(n211) );
  XOR U1397 ( .A(n214), .B(n215), .Z(n213) );
  XOR U1398 ( .A(n216), .B(n217), .Z(n215) );
  XOR U1399 ( .A(n141), .B(n218), .Z(n217) );
  XOR U1400 ( .A(n219), .B(n142), .Z(n218) );
  XOR U1401 ( .A(n220), .B(n221), .Z(n142) );
  XOR U1402 ( .A(n140), .B(n222), .Z(n221) );
  XOR U1403 ( .A(n223), .B(n224), .Z(n222) );
  XOR U1404 ( .A(n225), .B(n226), .Z(n224) );
  XOR U1405 ( .A(n227), .B(n228), .Z(n226) );
  XOR U1406 ( .A(n229), .B(n230), .Z(n228) );
  XOR U1407 ( .A(n231), .B(n232), .Z(n230) );
  XOR U1408 ( .A(n233), .B(n234), .Z(n232) );
  XOR U1409 ( .A(n235), .B(n236), .Z(n234) );
  XOR U1410 ( .A(n237), .B(n238), .Z(n236) );
  XOR U1411 ( .A(n130), .B(n239), .Z(n238) );
  XOR U1412 ( .A(n240), .B(n131), .Z(n239) );
  XOR U1413 ( .A(n241), .B(n242), .Z(n131) );
  XOR U1414 ( .A(n129), .B(n243), .Z(n242) );
  XOR U1415 ( .A(n244), .B(n245), .Z(n243) );
  XOR U1416 ( .A(n246), .B(n247), .Z(n245) );
  XOR U1417 ( .A(n248), .B(n249), .Z(n247) );
  XOR U1418 ( .A(n250), .B(n251), .Z(n249) );
  XOR U1419 ( .A(n252), .B(n253), .Z(n251) );
  XOR U1420 ( .A(n254), .B(n255), .Z(n253) );
  XOR U1421 ( .A(n127), .B(n256), .Z(n255) );
  XNOR U1422 ( .A(n257), .B(n126), .Z(n256) );
  XOR U1423 ( .A(n125), .B(n115), .Z(n258) );
  XOR U1424 ( .A(n259), .B(n260), .Z(n115) );
  XOR U1425 ( .A(n113), .B(n261), .Z(n260) );
  XOR U1426 ( .A(n262), .B(n263), .Z(n261) );
  XOR U1427 ( .A(n264), .B(n265), .Z(n263) );
  XOR U1428 ( .A(n266), .B(n267), .Z(n265) );
  XOR U1429 ( .A(n268), .B(n269), .Z(n267) );
  XOR U1430 ( .A(n270), .B(n271), .Z(n269) );
  XOR U1431 ( .A(n272), .B(n273), .Z(n271) );
  XOR U1432 ( .A(n274), .B(n275), .Z(n273) );
  XOR U1433 ( .A(n276), .B(n277), .Z(n275) );
  XOR U1434 ( .A(n278), .B(n279), .Z(n277) );
  XOR U1435 ( .A(n280), .B(n281), .Z(n279) );
  NAND U1436 ( .A(b[30]), .B(a[31]), .Z(n281) );
  AND U1437 ( .A(a[30]), .B(b[31]), .Z(n280) );
  XOR U1438 ( .A(n282), .B(n278), .Z(n274) );
  XOR U1439 ( .A(n283), .B(n284), .Z(n278) );
  NOR U1440 ( .A(n285), .B(n286), .Z(n283) );
  AND U1441 ( .A(a[32]), .B(b[29]), .Z(n282) );
  XOR U1442 ( .A(n287), .B(n276), .Z(n270) );
  XOR U1443 ( .A(n288), .B(n289), .Z(n276) );
  ANDN U1444 ( .B(n290), .A(n291), .Z(n288) );
  AND U1445 ( .A(b[28]), .B(a[33]), .Z(n287) );
  XOR U1446 ( .A(n292), .B(n272), .Z(n266) );
  XOR U1447 ( .A(n293), .B(n294), .Z(n272) );
  ANDN U1448 ( .B(n295), .A(n296), .Z(n293) );
  AND U1449 ( .A(a[34]), .B(b[27]), .Z(n292) );
  XOR U1450 ( .A(n297), .B(n268), .Z(n262) );
  XOR U1451 ( .A(n298), .B(n299), .Z(n268) );
  ANDN U1452 ( .B(n300), .A(n301), .Z(n298) );
  AND U1453 ( .A(b[26]), .B(a[35]), .Z(n297) );
  XOR U1454 ( .A(n302), .B(n264), .Z(n259) );
  XOR U1455 ( .A(n303), .B(n304), .Z(n264) );
  ANDN U1456 ( .B(n305), .A(n306), .Z(n303) );
  AND U1457 ( .A(a[36]), .B(b[25]), .Z(n302) );
  XNOR U1458 ( .A(n307), .B(n113), .Z(n114) );
  XOR U1459 ( .A(n308), .B(n309), .Z(n113) );
  ANDN U1460 ( .B(n310), .A(n311), .Z(n308) );
  AND U1461 ( .A(b[24]), .B(a[37]), .Z(n307) );
  XOR U1462 ( .A(n312), .B(n125), .Z(n127) );
  XOR U1463 ( .A(n313), .B(n314), .Z(n125) );
  ANDN U1464 ( .B(n315), .A(n316), .Z(n313) );
  AND U1465 ( .A(a[38]), .B(b[23]), .Z(n312) );
  XOR U1466 ( .A(n317), .B(n257), .Z(n252) );
  XOR U1467 ( .A(n318), .B(n319), .Z(n257) );
  ANDN U1468 ( .B(n320), .A(n321), .Z(n318) );
  AND U1469 ( .A(b[22]), .B(a[39]), .Z(n317) );
  XOR U1470 ( .A(n322), .B(n254), .Z(n248) );
  XOR U1471 ( .A(n323), .B(n324), .Z(n254) );
  ANDN U1472 ( .B(n325), .A(n326), .Z(n323) );
  AND U1473 ( .A(a[40]), .B(b[21]), .Z(n322) );
  XOR U1474 ( .A(n327), .B(n250), .Z(n244) );
  XOR U1475 ( .A(n328), .B(n329), .Z(n250) );
  ANDN U1476 ( .B(n330), .A(n331), .Z(n328) );
  AND U1477 ( .A(b[20]), .B(a[41]), .Z(n327) );
  XOR U1478 ( .A(n332), .B(n246), .Z(n241) );
  XOR U1479 ( .A(n333), .B(n334), .Z(n246) );
  ANDN U1480 ( .B(n335), .A(n336), .Z(n333) );
  AND U1481 ( .A(a[42]), .B(b[19]), .Z(n332) );
  XOR U1482 ( .A(n337), .B(n129), .Z(n130) );
  XOR U1483 ( .A(n338), .B(n339), .Z(n129) );
  ANDN U1484 ( .B(n340), .A(n341), .Z(n338) );
  AND U1485 ( .A(b[18]), .B(a[43]), .Z(n337) );
  XOR U1486 ( .A(n342), .B(n240), .Z(n235) );
  XOR U1487 ( .A(n343), .B(n344), .Z(n240) );
  ANDN U1488 ( .B(n345), .A(n346), .Z(n343) );
  AND U1489 ( .A(a[44]), .B(b[17]), .Z(n342) );
  XOR U1490 ( .A(n347), .B(n237), .Z(n231) );
  XOR U1491 ( .A(n348), .B(n349), .Z(n237) );
  ANDN U1492 ( .B(n350), .A(n351), .Z(n348) );
  AND U1493 ( .A(b[16]), .B(a[45]), .Z(n347) );
  XOR U1494 ( .A(n352), .B(n233), .Z(n227) );
  XOR U1495 ( .A(n353), .B(n354), .Z(n233) );
  ANDN U1496 ( .B(n355), .A(n356), .Z(n353) );
  AND U1497 ( .A(a[46]), .B(b[15]), .Z(n352) );
  XOR U1498 ( .A(n357), .B(n229), .Z(n223) );
  XOR U1499 ( .A(n358), .B(n359), .Z(n229) );
  ANDN U1500 ( .B(n360), .A(n361), .Z(n358) );
  AND U1501 ( .A(b[14]), .B(a[47]), .Z(n357) );
  XOR U1502 ( .A(n362), .B(n225), .Z(n220) );
  XOR U1503 ( .A(n363), .B(n364), .Z(n225) );
  ANDN U1504 ( .B(n365), .A(n366), .Z(n363) );
  AND U1505 ( .A(a[48]), .B(b[13]), .Z(n362) );
  XOR U1506 ( .A(n367), .B(n140), .Z(n141) );
  XOR U1507 ( .A(n368), .B(n369), .Z(n140) );
  ANDN U1508 ( .B(n370), .A(n371), .Z(n368) );
  AND U1509 ( .A(b[12]), .B(a[49]), .Z(n367) );
  XOR U1510 ( .A(n372), .B(n219), .Z(n214) );
  XOR U1511 ( .A(n373), .B(n374), .Z(n219) );
  ANDN U1512 ( .B(n375), .A(n376), .Z(n373) );
  AND U1513 ( .A(a[50]), .B(b[11]), .Z(n372) );
  XOR U1514 ( .A(n377), .B(n216), .Z(n210) );
  XOR U1515 ( .A(n378), .B(n379), .Z(n216) );
  ANDN U1516 ( .B(n380), .A(n381), .Z(n378) );
  AND U1517 ( .A(b[10]), .B(a[51]), .Z(n377) );
  XOR U1518 ( .A(n382), .B(n212), .Z(n206) );
  XOR U1519 ( .A(n383), .B(n384), .Z(n212) );
  ANDN U1520 ( .B(n385), .A(n386), .Z(n383) );
  AND U1521 ( .A(a[52]), .B(b[9]), .Z(n382) );
  XOR U1522 ( .A(n387), .B(n208), .Z(n202) );
  XOR U1523 ( .A(n388), .B(n389), .Z(n208) );
  ANDN U1524 ( .B(n390), .A(n391), .Z(n388) );
  AND U1525 ( .A(b[8]), .B(a[53]), .Z(n387) );
  XOR U1526 ( .A(n392), .B(n204), .Z(n199) );
  XOR U1527 ( .A(n393), .B(n394), .Z(n204) );
  ANDN U1528 ( .B(n395), .A(n396), .Z(n393) );
  AND U1529 ( .A(a[54]), .B(b[7]), .Z(n392) );
  XOR U1530 ( .A(n397), .B(n151), .Z(n152) );
  XOR U1531 ( .A(n398), .B(n399), .Z(n151) );
  ANDN U1532 ( .B(n400), .A(n401), .Z(n398) );
  AND U1533 ( .A(b[6]), .B(a[55]), .Z(n397) );
  XOR U1534 ( .A(n402), .B(n198), .Z(n193) );
  XOR U1535 ( .A(n403), .B(n404), .Z(n198) );
  ANDN U1536 ( .B(n405), .A(n406), .Z(n403) );
  AND U1537 ( .A(b[5]), .B(a[56]), .Z(n402) );
  XOR U1538 ( .A(n407), .B(n195), .Z(n189) );
  XOR U1539 ( .A(n408), .B(n409), .Z(n195) );
  ANDN U1540 ( .B(n410), .A(n411), .Z(n408) );
  AND U1541 ( .A(a[57]), .B(b[4]), .Z(n407) );
  XNOR U1542 ( .A(n412), .B(n413), .Z(n183) );
  NANDN U1543 ( .A(n414), .B(n415), .Z(n413) );
  XOR U1544 ( .A(n416), .B(n191), .Z(n186) );
  XNOR U1545 ( .A(n417), .B(n418), .Z(n191) );
  AND U1546 ( .A(n419), .B(n420), .Z(n417) );
  AND U1547 ( .A(a[58]), .B(b[3]), .Z(n416) );
  XNOR U1548 ( .A(n421), .B(n422), .Z(swire[60]) );
  XOR U1549 ( .A(n184), .B(n423), .Z(n422) );
  XOR U1550 ( .A(n185), .B(n421), .Z(n423) );
  NAND U1551 ( .A(a[60]), .B(b[0]), .Z(n185) );
  XNOR U1552 ( .A(n414), .B(n415), .Z(n184) );
  XOR U1553 ( .A(n412), .B(n424), .Z(n415) );
  NAND U1554 ( .A(a[59]), .B(b[1]), .Z(n424) );
  XOR U1555 ( .A(n420), .B(n425), .Z(n414) );
  XOR U1556 ( .A(n412), .B(n419), .Z(n425) );
  XNOR U1557 ( .A(n426), .B(n418), .Z(n419) );
  AND U1558 ( .A(a[58]), .B(b[2]), .Z(n426) );
  NANDN U1559 ( .A(n427), .B(n428), .Z(n412) );
  XOR U1560 ( .A(n418), .B(n410), .Z(n429) );
  XNOR U1561 ( .A(n409), .B(n405), .Z(n430) );
  XNOR U1562 ( .A(n404), .B(n400), .Z(n431) );
  XNOR U1563 ( .A(n399), .B(n395), .Z(n432) );
  XNOR U1564 ( .A(n394), .B(n390), .Z(n433) );
  XNOR U1565 ( .A(n389), .B(n385), .Z(n434) );
  XNOR U1566 ( .A(n384), .B(n380), .Z(n435) );
  XNOR U1567 ( .A(n379), .B(n375), .Z(n436) );
  XNOR U1568 ( .A(n374), .B(n370), .Z(n437) );
  XNOR U1569 ( .A(n369), .B(n365), .Z(n438) );
  XNOR U1570 ( .A(n364), .B(n360), .Z(n439) );
  XNOR U1571 ( .A(n359), .B(n355), .Z(n440) );
  XNOR U1572 ( .A(n354), .B(n350), .Z(n441) );
  XNOR U1573 ( .A(n349), .B(n345), .Z(n442) );
  XNOR U1574 ( .A(n344), .B(n340), .Z(n443) );
  XNOR U1575 ( .A(n339), .B(n335), .Z(n444) );
  XNOR U1576 ( .A(n334), .B(n330), .Z(n445) );
  XNOR U1577 ( .A(n329), .B(n325), .Z(n446) );
  XNOR U1578 ( .A(n324), .B(n320), .Z(n447) );
  XNOR U1579 ( .A(n319), .B(n315), .Z(n448) );
  XNOR U1580 ( .A(n314), .B(n310), .Z(n449) );
  XNOR U1581 ( .A(n309), .B(n305), .Z(n450) );
  XNOR U1582 ( .A(n304), .B(n300), .Z(n451) );
  XNOR U1583 ( .A(n299), .B(n295), .Z(n452) );
  XNOR U1584 ( .A(n294), .B(n290), .Z(n453) );
  XOR U1585 ( .A(n289), .B(n286), .Z(n454) );
  XOR U1586 ( .A(n455), .B(n456), .Z(n286) );
  XOR U1587 ( .A(n284), .B(n457), .Z(n456) );
  XOR U1588 ( .A(n458), .B(n459), .Z(n457) );
  XOR U1589 ( .A(n460), .B(n461), .Z(n459) );
  NAND U1590 ( .A(a[30]), .B(b[30]), .Z(n461) );
  AND U1591 ( .A(a[29]), .B(b[31]), .Z(n460) );
  XOR U1592 ( .A(n462), .B(n458), .Z(n455) );
  XOR U1593 ( .A(n463), .B(n464), .Z(n458) );
  NOR U1594 ( .A(n465), .B(n466), .Z(n463) );
  AND U1595 ( .A(b[29]), .B(a[31]), .Z(n462) );
  XNOR U1596 ( .A(n467), .B(n284), .Z(n285) );
  XOR U1597 ( .A(n468), .B(n469), .Z(n284) );
  ANDN U1598 ( .B(n470), .A(n471), .Z(n468) );
  AND U1599 ( .A(a[32]), .B(b[28]), .Z(n467) );
  XNOR U1600 ( .A(n472), .B(n289), .Z(n291) );
  XOR U1601 ( .A(n473), .B(n474), .Z(n289) );
  ANDN U1602 ( .B(n475), .A(n476), .Z(n473) );
  AND U1603 ( .A(b[27]), .B(a[33]), .Z(n472) );
  XNOR U1604 ( .A(n477), .B(n294), .Z(n296) );
  XOR U1605 ( .A(n478), .B(n479), .Z(n294) );
  ANDN U1606 ( .B(n480), .A(n481), .Z(n478) );
  AND U1607 ( .A(a[34]), .B(b[26]), .Z(n477) );
  XNOR U1608 ( .A(n482), .B(n299), .Z(n301) );
  XOR U1609 ( .A(n483), .B(n484), .Z(n299) );
  ANDN U1610 ( .B(n485), .A(n486), .Z(n483) );
  AND U1611 ( .A(b[25]), .B(a[35]), .Z(n482) );
  XNOR U1612 ( .A(n487), .B(n304), .Z(n306) );
  XOR U1613 ( .A(n488), .B(n489), .Z(n304) );
  ANDN U1614 ( .B(n490), .A(n491), .Z(n488) );
  AND U1615 ( .A(a[36]), .B(b[24]), .Z(n487) );
  XNOR U1616 ( .A(n492), .B(n309), .Z(n311) );
  XOR U1617 ( .A(n493), .B(n494), .Z(n309) );
  ANDN U1618 ( .B(n495), .A(n496), .Z(n493) );
  AND U1619 ( .A(b[23]), .B(a[37]), .Z(n492) );
  XNOR U1620 ( .A(n497), .B(n314), .Z(n316) );
  XOR U1621 ( .A(n498), .B(n499), .Z(n314) );
  ANDN U1622 ( .B(n500), .A(n501), .Z(n498) );
  AND U1623 ( .A(a[38]), .B(b[22]), .Z(n497) );
  XNOR U1624 ( .A(n502), .B(n319), .Z(n321) );
  XOR U1625 ( .A(n503), .B(n504), .Z(n319) );
  ANDN U1626 ( .B(n505), .A(n506), .Z(n503) );
  AND U1627 ( .A(b[21]), .B(a[39]), .Z(n502) );
  XNOR U1628 ( .A(n507), .B(n324), .Z(n326) );
  XOR U1629 ( .A(n508), .B(n509), .Z(n324) );
  ANDN U1630 ( .B(n510), .A(n511), .Z(n508) );
  AND U1631 ( .A(a[40]), .B(b[20]), .Z(n507) );
  XNOR U1632 ( .A(n512), .B(n329), .Z(n331) );
  XOR U1633 ( .A(n513), .B(n514), .Z(n329) );
  ANDN U1634 ( .B(n515), .A(n516), .Z(n513) );
  AND U1635 ( .A(b[19]), .B(a[41]), .Z(n512) );
  XNOR U1636 ( .A(n517), .B(n334), .Z(n336) );
  XOR U1637 ( .A(n518), .B(n519), .Z(n334) );
  ANDN U1638 ( .B(n520), .A(n521), .Z(n518) );
  AND U1639 ( .A(a[42]), .B(b[18]), .Z(n517) );
  XNOR U1640 ( .A(n522), .B(n339), .Z(n341) );
  XOR U1641 ( .A(n523), .B(n524), .Z(n339) );
  ANDN U1642 ( .B(n525), .A(n526), .Z(n523) );
  AND U1643 ( .A(b[17]), .B(a[43]), .Z(n522) );
  XNOR U1644 ( .A(n527), .B(n344), .Z(n346) );
  XOR U1645 ( .A(n528), .B(n529), .Z(n344) );
  ANDN U1646 ( .B(n530), .A(n531), .Z(n528) );
  AND U1647 ( .A(a[44]), .B(b[16]), .Z(n527) );
  XNOR U1648 ( .A(n532), .B(n349), .Z(n351) );
  XOR U1649 ( .A(n533), .B(n534), .Z(n349) );
  ANDN U1650 ( .B(n535), .A(n536), .Z(n533) );
  AND U1651 ( .A(b[15]), .B(a[45]), .Z(n532) );
  XNOR U1652 ( .A(n537), .B(n354), .Z(n356) );
  XOR U1653 ( .A(n538), .B(n539), .Z(n354) );
  ANDN U1654 ( .B(n540), .A(n541), .Z(n538) );
  AND U1655 ( .A(a[46]), .B(b[14]), .Z(n537) );
  XNOR U1656 ( .A(n542), .B(n359), .Z(n361) );
  XOR U1657 ( .A(n543), .B(n544), .Z(n359) );
  ANDN U1658 ( .B(n545), .A(n546), .Z(n543) );
  AND U1659 ( .A(b[13]), .B(a[47]), .Z(n542) );
  XNOR U1660 ( .A(n547), .B(n364), .Z(n366) );
  XOR U1661 ( .A(n548), .B(n549), .Z(n364) );
  ANDN U1662 ( .B(n550), .A(n551), .Z(n548) );
  AND U1663 ( .A(a[48]), .B(b[12]), .Z(n547) );
  XNOR U1664 ( .A(n552), .B(n369), .Z(n371) );
  XOR U1665 ( .A(n553), .B(n554), .Z(n369) );
  ANDN U1666 ( .B(n555), .A(n556), .Z(n553) );
  AND U1667 ( .A(b[11]), .B(a[49]), .Z(n552) );
  XNOR U1668 ( .A(n557), .B(n374), .Z(n376) );
  XOR U1669 ( .A(n558), .B(n559), .Z(n374) );
  ANDN U1670 ( .B(n560), .A(n561), .Z(n558) );
  AND U1671 ( .A(a[50]), .B(b[10]), .Z(n557) );
  XNOR U1672 ( .A(n562), .B(n379), .Z(n381) );
  XOR U1673 ( .A(n563), .B(n564), .Z(n379) );
  ANDN U1674 ( .B(n565), .A(n566), .Z(n563) );
  AND U1675 ( .A(b[9]), .B(a[51]), .Z(n562) );
  XNOR U1676 ( .A(n567), .B(n384), .Z(n386) );
  XOR U1677 ( .A(n568), .B(n569), .Z(n384) );
  ANDN U1678 ( .B(n570), .A(n571), .Z(n568) );
  AND U1679 ( .A(a[52]), .B(b[8]), .Z(n567) );
  XNOR U1680 ( .A(n572), .B(n389), .Z(n391) );
  XOR U1681 ( .A(n573), .B(n574), .Z(n389) );
  ANDN U1682 ( .B(n575), .A(n576), .Z(n573) );
  AND U1683 ( .A(b[7]), .B(a[53]), .Z(n572) );
  XNOR U1684 ( .A(n577), .B(n394), .Z(n396) );
  XOR U1685 ( .A(n578), .B(n579), .Z(n394) );
  ANDN U1686 ( .B(n580), .A(n581), .Z(n578) );
  AND U1687 ( .A(b[6]), .B(a[54]), .Z(n577) );
  XNOR U1688 ( .A(n582), .B(n399), .Z(n401) );
  XOR U1689 ( .A(n583), .B(n584), .Z(n399) );
  ANDN U1690 ( .B(n585), .A(n586), .Z(n583) );
  AND U1691 ( .A(b[5]), .B(a[55]), .Z(n582) );
  XNOR U1692 ( .A(n587), .B(n404), .Z(n406) );
  XOR U1693 ( .A(n588), .B(n589), .Z(n404) );
  ANDN U1694 ( .B(n590), .A(n591), .Z(n588) );
  AND U1695 ( .A(b[4]), .B(a[56]), .Z(n587) );
  XNOR U1696 ( .A(n592), .B(n593), .Z(n418) );
  NANDN U1697 ( .A(n594), .B(n595), .Z(n593) );
  XNOR U1698 ( .A(n596), .B(n409), .Z(n411) );
  XNOR U1699 ( .A(n597), .B(n598), .Z(n409) );
  AND U1700 ( .A(n599), .B(n600), .Z(n597) );
  AND U1701 ( .A(a[57]), .B(b[3]), .Z(n596) );
  XNOR U1702 ( .A(n601), .B(n602), .Z(swire[59]) );
  XOR U1703 ( .A(n428), .B(n603), .Z(n602) );
  XOR U1704 ( .A(n427), .B(n601), .Z(n603) );
  NAND U1705 ( .A(a[59]), .B(b[0]), .Z(n427) );
  XNOR U1706 ( .A(n594), .B(n595), .Z(n428) );
  XOR U1707 ( .A(n592), .B(n604), .Z(n595) );
  NAND U1708 ( .A(a[58]), .B(b[1]), .Z(n604) );
  XOR U1709 ( .A(n600), .B(n605), .Z(n594) );
  XOR U1710 ( .A(n592), .B(n599), .Z(n605) );
  XNOR U1711 ( .A(n606), .B(n598), .Z(n599) );
  AND U1712 ( .A(a[57]), .B(b[2]), .Z(n606) );
  NANDN U1713 ( .A(n607), .B(n608), .Z(n592) );
  XOR U1714 ( .A(n598), .B(n590), .Z(n609) );
  XNOR U1715 ( .A(n589), .B(n585), .Z(n610) );
  XNOR U1716 ( .A(n584), .B(n580), .Z(n611) );
  XNOR U1717 ( .A(n579), .B(n575), .Z(n612) );
  XNOR U1718 ( .A(n574), .B(n570), .Z(n613) );
  XNOR U1719 ( .A(n569), .B(n565), .Z(n614) );
  XNOR U1720 ( .A(n564), .B(n560), .Z(n615) );
  XNOR U1721 ( .A(n616), .B(n617), .Z(n560) );
  XNOR U1722 ( .A(n559), .B(n555), .Z(n617) );
  XNOR U1723 ( .A(n554), .B(n550), .Z(n618) );
  XNOR U1724 ( .A(n549), .B(n545), .Z(n619) );
  XNOR U1725 ( .A(n544), .B(n540), .Z(n620) );
  XNOR U1726 ( .A(n539), .B(n535), .Z(n621) );
  XNOR U1727 ( .A(n534), .B(n530), .Z(n622) );
  XNOR U1728 ( .A(n529), .B(n525), .Z(n623) );
  XNOR U1729 ( .A(n524), .B(n520), .Z(n624) );
  XNOR U1730 ( .A(n519), .B(n515), .Z(n625) );
  XNOR U1731 ( .A(n514), .B(n510), .Z(n626) );
  XNOR U1732 ( .A(n509), .B(n505), .Z(n627) );
  XNOR U1733 ( .A(n504), .B(n500), .Z(n628) );
  XNOR U1734 ( .A(n499), .B(n495), .Z(n629) );
  XNOR U1735 ( .A(n494), .B(n490), .Z(n630) );
  XNOR U1736 ( .A(n489), .B(n485), .Z(n631) );
  XNOR U1737 ( .A(n484), .B(n480), .Z(n632) );
  XNOR U1738 ( .A(n479), .B(n475), .Z(n633) );
  XNOR U1739 ( .A(n474), .B(n470), .Z(n634) );
  XOR U1740 ( .A(n469), .B(n466), .Z(n635) );
  XOR U1741 ( .A(n636), .B(n637), .Z(n466) );
  XOR U1742 ( .A(n464), .B(n638), .Z(n637) );
  XOR U1743 ( .A(n639), .B(n640), .Z(n638) );
  XOR U1744 ( .A(n641), .B(n642), .Z(n640) );
  NAND U1745 ( .A(a[29]), .B(b[30]), .Z(n642) );
  AND U1746 ( .A(a[28]), .B(b[31]), .Z(n641) );
  XOR U1747 ( .A(n643), .B(n639), .Z(n636) );
  XOR U1748 ( .A(n644), .B(n645), .Z(n639) );
  NOR U1749 ( .A(n646), .B(n647), .Z(n644) );
  AND U1750 ( .A(a[30]), .B(b[29]), .Z(n643) );
  XNOR U1751 ( .A(n648), .B(n464), .Z(n465) );
  XOR U1752 ( .A(n649), .B(n650), .Z(n464) );
  ANDN U1753 ( .B(n651), .A(n652), .Z(n649) );
  AND U1754 ( .A(b[28]), .B(a[31]), .Z(n648) );
  XNOR U1755 ( .A(n653), .B(n469), .Z(n471) );
  XOR U1756 ( .A(n654), .B(n655), .Z(n469) );
  ANDN U1757 ( .B(n656), .A(n657), .Z(n654) );
  AND U1758 ( .A(a[32]), .B(b[27]), .Z(n653) );
  XNOR U1759 ( .A(n658), .B(n474), .Z(n476) );
  XOR U1760 ( .A(n659), .B(n660), .Z(n474) );
  ANDN U1761 ( .B(n661), .A(n662), .Z(n659) );
  AND U1762 ( .A(b[26]), .B(a[33]), .Z(n658) );
  XNOR U1763 ( .A(n663), .B(n479), .Z(n481) );
  XOR U1764 ( .A(n664), .B(n665), .Z(n479) );
  ANDN U1765 ( .B(n666), .A(n667), .Z(n664) );
  AND U1766 ( .A(a[34]), .B(b[25]), .Z(n663) );
  XNOR U1767 ( .A(n668), .B(n484), .Z(n486) );
  XOR U1768 ( .A(n669), .B(n670), .Z(n484) );
  ANDN U1769 ( .B(n671), .A(n672), .Z(n669) );
  AND U1770 ( .A(b[24]), .B(a[35]), .Z(n668) );
  XNOR U1771 ( .A(n673), .B(n489), .Z(n491) );
  XOR U1772 ( .A(n674), .B(n675), .Z(n489) );
  ANDN U1773 ( .B(n676), .A(n677), .Z(n674) );
  AND U1774 ( .A(a[36]), .B(b[23]), .Z(n673) );
  XNOR U1775 ( .A(n678), .B(n494), .Z(n496) );
  XOR U1776 ( .A(n679), .B(n680), .Z(n494) );
  ANDN U1777 ( .B(n681), .A(n682), .Z(n679) );
  AND U1778 ( .A(b[22]), .B(a[37]), .Z(n678) );
  XNOR U1779 ( .A(n683), .B(n499), .Z(n501) );
  XOR U1780 ( .A(n684), .B(n685), .Z(n499) );
  ANDN U1781 ( .B(n686), .A(n687), .Z(n684) );
  AND U1782 ( .A(a[38]), .B(b[21]), .Z(n683) );
  XNOR U1783 ( .A(n688), .B(n504), .Z(n506) );
  XOR U1784 ( .A(n689), .B(n690), .Z(n504) );
  ANDN U1785 ( .B(n691), .A(n692), .Z(n689) );
  AND U1786 ( .A(b[20]), .B(a[39]), .Z(n688) );
  XNOR U1787 ( .A(n693), .B(n509), .Z(n511) );
  XOR U1788 ( .A(n694), .B(n695), .Z(n509) );
  ANDN U1789 ( .B(n696), .A(n697), .Z(n694) );
  AND U1790 ( .A(a[40]), .B(b[19]), .Z(n693) );
  XNOR U1791 ( .A(n698), .B(n514), .Z(n516) );
  XOR U1792 ( .A(n699), .B(n700), .Z(n514) );
  ANDN U1793 ( .B(n701), .A(n702), .Z(n699) );
  AND U1794 ( .A(b[18]), .B(a[41]), .Z(n698) );
  XNOR U1795 ( .A(n703), .B(n519), .Z(n521) );
  XOR U1796 ( .A(n704), .B(n705), .Z(n519) );
  ANDN U1797 ( .B(n706), .A(n707), .Z(n704) );
  AND U1798 ( .A(a[42]), .B(b[17]), .Z(n703) );
  XNOR U1799 ( .A(n708), .B(n524), .Z(n526) );
  XOR U1800 ( .A(n709), .B(n710), .Z(n524) );
  ANDN U1801 ( .B(n711), .A(n712), .Z(n709) );
  AND U1802 ( .A(b[16]), .B(a[43]), .Z(n708) );
  XNOR U1803 ( .A(n713), .B(n529), .Z(n531) );
  XOR U1804 ( .A(n714), .B(n715), .Z(n529) );
  ANDN U1805 ( .B(n716), .A(n717), .Z(n714) );
  AND U1806 ( .A(a[44]), .B(b[15]), .Z(n713) );
  XNOR U1807 ( .A(n718), .B(n534), .Z(n536) );
  XOR U1808 ( .A(n719), .B(n720), .Z(n534) );
  ANDN U1809 ( .B(n721), .A(n722), .Z(n719) );
  AND U1810 ( .A(b[14]), .B(a[45]), .Z(n718) );
  XNOR U1811 ( .A(n723), .B(n539), .Z(n541) );
  XOR U1812 ( .A(n724), .B(n725), .Z(n539) );
  ANDN U1813 ( .B(n726), .A(n727), .Z(n724) );
  AND U1814 ( .A(a[46]), .B(b[13]), .Z(n723) );
  XNOR U1815 ( .A(n728), .B(n544), .Z(n546) );
  XOR U1816 ( .A(n729), .B(n730), .Z(n544) );
  ANDN U1817 ( .B(n731), .A(n732), .Z(n729) );
  AND U1818 ( .A(b[12]), .B(a[47]), .Z(n728) );
  XNOR U1819 ( .A(n733), .B(n549), .Z(n551) );
  XOR U1820 ( .A(n734), .B(n735), .Z(n549) );
  ANDN U1821 ( .B(n736), .A(n737), .Z(n734) );
  AND U1822 ( .A(a[48]), .B(b[11]), .Z(n733) );
  IV U1823 ( .A(n556), .Z(n616) );
  XNOR U1824 ( .A(n738), .B(n554), .Z(n556) );
  XOR U1825 ( .A(n739), .B(n740), .Z(n554) );
  ANDN U1826 ( .B(n741), .A(n742), .Z(n739) );
  AND U1827 ( .A(b[10]), .B(a[49]), .Z(n738) );
  XNOR U1828 ( .A(n743), .B(n559), .Z(n561) );
  XOR U1829 ( .A(n744), .B(n745), .Z(n559) );
  ANDN U1830 ( .B(n746), .A(n747), .Z(n744) );
  AND U1831 ( .A(a[50]), .B(b[9]), .Z(n743) );
  XNOR U1832 ( .A(n748), .B(n564), .Z(n566) );
  XOR U1833 ( .A(n749), .B(n750), .Z(n564) );
  ANDN U1834 ( .B(n751), .A(n752), .Z(n749) );
  AND U1835 ( .A(b[8]), .B(a[51]), .Z(n748) );
  XNOR U1836 ( .A(n753), .B(n569), .Z(n571) );
  XOR U1837 ( .A(n754), .B(n755), .Z(n569) );
  ANDN U1838 ( .B(n756), .A(n757), .Z(n754) );
  AND U1839 ( .A(a[52]), .B(b[7]), .Z(n753) );
  XNOR U1840 ( .A(n758), .B(n574), .Z(n576) );
  XOR U1841 ( .A(n759), .B(n760), .Z(n574) );
  ANDN U1842 ( .B(n761), .A(n762), .Z(n759) );
  AND U1843 ( .A(b[6]), .B(a[53]), .Z(n758) );
  XNOR U1844 ( .A(n763), .B(n579), .Z(n581) );
  XOR U1845 ( .A(n764), .B(n765), .Z(n579) );
  ANDN U1846 ( .B(n766), .A(n767), .Z(n764) );
  AND U1847 ( .A(b[5]), .B(a[54]), .Z(n763) );
  XNOR U1848 ( .A(n768), .B(n584), .Z(n586) );
  XOR U1849 ( .A(n769), .B(n770), .Z(n584) );
  ANDN U1850 ( .B(n771), .A(n772), .Z(n769) );
  AND U1851 ( .A(b[4]), .B(a[55]), .Z(n768) );
  XNOR U1852 ( .A(n773), .B(n774), .Z(n598) );
  NANDN U1853 ( .A(n775), .B(n776), .Z(n774) );
  XNOR U1854 ( .A(n777), .B(n589), .Z(n591) );
  XNOR U1855 ( .A(n778), .B(n779), .Z(n589) );
  AND U1856 ( .A(n780), .B(n781), .Z(n778) );
  AND U1857 ( .A(b[3]), .B(a[56]), .Z(n777) );
  XNOR U1858 ( .A(n782), .B(n783), .Z(swire[58]) );
  XOR U1859 ( .A(n608), .B(n785), .Z(n783) );
  XNOR U1860 ( .A(n607), .B(n784), .Z(n785) );
  IV U1861 ( .A(n782), .Z(n784) );
  NAND U1862 ( .A(a[58]), .B(b[0]), .Z(n607) );
  XNOR U1863 ( .A(n775), .B(n776), .Z(n608) );
  XOR U1864 ( .A(n773), .B(n786), .Z(n776) );
  NAND U1865 ( .A(a[57]), .B(b[1]), .Z(n786) );
  XOR U1866 ( .A(n781), .B(n787), .Z(n775) );
  XOR U1867 ( .A(n773), .B(n780), .Z(n787) );
  XNOR U1868 ( .A(n788), .B(n779), .Z(n780) );
  AND U1869 ( .A(b[2]), .B(a[56]), .Z(n788) );
  NANDN U1870 ( .A(n789), .B(n790), .Z(n773) );
  XOR U1871 ( .A(n779), .B(n771), .Z(n791) );
  XNOR U1872 ( .A(n770), .B(n766), .Z(n792) );
  XNOR U1873 ( .A(n765), .B(n761), .Z(n793) );
  XNOR U1874 ( .A(n760), .B(n756), .Z(n794) );
  XNOR U1875 ( .A(n755), .B(n751), .Z(n795) );
  XNOR U1876 ( .A(n750), .B(n746), .Z(n796) );
  XNOR U1877 ( .A(n745), .B(n741), .Z(n797) );
  XNOR U1878 ( .A(n740), .B(n736), .Z(n798) );
  XNOR U1879 ( .A(n735), .B(n731), .Z(n799) );
  XNOR U1880 ( .A(n730), .B(n726), .Z(n800) );
  XNOR U1881 ( .A(n725), .B(n721), .Z(n801) );
  XNOR U1882 ( .A(n720), .B(n716), .Z(n802) );
  XNOR U1883 ( .A(n803), .B(n804), .Z(n716) );
  XNOR U1884 ( .A(n715), .B(n711), .Z(n804) );
  XNOR U1885 ( .A(n710), .B(n706), .Z(n805) );
  XNOR U1886 ( .A(n705), .B(n701), .Z(n806) );
  XNOR U1887 ( .A(n700), .B(n696), .Z(n807) );
  XNOR U1888 ( .A(n695), .B(n691), .Z(n808) );
  XNOR U1889 ( .A(n690), .B(n686), .Z(n809) );
  XNOR U1890 ( .A(n685), .B(n681), .Z(n810) );
  XNOR U1891 ( .A(n680), .B(n676), .Z(n811) );
  XNOR U1892 ( .A(n675), .B(n671), .Z(n812) );
  XNOR U1893 ( .A(n670), .B(n666), .Z(n813) );
  XNOR U1894 ( .A(n665), .B(n661), .Z(n814) );
  XNOR U1895 ( .A(n660), .B(n656), .Z(n815) );
  XNOR U1896 ( .A(n655), .B(n651), .Z(n816) );
  XOR U1897 ( .A(n650), .B(n647), .Z(n817) );
  XOR U1898 ( .A(n818), .B(n819), .Z(n647) );
  XOR U1899 ( .A(n645), .B(n820), .Z(n819) );
  XOR U1900 ( .A(n821), .B(n822), .Z(n820) );
  XOR U1901 ( .A(n823), .B(n824), .Z(n822) );
  NAND U1902 ( .A(a[28]), .B(b[30]), .Z(n824) );
  AND U1903 ( .A(a[27]), .B(b[31]), .Z(n823) );
  XOR U1904 ( .A(n825), .B(n821), .Z(n818) );
  XOR U1905 ( .A(n826), .B(n827), .Z(n821) );
  NOR U1906 ( .A(n828), .B(n829), .Z(n826) );
  AND U1907 ( .A(b[29]), .B(a[29]), .Z(n825) );
  XNOR U1908 ( .A(n830), .B(n645), .Z(n646) );
  XOR U1909 ( .A(n831), .B(n832), .Z(n645) );
  ANDN U1910 ( .B(n833), .A(n834), .Z(n831) );
  AND U1911 ( .A(a[30]), .B(b[28]), .Z(n830) );
  XNOR U1912 ( .A(n835), .B(n650), .Z(n652) );
  XOR U1913 ( .A(n836), .B(n837), .Z(n650) );
  ANDN U1914 ( .B(n838), .A(n839), .Z(n836) );
  AND U1915 ( .A(b[27]), .B(a[31]), .Z(n835) );
  XNOR U1916 ( .A(n840), .B(n655), .Z(n657) );
  XOR U1917 ( .A(n841), .B(n842), .Z(n655) );
  ANDN U1918 ( .B(n843), .A(n844), .Z(n841) );
  AND U1919 ( .A(a[32]), .B(b[26]), .Z(n840) );
  XNOR U1920 ( .A(n845), .B(n660), .Z(n662) );
  XOR U1921 ( .A(n846), .B(n847), .Z(n660) );
  ANDN U1922 ( .B(n848), .A(n849), .Z(n846) );
  AND U1923 ( .A(b[25]), .B(a[33]), .Z(n845) );
  XNOR U1924 ( .A(n850), .B(n665), .Z(n667) );
  XOR U1925 ( .A(n851), .B(n852), .Z(n665) );
  ANDN U1926 ( .B(n853), .A(n854), .Z(n851) );
  AND U1927 ( .A(a[34]), .B(b[24]), .Z(n850) );
  XNOR U1928 ( .A(n855), .B(n670), .Z(n672) );
  XOR U1929 ( .A(n856), .B(n857), .Z(n670) );
  ANDN U1930 ( .B(n858), .A(n859), .Z(n856) );
  AND U1931 ( .A(b[23]), .B(a[35]), .Z(n855) );
  XNOR U1932 ( .A(n860), .B(n675), .Z(n677) );
  XOR U1933 ( .A(n861), .B(n862), .Z(n675) );
  ANDN U1934 ( .B(n863), .A(n864), .Z(n861) );
  AND U1935 ( .A(a[36]), .B(b[22]), .Z(n860) );
  XNOR U1936 ( .A(n865), .B(n680), .Z(n682) );
  XOR U1937 ( .A(n866), .B(n867), .Z(n680) );
  ANDN U1938 ( .B(n868), .A(n869), .Z(n866) );
  AND U1939 ( .A(b[21]), .B(a[37]), .Z(n865) );
  XNOR U1940 ( .A(n870), .B(n685), .Z(n687) );
  XOR U1941 ( .A(n871), .B(n872), .Z(n685) );
  ANDN U1942 ( .B(n873), .A(n874), .Z(n871) );
  AND U1943 ( .A(a[38]), .B(b[20]), .Z(n870) );
  XNOR U1944 ( .A(n875), .B(n690), .Z(n692) );
  XOR U1945 ( .A(n876), .B(n877), .Z(n690) );
  ANDN U1946 ( .B(n878), .A(n879), .Z(n876) );
  AND U1947 ( .A(b[19]), .B(a[39]), .Z(n875) );
  XNOR U1948 ( .A(n880), .B(n695), .Z(n697) );
  XOR U1949 ( .A(n881), .B(n882), .Z(n695) );
  ANDN U1950 ( .B(n883), .A(n884), .Z(n881) );
  AND U1951 ( .A(a[40]), .B(b[18]), .Z(n880) );
  XNOR U1952 ( .A(n885), .B(n700), .Z(n702) );
  XOR U1953 ( .A(n886), .B(n887), .Z(n700) );
  ANDN U1954 ( .B(n888), .A(n889), .Z(n886) );
  AND U1955 ( .A(b[17]), .B(a[41]), .Z(n885) );
  XNOR U1956 ( .A(n890), .B(n705), .Z(n707) );
  XOR U1957 ( .A(n891), .B(n892), .Z(n705) );
  ANDN U1958 ( .B(n893), .A(n894), .Z(n891) );
  AND U1959 ( .A(a[42]), .B(b[16]), .Z(n890) );
  IV U1960 ( .A(n712), .Z(n803) );
  XNOR U1961 ( .A(n895), .B(n710), .Z(n712) );
  XOR U1962 ( .A(n896), .B(n897), .Z(n710) );
  ANDN U1963 ( .B(n898), .A(n899), .Z(n896) );
  AND U1964 ( .A(b[15]), .B(a[43]), .Z(n895) );
  XNOR U1965 ( .A(n900), .B(n715), .Z(n717) );
  XOR U1966 ( .A(n901), .B(n902), .Z(n715) );
  ANDN U1967 ( .B(n903), .A(n904), .Z(n901) );
  AND U1968 ( .A(a[44]), .B(b[14]), .Z(n900) );
  XNOR U1969 ( .A(n905), .B(n720), .Z(n722) );
  XOR U1970 ( .A(n906), .B(n907), .Z(n720) );
  ANDN U1971 ( .B(n908), .A(n909), .Z(n906) );
  AND U1972 ( .A(b[13]), .B(a[45]), .Z(n905) );
  XNOR U1973 ( .A(n910), .B(n725), .Z(n727) );
  XOR U1974 ( .A(n911), .B(n912), .Z(n725) );
  ANDN U1975 ( .B(n913), .A(n914), .Z(n911) );
  AND U1976 ( .A(a[46]), .B(b[12]), .Z(n910) );
  XNOR U1977 ( .A(n915), .B(n730), .Z(n732) );
  XOR U1978 ( .A(n916), .B(n917), .Z(n730) );
  ANDN U1979 ( .B(n918), .A(n919), .Z(n916) );
  AND U1980 ( .A(b[11]), .B(a[47]), .Z(n915) );
  XNOR U1981 ( .A(n920), .B(n735), .Z(n737) );
  XOR U1982 ( .A(n921), .B(n922), .Z(n735) );
  ANDN U1983 ( .B(n923), .A(n924), .Z(n921) );
  AND U1984 ( .A(a[48]), .B(b[10]), .Z(n920) );
  XNOR U1985 ( .A(n925), .B(n740), .Z(n742) );
  XOR U1986 ( .A(n926), .B(n927), .Z(n740) );
  ANDN U1987 ( .B(n928), .A(n929), .Z(n926) );
  AND U1988 ( .A(b[9]), .B(a[49]), .Z(n925) );
  XNOR U1989 ( .A(n930), .B(n745), .Z(n747) );
  XOR U1990 ( .A(n931), .B(n932), .Z(n745) );
  ANDN U1991 ( .B(n933), .A(n934), .Z(n931) );
  AND U1992 ( .A(a[50]), .B(b[8]), .Z(n930) );
  XNOR U1993 ( .A(n935), .B(n750), .Z(n752) );
  XOR U1994 ( .A(n936), .B(n937), .Z(n750) );
  ANDN U1995 ( .B(n938), .A(n939), .Z(n936) );
  AND U1996 ( .A(b[7]), .B(a[51]), .Z(n935) );
  XNOR U1997 ( .A(n940), .B(n755), .Z(n757) );
  XOR U1998 ( .A(n941), .B(n942), .Z(n755) );
  ANDN U1999 ( .B(n943), .A(n944), .Z(n941) );
  AND U2000 ( .A(b[6]), .B(a[52]), .Z(n940) );
  XNOR U2001 ( .A(n945), .B(n760), .Z(n762) );
  XOR U2002 ( .A(n946), .B(n947), .Z(n760) );
  ANDN U2003 ( .B(n948), .A(n949), .Z(n946) );
  AND U2004 ( .A(b[5]), .B(a[53]), .Z(n945) );
  XNOR U2005 ( .A(n950), .B(n765), .Z(n767) );
  XOR U2006 ( .A(n951), .B(n952), .Z(n765) );
  ANDN U2007 ( .B(n953), .A(n954), .Z(n951) );
  AND U2008 ( .A(b[4]), .B(a[54]), .Z(n950) );
  XNOR U2009 ( .A(n955), .B(n956), .Z(n779) );
  NANDN U2010 ( .A(n957), .B(n958), .Z(n956) );
  XNOR U2011 ( .A(n959), .B(n770), .Z(n772) );
  XNOR U2012 ( .A(n960), .B(n961), .Z(n770) );
  AND U2013 ( .A(n962), .B(n963), .Z(n960) );
  AND U2014 ( .A(b[3]), .B(a[55]), .Z(n959) );
  XNOR U2015 ( .A(n964), .B(n965), .Z(swire[57]) );
  XOR U2016 ( .A(n790), .B(n966), .Z(n965) );
  XOR U2017 ( .A(n789), .B(n964), .Z(n966) );
  NAND U2018 ( .A(a[57]), .B(b[0]), .Z(n789) );
  XNOR U2019 ( .A(n957), .B(n958), .Z(n790) );
  XOR U2020 ( .A(n955), .B(n967), .Z(n958) );
  NAND U2021 ( .A(a[56]), .B(b[1]), .Z(n967) );
  XOR U2022 ( .A(n963), .B(n968), .Z(n957) );
  XOR U2023 ( .A(n955), .B(n962), .Z(n968) );
  XNOR U2024 ( .A(n969), .B(n961), .Z(n962) );
  AND U2025 ( .A(b[2]), .B(a[55]), .Z(n969) );
  NANDN U2026 ( .A(n970), .B(n971), .Z(n955) );
  XOR U2027 ( .A(n961), .B(n953), .Z(n972) );
  XNOR U2028 ( .A(n952), .B(n948), .Z(n973) );
  XNOR U2029 ( .A(n947), .B(n943), .Z(n974) );
  XNOR U2030 ( .A(n942), .B(n938), .Z(n975) );
  XNOR U2031 ( .A(n937), .B(n933), .Z(n976) );
  XNOR U2032 ( .A(n932), .B(n928), .Z(n977) );
  XNOR U2033 ( .A(n927), .B(n923), .Z(n978) );
  XNOR U2034 ( .A(n979), .B(n980), .Z(n923) );
  XNOR U2035 ( .A(n922), .B(n918), .Z(n980) );
  XNOR U2036 ( .A(n917), .B(n913), .Z(n981) );
  XNOR U2037 ( .A(n912), .B(n908), .Z(n982) );
  XNOR U2038 ( .A(n983), .B(n984), .Z(n908) );
  XNOR U2039 ( .A(n907), .B(n903), .Z(n984) );
  XNOR U2040 ( .A(n902), .B(n898), .Z(n985) );
  XNOR U2041 ( .A(n897), .B(n893), .Z(n986) );
  XNOR U2042 ( .A(n892), .B(n888), .Z(n987) );
  XNOR U2043 ( .A(n887), .B(n883), .Z(n988) );
  XNOR U2044 ( .A(n882), .B(n878), .Z(n989) );
  XNOR U2045 ( .A(n877), .B(n873), .Z(n990) );
  XNOR U2046 ( .A(n872), .B(n868), .Z(n991) );
  XNOR U2047 ( .A(n867), .B(n863), .Z(n992) );
  XNOR U2048 ( .A(n862), .B(n858), .Z(n993) );
  XNOR U2049 ( .A(n857), .B(n853), .Z(n994) );
  XNOR U2050 ( .A(n852), .B(n848), .Z(n995) );
  XNOR U2051 ( .A(n847), .B(n843), .Z(n996) );
  XNOR U2052 ( .A(n842), .B(n838), .Z(n997) );
  XNOR U2053 ( .A(n837), .B(n833), .Z(n998) );
  XOR U2054 ( .A(n832), .B(n829), .Z(n999) );
  XOR U2055 ( .A(n1000), .B(n1001), .Z(n829) );
  XOR U2056 ( .A(n827), .B(n1002), .Z(n1001) );
  XOR U2057 ( .A(n1003), .B(n1004), .Z(n1002) );
  XOR U2058 ( .A(n1005), .B(n1006), .Z(n1004) );
  NAND U2059 ( .A(a[27]), .B(b[30]), .Z(n1006) );
  AND U2060 ( .A(a[26]), .B(b[31]), .Z(n1005) );
  XOR U2061 ( .A(n1007), .B(n1003), .Z(n1000) );
  XOR U2062 ( .A(n1008), .B(n1009), .Z(n1003) );
  NOR U2063 ( .A(n1010), .B(n1011), .Z(n1008) );
  AND U2064 ( .A(a[28]), .B(b[29]), .Z(n1007) );
  XNOR U2065 ( .A(n1012), .B(n827), .Z(n828) );
  XOR U2066 ( .A(n1013), .B(n1014), .Z(n827) );
  ANDN U2067 ( .B(n1015), .A(n1016), .Z(n1013) );
  AND U2068 ( .A(b[28]), .B(a[29]), .Z(n1012) );
  XNOR U2069 ( .A(n1017), .B(n832), .Z(n834) );
  XOR U2070 ( .A(n1018), .B(n1019), .Z(n832) );
  ANDN U2071 ( .B(n1020), .A(n1021), .Z(n1018) );
  AND U2072 ( .A(a[30]), .B(b[27]), .Z(n1017) );
  XNOR U2073 ( .A(n1022), .B(n837), .Z(n839) );
  XOR U2074 ( .A(n1023), .B(n1024), .Z(n837) );
  ANDN U2075 ( .B(n1025), .A(n1026), .Z(n1023) );
  AND U2076 ( .A(b[26]), .B(a[31]), .Z(n1022) );
  XNOR U2077 ( .A(n1027), .B(n842), .Z(n844) );
  XOR U2078 ( .A(n1028), .B(n1029), .Z(n842) );
  ANDN U2079 ( .B(n1030), .A(n1031), .Z(n1028) );
  AND U2080 ( .A(a[32]), .B(b[25]), .Z(n1027) );
  XNOR U2081 ( .A(n1032), .B(n847), .Z(n849) );
  XOR U2082 ( .A(n1033), .B(n1034), .Z(n847) );
  ANDN U2083 ( .B(n1035), .A(n1036), .Z(n1033) );
  AND U2084 ( .A(b[24]), .B(a[33]), .Z(n1032) );
  XNOR U2085 ( .A(n1037), .B(n852), .Z(n854) );
  XOR U2086 ( .A(n1038), .B(n1039), .Z(n852) );
  ANDN U2087 ( .B(n1040), .A(n1041), .Z(n1038) );
  AND U2088 ( .A(a[34]), .B(b[23]), .Z(n1037) );
  XNOR U2089 ( .A(n1042), .B(n857), .Z(n859) );
  XOR U2090 ( .A(n1043), .B(n1044), .Z(n857) );
  ANDN U2091 ( .B(n1045), .A(n1046), .Z(n1043) );
  AND U2092 ( .A(b[22]), .B(a[35]), .Z(n1042) );
  XNOR U2093 ( .A(n1047), .B(n862), .Z(n864) );
  XOR U2094 ( .A(n1048), .B(n1049), .Z(n862) );
  ANDN U2095 ( .B(n1050), .A(n1051), .Z(n1048) );
  AND U2096 ( .A(a[36]), .B(b[21]), .Z(n1047) );
  XNOR U2097 ( .A(n1052), .B(n867), .Z(n869) );
  XOR U2098 ( .A(n1053), .B(n1054), .Z(n867) );
  ANDN U2099 ( .B(n1055), .A(n1056), .Z(n1053) );
  AND U2100 ( .A(b[20]), .B(a[37]), .Z(n1052) );
  XNOR U2101 ( .A(n1057), .B(n872), .Z(n874) );
  XOR U2102 ( .A(n1058), .B(n1059), .Z(n872) );
  ANDN U2103 ( .B(n1060), .A(n1061), .Z(n1058) );
  AND U2104 ( .A(a[38]), .B(b[19]), .Z(n1057) );
  XNOR U2105 ( .A(n1062), .B(n877), .Z(n879) );
  XOR U2106 ( .A(n1063), .B(n1064), .Z(n877) );
  ANDN U2107 ( .B(n1065), .A(n1066), .Z(n1063) );
  AND U2108 ( .A(b[18]), .B(a[39]), .Z(n1062) );
  XNOR U2109 ( .A(n1067), .B(n882), .Z(n884) );
  XOR U2110 ( .A(n1068), .B(n1069), .Z(n882) );
  ANDN U2111 ( .B(n1070), .A(n1071), .Z(n1068) );
  AND U2112 ( .A(a[40]), .B(b[17]), .Z(n1067) );
  XNOR U2113 ( .A(n1072), .B(n887), .Z(n889) );
  XOR U2114 ( .A(n1073), .B(n1074), .Z(n887) );
  ANDN U2115 ( .B(n1075), .A(n1076), .Z(n1073) );
  AND U2116 ( .A(b[16]), .B(a[41]), .Z(n1072) );
  XNOR U2117 ( .A(n1077), .B(n892), .Z(n894) );
  XOR U2118 ( .A(n1078), .B(n1079), .Z(n892) );
  ANDN U2119 ( .B(n1080), .A(n1081), .Z(n1078) );
  AND U2120 ( .A(a[42]), .B(b[15]), .Z(n1077) );
  XNOR U2121 ( .A(n1082), .B(n897), .Z(n899) );
  XOR U2122 ( .A(n1083), .B(n1084), .Z(n897) );
  ANDN U2123 ( .B(n1085), .A(n1086), .Z(n1083) );
  AND U2124 ( .A(b[14]), .B(a[43]), .Z(n1082) );
  IV U2125 ( .A(n904), .Z(n983) );
  XNOR U2126 ( .A(n1087), .B(n902), .Z(n904) );
  XOR U2127 ( .A(n1088), .B(n1089), .Z(n902) );
  ANDN U2128 ( .B(n1090), .A(n1091), .Z(n1088) );
  AND U2129 ( .A(a[44]), .B(b[13]), .Z(n1087) );
  XNOR U2130 ( .A(n1092), .B(n907), .Z(n909) );
  XOR U2131 ( .A(n1093), .B(n1094), .Z(n907) );
  ANDN U2132 ( .B(n1095), .A(n1096), .Z(n1093) );
  AND U2133 ( .A(b[12]), .B(a[45]), .Z(n1092) );
  XNOR U2134 ( .A(n1097), .B(n912), .Z(n914) );
  XOR U2135 ( .A(n1098), .B(n1099), .Z(n912) );
  ANDN U2136 ( .B(n1100), .A(n1101), .Z(n1098) );
  AND U2137 ( .A(a[46]), .B(b[11]), .Z(n1097) );
  IV U2138 ( .A(n919), .Z(n979) );
  XNOR U2139 ( .A(n1102), .B(n917), .Z(n919) );
  XOR U2140 ( .A(n1103), .B(n1104), .Z(n917) );
  ANDN U2141 ( .B(n1105), .A(n1106), .Z(n1103) );
  AND U2142 ( .A(b[10]), .B(a[47]), .Z(n1102) );
  XNOR U2143 ( .A(n1107), .B(n922), .Z(n924) );
  XOR U2144 ( .A(n1108), .B(n1109), .Z(n922) );
  ANDN U2145 ( .B(n1110), .A(n1111), .Z(n1108) );
  AND U2146 ( .A(a[48]), .B(b[9]), .Z(n1107) );
  XNOR U2147 ( .A(n1112), .B(n927), .Z(n929) );
  XOR U2148 ( .A(n1113), .B(n1114), .Z(n927) );
  ANDN U2149 ( .B(n1115), .A(n1116), .Z(n1113) );
  AND U2150 ( .A(b[8]), .B(a[49]), .Z(n1112) );
  XNOR U2151 ( .A(n1117), .B(n932), .Z(n934) );
  XOR U2152 ( .A(n1118), .B(n1119), .Z(n932) );
  ANDN U2153 ( .B(n1120), .A(n1121), .Z(n1118) );
  AND U2154 ( .A(a[50]), .B(b[7]), .Z(n1117) );
  XNOR U2155 ( .A(n1122), .B(n937), .Z(n939) );
  XOR U2156 ( .A(n1123), .B(n1124), .Z(n937) );
  ANDN U2157 ( .B(n1125), .A(n1126), .Z(n1123) );
  AND U2158 ( .A(b[6]), .B(a[51]), .Z(n1122) );
  XNOR U2159 ( .A(n1127), .B(n942), .Z(n944) );
  XOR U2160 ( .A(n1128), .B(n1129), .Z(n942) );
  ANDN U2161 ( .B(n1130), .A(n1131), .Z(n1128) );
  AND U2162 ( .A(b[5]), .B(a[52]), .Z(n1127) );
  XNOR U2163 ( .A(n1132), .B(n947), .Z(n949) );
  XOR U2164 ( .A(n1133), .B(n1134), .Z(n947) );
  ANDN U2165 ( .B(n1135), .A(n1136), .Z(n1133) );
  AND U2166 ( .A(b[4]), .B(a[53]), .Z(n1132) );
  XNOR U2167 ( .A(n1137), .B(n1138), .Z(n961) );
  NANDN U2168 ( .A(n1139), .B(n1140), .Z(n1138) );
  XNOR U2169 ( .A(n1141), .B(n952), .Z(n954) );
  XNOR U2170 ( .A(n1142), .B(n1143), .Z(n952) );
  AND U2171 ( .A(n1144), .B(n1145), .Z(n1142) );
  AND U2172 ( .A(b[3]), .B(a[54]), .Z(n1141) );
  XNOR U2173 ( .A(n1146), .B(n1147), .Z(swire[56]) );
  XOR U2174 ( .A(n971), .B(n1149), .Z(n1147) );
  XNOR U2175 ( .A(n970), .B(n1148), .Z(n1149) );
  IV U2176 ( .A(n1146), .Z(n1148) );
  NAND U2177 ( .A(a[56]), .B(b[0]), .Z(n970) );
  XNOR U2178 ( .A(n1139), .B(n1140), .Z(n971) );
  XOR U2179 ( .A(n1137), .B(n1150), .Z(n1140) );
  NAND U2180 ( .A(b[1]), .B(a[55]), .Z(n1150) );
  XOR U2181 ( .A(n1145), .B(n1151), .Z(n1139) );
  XOR U2182 ( .A(n1137), .B(n1144), .Z(n1151) );
  XNOR U2183 ( .A(n1152), .B(n1143), .Z(n1144) );
  AND U2184 ( .A(b[2]), .B(a[54]), .Z(n1152) );
  NANDN U2185 ( .A(n1153), .B(n1154), .Z(n1137) );
  XOR U2186 ( .A(n1143), .B(n1135), .Z(n1155) );
  XNOR U2187 ( .A(n1134), .B(n1130), .Z(n1156) );
  XNOR U2188 ( .A(n1129), .B(n1125), .Z(n1157) );
  XNOR U2189 ( .A(n1124), .B(n1120), .Z(n1158) );
  XNOR U2190 ( .A(n1119), .B(n1115), .Z(n1159) );
  XNOR U2191 ( .A(n1114), .B(n1110), .Z(n1160) );
  XNOR U2192 ( .A(n1109), .B(n1105), .Z(n1161) );
  XNOR U2193 ( .A(n1104), .B(n1100), .Z(n1162) );
  XNOR U2194 ( .A(n1099), .B(n1095), .Z(n1163) );
  XNOR U2195 ( .A(n1094), .B(n1090), .Z(n1164) );
  XNOR U2196 ( .A(n1089), .B(n1085), .Z(n1165) );
  XNOR U2197 ( .A(n1084), .B(n1080), .Z(n1166) );
  XNOR U2198 ( .A(n1079), .B(n1075), .Z(n1167) );
  XNOR U2199 ( .A(n1074), .B(n1070), .Z(n1168) );
  XNOR U2200 ( .A(n1069), .B(n1065), .Z(n1169) );
  XNOR U2201 ( .A(n1170), .B(n1171), .Z(n1065) );
  XNOR U2202 ( .A(n1064), .B(n1060), .Z(n1171) );
  XNOR U2203 ( .A(n1059), .B(n1055), .Z(n1172) );
  XNOR U2204 ( .A(n1054), .B(n1050), .Z(n1173) );
  XNOR U2205 ( .A(n1049), .B(n1045), .Z(n1174) );
  XNOR U2206 ( .A(n1044), .B(n1040), .Z(n1175) );
  XNOR U2207 ( .A(n1039), .B(n1035), .Z(n1176) );
  XNOR U2208 ( .A(n1034), .B(n1030), .Z(n1177) );
  XNOR U2209 ( .A(n1029), .B(n1025), .Z(n1178) );
  XNOR U2210 ( .A(n1024), .B(n1020), .Z(n1179) );
  XNOR U2211 ( .A(n1019), .B(n1015), .Z(n1180) );
  XOR U2212 ( .A(n1014), .B(n1011), .Z(n1181) );
  XOR U2213 ( .A(n1182), .B(n1183), .Z(n1011) );
  XOR U2214 ( .A(n1009), .B(n1184), .Z(n1183) );
  XOR U2215 ( .A(n1185), .B(n1186), .Z(n1184) );
  XOR U2216 ( .A(n1187), .B(n1188), .Z(n1186) );
  NAND U2217 ( .A(a[26]), .B(b[30]), .Z(n1188) );
  AND U2218 ( .A(a[25]), .B(b[31]), .Z(n1187) );
  XOR U2219 ( .A(n1189), .B(n1185), .Z(n1182) );
  XOR U2220 ( .A(n1190), .B(n1191), .Z(n1185) );
  NOR U2221 ( .A(n1192), .B(n1193), .Z(n1190) );
  AND U2222 ( .A(a[27]), .B(b[29]), .Z(n1189) );
  XNOR U2223 ( .A(n1194), .B(n1009), .Z(n1010) );
  XOR U2224 ( .A(n1195), .B(n1196), .Z(n1009) );
  ANDN U2225 ( .B(n1197), .A(n1198), .Z(n1195) );
  AND U2226 ( .A(a[28]), .B(b[28]), .Z(n1194) );
  XNOR U2227 ( .A(n1199), .B(n1014), .Z(n1016) );
  XOR U2228 ( .A(n1200), .B(n1201), .Z(n1014) );
  ANDN U2229 ( .B(n1202), .A(n1203), .Z(n1200) );
  AND U2230 ( .A(b[27]), .B(a[29]), .Z(n1199) );
  XNOR U2231 ( .A(n1204), .B(n1019), .Z(n1021) );
  XOR U2232 ( .A(n1205), .B(n1206), .Z(n1019) );
  ANDN U2233 ( .B(n1207), .A(n1208), .Z(n1205) );
  AND U2234 ( .A(a[30]), .B(b[26]), .Z(n1204) );
  XNOR U2235 ( .A(n1209), .B(n1024), .Z(n1026) );
  XOR U2236 ( .A(n1210), .B(n1211), .Z(n1024) );
  ANDN U2237 ( .B(n1212), .A(n1213), .Z(n1210) );
  AND U2238 ( .A(b[25]), .B(a[31]), .Z(n1209) );
  XNOR U2239 ( .A(n1214), .B(n1029), .Z(n1031) );
  XOR U2240 ( .A(n1215), .B(n1216), .Z(n1029) );
  ANDN U2241 ( .B(n1217), .A(n1218), .Z(n1215) );
  AND U2242 ( .A(a[32]), .B(b[24]), .Z(n1214) );
  XNOR U2243 ( .A(n1219), .B(n1034), .Z(n1036) );
  XOR U2244 ( .A(n1220), .B(n1221), .Z(n1034) );
  ANDN U2245 ( .B(n1222), .A(n1223), .Z(n1220) );
  AND U2246 ( .A(b[23]), .B(a[33]), .Z(n1219) );
  XNOR U2247 ( .A(n1224), .B(n1039), .Z(n1041) );
  XOR U2248 ( .A(n1225), .B(n1226), .Z(n1039) );
  ANDN U2249 ( .B(n1227), .A(n1228), .Z(n1225) );
  AND U2250 ( .A(a[34]), .B(b[22]), .Z(n1224) );
  XNOR U2251 ( .A(n1229), .B(n1044), .Z(n1046) );
  XOR U2252 ( .A(n1230), .B(n1231), .Z(n1044) );
  ANDN U2253 ( .B(n1232), .A(n1233), .Z(n1230) );
  AND U2254 ( .A(b[21]), .B(a[35]), .Z(n1229) );
  XNOR U2255 ( .A(n1234), .B(n1049), .Z(n1051) );
  XOR U2256 ( .A(n1235), .B(n1236), .Z(n1049) );
  ANDN U2257 ( .B(n1237), .A(n1238), .Z(n1235) );
  AND U2258 ( .A(a[36]), .B(b[20]), .Z(n1234) );
  XNOR U2259 ( .A(n1239), .B(n1054), .Z(n1056) );
  XOR U2260 ( .A(n1240), .B(n1241), .Z(n1054) );
  ANDN U2261 ( .B(n1242), .A(n1243), .Z(n1240) );
  AND U2262 ( .A(b[19]), .B(a[37]), .Z(n1239) );
  IV U2263 ( .A(n1061), .Z(n1170) );
  XNOR U2264 ( .A(n1244), .B(n1059), .Z(n1061) );
  XOR U2265 ( .A(n1245), .B(n1246), .Z(n1059) );
  ANDN U2266 ( .B(n1247), .A(n1248), .Z(n1245) );
  AND U2267 ( .A(a[38]), .B(b[18]), .Z(n1244) );
  XNOR U2268 ( .A(n1249), .B(n1064), .Z(n1066) );
  XOR U2269 ( .A(n1250), .B(n1251), .Z(n1064) );
  ANDN U2270 ( .B(n1252), .A(n1253), .Z(n1250) );
  AND U2271 ( .A(b[17]), .B(a[39]), .Z(n1249) );
  XNOR U2272 ( .A(n1254), .B(n1069), .Z(n1071) );
  XOR U2273 ( .A(n1255), .B(n1256), .Z(n1069) );
  ANDN U2274 ( .B(n1257), .A(n1258), .Z(n1255) );
  AND U2275 ( .A(a[40]), .B(b[16]), .Z(n1254) );
  XNOR U2276 ( .A(n1259), .B(n1074), .Z(n1076) );
  XOR U2277 ( .A(n1260), .B(n1261), .Z(n1074) );
  ANDN U2278 ( .B(n1262), .A(n1263), .Z(n1260) );
  AND U2279 ( .A(b[15]), .B(a[41]), .Z(n1259) );
  XNOR U2280 ( .A(n1264), .B(n1079), .Z(n1081) );
  XOR U2281 ( .A(n1265), .B(n1266), .Z(n1079) );
  ANDN U2282 ( .B(n1267), .A(n1268), .Z(n1265) );
  AND U2283 ( .A(a[42]), .B(b[14]), .Z(n1264) );
  XNOR U2284 ( .A(n1269), .B(n1084), .Z(n1086) );
  XOR U2285 ( .A(n1270), .B(n1271), .Z(n1084) );
  ANDN U2286 ( .B(n1272), .A(n1273), .Z(n1270) );
  AND U2287 ( .A(b[13]), .B(a[43]), .Z(n1269) );
  XNOR U2288 ( .A(n1274), .B(n1089), .Z(n1091) );
  XOR U2289 ( .A(n1275), .B(n1276), .Z(n1089) );
  ANDN U2290 ( .B(n1277), .A(n1278), .Z(n1275) );
  AND U2291 ( .A(a[44]), .B(b[12]), .Z(n1274) );
  XNOR U2292 ( .A(n1279), .B(n1094), .Z(n1096) );
  XOR U2293 ( .A(n1280), .B(n1281), .Z(n1094) );
  ANDN U2294 ( .B(n1282), .A(n1283), .Z(n1280) );
  AND U2295 ( .A(b[11]), .B(a[45]), .Z(n1279) );
  XNOR U2296 ( .A(n1284), .B(n1099), .Z(n1101) );
  XOR U2297 ( .A(n1285), .B(n1286), .Z(n1099) );
  ANDN U2298 ( .B(n1287), .A(n1288), .Z(n1285) );
  AND U2299 ( .A(a[46]), .B(b[10]), .Z(n1284) );
  XNOR U2300 ( .A(n1289), .B(n1104), .Z(n1106) );
  XOR U2301 ( .A(n1290), .B(n1291), .Z(n1104) );
  ANDN U2302 ( .B(n1292), .A(n1293), .Z(n1290) );
  AND U2303 ( .A(b[9]), .B(a[47]), .Z(n1289) );
  XNOR U2304 ( .A(n1294), .B(n1109), .Z(n1111) );
  XOR U2305 ( .A(n1295), .B(n1296), .Z(n1109) );
  ANDN U2306 ( .B(n1297), .A(n1298), .Z(n1295) );
  AND U2307 ( .A(a[48]), .B(b[8]), .Z(n1294) );
  XNOR U2308 ( .A(n1299), .B(n1114), .Z(n1116) );
  XOR U2309 ( .A(n1300), .B(n1301), .Z(n1114) );
  ANDN U2310 ( .B(n1302), .A(n1303), .Z(n1300) );
  AND U2311 ( .A(b[7]), .B(a[49]), .Z(n1299) );
  XNOR U2312 ( .A(n1304), .B(n1119), .Z(n1121) );
  XOR U2313 ( .A(n1305), .B(n1306), .Z(n1119) );
  ANDN U2314 ( .B(n1307), .A(n1308), .Z(n1305) );
  AND U2315 ( .A(b[6]), .B(a[50]), .Z(n1304) );
  XNOR U2316 ( .A(n1309), .B(n1124), .Z(n1126) );
  XOR U2317 ( .A(n1310), .B(n1311), .Z(n1124) );
  ANDN U2318 ( .B(n1312), .A(n1313), .Z(n1310) );
  AND U2319 ( .A(b[5]), .B(a[51]), .Z(n1309) );
  XNOR U2320 ( .A(n1314), .B(n1129), .Z(n1131) );
  XOR U2321 ( .A(n1315), .B(n1316), .Z(n1129) );
  ANDN U2322 ( .B(n1317), .A(n1318), .Z(n1315) );
  AND U2323 ( .A(b[4]), .B(a[52]), .Z(n1314) );
  XNOR U2324 ( .A(n1319), .B(n1320), .Z(n1143) );
  NANDN U2325 ( .A(n1321), .B(n1322), .Z(n1320) );
  XNOR U2326 ( .A(n1323), .B(n1134), .Z(n1136) );
  XNOR U2327 ( .A(n1324), .B(n1325), .Z(n1134) );
  AND U2328 ( .A(n1326), .B(n1327), .Z(n1324) );
  AND U2329 ( .A(b[3]), .B(a[53]), .Z(n1323) );
  XNOR U2330 ( .A(n1328), .B(n1329), .Z(swire[55]) );
  XOR U2331 ( .A(n1154), .B(n1330), .Z(n1329) );
  XOR U2332 ( .A(n1153), .B(n1328), .Z(n1330) );
  NAND U2333 ( .A(a[55]), .B(b[0]), .Z(n1153) );
  XNOR U2334 ( .A(n1321), .B(n1322), .Z(n1154) );
  XOR U2335 ( .A(n1319), .B(n1331), .Z(n1322) );
  NAND U2336 ( .A(a[54]), .B(b[1]), .Z(n1331) );
  XOR U2337 ( .A(n1327), .B(n1332), .Z(n1321) );
  XOR U2338 ( .A(n1319), .B(n1326), .Z(n1332) );
  XNOR U2339 ( .A(n1333), .B(n1325), .Z(n1326) );
  AND U2340 ( .A(b[2]), .B(a[53]), .Z(n1333) );
  NANDN U2341 ( .A(n1334), .B(n1335), .Z(n1319) );
  XOR U2342 ( .A(n1325), .B(n1317), .Z(n1336) );
  XNOR U2343 ( .A(n1316), .B(n1312), .Z(n1337) );
  XNOR U2344 ( .A(n1311), .B(n1307), .Z(n1338) );
  XNOR U2345 ( .A(n1306), .B(n1302), .Z(n1339) );
  XNOR U2346 ( .A(n1301), .B(n1297), .Z(n1340) );
  XNOR U2347 ( .A(n1296), .B(n1292), .Z(n1341) );
  XNOR U2348 ( .A(n1291), .B(n1287), .Z(n1342) );
  XNOR U2349 ( .A(n1286), .B(n1282), .Z(n1343) );
  XNOR U2350 ( .A(n1281), .B(n1277), .Z(n1344) );
  XNOR U2351 ( .A(n1276), .B(n1272), .Z(n1345) );
  XNOR U2352 ( .A(n1271), .B(n1267), .Z(n1346) );
  XNOR U2353 ( .A(n1266), .B(n1262), .Z(n1347) );
  XNOR U2354 ( .A(n1348), .B(n1349), .Z(n1262) );
  XNOR U2355 ( .A(n1261), .B(n1257), .Z(n1349) );
  XNOR U2356 ( .A(n1256), .B(n1252), .Z(n1350) );
  XNOR U2357 ( .A(n1251), .B(n1247), .Z(n1351) );
  XNOR U2358 ( .A(n1246), .B(n1242), .Z(n1352) );
  XNOR U2359 ( .A(n1241), .B(n1237), .Z(n1353) );
  XNOR U2360 ( .A(n1236), .B(n1232), .Z(n1354) );
  XNOR U2361 ( .A(n1231), .B(n1227), .Z(n1355) );
  XNOR U2362 ( .A(n1226), .B(n1222), .Z(n1356) );
  XNOR U2363 ( .A(n1221), .B(n1217), .Z(n1357) );
  XNOR U2364 ( .A(n1216), .B(n1212), .Z(n1358) );
  XNOR U2365 ( .A(n1211), .B(n1207), .Z(n1359) );
  XNOR U2366 ( .A(n1206), .B(n1202), .Z(n1360) );
  XNOR U2367 ( .A(n1201), .B(n1197), .Z(n1361) );
  XOR U2368 ( .A(n1196), .B(n1193), .Z(n1362) );
  XOR U2369 ( .A(n1363), .B(n1364), .Z(n1193) );
  XOR U2370 ( .A(n1191), .B(n1365), .Z(n1364) );
  XOR U2371 ( .A(n1366), .B(n1367), .Z(n1365) );
  XOR U2372 ( .A(n1368), .B(n1369), .Z(n1367) );
  NAND U2373 ( .A(a[25]), .B(b[30]), .Z(n1369) );
  AND U2374 ( .A(a[24]), .B(b[31]), .Z(n1368) );
  XOR U2375 ( .A(n1370), .B(n1366), .Z(n1363) );
  XOR U2376 ( .A(n1371), .B(n1372), .Z(n1366) );
  NOR U2377 ( .A(n1373), .B(n1374), .Z(n1371) );
  AND U2378 ( .A(a[26]), .B(b[29]), .Z(n1370) );
  XNOR U2379 ( .A(n1375), .B(n1191), .Z(n1192) );
  XOR U2380 ( .A(n1376), .B(n1377), .Z(n1191) );
  ANDN U2381 ( .B(n1378), .A(n1379), .Z(n1376) );
  AND U2382 ( .A(a[27]), .B(b[28]), .Z(n1375) );
  XNOR U2383 ( .A(n1380), .B(n1196), .Z(n1198) );
  XOR U2384 ( .A(n1381), .B(n1382), .Z(n1196) );
  ANDN U2385 ( .B(n1383), .A(n1384), .Z(n1381) );
  AND U2386 ( .A(a[28]), .B(b[27]), .Z(n1380) );
  XNOR U2387 ( .A(n1385), .B(n1201), .Z(n1203) );
  XOR U2388 ( .A(n1386), .B(n1387), .Z(n1201) );
  ANDN U2389 ( .B(n1388), .A(n1389), .Z(n1386) );
  AND U2390 ( .A(b[26]), .B(a[29]), .Z(n1385) );
  XNOR U2391 ( .A(n1390), .B(n1206), .Z(n1208) );
  XOR U2392 ( .A(n1391), .B(n1392), .Z(n1206) );
  ANDN U2393 ( .B(n1393), .A(n1394), .Z(n1391) );
  AND U2394 ( .A(a[30]), .B(b[25]), .Z(n1390) );
  XNOR U2395 ( .A(n1395), .B(n1211), .Z(n1213) );
  XOR U2396 ( .A(n1396), .B(n1397), .Z(n1211) );
  ANDN U2397 ( .B(n1398), .A(n1399), .Z(n1396) );
  AND U2398 ( .A(b[24]), .B(a[31]), .Z(n1395) );
  XNOR U2399 ( .A(n1400), .B(n1216), .Z(n1218) );
  XOR U2400 ( .A(n1401), .B(n1402), .Z(n1216) );
  ANDN U2401 ( .B(n1403), .A(n1404), .Z(n1401) );
  AND U2402 ( .A(a[32]), .B(b[23]), .Z(n1400) );
  XNOR U2403 ( .A(n1405), .B(n1221), .Z(n1223) );
  XOR U2404 ( .A(n1406), .B(n1407), .Z(n1221) );
  ANDN U2405 ( .B(n1408), .A(n1409), .Z(n1406) );
  AND U2406 ( .A(b[22]), .B(a[33]), .Z(n1405) );
  XNOR U2407 ( .A(n1410), .B(n1226), .Z(n1228) );
  XOR U2408 ( .A(n1411), .B(n1412), .Z(n1226) );
  ANDN U2409 ( .B(n1413), .A(n1414), .Z(n1411) );
  AND U2410 ( .A(a[34]), .B(b[21]), .Z(n1410) );
  XNOR U2411 ( .A(n1415), .B(n1231), .Z(n1233) );
  XOR U2412 ( .A(n1416), .B(n1417), .Z(n1231) );
  ANDN U2413 ( .B(n1418), .A(n1419), .Z(n1416) );
  AND U2414 ( .A(b[20]), .B(a[35]), .Z(n1415) );
  XNOR U2415 ( .A(n1420), .B(n1236), .Z(n1238) );
  XOR U2416 ( .A(n1421), .B(n1422), .Z(n1236) );
  ANDN U2417 ( .B(n1423), .A(n1424), .Z(n1421) );
  AND U2418 ( .A(a[36]), .B(b[19]), .Z(n1420) );
  XNOR U2419 ( .A(n1425), .B(n1241), .Z(n1243) );
  XOR U2420 ( .A(n1426), .B(n1427), .Z(n1241) );
  ANDN U2421 ( .B(n1428), .A(n1429), .Z(n1426) );
  AND U2422 ( .A(b[18]), .B(a[37]), .Z(n1425) );
  XNOR U2423 ( .A(n1430), .B(n1246), .Z(n1248) );
  XOR U2424 ( .A(n1431), .B(n1432), .Z(n1246) );
  ANDN U2425 ( .B(n1433), .A(n1434), .Z(n1431) );
  AND U2426 ( .A(a[38]), .B(b[17]), .Z(n1430) );
  XNOR U2427 ( .A(n1435), .B(n1251), .Z(n1253) );
  XOR U2428 ( .A(n1436), .B(n1437), .Z(n1251) );
  ANDN U2429 ( .B(n1438), .A(n1439), .Z(n1436) );
  AND U2430 ( .A(b[16]), .B(a[39]), .Z(n1435) );
  IV U2431 ( .A(n1258), .Z(n1348) );
  XNOR U2432 ( .A(n1440), .B(n1256), .Z(n1258) );
  XOR U2433 ( .A(n1441), .B(n1442), .Z(n1256) );
  ANDN U2434 ( .B(n1443), .A(n1444), .Z(n1441) );
  AND U2435 ( .A(a[40]), .B(b[15]), .Z(n1440) );
  XNOR U2436 ( .A(n1445), .B(n1261), .Z(n1263) );
  XOR U2437 ( .A(n1446), .B(n1447), .Z(n1261) );
  ANDN U2438 ( .B(n1448), .A(n1449), .Z(n1446) );
  AND U2439 ( .A(b[14]), .B(a[41]), .Z(n1445) );
  XNOR U2440 ( .A(n1450), .B(n1266), .Z(n1268) );
  XOR U2441 ( .A(n1451), .B(n1452), .Z(n1266) );
  ANDN U2442 ( .B(n1453), .A(n1454), .Z(n1451) );
  AND U2443 ( .A(a[42]), .B(b[13]), .Z(n1450) );
  XNOR U2444 ( .A(n1455), .B(n1271), .Z(n1273) );
  XOR U2445 ( .A(n1456), .B(n1457), .Z(n1271) );
  ANDN U2446 ( .B(n1458), .A(n1459), .Z(n1456) );
  AND U2447 ( .A(b[12]), .B(a[43]), .Z(n1455) );
  XNOR U2448 ( .A(n1460), .B(n1276), .Z(n1278) );
  XOR U2449 ( .A(n1461), .B(n1462), .Z(n1276) );
  ANDN U2450 ( .B(n1463), .A(n1464), .Z(n1461) );
  AND U2451 ( .A(a[44]), .B(b[11]), .Z(n1460) );
  XNOR U2452 ( .A(n1465), .B(n1281), .Z(n1283) );
  XOR U2453 ( .A(n1466), .B(n1467), .Z(n1281) );
  ANDN U2454 ( .B(n1468), .A(n1469), .Z(n1466) );
  AND U2455 ( .A(b[10]), .B(a[45]), .Z(n1465) );
  XNOR U2456 ( .A(n1470), .B(n1286), .Z(n1288) );
  XOR U2457 ( .A(n1471), .B(n1472), .Z(n1286) );
  ANDN U2458 ( .B(n1473), .A(n1474), .Z(n1471) );
  AND U2459 ( .A(a[46]), .B(b[9]), .Z(n1470) );
  XNOR U2460 ( .A(n1475), .B(n1291), .Z(n1293) );
  XOR U2461 ( .A(n1476), .B(n1477), .Z(n1291) );
  ANDN U2462 ( .B(n1478), .A(n1479), .Z(n1476) );
  AND U2463 ( .A(b[8]), .B(a[47]), .Z(n1475) );
  XNOR U2464 ( .A(n1480), .B(n1296), .Z(n1298) );
  XOR U2465 ( .A(n1481), .B(n1482), .Z(n1296) );
  ANDN U2466 ( .B(n1483), .A(n1484), .Z(n1481) );
  AND U2467 ( .A(a[48]), .B(b[7]), .Z(n1480) );
  XNOR U2468 ( .A(n1485), .B(n1301), .Z(n1303) );
  XOR U2469 ( .A(n1486), .B(n1487), .Z(n1301) );
  ANDN U2470 ( .B(n1488), .A(n1489), .Z(n1486) );
  AND U2471 ( .A(b[6]), .B(a[49]), .Z(n1485) );
  XNOR U2472 ( .A(n1490), .B(n1306), .Z(n1308) );
  XOR U2473 ( .A(n1491), .B(n1492), .Z(n1306) );
  ANDN U2474 ( .B(n1493), .A(n1494), .Z(n1491) );
  AND U2475 ( .A(b[5]), .B(a[50]), .Z(n1490) );
  XNOR U2476 ( .A(n1495), .B(n1311), .Z(n1313) );
  XOR U2477 ( .A(n1496), .B(n1497), .Z(n1311) );
  ANDN U2478 ( .B(n1498), .A(n1499), .Z(n1496) );
  AND U2479 ( .A(b[4]), .B(a[51]), .Z(n1495) );
  XNOR U2480 ( .A(n1500), .B(n1501), .Z(n1325) );
  NANDN U2481 ( .A(n1502), .B(n1503), .Z(n1501) );
  XNOR U2482 ( .A(n1504), .B(n1316), .Z(n1318) );
  XNOR U2483 ( .A(n1505), .B(n1506), .Z(n1316) );
  AND U2484 ( .A(n1507), .B(n1508), .Z(n1505) );
  AND U2485 ( .A(b[3]), .B(a[52]), .Z(n1504) );
  XNOR U2486 ( .A(n1509), .B(n1510), .Z(swire[54]) );
  XOR U2487 ( .A(n1335), .B(n1512), .Z(n1510) );
  XNOR U2488 ( .A(n1334), .B(n1511), .Z(n1512) );
  IV U2489 ( .A(n1509), .Z(n1511) );
  NAND U2490 ( .A(a[54]), .B(b[0]), .Z(n1334) );
  XNOR U2491 ( .A(n1502), .B(n1503), .Z(n1335) );
  XOR U2492 ( .A(n1500), .B(n1513), .Z(n1503) );
  NAND U2493 ( .A(b[1]), .B(a[53]), .Z(n1513) );
  XOR U2494 ( .A(n1508), .B(n1514), .Z(n1502) );
  XOR U2495 ( .A(n1500), .B(n1507), .Z(n1514) );
  XNOR U2496 ( .A(n1515), .B(n1506), .Z(n1507) );
  AND U2497 ( .A(b[2]), .B(a[52]), .Z(n1515) );
  NANDN U2498 ( .A(n1516), .B(n1517), .Z(n1500) );
  XOR U2499 ( .A(n1506), .B(n1498), .Z(n1518) );
  XNOR U2500 ( .A(n1497), .B(n1493), .Z(n1519) );
  XNOR U2501 ( .A(n1492), .B(n1488), .Z(n1520) );
  XNOR U2502 ( .A(n1487), .B(n1483), .Z(n1521) );
  XNOR U2503 ( .A(n1482), .B(n1478), .Z(n1522) );
  XNOR U2504 ( .A(n1477), .B(n1473), .Z(n1523) );
  XNOR U2505 ( .A(n1472), .B(n1468), .Z(n1524) );
  XNOR U2506 ( .A(n1467), .B(n1463), .Z(n1525) );
  XNOR U2507 ( .A(n1462), .B(n1458), .Z(n1526) );
  XNOR U2508 ( .A(n1457), .B(n1453), .Z(n1527) );
  XNOR U2509 ( .A(n1452), .B(n1448), .Z(n1528) );
  XNOR U2510 ( .A(n1447), .B(n1443), .Z(n1529) );
  XNOR U2511 ( .A(n1442), .B(n1438), .Z(n1530) );
  XNOR U2512 ( .A(n1437), .B(n1433), .Z(n1531) );
  XNOR U2513 ( .A(n1432), .B(n1428), .Z(n1532) );
  XNOR U2514 ( .A(n1427), .B(n1423), .Z(n1533) );
  XNOR U2515 ( .A(n1422), .B(n1418), .Z(n1534) );
  XNOR U2516 ( .A(n1417), .B(n1413), .Z(n1535) );
  XNOR U2517 ( .A(n1412), .B(n1408), .Z(n1536) );
  XNOR U2518 ( .A(n1537), .B(n1538), .Z(n1408) );
  XNOR U2519 ( .A(n1407), .B(n1403), .Z(n1538) );
  XNOR U2520 ( .A(n1402), .B(n1398), .Z(n1539) );
  XNOR U2521 ( .A(n1397), .B(n1393), .Z(n1540) );
  XNOR U2522 ( .A(n1392), .B(n1388), .Z(n1541) );
  XNOR U2523 ( .A(n1387), .B(n1383), .Z(n1542) );
  XNOR U2524 ( .A(n1382), .B(n1378), .Z(n1543) );
  XOR U2525 ( .A(n1377), .B(n1374), .Z(n1544) );
  XOR U2526 ( .A(n1545), .B(n1546), .Z(n1374) );
  XOR U2527 ( .A(n1372), .B(n1547), .Z(n1546) );
  XOR U2528 ( .A(n1548), .B(n1549), .Z(n1547) );
  XOR U2529 ( .A(n1550), .B(n1551), .Z(n1549) );
  NAND U2530 ( .A(a[24]), .B(b[30]), .Z(n1551) );
  AND U2531 ( .A(a[23]), .B(b[31]), .Z(n1550) );
  XOR U2532 ( .A(n1552), .B(n1548), .Z(n1545) );
  XOR U2533 ( .A(n1553), .B(n1554), .Z(n1548) );
  NOR U2534 ( .A(n1555), .B(n1556), .Z(n1553) );
  AND U2535 ( .A(a[25]), .B(b[29]), .Z(n1552) );
  XNOR U2536 ( .A(n1557), .B(n1372), .Z(n1373) );
  XOR U2537 ( .A(n1558), .B(n1559), .Z(n1372) );
  ANDN U2538 ( .B(n1560), .A(n1561), .Z(n1558) );
  AND U2539 ( .A(a[26]), .B(b[28]), .Z(n1557) );
  XNOR U2540 ( .A(n1562), .B(n1377), .Z(n1379) );
  XOR U2541 ( .A(n1563), .B(n1564), .Z(n1377) );
  ANDN U2542 ( .B(n1565), .A(n1566), .Z(n1563) );
  AND U2543 ( .A(b[27]), .B(a[27]), .Z(n1562) );
  XNOR U2544 ( .A(n1567), .B(n1382), .Z(n1384) );
  XOR U2545 ( .A(n1568), .B(n1569), .Z(n1382) );
  ANDN U2546 ( .B(n1570), .A(n1571), .Z(n1568) );
  AND U2547 ( .A(a[28]), .B(b[26]), .Z(n1567) );
  XNOR U2548 ( .A(n1572), .B(n1387), .Z(n1389) );
  XOR U2549 ( .A(n1573), .B(n1574), .Z(n1387) );
  ANDN U2550 ( .B(n1575), .A(n1576), .Z(n1573) );
  AND U2551 ( .A(b[25]), .B(a[29]), .Z(n1572) );
  XNOR U2552 ( .A(n1577), .B(n1392), .Z(n1394) );
  XOR U2553 ( .A(n1578), .B(n1579), .Z(n1392) );
  ANDN U2554 ( .B(n1580), .A(n1581), .Z(n1578) );
  AND U2555 ( .A(a[30]), .B(b[24]), .Z(n1577) );
  XNOR U2556 ( .A(n1582), .B(n1397), .Z(n1399) );
  XOR U2557 ( .A(n1583), .B(n1584), .Z(n1397) );
  ANDN U2558 ( .B(n1585), .A(n1586), .Z(n1583) );
  AND U2559 ( .A(b[23]), .B(a[31]), .Z(n1582) );
  IV U2560 ( .A(n1404), .Z(n1537) );
  XNOR U2561 ( .A(n1587), .B(n1402), .Z(n1404) );
  XOR U2562 ( .A(n1588), .B(n1589), .Z(n1402) );
  ANDN U2563 ( .B(n1590), .A(n1591), .Z(n1588) );
  AND U2564 ( .A(a[32]), .B(b[22]), .Z(n1587) );
  XNOR U2565 ( .A(n1592), .B(n1407), .Z(n1409) );
  XOR U2566 ( .A(n1593), .B(n1594), .Z(n1407) );
  ANDN U2567 ( .B(n1595), .A(n1596), .Z(n1593) );
  AND U2568 ( .A(b[21]), .B(a[33]), .Z(n1592) );
  XNOR U2569 ( .A(n1597), .B(n1412), .Z(n1414) );
  XOR U2570 ( .A(n1598), .B(n1599), .Z(n1412) );
  ANDN U2571 ( .B(n1600), .A(n1601), .Z(n1598) );
  AND U2572 ( .A(a[34]), .B(b[20]), .Z(n1597) );
  XNOR U2573 ( .A(n1602), .B(n1417), .Z(n1419) );
  XOR U2574 ( .A(n1603), .B(n1604), .Z(n1417) );
  ANDN U2575 ( .B(n1605), .A(n1606), .Z(n1603) );
  AND U2576 ( .A(b[19]), .B(a[35]), .Z(n1602) );
  XNOR U2577 ( .A(n1607), .B(n1422), .Z(n1424) );
  XOR U2578 ( .A(n1608), .B(n1609), .Z(n1422) );
  ANDN U2579 ( .B(n1610), .A(n1611), .Z(n1608) );
  AND U2580 ( .A(a[36]), .B(b[18]), .Z(n1607) );
  XNOR U2581 ( .A(n1612), .B(n1427), .Z(n1429) );
  XOR U2582 ( .A(n1613), .B(n1614), .Z(n1427) );
  ANDN U2583 ( .B(n1615), .A(n1616), .Z(n1613) );
  AND U2584 ( .A(b[17]), .B(a[37]), .Z(n1612) );
  XNOR U2585 ( .A(n1617), .B(n1432), .Z(n1434) );
  XOR U2586 ( .A(n1618), .B(n1619), .Z(n1432) );
  ANDN U2587 ( .B(n1620), .A(n1621), .Z(n1618) );
  AND U2588 ( .A(a[38]), .B(b[16]), .Z(n1617) );
  XNOR U2589 ( .A(n1622), .B(n1437), .Z(n1439) );
  XOR U2590 ( .A(n1623), .B(n1624), .Z(n1437) );
  ANDN U2591 ( .B(n1625), .A(n1626), .Z(n1623) );
  AND U2592 ( .A(b[15]), .B(a[39]), .Z(n1622) );
  XNOR U2593 ( .A(n1627), .B(n1442), .Z(n1444) );
  XOR U2594 ( .A(n1628), .B(n1629), .Z(n1442) );
  ANDN U2595 ( .B(n1630), .A(n1631), .Z(n1628) );
  AND U2596 ( .A(a[40]), .B(b[14]), .Z(n1627) );
  XNOR U2597 ( .A(n1632), .B(n1447), .Z(n1449) );
  XOR U2598 ( .A(n1633), .B(n1634), .Z(n1447) );
  ANDN U2599 ( .B(n1635), .A(n1636), .Z(n1633) );
  AND U2600 ( .A(b[13]), .B(a[41]), .Z(n1632) );
  XNOR U2601 ( .A(n1637), .B(n1452), .Z(n1454) );
  XOR U2602 ( .A(n1638), .B(n1639), .Z(n1452) );
  ANDN U2603 ( .B(n1640), .A(n1641), .Z(n1638) );
  AND U2604 ( .A(a[42]), .B(b[12]), .Z(n1637) );
  XNOR U2605 ( .A(n1642), .B(n1457), .Z(n1459) );
  XOR U2606 ( .A(n1643), .B(n1644), .Z(n1457) );
  ANDN U2607 ( .B(n1645), .A(n1646), .Z(n1643) );
  AND U2608 ( .A(b[11]), .B(a[43]), .Z(n1642) );
  XNOR U2609 ( .A(n1647), .B(n1462), .Z(n1464) );
  XOR U2610 ( .A(n1648), .B(n1649), .Z(n1462) );
  ANDN U2611 ( .B(n1650), .A(n1651), .Z(n1648) );
  AND U2612 ( .A(a[44]), .B(b[10]), .Z(n1647) );
  XNOR U2613 ( .A(n1652), .B(n1467), .Z(n1469) );
  XOR U2614 ( .A(n1653), .B(n1654), .Z(n1467) );
  ANDN U2615 ( .B(n1655), .A(n1656), .Z(n1653) );
  AND U2616 ( .A(b[9]), .B(a[45]), .Z(n1652) );
  XNOR U2617 ( .A(n1657), .B(n1472), .Z(n1474) );
  XOR U2618 ( .A(n1658), .B(n1659), .Z(n1472) );
  ANDN U2619 ( .B(n1660), .A(n1661), .Z(n1658) );
  AND U2620 ( .A(a[46]), .B(b[8]), .Z(n1657) );
  XNOR U2621 ( .A(n1662), .B(n1477), .Z(n1479) );
  XOR U2622 ( .A(n1663), .B(n1664), .Z(n1477) );
  ANDN U2623 ( .B(n1665), .A(n1666), .Z(n1663) );
  AND U2624 ( .A(b[7]), .B(a[47]), .Z(n1662) );
  XNOR U2625 ( .A(n1667), .B(n1482), .Z(n1484) );
  XOR U2626 ( .A(n1668), .B(n1669), .Z(n1482) );
  ANDN U2627 ( .B(n1670), .A(n1671), .Z(n1668) );
  AND U2628 ( .A(b[6]), .B(a[48]), .Z(n1667) );
  XNOR U2629 ( .A(n1672), .B(n1487), .Z(n1489) );
  XOR U2630 ( .A(n1673), .B(n1674), .Z(n1487) );
  ANDN U2631 ( .B(n1675), .A(n1676), .Z(n1673) );
  AND U2632 ( .A(b[5]), .B(a[49]), .Z(n1672) );
  XNOR U2633 ( .A(n1677), .B(n1492), .Z(n1494) );
  XOR U2634 ( .A(n1678), .B(n1679), .Z(n1492) );
  ANDN U2635 ( .B(n1680), .A(n1681), .Z(n1678) );
  AND U2636 ( .A(b[4]), .B(a[50]), .Z(n1677) );
  XNOR U2637 ( .A(n1682), .B(n1683), .Z(n1506) );
  NANDN U2638 ( .A(n1684), .B(n1685), .Z(n1683) );
  XNOR U2639 ( .A(n1686), .B(n1497), .Z(n1499) );
  XNOR U2640 ( .A(n1687), .B(n1688), .Z(n1497) );
  AND U2641 ( .A(n1689), .B(n1690), .Z(n1687) );
  AND U2642 ( .A(b[3]), .B(a[51]), .Z(n1686) );
  XNOR U2643 ( .A(n1691), .B(n1692), .Z(swire[53]) );
  XOR U2644 ( .A(n1517), .B(n1693), .Z(n1692) );
  XOR U2645 ( .A(n1516), .B(n1691), .Z(n1693) );
  NAND U2646 ( .A(a[53]), .B(b[0]), .Z(n1516) );
  XNOR U2647 ( .A(n1684), .B(n1685), .Z(n1517) );
  XOR U2648 ( .A(n1682), .B(n1694), .Z(n1685) );
  NAND U2649 ( .A(a[52]), .B(b[1]), .Z(n1694) );
  XOR U2650 ( .A(n1690), .B(n1695), .Z(n1684) );
  XOR U2651 ( .A(n1682), .B(n1689), .Z(n1695) );
  XNOR U2652 ( .A(n1696), .B(n1688), .Z(n1689) );
  AND U2653 ( .A(b[2]), .B(a[51]), .Z(n1696) );
  NANDN U2654 ( .A(n1697), .B(n1698), .Z(n1682) );
  XOR U2655 ( .A(n1688), .B(n1680), .Z(n1699) );
  XNOR U2656 ( .A(n1679), .B(n1675), .Z(n1700) );
  XNOR U2657 ( .A(n1674), .B(n1670), .Z(n1701) );
  XNOR U2658 ( .A(n1669), .B(n1665), .Z(n1702) );
  XNOR U2659 ( .A(n1664), .B(n1660), .Z(n1703) );
  XNOR U2660 ( .A(n1659), .B(n1655), .Z(n1704) );
  XNOR U2661 ( .A(n1654), .B(n1650), .Z(n1705) );
  XNOR U2662 ( .A(n1649), .B(n1645), .Z(n1706) );
  XNOR U2663 ( .A(n1644), .B(n1640), .Z(n1707) );
  XNOR U2664 ( .A(n1639), .B(n1635), .Z(n1708) );
  XNOR U2665 ( .A(n1634), .B(n1630), .Z(n1709) );
  XNOR U2666 ( .A(n1629), .B(n1625), .Z(n1710) );
  XNOR U2667 ( .A(n1624), .B(n1620), .Z(n1711) );
  XNOR U2668 ( .A(n1619), .B(n1615), .Z(n1712) );
  XNOR U2669 ( .A(n1614), .B(n1610), .Z(n1713) );
  XNOR U2670 ( .A(n1714), .B(n1715), .Z(n1610) );
  XNOR U2671 ( .A(n1609), .B(n1605), .Z(n1715) );
  XNOR U2672 ( .A(n1604), .B(n1600), .Z(n1716) );
  XNOR U2673 ( .A(n1599), .B(n1595), .Z(n1717) );
  XNOR U2674 ( .A(n1594), .B(n1590), .Z(n1718) );
  XNOR U2675 ( .A(n1589), .B(n1585), .Z(n1719) );
  XNOR U2676 ( .A(n1720), .B(n1721), .Z(n1585) );
  XNOR U2677 ( .A(n1584), .B(n1580), .Z(n1721) );
  XNOR U2678 ( .A(n1579), .B(n1575), .Z(n1722) );
  XNOR U2679 ( .A(n1574), .B(n1570), .Z(n1723) );
  XNOR U2680 ( .A(n1569), .B(n1565), .Z(n1724) );
  XNOR U2681 ( .A(n1564), .B(n1560), .Z(n1725) );
  XOR U2682 ( .A(n1559), .B(n1556), .Z(n1726) );
  XOR U2683 ( .A(n1727), .B(n1728), .Z(n1556) );
  XOR U2684 ( .A(n1554), .B(n1729), .Z(n1728) );
  XOR U2685 ( .A(n1730), .B(n1731), .Z(n1729) );
  XOR U2686 ( .A(n1732), .B(n1733), .Z(n1731) );
  NAND U2687 ( .A(a[23]), .B(b[30]), .Z(n1733) );
  AND U2688 ( .A(a[22]), .B(b[31]), .Z(n1732) );
  XOR U2689 ( .A(n1734), .B(n1730), .Z(n1727) );
  XOR U2690 ( .A(n1735), .B(n1736), .Z(n1730) );
  NOR U2691 ( .A(n1737), .B(n1738), .Z(n1735) );
  AND U2692 ( .A(a[24]), .B(b[29]), .Z(n1734) );
  XNOR U2693 ( .A(n1739), .B(n1554), .Z(n1555) );
  XOR U2694 ( .A(n1740), .B(n1741), .Z(n1554) );
  ANDN U2695 ( .B(n1742), .A(n1743), .Z(n1740) );
  AND U2696 ( .A(a[25]), .B(b[28]), .Z(n1739) );
  XNOR U2697 ( .A(n1744), .B(n1559), .Z(n1561) );
  XOR U2698 ( .A(n1745), .B(n1746), .Z(n1559) );
  ANDN U2699 ( .B(n1747), .A(n1748), .Z(n1745) );
  AND U2700 ( .A(a[26]), .B(b[27]), .Z(n1744) );
  XNOR U2701 ( .A(n1749), .B(n1564), .Z(n1566) );
  XOR U2702 ( .A(n1750), .B(n1751), .Z(n1564) );
  ANDN U2703 ( .B(n1752), .A(n1753), .Z(n1750) );
  AND U2704 ( .A(b[26]), .B(a[27]), .Z(n1749) );
  XNOR U2705 ( .A(n1754), .B(n1569), .Z(n1571) );
  XOR U2706 ( .A(n1755), .B(n1756), .Z(n1569) );
  ANDN U2707 ( .B(n1757), .A(n1758), .Z(n1755) );
  AND U2708 ( .A(a[28]), .B(b[25]), .Z(n1754) );
  XNOR U2709 ( .A(n1759), .B(n1574), .Z(n1576) );
  XOR U2710 ( .A(n1760), .B(n1761), .Z(n1574) );
  ANDN U2711 ( .B(n1762), .A(n1763), .Z(n1760) );
  AND U2712 ( .A(b[24]), .B(a[29]), .Z(n1759) );
  IV U2713 ( .A(n1581), .Z(n1720) );
  XNOR U2714 ( .A(n1764), .B(n1579), .Z(n1581) );
  XOR U2715 ( .A(n1765), .B(n1766), .Z(n1579) );
  ANDN U2716 ( .B(n1767), .A(n1768), .Z(n1765) );
  AND U2717 ( .A(a[30]), .B(b[23]), .Z(n1764) );
  XNOR U2718 ( .A(n1769), .B(n1584), .Z(n1586) );
  XOR U2719 ( .A(n1770), .B(n1771), .Z(n1584) );
  ANDN U2720 ( .B(n1772), .A(n1773), .Z(n1770) );
  AND U2721 ( .A(b[22]), .B(a[31]), .Z(n1769) );
  XNOR U2722 ( .A(n1774), .B(n1589), .Z(n1591) );
  XOR U2723 ( .A(n1775), .B(n1776), .Z(n1589) );
  ANDN U2724 ( .B(n1777), .A(n1778), .Z(n1775) );
  AND U2725 ( .A(a[32]), .B(b[21]), .Z(n1774) );
  XNOR U2726 ( .A(n1779), .B(n1594), .Z(n1596) );
  XOR U2727 ( .A(n1780), .B(n1781), .Z(n1594) );
  ANDN U2728 ( .B(n1782), .A(n1783), .Z(n1780) );
  AND U2729 ( .A(b[20]), .B(a[33]), .Z(n1779) );
  XNOR U2730 ( .A(n1784), .B(n1599), .Z(n1601) );
  XOR U2731 ( .A(n1785), .B(n1786), .Z(n1599) );
  ANDN U2732 ( .B(n1787), .A(n1788), .Z(n1785) );
  AND U2733 ( .A(a[34]), .B(b[19]), .Z(n1784) );
  IV U2734 ( .A(n1606), .Z(n1714) );
  XNOR U2735 ( .A(n1789), .B(n1604), .Z(n1606) );
  XOR U2736 ( .A(n1790), .B(n1791), .Z(n1604) );
  ANDN U2737 ( .B(n1792), .A(n1793), .Z(n1790) );
  AND U2738 ( .A(b[18]), .B(a[35]), .Z(n1789) );
  XNOR U2739 ( .A(n1794), .B(n1609), .Z(n1611) );
  XOR U2740 ( .A(n1795), .B(n1796), .Z(n1609) );
  ANDN U2741 ( .B(n1797), .A(n1798), .Z(n1795) );
  AND U2742 ( .A(a[36]), .B(b[17]), .Z(n1794) );
  XNOR U2743 ( .A(n1799), .B(n1614), .Z(n1616) );
  XOR U2744 ( .A(n1800), .B(n1801), .Z(n1614) );
  ANDN U2745 ( .B(n1802), .A(n1803), .Z(n1800) );
  AND U2746 ( .A(b[16]), .B(a[37]), .Z(n1799) );
  XNOR U2747 ( .A(n1804), .B(n1619), .Z(n1621) );
  XOR U2748 ( .A(n1805), .B(n1806), .Z(n1619) );
  ANDN U2749 ( .B(n1807), .A(n1808), .Z(n1805) );
  AND U2750 ( .A(a[38]), .B(b[15]), .Z(n1804) );
  XNOR U2751 ( .A(n1809), .B(n1624), .Z(n1626) );
  XOR U2752 ( .A(n1810), .B(n1811), .Z(n1624) );
  ANDN U2753 ( .B(n1812), .A(n1813), .Z(n1810) );
  AND U2754 ( .A(b[14]), .B(a[39]), .Z(n1809) );
  XNOR U2755 ( .A(n1814), .B(n1629), .Z(n1631) );
  XOR U2756 ( .A(n1815), .B(n1816), .Z(n1629) );
  ANDN U2757 ( .B(n1817), .A(n1818), .Z(n1815) );
  AND U2758 ( .A(a[40]), .B(b[13]), .Z(n1814) );
  XNOR U2759 ( .A(n1819), .B(n1634), .Z(n1636) );
  XOR U2760 ( .A(n1820), .B(n1821), .Z(n1634) );
  ANDN U2761 ( .B(n1822), .A(n1823), .Z(n1820) );
  AND U2762 ( .A(b[12]), .B(a[41]), .Z(n1819) );
  XNOR U2763 ( .A(n1824), .B(n1639), .Z(n1641) );
  XOR U2764 ( .A(n1825), .B(n1826), .Z(n1639) );
  ANDN U2765 ( .B(n1827), .A(n1828), .Z(n1825) );
  AND U2766 ( .A(a[42]), .B(b[11]), .Z(n1824) );
  XNOR U2767 ( .A(n1829), .B(n1644), .Z(n1646) );
  XOR U2768 ( .A(n1830), .B(n1831), .Z(n1644) );
  ANDN U2769 ( .B(n1832), .A(n1833), .Z(n1830) );
  AND U2770 ( .A(b[10]), .B(a[43]), .Z(n1829) );
  XNOR U2771 ( .A(n1834), .B(n1649), .Z(n1651) );
  XOR U2772 ( .A(n1835), .B(n1836), .Z(n1649) );
  ANDN U2773 ( .B(n1837), .A(n1838), .Z(n1835) );
  AND U2774 ( .A(a[44]), .B(b[9]), .Z(n1834) );
  XNOR U2775 ( .A(n1839), .B(n1654), .Z(n1656) );
  XOR U2776 ( .A(n1840), .B(n1841), .Z(n1654) );
  ANDN U2777 ( .B(n1842), .A(n1843), .Z(n1840) );
  AND U2778 ( .A(b[8]), .B(a[45]), .Z(n1839) );
  XNOR U2779 ( .A(n1844), .B(n1659), .Z(n1661) );
  XOR U2780 ( .A(n1845), .B(n1846), .Z(n1659) );
  ANDN U2781 ( .B(n1847), .A(n1848), .Z(n1845) );
  AND U2782 ( .A(a[46]), .B(b[7]), .Z(n1844) );
  XNOR U2783 ( .A(n1849), .B(n1664), .Z(n1666) );
  XOR U2784 ( .A(n1850), .B(n1851), .Z(n1664) );
  ANDN U2785 ( .B(n1852), .A(n1853), .Z(n1850) );
  AND U2786 ( .A(b[6]), .B(a[47]), .Z(n1849) );
  XNOR U2787 ( .A(n1854), .B(n1669), .Z(n1671) );
  XOR U2788 ( .A(n1855), .B(n1856), .Z(n1669) );
  ANDN U2789 ( .B(n1857), .A(n1858), .Z(n1855) );
  AND U2790 ( .A(b[5]), .B(a[48]), .Z(n1854) );
  XNOR U2791 ( .A(n1859), .B(n1674), .Z(n1676) );
  XOR U2792 ( .A(n1860), .B(n1861), .Z(n1674) );
  ANDN U2793 ( .B(n1862), .A(n1863), .Z(n1860) );
  AND U2794 ( .A(b[4]), .B(a[49]), .Z(n1859) );
  XNOR U2795 ( .A(n1864), .B(n1865), .Z(n1688) );
  NANDN U2796 ( .A(n1866), .B(n1867), .Z(n1865) );
  XNOR U2797 ( .A(n1868), .B(n1679), .Z(n1681) );
  XNOR U2798 ( .A(n1869), .B(n1870), .Z(n1679) );
  AND U2799 ( .A(n1871), .B(n1872), .Z(n1869) );
  AND U2800 ( .A(b[3]), .B(a[50]), .Z(n1868) );
  XNOR U2801 ( .A(n1873), .B(n1874), .Z(swire[52]) );
  XOR U2802 ( .A(n1698), .B(n1876), .Z(n1874) );
  XNOR U2803 ( .A(n1697), .B(n1875), .Z(n1876) );
  IV U2804 ( .A(n1873), .Z(n1875) );
  NAND U2805 ( .A(a[52]), .B(b[0]), .Z(n1697) );
  XNOR U2806 ( .A(n1866), .B(n1867), .Z(n1698) );
  XOR U2807 ( .A(n1864), .B(n1877), .Z(n1867) );
  NAND U2808 ( .A(b[1]), .B(a[51]), .Z(n1877) );
  XOR U2809 ( .A(n1872), .B(n1878), .Z(n1866) );
  XOR U2810 ( .A(n1864), .B(n1871), .Z(n1878) );
  XNOR U2811 ( .A(n1879), .B(n1870), .Z(n1871) );
  AND U2812 ( .A(b[2]), .B(a[50]), .Z(n1879) );
  NANDN U2813 ( .A(n1880), .B(n1881), .Z(n1864) );
  XOR U2814 ( .A(n1870), .B(n1862), .Z(n1882) );
  XNOR U2815 ( .A(n1861), .B(n1857), .Z(n1883) );
  XNOR U2816 ( .A(n1856), .B(n1852), .Z(n1884) );
  XNOR U2817 ( .A(n1851), .B(n1847), .Z(n1885) );
  XNOR U2818 ( .A(n1846), .B(n1842), .Z(n1886) );
  XNOR U2819 ( .A(n1841), .B(n1837), .Z(n1887) );
  XNOR U2820 ( .A(n1836), .B(n1832), .Z(n1888) );
  XNOR U2821 ( .A(n1831), .B(n1827), .Z(n1889) );
  XNOR U2822 ( .A(n1826), .B(n1822), .Z(n1890) );
  XNOR U2823 ( .A(n1821), .B(n1817), .Z(n1891) );
  XNOR U2824 ( .A(n1816), .B(n1812), .Z(n1892) );
  XNOR U2825 ( .A(n1811), .B(n1807), .Z(n1893) );
  XNOR U2826 ( .A(n1806), .B(n1802), .Z(n1894) );
  XNOR U2827 ( .A(n1801), .B(n1797), .Z(n1895) );
  XNOR U2828 ( .A(n1796), .B(n1792), .Z(n1896) );
  XNOR U2829 ( .A(n1791), .B(n1787), .Z(n1897) );
  XNOR U2830 ( .A(n1786), .B(n1782), .Z(n1898) );
  XNOR U2831 ( .A(n1781), .B(n1777), .Z(n1899) );
  XNOR U2832 ( .A(n1776), .B(n1772), .Z(n1900) );
  XNOR U2833 ( .A(n1771), .B(n1767), .Z(n1901) );
  XNOR U2834 ( .A(n1766), .B(n1762), .Z(n1902) );
  XNOR U2835 ( .A(n1761), .B(n1757), .Z(n1903) );
  XNOR U2836 ( .A(n1756), .B(n1752), .Z(n1904) );
  XNOR U2837 ( .A(n1751), .B(n1747), .Z(n1905) );
  XNOR U2838 ( .A(n1746), .B(n1742), .Z(n1906) );
  XOR U2839 ( .A(n1741), .B(n1738), .Z(n1907) );
  XOR U2840 ( .A(n1908), .B(n1909), .Z(n1738) );
  XOR U2841 ( .A(n1736), .B(n1910), .Z(n1909) );
  XOR U2842 ( .A(n1911), .B(n1912), .Z(n1910) );
  XOR U2843 ( .A(n1913), .B(n1914), .Z(n1912) );
  NAND U2844 ( .A(a[22]), .B(b[30]), .Z(n1914) );
  AND U2845 ( .A(a[21]), .B(b[31]), .Z(n1913) );
  XOR U2846 ( .A(n1915), .B(n1911), .Z(n1908) );
  XOR U2847 ( .A(n1916), .B(n1917), .Z(n1911) );
  NOR U2848 ( .A(n1918), .B(n1919), .Z(n1916) );
  AND U2849 ( .A(a[23]), .B(b[29]), .Z(n1915) );
  XNOR U2850 ( .A(n1920), .B(n1736), .Z(n1737) );
  XOR U2851 ( .A(n1921), .B(n1922), .Z(n1736) );
  ANDN U2852 ( .B(n1923), .A(n1924), .Z(n1921) );
  AND U2853 ( .A(a[24]), .B(b[28]), .Z(n1920) );
  XNOR U2854 ( .A(n1925), .B(n1741), .Z(n1743) );
  XOR U2855 ( .A(n1926), .B(n1927), .Z(n1741) );
  ANDN U2856 ( .B(n1928), .A(n1929), .Z(n1926) );
  AND U2857 ( .A(a[25]), .B(b[27]), .Z(n1925) );
  XNOR U2858 ( .A(n1930), .B(n1746), .Z(n1748) );
  XOR U2859 ( .A(n1931), .B(n1932), .Z(n1746) );
  ANDN U2860 ( .B(n1933), .A(n1934), .Z(n1931) );
  AND U2861 ( .A(a[26]), .B(b[26]), .Z(n1930) );
  XNOR U2862 ( .A(n1935), .B(n1751), .Z(n1753) );
  XOR U2863 ( .A(n1936), .B(n1937), .Z(n1751) );
  ANDN U2864 ( .B(n1938), .A(n1939), .Z(n1936) );
  AND U2865 ( .A(b[25]), .B(a[27]), .Z(n1935) );
  XNOR U2866 ( .A(n1940), .B(n1756), .Z(n1758) );
  XOR U2867 ( .A(n1941), .B(n1942), .Z(n1756) );
  ANDN U2868 ( .B(n1943), .A(n1944), .Z(n1941) );
  AND U2869 ( .A(a[28]), .B(b[24]), .Z(n1940) );
  XNOR U2870 ( .A(n1945), .B(n1761), .Z(n1763) );
  XOR U2871 ( .A(n1946), .B(n1947), .Z(n1761) );
  ANDN U2872 ( .B(n1948), .A(n1949), .Z(n1946) );
  AND U2873 ( .A(b[23]), .B(a[29]), .Z(n1945) );
  XNOR U2874 ( .A(n1950), .B(n1766), .Z(n1768) );
  XOR U2875 ( .A(n1951), .B(n1952), .Z(n1766) );
  ANDN U2876 ( .B(n1953), .A(n1954), .Z(n1951) );
  AND U2877 ( .A(a[30]), .B(b[22]), .Z(n1950) );
  XNOR U2878 ( .A(n1955), .B(n1771), .Z(n1773) );
  XOR U2879 ( .A(n1956), .B(n1957), .Z(n1771) );
  ANDN U2880 ( .B(n1958), .A(n1959), .Z(n1956) );
  AND U2881 ( .A(b[21]), .B(a[31]), .Z(n1955) );
  XNOR U2882 ( .A(n1960), .B(n1776), .Z(n1778) );
  XOR U2883 ( .A(n1961), .B(n1962), .Z(n1776) );
  ANDN U2884 ( .B(n1963), .A(n1964), .Z(n1961) );
  AND U2885 ( .A(a[32]), .B(b[20]), .Z(n1960) );
  XNOR U2886 ( .A(n1965), .B(n1781), .Z(n1783) );
  XOR U2887 ( .A(n1966), .B(n1967), .Z(n1781) );
  ANDN U2888 ( .B(n1968), .A(n1969), .Z(n1966) );
  AND U2889 ( .A(b[19]), .B(a[33]), .Z(n1965) );
  XNOR U2890 ( .A(n1970), .B(n1786), .Z(n1788) );
  XOR U2891 ( .A(n1971), .B(n1972), .Z(n1786) );
  ANDN U2892 ( .B(n1973), .A(n1974), .Z(n1971) );
  AND U2893 ( .A(a[34]), .B(b[18]), .Z(n1970) );
  XNOR U2894 ( .A(n1975), .B(n1791), .Z(n1793) );
  XOR U2895 ( .A(n1976), .B(n1977), .Z(n1791) );
  ANDN U2896 ( .B(n1978), .A(n1979), .Z(n1976) );
  AND U2897 ( .A(b[17]), .B(a[35]), .Z(n1975) );
  XNOR U2898 ( .A(n1980), .B(n1796), .Z(n1798) );
  XOR U2899 ( .A(n1981), .B(n1982), .Z(n1796) );
  ANDN U2900 ( .B(n1983), .A(n1984), .Z(n1981) );
  AND U2901 ( .A(a[36]), .B(b[16]), .Z(n1980) );
  XNOR U2902 ( .A(n1985), .B(n1801), .Z(n1803) );
  XOR U2903 ( .A(n1986), .B(n1987), .Z(n1801) );
  ANDN U2904 ( .B(n1988), .A(n1989), .Z(n1986) );
  AND U2905 ( .A(b[15]), .B(a[37]), .Z(n1985) );
  XNOR U2906 ( .A(n1990), .B(n1806), .Z(n1808) );
  XOR U2907 ( .A(n1991), .B(n1992), .Z(n1806) );
  ANDN U2908 ( .B(n1993), .A(n1994), .Z(n1991) );
  AND U2909 ( .A(a[38]), .B(b[14]), .Z(n1990) );
  XNOR U2910 ( .A(n1995), .B(n1811), .Z(n1813) );
  XOR U2911 ( .A(n1996), .B(n1997), .Z(n1811) );
  ANDN U2912 ( .B(n1998), .A(n1999), .Z(n1996) );
  AND U2913 ( .A(b[13]), .B(a[39]), .Z(n1995) );
  XNOR U2914 ( .A(n2000), .B(n1816), .Z(n1818) );
  XOR U2915 ( .A(n2001), .B(n2002), .Z(n1816) );
  ANDN U2916 ( .B(n2003), .A(n2004), .Z(n2001) );
  AND U2917 ( .A(a[40]), .B(b[12]), .Z(n2000) );
  XNOR U2918 ( .A(n2005), .B(n1821), .Z(n1823) );
  XOR U2919 ( .A(n2006), .B(n2007), .Z(n1821) );
  ANDN U2920 ( .B(n2008), .A(n2009), .Z(n2006) );
  AND U2921 ( .A(b[11]), .B(a[41]), .Z(n2005) );
  XNOR U2922 ( .A(n2010), .B(n1826), .Z(n1828) );
  XOR U2923 ( .A(n2011), .B(n2012), .Z(n1826) );
  ANDN U2924 ( .B(n2013), .A(n2014), .Z(n2011) );
  AND U2925 ( .A(a[42]), .B(b[10]), .Z(n2010) );
  XNOR U2926 ( .A(n2015), .B(n1831), .Z(n1833) );
  XOR U2927 ( .A(n2016), .B(n2017), .Z(n1831) );
  ANDN U2928 ( .B(n2018), .A(n2019), .Z(n2016) );
  AND U2929 ( .A(b[9]), .B(a[43]), .Z(n2015) );
  XNOR U2930 ( .A(n2020), .B(n1836), .Z(n1838) );
  XOR U2931 ( .A(n2021), .B(n2022), .Z(n1836) );
  ANDN U2932 ( .B(n2023), .A(n2024), .Z(n2021) );
  AND U2933 ( .A(a[44]), .B(b[8]), .Z(n2020) );
  XNOR U2934 ( .A(n2025), .B(n1841), .Z(n1843) );
  XOR U2935 ( .A(n2026), .B(n2027), .Z(n1841) );
  ANDN U2936 ( .B(n2028), .A(n2029), .Z(n2026) );
  AND U2937 ( .A(b[7]), .B(a[45]), .Z(n2025) );
  XNOR U2938 ( .A(n2030), .B(n1846), .Z(n1848) );
  XOR U2939 ( .A(n2031), .B(n2032), .Z(n1846) );
  ANDN U2940 ( .B(n2033), .A(n2034), .Z(n2031) );
  AND U2941 ( .A(b[6]), .B(a[46]), .Z(n2030) );
  XNOR U2942 ( .A(n2035), .B(n1851), .Z(n1853) );
  XOR U2943 ( .A(n2036), .B(n2037), .Z(n1851) );
  ANDN U2944 ( .B(n2038), .A(n2039), .Z(n2036) );
  AND U2945 ( .A(b[5]), .B(a[47]), .Z(n2035) );
  XNOR U2946 ( .A(n2040), .B(n1856), .Z(n1858) );
  XOR U2947 ( .A(n2041), .B(n2042), .Z(n1856) );
  ANDN U2948 ( .B(n2043), .A(n2044), .Z(n2041) );
  AND U2949 ( .A(b[4]), .B(a[48]), .Z(n2040) );
  XNOR U2950 ( .A(n2045), .B(n2046), .Z(n1870) );
  NANDN U2951 ( .A(n2047), .B(n2048), .Z(n2046) );
  XNOR U2952 ( .A(n2049), .B(n1861), .Z(n1863) );
  XNOR U2953 ( .A(n2050), .B(n2051), .Z(n1861) );
  AND U2954 ( .A(n2052), .B(n2053), .Z(n2050) );
  AND U2955 ( .A(b[3]), .B(a[49]), .Z(n2049) );
  XNOR U2956 ( .A(n2054), .B(n2055), .Z(swire[51]) );
  XOR U2957 ( .A(n1881), .B(n2056), .Z(n2055) );
  XOR U2958 ( .A(n1880), .B(n2054), .Z(n2056) );
  NAND U2959 ( .A(a[51]), .B(b[0]), .Z(n1880) );
  XNOR U2960 ( .A(n2047), .B(n2048), .Z(n1881) );
  XOR U2961 ( .A(n2045), .B(n2057), .Z(n2048) );
  NAND U2962 ( .A(a[50]), .B(b[1]), .Z(n2057) );
  XOR U2963 ( .A(n2053), .B(n2058), .Z(n2047) );
  XOR U2964 ( .A(n2045), .B(n2052), .Z(n2058) );
  XNOR U2965 ( .A(n2059), .B(n2051), .Z(n2052) );
  AND U2966 ( .A(b[2]), .B(a[49]), .Z(n2059) );
  NANDN U2967 ( .A(n2060), .B(n2061), .Z(n2045) );
  XOR U2968 ( .A(n2051), .B(n2043), .Z(n2062) );
  XNOR U2969 ( .A(n2042), .B(n2038), .Z(n2063) );
  XNOR U2970 ( .A(n2037), .B(n2033), .Z(n2064) );
  XNOR U2971 ( .A(n2032), .B(n2028), .Z(n2065) );
  XNOR U2972 ( .A(n2027), .B(n2023), .Z(n2066) );
  XNOR U2973 ( .A(n2022), .B(n2018), .Z(n2067) );
  XNOR U2974 ( .A(n2017), .B(n2013), .Z(n2068) );
  XNOR U2975 ( .A(n2012), .B(n2008), .Z(n2069) );
  XNOR U2976 ( .A(n2007), .B(n2003), .Z(n2070) );
  XNOR U2977 ( .A(n2002), .B(n1998), .Z(n2071) );
  XNOR U2978 ( .A(n1997), .B(n1993), .Z(n2072) );
  XNOR U2979 ( .A(n1992), .B(n1988), .Z(n2073) );
  XNOR U2980 ( .A(n1987), .B(n1983), .Z(n2074) );
  XNOR U2981 ( .A(n1982), .B(n1978), .Z(n2075) );
  XNOR U2982 ( .A(n1977), .B(n1973), .Z(n2076) );
  XNOR U2983 ( .A(n1972), .B(n1968), .Z(n2077) );
  XNOR U2984 ( .A(n1967), .B(n1963), .Z(n2078) );
  XNOR U2985 ( .A(n1962), .B(n1958), .Z(n2079) );
  XNOR U2986 ( .A(n1957), .B(n1953), .Z(n2080) );
  XNOR U2987 ( .A(n1952), .B(n1948), .Z(n2081) );
  XNOR U2988 ( .A(n1947), .B(n1943), .Z(n2082) );
  XNOR U2989 ( .A(n1942), .B(n1938), .Z(n2083) );
  XNOR U2990 ( .A(n1937), .B(n1933), .Z(n2084) );
  XNOR U2991 ( .A(n1932), .B(n1928), .Z(n2085) );
  XNOR U2992 ( .A(n1927), .B(n1923), .Z(n2086) );
  XOR U2993 ( .A(n1922), .B(n1919), .Z(n2087) );
  XOR U2994 ( .A(n2088), .B(n2089), .Z(n1919) );
  XOR U2995 ( .A(n1917), .B(n2090), .Z(n2089) );
  XOR U2996 ( .A(n2091), .B(n2092), .Z(n2090) );
  XOR U2997 ( .A(n2093), .B(n2094), .Z(n2092) );
  NAND U2998 ( .A(a[21]), .B(b[30]), .Z(n2094) );
  AND U2999 ( .A(a[20]), .B(b[31]), .Z(n2093) );
  XOR U3000 ( .A(n2095), .B(n2091), .Z(n2088) );
  XOR U3001 ( .A(n2096), .B(n2097), .Z(n2091) );
  NOR U3002 ( .A(n2098), .B(n2099), .Z(n2096) );
  AND U3003 ( .A(a[22]), .B(b[29]), .Z(n2095) );
  XNOR U3004 ( .A(n2100), .B(n1917), .Z(n1918) );
  XOR U3005 ( .A(n2101), .B(n2102), .Z(n1917) );
  ANDN U3006 ( .B(n2103), .A(n2104), .Z(n2101) );
  AND U3007 ( .A(a[23]), .B(b[28]), .Z(n2100) );
  XNOR U3008 ( .A(n2105), .B(n1922), .Z(n1924) );
  XOR U3009 ( .A(n2106), .B(n2107), .Z(n1922) );
  ANDN U3010 ( .B(n2108), .A(n2109), .Z(n2106) );
  AND U3011 ( .A(a[24]), .B(b[27]), .Z(n2105) );
  XNOR U3012 ( .A(n2110), .B(n1927), .Z(n1929) );
  XOR U3013 ( .A(n2111), .B(n2112), .Z(n1927) );
  ANDN U3014 ( .B(n2113), .A(n2114), .Z(n2111) );
  AND U3015 ( .A(a[25]), .B(b[26]), .Z(n2110) );
  XNOR U3016 ( .A(n2115), .B(n1932), .Z(n1934) );
  XOR U3017 ( .A(n2116), .B(n2117), .Z(n1932) );
  ANDN U3018 ( .B(n2118), .A(n2119), .Z(n2116) );
  AND U3019 ( .A(a[26]), .B(b[25]), .Z(n2115) );
  XNOR U3020 ( .A(n2120), .B(n1937), .Z(n1939) );
  XOR U3021 ( .A(n2121), .B(n2122), .Z(n1937) );
  ANDN U3022 ( .B(n2123), .A(n2124), .Z(n2121) );
  AND U3023 ( .A(b[24]), .B(a[27]), .Z(n2120) );
  XNOR U3024 ( .A(n2125), .B(n1942), .Z(n1944) );
  XOR U3025 ( .A(n2126), .B(n2127), .Z(n1942) );
  ANDN U3026 ( .B(n2128), .A(n2129), .Z(n2126) );
  AND U3027 ( .A(a[28]), .B(b[23]), .Z(n2125) );
  XNOR U3028 ( .A(n2130), .B(n1947), .Z(n1949) );
  XOR U3029 ( .A(n2131), .B(n2132), .Z(n1947) );
  ANDN U3030 ( .B(n2133), .A(n2134), .Z(n2131) );
  AND U3031 ( .A(b[22]), .B(a[29]), .Z(n2130) );
  XNOR U3032 ( .A(n2135), .B(n1952), .Z(n1954) );
  XOR U3033 ( .A(n2136), .B(n2137), .Z(n1952) );
  ANDN U3034 ( .B(n2138), .A(n2139), .Z(n2136) );
  AND U3035 ( .A(a[30]), .B(b[21]), .Z(n2135) );
  XNOR U3036 ( .A(n2140), .B(n1957), .Z(n1959) );
  XOR U3037 ( .A(n2141), .B(n2142), .Z(n1957) );
  ANDN U3038 ( .B(n2143), .A(n2144), .Z(n2141) );
  AND U3039 ( .A(b[20]), .B(a[31]), .Z(n2140) );
  XNOR U3040 ( .A(n2145), .B(n1962), .Z(n1964) );
  XOR U3041 ( .A(n2146), .B(n2147), .Z(n1962) );
  ANDN U3042 ( .B(n2148), .A(n2149), .Z(n2146) );
  AND U3043 ( .A(a[32]), .B(b[19]), .Z(n2145) );
  XNOR U3044 ( .A(n2150), .B(n1967), .Z(n1969) );
  XOR U3045 ( .A(n2151), .B(n2152), .Z(n1967) );
  ANDN U3046 ( .B(n2153), .A(n2154), .Z(n2151) );
  AND U3047 ( .A(b[18]), .B(a[33]), .Z(n2150) );
  XNOR U3048 ( .A(n2155), .B(n1972), .Z(n1974) );
  XOR U3049 ( .A(n2156), .B(n2157), .Z(n1972) );
  ANDN U3050 ( .B(n2158), .A(n2159), .Z(n2156) );
  AND U3051 ( .A(a[34]), .B(b[17]), .Z(n2155) );
  XNOR U3052 ( .A(n2160), .B(n1977), .Z(n1979) );
  XOR U3053 ( .A(n2161), .B(n2162), .Z(n1977) );
  ANDN U3054 ( .B(n2163), .A(n2164), .Z(n2161) );
  AND U3055 ( .A(b[16]), .B(a[35]), .Z(n2160) );
  XNOR U3056 ( .A(n2165), .B(n1982), .Z(n1984) );
  XOR U3057 ( .A(n2166), .B(n2167), .Z(n1982) );
  ANDN U3058 ( .B(n2168), .A(n2169), .Z(n2166) );
  AND U3059 ( .A(a[36]), .B(b[15]), .Z(n2165) );
  XNOR U3060 ( .A(n2170), .B(n1987), .Z(n1989) );
  XOR U3061 ( .A(n2171), .B(n2172), .Z(n1987) );
  ANDN U3062 ( .B(n2173), .A(n2174), .Z(n2171) );
  AND U3063 ( .A(b[14]), .B(a[37]), .Z(n2170) );
  XNOR U3064 ( .A(n2175), .B(n1992), .Z(n1994) );
  XOR U3065 ( .A(n2176), .B(n2177), .Z(n1992) );
  ANDN U3066 ( .B(n2178), .A(n2179), .Z(n2176) );
  AND U3067 ( .A(a[38]), .B(b[13]), .Z(n2175) );
  XNOR U3068 ( .A(n2180), .B(n1997), .Z(n1999) );
  XOR U3069 ( .A(n2181), .B(n2182), .Z(n1997) );
  ANDN U3070 ( .B(n2183), .A(n2184), .Z(n2181) );
  AND U3071 ( .A(b[12]), .B(a[39]), .Z(n2180) );
  XNOR U3072 ( .A(n2185), .B(n2002), .Z(n2004) );
  XOR U3073 ( .A(n2186), .B(n2187), .Z(n2002) );
  ANDN U3074 ( .B(n2188), .A(n2189), .Z(n2186) );
  AND U3075 ( .A(a[40]), .B(b[11]), .Z(n2185) );
  XNOR U3076 ( .A(n2190), .B(n2007), .Z(n2009) );
  XOR U3077 ( .A(n2191), .B(n2192), .Z(n2007) );
  ANDN U3078 ( .B(n2193), .A(n2194), .Z(n2191) );
  AND U3079 ( .A(b[10]), .B(a[41]), .Z(n2190) );
  XNOR U3080 ( .A(n2195), .B(n2012), .Z(n2014) );
  XOR U3081 ( .A(n2196), .B(n2197), .Z(n2012) );
  ANDN U3082 ( .B(n2198), .A(n2199), .Z(n2196) );
  AND U3083 ( .A(a[42]), .B(b[9]), .Z(n2195) );
  XNOR U3084 ( .A(n2200), .B(n2017), .Z(n2019) );
  XOR U3085 ( .A(n2201), .B(n2202), .Z(n2017) );
  ANDN U3086 ( .B(n2203), .A(n2204), .Z(n2201) );
  AND U3087 ( .A(b[8]), .B(a[43]), .Z(n2200) );
  XNOR U3088 ( .A(n2205), .B(n2022), .Z(n2024) );
  XOR U3089 ( .A(n2206), .B(n2207), .Z(n2022) );
  ANDN U3090 ( .B(n2208), .A(n2209), .Z(n2206) );
  AND U3091 ( .A(a[44]), .B(b[7]), .Z(n2205) );
  XNOR U3092 ( .A(n2210), .B(n2027), .Z(n2029) );
  XOR U3093 ( .A(n2211), .B(n2212), .Z(n2027) );
  ANDN U3094 ( .B(n2213), .A(n2214), .Z(n2211) );
  AND U3095 ( .A(b[6]), .B(a[45]), .Z(n2210) );
  XNOR U3096 ( .A(n2215), .B(n2032), .Z(n2034) );
  XOR U3097 ( .A(n2216), .B(n2217), .Z(n2032) );
  ANDN U3098 ( .B(n2218), .A(n2219), .Z(n2216) );
  AND U3099 ( .A(b[5]), .B(a[46]), .Z(n2215) );
  XNOR U3100 ( .A(n2220), .B(n2037), .Z(n2039) );
  XOR U3101 ( .A(n2221), .B(n2222), .Z(n2037) );
  ANDN U3102 ( .B(n2223), .A(n2224), .Z(n2221) );
  AND U3103 ( .A(b[4]), .B(a[47]), .Z(n2220) );
  XNOR U3104 ( .A(n2225), .B(n2226), .Z(n2051) );
  NANDN U3105 ( .A(n2227), .B(n2228), .Z(n2226) );
  XNOR U3106 ( .A(n2229), .B(n2042), .Z(n2044) );
  XNOR U3107 ( .A(n2230), .B(n2231), .Z(n2042) );
  AND U3108 ( .A(n2232), .B(n2233), .Z(n2230) );
  AND U3109 ( .A(b[3]), .B(a[48]), .Z(n2229) );
  XNOR U3110 ( .A(n2234), .B(n2235), .Z(swire[50]) );
  XOR U3111 ( .A(n2061), .B(n2237), .Z(n2235) );
  XNOR U3112 ( .A(n2060), .B(n2236), .Z(n2237) );
  IV U3113 ( .A(n2234), .Z(n2236) );
  NAND U3114 ( .A(a[50]), .B(b[0]), .Z(n2060) );
  XNOR U3115 ( .A(n2227), .B(n2228), .Z(n2061) );
  XOR U3116 ( .A(n2225), .B(n2238), .Z(n2228) );
  NAND U3117 ( .A(b[1]), .B(a[49]), .Z(n2238) );
  XOR U3118 ( .A(n2233), .B(n2239), .Z(n2227) );
  XOR U3119 ( .A(n2225), .B(n2232), .Z(n2239) );
  XNOR U3120 ( .A(n2240), .B(n2231), .Z(n2232) );
  AND U3121 ( .A(b[2]), .B(a[48]), .Z(n2240) );
  NANDN U3122 ( .A(n2241), .B(n2242), .Z(n2225) );
  XOR U3123 ( .A(n2231), .B(n2223), .Z(n2243) );
  XNOR U3124 ( .A(n2222), .B(n2218), .Z(n2244) );
  XNOR U3125 ( .A(n2217), .B(n2213), .Z(n2245) );
  XNOR U3126 ( .A(n2212), .B(n2208), .Z(n2246) );
  XNOR U3127 ( .A(n2207), .B(n2203), .Z(n2247) );
  XNOR U3128 ( .A(n2202), .B(n2198), .Z(n2248) );
  XNOR U3129 ( .A(n2197), .B(n2193), .Z(n2249) );
  XNOR U3130 ( .A(n2192), .B(n2188), .Z(n2250) );
  XNOR U3131 ( .A(n2187), .B(n2183), .Z(n2251) );
  XNOR U3132 ( .A(n2182), .B(n2178), .Z(n2252) );
  XNOR U3133 ( .A(n2177), .B(n2173), .Z(n2253) );
  XNOR U3134 ( .A(n2172), .B(n2168), .Z(n2254) );
  XNOR U3135 ( .A(n2167), .B(n2163), .Z(n2255) );
  XNOR U3136 ( .A(n2162), .B(n2158), .Z(n2256) );
  XNOR U3137 ( .A(n2157), .B(n2153), .Z(n2257) );
  XNOR U3138 ( .A(n2152), .B(n2148), .Z(n2258) );
  XNOR U3139 ( .A(n2147), .B(n2143), .Z(n2259) );
  XNOR U3140 ( .A(n2142), .B(n2138), .Z(n2260) );
  XNOR U3141 ( .A(n2137), .B(n2133), .Z(n2261) );
  XNOR U3142 ( .A(n2132), .B(n2128), .Z(n2262) );
  XNOR U3143 ( .A(n2127), .B(n2123), .Z(n2263) );
  XNOR U3144 ( .A(n2122), .B(n2118), .Z(n2264) );
  XNOR U3145 ( .A(n2117), .B(n2113), .Z(n2265) );
  XNOR U3146 ( .A(n2112), .B(n2108), .Z(n2266) );
  XNOR U3147 ( .A(n2107), .B(n2103), .Z(n2267) );
  XOR U3148 ( .A(n2102), .B(n2099), .Z(n2268) );
  XOR U3149 ( .A(n2269), .B(n2270), .Z(n2099) );
  XOR U3150 ( .A(n2097), .B(n2271), .Z(n2270) );
  XOR U3151 ( .A(n2272), .B(n2273), .Z(n2271) );
  XOR U3152 ( .A(n2274), .B(n2275), .Z(n2273) );
  NAND U3153 ( .A(a[20]), .B(b[30]), .Z(n2275) );
  AND U3154 ( .A(a[19]), .B(b[31]), .Z(n2274) );
  XOR U3155 ( .A(n2276), .B(n2272), .Z(n2269) );
  XOR U3156 ( .A(n2277), .B(n2278), .Z(n2272) );
  NOR U3157 ( .A(n2279), .B(n2280), .Z(n2277) );
  AND U3158 ( .A(a[21]), .B(b[29]), .Z(n2276) );
  XNOR U3159 ( .A(n2281), .B(n2097), .Z(n2098) );
  XOR U3160 ( .A(n2282), .B(n2283), .Z(n2097) );
  ANDN U3161 ( .B(n2284), .A(n2285), .Z(n2282) );
  AND U3162 ( .A(a[22]), .B(b[28]), .Z(n2281) );
  XNOR U3163 ( .A(n2286), .B(n2102), .Z(n2104) );
  XOR U3164 ( .A(n2287), .B(n2288), .Z(n2102) );
  ANDN U3165 ( .B(n2289), .A(n2290), .Z(n2287) );
  AND U3166 ( .A(a[23]), .B(b[27]), .Z(n2286) );
  XNOR U3167 ( .A(n2291), .B(n2107), .Z(n2109) );
  XOR U3168 ( .A(n2292), .B(n2293), .Z(n2107) );
  ANDN U3169 ( .B(n2294), .A(n2295), .Z(n2292) );
  AND U3170 ( .A(a[24]), .B(b[26]), .Z(n2291) );
  XNOR U3171 ( .A(n2296), .B(n2112), .Z(n2114) );
  XOR U3172 ( .A(n2297), .B(n2298), .Z(n2112) );
  ANDN U3173 ( .B(n2299), .A(n2300), .Z(n2297) );
  AND U3174 ( .A(b[25]), .B(a[25]), .Z(n2296) );
  XNOR U3175 ( .A(n2301), .B(n2117), .Z(n2119) );
  XOR U3176 ( .A(n2302), .B(n2303), .Z(n2117) );
  ANDN U3177 ( .B(n2304), .A(n2305), .Z(n2302) );
  AND U3178 ( .A(a[26]), .B(b[24]), .Z(n2301) );
  XNOR U3179 ( .A(n2306), .B(n2122), .Z(n2124) );
  XOR U3180 ( .A(n2307), .B(n2308), .Z(n2122) );
  ANDN U3181 ( .B(n2309), .A(n2310), .Z(n2307) );
  AND U3182 ( .A(b[23]), .B(a[27]), .Z(n2306) );
  XNOR U3183 ( .A(n2311), .B(n2127), .Z(n2129) );
  XOR U3184 ( .A(n2312), .B(n2313), .Z(n2127) );
  ANDN U3185 ( .B(n2314), .A(n2315), .Z(n2312) );
  AND U3186 ( .A(a[28]), .B(b[22]), .Z(n2311) );
  XNOR U3187 ( .A(n2316), .B(n2132), .Z(n2134) );
  XOR U3188 ( .A(n2317), .B(n2318), .Z(n2132) );
  ANDN U3189 ( .B(n2319), .A(n2320), .Z(n2317) );
  AND U3190 ( .A(b[21]), .B(a[29]), .Z(n2316) );
  XNOR U3191 ( .A(n2321), .B(n2137), .Z(n2139) );
  XOR U3192 ( .A(n2322), .B(n2323), .Z(n2137) );
  ANDN U3193 ( .B(n2324), .A(n2325), .Z(n2322) );
  AND U3194 ( .A(a[30]), .B(b[20]), .Z(n2321) );
  XNOR U3195 ( .A(n2326), .B(n2142), .Z(n2144) );
  XOR U3196 ( .A(n2327), .B(n2328), .Z(n2142) );
  ANDN U3197 ( .B(n2329), .A(n2330), .Z(n2327) );
  AND U3198 ( .A(b[19]), .B(a[31]), .Z(n2326) );
  XNOR U3199 ( .A(n2331), .B(n2147), .Z(n2149) );
  XOR U3200 ( .A(n2332), .B(n2333), .Z(n2147) );
  ANDN U3201 ( .B(n2334), .A(n2335), .Z(n2332) );
  AND U3202 ( .A(a[32]), .B(b[18]), .Z(n2331) );
  XNOR U3203 ( .A(n2336), .B(n2152), .Z(n2154) );
  XOR U3204 ( .A(n2337), .B(n2338), .Z(n2152) );
  ANDN U3205 ( .B(n2339), .A(n2340), .Z(n2337) );
  AND U3206 ( .A(b[17]), .B(a[33]), .Z(n2336) );
  XNOR U3207 ( .A(n2341), .B(n2157), .Z(n2159) );
  XOR U3208 ( .A(n2342), .B(n2343), .Z(n2157) );
  ANDN U3209 ( .B(n2344), .A(n2345), .Z(n2342) );
  AND U3210 ( .A(a[34]), .B(b[16]), .Z(n2341) );
  XNOR U3211 ( .A(n2346), .B(n2162), .Z(n2164) );
  XOR U3212 ( .A(n2347), .B(n2348), .Z(n2162) );
  ANDN U3213 ( .B(n2349), .A(n2350), .Z(n2347) );
  AND U3214 ( .A(b[15]), .B(a[35]), .Z(n2346) );
  XNOR U3215 ( .A(n2351), .B(n2167), .Z(n2169) );
  XOR U3216 ( .A(n2352), .B(n2353), .Z(n2167) );
  ANDN U3217 ( .B(n2354), .A(n2355), .Z(n2352) );
  AND U3218 ( .A(a[36]), .B(b[14]), .Z(n2351) );
  XNOR U3219 ( .A(n2356), .B(n2172), .Z(n2174) );
  XOR U3220 ( .A(n2357), .B(n2358), .Z(n2172) );
  ANDN U3221 ( .B(n2359), .A(n2360), .Z(n2357) );
  AND U3222 ( .A(b[13]), .B(a[37]), .Z(n2356) );
  XNOR U3223 ( .A(n2361), .B(n2177), .Z(n2179) );
  XOR U3224 ( .A(n2362), .B(n2363), .Z(n2177) );
  ANDN U3225 ( .B(n2364), .A(n2365), .Z(n2362) );
  AND U3226 ( .A(a[38]), .B(b[12]), .Z(n2361) );
  XNOR U3227 ( .A(n2366), .B(n2182), .Z(n2184) );
  XOR U3228 ( .A(n2367), .B(n2368), .Z(n2182) );
  ANDN U3229 ( .B(n2369), .A(n2370), .Z(n2367) );
  AND U3230 ( .A(b[11]), .B(a[39]), .Z(n2366) );
  XNOR U3231 ( .A(n2371), .B(n2187), .Z(n2189) );
  XOR U3232 ( .A(n2372), .B(n2373), .Z(n2187) );
  ANDN U3233 ( .B(n2374), .A(n2375), .Z(n2372) );
  AND U3234 ( .A(a[40]), .B(b[10]), .Z(n2371) );
  XNOR U3235 ( .A(n2376), .B(n2192), .Z(n2194) );
  XOR U3236 ( .A(n2377), .B(n2378), .Z(n2192) );
  ANDN U3237 ( .B(n2379), .A(n2380), .Z(n2377) );
  AND U3238 ( .A(b[9]), .B(a[41]), .Z(n2376) );
  XNOR U3239 ( .A(n2381), .B(n2197), .Z(n2199) );
  XOR U3240 ( .A(n2382), .B(n2383), .Z(n2197) );
  ANDN U3241 ( .B(n2384), .A(n2385), .Z(n2382) );
  AND U3242 ( .A(a[42]), .B(b[8]), .Z(n2381) );
  XNOR U3243 ( .A(n2386), .B(n2202), .Z(n2204) );
  XOR U3244 ( .A(n2387), .B(n2388), .Z(n2202) );
  ANDN U3245 ( .B(n2389), .A(n2390), .Z(n2387) );
  AND U3246 ( .A(b[7]), .B(a[43]), .Z(n2386) );
  XNOR U3247 ( .A(n2391), .B(n2207), .Z(n2209) );
  XOR U3248 ( .A(n2392), .B(n2393), .Z(n2207) );
  ANDN U3249 ( .B(n2394), .A(n2395), .Z(n2392) );
  AND U3250 ( .A(b[6]), .B(a[44]), .Z(n2391) );
  XNOR U3251 ( .A(n2396), .B(n2212), .Z(n2214) );
  XOR U3252 ( .A(n2397), .B(n2398), .Z(n2212) );
  ANDN U3253 ( .B(n2399), .A(n2400), .Z(n2397) );
  AND U3254 ( .A(b[5]), .B(a[45]), .Z(n2396) );
  XNOR U3255 ( .A(n2401), .B(n2217), .Z(n2219) );
  XOR U3256 ( .A(n2402), .B(n2403), .Z(n2217) );
  ANDN U3257 ( .B(n2404), .A(n2405), .Z(n2402) );
  AND U3258 ( .A(b[4]), .B(a[46]), .Z(n2401) );
  XNOR U3259 ( .A(n2406), .B(n2407), .Z(n2231) );
  NANDN U3260 ( .A(n2408), .B(n2409), .Z(n2407) );
  XNOR U3261 ( .A(n2410), .B(n2222), .Z(n2224) );
  XNOR U3262 ( .A(n2411), .B(n2412), .Z(n2222) );
  AND U3263 ( .A(n2413), .B(n2414), .Z(n2411) );
  AND U3264 ( .A(b[3]), .B(a[47]), .Z(n2410) );
  XNOR U3265 ( .A(n2415), .B(n2416), .Z(swire[49]) );
  XOR U3266 ( .A(n2242), .B(n2417), .Z(n2416) );
  XOR U3267 ( .A(n2241), .B(n2415), .Z(n2417) );
  NAND U3268 ( .A(a[49]), .B(b[0]), .Z(n2241) );
  XNOR U3269 ( .A(n2408), .B(n2409), .Z(n2242) );
  XOR U3270 ( .A(n2406), .B(n2418), .Z(n2409) );
  NAND U3271 ( .A(a[48]), .B(b[1]), .Z(n2418) );
  XOR U3272 ( .A(n2414), .B(n2419), .Z(n2408) );
  XOR U3273 ( .A(n2406), .B(n2413), .Z(n2419) );
  XNOR U3274 ( .A(n2420), .B(n2412), .Z(n2413) );
  AND U3275 ( .A(b[2]), .B(a[47]), .Z(n2420) );
  NANDN U3276 ( .A(n2421), .B(n2422), .Z(n2406) );
  XOR U3277 ( .A(n2412), .B(n2404), .Z(n2423) );
  XNOR U3278 ( .A(n2403), .B(n2399), .Z(n2424) );
  XNOR U3279 ( .A(n2398), .B(n2394), .Z(n2425) );
  XNOR U3280 ( .A(n2393), .B(n2389), .Z(n2426) );
  XNOR U3281 ( .A(n2388), .B(n2384), .Z(n2427) );
  XNOR U3282 ( .A(n2383), .B(n2379), .Z(n2428) );
  XNOR U3283 ( .A(n2378), .B(n2374), .Z(n2429) );
  XNOR U3284 ( .A(n2373), .B(n2369), .Z(n2430) );
  XNOR U3285 ( .A(n2368), .B(n2364), .Z(n2431) );
  XNOR U3286 ( .A(n2363), .B(n2359), .Z(n2432) );
  XNOR U3287 ( .A(n2358), .B(n2354), .Z(n2433) );
  XNOR U3288 ( .A(n2353), .B(n2349), .Z(n2434) );
  XNOR U3289 ( .A(n2348), .B(n2344), .Z(n2435) );
  XNOR U3290 ( .A(n2343), .B(n2339), .Z(n2436) );
  XNOR U3291 ( .A(n2338), .B(n2334), .Z(n2437) );
  XNOR U3292 ( .A(n2333), .B(n2329), .Z(n2438) );
  XNOR U3293 ( .A(n2328), .B(n2324), .Z(n2439) );
  XNOR U3294 ( .A(n2323), .B(n2319), .Z(n2440) );
  XNOR U3295 ( .A(n2318), .B(n2314), .Z(n2441) );
  XNOR U3296 ( .A(n2313), .B(n2309), .Z(n2442) );
  XNOR U3297 ( .A(n2308), .B(n2304), .Z(n2443) );
  XNOR U3298 ( .A(n2303), .B(n2299), .Z(n2444) );
  XNOR U3299 ( .A(n2298), .B(n2294), .Z(n2445) );
  XNOR U3300 ( .A(n2293), .B(n2289), .Z(n2446) );
  XNOR U3301 ( .A(n2288), .B(n2284), .Z(n2447) );
  XOR U3302 ( .A(n2283), .B(n2280), .Z(n2448) );
  XOR U3303 ( .A(n2449), .B(n2450), .Z(n2280) );
  XOR U3304 ( .A(n2278), .B(n2451), .Z(n2450) );
  XOR U3305 ( .A(n2452), .B(n2453), .Z(n2451) );
  XOR U3306 ( .A(n2454), .B(n2455), .Z(n2453) );
  NAND U3307 ( .A(a[19]), .B(b[30]), .Z(n2455) );
  AND U3308 ( .A(a[18]), .B(b[31]), .Z(n2454) );
  XOR U3309 ( .A(n2456), .B(n2452), .Z(n2449) );
  XOR U3310 ( .A(n2457), .B(n2458), .Z(n2452) );
  NOR U3311 ( .A(n2459), .B(n2460), .Z(n2457) );
  AND U3312 ( .A(a[20]), .B(b[29]), .Z(n2456) );
  XNOR U3313 ( .A(n2461), .B(n2278), .Z(n2279) );
  XOR U3314 ( .A(n2462), .B(n2463), .Z(n2278) );
  ANDN U3315 ( .B(n2464), .A(n2465), .Z(n2462) );
  AND U3316 ( .A(a[21]), .B(b[28]), .Z(n2461) );
  XNOR U3317 ( .A(n2466), .B(n2283), .Z(n2285) );
  XOR U3318 ( .A(n2467), .B(n2468), .Z(n2283) );
  ANDN U3319 ( .B(n2469), .A(n2470), .Z(n2467) );
  AND U3320 ( .A(a[22]), .B(b[27]), .Z(n2466) );
  XNOR U3321 ( .A(n2471), .B(n2288), .Z(n2290) );
  XOR U3322 ( .A(n2472), .B(n2473), .Z(n2288) );
  ANDN U3323 ( .B(n2474), .A(n2475), .Z(n2472) );
  AND U3324 ( .A(a[23]), .B(b[26]), .Z(n2471) );
  XNOR U3325 ( .A(n2476), .B(n2293), .Z(n2295) );
  XOR U3326 ( .A(n2477), .B(n2478), .Z(n2293) );
  ANDN U3327 ( .B(n2479), .A(n2480), .Z(n2477) );
  AND U3328 ( .A(a[24]), .B(b[25]), .Z(n2476) );
  XNOR U3329 ( .A(n2481), .B(n2298), .Z(n2300) );
  XOR U3330 ( .A(n2482), .B(n2483), .Z(n2298) );
  ANDN U3331 ( .B(n2484), .A(n2485), .Z(n2482) );
  AND U3332 ( .A(b[24]), .B(a[25]), .Z(n2481) );
  XNOR U3333 ( .A(n2486), .B(n2303), .Z(n2305) );
  XOR U3334 ( .A(n2487), .B(n2488), .Z(n2303) );
  ANDN U3335 ( .B(n2489), .A(n2490), .Z(n2487) );
  AND U3336 ( .A(a[26]), .B(b[23]), .Z(n2486) );
  XNOR U3337 ( .A(n2491), .B(n2308), .Z(n2310) );
  XOR U3338 ( .A(n2492), .B(n2493), .Z(n2308) );
  ANDN U3339 ( .B(n2494), .A(n2495), .Z(n2492) );
  AND U3340 ( .A(b[22]), .B(a[27]), .Z(n2491) );
  XNOR U3341 ( .A(n2496), .B(n2313), .Z(n2315) );
  XOR U3342 ( .A(n2497), .B(n2498), .Z(n2313) );
  ANDN U3343 ( .B(n2499), .A(n2500), .Z(n2497) );
  AND U3344 ( .A(a[28]), .B(b[21]), .Z(n2496) );
  XNOR U3345 ( .A(n2501), .B(n2318), .Z(n2320) );
  XOR U3346 ( .A(n2502), .B(n2503), .Z(n2318) );
  ANDN U3347 ( .B(n2504), .A(n2505), .Z(n2502) );
  AND U3348 ( .A(b[20]), .B(a[29]), .Z(n2501) );
  XNOR U3349 ( .A(n2506), .B(n2323), .Z(n2325) );
  XOR U3350 ( .A(n2507), .B(n2508), .Z(n2323) );
  ANDN U3351 ( .B(n2509), .A(n2510), .Z(n2507) );
  AND U3352 ( .A(a[30]), .B(b[19]), .Z(n2506) );
  XNOR U3353 ( .A(n2511), .B(n2328), .Z(n2330) );
  XOR U3354 ( .A(n2512), .B(n2513), .Z(n2328) );
  ANDN U3355 ( .B(n2514), .A(n2515), .Z(n2512) );
  AND U3356 ( .A(b[18]), .B(a[31]), .Z(n2511) );
  XNOR U3357 ( .A(n2516), .B(n2333), .Z(n2335) );
  XOR U3358 ( .A(n2517), .B(n2518), .Z(n2333) );
  ANDN U3359 ( .B(n2519), .A(n2520), .Z(n2517) );
  AND U3360 ( .A(a[32]), .B(b[17]), .Z(n2516) );
  XNOR U3361 ( .A(n2521), .B(n2338), .Z(n2340) );
  XOR U3362 ( .A(n2522), .B(n2523), .Z(n2338) );
  ANDN U3363 ( .B(n2524), .A(n2525), .Z(n2522) );
  AND U3364 ( .A(b[16]), .B(a[33]), .Z(n2521) );
  XNOR U3365 ( .A(n2526), .B(n2343), .Z(n2345) );
  XOR U3366 ( .A(n2527), .B(n2528), .Z(n2343) );
  ANDN U3367 ( .B(n2529), .A(n2530), .Z(n2527) );
  AND U3368 ( .A(a[34]), .B(b[15]), .Z(n2526) );
  XNOR U3369 ( .A(n2531), .B(n2348), .Z(n2350) );
  XOR U3370 ( .A(n2532), .B(n2533), .Z(n2348) );
  ANDN U3371 ( .B(n2534), .A(n2535), .Z(n2532) );
  AND U3372 ( .A(b[14]), .B(a[35]), .Z(n2531) );
  XNOR U3373 ( .A(n2536), .B(n2353), .Z(n2355) );
  XOR U3374 ( .A(n2537), .B(n2538), .Z(n2353) );
  ANDN U3375 ( .B(n2539), .A(n2540), .Z(n2537) );
  AND U3376 ( .A(a[36]), .B(b[13]), .Z(n2536) );
  XNOR U3377 ( .A(n2541), .B(n2358), .Z(n2360) );
  XOR U3378 ( .A(n2542), .B(n2543), .Z(n2358) );
  ANDN U3379 ( .B(n2544), .A(n2545), .Z(n2542) );
  AND U3380 ( .A(b[12]), .B(a[37]), .Z(n2541) );
  XNOR U3381 ( .A(n2546), .B(n2363), .Z(n2365) );
  XOR U3382 ( .A(n2547), .B(n2548), .Z(n2363) );
  ANDN U3383 ( .B(n2549), .A(n2550), .Z(n2547) );
  AND U3384 ( .A(a[38]), .B(b[11]), .Z(n2546) );
  XNOR U3385 ( .A(n2551), .B(n2368), .Z(n2370) );
  XOR U3386 ( .A(n2552), .B(n2553), .Z(n2368) );
  ANDN U3387 ( .B(n2554), .A(n2555), .Z(n2552) );
  AND U3388 ( .A(b[10]), .B(a[39]), .Z(n2551) );
  XNOR U3389 ( .A(n2556), .B(n2373), .Z(n2375) );
  XOR U3390 ( .A(n2557), .B(n2558), .Z(n2373) );
  ANDN U3391 ( .B(n2559), .A(n2560), .Z(n2557) );
  AND U3392 ( .A(a[40]), .B(b[9]), .Z(n2556) );
  XNOR U3393 ( .A(n2561), .B(n2378), .Z(n2380) );
  XOR U3394 ( .A(n2562), .B(n2563), .Z(n2378) );
  ANDN U3395 ( .B(n2564), .A(n2565), .Z(n2562) );
  AND U3396 ( .A(b[8]), .B(a[41]), .Z(n2561) );
  XNOR U3397 ( .A(n2566), .B(n2383), .Z(n2385) );
  XOR U3398 ( .A(n2567), .B(n2568), .Z(n2383) );
  ANDN U3399 ( .B(n2569), .A(n2570), .Z(n2567) );
  AND U3400 ( .A(a[42]), .B(b[7]), .Z(n2566) );
  XNOR U3401 ( .A(n2571), .B(n2388), .Z(n2390) );
  XOR U3402 ( .A(n2572), .B(n2573), .Z(n2388) );
  ANDN U3403 ( .B(n2574), .A(n2575), .Z(n2572) );
  AND U3404 ( .A(b[6]), .B(a[43]), .Z(n2571) );
  XNOR U3405 ( .A(n2576), .B(n2393), .Z(n2395) );
  XOR U3406 ( .A(n2577), .B(n2578), .Z(n2393) );
  ANDN U3407 ( .B(n2579), .A(n2580), .Z(n2577) );
  AND U3408 ( .A(b[5]), .B(a[44]), .Z(n2576) );
  XNOR U3409 ( .A(n2581), .B(n2398), .Z(n2400) );
  XOR U3410 ( .A(n2582), .B(n2583), .Z(n2398) );
  ANDN U3411 ( .B(n2584), .A(n2585), .Z(n2582) );
  AND U3412 ( .A(b[4]), .B(a[45]), .Z(n2581) );
  XNOR U3413 ( .A(n2586), .B(n2587), .Z(n2412) );
  NANDN U3414 ( .A(n2588), .B(n2589), .Z(n2587) );
  XNOR U3415 ( .A(n2590), .B(n2403), .Z(n2405) );
  XNOR U3416 ( .A(n2591), .B(n2592), .Z(n2403) );
  AND U3417 ( .A(n2593), .B(n2594), .Z(n2591) );
  AND U3418 ( .A(b[3]), .B(a[46]), .Z(n2590) );
  XNOR U3419 ( .A(n2595), .B(n2596), .Z(swire[48]) );
  XOR U3420 ( .A(n2422), .B(n2598), .Z(n2596) );
  XNOR U3421 ( .A(n2421), .B(n2597), .Z(n2598) );
  IV U3422 ( .A(n2595), .Z(n2597) );
  NAND U3423 ( .A(a[48]), .B(b[0]), .Z(n2421) );
  XNOR U3424 ( .A(n2588), .B(n2589), .Z(n2422) );
  XOR U3425 ( .A(n2586), .B(n2599), .Z(n2589) );
  NAND U3426 ( .A(b[1]), .B(a[47]), .Z(n2599) );
  XOR U3427 ( .A(n2594), .B(n2600), .Z(n2588) );
  XOR U3428 ( .A(n2586), .B(n2593), .Z(n2600) );
  XNOR U3429 ( .A(n2601), .B(n2592), .Z(n2593) );
  AND U3430 ( .A(b[2]), .B(a[46]), .Z(n2601) );
  NANDN U3431 ( .A(n2602), .B(n2603), .Z(n2586) );
  XOR U3432 ( .A(n2592), .B(n2584), .Z(n2604) );
  XNOR U3433 ( .A(n2583), .B(n2579), .Z(n2605) );
  XNOR U3434 ( .A(n2578), .B(n2574), .Z(n2606) );
  XNOR U3435 ( .A(n2573), .B(n2569), .Z(n2607) );
  XNOR U3436 ( .A(n2568), .B(n2564), .Z(n2608) );
  XNOR U3437 ( .A(n2563), .B(n2559), .Z(n2609) );
  XNOR U3438 ( .A(n2558), .B(n2554), .Z(n2610) );
  XNOR U3439 ( .A(n2553), .B(n2549), .Z(n2611) );
  XNOR U3440 ( .A(n2548), .B(n2544), .Z(n2612) );
  XNOR U3441 ( .A(n2543), .B(n2539), .Z(n2613) );
  XNOR U3442 ( .A(n2538), .B(n2534), .Z(n2614) );
  XNOR U3443 ( .A(n2533), .B(n2529), .Z(n2615) );
  XNOR U3444 ( .A(n2528), .B(n2524), .Z(n2616) );
  XNOR U3445 ( .A(n2523), .B(n2519), .Z(n2617) );
  XNOR U3446 ( .A(n2518), .B(n2514), .Z(n2618) );
  XNOR U3447 ( .A(n2513), .B(n2509), .Z(n2619) );
  XNOR U3448 ( .A(n2508), .B(n2504), .Z(n2620) );
  XNOR U3449 ( .A(n2503), .B(n2499), .Z(n2621) );
  XNOR U3450 ( .A(n2498), .B(n2494), .Z(n2622) );
  XNOR U3451 ( .A(n2493), .B(n2489), .Z(n2623) );
  XNOR U3452 ( .A(n2488), .B(n2484), .Z(n2624) );
  XNOR U3453 ( .A(n2483), .B(n2479), .Z(n2625) );
  XNOR U3454 ( .A(n2478), .B(n2474), .Z(n2626) );
  XNOR U3455 ( .A(n2473), .B(n2469), .Z(n2627) );
  XNOR U3456 ( .A(n2468), .B(n2464), .Z(n2628) );
  XOR U3457 ( .A(n2463), .B(n2460), .Z(n2629) );
  XOR U3458 ( .A(n2630), .B(n2631), .Z(n2460) );
  XOR U3459 ( .A(n2458), .B(n2632), .Z(n2631) );
  XOR U3460 ( .A(n2633), .B(n2634), .Z(n2632) );
  XOR U3461 ( .A(n2635), .B(n2636), .Z(n2634) );
  NAND U3462 ( .A(a[18]), .B(b[30]), .Z(n2636) );
  AND U3463 ( .A(a[17]), .B(b[31]), .Z(n2635) );
  XOR U3464 ( .A(n2637), .B(n2633), .Z(n2630) );
  XOR U3465 ( .A(n2638), .B(n2639), .Z(n2633) );
  NOR U3466 ( .A(n2640), .B(n2641), .Z(n2638) );
  AND U3467 ( .A(a[19]), .B(b[29]), .Z(n2637) );
  XNOR U3468 ( .A(n2642), .B(n2458), .Z(n2459) );
  XOR U3469 ( .A(n2643), .B(n2644), .Z(n2458) );
  ANDN U3470 ( .B(n2645), .A(n2646), .Z(n2643) );
  AND U3471 ( .A(a[20]), .B(b[28]), .Z(n2642) );
  XNOR U3472 ( .A(n2647), .B(n2463), .Z(n2465) );
  XOR U3473 ( .A(n2648), .B(n2649), .Z(n2463) );
  ANDN U3474 ( .B(n2650), .A(n2651), .Z(n2648) );
  AND U3475 ( .A(a[21]), .B(b[27]), .Z(n2647) );
  XNOR U3476 ( .A(n2652), .B(n2468), .Z(n2470) );
  XOR U3477 ( .A(n2653), .B(n2654), .Z(n2468) );
  ANDN U3478 ( .B(n2655), .A(n2656), .Z(n2653) );
  AND U3479 ( .A(a[22]), .B(b[26]), .Z(n2652) );
  XNOR U3480 ( .A(n2657), .B(n2473), .Z(n2475) );
  XOR U3481 ( .A(n2658), .B(n2659), .Z(n2473) );
  ANDN U3482 ( .B(n2660), .A(n2661), .Z(n2658) );
  AND U3483 ( .A(a[23]), .B(b[25]), .Z(n2657) );
  XNOR U3484 ( .A(n2662), .B(n2478), .Z(n2480) );
  XOR U3485 ( .A(n2663), .B(n2664), .Z(n2478) );
  ANDN U3486 ( .B(n2665), .A(n2666), .Z(n2663) );
  AND U3487 ( .A(a[24]), .B(b[24]), .Z(n2662) );
  XNOR U3488 ( .A(n2667), .B(n2483), .Z(n2485) );
  XOR U3489 ( .A(n2668), .B(n2669), .Z(n2483) );
  ANDN U3490 ( .B(n2670), .A(n2671), .Z(n2668) );
  AND U3491 ( .A(b[23]), .B(a[25]), .Z(n2667) );
  XNOR U3492 ( .A(n2672), .B(n2488), .Z(n2490) );
  XOR U3493 ( .A(n2673), .B(n2674), .Z(n2488) );
  ANDN U3494 ( .B(n2675), .A(n2676), .Z(n2673) );
  AND U3495 ( .A(a[26]), .B(b[22]), .Z(n2672) );
  XNOR U3496 ( .A(n2677), .B(n2493), .Z(n2495) );
  XOR U3497 ( .A(n2678), .B(n2679), .Z(n2493) );
  ANDN U3498 ( .B(n2680), .A(n2681), .Z(n2678) );
  AND U3499 ( .A(b[21]), .B(a[27]), .Z(n2677) );
  XNOR U3500 ( .A(n2682), .B(n2498), .Z(n2500) );
  XOR U3501 ( .A(n2683), .B(n2684), .Z(n2498) );
  ANDN U3502 ( .B(n2685), .A(n2686), .Z(n2683) );
  AND U3503 ( .A(a[28]), .B(b[20]), .Z(n2682) );
  XNOR U3504 ( .A(n2687), .B(n2503), .Z(n2505) );
  XOR U3505 ( .A(n2688), .B(n2689), .Z(n2503) );
  ANDN U3506 ( .B(n2690), .A(n2691), .Z(n2688) );
  AND U3507 ( .A(b[19]), .B(a[29]), .Z(n2687) );
  XNOR U3508 ( .A(n2692), .B(n2508), .Z(n2510) );
  XOR U3509 ( .A(n2693), .B(n2694), .Z(n2508) );
  ANDN U3510 ( .B(n2695), .A(n2696), .Z(n2693) );
  AND U3511 ( .A(a[30]), .B(b[18]), .Z(n2692) );
  XNOR U3512 ( .A(n2697), .B(n2513), .Z(n2515) );
  XOR U3513 ( .A(n2698), .B(n2699), .Z(n2513) );
  ANDN U3514 ( .B(n2700), .A(n2701), .Z(n2698) );
  AND U3515 ( .A(b[17]), .B(a[31]), .Z(n2697) );
  XNOR U3516 ( .A(n2702), .B(n2518), .Z(n2520) );
  XOR U3517 ( .A(n2703), .B(n2704), .Z(n2518) );
  ANDN U3518 ( .B(n2705), .A(n2706), .Z(n2703) );
  AND U3519 ( .A(a[32]), .B(b[16]), .Z(n2702) );
  XNOR U3520 ( .A(n2707), .B(n2523), .Z(n2525) );
  XOR U3521 ( .A(n2708), .B(n2709), .Z(n2523) );
  ANDN U3522 ( .B(n2710), .A(n2711), .Z(n2708) );
  AND U3523 ( .A(b[15]), .B(a[33]), .Z(n2707) );
  XNOR U3524 ( .A(n2712), .B(n2528), .Z(n2530) );
  XOR U3525 ( .A(n2713), .B(n2714), .Z(n2528) );
  ANDN U3526 ( .B(n2715), .A(n2716), .Z(n2713) );
  AND U3527 ( .A(a[34]), .B(b[14]), .Z(n2712) );
  XNOR U3528 ( .A(n2717), .B(n2533), .Z(n2535) );
  XOR U3529 ( .A(n2718), .B(n2719), .Z(n2533) );
  ANDN U3530 ( .B(n2720), .A(n2721), .Z(n2718) );
  AND U3531 ( .A(b[13]), .B(a[35]), .Z(n2717) );
  XNOR U3532 ( .A(n2722), .B(n2538), .Z(n2540) );
  XOR U3533 ( .A(n2723), .B(n2724), .Z(n2538) );
  ANDN U3534 ( .B(n2725), .A(n2726), .Z(n2723) );
  AND U3535 ( .A(a[36]), .B(b[12]), .Z(n2722) );
  XNOR U3536 ( .A(n2727), .B(n2543), .Z(n2545) );
  XOR U3537 ( .A(n2728), .B(n2729), .Z(n2543) );
  ANDN U3538 ( .B(n2730), .A(n2731), .Z(n2728) );
  AND U3539 ( .A(b[11]), .B(a[37]), .Z(n2727) );
  XNOR U3540 ( .A(n2732), .B(n2548), .Z(n2550) );
  XOR U3541 ( .A(n2733), .B(n2734), .Z(n2548) );
  ANDN U3542 ( .B(n2735), .A(n2736), .Z(n2733) );
  AND U3543 ( .A(a[38]), .B(b[10]), .Z(n2732) );
  XNOR U3544 ( .A(n2737), .B(n2553), .Z(n2555) );
  XOR U3545 ( .A(n2738), .B(n2739), .Z(n2553) );
  ANDN U3546 ( .B(n2740), .A(n2741), .Z(n2738) );
  AND U3547 ( .A(b[9]), .B(a[39]), .Z(n2737) );
  XNOR U3548 ( .A(n2742), .B(n2558), .Z(n2560) );
  XOR U3549 ( .A(n2743), .B(n2744), .Z(n2558) );
  ANDN U3550 ( .B(n2745), .A(n2746), .Z(n2743) );
  AND U3551 ( .A(a[40]), .B(b[8]), .Z(n2742) );
  XNOR U3552 ( .A(n2747), .B(n2563), .Z(n2565) );
  XOR U3553 ( .A(n2748), .B(n2749), .Z(n2563) );
  ANDN U3554 ( .B(n2750), .A(n2751), .Z(n2748) );
  AND U3555 ( .A(b[7]), .B(a[41]), .Z(n2747) );
  XNOR U3556 ( .A(n2752), .B(n2568), .Z(n2570) );
  XOR U3557 ( .A(n2753), .B(n2754), .Z(n2568) );
  ANDN U3558 ( .B(n2755), .A(n2756), .Z(n2753) );
  AND U3559 ( .A(b[6]), .B(a[42]), .Z(n2752) );
  XNOR U3560 ( .A(n2757), .B(n2573), .Z(n2575) );
  XOR U3561 ( .A(n2758), .B(n2759), .Z(n2573) );
  ANDN U3562 ( .B(n2760), .A(n2761), .Z(n2758) );
  AND U3563 ( .A(b[5]), .B(a[43]), .Z(n2757) );
  XNOR U3564 ( .A(n2762), .B(n2578), .Z(n2580) );
  XOR U3565 ( .A(n2763), .B(n2764), .Z(n2578) );
  ANDN U3566 ( .B(n2765), .A(n2766), .Z(n2763) );
  AND U3567 ( .A(b[4]), .B(a[44]), .Z(n2762) );
  XNOR U3568 ( .A(n2767), .B(n2768), .Z(n2592) );
  NANDN U3569 ( .A(n2769), .B(n2770), .Z(n2768) );
  XNOR U3570 ( .A(n2771), .B(n2583), .Z(n2585) );
  XNOR U3571 ( .A(n2772), .B(n2773), .Z(n2583) );
  AND U3572 ( .A(n2774), .B(n2775), .Z(n2772) );
  AND U3573 ( .A(b[3]), .B(a[45]), .Z(n2771) );
  XNOR U3574 ( .A(n2776), .B(n2777), .Z(swire[47]) );
  XOR U3575 ( .A(n2603), .B(n2778), .Z(n2777) );
  XOR U3576 ( .A(n2602), .B(n2776), .Z(n2778) );
  NAND U3577 ( .A(a[47]), .B(b[0]), .Z(n2602) );
  XNOR U3578 ( .A(n2769), .B(n2770), .Z(n2603) );
  XOR U3579 ( .A(n2767), .B(n2779), .Z(n2770) );
  NAND U3580 ( .A(a[46]), .B(b[1]), .Z(n2779) );
  XOR U3581 ( .A(n2775), .B(n2780), .Z(n2769) );
  XOR U3582 ( .A(n2767), .B(n2774), .Z(n2780) );
  XNOR U3583 ( .A(n2781), .B(n2773), .Z(n2774) );
  AND U3584 ( .A(b[2]), .B(a[45]), .Z(n2781) );
  NANDN U3585 ( .A(n2782), .B(n2783), .Z(n2767) );
  XOR U3586 ( .A(n2773), .B(n2765), .Z(n2784) );
  XNOR U3587 ( .A(n2764), .B(n2760), .Z(n2785) );
  XNOR U3588 ( .A(n2759), .B(n2755), .Z(n2786) );
  XNOR U3589 ( .A(n2754), .B(n2750), .Z(n2787) );
  XNOR U3590 ( .A(n2749), .B(n2745), .Z(n2788) );
  XNOR U3591 ( .A(n2744), .B(n2740), .Z(n2789) );
  XNOR U3592 ( .A(n2739), .B(n2735), .Z(n2790) );
  XNOR U3593 ( .A(n2734), .B(n2730), .Z(n2791) );
  XNOR U3594 ( .A(n2729), .B(n2725), .Z(n2792) );
  XNOR U3595 ( .A(n2724), .B(n2720), .Z(n2793) );
  XNOR U3596 ( .A(n2719), .B(n2715), .Z(n2794) );
  XNOR U3597 ( .A(n2714), .B(n2710), .Z(n2795) );
  XNOR U3598 ( .A(n2709), .B(n2705), .Z(n2796) );
  XNOR U3599 ( .A(n2704), .B(n2700), .Z(n2797) );
  XNOR U3600 ( .A(n2699), .B(n2695), .Z(n2798) );
  XNOR U3601 ( .A(n2694), .B(n2690), .Z(n2799) );
  XNOR U3602 ( .A(n2689), .B(n2685), .Z(n2800) );
  XNOR U3603 ( .A(n2684), .B(n2680), .Z(n2801) );
  XNOR U3604 ( .A(n2679), .B(n2675), .Z(n2802) );
  XNOR U3605 ( .A(n2674), .B(n2670), .Z(n2803) );
  XNOR U3606 ( .A(n2669), .B(n2665), .Z(n2804) );
  XNOR U3607 ( .A(n2664), .B(n2660), .Z(n2805) );
  XNOR U3608 ( .A(n2659), .B(n2655), .Z(n2806) );
  XNOR U3609 ( .A(n2654), .B(n2650), .Z(n2807) );
  XNOR U3610 ( .A(n2649), .B(n2645), .Z(n2808) );
  XOR U3611 ( .A(n2644), .B(n2641), .Z(n2809) );
  XOR U3612 ( .A(n2810), .B(n2811), .Z(n2641) );
  XOR U3613 ( .A(n2639), .B(n2812), .Z(n2811) );
  XOR U3614 ( .A(n2813), .B(n2814), .Z(n2812) );
  XOR U3615 ( .A(n2815), .B(n2816), .Z(n2814) );
  NAND U3616 ( .A(a[17]), .B(b[30]), .Z(n2816) );
  AND U3617 ( .A(a[16]), .B(b[31]), .Z(n2815) );
  XOR U3618 ( .A(n2817), .B(n2813), .Z(n2810) );
  XOR U3619 ( .A(n2818), .B(n2819), .Z(n2813) );
  NOR U3620 ( .A(n2820), .B(n2821), .Z(n2818) );
  AND U3621 ( .A(a[18]), .B(b[29]), .Z(n2817) );
  XNOR U3622 ( .A(n2822), .B(n2639), .Z(n2640) );
  XOR U3623 ( .A(n2823), .B(n2824), .Z(n2639) );
  ANDN U3624 ( .B(n2825), .A(n2826), .Z(n2823) );
  AND U3625 ( .A(a[19]), .B(b[28]), .Z(n2822) );
  XNOR U3626 ( .A(n2827), .B(n2644), .Z(n2646) );
  XOR U3627 ( .A(n2828), .B(n2829), .Z(n2644) );
  ANDN U3628 ( .B(n2830), .A(n2831), .Z(n2828) );
  AND U3629 ( .A(a[20]), .B(b[27]), .Z(n2827) );
  XNOR U3630 ( .A(n2832), .B(n2649), .Z(n2651) );
  XOR U3631 ( .A(n2833), .B(n2834), .Z(n2649) );
  ANDN U3632 ( .B(n2835), .A(n2836), .Z(n2833) );
  AND U3633 ( .A(a[21]), .B(b[26]), .Z(n2832) );
  XNOR U3634 ( .A(n2837), .B(n2654), .Z(n2656) );
  XOR U3635 ( .A(n2838), .B(n2839), .Z(n2654) );
  ANDN U3636 ( .B(n2840), .A(n2841), .Z(n2838) );
  AND U3637 ( .A(a[22]), .B(b[25]), .Z(n2837) );
  XNOR U3638 ( .A(n2842), .B(n2659), .Z(n2661) );
  XOR U3639 ( .A(n2843), .B(n2844), .Z(n2659) );
  ANDN U3640 ( .B(n2845), .A(n2846), .Z(n2843) );
  AND U3641 ( .A(a[23]), .B(b[24]), .Z(n2842) );
  XNOR U3642 ( .A(n2847), .B(n2664), .Z(n2666) );
  XOR U3643 ( .A(n2848), .B(n2849), .Z(n2664) );
  ANDN U3644 ( .B(n2850), .A(n2851), .Z(n2848) );
  AND U3645 ( .A(a[24]), .B(b[23]), .Z(n2847) );
  XNOR U3646 ( .A(n2852), .B(n2669), .Z(n2671) );
  XOR U3647 ( .A(n2853), .B(n2854), .Z(n2669) );
  ANDN U3648 ( .B(n2855), .A(n2856), .Z(n2853) );
  AND U3649 ( .A(b[22]), .B(a[25]), .Z(n2852) );
  XNOR U3650 ( .A(n2857), .B(n2674), .Z(n2676) );
  XOR U3651 ( .A(n2858), .B(n2859), .Z(n2674) );
  ANDN U3652 ( .B(n2860), .A(n2861), .Z(n2858) );
  AND U3653 ( .A(a[26]), .B(b[21]), .Z(n2857) );
  XNOR U3654 ( .A(n2862), .B(n2679), .Z(n2681) );
  XOR U3655 ( .A(n2863), .B(n2864), .Z(n2679) );
  ANDN U3656 ( .B(n2865), .A(n2866), .Z(n2863) );
  AND U3657 ( .A(b[20]), .B(a[27]), .Z(n2862) );
  XNOR U3658 ( .A(n2867), .B(n2684), .Z(n2686) );
  XOR U3659 ( .A(n2868), .B(n2869), .Z(n2684) );
  ANDN U3660 ( .B(n2870), .A(n2871), .Z(n2868) );
  AND U3661 ( .A(a[28]), .B(b[19]), .Z(n2867) );
  XNOR U3662 ( .A(n2872), .B(n2689), .Z(n2691) );
  XOR U3663 ( .A(n2873), .B(n2874), .Z(n2689) );
  ANDN U3664 ( .B(n2875), .A(n2876), .Z(n2873) );
  AND U3665 ( .A(b[18]), .B(a[29]), .Z(n2872) );
  XNOR U3666 ( .A(n2877), .B(n2694), .Z(n2696) );
  XOR U3667 ( .A(n2878), .B(n2879), .Z(n2694) );
  ANDN U3668 ( .B(n2880), .A(n2881), .Z(n2878) );
  AND U3669 ( .A(a[30]), .B(b[17]), .Z(n2877) );
  XNOR U3670 ( .A(n2882), .B(n2699), .Z(n2701) );
  XOR U3671 ( .A(n2883), .B(n2884), .Z(n2699) );
  ANDN U3672 ( .B(n2885), .A(n2886), .Z(n2883) );
  AND U3673 ( .A(b[16]), .B(a[31]), .Z(n2882) );
  XNOR U3674 ( .A(n2887), .B(n2704), .Z(n2706) );
  XOR U3675 ( .A(n2888), .B(n2889), .Z(n2704) );
  ANDN U3676 ( .B(n2890), .A(n2891), .Z(n2888) );
  AND U3677 ( .A(a[32]), .B(b[15]), .Z(n2887) );
  XNOR U3678 ( .A(n2892), .B(n2709), .Z(n2711) );
  XOR U3679 ( .A(n2893), .B(n2894), .Z(n2709) );
  ANDN U3680 ( .B(n2895), .A(n2896), .Z(n2893) );
  AND U3681 ( .A(b[14]), .B(a[33]), .Z(n2892) );
  XNOR U3682 ( .A(n2897), .B(n2714), .Z(n2716) );
  XOR U3683 ( .A(n2898), .B(n2899), .Z(n2714) );
  ANDN U3684 ( .B(n2900), .A(n2901), .Z(n2898) );
  AND U3685 ( .A(a[34]), .B(b[13]), .Z(n2897) );
  XNOR U3686 ( .A(n2902), .B(n2719), .Z(n2721) );
  XOR U3687 ( .A(n2903), .B(n2904), .Z(n2719) );
  ANDN U3688 ( .B(n2905), .A(n2906), .Z(n2903) );
  AND U3689 ( .A(b[12]), .B(a[35]), .Z(n2902) );
  XNOR U3690 ( .A(n2907), .B(n2724), .Z(n2726) );
  XOR U3691 ( .A(n2908), .B(n2909), .Z(n2724) );
  ANDN U3692 ( .B(n2910), .A(n2911), .Z(n2908) );
  AND U3693 ( .A(a[36]), .B(b[11]), .Z(n2907) );
  XNOR U3694 ( .A(n2912), .B(n2729), .Z(n2731) );
  XOR U3695 ( .A(n2913), .B(n2914), .Z(n2729) );
  ANDN U3696 ( .B(n2915), .A(n2916), .Z(n2913) );
  AND U3697 ( .A(b[10]), .B(a[37]), .Z(n2912) );
  XNOR U3698 ( .A(n2917), .B(n2734), .Z(n2736) );
  XOR U3699 ( .A(n2918), .B(n2919), .Z(n2734) );
  ANDN U3700 ( .B(n2920), .A(n2921), .Z(n2918) );
  AND U3701 ( .A(a[38]), .B(b[9]), .Z(n2917) );
  XNOR U3702 ( .A(n2922), .B(n2739), .Z(n2741) );
  XOR U3703 ( .A(n2923), .B(n2924), .Z(n2739) );
  ANDN U3704 ( .B(n2925), .A(n2926), .Z(n2923) );
  AND U3705 ( .A(b[8]), .B(a[39]), .Z(n2922) );
  XNOR U3706 ( .A(n2927), .B(n2744), .Z(n2746) );
  XOR U3707 ( .A(n2928), .B(n2929), .Z(n2744) );
  ANDN U3708 ( .B(n2930), .A(n2931), .Z(n2928) );
  AND U3709 ( .A(a[40]), .B(b[7]), .Z(n2927) );
  XNOR U3710 ( .A(n2932), .B(n2749), .Z(n2751) );
  XOR U3711 ( .A(n2933), .B(n2934), .Z(n2749) );
  ANDN U3712 ( .B(n2935), .A(n2936), .Z(n2933) );
  AND U3713 ( .A(b[6]), .B(a[41]), .Z(n2932) );
  XNOR U3714 ( .A(n2937), .B(n2754), .Z(n2756) );
  XOR U3715 ( .A(n2938), .B(n2939), .Z(n2754) );
  ANDN U3716 ( .B(n2940), .A(n2941), .Z(n2938) );
  AND U3717 ( .A(b[5]), .B(a[42]), .Z(n2937) );
  XNOR U3718 ( .A(n2942), .B(n2759), .Z(n2761) );
  XOR U3719 ( .A(n2943), .B(n2944), .Z(n2759) );
  ANDN U3720 ( .B(n2945), .A(n2946), .Z(n2943) );
  AND U3721 ( .A(b[4]), .B(a[43]), .Z(n2942) );
  XNOR U3722 ( .A(n2947), .B(n2948), .Z(n2773) );
  NANDN U3723 ( .A(n2949), .B(n2950), .Z(n2948) );
  XNOR U3724 ( .A(n2951), .B(n2764), .Z(n2766) );
  XNOR U3725 ( .A(n2952), .B(n2953), .Z(n2764) );
  AND U3726 ( .A(n2954), .B(n2955), .Z(n2952) );
  AND U3727 ( .A(b[3]), .B(a[44]), .Z(n2951) );
  XNOR U3728 ( .A(n2956), .B(n2957), .Z(swire[46]) );
  XOR U3729 ( .A(n2783), .B(n2959), .Z(n2957) );
  XNOR U3730 ( .A(n2782), .B(n2958), .Z(n2959) );
  IV U3731 ( .A(n2956), .Z(n2958) );
  NAND U3732 ( .A(a[46]), .B(b[0]), .Z(n2782) );
  XNOR U3733 ( .A(n2949), .B(n2950), .Z(n2783) );
  XOR U3734 ( .A(n2947), .B(n2960), .Z(n2950) );
  NAND U3735 ( .A(b[1]), .B(a[45]), .Z(n2960) );
  XOR U3736 ( .A(n2955), .B(n2961), .Z(n2949) );
  XOR U3737 ( .A(n2947), .B(n2954), .Z(n2961) );
  XNOR U3738 ( .A(n2962), .B(n2953), .Z(n2954) );
  AND U3739 ( .A(b[2]), .B(a[44]), .Z(n2962) );
  NANDN U3740 ( .A(n2963), .B(n2964), .Z(n2947) );
  XOR U3741 ( .A(n2953), .B(n2945), .Z(n2965) );
  XNOR U3742 ( .A(n2944), .B(n2940), .Z(n2966) );
  XNOR U3743 ( .A(n2939), .B(n2935), .Z(n2967) );
  XNOR U3744 ( .A(n2934), .B(n2930), .Z(n2968) );
  XNOR U3745 ( .A(n2929), .B(n2925), .Z(n2969) );
  XNOR U3746 ( .A(n2924), .B(n2920), .Z(n2970) );
  XNOR U3747 ( .A(n2919), .B(n2915), .Z(n2971) );
  XNOR U3748 ( .A(n2914), .B(n2910), .Z(n2972) );
  XNOR U3749 ( .A(n2909), .B(n2905), .Z(n2973) );
  XNOR U3750 ( .A(n2904), .B(n2900), .Z(n2974) );
  XNOR U3751 ( .A(n2899), .B(n2895), .Z(n2975) );
  XNOR U3752 ( .A(n2894), .B(n2890), .Z(n2976) );
  XNOR U3753 ( .A(n2889), .B(n2885), .Z(n2977) );
  XNOR U3754 ( .A(n2884), .B(n2880), .Z(n2978) );
  XNOR U3755 ( .A(n2879), .B(n2875), .Z(n2979) );
  XNOR U3756 ( .A(n2874), .B(n2870), .Z(n2980) );
  XNOR U3757 ( .A(n2869), .B(n2865), .Z(n2981) );
  XNOR U3758 ( .A(n2864), .B(n2860), .Z(n2982) );
  XNOR U3759 ( .A(n2859), .B(n2855), .Z(n2983) );
  XNOR U3760 ( .A(n2854), .B(n2850), .Z(n2984) );
  XNOR U3761 ( .A(n2849), .B(n2845), .Z(n2985) );
  XNOR U3762 ( .A(n2844), .B(n2840), .Z(n2986) );
  XNOR U3763 ( .A(n2839), .B(n2835), .Z(n2987) );
  XNOR U3764 ( .A(n2834), .B(n2830), .Z(n2988) );
  XNOR U3765 ( .A(n2829), .B(n2825), .Z(n2989) );
  XOR U3766 ( .A(n2824), .B(n2821), .Z(n2990) );
  XOR U3767 ( .A(n2991), .B(n2992), .Z(n2821) );
  XOR U3768 ( .A(n2819), .B(n2993), .Z(n2992) );
  XOR U3769 ( .A(n2994), .B(n2995), .Z(n2993) );
  XOR U3770 ( .A(n2996), .B(n2997), .Z(n2995) );
  NAND U3771 ( .A(a[16]), .B(b[30]), .Z(n2997) );
  AND U3772 ( .A(a[15]), .B(b[31]), .Z(n2996) );
  XOR U3773 ( .A(n2998), .B(n2994), .Z(n2991) );
  XOR U3774 ( .A(n2999), .B(n3000), .Z(n2994) );
  NOR U3775 ( .A(n3001), .B(n3002), .Z(n2999) );
  AND U3776 ( .A(a[17]), .B(b[29]), .Z(n2998) );
  XNOR U3777 ( .A(n3003), .B(n2819), .Z(n2820) );
  XOR U3778 ( .A(n3004), .B(n3005), .Z(n2819) );
  ANDN U3779 ( .B(n3006), .A(n3007), .Z(n3004) );
  AND U3780 ( .A(a[18]), .B(b[28]), .Z(n3003) );
  XNOR U3781 ( .A(n3008), .B(n2824), .Z(n2826) );
  XOR U3782 ( .A(n3009), .B(n3010), .Z(n2824) );
  ANDN U3783 ( .B(n3011), .A(n3012), .Z(n3009) );
  AND U3784 ( .A(a[19]), .B(b[27]), .Z(n3008) );
  XNOR U3785 ( .A(n3013), .B(n2829), .Z(n2831) );
  XOR U3786 ( .A(n3014), .B(n3015), .Z(n2829) );
  ANDN U3787 ( .B(n3016), .A(n3017), .Z(n3014) );
  AND U3788 ( .A(a[20]), .B(b[26]), .Z(n3013) );
  XNOR U3789 ( .A(n3018), .B(n2834), .Z(n2836) );
  XOR U3790 ( .A(n3019), .B(n3020), .Z(n2834) );
  ANDN U3791 ( .B(n3021), .A(n3022), .Z(n3019) );
  AND U3792 ( .A(a[21]), .B(b[25]), .Z(n3018) );
  XNOR U3793 ( .A(n3023), .B(n2839), .Z(n2841) );
  XOR U3794 ( .A(n3024), .B(n3025), .Z(n2839) );
  ANDN U3795 ( .B(n3026), .A(n3027), .Z(n3024) );
  AND U3796 ( .A(a[22]), .B(b[24]), .Z(n3023) );
  XNOR U3797 ( .A(n3028), .B(n2844), .Z(n2846) );
  XOR U3798 ( .A(n3029), .B(n3030), .Z(n2844) );
  ANDN U3799 ( .B(n3031), .A(n3032), .Z(n3029) );
  AND U3800 ( .A(b[23]), .B(a[23]), .Z(n3028) );
  XNOR U3801 ( .A(n3033), .B(n2849), .Z(n2851) );
  XOR U3802 ( .A(n3034), .B(n3035), .Z(n2849) );
  ANDN U3803 ( .B(n3036), .A(n3037), .Z(n3034) );
  AND U3804 ( .A(a[24]), .B(b[22]), .Z(n3033) );
  XNOR U3805 ( .A(n3038), .B(n2854), .Z(n2856) );
  XOR U3806 ( .A(n3039), .B(n3040), .Z(n2854) );
  ANDN U3807 ( .B(n3041), .A(n3042), .Z(n3039) );
  AND U3808 ( .A(b[21]), .B(a[25]), .Z(n3038) );
  XNOR U3809 ( .A(n3043), .B(n2859), .Z(n2861) );
  XOR U3810 ( .A(n3044), .B(n3045), .Z(n2859) );
  ANDN U3811 ( .B(n3046), .A(n3047), .Z(n3044) );
  AND U3812 ( .A(a[26]), .B(b[20]), .Z(n3043) );
  XNOR U3813 ( .A(n3048), .B(n2864), .Z(n2866) );
  XOR U3814 ( .A(n3049), .B(n3050), .Z(n2864) );
  ANDN U3815 ( .B(n3051), .A(n3052), .Z(n3049) );
  AND U3816 ( .A(b[19]), .B(a[27]), .Z(n3048) );
  XNOR U3817 ( .A(n3053), .B(n2869), .Z(n2871) );
  XOR U3818 ( .A(n3054), .B(n3055), .Z(n2869) );
  ANDN U3819 ( .B(n3056), .A(n3057), .Z(n3054) );
  AND U3820 ( .A(a[28]), .B(b[18]), .Z(n3053) );
  XNOR U3821 ( .A(n3058), .B(n2874), .Z(n2876) );
  XOR U3822 ( .A(n3059), .B(n3060), .Z(n2874) );
  ANDN U3823 ( .B(n3061), .A(n3062), .Z(n3059) );
  AND U3824 ( .A(b[17]), .B(a[29]), .Z(n3058) );
  XNOR U3825 ( .A(n3063), .B(n2879), .Z(n2881) );
  XOR U3826 ( .A(n3064), .B(n3065), .Z(n2879) );
  ANDN U3827 ( .B(n3066), .A(n3067), .Z(n3064) );
  AND U3828 ( .A(a[30]), .B(b[16]), .Z(n3063) );
  XNOR U3829 ( .A(n3068), .B(n2884), .Z(n2886) );
  XOR U3830 ( .A(n3069), .B(n3070), .Z(n2884) );
  ANDN U3831 ( .B(n3071), .A(n3072), .Z(n3069) );
  AND U3832 ( .A(b[15]), .B(a[31]), .Z(n3068) );
  XNOR U3833 ( .A(n3073), .B(n2889), .Z(n2891) );
  XOR U3834 ( .A(n3074), .B(n3075), .Z(n2889) );
  ANDN U3835 ( .B(n3076), .A(n3077), .Z(n3074) );
  AND U3836 ( .A(a[32]), .B(b[14]), .Z(n3073) );
  XNOR U3837 ( .A(n3078), .B(n2894), .Z(n2896) );
  XOR U3838 ( .A(n3079), .B(n3080), .Z(n2894) );
  ANDN U3839 ( .B(n3081), .A(n3082), .Z(n3079) );
  AND U3840 ( .A(b[13]), .B(a[33]), .Z(n3078) );
  XNOR U3841 ( .A(n3083), .B(n2899), .Z(n2901) );
  XOR U3842 ( .A(n3084), .B(n3085), .Z(n2899) );
  ANDN U3843 ( .B(n3086), .A(n3087), .Z(n3084) );
  AND U3844 ( .A(a[34]), .B(b[12]), .Z(n3083) );
  XNOR U3845 ( .A(n3088), .B(n2904), .Z(n2906) );
  XOR U3846 ( .A(n3089), .B(n3090), .Z(n2904) );
  ANDN U3847 ( .B(n3091), .A(n3092), .Z(n3089) );
  AND U3848 ( .A(b[11]), .B(a[35]), .Z(n3088) );
  XNOR U3849 ( .A(n3093), .B(n2909), .Z(n2911) );
  XOR U3850 ( .A(n3094), .B(n3095), .Z(n2909) );
  ANDN U3851 ( .B(n3096), .A(n3097), .Z(n3094) );
  AND U3852 ( .A(a[36]), .B(b[10]), .Z(n3093) );
  XNOR U3853 ( .A(n3098), .B(n2914), .Z(n2916) );
  XOR U3854 ( .A(n3099), .B(n3100), .Z(n2914) );
  ANDN U3855 ( .B(n3101), .A(n3102), .Z(n3099) );
  AND U3856 ( .A(b[9]), .B(a[37]), .Z(n3098) );
  XNOR U3857 ( .A(n3103), .B(n2919), .Z(n2921) );
  XOR U3858 ( .A(n3104), .B(n3105), .Z(n2919) );
  ANDN U3859 ( .B(n3106), .A(n3107), .Z(n3104) );
  AND U3860 ( .A(a[38]), .B(b[8]), .Z(n3103) );
  XNOR U3861 ( .A(n3108), .B(n2924), .Z(n2926) );
  XOR U3862 ( .A(n3109), .B(n3110), .Z(n2924) );
  ANDN U3863 ( .B(n3111), .A(n3112), .Z(n3109) );
  AND U3864 ( .A(b[7]), .B(a[39]), .Z(n3108) );
  XNOR U3865 ( .A(n3113), .B(n2929), .Z(n2931) );
  XOR U3866 ( .A(n3114), .B(n3115), .Z(n2929) );
  ANDN U3867 ( .B(n3116), .A(n3117), .Z(n3114) );
  AND U3868 ( .A(b[6]), .B(a[40]), .Z(n3113) );
  XNOR U3869 ( .A(n3118), .B(n2934), .Z(n2936) );
  XOR U3870 ( .A(n3119), .B(n3120), .Z(n2934) );
  ANDN U3871 ( .B(n3121), .A(n3122), .Z(n3119) );
  AND U3872 ( .A(b[5]), .B(a[41]), .Z(n3118) );
  XNOR U3873 ( .A(n3123), .B(n2939), .Z(n2941) );
  XOR U3874 ( .A(n3124), .B(n3125), .Z(n2939) );
  ANDN U3875 ( .B(n3126), .A(n3127), .Z(n3124) );
  AND U3876 ( .A(b[4]), .B(a[42]), .Z(n3123) );
  XNOR U3877 ( .A(n3128), .B(n3129), .Z(n2953) );
  NANDN U3878 ( .A(n3130), .B(n3131), .Z(n3129) );
  XNOR U3879 ( .A(n3132), .B(n2944), .Z(n2946) );
  XNOR U3880 ( .A(n3133), .B(n3134), .Z(n2944) );
  AND U3881 ( .A(n3135), .B(n3136), .Z(n3133) );
  AND U3882 ( .A(b[3]), .B(a[43]), .Z(n3132) );
  XNOR U3883 ( .A(n3137), .B(n3138), .Z(swire[45]) );
  XOR U3884 ( .A(n2964), .B(n3139), .Z(n3138) );
  XOR U3885 ( .A(n2963), .B(n3137), .Z(n3139) );
  NAND U3886 ( .A(a[45]), .B(b[0]), .Z(n2963) );
  XNOR U3887 ( .A(n3130), .B(n3131), .Z(n2964) );
  XOR U3888 ( .A(n3128), .B(n3140), .Z(n3131) );
  NAND U3889 ( .A(a[44]), .B(b[1]), .Z(n3140) );
  XOR U3890 ( .A(n3136), .B(n3141), .Z(n3130) );
  XOR U3891 ( .A(n3128), .B(n3135), .Z(n3141) );
  XNOR U3892 ( .A(n3142), .B(n3134), .Z(n3135) );
  AND U3893 ( .A(b[2]), .B(a[43]), .Z(n3142) );
  NANDN U3894 ( .A(n3143), .B(n3144), .Z(n3128) );
  XOR U3895 ( .A(n3134), .B(n3126), .Z(n3145) );
  XNOR U3896 ( .A(n3125), .B(n3121), .Z(n3146) );
  XNOR U3897 ( .A(n3120), .B(n3116), .Z(n3147) );
  XNOR U3898 ( .A(n3115), .B(n3111), .Z(n3148) );
  XNOR U3899 ( .A(n3110), .B(n3106), .Z(n3149) );
  XNOR U3900 ( .A(n3105), .B(n3101), .Z(n3150) );
  XNOR U3901 ( .A(n3100), .B(n3096), .Z(n3151) );
  XNOR U3902 ( .A(n3095), .B(n3091), .Z(n3152) );
  XNOR U3903 ( .A(n3090), .B(n3086), .Z(n3153) );
  XNOR U3904 ( .A(n3085), .B(n3081), .Z(n3154) );
  XNOR U3905 ( .A(n3080), .B(n3076), .Z(n3155) );
  XNOR U3906 ( .A(n3075), .B(n3071), .Z(n3156) );
  XNOR U3907 ( .A(n3070), .B(n3066), .Z(n3157) );
  XNOR U3908 ( .A(n3065), .B(n3061), .Z(n3158) );
  XNOR U3909 ( .A(n3060), .B(n3056), .Z(n3159) );
  XNOR U3910 ( .A(n3055), .B(n3051), .Z(n3160) );
  XNOR U3911 ( .A(n3050), .B(n3046), .Z(n3161) );
  XNOR U3912 ( .A(n3045), .B(n3041), .Z(n3162) );
  XNOR U3913 ( .A(n3040), .B(n3036), .Z(n3163) );
  XNOR U3914 ( .A(n3035), .B(n3031), .Z(n3164) );
  XNOR U3915 ( .A(n3030), .B(n3026), .Z(n3165) );
  XNOR U3916 ( .A(n3025), .B(n3021), .Z(n3166) );
  XNOR U3917 ( .A(n3020), .B(n3016), .Z(n3167) );
  XNOR U3918 ( .A(n3015), .B(n3011), .Z(n3168) );
  XNOR U3919 ( .A(n3010), .B(n3006), .Z(n3169) );
  XOR U3920 ( .A(n3005), .B(n3002), .Z(n3170) );
  XOR U3921 ( .A(n3171), .B(n3172), .Z(n3002) );
  XOR U3922 ( .A(n3000), .B(n3173), .Z(n3172) );
  XOR U3923 ( .A(n3174), .B(n3175), .Z(n3173) );
  XOR U3924 ( .A(n3176), .B(n3177), .Z(n3175) );
  NAND U3925 ( .A(a[15]), .B(b[30]), .Z(n3177) );
  AND U3926 ( .A(a[14]), .B(b[31]), .Z(n3176) );
  XOR U3927 ( .A(n3178), .B(n3174), .Z(n3171) );
  XOR U3928 ( .A(n3179), .B(n3180), .Z(n3174) );
  NOR U3929 ( .A(n3181), .B(n3182), .Z(n3179) );
  AND U3930 ( .A(a[16]), .B(b[29]), .Z(n3178) );
  XNOR U3931 ( .A(n3183), .B(n3000), .Z(n3001) );
  XOR U3932 ( .A(n3184), .B(n3185), .Z(n3000) );
  ANDN U3933 ( .B(n3186), .A(n3187), .Z(n3184) );
  AND U3934 ( .A(a[17]), .B(b[28]), .Z(n3183) );
  XNOR U3935 ( .A(n3188), .B(n3005), .Z(n3007) );
  XOR U3936 ( .A(n3189), .B(n3190), .Z(n3005) );
  ANDN U3937 ( .B(n3191), .A(n3192), .Z(n3189) );
  AND U3938 ( .A(a[18]), .B(b[27]), .Z(n3188) );
  XNOR U3939 ( .A(n3193), .B(n3010), .Z(n3012) );
  XOR U3940 ( .A(n3194), .B(n3195), .Z(n3010) );
  ANDN U3941 ( .B(n3196), .A(n3197), .Z(n3194) );
  AND U3942 ( .A(a[19]), .B(b[26]), .Z(n3193) );
  XNOR U3943 ( .A(n3198), .B(n3015), .Z(n3017) );
  XOR U3944 ( .A(n3199), .B(n3200), .Z(n3015) );
  ANDN U3945 ( .B(n3201), .A(n3202), .Z(n3199) );
  AND U3946 ( .A(a[20]), .B(b[25]), .Z(n3198) );
  XNOR U3947 ( .A(n3203), .B(n3020), .Z(n3022) );
  XOR U3948 ( .A(n3204), .B(n3205), .Z(n3020) );
  ANDN U3949 ( .B(n3206), .A(n3207), .Z(n3204) );
  AND U3950 ( .A(a[21]), .B(b[24]), .Z(n3203) );
  XNOR U3951 ( .A(n3208), .B(n3025), .Z(n3027) );
  XOR U3952 ( .A(n3209), .B(n3210), .Z(n3025) );
  ANDN U3953 ( .B(n3211), .A(n3212), .Z(n3209) );
  AND U3954 ( .A(a[22]), .B(b[23]), .Z(n3208) );
  XNOR U3955 ( .A(n3213), .B(n3030), .Z(n3032) );
  XOR U3956 ( .A(n3214), .B(n3215), .Z(n3030) );
  ANDN U3957 ( .B(n3216), .A(n3217), .Z(n3214) );
  AND U3958 ( .A(b[22]), .B(a[23]), .Z(n3213) );
  XNOR U3959 ( .A(n3218), .B(n3035), .Z(n3037) );
  XOR U3960 ( .A(n3219), .B(n3220), .Z(n3035) );
  ANDN U3961 ( .B(n3221), .A(n3222), .Z(n3219) );
  AND U3962 ( .A(a[24]), .B(b[21]), .Z(n3218) );
  XNOR U3963 ( .A(n3223), .B(n3040), .Z(n3042) );
  XOR U3964 ( .A(n3224), .B(n3225), .Z(n3040) );
  ANDN U3965 ( .B(n3226), .A(n3227), .Z(n3224) );
  AND U3966 ( .A(b[20]), .B(a[25]), .Z(n3223) );
  XNOR U3967 ( .A(n3228), .B(n3045), .Z(n3047) );
  XOR U3968 ( .A(n3229), .B(n3230), .Z(n3045) );
  ANDN U3969 ( .B(n3231), .A(n3232), .Z(n3229) );
  AND U3970 ( .A(a[26]), .B(b[19]), .Z(n3228) );
  XNOR U3971 ( .A(n3233), .B(n3050), .Z(n3052) );
  XOR U3972 ( .A(n3234), .B(n3235), .Z(n3050) );
  ANDN U3973 ( .B(n3236), .A(n3237), .Z(n3234) );
  AND U3974 ( .A(b[18]), .B(a[27]), .Z(n3233) );
  XNOR U3975 ( .A(n3238), .B(n3055), .Z(n3057) );
  XOR U3976 ( .A(n3239), .B(n3240), .Z(n3055) );
  ANDN U3977 ( .B(n3241), .A(n3242), .Z(n3239) );
  AND U3978 ( .A(a[28]), .B(b[17]), .Z(n3238) );
  XNOR U3979 ( .A(n3243), .B(n3060), .Z(n3062) );
  XOR U3980 ( .A(n3244), .B(n3245), .Z(n3060) );
  ANDN U3981 ( .B(n3246), .A(n3247), .Z(n3244) );
  AND U3982 ( .A(b[16]), .B(a[29]), .Z(n3243) );
  XNOR U3983 ( .A(n3248), .B(n3065), .Z(n3067) );
  XOR U3984 ( .A(n3249), .B(n3250), .Z(n3065) );
  ANDN U3985 ( .B(n3251), .A(n3252), .Z(n3249) );
  AND U3986 ( .A(a[30]), .B(b[15]), .Z(n3248) );
  XNOR U3987 ( .A(n3253), .B(n3070), .Z(n3072) );
  XOR U3988 ( .A(n3254), .B(n3255), .Z(n3070) );
  ANDN U3989 ( .B(n3256), .A(n3257), .Z(n3254) );
  AND U3990 ( .A(b[14]), .B(a[31]), .Z(n3253) );
  XNOR U3991 ( .A(n3258), .B(n3075), .Z(n3077) );
  XOR U3992 ( .A(n3259), .B(n3260), .Z(n3075) );
  ANDN U3993 ( .B(n3261), .A(n3262), .Z(n3259) );
  AND U3994 ( .A(a[32]), .B(b[13]), .Z(n3258) );
  XNOR U3995 ( .A(n3263), .B(n3080), .Z(n3082) );
  XOR U3996 ( .A(n3264), .B(n3265), .Z(n3080) );
  ANDN U3997 ( .B(n3266), .A(n3267), .Z(n3264) );
  AND U3998 ( .A(b[12]), .B(a[33]), .Z(n3263) );
  XNOR U3999 ( .A(n3268), .B(n3085), .Z(n3087) );
  XOR U4000 ( .A(n3269), .B(n3270), .Z(n3085) );
  ANDN U4001 ( .B(n3271), .A(n3272), .Z(n3269) );
  AND U4002 ( .A(a[34]), .B(b[11]), .Z(n3268) );
  XNOR U4003 ( .A(n3273), .B(n3090), .Z(n3092) );
  XOR U4004 ( .A(n3274), .B(n3275), .Z(n3090) );
  ANDN U4005 ( .B(n3276), .A(n3277), .Z(n3274) );
  AND U4006 ( .A(b[10]), .B(a[35]), .Z(n3273) );
  XNOR U4007 ( .A(n3278), .B(n3095), .Z(n3097) );
  XOR U4008 ( .A(n3279), .B(n3280), .Z(n3095) );
  ANDN U4009 ( .B(n3281), .A(n3282), .Z(n3279) );
  AND U4010 ( .A(a[36]), .B(b[9]), .Z(n3278) );
  XNOR U4011 ( .A(n3283), .B(n3100), .Z(n3102) );
  XOR U4012 ( .A(n3284), .B(n3285), .Z(n3100) );
  ANDN U4013 ( .B(n3286), .A(n3287), .Z(n3284) );
  AND U4014 ( .A(b[8]), .B(a[37]), .Z(n3283) );
  XNOR U4015 ( .A(n3288), .B(n3105), .Z(n3107) );
  XOR U4016 ( .A(n3289), .B(n3290), .Z(n3105) );
  ANDN U4017 ( .B(n3291), .A(n3292), .Z(n3289) );
  AND U4018 ( .A(a[38]), .B(b[7]), .Z(n3288) );
  XNOR U4019 ( .A(n3293), .B(n3110), .Z(n3112) );
  XOR U4020 ( .A(n3294), .B(n3295), .Z(n3110) );
  ANDN U4021 ( .B(n3296), .A(n3297), .Z(n3294) );
  AND U4022 ( .A(b[6]), .B(a[39]), .Z(n3293) );
  XNOR U4023 ( .A(n3298), .B(n3115), .Z(n3117) );
  XOR U4024 ( .A(n3299), .B(n3300), .Z(n3115) );
  ANDN U4025 ( .B(n3301), .A(n3302), .Z(n3299) );
  AND U4026 ( .A(b[5]), .B(a[40]), .Z(n3298) );
  XNOR U4027 ( .A(n3303), .B(n3120), .Z(n3122) );
  XOR U4028 ( .A(n3304), .B(n3305), .Z(n3120) );
  ANDN U4029 ( .B(n3306), .A(n3307), .Z(n3304) );
  AND U4030 ( .A(b[4]), .B(a[41]), .Z(n3303) );
  XNOR U4031 ( .A(n3308), .B(n3309), .Z(n3134) );
  NANDN U4032 ( .A(n3310), .B(n3311), .Z(n3309) );
  XNOR U4033 ( .A(n3312), .B(n3125), .Z(n3127) );
  XNOR U4034 ( .A(n3313), .B(n3314), .Z(n3125) );
  AND U4035 ( .A(n3315), .B(n3316), .Z(n3313) );
  AND U4036 ( .A(b[3]), .B(a[42]), .Z(n3312) );
  XNOR U4037 ( .A(n3317), .B(n3318), .Z(swire[44]) );
  XOR U4038 ( .A(n3144), .B(n3320), .Z(n3318) );
  XNOR U4039 ( .A(n3143), .B(n3319), .Z(n3320) );
  IV U4040 ( .A(n3317), .Z(n3319) );
  NAND U4041 ( .A(a[44]), .B(b[0]), .Z(n3143) );
  XNOR U4042 ( .A(n3310), .B(n3311), .Z(n3144) );
  XOR U4043 ( .A(n3308), .B(n3321), .Z(n3311) );
  NAND U4044 ( .A(b[1]), .B(a[43]), .Z(n3321) );
  XOR U4045 ( .A(n3316), .B(n3322), .Z(n3310) );
  XOR U4046 ( .A(n3308), .B(n3315), .Z(n3322) );
  XNOR U4047 ( .A(n3323), .B(n3314), .Z(n3315) );
  AND U4048 ( .A(b[2]), .B(a[42]), .Z(n3323) );
  NANDN U4049 ( .A(n3324), .B(n3325), .Z(n3308) );
  XOR U4050 ( .A(n3314), .B(n3306), .Z(n3326) );
  XNOR U4051 ( .A(n3305), .B(n3301), .Z(n3327) );
  XNOR U4052 ( .A(n3300), .B(n3296), .Z(n3328) );
  XNOR U4053 ( .A(n3295), .B(n3291), .Z(n3329) );
  XNOR U4054 ( .A(n3290), .B(n3286), .Z(n3330) );
  XNOR U4055 ( .A(n3285), .B(n3281), .Z(n3331) );
  XNOR U4056 ( .A(n3280), .B(n3276), .Z(n3332) );
  XNOR U4057 ( .A(n3275), .B(n3271), .Z(n3333) );
  XNOR U4058 ( .A(n3270), .B(n3266), .Z(n3334) );
  XNOR U4059 ( .A(n3265), .B(n3261), .Z(n3335) );
  XNOR U4060 ( .A(n3260), .B(n3256), .Z(n3336) );
  XNOR U4061 ( .A(n3255), .B(n3251), .Z(n3337) );
  XNOR U4062 ( .A(n3250), .B(n3246), .Z(n3338) );
  XNOR U4063 ( .A(n3245), .B(n3241), .Z(n3339) );
  XNOR U4064 ( .A(n3240), .B(n3236), .Z(n3340) );
  XNOR U4065 ( .A(n3235), .B(n3231), .Z(n3341) );
  XNOR U4066 ( .A(n3230), .B(n3226), .Z(n3342) );
  XNOR U4067 ( .A(n3225), .B(n3221), .Z(n3343) );
  XNOR U4068 ( .A(n3220), .B(n3216), .Z(n3344) );
  XNOR U4069 ( .A(n3215), .B(n3211), .Z(n3345) );
  XNOR U4070 ( .A(n3210), .B(n3206), .Z(n3346) );
  XNOR U4071 ( .A(n3205), .B(n3201), .Z(n3347) );
  XNOR U4072 ( .A(n3200), .B(n3196), .Z(n3348) );
  XNOR U4073 ( .A(n3195), .B(n3191), .Z(n3349) );
  XNOR U4074 ( .A(n3190), .B(n3186), .Z(n3350) );
  XOR U4075 ( .A(n3185), .B(n3182), .Z(n3351) );
  XOR U4076 ( .A(n3352), .B(n3353), .Z(n3182) );
  XOR U4077 ( .A(n3180), .B(n3354), .Z(n3353) );
  XOR U4078 ( .A(n3355), .B(n3356), .Z(n3354) );
  XOR U4079 ( .A(n3357), .B(n3358), .Z(n3356) );
  NAND U4080 ( .A(a[14]), .B(b[30]), .Z(n3358) );
  AND U4081 ( .A(a[13]), .B(b[31]), .Z(n3357) );
  XOR U4082 ( .A(n3359), .B(n3355), .Z(n3352) );
  XOR U4083 ( .A(n3360), .B(n3361), .Z(n3355) );
  NOR U4084 ( .A(n3362), .B(n3363), .Z(n3360) );
  AND U4085 ( .A(a[15]), .B(b[29]), .Z(n3359) );
  XNOR U4086 ( .A(n3364), .B(n3180), .Z(n3181) );
  XOR U4087 ( .A(n3365), .B(n3366), .Z(n3180) );
  ANDN U4088 ( .B(n3367), .A(n3368), .Z(n3365) );
  AND U4089 ( .A(a[16]), .B(b[28]), .Z(n3364) );
  XNOR U4090 ( .A(n3369), .B(n3185), .Z(n3187) );
  XOR U4091 ( .A(n3370), .B(n3371), .Z(n3185) );
  ANDN U4092 ( .B(n3372), .A(n3373), .Z(n3370) );
  AND U4093 ( .A(a[17]), .B(b[27]), .Z(n3369) );
  XNOR U4094 ( .A(n3374), .B(n3190), .Z(n3192) );
  XOR U4095 ( .A(n3375), .B(n3376), .Z(n3190) );
  ANDN U4096 ( .B(n3377), .A(n3378), .Z(n3375) );
  AND U4097 ( .A(a[18]), .B(b[26]), .Z(n3374) );
  XNOR U4098 ( .A(n3379), .B(n3195), .Z(n3197) );
  XOR U4099 ( .A(n3380), .B(n3381), .Z(n3195) );
  ANDN U4100 ( .B(n3382), .A(n3383), .Z(n3380) );
  AND U4101 ( .A(a[19]), .B(b[25]), .Z(n3379) );
  XNOR U4102 ( .A(n3384), .B(n3200), .Z(n3202) );
  XOR U4103 ( .A(n3385), .B(n3386), .Z(n3200) );
  ANDN U4104 ( .B(n3387), .A(n3388), .Z(n3385) );
  AND U4105 ( .A(a[20]), .B(b[24]), .Z(n3384) );
  XNOR U4106 ( .A(n3389), .B(n3205), .Z(n3207) );
  XOR U4107 ( .A(n3390), .B(n3391), .Z(n3205) );
  ANDN U4108 ( .B(n3392), .A(n3393), .Z(n3390) );
  AND U4109 ( .A(a[21]), .B(b[23]), .Z(n3389) );
  XNOR U4110 ( .A(n3394), .B(n3210), .Z(n3212) );
  XOR U4111 ( .A(n3395), .B(n3396), .Z(n3210) );
  ANDN U4112 ( .B(n3397), .A(n3398), .Z(n3395) );
  AND U4113 ( .A(a[22]), .B(b[22]), .Z(n3394) );
  XNOR U4114 ( .A(n3399), .B(n3215), .Z(n3217) );
  XOR U4115 ( .A(n3400), .B(n3401), .Z(n3215) );
  ANDN U4116 ( .B(n3402), .A(n3403), .Z(n3400) );
  AND U4117 ( .A(b[21]), .B(a[23]), .Z(n3399) );
  XNOR U4118 ( .A(n3404), .B(n3220), .Z(n3222) );
  XOR U4119 ( .A(n3405), .B(n3406), .Z(n3220) );
  ANDN U4120 ( .B(n3407), .A(n3408), .Z(n3405) );
  AND U4121 ( .A(a[24]), .B(b[20]), .Z(n3404) );
  XNOR U4122 ( .A(n3409), .B(n3225), .Z(n3227) );
  XOR U4123 ( .A(n3410), .B(n3411), .Z(n3225) );
  ANDN U4124 ( .B(n3412), .A(n3413), .Z(n3410) );
  AND U4125 ( .A(b[19]), .B(a[25]), .Z(n3409) );
  XNOR U4126 ( .A(n3414), .B(n3230), .Z(n3232) );
  XOR U4127 ( .A(n3415), .B(n3416), .Z(n3230) );
  ANDN U4128 ( .B(n3417), .A(n3418), .Z(n3415) );
  AND U4129 ( .A(a[26]), .B(b[18]), .Z(n3414) );
  XNOR U4130 ( .A(n3419), .B(n3235), .Z(n3237) );
  XOR U4131 ( .A(n3420), .B(n3421), .Z(n3235) );
  ANDN U4132 ( .B(n3422), .A(n3423), .Z(n3420) );
  AND U4133 ( .A(b[17]), .B(a[27]), .Z(n3419) );
  XNOR U4134 ( .A(n3424), .B(n3240), .Z(n3242) );
  XOR U4135 ( .A(n3425), .B(n3426), .Z(n3240) );
  ANDN U4136 ( .B(n3427), .A(n3428), .Z(n3425) );
  AND U4137 ( .A(a[28]), .B(b[16]), .Z(n3424) );
  XNOR U4138 ( .A(n3429), .B(n3245), .Z(n3247) );
  XOR U4139 ( .A(n3430), .B(n3431), .Z(n3245) );
  ANDN U4140 ( .B(n3432), .A(n3433), .Z(n3430) );
  AND U4141 ( .A(b[15]), .B(a[29]), .Z(n3429) );
  XNOR U4142 ( .A(n3434), .B(n3250), .Z(n3252) );
  XOR U4143 ( .A(n3435), .B(n3436), .Z(n3250) );
  ANDN U4144 ( .B(n3437), .A(n3438), .Z(n3435) );
  AND U4145 ( .A(a[30]), .B(b[14]), .Z(n3434) );
  XNOR U4146 ( .A(n3439), .B(n3255), .Z(n3257) );
  XOR U4147 ( .A(n3440), .B(n3441), .Z(n3255) );
  ANDN U4148 ( .B(n3442), .A(n3443), .Z(n3440) );
  AND U4149 ( .A(b[13]), .B(a[31]), .Z(n3439) );
  XNOR U4150 ( .A(n3444), .B(n3260), .Z(n3262) );
  XOR U4151 ( .A(n3445), .B(n3446), .Z(n3260) );
  ANDN U4152 ( .B(n3447), .A(n3448), .Z(n3445) );
  AND U4153 ( .A(a[32]), .B(b[12]), .Z(n3444) );
  XNOR U4154 ( .A(n3449), .B(n3265), .Z(n3267) );
  XOR U4155 ( .A(n3450), .B(n3451), .Z(n3265) );
  ANDN U4156 ( .B(n3452), .A(n3453), .Z(n3450) );
  AND U4157 ( .A(b[11]), .B(a[33]), .Z(n3449) );
  XNOR U4158 ( .A(n3454), .B(n3270), .Z(n3272) );
  XOR U4159 ( .A(n3455), .B(n3456), .Z(n3270) );
  ANDN U4160 ( .B(n3457), .A(n3458), .Z(n3455) );
  AND U4161 ( .A(a[34]), .B(b[10]), .Z(n3454) );
  XNOR U4162 ( .A(n3459), .B(n3275), .Z(n3277) );
  XOR U4163 ( .A(n3460), .B(n3461), .Z(n3275) );
  ANDN U4164 ( .B(n3462), .A(n3463), .Z(n3460) );
  AND U4165 ( .A(b[9]), .B(a[35]), .Z(n3459) );
  XNOR U4166 ( .A(n3464), .B(n3280), .Z(n3282) );
  XOR U4167 ( .A(n3465), .B(n3466), .Z(n3280) );
  ANDN U4168 ( .B(n3467), .A(n3468), .Z(n3465) );
  AND U4169 ( .A(a[36]), .B(b[8]), .Z(n3464) );
  XNOR U4170 ( .A(n3469), .B(n3285), .Z(n3287) );
  XOR U4171 ( .A(n3470), .B(n3471), .Z(n3285) );
  ANDN U4172 ( .B(n3472), .A(n3473), .Z(n3470) );
  AND U4173 ( .A(b[7]), .B(a[37]), .Z(n3469) );
  XNOR U4174 ( .A(n3474), .B(n3290), .Z(n3292) );
  XOR U4175 ( .A(n3475), .B(n3476), .Z(n3290) );
  ANDN U4176 ( .B(n3477), .A(n3478), .Z(n3475) );
  AND U4177 ( .A(b[6]), .B(a[38]), .Z(n3474) );
  XNOR U4178 ( .A(n3479), .B(n3295), .Z(n3297) );
  XOR U4179 ( .A(n3480), .B(n3481), .Z(n3295) );
  ANDN U4180 ( .B(n3482), .A(n3483), .Z(n3480) );
  AND U4181 ( .A(b[5]), .B(a[39]), .Z(n3479) );
  XNOR U4182 ( .A(n3484), .B(n3300), .Z(n3302) );
  XOR U4183 ( .A(n3485), .B(n3486), .Z(n3300) );
  ANDN U4184 ( .B(n3487), .A(n3488), .Z(n3485) );
  AND U4185 ( .A(b[4]), .B(a[40]), .Z(n3484) );
  XNOR U4186 ( .A(n3489), .B(n3490), .Z(n3314) );
  NANDN U4187 ( .A(n3491), .B(n3492), .Z(n3490) );
  XNOR U4188 ( .A(n3493), .B(n3305), .Z(n3307) );
  XNOR U4189 ( .A(n3494), .B(n3495), .Z(n3305) );
  AND U4190 ( .A(n3496), .B(n3497), .Z(n3494) );
  AND U4191 ( .A(b[3]), .B(a[41]), .Z(n3493) );
  XNOR U4192 ( .A(n3498), .B(n3499), .Z(swire[43]) );
  XOR U4193 ( .A(n3325), .B(n3500), .Z(n3499) );
  XOR U4194 ( .A(n3324), .B(n3498), .Z(n3500) );
  NAND U4195 ( .A(a[43]), .B(b[0]), .Z(n3324) );
  XNOR U4196 ( .A(n3491), .B(n3492), .Z(n3325) );
  XOR U4197 ( .A(n3489), .B(n3501), .Z(n3492) );
  NAND U4198 ( .A(a[42]), .B(b[1]), .Z(n3501) );
  XOR U4199 ( .A(n3497), .B(n3502), .Z(n3491) );
  XOR U4200 ( .A(n3489), .B(n3496), .Z(n3502) );
  XNOR U4201 ( .A(n3503), .B(n3495), .Z(n3496) );
  AND U4202 ( .A(b[2]), .B(a[41]), .Z(n3503) );
  NANDN U4203 ( .A(n3504), .B(n3505), .Z(n3489) );
  XOR U4204 ( .A(n3495), .B(n3487), .Z(n3506) );
  XNOR U4205 ( .A(n3486), .B(n3482), .Z(n3507) );
  XNOR U4206 ( .A(n3481), .B(n3477), .Z(n3508) );
  XNOR U4207 ( .A(n3476), .B(n3472), .Z(n3509) );
  XNOR U4208 ( .A(n3471), .B(n3467), .Z(n3510) );
  XNOR U4209 ( .A(n3466), .B(n3462), .Z(n3511) );
  XNOR U4210 ( .A(n3461), .B(n3457), .Z(n3512) );
  XNOR U4211 ( .A(n3456), .B(n3452), .Z(n3513) );
  XNOR U4212 ( .A(n3451), .B(n3447), .Z(n3514) );
  XNOR U4213 ( .A(n3446), .B(n3442), .Z(n3515) );
  XNOR U4214 ( .A(n3441), .B(n3437), .Z(n3516) );
  XNOR U4215 ( .A(n3436), .B(n3432), .Z(n3517) );
  XNOR U4216 ( .A(n3431), .B(n3427), .Z(n3518) );
  XNOR U4217 ( .A(n3426), .B(n3422), .Z(n3519) );
  XNOR U4218 ( .A(n3421), .B(n3417), .Z(n3520) );
  XNOR U4219 ( .A(n3416), .B(n3412), .Z(n3521) );
  XNOR U4220 ( .A(n3411), .B(n3407), .Z(n3522) );
  XNOR U4221 ( .A(n3406), .B(n3402), .Z(n3523) );
  XNOR U4222 ( .A(n3401), .B(n3397), .Z(n3524) );
  XNOR U4223 ( .A(n3396), .B(n3392), .Z(n3525) );
  XNOR U4224 ( .A(n3391), .B(n3387), .Z(n3526) );
  XNOR U4225 ( .A(n3386), .B(n3382), .Z(n3527) );
  XNOR U4226 ( .A(n3381), .B(n3377), .Z(n3528) );
  XNOR U4227 ( .A(n3376), .B(n3372), .Z(n3529) );
  XNOR U4228 ( .A(n3371), .B(n3367), .Z(n3530) );
  XOR U4229 ( .A(n3366), .B(n3363), .Z(n3531) );
  XOR U4230 ( .A(n3532), .B(n3533), .Z(n3363) );
  XOR U4231 ( .A(n3361), .B(n3534), .Z(n3533) );
  XOR U4232 ( .A(n3535), .B(n3536), .Z(n3534) );
  XOR U4233 ( .A(n3537), .B(n3538), .Z(n3536) );
  NAND U4234 ( .A(a[13]), .B(b[30]), .Z(n3538) );
  AND U4235 ( .A(a[12]), .B(b[31]), .Z(n3537) );
  XOR U4236 ( .A(n3539), .B(n3535), .Z(n3532) );
  XOR U4237 ( .A(n3540), .B(n3541), .Z(n3535) );
  NOR U4238 ( .A(n3542), .B(n3543), .Z(n3540) );
  AND U4239 ( .A(a[14]), .B(b[29]), .Z(n3539) );
  XNOR U4240 ( .A(n3544), .B(n3361), .Z(n3362) );
  XOR U4241 ( .A(n3545), .B(n3546), .Z(n3361) );
  ANDN U4242 ( .B(n3547), .A(n3548), .Z(n3545) );
  AND U4243 ( .A(a[15]), .B(b[28]), .Z(n3544) );
  XNOR U4244 ( .A(n3549), .B(n3366), .Z(n3368) );
  XOR U4245 ( .A(n3550), .B(n3551), .Z(n3366) );
  ANDN U4246 ( .B(n3552), .A(n3553), .Z(n3550) );
  AND U4247 ( .A(a[16]), .B(b[27]), .Z(n3549) );
  XNOR U4248 ( .A(n3554), .B(n3371), .Z(n3373) );
  XOR U4249 ( .A(n3555), .B(n3556), .Z(n3371) );
  ANDN U4250 ( .B(n3557), .A(n3558), .Z(n3555) );
  AND U4251 ( .A(a[17]), .B(b[26]), .Z(n3554) );
  XNOR U4252 ( .A(n3559), .B(n3376), .Z(n3378) );
  XOR U4253 ( .A(n3560), .B(n3561), .Z(n3376) );
  ANDN U4254 ( .B(n3562), .A(n3563), .Z(n3560) );
  AND U4255 ( .A(a[18]), .B(b[25]), .Z(n3559) );
  XNOR U4256 ( .A(n3564), .B(n3381), .Z(n3383) );
  XOR U4257 ( .A(n3565), .B(n3566), .Z(n3381) );
  ANDN U4258 ( .B(n3567), .A(n3568), .Z(n3565) );
  AND U4259 ( .A(a[19]), .B(b[24]), .Z(n3564) );
  XNOR U4260 ( .A(n3569), .B(n3386), .Z(n3388) );
  XOR U4261 ( .A(n3570), .B(n3571), .Z(n3386) );
  ANDN U4262 ( .B(n3572), .A(n3573), .Z(n3570) );
  AND U4263 ( .A(a[20]), .B(b[23]), .Z(n3569) );
  XNOR U4264 ( .A(n3574), .B(n3391), .Z(n3393) );
  XOR U4265 ( .A(n3575), .B(n3576), .Z(n3391) );
  ANDN U4266 ( .B(n3577), .A(n3578), .Z(n3575) );
  AND U4267 ( .A(a[21]), .B(b[22]), .Z(n3574) );
  XNOR U4268 ( .A(n3579), .B(n3396), .Z(n3398) );
  XOR U4269 ( .A(n3580), .B(n3581), .Z(n3396) );
  ANDN U4270 ( .B(n3582), .A(n3583), .Z(n3580) );
  AND U4271 ( .A(a[22]), .B(b[21]), .Z(n3579) );
  XNOR U4272 ( .A(n3584), .B(n3401), .Z(n3403) );
  XOR U4273 ( .A(n3585), .B(n3586), .Z(n3401) );
  ANDN U4274 ( .B(n3587), .A(n3588), .Z(n3585) );
  AND U4275 ( .A(b[20]), .B(a[23]), .Z(n3584) );
  XNOR U4276 ( .A(n3589), .B(n3406), .Z(n3408) );
  XOR U4277 ( .A(n3590), .B(n3591), .Z(n3406) );
  ANDN U4278 ( .B(n3592), .A(n3593), .Z(n3590) );
  AND U4279 ( .A(a[24]), .B(b[19]), .Z(n3589) );
  XNOR U4280 ( .A(n3594), .B(n3411), .Z(n3413) );
  XOR U4281 ( .A(n3595), .B(n3596), .Z(n3411) );
  ANDN U4282 ( .B(n3597), .A(n3598), .Z(n3595) );
  AND U4283 ( .A(b[18]), .B(a[25]), .Z(n3594) );
  XNOR U4284 ( .A(n3599), .B(n3416), .Z(n3418) );
  XOR U4285 ( .A(n3600), .B(n3601), .Z(n3416) );
  ANDN U4286 ( .B(n3602), .A(n3603), .Z(n3600) );
  AND U4287 ( .A(a[26]), .B(b[17]), .Z(n3599) );
  XNOR U4288 ( .A(n3604), .B(n3421), .Z(n3423) );
  XOR U4289 ( .A(n3605), .B(n3606), .Z(n3421) );
  ANDN U4290 ( .B(n3607), .A(n3608), .Z(n3605) );
  AND U4291 ( .A(b[16]), .B(a[27]), .Z(n3604) );
  XNOR U4292 ( .A(n3609), .B(n3426), .Z(n3428) );
  XOR U4293 ( .A(n3610), .B(n3611), .Z(n3426) );
  ANDN U4294 ( .B(n3612), .A(n3613), .Z(n3610) );
  AND U4295 ( .A(a[28]), .B(b[15]), .Z(n3609) );
  XNOR U4296 ( .A(n3614), .B(n3431), .Z(n3433) );
  XOR U4297 ( .A(n3615), .B(n3616), .Z(n3431) );
  ANDN U4298 ( .B(n3617), .A(n3618), .Z(n3615) );
  AND U4299 ( .A(b[14]), .B(a[29]), .Z(n3614) );
  XNOR U4300 ( .A(n3619), .B(n3436), .Z(n3438) );
  XOR U4301 ( .A(n3620), .B(n3621), .Z(n3436) );
  ANDN U4302 ( .B(n3622), .A(n3623), .Z(n3620) );
  AND U4303 ( .A(a[30]), .B(b[13]), .Z(n3619) );
  XNOR U4304 ( .A(n3624), .B(n3441), .Z(n3443) );
  XOR U4305 ( .A(n3625), .B(n3626), .Z(n3441) );
  ANDN U4306 ( .B(n3627), .A(n3628), .Z(n3625) );
  AND U4307 ( .A(b[12]), .B(a[31]), .Z(n3624) );
  XNOR U4308 ( .A(n3629), .B(n3446), .Z(n3448) );
  XOR U4309 ( .A(n3630), .B(n3631), .Z(n3446) );
  ANDN U4310 ( .B(n3632), .A(n3633), .Z(n3630) );
  AND U4311 ( .A(a[32]), .B(b[11]), .Z(n3629) );
  XNOR U4312 ( .A(n3634), .B(n3451), .Z(n3453) );
  XOR U4313 ( .A(n3635), .B(n3636), .Z(n3451) );
  ANDN U4314 ( .B(n3637), .A(n3638), .Z(n3635) );
  AND U4315 ( .A(b[10]), .B(a[33]), .Z(n3634) );
  XNOR U4316 ( .A(n3639), .B(n3456), .Z(n3458) );
  XOR U4317 ( .A(n3640), .B(n3641), .Z(n3456) );
  ANDN U4318 ( .B(n3642), .A(n3643), .Z(n3640) );
  AND U4319 ( .A(a[34]), .B(b[9]), .Z(n3639) );
  XNOR U4320 ( .A(n3644), .B(n3461), .Z(n3463) );
  XOR U4321 ( .A(n3645), .B(n3646), .Z(n3461) );
  ANDN U4322 ( .B(n3647), .A(n3648), .Z(n3645) );
  AND U4323 ( .A(b[8]), .B(a[35]), .Z(n3644) );
  XNOR U4324 ( .A(n3649), .B(n3466), .Z(n3468) );
  XOR U4325 ( .A(n3650), .B(n3651), .Z(n3466) );
  ANDN U4326 ( .B(n3652), .A(n3653), .Z(n3650) );
  AND U4327 ( .A(a[36]), .B(b[7]), .Z(n3649) );
  XNOR U4328 ( .A(n3654), .B(n3471), .Z(n3473) );
  XOR U4329 ( .A(n3655), .B(n3656), .Z(n3471) );
  ANDN U4330 ( .B(n3657), .A(n3658), .Z(n3655) );
  AND U4331 ( .A(b[6]), .B(a[37]), .Z(n3654) );
  XNOR U4332 ( .A(n3659), .B(n3476), .Z(n3478) );
  XOR U4333 ( .A(n3660), .B(n3661), .Z(n3476) );
  ANDN U4334 ( .B(n3662), .A(n3663), .Z(n3660) );
  AND U4335 ( .A(b[5]), .B(a[38]), .Z(n3659) );
  XNOR U4336 ( .A(n3664), .B(n3481), .Z(n3483) );
  XOR U4337 ( .A(n3665), .B(n3666), .Z(n3481) );
  ANDN U4338 ( .B(n3667), .A(n3668), .Z(n3665) );
  AND U4339 ( .A(b[4]), .B(a[39]), .Z(n3664) );
  XNOR U4340 ( .A(n3669), .B(n3670), .Z(n3495) );
  NANDN U4341 ( .A(n3671), .B(n3672), .Z(n3670) );
  XNOR U4342 ( .A(n3673), .B(n3486), .Z(n3488) );
  XNOR U4343 ( .A(n3674), .B(n3675), .Z(n3486) );
  AND U4344 ( .A(n3676), .B(n3677), .Z(n3674) );
  AND U4345 ( .A(b[3]), .B(a[40]), .Z(n3673) );
  XNOR U4346 ( .A(n3678), .B(n3679), .Z(swire[42]) );
  XOR U4347 ( .A(n3505), .B(n3681), .Z(n3679) );
  XNOR U4348 ( .A(n3504), .B(n3680), .Z(n3681) );
  IV U4349 ( .A(n3678), .Z(n3680) );
  NAND U4350 ( .A(a[42]), .B(b[0]), .Z(n3504) );
  XNOR U4351 ( .A(n3671), .B(n3672), .Z(n3505) );
  XOR U4352 ( .A(n3669), .B(n3682), .Z(n3672) );
  NAND U4353 ( .A(b[1]), .B(a[41]), .Z(n3682) );
  XOR U4354 ( .A(n3677), .B(n3683), .Z(n3671) );
  XOR U4355 ( .A(n3669), .B(n3676), .Z(n3683) );
  XNOR U4356 ( .A(n3684), .B(n3675), .Z(n3676) );
  AND U4357 ( .A(b[2]), .B(a[40]), .Z(n3684) );
  NANDN U4358 ( .A(n3685), .B(n3686), .Z(n3669) );
  XOR U4359 ( .A(n3675), .B(n3667), .Z(n3687) );
  XNOR U4360 ( .A(n3666), .B(n3662), .Z(n3688) );
  XNOR U4361 ( .A(n3661), .B(n3657), .Z(n3689) );
  XNOR U4362 ( .A(n3656), .B(n3652), .Z(n3690) );
  XNOR U4363 ( .A(n3651), .B(n3647), .Z(n3691) );
  XNOR U4364 ( .A(n3646), .B(n3642), .Z(n3692) );
  XNOR U4365 ( .A(n3641), .B(n3637), .Z(n3693) );
  XNOR U4366 ( .A(n3636), .B(n3632), .Z(n3694) );
  XNOR U4367 ( .A(n3631), .B(n3627), .Z(n3695) );
  XNOR U4368 ( .A(n3626), .B(n3622), .Z(n3696) );
  XNOR U4369 ( .A(n3621), .B(n3617), .Z(n3697) );
  XNOR U4370 ( .A(n3616), .B(n3612), .Z(n3698) );
  XNOR U4371 ( .A(n3611), .B(n3607), .Z(n3699) );
  XNOR U4372 ( .A(n3606), .B(n3602), .Z(n3700) );
  XNOR U4373 ( .A(n3601), .B(n3597), .Z(n3701) );
  XNOR U4374 ( .A(n3596), .B(n3592), .Z(n3702) );
  XNOR U4375 ( .A(n3591), .B(n3587), .Z(n3703) );
  XNOR U4376 ( .A(n3586), .B(n3582), .Z(n3704) );
  XNOR U4377 ( .A(n3581), .B(n3577), .Z(n3705) );
  XNOR U4378 ( .A(n3576), .B(n3572), .Z(n3706) );
  XNOR U4379 ( .A(n3571), .B(n3567), .Z(n3707) );
  XNOR U4380 ( .A(n3566), .B(n3562), .Z(n3708) );
  XNOR U4381 ( .A(n3561), .B(n3557), .Z(n3709) );
  XNOR U4382 ( .A(n3556), .B(n3552), .Z(n3710) );
  XNOR U4383 ( .A(n3551), .B(n3547), .Z(n3711) );
  XOR U4384 ( .A(n3546), .B(n3543), .Z(n3712) );
  XOR U4385 ( .A(n3713), .B(n3714), .Z(n3543) );
  XOR U4386 ( .A(n3541), .B(n3715), .Z(n3714) );
  XOR U4387 ( .A(n3716), .B(n3717), .Z(n3715) );
  XOR U4388 ( .A(n3718), .B(n3719), .Z(n3717) );
  NAND U4389 ( .A(a[12]), .B(b[30]), .Z(n3719) );
  AND U4390 ( .A(a[11]), .B(b[31]), .Z(n3718) );
  XOR U4391 ( .A(n3720), .B(n3716), .Z(n3713) );
  XOR U4392 ( .A(n3721), .B(n3722), .Z(n3716) );
  NOR U4393 ( .A(n3723), .B(n3724), .Z(n3721) );
  AND U4394 ( .A(a[13]), .B(b[29]), .Z(n3720) );
  XNOR U4395 ( .A(n3725), .B(n3541), .Z(n3542) );
  XOR U4396 ( .A(n3726), .B(n3727), .Z(n3541) );
  ANDN U4397 ( .B(n3728), .A(n3729), .Z(n3726) );
  AND U4398 ( .A(a[14]), .B(b[28]), .Z(n3725) );
  XNOR U4399 ( .A(n3730), .B(n3546), .Z(n3548) );
  XOR U4400 ( .A(n3731), .B(n3732), .Z(n3546) );
  ANDN U4401 ( .B(n3733), .A(n3734), .Z(n3731) );
  AND U4402 ( .A(a[15]), .B(b[27]), .Z(n3730) );
  XNOR U4403 ( .A(n3735), .B(n3551), .Z(n3553) );
  XOR U4404 ( .A(n3736), .B(n3737), .Z(n3551) );
  ANDN U4405 ( .B(n3738), .A(n3739), .Z(n3736) );
  AND U4406 ( .A(a[16]), .B(b[26]), .Z(n3735) );
  XNOR U4407 ( .A(n3740), .B(n3556), .Z(n3558) );
  XOR U4408 ( .A(n3741), .B(n3742), .Z(n3556) );
  ANDN U4409 ( .B(n3743), .A(n3744), .Z(n3741) );
  AND U4410 ( .A(a[17]), .B(b[25]), .Z(n3740) );
  XNOR U4411 ( .A(n3745), .B(n3561), .Z(n3563) );
  XOR U4412 ( .A(n3746), .B(n3747), .Z(n3561) );
  ANDN U4413 ( .B(n3748), .A(n3749), .Z(n3746) );
  AND U4414 ( .A(a[18]), .B(b[24]), .Z(n3745) );
  XNOR U4415 ( .A(n3750), .B(n3566), .Z(n3568) );
  XOR U4416 ( .A(n3751), .B(n3752), .Z(n3566) );
  ANDN U4417 ( .B(n3753), .A(n3754), .Z(n3751) );
  AND U4418 ( .A(a[19]), .B(b[23]), .Z(n3750) );
  XNOR U4419 ( .A(n3755), .B(n3571), .Z(n3573) );
  XOR U4420 ( .A(n3756), .B(n3757), .Z(n3571) );
  ANDN U4421 ( .B(n3758), .A(n3759), .Z(n3756) );
  AND U4422 ( .A(a[20]), .B(b[22]), .Z(n3755) );
  XNOR U4423 ( .A(n3760), .B(n3576), .Z(n3578) );
  XOR U4424 ( .A(n3761), .B(n3762), .Z(n3576) );
  ANDN U4425 ( .B(n3763), .A(n3764), .Z(n3761) );
  AND U4426 ( .A(b[21]), .B(a[21]), .Z(n3760) );
  XNOR U4427 ( .A(n3765), .B(n3581), .Z(n3583) );
  XOR U4428 ( .A(n3766), .B(n3767), .Z(n3581) );
  ANDN U4429 ( .B(n3768), .A(n3769), .Z(n3766) );
  AND U4430 ( .A(a[22]), .B(b[20]), .Z(n3765) );
  XNOR U4431 ( .A(n3770), .B(n3586), .Z(n3588) );
  XOR U4432 ( .A(n3771), .B(n3772), .Z(n3586) );
  ANDN U4433 ( .B(n3773), .A(n3774), .Z(n3771) );
  AND U4434 ( .A(b[19]), .B(a[23]), .Z(n3770) );
  XNOR U4435 ( .A(n3775), .B(n3591), .Z(n3593) );
  XOR U4436 ( .A(n3776), .B(n3777), .Z(n3591) );
  ANDN U4437 ( .B(n3778), .A(n3779), .Z(n3776) );
  AND U4438 ( .A(a[24]), .B(b[18]), .Z(n3775) );
  XNOR U4439 ( .A(n3780), .B(n3596), .Z(n3598) );
  XOR U4440 ( .A(n3781), .B(n3782), .Z(n3596) );
  ANDN U4441 ( .B(n3783), .A(n3784), .Z(n3781) );
  AND U4442 ( .A(b[17]), .B(a[25]), .Z(n3780) );
  XNOR U4443 ( .A(n3785), .B(n3601), .Z(n3603) );
  XOR U4444 ( .A(n3786), .B(n3787), .Z(n3601) );
  ANDN U4445 ( .B(n3788), .A(n3789), .Z(n3786) );
  AND U4446 ( .A(a[26]), .B(b[16]), .Z(n3785) );
  XNOR U4447 ( .A(n3790), .B(n3606), .Z(n3608) );
  XOR U4448 ( .A(n3791), .B(n3792), .Z(n3606) );
  ANDN U4449 ( .B(n3793), .A(n3794), .Z(n3791) );
  AND U4450 ( .A(b[15]), .B(a[27]), .Z(n3790) );
  XNOR U4451 ( .A(n3795), .B(n3611), .Z(n3613) );
  XOR U4452 ( .A(n3796), .B(n3797), .Z(n3611) );
  ANDN U4453 ( .B(n3798), .A(n3799), .Z(n3796) );
  AND U4454 ( .A(a[28]), .B(b[14]), .Z(n3795) );
  XNOR U4455 ( .A(n3800), .B(n3616), .Z(n3618) );
  XOR U4456 ( .A(n3801), .B(n3802), .Z(n3616) );
  ANDN U4457 ( .B(n3803), .A(n3804), .Z(n3801) );
  AND U4458 ( .A(b[13]), .B(a[29]), .Z(n3800) );
  XNOR U4459 ( .A(n3805), .B(n3621), .Z(n3623) );
  XOR U4460 ( .A(n3806), .B(n3807), .Z(n3621) );
  ANDN U4461 ( .B(n3808), .A(n3809), .Z(n3806) );
  AND U4462 ( .A(a[30]), .B(b[12]), .Z(n3805) );
  XNOR U4463 ( .A(n3810), .B(n3626), .Z(n3628) );
  XOR U4464 ( .A(n3811), .B(n3812), .Z(n3626) );
  ANDN U4465 ( .B(n3813), .A(n3814), .Z(n3811) );
  AND U4466 ( .A(b[11]), .B(a[31]), .Z(n3810) );
  XNOR U4467 ( .A(n3815), .B(n3631), .Z(n3633) );
  XOR U4468 ( .A(n3816), .B(n3817), .Z(n3631) );
  ANDN U4469 ( .B(n3818), .A(n3819), .Z(n3816) );
  AND U4470 ( .A(a[32]), .B(b[10]), .Z(n3815) );
  XNOR U4471 ( .A(n3820), .B(n3636), .Z(n3638) );
  XOR U4472 ( .A(n3821), .B(n3822), .Z(n3636) );
  ANDN U4473 ( .B(n3823), .A(n3824), .Z(n3821) );
  AND U4474 ( .A(b[9]), .B(a[33]), .Z(n3820) );
  XNOR U4475 ( .A(n3825), .B(n3641), .Z(n3643) );
  XOR U4476 ( .A(n3826), .B(n3827), .Z(n3641) );
  ANDN U4477 ( .B(n3828), .A(n3829), .Z(n3826) );
  AND U4478 ( .A(a[34]), .B(b[8]), .Z(n3825) );
  XNOR U4479 ( .A(n3830), .B(n3646), .Z(n3648) );
  XOR U4480 ( .A(n3831), .B(n3832), .Z(n3646) );
  ANDN U4481 ( .B(n3833), .A(n3834), .Z(n3831) );
  AND U4482 ( .A(b[7]), .B(a[35]), .Z(n3830) );
  XNOR U4483 ( .A(n3835), .B(n3651), .Z(n3653) );
  XOR U4484 ( .A(n3836), .B(n3837), .Z(n3651) );
  ANDN U4485 ( .B(n3838), .A(n3839), .Z(n3836) );
  AND U4486 ( .A(b[6]), .B(a[36]), .Z(n3835) );
  XNOR U4487 ( .A(n3840), .B(n3656), .Z(n3658) );
  XOR U4488 ( .A(n3841), .B(n3842), .Z(n3656) );
  ANDN U4489 ( .B(n3843), .A(n3844), .Z(n3841) );
  AND U4490 ( .A(b[5]), .B(a[37]), .Z(n3840) );
  XNOR U4491 ( .A(n3845), .B(n3661), .Z(n3663) );
  XOR U4492 ( .A(n3846), .B(n3847), .Z(n3661) );
  ANDN U4493 ( .B(n3848), .A(n3849), .Z(n3846) );
  AND U4494 ( .A(b[4]), .B(a[38]), .Z(n3845) );
  XNOR U4495 ( .A(n3850), .B(n3851), .Z(n3675) );
  NANDN U4496 ( .A(n3852), .B(n3853), .Z(n3851) );
  XNOR U4497 ( .A(n3854), .B(n3666), .Z(n3668) );
  XNOR U4498 ( .A(n3855), .B(n3856), .Z(n3666) );
  AND U4499 ( .A(n3857), .B(n3858), .Z(n3855) );
  AND U4500 ( .A(b[3]), .B(a[39]), .Z(n3854) );
  XNOR U4501 ( .A(n3859), .B(n3860), .Z(swire[41]) );
  XOR U4502 ( .A(n3686), .B(n3861), .Z(n3860) );
  XOR U4503 ( .A(n3685), .B(n3859), .Z(n3861) );
  NAND U4504 ( .A(a[41]), .B(b[0]), .Z(n3685) );
  XNOR U4505 ( .A(n3852), .B(n3853), .Z(n3686) );
  XOR U4506 ( .A(n3850), .B(n3862), .Z(n3853) );
  NAND U4507 ( .A(a[40]), .B(b[1]), .Z(n3862) );
  XOR U4508 ( .A(n3858), .B(n3863), .Z(n3852) );
  XOR U4509 ( .A(n3850), .B(n3857), .Z(n3863) );
  XNOR U4510 ( .A(n3864), .B(n3856), .Z(n3857) );
  AND U4511 ( .A(b[2]), .B(a[39]), .Z(n3864) );
  NANDN U4512 ( .A(n3865), .B(n3866), .Z(n3850) );
  XOR U4513 ( .A(n3856), .B(n3848), .Z(n3867) );
  XNOR U4514 ( .A(n3847), .B(n3843), .Z(n3868) );
  XNOR U4515 ( .A(n3842), .B(n3838), .Z(n3869) );
  XNOR U4516 ( .A(n3837), .B(n3833), .Z(n3870) );
  XNOR U4517 ( .A(n3832), .B(n3828), .Z(n3871) );
  XNOR U4518 ( .A(n3827), .B(n3823), .Z(n3872) );
  XNOR U4519 ( .A(n3822), .B(n3818), .Z(n3873) );
  XNOR U4520 ( .A(n3817), .B(n3813), .Z(n3874) );
  XNOR U4521 ( .A(n3812), .B(n3808), .Z(n3875) );
  XNOR U4522 ( .A(n3807), .B(n3803), .Z(n3876) );
  XNOR U4523 ( .A(n3802), .B(n3798), .Z(n3877) );
  XNOR U4524 ( .A(n3797), .B(n3793), .Z(n3878) );
  XNOR U4525 ( .A(n3792), .B(n3788), .Z(n3879) );
  XNOR U4526 ( .A(n3787), .B(n3783), .Z(n3880) );
  XNOR U4527 ( .A(n3782), .B(n3778), .Z(n3881) );
  XNOR U4528 ( .A(n3777), .B(n3773), .Z(n3882) );
  XNOR U4529 ( .A(n3772), .B(n3768), .Z(n3883) );
  XNOR U4530 ( .A(n3767), .B(n3763), .Z(n3884) );
  XNOR U4531 ( .A(n3762), .B(n3758), .Z(n3885) );
  XNOR U4532 ( .A(n3757), .B(n3753), .Z(n3886) );
  XNOR U4533 ( .A(n3752), .B(n3748), .Z(n3887) );
  XNOR U4534 ( .A(n3747), .B(n3743), .Z(n3888) );
  XNOR U4535 ( .A(n3742), .B(n3738), .Z(n3889) );
  XNOR U4536 ( .A(n3737), .B(n3733), .Z(n3890) );
  XNOR U4537 ( .A(n3732), .B(n3728), .Z(n3891) );
  XOR U4538 ( .A(n3727), .B(n3724), .Z(n3892) );
  XOR U4539 ( .A(n3893), .B(n3894), .Z(n3724) );
  XOR U4540 ( .A(n3722), .B(n3895), .Z(n3894) );
  XOR U4541 ( .A(n3896), .B(n3897), .Z(n3895) );
  XOR U4542 ( .A(n3898), .B(n3899), .Z(n3897) );
  NAND U4543 ( .A(a[11]), .B(b[30]), .Z(n3899) );
  AND U4544 ( .A(a[10]), .B(b[31]), .Z(n3898) );
  XOR U4545 ( .A(n3900), .B(n3896), .Z(n3893) );
  XOR U4546 ( .A(n3901), .B(n3902), .Z(n3896) );
  NOR U4547 ( .A(n3903), .B(n3904), .Z(n3901) );
  AND U4548 ( .A(a[12]), .B(b[29]), .Z(n3900) );
  XNOR U4549 ( .A(n3905), .B(n3722), .Z(n3723) );
  XOR U4550 ( .A(n3906), .B(n3907), .Z(n3722) );
  ANDN U4551 ( .B(n3908), .A(n3909), .Z(n3906) );
  AND U4552 ( .A(a[13]), .B(b[28]), .Z(n3905) );
  XNOR U4553 ( .A(n3910), .B(n3727), .Z(n3729) );
  XOR U4554 ( .A(n3911), .B(n3912), .Z(n3727) );
  ANDN U4555 ( .B(n3913), .A(n3914), .Z(n3911) );
  AND U4556 ( .A(a[14]), .B(b[27]), .Z(n3910) );
  XNOR U4557 ( .A(n3915), .B(n3732), .Z(n3734) );
  XOR U4558 ( .A(n3916), .B(n3917), .Z(n3732) );
  ANDN U4559 ( .B(n3918), .A(n3919), .Z(n3916) );
  AND U4560 ( .A(a[15]), .B(b[26]), .Z(n3915) );
  XNOR U4561 ( .A(n3920), .B(n3737), .Z(n3739) );
  XOR U4562 ( .A(n3921), .B(n3922), .Z(n3737) );
  ANDN U4563 ( .B(n3923), .A(n3924), .Z(n3921) );
  AND U4564 ( .A(a[16]), .B(b[25]), .Z(n3920) );
  XNOR U4565 ( .A(n3925), .B(n3742), .Z(n3744) );
  XOR U4566 ( .A(n3926), .B(n3927), .Z(n3742) );
  ANDN U4567 ( .B(n3928), .A(n3929), .Z(n3926) );
  AND U4568 ( .A(a[17]), .B(b[24]), .Z(n3925) );
  XNOR U4569 ( .A(n3930), .B(n3747), .Z(n3749) );
  XOR U4570 ( .A(n3931), .B(n3932), .Z(n3747) );
  ANDN U4571 ( .B(n3933), .A(n3934), .Z(n3931) );
  AND U4572 ( .A(a[18]), .B(b[23]), .Z(n3930) );
  XNOR U4573 ( .A(n3935), .B(n3752), .Z(n3754) );
  XOR U4574 ( .A(n3936), .B(n3937), .Z(n3752) );
  ANDN U4575 ( .B(n3938), .A(n3939), .Z(n3936) );
  AND U4576 ( .A(a[19]), .B(b[22]), .Z(n3935) );
  XNOR U4577 ( .A(n3940), .B(n3757), .Z(n3759) );
  XOR U4578 ( .A(n3941), .B(n3942), .Z(n3757) );
  ANDN U4579 ( .B(n3943), .A(n3944), .Z(n3941) );
  AND U4580 ( .A(a[20]), .B(b[21]), .Z(n3940) );
  XNOR U4581 ( .A(n3945), .B(n3762), .Z(n3764) );
  XOR U4582 ( .A(n3946), .B(n3947), .Z(n3762) );
  ANDN U4583 ( .B(n3948), .A(n3949), .Z(n3946) );
  AND U4584 ( .A(b[20]), .B(a[21]), .Z(n3945) );
  XNOR U4585 ( .A(n3950), .B(n3767), .Z(n3769) );
  XOR U4586 ( .A(n3951), .B(n3952), .Z(n3767) );
  ANDN U4587 ( .B(n3953), .A(n3954), .Z(n3951) );
  AND U4588 ( .A(a[22]), .B(b[19]), .Z(n3950) );
  XNOR U4589 ( .A(n3955), .B(n3772), .Z(n3774) );
  XOR U4590 ( .A(n3956), .B(n3957), .Z(n3772) );
  ANDN U4591 ( .B(n3958), .A(n3959), .Z(n3956) );
  AND U4592 ( .A(b[18]), .B(a[23]), .Z(n3955) );
  XNOR U4593 ( .A(n3960), .B(n3777), .Z(n3779) );
  XOR U4594 ( .A(n3961), .B(n3962), .Z(n3777) );
  ANDN U4595 ( .B(n3963), .A(n3964), .Z(n3961) );
  AND U4596 ( .A(a[24]), .B(b[17]), .Z(n3960) );
  XNOR U4597 ( .A(n3965), .B(n3782), .Z(n3784) );
  XOR U4598 ( .A(n3966), .B(n3967), .Z(n3782) );
  ANDN U4599 ( .B(n3968), .A(n3969), .Z(n3966) );
  AND U4600 ( .A(b[16]), .B(a[25]), .Z(n3965) );
  XNOR U4601 ( .A(n3970), .B(n3787), .Z(n3789) );
  XOR U4602 ( .A(n3971), .B(n3972), .Z(n3787) );
  ANDN U4603 ( .B(n3973), .A(n3974), .Z(n3971) );
  AND U4604 ( .A(a[26]), .B(b[15]), .Z(n3970) );
  XNOR U4605 ( .A(n3975), .B(n3792), .Z(n3794) );
  XOR U4606 ( .A(n3976), .B(n3977), .Z(n3792) );
  ANDN U4607 ( .B(n3978), .A(n3979), .Z(n3976) );
  AND U4608 ( .A(b[14]), .B(a[27]), .Z(n3975) );
  XNOR U4609 ( .A(n3980), .B(n3797), .Z(n3799) );
  XOR U4610 ( .A(n3981), .B(n3982), .Z(n3797) );
  ANDN U4611 ( .B(n3983), .A(n3984), .Z(n3981) );
  AND U4612 ( .A(a[28]), .B(b[13]), .Z(n3980) );
  XNOR U4613 ( .A(n3985), .B(n3802), .Z(n3804) );
  XOR U4614 ( .A(n3986), .B(n3987), .Z(n3802) );
  ANDN U4615 ( .B(n3988), .A(n3989), .Z(n3986) );
  AND U4616 ( .A(b[12]), .B(a[29]), .Z(n3985) );
  XNOR U4617 ( .A(n3990), .B(n3807), .Z(n3809) );
  XOR U4618 ( .A(n3991), .B(n3992), .Z(n3807) );
  ANDN U4619 ( .B(n3993), .A(n3994), .Z(n3991) );
  AND U4620 ( .A(a[30]), .B(b[11]), .Z(n3990) );
  XNOR U4621 ( .A(n3995), .B(n3812), .Z(n3814) );
  XOR U4622 ( .A(n3996), .B(n3997), .Z(n3812) );
  ANDN U4623 ( .B(n3998), .A(n3999), .Z(n3996) );
  AND U4624 ( .A(b[10]), .B(a[31]), .Z(n3995) );
  XNOR U4625 ( .A(n4000), .B(n3817), .Z(n3819) );
  XOR U4626 ( .A(n4001), .B(n4002), .Z(n3817) );
  ANDN U4627 ( .B(n4003), .A(n4004), .Z(n4001) );
  AND U4628 ( .A(a[32]), .B(b[9]), .Z(n4000) );
  XNOR U4629 ( .A(n4005), .B(n3822), .Z(n3824) );
  XOR U4630 ( .A(n4006), .B(n4007), .Z(n3822) );
  ANDN U4631 ( .B(n4008), .A(n4009), .Z(n4006) );
  AND U4632 ( .A(b[8]), .B(a[33]), .Z(n4005) );
  XNOR U4633 ( .A(n4010), .B(n3827), .Z(n3829) );
  XOR U4634 ( .A(n4011), .B(n4012), .Z(n3827) );
  ANDN U4635 ( .B(n4013), .A(n4014), .Z(n4011) );
  AND U4636 ( .A(a[34]), .B(b[7]), .Z(n4010) );
  XNOR U4637 ( .A(n4015), .B(n3832), .Z(n3834) );
  XOR U4638 ( .A(n4016), .B(n4017), .Z(n3832) );
  ANDN U4639 ( .B(n4018), .A(n4019), .Z(n4016) );
  AND U4640 ( .A(b[6]), .B(a[35]), .Z(n4015) );
  XNOR U4641 ( .A(n4020), .B(n3837), .Z(n3839) );
  XOR U4642 ( .A(n4021), .B(n4022), .Z(n3837) );
  ANDN U4643 ( .B(n4023), .A(n4024), .Z(n4021) );
  AND U4644 ( .A(b[5]), .B(a[36]), .Z(n4020) );
  XNOR U4645 ( .A(n4025), .B(n3842), .Z(n3844) );
  XOR U4646 ( .A(n4026), .B(n4027), .Z(n3842) );
  ANDN U4647 ( .B(n4028), .A(n4029), .Z(n4026) );
  AND U4648 ( .A(b[4]), .B(a[37]), .Z(n4025) );
  XNOR U4649 ( .A(n4030), .B(n4031), .Z(n3856) );
  NANDN U4650 ( .A(n4032), .B(n4033), .Z(n4031) );
  XNOR U4651 ( .A(n4034), .B(n3847), .Z(n3849) );
  XNOR U4652 ( .A(n4035), .B(n4036), .Z(n3847) );
  AND U4653 ( .A(n4037), .B(n4038), .Z(n4035) );
  AND U4654 ( .A(b[3]), .B(a[38]), .Z(n4034) );
  XNOR U4655 ( .A(n4039), .B(n4040), .Z(swire[40]) );
  XOR U4656 ( .A(n3866), .B(n4042), .Z(n4040) );
  XNOR U4657 ( .A(n3865), .B(n4041), .Z(n4042) );
  IV U4658 ( .A(n4039), .Z(n4041) );
  NAND U4659 ( .A(a[40]), .B(b[0]), .Z(n3865) );
  XNOR U4660 ( .A(n4032), .B(n4033), .Z(n3866) );
  XOR U4661 ( .A(n4030), .B(n4043), .Z(n4033) );
  NAND U4662 ( .A(b[1]), .B(a[39]), .Z(n4043) );
  XOR U4663 ( .A(n4038), .B(n4044), .Z(n4032) );
  XOR U4664 ( .A(n4030), .B(n4037), .Z(n4044) );
  XNOR U4665 ( .A(n4045), .B(n4036), .Z(n4037) );
  AND U4666 ( .A(b[2]), .B(a[38]), .Z(n4045) );
  NANDN U4667 ( .A(n4046), .B(n4047), .Z(n4030) );
  XOR U4668 ( .A(n4036), .B(n4028), .Z(n4048) );
  XNOR U4669 ( .A(n4027), .B(n4023), .Z(n4049) );
  XNOR U4670 ( .A(n4022), .B(n4018), .Z(n4050) );
  XNOR U4671 ( .A(n4017), .B(n4013), .Z(n4051) );
  XNOR U4672 ( .A(n4012), .B(n4008), .Z(n4052) );
  XNOR U4673 ( .A(n4007), .B(n4003), .Z(n4053) );
  XNOR U4674 ( .A(n4002), .B(n3998), .Z(n4054) );
  XNOR U4675 ( .A(n3997), .B(n3993), .Z(n4055) );
  XNOR U4676 ( .A(n3992), .B(n3988), .Z(n4056) );
  XNOR U4677 ( .A(n3987), .B(n3983), .Z(n4057) );
  XNOR U4678 ( .A(n3982), .B(n3978), .Z(n4058) );
  XNOR U4679 ( .A(n3977), .B(n3973), .Z(n4059) );
  XNOR U4680 ( .A(n3972), .B(n3968), .Z(n4060) );
  XNOR U4681 ( .A(n3967), .B(n3963), .Z(n4061) );
  XNOR U4682 ( .A(n3962), .B(n3958), .Z(n4062) );
  XNOR U4683 ( .A(n3957), .B(n3953), .Z(n4063) );
  XNOR U4684 ( .A(n3952), .B(n3948), .Z(n4064) );
  XNOR U4685 ( .A(n3947), .B(n3943), .Z(n4065) );
  XNOR U4686 ( .A(n3942), .B(n3938), .Z(n4066) );
  XNOR U4687 ( .A(n3937), .B(n3933), .Z(n4067) );
  XNOR U4688 ( .A(n3932), .B(n3928), .Z(n4068) );
  XNOR U4689 ( .A(n3927), .B(n3923), .Z(n4069) );
  XNOR U4690 ( .A(n3922), .B(n3918), .Z(n4070) );
  XNOR U4691 ( .A(n3917), .B(n3913), .Z(n4071) );
  XNOR U4692 ( .A(n3912), .B(n3908), .Z(n4072) );
  XOR U4693 ( .A(n3907), .B(n3904), .Z(n4073) );
  XOR U4694 ( .A(n4074), .B(n4075), .Z(n3904) );
  XOR U4695 ( .A(n3902), .B(n4076), .Z(n4075) );
  XOR U4696 ( .A(n4077), .B(n4078), .Z(n4076) );
  XOR U4697 ( .A(n4079), .B(n4080), .Z(n4078) );
  NAND U4698 ( .A(a[10]), .B(b[30]), .Z(n4080) );
  AND U4699 ( .A(a[9]), .B(b[31]), .Z(n4079) );
  XOR U4700 ( .A(n4081), .B(n4077), .Z(n4074) );
  XOR U4701 ( .A(n4082), .B(n4083), .Z(n4077) );
  NOR U4702 ( .A(n4084), .B(n4085), .Z(n4082) );
  AND U4703 ( .A(a[11]), .B(b[29]), .Z(n4081) );
  XNOR U4704 ( .A(n4086), .B(n3902), .Z(n3903) );
  XOR U4705 ( .A(n4087), .B(n4088), .Z(n3902) );
  ANDN U4706 ( .B(n4089), .A(n4090), .Z(n4087) );
  AND U4707 ( .A(a[12]), .B(b[28]), .Z(n4086) );
  XNOR U4708 ( .A(n4091), .B(n3907), .Z(n3909) );
  XOR U4709 ( .A(n4092), .B(n4093), .Z(n3907) );
  ANDN U4710 ( .B(n4094), .A(n4095), .Z(n4092) );
  AND U4711 ( .A(a[13]), .B(b[27]), .Z(n4091) );
  XNOR U4712 ( .A(n4096), .B(n3912), .Z(n3914) );
  XOR U4713 ( .A(n4097), .B(n4098), .Z(n3912) );
  ANDN U4714 ( .B(n4099), .A(n4100), .Z(n4097) );
  AND U4715 ( .A(a[14]), .B(b[26]), .Z(n4096) );
  XNOR U4716 ( .A(n4101), .B(n3917), .Z(n3919) );
  XOR U4717 ( .A(n4102), .B(n4103), .Z(n3917) );
  ANDN U4718 ( .B(n4104), .A(n4105), .Z(n4102) );
  AND U4719 ( .A(a[15]), .B(b[25]), .Z(n4101) );
  XNOR U4720 ( .A(n4106), .B(n3922), .Z(n3924) );
  XOR U4721 ( .A(n4107), .B(n4108), .Z(n3922) );
  ANDN U4722 ( .B(n4109), .A(n4110), .Z(n4107) );
  AND U4723 ( .A(a[16]), .B(b[24]), .Z(n4106) );
  XNOR U4724 ( .A(n4111), .B(n3927), .Z(n3929) );
  XOR U4725 ( .A(n4112), .B(n4113), .Z(n3927) );
  ANDN U4726 ( .B(n4114), .A(n4115), .Z(n4112) );
  AND U4727 ( .A(a[17]), .B(b[23]), .Z(n4111) );
  XNOR U4728 ( .A(n4116), .B(n3932), .Z(n3934) );
  XOR U4729 ( .A(n4117), .B(n4118), .Z(n3932) );
  ANDN U4730 ( .B(n4119), .A(n4120), .Z(n4117) );
  AND U4731 ( .A(a[18]), .B(b[22]), .Z(n4116) );
  XNOR U4732 ( .A(n4121), .B(n3937), .Z(n3939) );
  XOR U4733 ( .A(n4122), .B(n4123), .Z(n3937) );
  ANDN U4734 ( .B(n4124), .A(n4125), .Z(n4122) );
  AND U4735 ( .A(a[19]), .B(b[21]), .Z(n4121) );
  XNOR U4736 ( .A(n4126), .B(n3942), .Z(n3944) );
  XOR U4737 ( .A(n4127), .B(n4128), .Z(n3942) );
  ANDN U4738 ( .B(n4129), .A(n4130), .Z(n4127) );
  AND U4739 ( .A(a[20]), .B(b[20]), .Z(n4126) );
  XNOR U4740 ( .A(n4131), .B(n3947), .Z(n3949) );
  XOR U4741 ( .A(n4132), .B(n4133), .Z(n3947) );
  ANDN U4742 ( .B(n4134), .A(n4135), .Z(n4132) );
  AND U4743 ( .A(b[19]), .B(a[21]), .Z(n4131) );
  XNOR U4744 ( .A(n4136), .B(n3952), .Z(n3954) );
  XOR U4745 ( .A(n4137), .B(n4138), .Z(n3952) );
  ANDN U4746 ( .B(n4139), .A(n4140), .Z(n4137) );
  AND U4747 ( .A(a[22]), .B(b[18]), .Z(n4136) );
  XNOR U4748 ( .A(n4141), .B(n3957), .Z(n3959) );
  XOR U4749 ( .A(n4142), .B(n4143), .Z(n3957) );
  ANDN U4750 ( .B(n4144), .A(n4145), .Z(n4142) );
  AND U4751 ( .A(b[17]), .B(a[23]), .Z(n4141) );
  XNOR U4752 ( .A(n4146), .B(n3962), .Z(n3964) );
  XOR U4753 ( .A(n4147), .B(n4148), .Z(n3962) );
  ANDN U4754 ( .B(n4149), .A(n4150), .Z(n4147) );
  AND U4755 ( .A(a[24]), .B(b[16]), .Z(n4146) );
  XNOR U4756 ( .A(n4151), .B(n3967), .Z(n3969) );
  XOR U4757 ( .A(n4152), .B(n4153), .Z(n3967) );
  ANDN U4758 ( .B(n4154), .A(n4155), .Z(n4152) );
  AND U4759 ( .A(b[15]), .B(a[25]), .Z(n4151) );
  XNOR U4760 ( .A(n4156), .B(n3972), .Z(n3974) );
  XOR U4761 ( .A(n4157), .B(n4158), .Z(n3972) );
  ANDN U4762 ( .B(n4159), .A(n4160), .Z(n4157) );
  AND U4763 ( .A(a[26]), .B(b[14]), .Z(n4156) );
  XNOR U4764 ( .A(n4161), .B(n3977), .Z(n3979) );
  XOR U4765 ( .A(n4162), .B(n4163), .Z(n3977) );
  ANDN U4766 ( .B(n4164), .A(n4165), .Z(n4162) );
  AND U4767 ( .A(b[13]), .B(a[27]), .Z(n4161) );
  XNOR U4768 ( .A(n4166), .B(n3982), .Z(n3984) );
  XOR U4769 ( .A(n4167), .B(n4168), .Z(n3982) );
  ANDN U4770 ( .B(n4169), .A(n4170), .Z(n4167) );
  AND U4771 ( .A(a[28]), .B(b[12]), .Z(n4166) );
  XNOR U4772 ( .A(n4171), .B(n3987), .Z(n3989) );
  XOR U4773 ( .A(n4172), .B(n4173), .Z(n3987) );
  ANDN U4774 ( .B(n4174), .A(n4175), .Z(n4172) );
  AND U4775 ( .A(b[11]), .B(a[29]), .Z(n4171) );
  XNOR U4776 ( .A(n4176), .B(n3992), .Z(n3994) );
  XOR U4777 ( .A(n4177), .B(n4178), .Z(n3992) );
  ANDN U4778 ( .B(n4179), .A(n4180), .Z(n4177) );
  AND U4779 ( .A(a[30]), .B(b[10]), .Z(n4176) );
  XNOR U4780 ( .A(n4181), .B(n3997), .Z(n3999) );
  XOR U4781 ( .A(n4182), .B(n4183), .Z(n3997) );
  ANDN U4782 ( .B(n4184), .A(n4185), .Z(n4182) );
  AND U4783 ( .A(b[9]), .B(a[31]), .Z(n4181) );
  XNOR U4784 ( .A(n4186), .B(n4002), .Z(n4004) );
  XOR U4785 ( .A(n4187), .B(n4188), .Z(n4002) );
  ANDN U4786 ( .B(n4189), .A(n4190), .Z(n4187) );
  AND U4787 ( .A(a[32]), .B(b[8]), .Z(n4186) );
  XNOR U4788 ( .A(n4191), .B(n4007), .Z(n4009) );
  XOR U4789 ( .A(n4192), .B(n4193), .Z(n4007) );
  ANDN U4790 ( .B(n4194), .A(n4195), .Z(n4192) );
  AND U4791 ( .A(b[7]), .B(a[33]), .Z(n4191) );
  XNOR U4792 ( .A(n4196), .B(n4012), .Z(n4014) );
  XOR U4793 ( .A(n4197), .B(n4198), .Z(n4012) );
  ANDN U4794 ( .B(n4199), .A(n4200), .Z(n4197) );
  AND U4795 ( .A(b[6]), .B(a[34]), .Z(n4196) );
  XNOR U4796 ( .A(n4201), .B(n4017), .Z(n4019) );
  XOR U4797 ( .A(n4202), .B(n4203), .Z(n4017) );
  ANDN U4798 ( .B(n4204), .A(n4205), .Z(n4202) );
  AND U4799 ( .A(b[5]), .B(a[35]), .Z(n4201) );
  XNOR U4800 ( .A(n4206), .B(n4022), .Z(n4024) );
  XOR U4801 ( .A(n4207), .B(n4208), .Z(n4022) );
  ANDN U4802 ( .B(n4209), .A(n4210), .Z(n4207) );
  AND U4803 ( .A(b[4]), .B(a[36]), .Z(n4206) );
  XNOR U4804 ( .A(n4211), .B(n4212), .Z(n4036) );
  NANDN U4805 ( .A(n4213), .B(n4214), .Z(n4212) );
  XNOR U4806 ( .A(n4215), .B(n4027), .Z(n4029) );
  XNOR U4807 ( .A(n4216), .B(n4217), .Z(n4027) );
  AND U4808 ( .A(n4218), .B(n4219), .Z(n4216) );
  AND U4809 ( .A(b[3]), .B(a[37]), .Z(n4215) );
  XNOR U4810 ( .A(n4220), .B(n4221), .Z(swire[39]) );
  XOR U4811 ( .A(n4047), .B(n4222), .Z(n4221) );
  XOR U4812 ( .A(n4046), .B(n4220), .Z(n4222) );
  NAND U4813 ( .A(a[39]), .B(b[0]), .Z(n4046) );
  XNOR U4814 ( .A(n4213), .B(n4214), .Z(n4047) );
  XOR U4815 ( .A(n4211), .B(n4223), .Z(n4214) );
  NAND U4816 ( .A(a[38]), .B(b[1]), .Z(n4223) );
  XOR U4817 ( .A(n4219), .B(n4224), .Z(n4213) );
  XOR U4818 ( .A(n4211), .B(n4218), .Z(n4224) );
  XNOR U4819 ( .A(n4225), .B(n4217), .Z(n4218) );
  AND U4820 ( .A(b[2]), .B(a[37]), .Z(n4225) );
  NANDN U4821 ( .A(n4226), .B(n4227), .Z(n4211) );
  XOR U4822 ( .A(n4217), .B(n4209), .Z(n4228) );
  XNOR U4823 ( .A(n4208), .B(n4204), .Z(n4229) );
  XNOR U4824 ( .A(n4203), .B(n4199), .Z(n4230) );
  XNOR U4825 ( .A(n4198), .B(n4194), .Z(n4231) );
  XNOR U4826 ( .A(n4193), .B(n4189), .Z(n4232) );
  XNOR U4827 ( .A(n4188), .B(n4184), .Z(n4233) );
  XNOR U4828 ( .A(n4183), .B(n4179), .Z(n4234) );
  XNOR U4829 ( .A(n4178), .B(n4174), .Z(n4235) );
  XNOR U4830 ( .A(n4173), .B(n4169), .Z(n4236) );
  XNOR U4831 ( .A(n4168), .B(n4164), .Z(n4237) );
  XNOR U4832 ( .A(n4163), .B(n4159), .Z(n4238) );
  XNOR U4833 ( .A(n4158), .B(n4154), .Z(n4239) );
  XNOR U4834 ( .A(n4153), .B(n4149), .Z(n4240) );
  XNOR U4835 ( .A(n4148), .B(n4144), .Z(n4241) );
  XNOR U4836 ( .A(n4143), .B(n4139), .Z(n4242) );
  XNOR U4837 ( .A(n4138), .B(n4134), .Z(n4243) );
  XNOR U4838 ( .A(n4133), .B(n4129), .Z(n4244) );
  XNOR U4839 ( .A(n4128), .B(n4124), .Z(n4245) );
  XNOR U4840 ( .A(n4123), .B(n4119), .Z(n4246) );
  XNOR U4841 ( .A(n4118), .B(n4114), .Z(n4247) );
  XNOR U4842 ( .A(n4113), .B(n4109), .Z(n4248) );
  XNOR U4843 ( .A(n4108), .B(n4104), .Z(n4249) );
  XNOR U4844 ( .A(n4103), .B(n4099), .Z(n4250) );
  XNOR U4845 ( .A(n4098), .B(n4094), .Z(n4251) );
  XNOR U4846 ( .A(n4093), .B(n4089), .Z(n4252) );
  XOR U4847 ( .A(n4088), .B(n4085), .Z(n4253) );
  XOR U4848 ( .A(n4254), .B(n4255), .Z(n4085) );
  XOR U4849 ( .A(n4083), .B(n4256), .Z(n4255) );
  XOR U4850 ( .A(n4257), .B(n4258), .Z(n4256) );
  XOR U4851 ( .A(n4259), .B(n4260), .Z(n4258) );
  NAND U4852 ( .A(a[9]), .B(b[30]), .Z(n4260) );
  AND U4853 ( .A(a[8]), .B(b[31]), .Z(n4259) );
  XOR U4854 ( .A(n4261), .B(n4257), .Z(n4254) );
  XOR U4855 ( .A(n4262), .B(n4263), .Z(n4257) );
  NOR U4856 ( .A(n4264), .B(n4265), .Z(n4262) );
  AND U4857 ( .A(a[10]), .B(b[29]), .Z(n4261) );
  XNOR U4858 ( .A(n4266), .B(n4083), .Z(n4084) );
  XOR U4859 ( .A(n4267), .B(n4268), .Z(n4083) );
  ANDN U4860 ( .B(n4269), .A(n4270), .Z(n4267) );
  AND U4861 ( .A(a[11]), .B(b[28]), .Z(n4266) );
  XNOR U4862 ( .A(n4271), .B(n4088), .Z(n4090) );
  XOR U4863 ( .A(n4272), .B(n4273), .Z(n4088) );
  ANDN U4864 ( .B(n4274), .A(n4275), .Z(n4272) );
  AND U4865 ( .A(a[12]), .B(b[27]), .Z(n4271) );
  XNOR U4866 ( .A(n4276), .B(n4093), .Z(n4095) );
  XOR U4867 ( .A(n4277), .B(n4278), .Z(n4093) );
  ANDN U4868 ( .B(n4279), .A(n4280), .Z(n4277) );
  AND U4869 ( .A(a[13]), .B(b[26]), .Z(n4276) );
  XNOR U4870 ( .A(n4281), .B(n4098), .Z(n4100) );
  XOR U4871 ( .A(n4282), .B(n4283), .Z(n4098) );
  ANDN U4872 ( .B(n4284), .A(n4285), .Z(n4282) );
  AND U4873 ( .A(a[14]), .B(b[25]), .Z(n4281) );
  XNOR U4874 ( .A(n4286), .B(n4103), .Z(n4105) );
  XOR U4875 ( .A(n4287), .B(n4288), .Z(n4103) );
  ANDN U4876 ( .B(n4289), .A(n4290), .Z(n4287) );
  AND U4877 ( .A(a[15]), .B(b[24]), .Z(n4286) );
  XNOR U4878 ( .A(n4291), .B(n4108), .Z(n4110) );
  XOR U4879 ( .A(n4292), .B(n4293), .Z(n4108) );
  ANDN U4880 ( .B(n4294), .A(n4295), .Z(n4292) );
  AND U4881 ( .A(a[16]), .B(b[23]), .Z(n4291) );
  XNOR U4882 ( .A(n4296), .B(n4113), .Z(n4115) );
  XOR U4883 ( .A(n4297), .B(n4298), .Z(n4113) );
  ANDN U4884 ( .B(n4299), .A(n4300), .Z(n4297) );
  AND U4885 ( .A(a[17]), .B(b[22]), .Z(n4296) );
  XNOR U4886 ( .A(n4301), .B(n4118), .Z(n4120) );
  XOR U4887 ( .A(n4302), .B(n4303), .Z(n4118) );
  ANDN U4888 ( .B(n4304), .A(n4305), .Z(n4302) );
  AND U4889 ( .A(a[18]), .B(b[21]), .Z(n4301) );
  XNOR U4890 ( .A(n4306), .B(n4123), .Z(n4125) );
  XOR U4891 ( .A(n4307), .B(n4308), .Z(n4123) );
  ANDN U4892 ( .B(n4309), .A(n4310), .Z(n4307) );
  AND U4893 ( .A(a[19]), .B(b[20]), .Z(n4306) );
  XNOR U4894 ( .A(n4311), .B(n4128), .Z(n4130) );
  XOR U4895 ( .A(n4312), .B(n4313), .Z(n4128) );
  ANDN U4896 ( .B(n4314), .A(n4315), .Z(n4312) );
  AND U4897 ( .A(a[20]), .B(b[19]), .Z(n4311) );
  XNOR U4898 ( .A(n4316), .B(n4133), .Z(n4135) );
  XOR U4899 ( .A(n4317), .B(n4318), .Z(n4133) );
  ANDN U4900 ( .B(n4319), .A(n4320), .Z(n4317) );
  AND U4901 ( .A(b[18]), .B(a[21]), .Z(n4316) );
  XNOR U4902 ( .A(n4321), .B(n4138), .Z(n4140) );
  XOR U4903 ( .A(n4322), .B(n4323), .Z(n4138) );
  ANDN U4904 ( .B(n4324), .A(n4325), .Z(n4322) );
  AND U4905 ( .A(a[22]), .B(b[17]), .Z(n4321) );
  XNOR U4906 ( .A(n4326), .B(n4143), .Z(n4145) );
  XOR U4907 ( .A(n4327), .B(n4328), .Z(n4143) );
  ANDN U4908 ( .B(n4329), .A(n4330), .Z(n4327) );
  AND U4909 ( .A(b[16]), .B(a[23]), .Z(n4326) );
  XNOR U4910 ( .A(n4331), .B(n4148), .Z(n4150) );
  XOR U4911 ( .A(n4332), .B(n4333), .Z(n4148) );
  ANDN U4912 ( .B(n4334), .A(n4335), .Z(n4332) );
  AND U4913 ( .A(a[24]), .B(b[15]), .Z(n4331) );
  XNOR U4914 ( .A(n4336), .B(n4153), .Z(n4155) );
  XOR U4915 ( .A(n4337), .B(n4338), .Z(n4153) );
  ANDN U4916 ( .B(n4339), .A(n4340), .Z(n4337) );
  AND U4917 ( .A(b[14]), .B(a[25]), .Z(n4336) );
  XNOR U4918 ( .A(n4341), .B(n4158), .Z(n4160) );
  XOR U4919 ( .A(n4342), .B(n4343), .Z(n4158) );
  ANDN U4920 ( .B(n4344), .A(n4345), .Z(n4342) );
  AND U4921 ( .A(a[26]), .B(b[13]), .Z(n4341) );
  XNOR U4922 ( .A(n4346), .B(n4163), .Z(n4165) );
  XOR U4923 ( .A(n4347), .B(n4348), .Z(n4163) );
  ANDN U4924 ( .B(n4349), .A(n4350), .Z(n4347) );
  AND U4925 ( .A(b[12]), .B(a[27]), .Z(n4346) );
  XNOR U4926 ( .A(n4351), .B(n4168), .Z(n4170) );
  XOR U4927 ( .A(n4352), .B(n4353), .Z(n4168) );
  ANDN U4928 ( .B(n4354), .A(n4355), .Z(n4352) );
  AND U4929 ( .A(a[28]), .B(b[11]), .Z(n4351) );
  XNOR U4930 ( .A(n4356), .B(n4173), .Z(n4175) );
  XOR U4931 ( .A(n4357), .B(n4358), .Z(n4173) );
  ANDN U4932 ( .B(n4359), .A(n4360), .Z(n4357) );
  AND U4933 ( .A(b[10]), .B(a[29]), .Z(n4356) );
  XNOR U4934 ( .A(n4361), .B(n4178), .Z(n4180) );
  XOR U4935 ( .A(n4362), .B(n4363), .Z(n4178) );
  ANDN U4936 ( .B(n4364), .A(n4365), .Z(n4362) );
  AND U4937 ( .A(a[30]), .B(b[9]), .Z(n4361) );
  XNOR U4938 ( .A(n4366), .B(n4183), .Z(n4185) );
  XOR U4939 ( .A(n4367), .B(n4368), .Z(n4183) );
  ANDN U4940 ( .B(n4369), .A(n4370), .Z(n4367) );
  AND U4941 ( .A(b[8]), .B(a[31]), .Z(n4366) );
  XNOR U4942 ( .A(n4371), .B(n4188), .Z(n4190) );
  XOR U4943 ( .A(n4372), .B(n4373), .Z(n4188) );
  ANDN U4944 ( .B(n4374), .A(n4375), .Z(n4372) );
  AND U4945 ( .A(a[32]), .B(b[7]), .Z(n4371) );
  XNOR U4946 ( .A(n4376), .B(n4193), .Z(n4195) );
  XOR U4947 ( .A(n4377), .B(n4378), .Z(n4193) );
  ANDN U4948 ( .B(n4379), .A(n4380), .Z(n4377) );
  AND U4949 ( .A(b[6]), .B(a[33]), .Z(n4376) );
  XNOR U4950 ( .A(n4381), .B(n4198), .Z(n4200) );
  XOR U4951 ( .A(n4382), .B(n4383), .Z(n4198) );
  ANDN U4952 ( .B(n4384), .A(n4385), .Z(n4382) );
  AND U4953 ( .A(b[5]), .B(a[34]), .Z(n4381) );
  XNOR U4954 ( .A(n4386), .B(n4203), .Z(n4205) );
  XOR U4955 ( .A(n4387), .B(n4388), .Z(n4203) );
  ANDN U4956 ( .B(n4389), .A(n4390), .Z(n4387) );
  AND U4957 ( .A(b[4]), .B(a[35]), .Z(n4386) );
  XNOR U4958 ( .A(n4391), .B(n4392), .Z(n4217) );
  NANDN U4959 ( .A(n4393), .B(n4394), .Z(n4392) );
  XNOR U4960 ( .A(n4395), .B(n4208), .Z(n4210) );
  XNOR U4961 ( .A(n4396), .B(n4397), .Z(n4208) );
  AND U4962 ( .A(n4398), .B(n4399), .Z(n4396) );
  AND U4963 ( .A(b[3]), .B(a[36]), .Z(n4395) );
  XNOR U4964 ( .A(n4400), .B(n4401), .Z(swire[38]) );
  XOR U4965 ( .A(n4227), .B(n4403), .Z(n4401) );
  XNOR U4966 ( .A(n4226), .B(n4402), .Z(n4403) );
  IV U4967 ( .A(n4400), .Z(n4402) );
  NAND U4968 ( .A(a[38]), .B(b[0]), .Z(n4226) );
  XNOR U4969 ( .A(n4393), .B(n4394), .Z(n4227) );
  XOR U4970 ( .A(n4391), .B(n4404), .Z(n4394) );
  NAND U4971 ( .A(b[1]), .B(a[37]), .Z(n4404) );
  XOR U4972 ( .A(n4399), .B(n4405), .Z(n4393) );
  XOR U4973 ( .A(n4391), .B(n4398), .Z(n4405) );
  XNOR U4974 ( .A(n4406), .B(n4397), .Z(n4398) );
  AND U4975 ( .A(b[2]), .B(a[36]), .Z(n4406) );
  NANDN U4976 ( .A(n4407), .B(n4408), .Z(n4391) );
  XOR U4977 ( .A(n4397), .B(n4389), .Z(n4409) );
  XNOR U4978 ( .A(n4388), .B(n4384), .Z(n4410) );
  XNOR U4979 ( .A(n4383), .B(n4379), .Z(n4411) );
  XNOR U4980 ( .A(n4378), .B(n4374), .Z(n4412) );
  XNOR U4981 ( .A(n4373), .B(n4369), .Z(n4413) );
  XNOR U4982 ( .A(n4368), .B(n4364), .Z(n4414) );
  XNOR U4983 ( .A(n4363), .B(n4359), .Z(n4415) );
  XNOR U4984 ( .A(n4358), .B(n4354), .Z(n4416) );
  XNOR U4985 ( .A(n4353), .B(n4349), .Z(n4417) );
  XNOR U4986 ( .A(n4348), .B(n4344), .Z(n4418) );
  XNOR U4987 ( .A(n4343), .B(n4339), .Z(n4419) );
  XNOR U4988 ( .A(n4338), .B(n4334), .Z(n4420) );
  XNOR U4989 ( .A(n4333), .B(n4329), .Z(n4421) );
  XNOR U4990 ( .A(n4328), .B(n4324), .Z(n4422) );
  XNOR U4991 ( .A(n4323), .B(n4319), .Z(n4423) );
  XNOR U4992 ( .A(n4318), .B(n4314), .Z(n4424) );
  XNOR U4993 ( .A(n4313), .B(n4309), .Z(n4425) );
  XNOR U4994 ( .A(n4308), .B(n4304), .Z(n4426) );
  XNOR U4995 ( .A(n4303), .B(n4299), .Z(n4427) );
  XNOR U4996 ( .A(n4298), .B(n4294), .Z(n4428) );
  XNOR U4997 ( .A(n4293), .B(n4289), .Z(n4429) );
  XNOR U4998 ( .A(n4288), .B(n4284), .Z(n4430) );
  XNOR U4999 ( .A(n4283), .B(n4279), .Z(n4431) );
  XNOR U5000 ( .A(n4278), .B(n4274), .Z(n4432) );
  XNOR U5001 ( .A(n4273), .B(n4269), .Z(n4433) );
  XOR U5002 ( .A(n4268), .B(n4265), .Z(n4434) );
  XOR U5003 ( .A(n4435), .B(n4436), .Z(n4265) );
  XOR U5004 ( .A(n4263), .B(n4437), .Z(n4436) );
  XOR U5005 ( .A(n4438), .B(n4439), .Z(n4437) );
  XOR U5006 ( .A(n4440), .B(n4441), .Z(n4439) );
  NAND U5007 ( .A(a[8]), .B(b[30]), .Z(n4441) );
  AND U5008 ( .A(a[7]), .B(b[31]), .Z(n4440) );
  XOR U5009 ( .A(n4442), .B(n4438), .Z(n4435) );
  XOR U5010 ( .A(n4443), .B(n4444), .Z(n4438) );
  NOR U5011 ( .A(n4445), .B(n4446), .Z(n4443) );
  AND U5012 ( .A(a[9]), .B(b[29]), .Z(n4442) );
  XNOR U5013 ( .A(n4447), .B(n4263), .Z(n4264) );
  XOR U5014 ( .A(n4448), .B(n4449), .Z(n4263) );
  ANDN U5015 ( .B(n4450), .A(n4451), .Z(n4448) );
  AND U5016 ( .A(a[10]), .B(b[28]), .Z(n4447) );
  XNOR U5017 ( .A(n4452), .B(n4268), .Z(n4270) );
  XOR U5018 ( .A(n4453), .B(n4454), .Z(n4268) );
  ANDN U5019 ( .B(n4455), .A(n4456), .Z(n4453) );
  AND U5020 ( .A(a[11]), .B(b[27]), .Z(n4452) );
  XNOR U5021 ( .A(n4457), .B(n4273), .Z(n4275) );
  XOR U5022 ( .A(n4458), .B(n4459), .Z(n4273) );
  ANDN U5023 ( .B(n4460), .A(n4461), .Z(n4458) );
  AND U5024 ( .A(a[12]), .B(b[26]), .Z(n4457) );
  XNOR U5025 ( .A(n4462), .B(n4278), .Z(n4280) );
  XOR U5026 ( .A(n4463), .B(n4464), .Z(n4278) );
  ANDN U5027 ( .B(n4465), .A(n4466), .Z(n4463) );
  AND U5028 ( .A(a[13]), .B(b[25]), .Z(n4462) );
  XNOR U5029 ( .A(n4467), .B(n4283), .Z(n4285) );
  XOR U5030 ( .A(n4468), .B(n4469), .Z(n4283) );
  ANDN U5031 ( .B(n4470), .A(n4471), .Z(n4468) );
  AND U5032 ( .A(a[14]), .B(b[24]), .Z(n4467) );
  XNOR U5033 ( .A(n4472), .B(n4288), .Z(n4290) );
  XOR U5034 ( .A(n4473), .B(n4474), .Z(n4288) );
  ANDN U5035 ( .B(n4475), .A(n4476), .Z(n4473) );
  AND U5036 ( .A(a[15]), .B(b[23]), .Z(n4472) );
  XNOR U5037 ( .A(n4477), .B(n4293), .Z(n4295) );
  XOR U5038 ( .A(n4478), .B(n4479), .Z(n4293) );
  ANDN U5039 ( .B(n4480), .A(n4481), .Z(n4478) );
  AND U5040 ( .A(a[16]), .B(b[22]), .Z(n4477) );
  XNOR U5041 ( .A(n4482), .B(n4298), .Z(n4300) );
  XOR U5042 ( .A(n4483), .B(n4484), .Z(n4298) );
  ANDN U5043 ( .B(n4485), .A(n4486), .Z(n4483) );
  AND U5044 ( .A(a[17]), .B(b[21]), .Z(n4482) );
  XNOR U5045 ( .A(n4487), .B(n4303), .Z(n4305) );
  XOR U5046 ( .A(n4488), .B(n4489), .Z(n4303) );
  ANDN U5047 ( .B(n4490), .A(n4491), .Z(n4488) );
  AND U5048 ( .A(a[18]), .B(b[20]), .Z(n4487) );
  XNOR U5049 ( .A(n4492), .B(n4308), .Z(n4310) );
  XOR U5050 ( .A(n4493), .B(n4494), .Z(n4308) );
  ANDN U5051 ( .B(n4495), .A(n4496), .Z(n4493) );
  AND U5052 ( .A(b[19]), .B(a[19]), .Z(n4492) );
  XNOR U5053 ( .A(n4497), .B(n4313), .Z(n4315) );
  XOR U5054 ( .A(n4498), .B(n4499), .Z(n4313) );
  ANDN U5055 ( .B(n4500), .A(n4501), .Z(n4498) );
  AND U5056 ( .A(a[20]), .B(b[18]), .Z(n4497) );
  XNOR U5057 ( .A(n4502), .B(n4318), .Z(n4320) );
  XOR U5058 ( .A(n4503), .B(n4504), .Z(n4318) );
  ANDN U5059 ( .B(n4505), .A(n4506), .Z(n4503) );
  AND U5060 ( .A(b[17]), .B(a[21]), .Z(n4502) );
  XNOR U5061 ( .A(n4507), .B(n4323), .Z(n4325) );
  XOR U5062 ( .A(n4508), .B(n4509), .Z(n4323) );
  ANDN U5063 ( .B(n4510), .A(n4511), .Z(n4508) );
  AND U5064 ( .A(a[22]), .B(b[16]), .Z(n4507) );
  XNOR U5065 ( .A(n4512), .B(n4328), .Z(n4330) );
  XOR U5066 ( .A(n4513), .B(n4514), .Z(n4328) );
  ANDN U5067 ( .B(n4515), .A(n4516), .Z(n4513) );
  AND U5068 ( .A(b[15]), .B(a[23]), .Z(n4512) );
  XNOR U5069 ( .A(n4517), .B(n4333), .Z(n4335) );
  XOR U5070 ( .A(n4518), .B(n4519), .Z(n4333) );
  ANDN U5071 ( .B(n4520), .A(n4521), .Z(n4518) );
  AND U5072 ( .A(a[24]), .B(b[14]), .Z(n4517) );
  XNOR U5073 ( .A(n4522), .B(n4338), .Z(n4340) );
  XOR U5074 ( .A(n4523), .B(n4524), .Z(n4338) );
  ANDN U5075 ( .B(n4525), .A(n4526), .Z(n4523) );
  AND U5076 ( .A(b[13]), .B(a[25]), .Z(n4522) );
  XNOR U5077 ( .A(n4527), .B(n4343), .Z(n4345) );
  XOR U5078 ( .A(n4528), .B(n4529), .Z(n4343) );
  ANDN U5079 ( .B(n4530), .A(n4531), .Z(n4528) );
  AND U5080 ( .A(a[26]), .B(b[12]), .Z(n4527) );
  XNOR U5081 ( .A(n4532), .B(n4348), .Z(n4350) );
  XOR U5082 ( .A(n4533), .B(n4534), .Z(n4348) );
  ANDN U5083 ( .B(n4535), .A(n4536), .Z(n4533) );
  AND U5084 ( .A(b[11]), .B(a[27]), .Z(n4532) );
  XNOR U5085 ( .A(n4537), .B(n4353), .Z(n4355) );
  XOR U5086 ( .A(n4538), .B(n4539), .Z(n4353) );
  ANDN U5087 ( .B(n4540), .A(n4541), .Z(n4538) );
  AND U5088 ( .A(a[28]), .B(b[10]), .Z(n4537) );
  XNOR U5089 ( .A(n4542), .B(n4358), .Z(n4360) );
  XOR U5090 ( .A(n4543), .B(n4544), .Z(n4358) );
  ANDN U5091 ( .B(n4545), .A(n4546), .Z(n4543) );
  AND U5092 ( .A(b[9]), .B(a[29]), .Z(n4542) );
  XNOR U5093 ( .A(n4547), .B(n4363), .Z(n4365) );
  XOR U5094 ( .A(n4548), .B(n4549), .Z(n4363) );
  ANDN U5095 ( .B(n4550), .A(n4551), .Z(n4548) );
  AND U5096 ( .A(a[30]), .B(b[8]), .Z(n4547) );
  XNOR U5097 ( .A(n4552), .B(n4368), .Z(n4370) );
  XOR U5098 ( .A(n4553), .B(n4554), .Z(n4368) );
  ANDN U5099 ( .B(n4555), .A(n4556), .Z(n4553) );
  AND U5100 ( .A(b[7]), .B(a[31]), .Z(n4552) );
  XNOR U5101 ( .A(n4557), .B(n4373), .Z(n4375) );
  XOR U5102 ( .A(n4558), .B(n4559), .Z(n4373) );
  ANDN U5103 ( .B(n4560), .A(n4561), .Z(n4558) );
  AND U5104 ( .A(b[6]), .B(a[32]), .Z(n4557) );
  XNOR U5105 ( .A(n4562), .B(n4378), .Z(n4380) );
  XOR U5106 ( .A(n4563), .B(n4564), .Z(n4378) );
  ANDN U5107 ( .B(n4565), .A(n4566), .Z(n4563) );
  AND U5108 ( .A(b[5]), .B(a[33]), .Z(n4562) );
  XNOR U5109 ( .A(n4567), .B(n4383), .Z(n4385) );
  XOR U5110 ( .A(n4568), .B(n4569), .Z(n4383) );
  ANDN U5111 ( .B(n4570), .A(n4571), .Z(n4568) );
  AND U5112 ( .A(b[4]), .B(a[34]), .Z(n4567) );
  XNOR U5113 ( .A(n4572), .B(n4573), .Z(n4397) );
  NANDN U5114 ( .A(n4574), .B(n4575), .Z(n4573) );
  XNOR U5115 ( .A(n4576), .B(n4388), .Z(n4390) );
  XNOR U5116 ( .A(n4577), .B(n4578), .Z(n4388) );
  AND U5117 ( .A(n4579), .B(n4580), .Z(n4577) );
  AND U5118 ( .A(b[3]), .B(a[35]), .Z(n4576) );
  XNOR U5119 ( .A(n4581), .B(n4582), .Z(swire[37]) );
  XOR U5120 ( .A(n4408), .B(n4583), .Z(n4582) );
  XOR U5121 ( .A(n4407), .B(n4581), .Z(n4583) );
  NAND U5122 ( .A(a[37]), .B(b[0]), .Z(n4407) );
  XNOR U5123 ( .A(n4574), .B(n4575), .Z(n4408) );
  XOR U5124 ( .A(n4572), .B(n4584), .Z(n4575) );
  NAND U5125 ( .A(a[36]), .B(b[1]), .Z(n4584) );
  XOR U5126 ( .A(n4580), .B(n4585), .Z(n4574) );
  XOR U5127 ( .A(n4572), .B(n4579), .Z(n4585) );
  XNOR U5128 ( .A(n4586), .B(n4578), .Z(n4579) );
  AND U5129 ( .A(b[2]), .B(a[35]), .Z(n4586) );
  NANDN U5130 ( .A(n4587), .B(n4588), .Z(n4572) );
  XOR U5131 ( .A(n4578), .B(n4570), .Z(n4589) );
  XNOR U5132 ( .A(n4569), .B(n4565), .Z(n4590) );
  XNOR U5133 ( .A(n4564), .B(n4560), .Z(n4591) );
  XNOR U5134 ( .A(n4559), .B(n4555), .Z(n4592) );
  XNOR U5135 ( .A(n4554), .B(n4550), .Z(n4593) );
  XNOR U5136 ( .A(n4549), .B(n4545), .Z(n4594) );
  XNOR U5137 ( .A(n4544), .B(n4540), .Z(n4595) );
  XNOR U5138 ( .A(n4539), .B(n4535), .Z(n4596) );
  XNOR U5139 ( .A(n4534), .B(n4530), .Z(n4597) );
  XNOR U5140 ( .A(n4529), .B(n4525), .Z(n4598) );
  XNOR U5141 ( .A(n4524), .B(n4520), .Z(n4599) );
  XNOR U5142 ( .A(n4519), .B(n4515), .Z(n4600) );
  XNOR U5143 ( .A(n4514), .B(n4510), .Z(n4601) );
  XNOR U5144 ( .A(n4509), .B(n4505), .Z(n4602) );
  XNOR U5145 ( .A(n4504), .B(n4500), .Z(n4603) );
  XNOR U5146 ( .A(n4499), .B(n4495), .Z(n4604) );
  XNOR U5147 ( .A(n4494), .B(n4490), .Z(n4605) );
  XNOR U5148 ( .A(n4489), .B(n4485), .Z(n4606) );
  XNOR U5149 ( .A(n4484), .B(n4480), .Z(n4607) );
  XNOR U5150 ( .A(n4479), .B(n4475), .Z(n4608) );
  XNOR U5151 ( .A(n4474), .B(n4470), .Z(n4609) );
  XNOR U5152 ( .A(n4469), .B(n4465), .Z(n4610) );
  XNOR U5153 ( .A(n4464), .B(n4460), .Z(n4611) );
  XNOR U5154 ( .A(n4459), .B(n4455), .Z(n4612) );
  XNOR U5155 ( .A(n4454), .B(n4450), .Z(n4613) );
  XOR U5156 ( .A(n4449), .B(n4446), .Z(n4614) );
  XOR U5157 ( .A(n4615), .B(n4616), .Z(n4446) );
  XOR U5158 ( .A(n4444), .B(n4617), .Z(n4616) );
  XOR U5159 ( .A(n4618), .B(n4619), .Z(n4617) );
  XOR U5160 ( .A(n4620), .B(n4621), .Z(n4619) );
  NAND U5161 ( .A(a[7]), .B(b[30]), .Z(n4621) );
  AND U5162 ( .A(a[6]), .B(b[31]), .Z(n4620) );
  XOR U5163 ( .A(n4622), .B(n4618), .Z(n4615) );
  XOR U5164 ( .A(n4623), .B(n4624), .Z(n4618) );
  NOR U5165 ( .A(n4625), .B(n4626), .Z(n4623) );
  AND U5166 ( .A(a[8]), .B(b[29]), .Z(n4622) );
  XNOR U5167 ( .A(n4627), .B(n4444), .Z(n4445) );
  XOR U5168 ( .A(n4628), .B(n4629), .Z(n4444) );
  ANDN U5169 ( .B(n4630), .A(n4631), .Z(n4628) );
  AND U5170 ( .A(a[9]), .B(b[28]), .Z(n4627) );
  XNOR U5171 ( .A(n4632), .B(n4449), .Z(n4451) );
  XOR U5172 ( .A(n4633), .B(n4634), .Z(n4449) );
  ANDN U5173 ( .B(n4635), .A(n4636), .Z(n4633) );
  AND U5174 ( .A(a[10]), .B(b[27]), .Z(n4632) );
  XNOR U5175 ( .A(n4637), .B(n4454), .Z(n4456) );
  XOR U5176 ( .A(n4638), .B(n4639), .Z(n4454) );
  ANDN U5177 ( .B(n4640), .A(n4641), .Z(n4638) );
  AND U5178 ( .A(a[11]), .B(b[26]), .Z(n4637) );
  XNOR U5179 ( .A(n4642), .B(n4459), .Z(n4461) );
  XOR U5180 ( .A(n4643), .B(n4644), .Z(n4459) );
  ANDN U5181 ( .B(n4645), .A(n4646), .Z(n4643) );
  AND U5182 ( .A(a[12]), .B(b[25]), .Z(n4642) );
  XNOR U5183 ( .A(n4647), .B(n4464), .Z(n4466) );
  XOR U5184 ( .A(n4648), .B(n4649), .Z(n4464) );
  ANDN U5185 ( .B(n4650), .A(n4651), .Z(n4648) );
  AND U5186 ( .A(a[13]), .B(b[24]), .Z(n4647) );
  XNOR U5187 ( .A(n4652), .B(n4469), .Z(n4471) );
  XOR U5188 ( .A(n4653), .B(n4654), .Z(n4469) );
  ANDN U5189 ( .B(n4655), .A(n4656), .Z(n4653) );
  AND U5190 ( .A(a[14]), .B(b[23]), .Z(n4652) );
  XNOR U5191 ( .A(n4657), .B(n4474), .Z(n4476) );
  XOR U5192 ( .A(n4658), .B(n4659), .Z(n4474) );
  ANDN U5193 ( .B(n4660), .A(n4661), .Z(n4658) );
  AND U5194 ( .A(a[15]), .B(b[22]), .Z(n4657) );
  XNOR U5195 ( .A(n4662), .B(n4479), .Z(n4481) );
  XOR U5196 ( .A(n4663), .B(n4664), .Z(n4479) );
  ANDN U5197 ( .B(n4665), .A(n4666), .Z(n4663) );
  AND U5198 ( .A(a[16]), .B(b[21]), .Z(n4662) );
  XNOR U5199 ( .A(n4667), .B(n4484), .Z(n4486) );
  XOR U5200 ( .A(n4668), .B(n4669), .Z(n4484) );
  ANDN U5201 ( .B(n4670), .A(n4671), .Z(n4668) );
  AND U5202 ( .A(a[17]), .B(b[20]), .Z(n4667) );
  XNOR U5203 ( .A(n4672), .B(n4489), .Z(n4491) );
  XOR U5204 ( .A(n4673), .B(n4674), .Z(n4489) );
  ANDN U5205 ( .B(n4675), .A(n4676), .Z(n4673) );
  AND U5206 ( .A(a[18]), .B(b[19]), .Z(n4672) );
  XNOR U5207 ( .A(n4677), .B(n4494), .Z(n4496) );
  XOR U5208 ( .A(n4678), .B(n4679), .Z(n4494) );
  ANDN U5209 ( .B(n4680), .A(n4681), .Z(n4678) );
  AND U5210 ( .A(b[18]), .B(a[19]), .Z(n4677) );
  XNOR U5211 ( .A(n4682), .B(n4499), .Z(n4501) );
  XOR U5212 ( .A(n4683), .B(n4684), .Z(n4499) );
  ANDN U5213 ( .B(n4685), .A(n4686), .Z(n4683) );
  AND U5214 ( .A(a[20]), .B(b[17]), .Z(n4682) );
  XNOR U5215 ( .A(n4687), .B(n4504), .Z(n4506) );
  XOR U5216 ( .A(n4688), .B(n4689), .Z(n4504) );
  ANDN U5217 ( .B(n4690), .A(n4691), .Z(n4688) );
  AND U5218 ( .A(b[16]), .B(a[21]), .Z(n4687) );
  XNOR U5219 ( .A(n4692), .B(n4509), .Z(n4511) );
  XOR U5220 ( .A(n4693), .B(n4694), .Z(n4509) );
  ANDN U5221 ( .B(n4695), .A(n4696), .Z(n4693) );
  AND U5222 ( .A(a[22]), .B(b[15]), .Z(n4692) );
  XNOR U5223 ( .A(n4697), .B(n4514), .Z(n4516) );
  XOR U5224 ( .A(n4698), .B(n4699), .Z(n4514) );
  ANDN U5225 ( .B(n4700), .A(n4701), .Z(n4698) );
  AND U5226 ( .A(b[14]), .B(a[23]), .Z(n4697) );
  XNOR U5227 ( .A(n4702), .B(n4519), .Z(n4521) );
  XOR U5228 ( .A(n4703), .B(n4704), .Z(n4519) );
  ANDN U5229 ( .B(n4705), .A(n4706), .Z(n4703) );
  AND U5230 ( .A(a[24]), .B(b[13]), .Z(n4702) );
  XNOR U5231 ( .A(n4707), .B(n4524), .Z(n4526) );
  XOR U5232 ( .A(n4708), .B(n4709), .Z(n4524) );
  ANDN U5233 ( .B(n4710), .A(n4711), .Z(n4708) );
  AND U5234 ( .A(b[12]), .B(a[25]), .Z(n4707) );
  XNOR U5235 ( .A(n4712), .B(n4529), .Z(n4531) );
  XOR U5236 ( .A(n4713), .B(n4714), .Z(n4529) );
  ANDN U5237 ( .B(n4715), .A(n4716), .Z(n4713) );
  AND U5238 ( .A(a[26]), .B(b[11]), .Z(n4712) );
  XNOR U5239 ( .A(n4717), .B(n4534), .Z(n4536) );
  XOR U5240 ( .A(n4718), .B(n4719), .Z(n4534) );
  ANDN U5241 ( .B(n4720), .A(n4721), .Z(n4718) );
  AND U5242 ( .A(b[10]), .B(a[27]), .Z(n4717) );
  XNOR U5243 ( .A(n4722), .B(n4539), .Z(n4541) );
  XOR U5244 ( .A(n4723), .B(n4724), .Z(n4539) );
  ANDN U5245 ( .B(n4725), .A(n4726), .Z(n4723) );
  AND U5246 ( .A(a[28]), .B(b[9]), .Z(n4722) );
  XNOR U5247 ( .A(n4727), .B(n4544), .Z(n4546) );
  XOR U5248 ( .A(n4728), .B(n4729), .Z(n4544) );
  ANDN U5249 ( .B(n4730), .A(n4731), .Z(n4728) );
  AND U5250 ( .A(b[8]), .B(a[29]), .Z(n4727) );
  XNOR U5251 ( .A(n4732), .B(n4549), .Z(n4551) );
  XOR U5252 ( .A(n4733), .B(n4734), .Z(n4549) );
  ANDN U5253 ( .B(n4735), .A(n4736), .Z(n4733) );
  AND U5254 ( .A(a[30]), .B(b[7]), .Z(n4732) );
  XNOR U5255 ( .A(n4737), .B(n4554), .Z(n4556) );
  XOR U5256 ( .A(n4738), .B(n4739), .Z(n4554) );
  ANDN U5257 ( .B(n4740), .A(n4741), .Z(n4738) );
  AND U5258 ( .A(b[6]), .B(a[31]), .Z(n4737) );
  XNOR U5259 ( .A(n4742), .B(n4559), .Z(n4561) );
  XOR U5260 ( .A(n4743), .B(n4744), .Z(n4559) );
  ANDN U5261 ( .B(n4745), .A(n4746), .Z(n4743) );
  AND U5262 ( .A(b[5]), .B(a[32]), .Z(n4742) );
  XNOR U5263 ( .A(n4747), .B(n4564), .Z(n4566) );
  XOR U5264 ( .A(n4748), .B(n4749), .Z(n4564) );
  ANDN U5265 ( .B(n4750), .A(n4751), .Z(n4748) );
  AND U5266 ( .A(b[4]), .B(a[33]), .Z(n4747) );
  XNOR U5267 ( .A(n4752), .B(n4753), .Z(n4578) );
  NANDN U5268 ( .A(n4754), .B(n4755), .Z(n4753) );
  XNOR U5269 ( .A(n4756), .B(n4569), .Z(n4571) );
  XNOR U5270 ( .A(n4757), .B(n4758), .Z(n4569) );
  AND U5271 ( .A(n4759), .B(n4760), .Z(n4757) );
  AND U5272 ( .A(b[3]), .B(a[34]), .Z(n4756) );
  XNOR U5273 ( .A(n4761), .B(n4762), .Z(swire[36]) );
  XOR U5274 ( .A(n4588), .B(n4764), .Z(n4762) );
  XNOR U5275 ( .A(n4587), .B(n4763), .Z(n4764) );
  IV U5276 ( .A(n4761), .Z(n4763) );
  NAND U5277 ( .A(a[36]), .B(b[0]), .Z(n4587) );
  XNOR U5278 ( .A(n4754), .B(n4755), .Z(n4588) );
  XOR U5279 ( .A(n4752), .B(n4765), .Z(n4755) );
  NAND U5280 ( .A(b[1]), .B(a[35]), .Z(n4765) );
  XOR U5281 ( .A(n4760), .B(n4766), .Z(n4754) );
  XOR U5282 ( .A(n4752), .B(n4759), .Z(n4766) );
  XNOR U5283 ( .A(n4767), .B(n4758), .Z(n4759) );
  AND U5284 ( .A(b[2]), .B(a[34]), .Z(n4767) );
  NANDN U5285 ( .A(n4768), .B(n4769), .Z(n4752) );
  XOR U5286 ( .A(n4758), .B(n4750), .Z(n4770) );
  XNOR U5287 ( .A(n4749), .B(n4745), .Z(n4771) );
  XNOR U5288 ( .A(n4744), .B(n4740), .Z(n4772) );
  XNOR U5289 ( .A(n4739), .B(n4735), .Z(n4773) );
  XNOR U5290 ( .A(n4734), .B(n4730), .Z(n4774) );
  XNOR U5291 ( .A(n4729), .B(n4725), .Z(n4775) );
  XNOR U5292 ( .A(n4724), .B(n4720), .Z(n4776) );
  XNOR U5293 ( .A(n4719), .B(n4715), .Z(n4777) );
  XNOR U5294 ( .A(n4714), .B(n4710), .Z(n4778) );
  XNOR U5295 ( .A(n4709), .B(n4705), .Z(n4779) );
  XNOR U5296 ( .A(n4704), .B(n4700), .Z(n4780) );
  XNOR U5297 ( .A(n4699), .B(n4695), .Z(n4781) );
  XNOR U5298 ( .A(n4694), .B(n4690), .Z(n4782) );
  XNOR U5299 ( .A(n4689), .B(n4685), .Z(n4783) );
  XNOR U5300 ( .A(n4684), .B(n4680), .Z(n4784) );
  XNOR U5301 ( .A(n4679), .B(n4675), .Z(n4785) );
  XNOR U5302 ( .A(n4674), .B(n4670), .Z(n4786) );
  XNOR U5303 ( .A(n4669), .B(n4665), .Z(n4787) );
  XNOR U5304 ( .A(n4664), .B(n4660), .Z(n4788) );
  XNOR U5305 ( .A(n4659), .B(n4655), .Z(n4789) );
  XNOR U5306 ( .A(n4654), .B(n4650), .Z(n4790) );
  XNOR U5307 ( .A(n4649), .B(n4645), .Z(n4791) );
  XNOR U5308 ( .A(n4644), .B(n4640), .Z(n4792) );
  XNOR U5309 ( .A(n4639), .B(n4635), .Z(n4793) );
  XNOR U5310 ( .A(n4634), .B(n4630), .Z(n4794) );
  XOR U5311 ( .A(n4629), .B(n4626), .Z(n4795) );
  XOR U5312 ( .A(n4796), .B(n4797), .Z(n4626) );
  XOR U5313 ( .A(n4624), .B(n4798), .Z(n4797) );
  XOR U5314 ( .A(n4799), .B(n4800), .Z(n4798) );
  XOR U5315 ( .A(n4801), .B(n4802), .Z(n4800) );
  NAND U5316 ( .A(a[6]), .B(b[30]), .Z(n4802) );
  AND U5317 ( .A(a[5]), .B(b[31]), .Z(n4801) );
  XOR U5318 ( .A(n4803), .B(n4799), .Z(n4796) );
  XOR U5319 ( .A(n4804), .B(n4805), .Z(n4799) );
  NOR U5320 ( .A(n4806), .B(n4807), .Z(n4804) );
  AND U5321 ( .A(a[7]), .B(b[29]), .Z(n4803) );
  XNOR U5322 ( .A(n4808), .B(n4624), .Z(n4625) );
  XOR U5323 ( .A(n4809), .B(n4810), .Z(n4624) );
  ANDN U5324 ( .B(n4811), .A(n4812), .Z(n4809) );
  AND U5325 ( .A(a[8]), .B(b[28]), .Z(n4808) );
  XNOR U5326 ( .A(n4813), .B(n4629), .Z(n4631) );
  XOR U5327 ( .A(n4814), .B(n4815), .Z(n4629) );
  ANDN U5328 ( .B(n4816), .A(n4817), .Z(n4814) );
  AND U5329 ( .A(a[9]), .B(b[27]), .Z(n4813) );
  XNOR U5330 ( .A(n4818), .B(n4634), .Z(n4636) );
  XOR U5331 ( .A(n4819), .B(n4820), .Z(n4634) );
  ANDN U5332 ( .B(n4821), .A(n4822), .Z(n4819) );
  AND U5333 ( .A(a[10]), .B(b[26]), .Z(n4818) );
  XNOR U5334 ( .A(n4823), .B(n4639), .Z(n4641) );
  XOR U5335 ( .A(n4824), .B(n4825), .Z(n4639) );
  ANDN U5336 ( .B(n4826), .A(n4827), .Z(n4824) );
  AND U5337 ( .A(a[11]), .B(b[25]), .Z(n4823) );
  XNOR U5338 ( .A(n4828), .B(n4644), .Z(n4646) );
  XOR U5339 ( .A(n4829), .B(n4830), .Z(n4644) );
  ANDN U5340 ( .B(n4831), .A(n4832), .Z(n4829) );
  AND U5341 ( .A(a[12]), .B(b[24]), .Z(n4828) );
  XNOR U5342 ( .A(n4833), .B(n4649), .Z(n4651) );
  XOR U5343 ( .A(n4834), .B(n4835), .Z(n4649) );
  ANDN U5344 ( .B(n4836), .A(n4837), .Z(n4834) );
  AND U5345 ( .A(a[13]), .B(b[23]), .Z(n4833) );
  XNOR U5346 ( .A(n4838), .B(n4654), .Z(n4656) );
  XOR U5347 ( .A(n4839), .B(n4840), .Z(n4654) );
  ANDN U5348 ( .B(n4841), .A(n4842), .Z(n4839) );
  AND U5349 ( .A(a[14]), .B(b[22]), .Z(n4838) );
  XNOR U5350 ( .A(n4843), .B(n4659), .Z(n4661) );
  XOR U5351 ( .A(n4844), .B(n4845), .Z(n4659) );
  ANDN U5352 ( .B(n4846), .A(n4847), .Z(n4844) );
  AND U5353 ( .A(a[15]), .B(b[21]), .Z(n4843) );
  XNOR U5354 ( .A(n4848), .B(n4664), .Z(n4666) );
  XOR U5355 ( .A(n4849), .B(n4850), .Z(n4664) );
  ANDN U5356 ( .B(n4851), .A(n4852), .Z(n4849) );
  AND U5357 ( .A(a[16]), .B(b[20]), .Z(n4848) );
  XNOR U5358 ( .A(n4853), .B(n4669), .Z(n4671) );
  XOR U5359 ( .A(n4854), .B(n4855), .Z(n4669) );
  ANDN U5360 ( .B(n4856), .A(n4857), .Z(n4854) );
  AND U5361 ( .A(a[17]), .B(b[19]), .Z(n4853) );
  XNOR U5362 ( .A(n4858), .B(n4674), .Z(n4676) );
  XOR U5363 ( .A(n4859), .B(n4860), .Z(n4674) );
  ANDN U5364 ( .B(n4861), .A(n4862), .Z(n4859) );
  AND U5365 ( .A(a[18]), .B(b[18]), .Z(n4858) );
  XNOR U5366 ( .A(n4863), .B(n4679), .Z(n4681) );
  XOR U5367 ( .A(n4864), .B(n4865), .Z(n4679) );
  ANDN U5368 ( .B(n4866), .A(n4867), .Z(n4864) );
  AND U5369 ( .A(b[17]), .B(a[19]), .Z(n4863) );
  XNOR U5370 ( .A(n4868), .B(n4684), .Z(n4686) );
  XOR U5371 ( .A(n4869), .B(n4870), .Z(n4684) );
  ANDN U5372 ( .B(n4871), .A(n4872), .Z(n4869) );
  AND U5373 ( .A(a[20]), .B(b[16]), .Z(n4868) );
  XNOR U5374 ( .A(n4873), .B(n4689), .Z(n4691) );
  XOR U5375 ( .A(n4874), .B(n4875), .Z(n4689) );
  ANDN U5376 ( .B(n4876), .A(n4877), .Z(n4874) );
  AND U5377 ( .A(b[15]), .B(a[21]), .Z(n4873) );
  XNOR U5378 ( .A(n4878), .B(n4694), .Z(n4696) );
  XOR U5379 ( .A(n4879), .B(n4880), .Z(n4694) );
  ANDN U5380 ( .B(n4881), .A(n4882), .Z(n4879) );
  AND U5381 ( .A(a[22]), .B(b[14]), .Z(n4878) );
  XNOR U5382 ( .A(n4883), .B(n4699), .Z(n4701) );
  XOR U5383 ( .A(n4884), .B(n4885), .Z(n4699) );
  ANDN U5384 ( .B(n4886), .A(n4887), .Z(n4884) );
  AND U5385 ( .A(b[13]), .B(a[23]), .Z(n4883) );
  XNOR U5386 ( .A(n4888), .B(n4704), .Z(n4706) );
  XOR U5387 ( .A(n4889), .B(n4890), .Z(n4704) );
  ANDN U5388 ( .B(n4891), .A(n4892), .Z(n4889) );
  AND U5389 ( .A(a[24]), .B(b[12]), .Z(n4888) );
  XNOR U5390 ( .A(n4893), .B(n4709), .Z(n4711) );
  XOR U5391 ( .A(n4894), .B(n4895), .Z(n4709) );
  ANDN U5392 ( .B(n4896), .A(n4897), .Z(n4894) );
  AND U5393 ( .A(b[11]), .B(a[25]), .Z(n4893) );
  XNOR U5394 ( .A(n4898), .B(n4714), .Z(n4716) );
  XOR U5395 ( .A(n4899), .B(n4900), .Z(n4714) );
  ANDN U5396 ( .B(n4901), .A(n4902), .Z(n4899) );
  AND U5397 ( .A(a[26]), .B(b[10]), .Z(n4898) );
  XNOR U5398 ( .A(n4903), .B(n4719), .Z(n4721) );
  XOR U5399 ( .A(n4904), .B(n4905), .Z(n4719) );
  ANDN U5400 ( .B(n4906), .A(n4907), .Z(n4904) );
  AND U5401 ( .A(b[9]), .B(a[27]), .Z(n4903) );
  XNOR U5402 ( .A(n4908), .B(n4724), .Z(n4726) );
  XOR U5403 ( .A(n4909), .B(n4910), .Z(n4724) );
  ANDN U5404 ( .B(n4911), .A(n4912), .Z(n4909) );
  AND U5405 ( .A(a[28]), .B(b[8]), .Z(n4908) );
  XNOR U5406 ( .A(n4913), .B(n4729), .Z(n4731) );
  XOR U5407 ( .A(n4914), .B(n4915), .Z(n4729) );
  ANDN U5408 ( .B(n4916), .A(n4917), .Z(n4914) );
  AND U5409 ( .A(b[7]), .B(a[29]), .Z(n4913) );
  XNOR U5410 ( .A(n4918), .B(n4734), .Z(n4736) );
  XOR U5411 ( .A(n4919), .B(n4920), .Z(n4734) );
  ANDN U5412 ( .B(n4921), .A(n4922), .Z(n4919) );
  AND U5413 ( .A(b[6]), .B(a[30]), .Z(n4918) );
  XNOR U5414 ( .A(n4923), .B(n4739), .Z(n4741) );
  XOR U5415 ( .A(n4924), .B(n4925), .Z(n4739) );
  ANDN U5416 ( .B(n4926), .A(n4927), .Z(n4924) );
  AND U5417 ( .A(b[5]), .B(a[31]), .Z(n4923) );
  XNOR U5418 ( .A(n4928), .B(n4744), .Z(n4746) );
  XOR U5419 ( .A(n4929), .B(n4930), .Z(n4744) );
  ANDN U5420 ( .B(n4931), .A(n4932), .Z(n4929) );
  AND U5421 ( .A(b[4]), .B(a[32]), .Z(n4928) );
  XNOR U5422 ( .A(n4933), .B(n4934), .Z(n4758) );
  NANDN U5423 ( .A(n4935), .B(n4936), .Z(n4934) );
  XNOR U5424 ( .A(n4937), .B(n4749), .Z(n4751) );
  XNOR U5425 ( .A(n4938), .B(n4939), .Z(n4749) );
  AND U5426 ( .A(n4940), .B(n4941), .Z(n4938) );
  AND U5427 ( .A(b[3]), .B(a[33]), .Z(n4937) );
  XNOR U5428 ( .A(n4942), .B(n4943), .Z(swire[35]) );
  XOR U5429 ( .A(n4769), .B(n4944), .Z(n4943) );
  XOR U5430 ( .A(n4768), .B(n4942), .Z(n4944) );
  NAND U5431 ( .A(a[35]), .B(b[0]), .Z(n4768) );
  XNOR U5432 ( .A(n4935), .B(n4936), .Z(n4769) );
  XOR U5433 ( .A(n4933), .B(n4945), .Z(n4936) );
  NAND U5434 ( .A(a[34]), .B(b[1]), .Z(n4945) );
  XOR U5435 ( .A(n4941), .B(n4946), .Z(n4935) );
  XOR U5436 ( .A(n4933), .B(n4940), .Z(n4946) );
  XNOR U5437 ( .A(n4947), .B(n4939), .Z(n4940) );
  AND U5438 ( .A(b[2]), .B(a[33]), .Z(n4947) );
  NANDN U5439 ( .A(n4948), .B(n4949), .Z(n4933) );
  XOR U5440 ( .A(n4939), .B(n4931), .Z(n4950) );
  XNOR U5441 ( .A(n4930), .B(n4926), .Z(n4951) );
  XNOR U5442 ( .A(n4925), .B(n4921), .Z(n4952) );
  XNOR U5443 ( .A(n4920), .B(n4916), .Z(n4953) );
  XNOR U5444 ( .A(n4915), .B(n4911), .Z(n4954) );
  XNOR U5445 ( .A(n4910), .B(n4906), .Z(n4955) );
  XNOR U5446 ( .A(n4905), .B(n4901), .Z(n4956) );
  XNOR U5447 ( .A(n4900), .B(n4896), .Z(n4957) );
  XNOR U5448 ( .A(n4895), .B(n4891), .Z(n4958) );
  XNOR U5449 ( .A(n4890), .B(n4886), .Z(n4959) );
  XNOR U5450 ( .A(n4885), .B(n4881), .Z(n4960) );
  XNOR U5451 ( .A(n4880), .B(n4876), .Z(n4961) );
  XNOR U5452 ( .A(n4875), .B(n4871), .Z(n4962) );
  XNOR U5453 ( .A(n4870), .B(n4866), .Z(n4963) );
  XNOR U5454 ( .A(n4865), .B(n4861), .Z(n4964) );
  XNOR U5455 ( .A(n4860), .B(n4856), .Z(n4965) );
  XNOR U5456 ( .A(n4855), .B(n4851), .Z(n4966) );
  XNOR U5457 ( .A(n4850), .B(n4846), .Z(n4967) );
  XNOR U5458 ( .A(n4845), .B(n4841), .Z(n4968) );
  XNOR U5459 ( .A(n4840), .B(n4836), .Z(n4969) );
  XNOR U5460 ( .A(n4835), .B(n4831), .Z(n4970) );
  XNOR U5461 ( .A(n4830), .B(n4826), .Z(n4971) );
  XNOR U5462 ( .A(n4825), .B(n4821), .Z(n4972) );
  XNOR U5463 ( .A(n4820), .B(n4816), .Z(n4973) );
  XNOR U5464 ( .A(n4815), .B(n4811), .Z(n4974) );
  XOR U5465 ( .A(n4810), .B(n4807), .Z(n4975) );
  XOR U5466 ( .A(n4976), .B(n4977), .Z(n4807) );
  XOR U5467 ( .A(n4805), .B(n4978), .Z(n4977) );
  XOR U5468 ( .A(n4979), .B(n4980), .Z(n4978) );
  XOR U5469 ( .A(n4981), .B(n4982), .Z(n4980) );
  NAND U5470 ( .A(a[5]), .B(b[30]), .Z(n4982) );
  AND U5471 ( .A(a[4]), .B(b[31]), .Z(n4981) );
  XOR U5472 ( .A(n4983), .B(n4979), .Z(n4976) );
  XOR U5473 ( .A(n4984), .B(n4985), .Z(n4979) );
  NOR U5474 ( .A(n4986), .B(n4987), .Z(n4984) );
  AND U5475 ( .A(a[6]), .B(b[29]), .Z(n4983) );
  XNOR U5476 ( .A(n4988), .B(n4805), .Z(n4806) );
  XOR U5477 ( .A(n4989), .B(n4990), .Z(n4805) );
  ANDN U5478 ( .B(n4991), .A(n4992), .Z(n4989) );
  AND U5479 ( .A(a[7]), .B(b[28]), .Z(n4988) );
  XNOR U5480 ( .A(n4993), .B(n4810), .Z(n4812) );
  XOR U5481 ( .A(n4994), .B(n4995), .Z(n4810) );
  ANDN U5482 ( .B(n4996), .A(n4997), .Z(n4994) );
  AND U5483 ( .A(a[8]), .B(b[27]), .Z(n4993) );
  XNOR U5484 ( .A(n4998), .B(n4815), .Z(n4817) );
  XOR U5485 ( .A(n4999), .B(n5000), .Z(n4815) );
  ANDN U5486 ( .B(n5001), .A(n5002), .Z(n4999) );
  AND U5487 ( .A(a[9]), .B(b[26]), .Z(n4998) );
  XNOR U5488 ( .A(n5003), .B(n4820), .Z(n4822) );
  XOR U5489 ( .A(n5004), .B(n5005), .Z(n4820) );
  ANDN U5490 ( .B(n5006), .A(n5007), .Z(n5004) );
  AND U5491 ( .A(a[10]), .B(b[25]), .Z(n5003) );
  XNOR U5492 ( .A(n5008), .B(n4825), .Z(n4827) );
  XOR U5493 ( .A(n5009), .B(n5010), .Z(n4825) );
  ANDN U5494 ( .B(n5011), .A(n5012), .Z(n5009) );
  AND U5495 ( .A(a[11]), .B(b[24]), .Z(n5008) );
  XNOR U5496 ( .A(n5013), .B(n4830), .Z(n4832) );
  XOR U5497 ( .A(n5014), .B(n5015), .Z(n4830) );
  ANDN U5498 ( .B(n5016), .A(n5017), .Z(n5014) );
  AND U5499 ( .A(a[12]), .B(b[23]), .Z(n5013) );
  XNOR U5500 ( .A(n5018), .B(n4835), .Z(n4837) );
  XOR U5501 ( .A(n5019), .B(n5020), .Z(n4835) );
  ANDN U5502 ( .B(n5021), .A(n5022), .Z(n5019) );
  AND U5503 ( .A(a[13]), .B(b[22]), .Z(n5018) );
  XNOR U5504 ( .A(n5023), .B(n4840), .Z(n4842) );
  XOR U5505 ( .A(n5024), .B(n5025), .Z(n4840) );
  ANDN U5506 ( .B(n5026), .A(n5027), .Z(n5024) );
  AND U5507 ( .A(a[14]), .B(b[21]), .Z(n5023) );
  XNOR U5508 ( .A(n5028), .B(n4845), .Z(n4847) );
  XOR U5509 ( .A(n5029), .B(n5030), .Z(n4845) );
  ANDN U5510 ( .B(n5031), .A(n5032), .Z(n5029) );
  AND U5511 ( .A(a[15]), .B(b[20]), .Z(n5028) );
  XNOR U5512 ( .A(n5033), .B(n4850), .Z(n4852) );
  XOR U5513 ( .A(n5034), .B(n5035), .Z(n4850) );
  ANDN U5514 ( .B(n5036), .A(n5037), .Z(n5034) );
  AND U5515 ( .A(a[16]), .B(b[19]), .Z(n5033) );
  XNOR U5516 ( .A(n5038), .B(n4855), .Z(n4857) );
  XOR U5517 ( .A(n5039), .B(n5040), .Z(n4855) );
  ANDN U5518 ( .B(n5041), .A(n5042), .Z(n5039) );
  AND U5519 ( .A(a[17]), .B(b[18]), .Z(n5038) );
  XNOR U5520 ( .A(n5043), .B(n4860), .Z(n4862) );
  XOR U5521 ( .A(n5044), .B(n5045), .Z(n4860) );
  ANDN U5522 ( .B(n5046), .A(n5047), .Z(n5044) );
  AND U5523 ( .A(a[18]), .B(b[17]), .Z(n5043) );
  XNOR U5524 ( .A(n5048), .B(n4865), .Z(n4867) );
  XOR U5525 ( .A(n5049), .B(n5050), .Z(n4865) );
  ANDN U5526 ( .B(n5051), .A(n5052), .Z(n5049) );
  AND U5527 ( .A(b[16]), .B(a[19]), .Z(n5048) );
  XNOR U5528 ( .A(n5053), .B(n4870), .Z(n4872) );
  XOR U5529 ( .A(n5054), .B(n5055), .Z(n4870) );
  ANDN U5530 ( .B(n5056), .A(n5057), .Z(n5054) );
  AND U5531 ( .A(a[20]), .B(b[15]), .Z(n5053) );
  XNOR U5532 ( .A(n5058), .B(n4875), .Z(n4877) );
  XOR U5533 ( .A(n5059), .B(n5060), .Z(n4875) );
  ANDN U5534 ( .B(n5061), .A(n5062), .Z(n5059) );
  AND U5535 ( .A(b[14]), .B(a[21]), .Z(n5058) );
  XNOR U5536 ( .A(n5063), .B(n4880), .Z(n4882) );
  XOR U5537 ( .A(n5064), .B(n5065), .Z(n4880) );
  ANDN U5538 ( .B(n5066), .A(n5067), .Z(n5064) );
  AND U5539 ( .A(a[22]), .B(b[13]), .Z(n5063) );
  XNOR U5540 ( .A(n5068), .B(n4885), .Z(n4887) );
  XOR U5541 ( .A(n5069), .B(n5070), .Z(n4885) );
  ANDN U5542 ( .B(n5071), .A(n5072), .Z(n5069) );
  AND U5543 ( .A(b[12]), .B(a[23]), .Z(n5068) );
  XNOR U5544 ( .A(n5073), .B(n4890), .Z(n4892) );
  XOR U5545 ( .A(n5074), .B(n5075), .Z(n4890) );
  ANDN U5546 ( .B(n5076), .A(n5077), .Z(n5074) );
  AND U5547 ( .A(a[24]), .B(b[11]), .Z(n5073) );
  XNOR U5548 ( .A(n5078), .B(n4895), .Z(n4897) );
  XOR U5549 ( .A(n5079), .B(n5080), .Z(n4895) );
  ANDN U5550 ( .B(n5081), .A(n5082), .Z(n5079) );
  AND U5551 ( .A(b[10]), .B(a[25]), .Z(n5078) );
  XNOR U5552 ( .A(n5083), .B(n4900), .Z(n4902) );
  XOR U5553 ( .A(n5084), .B(n5085), .Z(n4900) );
  ANDN U5554 ( .B(n5086), .A(n5087), .Z(n5084) );
  AND U5555 ( .A(a[26]), .B(b[9]), .Z(n5083) );
  XNOR U5556 ( .A(n5088), .B(n4905), .Z(n4907) );
  XOR U5557 ( .A(n5089), .B(n5090), .Z(n4905) );
  ANDN U5558 ( .B(n5091), .A(n5092), .Z(n5089) );
  AND U5559 ( .A(b[8]), .B(a[27]), .Z(n5088) );
  XNOR U5560 ( .A(n5093), .B(n4910), .Z(n4912) );
  XOR U5561 ( .A(n5094), .B(n5095), .Z(n4910) );
  ANDN U5562 ( .B(n5096), .A(n5097), .Z(n5094) );
  AND U5563 ( .A(a[28]), .B(b[7]), .Z(n5093) );
  XNOR U5564 ( .A(n5098), .B(n4915), .Z(n4917) );
  XOR U5565 ( .A(n5099), .B(n5100), .Z(n4915) );
  ANDN U5566 ( .B(n5101), .A(n5102), .Z(n5099) );
  AND U5567 ( .A(b[6]), .B(a[29]), .Z(n5098) );
  XNOR U5568 ( .A(n5103), .B(n4920), .Z(n4922) );
  XOR U5569 ( .A(n5104), .B(n5105), .Z(n4920) );
  ANDN U5570 ( .B(n5106), .A(n5107), .Z(n5104) );
  AND U5571 ( .A(b[5]), .B(a[30]), .Z(n5103) );
  XNOR U5572 ( .A(n5108), .B(n4925), .Z(n4927) );
  XOR U5573 ( .A(n5109), .B(n5110), .Z(n4925) );
  ANDN U5574 ( .B(n5111), .A(n5112), .Z(n5109) );
  AND U5575 ( .A(b[4]), .B(a[31]), .Z(n5108) );
  XNOR U5576 ( .A(n5113), .B(n5114), .Z(n4939) );
  NANDN U5577 ( .A(n5115), .B(n5116), .Z(n5114) );
  XNOR U5578 ( .A(n5117), .B(n4930), .Z(n4932) );
  XNOR U5579 ( .A(n5118), .B(n5119), .Z(n4930) );
  AND U5580 ( .A(n5120), .B(n5121), .Z(n5118) );
  AND U5581 ( .A(b[3]), .B(a[32]), .Z(n5117) );
  XNOR U5582 ( .A(n5122), .B(n5123), .Z(swire[34]) );
  XOR U5583 ( .A(n4949), .B(n5125), .Z(n5123) );
  XNOR U5584 ( .A(n4948), .B(n5124), .Z(n5125) );
  IV U5585 ( .A(n5122), .Z(n5124) );
  NAND U5586 ( .A(a[34]), .B(b[0]), .Z(n4948) );
  XNOR U5587 ( .A(n5115), .B(n5116), .Z(n4949) );
  XOR U5588 ( .A(n5113), .B(n5126), .Z(n5116) );
  NAND U5589 ( .A(b[1]), .B(a[33]), .Z(n5126) );
  XOR U5590 ( .A(n5121), .B(n5127), .Z(n5115) );
  XOR U5591 ( .A(n5113), .B(n5120), .Z(n5127) );
  XNOR U5592 ( .A(n5128), .B(n5119), .Z(n5120) );
  AND U5593 ( .A(b[2]), .B(a[32]), .Z(n5128) );
  NANDN U5594 ( .A(n5129), .B(n5130), .Z(n5113) );
  XOR U5595 ( .A(n5119), .B(n5111), .Z(n5131) );
  XNOR U5596 ( .A(n5110), .B(n5106), .Z(n5132) );
  XNOR U5597 ( .A(n5105), .B(n5101), .Z(n5133) );
  XNOR U5598 ( .A(n5100), .B(n5096), .Z(n5134) );
  XNOR U5599 ( .A(n5095), .B(n5091), .Z(n5135) );
  XNOR U5600 ( .A(n5090), .B(n5086), .Z(n5136) );
  XNOR U5601 ( .A(n5085), .B(n5081), .Z(n5137) );
  XNOR U5602 ( .A(n5080), .B(n5076), .Z(n5138) );
  XNOR U5603 ( .A(n5075), .B(n5071), .Z(n5139) );
  XNOR U5604 ( .A(n5070), .B(n5066), .Z(n5140) );
  XNOR U5605 ( .A(n5065), .B(n5061), .Z(n5141) );
  XNOR U5606 ( .A(n5060), .B(n5056), .Z(n5142) );
  XNOR U5607 ( .A(n5055), .B(n5051), .Z(n5143) );
  XNOR U5608 ( .A(n5050), .B(n5046), .Z(n5144) );
  XNOR U5609 ( .A(n5045), .B(n5041), .Z(n5145) );
  XNOR U5610 ( .A(n5040), .B(n5036), .Z(n5146) );
  XNOR U5611 ( .A(n5035), .B(n5031), .Z(n5147) );
  XNOR U5612 ( .A(n5030), .B(n5026), .Z(n5148) );
  XNOR U5613 ( .A(n5025), .B(n5021), .Z(n5149) );
  XNOR U5614 ( .A(n5020), .B(n5016), .Z(n5150) );
  XNOR U5615 ( .A(n5015), .B(n5011), .Z(n5151) );
  XNOR U5616 ( .A(n5010), .B(n5006), .Z(n5152) );
  XNOR U5617 ( .A(n5005), .B(n5001), .Z(n5153) );
  XNOR U5618 ( .A(n5000), .B(n4996), .Z(n5154) );
  XNOR U5619 ( .A(n4995), .B(n4991), .Z(n5155) );
  XOR U5620 ( .A(n4990), .B(n4987), .Z(n5156) );
  XOR U5621 ( .A(n5157), .B(n5158), .Z(n4987) );
  XOR U5622 ( .A(n4985), .B(n5159), .Z(n5158) );
  XOR U5623 ( .A(n5160), .B(n5161), .Z(n5159) );
  XOR U5624 ( .A(n5162), .B(n5163), .Z(n5161) );
  NAND U5625 ( .A(a[4]), .B(b[30]), .Z(n5163) );
  AND U5626 ( .A(a[3]), .B(b[31]), .Z(n5162) );
  XOR U5627 ( .A(n5164), .B(n5160), .Z(n5157) );
  XOR U5628 ( .A(n5165), .B(n5166), .Z(n5160) );
  NOR U5629 ( .A(n5167), .B(n5168), .Z(n5165) );
  AND U5630 ( .A(a[5]), .B(b[29]), .Z(n5164) );
  XNOR U5631 ( .A(n5169), .B(n4985), .Z(n4986) );
  XOR U5632 ( .A(n5170), .B(n5171), .Z(n4985) );
  ANDN U5633 ( .B(n5172), .A(n5173), .Z(n5170) );
  AND U5634 ( .A(a[6]), .B(b[28]), .Z(n5169) );
  XNOR U5635 ( .A(n5174), .B(n4990), .Z(n4992) );
  XOR U5636 ( .A(n5175), .B(n5176), .Z(n4990) );
  ANDN U5637 ( .B(n5177), .A(n5178), .Z(n5175) );
  AND U5638 ( .A(a[7]), .B(b[27]), .Z(n5174) );
  XNOR U5639 ( .A(n5179), .B(n4995), .Z(n4997) );
  XOR U5640 ( .A(n5180), .B(n5181), .Z(n4995) );
  ANDN U5641 ( .B(n5182), .A(n5183), .Z(n5180) );
  AND U5642 ( .A(a[8]), .B(b[26]), .Z(n5179) );
  XNOR U5643 ( .A(n5184), .B(n5000), .Z(n5002) );
  XOR U5644 ( .A(n5185), .B(n5186), .Z(n5000) );
  ANDN U5645 ( .B(n5187), .A(n5188), .Z(n5185) );
  AND U5646 ( .A(a[9]), .B(b[25]), .Z(n5184) );
  XNOR U5647 ( .A(n5189), .B(n5005), .Z(n5007) );
  XOR U5648 ( .A(n5190), .B(n5191), .Z(n5005) );
  ANDN U5649 ( .B(n5192), .A(n5193), .Z(n5190) );
  AND U5650 ( .A(a[10]), .B(b[24]), .Z(n5189) );
  XNOR U5651 ( .A(n5194), .B(n5010), .Z(n5012) );
  XOR U5652 ( .A(n5195), .B(n5196), .Z(n5010) );
  ANDN U5653 ( .B(n5197), .A(n5198), .Z(n5195) );
  AND U5654 ( .A(a[11]), .B(b[23]), .Z(n5194) );
  XNOR U5655 ( .A(n5199), .B(n5015), .Z(n5017) );
  XOR U5656 ( .A(n5200), .B(n5201), .Z(n5015) );
  ANDN U5657 ( .B(n5202), .A(n5203), .Z(n5200) );
  AND U5658 ( .A(a[12]), .B(b[22]), .Z(n5199) );
  XNOR U5659 ( .A(n5204), .B(n5020), .Z(n5022) );
  XOR U5660 ( .A(n5205), .B(n5206), .Z(n5020) );
  ANDN U5661 ( .B(n5207), .A(n5208), .Z(n5205) );
  AND U5662 ( .A(a[13]), .B(b[21]), .Z(n5204) );
  XNOR U5663 ( .A(n5209), .B(n5025), .Z(n5027) );
  XOR U5664 ( .A(n5210), .B(n5211), .Z(n5025) );
  ANDN U5665 ( .B(n5212), .A(n5213), .Z(n5210) );
  AND U5666 ( .A(a[14]), .B(b[20]), .Z(n5209) );
  XNOR U5667 ( .A(n5214), .B(n5030), .Z(n5032) );
  XOR U5668 ( .A(n5215), .B(n5216), .Z(n5030) );
  ANDN U5669 ( .B(n5217), .A(n5218), .Z(n5215) );
  AND U5670 ( .A(a[15]), .B(b[19]), .Z(n5214) );
  XNOR U5671 ( .A(n5219), .B(n5035), .Z(n5037) );
  XOR U5672 ( .A(n5220), .B(n5221), .Z(n5035) );
  ANDN U5673 ( .B(n5222), .A(n5223), .Z(n5220) );
  AND U5674 ( .A(a[16]), .B(b[18]), .Z(n5219) );
  XNOR U5675 ( .A(n5224), .B(n5040), .Z(n5042) );
  XOR U5676 ( .A(n5225), .B(n5226), .Z(n5040) );
  ANDN U5677 ( .B(n5227), .A(n5228), .Z(n5225) );
  AND U5678 ( .A(b[17]), .B(a[17]), .Z(n5224) );
  XNOR U5679 ( .A(n5229), .B(n5045), .Z(n5047) );
  XOR U5680 ( .A(n5230), .B(n5231), .Z(n5045) );
  ANDN U5681 ( .B(n5232), .A(n5233), .Z(n5230) );
  AND U5682 ( .A(a[18]), .B(b[16]), .Z(n5229) );
  XNOR U5683 ( .A(n5234), .B(n5050), .Z(n5052) );
  XOR U5684 ( .A(n5235), .B(n5236), .Z(n5050) );
  ANDN U5685 ( .B(n5237), .A(n5238), .Z(n5235) );
  AND U5686 ( .A(b[15]), .B(a[19]), .Z(n5234) );
  XNOR U5687 ( .A(n5239), .B(n5055), .Z(n5057) );
  XOR U5688 ( .A(n5240), .B(n5241), .Z(n5055) );
  ANDN U5689 ( .B(n5242), .A(n5243), .Z(n5240) );
  AND U5690 ( .A(a[20]), .B(b[14]), .Z(n5239) );
  XNOR U5691 ( .A(n5244), .B(n5060), .Z(n5062) );
  XOR U5692 ( .A(n5245), .B(n5246), .Z(n5060) );
  ANDN U5693 ( .B(n5247), .A(n5248), .Z(n5245) );
  AND U5694 ( .A(b[13]), .B(a[21]), .Z(n5244) );
  XNOR U5695 ( .A(n5249), .B(n5065), .Z(n5067) );
  XOR U5696 ( .A(n5250), .B(n5251), .Z(n5065) );
  ANDN U5697 ( .B(n5252), .A(n5253), .Z(n5250) );
  AND U5698 ( .A(a[22]), .B(b[12]), .Z(n5249) );
  XNOR U5699 ( .A(n5254), .B(n5070), .Z(n5072) );
  XOR U5700 ( .A(n5255), .B(n5256), .Z(n5070) );
  ANDN U5701 ( .B(n5257), .A(n5258), .Z(n5255) );
  AND U5702 ( .A(b[11]), .B(a[23]), .Z(n5254) );
  XNOR U5703 ( .A(n5259), .B(n5075), .Z(n5077) );
  XOR U5704 ( .A(n5260), .B(n5261), .Z(n5075) );
  ANDN U5705 ( .B(n5262), .A(n5263), .Z(n5260) );
  AND U5706 ( .A(a[24]), .B(b[10]), .Z(n5259) );
  XNOR U5707 ( .A(n5264), .B(n5080), .Z(n5082) );
  XOR U5708 ( .A(n5265), .B(n5266), .Z(n5080) );
  ANDN U5709 ( .B(n5267), .A(n5268), .Z(n5265) );
  AND U5710 ( .A(b[9]), .B(a[25]), .Z(n5264) );
  XNOR U5711 ( .A(n5269), .B(n5085), .Z(n5087) );
  XOR U5712 ( .A(n5270), .B(n5271), .Z(n5085) );
  ANDN U5713 ( .B(n5272), .A(n5273), .Z(n5270) );
  AND U5714 ( .A(a[26]), .B(b[8]), .Z(n5269) );
  XNOR U5715 ( .A(n5274), .B(n5090), .Z(n5092) );
  XOR U5716 ( .A(n5275), .B(n5276), .Z(n5090) );
  ANDN U5717 ( .B(n5277), .A(n5278), .Z(n5275) );
  AND U5718 ( .A(b[7]), .B(a[27]), .Z(n5274) );
  XNOR U5719 ( .A(n5279), .B(n5095), .Z(n5097) );
  XOR U5720 ( .A(n5280), .B(n5281), .Z(n5095) );
  ANDN U5721 ( .B(n5282), .A(n5283), .Z(n5280) );
  AND U5722 ( .A(b[6]), .B(a[28]), .Z(n5279) );
  XNOR U5723 ( .A(n5284), .B(n5100), .Z(n5102) );
  XOR U5724 ( .A(n5285), .B(n5286), .Z(n5100) );
  ANDN U5725 ( .B(n5287), .A(n5288), .Z(n5285) );
  AND U5726 ( .A(b[5]), .B(a[29]), .Z(n5284) );
  XNOR U5727 ( .A(n5289), .B(n5105), .Z(n5107) );
  XOR U5728 ( .A(n5290), .B(n5291), .Z(n5105) );
  ANDN U5729 ( .B(n5292), .A(n5293), .Z(n5290) );
  AND U5730 ( .A(b[4]), .B(a[30]), .Z(n5289) );
  XNOR U5731 ( .A(n5294), .B(n5295), .Z(n5119) );
  NANDN U5732 ( .A(n5296), .B(n5297), .Z(n5295) );
  XNOR U5733 ( .A(n5298), .B(n5110), .Z(n5112) );
  XNOR U5734 ( .A(n5299), .B(n5300), .Z(n5110) );
  AND U5735 ( .A(n5301), .B(n5302), .Z(n5299) );
  AND U5736 ( .A(b[3]), .B(a[31]), .Z(n5298) );
  XNOR U5737 ( .A(n5303), .B(n5304), .Z(swire[33]) );
  XOR U5738 ( .A(n5130), .B(n5305), .Z(n5304) );
  XOR U5739 ( .A(n5129), .B(n5303), .Z(n5305) );
  NAND U5740 ( .A(a[33]), .B(b[0]), .Z(n5129) );
  XNOR U5741 ( .A(n5296), .B(n5297), .Z(n5130) );
  XOR U5742 ( .A(n5294), .B(n5306), .Z(n5297) );
  NAND U5743 ( .A(a[32]), .B(b[1]), .Z(n5306) );
  XOR U5744 ( .A(n5302), .B(n5307), .Z(n5296) );
  XOR U5745 ( .A(n5294), .B(n5301), .Z(n5307) );
  XNOR U5746 ( .A(n5308), .B(n5300), .Z(n5301) );
  AND U5747 ( .A(b[2]), .B(a[31]), .Z(n5308) );
  NANDN U5748 ( .A(n5309), .B(n5310), .Z(n5294) );
  XOR U5749 ( .A(n5300), .B(n5292), .Z(n5311) );
  XNOR U5750 ( .A(n5291), .B(n5287), .Z(n5312) );
  XNOR U5751 ( .A(n5286), .B(n5282), .Z(n5313) );
  XNOR U5752 ( .A(n5281), .B(n5277), .Z(n5314) );
  XNOR U5753 ( .A(n5276), .B(n5272), .Z(n5315) );
  XNOR U5754 ( .A(n5271), .B(n5267), .Z(n5316) );
  XNOR U5755 ( .A(n5266), .B(n5262), .Z(n5317) );
  XNOR U5756 ( .A(n5261), .B(n5257), .Z(n5318) );
  XNOR U5757 ( .A(n5256), .B(n5252), .Z(n5319) );
  XNOR U5758 ( .A(n5251), .B(n5247), .Z(n5320) );
  XNOR U5759 ( .A(n5246), .B(n5242), .Z(n5321) );
  XNOR U5760 ( .A(n5241), .B(n5237), .Z(n5322) );
  XNOR U5761 ( .A(n5236), .B(n5232), .Z(n5323) );
  XNOR U5762 ( .A(n5231), .B(n5227), .Z(n5324) );
  XNOR U5763 ( .A(n5226), .B(n5222), .Z(n5325) );
  XNOR U5764 ( .A(n5221), .B(n5217), .Z(n5326) );
  XNOR U5765 ( .A(n5216), .B(n5212), .Z(n5327) );
  XNOR U5766 ( .A(n5211), .B(n5207), .Z(n5328) );
  XNOR U5767 ( .A(n5206), .B(n5202), .Z(n5329) );
  XNOR U5768 ( .A(n5201), .B(n5197), .Z(n5330) );
  XNOR U5769 ( .A(n5196), .B(n5192), .Z(n5331) );
  XNOR U5770 ( .A(n5191), .B(n5187), .Z(n5332) );
  XNOR U5771 ( .A(n5186), .B(n5182), .Z(n5333) );
  XNOR U5772 ( .A(n5181), .B(n5177), .Z(n5334) );
  XNOR U5773 ( .A(n5176), .B(n5172), .Z(n5335) );
  XOR U5774 ( .A(n5171), .B(n5168), .Z(n5336) );
  XOR U5775 ( .A(n5337), .B(n5338), .Z(n5168) );
  XOR U5776 ( .A(n5166), .B(n5339), .Z(n5338) );
  XOR U5777 ( .A(n5340), .B(n5341), .Z(n5339) );
  XOR U5778 ( .A(n5342), .B(n5343), .Z(n5341) );
  NAND U5779 ( .A(a[3]), .B(b[30]), .Z(n5343) );
  AND U5780 ( .A(a[2]), .B(b[31]), .Z(n5342) );
  XOR U5781 ( .A(n5344), .B(n5340), .Z(n5337) );
  XOR U5782 ( .A(n5345), .B(n5346), .Z(n5340) );
  NOR U5783 ( .A(n5347), .B(n5348), .Z(n5345) );
  AND U5784 ( .A(a[4]), .B(b[29]), .Z(n5344) );
  XNOR U5785 ( .A(n5349), .B(n5166), .Z(n5167) );
  XOR U5786 ( .A(n5350), .B(n5351), .Z(n5166) );
  ANDN U5787 ( .B(n5352), .A(n5353), .Z(n5350) );
  AND U5788 ( .A(a[5]), .B(b[28]), .Z(n5349) );
  XNOR U5789 ( .A(n5354), .B(n5171), .Z(n5173) );
  XOR U5790 ( .A(n5355), .B(n5356), .Z(n5171) );
  ANDN U5791 ( .B(n5357), .A(n5358), .Z(n5355) );
  AND U5792 ( .A(a[6]), .B(b[27]), .Z(n5354) );
  XNOR U5793 ( .A(n5359), .B(n5176), .Z(n5178) );
  XOR U5794 ( .A(n5360), .B(n5361), .Z(n5176) );
  ANDN U5795 ( .B(n5362), .A(n5363), .Z(n5360) );
  AND U5796 ( .A(a[7]), .B(b[26]), .Z(n5359) );
  XNOR U5797 ( .A(n5364), .B(n5181), .Z(n5183) );
  XOR U5798 ( .A(n5365), .B(n5366), .Z(n5181) );
  ANDN U5799 ( .B(n5367), .A(n5368), .Z(n5365) );
  AND U5800 ( .A(a[8]), .B(b[25]), .Z(n5364) );
  XNOR U5801 ( .A(n5369), .B(n5186), .Z(n5188) );
  XOR U5802 ( .A(n5370), .B(n5371), .Z(n5186) );
  ANDN U5803 ( .B(n5372), .A(n5373), .Z(n5370) );
  AND U5804 ( .A(a[9]), .B(b[24]), .Z(n5369) );
  XNOR U5805 ( .A(n5374), .B(n5191), .Z(n5193) );
  XOR U5806 ( .A(n5375), .B(n5376), .Z(n5191) );
  ANDN U5807 ( .B(n5377), .A(n5378), .Z(n5375) );
  AND U5808 ( .A(a[10]), .B(b[23]), .Z(n5374) );
  XNOR U5809 ( .A(n5379), .B(n5196), .Z(n5198) );
  XOR U5810 ( .A(n5380), .B(n5381), .Z(n5196) );
  ANDN U5811 ( .B(n5382), .A(n5383), .Z(n5380) );
  AND U5812 ( .A(a[11]), .B(b[22]), .Z(n5379) );
  XNOR U5813 ( .A(n5384), .B(n5201), .Z(n5203) );
  XOR U5814 ( .A(n5385), .B(n5386), .Z(n5201) );
  ANDN U5815 ( .B(n5387), .A(n5388), .Z(n5385) );
  AND U5816 ( .A(a[12]), .B(b[21]), .Z(n5384) );
  XNOR U5817 ( .A(n5389), .B(n5206), .Z(n5208) );
  XOR U5818 ( .A(n5390), .B(n5391), .Z(n5206) );
  ANDN U5819 ( .B(n5392), .A(n5393), .Z(n5390) );
  AND U5820 ( .A(a[13]), .B(b[20]), .Z(n5389) );
  XNOR U5821 ( .A(n5394), .B(n5211), .Z(n5213) );
  XOR U5822 ( .A(n5395), .B(n5396), .Z(n5211) );
  ANDN U5823 ( .B(n5397), .A(n5398), .Z(n5395) );
  AND U5824 ( .A(a[14]), .B(b[19]), .Z(n5394) );
  XNOR U5825 ( .A(n5399), .B(n5216), .Z(n5218) );
  XOR U5826 ( .A(n5400), .B(n5401), .Z(n5216) );
  ANDN U5827 ( .B(n5402), .A(n5403), .Z(n5400) );
  AND U5828 ( .A(a[15]), .B(b[18]), .Z(n5399) );
  XNOR U5829 ( .A(n5404), .B(n5221), .Z(n5223) );
  XOR U5830 ( .A(n5405), .B(n5406), .Z(n5221) );
  ANDN U5831 ( .B(n5407), .A(n5408), .Z(n5405) );
  AND U5832 ( .A(a[16]), .B(b[17]), .Z(n5404) );
  XNOR U5833 ( .A(n5409), .B(n5226), .Z(n5228) );
  XOR U5834 ( .A(n5410), .B(n5411), .Z(n5226) );
  ANDN U5835 ( .B(n5412), .A(n5413), .Z(n5410) );
  AND U5836 ( .A(b[16]), .B(a[17]), .Z(n5409) );
  XNOR U5837 ( .A(n5414), .B(n5231), .Z(n5233) );
  XOR U5838 ( .A(n5415), .B(n5416), .Z(n5231) );
  ANDN U5839 ( .B(n5417), .A(n5418), .Z(n5415) );
  AND U5840 ( .A(a[18]), .B(b[15]), .Z(n5414) );
  XNOR U5841 ( .A(n5419), .B(n5236), .Z(n5238) );
  XOR U5842 ( .A(n5420), .B(n5421), .Z(n5236) );
  ANDN U5843 ( .B(n5422), .A(n5423), .Z(n5420) );
  AND U5844 ( .A(b[14]), .B(a[19]), .Z(n5419) );
  XNOR U5845 ( .A(n5424), .B(n5241), .Z(n5243) );
  XOR U5846 ( .A(n5425), .B(n5426), .Z(n5241) );
  ANDN U5847 ( .B(n5427), .A(n5428), .Z(n5425) );
  AND U5848 ( .A(a[20]), .B(b[13]), .Z(n5424) );
  XNOR U5849 ( .A(n5429), .B(n5246), .Z(n5248) );
  XOR U5850 ( .A(n5430), .B(n5431), .Z(n5246) );
  ANDN U5851 ( .B(n5432), .A(n5433), .Z(n5430) );
  AND U5852 ( .A(b[12]), .B(a[21]), .Z(n5429) );
  XNOR U5853 ( .A(n5434), .B(n5251), .Z(n5253) );
  XOR U5854 ( .A(n5435), .B(n5436), .Z(n5251) );
  ANDN U5855 ( .B(n5437), .A(n5438), .Z(n5435) );
  AND U5856 ( .A(a[22]), .B(b[11]), .Z(n5434) );
  XNOR U5857 ( .A(n5439), .B(n5256), .Z(n5258) );
  XOR U5858 ( .A(n5440), .B(n5441), .Z(n5256) );
  ANDN U5859 ( .B(n5442), .A(n5443), .Z(n5440) );
  AND U5860 ( .A(b[10]), .B(a[23]), .Z(n5439) );
  XNOR U5861 ( .A(n5444), .B(n5261), .Z(n5263) );
  XOR U5862 ( .A(n5445), .B(n5446), .Z(n5261) );
  ANDN U5863 ( .B(n5447), .A(n5448), .Z(n5445) );
  AND U5864 ( .A(a[24]), .B(b[9]), .Z(n5444) );
  XNOR U5865 ( .A(n5449), .B(n5266), .Z(n5268) );
  XOR U5866 ( .A(n5450), .B(n5451), .Z(n5266) );
  ANDN U5867 ( .B(n5452), .A(n5453), .Z(n5450) );
  AND U5868 ( .A(b[8]), .B(a[25]), .Z(n5449) );
  XNOR U5869 ( .A(n5454), .B(n5271), .Z(n5273) );
  XOR U5870 ( .A(n5455), .B(n5456), .Z(n5271) );
  ANDN U5871 ( .B(n5457), .A(n5458), .Z(n5455) );
  AND U5872 ( .A(a[26]), .B(b[7]), .Z(n5454) );
  XNOR U5873 ( .A(n5459), .B(n5276), .Z(n5278) );
  XOR U5874 ( .A(n5460), .B(n5461), .Z(n5276) );
  ANDN U5875 ( .B(n5462), .A(n5463), .Z(n5460) );
  AND U5876 ( .A(b[6]), .B(a[27]), .Z(n5459) );
  XNOR U5877 ( .A(n5464), .B(n5281), .Z(n5283) );
  XOR U5878 ( .A(n5465), .B(n5466), .Z(n5281) );
  ANDN U5879 ( .B(n5467), .A(n5468), .Z(n5465) );
  AND U5880 ( .A(b[5]), .B(a[28]), .Z(n5464) );
  XNOR U5881 ( .A(n5469), .B(n5286), .Z(n5288) );
  XOR U5882 ( .A(n5470), .B(n5471), .Z(n5286) );
  ANDN U5883 ( .B(n5472), .A(n5473), .Z(n5470) );
  AND U5884 ( .A(b[4]), .B(a[29]), .Z(n5469) );
  XNOR U5885 ( .A(n5474), .B(n5475), .Z(n5300) );
  NANDN U5886 ( .A(n5476), .B(n5477), .Z(n5475) );
  XNOR U5887 ( .A(n5478), .B(n5291), .Z(n5293) );
  XNOR U5888 ( .A(n5479), .B(n5480), .Z(n5291) );
  AND U5889 ( .A(n5481), .B(n5482), .Z(n5479) );
  AND U5890 ( .A(b[3]), .B(a[30]), .Z(n5478) );
  XOR U5891 ( .A(n5483), .B(n5485), .Z(swire[32]) );
  XNOR U5892 ( .A(n5483), .B(n5486), .Z(n5485) );
  XOR U5893 ( .A(n5309), .B(n5310), .Z(n5486) );
  XNOR U5894 ( .A(n5476), .B(n5477), .Z(n5310) );
  XOR U5895 ( .A(n5474), .B(n5487), .Z(n5477) );
  NAND U5896 ( .A(b[1]), .B(a[31]), .Z(n5487) );
  XOR U5897 ( .A(n5482), .B(n5488), .Z(n5476) );
  XOR U5898 ( .A(n5474), .B(n5481), .Z(n5488) );
  XNOR U5899 ( .A(n5489), .B(n5480), .Z(n5481) );
  AND U5900 ( .A(b[2]), .B(a[30]), .Z(n5489) );
  NANDN U5901 ( .A(n5490), .B(n5491), .Z(n5474) );
  XOR U5902 ( .A(n5480), .B(n5472), .Z(n5492) );
  XNOR U5903 ( .A(n5471), .B(n5467), .Z(n5493) );
  XNOR U5904 ( .A(n5466), .B(n5462), .Z(n5494) );
  XNOR U5905 ( .A(n5461), .B(n5457), .Z(n5495) );
  XNOR U5906 ( .A(n5456), .B(n5452), .Z(n5496) );
  XNOR U5907 ( .A(n5451), .B(n5447), .Z(n5497) );
  XNOR U5908 ( .A(n5446), .B(n5442), .Z(n5498) );
  XNOR U5909 ( .A(n5441), .B(n5437), .Z(n5499) );
  XNOR U5910 ( .A(n5436), .B(n5432), .Z(n5500) );
  XNOR U5911 ( .A(n5431), .B(n5427), .Z(n5501) );
  XNOR U5912 ( .A(n5426), .B(n5422), .Z(n5502) );
  XNOR U5913 ( .A(n5421), .B(n5417), .Z(n5503) );
  XNOR U5914 ( .A(n5416), .B(n5412), .Z(n5504) );
  XNOR U5915 ( .A(n5411), .B(n5407), .Z(n5505) );
  XNOR U5916 ( .A(n5406), .B(n5402), .Z(n5506) );
  XNOR U5917 ( .A(n5401), .B(n5397), .Z(n5507) );
  XNOR U5918 ( .A(n5396), .B(n5392), .Z(n5508) );
  XNOR U5919 ( .A(n5391), .B(n5387), .Z(n5509) );
  XNOR U5920 ( .A(n5386), .B(n5382), .Z(n5510) );
  XNOR U5921 ( .A(n5381), .B(n5377), .Z(n5511) );
  XNOR U5922 ( .A(n5376), .B(n5372), .Z(n5512) );
  XNOR U5923 ( .A(n5371), .B(n5367), .Z(n5513) );
  XNOR U5924 ( .A(n5366), .B(n5362), .Z(n5514) );
  XNOR U5925 ( .A(n5361), .B(n5357), .Z(n5515) );
  XNOR U5926 ( .A(n5356), .B(n5352), .Z(n5516) );
  XOR U5927 ( .A(n5351), .B(n5348), .Z(n5517) );
  XOR U5928 ( .A(n5518), .B(n5519), .Z(n5348) );
  XOR U5929 ( .A(n5346), .B(n5520), .Z(n5519) );
  XOR U5930 ( .A(n5521), .B(n5522), .Z(n5520) );
  XOR U5931 ( .A(n5523), .B(n5524), .Z(n5522) );
  NAND U5932 ( .A(a[2]), .B(b[30]), .Z(n5524) );
  AND U5933 ( .A(a[1]), .B(b[31]), .Z(n5523) );
  XOR U5934 ( .A(n5525), .B(n5521), .Z(n5518) );
  XOR U5935 ( .A(n5526), .B(n5527), .Z(n5521) );
  NOR U5936 ( .A(n5528), .B(n5529), .Z(n5526) );
  AND U5937 ( .A(a[3]), .B(b[29]), .Z(n5525) );
  XNOR U5938 ( .A(n5530), .B(n5346), .Z(n5347) );
  XOR U5939 ( .A(n5531), .B(n5532), .Z(n5346) );
  ANDN U5940 ( .B(n5533), .A(n5534), .Z(n5531) );
  AND U5941 ( .A(a[4]), .B(b[28]), .Z(n5530) );
  XNOR U5942 ( .A(n5535), .B(n5351), .Z(n5353) );
  XOR U5943 ( .A(n5536), .B(n5537), .Z(n5351) );
  ANDN U5944 ( .B(n5538), .A(n5539), .Z(n5536) );
  AND U5945 ( .A(a[5]), .B(b[27]), .Z(n5535) );
  XNOR U5946 ( .A(n5540), .B(n5356), .Z(n5358) );
  XOR U5947 ( .A(n5541), .B(n5542), .Z(n5356) );
  ANDN U5948 ( .B(n5543), .A(n5544), .Z(n5541) );
  AND U5949 ( .A(a[6]), .B(b[26]), .Z(n5540) );
  XNOR U5950 ( .A(n5545), .B(n5361), .Z(n5363) );
  XOR U5951 ( .A(n5546), .B(n5547), .Z(n5361) );
  ANDN U5952 ( .B(n5548), .A(n5549), .Z(n5546) );
  AND U5953 ( .A(a[7]), .B(b[25]), .Z(n5545) );
  XNOR U5954 ( .A(n5550), .B(n5366), .Z(n5368) );
  XOR U5955 ( .A(n5551), .B(n5552), .Z(n5366) );
  ANDN U5956 ( .B(n5553), .A(n5554), .Z(n5551) );
  AND U5957 ( .A(a[8]), .B(b[24]), .Z(n5550) );
  XNOR U5958 ( .A(n5555), .B(n5371), .Z(n5373) );
  XOR U5959 ( .A(n5556), .B(n5557), .Z(n5371) );
  ANDN U5960 ( .B(n5558), .A(n5559), .Z(n5556) );
  AND U5961 ( .A(a[9]), .B(b[23]), .Z(n5555) );
  XNOR U5962 ( .A(n5560), .B(n5376), .Z(n5378) );
  XOR U5963 ( .A(n5561), .B(n5562), .Z(n5376) );
  ANDN U5964 ( .B(n5563), .A(n5564), .Z(n5561) );
  AND U5965 ( .A(a[10]), .B(b[22]), .Z(n5560) );
  XNOR U5966 ( .A(n5565), .B(n5381), .Z(n5383) );
  XOR U5967 ( .A(n5566), .B(n5567), .Z(n5381) );
  ANDN U5968 ( .B(n5568), .A(n5569), .Z(n5566) );
  AND U5969 ( .A(a[11]), .B(b[21]), .Z(n5565) );
  XNOR U5970 ( .A(n5570), .B(n5386), .Z(n5388) );
  XOR U5971 ( .A(n5571), .B(n5572), .Z(n5386) );
  ANDN U5972 ( .B(n5573), .A(n5574), .Z(n5571) );
  AND U5973 ( .A(a[12]), .B(b[20]), .Z(n5570) );
  XNOR U5974 ( .A(n5575), .B(n5391), .Z(n5393) );
  XOR U5975 ( .A(n5576), .B(n5577), .Z(n5391) );
  ANDN U5976 ( .B(n5578), .A(n5579), .Z(n5576) );
  AND U5977 ( .A(a[13]), .B(b[19]), .Z(n5575) );
  XNOR U5978 ( .A(n5580), .B(n5396), .Z(n5398) );
  XOR U5979 ( .A(n5581), .B(n5582), .Z(n5396) );
  ANDN U5980 ( .B(n5583), .A(n5584), .Z(n5581) );
  AND U5981 ( .A(a[14]), .B(b[18]), .Z(n5580) );
  XNOR U5982 ( .A(n5585), .B(n5401), .Z(n5403) );
  XOR U5983 ( .A(n5586), .B(n5587), .Z(n5401) );
  ANDN U5984 ( .B(n5588), .A(n5589), .Z(n5586) );
  AND U5985 ( .A(a[15]), .B(b[17]), .Z(n5585) );
  XNOR U5986 ( .A(n5590), .B(n5406), .Z(n5408) );
  XOR U5987 ( .A(n5591), .B(n5592), .Z(n5406) );
  ANDN U5988 ( .B(n5593), .A(n5594), .Z(n5591) );
  AND U5989 ( .A(a[16]), .B(b[16]), .Z(n5590) );
  XNOR U5990 ( .A(n5595), .B(n5411), .Z(n5413) );
  XOR U5991 ( .A(n5596), .B(n5597), .Z(n5411) );
  ANDN U5992 ( .B(n5598), .A(n5599), .Z(n5596) );
  AND U5993 ( .A(b[15]), .B(a[17]), .Z(n5595) );
  XNOR U5994 ( .A(n5600), .B(n5416), .Z(n5418) );
  XOR U5995 ( .A(n5601), .B(n5602), .Z(n5416) );
  ANDN U5996 ( .B(n5603), .A(n5604), .Z(n5601) );
  AND U5997 ( .A(a[18]), .B(b[14]), .Z(n5600) );
  XNOR U5998 ( .A(n5605), .B(n5421), .Z(n5423) );
  XOR U5999 ( .A(n5606), .B(n5607), .Z(n5421) );
  ANDN U6000 ( .B(n5608), .A(n5609), .Z(n5606) );
  AND U6001 ( .A(b[13]), .B(a[19]), .Z(n5605) );
  XNOR U6002 ( .A(n5610), .B(n5426), .Z(n5428) );
  XOR U6003 ( .A(n5611), .B(n5612), .Z(n5426) );
  ANDN U6004 ( .B(n5613), .A(n5614), .Z(n5611) );
  AND U6005 ( .A(a[20]), .B(b[12]), .Z(n5610) );
  XNOR U6006 ( .A(n5615), .B(n5431), .Z(n5433) );
  XOR U6007 ( .A(n5616), .B(n5617), .Z(n5431) );
  ANDN U6008 ( .B(n5618), .A(n5619), .Z(n5616) );
  AND U6009 ( .A(b[11]), .B(a[21]), .Z(n5615) );
  XNOR U6010 ( .A(n5620), .B(n5436), .Z(n5438) );
  XOR U6011 ( .A(n5621), .B(n5622), .Z(n5436) );
  ANDN U6012 ( .B(n5623), .A(n5624), .Z(n5621) );
  AND U6013 ( .A(a[22]), .B(b[10]), .Z(n5620) );
  XNOR U6014 ( .A(n5625), .B(n5441), .Z(n5443) );
  XOR U6015 ( .A(n5626), .B(n5627), .Z(n5441) );
  ANDN U6016 ( .B(n5628), .A(n5629), .Z(n5626) );
  AND U6017 ( .A(b[9]), .B(a[23]), .Z(n5625) );
  XNOR U6018 ( .A(n5630), .B(n5446), .Z(n5448) );
  XOR U6019 ( .A(n5631), .B(n5632), .Z(n5446) );
  ANDN U6020 ( .B(n5633), .A(n5634), .Z(n5631) );
  AND U6021 ( .A(a[24]), .B(b[8]), .Z(n5630) );
  XNOR U6022 ( .A(n5635), .B(n5451), .Z(n5453) );
  XOR U6023 ( .A(n5636), .B(n5637), .Z(n5451) );
  ANDN U6024 ( .B(n5638), .A(n5639), .Z(n5636) );
  AND U6025 ( .A(b[7]), .B(a[25]), .Z(n5635) );
  XNOR U6026 ( .A(n5640), .B(n5456), .Z(n5458) );
  XOR U6027 ( .A(n5641), .B(n5642), .Z(n5456) );
  ANDN U6028 ( .B(n5643), .A(n5644), .Z(n5641) );
  AND U6029 ( .A(b[6]), .B(a[26]), .Z(n5640) );
  XNOR U6030 ( .A(n5645), .B(n5461), .Z(n5463) );
  XOR U6031 ( .A(n5646), .B(n5647), .Z(n5461) );
  ANDN U6032 ( .B(n5648), .A(n5649), .Z(n5646) );
  AND U6033 ( .A(b[5]), .B(a[27]), .Z(n5645) );
  XNOR U6034 ( .A(n5650), .B(n5466), .Z(n5468) );
  XOR U6035 ( .A(n5651), .B(n5652), .Z(n5466) );
  ANDN U6036 ( .B(n5653), .A(n5654), .Z(n5651) );
  AND U6037 ( .A(b[4]), .B(a[28]), .Z(n5650) );
  XNOR U6038 ( .A(n5655), .B(n5656), .Z(n5480) );
  NANDN U6039 ( .A(n5657), .B(n5658), .Z(n5656) );
  XNOR U6040 ( .A(n5659), .B(n5471), .Z(n5473) );
  XNOR U6041 ( .A(n5660), .B(n5661), .Z(n5471) );
  AND U6042 ( .A(n5662), .B(n5663), .Z(n5660) );
  AND U6043 ( .A(b[3]), .B(a[29]), .Z(n5659) );
  NAND U6044 ( .A(a[32]), .B(b[0]), .Z(n5309) );
  IV U6045 ( .A(n5484), .Z(n5483) );
  XOR U6046 ( .A(n5664), .B(n5665), .Z(n5484) );
  ANDN U6047 ( .B(n5666), .A(n5667), .Z(n5664) );
  XNOR U6048 ( .A(n5666), .B(n5667), .Z(c[63]) );
  XNOR U6049 ( .A(sreg[95]), .B(n5668), .Z(n5667) );
  XNOR U6050 ( .A(n5668), .B(n5669), .Z(n5666) );
  XOR U6051 ( .A(n5490), .B(n5491), .Z(n5669) );
  XNOR U6052 ( .A(n5657), .B(n5658), .Z(n5491) );
  XOR U6053 ( .A(n5655), .B(n5670), .Z(n5658) );
  NAND U6054 ( .A(a[30]), .B(b[1]), .Z(n5670) );
  XOR U6055 ( .A(n5663), .B(n5671), .Z(n5657) );
  XOR U6056 ( .A(n5655), .B(n5662), .Z(n5671) );
  XNOR U6057 ( .A(n5672), .B(n5661), .Z(n5662) );
  AND U6058 ( .A(b[2]), .B(a[29]), .Z(n5672) );
  NANDN U6059 ( .A(n5673), .B(n5674), .Z(n5655) );
  XOR U6060 ( .A(n5661), .B(n5653), .Z(n5675) );
  XNOR U6061 ( .A(n5652), .B(n5648), .Z(n5676) );
  XNOR U6062 ( .A(n5647), .B(n5643), .Z(n5677) );
  XNOR U6063 ( .A(n5642), .B(n5638), .Z(n5678) );
  XNOR U6064 ( .A(n5637), .B(n5633), .Z(n5679) );
  XNOR U6065 ( .A(n5632), .B(n5628), .Z(n5680) );
  XNOR U6066 ( .A(n5627), .B(n5623), .Z(n5681) );
  XNOR U6067 ( .A(n5622), .B(n5618), .Z(n5682) );
  XNOR U6068 ( .A(n5617), .B(n5613), .Z(n5683) );
  XNOR U6069 ( .A(n5612), .B(n5608), .Z(n5684) );
  XNOR U6070 ( .A(n5607), .B(n5603), .Z(n5685) );
  XNOR U6071 ( .A(n5602), .B(n5598), .Z(n5686) );
  XNOR U6072 ( .A(n5597), .B(n5593), .Z(n5687) );
  XNOR U6073 ( .A(n5592), .B(n5588), .Z(n5688) );
  XNOR U6074 ( .A(n5587), .B(n5583), .Z(n5689) );
  XNOR U6075 ( .A(n5582), .B(n5578), .Z(n5690) );
  XNOR U6076 ( .A(n5577), .B(n5573), .Z(n5691) );
  XNOR U6077 ( .A(n5572), .B(n5568), .Z(n5692) );
  XNOR U6078 ( .A(n5567), .B(n5563), .Z(n5693) );
  XNOR U6079 ( .A(n5562), .B(n5558), .Z(n5694) );
  XNOR U6080 ( .A(n5557), .B(n5553), .Z(n5695) );
  XNOR U6081 ( .A(n5552), .B(n5548), .Z(n5696) );
  XNOR U6082 ( .A(n5547), .B(n5543), .Z(n5697) );
  XNOR U6083 ( .A(n5542), .B(n5538), .Z(n5698) );
  XNOR U6084 ( .A(n5537), .B(n5533), .Z(n5699) );
  XOR U6085 ( .A(n5532), .B(n5529), .Z(n5700) );
  XOR U6086 ( .A(n5701), .B(n5702), .Z(n5529) );
  XOR U6087 ( .A(n5527), .B(n5703), .Z(n5702) );
  XOR U6088 ( .A(n5704), .B(n5705), .Z(n5703) );
  XOR U6089 ( .A(n5706), .B(n5707), .Z(n5705) );
  NAND U6090 ( .A(a[1]), .B(b[30]), .Z(n5707) );
  AND U6091 ( .A(a[0]), .B(b[31]), .Z(n5706) );
  XOR U6092 ( .A(n5708), .B(n5704), .Z(n5701) );
  XOR U6093 ( .A(n5709), .B(n5710), .Z(n5704) );
  NOR U6094 ( .A(n5711), .B(n5712), .Z(n5709) );
  AND U6095 ( .A(a[2]), .B(b[29]), .Z(n5708) );
  XNOR U6096 ( .A(n5713), .B(n5527), .Z(n5528) );
  XOR U6097 ( .A(n5714), .B(n5715), .Z(n5527) );
  ANDN U6098 ( .B(n5716), .A(n5717), .Z(n5714) );
  AND U6099 ( .A(a[3]), .B(b[28]), .Z(n5713) );
  XNOR U6100 ( .A(n5718), .B(n5532), .Z(n5534) );
  XOR U6101 ( .A(n5719), .B(n5720), .Z(n5532) );
  ANDN U6102 ( .B(n5721), .A(n5722), .Z(n5719) );
  AND U6103 ( .A(a[4]), .B(b[27]), .Z(n5718) );
  XNOR U6104 ( .A(n5723), .B(n5537), .Z(n5539) );
  XOR U6105 ( .A(n5724), .B(n5725), .Z(n5537) );
  ANDN U6106 ( .B(n5726), .A(n5727), .Z(n5724) );
  AND U6107 ( .A(a[5]), .B(b[26]), .Z(n5723) );
  XNOR U6108 ( .A(n5728), .B(n5542), .Z(n5544) );
  XOR U6109 ( .A(n5729), .B(n5730), .Z(n5542) );
  ANDN U6110 ( .B(n5731), .A(n5732), .Z(n5729) );
  AND U6111 ( .A(a[6]), .B(b[25]), .Z(n5728) );
  XNOR U6112 ( .A(n5733), .B(n5547), .Z(n5549) );
  XOR U6113 ( .A(n5734), .B(n5735), .Z(n5547) );
  ANDN U6114 ( .B(n5736), .A(n5737), .Z(n5734) );
  AND U6115 ( .A(a[7]), .B(b[24]), .Z(n5733) );
  XNOR U6116 ( .A(n5738), .B(n5552), .Z(n5554) );
  XOR U6117 ( .A(n5739), .B(n5740), .Z(n5552) );
  ANDN U6118 ( .B(n5741), .A(n5742), .Z(n5739) );
  AND U6119 ( .A(a[8]), .B(b[23]), .Z(n5738) );
  XNOR U6120 ( .A(n5743), .B(n5557), .Z(n5559) );
  XOR U6121 ( .A(n5744), .B(n5745), .Z(n5557) );
  ANDN U6122 ( .B(n5746), .A(n5747), .Z(n5744) );
  AND U6123 ( .A(a[9]), .B(b[22]), .Z(n5743) );
  XNOR U6124 ( .A(n5748), .B(n5562), .Z(n5564) );
  XOR U6125 ( .A(n5749), .B(n5750), .Z(n5562) );
  ANDN U6126 ( .B(n5751), .A(n5752), .Z(n5749) );
  AND U6127 ( .A(a[10]), .B(b[21]), .Z(n5748) );
  XNOR U6128 ( .A(n5753), .B(n5567), .Z(n5569) );
  XOR U6129 ( .A(n5754), .B(n5755), .Z(n5567) );
  ANDN U6130 ( .B(n5756), .A(n5757), .Z(n5754) );
  AND U6131 ( .A(a[11]), .B(b[20]), .Z(n5753) );
  XNOR U6132 ( .A(n5758), .B(n5572), .Z(n5574) );
  XOR U6133 ( .A(n5759), .B(n5760), .Z(n5572) );
  ANDN U6134 ( .B(n5761), .A(n5762), .Z(n5759) );
  AND U6135 ( .A(a[12]), .B(b[19]), .Z(n5758) );
  XNOR U6136 ( .A(n5763), .B(n5577), .Z(n5579) );
  XOR U6137 ( .A(n5764), .B(n5765), .Z(n5577) );
  ANDN U6138 ( .B(n5766), .A(n5767), .Z(n5764) );
  AND U6139 ( .A(a[13]), .B(b[18]), .Z(n5763) );
  XNOR U6140 ( .A(n5768), .B(n5582), .Z(n5584) );
  XOR U6141 ( .A(n5769), .B(n5770), .Z(n5582) );
  ANDN U6142 ( .B(n5771), .A(n5772), .Z(n5769) );
  AND U6143 ( .A(a[14]), .B(b[17]), .Z(n5768) );
  XNOR U6144 ( .A(n5773), .B(n5587), .Z(n5589) );
  XOR U6145 ( .A(n5774), .B(n5775), .Z(n5587) );
  ANDN U6146 ( .B(n5776), .A(n5777), .Z(n5774) );
  AND U6147 ( .A(a[15]), .B(b[16]), .Z(n5773) );
  XNOR U6148 ( .A(n5778), .B(n5592), .Z(n5594) );
  XOR U6149 ( .A(n5779), .B(n5780), .Z(n5592) );
  ANDN U6150 ( .B(n5781), .A(n5782), .Z(n5779) );
  AND U6151 ( .A(a[16]), .B(b[15]), .Z(n5778) );
  XNOR U6152 ( .A(n5783), .B(n5597), .Z(n5599) );
  XOR U6153 ( .A(n5784), .B(n5785), .Z(n5597) );
  ANDN U6154 ( .B(n5786), .A(n5787), .Z(n5784) );
  AND U6155 ( .A(b[14]), .B(a[17]), .Z(n5783) );
  XNOR U6156 ( .A(n5788), .B(n5602), .Z(n5604) );
  XOR U6157 ( .A(n5789), .B(n5790), .Z(n5602) );
  ANDN U6158 ( .B(n5791), .A(n5792), .Z(n5789) );
  AND U6159 ( .A(a[18]), .B(b[13]), .Z(n5788) );
  XNOR U6160 ( .A(n5793), .B(n5607), .Z(n5609) );
  XOR U6161 ( .A(n5794), .B(n5795), .Z(n5607) );
  ANDN U6162 ( .B(n5796), .A(n5797), .Z(n5794) );
  AND U6163 ( .A(b[12]), .B(a[19]), .Z(n5793) );
  XNOR U6164 ( .A(n5798), .B(n5612), .Z(n5614) );
  XOR U6165 ( .A(n5799), .B(n5800), .Z(n5612) );
  ANDN U6166 ( .B(n5801), .A(n5802), .Z(n5799) );
  AND U6167 ( .A(a[20]), .B(b[11]), .Z(n5798) );
  XNOR U6168 ( .A(n5803), .B(n5617), .Z(n5619) );
  XOR U6169 ( .A(n5804), .B(n5805), .Z(n5617) );
  ANDN U6170 ( .B(n5806), .A(n5807), .Z(n5804) );
  AND U6171 ( .A(b[10]), .B(a[21]), .Z(n5803) );
  XNOR U6172 ( .A(n5808), .B(n5622), .Z(n5624) );
  XOR U6173 ( .A(n5809), .B(n5810), .Z(n5622) );
  ANDN U6174 ( .B(n5811), .A(n5812), .Z(n5809) );
  AND U6175 ( .A(a[22]), .B(b[9]), .Z(n5808) );
  XNOR U6176 ( .A(n5813), .B(n5627), .Z(n5629) );
  XOR U6177 ( .A(n5814), .B(n5815), .Z(n5627) );
  ANDN U6178 ( .B(n5816), .A(n5817), .Z(n5814) );
  AND U6179 ( .A(b[8]), .B(a[23]), .Z(n5813) );
  XNOR U6180 ( .A(n5818), .B(n5632), .Z(n5634) );
  XOR U6181 ( .A(n5819), .B(n5820), .Z(n5632) );
  ANDN U6182 ( .B(n5821), .A(n5822), .Z(n5819) );
  AND U6183 ( .A(a[24]), .B(b[7]), .Z(n5818) );
  XNOR U6184 ( .A(n5823), .B(n5637), .Z(n5639) );
  XOR U6185 ( .A(n5824), .B(n5825), .Z(n5637) );
  ANDN U6186 ( .B(n5826), .A(n5827), .Z(n5824) );
  AND U6187 ( .A(b[6]), .B(a[25]), .Z(n5823) );
  XNOR U6188 ( .A(n5828), .B(n5642), .Z(n5644) );
  XOR U6189 ( .A(n5829), .B(n5830), .Z(n5642) );
  ANDN U6190 ( .B(n5831), .A(n5832), .Z(n5829) );
  AND U6191 ( .A(b[5]), .B(a[26]), .Z(n5828) );
  XNOR U6192 ( .A(n5833), .B(n5647), .Z(n5649) );
  XOR U6193 ( .A(n5834), .B(n5835), .Z(n5647) );
  ANDN U6194 ( .B(n5836), .A(n5837), .Z(n5834) );
  AND U6195 ( .A(b[4]), .B(a[27]), .Z(n5833) );
  XNOR U6196 ( .A(n5838), .B(n5839), .Z(n5661) );
  NANDN U6197 ( .A(n5840), .B(n5841), .Z(n5839) );
  XNOR U6198 ( .A(n5842), .B(n5652), .Z(n5654) );
  XNOR U6199 ( .A(n5843), .B(n5844), .Z(n5652) );
  AND U6200 ( .A(n5845), .B(n5846), .Z(n5843) );
  AND U6201 ( .A(b[3]), .B(a[28]), .Z(n5842) );
  NAND U6202 ( .A(a[31]), .B(b[0]), .Z(n5490) );
  IV U6203 ( .A(n5665), .Z(n5668) );
  XOR U6204 ( .A(n5847), .B(n5848), .Z(n5665) );
  ANDN U6205 ( .B(n5849), .A(n5850), .Z(n5847) );
  XNOR U6206 ( .A(n5849), .B(n5850), .Z(c[62]) );
  XNOR U6207 ( .A(sreg[94]), .B(n5851), .Z(n5850) );
  XNOR U6208 ( .A(n5851), .B(n5852), .Z(n5849) );
  XOR U6209 ( .A(n5673), .B(n5674), .Z(n5852) );
  XNOR U6210 ( .A(n5840), .B(n5841), .Z(n5674) );
  XOR U6211 ( .A(n5838), .B(n5853), .Z(n5841) );
  NAND U6212 ( .A(b[1]), .B(a[29]), .Z(n5853) );
  XOR U6213 ( .A(n5846), .B(n5854), .Z(n5840) );
  XOR U6214 ( .A(n5838), .B(n5845), .Z(n5854) );
  XNOR U6215 ( .A(n5855), .B(n5844), .Z(n5845) );
  AND U6216 ( .A(b[2]), .B(a[28]), .Z(n5855) );
  NANDN U6217 ( .A(n5856), .B(n5857), .Z(n5838) );
  XOR U6218 ( .A(n5844), .B(n5836), .Z(n5858) );
  XNOR U6219 ( .A(n5835), .B(n5831), .Z(n5859) );
  XNOR U6220 ( .A(n5830), .B(n5826), .Z(n5860) );
  XNOR U6221 ( .A(n5825), .B(n5821), .Z(n5861) );
  XNOR U6222 ( .A(n5820), .B(n5816), .Z(n5862) );
  XNOR U6223 ( .A(n5815), .B(n5811), .Z(n5863) );
  XNOR U6224 ( .A(n5810), .B(n5806), .Z(n5864) );
  XNOR U6225 ( .A(n5805), .B(n5801), .Z(n5865) );
  XNOR U6226 ( .A(n5800), .B(n5796), .Z(n5866) );
  XNOR U6227 ( .A(n5795), .B(n5791), .Z(n5867) );
  XNOR U6228 ( .A(n5790), .B(n5786), .Z(n5868) );
  XNOR U6229 ( .A(n5785), .B(n5781), .Z(n5869) );
  XNOR U6230 ( .A(n5780), .B(n5776), .Z(n5870) );
  XNOR U6231 ( .A(n5775), .B(n5771), .Z(n5871) );
  XNOR U6232 ( .A(n5770), .B(n5766), .Z(n5872) );
  XNOR U6233 ( .A(n5765), .B(n5761), .Z(n5873) );
  XNOR U6234 ( .A(n5760), .B(n5756), .Z(n5874) );
  XNOR U6235 ( .A(n5755), .B(n5751), .Z(n5875) );
  XNOR U6236 ( .A(n5750), .B(n5746), .Z(n5876) );
  XNOR U6237 ( .A(n5745), .B(n5741), .Z(n5877) );
  XNOR U6238 ( .A(n5740), .B(n5736), .Z(n5878) );
  XNOR U6239 ( .A(n5735), .B(n5731), .Z(n5879) );
  XNOR U6240 ( .A(n5730), .B(n5726), .Z(n5880) );
  XNOR U6241 ( .A(n5725), .B(n5721), .Z(n5881) );
  XNOR U6242 ( .A(n5720), .B(n5716), .Z(n5882) );
  XOR U6243 ( .A(n5715), .B(n5712), .Z(n5883) );
  XOR U6244 ( .A(n5884), .B(n5885), .Z(n5712) );
  XOR U6245 ( .A(n5710), .B(n5886), .Z(n5885) );
  XOR U6246 ( .A(n5887), .B(n5888), .Z(n5886) );
  AND U6247 ( .A(a[0]), .B(b[30]), .Z(n5887) );
  XNOR U6248 ( .A(n5889), .B(n5888), .Z(n5884) );
  XNOR U6249 ( .A(n5890), .B(n5891), .Z(n5888) );
  ANDN U6250 ( .B(n5892), .A(n5893), .Z(n5890) );
  AND U6251 ( .A(a[1]), .B(b[29]), .Z(n5889) );
  XNOR U6252 ( .A(n5894), .B(n5710), .Z(n5711) );
  XOR U6253 ( .A(n5895), .B(n5896), .Z(n5710) );
  ANDN U6254 ( .B(n5897), .A(n5898), .Z(n5895) );
  AND U6255 ( .A(a[2]), .B(b[28]), .Z(n5894) );
  XNOR U6256 ( .A(n5899), .B(n5715), .Z(n5717) );
  XOR U6257 ( .A(n5900), .B(n5901), .Z(n5715) );
  ANDN U6258 ( .B(n5902), .A(n5903), .Z(n5900) );
  AND U6259 ( .A(a[3]), .B(b[27]), .Z(n5899) );
  XNOR U6260 ( .A(n5904), .B(n5720), .Z(n5722) );
  XOR U6261 ( .A(n5905), .B(n5906), .Z(n5720) );
  ANDN U6262 ( .B(n5907), .A(n5908), .Z(n5905) );
  AND U6263 ( .A(a[4]), .B(b[26]), .Z(n5904) );
  XNOR U6264 ( .A(n5909), .B(n5725), .Z(n5727) );
  XOR U6265 ( .A(n5910), .B(n5911), .Z(n5725) );
  ANDN U6266 ( .B(n5912), .A(n5913), .Z(n5910) );
  AND U6267 ( .A(a[5]), .B(b[25]), .Z(n5909) );
  XNOR U6268 ( .A(n5914), .B(n5730), .Z(n5732) );
  XOR U6269 ( .A(n5915), .B(n5916), .Z(n5730) );
  ANDN U6270 ( .B(n5917), .A(n5918), .Z(n5915) );
  AND U6271 ( .A(a[6]), .B(b[24]), .Z(n5914) );
  XNOR U6272 ( .A(n5919), .B(n5735), .Z(n5737) );
  XOR U6273 ( .A(n5920), .B(n5921), .Z(n5735) );
  ANDN U6274 ( .B(n5922), .A(n5923), .Z(n5920) );
  AND U6275 ( .A(a[7]), .B(b[23]), .Z(n5919) );
  XNOR U6276 ( .A(n5924), .B(n5740), .Z(n5742) );
  XOR U6277 ( .A(n5925), .B(n5926), .Z(n5740) );
  ANDN U6278 ( .B(n5927), .A(n5928), .Z(n5925) );
  AND U6279 ( .A(a[8]), .B(b[22]), .Z(n5924) );
  XNOR U6280 ( .A(n5929), .B(n5745), .Z(n5747) );
  XOR U6281 ( .A(n5930), .B(n5931), .Z(n5745) );
  ANDN U6282 ( .B(n5932), .A(n5933), .Z(n5930) );
  AND U6283 ( .A(a[9]), .B(b[21]), .Z(n5929) );
  XNOR U6284 ( .A(n5934), .B(n5750), .Z(n5752) );
  XOR U6285 ( .A(n5935), .B(n5936), .Z(n5750) );
  ANDN U6286 ( .B(n5937), .A(n5938), .Z(n5935) );
  AND U6287 ( .A(a[10]), .B(b[20]), .Z(n5934) );
  XNOR U6288 ( .A(n5939), .B(n5755), .Z(n5757) );
  XOR U6289 ( .A(n5940), .B(n5941), .Z(n5755) );
  ANDN U6290 ( .B(n5942), .A(n5943), .Z(n5940) );
  AND U6291 ( .A(a[11]), .B(b[19]), .Z(n5939) );
  XNOR U6292 ( .A(n5944), .B(n5760), .Z(n5762) );
  XOR U6293 ( .A(n5945), .B(n5946), .Z(n5760) );
  ANDN U6294 ( .B(n5947), .A(n5948), .Z(n5945) );
  AND U6295 ( .A(a[12]), .B(b[18]), .Z(n5944) );
  XNOR U6296 ( .A(n5949), .B(n5765), .Z(n5767) );
  XOR U6297 ( .A(n5950), .B(n5951), .Z(n5765) );
  ANDN U6298 ( .B(n5952), .A(n5953), .Z(n5950) );
  AND U6299 ( .A(a[13]), .B(b[17]), .Z(n5949) );
  XNOR U6300 ( .A(n5954), .B(n5770), .Z(n5772) );
  XOR U6301 ( .A(n5955), .B(n5956), .Z(n5770) );
  ANDN U6302 ( .B(n5957), .A(n5958), .Z(n5955) );
  AND U6303 ( .A(a[14]), .B(b[16]), .Z(n5954) );
  XNOR U6304 ( .A(n5959), .B(n5775), .Z(n5777) );
  XOR U6305 ( .A(n5960), .B(n5961), .Z(n5775) );
  ANDN U6306 ( .B(n5962), .A(n5963), .Z(n5960) );
  AND U6307 ( .A(b[15]), .B(a[15]), .Z(n5959) );
  XNOR U6308 ( .A(n5964), .B(n5780), .Z(n5782) );
  XOR U6309 ( .A(n5965), .B(n5966), .Z(n5780) );
  ANDN U6310 ( .B(n5967), .A(n5968), .Z(n5965) );
  AND U6311 ( .A(a[16]), .B(b[14]), .Z(n5964) );
  XNOR U6312 ( .A(n5969), .B(n5785), .Z(n5787) );
  XOR U6313 ( .A(n5970), .B(n5971), .Z(n5785) );
  ANDN U6314 ( .B(n5972), .A(n5973), .Z(n5970) );
  AND U6315 ( .A(b[13]), .B(a[17]), .Z(n5969) );
  XNOR U6316 ( .A(n5974), .B(n5790), .Z(n5792) );
  XOR U6317 ( .A(n5975), .B(n5976), .Z(n5790) );
  ANDN U6318 ( .B(n5977), .A(n5978), .Z(n5975) );
  AND U6319 ( .A(a[18]), .B(b[12]), .Z(n5974) );
  XNOR U6320 ( .A(n5979), .B(n5795), .Z(n5797) );
  XOR U6321 ( .A(n5980), .B(n5981), .Z(n5795) );
  ANDN U6322 ( .B(n5982), .A(n5983), .Z(n5980) );
  AND U6323 ( .A(b[11]), .B(a[19]), .Z(n5979) );
  XNOR U6324 ( .A(n5984), .B(n5800), .Z(n5802) );
  XOR U6325 ( .A(n5985), .B(n5986), .Z(n5800) );
  ANDN U6326 ( .B(n5987), .A(n5988), .Z(n5985) );
  AND U6327 ( .A(a[20]), .B(b[10]), .Z(n5984) );
  XNOR U6328 ( .A(n5989), .B(n5805), .Z(n5807) );
  XOR U6329 ( .A(n5990), .B(n5991), .Z(n5805) );
  ANDN U6330 ( .B(n5992), .A(n5993), .Z(n5990) );
  AND U6331 ( .A(b[9]), .B(a[21]), .Z(n5989) );
  XNOR U6332 ( .A(n5994), .B(n5810), .Z(n5812) );
  XOR U6333 ( .A(n5995), .B(n5996), .Z(n5810) );
  ANDN U6334 ( .B(n5997), .A(n5998), .Z(n5995) );
  AND U6335 ( .A(a[22]), .B(b[8]), .Z(n5994) );
  XNOR U6336 ( .A(n5999), .B(n5815), .Z(n5817) );
  XOR U6337 ( .A(n6000), .B(n6001), .Z(n5815) );
  ANDN U6338 ( .B(n6002), .A(n6003), .Z(n6000) );
  AND U6339 ( .A(b[7]), .B(a[23]), .Z(n5999) );
  XNOR U6340 ( .A(n6004), .B(n5820), .Z(n5822) );
  XOR U6341 ( .A(n6005), .B(n6006), .Z(n5820) );
  ANDN U6342 ( .B(n6007), .A(n6008), .Z(n6005) );
  AND U6343 ( .A(b[6]), .B(a[24]), .Z(n6004) );
  XNOR U6344 ( .A(n6009), .B(n5825), .Z(n5827) );
  XOR U6345 ( .A(n6010), .B(n6011), .Z(n5825) );
  ANDN U6346 ( .B(n6012), .A(n6013), .Z(n6010) );
  AND U6347 ( .A(b[5]), .B(a[25]), .Z(n6009) );
  XNOR U6348 ( .A(n6014), .B(n5830), .Z(n5832) );
  XOR U6349 ( .A(n6015), .B(n6016), .Z(n5830) );
  ANDN U6350 ( .B(n6017), .A(n6018), .Z(n6015) );
  AND U6351 ( .A(b[4]), .B(a[26]), .Z(n6014) );
  XNOR U6352 ( .A(n6019), .B(n6020), .Z(n5844) );
  NANDN U6353 ( .A(n6021), .B(n6022), .Z(n6020) );
  XNOR U6354 ( .A(n6023), .B(n5835), .Z(n5837) );
  XNOR U6355 ( .A(n6024), .B(n6025), .Z(n5835) );
  AND U6356 ( .A(n6026), .B(n6027), .Z(n6024) );
  AND U6357 ( .A(b[3]), .B(a[27]), .Z(n6023) );
  NAND U6358 ( .A(a[30]), .B(b[0]), .Z(n5673) );
  IV U6359 ( .A(n5848), .Z(n5851) );
  XOR U6360 ( .A(n6028), .B(n6029), .Z(n5848) );
  ANDN U6361 ( .B(n6030), .A(n6031), .Z(n6028) );
  XNOR U6362 ( .A(n6030), .B(n6031), .Z(c[61]) );
  XNOR U6363 ( .A(sreg[93]), .B(n6032), .Z(n6031) );
  XNOR U6364 ( .A(n6032), .B(n6033), .Z(n6030) );
  XOR U6365 ( .A(n5856), .B(n5857), .Z(n6033) );
  XNOR U6366 ( .A(n6021), .B(n6022), .Z(n5857) );
  XOR U6367 ( .A(n6019), .B(n6034), .Z(n6022) );
  NAND U6368 ( .A(a[28]), .B(b[1]), .Z(n6034) );
  XOR U6369 ( .A(n6027), .B(n6035), .Z(n6021) );
  XOR U6370 ( .A(n6019), .B(n6026), .Z(n6035) );
  XNOR U6371 ( .A(n6036), .B(n6025), .Z(n6026) );
  AND U6372 ( .A(b[2]), .B(a[27]), .Z(n6036) );
  NANDN U6373 ( .A(n6037), .B(n6038), .Z(n6019) );
  XOR U6374 ( .A(n6025), .B(n6017), .Z(n6039) );
  XNOR U6375 ( .A(n6016), .B(n6012), .Z(n6040) );
  XNOR U6376 ( .A(n6011), .B(n6007), .Z(n6041) );
  XNOR U6377 ( .A(n6006), .B(n6002), .Z(n6042) );
  XNOR U6378 ( .A(n6001), .B(n5997), .Z(n6043) );
  XNOR U6379 ( .A(n5996), .B(n5992), .Z(n6044) );
  XNOR U6380 ( .A(n5991), .B(n5987), .Z(n6045) );
  XNOR U6381 ( .A(n5986), .B(n5982), .Z(n6046) );
  XNOR U6382 ( .A(n5981), .B(n5977), .Z(n6047) );
  XNOR U6383 ( .A(n5976), .B(n5972), .Z(n6048) );
  XNOR U6384 ( .A(n5971), .B(n5967), .Z(n6049) );
  XNOR U6385 ( .A(n5966), .B(n5962), .Z(n6050) );
  XNOR U6386 ( .A(n5961), .B(n5957), .Z(n6051) );
  XNOR U6387 ( .A(n5956), .B(n5952), .Z(n6052) );
  XNOR U6388 ( .A(n5951), .B(n5947), .Z(n6053) );
  XNOR U6389 ( .A(n5946), .B(n5942), .Z(n6054) );
  XNOR U6390 ( .A(n5941), .B(n5937), .Z(n6055) );
  XNOR U6391 ( .A(n5936), .B(n5932), .Z(n6056) );
  XNOR U6392 ( .A(n5931), .B(n5927), .Z(n6057) );
  XNOR U6393 ( .A(n5926), .B(n5922), .Z(n6058) );
  XNOR U6394 ( .A(n5921), .B(n5917), .Z(n6059) );
  XNOR U6395 ( .A(n5916), .B(n5912), .Z(n6060) );
  XNOR U6396 ( .A(n5911), .B(n5907), .Z(n6061) );
  XNOR U6397 ( .A(n5906), .B(n5902), .Z(n6062) );
  XNOR U6398 ( .A(n5901), .B(n5897), .Z(n6063) );
  XNOR U6399 ( .A(n5896), .B(n5892), .Z(n6064) );
  XOR U6400 ( .A(n6065), .B(n5891), .Z(n5892) );
  AND U6401 ( .A(a[0]), .B(b[29]), .Z(n6065) );
  XNOR U6402 ( .A(n6066), .B(n5891), .Z(n5893) );
  XNOR U6403 ( .A(n6067), .B(n6068), .Z(n5891) );
  ANDN U6404 ( .B(n6069), .A(n6070), .Z(n6067) );
  AND U6405 ( .A(a[1]), .B(b[28]), .Z(n6066) );
  XNOR U6406 ( .A(n6071), .B(n5896), .Z(n5898) );
  XOR U6407 ( .A(n6072), .B(n6073), .Z(n5896) );
  ANDN U6408 ( .B(n6074), .A(n6075), .Z(n6072) );
  AND U6409 ( .A(a[2]), .B(b[27]), .Z(n6071) );
  XNOR U6410 ( .A(n6076), .B(n5901), .Z(n5903) );
  XOR U6411 ( .A(n6077), .B(n6078), .Z(n5901) );
  ANDN U6412 ( .B(n6079), .A(n6080), .Z(n6077) );
  AND U6413 ( .A(a[3]), .B(b[26]), .Z(n6076) );
  XNOR U6414 ( .A(n6081), .B(n5906), .Z(n5908) );
  XOR U6415 ( .A(n6082), .B(n6083), .Z(n5906) );
  ANDN U6416 ( .B(n6084), .A(n6085), .Z(n6082) );
  AND U6417 ( .A(a[4]), .B(b[25]), .Z(n6081) );
  XNOR U6418 ( .A(n6086), .B(n5911), .Z(n5913) );
  XOR U6419 ( .A(n6087), .B(n6088), .Z(n5911) );
  ANDN U6420 ( .B(n6089), .A(n6090), .Z(n6087) );
  AND U6421 ( .A(a[5]), .B(b[24]), .Z(n6086) );
  XNOR U6422 ( .A(n6091), .B(n5916), .Z(n5918) );
  XOR U6423 ( .A(n6092), .B(n6093), .Z(n5916) );
  ANDN U6424 ( .B(n6094), .A(n6095), .Z(n6092) );
  AND U6425 ( .A(a[6]), .B(b[23]), .Z(n6091) );
  XNOR U6426 ( .A(n6096), .B(n5921), .Z(n5923) );
  XOR U6427 ( .A(n6097), .B(n6098), .Z(n5921) );
  ANDN U6428 ( .B(n6099), .A(n6100), .Z(n6097) );
  AND U6429 ( .A(a[7]), .B(b[22]), .Z(n6096) );
  XNOR U6430 ( .A(n6101), .B(n5926), .Z(n5928) );
  XOR U6431 ( .A(n6102), .B(n6103), .Z(n5926) );
  ANDN U6432 ( .B(n6104), .A(n6105), .Z(n6102) );
  AND U6433 ( .A(a[8]), .B(b[21]), .Z(n6101) );
  XNOR U6434 ( .A(n6106), .B(n5931), .Z(n5933) );
  XOR U6435 ( .A(n6107), .B(n6108), .Z(n5931) );
  ANDN U6436 ( .B(n6109), .A(n6110), .Z(n6107) );
  AND U6437 ( .A(a[9]), .B(b[20]), .Z(n6106) );
  XNOR U6438 ( .A(n6111), .B(n5936), .Z(n5938) );
  XOR U6439 ( .A(n6112), .B(n6113), .Z(n5936) );
  ANDN U6440 ( .B(n6114), .A(n6115), .Z(n6112) );
  AND U6441 ( .A(a[10]), .B(b[19]), .Z(n6111) );
  XNOR U6442 ( .A(n6116), .B(n5941), .Z(n5943) );
  XOR U6443 ( .A(n6117), .B(n6118), .Z(n5941) );
  ANDN U6444 ( .B(n6119), .A(n6120), .Z(n6117) );
  AND U6445 ( .A(a[11]), .B(b[18]), .Z(n6116) );
  XNOR U6446 ( .A(n6121), .B(n5946), .Z(n5948) );
  XOR U6447 ( .A(n6122), .B(n6123), .Z(n5946) );
  ANDN U6448 ( .B(n6124), .A(n6125), .Z(n6122) );
  AND U6449 ( .A(a[12]), .B(b[17]), .Z(n6121) );
  XNOR U6450 ( .A(n6126), .B(n5951), .Z(n5953) );
  XOR U6451 ( .A(n6127), .B(n6128), .Z(n5951) );
  ANDN U6452 ( .B(n6129), .A(n6130), .Z(n6127) );
  AND U6453 ( .A(a[13]), .B(b[16]), .Z(n6126) );
  XNOR U6454 ( .A(n6131), .B(n5956), .Z(n5958) );
  XOR U6455 ( .A(n6132), .B(n6133), .Z(n5956) );
  ANDN U6456 ( .B(n6134), .A(n6135), .Z(n6132) );
  AND U6457 ( .A(a[14]), .B(b[15]), .Z(n6131) );
  XNOR U6458 ( .A(n6136), .B(n5961), .Z(n5963) );
  XOR U6459 ( .A(n6137), .B(n6138), .Z(n5961) );
  ANDN U6460 ( .B(n6139), .A(n6140), .Z(n6137) );
  AND U6461 ( .A(b[14]), .B(a[15]), .Z(n6136) );
  XNOR U6462 ( .A(n6141), .B(n5966), .Z(n5968) );
  XOR U6463 ( .A(n6142), .B(n6143), .Z(n5966) );
  ANDN U6464 ( .B(n6144), .A(n6145), .Z(n6142) );
  AND U6465 ( .A(a[16]), .B(b[13]), .Z(n6141) );
  XNOR U6466 ( .A(n6146), .B(n5971), .Z(n5973) );
  XOR U6467 ( .A(n6147), .B(n6148), .Z(n5971) );
  ANDN U6468 ( .B(n6149), .A(n6150), .Z(n6147) );
  AND U6469 ( .A(b[12]), .B(a[17]), .Z(n6146) );
  XNOR U6470 ( .A(n6151), .B(n5976), .Z(n5978) );
  XOR U6471 ( .A(n6152), .B(n6153), .Z(n5976) );
  ANDN U6472 ( .B(n6154), .A(n6155), .Z(n6152) );
  AND U6473 ( .A(a[18]), .B(b[11]), .Z(n6151) );
  XNOR U6474 ( .A(n6156), .B(n5981), .Z(n5983) );
  XOR U6475 ( .A(n6157), .B(n6158), .Z(n5981) );
  ANDN U6476 ( .B(n6159), .A(n6160), .Z(n6157) );
  AND U6477 ( .A(b[10]), .B(a[19]), .Z(n6156) );
  XNOR U6478 ( .A(n6161), .B(n5986), .Z(n5988) );
  XOR U6479 ( .A(n6162), .B(n6163), .Z(n5986) );
  ANDN U6480 ( .B(n6164), .A(n6165), .Z(n6162) );
  AND U6481 ( .A(a[20]), .B(b[9]), .Z(n6161) );
  XNOR U6482 ( .A(n6166), .B(n5991), .Z(n5993) );
  XOR U6483 ( .A(n6167), .B(n6168), .Z(n5991) );
  ANDN U6484 ( .B(n6169), .A(n6170), .Z(n6167) );
  AND U6485 ( .A(b[8]), .B(a[21]), .Z(n6166) );
  XNOR U6486 ( .A(n6171), .B(n5996), .Z(n5998) );
  XOR U6487 ( .A(n6172), .B(n6173), .Z(n5996) );
  ANDN U6488 ( .B(n6174), .A(n6175), .Z(n6172) );
  AND U6489 ( .A(a[22]), .B(b[7]), .Z(n6171) );
  XNOR U6490 ( .A(n6176), .B(n6001), .Z(n6003) );
  XOR U6491 ( .A(n6177), .B(n6178), .Z(n6001) );
  ANDN U6492 ( .B(n6179), .A(n6180), .Z(n6177) );
  AND U6493 ( .A(b[6]), .B(a[23]), .Z(n6176) );
  XNOR U6494 ( .A(n6181), .B(n6006), .Z(n6008) );
  XOR U6495 ( .A(n6182), .B(n6183), .Z(n6006) );
  ANDN U6496 ( .B(n6184), .A(n6185), .Z(n6182) );
  AND U6497 ( .A(b[5]), .B(a[24]), .Z(n6181) );
  XNOR U6498 ( .A(n6186), .B(n6011), .Z(n6013) );
  XOR U6499 ( .A(n6187), .B(n6188), .Z(n6011) );
  ANDN U6500 ( .B(n6189), .A(n6190), .Z(n6187) );
  AND U6501 ( .A(b[4]), .B(a[25]), .Z(n6186) );
  XNOR U6502 ( .A(n6191), .B(n6192), .Z(n6025) );
  NANDN U6503 ( .A(n6193), .B(n6194), .Z(n6192) );
  XNOR U6504 ( .A(n6195), .B(n6016), .Z(n6018) );
  XNOR U6505 ( .A(n6196), .B(n6197), .Z(n6016) );
  AND U6506 ( .A(n6198), .B(n6199), .Z(n6196) );
  AND U6507 ( .A(b[3]), .B(a[26]), .Z(n6195) );
  NAND U6508 ( .A(a[29]), .B(b[0]), .Z(n5856) );
  IV U6509 ( .A(n6029), .Z(n6032) );
  XOR U6510 ( .A(n6200), .B(n6201), .Z(n6029) );
  ANDN U6511 ( .B(n6202), .A(n6203), .Z(n6200) );
  XNOR U6512 ( .A(n6202), .B(n6203), .Z(c[60]) );
  XNOR U6513 ( .A(sreg[92]), .B(n6204), .Z(n6203) );
  XNOR U6514 ( .A(n6204), .B(n6205), .Z(n6202) );
  XOR U6515 ( .A(n6037), .B(n6038), .Z(n6205) );
  XNOR U6516 ( .A(n6193), .B(n6194), .Z(n6038) );
  XOR U6517 ( .A(n6191), .B(n6206), .Z(n6194) );
  NAND U6518 ( .A(b[1]), .B(a[27]), .Z(n6206) );
  XOR U6519 ( .A(n6199), .B(n6207), .Z(n6193) );
  XOR U6520 ( .A(n6191), .B(n6198), .Z(n6207) );
  XNOR U6521 ( .A(n6208), .B(n6197), .Z(n6198) );
  AND U6522 ( .A(b[2]), .B(a[26]), .Z(n6208) );
  NANDN U6523 ( .A(n6209), .B(n6210), .Z(n6191) );
  XOR U6524 ( .A(n6197), .B(n6189), .Z(n6211) );
  XNOR U6525 ( .A(n6188), .B(n6184), .Z(n6212) );
  XNOR U6526 ( .A(n6183), .B(n6179), .Z(n6213) );
  XNOR U6527 ( .A(n6178), .B(n6174), .Z(n6214) );
  XNOR U6528 ( .A(n6173), .B(n6169), .Z(n6215) );
  XNOR U6529 ( .A(n6168), .B(n6164), .Z(n6216) );
  XNOR U6530 ( .A(n6163), .B(n6159), .Z(n6217) );
  XNOR U6531 ( .A(n6158), .B(n6154), .Z(n6218) );
  XNOR U6532 ( .A(n6153), .B(n6149), .Z(n6219) );
  XNOR U6533 ( .A(n6148), .B(n6144), .Z(n6220) );
  XNOR U6534 ( .A(n6143), .B(n6139), .Z(n6221) );
  XNOR U6535 ( .A(n6138), .B(n6134), .Z(n6222) );
  XNOR U6536 ( .A(n6133), .B(n6129), .Z(n6223) );
  XNOR U6537 ( .A(n6128), .B(n6124), .Z(n6224) );
  XNOR U6538 ( .A(n6123), .B(n6119), .Z(n6225) );
  XNOR U6539 ( .A(n6118), .B(n6114), .Z(n6226) );
  XNOR U6540 ( .A(n6113), .B(n6109), .Z(n6227) );
  XNOR U6541 ( .A(n6108), .B(n6104), .Z(n6228) );
  XNOR U6542 ( .A(n6103), .B(n6099), .Z(n6229) );
  XNOR U6543 ( .A(n6098), .B(n6094), .Z(n6230) );
  XNOR U6544 ( .A(n6093), .B(n6089), .Z(n6231) );
  XNOR U6545 ( .A(n6088), .B(n6084), .Z(n6232) );
  XNOR U6546 ( .A(n6083), .B(n6079), .Z(n6233) );
  XNOR U6547 ( .A(n6078), .B(n6074), .Z(n6234) );
  XNOR U6548 ( .A(n6073), .B(n6069), .Z(n6235) );
  XNOR U6549 ( .A(n6236), .B(n6068), .Z(n6069) );
  AND U6550 ( .A(a[0]), .B(b[28]), .Z(n6236) );
  XOR U6551 ( .A(n6237), .B(n6068), .Z(n6070) );
  XNOR U6552 ( .A(n6238), .B(n6239), .Z(n6068) );
  ANDN U6553 ( .B(n6240), .A(n6241), .Z(n6238) );
  AND U6554 ( .A(a[1]), .B(b[27]), .Z(n6237) );
  XNOR U6555 ( .A(n6242), .B(n6073), .Z(n6075) );
  XOR U6556 ( .A(n6243), .B(n6244), .Z(n6073) );
  ANDN U6557 ( .B(n6245), .A(n6246), .Z(n6243) );
  AND U6558 ( .A(a[2]), .B(b[26]), .Z(n6242) );
  XNOR U6559 ( .A(n6247), .B(n6078), .Z(n6080) );
  XOR U6560 ( .A(n6248), .B(n6249), .Z(n6078) );
  ANDN U6561 ( .B(n6250), .A(n6251), .Z(n6248) );
  AND U6562 ( .A(a[3]), .B(b[25]), .Z(n6247) );
  XNOR U6563 ( .A(n6252), .B(n6083), .Z(n6085) );
  XOR U6564 ( .A(n6253), .B(n6254), .Z(n6083) );
  ANDN U6565 ( .B(n6255), .A(n6256), .Z(n6253) );
  AND U6566 ( .A(a[4]), .B(b[24]), .Z(n6252) );
  XNOR U6567 ( .A(n6257), .B(n6088), .Z(n6090) );
  XOR U6568 ( .A(n6258), .B(n6259), .Z(n6088) );
  ANDN U6569 ( .B(n6260), .A(n6261), .Z(n6258) );
  AND U6570 ( .A(a[5]), .B(b[23]), .Z(n6257) );
  XNOR U6571 ( .A(n6262), .B(n6093), .Z(n6095) );
  XOR U6572 ( .A(n6263), .B(n6264), .Z(n6093) );
  ANDN U6573 ( .B(n6265), .A(n6266), .Z(n6263) );
  AND U6574 ( .A(a[6]), .B(b[22]), .Z(n6262) );
  XNOR U6575 ( .A(n6267), .B(n6098), .Z(n6100) );
  XOR U6576 ( .A(n6268), .B(n6269), .Z(n6098) );
  ANDN U6577 ( .B(n6270), .A(n6271), .Z(n6268) );
  AND U6578 ( .A(a[7]), .B(b[21]), .Z(n6267) );
  XNOR U6579 ( .A(n6272), .B(n6103), .Z(n6105) );
  XOR U6580 ( .A(n6273), .B(n6274), .Z(n6103) );
  ANDN U6581 ( .B(n6275), .A(n6276), .Z(n6273) );
  AND U6582 ( .A(a[8]), .B(b[20]), .Z(n6272) );
  XNOR U6583 ( .A(n6277), .B(n6108), .Z(n6110) );
  XOR U6584 ( .A(n6278), .B(n6279), .Z(n6108) );
  ANDN U6585 ( .B(n6280), .A(n6281), .Z(n6278) );
  AND U6586 ( .A(a[9]), .B(b[19]), .Z(n6277) );
  XNOR U6587 ( .A(n6282), .B(n6113), .Z(n6115) );
  XOR U6588 ( .A(n6283), .B(n6284), .Z(n6113) );
  ANDN U6589 ( .B(n6285), .A(n6286), .Z(n6283) );
  AND U6590 ( .A(a[10]), .B(b[18]), .Z(n6282) );
  XNOR U6591 ( .A(n6287), .B(n6118), .Z(n6120) );
  XOR U6592 ( .A(n6288), .B(n6289), .Z(n6118) );
  ANDN U6593 ( .B(n6290), .A(n6291), .Z(n6288) );
  AND U6594 ( .A(a[11]), .B(b[17]), .Z(n6287) );
  XNOR U6595 ( .A(n6292), .B(n6123), .Z(n6125) );
  XOR U6596 ( .A(n6293), .B(n6294), .Z(n6123) );
  ANDN U6597 ( .B(n6295), .A(n6296), .Z(n6293) );
  AND U6598 ( .A(a[12]), .B(b[16]), .Z(n6292) );
  XNOR U6599 ( .A(n6297), .B(n6128), .Z(n6130) );
  XOR U6600 ( .A(n6298), .B(n6299), .Z(n6128) );
  ANDN U6601 ( .B(n6300), .A(n6301), .Z(n6298) );
  AND U6602 ( .A(a[13]), .B(b[15]), .Z(n6297) );
  XNOR U6603 ( .A(n6302), .B(n6133), .Z(n6135) );
  XOR U6604 ( .A(n6303), .B(n6304), .Z(n6133) );
  ANDN U6605 ( .B(n6305), .A(n6306), .Z(n6303) );
  AND U6606 ( .A(a[14]), .B(b[14]), .Z(n6302) );
  XNOR U6607 ( .A(n6307), .B(n6138), .Z(n6140) );
  XOR U6608 ( .A(n6308), .B(n6309), .Z(n6138) );
  ANDN U6609 ( .B(n6310), .A(n6311), .Z(n6308) );
  AND U6610 ( .A(b[13]), .B(a[15]), .Z(n6307) );
  XNOR U6611 ( .A(n6312), .B(n6143), .Z(n6145) );
  XOR U6612 ( .A(n6313), .B(n6314), .Z(n6143) );
  ANDN U6613 ( .B(n6315), .A(n6316), .Z(n6313) );
  AND U6614 ( .A(a[16]), .B(b[12]), .Z(n6312) );
  XNOR U6615 ( .A(n6317), .B(n6148), .Z(n6150) );
  XOR U6616 ( .A(n6318), .B(n6319), .Z(n6148) );
  ANDN U6617 ( .B(n6320), .A(n6321), .Z(n6318) );
  AND U6618 ( .A(b[11]), .B(a[17]), .Z(n6317) );
  XNOR U6619 ( .A(n6322), .B(n6153), .Z(n6155) );
  XOR U6620 ( .A(n6323), .B(n6324), .Z(n6153) );
  ANDN U6621 ( .B(n6325), .A(n6326), .Z(n6323) );
  AND U6622 ( .A(a[18]), .B(b[10]), .Z(n6322) );
  XNOR U6623 ( .A(n6327), .B(n6158), .Z(n6160) );
  XOR U6624 ( .A(n6328), .B(n6329), .Z(n6158) );
  ANDN U6625 ( .B(n6330), .A(n6331), .Z(n6328) );
  AND U6626 ( .A(b[9]), .B(a[19]), .Z(n6327) );
  XNOR U6627 ( .A(n6332), .B(n6163), .Z(n6165) );
  XOR U6628 ( .A(n6333), .B(n6334), .Z(n6163) );
  ANDN U6629 ( .B(n6335), .A(n6336), .Z(n6333) );
  AND U6630 ( .A(a[20]), .B(b[8]), .Z(n6332) );
  XNOR U6631 ( .A(n6337), .B(n6168), .Z(n6170) );
  XOR U6632 ( .A(n6338), .B(n6339), .Z(n6168) );
  ANDN U6633 ( .B(n6340), .A(n6341), .Z(n6338) );
  AND U6634 ( .A(b[7]), .B(a[21]), .Z(n6337) );
  XNOR U6635 ( .A(n6342), .B(n6173), .Z(n6175) );
  XOR U6636 ( .A(n6343), .B(n6344), .Z(n6173) );
  ANDN U6637 ( .B(n6345), .A(n6346), .Z(n6343) );
  AND U6638 ( .A(b[6]), .B(a[22]), .Z(n6342) );
  XNOR U6639 ( .A(n6347), .B(n6178), .Z(n6180) );
  XOR U6640 ( .A(n6348), .B(n6349), .Z(n6178) );
  ANDN U6641 ( .B(n6350), .A(n6351), .Z(n6348) );
  AND U6642 ( .A(b[5]), .B(a[23]), .Z(n6347) );
  XNOR U6643 ( .A(n6352), .B(n6183), .Z(n6185) );
  XOR U6644 ( .A(n6353), .B(n6354), .Z(n6183) );
  ANDN U6645 ( .B(n6355), .A(n6356), .Z(n6353) );
  AND U6646 ( .A(b[4]), .B(a[24]), .Z(n6352) );
  XNOR U6647 ( .A(n6357), .B(n6358), .Z(n6197) );
  NANDN U6648 ( .A(n6359), .B(n6360), .Z(n6358) );
  XNOR U6649 ( .A(n6361), .B(n6188), .Z(n6190) );
  XNOR U6650 ( .A(n6362), .B(n6363), .Z(n6188) );
  AND U6651 ( .A(n6364), .B(n6365), .Z(n6362) );
  AND U6652 ( .A(b[3]), .B(a[25]), .Z(n6361) );
  NAND U6653 ( .A(a[28]), .B(b[0]), .Z(n6037) );
  IV U6654 ( .A(n6201), .Z(n6204) );
  XOR U6655 ( .A(n6366), .B(n6367), .Z(n6201) );
  ANDN U6656 ( .B(n6368), .A(n6369), .Z(n6366) );
  XNOR U6657 ( .A(n6368), .B(n6369), .Z(c[59]) );
  XNOR U6658 ( .A(sreg[91]), .B(n6370), .Z(n6369) );
  XNOR U6659 ( .A(n6370), .B(n6371), .Z(n6368) );
  XOR U6660 ( .A(n6209), .B(n6210), .Z(n6371) );
  XNOR U6661 ( .A(n6359), .B(n6360), .Z(n6210) );
  XOR U6662 ( .A(n6357), .B(n6372), .Z(n6360) );
  NAND U6663 ( .A(a[26]), .B(b[1]), .Z(n6372) );
  XOR U6664 ( .A(n6365), .B(n6373), .Z(n6359) );
  XOR U6665 ( .A(n6357), .B(n6364), .Z(n6373) );
  XNOR U6666 ( .A(n6374), .B(n6363), .Z(n6364) );
  AND U6667 ( .A(b[2]), .B(a[25]), .Z(n6374) );
  NANDN U6668 ( .A(n6375), .B(n6376), .Z(n6357) );
  XOR U6669 ( .A(n6363), .B(n6355), .Z(n6377) );
  XNOR U6670 ( .A(n6354), .B(n6350), .Z(n6378) );
  XNOR U6671 ( .A(n6349), .B(n6345), .Z(n6379) );
  XNOR U6672 ( .A(n6344), .B(n6340), .Z(n6380) );
  XNOR U6673 ( .A(n6339), .B(n6335), .Z(n6381) );
  XNOR U6674 ( .A(n6334), .B(n6330), .Z(n6382) );
  XNOR U6675 ( .A(n6329), .B(n6325), .Z(n6383) );
  XNOR U6676 ( .A(n6324), .B(n6320), .Z(n6384) );
  XNOR U6677 ( .A(n6319), .B(n6315), .Z(n6385) );
  XNOR U6678 ( .A(n6314), .B(n6310), .Z(n6386) );
  XNOR U6679 ( .A(n6309), .B(n6305), .Z(n6387) );
  XNOR U6680 ( .A(n6304), .B(n6300), .Z(n6388) );
  XNOR U6681 ( .A(n6299), .B(n6295), .Z(n6389) );
  XNOR U6682 ( .A(n6294), .B(n6290), .Z(n6390) );
  XNOR U6683 ( .A(n6289), .B(n6285), .Z(n6391) );
  XNOR U6684 ( .A(n6284), .B(n6280), .Z(n6392) );
  XNOR U6685 ( .A(n6279), .B(n6275), .Z(n6393) );
  XNOR U6686 ( .A(n6274), .B(n6270), .Z(n6394) );
  XNOR U6687 ( .A(n6269), .B(n6265), .Z(n6395) );
  XNOR U6688 ( .A(n6264), .B(n6260), .Z(n6396) );
  XNOR U6689 ( .A(n6259), .B(n6255), .Z(n6397) );
  XNOR U6690 ( .A(n6254), .B(n6250), .Z(n6398) );
  XNOR U6691 ( .A(n6249), .B(n6245), .Z(n6399) );
  XNOR U6692 ( .A(n6244), .B(n6240), .Z(n6400) );
  XOR U6693 ( .A(n6401), .B(n6239), .Z(n6240) );
  AND U6694 ( .A(a[0]), .B(b[27]), .Z(n6401) );
  XNOR U6695 ( .A(n6402), .B(n6239), .Z(n6241) );
  XNOR U6696 ( .A(n6403), .B(n6404), .Z(n6239) );
  ANDN U6697 ( .B(n6405), .A(n6406), .Z(n6403) );
  AND U6698 ( .A(a[1]), .B(b[26]), .Z(n6402) );
  XNOR U6699 ( .A(n6407), .B(n6244), .Z(n6246) );
  XOR U6700 ( .A(n6408), .B(n6409), .Z(n6244) );
  ANDN U6701 ( .B(n6410), .A(n6411), .Z(n6408) );
  AND U6702 ( .A(a[2]), .B(b[25]), .Z(n6407) );
  XNOR U6703 ( .A(n6412), .B(n6249), .Z(n6251) );
  XOR U6704 ( .A(n6413), .B(n6414), .Z(n6249) );
  ANDN U6705 ( .B(n6415), .A(n6416), .Z(n6413) );
  AND U6706 ( .A(a[3]), .B(b[24]), .Z(n6412) );
  XNOR U6707 ( .A(n6417), .B(n6254), .Z(n6256) );
  XOR U6708 ( .A(n6418), .B(n6419), .Z(n6254) );
  ANDN U6709 ( .B(n6420), .A(n6421), .Z(n6418) );
  AND U6710 ( .A(a[4]), .B(b[23]), .Z(n6417) );
  XNOR U6711 ( .A(n6422), .B(n6259), .Z(n6261) );
  XOR U6712 ( .A(n6423), .B(n6424), .Z(n6259) );
  ANDN U6713 ( .B(n6425), .A(n6426), .Z(n6423) );
  AND U6714 ( .A(a[5]), .B(b[22]), .Z(n6422) );
  XNOR U6715 ( .A(n6427), .B(n6264), .Z(n6266) );
  XOR U6716 ( .A(n6428), .B(n6429), .Z(n6264) );
  ANDN U6717 ( .B(n6430), .A(n6431), .Z(n6428) );
  AND U6718 ( .A(a[6]), .B(b[21]), .Z(n6427) );
  XNOR U6719 ( .A(n6432), .B(n6269), .Z(n6271) );
  XOR U6720 ( .A(n6433), .B(n6434), .Z(n6269) );
  ANDN U6721 ( .B(n6435), .A(n6436), .Z(n6433) );
  AND U6722 ( .A(a[7]), .B(b[20]), .Z(n6432) );
  XNOR U6723 ( .A(n6437), .B(n6274), .Z(n6276) );
  XOR U6724 ( .A(n6438), .B(n6439), .Z(n6274) );
  ANDN U6725 ( .B(n6440), .A(n6441), .Z(n6438) );
  AND U6726 ( .A(a[8]), .B(b[19]), .Z(n6437) );
  XNOR U6727 ( .A(n6442), .B(n6279), .Z(n6281) );
  XOR U6728 ( .A(n6443), .B(n6444), .Z(n6279) );
  ANDN U6729 ( .B(n6445), .A(n6446), .Z(n6443) );
  AND U6730 ( .A(a[9]), .B(b[18]), .Z(n6442) );
  XNOR U6731 ( .A(n6447), .B(n6284), .Z(n6286) );
  XOR U6732 ( .A(n6448), .B(n6449), .Z(n6284) );
  ANDN U6733 ( .B(n6450), .A(n6451), .Z(n6448) );
  AND U6734 ( .A(a[10]), .B(b[17]), .Z(n6447) );
  XNOR U6735 ( .A(n6452), .B(n6289), .Z(n6291) );
  XOR U6736 ( .A(n6453), .B(n6454), .Z(n6289) );
  ANDN U6737 ( .B(n6455), .A(n6456), .Z(n6453) );
  AND U6738 ( .A(a[11]), .B(b[16]), .Z(n6452) );
  XNOR U6739 ( .A(n6457), .B(n6294), .Z(n6296) );
  XOR U6740 ( .A(n6458), .B(n6459), .Z(n6294) );
  ANDN U6741 ( .B(n6460), .A(n6461), .Z(n6458) );
  AND U6742 ( .A(a[12]), .B(b[15]), .Z(n6457) );
  XNOR U6743 ( .A(n6462), .B(n6299), .Z(n6301) );
  XOR U6744 ( .A(n6463), .B(n6464), .Z(n6299) );
  ANDN U6745 ( .B(n6465), .A(n6466), .Z(n6463) );
  AND U6746 ( .A(a[13]), .B(b[14]), .Z(n6462) );
  XNOR U6747 ( .A(n6467), .B(n6304), .Z(n6306) );
  XOR U6748 ( .A(n6468), .B(n6469), .Z(n6304) );
  ANDN U6749 ( .B(n6470), .A(n6471), .Z(n6468) );
  AND U6750 ( .A(a[14]), .B(b[13]), .Z(n6467) );
  XNOR U6751 ( .A(n6472), .B(n6309), .Z(n6311) );
  XOR U6752 ( .A(n6473), .B(n6474), .Z(n6309) );
  ANDN U6753 ( .B(n6475), .A(n6476), .Z(n6473) );
  AND U6754 ( .A(b[12]), .B(a[15]), .Z(n6472) );
  XNOR U6755 ( .A(n6477), .B(n6314), .Z(n6316) );
  XOR U6756 ( .A(n6478), .B(n6479), .Z(n6314) );
  ANDN U6757 ( .B(n6480), .A(n6481), .Z(n6478) );
  AND U6758 ( .A(a[16]), .B(b[11]), .Z(n6477) );
  XNOR U6759 ( .A(n6482), .B(n6319), .Z(n6321) );
  XOR U6760 ( .A(n6483), .B(n6484), .Z(n6319) );
  ANDN U6761 ( .B(n6485), .A(n6486), .Z(n6483) );
  AND U6762 ( .A(b[10]), .B(a[17]), .Z(n6482) );
  XNOR U6763 ( .A(n6487), .B(n6324), .Z(n6326) );
  XOR U6764 ( .A(n6488), .B(n6489), .Z(n6324) );
  ANDN U6765 ( .B(n6490), .A(n6491), .Z(n6488) );
  AND U6766 ( .A(a[18]), .B(b[9]), .Z(n6487) );
  XNOR U6767 ( .A(n6492), .B(n6329), .Z(n6331) );
  XOR U6768 ( .A(n6493), .B(n6494), .Z(n6329) );
  ANDN U6769 ( .B(n6495), .A(n6496), .Z(n6493) );
  AND U6770 ( .A(b[8]), .B(a[19]), .Z(n6492) );
  XNOR U6771 ( .A(n6497), .B(n6334), .Z(n6336) );
  XOR U6772 ( .A(n6498), .B(n6499), .Z(n6334) );
  ANDN U6773 ( .B(n6500), .A(n6501), .Z(n6498) );
  AND U6774 ( .A(a[20]), .B(b[7]), .Z(n6497) );
  XNOR U6775 ( .A(n6502), .B(n6339), .Z(n6341) );
  XOR U6776 ( .A(n6503), .B(n6504), .Z(n6339) );
  ANDN U6777 ( .B(n6505), .A(n6506), .Z(n6503) );
  AND U6778 ( .A(b[6]), .B(a[21]), .Z(n6502) );
  XNOR U6779 ( .A(n6507), .B(n6344), .Z(n6346) );
  XOR U6780 ( .A(n6508), .B(n6509), .Z(n6344) );
  ANDN U6781 ( .B(n6510), .A(n6511), .Z(n6508) );
  AND U6782 ( .A(b[5]), .B(a[22]), .Z(n6507) );
  XNOR U6783 ( .A(n6512), .B(n6349), .Z(n6351) );
  XOR U6784 ( .A(n6513), .B(n6514), .Z(n6349) );
  ANDN U6785 ( .B(n6515), .A(n6516), .Z(n6513) );
  AND U6786 ( .A(b[4]), .B(a[23]), .Z(n6512) );
  XNOR U6787 ( .A(n6517), .B(n6518), .Z(n6363) );
  NANDN U6788 ( .A(n6519), .B(n6520), .Z(n6518) );
  XNOR U6789 ( .A(n6521), .B(n6354), .Z(n6356) );
  XNOR U6790 ( .A(n6522), .B(n6523), .Z(n6354) );
  AND U6791 ( .A(n6524), .B(n6525), .Z(n6522) );
  AND U6792 ( .A(b[3]), .B(a[24]), .Z(n6521) );
  NAND U6793 ( .A(a[27]), .B(b[0]), .Z(n6209) );
  IV U6794 ( .A(n6367), .Z(n6370) );
  XOR U6795 ( .A(n6526), .B(n6527), .Z(n6367) );
  ANDN U6796 ( .B(n6528), .A(n6529), .Z(n6526) );
  XNOR U6797 ( .A(n6528), .B(n6529), .Z(c[58]) );
  XNOR U6798 ( .A(sreg[90]), .B(n6530), .Z(n6529) );
  XNOR U6799 ( .A(n6530), .B(n6531), .Z(n6528) );
  XOR U6800 ( .A(n6375), .B(n6376), .Z(n6531) );
  XNOR U6801 ( .A(n6519), .B(n6520), .Z(n6376) );
  XOR U6802 ( .A(n6517), .B(n6532), .Z(n6520) );
  NAND U6803 ( .A(b[1]), .B(a[25]), .Z(n6532) );
  XOR U6804 ( .A(n6525), .B(n6533), .Z(n6519) );
  XOR U6805 ( .A(n6517), .B(n6524), .Z(n6533) );
  XNOR U6806 ( .A(n6534), .B(n6523), .Z(n6524) );
  AND U6807 ( .A(b[2]), .B(a[24]), .Z(n6534) );
  NANDN U6808 ( .A(n6535), .B(n6536), .Z(n6517) );
  XOR U6809 ( .A(n6523), .B(n6515), .Z(n6537) );
  XNOR U6810 ( .A(n6514), .B(n6510), .Z(n6538) );
  XNOR U6811 ( .A(n6509), .B(n6505), .Z(n6539) );
  XNOR U6812 ( .A(n6504), .B(n6500), .Z(n6540) );
  XNOR U6813 ( .A(n6499), .B(n6495), .Z(n6541) );
  XNOR U6814 ( .A(n6494), .B(n6490), .Z(n6542) );
  XNOR U6815 ( .A(n6489), .B(n6485), .Z(n6543) );
  XNOR U6816 ( .A(n6484), .B(n6480), .Z(n6544) );
  XNOR U6817 ( .A(n6479), .B(n6475), .Z(n6545) );
  XNOR U6818 ( .A(n6474), .B(n6470), .Z(n6546) );
  XNOR U6819 ( .A(n6469), .B(n6465), .Z(n6547) );
  XNOR U6820 ( .A(n6464), .B(n6460), .Z(n6548) );
  XNOR U6821 ( .A(n6459), .B(n6455), .Z(n6549) );
  XNOR U6822 ( .A(n6454), .B(n6450), .Z(n6550) );
  XNOR U6823 ( .A(n6449), .B(n6445), .Z(n6551) );
  XNOR U6824 ( .A(n6444), .B(n6440), .Z(n6552) );
  XNOR U6825 ( .A(n6439), .B(n6435), .Z(n6553) );
  XNOR U6826 ( .A(n6434), .B(n6430), .Z(n6554) );
  XNOR U6827 ( .A(n6429), .B(n6425), .Z(n6555) );
  XNOR U6828 ( .A(n6424), .B(n6420), .Z(n6556) );
  XNOR U6829 ( .A(n6419), .B(n6415), .Z(n6557) );
  XNOR U6830 ( .A(n6414), .B(n6410), .Z(n6558) );
  XNOR U6831 ( .A(n6409), .B(n6405), .Z(n6559) );
  XNOR U6832 ( .A(n6560), .B(n6404), .Z(n6405) );
  AND U6833 ( .A(a[0]), .B(b[26]), .Z(n6560) );
  XOR U6834 ( .A(n6561), .B(n6404), .Z(n6406) );
  XNOR U6835 ( .A(n6562), .B(n6563), .Z(n6404) );
  ANDN U6836 ( .B(n6564), .A(n6565), .Z(n6562) );
  AND U6837 ( .A(a[1]), .B(b[25]), .Z(n6561) );
  XNOR U6838 ( .A(n6566), .B(n6409), .Z(n6411) );
  XOR U6839 ( .A(n6567), .B(n6568), .Z(n6409) );
  ANDN U6840 ( .B(n6569), .A(n6570), .Z(n6567) );
  AND U6841 ( .A(a[2]), .B(b[24]), .Z(n6566) );
  XNOR U6842 ( .A(n6571), .B(n6414), .Z(n6416) );
  XOR U6843 ( .A(n6572), .B(n6573), .Z(n6414) );
  ANDN U6844 ( .B(n6574), .A(n6575), .Z(n6572) );
  AND U6845 ( .A(a[3]), .B(b[23]), .Z(n6571) );
  XNOR U6846 ( .A(n6576), .B(n6419), .Z(n6421) );
  XOR U6847 ( .A(n6577), .B(n6578), .Z(n6419) );
  ANDN U6848 ( .B(n6579), .A(n6580), .Z(n6577) );
  AND U6849 ( .A(a[4]), .B(b[22]), .Z(n6576) );
  XNOR U6850 ( .A(n6581), .B(n6424), .Z(n6426) );
  XOR U6851 ( .A(n6582), .B(n6583), .Z(n6424) );
  ANDN U6852 ( .B(n6584), .A(n6585), .Z(n6582) );
  AND U6853 ( .A(a[5]), .B(b[21]), .Z(n6581) );
  XNOR U6854 ( .A(n6586), .B(n6429), .Z(n6431) );
  XOR U6855 ( .A(n6587), .B(n6588), .Z(n6429) );
  ANDN U6856 ( .B(n6589), .A(n6590), .Z(n6587) );
  AND U6857 ( .A(a[6]), .B(b[20]), .Z(n6586) );
  XNOR U6858 ( .A(n6591), .B(n6434), .Z(n6436) );
  XOR U6859 ( .A(n6592), .B(n6593), .Z(n6434) );
  ANDN U6860 ( .B(n6594), .A(n6595), .Z(n6592) );
  AND U6861 ( .A(a[7]), .B(b[19]), .Z(n6591) );
  XNOR U6862 ( .A(n6596), .B(n6439), .Z(n6441) );
  XOR U6863 ( .A(n6597), .B(n6598), .Z(n6439) );
  ANDN U6864 ( .B(n6599), .A(n6600), .Z(n6597) );
  AND U6865 ( .A(a[8]), .B(b[18]), .Z(n6596) );
  XNOR U6866 ( .A(n6601), .B(n6444), .Z(n6446) );
  XOR U6867 ( .A(n6602), .B(n6603), .Z(n6444) );
  ANDN U6868 ( .B(n6604), .A(n6605), .Z(n6602) );
  AND U6869 ( .A(a[9]), .B(b[17]), .Z(n6601) );
  XNOR U6870 ( .A(n6606), .B(n6449), .Z(n6451) );
  XOR U6871 ( .A(n6607), .B(n6608), .Z(n6449) );
  ANDN U6872 ( .B(n6609), .A(n6610), .Z(n6607) );
  AND U6873 ( .A(a[10]), .B(b[16]), .Z(n6606) );
  XNOR U6874 ( .A(n6611), .B(n6454), .Z(n6456) );
  XOR U6875 ( .A(n6612), .B(n6613), .Z(n6454) );
  ANDN U6876 ( .B(n6614), .A(n6615), .Z(n6612) );
  AND U6877 ( .A(a[11]), .B(b[15]), .Z(n6611) );
  XNOR U6878 ( .A(n6616), .B(n6459), .Z(n6461) );
  XOR U6879 ( .A(n6617), .B(n6618), .Z(n6459) );
  ANDN U6880 ( .B(n6619), .A(n6620), .Z(n6617) );
  AND U6881 ( .A(a[12]), .B(b[14]), .Z(n6616) );
  XNOR U6882 ( .A(n6621), .B(n6464), .Z(n6466) );
  XOR U6883 ( .A(n6622), .B(n6623), .Z(n6464) );
  ANDN U6884 ( .B(n6624), .A(n6625), .Z(n6622) );
  AND U6885 ( .A(b[13]), .B(a[13]), .Z(n6621) );
  XNOR U6886 ( .A(n6626), .B(n6469), .Z(n6471) );
  XOR U6887 ( .A(n6627), .B(n6628), .Z(n6469) );
  ANDN U6888 ( .B(n6629), .A(n6630), .Z(n6627) );
  AND U6889 ( .A(a[14]), .B(b[12]), .Z(n6626) );
  XNOR U6890 ( .A(n6631), .B(n6474), .Z(n6476) );
  XOR U6891 ( .A(n6632), .B(n6633), .Z(n6474) );
  ANDN U6892 ( .B(n6634), .A(n6635), .Z(n6632) );
  AND U6893 ( .A(b[11]), .B(a[15]), .Z(n6631) );
  XNOR U6894 ( .A(n6636), .B(n6479), .Z(n6481) );
  XOR U6895 ( .A(n6637), .B(n6638), .Z(n6479) );
  ANDN U6896 ( .B(n6639), .A(n6640), .Z(n6637) );
  AND U6897 ( .A(a[16]), .B(b[10]), .Z(n6636) );
  XNOR U6898 ( .A(n6641), .B(n6484), .Z(n6486) );
  XOR U6899 ( .A(n6642), .B(n6643), .Z(n6484) );
  ANDN U6900 ( .B(n6644), .A(n6645), .Z(n6642) );
  AND U6901 ( .A(b[9]), .B(a[17]), .Z(n6641) );
  XNOR U6902 ( .A(n6646), .B(n6489), .Z(n6491) );
  XOR U6903 ( .A(n6647), .B(n6648), .Z(n6489) );
  ANDN U6904 ( .B(n6649), .A(n6650), .Z(n6647) );
  AND U6905 ( .A(a[18]), .B(b[8]), .Z(n6646) );
  XNOR U6906 ( .A(n6651), .B(n6494), .Z(n6496) );
  XOR U6907 ( .A(n6652), .B(n6653), .Z(n6494) );
  ANDN U6908 ( .B(n6654), .A(n6655), .Z(n6652) );
  AND U6909 ( .A(b[7]), .B(a[19]), .Z(n6651) );
  XNOR U6910 ( .A(n6656), .B(n6499), .Z(n6501) );
  XOR U6911 ( .A(n6657), .B(n6658), .Z(n6499) );
  ANDN U6912 ( .B(n6659), .A(n6660), .Z(n6657) );
  AND U6913 ( .A(b[6]), .B(a[20]), .Z(n6656) );
  XNOR U6914 ( .A(n6661), .B(n6504), .Z(n6506) );
  XOR U6915 ( .A(n6662), .B(n6663), .Z(n6504) );
  ANDN U6916 ( .B(n6664), .A(n6665), .Z(n6662) );
  AND U6917 ( .A(b[5]), .B(a[21]), .Z(n6661) );
  XNOR U6918 ( .A(n6666), .B(n6509), .Z(n6511) );
  XOR U6919 ( .A(n6667), .B(n6668), .Z(n6509) );
  ANDN U6920 ( .B(n6669), .A(n6670), .Z(n6667) );
  AND U6921 ( .A(b[4]), .B(a[22]), .Z(n6666) );
  XNOR U6922 ( .A(n6671), .B(n6672), .Z(n6523) );
  NANDN U6923 ( .A(n6673), .B(n6674), .Z(n6672) );
  XNOR U6924 ( .A(n6675), .B(n6514), .Z(n6516) );
  XNOR U6925 ( .A(n6676), .B(n6677), .Z(n6514) );
  AND U6926 ( .A(n6678), .B(n6679), .Z(n6676) );
  AND U6927 ( .A(b[3]), .B(a[23]), .Z(n6675) );
  NAND U6928 ( .A(a[26]), .B(b[0]), .Z(n6375) );
  IV U6929 ( .A(n6527), .Z(n6530) );
  XOR U6930 ( .A(n6680), .B(n6681), .Z(n6527) );
  ANDN U6931 ( .B(n6682), .A(n6683), .Z(n6680) );
  XNOR U6932 ( .A(n6682), .B(n6683), .Z(c[57]) );
  XNOR U6933 ( .A(sreg[89]), .B(n6684), .Z(n6683) );
  XNOR U6934 ( .A(n6684), .B(n6685), .Z(n6682) );
  XOR U6935 ( .A(n6535), .B(n6536), .Z(n6685) );
  XNOR U6936 ( .A(n6673), .B(n6674), .Z(n6536) );
  XOR U6937 ( .A(n6671), .B(n6686), .Z(n6674) );
  NAND U6938 ( .A(a[24]), .B(b[1]), .Z(n6686) );
  XOR U6939 ( .A(n6679), .B(n6687), .Z(n6673) );
  XOR U6940 ( .A(n6671), .B(n6678), .Z(n6687) );
  XNOR U6941 ( .A(n6688), .B(n6677), .Z(n6678) );
  AND U6942 ( .A(b[2]), .B(a[23]), .Z(n6688) );
  NANDN U6943 ( .A(n6689), .B(n6690), .Z(n6671) );
  XOR U6944 ( .A(n6677), .B(n6669), .Z(n6691) );
  XNOR U6945 ( .A(n6668), .B(n6664), .Z(n6692) );
  XNOR U6946 ( .A(n6663), .B(n6659), .Z(n6693) );
  XNOR U6947 ( .A(n6658), .B(n6654), .Z(n6694) );
  XNOR U6948 ( .A(n6653), .B(n6649), .Z(n6695) );
  XNOR U6949 ( .A(n6648), .B(n6644), .Z(n6696) );
  XNOR U6950 ( .A(n6643), .B(n6639), .Z(n6697) );
  XNOR U6951 ( .A(n6638), .B(n6634), .Z(n6698) );
  XNOR U6952 ( .A(n6633), .B(n6629), .Z(n6699) );
  XNOR U6953 ( .A(n6628), .B(n6624), .Z(n6700) );
  XNOR U6954 ( .A(n6623), .B(n6619), .Z(n6701) );
  XNOR U6955 ( .A(n6618), .B(n6614), .Z(n6702) );
  XNOR U6956 ( .A(n6613), .B(n6609), .Z(n6703) );
  XNOR U6957 ( .A(n6608), .B(n6604), .Z(n6704) );
  XNOR U6958 ( .A(n6603), .B(n6599), .Z(n6705) );
  XNOR U6959 ( .A(n6598), .B(n6594), .Z(n6706) );
  XNOR U6960 ( .A(n6593), .B(n6589), .Z(n6707) );
  XNOR U6961 ( .A(n6588), .B(n6584), .Z(n6708) );
  XNOR U6962 ( .A(n6583), .B(n6579), .Z(n6709) );
  XNOR U6963 ( .A(n6578), .B(n6574), .Z(n6710) );
  XNOR U6964 ( .A(n6573), .B(n6569), .Z(n6711) );
  XNOR U6965 ( .A(n6568), .B(n6564), .Z(n6712) );
  XOR U6966 ( .A(n6713), .B(n6563), .Z(n6564) );
  AND U6967 ( .A(a[0]), .B(b[25]), .Z(n6713) );
  XNOR U6968 ( .A(n6714), .B(n6563), .Z(n6565) );
  XNOR U6969 ( .A(n6715), .B(n6716), .Z(n6563) );
  ANDN U6970 ( .B(n6717), .A(n6718), .Z(n6715) );
  AND U6971 ( .A(a[1]), .B(b[24]), .Z(n6714) );
  XNOR U6972 ( .A(n6719), .B(n6568), .Z(n6570) );
  XOR U6973 ( .A(n6720), .B(n6721), .Z(n6568) );
  ANDN U6974 ( .B(n6722), .A(n6723), .Z(n6720) );
  AND U6975 ( .A(a[2]), .B(b[23]), .Z(n6719) );
  XNOR U6976 ( .A(n6724), .B(n6573), .Z(n6575) );
  XOR U6977 ( .A(n6725), .B(n6726), .Z(n6573) );
  ANDN U6978 ( .B(n6727), .A(n6728), .Z(n6725) );
  AND U6979 ( .A(a[3]), .B(b[22]), .Z(n6724) );
  XNOR U6980 ( .A(n6729), .B(n6578), .Z(n6580) );
  XOR U6981 ( .A(n6730), .B(n6731), .Z(n6578) );
  ANDN U6982 ( .B(n6732), .A(n6733), .Z(n6730) );
  AND U6983 ( .A(a[4]), .B(b[21]), .Z(n6729) );
  XNOR U6984 ( .A(n6734), .B(n6583), .Z(n6585) );
  XOR U6985 ( .A(n6735), .B(n6736), .Z(n6583) );
  ANDN U6986 ( .B(n6737), .A(n6738), .Z(n6735) );
  AND U6987 ( .A(a[5]), .B(b[20]), .Z(n6734) );
  XNOR U6988 ( .A(n6739), .B(n6588), .Z(n6590) );
  XOR U6989 ( .A(n6740), .B(n6741), .Z(n6588) );
  ANDN U6990 ( .B(n6742), .A(n6743), .Z(n6740) );
  AND U6991 ( .A(a[6]), .B(b[19]), .Z(n6739) );
  XNOR U6992 ( .A(n6744), .B(n6593), .Z(n6595) );
  XOR U6993 ( .A(n6745), .B(n6746), .Z(n6593) );
  ANDN U6994 ( .B(n6747), .A(n6748), .Z(n6745) );
  AND U6995 ( .A(a[7]), .B(b[18]), .Z(n6744) );
  XNOR U6996 ( .A(n6749), .B(n6598), .Z(n6600) );
  XOR U6997 ( .A(n6750), .B(n6751), .Z(n6598) );
  ANDN U6998 ( .B(n6752), .A(n6753), .Z(n6750) );
  AND U6999 ( .A(a[8]), .B(b[17]), .Z(n6749) );
  XNOR U7000 ( .A(n6754), .B(n6603), .Z(n6605) );
  XOR U7001 ( .A(n6755), .B(n6756), .Z(n6603) );
  ANDN U7002 ( .B(n6757), .A(n6758), .Z(n6755) );
  AND U7003 ( .A(a[9]), .B(b[16]), .Z(n6754) );
  XNOR U7004 ( .A(n6759), .B(n6608), .Z(n6610) );
  XOR U7005 ( .A(n6760), .B(n6761), .Z(n6608) );
  ANDN U7006 ( .B(n6762), .A(n6763), .Z(n6760) );
  AND U7007 ( .A(a[10]), .B(b[15]), .Z(n6759) );
  XNOR U7008 ( .A(n6764), .B(n6613), .Z(n6615) );
  XOR U7009 ( .A(n6765), .B(n6766), .Z(n6613) );
  ANDN U7010 ( .B(n6767), .A(n6768), .Z(n6765) );
  AND U7011 ( .A(a[11]), .B(b[14]), .Z(n6764) );
  XNOR U7012 ( .A(n6769), .B(n6618), .Z(n6620) );
  XOR U7013 ( .A(n6770), .B(n6771), .Z(n6618) );
  ANDN U7014 ( .B(n6772), .A(n6773), .Z(n6770) );
  AND U7015 ( .A(a[12]), .B(b[13]), .Z(n6769) );
  XNOR U7016 ( .A(n6774), .B(n6623), .Z(n6625) );
  XOR U7017 ( .A(n6775), .B(n6776), .Z(n6623) );
  ANDN U7018 ( .B(n6777), .A(n6778), .Z(n6775) );
  AND U7019 ( .A(b[12]), .B(a[13]), .Z(n6774) );
  XNOR U7020 ( .A(n6779), .B(n6628), .Z(n6630) );
  XOR U7021 ( .A(n6780), .B(n6781), .Z(n6628) );
  ANDN U7022 ( .B(n6782), .A(n6783), .Z(n6780) );
  AND U7023 ( .A(a[14]), .B(b[11]), .Z(n6779) );
  XNOR U7024 ( .A(n6784), .B(n6633), .Z(n6635) );
  XOR U7025 ( .A(n6785), .B(n6786), .Z(n6633) );
  ANDN U7026 ( .B(n6787), .A(n6788), .Z(n6785) );
  AND U7027 ( .A(b[10]), .B(a[15]), .Z(n6784) );
  XNOR U7028 ( .A(n6789), .B(n6638), .Z(n6640) );
  XOR U7029 ( .A(n6790), .B(n6791), .Z(n6638) );
  ANDN U7030 ( .B(n6792), .A(n6793), .Z(n6790) );
  AND U7031 ( .A(a[16]), .B(b[9]), .Z(n6789) );
  XNOR U7032 ( .A(n6794), .B(n6643), .Z(n6645) );
  XOR U7033 ( .A(n6795), .B(n6796), .Z(n6643) );
  ANDN U7034 ( .B(n6797), .A(n6798), .Z(n6795) );
  AND U7035 ( .A(b[8]), .B(a[17]), .Z(n6794) );
  XNOR U7036 ( .A(n6799), .B(n6648), .Z(n6650) );
  XOR U7037 ( .A(n6800), .B(n6801), .Z(n6648) );
  ANDN U7038 ( .B(n6802), .A(n6803), .Z(n6800) );
  AND U7039 ( .A(a[18]), .B(b[7]), .Z(n6799) );
  XNOR U7040 ( .A(n6804), .B(n6653), .Z(n6655) );
  XOR U7041 ( .A(n6805), .B(n6806), .Z(n6653) );
  ANDN U7042 ( .B(n6807), .A(n6808), .Z(n6805) );
  AND U7043 ( .A(b[6]), .B(a[19]), .Z(n6804) );
  XNOR U7044 ( .A(n6809), .B(n6658), .Z(n6660) );
  XOR U7045 ( .A(n6810), .B(n6811), .Z(n6658) );
  ANDN U7046 ( .B(n6812), .A(n6813), .Z(n6810) );
  AND U7047 ( .A(b[5]), .B(a[20]), .Z(n6809) );
  XNOR U7048 ( .A(n6814), .B(n6663), .Z(n6665) );
  XOR U7049 ( .A(n6815), .B(n6816), .Z(n6663) );
  ANDN U7050 ( .B(n6817), .A(n6818), .Z(n6815) );
  AND U7051 ( .A(b[4]), .B(a[21]), .Z(n6814) );
  XNOR U7052 ( .A(n6819), .B(n6820), .Z(n6677) );
  NANDN U7053 ( .A(n6821), .B(n6822), .Z(n6820) );
  XNOR U7054 ( .A(n6823), .B(n6668), .Z(n6670) );
  XNOR U7055 ( .A(n6824), .B(n6825), .Z(n6668) );
  AND U7056 ( .A(n6826), .B(n6827), .Z(n6824) );
  AND U7057 ( .A(b[3]), .B(a[22]), .Z(n6823) );
  NAND U7058 ( .A(a[25]), .B(b[0]), .Z(n6535) );
  IV U7059 ( .A(n6681), .Z(n6684) );
  XOR U7060 ( .A(n6828), .B(n6829), .Z(n6681) );
  ANDN U7061 ( .B(n6830), .A(n6831), .Z(n6828) );
  XNOR U7062 ( .A(n6830), .B(n6831), .Z(c[56]) );
  XNOR U7063 ( .A(sreg[88]), .B(n6832), .Z(n6831) );
  XNOR U7064 ( .A(n6832), .B(n6833), .Z(n6830) );
  XOR U7065 ( .A(n6689), .B(n6690), .Z(n6833) );
  XNOR U7066 ( .A(n6821), .B(n6822), .Z(n6690) );
  XOR U7067 ( .A(n6819), .B(n6834), .Z(n6822) );
  NAND U7068 ( .A(b[1]), .B(a[23]), .Z(n6834) );
  XOR U7069 ( .A(n6827), .B(n6835), .Z(n6821) );
  XOR U7070 ( .A(n6819), .B(n6826), .Z(n6835) );
  XNOR U7071 ( .A(n6836), .B(n6825), .Z(n6826) );
  AND U7072 ( .A(b[2]), .B(a[22]), .Z(n6836) );
  NANDN U7073 ( .A(n6837), .B(n6838), .Z(n6819) );
  XOR U7074 ( .A(n6825), .B(n6817), .Z(n6839) );
  XNOR U7075 ( .A(n6816), .B(n6812), .Z(n6840) );
  XNOR U7076 ( .A(n6811), .B(n6807), .Z(n6841) );
  XNOR U7077 ( .A(n6806), .B(n6802), .Z(n6842) );
  XNOR U7078 ( .A(n6801), .B(n6797), .Z(n6843) );
  XNOR U7079 ( .A(n6796), .B(n6792), .Z(n6844) );
  XNOR U7080 ( .A(n6791), .B(n6787), .Z(n6845) );
  XNOR U7081 ( .A(n6786), .B(n6782), .Z(n6846) );
  XNOR U7082 ( .A(n6781), .B(n6777), .Z(n6847) );
  XNOR U7083 ( .A(n6776), .B(n6772), .Z(n6848) );
  XNOR U7084 ( .A(n6771), .B(n6767), .Z(n6849) );
  XNOR U7085 ( .A(n6766), .B(n6762), .Z(n6850) );
  XNOR U7086 ( .A(n6761), .B(n6757), .Z(n6851) );
  XNOR U7087 ( .A(n6756), .B(n6752), .Z(n6852) );
  XNOR U7088 ( .A(n6751), .B(n6747), .Z(n6853) );
  XNOR U7089 ( .A(n6746), .B(n6742), .Z(n6854) );
  XNOR U7090 ( .A(n6741), .B(n6737), .Z(n6855) );
  XNOR U7091 ( .A(n6736), .B(n6732), .Z(n6856) );
  XNOR U7092 ( .A(n6731), .B(n6727), .Z(n6857) );
  XNOR U7093 ( .A(n6726), .B(n6722), .Z(n6858) );
  XNOR U7094 ( .A(n6721), .B(n6717), .Z(n6859) );
  XNOR U7095 ( .A(n6860), .B(n6716), .Z(n6717) );
  AND U7096 ( .A(a[0]), .B(b[24]), .Z(n6860) );
  XOR U7097 ( .A(n6861), .B(n6716), .Z(n6718) );
  XNOR U7098 ( .A(n6862), .B(n6863), .Z(n6716) );
  ANDN U7099 ( .B(n6864), .A(n6865), .Z(n6862) );
  AND U7100 ( .A(a[1]), .B(b[23]), .Z(n6861) );
  XNOR U7101 ( .A(n6866), .B(n6721), .Z(n6723) );
  XOR U7102 ( .A(n6867), .B(n6868), .Z(n6721) );
  ANDN U7103 ( .B(n6869), .A(n6870), .Z(n6867) );
  AND U7104 ( .A(a[2]), .B(b[22]), .Z(n6866) );
  XNOR U7105 ( .A(n6871), .B(n6726), .Z(n6728) );
  XOR U7106 ( .A(n6872), .B(n6873), .Z(n6726) );
  ANDN U7107 ( .B(n6874), .A(n6875), .Z(n6872) );
  AND U7108 ( .A(a[3]), .B(b[21]), .Z(n6871) );
  XNOR U7109 ( .A(n6876), .B(n6731), .Z(n6733) );
  XOR U7110 ( .A(n6877), .B(n6878), .Z(n6731) );
  ANDN U7111 ( .B(n6879), .A(n6880), .Z(n6877) );
  AND U7112 ( .A(a[4]), .B(b[20]), .Z(n6876) );
  XNOR U7113 ( .A(n6881), .B(n6736), .Z(n6738) );
  XOR U7114 ( .A(n6882), .B(n6883), .Z(n6736) );
  ANDN U7115 ( .B(n6884), .A(n6885), .Z(n6882) );
  AND U7116 ( .A(a[5]), .B(b[19]), .Z(n6881) );
  XNOR U7117 ( .A(n6886), .B(n6741), .Z(n6743) );
  XOR U7118 ( .A(n6887), .B(n6888), .Z(n6741) );
  ANDN U7119 ( .B(n6889), .A(n6890), .Z(n6887) );
  AND U7120 ( .A(a[6]), .B(b[18]), .Z(n6886) );
  XNOR U7121 ( .A(n6891), .B(n6746), .Z(n6748) );
  XOR U7122 ( .A(n6892), .B(n6893), .Z(n6746) );
  ANDN U7123 ( .B(n6894), .A(n6895), .Z(n6892) );
  AND U7124 ( .A(a[7]), .B(b[17]), .Z(n6891) );
  XNOR U7125 ( .A(n6896), .B(n6751), .Z(n6753) );
  XOR U7126 ( .A(n6897), .B(n6898), .Z(n6751) );
  ANDN U7127 ( .B(n6899), .A(n6900), .Z(n6897) );
  AND U7128 ( .A(a[8]), .B(b[16]), .Z(n6896) );
  XNOR U7129 ( .A(n6901), .B(n6756), .Z(n6758) );
  XOR U7130 ( .A(n6902), .B(n6903), .Z(n6756) );
  ANDN U7131 ( .B(n6904), .A(n6905), .Z(n6902) );
  AND U7132 ( .A(a[9]), .B(b[15]), .Z(n6901) );
  XNOR U7133 ( .A(n6906), .B(n6761), .Z(n6763) );
  XOR U7134 ( .A(n6907), .B(n6908), .Z(n6761) );
  ANDN U7135 ( .B(n6909), .A(n6910), .Z(n6907) );
  AND U7136 ( .A(a[10]), .B(b[14]), .Z(n6906) );
  XNOR U7137 ( .A(n6911), .B(n6766), .Z(n6768) );
  XOR U7138 ( .A(n6912), .B(n6913), .Z(n6766) );
  ANDN U7139 ( .B(n6914), .A(n6915), .Z(n6912) );
  AND U7140 ( .A(a[11]), .B(b[13]), .Z(n6911) );
  XNOR U7141 ( .A(n6916), .B(n6771), .Z(n6773) );
  XOR U7142 ( .A(n6917), .B(n6918), .Z(n6771) );
  ANDN U7143 ( .B(n6919), .A(n6920), .Z(n6917) );
  AND U7144 ( .A(a[12]), .B(b[12]), .Z(n6916) );
  XNOR U7145 ( .A(n6921), .B(n6776), .Z(n6778) );
  XOR U7146 ( .A(n6922), .B(n6923), .Z(n6776) );
  ANDN U7147 ( .B(n6924), .A(n6925), .Z(n6922) );
  AND U7148 ( .A(b[11]), .B(a[13]), .Z(n6921) );
  XNOR U7149 ( .A(n6926), .B(n6781), .Z(n6783) );
  XOR U7150 ( .A(n6927), .B(n6928), .Z(n6781) );
  ANDN U7151 ( .B(n6929), .A(n6930), .Z(n6927) );
  AND U7152 ( .A(a[14]), .B(b[10]), .Z(n6926) );
  XNOR U7153 ( .A(n6931), .B(n6786), .Z(n6788) );
  XOR U7154 ( .A(n6932), .B(n6933), .Z(n6786) );
  ANDN U7155 ( .B(n6934), .A(n6935), .Z(n6932) );
  AND U7156 ( .A(b[9]), .B(a[15]), .Z(n6931) );
  XNOR U7157 ( .A(n6936), .B(n6791), .Z(n6793) );
  XOR U7158 ( .A(n6937), .B(n6938), .Z(n6791) );
  ANDN U7159 ( .B(n6939), .A(n6940), .Z(n6937) );
  AND U7160 ( .A(a[16]), .B(b[8]), .Z(n6936) );
  XNOR U7161 ( .A(n6941), .B(n6796), .Z(n6798) );
  XOR U7162 ( .A(n6942), .B(n6943), .Z(n6796) );
  ANDN U7163 ( .B(n6944), .A(n6945), .Z(n6942) );
  AND U7164 ( .A(b[7]), .B(a[17]), .Z(n6941) );
  XNOR U7165 ( .A(n6946), .B(n6801), .Z(n6803) );
  XOR U7166 ( .A(n6947), .B(n6948), .Z(n6801) );
  ANDN U7167 ( .B(n6949), .A(n6950), .Z(n6947) );
  AND U7168 ( .A(b[6]), .B(a[18]), .Z(n6946) );
  XNOR U7169 ( .A(n6951), .B(n6806), .Z(n6808) );
  XOR U7170 ( .A(n6952), .B(n6953), .Z(n6806) );
  ANDN U7171 ( .B(n6954), .A(n6955), .Z(n6952) );
  AND U7172 ( .A(b[5]), .B(a[19]), .Z(n6951) );
  XNOR U7173 ( .A(n6956), .B(n6811), .Z(n6813) );
  XOR U7174 ( .A(n6957), .B(n6958), .Z(n6811) );
  ANDN U7175 ( .B(n6959), .A(n6960), .Z(n6957) );
  AND U7176 ( .A(b[4]), .B(a[20]), .Z(n6956) );
  XNOR U7177 ( .A(n6961), .B(n6962), .Z(n6825) );
  NANDN U7178 ( .A(n6963), .B(n6964), .Z(n6962) );
  XNOR U7179 ( .A(n6965), .B(n6816), .Z(n6818) );
  XNOR U7180 ( .A(n6966), .B(n6967), .Z(n6816) );
  AND U7181 ( .A(n6968), .B(n6969), .Z(n6966) );
  AND U7182 ( .A(b[3]), .B(a[21]), .Z(n6965) );
  NAND U7183 ( .A(a[24]), .B(b[0]), .Z(n6689) );
  IV U7184 ( .A(n6829), .Z(n6832) );
  XOR U7185 ( .A(n6970), .B(n6971), .Z(n6829) );
  ANDN U7186 ( .B(n6972), .A(n6973), .Z(n6970) );
  XNOR U7187 ( .A(n6972), .B(n6973), .Z(c[55]) );
  XNOR U7188 ( .A(sreg[87]), .B(n6974), .Z(n6973) );
  XNOR U7189 ( .A(n6974), .B(n6975), .Z(n6972) );
  XOR U7190 ( .A(n6837), .B(n6838), .Z(n6975) );
  XNOR U7191 ( .A(n6963), .B(n6964), .Z(n6838) );
  XOR U7192 ( .A(n6961), .B(n6976), .Z(n6964) );
  NAND U7193 ( .A(a[22]), .B(b[1]), .Z(n6976) );
  XOR U7194 ( .A(n6969), .B(n6977), .Z(n6963) );
  XOR U7195 ( .A(n6961), .B(n6968), .Z(n6977) );
  XNOR U7196 ( .A(n6978), .B(n6967), .Z(n6968) );
  AND U7197 ( .A(b[2]), .B(a[21]), .Z(n6978) );
  NANDN U7198 ( .A(n6979), .B(n6980), .Z(n6961) );
  XOR U7199 ( .A(n6967), .B(n6959), .Z(n6981) );
  XNOR U7200 ( .A(n6958), .B(n6954), .Z(n6982) );
  XNOR U7201 ( .A(n6953), .B(n6949), .Z(n6983) );
  XNOR U7202 ( .A(n6948), .B(n6944), .Z(n6984) );
  XNOR U7203 ( .A(n6943), .B(n6939), .Z(n6985) );
  XNOR U7204 ( .A(n6938), .B(n6934), .Z(n6986) );
  XNOR U7205 ( .A(n6933), .B(n6929), .Z(n6987) );
  XNOR U7206 ( .A(n6928), .B(n6924), .Z(n6988) );
  XNOR U7207 ( .A(n6923), .B(n6919), .Z(n6989) );
  XNOR U7208 ( .A(n6918), .B(n6914), .Z(n6990) );
  XNOR U7209 ( .A(n6913), .B(n6909), .Z(n6991) );
  XNOR U7210 ( .A(n6908), .B(n6904), .Z(n6992) );
  XNOR U7211 ( .A(n6903), .B(n6899), .Z(n6993) );
  XNOR U7212 ( .A(n6898), .B(n6894), .Z(n6994) );
  XNOR U7213 ( .A(n6893), .B(n6889), .Z(n6995) );
  XNOR U7214 ( .A(n6888), .B(n6884), .Z(n6996) );
  XNOR U7215 ( .A(n6883), .B(n6879), .Z(n6997) );
  XNOR U7216 ( .A(n6878), .B(n6874), .Z(n6998) );
  XNOR U7217 ( .A(n6873), .B(n6869), .Z(n6999) );
  XNOR U7218 ( .A(n6868), .B(n6864), .Z(n7000) );
  XOR U7219 ( .A(n7001), .B(n6863), .Z(n6864) );
  AND U7220 ( .A(a[0]), .B(b[23]), .Z(n7001) );
  XNOR U7221 ( .A(n7002), .B(n6863), .Z(n6865) );
  XNOR U7222 ( .A(n7003), .B(n7004), .Z(n6863) );
  ANDN U7223 ( .B(n7005), .A(n7006), .Z(n7003) );
  AND U7224 ( .A(a[1]), .B(b[22]), .Z(n7002) );
  XNOR U7225 ( .A(n7007), .B(n6868), .Z(n6870) );
  XOR U7226 ( .A(n7008), .B(n7009), .Z(n6868) );
  ANDN U7227 ( .B(n7010), .A(n7011), .Z(n7008) );
  AND U7228 ( .A(a[2]), .B(b[21]), .Z(n7007) );
  XNOR U7229 ( .A(n7012), .B(n6873), .Z(n6875) );
  XOR U7230 ( .A(n7013), .B(n7014), .Z(n6873) );
  ANDN U7231 ( .B(n7015), .A(n7016), .Z(n7013) );
  AND U7232 ( .A(a[3]), .B(b[20]), .Z(n7012) );
  XNOR U7233 ( .A(n7017), .B(n6878), .Z(n6880) );
  XOR U7234 ( .A(n7018), .B(n7019), .Z(n6878) );
  ANDN U7235 ( .B(n7020), .A(n7021), .Z(n7018) );
  AND U7236 ( .A(a[4]), .B(b[19]), .Z(n7017) );
  XNOR U7237 ( .A(n7022), .B(n6883), .Z(n6885) );
  XOR U7238 ( .A(n7023), .B(n7024), .Z(n6883) );
  ANDN U7239 ( .B(n7025), .A(n7026), .Z(n7023) );
  AND U7240 ( .A(a[5]), .B(b[18]), .Z(n7022) );
  XNOR U7241 ( .A(n7027), .B(n6888), .Z(n6890) );
  XOR U7242 ( .A(n7028), .B(n7029), .Z(n6888) );
  ANDN U7243 ( .B(n7030), .A(n7031), .Z(n7028) );
  AND U7244 ( .A(a[6]), .B(b[17]), .Z(n7027) );
  XNOR U7245 ( .A(n7032), .B(n6893), .Z(n6895) );
  XOR U7246 ( .A(n7033), .B(n7034), .Z(n6893) );
  ANDN U7247 ( .B(n7035), .A(n7036), .Z(n7033) );
  AND U7248 ( .A(a[7]), .B(b[16]), .Z(n7032) );
  XNOR U7249 ( .A(n7037), .B(n6898), .Z(n6900) );
  XOR U7250 ( .A(n7038), .B(n7039), .Z(n6898) );
  ANDN U7251 ( .B(n7040), .A(n7041), .Z(n7038) );
  AND U7252 ( .A(a[8]), .B(b[15]), .Z(n7037) );
  XNOR U7253 ( .A(n7042), .B(n6903), .Z(n6905) );
  XOR U7254 ( .A(n7043), .B(n7044), .Z(n6903) );
  ANDN U7255 ( .B(n7045), .A(n7046), .Z(n7043) );
  AND U7256 ( .A(a[9]), .B(b[14]), .Z(n7042) );
  XNOR U7257 ( .A(n7047), .B(n6908), .Z(n6910) );
  XOR U7258 ( .A(n7048), .B(n7049), .Z(n6908) );
  ANDN U7259 ( .B(n7050), .A(n7051), .Z(n7048) );
  AND U7260 ( .A(a[10]), .B(b[13]), .Z(n7047) );
  XNOR U7261 ( .A(n7052), .B(n6913), .Z(n6915) );
  XOR U7262 ( .A(n7053), .B(n7054), .Z(n6913) );
  ANDN U7263 ( .B(n7055), .A(n7056), .Z(n7053) );
  AND U7264 ( .A(a[11]), .B(b[12]), .Z(n7052) );
  XNOR U7265 ( .A(n7057), .B(n6918), .Z(n6920) );
  XOR U7266 ( .A(n7058), .B(n7059), .Z(n6918) );
  ANDN U7267 ( .B(n7060), .A(n7061), .Z(n7058) );
  AND U7268 ( .A(a[12]), .B(b[11]), .Z(n7057) );
  XNOR U7269 ( .A(n7062), .B(n6923), .Z(n6925) );
  XOR U7270 ( .A(n7063), .B(n7064), .Z(n6923) );
  ANDN U7271 ( .B(n7065), .A(n7066), .Z(n7063) );
  AND U7272 ( .A(b[10]), .B(a[13]), .Z(n7062) );
  XNOR U7273 ( .A(n7067), .B(n6928), .Z(n6930) );
  XOR U7274 ( .A(n7068), .B(n7069), .Z(n6928) );
  ANDN U7275 ( .B(n7070), .A(n7071), .Z(n7068) );
  AND U7276 ( .A(a[14]), .B(b[9]), .Z(n7067) );
  XNOR U7277 ( .A(n7072), .B(n6933), .Z(n6935) );
  XOR U7278 ( .A(n7073), .B(n7074), .Z(n6933) );
  ANDN U7279 ( .B(n7075), .A(n7076), .Z(n7073) );
  AND U7280 ( .A(b[8]), .B(a[15]), .Z(n7072) );
  XNOR U7281 ( .A(n7077), .B(n6938), .Z(n6940) );
  XOR U7282 ( .A(n7078), .B(n7079), .Z(n6938) );
  ANDN U7283 ( .B(n7080), .A(n7081), .Z(n7078) );
  AND U7284 ( .A(a[16]), .B(b[7]), .Z(n7077) );
  XNOR U7285 ( .A(n7082), .B(n6943), .Z(n6945) );
  XOR U7286 ( .A(n7083), .B(n7084), .Z(n6943) );
  ANDN U7287 ( .B(n7085), .A(n7086), .Z(n7083) );
  AND U7288 ( .A(b[6]), .B(a[17]), .Z(n7082) );
  XNOR U7289 ( .A(n7087), .B(n6948), .Z(n6950) );
  XOR U7290 ( .A(n7088), .B(n7089), .Z(n6948) );
  ANDN U7291 ( .B(n7090), .A(n7091), .Z(n7088) );
  AND U7292 ( .A(b[5]), .B(a[18]), .Z(n7087) );
  XNOR U7293 ( .A(n7092), .B(n6953), .Z(n6955) );
  XOR U7294 ( .A(n7093), .B(n7094), .Z(n6953) );
  ANDN U7295 ( .B(n7095), .A(n7096), .Z(n7093) );
  AND U7296 ( .A(b[4]), .B(a[19]), .Z(n7092) );
  XNOR U7297 ( .A(n7097), .B(n7098), .Z(n6967) );
  NANDN U7298 ( .A(n7099), .B(n7100), .Z(n7098) );
  XNOR U7299 ( .A(n7101), .B(n6958), .Z(n6960) );
  XNOR U7300 ( .A(n7102), .B(n7103), .Z(n6958) );
  AND U7301 ( .A(n7104), .B(n7105), .Z(n7102) );
  AND U7302 ( .A(b[3]), .B(a[20]), .Z(n7101) );
  NAND U7303 ( .A(a[23]), .B(b[0]), .Z(n6837) );
  IV U7304 ( .A(n6971), .Z(n6974) );
  XOR U7305 ( .A(n7106), .B(n7107), .Z(n6971) );
  ANDN U7306 ( .B(n7108), .A(n7109), .Z(n7106) );
  XNOR U7307 ( .A(n7108), .B(n7109), .Z(c[54]) );
  XNOR U7308 ( .A(sreg[86]), .B(n7110), .Z(n7109) );
  XNOR U7309 ( .A(n7110), .B(n7111), .Z(n7108) );
  XOR U7310 ( .A(n6979), .B(n6980), .Z(n7111) );
  XNOR U7311 ( .A(n7099), .B(n7100), .Z(n6980) );
  XOR U7312 ( .A(n7097), .B(n7112), .Z(n7100) );
  NAND U7313 ( .A(b[1]), .B(a[21]), .Z(n7112) );
  XOR U7314 ( .A(n7105), .B(n7113), .Z(n7099) );
  XOR U7315 ( .A(n7097), .B(n7104), .Z(n7113) );
  XNOR U7316 ( .A(n7114), .B(n7103), .Z(n7104) );
  AND U7317 ( .A(b[2]), .B(a[20]), .Z(n7114) );
  NANDN U7318 ( .A(n7115), .B(n7116), .Z(n7097) );
  XOR U7319 ( .A(n7103), .B(n7095), .Z(n7117) );
  XNOR U7320 ( .A(n7094), .B(n7090), .Z(n7118) );
  XNOR U7321 ( .A(n7089), .B(n7085), .Z(n7119) );
  XNOR U7322 ( .A(n7084), .B(n7080), .Z(n7120) );
  XNOR U7323 ( .A(n7079), .B(n7075), .Z(n7121) );
  XNOR U7324 ( .A(n7074), .B(n7070), .Z(n7122) );
  XNOR U7325 ( .A(n7069), .B(n7065), .Z(n7123) );
  XNOR U7326 ( .A(n7064), .B(n7060), .Z(n7124) );
  XNOR U7327 ( .A(n7059), .B(n7055), .Z(n7125) );
  XNOR U7328 ( .A(n7054), .B(n7050), .Z(n7126) );
  XNOR U7329 ( .A(n7049), .B(n7045), .Z(n7127) );
  XNOR U7330 ( .A(n7044), .B(n7040), .Z(n7128) );
  XNOR U7331 ( .A(n7039), .B(n7035), .Z(n7129) );
  XNOR U7332 ( .A(n7034), .B(n7030), .Z(n7130) );
  XNOR U7333 ( .A(n7029), .B(n7025), .Z(n7131) );
  XNOR U7334 ( .A(n7024), .B(n7020), .Z(n7132) );
  XNOR U7335 ( .A(n7019), .B(n7015), .Z(n7133) );
  XNOR U7336 ( .A(n7014), .B(n7010), .Z(n7134) );
  XNOR U7337 ( .A(n7009), .B(n7005), .Z(n7135) );
  XNOR U7338 ( .A(n7136), .B(n7004), .Z(n7005) );
  AND U7339 ( .A(a[0]), .B(b[22]), .Z(n7136) );
  XOR U7340 ( .A(n7137), .B(n7004), .Z(n7006) );
  XNOR U7341 ( .A(n7138), .B(n7139), .Z(n7004) );
  ANDN U7342 ( .B(n7140), .A(n7141), .Z(n7138) );
  AND U7343 ( .A(a[1]), .B(b[21]), .Z(n7137) );
  XNOR U7344 ( .A(n7142), .B(n7009), .Z(n7011) );
  XOR U7345 ( .A(n7143), .B(n7144), .Z(n7009) );
  ANDN U7346 ( .B(n7145), .A(n7146), .Z(n7143) );
  AND U7347 ( .A(a[2]), .B(b[20]), .Z(n7142) );
  XNOR U7348 ( .A(n7147), .B(n7014), .Z(n7016) );
  XOR U7349 ( .A(n7148), .B(n7149), .Z(n7014) );
  ANDN U7350 ( .B(n7150), .A(n7151), .Z(n7148) );
  AND U7351 ( .A(a[3]), .B(b[19]), .Z(n7147) );
  XNOR U7352 ( .A(n7152), .B(n7019), .Z(n7021) );
  XOR U7353 ( .A(n7153), .B(n7154), .Z(n7019) );
  ANDN U7354 ( .B(n7155), .A(n7156), .Z(n7153) );
  AND U7355 ( .A(a[4]), .B(b[18]), .Z(n7152) );
  XNOR U7356 ( .A(n7157), .B(n7024), .Z(n7026) );
  XOR U7357 ( .A(n7158), .B(n7159), .Z(n7024) );
  ANDN U7358 ( .B(n7160), .A(n7161), .Z(n7158) );
  AND U7359 ( .A(a[5]), .B(b[17]), .Z(n7157) );
  XNOR U7360 ( .A(n7162), .B(n7029), .Z(n7031) );
  XOR U7361 ( .A(n7163), .B(n7164), .Z(n7029) );
  ANDN U7362 ( .B(n7165), .A(n7166), .Z(n7163) );
  AND U7363 ( .A(a[6]), .B(b[16]), .Z(n7162) );
  XNOR U7364 ( .A(n7167), .B(n7034), .Z(n7036) );
  XOR U7365 ( .A(n7168), .B(n7169), .Z(n7034) );
  ANDN U7366 ( .B(n7170), .A(n7171), .Z(n7168) );
  AND U7367 ( .A(a[7]), .B(b[15]), .Z(n7167) );
  XNOR U7368 ( .A(n7172), .B(n7039), .Z(n7041) );
  XOR U7369 ( .A(n7173), .B(n7174), .Z(n7039) );
  ANDN U7370 ( .B(n7175), .A(n7176), .Z(n7173) );
  AND U7371 ( .A(a[8]), .B(b[14]), .Z(n7172) );
  XNOR U7372 ( .A(n7177), .B(n7044), .Z(n7046) );
  XOR U7373 ( .A(n7178), .B(n7179), .Z(n7044) );
  ANDN U7374 ( .B(n7180), .A(n7181), .Z(n7178) );
  AND U7375 ( .A(a[9]), .B(b[13]), .Z(n7177) );
  XNOR U7376 ( .A(n7182), .B(n7049), .Z(n7051) );
  XOR U7377 ( .A(n7183), .B(n7184), .Z(n7049) );
  ANDN U7378 ( .B(n7185), .A(n7186), .Z(n7183) );
  AND U7379 ( .A(a[10]), .B(b[12]), .Z(n7182) );
  XNOR U7380 ( .A(n7187), .B(n7054), .Z(n7056) );
  XOR U7381 ( .A(n7188), .B(n7189), .Z(n7054) );
  ANDN U7382 ( .B(n7190), .A(n7191), .Z(n7188) );
  AND U7383 ( .A(b[11]), .B(a[11]), .Z(n7187) );
  XNOR U7384 ( .A(n7192), .B(n7059), .Z(n7061) );
  XOR U7385 ( .A(n7193), .B(n7194), .Z(n7059) );
  ANDN U7386 ( .B(n7195), .A(n7196), .Z(n7193) );
  AND U7387 ( .A(a[12]), .B(b[10]), .Z(n7192) );
  XNOR U7388 ( .A(n7197), .B(n7064), .Z(n7066) );
  XOR U7389 ( .A(n7198), .B(n7199), .Z(n7064) );
  ANDN U7390 ( .B(n7200), .A(n7201), .Z(n7198) );
  AND U7391 ( .A(b[9]), .B(a[13]), .Z(n7197) );
  XNOR U7392 ( .A(n7202), .B(n7069), .Z(n7071) );
  XOR U7393 ( .A(n7203), .B(n7204), .Z(n7069) );
  ANDN U7394 ( .B(n7205), .A(n7206), .Z(n7203) );
  AND U7395 ( .A(a[14]), .B(b[8]), .Z(n7202) );
  XNOR U7396 ( .A(n7207), .B(n7074), .Z(n7076) );
  XOR U7397 ( .A(n7208), .B(n7209), .Z(n7074) );
  ANDN U7398 ( .B(n7210), .A(n7211), .Z(n7208) );
  AND U7399 ( .A(b[7]), .B(a[15]), .Z(n7207) );
  XNOR U7400 ( .A(n7212), .B(n7079), .Z(n7081) );
  XOR U7401 ( .A(n7213), .B(n7214), .Z(n7079) );
  ANDN U7402 ( .B(n7215), .A(n7216), .Z(n7213) );
  AND U7403 ( .A(b[6]), .B(a[16]), .Z(n7212) );
  XNOR U7404 ( .A(n7217), .B(n7084), .Z(n7086) );
  XOR U7405 ( .A(n7218), .B(n7219), .Z(n7084) );
  ANDN U7406 ( .B(n7220), .A(n7221), .Z(n7218) );
  AND U7407 ( .A(b[5]), .B(a[17]), .Z(n7217) );
  XNOR U7408 ( .A(n7222), .B(n7089), .Z(n7091) );
  XOR U7409 ( .A(n7223), .B(n7224), .Z(n7089) );
  ANDN U7410 ( .B(n7225), .A(n7226), .Z(n7223) );
  AND U7411 ( .A(b[4]), .B(a[18]), .Z(n7222) );
  XNOR U7412 ( .A(n7227), .B(n7228), .Z(n7103) );
  NANDN U7413 ( .A(n7229), .B(n7230), .Z(n7228) );
  XNOR U7414 ( .A(n7231), .B(n7094), .Z(n7096) );
  XNOR U7415 ( .A(n7232), .B(n7233), .Z(n7094) );
  AND U7416 ( .A(n7234), .B(n7235), .Z(n7232) );
  AND U7417 ( .A(b[3]), .B(a[19]), .Z(n7231) );
  NAND U7418 ( .A(a[22]), .B(b[0]), .Z(n6979) );
  IV U7419 ( .A(n7107), .Z(n7110) );
  XOR U7420 ( .A(n7236), .B(n7237), .Z(n7107) );
  ANDN U7421 ( .B(n7238), .A(n7239), .Z(n7236) );
  XNOR U7422 ( .A(n7238), .B(n7239), .Z(c[53]) );
  XNOR U7423 ( .A(sreg[85]), .B(n7240), .Z(n7239) );
  XNOR U7424 ( .A(n7240), .B(n7241), .Z(n7238) );
  XOR U7425 ( .A(n7115), .B(n7116), .Z(n7241) );
  XNOR U7426 ( .A(n7229), .B(n7230), .Z(n7116) );
  XOR U7427 ( .A(n7227), .B(n7242), .Z(n7230) );
  NAND U7428 ( .A(a[20]), .B(b[1]), .Z(n7242) );
  XOR U7429 ( .A(n7235), .B(n7243), .Z(n7229) );
  XOR U7430 ( .A(n7227), .B(n7234), .Z(n7243) );
  XNOR U7431 ( .A(n7244), .B(n7233), .Z(n7234) );
  AND U7432 ( .A(b[2]), .B(a[19]), .Z(n7244) );
  NANDN U7433 ( .A(n7245), .B(n7246), .Z(n7227) );
  XOR U7434 ( .A(n7233), .B(n7225), .Z(n7247) );
  XNOR U7435 ( .A(n7224), .B(n7220), .Z(n7248) );
  XNOR U7436 ( .A(n7219), .B(n7215), .Z(n7249) );
  XNOR U7437 ( .A(n7214), .B(n7210), .Z(n7250) );
  XNOR U7438 ( .A(n7209), .B(n7205), .Z(n7251) );
  XNOR U7439 ( .A(n7204), .B(n7200), .Z(n7252) );
  XNOR U7440 ( .A(n7199), .B(n7195), .Z(n7253) );
  XNOR U7441 ( .A(n7194), .B(n7190), .Z(n7254) );
  XNOR U7442 ( .A(n7189), .B(n7185), .Z(n7255) );
  XNOR U7443 ( .A(n7184), .B(n7180), .Z(n7256) );
  XNOR U7444 ( .A(n7179), .B(n7175), .Z(n7257) );
  XNOR U7445 ( .A(n7174), .B(n7170), .Z(n7258) );
  XNOR U7446 ( .A(n7169), .B(n7165), .Z(n7259) );
  XNOR U7447 ( .A(n7164), .B(n7160), .Z(n7260) );
  XNOR U7448 ( .A(n7159), .B(n7155), .Z(n7261) );
  XNOR U7449 ( .A(n7154), .B(n7150), .Z(n7262) );
  XNOR U7450 ( .A(n7149), .B(n7145), .Z(n7263) );
  XNOR U7451 ( .A(n7144), .B(n7140), .Z(n7264) );
  XOR U7452 ( .A(n7265), .B(n7139), .Z(n7140) );
  AND U7453 ( .A(a[0]), .B(b[21]), .Z(n7265) );
  XNOR U7454 ( .A(n7266), .B(n7139), .Z(n7141) );
  XNOR U7455 ( .A(n7267), .B(n7268), .Z(n7139) );
  ANDN U7456 ( .B(n7269), .A(n7270), .Z(n7267) );
  AND U7457 ( .A(a[1]), .B(b[20]), .Z(n7266) );
  XNOR U7458 ( .A(n7271), .B(n7144), .Z(n7146) );
  XOR U7459 ( .A(n7272), .B(n7273), .Z(n7144) );
  ANDN U7460 ( .B(n7274), .A(n7275), .Z(n7272) );
  AND U7461 ( .A(a[2]), .B(b[19]), .Z(n7271) );
  XNOR U7462 ( .A(n7276), .B(n7149), .Z(n7151) );
  XOR U7463 ( .A(n7277), .B(n7278), .Z(n7149) );
  ANDN U7464 ( .B(n7279), .A(n7280), .Z(n7277) );
  AND U7465 ( .A(a[3]), .B(b[18]), .Z(n7276) );
  XNOR U7466 ( .A(n7281), .B(n7154), .Z(n7156) );
  XOR U7467 ( .A(n7282), .B(n7283), .Z(n7154) );
  ANDN U7468 ( .B(n7284), .A(n7285), .Z(n7282) );
  AND U7469 ( .A(a[4]), .B(b[17]), .Z(n7281) );
  XNOR U7470 ( .A(n7286), .B(n7159), .Z(n7161) );
  XOR U7471 ( .A(n7287), .B(n7288), .Z(n7159) );
  ANDN U7472 ( .B(n7289), .A(n7290), .Z(n7287) );
  AND U7473 ( .A(a[5]), .B(b[16]), .Z(n7286) );
  XNOR U7474 ( .A(n7291), .B(n7164), .Z(n7166) );
  XOR U7475 ( .A(n7292), .B(n7293), .Z(n7164) );
  ANDN U7476 ( .B(n7294), .A(n7295), .Z(n7292) );
  AND U7477 ( .A(a[6]), .B(b[15]), .Z(n7291) );
  XNOR U7478 ( .A(n7296), .B(n7169), .Z(n7171) );
  XOR U7479 ( .A(n7297), .B(n7298), .Z(n7169) );
  ANDN U7480 ( .B(n7299), .A(n7300), .Z(n7297) );
  AND U7481 ( .A(a[7]), .B(b[14]), .Z(n7296) );
  XNOR U7482 ( .A(n7301), .B(n7174), .Z(n7176) );
  XOR U7483 ( .A(n7302), .B(n7303), .Z(n7174) );
  ANDN U7484 ( .B(n7304), .A(n7305), .Z(n7302) );
  AND U7485 ( .A(a[8]), .B(b[13]), .Z(n7301) );
  XNOR U7486 ( .A(n7306), .B(n7179), .Z(n7181) );
  XOR U7487 ( .A(n7307), .B(n7308), .Z(n7179) );
  ANDN U7488 ( .B(n7309), .A(n7310), .Z(n7307) );
  AND U7489 ( .A(a[9]), .B(b[12]), .Z(n7306) );
  XNOR U7490 ( .A(n7311), .B(n7184), .Z(n7186) );
  XOR U7491 ( .A(n7312), .B(n7313), .Z(n7184) );
  ANDN U7492 ( .B(n7314), .A(n7315), .Z(n7312) );
  AND U7493 ( .A(a[10]), .B(b[11]), .Z(n7311) );
  XNOR U7494 ( .A(n7316), .B(n7189), .Z(n7191) );
  XOR U7495 ( .A(n7317), .B(n7318), .Z(n7189) );
  ANDN U7496 ( .B(n7319), .A(n7320), .Z(n7317) );
  AND U7497 ( .A(b[10]), .B(a[11]), .Z(n7316) );
  XNOR U7498 ( .A(n7321), .B(n7194), .Z(n7196) );
  XOR U7499 ( .A(n7322), .B(n7323), .Z(n7194) );
  ANDN U7500 ( .B(n7324), .A(n7325), .Z(n7322) );
  AND U7501 ( .A(a[12]), .B(b[9]), .Z(n7321) );
  XNOR U7502 ( .A(n7326), .B(n7199), .Z(n7201) );
  XOR U7503 ( .A(n7327), .B(n7328), .Z(n7199) );
  ANDN U7504 ( .B(n7329), .A(n7330), .Z(n7327) );
  AND U7505 ( .A(b[8]), .B(a[13]), .Z(n7326) );
  XNOR U7506 ( .A(n7331), .B(n7204), .Z(n7206) );
  XOR U7507 ( .A(n7332), .B(n7333), .Z(n7204) );
  ANDN U7508 ( .B(n7334), .A(n7335), .Z(n7332) );
  AND U7509 ( .A(a[14]), .B(b[7]), .Z(n7331) );
  XNOR U7510 ( .A(n7336), .B(n7209), .Z(n7211) );
  XOR U7511 ( .A(n7337), .B(n7338), .Z(n7209) );
  ANDN U7512 ( .B(n7339), .A(n7340), .Z(n7337) );
  AND U7513 ( .A(b[6]), .B(a[15]), .Z(n7336) );
  XNOR U7514 ( .A(n7341), .B(n7214), .Z(n7216) );
  XOR U7515 ( .A(n7342), .B(n7343), .Z(n7214) );
  ANDN U7516 ( .B(n7344), .A(n7345), .Z(n7342) );
  AND U7517 ( .A(b[5]), .B(a[16]), .Z(n7341) );
  XNOR U7518 ( .A(n7346), .B(n7219), .Z(n7221) );
  XOR U7519 ( .A(n7347), .B(n7348), .Z(n7219) );
  ANDN U7520 ( .B(n7349), .A(n7350), .Z(n7347) );
  AND U7521 ( .A(b[4]), .B(a[17]), .Z(n7346) );
  XNOR U7522 ( .A(n7351), .B(n7352), .Z(n7233) );
  NANDN U7523 ( .A(n7353), .B(n7354), .Z(n7352) );
  XNOR U7524 ( .A(n7355), .B(n7224), .Z(n7226) );
  XNOR U7525 ( .A(n7356), .B(n7357), .Z(n7224) );
  AND U7526 ( .A(n7358), .B(n7359), .Z(n7356) );
  AND U7527 ( .A(b[3]), .B(a[18]), .Z(n7355) );
  NAND U7528 ( .A(a[21]), .B(b[0]), .Z(n7115) );
  IV U7529 ( .A(n7237), .Z(n7240) );
  XOR U7530 ( .A(n7360), .B(n7361), .Z(n7237) );
  ANDN U7531 ( .B(n7362), .A(n7363), .Z(n7360) );
  XNOR U7532 ( .A(n7362), .B(n7363), .Z(c[52]) );
  XNOR U7533 ( .A(sreg[84]), .B(n7364), .Z(n7363) );
  XNOR U7534 ( .A(n7364), .B(n7365), .Z(n7362) );
  XOR U7535 ( .A(n7245), .B(n7246), .Z(n7365) );
  XNOR U7536 ( .A(n7353), .B(n7354), .Z(n7246) );
  XOR U7537 ( .A(n7351), .B(n7366), .Z(n7354) );
  NAND U7538 ( .A(b[1]), .B(a[19]), .Z(n7366) );
  XOR U7539 ( .A(n7359), .B(n7367), .Z(n7353) );
  XOR U7540 ( .A(n7351), .B(n7358), .Z(n7367) );
  XNOR U7541 ( .A(n7368), .B(n7357), .Z(n7358) );
  AND U7542 ( .A(b[2]), .B(a[18]), .Z(n7368) );
  NANDN U7543 ( .A(n7369), .B(n7370), .Z(n7351) );
  XOR U7544 ( .A(n7357), .B(n7349), .Z(n7371) );
  XNOR U7545 ( .A(n7348), .B(n7344), .Z(n7372) );
  XNOR U7546 ( .A(n7343), .B(n7339), .Z(n7373) );
  XNOR U7547 ( .A(n7338), .B(n7334), .Z(n7374) );
  XNOR U7548 ( .A(n7333), .B(n7329), .Z(n7375) );
  XNOR U7549 ( .A(n7328), .B(n7324), .Z(n7376) );
  XNOR U7550 ( .A(n7323), .B(n7319), .Z(n7377) );
  XNOR U7551 ( .A(n7318), .B(n7314), .Z(n7378) );
  XNOR U7552 ( .A(n7313), .B(n7309), .Z(n7379) );
  XNOR U7553 ( .A(n7308), .B(n7304), .Z(n7380) );
  XNOR U7554 ( .A(n7303), .B(n7299), .Z(n7381) );
  XNOR U7555 ( .A(n7298), .B(n7294), .Z(n7382) );
  XNOR U7556 ( .A(n7293), .B(n7289), .Z(n7383) );
  XNOR U7557 ( .A(n7288), .B(n7284), .Z(n7384) );
  XNOR U7558 ( .A(n7283), .B(n7279), .Z(n7385) );
  XNOR U7559 ( .A(n7278), .B(n7274), .Z(n7386) );
  XNOR U7560 ( .A(n7273), .B(n7269), .Z(n7387) );
  XNOR U7561 ( .A(n7388), .B(n7268), .Z(n7269) );
  AND U7562 ( .A(a[0]), .B(b[20]), .Z(n7388) );
  XOR U7563 ( .A(n7389), .B(n7268), .Z(n7270) );
  XNOR U7564 ( .A(n7390), .B(n7391), .Z(n7268) );
  ANDN U7565 ( .B(n7392), .A(n7393), .Z(n7390) );
  AND U7566 ( .A(a[1]), .B(b[19]), .Z(n7389) );
  XNOR U7567 ( .A(n7394), .B(n7273), .Z(n7275) );
  XOR U7568 ( .A(n7395), .B(n7396), .Z(n7273) );
  ANDN U7569 ( .B(n7397), .A(n7398), .Z(n7395) );
  AND U7570 ( .A(a[2]), .B(b[18]), .Z(n7394) );
  XNOR U7571 ( .A(n7399), .B(n7278), .Z(n7280) );
  XOR U7572 ( .A(n7400), .B(n7401), .Z(n7278) );
  ANDN U7573 ( .B(n7402), .A(n7403), .Z(n7400) );
  AND U7574 ( .A(a[3]), .B(b[17]), .Z(n7399) );
  XNOR U7575 ( .A(n7404), .B(n7283), .Z(n7285) );
  XOR U7576 ( .A(n7405), .B(n7406), .Z(n7283) );
  ANDN U7577 ( .B(n7407), .A(n7408), .Z(n7405) );
  AND U7578 ( .A(a[4]), .B(b[16]), .Z(n7404) );
  XNOR U7579 ( .A(n7409), .B(n7288), .Z(n7290) );
  XOR U7580 ( .A(n7410), .B(n7411), .Z(n7288) );
  ANDN U7581 ( .B(n7412), .A(n7413), .Z(n7410) );
  AND U7582 ( .A(a[5]), .B(b[15]), .Z(n7409) );
  XNOR U7583 ( .A(n7414), .B(n7293), .Z(n7295) );
  XOR U7584 ( .A(n7415), .B(n7416), .Z(n7293) );
  ANDN U7585 ( .B(n7417), .A(n7418), .Z(n7415) );
  AND U7586 ( .A(a[6]), .B(b[14]), .Z(n7414) );
  XNOR U7587 ( .A(n7419), .B(n7298), .Z(n7300) );
  XOR U7588 ( .A(n7420), .B(n7421), .Z(n7298) );
  ANDN U7589 ( .B(n7422), .A(n7423), .Z(n7420) );
  AND U7590 ( .A(a[7]), .B(b[13]), .Z(n7419) );
  XNOR U7591 ( .A(n7424), .B(n7303), .Z(n7305) );
  XOR U7592 ( .A(n7425), .B(n7426), .Z(n7303) );
  ANDN U7593 ( .B(n7427), .A(n7428), .Z(n7425) );
  AND U7594 ( .A(a[8]), .B(b[12]), .Z(n7424) );
  XNOR U7595 ( .A(n7429), .B(n7308), .Z(n7310) );
  XOR U7596 ( .A(n7430), .B(n7431), .Z(n7308) );
  ANDN U7597 ( .B(n7432), .A(n7433), .Z(n7430) );
  AND U7598 ( .A(a[9]), .B(b[11]), .Z(n7429) );
  XNOR U7599 ( .A(n7434), .B(n7313), .Z(n7315) );
  XOR U7600 ( .A(n7435), .B(n7436), .Z(n7313) );
  ANDN U7601 ( .B(n7437), .A(n7438), .Z(n7435) );
  AND U7602 ( .A(a[10]), .B(b[10]), .Z(n7434) );
  XNOR U7603 ( .A(n7439), .B(n7318), .Z(n7320) );
  XOR U7604 ( .A(n7440), .B(n7441), .Z(n7318) );
  ANDN U7605 ( .B(n7442), .A(n7443), .Z(n7440) );
  AND U7606 ( .A(b[9]), .B(a[11]), .Z(n7439) );
  XNOR U7607 ( .A(n7444), .B(n7323), .Z(n7325) );
  XOR U7608 ( .A(n7445), .B(n7446), .Z(n7323) );
  ANDN U7609 ( .B(n7447), .A(n7448), .Z(n7445) );
  AND U7610 ( .A(a[12]), .B(b[8]), .Z(n7444) );
  XNOR U7611 ( .A(n7449), .B(n7328), .Z(n7330) );
  XOR U7612 ( .A(n7450), .B(n7451), .Z(n7328) );
  ANDN U7613 ( .B(n7452), .A(n7453), .Z(n7450) );
  AND U7614 ( .A(b[7]), .B(a[13]), .Z(n7449) );
  XNOR U7615 ( .A(n7454), .B(n7333), .Z(n7335) );
  XOR U7616 ( .A(n7455), .B(n7456), .Z(n7333) );
  ANDN U7617 ( .B(n7457), .A(n7458), .Z(n7455) );
  AND U7618 ( .A(b[6]), .B(a[14]), .Z(n7454) );
  XNOR U7619 ( .A(n7459), .B(n7338), .Z(n7340) );
  XOR U7620 ( .A(n7460), .B(n7461), .Z(n7338) );
  ANDN U7621 ( .B(n7462), .A(n7463), .Z(n7460) );
  AND U7622 ( .A(b[5]), .B(a[15]), .Z(n7459) );
  XNOR U7623 ( .A(n7464), .B(n7343), .Z(n7345) );
  XOR U7624 ( .A(n7465), .B(n7466), .Z(n7343) );
  ANDN U7625 ( .B(n7467), .A(n7468), .Z(n7465) );
  AND U7626 ( .A(b[4]), .B(a[16]), .Z(n7464) );
  XNOR U7627 ( .A(n7469), .B(n7470), .Z(n7357) );
  NANDN U7628 ( .A(n7471), .B(n7472), .Z(n7470) );
  XNOR U7629 ( .A(n7473), .B(n7348), .Z(n7350) );
  XNOR U7630 ( .A(n7474), .B(n7475), .Z(n7348) );
  AND U7631 ( .A(n7476), .B(n7477), .Z(n7474) );
  AND U7632 ( .A(b[3]), .B(a[17]), .Z(n7473) );
  NAND U7633 ( .A(a[20]), .B(b[0]), .Z(n7245) );
  IV U7634 ( .A(n7361), .Z(n7364) );
  XOR U7635 ( .A(n7478), .B(n7479), .Z(n7361) );
  ANDN U7636 ( .B(n7480), .A(n7481), .Z(n7478) );
  XNOR U7637 ( .A(n7480), .B(n7481), .Z(c[51]) );
  XNOR U7638 ( .A(sreg[83]), .B(n7482), .Z(n7481) );
  XNOR U7639 ( .A(n7482), .B(n7483), .Z(n7480) );
  XOR U7640 ( .A(n7369), .B(n7370), .Z(n7483) );
  XNOR U7641 ( .A(n7471), .B(n7472), .Z(n7370) );
  XOR U7642 ( .A(n7469), .B(n7484), .Z(n7472) );
  NAND U7643 ( .A(a[18]), .B(b[1]), .Z(n7484) );
  XOR U7644 ( .A(n7477), .B(n7485), .Z(n7471) );
  XOR U7645 ( .A(n7469), .B(n7476), .Z(n7485) );
  XNOR U7646 ( .A(n7486), .B(n7475), .Z(n7476) );
  AND U7647 ( .A(b[2]), .B(a[17]), .Z(n7486) );
  NANDN U7648 ( .A(n7487), .B(n7488), .Z(n7469) );
  XOR U7649 ( .A(n7475), .B(n7467), .Z(n7489) );
  XNOR U7650 ( .A(n7466), .B(n7462), .Z(n7490) );
  XNOR U7651 ( .A(n7461), .B(n7457), .Z(n7491) );
  XNOR U7652 ( .A(n7456), .B(n7452), .Z(n7492) );
  XNOR U7653 ( .A(n7451), .B(n7447), .Z(n7493) );
  XNOR U7654 ( .A(n7446), .B(n7442), .Z(n7494) );
  XNOR U7655 ( .A(n7441), .B(n7437), .Z(n7495) );
  XNOR U7656 ( .A(n7436), .B(n7432), .Z(n7496) );
  XNOR U7657 ( .A(n7431), .B(n7427), .Z(n7497) );
  XNOR U7658 ( .A(n7426), .B(n7422), .Z(n7498) );
  XNOR U7659 ( .A(n7421), .B(n7417), .Z(n7499) );
  XNOR U7660 ( .A(n7416), .B(n7412), .Z(n7500) );
  XNOR U7661 ( .A(n7411), .B(n7407), .Z(n7501) );
  XNOR U7662 ( .A(n7406), .B(n7402), .Z(n7502) );
  XNOR U7663 ( .A(n7401), .B(n7397), .Z(n7503) );
  XNOR U7664 ( .A(n7396), .B(n7392), .Z(n7504) );
  XOR U7665 ( .A(n7505), .B(n7391), .Z(n7392) );
  AND U7666 ( .A(a[0]), .B(b[19]), .Z(n7505) );
  XNOR U7667 ( .A(n7506), .B(n7391), .Z(n7393) );
  XNOR U7668 ( .A(n7507), .B(n7508), .Z(n7391) );
  ANDN U7669 ( .B(n7509), .A(n7510), .Z(n7507) );
  AND U7670 ( .A(a[1]), .B(b[18]), .Z(n7506) );
  XNOR U7671 ( .A(n7511), .B(n7396), .Z(n7398) );
  XOR U7672 ( .A(n7512), .B(n7513), .Z(n7396) );
  ANDN U7673 ( .B(n7514), .A(n7515), .Z(n7512) );
  AND U7674 ( .A(a[2]), .B(b[17]), .Z(n7511) );
  XNOR U7675 ( .A(n7516), .B(n7401), .Z(n7403) );
  XOR U7676 ( .A(n7517), .B(n7518), .Z(n7401) );
  ANDN U7677 ( .B(n7519), .A(n7520), .Z(n7517) );
  AND U7678 ( .A(a[3]), .B(b[16]), .Z(n7516) );
  XNOR U7679 ( .A(n7521), .B(n7406), .Z(n7408) );
  XOR U7680 ( .A(n7522), .B(n7523), .Z(n7406) );
  ANDN U7681 ( .B(n7524), .A(n7525), .Z(n7522) );
  AND U7682 ( .A(a[4]), .B(b[15]), .Z(n7521) );
  XNOR U7683 ( .A(n7526), .B(n7411), .Z(n7413) );
  XOR U7684 ( .A(n7527), .B(n7528), .Z(n7411) );
  ANDN U7685 ( .B(n7529), .A(n7530), .Z(n7527) );
  AND U7686 ( .A(a[5]), .B(b[14]), .Z(n7526) );
  XNOR U7687 ( .A(n7531), .B(n7416), .Z(n7418) );
  XOR U7688 ( .A(n7532), .B(n7533), .Z(n7416) );
  ANDN U7689 ( .B(n7534), .A(n7535), .Z(n7532) );
  AND U7690 ( .A(a[6]), .B(b[13]), .Z(n7531) );
  XNOR U7691 ( .A(n7536), .B(n7421), .Z(n7423) );
  XOR U7692 ( .A(n7537), .B(n7538), .Z(n7421) );
  ANDN U7693 ( .B(n7539), .A(n7540), .Z(n7537) );
  AND U7694 ( .A(a[7]), .B(b[12]), .Z(n7536) );
  XNOR U7695 ( .A(n7541), .B(n7426), .Z(n7428) );
  XOR U7696 ( .A(n7542), .B(n7543), .Z(n7426) );
  ANDN U7697 ( .B(n7544), .A(n7545), .Z(n7542) );
  AND U7698 ( .A(a[8]), .B(b[11]), .Z(n7541) );
  XNOR U7699 ( .A(n7546), .B(n7431), .Z(n7433) );
  XOR U7700 ( .A(n7547), .B(n7548), .Z(n7431) );
  ANDN U7701 ( .B(n7549), .A(n7550), .Z(n7547) );
  AND U7702 ( .A(a[9]), .B(b[10]), .Z(n7546) );
  XNOR U7703 ( .A(n7551), .B(n7436), .Z(n7438) );
  XOR U7704 ( .A(n7552), .B(n7553), .Z(n7436) );
  ANDN U7705 ( .B(n7554), .A(n7555), .Z(n7552) );
  AND U7706 ( .A(a[10]), .B(b[9]), .Z(n7551) );
  XNOR U7707 ( .A(n7556), .B(n7441), .Z(n7443) );
  XOR U7708 ( .A(n7557), .B(n7558), .Z(n7441) );
  ANDN U7709 ( .B(n7559), .A(n7560), .Z(n7557) );
  AND U7710 ( .A(b[8]), .B(a[11]), .Z(n7556) );
  XNOR U7711 ( .A(n7561), .B(n7446), .Z(n7448) );
  XOR U7712 ( .A(n7562), .B(n7563), .Z(n7446) );
  ANDN U7713 ( .B(n7564), .A(n7565), .Z(n7562) );
  AND U7714 ( .A(a[12]), .B(b[7]), .Z(n7561) );
  XNOR U7715 ( .A(n7566), .B(n7451), .Z(n7453) );
  XOR U7716 ( .A(n7567), .B(n7568), .Z(n7451) );
  ANDN U7717 ( .B(n7569), .A(n7570), .Z(n7567) );
  AND U7718 ( .A(b[6]), .B(a[13]), .Z(n7566) );
  XNOR U7719 ( .A(n7571), .B(n7456), .Z(n7458) );
  XOR U7720 ( .A(n7572), .B(n7573), .Z(n7456) );
  ANDN U7721 ( .B(n7574), .A(n7575), .Z(n7572) );
  AND U7722 ( .A(b[5]), .B(a[14]), .Z(n7571) );
  XNOR U7723 ( .A(n7576), .B(n7461), .Z(n7463) );
  XOR U7724 ( .A(n7577), .B(n7578), .Z(n7461) );
  ANDN U7725 ( .B(n7579), .A(n7580), .Z(n7577) );
  AND U7726 ( .A(b[4]), .B(a[15]), .Z(n7576) );
  XNOR U7727 ( .A(n7581), .B(n7582), .Z(n7475) );
  NANDN U7728 ( .A(n7583), .B(n7584), .Z(n7582) );
  XNOR U7729 ( .A(n7585), .B(n7466), .Z(n7468) );
  XNOR U7730 ( .A(n7586), .B(n7587), .Z(n7466) );
  AND U7731 ( .A(n7588), .B(n7589), .Z(n7586) );
  AND U7732 ( .A(b[3]), .B(a[16]), .Z(n7585) );
  NAND U7733 ( .A(a[19]), .B(b[0]), .Z(n7369) );
  IV U7734 ( .A(n7479), .Z(n7482) );
  XOR U7735 ( .A(n7590), .B(n7591), .Z(n7479) );
  ANDN U7736 ( .B(n7592), .A(n7593), .Z(n7590) );
  XNOR U7737 ( .A(n7592), .B(n7593), .Z(c[50]) );
  XNOR U7738 ( .A(sreg[82]), .B(n7594), .Z(n7593) );
  XNOR U7739 ( .A(n7594), .B(n7595), .Z(n7592) );
  XOR U7740 ( .A(n7487), .B(n7488), .Z(n7595) );
  XNOR U7741 ( .A(n7583), .B(n7584), .Z(n7488) );
  XOR U7742 ( .A(n7581), .B(n7596), .Z(n7584) );
  NAND U7743 ( .A(b[1]), .B(a[17]), .Z(n7596) );
  XOR U7744 ( .A(n7589), .B(n7597), .Z(n7583) );
  XOR U7745 ( .A(n7581), .B(n7588), .Z(n7597) );
  XNOR U7746 ( .A(n7598), .B(n7587), .Z(n7588) );
  AND U7747 ( .A(b[2]), .B(a[16]), .Z(n7598) );
  NANDN U7748 ( .A(n7599), .B(n7600), .Z(n7581) );
  XOR U7749 ( .A(n7587), .B(n7579), .Z(n7601) );
  XNOR U7750 ( .A(n7578), .B(n7574), .Z(n7602) );
  XNOR U7751 ( .A(n7573), .B(n7569), .Z(n7603) );
  XNOR U7752 ( .A(n7568), .B(n7564), .Z(n7604) );
  XNOR U7753 ( .A(n7563), .B(n7559), .Z(n7605) );
  XNOR U7754 ( .A(n7558), .B(n7554), .Z(n7606) );
  XNOR U7755 ( .A(n7553), .B(n7549), .Z(n7607) );
  XNOR U7756 ( .A(n7548), .B(n7544), .Z(n7608) );
  XNOR U7757 ( .A(n7543), .B(n7539), .Z(n7609) );
  XNOR U7758 ( .A(n7538), .B(n7534), .Z(n7610) );
  XNOR U7759 ( .A(n7533), .B(n7529), .Z(n7611) );
  XNOR U7760 ( .A(n7528), .B(n7524), .Z(n7612) );
  XNOR U7761 ( .A(n7523), .B(n7519), .Z(n7613) );
  XNOR U7762 ( .A(n7518), .B(n7514), .Z(n7614) );
  XNOR U7763 ( .A(n7513), .B(n7509), .Z(n7615) );
  XNOR U7764 ( .A(n7616), .B(n7508), .Z(n7509) );
  AND U7765 ( .A(a[0]), .B(b[18]), .Z(n7616) );
  XOR U7766 ( .A(n7617), .B(n7508), .Z(n7510) );
  XNOR U7767 ( .A(n7618), .B(n7619), .Z(n7508) );
  ANDN U7768 ( .B(n7620), .A(n7621), .Z(n7618) );
  AND U7769 ( .A(a[1]), .B(b[17]), .Z(n7617) );
  XNOR U7770 ( .A(n7622), .B(n7513), .Z(n7515) );
  XOR U7771 ( .A(n7623), .B(n7624), .Z(n7513) );
  ANDN U7772 ( .B(n7625), .A(n7626), .Z(n7623) );
  AND U7773 ( .A(a[2]), .B(b[16]), .Z(n7622) );
  XNOR U7774 ( .A(n7627), .B(n7518), .Z(n7520) );
  XOR U7775 ( .A(n7628), .B(n7629), .Z(n7518) );
  ANDN U7776 ( .B(n7630), .A(n7631), .Z(n7628) );
  AND U7777 ( .A(a[3]), .B(b[15]), .Z(n7627) );
  XNOR U7778 ( .A(n7632), .B(n7523), .Z(n7525) );
  XOR U7779 ( .A(n7633), .B(n7634), .Z(n7523) );
  ANDN U7780 ( .B(n7635), .A(n7636), .Z(n7633) );
  AND U7781 ( .A(a[4]), .B(b[14]), .Z(n7632) );
  XNOR U7782 ( .A(n7637), .B(n7528), .Z(n7530) );
  XOR U7783 ( .A(n7638), .B(n7639), .Z(n7528) );
  ANDN U7784 ( .B(n7640), .A(n7641), .Z(n7638) );
  AND U7785 ( .A(a[5]), .B(b[13]), .Z(n7637) );
  XNOR U7786 ( .A(n7642), .B(n7533), .Z(n7535) );
  XOR U7787 ( .A(n7643), .B(n7644), .Z(n7533) );
  ANDN U7788 ( .B(n7645), .A(n7646), .Z(n7643) );
  AND U7789 ( .A(a[6]), .B(b[12]), .Z(n7642) );
  XNOR U7790 ( .A(n7647), .B(n7538), .Z(n7540) );
  XOR U7791 ( .A(n7648), .B(n7649), .Z(n7538) );
  ANDN U7792 ( .B(n7650), .A(n7651), .Z(n7648) );
  AND U7793 ( .A(a[7]), .B(b[11]), .Z(n7647) );
  XNOR U7794 ( .A(n7652), .B(n7543), .Z(n7545) );
  XOR U7795 ( .A(n7653), .B(n7654), .Z(n7543) );
  ANDN U7796 ( .B(n7655), .A(n7656), .Z(n7653) );
  AND U7797 ( .A(a[8]), .B(b[10]), .Z(n7652) );
  XNOR U7798 ( .A(n7657), .B(n7548), .Z(n7550) );
  XOR U7799 ( .A(n7658), .B(n7659), .Z(n7548) );
  ANDN U7800 ( .B(n7660), .A(n7661), .Z(n7658) );
  AND U7801 ( .A(b[9]), .B(a[9]), .Z(n7657) );
  XNOR U7802 ( .A(n7662), .B(n7553), .Z(n7555) );
  XOR U7803 ( .A(n7663), .B(n7664), .Z(n7553) );
  ANDN U7804 ( .B(n7665), .A(n7666), .Z(n7663) );
  AND U7805 ( .A(a[10]), .B(b[8]), .Z(n7662) );
  XNOR U7806 ( .A(n7667), .B(n7558), .Z(n7560) );
  XOR U7807 ( .A(n7668), .B(n7669), .Z(n7558) );
  ANDN U7808 ( .B(n7670), .A(n7671), .Z(n7668) );
  AND U7809 ( .A(b[7]), .B(a[11]), .Z(n7667) );
  XNOR U7810 ( .A(n7672), .B(n7563), .Z(n7565) );
  XOR U7811 ( .A(n7673), .B(n7674), .Z(n7563) );
  ANDN U7812 ( .B(n7675), .A(n7676), .Z(n7673) );
  AND U7813 ( .A(b[6]), .B(a[12]), .Z(n7672) );
  XNOR U7814 ( .A(n7677), .B(n7568), .Z(n7570) );
  XOR U7815 ( .A(n7678), .B(n7679), .Z(n7568) );
  ANDN U7816 ( .B(n7680), .A(n7681), .Z(n7678) );
  AND U7817 ( .A(b[5]), .B(a[13]), .Z(n7677) );
  XNOR U7818 ( .A(n7682), .B(n7573), .Z(n7575) );
  XOR U7819 ( .A(n7683), .B(n7684), .Z(n7573) );
  ANDN U7820 ( .B(n7685), .A(n7686), .Z(n7683) );
  AND U7821 ( .A(b[4]), .B(a[14]), .Z(n7682) );
  XNOR U7822 ( .A(n7687), .B(n7688), .Z(n7587) );
  NANDN U7823 ( .A(n7689), .B(n7690), .Z(n7688) );
  XNOR U7824 ( .A(n7691), .B(n7578), .Z(n7580) );
  XNOR U7825 ( .A(n7692), .B(n7693), .Z(n7578) );
  AND U7826 ( .A(n7694), .B(n7695), .Z(n7692) );
  AND U7827 ( .A(b[3]), .B(a[15]), .Z(n7691) );
  NAND U7828 ( .A(a[18]), .B(b[0]), .Z(n7487) );
  IV U7829 ( .A(n7591), .Z(n7594) );
  XOR U7830 ( .A(n7696), .B(n7697), .Z(n7591) );
  ANDN U7831 ( .B(n7698), .A(n7699), .Z(n7696) );
  XNOR U7832 ( .A(n7698), .B(n7699), .Z(c[49]) );
  XNOR U7833 ( .A(sreg[81]), .B(n7700), .Z(n7699) );
  XNOR U7834 ( .A(n7700), .B(n7701), .Z(n7698) );
  XOR U7835 ( .A(n7599), .B(n7600), .Z(n7701) );
  XNOR U7836 ( .A(n7689), .B(n7690), .Z(n7600) );
  XOR U7837 ( .A(n7687), .B(n7702), .Z(n7690) );
  NAND U7838 ( .A(a[16]), .B(b[1]), .Z(n7702) );
  XOR U7839 ( .A(n7695), .B(n7703), .Z(n7689) );
  XOR U7840 ( .A(n7687), .B(n7694), .Z(n7703) );
  XNOR U7841 ( .A(n7704), .B(n7693), .Z(n7694) );
  AND U7842 ( .A(b[2]), .B(a[15]), .Z(n7704) );
  NANDN U7843 ( .A(n7705), .B(n7706), .Z(n7687) );
  XOR U7844 ( .A(n7693), .B(n7685), .Z(n7707) );
  XNOR U7845 ( .A(n7684), .B(n7680), .Z(n7708) );
  XNOR U7846 ( .A(n7679), .B(n7675), .Z(n7709) );
  XNOR U7847 ( .A(n7674), .B(n7670), .Z(n7710) );
  XNOR U7848 ( .A(n7669), .B(n7665), .Z(n7711) );
  XNOR U7849 ( .A(n7664), .B(n7660), .Z(n7712) );
  XNOR U7850 ( .A(n7659), .B(n7655), .Z(n7713) );
  XNOR U7851 ( .A(n7654), .B(n7650), .Z(n7714) );
  XNOR U7852 ( .A(n7649), .B(n7645), .Z(n7715) );
  XNOR U7853 ( .A(n7644), .B(n7640), .Z(n7716) );
  XNOR U7854 ( .A(n7639), .B(n7635), .Z(n7717) );
  XNOR U7855 ( .A(n7634), .B(n7630), .Z(n7718) );
  XNOR U7856 ( .A(n7629), .B(n7625), .Z(n7719) );
  XNOR U7857 ( .A(n7624), .B(n7620), .Z(n7720) );
  XOR U7858 ( .A(n7721), .B(n7619), .Z(n7620) );
  AND U7859 ( .A(a[0]), .B(b[17]), .Z(n7721) );
  XNOR U7860 ( .A(n7722), .B(n7619), .Z(n7621) );
  XNOR U7861 ( .A(n7723), .B(n7724), .Z(n7619) );
  ANDN U7862 ( .B(n7725), .A(n7726), .Z(n7723) );
  AND U7863 ( .A(a[1]), .B(b[16]), .Z(n7722) );
  XNOR U7864 ( .A(n7727), .B(n7624), .Z(n7626) );
  XOR U7865 ( .A(n7728), .B(n7729), .Z(n7624) );
  ANDN U7866 ( .B(n7730), .A(n7731), .Z(n7728) );
  AND U7867 ( .A(a[2]), .B(b[15]), .Z(n7727) );
  XNOR U7868 ( .A(n7732), .B(n7629), .Z(n7631) );
  XOR U7869 ( .A(n7733), .B(n7734), .Z(n7629) );
  ANDN U7870 ( .B(n7735), .A(n7736), .Z(n7733) );
  AND U7871 ( .A(a[3]), .B(b[14]), .Z(n7732) );
  XNOR U7872 ( .A(n7737), .B(n7634), .Z(n7636) );
  XOR U7873 ( .A(n7738), .B(n7739), .Z(n7634) );
  ANDN U7874 ( .B(n7740), .A(n7741), .Z(n7738) );
  AND U7875 ( .A(a[4]), .B(b[13]), .Z(n7737) );
  XNOR U7876 ( .A(n7742), .B(n7639), .Z(n7641) );
  XOR U7877 ( .A(n7743), .B(n7744), .Z(n7639) );
  ANDN U7878 ( .B(n7745), .A(n7746), .Z(n7743) );
  AND U7879 ( .A(a[5]), .B(b[12]), .Z(n7742) );
  XNOR U7880 ( .A(n7747), .B(n7644), .Z(n7646) );
  XOR U7881 ( .A(n7748), .B(n7749), .Z(n7644) );
  ANDN U7882 ( .B(n7750), .A(n7751), .Z(n7748) );
  AND U7883 ( .A(a[6]), .B(b[11]), .Z(n7747) );
  XNOR U7884 ( .A(n7752), .B(n7649), .Z(n7651) );
  XOR U7885 ( .A(n7753), .B(n7754), .Z(n7649) );
  ANDN U7886 ( .B(n7755), .A(n7756), .Z(n7753) );
  AND U7887 ( .A(a[7]), .B(b[10]), .Z(n7752) );
  XNOR U7888 ( .A(n7757), .B(n7654), .Z(n7656) );
  XOR U7889 ( .A(n7758), .B(n7759), .Z(n7654) );
  ANDN U7890 ( .B(n7760), .A(n7761), .Z(n7758) );
  AND U7891 ( .A(a[8]), .B(b[9]), .Z(n7757) );
  XNOR U7892 ( .A(n7762), .B(n7659), .Z(n7661) );
  XOR U7893 ( .A(n7763), .B(n7764), .Z(n7659) );
  ANDN U7894 ( .B(n7765), .A(n7766), .Z(n7763) );
  AND U7895 ( .A(b[8]), .B(a[9]), .Z(n7762) );
  XNOR U7896 ( .A(n7767), .B(n7664), .Z(n7666) );
  XOR U7897 ( .A(n7768), .B(n7769), .Z(n7664) );
  ANDN U7898 ( .B(n7770), .A(n7771), .Z(n7768) );
  AND U7899 ( .A(a[10]), .B(b[7]), .Z(n7767) );
  XNOR U7900 ( .A(n7772), .B(n7669), .Z(n7671) );
  XOR U7901 ( .A(n7773), .B(n7774), .Z(n7669) );
  ANDN U7902 ( .B(n7775), .A(n7776), .Z(n7773) );
  AND U7903 ( .A(b[6]), .B(a[11]), .Z(n7772) );
  XNOR U7904 ( .A(n7777), .B(n7674), .Z(n7676) );
  XOR U7905 ( .A(n7778), .B(n7779), .Z(n7674) );
  ANDN U7906 ( .B(n7780), .A(n7781), .Z(n7778) );
  AND U7907 ( .A(b[5]), .B(a[12]), .Z(n7777) );
  XNOR U7908 ( .A(n7782), .B(n7679), .Z(n7681) );
  XOR U7909 ( .A(n7783), .B(n7784), .Z(n7679) );
  ANDN U7910 ( .B(n7785), .A(n7786), .Z(n7783) );
  AND U7911 ( .A(b[4]), .B(a[13]), .Z(n7782) );
  XNOR U7912 ( .A(n7787), .B(n7788), .Z(n7693) );
  NANDN U7913 ( .A(n7789), .B(n7790), .Z(n7788) );
  XNOR U7914 ( .A(n7791), .B(n7684), .Z(n7686) );
  XNOR U7915 ( .A(n7792), .B(n7793), .Z(n7684) );
  AND U7916 ( .A(n7794), .B(n7795), .Z(n7792) );
  AND U7917 ( .A(b[3]), .B(a[14]), .Z(n7791) );
  NAND U7918 ( .A(a[17]), .B(b[0]), .Z(n7599) );
  IV U7919 ( .A(n7697), .Z(n7700) );
  XOR U7920 ( .A(n7796), .B(n7797), .Z(n7697) );
  ANDN U7921 ( .B(n7798), .A(n7799), .Z(n7796) );
  XNOR U7922 ( .A(n7798), .B(n7799), .Z(c[48]) );
  XNOR U7923 ( .A(sreg[80]), .B(n7800), .Z(n7799) );
  XNOR U7924 ( .A(n7800), .B(n7801), .Z(n7798) );
  XOR U7925 ( .A(n7705), .B(n7706), .Z(n7801) );
  XNOR U7926 ( .A(n7789), .B(n7790), .Z(n7706) );
  XOR U7927 ( .A(n7787), .B(n7802), .Z(n7790) );
  NAND U7928 ( .A(b[1]), .B(a[15]), .Z(n7802) );
  XOR U7929 ( .A(n7795), .B(n7803), .Z(n7789) );
  XOR U7930 ( .A(n7787), .B(n7794), .Z(n7803) );
  XNOR U7931 ( .A(n7804), .B(n7793), .Z(n7794) );
  AND U7932 ( .A(b[2]), .B(a[14]), .Z(n7804) );
  NANDN U7933 ( .A(n7805), .B(n7806), .Z(n7787) );
  XOR U7934 ( .A(n7793), .B(n7785), .Z(n7807) );
  XNOR U7935 ( .A(n7784), .B(n7780), .Z(n7808) );
  XNOR U7936 ( .A(n7779), .B(n7775), .Z(n7809) );
  XNOR U7937 ( .A(n7774), .B(n7770), .Z(n7810) );
  XNOR U7938 ( .A(n7769), .B(n7765), .Z(n7811) );
  XNOR U7939 ( .A(n7764), .B(n7760), .Z(n7812) );
  XNOR U7940 ( .A(n7759), .B(n7755), .Z(n7813) );
  XNOR U7941 ( .A(n7754), .B(n7750), .Z(n7814) );
  XNOR U7942 ( .A(n7749), .B(n7745), .Z(n7815) );
  XNOR U7943 ( .A(n7744), .B(n7740), .Z(n7816) );
  XNOR U7944 ( .A(n7739), .B(n7735), .Z(n7817) );
  XNOR U7945 ( .A(n7734), .B(n7730), .Z(n7818) );
  XNOR U7946 ( .A(n7729), .B(n7725), .Z(n7819) );
  XNOR U7947 ( .A(n7820), .B(n7724), .Z(n7725) );
  AND U7948 ( .A(a[0]), .B(b[16]), .Z(n7820) );
  XOR U7949 ( .A(n7821), .B(n7724), .Z(n7726) );
  XNOR U7950 ( .A(n7822), .B(n7823), .Z(n7724) );
  ANDN U7951 ( .B(n7824), .A(n7825), .Z(n7822) );
  AND U7952 ( .A(a[1]), .B(b[15]), .Z(n7821) );
  XNOR U7953 ( .A(n7826), .B(n7729), .Z(n7731) );
  XOR U7954 ( .A(n7827), .B(n7828), .Z(n7729) );
  ANDN U7955 ( .B(n7829), .A(n7830), .Z(n7827) );
  AND U7956 ( .A(a[2]), .B(b[14]), .Z(n7826) );
  XNOR U7957 ( .A(n7831), .B(n7734), .Z(n7736) );
  XOR U7958 ( .A(n7832), .B(n7833), .Z(n7734) );
  ANDN U7959 ( .B(n7834), .A(n7835), .Z(n7832) );
  AND U7960 ( .A(a[3]), .B(b[13]), .Z(n7831) );
  XNOR U7961 ( .A(n7836), .B(n7739), .Z(n7741) );
  XOR U7962 ( .A(n7837), .B(n7838), .Z(n7739) );
  ANDN U7963 ( .B(n7839), .A(n7840), .Z(n7837) );
  AND U7964 ( .A(a[4]), .B(b[12]), .Z(n7836) );
  XNOR U7965 ( .A(n7841), .B(n7744), .Z(n7746) );
  XOR U7966 ( .A(n7842), .B(n7843), .Z(n7744) );
  ANDN U7967 ( .B(n7844), .A(n7845), .Z(n7842) );
  AND U7968 ( .A(a[5]), .B(b[11]), .Z(n7841) );
  XNOR U7969 ( .A(n7846), .B(n7749), .Z(n7751) );
  XOR U7970 ( .A(n7847), .B(n7848), .Z(n7749) );
  ANDN U7971 ( .B(n7849), .A(n7850), .Z(n7847) );
  AND U7972 ( .A(a[6]), .B(b[10]), .Z(n7846) );
  XNOR U7973 ( .A(n7851), .B(n7754), .Z(n7756) );
  XOR U7974 ( .A(n7852), .B(n7853), .Z(n7754) );
  ANDN U7975 ( .B(n7854), .A(n7855), .Z(n7852) );
  AND U7976 ( .A(a[7]), .B(b[9]), .Z(n7851) );
  XNOR U7977 ( .A(n7856), .B(n7759), .Z(n7761) );
  XOR U7978 ( .A(n7857), .B(n7858), .Z(n7759) );
  ANDN U7979 ( .B(n7859), .A(n7860), .Z(n7857) );
  AND U7980 ( .A(a[8]), .B(b[8]), .Z(n7856) );
  XNOR U7981 ( .A(n7861), .B(n7764), .Z(n7766) );
  XOR U7982 ( .A(n7862), .B(n7863), .Z(n7764) );
  ANDN U7983 ( .B(n7864), .A(n7865), .Z(n7862) );
  AND U7984 ( .A(b[7]), .B(a[9]), .Z(n7861) );
  XNOR U7985 ( .A(n7866), .B(n7769), .Z(n7771) );
  XOR U7986 ( .A(n7867), .B(n7868), .Z(n7769) );
  ANDN U7987 ( .B(n7869), .A(n7870), .Z(n7867) );
  AND U7988 ( .A(b[6]), .B(a[10]), .Z(n7866) );
  XNOR U7989 ( .A(n7871), .B(n7774), .Z(n7776) );
  XOR U7990 ( .A(n7872), .B(n7873), .Z(n7774) );
  ANDN U7991 ( .B(n7874), .A(n7875), .Z(n7872) );
  AND U7992 ( .A(b[5]), .B(a[11]), .Z(n7871) );
  XNOR U7993 ( .A(n7876), .B(n7779), .Z(n7781) );
  XOR U7994 ( .A(n7877), .B(n7878), .Z(n7779) );
  ANDN U7995 ( .B(n7879), .A(n7880), .Z(n7877) );
  AND U7996 ( .A(b[4]), .B(a[12]), .Z(n7876) );
  XNOR U7997 ( .A(n7881), .B(n7882), .Z(n7793) );
  NANDN U7998 ( .A(n7883), .B(n7884), .Z(n7882) );
  XNOR U7999 ( .A(n7885), .B(n7784), .Z(n7786) );
  XNOR U8000 ( .A(n7886), .B(n7887), .Z(n7784) );
  AND U8001 ( .A(n7888), .B(n7889), .Z(n7886) );
  AND U8002 ( .A(b[3]), .B(a[13]), .Z(n7885) );
  NAND U8003 ( .A(a[16]), .B(b[0]), .Z(n7705) );
  IV U8004 ( .A(n7797), .Z(n7800) );
  XOR U8005 ( .A(n7890), .B(n7891), .Z(n7797) );
  ANDN U8006 ( .B(n7892), .A(n7893), .Z(n7890) );
  XNOR U8007 ( .A(n7892), .B(n7893), .Z(c[47]) );
  XNOR U8008 ( .A(sreg[79]), .B(n7894), .Z(n7893) );
  XNOR U8009 ( .A(n7894), .B(n7895), .Z(n7892) );
  XOR U8010 ( .A(n7805), .B(n7806), .Z(n7895) );
  XNOR U8011 ( .A(n7883), .B(n7884), .Z(n7806) );
  XOR U8012 ( .A(n7881), .B(n7896), .Z(n7884) );
  NAND U8013 ( .A(a[14]), .B(b[1]), .Z(n7896) );
  XOR U8014 ( .A(n7889), .B(n7897), .Z(n7883) );
  XOR U8015 ( .A(n7881), .B(n7888), .Z(n7897) );
  XNOR U8016 ( .A(n7898), .B(n7887), .Z(n7888) );
  AND U8017 ( .A(b[2]), .B(a[13]), .Z(n7898) );
  NANDN U8018 ( .A(n7899), .B(n7900), .Z(n7881) );
  XOR U8019 ( .A(n7887), .B(n7879), .Z(n7901) );
  XNOR U8020 ( .A(n7878), .B(n7874), .Z(n7902) );
  XNOR U8021 ( .A(n7873), .B(n7869), .Z(n7903) );
  XNOR U8022 ( .A(n7868), .B(n7864), .Z(n7904) );
  XNOR U8023 ( .A(n7863), .B(n7859), .Z(n7905) );
  XNOR U8024 ( .A(n7858), .B(n7854), .Z(n7906) );
  XNOR U8025 ( .A(n7853), .B(n7849), .Z(n7907) );
  XNOR U8026 ( .A(n7848), .B(n7844), .Z(n7908) );
  XNOR U8027 ( .A(n7843), .B(n7839), .Z(n7909) );
  XNOR U8028 ( .A(n7838), .B(n7834), .Z(n7910) );
  XNOR U8029 ( .A(n7833), .B(n7829), .Z(n7911) );
  XNOR U8030 ( .A(n7828), .B(n7824), .Z(n7912) );
  XOR U8031 ( .A(n7913), .B(n7823), .Z(n7824) );
  AND U8032 ( .A(a[0]), .B(b[15]), .Z(n7913) );
  XNOR U8033 ( .A(n7914), .B(n7823), .Z(n7825) );
  XNOR U8034 ( .A(n7915), .B(n7916), .Z(n7823) );
  ANDN U8035 ( .B(n7917), .A(n7918), .Z(n7915) );
  AND U8036 ( .A(a[1]), .B(b[14]), .Z(n7914) );
  XNOR U8037 ( .A(n7919), .B(n7828), .Z(n7830) );
  XOR U8038 ( .A(n7920), .B(n7921), .Z(n7828) );
  ANDN U8039 ( .B(n7922), .A(n7923), .Z(n7920) );
  AND U8040 ( .A(a[2]), .B(b[13]), .Z(n7919) );
  XNOR U8041 ( .A(n7924), .B(n7833), .Z(n7835) );
  XOR U8042 ( .A(n7925), .B(n7926), .Z(n7833) );
  ANDN U8043 ( .B(n7927), .A(n7928), .Z(n7925) );
  AND U8044 ( .A(a[3]), .B(b[12]), .Z(n7924) );
  XNOR U8045 ( .A(n7929), .B(n7838), .Z(n7840) );
  XOR U8046 ( .A(n7930), .B(n7931), .Z(n7838) );
  ANDN U8047 ( .B(n7932), .A(n7933), .Z(n7930) );
  AND U8048 ( .A(a[4]), .B(b[11]), .Z(n7929) );
  XNOR U8049 ( .A(n7934), .B(n7843), .Z(n7845) );
  XOR U8050 ( .A(n7935), .B(n7936), .Z(n7843) );
  ANDN U8051 ( .B(n7937), .A(n7938), .Z(n7935) );
  AND U8052 ( .A(a[5]), .B(b[10]), .Z(n7934) );
  XNOR U8053 ( .A(n7939), .B(n7848), .Z(n7850) );
  XOR U8054 ( .A(n7940), .B(n7941), .Z(n7848) );
  ANDN U8055 ( .B(n7942), .A(n7943), .Z(n7940) );
  AND U8056 ( .A(a[6]), .B(b[9]), .Z(n7939) );
  XNOR U8057 ( .A(n7944), .B(n7853), .Z(n7855) );
  XOR U8058 ( .A(n7945), .B(n7946), .Z(n7853) );
  ANDN U8059 ( .B(n7947), .A(n7948), .Z(n7945) );
  AND U8060 ( .A(a[7]), .B(b[8]), .Z(n7944) );
  XNOR U8061 ( .A(n7949), .B(n7858), .Z(n7860) );
  XOR U8062 ( .A(n7950), .B(n7951), .Z(n7858) );
  ANDN U8063 ( .B(n7952), .A(n7953), .Z(n7950) );
  AND U8064 ( .A(a[8]), .B(b[7]), .Z(n7949) );
  XNOR U8065 ( .A(n7954), .B(n7863), .Z(n7865) );
  XOR U8066 ( .A(n7955), .B(n7956), .Z(n7863) );
  ANDN U8067 ( .B(n7957), .A(n7958), .Z(n7955) );
  AND U8068 ( .A(b[6]), .B(a[9]), .Z(n7954) );
  XNOR U8069 ( .A(n7959), .B(n7868), .Z(n7870) );
  XOR U8070 ( .A(n7960), .B(n7961), .Z(n7868) );
  ANDN U8071 ( .B(n7962), .A(n7963), .Z(n7960) );
  AND U8072 ( .A(b[5]), .B(a[10]), .Z(n7959) );
  XNOR U8073 ( .A(n7964), .B(n7873), .Z(n7875) );
  XOR U8074 ( .A(n7965), .B(n7966), .Z(n7873) );
  ANDN U8075 ( .B(n7967), .A(n7968), .Z(n7965) );
  AND U8076 ( .A(b[4]), .B(a[11]), .Z(n7964) );
  XNOR U8077 ( .A(n7969), .B(n7970), .Z(n7887) );
  NANDN U8078 ( .A(n7971), .B(n7972), .Z(n7970) );
  XNOR U8079 ( .A(n7973), .B(n7878), .Z(n7880) );
  XNOR U8080 ( .A(n7974), .B(n7975), .Z(n7878) );
  AND U8081 ( .A(n7976), .B(n7977), .Z(n7974) );
  AND U8082 ( .A(b[3]), .B(a[12]), .Z(n7973) );
  NAND U8083 ( .A(a[15]), .B(b[0]), .Z(n7805) );
  IV U8084 ( .A(n7891), .Z(n7894) );
  XOR U8085 ( .A(n7978), .B(n7979), .Z(n7891) );
  ANDN U8086 ( .B(n7980), .A(n7981), .Z(n7978) );
  XNOR U8087 ( .A(n7980), .B(n7981), .Z(c[46]) );
  XNOR U8088 ( .A(sreg[78]), .B(n7982), .Z(n7981) );
  XNOR U8089 ( .A(n7982), .B(n7983), .Z(n7980) );
  XOR U8090 ( .A(n7899), .B(n7900), .Z(n7983) );
  XNOR U8091 ( .A(n7971), .B(n7972), .Z(n7900) );
  XOR U8092 ( .A(n7969), .B(n7984), .Z(n7972) );
  NAND U8093 ( .A(b[1]), .B(a[13]), .Z(n7984) );
  XOR U8094 ( .A(n7977), .B(n7985), .Z(n7971) );
  XOR U8095 ( .A(n7969), .B(n7976), .Z(n7985) );
  XNOR U8096 ( .A(n7986), .B(n7975), .Z(n7976) );
  AND U8097 ( .A(b[2]), .B(a[12]), .Z(n7986) );
  NANDN U8098 ( .A(n7987), .B(n7988), .Z(n7969) );
  XOR U8099 ( .A(n7975), .B(n7967), .Z(n7989) );
  XNOR U8100 ( .A(n7966), .B(n7962), .Z(n7990) );
  XNOR U8101 ( .A(n7961), .B(n7957), .Z(n7991) );
  XNOR U8102 ( .A(n7956), .B(n7952), .Z(n7992) );
  XNOR U8103 ( .A(n7951), .B(n7947), .Z(n7993) );
  XNOR U8104 ( .A(n7946), .B(n7942), .Z(n7994) );
  XNOR U8105 ( .A(n7941), .B(n7937), .Z(n7995) );
  XNOR U8106 ( .A(n7936), .B(n7932), .Z(n7996) );
  XNOR U8107 ( .A(n7931), .B(n7927), .Z(n7997) );
  XNOR U8108 ( .A(n7926), .B(n7922), .Z(n7998) );
  XNOR U8109 ( .A(n7921), .B(n7917), .Z(n7999) );
  XNOR U8110 ( .A(n8000), .B(n7916), .Z(n7917) );
  AND U8111 ( .A(a[0]), .B(b[14]), .Z(n8000) );
  XOR U8112 ( .A(n8001), .B(n7916), .Z(n7918) );
  XNOR U8113 ( .A(n8002), .B(n8003), .Z(n7916) );
  ANDN U8114 ( .B(n8004), .A(n8005), .Z(n8002) );
  AND U8115 ( .A(a[1]), .B(b[13]), .Z(n8001) );
  XNOR U8116 ( .A(n8006), .B(n7921), .Z(n7923) );
  XOR U8117 ( .A(n8007), .B(n8008), .Z(n7921) );
  ANDN U8118 ( .B(n8009), .A(n8010), .Z(n8007) );
  AND U8119 ( .A(a[2]), .B(b[12]), .Z(n8006) );
  XNOR U8120 ( .A(n8011), .B(n7926), .Z(n7928) );
  XOR U8121 ( .A(n8012), .B(n8013), .Z(n7926) );
  ANDN U8122 ( .B(n8014), .A(n8015), .Z(n8012) );
  AND U8123 ( .A(a[3]), .B(b[11]), .Z(n8011) );
  XNOR U8124 ( .A(n8016), .B(n7931), .Z(n7933) );
  XOR U8125 ( .A(n8017), .B(n8018), .Z(n7931) );
  ANDN U8126 ( .B(n8019), .A(n8020), .Z(n8017) );
  AND U8127 ( .A(a[4]), .B(b[10]), .Z(n8016) );
  XNOR U8128 ( .A(n8021), .B(n7936), .Z(n7938) );
  XOR U8129 ( .A(n8022), .B(n8023), .Z(n7936) );
  ANDN U8130 ( .B(n8024), .A(n8025), .Z(n8022) );
  AND U8131 ( .A(a[5]), .B(b[9]), .Z(n8021) );
  XNOR U8132 ( .A(n8026), .B(n7941), .Z(n7943) );
  XOR U8133 ( .A(n8027), .B(n8028), .Z(n7941) );
  ANDN U8134 ( .B(n8029), .A(n8030), .Z(n8027) );
  AND U8135 ( .A(a[6]), .B(b[8]), .Z(n8026) );
  XNOR U8136 ( .A(n8031), .B(n7946), .Z(n7948) );
  XOR U8137 ( .A(n8032), .B(n8033), .Z(n7946) );
  ANDN U8138 ( .B(n8034), .A(n8035), .Z(n8032) );
  AND U8139 ( .A(b[7]), .B(a[7]), .Z(n8031) );
  XNOR U8140 ( .A(n8036), .B(n7951), .Z(n7953) );
  XOR U8141 ( .A(n8037), .B(n8038), .Z(n7951) );
  ANDN U8142 ( .B(n8039), .A(n8040), .Z(n8037) );
  AND U8143 ( .A(b[6]), .B(a[8]), .Z(n8036) );
  XNOR U8144 ( .A(n8041), .B(n7956), .Z(n7958) );
  XOR U8145 ( .A(n8042), .B(n8043), .Z(n7956) );
  ANDN U8146 ( .B(n8044), .A(n8045), .Z(n8042) );
  AND U8147 ( .A(b[5]), .B(a[9]), .Z(n8041) );
  XNOR U8148 ( .A(n8046), .B(n7961), .Z(n7963) );
  XOR U8149 ( .A(n8047), .B(n8048), .Z(n7961) );
  ANDN U8150 ( .B(n8049), .A(n8050), .Z(n8047) );
  AND U8151 ( .A(b[4]), .B(a[10]), .Z(n8046) );
  XNOR U8152 ( .A(n8051), .B(n8052), .Z(n7975) );
  NANDN U8153 ( .A(n8053), .B(n8054), .Z(n8052) );
  XNOR U8154 ( .A(n8055), .B(n7966), .Z(n7968) );
  XNOR U8155 ( .A(n8056), .B(n8057), .Z(n7966) );
  AND U8156 ( .A(n8058), .B(n8059), .Z(n8056) );
  AND U8157 ( .A(b[3]), .B(a[11]), .Z(n8055) );
  NAND U8158 ( .A(a[14]), .B(b[0]), .Z(n7899) );
  IV U8159 ( .A(n7979), .Z(n7982) );
  XOR U8160 ( .A(n8060), .B(n8061), .Z(n7979) );
  ANDN U8161 ( .B(n8062), .A(n8063), .Z(n8060) );
  XNOR U8162 ( .A(n8062), .B(n8063), .Z(c[45]) );
  XNOR U8163 ( .A(sreg[77]), .B(n8064), .Z(n8063) );
  XNOR U8164 ( .A(n8064), .B(n8065), .Z(n8062) );
  XOR U8165 ( .A(n7987), .B(n7988), .Z(n8065) );
  XNOR U8166 ( .A(n8053), .B(n8054), .Z(n7988) );
  XOR U8167 ( .A(n8051), .B(n8066), .Z(n8054) );
  NAND U8168 ( .A(a[12]), .B(b[1]), .Z(n8066) );
  XOR U8169 ( .A(n8059), .B(n8067), .Z(n8053) );
  XOR U8170 ( .A(n8051), .B(n8058), .Z(n8067) );
  XNOR U8171 ( .A(n8068), .B(n8057), .Z(n8058) );
  AND U8172 ( .A(b[2]), .B(a[11]), .Z(n8068) );
  NANDN U8173 ( .A(n8069), .B(n8070), .Z(n8051) );
  XOR U8174 ( .A(n8057), .B(n8049), .Z(n8071) );
  XNOR U8175 ( .A(n8048), .B(n8044), .Z(n8072) );
  XNOR U8176 ( .A(n8043), .B(n8039), .Z(n8073) );
  XNOR U8177 ( .A(n8038), .B(n8034), .Z(n8074) );
  XNOR U8178 ( .A(n8033), .B(n8029), .Z(n8075) );
  XNOR U8179 ( .A(n8028), .B(n8024), .Z(n8076) );
  XNOR U8180 ( .A(n8023), .B(n8019), .Z(n8077) );
  XNOR U8181 ( .A(n8018), .B(n8014), .Z(n8078) );
  XNOR U8182 ( .A(n8013), .B(n8009), .Z(n8079) );
  XNOR U8183 ( .A(n8008), .B(n8004), .Z(n8080) );
  XOR U8184 ( .A(n8081), .B(n8003), .Z(n8004) );
  AND U8185 ( .A(a[0]), .B(b[13]), .Z(n8081) );
  XNOR U8186 ( .A(n8082), .B(n8003), .Z(n8005) );
  XNOR U8187 ( .A(n8083), .B(n8084), .Z(n8003) );
  ANDN U8188 ( .B(n8085), .A(n8086), .Z(n8083) );
  AND U8189 ( .A(a[1]), .B(b[12]), .Z(n8082) );
  XNOR U8190 ( .A(n8087), .B(n8008), .Z(n8010) );
  XOR U8191 ( .A(n8088), .B(n8089), .Z(n8008) );
  ANDN U8192 ( .B(n8090), .A(n8091), .Z(n8088) );
  AND U8193 ( .A(a[2]), .B(b[11]), .Z(n8087) );
  XNOR U8194 ( .A(n8092), .B(n8013), .Z(n8015) );
  XOR U8195 ( .A(n8093), .B(n8094), .Z(n8013) );
  ANDN U8196 ( .B(n8095), .A(n8096), .Z(n8093) );
  AND U8197 ( .A(a[3]), .B(b[10]), .Z(n8092) );
  XNOR U8198 ( .A(n8097), .B(n8018), .Z(n8020) );
  XOR U8199 ( .A(n8098), .B(n8099), .Z(n8018) );
  ANDN U8200 ( .B(n8100), .A(n8101), .Z(n8098) );
  AND U8201 ( .A(a[4]), .B(b[9]), .Z(n8097) );
  XNOR U8202 ( .A(n8102), .B(n8023), .Z(n8025) );
  XOR U8203 ( .A(n8103), .B(n8104), .Z(n8023) );
  ANDN U8204 ( .B(n8105), .A(n8106), .Z(n8103) );
  AND U8205 ( .A(a[5]), .B(b[8]), .Z(n8102) );
  XNOR U8206 ( .A(n8107), .B(n8028), .Z(n8030) );
  XOR U8207 ( .A(n8108), .B(n8109), .Z(n8028) );
  ANDN U8208 ( .B(n8110), .A(n8111), .Z(n8108) );
  AND U8209 ( .A(a[6]), .B(b[7]), .Z(n8107) );
  XNOR U8210 ( .A(n8112), .B(n8033), .Z(n8035) );
  XOR U8211 ( .A(n8113), .B(n8114), .Z(n8033) );
  ANDN U8212 ( .B(n8115), .A(n8116), .Z(n8113) );
  AND U8213 ( .A(b[6]), .B(a[7]), .Z(n8112) );
  XNOR U8214 ( .A(n8117), .B(n8038), .Z(n8040) );
  XOR U8215 ( .A(n8118), .B(n8119), .Z(n8038) );
  ANDN U8216 ( .B(n8120), .A(n8121), .Z(n8118) );
  AND U8217 ( .A(b[5]), .B(a[8]), .Z(n8117) );
  XNOR U8218 ( .A(n8122), .B(n8043), .Z(n8045) );
  XOR U8219 ( .A(n8123), .B(n8124), .Z(n8043) );
  ANDN U8220 ( .B(n8125), .A(n8126), .Z(n8123) );
  AND U8221 ( .A(b[4]), .B(a[9]), .Z(n8122) );
  XNOR U8222 ( .A(n8127), .B(n8128), .Z(n8057) );
  NANDN U8223 ( .A(n8129), .B(n8130), .Z(n8128) );
  XNOR U8224 ( .A(n8131), .B(n8048), .Z(n8050) );
  XNOR U8225 ( .A(n8132), .B(n8133), .Z(n8048) );
  AND U8226 ( .A(n8134), .B(n8135), .Z(n8132) );
  AND U8227 ( .A(b[3]), .B(a[10]), .Z(n8131) );
  NAND U8228 ( .A(a[13]), .B(b[0]), .Z(n7987) );
  IV U8229 ( .A(n8061), .Z(n8064) );
  XOR U8230 ( .A(n8136), .B(n8137), .Z(n8061) );
  ANDN U8231 ( .B(n8138), .A(n8139), .Z(n8136) );
  XNOR U8232 ( .A(n8138), .B(n8139), .Z(c[44]) );
  XNOR U8233 ( .A(sreg[76]), .B(n8140), .Z(n8139) );
  XNOR U8234 ( .A(n8140), .B(n8141), .Z(n8138) );
  XOR U8235 ( .A(n8069), .B(n8070), .Z(n8141) );
  XNOR U8236 ( .A(n8129), .B(n8130), .Z(n8070) );
  XOR U8237 ( .A(n8127), .B(n8142), .Z(n8130) );
  NAND U8238 ( .A(b[1]), .B(a[11]), .Z(n8142) );
  XOR U8239 ( .A(n8135), .B(n8143), .Z(n8129) );
  XOR U8240 ( .A(n8127), .B(n8134), .Z(n8143) );
  XNOR U8241 ( .A(n8144), .B(n8133), .Z(n8134) );
  AND U8242 ( .A(b[2]), .B(a[10]), .Z(n8144) );
  NANDN U8243 ( .A(n8145), .B(n8146), .Z(n8127) );
  XOR U8244 ( .A(n8133), .B(n8125), .Z(n8147) );
  XNOR U8245 ( .A(n8124), .B(n8120), .Z(n8148) );
  XNOR U8246 ( .A(n8119), .B(n8115), .Z(n8149) );
  XNOR U8247 ( .A(n8114), .B(n8110), .Z(n8150) );
  XNOR U8248 ( .A(n8109), .B(n8105), .Z(n8151) );
  XNOR U8249 ( .A(n8104), .B(n8100), .Z(n8152) );
  XNOR U8250 ( .A(n8099), .B(n8095), .Z(n8153) );
  XNOR U8251 ( .A(n8094), .B(n8090), .Z(n8154) );
  XNOR U8252 ( .A(n8089), .B(n8085), .Z(n8155) );
  XNOR U8253 ( .A(n8156), .B(n8084), .Z(n8085) );
  AND U8254 ( .A(a[0]), .B(b[12]), .Z(n8156) );
  XOR U8255 ( .A(n8157), .B(n8084), .Z(n8086) );
  XNOR U8256 ( .A(n8158), .B(n8159), .Z(n8084) );
  ANDN U8257 ( .B(n8160), .A(n8161), .Z(n8158) );
  AND U8258 ( .A(a[1]), .B(b[11]), .Z(n8157) );
  XNOR U8259 ( .A(n8162), .B(n8089), .Z(n8091) );
  XOR U8260 ( .A(n8163), .B(n8164), .Z(n8089) );
  ANDN U8261 ( .B(n8165), .A(n8166), .Z(n8163) );
  AND U8262 ( .A(a[2]), .B(b[10]), .Z(n8162) );
  XNOR U8263 ( .A(n8167), .B(n8094), .Z(n8096) );
  XOR U8264 ( .A(n8168), .B(n8169), .Z(n8094) );
  ANDN U8265 ( .B(n8170), .A(n8171), .Z(n8168) );
  AND U8266 ( .A(a[3]), .B(b[9]), .Z(n8167) );
  XNOR U8267 ( .A(n8172), .B(n8099), .Z(n8101) );
  XOR U8268 ( .A(n8173), .B(n8174), .Z(n8099) );
  ANDN U8269 ( .B(n8175), .A(n8176), .Z(n8173) );
  AND U8270 ( .A(a[4]), .B(b[8]), .Z(n8172) );
  XNOR U8271 ( .A(n8177), .B(n8104), .Z(n8106) );
  XOR U8272 ( .A(n8178), .B(n8179), .Z(n8104) );
  ANDN U8273 ( .B(n8180), .A(n8181), .Z(n8178) );
  AND U8274 ( .A(a[5]), .B(b[7]), .Z(n8177) );
  XNOR U8275 ( .A(n8182), .B(n8109), .Z(n8111) );
  XOR U8276 ( .A(n8183), .B(n8184), .Z(n8109) );
  ANDN U8277 ( .B(n8185), .A(n8186), .Z(n8183) );
  AND U8278 ( .A(b[6]), .B(a[6]), .Z(n8182) );
  XNOR U8279 ( .A(n8187), .B(n8114), .Z(n8116) );
  XOR U8280 ( .A(n8188), .B(n8189), .Z(n8114) );
  ANDN U8281 ( .B(n8190), .A(n8191), .Z(n8188) );
  AND U8282 ( .A(b[5]), .B(a[7]), .Z(n8187) );
  XNOR U8283 ( .A(n8192), .B(n8119), .Z(n8121) );
  XOR U8284 ( .A(n8193), .B(n8194), .Z(n8119) );
  ANDN U8285 ( .B(n8195), .A(n8196), .Z(n8193) );
  AND U8286 ( .A(b[4]), .B(a[8]), .Z(n8192) );
  XNOR U8287 ( .A(n8197), .B(n8198), .Z(n8133) );
  NANDN U8288 ( .A(n8199), .B(n8200), .Z(n8198) );
  XNOR U8289 ( .A(n8201), .B(n8124), .Z(n8126) );
  XNOR U8290 ( .A(n8202), .B(n8203), .Z(n8124) );
  AND U8291 ( .A(n8204), .B(n8205), .Z(n8202) );
  AND U8292 ( .A(b[3]), .B(a[9]), .Z(n8201) );
  NAND U8293 ( .A(a[12]), .B(b[0]), .Z(n8069) );
  IV U8294 ( .A(n8137), .Z(n8140) );
  XOR U8295 ( .A(n8206), .B(n8207), .Z(n8137) );
  ANDN U8296 ( .B(n8208), .A(n8209), .Z(n8206) );
  XNOR U8297 ( .A(n8208), .B(n8209), .Z(c[43]) );
  XNOR U8298 ( .A(sreg[75]), .B(n8210), .Z(n8209) );
  XNOR U8299 ( .A(n8210), .B(n8211), .Z(n8208) );
  XOR U8300 ( .A(n8145), .B(n8146), .Z(n8211) );
  XNOR U8301 ( .A(n8199), .B(n8200), .Z(n8146) );
  XOR U8302 ( .A(n8197), .B(n8212), .Z(n8200) );
  NAND U8303 ( .A(a[10]), .B(b[1]), .Z(n8212) );
  XOR U8304 ( .A(n8205), .B(n8213), .Z(n8199) );
  XOR U8305 ( .A(n8197), .B(n8204), .Z(n8213) );
  XNOR U8306 ( .A(n8214), .B(n8203), .Z(n8204) );
  AND U8307 ( .A(b[2]), .B(a[9]), .Z(n8214) );
  NANDN U8308 ( .A(n8215), .B(n8216), .Z(n8197) );
  XOR U8309 ( .A(n8203), .B(n8195), .Z(n8217) );
  XNOR U8310 ( .A(n8194), .B(n8190), .Z(n8218) );
  XNOR U8311 ( .A(n8189), .B(n8185), .Z(n8219) );
  XNOR U8312 ( .A(n8184), .B(n8180), .Z(n8220) );
  XNOR U8313 ( .A(n8179), .B(n8175), .Z(n8221) );
  XNOR U8314 ( .A(n8174), .B(n8170), .Z(n8222) );
  XNOR U8315 ( .A(n8169), .B(n8165), .Z(n8223) );
  XNOR U8316 ( .A(n8164), .B(n8160), .Z(n8224) );
  XOR U8317 ( .A(n8225), .B(n8159), .Z(n8160) );
  AND U8318 ( .A(a[0]), .B(b[11]), .Z(n8225) );
  XNOR U8319 ( .A(n8226), .B(n8159), .Z(n8161) );
  XNOR U8320 ( .A(n8227), .B(n8228), .Z(n8159) );
  ANDN U8321 ( .B(n8229), .A(n8230), .Z(n8227) );
  AND U8322 ( .A(a[1]), .B(b[10]), .Z(n8226) );
  XNOR U8323 ( .A(n8231), .B(n8164), .Z(n8166) );
  XOR U8324 ( .A(n8232), .B(n8233), .Z(n8164) );
  ANDN U8325 ( .B(n8234), .A(n8235), .Z(n8232) );
  AND U8326 ( .A(a[2]), .B(b[9]), .Z(n8231) );
  XNOR U8327 ( .A(n8236), .B(n8169), .Z(n8171) );
  XOR U8328 ( .A(n8237), .B(n8238), .Z(n8169) );
  ANDN U8329 ( .B(n8239), .A(n8240), .Z(n8237) );
  AND U8330 ( .A(a[3]), .B(b[8]), .Z(n8236) );
  XNOR U8331 ( .A(n8241), .B(n8174), .Z(n8176) );
  XOR U8332 ( .A(n8242), .B(n8243), .Z(n8174) );
  ANDN U8333 ( .B(n8244), .A(n8245), .Z(n8242) );
  AND U8334 ( .A(a[4]), .B(b[7]), .Z(n8241) );
  XNOR U8335 ( .A(n8246), .B(n8179), .Z(n8181) );
  XOR U8336 ( .A(n8247), .B(n8248), .Z(n8179) );
  ANDN U8337 ( .B(n8249), .A(n8250), .Z(n8247) );
  AND U8338 ( .A(b[6]), .B(a[5]), .Z(n8246) );
  XNOR U8339 ( .A(n8251), .B(n8184), .Z(n8186) );
  XOR U8340 ( .A(n8252), .B(n8253), .Z(n8184) );
  ANDN U8341 ( .B(n8254), .A(n8255), .Z(n8252) );
  AND U8342 ( .A(b[5]), .B(a[6]), .Z(n8251) );
  XNOR U8343 ( .A(n8256), .B(n8189), .Z(n8191) );
  XOR U8344 ( .A(n8257), .B(n8258), .Z(n8189) );
  ANDN U8345 ( .B(n8259), .A(n8260), .Z(n8257) );
  AND U8346 ( .A(b[4]), .B(a[7]), .Z(n8256) );
  XNOR U8347 ( .A(n8261), .B(n8262), .Z(n8203) );
  NANDN U8348 ( .A(n8263), .B(n8264), .Z(n8262) );
  XNOR U8349 ( .A(n8265), .B(n8194), .Z(n8196) );
  XNOR U8350 ( .A(n8266), .B(n8267), .Z(n8194) );
  AND U8351 ( .A(n8268), .B(n8269), .Z(n8266) );
  AND U8352 ( .A(b[3]), .B(a[8]), .Z(n8265) );
  NAND U8353 ( .A(a[11]), .B(b[0]), .Z(n8145) );
  IV U8354 ( .A(n8207), .Z(n8210) );
  XOR U8355 ( .A(n8270), .B(n8271), .Z(n8207) );
  ANDN U8356 ( .B(n8272), .A(n8273), .Z(n8270) );
  XNOR U8357 ( .A(n8272), .B(n8273), .Z(c[42]) );
  XNOR U8358 ( .A(sreg[74]), .B(n8274), .Z(n8273) );
  XNOR U8359 ( .A(n8274), .B(n8275), .Z(n8272) );
  XOR U8360 ( .A(n8215), .B(n8216), .Z(n8275) );
  XNOR U8361 ( .A(n8263), .B(n8264), .Z(n8216) );
  XOR U8362 ( .A(n8261), .B(n8276), .Z(n8264) );
  NAND U8363 ( .A(b[1]), .B(a[9]), .Z(n8276) );
  XOR U8364 ( .A(n8269), .B(n8277), .Z(n8263) );
  XOR U8365 ( .A(n8261), .B(n8268), .Z(n8277) );
  XNOR U8366 ( .A(n8278), .B(n8267), .Z(n8268) );
  AND U8367 ( .A(b[2]), .B(a[8]), .Z(n8278) );
  NANDN U8368 ( .A(n8279), .B(n8280), .Z(n8261) );
  XOR U8369 ( .A(n8267), .B(n8259), .Z(n8281) );
  XNOR U8370 ( .A(n8258), .B(n8254), .Z(n8282) );
  XNOR U8371 ( .A(n8253), .B(n8249), .Z(n8283) );
  XNOR U8372 ( .A(n8248), .B(n8244), .Z(n8284) );
  XNOR U8373 ( .A(n8243), .B(n8239), .Z(n8285) );
  XNOR U8374 ( .A(n8238), .B(n8234), .Z(n8286) );
  XNOR U8375 ( .A(n8233), .B(n8229), .Z(n8287) );
  XNOR U8376 ( .A(n8288), .B(n8228), .Z(n8229) );
  AND U8377 ( .A(a[0]), .B(b[10]), .Z(n8288) );
  XOR U8378 ( .A(n8289), .B(n8228), .Z(n8230) );
  XNOR U8379 ( .A(n8290), .B(n8291), .Z(n8228) );
  ANDN U8380 ( .B(n8292), .A(n8293), .Z(n8290) );
  AND U8381 ( .A(a[1]), .B(b[9]), .Z(n8289) );
  XNOR U8382 ( .A(n8294), .B(n8233), .Z(n8235) );
  XOR U8383 ( .A(n8295), .B(n8296), .Z(n8233) );
  ANDN U8384 ( .B(n8297), .A(n8298), .Z(n8295) );
  AND U8385 ( .A(a[2]), .B(b[8]), .Z(n8294) );
  XNOR U8386 ( .A(n8299), .B(n8238), .Z(n8240) );
  XOR U8387 ( .A(n8300), .B(n8301), .Z(n8238) );
  ANDN U8388 ( .B(n8302), .A(n8303), .Z(n8300) );
  AND U8389 ( .A(a[3]), .B(b[7]), .Z(n8299) );
  XNOR U8390 ( .A(n8304), .B(n8243), .Z(n8245) );
  XOR U8391 ( .A(n8305), .B(n8306), .Z(n8243) );
  ANDN U8392 ( .B(n8307), .A(n8308), .Z(n8305) );
  AND U8393 ( .A(b[6]), .B(a[4]), .Z(n8304) );
  XNOR U8394 ( .A(n8309), .B(n8248), .Z(n8250) );
  XOR U8395 ( .A(n8310), .B(n8311), .Z(n8248) );
  ANDN U8396 ( .B(n8312), .A(n8313), .Z(n8310) );
  AND U8397 ( .A(b[5]), .B(a[5]), .Z(n8309) );
  XNOR U8398 ( .A(n8314), .B(n8253), .Z(n8255) );
  XOR U8399 ( .A(n8315), .B(n8316), .Z(n8253) );
  ANDN U8400 ( .B(n8317), .A(n8318), .Z(n8315) );
  AND U8401 ( .A(b[4]), .B(a[6]), .Z(n8314) );
  XNOR U8402 ( .A(n8319), .B(n8320), .Z(n8267) );
  NANDN U8403 ( .A(n8321), .B(n8322), .Z(n8320) );
  XNOR U8404 ( .A(n8323), .B(n8258), .Z(n8260) );
  XNOR U8405 ( .A(n8324), .B(n8325), .Z(n8258) );
  AND U8406 ( .A(n8326), .B(n8327), .Z(n8324) );
  AND U8407 ( .A(b[3]), .B(a[7]), .Z(n8323) );
  NAND U8408 ( .A(a[10]), .B(b[0]), .Z(n8215) );
  IV U8409 ( .A(n8271), .Z(n8274) );
  XOR U8410 ( .A(n8328), .B(n8329), .Z(n8271) );
  ANDN U8411 ( .B(n8330), .A(n8331), .Z(n8328) );
  XNOR U8412 ( .A(n8330), .B(n8331), .Z(c[41]) );
  XNOR U8413 ( .A(sreg[73]), .B(n8332), .Z(n8331) );
  XNOR U8414 ( .A(n8332), .B(n8333), .Z(n8330) );
  XOR U8415 ( .A(n8279), .B(n8280), .Z(n8333) );
  XNOR U8416 ( .A(n8321), .B(n8322), .Z(n8280) );
  XOR U8417 ( .A(n8319), .B(n8334), .Z(n8322) );
  NAND U8418 ( .A(a[8]), .B(b[1]), .Z(n8334) );
  XOR U8419 ( .A(n8327), .B(n8335), .Z(n8321) );
  XOR U8420 ( .A(n8319), .B(n8326), .Z(n8335) );
  XNOR U8421 ( .A(n8336), .B(n8325), .Z(n8326) );
  AND U8422 ( .A(b[2]), .B(a[7]), .Z(n8336) );
  NANDN U8423 ( .A(n8337), .B(n8338), .Z(n8319) );
  XOR U8424 ( .A(n8325), .B(n8317), .Z(n8339) );
  XNOR U8425 ( .A(n8316), .B(n8312), .Z(n8340) );
  XNOR U8426 ( .A(n8311), .B(n8307), .Z(n8341) );
  XNOR U8427 ( .A(n8306), .B(n8302), .Z(n8342) );
  XNOR U8428 ( .A(n8301), .B(n8297), .Z(n8343) );
  XNOR U8429 ( .A(n8296), .B(n8292), .Z(n8344) );
  XOR U8430 ( .A(n8345), .B(n8291), .Z(n8292) );
  AND U8431 ( .A(a[0]), .B(b[9]), .Z(n8345) );
  XNOR U8432 ( .A(n8346), .B(n8291), .Z(n8293) );
  XNOR U8433 ( .A(n8347), .B(n8348), .Z(n8291) );
  ANDN U8434 ( .B(n8349), .A(n8350), .Z(n8347) );
  AND U8435 ( .A(a[1]), .B(b[8]), .Z(n8346) );
  XNOR U8436 ( .A(n8351), .B(n8296), .Z(n8298) );
  XOR U8437 ( .A(n8352), .B(n8353), .Z(n8296) );
  ANDN U8438 ( .B(n8354), .A(n8355), .Z(n8352) );
  AND U8439 ( .A(a[2]), .B(b[7]), .Z(n8351) );
  XNOR U8440 ( .A(n8356), .B(n8301), .Z(n8303) );
  XOR U8441 ( .A(n8357), .B(n8358), .Z(n8301) );
  ANDN U8442 ( .B(n8359), .A(n8360), .Z(n8357) );
  AND U8443 ( .A(b[6]), .B(a[3]), .Z(n8356) );
  XNOR U8444 ( .A(n8361), .B(n8306), .Z(n8308) );
  XOR U8445 ( .A(n8362), .B(n8363), .Z(n8306) );
  ANDN U8446 ( .B(n8364), .A(n8365), .Z(n8362) );
  AND U8447 ( .A(b[5]), .B(a[4]), .Z(n8361) );
  XNOR U8448 ( .A(n8366), .B(n8311), .Z(n8313) );
  XOR U8449 ( .A(n8367), .B(n8368), .Z(n8311) );
  ANDN U8450 ( .B(n8369), .A(n8370), .Z(n8367) );
  AND U8451 ( .A(b[4]), .B(a[5]), .Z(n8366) );
  XNOR U8452 ( .A(n8371), .B(n8372), .Z(n8325) );
  NANDN U8453 ( .A(n8373), .B(n8374), .Z(n8372) );
  XNOR U8454 ( .A(n8375), .B(n8316), .Z(n8318) );
  XNOR U8455 ( .A(n8376), .B(n8377), .Z(n8316) );
  AND U8456 ( .A(n8378), .B(n8379), .Z(n8376) );
  AND U8457 ( .A(b[3]), .B(a[6]), .Z(n8375) );
  NAND U8458 ( .A(a[9]), .B(b[0]), .Z(n8279) );
  IV U8459 ( .A(n8329), .Z(n8332) );
  XOR U8460 ( .A(n8380), .B(n8381), .Z(n8329) );
  ANDN U8461 ( .B(n8382), .A(n8383), .Z(n8380) );
  XNOR U8462 ( .A(n8382), .B(n8383), .Z(c[40]) );
  XNOR U8463 ( .A(sreg[72]), .B(n8384), .Z(n8383) );
  XNOR U8464 ( .A(n8384), .B(n8385), .Z(n8382) );
  XOR U8465 ( .A(n8337), .B(n8338), .Z(n8385) );
  XNOR U8466 ( .A(n8373), .B(n8374), .Z(n8338) );
  XOR U8467 ( .A(n8371), .B(n8386), .Z(n8374) );
  NAND U8468 ( .A(b[1]), .B(a[7]), .Z(n8386) );
  XOR U8469 ( .A(n8379), .B(n8387), .Z(n8373) );
  XOR U8470 ( .A(n8371), .B(n8378), .Z(n8387) );
  XNOR U8471 ( .A(n8388), .B(n8377), .Z(n8378) );
  AND U8472 ( .A(b[2]), .B(a[6]), .Z(n8388) );
  NANDN U8473 ( .A(n8389), .B(n8390), .Z(n8371) );
  XOR U8474 ( .A(n8377), .B(n8369), .Z(n8391) );
  XNOR U8475 ( .A(n8368), .B(n8364), .Z(n8392) );
  XNOR U8476 ( .A(n8363), .B(n8359), .Z(n8393) );
  XNOR U8477 ( .A(n8358), .B(n8354), .Z(n8394) );
  XNOR U8478 ( .A(n8353), .B(n8349), .Z(n8395) );
  XNOR U8479 ( .A(n8396), .B(n8348), .Z(n8349) );
  AND U8480 ( .A(a[0]), .B(b[8]), .Z(n8396) );
  XOR U8481 ( .A(n8397), .B(n8348), .Z(n8350) );
  XNOR U8482 ( .A(n8398), .B(n8399), .Z(n8348) );
  ANDN U8483 ( .B(n8400), .A(n8401), .Z(n8398) );
  AND U8484 ( .A(a[1]), .B(b[7]), .Z(n8397) );
  XNOR U8485 ( .A(n8402), .B(n8353), .Z(n8355) );
  XOR U8486 ( .A(n8403), .B(n8404), .Z(n8353) );
  ANDN U8487 ( .B(n8405), .A(n8406), .Z(n8403) );
  AND U8488 ( .A(b[6]), .B(a[2]), .Z(n8402) );
  XNOR U8489 ( .A(n8407), .B(n8358), .Z(n8360) );
  XOR U8490 ( .A(n8408), .B(n8409), .Z(n8358) );
  ANDN U8491 ( .B(n8410), .A(n8411), .Z(n8408) );
  AND U8492 ( .A(b[5]), .B(a[3]), .Z(n8407) );
  XNOR U8493 ( .A(n8412), .B(n8363), .Z(n8365) );
  XOR U8494 ( .A(n8413), .B(n8414), .Z(n8363) );
  ANDN U8495 ( .B(n8415), .A(n8416), .Z(n8413) );
  AND U8496 ( .A(b[4]), .B(a[4]), .Z(n8412) );
  XNOR U8497 ( .A(n8417), .B(n8418), .Z(n8377) );
  NANDN U8498 ( .A(n8419), .B(n8420), .Z(n8418) );
  XNOR U8499 ( .A(n8421), .B(n8368), .Z(n8370) );
  XNOR U8500 ( .A(n8422), .B(n8423), .Z(n8368) );
  AND U8501 ( .A(n8424), .B(n8425), .Z(n8422) );
  AND U8502 ( .A(b[3]), .B(a[5]), .Z(n8421) );
  NAND U8503 ( .A(a[8]), .B(b[0]), .Z(n8337) );
  IV U8504 ( .A(n8381), .Z(n8384) );
  XOR U8505 ( .A(n8426), .B(n8427), .Z(n8381) );
  ANDN U8506 ( .B(n8428), .A(n8429), .Z(n8426) );
  XNOR U8507 ( .A(n8428), .B(n8429), .Z(c[39]) );
  XNOR U8508 ( .A(sreg[71]), .B(n8430), .Z(n8429) );
  XNOR U8509 ( .A(n8430), .B(n8431), .Z(n8428) );
  XOR U8510 ( .A(n8389), .B(n8390), .Z(n8431) );
  XNOR U8511 ( .A(n8419), .B(n8420), .Z(n8390) );
  XOR U8512 ( .A(n8417), .B(n8432), .Z(n8420) );
  NAND U8513 ( .A(a[6]), .B(b[1]), .Z(n8432) );
  XOR U8514 ( .A(n8425), .B(n8433), .Z(n8419) );
  XOR U8515 ( .A(n8417), .B(n8424), .Z(n8433) );
  XNOR U8516 ( .A(n8434), .B(n8423), .Z(n8424) );
  AND U8517 ( .A(b[2]), .B(a[5]), .Z(n8434) );
  NANDN U8518 ( .A(n8435), .B(n8436), .Z(n8417) );
  XOR U8519 ( .A(n8423), .B(n8415), .Z(n8437) );
  XNOR U8520 ( .A(n8414), .B(n8410), .Z(n8438) );
  XNOR U8521 ( .A(n8409), .B(n8405), .Z(n8439) );
  XNOR U8522 ( .A(n8404), .B(n8400), .Z(n8440) );
  XOR U8523 ( .A(n8441), .B(n8399), .Z(n8400) );
  AND U8524 ( .A(a[0]), .B(b[7]), .Z(n8441) );
  XNOR U8525 ( .A(n8442), .B(n8399), .Z(n8401) );
  XNOR U8526 ( .A(n8443), .B(n8444), .Z(n8399) );
  ANDN U8527 ( .B(n8445), .A(n8446), .Z(n8443) );
  AND U8528 ( .A(b[6]), .B(a[1]), .Z(n8442) );
  XNOR U8529 ( .A(n8447), .B(n8404), .Z(n8406) );
  XOR U8530 ( .A(n8448), .B(n8449), .Z(n8404) );
  ANDN U8531 ( .B(n8450), .A(n8451), .Z(n8448) );
  AND U8532 ( .A(b[5]), .B(a[2]), .Z(n8447) );
  XNOR U8533 ( .A(n8452), .B(n8409), .Z(n8411) );
  XOR U8534 ( .A(n8453), .B(n8454), .Z(n8409) );
  ANDN U8535 ( .B(n8455), .A(n8456), .Z(n8453) );
  AND U8536 ( .A(b[4]), .B(a[3]), .Z(n8452) );
  XNOR U8537 ( .A(n8457), .B(n8458), .Z(n8423) );
  NANDN U8538 ( .A(n8459), .B(n8460), .Z(n8458) );
  XNOR U8539 ( .A(n8461), .B(n8414), .Z(n8416) );
  XNOR U8540 ( .A(n8462), .B(n8463), .Z(n8414) );
  AND U8541 ( .A(n8464), .B(n8465), .Z(n8462) );
  AND U8542 ( .A(b[3]), .B(a[4]), .Z(n8461) );
  NAND U8543 ( .A(a[7]), .B(b[0]), .Z(n8389) );
  IV U8544 ( .A(n8427), .Z(n8430) );
  XOR U8545 ( .A(n8466), .B(n8467), .Z(n8427) );
  ANDN U8546 ( .B(n8468), .A(n8469), .Z(n8466) );
  XNOR U8547 ( .A(n8468), .B(n8469), .Z(c[38]) );
  XNOR U8548 ( .A(sreg[70]), .B(n8470), .Z(n8469) );
  XNOR U8549 ( .A(n8470), .B(n8471), .Z(n8468) );
  XOR U8550 ( .A(n8435), .B(n8436), .Z(n8471) );
  XNOR U8551 ( .A(n8459), .B(n8460), .Z(n8436) );
  XOR U8552 ( .A(n8457), .B(n8472), .Z(n8460) );
  NAND U8553 ( .A(b[1]), .B(a[5]), .Z(n8472) );
  XOR U8554 ( .A(n8465), .B(n8473), .Z(n8459) );
  XOR U8555 ( .A(n8457), .B(n8464), .Z(n8473) );
  XNOR U8556 ( .A(n8474), .B(n8463), .Z(n8464) );
  AND U8557 ( .A(b[2]), .B(a[4]), .Z(n8474) );
  NANDN U8558 ( .A(n8475), .B(n8476), .Z(n8457) );
  XOR U8559 ( .A(n8463), .B(n8455), .Z(n8477) );
  XNOR U8560 ( .A(n8454), .B(n8450), .Z(n8478) );
  XNOR U8561 ( .A(n8449), .B(n8445), .Z(n8479) );
  XNOR U8562 ( .A(n8480), .B(n8444), .Z(n8445) );
  AND U8563 ( .A(b[6]), .B(a[0]), .Z(n8480) );
  XOR U8564 ( .A(n8481), .B(n8444), .Z(n8446) );
  XNOR U8565 ( .A(n8482), .B(n8483), .Z(n8444) );
  ANDN U8566 ( .B(n8484), .A(n8485), .Z(n8482) );
  AND U8567 ( .A(b[5]), .B(a[1]), .Z(n8481) );
  XNOR U8568 ( .A(n8486), .B(n8449), .Z(n8451) );
  XOR U8569 ( .A(n8487), .B(n8488), .Z(n8449) );
  ANDN U8570 ( .B(n8489), .A(n8490), .Z(n8487) );
  AND U8571 ( .A(b[4]), .B(a[2]), .Z(n8486) );
  XNOR U8572 ( .A(n8491), .B(n8492), .Z(n8463) );
  NANDN U8573 ( .A(n8493), .B(n8494), .Z(n8492) );
  XNOR U8574 ( .A(n8495), .B(n8454), .Z(n8456) );
  XNOR U8575 ( .A(n8496), .B(n8497), .Z(n8454) );
  AND U8576 ( .A(n8498), .B(n8499), .Z(n8496) );
  AND U8577 ( .A(b[3]), .B(a[3]), .Z(n8495) );
  NAND U8578 ( .A(a[6]), .B(b[0]), .Z(n8435) );
  IV U8579 ( .A(n8467), .Z(n8470) );
  XOR U8580 ( .A(n8500), .B(n8501), .Z(n8467) );
  ANDN U8581 ( .B(n8502), .A(n8503), .Z(n8500) );
  XNOR U8582 ( .A(n8502), .B(n8503), .Z(c[37]) );
  XNOR U8583 ( .A(sreg[69]), .B(n8504), .Z(n8503) );
  XNOR U8584 ( .A(n8504), .B(n8505), .Z(n8502) );
  XOR U8585 ( .A(n8475), .B(n8476), .Z(n8505) );
  XNOR U8586 ( .A(n8493), .B(n8494), .Z(n8476) );
  XOR U8587 ( .A(n8491), .B(n8506), .Z(n8494) );
  NAND U8588 ( .A(a[4]), .B(b[1]), .Z(n8506) );
  XOR U8589 ( .A(n8499), .B(n8507), .Z(n8493) );
  XOR U8590 ( .A(n8491), .B(n8498), .Z(n8507) );
  XNOR U8591 ( .A(n8508), .B(n8497), .Z(n8498) );
  AND U8592 ( .A(b[2]), .B(a[3]), .Z(n8508) );
  NANDN U8593 ( .A(n8509), .B(n8510), .Z(n8491) );
  XOR U8594 ( .A(n8497), .B(n8489), .Z(n8511) );
  XNOR U8595 ( .A(n8488), .B(n8484), .Z(n8512) );
  XOR U8596 ( .A(n8513), .B(n8483), .Z(n8484) );
  AND U8597 ( .A(b[5]), .B(a[0]), .Z(n8513) );
  XNOR U8598 ( .A(n8514), .B(n8483), .Z(n8485) );
  XNOR U8599 ( .A(n8515), .B(n8516), .Z(n8483) );
  ANDN U8600 ( .B(n8517), .A(n8518), .Z(n8515) );
  AND U8601 ( .A(b[4]), .B(a[1]), .Z(n8514) );
  XNOR U8602 ( .A(n8519), .B(n8520), .Z(n8497) );
  NANDN U8603 ( .A(n8521), .B(n8522), .Z(n8520) );
  XNOR U8604 ( .A(n8523), .B(n8488), .Z(n8490) );
  XNOR U8605 ( .A(n8524), .B(n8525), .Z(n8488) );
  AND U8606 ( .A(n8526), .B(n8527), .Z(n8524) );
  AND U8607 ( .A(b[3]), .B(a[2]), .Z(n8523) );
  NAND U8608 ( .A(a[5]), .B(b[0]), .Z(n8475) );
  IV U8609 ( .A(n8501), .Z(n8504) );
  XOR U8610 ( .A(n8528), .B(n8529), .Z(n8501) );
  ANDN U8611 ( .B(n8530), .A(n8531), .Z(n8528) );
  XNOR U8612 ( .A(n8530), .B(n8531), .Z(c[36]) );
  XNOR U8613 ( .A(sreg[68]), .B(n8532), .Z(n8531) );
  XNOR U8614 ( .A(n8532), .B(n8533), .Z(n8530) );
  XOR U8615 ( .A(n8509), .B(n8510), .Z(n8533) );
  XNOR U8616 ( .A(n8521), .B(n8522), .Z(n8510) );
  XOR U8617 ( .A(n8519), .B(n8534), .Z(n8522) );
  NAND U8618 ( .A(b[1]), .B(a[3]), .Z(n8534) );
  XOR U8619 ( .A(n8527), .B(n8535), .Z(n8521) );
  XOR U8620 ( .A(n8519), .B(n8526), .Z(n8535) );
  XNOR U8621 ( .A(n8536), .B(n8525), .Z(n8526) );
  AND U8622 ( .A(b[2]), .B(a[2]), .Z(n8536) );
  NANDN U8623 ( .A(n8537), .B(n8538), .Z(n8519) );
  XOR U8624 ( .A(n8525), .B(n8517), .Z(n8539) );
  XNOR U8625 ( .A(n8540), .B(n8516), .Z(n8517) );
  AND U8626 ( .A(b[4]), .B(a[0]), .Z(n8540) );
  XNOR U8627 ( .A(n8541), .B(n8542), .Z(n8525) );
  NANDN U8628 ( .A(n8543), .B(n8544), .Z(n8542) );
  XOR U8629 ( .A(n8545), .B(n8516), .Z(n8518) );
  XOR U8630 ( .A(n8546), .B(n8547), .Z(n8516) );
  AND U8631 ( .A(n8548), .B(n8549), .Z(n8546) );
  AND U8632 ( .A(b[3]), .B(a[1]), .Z(n8545) );
  NAND U8633 ( .A(a[4]), .B(b[0]), .Z(n8509) );
  IV U8634 ( .A(n8529), .Z(n8532) );
  XOR U8635 ( .A(n8550), .B(n8551), .Z(n8529) );
  ANDN U8636 ( .B(n8552), .A(n8553), .Z(n8550) );
  XNOR U8637 ( .A(n8552), .B(n8553), .Z(c[35]) );
  XNOR U8638 ( .A(sreg[67]), .B(n8554), .Z(n8553) );
  XNOR U8639 ( .A(n8554), .B(n8555), .Z(n8552) );
  XOR U8640 ( .A(n8537), .B(n8538), .Z(n8555) );
  XNOR U8641 ( .A(n8543), .B(n8544), .Z(n8538) );
  XOR U8642 ( .A(n8541), .B(n8556), .Z(n8544) );
  NAND U8643 ( .A(a[2]), .B(b[1]), .Z(n8556) );
  XOR U8644 ( .A(n8549), .B(n8557), .Z(n8543) );
  XOR U8645 ( .A(n8541), .B(n8548), .Z(n8557) );
  XNOR U8646 ( .A(n8558), .B(n8547), .Z(n8548) );
  AND U8647 ( .A(b[2]), .B(a[1]), .Z(n8558) );
  NANDN U8648 ( .A(n8559), .B(n8560), .Z(n8541) );
  XNOR U8649 ( .A(n8561), .B(n8547), .Z(n8549) );
  XOR U8650 ( .A(n8562), .B(n8563), .Z(n8547) );
  NAND U8651 ( .A(n8564), .B(n8565), .Z(n8563) );
  AND U8652 ( .A(b[3]), .B(a[0]), .Z(n8561) );
  NAND U8653 ( .A(a[3]), .B(b[0]), .Z(n8537) );
  IV U8654 ( .A(n8551), .Z(n8554) );
  XOR U8655 ( .A(n8566), .B(n8567), .Z(n8551) );
  ANDN U8656 ( .B(n8568), .A(n8569), .Z(n8566) );
  XNOR U8657 ( .A(n8568), .B(n8569), .Z(c[34]) );
  XOR U8658 ( .A(sreg[66]), .B(n8567), .Z(n8569) );
  XOR U8659 ( .A(n8567), .B(n8570), .Z(n8568) );
  XOR U8660 ( .A(n8559), .B(n8560), .Z(n8570) );
  XOR U8661 ( .A(n8564), .B(n8565), .Z(n8560) );
  XNOR U8662 ( .A(n8562), .B(n8571), .Z(n8565) );
  NAND U8663 ( .A(b[1]), .B(a[1]), .Z(n8571) );
  XOR U8664 ( .A(n8572), .B(n8562), .Z(n8564) );
  NOR U8665 ( .A(n8573), .B(n8574), .Z(n8562) );
  AND U8666 ( .A(b[2]), .B(a[0]), .Z(n8572) );
  NAND U8667 ( .A(a[2]), .B(b[0]), .Z(n8559) );
  XOR U8668 ( .A(n8575), .B(n8576), .Z(n8567) );
  NAND U8669 ( .A(n8577), .B(n8578), .Z(n8576) );
  XOR U8670 ( .A(n8577), .B(n8578), .Z(c[33]) );
  XOR U8671 ( .A(sreg[65]), .B(n8575), .Z(n8578) );
  XNOR U8672 ( .A(n8575), .B(n8579), .Z(n8577) );
  XNOR U8673 ( .A(n8573), .B(n8574), .Z(n8579) );
  NAND U8674 ( .A(b[0]), .B(a[1]), .Z(n8574) );
  NAND U8675 ( .A(b[1]), .B(a[0]), .Z(n8573) );
  ANDN U8676 ( .B(sreg[64]), .A(n8580), .Z(n8575) );
  XNOR U8677 ( .A(sreg[64]), .B(n8580), .Z(c[32]) );
  NAND U8678 ( .A(a[0]), .B(b[0]), .Z(n8580) );
endmodule

